// Benchmark "amba10c5y_cert" written by ABC on Sat Jul 29 22:48:07 2017

module amba10c5y_cert ( 
    n87, reg_i_hbusreq2_out, reg_controllable_hgrant8_out,
    reg_i_hbusreq3_out, reg_controllable_hgrant9_out, reg_i_hbusreq4_out,
    reg_i_hbusreq5_out, reg_i_hbusreq6_out, reg_controllable_nstart_out,
    reg_i_hbusreq7_out, reg_i_hbusreq8_out, reg_i_hbusreq9_out,
    reg_stateG3_0_out, reg_stateG3_1_out, reg_stateG3_2_out,
    reg_i_hlock9_out, reg_stateA1_out, reg_controllable_hmastlock_out,
    reg_i_hlock8_out, fair_cnt<0>_out , fair_cnt<1>_out ,
    fair_cnt<2>_out , reg_i_hlock7_out, reg_controllable_hmaster0_out,
    reg_stateG10_1_out, reg_i_hlock6_out, next_env_fair_out,
    reg_stateG10_2_out, reg_stateG2_out, reg_i_hlock5_out,
    reg_controllable_hmaster1_out, reg_stateG10_3_out, reg_i_hlock4_out,
    reg_controllable_hmaster2_out, reg_controllable_ndecide_out,
    reg_stateG10_4_out, reg_i_hready_out, reg_i_hlock3_out,
    reg_controllable_hmaster3_out, reg_stateG10_5_out,
    reg_controllable_hgrant1_out, reg_i_hlock2_out,
    reg_controllable_busreq_out, reg_i_hlock1_out, reg_stateG10_6_out,
    reg_controllable_hgrant2_out, reg_i_hlock0_out,
    reg_controllable_nhgrant0_out, reg_stateG10_7_out,
    reg_controllable_hgrant3_out, env_safe_err_happened_out,
    reg_stateG10_8_out, reg_controllable_hgrant4_out, reg_stateG10_9_out,
    reg_controllable_hgrant5_out, reg_i_hbusreq0_out,
    reg_controllable_hgrant6_out, next_sys_fair<0>_out ,
    next_sys_fair<1>_out , next_sys_fair<2>_out , next_sys_fair<3>_out ,
    next_sys_fair<4>_out , reg_i_hbusreq1_out,
    reg_controllable_hgrant7_out, reg_controllable_locked_out, i_hlock0,
    i_hlock1, i_hlock2, i_hlock3, i_hlock4, i_hlock5, i_hlock6, i_hlock7,
    i_hlock8, i_hlock9, i_hready, i_hburst1, i_hburst0, i_hbusreq0,
    i_hbusreq1, i_hbusreq2, i_hbusreq3, i_hbusreq4, i_hbusreq5, i_hbusreq6,
    i_hbusreq7, i_hbusreq8, i_hbusreq9, controllable_nhgrant0,
    controllable_hgrant1, controllable_locked, controllable_nstart,
    controllable_hgrant2, controllable_hgrant3, controllable_hgrant4,
    controllable_hgrant5, controllable_hgrant6, controllable_hgrant7,
    controllable_hgrant8, controllable_hgrant9, controllable_busreq,
    controllable_ndecide, controllable_hmaster3, controllable_hmaster2,
    controllable_hmaster1, controllable_hmaster0, controllable_hmastlock,
    inductivity_check   );
  input  n87, reg_i_hbusreq2_out, reg_controllable_hgrant8_out,
    reg_i_hbusreq3_out, reg_controllable_hgrant9_out, reg_i_hbusreq4_out,
    reg_i_hbusreq5_out, reg_i_hbusreq6_out, reg_controllable_nstart_out,
    reg_i_hbusreq7_out, reg_i_hbusreq8_out, reg_i_hbusreq9_out,
    reg_stateG3_0_out, reg_stateG3_1_out, reg_stateG3_2_out,
    reg_i_hlock9_out, reg_stateA1_out, reg_controllable_hmastlock_out,
    reg_i_hlock8_out, fair_cnt<0>_out , fair_cnt<1>_out ,
    fair_cnt<2>_out , reg_i_hlock7_out, reg_controllable_hmaster0_out,
    reg_stateG10_1_out, reg_i_hlock6_out, next_env_fair_out,
    reg_stateG10_2_out, reg_stateG2_out, reg_i_hlock5_out,
    reg_controllable_hmaster1_out, reg_stateG10_3_out, reg_i_hlock4_out,
    reg_controllable_hmaster2_out, reg_controllable_ndecide_out,
    reg_stateG10_4_out, reg_i_hready_out, reg_i_hlock3_out,
    reg_controllable_hmaster3_out, reg_stateG10_5_out,
    reg_controllable_hgrant1_out, reg_i_hlock2_out,
    reg_controllable_busreq_out, reg_i_hlock1_out, reg_stateG10_6_out,
    reg_controllable_hgrant2_out, reg_i_hlock0_out,
    reg_controllable_nhgrant0_out, reg_stateG10_7_out,
    reg_controllable_hgrant3_out, env_safe_err_happened_out,
    reg_stateG10_8_out, reg_controllable_hgrant4_out, reg_stateG10_9_out,
    reg_controllable_hgrant5_out, reg_i_hbusreq0_out,
    reg_controllable_hgrant6_out, next_sys_fair<0>_out ,
    next_sys_fair<1>_out , next_sys_fair<2>_out , next_sys_fair<3>_out ,
    next_sys_fair<4>_out , reg_i_hbusreq1_out,
    reg_controllable_hgrant7_out, reg_controllable_locked_out, i_hlock0,
    i_hlock1, i_hlock2, i_hlock3, i_hlock4, i_hlock5, i_hlock6, i_hlock7,
    i_hlock8, i_hlock9, i_hready, i_hburst1, i_hburst0, i_hbusreq0,
    i_hbusreq1, i_hbusreq2, i_hbusreq3, i_hbusreq4, i_hbusreq5, i_hbusreq6,
    i_hbusreq7, i_hbusreq8, i_hbusreq9, controllable_nhgrant0,
    controllable_hgrant1, controllable_locked, controllable_nstart,
    controllable_hgrant2, controllable_hgrant3, controllable_hgrant4,
    controllable_hgrant5, controllable_hgrant6, controllable_hgrant7,
    controllable_hgrant8, controllable_hgrant9, controllable_busreq,
    controllable_ndecide, controllable_hmaster3, controllable_hmaster2,
    controllable_hmaster1, controllable_hmaster0, controllable_hmastlock;
  output inductivity_check ;
  wire n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
    n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
    n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
    n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
    n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
    n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
    n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
    n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
    n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
    n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
    n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
    n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
    n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
    n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
    n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
    n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
    n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
    n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
    n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
    n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
    n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
    n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
    n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
    n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
    n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
    n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
    n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
    n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
    n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
    n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
    n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
    n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
    n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
    n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
    n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
    n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
    n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
    n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
    n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
    n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
    n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
    n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
    n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
    n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
    n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
    n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
    n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
    n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
    n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
    n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
    n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
    n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
    n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
    n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
    n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
    n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
    n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
    n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
    n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
    n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
    n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
    n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
    n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
    n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
    n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
    n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
    n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
    n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
    n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
    n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
    n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
    n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
    n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
    n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
    n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
    n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
    n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
    n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
    n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
    n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
    n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
    n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
    n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
    n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
    n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
    n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
    n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
    n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
    n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
    n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
    n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
    n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
    n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
    n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
    n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
    n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
    n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
    n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
    n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
    n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
    n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
    n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
    n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
    n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
    n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
    n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
    n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
    n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
    n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
    n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
    n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
    n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
    n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
    n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
    n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
    n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
    n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
    n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
    n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
    n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
    n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
    n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
    n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
    n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
    n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
    n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
    n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
    n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
    n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
    n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
    n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
    n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
    n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
    n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
    n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
    n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
    n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
    n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
    n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
    n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
    n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
    n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
    n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
    n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
    n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
    n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
    n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
    n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
    n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
    n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
    n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
    n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
    n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
    n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
    n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
    n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
    n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
    n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
    n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
    n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
    n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
    n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
    n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
    n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
    n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
    n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
    n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
    n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
    n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
    n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
    n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
    n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
    n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
    n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
    n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
    n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
    n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
    n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
    n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
    n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
    n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
    n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
    n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
    n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
    n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
    n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
    n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
    n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
    n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
    n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
    n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
    n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
    n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
    n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
    n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
    n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
    n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
    n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
    n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
    n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
    n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
    n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
    n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
    n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
    n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
    n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
    n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
    n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
    n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
    n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
    n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
    n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
    n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
    n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
    n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
    n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
    n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
    n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
    n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
    n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
    n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
    n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
    n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
    n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
    n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
    n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
    n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
    n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
    n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
    n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
    n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
    n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
    n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
    n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
    n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
    n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
    n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
    n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
    n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
    n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
    n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
    n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
    n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
    n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
    n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
    n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
    n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
    n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
    n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
    n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
    n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
    n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
    n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
    n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
    n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
    n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
    n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
    n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
    n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
    n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
    n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
    n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
    n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
    n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
    n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
    n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
    n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
    n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
    n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
    n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
    n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
    n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
    n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
    n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
    n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
    n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
    n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
    n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
    n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
    n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
    n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
    n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
    n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
    n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
    n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
    n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
    n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
    n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
    n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
    n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
    n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
    n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
    n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
    n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
    n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
    n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
    n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
    n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
    n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
    n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
    n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
    n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
    n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
    n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
    n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
    n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
    n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
    n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
    n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
    n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
    n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
    n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
    n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
    n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
    n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
    n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
    n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
    n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
    n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
    n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
    n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
    n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
    n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
    n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
    n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
    n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
    n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
    n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
    n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
    n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
    n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
    n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
    n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
    n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
    n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
    n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
    n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
    n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
    n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
    n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
    n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
    n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
    n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
    n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
    n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
    n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
    n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
    n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
    n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
    n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
    n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
    n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
    n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
    n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
    n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
    n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
    n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
    n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
    n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
    n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
    n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
    n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
    n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
    n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
    n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
    n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
    n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
    n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
    n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
    n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
    n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
    n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
    n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
    n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
    n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
    n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
    n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
    n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
    n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
    n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
    n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
    n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
    n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085,
    n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
    n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
    n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
    n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
    n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
    n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
    n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
    n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
    n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
    n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
    n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195,
    n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205,
    n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215,
    n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225,
    n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235,
    n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245,
    n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255,
    n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265,
    n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275,
    n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
    n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
    n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
    n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
    n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
    n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
    n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
    n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
    n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
    n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
    n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
    n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
    n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
    n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
    n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
    n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
    n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
    n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
    n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
    n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
    n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
    n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
    n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
    n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
    n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
    n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
    n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
    n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
    n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
    n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
    n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
    n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
    n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
    n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
    n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
    n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
    n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
    n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
    n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
    n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
    n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
    n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
    n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
    n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
    n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
    n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
    n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
    n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
    n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
    n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
    n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
    n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
    n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
    n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
    n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
    n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
    n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
    n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
    n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
    n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
    n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
    n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
    n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
    n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
    n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
    n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
    n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
    n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
    n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
    n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
    n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
    n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
    n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
    n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
    n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
    n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
    n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
    n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
    n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
    n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
    n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
    n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
    n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
    n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
    n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
    n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
    n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
    n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
    n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
    n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
    n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
    n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
    n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
    n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
    n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
    n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
    n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
    n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
    n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
    n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
    n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
    n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
    n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
    n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
    n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
    n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
    n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
    n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
    n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
    n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
    n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
    n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
    n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
    n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,
    n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
    n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,
    n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
    n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,
    n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
    n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
    n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485,
    n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495,
    n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505,
    n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515,
    n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525,
    n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,
    n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,
    n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555,
    n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565,
    n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575,
    n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
    n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595,
    n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
    n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
    n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
    n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,
    n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645,
    n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655,
    n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665,
    n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675,
    n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685,
    n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695,
    n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705,
    n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715,
    n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725,
    n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735,
    n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745,
    n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755,
    n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765,
    n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775,
    n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785,
    n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795,
    n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805,
    n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815,
    n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825,
    n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835,
    n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845,
    n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855,
    n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865,
    n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875,
    n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885,
    n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895,
    n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905,
    n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915,
    n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,
    n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,
    n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945,
    n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955,
    n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
    n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975,
    n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985,
    n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995,
    n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005,
    n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015,
    n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025,
    n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035,
    n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045,
    n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,
    n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
    n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
    n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085,
    n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095,
    n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105,
    n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115,
    n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125,
    n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135,
    n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145,
    n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155,
    n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165,
    n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175,
    n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185,
    n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195,
    n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205,
    n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215,
    n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225,
    n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235,
    n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245,
    n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255,
    n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265,
    n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275,
    n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285,
    n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295,
    n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305,
    n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315,
    n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325,
    n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335,
    n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345,
    n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355,
    n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365,
    n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375,
    n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385,
    n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395,
    n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405,
    n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415,
    n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425,
    n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435,
    n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445,
    n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455,
    n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465,
    n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475,
    n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485,
    n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495,
    n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505,
    n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515,
    n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
    n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535,
    n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545,
    n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
    n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
    n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
    n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
    n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
    n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
    n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
    n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
    n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
    n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
    n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
    n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
    n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
    n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
    n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
    n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
    n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
    n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
    n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
    n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
    n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
    n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
    n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
    n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
    n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
    n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
    n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
    n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
    n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
    n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
    n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
    n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
    n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
    n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
    n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
    n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
    n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
    n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
    n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
    n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
    n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
    n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
    n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
    n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
    n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
    n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
    n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
    n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
    n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
    n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
    n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
    n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
    n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
    n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
    n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
    n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
    n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
    n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
    n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
    n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
    n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
    n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
    n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
    n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
    n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
    n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
    n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
    n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
    n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
    n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
    n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
    n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
    n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
    n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
    n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
    n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
    n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
    n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
    n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
    n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
    n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
    n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
    n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
    n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
    n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
    n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
    n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
    n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
    n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
    n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
    n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
    n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
    n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
    n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
    n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
    n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
    n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
    n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
    n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
    n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
    n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
    n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
    n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
    n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
    n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
    n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
    n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
    n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
    n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
    n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
    n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
    n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
    n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
    n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
    n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
    n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705,
    n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715,
    n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
    n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735,
    n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745,
    n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755,
    n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
    n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
    n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
    n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
    n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
    n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
    n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
    n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
    n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
    n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
    n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
    n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
    n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
    n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
    n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
    n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
    n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
    n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
    n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
    n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
    n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
    n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
    n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
    n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
    n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
    n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
    n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
    n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
    n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
    n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
    n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
    n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
    n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
    n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
    n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
    n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
    n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
    n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
    n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
    n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
    n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
    n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
    n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
    n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
    n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
    n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
    n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
    n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
    n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
    n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
    n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
    n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
    n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
    n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
    n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
    n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315,
    n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325,
    n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335,
    n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345,
    n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355,
    n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365,
    n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375,
    n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385,
    n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395,
    n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
    n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415,
    n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
    n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
    n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
    n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
    n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
    n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
    n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
    n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
    n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
    n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515,
    n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
    n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
    n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545,
    n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
    n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
    n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
    n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
    n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595,
    n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605,
    n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615,
    n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
    n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635,
    n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645,
    n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655,
    n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665,
    n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675,
    n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685,
    n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695,
    n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705,
    n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715,
    n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725,
    n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735,
    n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745,
    n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755,
    n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765,
    n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775,
    n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
    n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795,
    n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805,
    n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815,
    n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
    n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
    n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
    n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
    n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
    n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
    n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
    n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
    n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
    n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
    n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
    n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
    n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
    n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
    n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
    n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
    n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
    n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
    n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
    n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
    n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
    n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035,
    n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
    n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055,
    n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
    n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
    n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
    n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
    n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
    n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
    n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
    n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
    n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
    n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
    n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
    n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
    n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
    n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
    n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
    n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
    n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
    n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
    n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
    n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
    n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
    n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
    n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
    n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
    n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
    n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
    n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
    n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
    n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
    n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355,
    n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
    n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
    n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
    n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
    n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
    n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
    n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
    n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
    n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
    n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
    n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
    n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
    n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
    n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
    n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
    n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
    n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
    n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
    n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545,
    n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555,
    n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565,
    n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575,
    n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585,
    n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595,
    n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605,
    n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615,
    n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625,
    n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635,
    n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645,
    n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655,
    n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665,
    n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675,
    n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685,
    n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
    n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705,
    n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715,
    n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
    n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
    n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
    n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
    n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
    n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
    n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
    n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
    n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
    n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
    n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
    n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
    n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
    n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
    n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
    n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
    n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
    n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
    n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
    n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
    n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
    n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
    n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
    n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
    n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
    n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
    n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
    n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
    n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
    n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
    n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022,
    n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
    n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
    n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
    n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
    n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
    n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076,
    n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
    n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094,
    n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
    n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
    n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
    n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
    n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
    n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148,
    n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157,
    n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166,
    n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
    n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
    n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
    n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
    n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
    n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220,
    n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229,
    n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238,
    n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
    n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
    n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
    n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
    n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283,
    n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292,
    n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301,
    n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310,
    n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
    n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
    n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
    n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
    n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355,
    n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364,
    n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373,
    n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382,
    n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
    n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
    n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
    n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
    n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427,
    n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436,
    n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445,
    n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454,
    n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
    n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
    n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
    n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
    n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499,
    n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508,
    n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517,
    n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526,
    n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
    n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
    n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
    n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562,
    n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571,
    n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580,
    n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589,
    n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598,
    n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
    n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
    n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
    n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634,
    n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643,
    n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652,
    n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661,
    n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670,
    n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
    n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
    n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
    n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706,
    n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715,
    n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724,
    n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733,
    n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742,
    n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
    n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
    n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
    n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778,
    n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787,
    n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796,
    n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805,
    n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814,
    n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
    n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
    n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
    n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850,
    n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859,
    n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868,
    n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877,
    n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886,
    n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
    n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
    n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
    n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922,
    n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931,
    n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940,
    n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949,
    n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958,
    n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
    n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
    n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
    n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994,
    n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003,
    n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012,
    n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021,
    n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030,
    n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
    n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
    n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
    n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066,
    n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075,
    n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084,
    n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093,
    n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102,
    n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
    n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
    n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
    n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138,
    n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147,
    n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156,
    n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165,
    n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174,
    n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
    n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
    n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
    n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210,
    n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219,
    n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228,
    n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237,
    n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246,
    n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
    n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
    n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
    n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282,
    n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291,
    n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300,
    n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309,
    n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318,
    n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
    n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
    n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
    n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354,
    n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363,
    n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372,
    n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381,
    n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390,
    n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
    n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
    n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
    n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426,
    n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435,
    n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444,
    n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453,
    n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462,
    n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
    n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
    n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
    n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498,
    n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507,
    n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516,
    n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525,
    n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534,
    n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
    n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
    n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
    n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570,
    n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579,
    n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588,
    n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597,
    n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606,
    n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
    n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
    n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
    n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642,
    n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651,
    n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660,
    n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669,
    n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678,
    n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
    n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
    n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
    n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714,
    n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723,
    n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732,
    n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741,
    n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750,
    n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
    n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
    n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
    n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786,
    n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795,
    n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804,
    n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813,
    n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822,
    n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
    n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
    n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
    n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858,
    n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867,
    n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876,
    n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885,
    n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894,
    n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
    n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
    n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
    n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930,
    n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939,
    n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948,
    n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957,
    n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966,
    n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
    n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
    n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
    n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002,
    n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011,
    n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020,
    n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029,
    n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038,
    n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
    n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
    n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
    n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074,
    n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083,
    n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092,
    n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101,
    n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110,
    n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
    n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
    n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
    n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146,
    n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155,
    n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164,
    n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173,
    n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182,
    n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
    n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
    n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
    n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218,
    n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227,
    n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236,
    n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245,
    n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254,
    n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
    n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
    n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
    n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
    n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299,
    n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308,
    n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317,
    n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326,
    n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
    n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
    n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
    n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362,
    n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371,
    n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380,
    n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389,
    n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398,
    n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
    n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
    n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
    n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434,
    n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443,
    n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452,
    n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461,
    n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470,
    n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
    n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
    n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
    n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506,
    n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515,
    n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524,
    n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533,
    n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542,
    n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
    n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
    n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
    n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578,
    n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587,
    n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596,
    n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605,
    n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614,
    n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
    n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
    n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
    n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650,
    n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659,
    n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668,
    n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677,
    n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686,
    n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
    n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
    n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
    n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722,
    n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731,
    n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740,
    n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749,
    n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758,
    n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
    n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
    n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
    n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794,
    n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803,
    n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812,
    n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821,
    n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830,
    n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
    n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
    n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
    n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866,
    n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875,
    n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884,
    n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893,
    n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902,
    n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
    n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
    n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
    n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938,
    n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947,
    n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956,
    n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965,
    n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974,
    n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
    n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
    n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
    n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010,
    n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019,
    n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028,
    n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037,
    n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046,
    n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055,
    n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
    n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
    n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082,
    n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091,
    n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100,
    n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109,
    n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118,
    n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127,
    n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
    n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
    n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154,
    n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163,
    n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172,
    n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181,
    n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190,
    n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199,
    n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
    n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
    n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226,
    n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235,
    n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244,
    n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253,
    n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262,
    n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271,
    n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
    n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
    n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298,
    n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307,
    n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316,
    n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325,
    n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334,
    n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343,
    n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
    n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
    n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370,
    n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379,
    n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388,
    n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397,
    n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406,
    n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415,
    n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
    n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
    n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
    n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451,
    n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460,
    n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469,
    n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478,
    n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487,
    n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
    n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
    n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
    n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523,
    n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532,
    n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541,
    n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550,
    n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559,
    n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
    n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
    n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
    n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595,
    n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604,
    n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613,
    n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622,
    n13623, n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631,
    n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
    n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
    n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
    n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667,
    n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676,
    n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685,
    n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694,
    n13695, n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703,
    n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
    n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
    n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730,
    n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739,
    n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748,
    n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757,
    n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766,
    n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775,
    n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
    n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
    n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802,
    n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811,
    n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820,
    n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829,
    n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837, n13838,
    n13839, n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847,
    n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
    n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
    n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
    n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883,
    n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892,
    n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901,
    n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909, n13910,
    n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919,
    n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
    n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
    n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
    n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955,
    n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964,
    n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973,
    n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982,
    n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991,
    n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
    n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
    n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
    n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027,
    n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036,
    n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045,
    n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053, n14054,
    n14055, n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063,
    n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
    n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
    n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,
    n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099,
    n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108,
    n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117,
    n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125, n14126,
    n14127, n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135,
    n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
    n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
    n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162,
    n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171,
    n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180,
    n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189,
    n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198,
    n14199, n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207,
    n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
    n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
    n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234,
    n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243,
    n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252,
    n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261,
    n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270,
    n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279,
    n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
    n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
    n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306,
    n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315,
    n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324,
    n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333,
    n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342,
    n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351,
    n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
    n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
    n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378,
    n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387,
    n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396,
    n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405,
    n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414,
    n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423,
    n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
    n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
    n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450,
    n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459,
    n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468,
    n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477,
    n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486,
    n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495,
    n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
    n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
    n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522,
    n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531,
    n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540,
    n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549,
    n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558,
    n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567,
    n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
    n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
    n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594,
    n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603,
    n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612,
    n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621,
    n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630,
    n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639,
    n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
    n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
    n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666,
    n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675,
    n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684,
    n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693,
    n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702,
    n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711,
    n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
    n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
    n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738,
    n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747,
    n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756,
    n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765,
    n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774,
    n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783,
    n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
    n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
    n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810,
    n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819,
    n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828,
    n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837,
    n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846,
    n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855,
    n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
    n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
    n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882,
    n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891,
    n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900,
    n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909,
    n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918,
    n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927,
    n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
    n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
    n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954,
    n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963,
    n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972,
    n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981,
    n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990,
    n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999,
    n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
    n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
    n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026,
    n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035,
    n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044,
    n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053,
    n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062,
    n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071,
    n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
    n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
    n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098,
    n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107,
    n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116,
    n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125,
    n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134,
    n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143,
    n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
    n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
    n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170,
    n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179,
    n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188,
    n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197,
    n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206,
    n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215,
    n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
    n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
    n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242,
    n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251,
    n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260,
    n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269,
    n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277, n15278,
    n15279, n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287,
    n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,
    n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
    n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314,
    n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323,
    n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331, n15332,
    n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341,
    n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349, n15350,
    n15351, n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359,
    n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,
    n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
    n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386,
    n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395,
    n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403, n15404,
    n15405, n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413,
    n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421, n15422,
    n15423, n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431,
    n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440,
    n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
    n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458,
    n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467,
    n15468, n15469, n15470, n15471, n15472, n15473, n15474, n15475, n15476,
    n15477, n15478, n15479, n15480, n15481, n15482, n15483, n15484, n15485,
    n15486, n15487, n15488, n15489, n15490, n15491, n15492, n15493, n15494,
    n15495, n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503,
    n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512,
    n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
    n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530,
    n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15539,
    n15540, n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548,
    n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15556, n15557,
    n15558, n15559, n15560, n15561, n15562, n15563, n15564, n15565, n15566,
    n15567, n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575,
    n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584,
    n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
    n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602,
    n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611,
    n15612, n15613, n15614, n15615, n15616, n15617, n15618, n15619, n15620,
    n15621, n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629,
    n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637, n15638,
    n15639, n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647,
    n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656,
    n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
    n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674,
    n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682, n15683,
    n15684, n15685, n15686, n15687, n15688, n15689, n15690, n15691, n15692,
    n15693, n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701,
    n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709, n15710,
    n15711, n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719,
    n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728,
    n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
    n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746,
    n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754, n15755,
    n15756, n15757, n15758, n15759, n15760, n15761, n15762, n15763, n15764,
    n15765, n15766, n15767, n15768, n15769, n15770, n15771, n15772, n15773,
    n15774, n15775, n15776, n15777, n15778, n15779, n15780, n15781, n15782,
    n15783, n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791,
    n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800,
    n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
    n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818,
    n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826, n15827,
    n15828, n15829, n15830, n15831, n15832, n15833, n15834, n15835, n15836,
    n15837, n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845,
    n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853, n15854,
    n15855, n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863,
    n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872,
    n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
    n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890,
    n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898, n15899,
    n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907, n15908,
    n15909, n15910, n15911, n15912, n15913, n15914, n15915, n15916, n15917,
    n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925, n15926,
    n15927, n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935,
    n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944,
    n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
    n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962,
    n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970, n15971,
    n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15979, n15980,
    n15981, n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15989,
    n15990, n15991, n15992, n15993, n15994, n15995, n15996, n15997, n15998,
    n15999, n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007,
    n16008, n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016,
    n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
    n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034,
    n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042, n16043,
    n16044, n16045, n16046, n16047, n16048, n16049, n16050, n16051, n16052,
    n16053, n16054, n16055, n16056, n16057, n16058, n16059, n16060, n16061,
    n16062, n16063, n16064, n16065, n16066, n16067, n16068, n16069, n16070,
    n16071, n16072, n16073, n16074, n16075, n16076, n16077, n16078, n16079,
    n16080, n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088,
    n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
    n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106,
    n16107, n16108, n16109, n16110, n16111, n16112, n16113, n16114, n16115,
    n16116, n16117, n16118, n16119, n16120, n16121, n16122, n16123, n16124,
    n16125, n16126, n16127, n16128, n16129, n16130, n16131, n16132, n16133,
    n16134, n16135, n16136, n16137, n16138, n16139, n16140, n16141, n16142,
    n16143, n16144, n16145, n16146, n16147, n16148, n16149, n16150, n16151,
    n16152, n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160,
    n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
    n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178,
    n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186, n16187,
    n16188, n16189, n16190, n16191, n16192, n16193, n16194, n16195, n16196,
    n16197, n16198, n16199, n16200, n16201, n16202, n16203, n16204, n16205,
    n16206, n16207, n16208, n16209, n16210, n16211, n16212, n16213, n16214,
    n16215, n16216, n16217, n16218, n16219, n16220, n16221, n16222, n16223,
    n16224, n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232,
    n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
    n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16250,
    n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258, n16259,
    n16260, n16261, n16262, n16263, n16264, n16265, n16266, n16267, n16268,
    n16269, n16270, n16271, n16272, n16273, n16274, n16275, n16276, n16277,
    n16278, n16279, n16280, n16281, n16282, n16283, n16284, n16285, n16286,
    n16287, n16288, n16289, n16290, n16291, n16292, n16293, n16294, n16295,
    n16296, n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304,
    n16305, n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
    n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322,
    n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330, n16331,
    n16332, n16333, n16334, n16335, n16336, n16337, n16338, n16339, n16340,
    n16341, n16342, n16343, n16344, n16345, n16346, n16347, n16348, n16349,
    n16350, n16351, n16352, n16353, n16354, n16355, n16356, n16357, n16358,
    n16359, n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16367,
    n16368, n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376,
    n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
    n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394,
    n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402, n16403,
    n16404, n16405, n16406, n16407, n16408, n16409, n16410, n16411, n16412,
    n16413, n16414, n16415, n16416, n16417, n16418, n16419, n16420, n16421,
    n16422, n16423, n16424, n16425, n16426, n16427, n16428, n16429, n16430,
    n16431, n16432, n16433, n16434, n16435, n16436, n16437, n16438, n16439,
    n16440, n16441, n16442, n16443, n16444, n16445, n16446, n16447, n16448,
    n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
    n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465, n16466,
    n16467, n16468, n16469, n16470, n16471, n16472, n16473, n16474, n16475,
    n16476, n16477, n16478, n16479, n16480, n16481, n16482, n16483, n16484,
    n16485, n16486, n16487, n16488, n16489, n16490, n16491, n16492, n16493,
    n16494, n16495, n16496, n16497, n16498, n16499, n16500, n16501, n16502,
    n16503, n16504, n16505, n16506, n16507, n16508, n16509, n16510, n16511,
    n16512, n16513, n16514, n16515, n16516, n16517, n16518, n16519, n16520,
    n16521, n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
    n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537, n16538,
    n16539, n16540, n16541, n16542, n16543, n16544, n16545, n16546, n16547,
    n16548, n16549, n16550, n16551, n16552, n16553, n16554, n16555, n16556,
    n16557, n16558, n16559, n16560, n16561, n16562, n16563, n16564, n16565,
    n16566, n16567, n16568, n16569, n16570, n16571, n16572, n16573, n16574,
    n16575, n16576, n16577, n16578, n16579, n16580, n16581, n16582, n16583,
    n16584, n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592,
    n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
    n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610,
    n16611, n16612, n16613, n16614, n16615, n16616, n16617, n16618, n16619,
    n16620, n16621, n16622, n16623, n16624, n16625, n16626, n16627, n16628,
    n16629, n16630, n16631, n16632, n16633, n16634, n16635, n16636, n16637,
    n16638, n16639, n16640, n16641, n16642, n16643, n16644, n16645, n16646,
    n16647, n16648, n16649, n16650, n16651, n16652, n16653, n16654, n16655,
    n16656, n16657, n16658, n16659, n16660, n16661, n16662, n16663, n16664,
    n16665, n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
    n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681, n16682,
    n16683, n16684, n16685, n16686, n16687, n16688, n16689, n16690, n16691,
    n16692, n16693, n16694, n16695, n16696, n16697, n16698, n16699, n16700,
    n16701, n16702, n16703, n16704, n16705, n16706, n16707, n16708, n16709,
    n16710, n16711, n16712, n16713, n16714, n16715, n16716, n16717, n16718,
    n16719, n16720, n16721, n16722, n16723, n16724, n16725, n16726, n16727,
    n16728, n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736,
    n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
    n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753, n16754,
    n16755, n16756, n16757, n16758, n16759, n16760, n16761, n16762, n16763,
    n16764, n16765, n16766, n16767, n16768, n16769, n16770, n16771, n16772,
    n16773, n16774, n16775, n16776, n16777, n16778, n16779, n16780, n16781,
    n16782, n16783, n16784, n16785, n16786, n16787, n16788, n16789, n16790,
    n16791, n16792, n16793, n16794, n16795, n16796, n16797, n16798, n16799,
    n16800, n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808,
    n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
    n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825, n16826,
    n16827, n16828, n16829, n16830, n16831, n16832, n16833, n16834, n16835,
    n16836, n16837, n16838, n16839, n16840, n16841, n16842, n16843, n16844,
    n16845, n16846, n16847, n16848, n16849, n16850, n16851, n16852, n16853,
    n16854, n16855, n16856, n16857, n16858, n16859, n16860, n16861, n16862,
    n16863, n16864, n16865, n16866, n16867, n16868, n16869, n16870, n16871,
    n16872, n16873, n16874, n16875, n16876, n16877, n16878, n16879, n16880,
    n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
    n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897, n16898,
    n16899, n16900, n16901, n16902, n16903, n16904, n16905, n16906, n16907,
    n16908, n16909, n16910, n16911, n16912, n16913, n16914, n16915, n16916,
    n16917, n16918, n16919, n16920, n16921, n16922, n16923, n16924, n16925,
    n16926, n16927, n16928, n16929, n16930, n16931, n16932, n16933, n16934,
    n16935, n16936, n16937, n16938, n16939, n16940, n16941, n16942, n16943,
    n16944, n16945, n16946, n16947, n16948, n16949, n16950, n16951, n16952,
    n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
    n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969, n16970,
    n16971, n16972, n16973, n16974, n16975, n16976, n16977, n16978, n16979,
    n16980, n16981, n16982, n16983, n16984, n16985, n16986, n16987, n16988,
    n16989, n16990, n16991, n16992, n16993, n16994, n16995, n16996, n16997,
    n16998, n16999, n17000, n17001, n17002, n17003, n17004, n17005, n17006,
    n17007, n17008, n17009, n17010, n17011, n17012, n17013, n17014, n17015,
    n17016, n17017, n17018, n17019, n17020, n17021, n17022, n17023, n17024,
    n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
    n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041, n17042,
    n17043, n17044, n17045, n17046, n17047, n17048, n17049, n17050, n17051,
    n17052, n17053, n17054, n17055, n17056, n17057, n17058, n17059, n17060,
    n17061, n17062, n17063, n17064, n17065, n17066, n17067, n17068, n17069,
    n17070, n17071, n17072, n17073, n17074, n17075, n17076, n17077, n17078,
    n17079, n17080, n17081, n17082, n17083, n17084, n17085, n17086, n17087,
    n17088, n17089, n17090, n17091, n17092, n17093, n17094, n17095, n17096,
    n17097, n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
    n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113, n17114,
    n17115, n17116, n17117, n17118, n17119, n17120, n17121, n17122, n17123,
    n17124, n17125, n17126, n17127, n17128, n17129, n17130, n17131, n17132,
    n17133, n17134, n17135, n17136, n17137, n17138, n17139, n17140, n17141,
    n17142, n17143, n17144, n17145, n17146, n17147, n17148, n17149, n17150,
    n17151, n17152, n17153, n17154, n17155, n17156, n17157, n17158, n17159,
    n17160, n17161, n17162, n17163, n17164, n17165, n17166, n17167, n17168,
    n17169, n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
    n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185, n17186,
    n17187, n17188, n17189, n17190, n17191, n17192, n17193, n17194, n17195,
    n17196, n17197, n17198, n17199, n17200, n17201, n17202, n17203, n17204,
    n17205, n17206, n17207, n17208, n17209, n17210, n17211, n17212, n17213,
    n17214, n17215, n17216, n17217, n17218, n17219, n17220, n17221, n17222,
    n17223, n17224, n17225, n17226, n17227, n17228, n17229, n17230, n17231,
    n17232, n17233, n17234, n17235, n17236, n17237, n17238, n17239, n17240,
    n17241, n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
    n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257, n17258,
    n17259, n17260, n17261, n17262, n17263, n17264, n17265, n17266, n17267,
    n17268, n17269, n17270, n17271, n17272, n17273, n17274, n17275, n17276,
    n17277, n17278, n17279, n17280, n17281, n17282, n17283, n17284, n17285,
    n17286, n17287, n17288, n17289, n17290, n17291, n17292, n17293, n17294,
    n17295, n17296, n17297, n17298, n17299, n17300, n17301, n17302, n17303,
    n17304, n17305, n17306, n17307, n17308, n17309, n17310, n17311, n17312,
    n17313, n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
    n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329, n17330,
    n17331, n17332, n17333, n17334, n17335, n17336, n17337, n17338, n17339,
    n17340, n17341, n17342, n17343, n17344, n17345, n17346, n17347, n17348,
    n17349, n17350, n17351, n17352, n17353, n17354, n17355, n17356, n17357,
    n17358, n17359, n17360, n17361, n17362, n17363, n17364, n17365, n17366,
    n17367, n17368, n17369, n17370, n17371, n17372, n17373, n17374, n17375,
    n17376, n17377, n17378, n17379, n17380, n17381, n17382, n17383, n17384,
    n17385, n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
    n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401, n17402,
    n17403, n17404, n17405, n17406, n17407, n17408, n17409, n17410, n17411,
    n17412, n17413, n17414, n17415, n17416, n17417, n17418, n17419, n17420,
    n17421, n17422, n17423, n17424, n17425, n17426, n17427, n17428, n17429,
    n17430, n17431, n17432, n17433, n17434, n17435, n17436, n17437, n17438,
    n17439, n17440, n17441, n17442, n17443, n17444, n17445, n17446, n17447,
    n17448, n17449, n17450, n17451, n17452, n17453, n17454, n17455, n17456,
    n17457, n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
    n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473, n17474,
    n17475, n17476, n17477, n17478, n17479, n17480, n17481, n17482, n17483,
    n17484, n17485, n17486, n17487, n17488, n17489, n17490, n17491, n17492,
    n17493, n17494, n17495, n17496, n17497, n17498, n17499, n17500, n17501,
    n17502, n17503, n17504, n17505, n17506, n17507, n17508, n17509, n17510,
    n17511, n17512, n17513, n17514, n17515, n17516, n17517, n17518, n17519,
    n17520, n17521, n17522, n17523, n17524, n17525, n17526, n17527, n17528,
    n17529, n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
    n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545, n17546,
    n17547, n17548, n17549, n17550, n17551, n17552, n17553, n17554, n17555,
    n17556, n17557, n17558, n17559, n17560, n17561, n17562, n17563, n17564,
    n17565, n17566, n17567, n17568, n17569, n17570, n17571, n17572, n17573,
    n17574, n17575, n17576, n17577, n17578, n17579, n17580, n17581, n17582,
    n17583, n17584, n17585, n17586, n17587, n17588, n17589, n17590, n17591,
    n17592, n17593, n17594, n17595, n17596, n17597, n17598, n17599, n17600,
    n17601, n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
    n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617, n17618,
    n17619, n17620, n17621, n17622, n17623, n17624, n17625, n17626, n17627,
    n17628, n17629, n17630, n17631, n17632, n17633, n17634, n17635, n17636,
    n17637, n17638, n17639, n17640, n17641, n17642, n17643, n17644, n17645,
    n17646, n17647, n17648, n17649, n17650, n17651, n17652, n17653, n17654,
    n17655, n17656, n17657, n17658, n17659, n17660, n17661, n17662, n17663,
    n17664, n17665, n17666, n17667, n17668, n17669, n17670, n17671, n17672,
    n17673, n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
    n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689, n17690,
    n17691, n17692, n17693, n17694, n17695, n17696, n17697, n17698, n17699,
    n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707, n17708,
    n17709, n17710, n17711, n17712, n17713, n17714, n17715, n17716, n17717,
    n17718, n17719, n17720, n17721, n17722, n17723, n17724, n17725, n17726,
    n17727, n17728, n17729, n17730, n17731, n17732, n17733, n17734, n17735,
    n17736, n17737, n17738, n17739, n17740, n17741, n17742, n17743, n17744,
    n17745, n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
    n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761, n17762,
    n17763, n17764, n17765, n17766, n17767, n17768, n17769, n17770, n17771,
    n17772, n17773, n17774, n17775, n17776, n17777, n17778, n17779, n17780,
    n17781, n17782, n17783, n17784, n17785, n17786, n17787, n17788, n17789,
    n17790, n17791, n17792, n17793, n17794, n17795, n17796, n17797, n17798,
    n17799, n17800, n17801, n17802, n17803, n17804, n17805, n17806, n17807,
    n17808, n17809, n17810, n17811, n17812, n17813, n17814, n17815, n17816,
    n17817, n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
    n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833, n17834,
    n17835, n17836, n17837, n17838, n17839, n17840, n17841, n17842, n17843,
    n17844, n17845, n17846, n17847, n17848, n17849, n17850, n17851, n17852,
    n17853, n17854, n17855, n17856, n17857, n17858, n17859, n17860, n17861,
    n17862, n17863, n17864, n17865, n17866, n17867, n17868, n17869, n17870,
    n17871, n17872, n17873, n17874, n17875, n17876, n17877, n17878, n17879,
    n17880, n17881, n17882, n17883, n17884, n17885, n17886, n17887, n17888,
    n17889, n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
    n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905, n17906,
    n17907, n17908, n17909, n17910, n17911, n17912, n17913, n17914, n17915,
    n17916, n17917, n17918, n17919, n17920, n17921, n17922, n17923, n17924,
    n17925, n17926, n17927, n17928, n17929, n17930, n17931, n17932, n17933,
    n17934, n17935, n17936, n17937, n17938, n17939, n17940, n17941, n17942,
    n17943, n17944, n17945, n17946, n17947, n17948, n17949, n17950, n17951,
    n17952, n17953, n17954, n17955, n17956, n17957, n17958, n17959, n17960,
    n17961, n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
    n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977, n17978,
    n17979, n17980, n17981, n17982, n17983, n17984, n17985, n17986, n17987,
    n17988, n17989, n17990, n17991, n17992, n17993, n17994, n17995, n17996,
    n17997, n17998, n17999, n18000, n18001, n18002, n18003, n18004, n18005,
    n18006, n18007, n18008, n18009, n18010, n18011, n18012, n18013, n18014,
    n18015, n18016, n18017, n18018, n18019, n18020, n18021, n18022, n18023,
    n18024, n18025, n18026, n18027, n18028, n18029, n18030, n18031, n18032,
    n18033, n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
    n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049, n18050,
    n18051, n18052, n18053, n18054, n18055, n18056, n18057, n18058, n18059,
    n18060, n18061, n18062, n18063, n18064, n18065, n18066, n18067, n18068,
    n18069, n18070, n18071, n18072, n18073, n18074, n18075, n18076, n18077,
    n18078, n18079, n18080, n18081, n18082, n18083, n18084, n18085, n18086,
    n18087, n18088, n18089, n18090, n18091, n18092, n18093, n18094, n18095,
    n18096, n18097, n18098, n18099, n18100, n18101, n18102, n18103, n18104,
    n18105, n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
    n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121, n18122,
    n18123, n18124, n18125, n18126, n18127, n18128, n18129, n18130, n18131,
    n18132, n18133, n18134, n18135, n18136, n18137, n18138, n18139, n18140,
    n18141, n18142, n18143, n18144, n18145, n18146, n18147, n18148, n18149,
    n18150, n18151, n18152, n18153, n18154, n18155, n18156, n18157, n18158,
    n18159, n18160, n18161, n18162, n18163, n18164, n18165, n18166, n18167,
    n18168, n18169, n18170, n18171, n18172, n18173, n18174, n18175, n18176,
    n18177, n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
    n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193, n18194,
    n18195, n18196, n18197, n18198, n18199, n18200, n18201, n18202, n18203,
    n18204, n18205, n18206, n18207, n18208, n18209, n18210, n18211, n18212,
    n18213, n18214, n18215, n18216, n18217, n18218, n18219, n18220, n18221,
    n18222, n18223, n18224, n18225, n18226, n18227, n18228, n18229, n18230,
    n18231, n18232, n18233, n18234, n18235, n18236, n18237, n18238, n18239,
    n18240, n18241, n18242, n18243, n18244, n18245, n18246, n18247, n18248,
    n18249, n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
    n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265, n18266,
    n18267, n18268, n18269, n18270, n18271, n18272, n18273, n18274, n18275,
    n18276, n18277, n18278, n18279, n18280, n18281, n18282, n18283, n18284,
    n18285, n18286, n18287, n18288, n18289, n18290, n18291, n18292, n18293,
    n18294, n18295, n18296, n18297, n18298, n18299, n18300, n18301, n18302,
    n18303, n18304, n18305, n18306, n18307, n18308, n18309, n18310, n18311,
    n18312, n18313, n18314, n18315, n18316, n18317, n18318, n18319, n18320,
    n18321, n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
    n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337, n18338,
    n18339, n18340, n18341, n18342, n18343, n18344, n18345, n18346, n18347,
    n18348, n18349, n18350, n18351, n18352, n18353, n18354, n18355, n18356,
    n18357, n18358, n18359, n18360, n18361, n18362, n18363, n18364, n18365,
    n18366, n18367, n18368, n18369, n18370, n18371, n18372, n18373, n18374,
    n18375, n18376, n18377, n18378, n18379, n18380, n18381, n18382, n18383,
    n18384, n18385, n18386, n18387, n18388, n18389, n18390, n18391, n18392,
    n18393, n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
    n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409, n18410,
    n18411, n18412, n18413, n18414, n18415, n18416, n18417, n18418, n18419,
    n18420, n18421, n18422, n18423, n18424, n18425, n18426, n18427, n18428,
    n18429, n18430, n18431, n18432, n18433, n18434, n18435, n18436, n18437,
    n18438, n18439, n18440, n18441, n18442, n18443, n18444, n18445, n18446,
    n18447, n18448, n18449, n18450, n18451, n18452, n18453, n18454, n18455,
    n18456, n18457, n18458, n18459, n18460, n18461, n18462, n18463, n18464,
    n18465, n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
    n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481, n18482,
    n18483, n18484, n18485, n18486, n18487, n18488, n18489, n18490, n18491,
    n18492, n18493, n18494, n18495, n18496, n18497, n18498, n18499, n18500,
    n18501, n18502, n18503, n18504, n18505, n18506, n18507, n18508, n18509,
    n18510, n18511, n18512, n18513, n18514, n18515, n18516, n18517, n18518,
    n18519, n18520, n18521, n18522, n18523, n18524, n18525, n18526, n18527,
    n18528, n18529, n18530, n18531, n18532, n18533, n18534, n18535, n18536,
    n18537, n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
    n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553, n18554,
    n18555, n18556, n18557, n18558, n18559, n18560, n18561, n18562, n18563,
    n18564, n18565, n18566, n18567, n18568, n18569, n18570, n18571, n18572,
    n18573, n18574, n18575, n18576, n18577, n18578, n18579, n18580, n18581,
    n18582, n18583, n18584, n18585, n18586, n18587, n18588, n18589, n18590,
    n18591, n18592, n18593, n18594, n18595, n18596, n18597, n18598, n18599,
    n18600, n18601, n18602, n18603, n18604, n18605, n18606, n18607, n18608,
    n18609, n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617,
    n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625, n18626,
    n18627, n18628, n18629, n18630, n18631, n18632, n18633, n18634, n18635,
    n18636, n18637, n18638, n18639, n18640, n18641, n18642, n18643, n18644,
    n18645, n18646, n18647, n18648, n18649, n18650, n18651, n18652, n18653,
    n18654, n18655, n18656, n18657, n18658, n18659, n18660, n18661, n18662,
    n18663, n18664, n18665, n18666, n18667, n18668, n18669, n18670, n18671,
    n18672, n18673, n18674, n18675, n18676, n18677, n18678, n18679, n18680,
    n18681, n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
    n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697, n18698,
    n18699, n18700, n18701, n18702, n18703, n18704, n18705, n18706, n18707,
    n18708, n18709, n18710, n18711, n18712, n18713, n18714, n18715, n18716,
    n18717, n18718, n18719, n18720, n18721, n18722, n18723, n18724, n18725,
    n18726, n18727, n18728, n18729, n18730, n18731, n18732, n18733, n18734,
    n18735, n18736, n18737, n18738, n18739, n18740, n18741, n18742, n18743,
    n18744, n18745, n18746, n18747, n18748, n18749, n18750, n18751, n18752,
    n18753, n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
    n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769, n18770,
    n18771, n18772, n18773, n18774, n18775, n18776, n18777, n18778, n18779,
    n18780, n18781, n18782, n18783, n18784, n18785, n18786, n18787, n18788,
    n18789, n18790, n18791, n18792, n18793, n18794, n18795, n18796, n18797,
    n18798, n18799, n18800, n18801, n18802, n18803, n18804, n18805, n18806,
    n18807, n18808, n18809, n18810, n18811, n18812, n18813, n18814, n18815,
    n18816, n18817, n18818, n18819, n18820, n18821, n18822, n18823, n18824,
    n18825, n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
    n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841, n18842,
    n18843, n18844, n18845, n18846, n18847, n18848, n18849, n18850, n18851,
    n18852, n18853, n18854, n18855, n18856, n18857, n18858, n18859, n18860,
    n18861, n18862, n18863, n18864, n18865, n18866, n18867, n18868, n18869,
    n18870, n18871, n18872, n18873, n18874, n18875, n18876, n18877, n18878,
    n18879, n18880, n18881, n18882, n18883, n18884, n18885, n18886, n18887,
    n18888, n18889, n18890, n18891, n18892, n18893, n18894, n18895, n18896,
    n18897, n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905,
    n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913, n18914,
    n18915, n18916, n18917, n18918, n18919, n18920, n18921, n18922, n18923,
    n18924, n18925, n18926, n18927, n18928, n18929, n18930, n18931, n18932,
    n18933, n18934, n18935, n18936, n18937, n18938, n18939, n18940, n18941,
    n18942, n18943, n18944, n18945, n18946, n18947, n18948, n18949, n18950,
    n18951, n18952, n18953, n18954, n18955, n18956, n18957, n18958, n18959,
    n18960, n18961, n18962, n18963, n18964, n18965, n18966, n18967, n18968,
    n18969, n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,
    n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985, n18986,
    n18987, n18988, n18989, n18990, n18991, n18992, n18993, n18994, n18995,
    n18996, n18997, n18998, n18999, n19000, n19001, n19002, n19003, n19004,
    n19005, n19006, n19007, n19008, n19009, n19010, n19011, n19012, n19013,
    n19014, n19015, n19016, n19017, n19018, n19019, n19020, n19021, n19022,
    n19023, n19024, n19025, n19026, n19027, n19028, n19029, n19030, n19031,
    n19032, n19033, n19034, n19035, n19036, n19037, n19038, n19039, n19040,
    n19041, n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
    n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057, n19058,
    n19059, n19060, n19061, n19062, n19063, n19064, n19065, n19066, n19067,
    n19068, n19069, n19070, n19071, n19072, n19073, n19074, n19075, n19076,
    n19077, n19078, n19079, n19080, n19081, n19082, n19083, n19084, n19085,
    n19086, n19087, n19088, n19089, n19090, n19091, n19092, n19093, n19094,
    n19095, n19096, n19097, n19098, n19099, n19100, n19101, n19102, n19103,
    n19104, n19105, n19106, n19107, n19108, n19109, n19110, n19111, n19112,
    n19113, n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
    n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129, n19130,
    n19131, n19132, n19133, n19134, n19135, n19136, n19137, n19138, n19139,
    n19140, n19141, n19142, n19143, n19144, n19145, n19146, n19147, n19148,
    n19149, n19150, n19151, n19152, n19153, n19154, n19155, n19156, n19157,
    n19158, n19159, n19160, n19161, n19162, n19163, n19164, n19165, n19166,
    n19167, n19168, n19169, n19170, n19171, n19172, n19173, n19174, n19175,
    n19176, n19177, n19178, n19179, n19180, n19181, n19182, n19183, n19184,
    n19185, n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
    n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201, n19202,
    n19203, n19204, n19205, n19206, n19207, n19208, n19209, n19210, n19211,
    n19212, n19213, n19214, n19215, n19216, n19217, n19218, n19219, n19220,
    n19221, n19222, n19223, n19224, n19225, n19226, n19227, n19228, n19229,
    n19230, n19231, n19232, n19233, n19234, n19235, n19236, n19237, n19238,
    n19239, n19240, n19241, n19242, n19243, n19244, n19245, n19246, n19247,
    n19248, n19249, n19250, n19251, n19252, n19253, n19254, n19255, n19256,
    n19257, n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
    n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273, n19274,
    n19275, n19276, n19277, n19278, n19279, n19280, n19281, n19282, n19283,
    n19284, n19285, n19286, n19287, n19288, n19289, n19290, n19291, n19292,
    n19293, n19294, n19295, n19296, n19297, n19298, n19299, n19300, n19301,
    n19302, n19303, n19304, n19305, n19306, n19307, n19308, n19309, n19310,
    n19311, n19312, n19313, n19314, n19315, n19316, n19317, n19318, n19319,
    n19320, n19321, n19322, n19323, n19324, n19325, n19326, n19327, n19328,
    n19329, n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
    n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345, n19346,
    n19347, n19348, n19349, n19350, n19351, n19352, n19353, n19354, n19355,
    n19356, n19357, n19358, n19359, n19360, n19361, n19362, n19363, n19364,
    n19365, n19366, n19367, n19368, n19369, n19370, n19371, n19372, n19373,
    n19374, n19375, n19376, n19377, n19378, n19379, n19380, n19381, n19382,
    n19383, n19384, n19385, n19386, n19387, n19388, n19389, n19390, n19391,
    n19392, n19393, n19394, n19395, n19396, n19397, n19398, n19399, n19400,
    n19401, n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
    n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417, n19418,
    n19419, n19420, n19421, n19422, n19423, n19424, n19425, n19426, n19427,
    n19428, n19429, n19430, n19431, n19432, n19433, n19434, n19435, n19436,
    n19437, n19438, n19439, n19440, n19441, n19442, n19443, n19444, n19445,
    n19446, n19447, n19448, n19449, n19450, n19451, n19452, n19453, n19454,
    n19455, n19456, n19457, n19458, n19459, n19460, n19461, n19462, n19463,
    n19464, n19465, n19466, n19467, n19468, n19469, n19470, n19471, n19472,
    n19473, n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
    n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489, n19490,
    n19491, n19492, n19493, n19494, n19495, n19496, n19497, n19498, n19499,
    n19500, n19501, n19502, n19503, n19504, n19505, n19506, n19507, n19508,
    n19509, n19510, n19511, n19512, n19513, n19514, n19515, n19516, n19517,
    n19518, n19519, n19520, n19521, n19522, n19523, n19524, n19525, n19526,
    n19527, n19528, n19529, n19530, n19531, n19532, n19533, n19534, n19535,
    n19536, n19537, n19538, n19539, n19540, n19541, n19542, n19543, n19544,
    n19545, n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
    n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561, n19562,
    n19563, n19564, n19565, n19566, n19567, n19568, n19569, n19570, n19571,
    n19572, n19573, n19574, n19575, n19576, n19577, n19578, n19579, n19580,
    n19581, n19582, n19583, n19584, n19585, n19586, n19587, n19588, n19589,
    n19590, n19591, n19592, n19593, n19594, n19595, n19596, n19597, n19598,
    n19599, n19600, n19601, n19602, n19603, n19604, n19605, n19606, n19607,
    n19608, n19609, n19610, n19611, n19612, n19613, n19614, n19615, n19616,
    n19617, n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
    n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633, n19634,
    n19635, n19636, n19637, n19638, n19639, n19640, n19641, n19642, n19643,
    n19644, n19645, n19646, n19647, n19648, n19649, n19650, n19651, n19652,
    n19653, n19654, n19655, n19656, n19657, n19658, n19659, n19660, n19661,
    n19662, n19663, n19664, n19665, n19666, n19667, n19668, n19669, n19670,
    n19671, n19672, n19673, n19674, n19675, n19676, n19677, n19678, n19679,
    n19680, n19681, n19682, n19683, n19684, n19685, n19686, n19687, n19688,
    n19689, n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
    n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705, n19706,
    n19707, n19708, n19709, n19710, n19711, n19712, n19713, n19714, n19715,
    n19716, n19717, n19718, n19719, n19720, n19721, n19722, n19723, n19724,
    n19725, n19726, n19727, n19728, n19729, n19730, n19731, n19732, n19733,
    n19734, n19735, n19736, n19737, n19738, n19739, n19740, n19741, n19742,
    n19743, n19744, n19745, n19746, n19747, n19748, n19749, n19750, n19751,
    n19752, n19753, n19754, n19755, n19756, n19757, n19758, n19759, n19760,
    n19761, n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769,
    n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777, n19778,
    n19779, n19780, n19781, n19782, n19783, n19784, n19785, n19786, n19787,
    n19788, n19789, n19790, n19791, n19792, n19793, n19794, n19795, n19796,
    n19797, n19798, n19799, n19800, n19801, n19802, n19803, n19804, n19805,
    n19806, n19807, n19808, n19809, n19810, n19811, n19812, n19813, n19814,
    n19815, n19816, n19817, n19818, n19819, n19820, n19821, n19822, n19823,
    n19824, n19825, n19826, n19827, n19828, n19829, n19830, n19831, n19832,
    n19833, n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841,
    n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849, n19850,
    n19851, n19852, n19853, n19854, n19855, n19856, n19857, n19858, n19859,
    n19860, n19861, n19862, n19863, n19864, n19865, n19866, n19867, n19868,
    n19869, n19870, n19871, n19872, n19873, n19874, n19875, n19876, n19877,
    n19878, n19879, n19880, n19881, n19882, n19883, n19884, n19885, n19886,
    n19887, n19888, n19889, n19890, n19891, n19892, n19893, n19894, n19895,
    n19896, n19897, n19898, n19899, n19900, n19901, n19902, n19903, n19904,
    n19905, n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913,
    n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921, n19922,
    n19923, n19924, n19925, n19926, n19927, n19928, n19929, n19930, n19931,
    n19932, n19933, n19934, n19935, n19936, n19937, n19938, n19939, n19940,
    n19941, n19942, n19943, n19944, n19945, n19946, n19947, n19948, n19949,
    n19950, n19951, n19952, n19953, n19954, n19955, n19956, n19957, n19958,
    n19959, n19960, n19961, n19962, n19963, n19964, n19965, n19966, n19967,
    n19968, n19969, n19970, n19971, n19972, n19973, n19974, n19975, n19976,
    n19977, n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985,
    n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993, n19994,
    n19995, n19996, n19997, n19998, n19999, n20000, n20001, n20002, n20003,
    n20004, n20005, n20006, n20007, n20008, n20009, n20010, n20011, n20012,
    n20013, n20014, n20015, n20016, n20017, n20018, n20019, n20020, n20021,
    n20022, n20023, n20024, n20025, n20026, n20027, n20028, n20029, n20030,
    n20031, n20032, n20033, n20034, n20035, n20036, n20037, n20038, n20039,
    n20040, n20041, n20042, n20043, n20044, n20045, n20046, n20047, n20048,
    n20049, n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057,
    n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065, n20066,
    n20067, n20068, n20069, n20070, n20071, n20072, n20073, n20074, n20075,
    n20076, n20077, n20078, n20079, n20080, n20081, n20082, n20083, n20084,
    n20085, n20086, n20087, n20088, n20089, n20090, n20091, n20092, n20093,
    n20094, n20095, n20096, n20097, n20098, n20099, n20100, n20101, n20102,
    n20103, n20104, n20105, n20106, n20107, n20108, n20109, n20110, n20111,
    n20112, n20113, n20114, n20115, n20116, n20117, n20118, n20119, n20120,
    n20121, n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129,
    n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137, n20138,
    n20139, n20140, n20141, n20142, n20143, n20144, n20145, n20146, n20147,
    n20148, n20149, n20150, n20151, n20152, n20153, n20154, n20155, n20156,
    n20157, n20158, n20159, n20160, n20161, n20162, n20163, n20164, n20165,
    n20166, n20167, n20168, n20169, n20170, n20171, n20172, n20173, n20174,
    n20175, n20176, n20177, n20178, n20179, n20180, n20181, n20182, n20183,
    n20184, n20185, n20186, n20187, n20188, n20189, n20190, n20191, n20192,
    n20193, n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201,
    n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209, n20210,
    n20211, n20212, n20213, n20214, n20215, n20216, n20217, n20218, n20219,
    n20220, n20221, n20222, n20223, n20224, n20225, n20226, n20227, n20228,
    n20229, n20230, n20231, n20232, n20233, n20234, n20235, n20236, n20237,
    n20238, n20239, n20240, n20241, n20242, n20243, n20244, n20245, n20246,
    n20247, n20248, n20249, n20250, n20251, n20252, n20253, n20254, n20255,
    n20256, n20257, n20258, n20259, n20260, n20261, n20262, n20263, n20264,
    n20265, n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273,
    n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281, n20282,
    n20283, n20284, n20285, n20286, n20287, n20288, n20289, n20290, n20291,
    n20292, n20293, n20294, n20295, n20296, n20297, n20298, n20299, n20300,
    n20301, n20302, n20303, n20304, n20305, n20306, n20307, n20308, n20309,
    n20310, n20311, n20312, n20313, n20314, n20315, n20316, n20317, n20318,
    n20319, n20320, n20321, n20322, n20323, n20324, n20325, n20326, n20327,
    n20328, n20329, n20330, n20331, n20332, n20333, n20334, n20335, n20336,
    n20337, n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345,
    n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353, n20354,
    n20355, n20356, n20357, n20358, n20359, n20360, n20361, n20362, n20363,
    n20364, n20365, n20366, n20367, n20368, n20369, n20370, n20371, n20372,
    n20373, n20374, n20375, n20376, n20377, n20378, n20379, n20380, n20381,
    n20382, n20383, n20384, n20385, n20386, n20387, n20388, n20389, n20390,
    n20391, n20392, n20393, n20394, n20395, n20396, n20397, n20398, n20399,
    n20400, n20401, n20402, n20403, n20404, n20405, n20406, n20407, n20408,
    n20409, n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417,
    n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425, n20426,
    n20427, n20428, n20429, n20430, n20431, n20432, n20433, n20434, n20435,
    n20436, n20437, n20438, n20439, n20440, n20441, n20442, n20443, n20444,
    n20445, n20446, n20447, n20448, n20449, n20450, n20451, n20452, n20453,
    n20454, n20455, n20456, n20457, n20458, n20459, n20460, n20461, n20462,
    n20463, n20464, n20465, n20466, n20467, n20468, n20469, n20470, n20471,
    n20472, n20473, n20474, n20475, n20476, n20477, n20478, n20479, n20480,
    n20481, n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489,
    n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497, n20498,
    n20499, n20500, n20501, n20502, n20503, n20504, n20505, n20506, n20507,
    n20508, n20509, n20510, n20511, n20512, n20513, n20514, n20515, n20516,
    n20517, n20518, n20519, n20520, n20521, n20522, n20523, n20524, n20525,
    n20526, n20527, n20528, n20529, n20530, n20531, n20532, n20533, n20534,
    n20535, n20536, n20537, n20538, n20539, n20540, n20541, n20542, n20543,
    n20544, n20545, n20546, n20547, n20548, n20549, n20550, n20551, n20552,
    n20553, n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561,
    n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569, n20570,
    n20571, n20572, n20573, n20574, n20575, n20576, n20577, n20578, n20579,
    n20580, n20581, n20582, n20583, n20584, n20585, n20586, n20587, n20588,
    n20589, n20590, n20591, n20592, n20593, n20594, n20595, n20596, n20597,
    n20598, n20599, n20600, n20601, n20602, n20603, n20604, n20605, n20606,
    n20607, n20608, n20609, n20610, n20611, n20612, n20613, n20614, n20615,
    n20616, n20617, n20618, n20619, n20620, n20621, n20622, n20623, n20624,
    n20625, n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633,
    n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641, n20642,
    n20643, n20644, n20645, n20646, n20647, n20648, n20649, n20650, n20651,
    n20652, n20653, n20654, n20655, n20656, n20657, n20658, n20659, n20660,
    n20661, n20662, n20663, n20664, n20665, n20666, n20667, n20668, n20669,
    n20670, n20671, n20672, n20673, n20674, n20675, n20676, n20677, n20678,
    n20679, n20680, n20681, n20682, n20683, n20684, n20685, n20686, n20687,
    n20688, n20689, n20690, n20691, n20692, n20693, n20694, n20695, n20696,
    n20697, n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705,
    n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713, n20714,
    n20715, n20716, n20717, n20718, n20719, n20720, n20721, n20722, n20723,
    n20724, n20725, n20726, n20727, n20728, n20729, n20730, n20731, n20732,
    n20733, n20734, n20735, n20736, n20737, n20738, n20739, n20740, n20741,
    n20742, n20743, n20744, n20745, n20746, n20747, n20748, n20749, n20750,
    n20751, n20752, n20753, n20754, n20755, n20756, n20757, n20758, n20759,
    n20760, n20761, n20762, n20763, n20764, n20765, n20766, n20767, n20768,
    n20769, n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777,
    n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785, n20786,
    n20787, n20788, n20789, n20790, n20791, n20792, n20793, n20794, n20795,
    n20796, n20797, n20798, n20799, n20800, n20801, n20802, n20803, n20804,
    n20805, n20806, n20807, n20808, n20809, n20810, n20811, n20812, n20813,
    n20814, n20815, n20816, n20817, n20818, n20819, n20820, n20821, n20822,
    n20823, n20824, n20825, n20826, n20827, n20828, n20829, n20830, n20831,
    n20832, n20833, n20834, n20835, n20836, n20837, n20838, n20839, n20840,
    n20841, n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849,
    n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857, n20858,
    n20859, n20860, n20861, n20862, n20863, n20864, n20865, n20866, n20867,
    n20868, n20869, n20870, n20871, n20872, n20873, n20874, n20875, n20876,
    n20877, n20878, n20879, n20880, n20881, n20882, n20883, n20884, n20885,
    n20886, n20887, n20888, n20889, n20890, n20891, n20892, n20893, n20894,
    n20895, n20896, n20897, n20898, n20899, n20900, n20901, n20902, n20903,
    n20904, n20905, n20906, n20907, n20908, n20909, n20910, n20911, n20912,
    n20913, n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921,
    n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929, n20930,
    n20931, n20932, n20933, n20934, n20935, n20936, n20937, n20938, n20939,
    n20940, n20941, n20942, n20943, n20944, n20945, n20946, n20947, n20948,
    n20949, n20950, n20951, n20952, n20953, n20954, n20955, n20956, n20957,
    n20958, n20959, n20960, n20961, n20962, n20963, n20964, n20965, n20966,
    n20967, n20968, n20969, n20970, n20971, n20972, n20973, n20974, n20975,
    n20976, n20977, n20978, n20979, n20980, n20981, n20982, n20983, n20984,
    n20985, n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993,
    n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001, n21002,
    n21003, n21004, n21005, n21006, n21007, n21008, n21009, n21010, n21011,
    n21012, n21013, n21014, n21015, n21016, n21017, n21018, n21019, n21020,
    n21021, n21022, n21023, n21024, n21025, n21026, n21027, n21028, n21029,
    n21030, n21031, n21032, n21033, n21034, n21035, n21036, n21037, n21038,
    n21039, n21040, n21041, n21042, n21043, n21044, n21045, n21046, n21047,
    n21048, n21049, n21050, n21051, n21052, n21053, n21054, n21055, n21056,
    n21057, n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065,
    n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073, n21074,
    n21075, n21076, n21077, n21078, n21079, n21080, n21081, n21082, n21083,
    n21084, n21085, n21086, n21087, n21088, n21089, n21090, n21091, n21092,
    n21093, n21094, n21095, n21096, n21097, n21098, n21099, n21100, n21101,
    n21102, n21103, n21104, n21105, n21106, n21107, n21108, n21109, n21110,
    n21111, n21112, n21113, n21114, n21115, n21116, n21117, n21118, n21119,
    n21120, n21121, n21122, n21123, n21124, n21125, n21126, n21127, n21128,
    n21129, n21130, n21131, n21132, n21133, n21134, n21135, n21136, n21137,
    n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145, n21146,
    n21147, n21148, n21149, n21150, n21151, n21152, n21153, n21154, n21155,
    n21156, n21157, n21158, n21159, n21160, n21161, n21162, n21163, n21164,
    n21165, n21166, n21167, n21168, n21169, n21170, n21171, n21172, n21173,
    n21174, n21175, n21176, n21177, n21178, n21179, n21180, n21181, n21182,
    n21183, n21184, n21185, n21186, n21187, n21188, n21189, n21190, n21191,
    n21192, n21193, n21194, n21195, n21196, n21197, n21198, n21199, n21200,
    n21201, n21202, n21203, n21204, n21205, n21206, n21207, n21208, n21209,
    n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217, n21218,
    n21219, n21220, n21221, n21222, n21223, n21224, n21225, n21226, n21227,
    n21228, n21229, n21230, n21231, n21232, n21233, n21234, n21235, n21236,
    n21237, n21238, n21239, n21240, n21241, n21242, n21243, n21244, n21245,
    n21246, n21247, n21248, n21249, n21250, n21251, n21252, n21253, n21254,
    n21255, n21256, n21257, n21258, n21259, n21260, n21261, n21262, n21263,
    n21264, n21265, n21266, n21267, n21268, n21269, n21270, n21271, n21272,
    n21273, n21274, n21275, n21276, n21277, n21278, n21279, n21280, n21281,
    n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289, n21290,
    n21291, n21292, n21293, n21294, n21295, n21296, n21297, n21298, n21299,
    n21300, n21301, n21302, n21303, n21304, n21305, n21306, n21307, n21308,
    n21309, n21310, n21311, n21312, n21313, n21314, n21315, n21316, n21317,
    n21318, n21319, n21320, n21321, n21322, n21323, n21324, n21325, n21326,
    n21327, n21328, n21329, n21330, n21331, n21332, n21333, n21334, n21335,
    n21336, n21337, n21338, n21339, n21340, n21341, n21342, n21343, n21344,
    n21345, n21346, n21347, n21348, n21349, n21350, n21351, n21352, n21353,
    n21354, n21355, n21356, n21357, n21358, n21359, n21360, n21361, n21362,
    n21363, n21364, n21365, n21366, n21367, n21368, n21369, n21370, n21371,
    n21372, n21373, n21374, n21375, n21376, n21377, n21378, n21379, n21380,
    n21381, n21382, n21383, n21384, n21385, n21386, n21387, n21388, n21389,
    n21390, n21391, n21392, n21393, n21394, n21395, n21396, n21397, n21398,
    n21399, n21400, n21401, n21402, n21403, n21404, n21405, n21406, n21407,
    n21408, n21409, n21410, n21411, n21412, n21413, n21414, n21415, n21416,
    n21417, n21418, n21419, n21420, n21421, n21422, n21423, n21424, n21425,
    n21426, n21427, n21428, n21429, n21430, n21431, n21432, n21433, n21434,
    n21435, n21436, n21437, n21438, n21439, n21440, n21441, n21442, n21443,
    n21444, n21445, n21446, n21447, n21448, n21449, n21450, n21451, n21452,
    n21453, n21454, n21455, n21456, n21457, n21458, n21459, n21460, n21461,
    n21462, n21463, n21464, n21465, n21466, n21467, n21468, n21469, n21470,
    n21471, n21472, n21473, n21474, n21475, n21476, n21477, n21478, n21479,
    n21480, n21481, n21482, n21483, n21484, n21485, n21486, n21487, n21488,
    n21489, n21490, n21491, n21492, n21493, n21494, n21495, n21496, n21497,
    n21498, n21499, n21500, n21501, n21502, n21503, n21504, n21505, n21506,
    n21507, n21508, n21509, n21510, n21511, n21512, n21513, n21514, n21515,
    n21516, n21517, n21518, n21519, n21520, n21521, n21522, n21523, n21524,
    n21525, n21526, n21527, n21528, n21529, n21530, n21531, n21532, n21533,
    n21534, n21535, n21536, n21537, n21538, n21539, n21540, n21541, n21542,
    n21543, n21544, n21545, n21546, n21547, n21548, n21549, n21550, n21551,
    n21552, n21553, n21554, n21555, n21556, n21557, n21558, n21559, n21560,
    n21561, n21562, n21563, n21564, n21565, n21566, n21567, n21568, n21569,
    n21570, n21571, n21572, n21573, n21574, n21575, n21576, n21577, n21578,
    n21579, n21580, n21581, n21582, n21583, n21584, n21585, n21586, n21587,
    n21588, n21589, n21590, n21591, n21592, n21593, n21594, n21595, n21596,
    n21597, n21598, n21599, n21600, n21601, n21602, n21603, n21604, n21605,
    n21606, n21607, n21608, n21609, n21610, n21611, n21612, n21613, n21614,
    n21615, n21616, n21617, n21618, n21619, n21620, n21621, n21622, n21623,
    n21624, n21625, n21626, n21627, n21628, n21629, n21630, n21631, n21632,
    n21633, n21634, n21635, n21636, n21637, n21638, n21639, n21640, n21641,
    n21642, n21643, n21644, n21645, n21646, n21647, n21648, n21649, n21650,
    n21651, n21652, n21653, n21654, n21655, n21656, n21657, n21658, n21659,
    n21660, n21661, n21662, n21663, n21664, n21665, n21666, n21667, n21668,
    n21669, n21670, n21671, n21672, n21673, n21674, n21675, n21676, n21677,
    n21678, n21679, n21680, n21681, n21682, n21683, n21684, n21685, n21686,
    n21687, n21688, n21689, n21690, n21691, n21692, n21693, n21694, n21695,
    n21696, n21697, n21698, n21699, n21700, n21701, n21702, n21703, n21704,
    n21705, n21706, n21707, n21708, n21709, n21710, n21711, n21712, n21713,
    n21714, n21715, n21716, n21717, n21718, n21719, n21720, n21721, n21722,
    n21723, n21724, n21725, n21726, n21727, n21728, n21729, n21730, n21731,
    n21732, n21733, n21734, n21735, n21736, n21737, n21738, n21739, n21740,
    n21741, n21742, n21743, n21744, n21745, n21746, n21747, n21748, n21749,
    n21750, n21751, n21752, n21753, n21754, n21755, n21756, n21757, n21758,
    n21759, n21760, n21761, n21762, n21763, n21764, n21765, n21766, n21767,
    n21768, n21769, n21770, n21771, n21772, n21773, n21774, n21775, n21776,
    n21777, n21778, n21779, n21780, n21781, n21782, n21783, n21784, n21785,
    n21786, n21787, n21788, n21789, n21790, n21791, n21792, n21793, n21794,
    n21795, n21796, n21797, n21798, n21799, n21800, n21801, n21802, n21803,
    n21804, n21805, n21806, n21807, n21808, n21809, n21810, n21811, n21812,
    n21813, n21814, n21815, n21816, n21817, n21818, n21819, n21820, n21821,
    n21822, n21823, n21824, n21825, n21826, n21827, n21828, n21829, n21830,
    n21831, n21832, n21833, n21834, n21835, n21836, n21837, n21838, n21839,
    n21840, n21841, n21842, n21843, n21844, n21845, n21846, n21847, n21848,
    n21849, n21850, n21851, n21852, n21853, n21854, n21855, n21856, n21857,
    n21858, n21859, n21860, n21861, n21862, n21863, n21864, n21865, n21866,
    n21867, n21868, n21869, n21870, n21871, n21872, n21873, n21874, n21875,
    n21876, n21877, n21878, n21879, n21880, n21881, n21882, n21883, n21884,
    n21885, n21886, n21887, n21888, n21889, n21890, n21891, n21892, n21893,
    n21894, n21895, n21896, n21897, n21898, n21899, n21900, n21901, n21902,
    n21903, n21904, n21905, n21906, n21907, n21908, n21909, n21910, n21911,
    n21912, n21913, n21914, n21915, n21916, n21917, n21918, n21919, n21920,
    n21921, n21922, n21923, n21924, n21925, n21926, n21927, n21928, n21929,
    n21930, n21931, n21932, n21933, n21934, n21935, n21936, n21937, n21938,
    n21939, n21940, n21941, n21942, n21943, n21944, n21945, n21946, n21947,
    n21948, n21949, n21950, n21951, n21952, n21953, n21954, n21955, n21956,
    n21957, n21958, n21959, n21960, n21961, n21962, n21963, n21964, n21965,
    n21966, n21967, n21968, n21969, n21970, n21971, n21972, n21973, n21974,
    n21975, n21976, n21977, n21978, n21979, n21980, n21981, n21982, n21983,
    n21984, n21985, n21986, n21987, n21988, n21989, n21990, n21991, n21992,
    n21993, n21994, n21995, n21996, n21997, n21998, n21999, n22000, n22001,
    n22002, n22003, n22004, n22005, n22006, n22007, n22008, n22009, n22010,
    n22011, n22012, n22013, n22014, n22015, n22016, n22017, n22018, n22019,
    n22020, n22021, n22022, n22023, n22024, n22025, n22026, n22027, n22028,
    n22029, n22030, n22031, n22032, n22033, n22034, n22035, n22036, n22037,
    n22038, n22039, n22040, n22041, n22042, n22043, n22044, n22045, n22046,
    n22047, n22048, n22049, n22050, n22051, n22052, n22053, n22054, n22055,
    n22056, n22057, n22058, n22059, n22060, n22061, n22062, n22063, n22064,
    n22065, n22066, n22067, n22068, n22069, n22070, n22071, n22072, n22073,
    n22074, n22075, n22076, n22077, n22078, n22079, n22080, n22081, n22082,
    n22083, n22084, n22085, n22086, n22087, n22088, n22089, n22090, n22091,
    n22092, n22093, n22094, n22095, n22096, n22097, n22098, n22099, n22100,
    n22101, n22102, n22103, n22104, n22105, n22106, n22107, n22108, n22109,
    n22110, n22111, n22112, n22113, n22114, n22115, n22116, n22117, n22118,
    n22119, n22120, n22121, n22122, n22123, n22124, n22125, n22126, n22127,
    n22128, n22129, n22130, n22131, n22132, n22133, n22134, n22135, n22136,
    n22137, n22138, n22139, n22140, n22141, n22142, n22143, n22144, n22145,
    n22146, n22147, n22148, n22149, n22150, n22151, n22152, n22153, n22154,
    n22155, n22156, n22157, n22158, n22159, n22160, n22161, n22162, n22163,
    n22164, n22165, n22166, n22167, n22168, n22169, n22170, n22171, n22172,
    n22173, n22174, n22175, n22176, n22177, n22178, n22179, n22180, n22181,
    n22182, n22183, n22184, n22185, n22186, n22187, n22188, n22189, n22190,
    n22191, n22192, n22193, n22194, n22195, n22196, n22197, n22198, n22199,
    n22200, n22201, n22202, n22203, n22204, n22205, n22206, n22207, n22208,
    n22209, n22210, n22211, n22212, n22213, n22214, n22215, n22216, n22217,
    n22218, n22219, n22220, n22221, n22222, n22223, n22224, n22225, n22226,
    n22227, n22228, n22229, n22230, n22231, n22232, n22233, n22234, n22235,
    n22236, n22237, n22238, n22239, n22240, n22241, n22242, n22243, n22244,
    n22245, n22246, n22247, n22248, n22249, n22250, n22251, n22252, n22253,
    n22254, n22255, n22256, n22257, n22258, n22259, n22260, n22261, n22262,
    n22263, n22264, n22265, n22266, n22267, n22268, n22269, n22270, n22271,
    n22272, n22273, n22274, n22275, n22276, n22277, n22278, n22279, n22280,
    n22281, n22282, n22283, n22284, n22285, n22286, n22287, n22288, n22289,
    n22290, n22291, n22292, n22293, n22294, n22295, n22296, n22297, n22298,
    n22299, n22300, n22301, n22302, n22303, n22304, n22305, n22306, n22307,
    n22308, n22309, n22310, n22311, n22312, n22313, n22314, n22315, n22316,
    n22317, n22318, n22319, n22320, n22321, n22322, n22323, n22324, n22325,
    n22326, n22327, n22328, n22329, n22330, n22331, n22332, n22333, n22334,
    n22335, n22336, n22337, n22338, n22339, n22340, n22341, n22342, n22343,
    n22344, n22345, n22346, n22347, n22348, n22349, n22350, n22351, n22352,
    n22353, n22354, n22355, n22356, n22357, n22358, n22359, n22360, n22361,
    n22362, n22363, n22364, n22365, n22366, n22367, n22368, n22369, n22370,
    n22371, n22372, n22373, n22374, n22375, n22376, n22377, n22378, n22379,
    n22380, n22381, n22382, n22383, n22384, n22385, n22386, n22387, n22388,
    n22389, n22390, n22391, n22392, n22393, n22394, n22395, n22396, n22397,
    n22398, n22399, n22400, n22401, n22402, n22403, n22404, n22405, n22406,
    n22407, n22408, n22409, n22410, n22411, n22412, n22413, n22414, n22415,
    n22416, n22417, n22418, n22419, n22420, n22421, n22422, n22423, n22424,
    n22425, n22426, n22427, n22428, n22429, n22430, n22431, n22432, n22433,
    n22434, n22435, n22436, n22437, n22438, n22439, n22440, n22441, n22442,
    n22443, n22444, n22445, n22446, n22447, n22448, n22449, n22450, n22451,
    n22452, n22453, n22454, n22455, n22456, n22457, n22458, n22459, n22460,
    n22461, n22462, n22463, n22464, n22465, n22466, n22467, n22468, n22469,
    n22470, n22471, n22472, n22473, n22474, n22475, n22476, n22477, n22478,
    n22479, n22480, n22481, n22482, n22483, n22484, n22485, n22486, n22487,
    n22488, n22489, n22490, n22491, n22492, n22493, n22494, n22495, n22496,
    n22497, n22498, n22499, n22500, n22501, n22502, n22503, n22504, n22505,
    n22506, n22507, n22508, n22509, n22510, n22511, n22512, n22513, n22514,
    n22515, n22516, n22517, n22518, n22519, n22520, n22521, n22522, n22523,
    n22524, n22525, n22526, n22527, n22528, n22529, n22530, n22531, n22532,
    n22533, n22534, n22535, n22536, n22537, n22538, n22539, n22540, n22541,
    n22542, n22543, n22544, n22545, n22546, n22547, n22548, n22549, n22550,
    n22551, n22552, n22553, n22554, n22555, n22556, n22557, n22558, n22559,
    n22560, n22561, n22562, n22563, n22564, n22565, n22566, n22567, n22568,
    n22569, n22570, n22571, n22572, n22573, n22574, n22575, n22576, n22577,
    n22578, n22579, n22580, n22581, n22582, n22583, n22584, n22585, n22586,
    n22587, n22588, n22589, n22590, n22591, n22592, n22593, n22594, n22595,
    n22596, n22597, n22598, n22599, n22600, n22601, n22602, n22603, n22604,
    n22605, n22606, n22607, n22608, n22609, n22610, n22611, n22612, n22613,
    n22614, n22615, n22616, n22617, n22618, n22619, n22620, n22621, n22622,
    n22623, n22624, n22625, n22626, n22627, n22628, n22629, n22630, n22631,
    n22632, n22633, n22634, n22635, n22636, n22637, n22638, n22639, n22640,
    n22641, n22642, n22643, n22644, n22645, n22646, n22647, n22648, n22649,
    n22650, n22651, n22652, n22653, n22654, n22655, n22656, n22657, n22658,
    n22659, n22660, n22661, n22662, n22663, n22664, n22665, n22666, n22667,
    n22668, n22669, n22670, n22671, n22672, n22673, n22674, n22675, n22676,
    n22677, n22678, n22679, n22680, n22681, n22682, n22683, n22684, n22685,
    n22686, n22687, n22688, n22689, n22690, n22691, n22692, n22693, n22694,
    n22695, n22696, n22697, n22698, n22699, n22700, n22701, n22702, n22703,
    n22704, n22705, n22706, n22707, n22708, n22709, n22710, n22711, n22712,
    n22713, n22714, n22715, n22716, n22717, n22718, n22719, n22720, n22721,
    n22722, n22723, n22724, n22725, n22726, n22727, n22728, n22729, n22730,
    n22731, n22732, n22733, n22734, n22735, n22736, n22737, n22738, n22739,
    n22740, n22741, n22742, n22743, n22744, n22745, n22746, n22747, n22748,
    n22749, n22750, n22751, n22752, n22753, n22754, n22755, n22756, n22757,
    n22758, n22759, n22760, n22761, n22762, n22763, n22764, n22765, n22766,
    n22767, n22768, n22769, n22770, n22771, n22772, n22773, n22774, n22775,
    n22776, n22777, n22778, n22779, n22780, n22781, n22782, n22783, n22784,
    n22785, n22786, n22787, n22788, n22789, n22790, n22791, n22792, n22793,
    n22794, n22795, n22796, n22797, n22798, n22799, n22800, n22801, n22802,
    n22803, n22804, n22805, n22806, n22807, n22808, n22809, n22810, n22811,
    n22812, n22813, n22814, n22815, n22816, n22817, n22818, n22819, n22820,
    n22821, n22822, n22823, n22824, n22825, n22826, n22827, n22828, n22829,
    n22830, n22831, n22832, n22833, n22834, n22835, n22836, n22837, n22838,
    n22839, n22840, n22841, n22842, n22843, n22844, n22845, n22846, n22847,
    n22848, n22849, n22850, n22851, n22852, n22853, n22854, n22855, n22856,
    n22857, n22858, n22859, n22860, n22861, n22862, n22863, n22864, n22865,
    n22866, n22867, n22868, n22869, n22870, n22871, n22872, n22873, n22874,
    n22875, n22876, n22877, n22878, n22879, n22880, n22881, n22882, n22883,
    n22884, n22885, n22886, n22887, n22888, n22889, n22890, n22891, n22892,
    n22893, n22894, n22895, n22896, n22897, n22898, n22899, n22900, n22901,
    n22902, n22903, n22904, n22905, n22906, n22907, n22908, n22909, n22910,
    n22911, n22912, n22913, n22914, n22915, n22916, n22917, n22918, n22919,
    n22920, n22921, n22922, n22923, n22924, n22925, n22926, n22927, n22928,
    n22929, n22930, n22931, n22932, n22933, n22934, n22935, n22936, n22937,
    n22938, n22939, n22940, n22941, n22942, n22943, n22944, n22945, n22946,
    n22947, n22948, n22949, n22950, n22951, n22952, n22953, n22954, n22955,
    n22956, n22957, n22958, n22959, n22960, n22961, n22962, n22963, n22964,
    n22965, n22966, n22967, n22968, n22969, n22970, n22971, n22972, n22973,
    n22974, n22975, n22976, n22977, n22978, n22979, n22980, n22981, n22982,
    n22983, n22984, n22985, n22986, n22987, n22988, n22989, n22990, n22991,
    n22992, n22993, n22994, n22995, n22996, n22997, n22998, n22999, n23000,
    n23001, n23002, n23003, n23004, n23005, n23006, n23007, n23008, n23009,
    n23010, n23011, n23012, n23013, n23014, n23015, n23016, n23017, n23018,
    n23019, n23020, n23021, n23022, n23023, n23024, n23025, n23026, n23027,
    n23028, n23029, n23030, n23031, n23032, n23033, n23034, n23035, n23036,
    n23037, n23038, n23039, n23040, n23041, n23042, n23043, n23044, n23045,
    n23046, n23047, n23048, n23049, n23050, n23051, n23052, n23053, n23054,
    n23055, n23056, n23057, n23058, n23059, n23060, n23061, n23062, n23063,
    n23064, n23065, n23066, n23067, n23068, n23069, n23070, n23071, n23072,
    n23073, n23074, n23075, n23076, n23077, n23078, n23079, n23080, n23081,
    n23082, n23083, n23084, n23085, n23086, n23087, n23088, n23089, n23090,
    n23091, n23092, n23093, n23094, n23095, n23096, n23097, n23098, n23099,
    n23100, n23101, n23102, n23103, n23104, n23105, n23106, n23107, n23108,
    n23109, n23110, n23111, n23112, n23113, n23114, n23115, n23116, n23117,
    n23118, n23119, n23120, n23121, n23122, n23123, n23124, n23125, n23126,
    n23127, n23128, n23129, n23130, n23131, n23132, n23133, n23134, n23135,
    n23136, n23137, n23138, n23139, n23140, n23141, n23142, n23143, n23144,
    n23145, n23146, n23147, n23148, n23149, n23150, n23151, n23152, n23153,
    n23154, n23155, n23156, n23157, n23158, n23159, n23160, n23161, n23162,
    n23163, n23164, n23165, n23166, n23167, n23168, n23169, n23170, n23171,
    n23172, n23173, n23174, n23175, n23176, n23177, n23178, n23179, n23180,
    n23181, n23182, n23183, n23184, n23185, n23186, n23187, n23188, n23189,
    n23190, n23191, n23192, n23193, n23194, n23195, n23196, n23197, n23198,
    n23199, n23200, n23201, n23202, n23203, n23204, n23205, n23206, n23207,
    n23208, n23209, n23210, n23211, n23212, n23213, n23214, n23215, n23216,
    n23217, n23218, n23219, n23220, n23221, n23222, n23223, n23224, n23225,
    n23226, n23227, n23228, n23229, n23230, n23231, n23232, n23233, n23234,
    n23235, n23236, n23237, n23238, n23239, n23240, n23241, n23242, n23243,
    n23244, n23245, n23246, n23247, n23248, n23249, n23250, n23251, n23252,
    n23253, n23254, n23255, n23256, n23257, n23258, n23259, n23260, n23261,
    n23262, n23263, n23264, n23265, n23266, n23267, n23268, n23269, n23270,
    n23271, n23272, n23273, n23274, n23275, n23276, n23277, n23278, n23279,
    n23280, n23281, n23282, n23283, n23284, n23285, n23286, n23287, n23288,
    n23289, n23290, n23291, n23292, n23293, n23294, n23295, n23296, n23297,
    n23298, n23299, n23300, n23301, n23302, n23303, n23304, n23305, n23306,
    n23307, n23308, n23309, n23310, n23311, n23312, n23313, n23314, n23315,
    n23316, n23317, n23318, n23319, n23320, n23321, n23322, n23323, n23324,
    n23325, n23326, n23327, n23328, n23329, n23330, n23331, n23332, n23333,
    n23334, n23335, n23336, n23337, n23338, n23339, n23340, n23341, n23342,
    n23343, n23344, n23345, n23346, n23347, n23348, n23349, n23350, n23351,
    n23352, n23353, n23354, n23355, n23356, n23357, n23358, n23359, n23360,
    n23361, n23362, n23363, n23364, n23365, n23366, n23367, n23368, n23369,
    n23370, n23371, n23372, n23373, n23374, n23375, n23376, n23377, n23378,
    n23379, n23380, n23381, n23382, n23383, n23384, n23385, n23386, n23387,
    n23388, n23389, n23390, n23391, n23392, n23393, n23394, n23395, n23396,
    n23397, n23398, n23399, n23400, n23401, n23402, n23403, n23404, n23405,
    n23406, n23407, n23408, n23409, n23410, n23411, n23412, n23413, n23414,
    n23415, n23416, n23417, n23418, n23419, n23420, n23421, n23422, n23423,
    n23424, n23425, n23426, n23427, n23428, n23429, n23430, n23431, n23432,
    n23433, n23434, n23435, n23436, n23437, n23438, n23439, n23440, n23441,
    n23442, n23443, n23444, n23445, n23446, n23447, n23448, n23449, n23450,
    n23451, n23452, n23453, n23454, n23455, n23456, n23457, n23458, n23459,
    n23460, n23461, n23462, n23463, n23464, n23465, n23466, n23467, n23468,
    n23469, n23470, n23471, n23472, n23473, n23474, n23475, n23476, n23477,
    n23478, n23479, n23480, n23481, n23482, n23483, n23484, n23485, n23486,
    n23487, n23488, n23489, n23490, n23491, n23492, n23493, n23494, n23495,
    n23496, n23497, n23498, n23499, n23500, n23501, n23502, n23503, n23504,
    n23505, n23506, n23507, n23508, n23509, n23510, n23511, n23512, n23513,
    n23514, n23515, n23516, n23517, n23518, n23519, n23520, n23521, n23522,
    n23523, n23524, n23525, n23526, n23527, n23528, n23529, n23530, n23531,
    n23532, n23533, n23534, n23535, n23536, n23537, n23538, n23539, n23540,
    n23541, n23542, n23543, n23544, n23545, n23546, n23547, n23548, n23549,
    n23550, n23551, n23552, n23553, n23554, n23555, n23556, n23557, n23558,
    n23559, n23560, n23561, n23562, n23563, n23564, n23565, n23566, n23567,
    n23568, n23569, n23570, n23571, n23572, n23573, n23574, n23575, n23576,
    n23577, n23578, n23579, n23580, n23581, n23582, n23583, n23584, n23585,
    n23586, n23587, n23588, n23589, n23590, n23591, n23592, n23593, n23594,
    n23595, n23596, n23597, n23598, n23599, n23600, n23601, n23602, n23603,
    n23604, n23605, n23606, n23607, n23608, n23609, n23610, n23611, n23612,
    n23613, n23614, n23615, n23616, n23617, n23618, n23619, n23620, n23621,
    n23622, n23623, n23624, n23625, n23626, n23627, n23628, n23629, n23630,
    n23631, n23632, n23633, n23634, n23635, n23636, n23637, n23638, n23639,
    n23640, n23641, n23642, n23643, n23644, n23645, n23646, n23647, n23648,
    n23649, n23650, n23651, n23652, n23653, n23654, n23655, n23656, n23657,
    n23658, n23659, n23660, n23661, n23662, n23663, n23664, n23665, n23666,
    n23667, n23668, n23669, n23670, n23671, n23672, n23673, n23674, n23675,
    n23676, n23677, n23678, n23679, n23680, n23681, n23682, n23683, n23684,
    n23685, n23686, n23687, n23688, n23689, n23690, n23691, n23692, n23693,
    n23694, n23695, n23696, n23697, n23698, n23699, n23700, n23701, n23702,
    n23703, n23704, n23705, n23706, n23707, n23708, n23709, n23710, n23711,
    n23712, n23713, n23714, n23715, n23716, n23717, n23718, n23719, n23720,
    n23721, n23722, n23723, n23724, n23725, n23726, n23727, n23728, n23729,
    n23730, n23731, n23732, n23733, n23734, n23735, n23736, n23737, n23738,
    n23739, n23740, n23741, n23742, n23743, n23744, n23745, n23746, n23747,
    n23748, n23749, n23750, n23751, n23752, n23753, n23754, n23755, n23756,
    n23757, n23758, n23759, n23760, n23761, n23762, n23763, n23764, n23765,
    n23766, n23767, n23768, n23769, n23770, n23771, n23772, n23773, n23774,
    n23775, n23776, n23777, n23778, n23779, n23780, n23781, n23782, n23783,
    n23784, n23785, n23786, n23787, n23788, n23789, n23790, n23791, n23792,
    n23793, n23794, n23795, n23796, n23797, n23798, n23799, n23800, n23801,
    n23802, n23803, n23804, n23805, n23806, n23807, n23808, n23809, n23810,
    n23811, n23812, n23813, n23814, n23815, n23816, n23817, n23818, n23819,
    n23820, n23821, n23822, n23823, n23824, n23825, n23826, n23827, n23828,
    n23829, n23830, n23831, n23832, n23833, n23834, n23835, n23836, n23837,
    n23838, n23839, n23840, n23841, n23842, n23843, n23844, n23845, n23846,
    n23847, n23848, n23849, n23850, n23851, n23852, n23853, n23854, n23855,
    n23856, n23857, n23858, n23859, n23860, n23861, n23862, n23863, n23864,
    n23865, n23866, n23867, n23868, n23869, n23870, n23871, n23872, n23873,
    n23874, n23875, n23876, n23877, n23878, n23879, n23880, n23881, n23882,
    n23883, n23884, n23885, n23886, n23887, n23888, n23889, n23890, n23891,
    n23892, n23893, n23894, n23895, n23896, n23897, n23898, n23899, n23900,
    n23901, n23902, n23903, n23904, n23905, n23906, n23907, n23908, n23909,
    n23910, n23911, n23912, n23913, n23914, n23915, n23916, n23917, n23918,
    n23919, n23920, n23921, n23922, n23923, n23924, n23925, n23926, n23927,
    n23928, n23929, n23930, n23931, n23932, n23933, n23934, n23935, n23936,
    n23937, n23938, n23939, n23940, n23941, n23942, n23943, n23944, n23945,
    n23946, n23947, n23948, n23949, n23950, n23951, n23952, n23953, n23954,
    n23955, n23956, n23957, n23958, n23959, n23960, n23961, n23962, n23963,
    n23964, n23965, n23966, n23967, n23968, n23969, n23970, n23971, n23972,
    n23973, n23974, n23975, n23976, n23977, n23978, n23979, n23980, n23981,
    n23982, n23983, n23984, n23985, n23986, n23987, n23988, n23989, n23990,
    n23991, n23992, n23993, n23994, n23995, n23996, n23997, n23998, n23999,
    n24000, n24001, n24002, n24003, n24004, n24005, n24006, n24007, n24008,
    n24009, n24010, n24011, n24012, n24013, n24014, n24015, n24016, n24017,
    n24018, n24019, n24020, n24021, n24022, n24023, n24024, n24025, n24026,
    n24027, n24028, n24029, n24030, n24031, n24032, n24033, n24034, n24035,
    n24036, n24037, n24038, n24039, n24040, n24041, n24042, n24043, n24044,
    n24045, n24046, n24047, n24048, n24049, n24050, n24051, n24052, n24053,
    n24054, n24055, n24056, n24057, n24058, n24059, n24060, n24061, n24062,
    n24063, n24064, n24065, n24066, n24067, n24068, n24069, n24070, n24071,
    n24072, n24073, n24074, n24075, n24076, n24077, n24078, n24079, n24080,
    n24081, n24082, n24083, n24084, n24085, n24086, n24087, n24088, n24089,
    n24090, n24091, n24092, n24093, n24094, n24095, n24096, n24097, n24098,
    n24099, n24100, n24101, n24102, n24103, n24104, n24105, n24106, n24107,
    n24108, n24109, n24110, n24111, n24112, n24113, n24114, n24115, n24116,
    n24117, n24118, n24119, n24120, n24121, n24122, n24123, n24124, n24125,
    n24126, n24127, n24128, n24129, n24130, n24131, n24132, n24133, n24134,
    n24135, n24136, n24137, n24138, n24139, n24140, n24141, n24142, n24143,
    n24144, n24145, n24146, n24147, n24148, n24149, n24150, n24151, n24152,
    n24153, n24154, n24155, n24156, n24157, n24158, n24159, n24160, n24161,
    n24162, n24163, n24164, n24165, n24166, n24167, n24168, n24169, n24170,
    n24171, n24172, n24173, n24174, n24175, n24176, n24177, n24178, n24179,
    n24180, n24181, n24182, n24183, n24184, n24185, n24186, n24187, n24188,
    n24189, n24190, n24191, n24192, n24193, n24194, n24195, n24196, n24197,
    n24198, n24199, n24200, n24201, n24202, n24203, n24204, n24205, n24206,
    n24207, n24208, n24209, n24210, n24211, n24212, n24213, n24214, n24215,
    n24216, n24217, n24218, n24219, n24220, n24221, n24222, n24223, n24224,
    n24225, n24226, n24227, n24228, n24229, n24230, n24231, n24232, n24233,
    n24234, n24235, n24236, n24237, n24238, n24239, n24240, n24241, n24242,
    n24243, n24244, n24245, n24246, n24247, n24248, n24249, n24250, n24251,
    n24252, n24253, n24254, n24255, n24256, n24257, n24258, n24259, n24260,
    n24261, n24262, n24263, n24264, n24265, n24266, n24267, n24268, n24269,
    n24270, n24271, n24272, n24273, n24274, n24275, n24276, n24277, n24278,
    n24279, n24280, n24281, n24282, n24283, n24284, n24285, n24286, n24287,
    n24288, n24289, n24290, n24291, n24292, n24293, n24294, n24295, n24296,
    n24297, n24298, n24299, n24300, n24301, n24302, n24303, n24304, n24305,
    n24306, n24307, n24308, n24309, n24310, n24311, n24312, n24313, n24314,
    n24315, n24316, n24317, n24318, n24319, n24320, n24321, n24322, n24323,
    n24324, n24325, n24326, n24327, n24328, n24329, n24330, n24331, n24332,
    n24333, n24334, n24335, n24336, n24337, n24338, n24339, n24340, n24341,
    n24342, n24343, n24344, n24345, n24346, n24347, n24348, n24349, n24350,
    n24351, n24352, n24353, n24354, n24355, n24356, n24357, n24358, n24359,
    n24360, n24361, n24362, n24363, n24364, n24365, n24366, n24367, n24368,
    n24369, n24370, n24371, n24372, n24373, n24374, n24375, n24376, n24377,
    n24378, n24379, n24380, n24381, n24382, n24383, n24384, n24385, n24386,
    n24387, n24388, n24389, n24390, n24391, n24392, n24393, n24394, n24395,
    n24396, n24397, n24398, n24399, n24400, n24401, n24402, n24403, n24404,
    n24405, n24406, n24407, n24408, n24409, n24410, n24411, n24412, n24413,
    n24414, n24415, n24416, n24417, n24418, n24419, n24420, n24421, n24422,
    n24423, n24424, n24425, n24426, n24427, n24428, n24429, n24430, n24431,
    n24432, n24433, n24434, n24435, n24436, n24437, n24438, n24439, n24440,
    n24441, n24442, n24443, n24444, n24445, n24446, n24447, n24448, n24449,
    n24450, n24451, n24452, n24453, n24454, n24455, n24456, n24457, n24458,
    n24459, n24460, n24461, n24462, n24463, n24464, n24465, n24466, n24467,
    n24468, n24469, n24470, n24471, n24472, n24473, n24474, n24475, n24476,
    n24477, n24478, n24479, n24480, n24481, n24482, n24483, n24484, n24485,
    n24486, n24487, n24488, n24489, n24490, n24491, n24492, n24493, n24494,
    n24495, n24496, n24497, n24498, n24499, n24500, n24501, n24502, n24503,
    n24504, n24505, n24506, n24507, n24508, n24509, n24510, n24511, n24512,
    n24513, n24514, n24515, n24516, n24517, n24518, n24519, n24520, n24521,
    n24522, n24523, n24524, n24525, n24526, n24527, n24528, n24529, n24530,
    n24531, n24532, n24533, n24534, n24535, n24536, n24537, n24538, n24539,
    n24540, n24541, n24542, n24543, n24544, n24545, n24546, n24547, n24548,
    n24549, n24550, n24551, n24552, n24553, n24554, n24555, n24556, n24557,
    n24558, n24559, n24560, n24561, n24562, n24563, n24564, n24565, n24566,
    n24567, n24568, n24569, n24570, n24571, n24572, n24573, n24574, n24575,
    n24576, n24577, n24578, n24579, n24580, n24581, n24582, n24583, n24584,
    n24585, n24586, n24587, n24588, n24589, n24590, n24591, n24592, n24593,
    n24594, n24595, n24596, n24597, n24598, n24599, n24600, n24601, n24602,
    n24603, n24604, n24605, n24606, n24607, n24608, n24609, n24610, n24611,
    n24612, n24613, n24614, n24615, n24616, n24617, n24618, n24619, n24620,
    n24621, n24622, n24623, n24624, n24625, n24626, n24627, n24628, n24629,
    n24630, n24631, n24632, n24633, n24634, n24635, n24636, n24637, n24638,
    n24639, n24640, n24641, n24642, n24643, n24644, n24645, n24646, n24647,
    n24648, n24649, n24650, n24651, n24652, n24653, n24654, n24655, n24656,
    n24657, n24658, n24659, n24660, n24661, n24662, n24663, n24664, n24665,
    n24666, n24667, n24668, n24669, n24670, n24671, n24672, n24673, n24674,
    n24675, n24676, n24677, n24678, n24679, n24680, n24681, n24682, n24683,
    n24684, n24685, n24686, n24687, n24688, n24689, n24690, n24691, n24692,
    n24693, n24694, n24695, n24696, n24697, n24698, n24699, n24700, n24701,
    n24702, n24703, n24704, n24705, n24706, n24707, n24708, n24709, n24710,
    n24711, n24712, n24713, n24714, n24715, n24716, n24717, n24718, n24719,
    n24720, n24721, n24722, n24723, n24724, n24725, n24726, n24727, n24728,
    n24729, n24730, n24731, n24732, n24733, n24734, n24735, n24736, n24737,
    n24738, n24739, n24740, n24741, n24742, n24743, n24744, n24745, n24746,
    n24747, n24748, n24749, n24750, n24751, n24752, n24753, n24754, n24755,
    n24756, n24757, n24758, n24759, n24760, n24761, n24762, n24763, n24764,
    n24765, n24766, n24767, n24768, n24769, n24770, n24771, n24772, n24773,
    n24774, n24775, n24776, n24777, n24778, n24779, n24780, n24781, n24782,
    n24783, n24784, n24785, n24786, n24787, n24788, n24789, n24790, n24791,
    n24792, n24793, n24794, n24795, n24796, n24797, n24798, n24799, n24800,
    n24801, n24802, n24803, n24804, n24805, n24806, n24807, n24808, n24809,
    n24810, n24811, n24812, n24813, n24814, n24815, n24816, n24817, n24818,
    n24819, n24820, n24821, n24822, n24823, n24824, n24825, n24826, n24827,
    n24828, n24829, n24830, n24831, n24832, n24833, n24834, n24835, n24836,
    n24837, n24838, n24839, n24840, n24841, n24842, n24843, n24844, n24845,
    n24846, n24847, n24848, n24849, n24850, n24851, n24852, n24853, n24854,
    n24855, n24856, n24857, n24858, n24859, n24860, n24861, n24862, n24863,
    n24864, n24865, n24866, n24867, n24868, n24869, n24870, n24871, n24872,
    n24873, n24874, n24875, n24876, n24877, n24878, n24879, n24880, n24881,
    n24882, n24883, n24884, n24885, n24886, n24887, n24888, n24889, n24890,
    n24891, n24892, n24893, n24894, n24895, n24896, n24897, n24898, n24899,
    n24900, n24901, n24902, n24903, n24904, n24905, n24906, n24907, n24908,
    n24909, n24910, n24911, n24912, n24913, n24914, n24915, n24916, n24917,
    n24918, n24919, n24920, n24921, n24922, n24923, n24924, n24925, n24926,
    n24927, n24928, n24929, n24930, n24931, n24932, n24933, n24934, n24935,
    n24936, n24937, n24938, n24939, n24940, n24941, n24942, n24943, n24944,
    n24945, n24946, n24947, n24948, n24949, n24950, n24951, n24952, n24953,
    n24954, n24955, n24956, n24957, n24958, n24959, n24960, n24961, n24962,
    n24963, n24964, n24965, n24966, n24967, n24968, n24969, n24970, n24971,
    n24972, n24973, n24974, n24975, n24976, n24977, n24978, n24979, n24980,
    n24981, n24982, n24983, n24984, n24985, n24986, n24987, n24988, n24989,
    n24990, n24991, n24992, n24993, n24994, n24995, n24996, n24997, n24998,
    n24999, n25000, n25001, n25002, n25003, n25004, n25005, n25006, n25007,
    n25008, n25009, n25010, n25011, n25012, n25013, n25014, n25015, n25016,
    n25017, n25018, n25019, n25020, n25021, n25022, n25023, n25024, n25025,
    n25026, n25027, n25028, n25029, n25030, n25031, n25032, n25033, n25034,
    n25035, n25036, n25037, n25038, n25039, n25040, n25041, n25042, n25043,
    n25044, n25045, n25046, n25047, n25048, n25049, n25050, n25051, n25052,
    n25053, n25054, n25055, n25056, n25057, n25058, n25059, n25060, n25061,
    n25062, n25063, n25064, n25065, n25066, n25067, n25068, n25069, n25070,
    n25071, n25072, n25073, n25074, n25075, n25076, n25077, n25078, n25079,
    n25080, n25081, n25082, n25083, n25084, n25085, n25086, n25087, n25088,
    n25089, n25090, n25091, n25092, n25093, n25094, n25095, n25096, n25097,
    n25098, n25099, n25100, n25101, n25102, n25103, n25104, n25105, n25106,
    n25107, n25108, n25109, n25110, n25111, n25112, n25113, n25114, n25115,
    n25116, n25117, n25118, n25119, n25120, n25121, n25122, n25123, n25124,
    n25125, n25126, n25127, n25128, n25129, n25130, n25131, n25132, n25133,
    n25134, n25135, n25136, n25137, n25138, n25139, n25140, n25141, n25142,
    n25143, n25144, n25145, n25146, n25147, n25148, n25149, n25150, n25151,
    n25152, n25153, n25154, n25155, n25156, n25157, n25158, n25159, n25160,
    n25161, n25162, n25163, n25164, n25165, n25166, n25167, n25168, n25169,
    n25170, n25171, n25172, n25173, n25174, n25175, n25176, n25177, n25178,
    n25179, n25180, n25181, n25182, n25183, n25184, n25185, n25186, n25187,
    n25188, n25189, n25190, n25191, n25192, n25193, n25194, n25195, n25196,
    n25197, n25198, n25199, n25200, n25201, n25202, n25203, n25204, n25205,
    n25206, n25207, n25208, n25209, n25210, n25211, n25212, n25213, n25214,
    n25215, n25216, n25217, n25218, n25219, n25220, n25221, n25222, n25223,
    n25224, n25225, n25226, n25227, n25228, n25229, n25230, n25231, n25232,
    n25233, n25234, n25235, n25236, n25237, n25238, n25239, n25240, n25241,
    n25242, n25243, n25244, n25245, n25246, n25247, n25248, n25249, n25250,
    n25251, n25252, n25253, n25254, n25255, n25256, n25257, n25258, n25259,
    n25260, n25261, n25262, n25263, n25264, n25265, n25266, n25267, n25268,
    n25269, n25270, n25271, n25272, n25273, n25274, n25275, n25276, n25277,
    n25278, n25279, n25280, n25281, n25282, n25283, n25284, n25285, n25286,
    n25287, n25288, n25289, n25290, n25291, n25292, n25293, n25294, n25295,
    n25296, n25297, n25298, n25299, n25300, n25301, n25302, n25303, n25304,
    n25305, n25306, n25307, n25308, n25309, n25310, n25311, n25312, n25313,
    n25314, n25315, n25316, n25317, n25318, n25319, n25320, n25321, n25322,
    n25323, n25324, n25325, n25326, n25327, n25328, n25329, n25330, n25331,
    n25332, n25333, n25334, n25335, n25336, n25337, n25338, n25339, n25340,
    n25341, n25342, n25343, n25344, n25345, n25346, n25347, n25348, n25349,
    n25350, n25351, n25352, n25353, n25354, n25355, n25356, n25357, n25358,
    n25359, n25360, n25361, n25362, n25363, n25364, n25365, n25366, n25367,
    n25368, n25369, n25370, n25371, n25372, n25373, n25374, n25375, n25376,
    n25377, n25378, n25379, n25380, n25381, n25382, n25383, n25384, n25385,
    n25386, n25387, n25388, n25389, n25390, n25391, n25392, n25393, n25394,
    n25395, n25396, n25397, n25398, n25399, n25400, n25401, n25402, n25403,
    n25404, n25405, n25406, n25407, n25408, n25409, n25410, n25411, n25412,
    n25413, n25414, n25415, n25416, n25417, n25418, n25419, n25420, n25421,
    n25422, n25423, n25424, n25425, n25426, n25427, n25428, n25429, n25430,
    n25431, n25432, n25433, n25434, n25435, n25436, n25437, n25438, n25439,
    n25440, n25441, n25442, n25443, n25444, n25445, n25446, n25447, n25448,
    n25449, n25450, n25451, n25452, n25453, n25454, n25455, n25456, n25457,
    n25458, n25459, n25460, n25461, n25462, n25463, n25464, n25465, n25466,
    n25467, n25468, n25469, n25470, n25471, n25472, n25473, n25474, n25475,
    n25476, n25477, n25478, n25479, n25480, n25481, n25482, n25483, n25484,
    n25485, n25486, n25487, n25488, n25489, n25490, n25491, n25492, n25493,
    n25494, n25495, n25496, n25497, n25498, n25499, n25500, n25501, n25502,
    n25503, n25504, n25505, n25506, n25507, n25508, n25509, n25510, n25511,
    n25512, n25513, n25514, n25515, n25516, n25517, n25518, n25519, n25520,
    n25521, n25522, n25523, n25524, n25525, n25526, n25527, n25528, n25529,
    n25530, n25531, n25532, n25533, n25534, n25535, n25536, n25537, n25538,
    n25539, n25540, n25541, n25542, n25543, n25544, n25545, n25546, n25547,
    n25548, n25549, n25550, n25551, n25552, n25553, n25554, n25555, n25556,
    n25557, n25558, n25559, n25560, n25561, n25562, n25563, n25564, n25565,
    n25566, n25567, n25568, n25569, n25570, n25571, n25572, n25573, n25574,
    n25575, n25576, n25577, n25578, n25579, n25580, n25581, n25582, n25583,
    n25584, n25585, n25586, n25587, n25588, n25589, n25590, n25591, n25592,
    n25593, n25594, n25595, n25596, n25597, n25598, n25599, n25600, n25601,
    n25602, n25603, n25604, n25605, n25606, n25607, n25608, n25609, n25610,
    n25611, n25612, n25613, n25614, n25615, n25616, n25617, n25618, n25619,
    n25620, n25621, n25622, n25623, n25624, n25625, n25626, n25627, n25628,
    n25629, n25630, n25631, n25632, n25633, n25634, n25635, n25636, n25637,
    n25638, n25639, n25640, n25641, n25642, n25643, n25644, n25645, n25646,
    n25647, n25648, n25649, n25650, n25651, n25652, n25653, n25654, n25655,
    n25656, n25657, n25658, n25659, n25660, n25661, n25662, n25663, n25664,
    n25665, n25666, n25667, n25668, n25669, n25670, n25671, n25672, n25673,
    n25674, n25675, n25676, n25677, n25678, n25679, n25680, n25681, n25682,
    n25683, n25684, n25685, n25686, n25687, n25688, n25689, n25690, n25691,
    n25692, n25693, n25694, n25695, n25696, n25697, n25698, n25699, n25700,
    n25701, n25702, n25703, n25704, n25705, n25706, n25707, n25708, n25709,
    n25710, n25711, n25712, n25713, n25714, n25715, n25716, n25717, n25718,
    n25719, n25720, n25721, n25722, n25723, n25724, n25725, n25726, n25727,
    n25728, n25729, n25730, n25731, n25732, n25733, n25734, n25735, n25736,
    n25737, n25738, n25739, n25740, n25741, n25742, n25743, n25744, n25745,
    n25746, n25747, n25748, n25749, n25750, n25751, n25752, n25753, n25754,
    n25755, n25756, n25757, n25758, n25759, n25760, n25761, n25762, n25763,
    n25764, n25765, n25766, n25767, n25768, n25769, n25770, n25771, n25772,
    n25773, n25774, n25775, n25776, n25777, n25778, n25779, n25780, n25781,
    n25782, n25783, n25784, n25785, n25786, n25787, n25788, n25789, n25790,
    n25791, n25792, n25793, n25794, n25795, n25796, n25797, n25798, n25799,
    n25800, n25801, n25802, n25803, n25804, n25805, n25806, n25807, n25808,
    n25809, n25810, n25811, n25812, n25813, n25814, n25815, n25816, n25817,
    n25818, n25819, n25820, n25821, n25822, n25823, n25824, n25825, n25826,
    n25827, n25828, n25829, n25830, n25831, n25832, n25833, n25834, n25835,
    n25836, n25837, n25838, n25839, n25840, n25841, n25842, n25843, n25844,
    n25845, n25846, n25847, n25848, n25849, n25850, n25851, n25852, n25853,
    n25854, n25855, n25856, n25857, n25858, n25859, n25860, n25861, n25862,
    n25863, n25864, n25865, n25866, n25867, n25868, n25869, n25870, n25871,
    n25872, n25873, n25874, n25875, n25876, n25877, n25878, n25879, n25880,
    n25881, n25882, n25883, n25884, n25885, n25886, n25887, n25888, n25889,
    n25890, n25891, n25892, n25893, n25894, n25895, n25896, n25897, n25898,
    n25899, n25900, n25901, n25902, n25903, n25904, n25905, n25906, n25907,
    n25908, n25909, n25910, n25911, n25912, n25913, n25914, n25915, n25916,
    n25917, n25918, n25919, n25920, n25921, n25922, n25923, n25924, n25925,
    n25926, n25927, n25928, n25929, n25930, n25931, n25932, n25933, n25934,
    n25935, n25936, n25937, n25938, n25939, n25940, n25941, n25942, n25943,
    n25944, n25945, n25946, n25947, n25948, n25949, n25950, n25951, n25952,
    n25953, n25954, n25955, n25956, n25957, n25958, n25959, n25960, n25961,
    n25962, n25963, n25964, n25965, n25966, n25967, n25968, n25969, n25970,
    n25971, n25972, n25973, n25974, n25975, n25976, n25977, n25978, n25979,
    n25980, n25981, n25982, n25983, n25984, n25985, n25986, n25987, n25988,
    n25989, n25990, n25991, n25992, n25993, n25994, n25995, n25996, n25997,
    n25998, n25999, n26000, n26001, n26002, n26003, n26004, n26005, n26006,
    n26007, n26008, n26009, n26010, n26011, n26012, n26013, n26014, n26015,
    n26016, n26017, n26018, n26019, n26020, n26021, n26022, n26023, n26024,
    n26025, n26026, n26027, n26028, n26029, n26030, n26031, n26032, n26033,
    n26034, n26035, n26036, n26037, n26038, n26039, n26040, n26041, n26042,
    n26043, n26044, n26045, n26046, n26047, n26048, n26049, n26050, n26051,
    n26052, n26053, n26054, n26055, n26056, n26057, n26058, n26059, n26060,
    n26061, n26062, n26063, n26064, n26065, n26066, n26067, n26068, n26069,
    n26070, n26071, n26072, n26073, n26074, n26075, n26076, n26077, n26078,
    n26079, n26080, n26081, n26082, n26083, n26084, n26085, n26086, n26087,
    n26088, n26089, n26090, n26091, n26092, n26093, n26094, n26095, n26096,
    n26097, n26098, n26099, n26100, n26101, n26102, n26103, n26104, n26105,
    n26106, n26107, n26108, n26109, n26110, n26111, n26112, n26113, n26114,
    n26115, n26116, n26117, n26118, n26119, n26120, n26121, n26122, n26123,
    n26124, n26125, n26126, n26127, n26128, n26129, n26130, n26131, n26132,
    n26133, n26134, n26135, n26136, n26137, n26138, n26139, n26140, n26141,
    n26142, n26143, n26144, n26145, n26146, n26147, n26148, n26149, n26150,
    n26151, n26152, n26153, n26154, n26155, n26156, n26157, n26158, n26159,
    n26160, n26161, n26162, n26163, n26164, n26165, n26166, n26167, n26168,
    n26169, n26170, n26171, n26172, n26173, n26174, n26175, n26176, n26177,
    n26178, n26179, n26180, n26181, n26182, n26183, n26184, n26185, n26186,
    n26187, n26188, n26189, n26190, n26191, n26192, n26193, n26194, n26195,
    n26196, n26197, n26198, n26199, n26200, n26201, n26202, n26203, n26204,
    n26205, n26206, n26207, n26208, n26209, n26210, n26211, n26212, n26213,
    n26214, n26215, n26216, n26217, n26218, n26219, n26220, n26221, n26222,
    n26223, n26224, n26225, n26226, n26227, n26228, n26229, n26230, n26231,
    n26232, n26233, n26234, n26235, n26236, n26237, n26238, n26239, n26240,
    n26241, n26242, n26243, n26244, n26245, n26246, n26247, n26248, n26249,
    n26250, n26251, n26252, n26253, n26254, n26255, n26256, n26257, n26258,
    n26259, n26260, n26261, n26262, n26263, n26264, n26265, n26266, n26267,
    n26268, n26269, n26270, n26271, n26272, n26273, n26274, n26275, n26276,
    n26277, n26278, n26279, n26280, n26281, n26282, n26283, n26284, n26285,
    n26286, n26287, n26288, n26289, n26290, n26291, n26292, n26293, n26294,
    n26295, n26296, n26297, n26298, n26299, n26300, n26301, n26302, n26303,
    n26304, n26305, n26306, n26307, n26308, n26309, n26310, n26311, n26312,
    n26313, n26314, n26315, n26316, n26317, n26318, n26319, n26320, n26321,
    n26322, n26323, n26324, n26325, n26326, n26327, n26328, n26329, n26330,
    n26331, n26332, n26333, n26334, n26335, n26336, n26337, n26338, n26339,
    n26340, n26341, n26342, n26343, n26344, n26345, n26346, n26347, n26348,
    n26349, n26350, n26351, n26352, n26353, n26354, n26355, n26356, n26357,
    n26358, n26359, n26360, n26361, n26362, n26363, n26364, n26365, n26366,
    n26367, n26368, n26369, n26370, n26371, n26372, n26373, n26374, n26375,
    n26376, n26377, n26378, n26379, n26380, n26381, n26382, n26383, n26384,
    n26385, n26386, n26387, n26388, n26389, n26390, n26391, n26392, n26393,
    n26394, n26395, n26396, n26397, n26398, n26399, n26400, n26401, n26402,
    n26403, n26404, n26405, n26406, n26407, n26408, n26409, n26410, n26411,
    n26412, n26413, n26414, n26415, n26416, n26417, n26418, n26419, n26420,
    n26421, n26422, n26423, n26424, n26425, n26426, n26427, n26428, n26429,
    n26430, n26431, n26432, n26433, n26434, n26435, n26436, n26437, n26438,
    n26439, n26440, n26441, n26442, n26443, n26444, n26445, n26446, n26447,
    n26448, n26449, n26450, n26451, n26452, n26453, n26454, n26455, n26456,
    n26457, n26458, n26459, n26460, n26461, n26462, n26463, n26464, n26465,
    n26466, n26467, n26468, n26469, n26470, n26471, n26472, n26473, n26474,
    n26475, n26476, n26477, n26478, n26479, n26480, n26481, n26482, n26483,
    n26484, n26485, n26486, n26487, n26488, n26489, n26490, n26491, n26492,
    n26493, n26494, n26495, n26496, n26497, n26498, n26499, n26500, n26501,
    n26502, n26503, n26504, n26505, n26506, n26507, n26508, n26509, n26510,
    n26511, n26512, n26513, n26514, n26515, n26516, n26517, n26518, n26519,
    n26520, n26521, n26522, n26523, n26524, n26525, n26526, n26527, n26528,
    n26529, n26530, n26531, n26532, n26533, n26534, n26535, n26536, n26537,
    n26538, n26539, n26540, n26541, n26542, n26543, n26544, n26545, n26546,
    n26547, n26548, n26549, n26550, n26551, n26552, n26553, n26554, n26555,
    n26556, n26557, n26558, n26559, n26560, n26561, n26562, n26563, n26564,
    n26565, n26566, n26567, n26568, n26569, n26570, n26571, n26572, n26573,
    n26574, n26575, n26576, n26577, n26578, n26579, n26580, n26581, n26582,
    n26583, n26584, n26585, n26586, n26587, n26588, n26589, n26590, n26591,
    n26592, n26593, n26594, n26595, n26596, n26597, n26598, n26599, n26600,
    n26601, n26602, n26603, n26604, n26605, n26606, n26607, n26608, n26609,
    n26610, n26611, n26612, n26613, n26614, n26615, n26616, n26617, n26618,
    n26619, n26620, n26621, n26622, n26623, n26624, n26625, n26626, n26627,
    n26628, n26629, n26630, n26631, n26632, n26633, n26634, n26635, n26636,
    n26637, n26638, n26639, n26640, n26641, n26642, n26643, n26644, n26645,
    n26646, n26647, n26648, n26649, n26650, n26651, n26652, n26653, n26654,
    n26655, n26656, n26657, n26658, n26659, n26660, n26661, n26662, n26663,
    n26664, n26665, n26666, n26667, n26668, n26669, n26670, n26671, n26672,
    n26673, n26674, n26675, n26676, n26677, n26678, n26679, n26680, n26681,
    n26682, n26683, n26684, n26685, n26686, n26687, n26688, n26689, n26690,
    n26691, n26692, n26693, n26694, n26695, n26696, n26697, n26698, n26699,
    n26700, n26701, n26702, n26703, n26704, n26705, n26706, n26707, n26708,
    n26709, n26710, n26711, n26712, n26713, n26714, n26715, n26716, n26717,
    n26718, n26719, n26720, n26721, n26722, n26723, n26724, n26725, n26726,
    n26727, n26728, n26729, n26730, n26731, n26732, n26733, n26734, n26735,
    n26736, n26737, n26738, n26739, n26740, n26741, n26742, n26743, n26744,
    n26745, n26746, n26747, n26748, n26749, n26750, n26751, n26752, n26753,
    n26754, n26755, n26756, n26757, n26758, n26759, n26760, n26761, n26762,
    n26763, n26764, n26765, n26766, n26767, n26768, n26769, n26770, n26771,
    n26772, n26773, n26774, n26775, n26776, n26777, n26778, n26779, n26780,
    n26781, n26782, n26783, n26784, n26785, n26786, n26787, n26788, n26789,
    n26790, n26791, n26792, n26793, n26794, n26795, n26796, n26797, n26798,
    n26799, n26800, n26801, n26802, n26803, n26804, n26805, n26806, n26807,
    n26808, n26809, n26810, n26811, n26812, n26813, n26814, n26815, n26816,
    n26817, n26818, n26819, n26820, n26821, n26822, n26823, n26824, n26825,
    n26826, n26827, n26828, n26829, n26830, n26831, n26832, n26833, n26834,
    n26835, n26836, n26837, n26838, n26839, n26840, n26841, n26842, n26843,
    n26844, n26845, n26846, n26847, n26848, n26849, n26850, n26851, n26852,
    n26853, n26854, n26855, n26856, n26857, n26858, n26859, n26860, n26861,
    n26862, n26863, n26864, n26865, n26866, n26867, n26868, n26869, n26870,
    n26871, n26872, n26873, n26874, n26875, n26876, n26877, n26878, n26879,
    n26880, n26881, n26882, n26883, n26884, n26885, n26886, n26887, n26888,
    n26889, n26890, n26891, n26892, n26893, n26894, n26895, n26896, n26897,
    n26898, n26899, n26900, n26901, n26902, n26903, n26904, n26905, n26906,
    n26907, n26908, n26909, n26910, n26911, n26912, n26913, n26914, n26915,
    n26916, n26917, n26918, n26919, n26920, n26921, n26922, n26923, n26924,
    n26925, n26926, n26927, n26928, n26929, n26930, n26931, n26932, n26933,
    n26934, n26935, n26936, n26937, n26938, n26939, n26940, n26941, n26942,
    n26943, n26944, n26945, n26946, n26947, n26948, n26949, n26950, n26951,
    n26952, n26953, n26954, n26955, n26956, n26957, n26958, n26959, n26960,
    n26961, n26962, n26963, n26964, n26965, n26966, n26967, n26968, n26969,
    n26970, n26971, n26972, n26973, n26974, n26975, n26976, n26977, n26978,
    n26979, n26980, n26981, n26982, n26983, n26984, n26985, n26986, n26987,
    n26988, n26989, n26990, n26991, n26992, n26993, n26994, n26995, n26996,
    n26997, n26998, n26999, n27000, n27001, n27002, n27003, n27004, n27005,
    n27006, n27007, n27008, n27009, n27010, n27011, n27012, n27013, n27014,
    n27015, n27016, n27017, n27018, n27019, n27020, n27021, n27022, n27023,
    n27024, n27025, n27026, n27027, n27028, n27029, n27030, n27031, n27032,
    n27033, n27034, n27035, n27036, n27037, n27038, n27039, n27040, n27041,
    n27042, n27043, n27044, n27045, n27046, n27047, n27048, n27049, n27050,
    n27051, n27052, n27053, n27054, n27055, n27056, n27057, n27058, n27059,
    n27060, n27061, n27062, n27063, n27064, n27065, n27066, n27067, n27068,
    n27069, n27070, n27071, n27072, n27073, n27074, n27075, n27076, n27077,
    n27078, n27079, n27080, n27081, n27082, n27083, n27084, n27085, n27086,
    n27087, n27088, n27089, n27090, n27091, n27092, n27093, n27094, n27095,
    n27096, n27097, n27098, n27099, n27100, n27101, n27102, n27103, n27104,
    n27105, n27106, n27107, n27108, n27109, n27110, n27111, n27112, n27113,
    n27114, n27115, n27116, n27117, n27118, n27119, n27120, n27121, n27122,
    n27123, n27124, n27125, n27126, n27127, n27128, n27129, n27130, n27131,
    n27132, n27133, n27134, n27135, n27136, n27137, n27138, n27139, n27140,
    n27141, n27142, n27143, n27144, n27145, n27146, n27147, n27148, n27149,
    n27150, n27151, n27152, n27153, n27154, n27155, n27156, n27157, n27158,
    n27159, n27160, n27161, n27162, n27163, n27164, n27165, n27166, n27167,
    n27168, n27169, n27170, n27171, n27172, n27173, n27174, n27175, n27176,
    n27177, n27178, n27179, n27180, n27181, n27182, n27183, n27184, n27185,
    n27186, n27187, n27188, n27189, n27190, n27191, n27192, n27193, n27194,
    n27195, n27196, n27197, n27198, n27199, n27200, n27201, n27202, n27203,
    n27204, n27205, n27206, n27207, n27208, n27209, n27210, n27211, n27212,
    n27213, n27214, n27215, n27216, n27217, n27218, n27219, n27220, n27221,
    n27222, n27223, n27224, n27225, n27226, n27227, n27228, n27229, n27230,
    n27231, n27232, n27233, n27234, n27235, n27236, n27237, n27238, n27239,
    n27240, n27241, n27242, n27243, n27244, n27245, n27246, n27247, n27248,
    n27249, n27250, n27251, n27252, n27253, n27254, n27255, n27256, n27257,
    n27258, n27259, n27260, n27261, n27262, n27263, n27264, n27265, n27266,
    n27267, n27268, n27269, n27270, n27271, n27272, n27273, n27274, n27275,
    n27276, n27277, n27278, n27279, n27280, n27281, n27282, n27283, n27284,
    n27285, n27286, n27287, n27288, n27289, n27290, n27291, n27292, n27293,
    n27294, n27295, n27296, n27297, n27298, n27299, n27300, n27301, n27302,
    n27303, n27304, n27305, n27306, n27307, n27308, n27309, n27310, n27311,
    n27312, n27313, n27314, n27315, n27316, n27317, n27318, n27319, n27320,
    n27321, n27322, n27323, n27324, n27325, n27326, n27327, n27328, n27329,
    n27330, n27331, n27332, n27333, n27334, n27335, n27336, n27337, n27338,
    n27339, n27340, n27341, n27342, n27343, n27344, n27345, n27346, n27347,
    n27348, n27349, n27350, n27351, n27352, n27353, n27354, n27355, n27356,
    n27357, n27358, n27359, n27360, n27361, n27362, n27363, n27364, n27365,
    n27366, n27367, n27368, n27369, n27370, n27371, n27372, n27373, n27374,
    n27375, n27376, n27377, n27378, n27379, n27380, n27381, n27382, n27383,
    n27384, n27385, n27386, n27387, n27388, n27389, n27390, n27391, n27392,
    n27393, n27394, n27395, n27396, n27397, n27398, n27399, n27400, n27401,
    n27402, n27403, n27404, n27405, n27406, n27407, n27408, n27409, n27410,
    n27411, n27412, n27413, n27414, n27415, n27416, n27417, n27418, n27419,
    n27420, n27421, n27422, n27423, n27424, n27425, n27426, n27427, n27428,
    n27429, n27430, n27431, n27432, n27433, n27434, n27435, n27436, n27437,
    n27438, n27439, n27440, n27441, n27442, n27443, n27444, n27445, n27446,
    n27447, n27448, n27449, n27450, n27451, n27452, n27453, n27454, n27455,
    n27456, n27457, n27458, n27459, n27460, n27461, n27462, n27463, n27464,
    n27465, n27466, n27467, n27468, n27469, n27470, n27471, n27472, n27473,
    n27474, n27475, n27476, n27477, n27478, n27479, n27480, n27481, n27482,
    n27483, n27484, n27485, n27486, n27487, n27488, n27489, n27490, n27491,
    n27492, n27493, n27494, n27495, n27496, n27497, n27498, n27499, n27500,
    n27501, n27502, n27503, n27504, n27505, n27506, n27507, n27508, n27509,
    n27510, n27511, n27512, n27513, n27514, n27515, n27516, n27517, n27518,
    n27519, n27520, n27521, n27522, n27523, n27524, n27525, n27526, n27527,
    n27528, n27529, n27530, n27531, n27532, n27533, n27534, n27535, n27536,
    n27537, n27538, n27539, n27540, n27541, n27542, n27543, n27544, n27545,
    n27546, n27547, n27548, n27549, n27550, n27551, n27552, n27553, n27554,
    n27555, n27556, n27557, n27558, n27559, n27560, n27561, n27562, n27563,
    n27564, n27565, n27566, n27567, n27568, n27569, n27570, n27571, n27572,
    n27573, n27574, n27575, n27576, n27577, n27578, n27579, n27580, n27581,
    n27582, n27583, n27584, n27585, n27586, n27587, n27588, n27589, n27590,
    n27591, n27592, n27593, n27594, n27595, n27596, n27597, n27598, n27599,
    n27600, n27601, n27602, n27603, n27604, n27605, n27606, n27607, n27608,
    n27609, n27610, n27611, n27612, n27613, n27614, n27615, n27616, n27617,
    n27618, n27619, n27620, n27621, n27622, n27623, n27624, n27625, n27626,
    n27627, n27628, n27629, n27630, n27631, n27632, n27633, n27634, n27635,
    n27636, n27637, n27638, n27639, n27640, n27641, n27642, n27643, n27644,
    n27645, n27646, n27647, n27648, n27649, n27650, n27651, n27652, n27653,
    n27654, n27655, n27656, n27657, n27658, n27659, n27660, n27661, n27662,
    n27663, n27664, n27665, n27666, n27667, n27668, n27669, n27670, n27671,
    n27672, n27673, n27674, n27675, n27676, n27677, n27678, n27679, n27680,
    n27681, n27682, n27683, n27684, n27685, n27686, n27687, n27688, n27689,
    n27690, n27691, n27692, n27693, n27694, n27695, n27696, n27697, n27698,
    n27699, n27700, n27701, n27702, n27703, n27704, n27705, n27706, n27707,
    n27708, n27709, n27710, n27711, n27712, n27713, n27714, n27715, n27716,
    n27717, n27718, n27719, n27720, n27721, n27722, n27723, n27724, n27725,
    n27726, n27727, n27728, n27729, n27730, n27731, n27732, n27733, n27734,
    n27735, n27736, n27737, n27738, n27739, n27740, n27741, n27742, n27743,
    n27744, n27745, n27746, n27747, n27748, n27749, n27750, n27751, n27752,
    n27753, n27754, n27755, n27756, n27757, n27758, n27759, n27760, n27761,
    n27762, n27763, n27764, n27765, n27766, n27767, n27768, n27769, n27770,
    n27771, n27772, n27773, n27774, n27775, n27776, n27777, n27778, n27779,
    n27780, n27781, n27782, n27783, n27784, n27785, n27786, n27787, n27788,
    n27789, n27790, n27791, n27792, n27793, n27794, n27795, n27796, n27797,
    n27798, n27799, n27800, n27801, n27802, n27803, n27804, n27805, n27806,
    n27807, n27808, n27809, n27810, n27811, n27812, n27813, n27814, n27815,
    n27816, n27817, n27818, n27819, n27820, n27821, n27822, n27823, n27824,
    n27825, n27826, n27827, n27828, n27829, n27830, n27831, n27832, n27833,
    n27834, n27835, n27836, n27837, n27838, n27839, n27840, n27841, n27842,
    n27843, n27844, n27845, n27846, n27847, n27848, n27849, n27850, n27851,
    n27852, n27853, n27854, n27855, n27856, n27857, n27858, n27859, n27860,
    n27861, n27862, n27863, n27864, n27865, n27866, n27867, n27868, n27869,
    n27870, n27871, n27872, n27873, n27874, n27875, n27876, n27877, n27878,
    n27879, n27880, n27881, n27882, n27883, n27884, n27885, n27886, n27887,
    n27888, n27889, n27890, n27891, n27892, n27893, n27894, n27895, n27896,
    n27897, n27898, n27899, n27900, n27901, n27902, n27903, n27904, n27905,
    n27906, n27907, n27908, n27909, n27910, n27911, n27912, n27913, n27914,
    n27915, n27916, n27917, n27918, n27919, n27920, n27921, n27922, n27923,
    n27924, n27925, n27926, n27927, n27928, n27929, n27930, n27931, n27932,
    n27933, n27934, n27935, n27936, n27937, n27938, n27939, n27940, n27941,
    n27942, n27943, n27944, n27945, n27946, n27947, n27948, n27949, n27950,
    n27951, n27952, n27953, n27954, n27955, n27956, n27957, n27958, n27959,
    n27960, n27961, n27962, n27963, n27964, n27965, n27966, n27967, n27968,
    n27969, n27970, n27971, n27972, n27973, n27974, n27975, n27976, n27977,
    n27978, n27979, n27980, n27981, n27982, n27983, n27984, n27985, n27986,
    n27987, n27988, n27989, n27990, n27991, n27992, n27993, n27994, n27995,
    n27996, n27997, n27998, n27999, n28000, n28001, n28002, n28003, n28004,
    n28005, n28006, n28007, n28008, n28009, n28010, n28011, n28012, n28013,
    n28014, n28015, n28016, n28017, n28018, n28019, n28020, n28021, n28022,
    n28023, n28024, n28025, n28026, n28027, n28028, n28029, n28030, n28031,
    n28032, n28033, n28034, n28035, n28036, n28037, n28038, n28039, n28040,
    n28041, n28042, n28043, n28044, n28045, n28046, n28047, n28048, n28049,
    n28050, n28051, n28052, n28053, n28054, n28055, n28056, n28057, n28058,
    n28059, n28060, n28061, n28062, n28063, n28064, n28065, n28066, n28067,
    n28068, n28069, n28070, n28071, n28072, n28073, n28074, n28075, n28076,
    n28077, n28078, n28079, n28080, n28081, n28082, n28083, n28084, n28085,
    n28086, n28087, n28088, n28089, n28090, n28091, n28092, n28093, n28094,
    n28095, n28096, n28097, n28098, n28099, n28100, n28101, n28102, n28103,
    n28104, n28105, n28106, n28107, n28108, n28109, n28110, n28111, n28112,
    n28113, n28114, n28115, n28116, n28117, n28118, n28119, n28120, n28121,
    n28122, n28123, n28124, n28125, n28126, n28127, n28128, n28129, n28130,
    n28131, n28132, n28133, n28134, n28135, n28136, n28137, n28138, n28139,
    n28140, n28141, n28142, n28143, n28144, n28145, n28146, n28147, n28148,
    n28149, n28150, n28151, n28152, n28153, n28154, n28155, n28156, n28157,
    n28158, n28159, n28160, n28161, n28162, n28163, n28164, n28165, n28166,
    n28167, n28168, n28169, n28170, n28171, n28172, n28173, n28174, n28175,
    n28176, n28177, n28178, n28179, n28180, n28181, n28182, n28183, n28184,
    n28185, n28186, n28187, n28188, n28189, n28190, n28191, n28192, n28193,
    n28194, n28195, n28196, n28197, n28198, n28199, n28200, n28201, n28202,
    n28203, n28204, n28205, n28206, n28207, n28208, n28209, n28210, n28211,
    n28212, n28213, n28214, n28215, n28216, n28217, n28218, n28219, n28220,
    n28221, n28222, n28223, n28224, n28225, n28226, n28227, n28228, n28229,
    n28230, n28231, n28232, n28233, n28234, n28235, n28236, n28237, n28238,
    n28239, n28240, n28241, n28242, n28243, n28244, n28245, n28246, n28247,
    n28248, n28249, n28250, n28251, n28252, n28253, n28254, n28255, n28256,
    n28257, n28258, n28259, n28260, n28261, n28262, n28263, n28264, n28265,
    n28266, n28267, n28268, n28269, n28270, n28271, n28272, n28273, n28274,
    n28275, n28276, n28277, n28278, n28279, n28280, n28281, n28282, n28283,
    n28284, n28285, n28286, n28287, n28288, n28289, n28290, n28291, n28292,
    n28293, n28294, n28295, n28296, n28297, n28298, n28299, n28300, n28301,
    n28302, n28303, n28304, n28305, n28306, n28307, n28308, n28309, n28310,
    n28311, n28312, n28313, n28314, n28315, n28316, n28317, n28318, n28319,
    n28320, n28321, n28322, n28323, n28324, n28325, n28326, n28327, n28328,
    n28329, n28330, n28331, n28332, n28333, n28334, n28335, n28336, n28337,
    n28338, n28339, n28340, n28341, n28342, n28343, n28344, n28345, n28346,
    n28347, n28348, n28349, n28350, n28351, n28352, n28353, n28354, n28355,
    n28356, n28357, n28358, n28359, n28360, n28361, n28362, n28363, n28364,
    n28365, n28366, n28367, n28368, n28369, n28370, n28371, n28372, n28373,
    n28374, n28375, n28376, n28377, n28378, n28379, n28380, n28381, n28382,
    n28383, n28384, n28385, n28386, n28387, n28388, n28389, n28390, n28391,
    n28392, n28393, n28394, n28395, n28396, n28397, n28398, n28399, n28400,
    n28401, n28402, n28403, n28404, n28405, n28406, n28407, n28408, n28409,
    n28410, n28411, n28412, n28413, n28414, n28415, n28416, n28417, n28418,
    n28419, n28420, n28421, n28422, n28423, n28424, n28425, n28426, n28427,
    n28428, n28429, n28430, n28431, n28432, n28433, n28434, n28435, n28436,
    n28437, n28438, n28439, n28440, n28441, n28442, n28443, n28444, n28445,
    n28446, n28447, n28448, n28449, n28450, n28451, n28452, n28453, n28454,
    n28455, n28456, n28457, n28458, n28459, n28460, n28461, n28462, n28463,
    n28464, n28465, n28466, n28467, n28468, n28469, n28470, n28471, n28472,
    n28473, n28474, n28475, n28476, n28477, n28478, n28479, n28480, n28481,
    n28482, n28483, n28484, n28485, n28486, n28487, n28488, n28489, n28490,
    n28491, n28492, n28493, n28494, n28495, n28496, n28497, n28498, n28499,
    n28500, n28501, n28502, n28503, n28504, n28505, n28506, n28507, n28508,
    n28509, n28510, n28511, n28512, n28513, n28514, n28515, n28516, n28517,
    n28518, n28519, n28520, n28521, n28522, n28523, n28524, n28525, n28526,
    n28527, n28528, n28529, n28530, n28531, n28532, n28533, n28534, n28535,
    n28536, n28537, n28538, n28539, n28540, n28541, n28542, n28543, n28544,
    n28545, n28546, n28547, n28548, n28549, n28550, n28551, n28552, n28553,
    n28554, n28555, n28556, n28557, n28558, n28559, n28560, n28561, n28562,
    n28563, n28564, n28565, n28566, n28567, n28568, n28569, n28570, n28571,
    n28572, n28573, n28574, n28575, n28576, n28577, n28578, n28579, n28580,
    n28581, n28582, n28583, n28584, n28585, n28586, n28587, n28588, n28589,
    n28590, n28591, n28592, n28593, n28594, n28595, n28596, n28597, n28598,
    n28599, n28600, n28601, n28602, n28603, n28604, n28605, n28606, n28607,
    n28608, n28609, n28610, n28611, n28612, n28613, n28614, n28615, n28616,
    n28617, n28618, n28619, n28620, n28621, n28622, n28623, n28624, n28625,
    n28626, n28627, n28628, n28629, n28630, n28631, n28632, n28633, n28634,
    n28635, n28636, n28637, n28638, n28639, n28640, n28641, n28642, n28643,
    n28644, n28645, n28646, n28647, n28648, n28649, n28650, n28651, n28652,
    n28653, n28654, n28655, n28656, n28657, n28658, n28659, n28660, n28661,
    n28662, n28663, n28664, n28665, n28666, n28667, n28668, n28669, n28670,
    n28671, n28672, n28673, n28674, n28675, n28676, n28677, n28678, n28679,
    n28680, n28681, n28682, n28683, n28684, n28685, n28686, n28687, n28688,
    n28689, n28690, n28691, n28692, n28693, n28694, n28695, n28696, n28697,
    n28698, n28699, n28700, n28701, n28702, n28703, n28704, n28705, n28706,
    n28707, n28708, n28709, n28710, n28711, n28712, n28713, n28714, n28715,
    n28716, n28717, n28718, n28719, n28720, n28721, n28722, n28723, n28724,
    n28725, n28726, n28727, n28728, n28729, n28730, n28731, n28732, n28733,
    n28734, n28735, n28736, n28737, n28738, n28739, n28740, n28741, n28742,
    n28743, n28744, n28745, n28746, n28747, n28748, n28749, n28750, n28751,
    n28752, n28753, n28754, n28755, n28756, n28757, n28758, n28759, n28760,
    n28761, n28762, n28763, n28764, n28765, n28766, n28767, n28768, n28769,
    n28770, n28771, n28772, n28773, n28774, n28775, n28776, n28777, n28778,
    n28779, n28780, n28781, n28782, n28783, n28784, n28785, n28786, n28787,
    n28788, n28789, n28790, n28791, n28792, n28793, n28794, n28795, n28796,
    n28797, n28798, n28799, n28800, n28801, n28802, n28803, n28804, n28805,
    n28806, n28807, n28808, n28809, n28810, n28811, n28812, n28813, n28814,
    n28815, n28816, n28817, n28818, n28819, n28820, n28821, n28822, n28823,
    n28824, n28825, n28826, n28827, n28828, n28829, n28830, n28831, n28832,
    n28833, n28834, n28835, n28836, n28837, n28838, n28839, n28840, n28841,
    n28842, n28843, n28844, n28845, n28846, n28847, n28848, n28849, n28850,
    n28851, n28852, n28853, n28854, n28855, n28856, n28857, n28858, n28859,
    n28860, n28861, n28862, n28863, n28864, n28865, n28866, n28867, n28868,
    n28869, n28870, n28871, n28872, n28873, n28874, n28875, n28876, n28877,
    n28878, n28879, n28880, n28881, n28882, n28883, n28884, n28885, n28886,
    n28887, n28888, n28889, n28890, n28891, n28892, n28893, n28894, n28895,
    n28896, n28897, n28898, n28899, n28900, n28901, n28902, n28903, n28904,
    n28905, n28906, n28907, n28908, n28909, n28910, n28911, n28912, n28913,
    n28914, n28915, n28916, n28917, n28918, n28919, n28920, n28921, n28922,
    n28923, n28924, n28925, n28926, n28927, n28928, n28929, n28930, n28931,
    n28932, n28933, n28934, n28935, n28936, n28937, n28938, n28939, n28940,
    n28941, n28942, n28943, n28944, n28945, n28946, n28947, n28948, n28949,
    n28950, n28951, n28952, n28953, n28954, n28955, n28956, n28957, n28958,
    n28959, n28960, n28961, n28962, n28963, n28964, n28965, n28966, n28967,
    n28968, n28969, n28970, n28971, n28972, n28973, n28974, n28975, n28976,
    n28977, n28978, n28979, n28980, n28981, n28982, n28983, n28984, n28985,
    n28986, n28987, n28988, n28989, n28990, n28991, n28992, n28993, n28994,
    n28995, n28996, n28997, n28998, n28999, n29000, n29001, n29002, n29003,
    n29004, n29005, n29006, n29007, n29008, n29009, n29010, n29011, n29012,
    n29013, n29014, n29015, n29016, n29017, n29018, n29019, n29020, n29021,
    n29022, n29023, n29024, n29025, n29026, n29027, n29028, n29029, n29030,
    n29031, n29032, n29033, n29034, n29035, n29036, n29037, n29038, n29039,
    n29040, n29041, n29042, n29043, n29044, n29045, n29046, n29047, n29048,
    n29049, n29050, n29051, n29052, n29053, n29054, n29055, n29056, n29057,
    n29058, n29059, n29060, n29061, n29062, n29063, n29064, n29065, n29066,
    n29067, n29068, n29069, n29070, n29071, n29072, n29073, n29074, n29075,
    n29076, n29077, n29078, n29079, n29080, n29081, n29082, n29083, n29084,
    n29085, n29086, n29087, n29088, n29089, n29090, n29091, n29092, n29093,
    n29094, n29095, n29096, n29097, n29098, n29099, n29100, n29101, n29102,
    n29103, n29104, n29105, n29106, n29107, n29108, n29109, n29110, n29111,
    n29112, n29113, n29114, n29115, n29116, n29117, n29118, n29119, n29120,
    n29121, n29122, n29123, n29124, n29125, n29126, n29127, n29128, n29129,
    n29130, n29131, n29132, n29133, n29134, n29135, n29136, n29137, n29138,
    n29139, n29140, n29141, n29142, n29143, n29144, n29145, n29146, n29147,
    n29148, n29149, n29150, n29151, n29152, n29153, n29154, n29155, n29156,
    n29157, n29158, n29159, n29160, n29161, n29162, n29163, n29164, n29165,
    n29166, n29167, n29168, n29169, n29170, n29171, n29172, n29173, n29174,
    n29175, n29176, n29177, n29178, n29179, n29180, n29181, n29182, n29183,
    n29184, n29185, n29186, n29187, n29188, n29189, n29190, n29191, n29192,
    n29193, n29194, n29195, n29196, n29197, n29198, n29199, n29200, n29201,
    n29202, n29203, n29204, n29205, n29206, n29207, n29208, n29209, n29210,
    n29211, n29212, n29213, n29214, n29215, n29216, n29217, n29218, n29219,
    n29220, n29221, n29222, n29223, n29224, n29225, n29226, n29227, n29228,
    n29229, n29230, n29231, n29232, n29233, n29234, n29235, n29236, n29237,
    n29238, n29239, n29240, n29241, n29242, n29243, n29244, n29245, n29246,
    n29247, n29248, n29249, n29250, n29251, n29252, n29253, n29254, n29255,
    n29256, n29257, n29258, n29259, n29260, n29261, n29262, n29263, n29264,
    n29265, n29266, n29267, n29268, n29269, n29270, n29271, n29272, n29273,
    n29274, n29275, n29276, n29277, n29278, n29279, n29280, n29281, n29282,
    n29283, n29284, n29285, n29286, n29287, n29288, n29289, n29290, n29291,
    n29292, n29293, n29294, n29295, n29296, n29297, n29298, n29299, n29300,
    n29301, n29302, n29303, n29304, n29305, n29306, n29307, n29308, n29309,
    n29310, n29311, n29312, n29313, n29314, n29315, n29316, n29317, n29318,
    n29319, n29320, n29321, n29322, n29323, n29324, n29325, n29326, n29327,
    n29328, n29329, n29330, n29331, n29332, n29333, n29334, n29335, n29336,
    n29337, n29338, n29339, n29340, n29341, n29342, n29343, n29344, n29345,
    n29346, n29347, n29348, n29349, n29350, n29351, n29352, n29353, n29354,
    n29355, n29356, n29357, n29358, n29359, n29360, n29361, n29362, n29363,
    n29364, n29365, n29366, n29367, n29368, n29369, n29370, n29371, n29372,
    n29373, n29374, n29375, n29376, n29377, n29378, n29379, n29380, n29381,
    n29382, n29383, n29384, n29385, n29386, n29387, n29388, n29389, n29390,
    n29391, n29392, n29393, n29394, n29395, n29396, n29397, n29398, n29399,
    n29400, n29401, n29402, n29403, n29404, n29405, n29406, n29407, n29408,
    n29409, n29410, n29411, n29412, n29413, n29414, n29415, n29416, n29417,
    n29418, n29419, n29420, n29421, n29422, n29423, n29424, n29425, n29426,
    n29427, n29428, n29429, n29430, n29431, n29432, n29433, n29434, n29435,
    n29436, n29437, n29438, n29439, n29440, n29441, n29442, n29443, n29444,
    n29445, n29446, n29447, n29448, n29449, n29450, n29451, n29452, n29453,
    n29454, n29455, n29456, n29457, n29458, n29459, n29460, n29461, n29462,
    n29463, n29464, n29465, n29466, n29467, n29468, n29469, n29470, n29471,
    n29472, n29473, n29474, n29475, n29476, n29477, n29478, n29479, n29480,
    n29481, n29482, n29483, n29484, n29485, n29486, n29487, n29488, n29489,
    n29490, n29491, n29492, n29493, n29494, n29495, n29496, n29497, n29498,
    n29499, n29500, n29501, n29502, n29503, n29504, n29505, n29506, n29507,
    n29508, n29509, n29510, n29511, n29512, n29513, n29514, n29515, n29516,
    n29517, n29518, n29519, n29520, n29521, n29522, n29523, n29524, n29525,
    n29526, n29527, n29528, n29529, n29530, n29531, n29532, n29533, n29534,
    n29535, n29536, n29537, n29538, n29539, n29540, n29541, n29542, n29543,
    n29544, n29545, n29546, n29547, n29548, n29549, n29550, n29551, n29552,
    n29553, n29554, n29555, n29556, n29557, n29558, n29559, n29560, n29561,
    n29562, n29563, n29564, n29565, n29566, n29567, n29568, n29569, n29570,
    n29571, n29572, n29573, n29574, n29575, n29576, n29577, n29578, n29579,
    n29580, n29581, n29582, n29583, n29584, n29585, n29586, n29587, n29588,
    n29589, n29590, n29591, n29592, n29593, n29594, n29595, n29596, n29597,
    n29598, n29599, n29600, n29601, n29602, n29603, n29604, n29605, n29606,
    n29607, n29608, n29609, n29610, n29611, n29612, n29613, n29614, n29615,
    n29616, n29617, n29618, n29619, n29620, n29621, n29622, n29623, n29624,
    n29625, n29626, n29627, n29628, n29629, n29630, n29631, n29632, n29633,
    n29634, n29635, n29636, n29637, n29638, n29639, n29640, n29641, n29642,
    n29643, n29644, n29645, n29646, n29647, n29648, n29649, n29650, n29651,
    n29652, n29653, n29654, n29655, n29656, n29657, n29658, n29659, n29660,
    n29661, n29662, n29663, n29664, n29665, n29666, n29667, n29668, n29669,
    n29670, n29671, n29672, n29673, n29674, n29675, n29676, n29677, n29678,
    n29679, n29680, n29681, n29682, n29683, n29684, n29685, n29686, n29687,
    n29688, n29689, n29690, n29691, n29692, n29693, n29694, n29695, n29696,
    n29697, n29698, n29699, n29700, n29701, n29702, n29703, n29704, n29705,
    n29706, n29707, n29708, n29709, n29710, n29711, n29712, n29713, n29714,
    n29715, n29716, n29717, n29718, n29719, n29720, n29721, n29722, n29723,
    n29724, n29725, n29726, n29727, n29728, n29729, n29730, n29731, n29732,
    n29733, n29734, n29735, n29736, n29737, n29738, n29739, n29740, n29741,
    n29742, n29743, n29744, n29745, n29746, n29747, n29748, n29749, n29750,
    n29751, n29752, n29753, n29754, n29755, n29756, n29757, n29758, n29759,
    n29760, n29761, n29762, n29763, n29764, n29765, n29766, n29767, n29768,
    n29769, n29770, n29771, n29772, n29773, n29774, n29775, n29776, n29777,
    n29778, n29779, n29780, n29781, n29782, n29783, n29784, n29785, n29786,
    n29787, n29788, n29789, n29790, n29791, n29792, n29793, n29794, n29795,
    n29796, n29797, n29798, n29799, n29800, n29801, n29802, n29803, n29804,
    n29805, n29806, n29807, n29808, n29809, n29810, n29811, n29812, n29813,
    n29814, n29815, n29816, n29817, n29818, n29819, n29820, n29821, n29822,
    n29823, n29824, n29825, n29826, n29827, n29828, n29829, n29830, n29831,
    n29832, n29833, n29834, n29835, n29836, n29837, n29838, n29839, n29840,
    n29841, n29842, n29843, n29844, n29845, n29846, n29847, n29848, n29849,
    n29850, n29851, n29852, n29853, n29854, n29855, n29856, n29857, n29858,
    n29859, n29860, n29861, n29862, n29863, n29864, n29865, n29866, n29867,
    n29868, n29869, n29870, n29871, n29872, n29873, n29874, n29875, n29876,
    n29877, n29878, n29879, n29880, n29881, n29882, n29883, n29884, n29885,
    n29886, n29887, n29888, n29889, n29890, n29891, n29892, n29893, n29894,
    n29895, n29896, n29897, n29898, n29899, n29900, n29901, n29902, n29903,
    n29904, n29905, n29906, n29907, n29908, n29909, n29910, n29911, n29912,
    n29913, n29914, n29915, n29916, n29917, n29918, n29919, n29920, n29921,
    n29922, n29923, n29924, n29925, n29926, n29927, n29928, n29929, n29930,
    n29931, n29932, n29933, n29934, n29935, n29936, n29937, n29938, n29939,
    n29940, n29941, n29942, n29943, n29944, n29945, n29946, n29947, n29948,
    n29949, n29950, n29951, n29952, n29953, n29954, n29955, n29956, n29957,
    n29958, n29959, n29960, n29961, n29962, n29963, n29964, n29965, n29966,
    n29967, n29968, n29969, n29970, n29971, n29972, n29973, n29974, n29975,
    n29976, n29977, n29978, n29979, n29980, n29981, n29982, n29983, n29984,
    n29985, n29986, n29987, n29988, n29989, n29990, n29991, n29992, n29993,
    n29994, n29995, n29996, n29997, n29998, n29999, n30000, n30001, n30002,
    n30003, n30004, n30005, n30006, n30007, n30008, n30009, n30010, n30011,
    n30012, n30013, n30014, n30015, n30016, n30017, n30018, n30019, n30020,
    n30021, n30022, n30023, n30024, n30025, n30026, n30027, n30028, n30029,
    n30030, n30031, n30032, n30033, n30034, n30035, n30036, n30037, n30038,
    n30039, n30040, n30041, n30042, n30043, n30044, n30045, n30046, n30047,
    n30048, n30049, n30050, n30051, n30052, n30053, n30054, n30055, n30056,
    n30057, n30058, n30059, n30060, n30061, n30062, n30063, n30064, n30065,
    n30066, n30067, n30068, n30069, n30070, n30071, n30072, n30073, n30074,
    n30075, n30076, n30077, n30078, n30079, n30080, n30081, n30082, n30083,
    n30084, n30085, n30086, n30087, n30088, n30089, n30090, n30091, n30092,
    n30093, n30094, n30095, n30096, n30097, n30098, n30099, n30100, n30101,
    n30102, n30103, n30104, n30105, n30106, n30107, n30108, n30109, n30110,
    n30111, n30112, n30113, n30114, n30115, n30116, n30117, n30118, n30119,
    n30120, n30121, n30122, n30123, n30124, n30125, n30126, n30127, n30128,
    n30129, n30130, n30131, n30132, n30133, n30134, n30135, n30136, n30137,
    n30138, n30139, n30140, n30141, n30142, n30143, n30144, n30145, n30146,
    n30147, n30148, n30149, n30150, n30151, n30152, n30153, n30154, n30155,
    n30156, n30157, n30158, n30159, n30160, n30161, n30162, n30163, n30164,
    n30165, n30166, n30167, n30168, n30169, n30170, n30171, n30172, n30173,
    n30174, n30175, n30176, n30177, n30178, n30179, n30180, n30181, n30182,
    n30183, n30184, n30185, n30186, n30187, n30188, n30189, n30190, n30191,
    n30192, n30193, n30194, n30195, n30196, n30197, n30198, n30199, n30200,
    n30201, n30202, n30203, n30204, n30205, n30206, n30207, n30208, n30209,
    n30210, n30211, n30212, n30213, n30214, n30215, n30216, n30217, n30218,
    n30219, n30220, n30221, n30222, n30223, n30224, n30225, n30226, n30227,
    n30228, n30229, n30230, n30231, n30232, n30233, n30234, n30235, n30236,
    n30237, n30238, n30239, n30240, n30241, n30242, n30243, n30244, n30245,
    n30246, n30247, n30248, n30249, n30250, n30251, n30252, n30253, n30254,
    n30255, n30256, n30257, n30258, n30259, n30260, n30261, n30262, n30263,
    n30264, n30265, n30266, n30267, n30268, n30269, n30270, n30271, n30272,
    n30273, n30274, n30275, n30276, n30277, n30278, n30279, n30280, n30281,
    n30282, n30283, n30284, n30285, n30286, n30287, n30288, n30289, n30290,
    n30291, n30292, n30293, n30294, n30295, n30296, n30297, n30298, n30299,
    n30300, n30301, n30302, n30303, n30304, n30305, n30306, n30307, n30308,
    n30309, n30310, n30311, n30312, n30313, n30314, n30315, n30316, n30317,
    n30318, n30319, n30320, n30321, n30322, n30323, n30324, n30325, n30326,
    n30327, n30328, n30329, n30330, n30331, n30332, n30333, n30334, n30335,
    n30336, n30337, n30338, n30339, n30340, n30341, n30342, n30343, n30344,
    n30345, n30346, n30347, n30348, n30349, n30350, n30351, n30352, n30353,
    n30354, n30355, n30356, n30357, n30358, n30359, n30360, n30361, n30362,
    n30363, n30364, n30365, n30366, n30367, n30368, n30369, n30370, n30371,
    n30372, n30373, n30374, n30375, n30376, n30377, n30378, n30379, n30380,
    n30381, n30382, n30383, n30384, n30385, n30386, n30387, n30388, n30389,
    n30390, n30391, n30392, n30393, n30394, n30395, n30396, n30397, n30398,
    n30399, n30400, n30401, n30402, n30403, n30404, n30405, n30406, n30407,
    n30408, n30409, n30410, n30411, n30412, n30413, n30414, n30415, n30416,
    n30417, n30418, n30419, n30420, n30421, n30422, n30423, n30424, n30425,
    n30426, n30427, n30428, n30429, n30430, n30431, n30432, n30433, n30434,
    n30435, n30436, n30437, n30438, n30439, n30440, n30441, n30442, n30443,
    n30444, n30445, n30446, n30447, n30448, n30449, n30450, n30451, n30452,
    n30453, n30454, n30455, n30456, n30457, n30458, n30459, n30460, n30461,
    n30462, n30463, n30464, n30465, n30466, n30467, n30468, n30469, n30470,
    n30471, n30472, n30473, n30474, n30475, n30476, n30477, n30478, n30479,
    n30480, n30481, n30482, n30483, n30484, n30485, n30486, n30487, n30488,
    n30489, n30490, n30491, n30492, n30493, n30494, n30495, n30496, n30497,
    n30498, n30499, n30500, n30501, n30502, n30503, n30504, n30505, n30506,
    n30507, n30508, n30509, n30510, n30511, n30512, n30513, n30514, n30515,
    n30516, n30517, n30518, n30519, n30520, n30521, n30522, n30523, n30524,
    n30525, n30526, n30527, n30528, n30529, n30530, n30531, n30532, n30533,
    n30534, n30535, n30536, n30537, n30538, n30539, n30540, n30541, n30542,
    n30543, n30544, n30545, n30546, n30547, n30548, n30549, n30550, n30551,
    n30552, n30553, n30554, n30555, n30556, n30557, n30558, n30559, n30560,
    n30561, n30562, n30563, n30564, n30565, n30566, n30567, n30568, n30569,
    n30570, n30571, n30572, n30573, n30574, n30575, n30576, n30577, n30578,
    n30579, n30580, n30581, n30582, n30583, n30584, n30585, n30586, n30587,
    n30588, n30589, n30590, n30591, n30592, n30593, n30594, n30595, n30596,
    n30597, n30598, n30599, n30600, n30601, n30602, n30603, n30604, n30605,
    n30606, n30607, n30608, n30609, n30610, n30611, n30612, n30613, n30614,
    n30615, n30616, n30617, n30618, n30619, n30620, n30621, n30622, n30623,
    n30624, n30625, n30626, n30627, n30628, n30629, n30630, n30631, n30632,
    n30633, n30634, n30635, n30636, n30637, n30638, n30639, n30640, n30641,
    n30642, n30643, n30644, n30645, n30646, n30647, n30648, n30649, n30650,
    n30651, n30652, n30653, n30654, n30655, n30656, n30657, n30658, n30659,
    n30660, n30661, n30662, n30663, n30664, n30665, n30666, n30667, n30668,
    n30669, n30670, n30671, n30672, n30673, n30674, n30675, n30676, n30677,
    n30678, n30679, n30680, n30681, n30682, n30683, n30684, n30685, n30686,
    n30687, n30688, n30689, n30690, n30691, n30692, n30693, n30694, n30695,
    n30696, n30697, n30698, n30699, n30700, n30701, n30702, n30703, n30704,
    n30705, n30706, n30707, n30708, n30709, n30710, n30711, n30712, n30713,
    n30714, n30715, n30716, n30717, n30718, n30719, n30720, n30721, n30722,
    n30723, n30724, n30725, n30726, n30727, n30728, n30729, n30730, n30731,
    n30732, n30733, n30734, n30735, n30736, n30737, n30738, n30739, n30740,
    n30741, n30742, n30743, n30744, n30745, n30746, n30747, n30748, n30749,
    n30750, n30751, n30752, n30753, n30754, n30755, n30756, n30757, n30758,
    n30759, n30760, n30761, n30762, n30763, n30764, n30765, n30766, n30767,
    n30768, n30769, n30770, n30771, n30772, n30773, n30774, n30775, n30776,
    n30777, n30778, n30779, n30780, n30781, n30782, n30783, n30784, n30785,
    n30786, n30787, n30788, n30789, n30790, n30791, n30792, n30793, n30794,
    n30795, n30796, n30797, n30798, n30799, n30800, n30801, n30802, n30803,
    n30804, n30805, n30806, n30807, n30808, n30809, n30810, n30811, n30812,
    n30813, n30814, n30815, n30816, n30817, n30818, n30819, n30820, n30821,
    n30822, n30823, n30824, n30825, n30826, n30827, n30828, n30829, n30830,
    n30831, n30832, n30833, n30834, n30835, n30836, n30837, n30838, n30839,
    n30840, n30841, n30842, n30843, n30844, n30845, n30846, n30847, n30848,
    n30849, n30850, n30851, n30852, n30853, n30854, n30855, n30856, n30857,
    n30858, n30859, n30860, n30861, n30862, n30863, n30864, n30865, n30866,
    n30867, n30868, n30869, n30870, n30871, n30872, n30873, n30874, n30875,
    n30876, n30877, n30878, n30879, n30880, n30881, n30882, n30883, n30884,
    n30885, n30886, n30887, n30888, n30889, n30890, n30891, n30892, n30893,
    n30894, n30895, n30896, n30897, n30898, n30899, n30900, n30901, n30902,
    n30903, n30904, n30905, n30906, n30907, n30908, n30909, n30910, n30911,
    n30912, n30913, n30914, n30915, n30916, n30917, n30918, n30919, n30920,
    n30921, n30922, n30923, n30924, n30925, n30926, n30927, n30928, n30929,
    n30930, n30931, n30932, n30933, n30934, n30935, n30936, n30937, n30938,
    n30939, n30940, n30941, n30942, n30943, n30944, n30945, n30946, n30947,
    n30948, n30949, n30950, n30951, n30952, n30953, n30954, n30955, n30956,
    n30957, n30958, n30959, n30960, n30961, n30962, n30963, n30964, n30965,
    n30966, n30967, n30968, n30969, n30970, n30971, n30972, n30973, n30974,
    n30975, n30976, n30977, n30978, n30979, n30980, n30981, n30982, n30983,
    n30984, n30985, n30986, n30987, n30988, n30989, n30990, n30991, n30992,
    n30993, n30994, n30995, n30996, n30997, n30998, n30999, n31000, n31001,
    n31002, n31003, n31004, n31005, n31006, n31007, n31008, n31009, n31010,
    n31011, n31012, n31013, n31014, n31015, n31016, n31017, n31018, n31019,
    n31020, n31021, n31022, n31023, n31024, n31025, n31026, n31027, n31028,
    n31029, n31030, n31031, n31032, n31033, n31034, n31035, n31036, n31037,
    n31038, n31039, n31040, n31041, n31042, n31043, n31044, n31045, n31046,
    n31047, n31048, n31049, n31050, n31051, n31052, n31053, n31054, n31055,
    n31056, n31057, n31058, n31059, n31060, n31061, n31062, n31063, n31064,
    n31065, n31066, n31067, n31068, n31069, n31070, n31071, n31072, n31073,
    n31074, n31075, n31076, n31077, n31078, n31079, n31080, n31081, n31082,
    n31083, n31084, n31085, n31086, n31087, n31088, n31089, n31090, n31091,
    n31092, n31093, n31094, n31095, n31096, n31097, n31098, n31099, n31100,
    n31101, n31102, n31103, n31104, n31105, n31106, n31107, n31108, n31109,
    n31110, n31111, n31112, n31113, n31114, n31115, n31116, n31117, n31118,
    n31119, n31120, n31121, n31122, n31123, n31124, n31125, n31126, n31127,
    n31128, n31129, n31130, n31131, n31132, n31133, n31134, n31135, n31136,
    n31137, n31138, n31139, n31140, n31141, n31142, n31143, n31144, n31145,
    n31146, n31147, n31148, n31149, n31150, n31151, n31152, n31153, n31154,
    n31155, n31156, n31157, n31158, n31159, n31160, n31161, n31162, n31163,
    n31164, n31165, n31166, n31167, n31168, n31169, n31170, n31171, n31172,
    n31173, n31174, n31175, n31176, n31177, n31178, n31179, n31180, n31181,
    n31182, n31183, n31184, n31185, n31186, n31187, n31188, n31189, n31190,
    n31191, n31192, n31193, n31194, n31195, n31196, n31197, n31198, n31199,
    n31200, n31201, n31202, n31203, n31204, n31205, n31206, n31207, n31208,
    n31209, n31210, n31211, n31212, n31213, n31214, n31215, n31216, n31217,
    n31218, n31219, n31220, n31221, n31222, n31223, n31224, n31225, n31226,
    n31227, n31228, n31229, n31230, n31231, n31232, n31233, n31234, n31235,
    n31236, n31237, n31238, n31239, n31240, n31241, n31242, n31243, n31244,
    n31245, n31246, n31247, n31248, n31249, n31250, n31251, n31252, n31253,
    n31254, n31255, n31256, n31257, n31258, n31259, n31260, n31261, n31262,
    n31263, n31264, n31265, n31266, n31267, n31268, n31269, n31270, n31271,
    n31272, n31273, n31274, n31275, n31276, n31277, n31278, n31279, n31280,
    n31281, n31282, n31283, n31284, n31285, n31286, n31287, n31288, n31289,
    n31290, n31291, n31292, n31293, n31294, n31295, n31296, n31297, n31298,
    n31299, n31300, n31301, n31302, n31303, n31304, n31305, n31306, n31307,
    n31308, n31309, n31310, n31311, n31312, n31313, n31314, n31315, n31316,
    n31317, n31318, n31319, n31320, n31321, n31322, n31323, n31324, n31325,
    n31326, n31327, n31328, n31329, n31330, n31331, n31332, n31333, n31334,
    n31335, n31336, n31337, n31338, n31339, n31340, n31341, n31342, n31343,
    n31344, n31345, n31346, n31347, n31348, n31349, n31350, n31351, n31352,
    n31353, n31354, n31355, n31356, n31357, n31358, n31359, n31360, n31361,
    n31362, n31363, n31364, n31365, n31366, n31367, n31368, n31369, n31370,
    n31371, n31372, n31373, n31374, n31375, n31376, n31377, n31378, n31379,
    n31380, n31381, n31382, n31383, n31384, n31385, n31386, n31387, n31388,
    n31389, n31390, n31391, n31392, n31393, n31394, n31395, n31396, n31397,
    n31398, n31399, n31400, n31401, n31402, n31403, n31404, n31405, n31406,
    n31407, n31408, n31409, n31410, n31411, n31412, n31413, n31414, n31415,
    n31416, n31417, n31418, n31419, n31420, n31421, n31422, n31423, n31424,
    n31425, n31426, n31427, n31428, n31429, n31430, n31431, n31432, n31433,
    n31434, n31435, n31436, n31437, n31438, n31439, n31440, n31441, n31442,
    n31443, n31444, n31445, n31446, n31447, n31448, n31449, n31450, n31451,
    n31452, n31453, n31454, n31455, n31456, n31457, n31458, n31459, n31460,
    n31461, n31462, n31463, n31464, n31465, n31466, n31467, n31468, n31469,
    n31470, n31471, n31472, n31473, n31474, n31475, n31476, n31477, n31478,
    n31479, n31480, n31481, n31482, n31483, n31484, n31485, n31486, n31487,
    n31488, n31489, n31490, n31491, n31492, n31493, n31494, n31495, n31496,
    n31497, n31498, n31499, n31500, n31501, n31502, n31503, n31504, n31505,
    n31506, n31507, n31508, n31509, n31510, n31511, n31512, n31513, n31514,
    n31515, n31516, n31517, n31518, n31519, n31520, n31521, n31522, n31523,
    n31524, n31525, n31526, n31527, n31528, n31529, n31530, n31531, n31532,
    n31533, n31534, n31535, n31536, n31537, n31538, n31539, n31540, n31541,
    n31542, n31543, n31544, n31545, n31546, n31547, n31548, n31549, n31550,
    n31551, n31552, n31553, n31554, n31555, n31556, n31557, n31558, n31559,
    n31560, n31561, n31562, n31563, n31564, n31565, n31566, n31567, n31568,
    n31569, n31570, n31571, n31572, n31573, n31574, n31575, n31576, n31577,
    n31578, n31579, n31580, n31581, n31582, n31583, n31584, n31585, n31586,
    n31587, n31588, n31589, n31590, n31591, n31592, n31593, n31594, n31595,
    n31596, n31597, n31598, n31599, n31600, n31601, n31602, n31603, n31604,
    n31605, n31606, n31607, n31608, n31609, n31610, n31611, n31612, n31613,
    n31614, n31615, n31616, n31617, n31618, n31619, n31620, n31621, n31622,
    n31623, n31624, n31625, n31626, n31627, n31628, n31629, n31630, n31631,
    n31632, n31633, n31634, n31635, n31636, n31637, n31638, n31639, n31640,
    n31641, n31642, n31643, n31644, n31645, n31646, n31647, n31648, n31649,
    n31650, n31651, n31652, n31653, n31654, n31655, n31656, n31657, n31658,
    n31659, n31660, n31661, n31662, n31663, n31664, n31665, n31666, n31667,
    n31668, n31669, n31670, n31671, n31672, n31673, n31674, n31675, n31676,
    n31677, n31678, n31679, n31680, n31681, n31682, n31683, n31684, n31685,
    n31686, n31687, n31688, n31689, n31690, n31691, n31692, n31693, n31694,
    n31695, n31696, n31697, n31698, n31699, n31700, n31701, n31702, n31703,
    n31704, n31705, n31706, n31707, n31708, n31709, n31710, n31711, n31712,
    n31713, n31714, n31715, n31716, n31717, n31718, n31719, n31720, n31721,
    n31722, n31723, n31724, n31725, n31726, n31727, n31728, n31729, n31730,
    n31731, n31732, n31733, n31734, n31735, n31736, n31737, n31738, n31739,
    n31740, n31741, n31742, n31743, n31744, n31745, n31746, n31747, n31748,
    n31749, n31750, n31751, n31752, n31753, n31754, n31755, n31756, n31757,
    n31758, n31759, n31760, n31761, n31762, n31763, n31764, n31765, n31766,
    n31767, n31768, n31769, n31770, n31771, n31772, n31773, n31774, n31775,
    n31776, n31777, n31778, n31779, n31780, n31781, n31782, n31783, n31784,
    n31785, n31786, n31787, n31788, n31789, n31790, n31791, n31792, n31793,
    n31794, n31795, n31796, n31797, n31798, n31799, n31800, n31801, n31802,
    n31803, n31804, n31805, n31806, n31807, n31808, n31809, n31810, n31811,
    n31812, n31813, n31814, n31815, n31816, n31817, n31818, n31819, n31820,
    n31821, n31822, n31823, n31824, n31825, n31826, n31827, n31828, n31829,
    n31830, n31831, n31832, n31833, n31834, n31835, n31836, n31837, n31838,
    n31839, n31840, n31841, n31842, n31843, n31844, n31845, n31846, n31847,
    n31848, n31849, n31850, n31851, n31852, n31853, n31854, n31855, n31856,
    n31857, n31858, n31859, n31860, n31861, n31862, n31863, n31864, n31865,
    n31866, n31867, n31868, n31869, n31870, n31871, n31872, n31873, n31874,
    n31875, n31876, n31877, n31878, n31879, n31880, n31881, n31882, n31883,
    n31884, n31885, n31886, n31887, n31888, n31889, n31890, n31891, n31892,
    n31893, n31894, n31895, n31896, n31897, n31898, n31899, n31900, n31901,
    n31902, n31903, n31904, n31905, n31906, n31907, n31908, n31909, n31910,
    n31911, n31912, n31913, n31914, n31915, n31916, n31917, n31918, n31919,
    n31920, n31921, n31922, n31923, n31924, n31925, n31926, n31927, n31928,
    n31929, n31930, n31931, n31932, n31933, n31934, n31935, n31936, n31937,
    n31938, n31939, n31940, n31941, n31942, n31943, n31944, n31945, n31946,
    n31947, n31948, n31949, n31950, n31951, n31952, n31953, n31954, n31955,
    n31956, n31957, n31958, n31959, n31960, n31961, n31962, n31963, n31964,
    n31965, n31966, n31967, n31968, n31969, n31970, n31971, n31972, n31973,
    n31974, n31975, n31976, n31977, n31978, n31979, n31980, n31981, n31982,
    n31983, n31984, n31985, n31986, n31987, n31988, n31989, n31990, n31991,
    n31992, n31993, n31994, n31995, n31996, n31997, n31998, n31999, n32000,
    n32001, n32002, n32003, n32004, n32005, n32006, n32007, n32008, n32009,
    n32010, n32011, n32012, n32013, n32014, n32015, n32016, n32017, n32018,
    n32019, n32020, n32021, n32022, n32023, n32024, n32025, n32026, n32027,
    n32028, n32029, n32030, n32031, n32032, n32033, n32034, n32035, n32036,
    n32037, n32038, n32039, n32040, n32041, n32042, n32043, n32044, n32045,
    n32046, n32047, n32048, n32049, n32050, n32051, n32052, n32053, n32054,
    n32055, n32056, n32057, n32058, n32059, n32060, n32061, n32062, n32063,
    n32064, n32065, n32066, n32067, n32068, n32069, n32070, n32071, n32072,
    n32073, n32074, n32075, n32076, n32077, n32078, n32079, n32080, n32081,
    n32082, n32083, n32084, n32085, n32086, n32087, n32088, n32089, n32090,
    n32091, n32092, n32093, n32094, n32095, n32096, n32097, n32098, n32099,
    n32100, n32101, n32102, n32103, n32104, n32105, n32106, n32107, n32108,
    n32109, n32110, n32111, n32112, n32113, n32114, n32115, n32116, n32117,
    n32118, n32119, n32120, n32121, n32122, n32123, n32124, n32125, n32126,
    n32127, n32128, n32129, n32130, n32131, n32132, n32133, n32134, n32135,
    n32136, n32137, n32138, n32139, n32140, n32141, n32142, n32143, n32144,
    n32145, n32146, n32147, n32148, n32149, n32150, n32151, n32152, n32153,
    n32154, n32155, n32156, n32157, n32158, n32159, n32160, n32161, n32162,
    n32163, n32164, n32165, n32166, n32167, n32168, n32169, n32170, n32171,
    n32172, n32173, n32174, n32175, n32176, n32177, n32178, n32179, n32180,
    n32181, n32182, n32183, n32184, n32185, n32186, n32187, n32188, n32189,
    n32190, n32191, n32192, n32193, n32194, n32195, n32196, n32197, n32198,
    n32199, n32200, n32201, n32202, n32203, n32204, n32205, n32206, n32207,
    n32208, n32209, n32210, n32211, n32212, n32213, n32214, n32215, n32216,
    n32217, n32218, n32219, n32220, n32221, n32222, n32223, n32224, n32225,
    n32226, n32227, n32228, n32229, n32230, n32231, n32232, n32233, n32234,
    n32235, n32236, n32237, n32238, n32239, n32240, n32241, n32242, n32243,
    n32244, n32245, n32246, n32247, n32248, n32249, n32250, n32251, n32252,
    n32253, n32254, n32255, n32256, n32257, n32258, n32259, n32260, n32261,
    n32262, n32263, n32264, n32265, n32266, n32267, n32268, n32269, n32270,
    n32271, n32272, n32273, n32274, n32275, n32276, n32277, n32278, n32279,
    n32280, n32281, n32282, n32283, n32284, n32285, n32286, n32287, n32288,
    n32289, n32290, n32291, n32292, n32293, n32294, n32295, n32296, n32297,
    n32298, n32299, n32300, n32301, n32302, n32303, n32304, n32305, n32306,
    n32307, n32308, n32309, n32310, n32311, n32312, n32313, n32314, n32315,
    n32316, n32317, n32318, n32319, n32320, n32321, n32322, n32323, n32324,
    n32325, n32326, n32327, n32328, n32329, n32330, n32331, n32332, n32333,
    n32334, n32335, n32336, n32337, n32338, n32339, n32340, n32341, n32342,
    n32343, n32344, n32345, n32346, n32347, n32348, n32349, n32350, n32351,
    n32352, n32353, n32354, n32355, n32356, n32357, n32358, n32359, n32360,
    n32361, n32362, n32363, n32364, n32365, n32366, n32367, n32368, n32369,
    n32370, n32371, n32372, n32373, n32374, n32375, n32376, n32377, n32378,
    n32379, n32380, n32381, n32382, n32383, n32384, n32385, n32386, n32387,
    n32388, n32389, n32390, n32391, n32392, n32393, n32394, n32395, n32396,
    n32397, n32398, n32399, n32400, n32401, n32402, n32403, n32404, n32405,
    n32406, n32407, n32408, n32409, n32410, n32411, n32412, n32413, n32414,
    n32415, n32416, n32417, n32418, n32419, n32420, n32421, n32422, n32423,
    n32424, n32425, n32426, n32427, n32428, n32429, n32430, n32431, n32432,
    n32433, n32434, n32435, n32436, n32437, n32438, n32439, n32440, n32441,
    n32442, n32443, n32444, n32445, n32446, n32447, n32448, n32449, n32450,
    n32451, n32452, n32453, n32454, n32455, n32456, n32457, n32458, n32459,
    n32460, n32461, n32462, n32463, n32464, n32465, n32466, n32467, n32468,
    n32469, n32470, n32471, n32472, n32473, n32474, n32475, n32476, n32477,
    n32478, n32479, n32480, n32481, n32482, n32483, n32484, n32485, n32486,
    n32487, n32488, n32489, n32490, n32491, n32492, n32493, n32494, n32495,
    n32496, n32497, n32498, n32499, n32500, n32501, n32502, n32503, n32504,
    n32505, n32506, n32507, n32508, n32509, n32510, n32511, n32512, n32513,
    n32514, n32515, n32516, n32517, n32518, n32519, n32520, n32521, n32522,
    n32523, n32524, n32525, n32526, n32527, n32528, n32529, n32530, n32531,
    n32532, n32533, n32534, n32535, n32536, n32537, n32538, n32539, n32540,
    n32541, n32542, n32543, n32544, n32545, n32546, n32547, n32548, n32549,
    n32550, n32551, n32552, n32553, n32554, n32555, n32556, n32557, n32558,
    n32559, n32560, n32561, n32562, n32563, n32564, n32565, n32566, n32567,
    n32568, n32569, n32570, n32571, n32572, n32573, n32574, n32575, n32576,
    n32577, n32578, n32579, n32580, n32581, n32582, n32583, n32584, n32585,
    n32586, n32587, n32588, n32589, n32590, n32591, n32592, n32593, n32594,
    n32595, n32596, n32597, n32598, n32599, n32600, n32601, n32602, n32603,
    n32604, n32605, n32606, n32607, n32608, n32609, n32610, n32611, n32612,
    n32613, n32614, n32615, n32616, n32617, n32618, n32619, n32620, n32621,
    n32622, n32623, n32624, n32625, n32626, n32627, n32628, n32629, n32630,
    n32631, n32632, n32633, n32634, n32635, n32636, n32637, n32638, n32639,
    n32640, n32641, n32642, n32643, n32644, n32645, n32646, n32647, n32648,
    n32649, n32650, n32651, n32652, n32653, n32654, n32655, n32656, n32657,
    n32658, n32659, n32660, n32661, n32662, n32663, n32664, n32665, n32666,
    n32667, n32668, n32669, n32670, n32671, n32672, n32673, n32674, n32675,
    n32676, n32677, n32678, n32679, n32680, n32681, n32682, n32683, n32684,
    n32685, n32686, n32687, n32688, n32689, n32690, n32691, n32692, n32693,
    n32694, n32695, n32696, n32697, n32698, n32699, n32700, n32701, n32702,
    n32703, n32704, n32705, n32706, n32707, n32708, n32709, n32710, n32711,
    n32712, n32713, n32714, n32715, n32716, n32717, n32718, n32719, n32720,
    n32721, n32722, n32723, n32724, n32725, n32726, n32727, n32728, n32729,
    n32730, n32731, n32732, n32733, n32734, n32735, n32736, n32737, n32738,
    n32739, n32740, n32741, n32742, n32743, n32744, n32745, n32746, n32747,
    n32748, n32749, n32750, n32751, n32752, n32753, n32754, n32755, n32756,
    n32757, n32758, n32759, n32760, n32761, n32762, n32763, n32764, n32765,
    n32766, n32767, n32768, n32769, n32770, n32771, n32772, n32773, n32774,
    n32775, n32776, n32777, n32778, n32779, n32780, n32781, n32782, n32783,
    n32784, n32785, n32786, n32787, n32788, n32789, n32790, n32791, n32792,
    n32793, n32794, n32795, n32796, n32797, n32798, n32799, n32800, n32801,
    n32802, n32803, n32804, n32805, n32806, n32807, n32808, n32809, n32810,
    n32811, n32812, n32813, n32814, n32815, n32816, n32817, n32818, n32819,
    n32820, n32821, n32822, n32823, n32824, n32825, n32826, n32827, n32828,
    n32829, n32830, n32831, n32832, n32833, n32834, n32835, n32836, n32837,
    n32838, n32839, n32840, n32841, n32842, n32843, n32844, n32845, n32846,
    n32847, n32848, n32849, n32850, n32851, n32852, n32853, n32854, n32855,
    n32856, n32857, n32858, n32859, n32860, n32861, n32862, n32863, n32864,
    n32865, n32866, n32867, n32868, n32869, n32870, n32871, n32872, n32873,
    n32874, n32875, n32876, n32877, n32878, n32879, n32880, n32881, n32882,
    n32883, n32884, n32885, n32886, n32887, n32888, n32889, n32890, n32891,
    n32892, n32893, n32894, n32895, n32896, n32897, n32898, n32899, n32900,
    n32901, n32902, n32903, n32904, n32905, n32906, n32907, n32908, n32909,
    n32910, n32911, n32912, n32913, n32914, n32915, n32916, n32917, n32918,
    n32919, n32920, n32921, n32922, n32923, n32924, n32925, n32926, n32927,
    n32928, n32929, n32930, n32931, n32932, n32933, n32934, n32935, n32936,
    n32937, n32938, n32939, n32940, n32941, n32942, n32943, n32944, n32945,
    n32946, n32947, n32948, n32949, n32950, n32951, n32952, n32953, n32954,
    n32955, n32956, n32957, n32958, n32959, n32960, n32961, n32962, n32963,
    n32964, n32965, n32966, n32967, n32968, n32969, n32970, n32971, n32972,
    n32973, n32974, n32975, n32976, n32977, n32978, n32979, n32980, n32981,
    n32982, n32983, n32984, n32985, n32986, n32987, n32988, n32989, n32990,
    n32991, n32992, n32993, n32994, n32995, n32996, n32997, n32998, n32999,
    n33000, n33001, n33002, n33003, n33004, n33005, n33006, n33007, n33008,
    n33009, n33010, n33011, n33012, n33013, n33014, n33015, n33016, n33017,
    n33018, n33019, n33020, n33021, n33022, n33023, n33024, n33025, n33026,
    n33027, n33028, n33029, n33030, n33031, n33032, n33033, n33034, n33035,
    n33036, n33037, n33038, n33039, n33040, n33041, n33042, n33043, n33044,
    n33045, n33046, n33047, n33048, n33049, n33050, n33051, n33052, n33053,
    n33054, n33055, n33056, n33057, n33058, n33059, n33060, n33061, n33062,
    n33063, n33064, n33065, n33066, n33067, n33068, n33069, n33070, n33071,
    n33072, n33073, n33074, n33075, n33076, n33077, n33078, n33079, n33080,
    n33081, n33082, n33083, n33084, n33085, n33086, n33087, n33088, n33089,
    n33090, n33091, n33092, n33093, n33094, n33095, n33096, n33097, n33098,
    n33099, n33100, n33101, n33102, n33103, n33104, n33105, n33106, n33107,
    n33108, n33109, n33110, n33111, n33112, n33113, n33114, n33115, n33116,
    n33117, n33118, n33119, n33120, n33121, n33122, n33123, n33124, n33125,
    n33126, n33127, n33128, n33129, n33130, n33131, n33132, n33133, n33134,
    n33135, n33136, n33137, n33138, n33139, n33140, n33141, n33142, n33143,
    n33144, n33145, n33146, n33147, n33148, n33149, n33150, n33151, n33152,
    n33153, n33154, n33155, n33156, n33157, n33158, n33159, n33160, n33161,
    n33162, n33163, n33164, n33165, n33166, n33167, n33168, n33169, n33170,
    n33171, n33172, n33173, n33174, n33175, n33176, n33177, n33178, n33179,
    n33180, n33181, n33182, n33183, n33184, n33185, n33186, n33187, n33188,
    n33189, n33190, n33191, n33192, n33193, n33194, n33195, n33196, n33197,
    n33198, n33199, n33200, n33201, n33202, n33203, n33204, n33205, n33206,
    n33207, n33208, n33209, n33210, n33211, n33212, n33213, n33214, n33215,
    n33216, n33217, n33218, n33219, n33220, n33221, n33222, n33223, n33224,
    n33225, n33226, n33227, n33228, n33229, n33230, n33231, n33232, n33233,
    n33234, n33235, n33236, n33237, n33238, n33239, n33240, n33241, n33242,
    n33243, n33244, n33245, n33246, n33247, n33248, n33249, n33250, n33251,
    n33252, n33253, n33254, n33255, n33256, n33257, n33258, n33259, n33260,
    n33261, n33262, n33263, n33264, n33265, n33266, n33267, n33268, n33269,
    n33270, n33271, n33272, n33273, n33274, n33275, n33276, n33277, n33278,
    n33279, n33280, n33281, n33282, n33283, n33284, n33285, n33286, n33287,
    n33288, n33289, n33290, n33291, n33292, n33293, n33294, n33295, n33296,
    n33297, n33298, n33299, n33300, n33301, n33302, n33303, n33304, n33305,
    n33306, n33307, n33308, n33309, n33310, n33311, n33312, n33313, n33314,
    n33315, n33316, n33317, n33318, n33319, n33320, n33321, n33322, n33323,
    n33324, n33325, n33326, n33327, n33328, n33329, n33330, n33331, n33332,
    n33333, n33334, n33335, n33336, n33337, n33338, n33339, n33340, n33341,
    n33342, n33343, n33344, n33345, n33346, n33347, n33348, n33349, n33350,
    n33351, n33352, n33353, n33354, n33355, n33356, n33357, n33358, n33359,
    n33360, n33361, n33362, n33363, n33364, n33365, n33366, n33367, n33368,
    n33369, n33370, n33371, n33372, n33373, n33374, n33375, n33376, n33377,
    n33378, n33379, n33380, n33381, n33382, n33383, n33384, n33385, n33386,
    n33387, n33388, n33389, n33390, n33391, n33392, n33393, n33394, n33395,
    n33396, n33397, n33398, n33399, n33400, n33401, n33402, n33403, n33404,
    n33405, n33406, n33407, n33408, n33409, n33410, n33411, n33412, n33413,
    n33414, n33415, n33416, n33417, n33418, n33419, n33420, n33421, n33422,
    n33423, n33424, n33425, n33426, n33427, n33428, n33429, n33430, n33431,
    n33432, n33433, n33434, n33435, n33436, n33437, n33438, n33439, n33440,
    n33441, n33442, n33443, n33444, n33445, n33446, n33447, n33448, n33449,
    n33450, n33451, n33452, n33453, n33454, n33455, n33456, n33457, n33458,
    n33459, n33460, n33461, n33462, n33463, n33464, n33465, n33466, n33467,
    n33468, n33469, n33470, n33471, n33472, n33473, n33474, n33475, n33476,
    n33477, n33478, n33479, n33480, n33481, n33482, n33483, n33484, n33485,
    n33486, n33487, n33488, n33489, n33490, n33491, n33492, n33493, n33494,
    n33495, n33496, n33497, n33498, n33499, n33500, n33501, n33502, n33503,
    n33504, n33505, n33506, n33507, n33508, n33509, n33510, n33511, n33512,
    n33513, n33514, n33515, n33516, n33517, n33518, n33519, n33520, n33521,
    n33522, n33523, n33524, n33525, n33526, n33527, n33528, n33529, n33530,
    n33531, n33532, n33533, n33534, n33535, n33536, n33537, n33538, n33539,
    n33540, n33541, n33542, n33543, n33544, n33545, n33546, n33547, n33548,
    n33549, n33550, n33551, n33552, n33553, n33554, n33555, n33556, n33557,
    n33558, n33559, n33560, n33561, n33562, n33563, n33564, n33565, n33566,
    n33567, n33568, n33569, n33570, n33571, n33572, n33573, n33574, n33575,
    n33576, n33577, n33578, n33579, n33580, n33581, n33582, n33583, n33584,
    n33585, n33586, n33587, n33588, n33589, n33590, n33591, n33592, n33593,
    n33594, n33595, n33596, n33597, n33598, n33599, n33600, n33601, n33602,
    n33603, n33604, n33605, n33606, n33607, n33608, n33609, n33610, n33611,
    n33612, n33613, n33614, n33615, n33616, n33617, n33618, n33619, n33620,
    n33621, n33622, n33623, n33624, n33625, n33626, n33627, n33628, n33629,
    n33630, n33631, n33632, n33633, n33634, n33635, n33636, n33637, n33638,
    n33639, n33640, n33641, n33642, n33643, n33644, n33645, n33646, n33647,
    n33648, n33649, n33650, n33651, n33652, n33653, n33654, n33655, n33656,
    n33657, n33658, n33659, n33660, n33661, n33662, n33663, n33664, n33665,
    n33666, n33667, n33668, n33669, n33670, n33671, n33672, n33673, n33674,
    n33675, n33676, n33677, n33678, n33679, n33680, n33681, n33682, n33683,
    n33684, n33685, n33686, n33687, n33688, n33689, n33690, n33691, n33692,
    n33693, n33694, n33695, n33696, n33697, n33698, n33699, n33700, n33701,
    n33702, n33703, n33704, n33705, n33706, n33707, n33708, n33709, n33710,
    n33711, n33712, n33713, n33714, n33715, n33716, n33717, n33718, n33719,
    n33720, n33721, n33722, n33723, n33724, n33725, n33726, n33727, n33728,
    n33729, n33730, n33731, n33732, n33733, n33734, n33735, n33736, n33737,
    n33738, n33739, n33740, n33741, n33742, n33743, n33744, n33745, n33746,
    n33747, n33748, n33749, n33750, n33751, n33752, n33753, n33754, n33755,
    n33756, n33757, n33758, n33759, n33760, n33761, n33762, n33763, n33764,
    n33765, n33766, n33767, n33768, n33769, n33770, n33771, n33772, n33773,
    n33774, n33775, n33776, n33777, n33778, n33779, n33780, n33781, n33782,
    n33783, n33784, n33785, n33786, n33787, n33788, n33789, n33790, n33791,
    n33792, n33793, n33794, n33795, n33796, n33797, n33798, n33799, n33800,
    n33801, n33802, n33803, n33804, n33805, n33806, n33807, n33808, n33809,
    n33810, n33811, n33812, n33813, n33814, n33815, n33816, n33817, n33818,
    n33819, n33820, n33821, n33822, n33823, n33824, n33825, n33826, n33827,
    n33828, n33829, n33830, n33831, n33832, n33833, n33834, n33835, n33836,
    n33837, n33838, n33839, n33840, n33841, n33842, n33843, n33844, n33845,
    n33846, n33847, n33848, n33849, n33850, n33851, n33852, n33853, n33854,
    n33855, n33856, n33857, n33858, n33859, n33860, n33861, n33862, n33863,
    n33864, n33865, n33866, n33867, n33868, n33869, n33870, n33871, n33872,
    n33873, n33874, n33875, n33876, n33877, n33878, n33879, n33880, n33881,
    n33882, n33883, n33884, n33885, n33886, n33887, n33888, n33889, n33890,
    n33891, n33892, n33893, n33894, n33895, n33896, n33897, n33898, n33899,
    n33900, n33901, n33902, n33903, n33904, n33905, n33906, n33907, n33908,
    n33909, n33910, n33911, n33912, n33913, n33914, n33915, n33916, n33917,
    n33918, n33919, n33920, n33921, n33922, n33923, n33924, n33925, n33926,
    n33927, n33928, n33929, n33930, n33931, n33932, n33933, n33934, n33935,
    n33936, n33937, n33938, n33939, n33940, n33941, n33942, n33943, n33944,
    n33945, n33946, n33947, n33948, n33949, n33950, n33951, n33952, n33953,
    n33954, n33955, n33956, n33957, n33958, n33959, n33960, n33961, n33962,
    n33963, n33964, n33965, n33966, n33967, n33968, n33969, n33970, n33971,
    n33972, n33973, n33974, n33975, n33976, n33977, n33978, n33979, n33980,
    n33981, n33982, n33983, n33984, n33985, n33986, n33987, n33988, n33989,
    n33990, n33991, n33992, n33993, n33994, n33995, n33996, n33997, n33998,
    n33999, n34000, n34001, n34002, n34003, n34004, n34005, n34006, n34007,
    n34008, n34009, n34010, n34011, n34012, n34013, n34014, n34015, n34016,
    n34017, n34018, n34019, n34020, n34021, n34022, n34023, n34024, n34025,
    n34026, n34027, n34028, n34029, n34030, n34031, n34032, n34033, n34034,
    n34035, n34036, n34037, n34038, n34039, n34040, n34041, n34042, n34043,
    n34044, n34045, n34046, n34047, n34048, n34049, n34050, n34051, n34052,
    n34053, n34054, n34055, n34056, n34057, n34058, n34059, n34060, n34061,
    n34062, n34063, n34064, n34065, n34066, n34067, n34068, n34069, n34070,
    n34071, n34072, n34073, n34074, n34075, n34076, n34077, n34078, n34079,
    n34080, n34081, n34082, n34083, n34084, n34085, n34086, n34087, n34088,
    n34089, n34090, n34091, n34092, n34093, n34094, n34095, n34096, n34097,
    n34098, n34099, n34100, n34101, n34102, n34103, n34104, n34105, n34106,
    n34107, n34108, n34109, n34110, n34111, n34112, n34113, n34114, n34115,
    n34116, n34117, n34118, n34119, n34120, n34121, n34122, n34123, n34124,
    n34125, n34126, n34127, n34128, n34129, n34130, n34131, n34132, n34133,
    n34134, n34135, n34136, n34137, n34138, n34139, n34140, n34141, n34142,
    n34143, n34144, n34145, n34146, n34147, n34148, n34149, n34150, n34151,
    n34152, n34153, n34154, n34155, n34156, n34157, n34158, n34159, n34160,
    n34161, n34162, n34163, n34164, n34165, n34166, n34167, n34168, n34169,
    n34170, n34171, n34172, n34173, n34174, n34175, n34176, n34177, n34178,
    n34179, n34180, n34181, n34182, n34183, n34184, n34185, n34186, n34187,
    n34188, n34189, n34190, n34191, n34192, n34193, n34194, n34195, n34196,
    n34197, n34198, n34199, n34200, n34201, n34202, n34203, n34204, n34205,
    n34206, n34207, n34208, n34209, n34210, n34211, n34212, n34213, n34214,
    n34215, n34216, n34217, n34218, n34219, n34220, n34221, n34222, n34223,
    n34224, n34225, n34226, n34227, n34228, n34229, n34230, n34231, n34232,
    n34233, n34234, n34235, n34236, n34237, n34238, n34239, n34240, n34241,
    n34242, n34243, n34244, n34245, n34246, n34247, n34248, n34249, n34250,
    n34251, n34252, n34253, n34254, n34255, n34256, n34257, n34258, n34259,
    n34260, n34261, n34262, n34263, n34264, n34265, n34266, n34267, n34268,
    n34269, n34270, n34271, n34272, n34273, n34274, n34275, n34276, n34277,
    n34278, n34279, n34280, n34281, n34282, n34283, n34284, n34285, n34286,
    n34287, n34288, n34289, n34290, n34291, n34292, n34293, n34294, n34295,
    n34296, n34297, n34298, n34299, n34300, n34301, n34302, n34303, n34304,
    n34305, n34306, n34307, n34308, n34309, n34310, n34311, n34312, n34313,
    n34314, n34315, n34316, n34317, n34318, n34319, n34320, n34321, n34322,
    n34323, n34324, n34325, n34326, n34327, n34328, n34329, n34330, n34331,
    n34332, n34333, n34334, n34335, n34336, n34337, n34338, n34339, n34340,
    n34341, n34342, n34343, n34344, n34345, n34346, n34347, n34348, n34349,
    n34350, n34351, n34352, n34353, n34354, n34355, n34356, n34357, n34358,
    n34359, n34360, n34361, n34362, n34363, n34364, n34365, n34366, n34367,
    n34368, n34369, n34370, n34371, n34372, n34373, n34374, n34375, n34376,
    n34377, n34378, n34379, n34380, n34381, n34382, n34383, n34384, n34385,
    n34386, n34387, n34388, n34389, n34390, n34391, n34392, n34393, n34394,
    n34395, n34396, n34397, n34398, n34399, n34400, n34401, n34402, n34403,
    n34404, n34405, n34406, n34407, n34408, n34409, n34410, n34411, n34412,
    n34413, n34414, n34415, n34416, n34417, n34418, n34419, n34420, n34421,
    n34422, n34423, n34424, n34425, n34426, n34427, n34428, n34429, n34430,
    n34431, n34432, n34433, n34434, n34435, n34436, n34437, n34438, n34439,
    n34440, n34441, n34442, n34443, n34444, n34445, n34446, n34447, n34448,
    n34449, n34450, n34451, n34452, n34453, n34454, n34455, n34456, n34457,
    n34458, n34459, n34460, n34461, n34462, n34463, n34464, n34465, n34466,
    n34467, n34468, n34469, n34470, n34471, n34472, n34473, n34474, n34475,
    n34476, n34477, n34478, n34479, n34480, n34481, n34482, n34483, n34484,
    n34485, n34486, n34487, n34488, n34489, n34490, n34491, n34492, n34493,
    n34494, n34495, n34496, n34497, n34498, n34499, n34500, n34501, n34502,
    n34503, n34504, n34505, n34506, n34507, n34508, n34509, n34510, n34511,
    n34512, n34513, n34514, n34515, n34516, n34517, n34518, n34519, n34520,
    n34521, n34522, n34523, n34524, n34525, n34526, n34527, n34528, n34529,
    n34530, n34531, n34532, n34533, n34534, n34535, n34536, n34537, n34538,
    n34539, n34540, n34541, n34542, n34543, n34544, n34545, n34546, n34547,
    n34548, n34549, n34550, n34551, n34552, n34553, n34554, n34555, n34556,
    n34557, n34558, n34559, n34560, n34561, n34562, n34563, n34564, n34565,
    n34566, n34567, n34568, n34569, n34570, n34571, n34572, n34573, n34574,
    n34575, n34576, n34577, n34578, n34579, n34580, n34581, n34582, n34583,
    n34584, n34585, n34586, n34587, n34588, n34589, n34590, n34591, n34592,
    n34593, n34594, n34595, n34596, n34597, n34598, n34599, n34600, n34601,
    n34602, n34603, n34604, n34605, n34606, n34607, n34608, n34609, n34610,
    n34611, n34612, n34613, n34614, n34615, n34616, n34617, n34618, n34619,
    n34620, n34621, n34622, n34623, n34624, n34625, n34626, n34627, n34628,
    n34629, n34630, n34631, n34632, n34633, n34634, n34635, n34636, n34637,
    n34638, n34639, n34640, n34641, n34642, n34643, n34644, n34645, n34646,
    n34647, n34648, n34649, n34650, n34651, n34652, n34653, n34654, n34655,
    n34656, n34657, n34658, n34659, n34660, n34661, n34662, n34663, n34664,
    n34665, n34666, n34667, n34668, n34669, n34670, n34671, n34672, n34673,
    n34674, n34675, n34676, n34677, n34678, n34679, n34680, n34681, n34682,
    n34683, n34684, n34685, n34686, n34687, n34688, n34689, n34690, n34691,
    n34692, n34693, n34694, n34695, n34696, n34697, n34698, n34699, n34700,
    n34701, n34702, n34703, n34704, n34705, n34706, n34707, n34708, n34709,
    n34710, n34711, n34712, n34713, n34714, n34715, n34716, n34717, n34718,
    n34719, n34720, n34721, n34722, n34723, n34724, n34725, n34726, n34727,
    n34728, n34729, n34730, n34731, n34732, n34733, n34734, n34735, n34736,
    n34737, n34738, n34739, n34740, n34741, n34742, n34743, n34744, n34745,
    n34746, n34747, n34748, n34749, n34750, n34751, n34752, n34753, n34754,
    n34755, n34756, n34757, n34758, n34759, n34760, n34761, n34762, n34763,
    n34764, n34765, n34766, n34767, n34768, n34769, n34770, n34771, n34772,
    n34773, n34774, n34775, n34776, n34777, n34778, n34779, n34780, n34781,
    n34782, n34783, n34784, n34785, n34786, n34787, n34788, n34789, n34790,
    n34791, n34792, n34793, n34794, n34795, n34796, n34797, n34798, n34799,
    n34800, n34801, n34802, n34803, n34804, n34805, n34806, n34807, n34808,
    n34809, n34810, n34811, n34812, n34813, n34814, n34815, n34816, n34817,
    n34818, n34819, n34820, n34821, n34822, n34823, n34824, n34825, n34826,
    n34827, n34828, n34829, n34830, n34831, n34832, n34833, n34834, n34835,
    n34836, n34837, n34838, n34839, n34840, n34841, n34842, n34843, n34844,
    n34845, n34846, n34847, n34848, n34849, n34850, n34851, n34852, n34853,
    n34854, n34855, n34856, n34857, n34858, n34859, n34860, n34861, n34862,
    n34863, n34864, n34865, n34866, n34867, n34868, n34869, n34870, n34871,
    n34872, n34873, n34874, n34875, n34876, n34877, n34878, n34879, n34880,
    n34881, n34882, n34883, n34884, n34885, n34886, n34887, n34888, n34889,
    n34890, n34891, n34892, n34893, n34894, n34895, n34896, n34897, n34898,
    n34899, n34900, n34901, n34902, n34903, n34904, n34905, n34906, n34907,
    n34908, n34909, n34910, n34911, n34912, n34913, n34914, n34915, n34916,
    n34917, n34918, n34919, n34920, n34921, n34922, n34923, n34924, n34925,
    n34926, n34927, n34928, n34929, n34930, n34931, n34932, n34933, n34934,
    n34935, n34936, n34937, n34938, n34939, n34940, n34941, n34942, n34943,
    n34944, n34945, n34946, n34947, n34948, n34949, n34950, n34951, n34952,
    n34953, n34954, n34955, n34956, n34957, n34958, n34959, n34960, n34961,
    n34962, n34963, n34964, n34965, n34966, n34967, n34968, n34969, n34970,
    n34971, n34972, n34973, n34974, n34975, n34976, n34977, n34978, n34979,
    n34980, n34981, n34982, n34983, n34984, n34985, n34986, n34987, n34988,
    n34989, n34990, n34991, n34992, n34993, n34994, n34995, n34996, n34997,
    n34998, n34999, n35000, n35001, n35002, n35003, n35004, n35005, n35006,
    n35007, n35008, n35009, n35010, n35011, n35012, n35013, n35014, n35015,
    n35016, n35017, n35018, n35019, n35020, n35021, n35022, n35023, n35024,
    n35025, n35026, n35027, n35028, n35029, n35030, n35031, n35032, n35033,
    n35034, n35035, n35036, n35037, n35038, n35039, n35040, n35041, n35042,
    n35043, n35044, n35045, n35046, n35047, n35048, n35049, n35050, n35051,
    n35052, n35053, n35054, n35055, n35056, n35057, n35058, n35059, n35060,
    n35061, n35062, n35063, n35064, n35065, n35066, n35067, n35068, n35069,
    n35070, n35071, n35072, n35073, n35074, n35075, n35076, n35077, n35078,
    n35079, n35080, n35081, n35082, n35083, n35084, n35085, n35086, n35087,
    n35088, n35089, n35090, n35091, n35092, n35093, n35094, n35095, n35096,
    n35097, n35098, n35099, n35100, n35101, n35102, n35103, n35104, n35105,
    n35106, n35107, n35108, n35109, n35110, n35111, n35112, n35113, n35114,
    n35115, n35116, n35117, n35118, n35119, n35120, n35121, n35122, n35123,
    n35124, n35125, n35126, n35127, n35128, n35129, n35130, n35131, n35132,
    n35133, n35134, n35135, n35136, n35137, n35138, n35139, n35140, n35141,
    n35142, n35143, n35144, n35145, n35146, n35147, n35148, n35149, n35150,
    n35151, n35152, n35153, n35154, n35155, n35156, n35157, n35158, n35159,
    n35160, n35161, n35162, n35163, n35164, n35165, n35166, n35167, n35168,
    n35169, n35170, n35171, n35172, n35173, n35174, n35175, n35176, n35177,
    n35178, n35179, n35180, n35181, n35182, n35183, n35184, n35185, n35186,
    n35187, n35188, n35189, n35190, n35191, n35192, n35193, n35194, n35195,
    n35196, n35197, n35198, n35199, n35200, n35201, n35202, n35203, n35204,
    n35205, n35206, n35207, n35208, n35209, n35210, n35211, n35212, n35213,
    n35214, n35215, n35216, n35217, n35218, n35219, n35220, n35221, n35222,
    n35223, n35224, n35225, n35226, n35227, n35228, n35229, n35230, n35231,
    n35232, n35233, n35234, n35235, n35236, n35237, n35238, n35239, n35240,
    n35241, n35242, n35243, n35244, n35245, n35246, n35247, n35248, n35249,
    n35250, n35251, n35252, n35253, n35254, n35255, n35256, n35257, n35258,
    n35259, n35260, n35261, n35262, n35263, n35264, n35265, n35266, n35267,
    n35268, n35269, n35270, n35271, n35272, n35273, n35274, n35275, n35276,
    n35277, n35278, n35279, n35280, n35281, n35282, n35283, n35284, n35285,
    n35286, n35287, n35288, n35289, n35290, n35291, n35292, n35293, n35294,
    n35295, n35296, n35297, n35298, n35299, n35300, n35301, n35302, n35303,
    n35304, n35305, n35306, n35307, n35308, n35309, n35310, n35311, n35312,
    n35313, n35314, n35315, n35316, n35317, n35318, n35319, n35320, n35321,
    n35322, n35323, n35324, n35325, n35326, n35327, n35328, n35329, n35330,
    n35331, n35332, n35333, n35334, n35335, n35336, n35337, n35338, n35339,
    n35340, n35341, n35342, n35343, n35344, n35345, n35346, n35347, n35348,
    n35349, n35350, n35351, n35352, n35353, n35354, n35355, n35356, n35357,
    n35358, n35359, n35360, n35361, n35362, n35363, n35364, n35365, n35366,
    n35367, n35368, n35369, n35370, n35371, n35372, n35373, n35374, n35375,
    n35376, n35377, n35378, n35379, n35380, n35381, n35382, n35383, n35384,
    n35385, n35386, n35387, n35388, n35389, n35390, n35391, n35392, n35393,
    n35394, n35395, n35396, n35397, n35398, n35399, n35400, n35401, n35402,
    n35403, n35404, n35405, n35406, n35407, n35408, n35409, n35410, n35411,
    n35412, n35413, n35414, n35415, n35416, n35417, n35418, n35419, n35420,
    n35421, n35422, n35423, n35424, n35425, n35426, n35427, n35428, n35429,
    n35430, n35431, n35432, n35433, n35434, n35435, n35436, n35437, n35438,
    n35439, n35440, n35441, n35442, n35443, n35444, n35445, n35446, n35447,
    n35448, n35449, n35450, n35451, n35452, n35453, n35454, n35455, n35456,
    n35457, n35458, n35459, n35460, n35461, n35462, n35463, n35464, n35465,
    n35466, n35467, n35468, n35469, n35470, n35471, n35472, n35473, n35474,
    n35475, n35476, n35477, n35478, n35479, n35480, n35481, n35482, n35483,
    n35484, n35485, n35486, n35487, n35488, n35489, n35490, n35491, n35492,
    n35493, n35494, n35495, n35496, n35497, n35498, n35499, n35500, n35501,
    n35502, n35503, n35504, n35505, n35506, n35507, n35508, n35509, n35510,
    n35511, n35512, n35513, n35514, n35515, n35516, n35517, n35518, n35519,
    n35520, n35521, n35522, n35523, n35524, n35525, n35526, n35527, n35528,
    n35529, n35530, n35531, n35532, n35533, n35534, n35535, n35536, n35537,
    n35538, n35539, n35540, n35541, n35542, n35543, n35544, n35545, n35546,
    n35547, n35548, n35549, n35550, n35551, n35552, n35553, n35554, n35555,
    n35556, n35557, n35558, n35559, n35560, n35561, n35562, n35563, n35564,
    n35565, n35566, n35567, n35568, n35569, n35570, n35571, n35572, n35573,
    n35574, n35575, n35576, n35577, n35578, n35579, n35580, n35581, n35582,
    n35583, n35584, n35585, n35586, n35587, n35588, n35589, n35590, n35591,
    n35592, n35593, n35594, n35595, n35596, n35597, n35598, n35599, n35600,
    n35601, n35602, n35603, n35604, n35605, n35606, n35607, n35608, n35609,
    n35610, n35611, n35612, n35613, n35614, n35615, n35616, n35617, n35618,
    n35619, n35620, n35621, n35622, n35623, n35624, n35625, n35626, n35627,
    n35628, n35629, n35630, n35631, n35632, n35633, n35634, n35635, n35636,
    n35637, n35638, n35639, n35640, n35641, n35642, n35643, n35644, n35645,
    n35646, n35647, n35648, n35649, n35650, n35651, n35652, n35653, n35654,
    n35655, n35656, n35657, n35658, n35659, n35660, n35661, n35662, n35663,
    n35664, n35665, n35666, n35667, n35668, n35669, n35670, n35671, n35672,
    n35673, n35674, n35675, n35676, n35677, n35678, n35679, n35680, n35681,
    n35682, n35683, n35684, n35685, n35686, n35687, n35688, n35689, n35690,
    n35691, n35692, n35693, n35694, n35695, n35696, n35697, n35698, n35699,
    n35700, n35701, n35702, n35703, n35704, n35705, n35706, n35707, n35708,
    n35709, n35710, n35711, n35712, n35713, n35714, n35715, n35716, n35717,
    n35718, n35719, n35720, n35721, n35722, n35723, n35724, n35725, n35726,
    n35727, n35728, n35729, n35730, n35731, n35732, n35733, n35734, n35735,
    n35736, n35737, n35738, n35739, n35740, n35741, n35742, n35743, n35744,
    n35745, n35746, n35747, n35748, n35749, n35750, n35751, n35752, n35753,
    n35754, n35755, n35756, n35757, n35758, n35759, n35760, n35761, n35762,
    n35763, n35764, n35765, n35766, n35767, n35768, n35769, n35770, n35771,
    n35772, n35773, n35774, n35775, n35776, n35777, n35778, n35779, n35780,
    n35781, n35782, n35783, n35784, n35785, n35786, n35787, n35788, n35789,
    n35790, n35791, n35792, n35793, n35794, n35795, n35796, n35797, n35798,
    n35799, n35800, n35801, n35802, n35803, n35804, n35805, n35806, n35807,
    n35808, n35809, n35810, n35811, n35812, n35813, n35814, n35815, n35816,
    n35817, n35818, n35819, n35820, n35821, n35822, n35823, n35824, n35825,
    n35826, n35827, n35828, n35829, n35830, n35831, n35832, n35833, n35834,
    n35835, n35836, n35837, n35838, n35839, n35840, n35841, n35842, n35843,
    n35844, n35845, n35846, n35847, n35848, n35849, n35850, n35851, n35852,
    n35853, n35854, n35855, n35856, n35857, n35858, n35859, n35860, n35861,
    n35862, n35863, n35864, n35865, n35866, n35867, n35868, n35869, n35870,
    n35871, n35872, n35873, n35874, n35875, n35876, n35877, n35878, n35879,
    n35880, n35881, n35882, n35883, n35884, n35885, n35886, n35887, n35888,
    n35889, n35890, n35891, n35892, n35893, n35894, n35895, n35896, n35897,
    n35898, n35899, n35900, n35901, n35902, n35903, n35904, n35905, n35906,
    n35907, n35908, n35909, n35910, n35911, n35912, n35913, n35914, n35915,
    n35916, n35917, n35918, n35919, n35920, n35921, n35922, n35923, n35924,
    n35925, n35926, n35927, n35928, n35929, n35930, n35931, n35932, n35933,
    n35934, n35935, n35936, n35937, n35938, n35939, n35940, n35941, n35942,
    n35943, n35944, n35945, n35946, n35947, n35948, n35949, n35950, n35951,
    n35952, n35953, n35954, n35955, n35956, n35957, n35958, n35959, n35960,
    n35961, n35962, n35963, n35964, n35965, n35966, n35967, n35968, n35969,
    n35970, n35971, n35972, n35973, n35974, n35975, n35976, n35977, n35978,
    n35979, n35980, n35981, n35982, n35983, n35984, n35985, n35986, n35987,
    n35988, n35989, n35990, n35991, n35992, n35993, n35994, n35995, n35996,
    n35997, n35998, n35999, n36000, n36001, n36002, n36003, n36004, n36005,
    n36006, n36007, n36008, n36009, n36010, n36011, n36012, n36013, n36014,
    n36015, n36016, n36017, n36018, n36019, n36020, n36021, n36022, n36023,
    n36024, n36025, n36026, n36027, n36028, n36029, n36030, n36031, n36032,
    n36033, n36034, n36035, n36036, n36037, n36038, n36039, n36040, n36041,
    n36042, n36043, n36044, n36045, n36046, n36047, n36048, n36049, n36050,
    n36051, n36052, n36053, n36054, n36055, n36056, n36057, n36058, n36059,
    n36060, n36061, n36062, n36063, n36064, n36065, n36066, n36067, n36068,
    n36069, n36070, n36071, n36072, n36073, n36074, n36075, n36076, n36077,
    n36078, n36079, n36080, n36081, n36082, n36083, n36084, n36085, n36086,
    n36087, n36088, n36089, n36090, n36091, n36092, n36093, n36094, n36095,
    n36096, n36097, n36098, n36099, n36100, n36101, n36102, n36103, n36104,
    n36105, n36106, n36107, n36108, n36109, n36110, n36111, n36112, n36113,
    n36114, n36115, n36116, n36117, n36118, n36119, n36120, n36121, n36122,
    n36123, n36124, n36125, n36126, n36127, n36128, n36129, n36130, n36131,
    n36132, n36133, n36134, n36135, n36136, n36137, n36138, n36139, n36140,
    n36141, n36142, n36143, n36144, n36145, n36146, n36147, n36148, n36149,
    n36150, n36151, n36152, n36153, n36154, n36155, n36156, n36157, n36158,
    n36159, n36160, n36161, n36162, n36163, n36164, n36165, n36166, n36167,
    n36168, n36169, n36170, n36171, n36172, n36173, n36174, n36175, n36176,
    n36177, n36178, n36179, n36180, n36181, n36182, n36183, n36184, n36185,
    n36186, n36187, n36188, n36189, n36190, n36191, n36192, n36193, n36194,
    n36195, n36196, n36197, n36198, n36199, n36200, n36201, n36202, n36203,
    n36204, n36205, n36206, n36207, n36208, n36209, n36210, n36211, n36212,
    n36213, n36214, n36215, n36216, n36217, n36218, n36219, n36220, n36221,
    n36222, n36223, n36224, n36225, n36226, n36227, n36228, n36229, n36230,
    n36231, n36232, n36233, n36234, n36235, n36236, n36237, n36238, n36239,
    n36240, n36241, n36242, n36243, n36244, n36245, n36246, n36247, n36248,
    n36249, n36250, n36251, n36252, n36253, n36254, n36255, n36256, n36257,
    n36258, n36259, n36260, n36261, n36262, n36263, n36264, n36265, n36266,
    n36267, n36268, n36269, n36270, n36271, n36272, n36273, n36274, n36275,
    n36276, n36277, n36278, n36279, n36280, n36281, n36282, n36283, n36284,
    n36285, n36286, n36287, n36288, n36289, n36290, n36291, n36292, n36293,
    n36294, n36295, n36296, n36297, n36298, n36299, n36300, n36301, n36302,
    n36303, n36304, n36305, n36306, n36307, n36308, n36309, n36310, n36311,
    n36312, n36313, n36314, n36315, n36316, n36317, n36318, n36319, n36320,
    n36321, n36322, n36323, n36324, n36325, n36326, n36327, n36328, n36329,
    n36330, n36331, n36332, n36333, n36334, n36335, n36336, n36337, n36338,
    n36339, n36340, n36341, n36342, n36343, n36344, n36345, n36346, n36347,
    n36348, n36349, n36350, n36351, n36352, n36353, n36354, n36355, n36356,
    n36357, n36358, n36359, n36360, n36361, n36362, n36363, n36364, n36365,
    n36366, n36367, n36368, n36369, n36370, n36371, n36372, n36373, n36374,
    n36375, n36376, n36377, n36378, n36379, n36380, n36381, n36382, n36383,
    n36384, n36385, n36386, n36387, n36388, n36389, n36390, n36391, n36392,
    n36393, n36394, n36395, n36396, n36397, n36398, n36399, n36400, n36401,
    n36402, n36403, n36404, n36405, n36406, n36407, n36408, n36409, n36410,
    n36411, n36412, n36413, n36414, n36415, n36416, n36417, n36418, n36419,
    n36420, n36421, n36422, n36423, n36424, n36425, n36426, n36427, n36428,
    n36429, n36430, n36431, n36432, n36433, n36434, n36435, n36436, n36437,
    n36438, n36439, n36440, n36441, n36442, n36443, n36444, n36445, n36446,
    n36447, n36448, n36449, n36450, n36451, n36452, n36453, n36454, n36455,
    n36456, n36457, n36458, n36459, n36460, n36461, n36462, n36463, n36464,
    n36465, n36466, n36467, n36468, n36469, n36470, n36471, n36472, n36473,
    n36474, n36475, n36476, n36477, n36478, n36479, n36480, n36481, n36482,
    n36483, n36484, n36485, n36486, n36487, n36488, n36489, n36490, n36491,
    n36492, n36493, n36494, n36495, n36496, n36497, n36498, n36499, n36500,
    n36501, n36502, n36503, n36504, n36505, n36506, n36507, n36508, n36509,
    n36510, n36511, n36512, n36513, n36514, n36515, n36516, n36517, n36518,
    n36519, n36520, n36521, n36522, n36523, n36524, n36525, n36526, n36527,
    n36528, n36529, n36530, n36531, n36532, n36533, n36534, n36535, n36536,
    n36537, n36538, n36539, n36540, n36541, n36542, n36543, n36544, n36545,
    n36546, n36547, n36548, n36549, n36550, n36551, n36552, n36553, n36554,
    n36555, n36556, n36557, n36558, n36559, n36560, n36561, n36562, n36563,
    n36564, n36565, n36566, n36567, n36568, n36569, n36570, n36571, n36572,
    n36573, n36574, n36575, n36576, n36577, n36578, n36579, n36580, n36581,
    n36582, n36583, n36584, n36585, n36586, n36587, n36588, n36589, n36590,
    n36591, n36592, n36593, n36594, n36595, n36596, n36597, n36598, n36599,
    n36600, n36601, n36602, n36603, n36604, n36605, n36606, n36607, n36608,
    n36609, n36610, n36611, n36612, n36613, n36614, n36615, n36616, n36617,
    n36618, n36619, n36620, n36621, n36622, n36623, n36624, n36625, n36626,
    n36627, n36628, n36629, n36630, n36631, n36632, n36633, n36634, n36635,
    n36636, n36637, n36638, n36639, n36640, n36641, n36642, n36643, n36644,
    n36645, n36646, n36647, n36648, n36649, n36650, n36651, n36652, n36653,
    n36654, n36655, n36656, n36657, n36658, n36659, n36660, n36661, n36662,
    n36663, n36664, n36665, n36666, n36667, n36668, n36669, n36670, n36671,
    n36672, n36673, n36674, n36675, n36676, n36677, n36678, n36679, n36680,
    n36681, n36682, n36683, n36684, n36685, n36686, n36687, n36688, n36689,
    n36690, n36691, n36692, n36693, n36694, n36695, n36696, n36697, n36698,
    n36699, n36700, n36701, n36702, n36703, n36704, n36705, n36706, n36707,
    n36708, n36709, n36710, n36711, n36712, n36713, n36714, n36715, n36716,
    n36717, n36718, n36719, n36720, n36721, n36722, n36723, n36724, n36725,
    n36726, n36727, n36728, n36729, n36730, n36731, n36732, n36733, n36734,
    n36735, n36736, n36737, n36738, n36739, n36740, n36741, n36742, n36743,
    n36744, n36745, n36746, n36747, n36748, n36749, n36750, n36751, n36752,
    n36753, n36754, n36755, n36756, n36757, n36758, n36759, n36760, n36761,
    n36762, n36763, n36764, n36765, n36766, n36767, n36768, n36769, n36770,
    n36771, n36772, n36773, n36774, n36775, n36776, n36777, n36778, n36779,
    n36780, n36781, n36782, n36783, n36784, n36785, n36786, n36787, n36788,
    n36789, n36790, n36791, n36792, n36793, n36794, n36795, n36796, n36797,
    n36798, n36799, n36800, n36801, n36802, n36803, n36804, n36805, n36806,
    n36807, n36808, n36809, n36810, n36811, n36812, n36813, n36814, n36815,
    n36816, n36817, n36818, n36819, n36820, n36821, n36822, n36823, n36824,
    n36825, n36826, n36827, n36828, n36829, n36830, n36831, n36832, n36833,
    n36834, n36835, n36836, n36837, n36838, n36839, n36840, n36841, n36842,
    n36843, n36844, n36845, n36846, n36847, n36848, n36849, n36850, n36851,
    n36852, n36853, n36854, n36855, n36856, n36857, n36858, n36859, n36860,
    n36861, n36862, n36863, n36864, n36865, n36866, n36867, n36868, n36869,
    n36870, n36871, n36872, n36873, n36874, n36875, n36876, n36877, n36878,
    n36879, n36880, n36881, n36882, n36883, n36884, n36885, n36886, n36887,
    n36888, n36889, n36890, n36891, n36892, n36893, n36894, n36895, n36896,
    n36897, n36898, n36899, n36900, n36901, n36902, n36903, n36904, n36905,
    n36906, n36907, n36908, n36909, n36910, n36911, n36912, n36913, n36914,
    n36915, n36916, n36917, n36918, n36919, n36920, n36921, n36922, n36923,
    n36924, n36925, n36926, n36927, n36928, n36929, n36930, n36931, n36932,
    n36933, n36934, n36935, n36936, n36937, n36938, n36939, n36940, n36941,
    n36942, n36943, n36944, n36945, n36946, n36947, n36948, n36949, n36950,
    n36951, n36952, n36953, n36954, n36955, n36956, n36957, n36958, n36959,
    n36960, n36961, n36962, n36963, n36964, n36965, n36966, n36967, n36968,
    n36969, n36970, n36971, n36972, n36973, n36974, n36975, n36976, n36977,
    n36978, n36979, n36980, n36981, n36982, n36983, n36984, n36985, n36986,
    n36987, n36988, n36989, n36990, n36991, n36992, n36993, n36994, n36995,
    n36996, n36997, n36998, n36999, n37000, n37001, n37002, n37003, n37004,
    n37005, n37006, n37007, n37008, n37009, n37010, n37011, n37012, n37013,
    n37014, n37015, n37016, n37017, n37018, n37019, n37020, n37021, n37022,
    n37023, n37024, n37025, n37026, n37027, n37028, n37029, n37030, n37031,
    n37032, n37033, n37034, n37035, n37036, n37037, n37038, n37039, n37040,
    n37041, n37042, n37043, n37044, n37045, n37046, n37047, n37048, n37049,
    n37050, n37051, n37052, n37053, n37054, n37055, n37056, n37057, n37058,
    n37059, n37060, n37061, n37062, n37063, n37064, n37065, n37066, n37067,
    n37068, n37069, n37070, n37071, n37072, n37073, n37074, n37075, n37076,
    n37077, n37078, n37079, n37080, n37081, n37082, n37083, n37084, n37085,
    n37086, n37087, n37088, n37089, n37090, n37091, n37092, n37093, n37094,
    n37095, n37096, n37097, n37098, n37099, n37100, n37101, n37102, n37103,
    n37104, n37105, n37106, n37107, n37108, n37109, n37110, n37111, n37112,
    n37113, n37114, n37115, n37116, n37117, n37118, n37119, n37120, n37121,
    n37122, n37123, n37124, n37125, n37126, n37127, n37128, n37129, n37130,
    n37131, n37132, n37133, n37134, n37135, n37136, n37137, n37138, n37139,
    n37140, n37141, n37142, n37143, n37144, n37145, n37146, n37147, n37148,
    n37149, n37150, n37151, n37152, n37153, n37154, n37155, n37156, n37157,
    n37158, n37159, n37160, n37161, n37162, n37163, n37164, n37165, n37166,
    n37167, n37168, n37169, n37170, n37171, n37172, n37173, n37174, n37175,
    n37176, n37177, n37178, n37179, n37180, n37181, n37182, n37183, n37184,
    n37185, n37186, n37187, n37188, n37189, n37190, n37191, n37192, n37193,
    n37194, n37195, n37196, n37197, n37198, n37199, n37200, n37201, n37202,
    n37203, n37204, n37205, n37206, n37207, n37208, n37209, n37210, n37211,
    n37212, n37213, n37214, n37215, n37216, n37217, n37218, n37219, n37220,
    n37221, n37222, n37223, n37224, n37225, n37226, n37227, n37228, n37229,
    n37230, n37231, n37232, n37233, n37234, n37235, n37236, n37237, n37238,
    n37239, n37240, n37241, n37242, n37243, n37244, n37245, n37246, n37247,
    n37248, n37249, n37250, n37251, n37252, n37253, n37254, n37255, n37256,
    n37257, n37258, n37259, n37260, n37261, n37262, n37263, n37264, n37265,
    n37266, n37267, n37268, n37269, n37270, n37271, n37272, n37273, n37274,
    n37275, n37276, n37277, n37278, n37279, n37280, n37281, n37282, n37283,
    n37284, n37285, n37286, n37287, n37288, n37289, n37290, n37291, n37292,
    n37293, n37294, n37295, n37296, n37297, n37298, n37299, n37300, n37301,
    n37302, n37303, n37304, n37305, n37306, n37307, n37308, n37309, n37310,
    n37311, n37312, n37313, n37314, n37315, n37316, n37317, n37318, n37319,
    n37320, n37321, n37322, n37323, n37324, n37325, n37326, n37327, n37328,
    n37329, n37330, n37331, n37332, n37333, n37334, n37335, n37336, n37337,
    n37338, n37339, n37340, n37341, n37342, n37343, n37344, n37345, n37346,
    n37347, n37348, n37349, n37350, n37351, n37352, n37353, n37354, n37355,
    n37356, n37357, n37358, n37359, n37360, n37361, n37362, n37363, n37364,
    n37365, n37366, n37367, n37368, n37369, n37370, n37371, n37372, n37373,
    n37374, n37375, n37376, n37377, n37378, n37379, n37380, n37381, n37382,
    n37383, n37384, n37385, n37386, n37387, n37388, n37389, n37390, n37391,
    n37392, n37393, n37394, n37395, n37396, n37397, n37398, n37399, n37400,
    n37401, n37402, n37403, n37404, n37405, n37406, n37407, n37408, n37409,
    n37410, n37411, n37412, n37413, n37414, n37415, n37416, n37417, n37418,
    n37419, n37420, n37421, n37422, n37423, n37424, n37425, n37426, n37427,
    n37428, n37429, n37430, n37431, n37432, n37433, n37434, n37435, n37436,
    n37437, n37438, n37439, n37440, n37441, n37442, n37443, n37444, n37445,
    n37446, n37447, n37448, n37449, n37450, n37451, n37452, n37453, n37454,
    n37455, n37456, n37457, n37458, n37459, n37460, n37461, n37462, n37463,
    n37464, n37465, n37466, n37467, n37468, n37469, n37470, n37471, n37472,
    n37473, n37474, n37475, n37476, n37477, n37478, n37479, n37480, n37481,
    n37482, n37483, n37484, n37485, n37486, n37487, n37488, n37489, n37490,
    n37491, n37492, n37493, n37494, n37495, n37496, n37497, n37498, n37499,
    n37500, n37501, n37502, n37503, n37504, n37505, n37506, n37507, n37508,
    n37509, n37510, n37511, n37512, n37513, n37514, n37515, n37516, n37517,
    n37518, n37519, n37520, n37521, n37522, n37523, n37524, n37525, n37526,
    n37527, n37528, n37529, n37530, n37531, n37532, n37533, n37534, n37535,
    n37536, n37537, n37538, n37539, n37540, n37541, n37542, n37543, n37544,
    n37545, n37546, n37547, n37548, n37549, n37550, n37551, n37552, n37553,
    n37554, n37555, n37556, n37557, n37558, n37559, n37560, n37561, n37562,
    n37563, n37564, n37565, n37566, n37567, n37568, n37569, n37570, n37571,
    n37572, n37573, n37574, n37575, n37576, n37577, n37578, n37579, n37580,
    n37581, n37582, n37583, n37584, n37585, n37586, n37587, n37588, n37589,
    n37590, n37591, n37592, n37593, n37594, n37595, n37596, n37597, n37598,
    n37599, n37600, n37601, n37602, n37603, n37604, n37605, n37606, n37607,
    n37608, n37609, n37610, n37611, n37612, n37613, n37614, n37615, n37616,
    n37617, n37618, n37619, n37620, n37621, n37622, n37623, n37624, n37625,
    n37626, n37627, n37628, n37629, n37630, n37631, n37632, n37633, n37634,
    n37635, n37636, n37637, n37638, n37639, n37640, n37641, n37642, n37643,
    n37644, n37645, n37646, n37647, n37648, n37649, n37650, n37651, n37652,
    n37653, n37654, n37655, n37656, n37657, n37658, n37659, n37660, n37661,
    n37662, n37663, n37664, n37665, n37666, n37667, n37668, n37669, n37670,
    n37671, n37672, n37673, n37674, n37675, n37676, n37677, n37678, n37679,
    n37680, n37681, n37682, n37683, n37684, n37685, n37686, n37687, n37688,
    n37689, n37690, n37691, n37692, n37693, n37694, n37695, n37696, n37697,
    n37698, n37699, n37700, n37701, n37702, n37703, n37704, n37705, n37706,
    n37707, n37708, n37709, n37710, n37711, n37712, n37713, n37714, n37715,
    n37716, n37717, n37718, n37719, n37720, n37721, n37722, n37723, n37724,
    n37725, n37726, n37727, n37728, n37729, n37730, n37731, n37732, n37733,
    n37734, n37735, n37736, n37737, n37738, n37739, n37740, n37741, n37742,
    n37743, n37744, n37745, n37746, n37747, n37748, n37749, n37750, n37751,
    n37752, n37753, n37754, n37755, n37756, n37757, n37758, n37759, n37760,
    n37761, n37762, n37763, n37764, n37765, n37766, n37767, n37768, n37769,
    n37770, n37771, n37772, n37773, n37774, n37775, n37776, n37777, n37778,
    n37779, n37780, n37781, n37782, n37783, n37784, n37785, n37786, n37787,
    n37788, n37789, n37790, n37791, n37792, n37793, n37794, n37795, n37796,
    n37797, n37798, n37799, n37800, n37801, n37802, n37803, n37804, n37805,
    n37806, n37807, n37808, n37809, n37810, n37811, n37812, n37813, n37814,
    n37815, n37816, n37817, n37818, n37819, n37820, n37821, n37822, n37823,
    n37824, n37825, n37826, n37827, n37828, n37829, n37830, n37831, n37832,
    n37833, n37834, n37835, n37836, n37837, n37838, n37839, n37840, n37841,
    n37842, n37843, n37844, n37845, n37846, n37847, n37848, n37849, n37850,
    n37851, n37852, n37853, n37854, n37855, n37856, n37857, n37858, n37859,
    n37860, n37861, n37862, n37863, n37864, n37865, n37866, n37867, n37868,
    n37869, n37870, n37871, n37872, n37873, n37874, n37875, n37876, n37877,
    n37878, n37879, n37880, n37881, n37882, n37883, n37884, n37885, n37886,
    n37887, n37888, n37889, n37890, n37891, n37892, n37893, n37894, n37895,
    n37896, n37897, n37898, n37899, n37900, n37901, n37902, n37903, n37904,
    n37905, n37906, n37907, n37908, n37909, n37910, n37911, n37912, n37913,
    n37914, n37915, n37916, n37917, n37918, n37919, n37920, n37921, n37922,
    n37923, n37924, n37925, n37926, n37927, n37928, n37929, n37930, n37931,
    n37932, n37933, n37934, n37935, n37936, n37937, n37938, n37939, n37940,
    n37941, n37942, n37943, n37944, n37945, n37946, n37947, n37948, n37949,
    n37950, n37951, n37952, n37953, n37954, n37955, n37956, n37957, n37958,
    n37959, n37960, n37961, n37962, n37963, n37964, n37965, n37966, n37967,
    n37968, n37969, n37970, n37971, n37972, n37973, n37974, n37975, n37976,
    n37977, n37978, n37979, n37980, n37981, n37982, n37983, n37984, n37985,
    n37986, n37987, n37988, n37989, n37990, n37991, n37992, n37993, n37994,
    n37995, n37996, n37997, n37998, n37999, n38000, n38001, n38002, n38003,
    n38004, n38005, n38006, n38007, n38008, n38009, n38010, n38011, n38012,
    n38013, n38014, n38015, n38016, n38017, n38018, n38019, n38020, n38021,
    n38022, n38023, n38024, n38025, n38026, n38027, n38028, n38029, n38030,
    n38031, n38032, n38033, n38034, n38035, n38036, n38037, n38038, n38039,
    n38040, n38041, n38042, n38043, n38044, n38045, n38046, n38047, n38048,
    n38049, n38050, n38051, n38052, n38053, n38054, n38055, n38056, n38057,
    n38058, n38059, n38060, n38061, n38062, n38063, n38064, n38065, n38066,
    n38067, n38068, n38069, n38070, n38071, n38072, n38073, n38074, n38075,
    n38076, n38077, n38078, n38079, n38080, n38081, n38082, n38083, n38084,
    n38085, n38086, n38087, n38088, n38089, n38090, n38091, n38092, n38093,
    n38094, n38095, n38096, n38097, n38098, n38099, n38100, n38101, n38102,
    n38103, n38104, n38105, n38106, n38107, n38108, n38109, n38110, n38111,
    n38112, n38113, n38114, n38115, n38116, n38117, n38118, n38119, n38120,
    n38121, n38122, n38123, n38124, n38125, n38126, n38127, n38128, n38129,
    n38130, n38131, n38132, n38133, n38134, n38135, n38136, n38137, n38138,
    n38139, n38140, n38141, n38142, n38143, n38144, n38145, n38146, n38147,
    n38148, n38149, n38150, n38151, n38152, n38153, n38154, n38155, n38156,
    n38157, n38158, n38159, n38160, n38161, n38162, n38163, n38164, n38165,
    n38166, n38167, n38168, n38169, n38170, n38171, n38172, n38173, n38174,
    n38175, n38176, n38177, n38178, n38179, n38180, n38181, n38182, n38183,
    n38184, n38185, n38186, n38187, n38188, n38189, n38190, n38191, n38192,
    n38193, n38194, n38195, n38196, n38197, n38198, n38199, n38200, n38201,
    n38202, n38203, n38204, n38205, n38206, n38207, n38208, n38209, n38210,
    n38211, n38212, n38213, n38214, n38215, n38216, n38217, n38218, n38219,
    n38220, n38221, n38222, n38223, n38224, n38225, n38226, n38227, n38228,
    n38229, n38230, n38231, n38232, n38233, n38234, n38235, n38236, n38237,
    n38238, n38239, n38240, n38241, n38242, n38243, n38244, n38245, n38246,
    n38247, n38248, n38249, n38250, n38251, n38252, n38253, n38254, n38255,
    n38256, n38257, n38258, n38259, n38260, n38261, n38262, n38263, n38264,
    n38265, n38266, n38267, n38268, n38269, n38270, n38271, n38272, n38273,
    n38274, n38275, n38276, n38277, n38278, n38279, n38280, n38281, n38282,
    n38283, n38284, n38285, n38286, n38287, n38288, n38289, n38290, n38291,
    n38292, n38293, n38294, n38295, n38296, n38297, n38298, n38299, n38300,
    n38301, n38302, n38303, n38304, n38305, n38306, n38307, n38308, n38309,
    n38310, n38311, n38312, n38313, n38314, n38315, n38316, n38317, n38318,
    n38319, n38320, n38321, n38322, n38323, n38324, n38325, n38326, n38327,
    n38328, n38329, n38330, n38331, n38332, n38333, n38334, n38335, n38336,
    n38337, n38338, n38339, n38340, n38341, n38342, n38343, n38344, n38345,
    n38346, n38347, n38348, n38349, n38350, n38351, n38352, n38353, n38354,
    n38355, n38356, n38357, n38358, n38359, n38360, n38361, n38362, n38363,
    n38364, n38365, n38366, n38367, n38368, n38369, n38370, n38371, n38372,
    n38373, n38374, n38375, n38376, n38377, n38378, n38379, n38380, n38381,
    n38382, n38383, n38384, n38385, n38386, n38387, n38388, n38389, n38390,
    n38391, n38392, n38393, n38394, n38395, n38396, n38397, n38398, n38399,
    n38400, n38401, n38402, n38403, n38404, n38405, n38406, n38407, n38408,
    n38409, n38410, n38411, n38412, n38413, n38414, n38415, n38416, n38417,
    n38418, n38419, n38420, n38421, n38422, n38423, n38424, n38425, n38426,
    n38427, n38428, n38429, n38430, n38431, n38432, n38433, n38434, n38435,
    n38436, n38437, n38438, n38439, n38440, n38441, n38442, n38443, n38444,
    n38445, n38446, n38447, n38448, n38449, n38450, n38451, n38452, n38453,
    n38454, n38455, n38456, n38457, n38458, n38459, n38460, n38461, n38462,
    n38463, n38464, n38465, n38466, n38467, n38468, n38469, n38470, n38471,
    n38472, n38473, n38474, n38475, n38476, n38477, n38478, n38479, n38480,
    n38481, n38482, n38483, n38484, n38485, n38486, n38487, n38488, n38489,
    n38490, n38491, n38492, n38493, n38494, n38495, n38496, n38497, n38498,
    n38499, n38500, n38501, n38502, n38503, n38504, n38505, n38506, n38507,
    n38508, n38509, n38510, n38511, n38512, n38513, n38514, n38515, n38516,
    n38517, n38518, n38519, n38520, n38521, n38522, n38523, n38524, n38525,
    n38526, n38527, n38528, n38529, n38530, n38531, n38532, n38533, n38534,
    n38535, n38536, n38537, n38538, n38539, n38540, n38541, n38542, n38543,
    n38544, n38545, n38546, n38547, n38548, n38549, n38550, n38551, n38552,
    n38553, n38554, n38555, n38556, n38557, n38558, n38559, n38560, n38561,
    n38562, n38563, n38564, n38565, n38566, n38567, n38568, n38569, n38570,
    n38571, n38572, n38573, n38574, n38575, n38576, n38577, n38578, n38579,
    n38580, n38581, n38582, n38583, n38584, n38585, n38586, n38587, n38588,
    n38589, n38590, n38591, n38592, n38593, n38594, n38595, n38596, n38597,
    n38598, n38599, n38600, n38601, n38602, n38603, n38604, n38605, n38606,
    n38607, n38608, n38609, n38610, n38611, n38612, n38613, n38614, n38615,
    n38616, n38617, n38618, n38619, n38620, n38621, n38622, n38623, n38624,
    n38625, n38626, n38627, n38628, n38629, n38630, n38631, n38632, n38633,
    n38634, n38635, n38636, n38637, n38638, n38639, n38640, n38641, n38642,
    n38643, n38644, n38645, n38646, n38647, n38648, n38649, n38650, n38651,
    n38652, n38653, n38654, n38655, n38656, n38657, n38658, n38659, n38660,
    n38661, n38662, n38663, n38664, n38665, n38666, n38667, n38668, n38669,
    n38670, n38671, n38672, n38673, n38674, n38675, n38676, n38677, n38678,
    n38679, n38680, n38681, n38682, n38683, n38684, n38685, n38686, n38687,
    n38688, n38689, n38690, n38691, n38692, n38693, n38694, n38695, n38696,
    n38697, n38698, n38699, n38700, n38701, n38702, n38703, n38704, n38705,
    n38706, n38707, n38708, n38709, n38710, n38711, n38712, n38713, n38714,
    n38715, n38716, n38717, n38718, n38719, n38720, n38721, n38722, n38723,
    n38724, n38725, n38726, n38727, n38728, n38729, n38730, n38731, n38732,
    n38733, n38734, n38735, n38736, n38737, n38738, n38739, n38740, n38741,
    n38742, n38743, n38744, n38745, n38746, n38747, n38748, n38749, n38750,
    n38751, n38752, n38753, n38754, n38755, n38756, n38757, n38758, n38759,
    n38760, n38761, n38762, n38763, n38764, n38765, n38766, n38767, n38768,
    n38769, n38770, n38771, n38772, n38773, n38774, n38775, n38776, n38777,
    n38778, n38779, n38780, n38781, n38782, n38783, n38784, n38785, n38786,
    n38787, n38788, n38789, n38790, n38791, n38792, n38793, n38794, n38795,
    n38796, n38797, n38798, n38799, n38800, n38801, n38802, n38803, n38804,
    n38805, n38806, n38807, n38808, n38809, n38810, n38811, n38812, n38813,
    n38814, n38815, n38816, n38817, n38818, n38819, n38820, n38821, n38822,
    n38823, n38824, n38825, n38826, n38827, n38828, n38829, n38830, n38831,
    n38832, n38833, n38834, n38835, n38836, n38837, n38838, n38839, n38840,
    n38841, n38842, n38843, n38844, n38845, n38846, n38847, n38848, n38849,
    n38850, n38851, n38852, n38853, n38854, n38855, n38856, n38857, n38858,
    n38859, n38860, n38861, n38862, n38863, n38864, n38865, n38866, n38867,
    n38868, n38869, n38870, n38871, n38872, n38873, n38874, n38875, n38876,
    n38877, n38878, n38879, n38880, n38881, n38882, n38883, n38884, n38885,
    n38886, n38887, n38888, n38889, n38890, n38891, n38892, n38893, n38894,
    n38895, n38896, n38897, n38898, n38899, n38900, n38901, n38902, n38903,
    n38904, n38905, n38906, n38907, n38908, n38909, n38910, n38911, n38912,
    n38913, n38914, n38915, n38916, n38917, n38918, n38919, n38920, n38921,
    n38922, n38923, n38924, n38925, n38926, n38927, n38928, n38929, n38930,
    n38931, n38932, n38933, n38934, n38935, n38936, n38937, n38938, n38939,
    n38940, n38941, n38942, n38943, n38944, n38945, n38946, n38947, n38948,
    n38949, n38950, n38951, n38952, n38953, n38954, n38955, n38956, n38957,
    n38958, n38959, n38960, n38961, n38962, n38963, n38964, n38965, n38966,
    n38967, n38968, n38969, n38970, n38971, n38972, n38973, n38974, n38975,
    n38976, n38977, n38978, n38979, n38980, n38981, n38982, n38983, n38984,
    n38985, n38986, n38987, n38988, n38989, n38990, n38991, n38992, n38993,
    n38994, n38995, n38996, n38997, n38998, n38999, n39000, n39001, n39002,
    n39003, n39004, n39005, n39006, n39007, n39008, n39009, n39010, n39011,
    n39012, n39013, n39014, n39015, n39016, n39017, n39018, n39019, n39020,
    n39021, n39022, n39023, n39024, n39025, n39026, n39027, n39028, n39029,
    n39030, n39031, n39032, n39033, n39034, n39035, n39036, n39037, n39038,
    n39039, n39040, n39041, n39042, n39043, n39044, n39045, n39046, n39047,
    n39048, n39049, n39050, n39051, n39052, n39053, n39054, n39055, n39056,
    n39057, n39058, n39059, n39060, n39061, n39062, n39063, n39064, n39065,
    n39066, n39067, n39068, n39069, n39070, n39071, n39072, n39073, n39074,
    n39075, n39076, n39077, n39078, n39079, n39080, n39081, n39082, n39083,
    n39084, n39085, n39086, n39087, n39088, n39089, n39090, n39091, n39092,
    n39093, n39094, n39095, n39096, n39097, n39098, n39099, n39100, n39101,
    n39102, n39103, n39104, n39105, n39106, n39107, n39108, n39109, n39110,
    n39111, n39112, n39113, n39114, n39115, n39116, n39117, n39118, n39119,
    n39120, n39121, n39122, n39123, n39124, n39125, n39126, n39127, n39128,
    n39129, n39130, n39131, n39132, n39133, n39134, n39135, n39136, n39137,
    n39138, n39139, n39140, n39141, n39142, n39143, n39144, n39145, n39146,
    n39147, n39148, n39149, n39150, n39151, n39152, n39153, n39154, n39155,
    n39156, n39157, n39158, n39159, n39160, n39161, n39162, n39163, n39164,
    n39165, n39166, n39167, n39168, n39169, n39170, n39171, n39172, n39173,
    n39174, n39175, n39176, n39177, n39178, n39179, n39180, n39181, n39182,
    n39183, n39184, n39185, n39186, n39187, n39188, n39189, n39190, n39191,
    n39192, n39193, n39194, n39195, n39196, n39197, n39198, n39199, n39200,
    n39201, n39202, n39203, n39204, n39205, n39206, n39207, n39208, n39209,
    n39210, n39211, n39212, n39213, n39214, n39215, n39216, n39217, n39218,
    n39219, n39220, n39221, n39222, n39223, n39224, n39225, n39226, n39227,
    n39228, n39229, n39230, n39231, n39232, n39233, n39234, n39235, n39236,
    n39237, n39238, n39239, n39240, n39241, n39242, n39243, n39244, n39245,
    n39246, n39247, n39248, n39249, n39250, n39251, n39252, n39253, n39254,
    n39255, n39256, n39257, n39258, n39259, n39260, n39261, n39262, n39263,
    n39264, n39265, n39266, n39267, n39268, n39269, n39270, n39271, n39272,
    n39273, n39274, n39275, n39276, n39277, n39278, n39279, n39280, n39281,
    n39282, n39283, n39284, n39285, n39286, n39287, n39288, n39289, n39290,
    n39291, n39292, n39293, n39294, n39295, n39296, n39297, n39298, n39299,
    n39300, n39301, n39302, n39303, n39304, n39305, n39306, n39307, n39308,
    n39309, n39310, n39311, n39312, n39313, n39314, n39315, n39316, n39317,
    n39318, n39319, n39320, n39321, n39322, n39323, n39324, n39325, n39326,
    n39327, n39328, n39329, n39330, n39331, n39332, n39333, n39334, n39335,
    n39336, n39337, n39338, n39339, n39340, n39341, n39342, n39343, n39344,
    n39345, n39346, n39347, n39348, n39349, n39350, n39351, n39352, n39353,
    n39354, n39355, n39356, n39357, n39358, n39359, n39360, n39361, n39362,
    n39363, n39364, n39365, n39366, n39367, n39368, n39369, n39370, n39371,
    n39372, n39373, n39374, n39375, n39376, n39377, n39378, n39379, n39380,
    n39381, n39382, n39383, n39384, n39385, n39386, n39387, n39388, n39389,
    n39390, n39391, n39392, n39393, n39394, n39395, n39396, n39397, n39398,
    n39399, n39400, n39401, n39402, n39403, n39404, n39405, n39406, n39407,
    n39408, n39409, n39410, n39411, n39412, n39413, n39414, n39415, n39416,
    n39417, n39418, n39419, n39420, n39421, n39422, n39423, n39424, n39425,
    n39426, n39427, n39428, n39429, n39430, n39431, n39432, n39433, n39434,
    n39435, n39436, n39437, n39438, n39439, n39440, n39441, n39442, n39443,
    n39444, n39445, n39446, n39447, n39448, n39449, n39450, n39451, n39452,
    n39453, n39454, n39455, n39456, n39457, n39458, n39459, n39460, n39461,
    n39462, n39463, n39464, n39465, n39466, n39467, n39468, n39469, n39470,
    n39471, n39472, n39473, n39474, n39475, n39476, n39477, n39478, n39479,
    n39480, n39481, n39482, n39483, n39484, n39485, n39486, n39487, n39488,
    n39489, n39490, n39491, n39492, n39493, n39494, n39495, n39496, n39497,
    n39498, n39499, n39500, n39501, n39502, n39503, n39504, n39505, n39506,
    n39507, n39508, n39509, n39510, n39511, n39512, n39513, n39514, n39515,
    n39516, n39517, n39518, n39519, n39520, n39521, n39522, n39523, n39524,
    n39525, n39526, n39527, n39528, n39529, n39530, n39531, n39532, n39533,
    n39534, n39535, n39536, n39537, n39538, n39539, n39540, n39541, n39542,
    n39543, n39544, n39545, n39546, n39547, n39548, n39549, n39550, n39551,
    n39552, n39553, n39554, n39555, n39556, n39557, n39558, n39559, n39560,
    n39561, n39562, n39563, n39564, n39565, n39566, n39567, n39568, n39569,
    n39570, n39571, n39572, n39573, n39574, n39575, n39576, n39577, n39578,
    n39579, n39580, n39581, n39582, n39583, n39584, n39585, n39586, n39587,
    n39588, n39589, n39590, n39591, n39592, n39593, n39594, n39595, n39596,
    n39597, n39598, n39599, n39600, n39601, n39602, n39603, n39604, n39605,
    n39606, n39607, n39608, n39609, n39610, n39611, n39612, n39613, n39614,
    n39615, n39616, n39617, n39618, n39619, n39620, n39621, n39622, n39623,
    n39624, n39625, n39626, n39627, n39628, n39629, n39630, n39631, n39632,
    n39633, n39634, n39635, n39636, n39637, n39638, n39639, n39640, n39641,
    n39642, n39643, n39644, n39645, n39646, n39647, n39648, n39649, n39650,
    n39651, n39652, n39653, n39654, n39655, n39656, n39657, n39658, n39659,
    n39660, n39661, n39662, n39663, n39664, n39665, n39666, n39667, n39668,
    n39669, n39670, n39671, n39672, n39673, n39674, n39675, n39676, n39677,
    n39678, n39679, n39680, n39681, n39682, n39683, n39684, n39685, n39686,
    n39687, n39688, n39689, n39690, n39691, n39692, n39693, n39694, n39695,
    n39696, n39697, n39698, n39699, n39700, n39701, n39702, n39703, n39704,
    n39705, n39706, n39707, n39708, n39709, n39710, n39711, n39712, n39713,
    n39714, n39715, n39716, n39717, n39718, n39719, n39720, n39721, n39722,
    n39723, n39724, n39725, n39726, n39727, n39728, n39729, n39730, n39731,
    n39732, n39733, n39734, n39735, n39736, n39737, n39738, n39739, n39740,
    n39741, n39742, n39743, n39744, n39745, n39746, n39747, n39748, n39749,
    n39750, n39751, n39752, n39753, n39754, n39755, n39756, n39757, n39758,
    n39759, n39760, n39761, n39762, n39763, n39764, n39765, n39766, n39767,
    n39768, n39769, n39770, n39771, n39772, n39773, n39774, n39775, n39776,
    n39777, n39778, n39779, n39780, n39781, n39782, n39783, n39784, n39785,
    n39786, n39787, n39788, n39789, n39790, n39791, n39792, n39793, n39794,
    n39795, n39796, n39797, n39798, n39799, n39800, n39801, n39802, n39803,
    n39804, n39805, n39806, n39807, n39808, n39809, n39810, n39811, n39812,
    n39813, n39814, n39815, n39816, n39817, n39818, n39819, n39820, n39821,
    n39822, n39823, n39824, n39825, n39826, n39827, n39828, n39829, n39830,
    n39831, n39832, n39833, n39834, n39835, n39836, n39837, n39838, n39839,
    n39840, n39841, n39842, n39843, n39844, n39845, n39846, n39847, n39848,
    n39849, n39850, n39851, n39852, n39853, n39854, n39855, n39856, n39857,
    n39858, n39859, n39860, n39861, n39862, n39863, n39864, n39865, n39866,
    n39867, n39868, n39869, n39870, n39871, n39872, n39873, n39874, n39875,
    n39876, n39877, n39878, n39879, n39880, n39881, n39882, n39883, n39884,
    n39885, n39886, n39887, n39888, n39889, n39890, n39891, n39892, n39893,
    n39894, n39895, n39896, n39897, n39898, n39899, n39900, n39901, n39902,
    n39903, n39904, n39905, n39906, n39907, n39908, n39909, n39910, n39911,
    n39912, n39913, n39914, n39915, n39916, n39917, n39918, n39919, n39920,
    n39921, n39922, n39923, n39924, n39925, n39926, n39927, n39928, n39929,
    n39930, n39931, n39932, n39933, n39934, n39935, n39936, n39937, n39938,
    n39939, n39940, n39941, n39942, n39943, n39944, n39945, n39946, n39947,
    n39948, n39949, n39950, n39951, n39952, n39953, n39954, n39955, n39956,
    n39957, n39958, n39959, n39960, n39961, n39962, n39963, n39964, n39965,
    n39966, n39967, n39968, n39969, n39970, n39971, n39972, n39973, n39974,
    n39975, n39976, n39977, n39978, n39979, n39980, n39981, n39982, n39983,
    n39984, n39985, n39986, n39987, n39988, n39989, n39990, n39991, n39992,
    n39993, n39994, n39995, n39996, n39997, n39998, n39999, n40000, n40001,
    n40002, n40003, n40004, n40005, n40006, n40007, n40008, n40009, n40010,
    n40011, n40012, n40013, n40014, n40015, n40016, n40017, n40018, n40019,
    n40020, n40021, n40022, n40023, n40024, n40025, n40026, n40027, n40028,
    n40029, n40030, n40031, n40032, n40033, n40034, n40035, n40036, n40037,
    n40038, n40039, n40040, n40041, n40042, n40043, n40044, n40045, n40046,
    n40047, n40048, n40049, n40050, n40051, n40052, n40053, n40054, n40055,
    n40056, n40057, n40058, n40059, n40060, n40061, n40062, n40063, n40064,
    n40065, n40066, n40067, n40068, n40069, n40070, n40071, n40072, n40073,
    n40074, n40075, n40076, n40077, n40078, n40079, n40080, n40081, n40082,
    n40083, n40084, n40085, n40086, n40087, n40088, n40089, n40090, n40091,
    n40092, n40093, n40094, n40095, n40096, n40097, n40098, n40099, n40100,
    n40101, n40102, n40103, n40104, n40105, n40106, n40107, n40108, n40109,
    n40110, n40111, n40112, n40113, n40114, n40115, n40116, n40117, n40118,
    n40119, n40120, n40121, n40122, n40123, n40124, n40125, n40126, n40127,
    n40128, n40129, n40130, n40131, n40132, n40133, n40134, n40135, n40136,
    n40137, n40138, n40139, n40140, n40141, n40142, n40143, n40144, n40145,
    n40146, n40147, n40148, n40149, n40150, n40151, n40152, n40153, n40154,
    n40155, n40156, n40157, n40158, n40159, n40160, n40161, n40162, n40163,
    n40164, n40165, n40166, n40167, n40168, n40169, n40170, n40171, n40172,
    n40173, n40174, n40175, n40176, n40177, n40178, n40179, n40180, n40181,
    n40182, n40183, n40184, n40185, n40186, n40187, n40188, n40189, n40190,
    n40191, n40192, n40193, n40194, n40195, n40196, n40197, n40198, n40199,
    n40200, n40201, n40202, n40203, n40204, n40205, n40206, n40207, n40208,
    n40209, n40210, n40211, n40212, n40213, n40214, n40215, n40216, n40217,
    n40218, n40219, n40220, n40221, n40222, n40223, n40224, n40225, n40226,
    n40227, n40228, n40229, n40230, n40231, n40232, n40233, n40234, n40235,
    n40236, n40237, n40238, n40239, n40240, n40241, n40242, n40243, n40244,
    n40245, n40246, n40247, n40248, n40249, n40250, n40251, n40252, n40253,
    n40254, n40255, n40256, n40257, n40258, n40259, n40260, n40261, n40262,
    n40263, n40264, n40265, n40266, n40267, n40268, n40269, n40270, n40271,
    n40272, n40273, n40274, n40275, n40276, n40277, n40278, n40279, n40280,
    n40281, n40282, n40283, n40284, n40285, n40286, n40287, n40288, n40289,
    n40290, n40291, n40292, n40293, n40294, n40295, n40296, n40297, n40298,
    n40299, n40300, n40301, n40302, n40303, n40304, n40305, n40306, n40307,
    n40308, n40309, n40310, n40311, n40312, n40313, n40314, n40315, n40316,
    n40317, n40318, n40319, n40320, n40321, n40322, n40323, n40324, n40325,
    n40326, n40327, n40328, n40329, n40330, n40331, n40332, n40333, n40334,
    n40335, n40336, n40337, n40338, n40339, n40340, n40341, n40342, n40343,
    n40344, n40345, n40346, n40347, n40348, n40349, n40350, n40351, n40352,
    n40353, n40354, n40355, n40356, n40357, n40358, n40359, n40360, n40361,
    n40362, n40363, n40364, n40365, n40366, n40367, n40368, n40369, n40370,
    n40371, n40372, n40373, n40374, n40375, n40376, n40377, n40378, n40379,
    n40380, n40381, n40382, n40383, n40384, n40385, n40386, n40387, n40388,
    n40389, n40390, n40391, n40392, n40393, n40394, n40395, n40396, n40397,
    n40398, n40399, n40400, n40401, n40402, n40403, n40404, n40405, n40406,
    n40407, n40408, n40409, n40410, n40411, n40412, n40413, n40414, n40415,
    n40416, n40417, n40418, n40419, n40420, n40421, n40422, n40423, n40424,
    n40425, n40426, n40427, n40428, n40429, n40430, n40431, n40432, n40433,
    n40434, n40435, n40436, n40437, n40438, n40439, n40440, n40441, n40442,
    n40443, n40444, n40445, n40446, n40447, n40448, n40449, n40450, n40451,
    n40452, n40453, n40454, n40455, n40456, n40457, n40458, n40459, n40460,
    n40461, n40462, n40463, n40464, n40465, n40466, n40467, n40468, n40469,
    n40470, n40471, n40472, n40473, n40474, n40475, n40476, n40477, n40478,
    n40479, n40480, n40481, n40482, n40483, n40484, n40485, n40486, n40487,
    n40488, n40489, n40490, n40491, n40492, n40493, n40494, n40495, n40496,
    n40497, n40498, n40499, n40500, n40501, n40502, n40503, n40504, n40505,
    n40506, n40507, n40508, n40509, n40510, n40511, n40512, n40513, n40514,
    n40515, n40516, n40517, n40518, n40519, n40520, n40521, n40522, n40523,
    n40524, n40525, n40526, n40527, n40528, n40529, n40530, n40531, n40532,
    n40533, n40534, n40535, n40536, n40537, n40538, n40539, n40540, n40541,
    n40542, n40543, n40544, n40545, n40546, n40547, n40548, n40549, n40550,
    n40551, n40552, n40553, n40554, n40555, n40556, n40557, n40558, n40559,
    n40560, n40561, n40562, n40563, n40564, n40565, n40566, n40567, n40568,
    n40569, n40570, n40571, n40572, n40573, n40574, n40575, n40576, n40577,
    n40578, n40579, n40580, n40581, n40582, n40583, n40584, n40585, n40586,
    n40587, n40588, n40589, n40590, n40591, n40592, n40593, n40594, n40595,
    n40596, n40597, n40598, n40599, n40600, n40601, n40602, n40603, n40604,
    n40605, n40606, n40607, n40608, n40609, n40610, n40611, n40612, n40613,
    n40614, n40615, n40616, n40617, n40618, n40619, n40620, n40621, n40622,
    n40623, n40624, n40625, n40626, n40627, n40628, n40629, n40630, n40631,
    n40632, n40633, n40634, n40635, n40636, n40637, n40638, n40639, n40640,
    n40641, n40642, n40643, n40644, n40645, n40646, n40647, n40648, n40649,
    n40650, n40651, n40652, n40653, n40654, n40655, n40656, n40657, n40658,
    n40659, n40660, n40661, n40662, n40663, n40664, n40665, n40666, n40667,
    n40668, n40669, n40670, n40671, n40672, n40673, n40674, n40675, n40676,
    n40677, n40678, n40679, n40680, n40681, n40682, n40683, n40684, n40685,
    n40686, n40687, n40688, n40689, n40690, n40691, n40692, n40693, n40694,
    n40695, n40696, n40697, n40698, n40699, n40700, n40701, n40702, n40703,
    n40704, n40705, n40706, n40707, n40708, n40709, n40710, n40711, n40712,
    n40713, n40714, n40715, n40716, n40717, n40718, n40719, n40720, n40721,
    n40722, n40723, n40724, n40725, n40726, n40727, n40728, n40729, n40730,
    n40731, n40732, n40733, n40734, n40735, n40736, n40737, n40738, n40739,
    n40740, n40741, n40742, n40743, n40744, n40745, n40746, n40747, n40748,
    n40749, n40750, n40751, n40752, n40753, n40754, n40755, n40756, n40757,
    n40758, n40759, n40760, n40761, n40762, n40763, n40764, n40765, n40766,
    n40767, n40768, n40769, n40770, n40771, n40772, n40773, n40774, n40775,
    n40776, n40777, n40778, n40779, n40780, n40781, n40782, n40783, n40784,
    n40785, n40786, n40787, n40788, n40789, n40790, n40791, n40792, n40793,
    n40794, n40795, n40796, n40797, n40798, n40799, n40800, n40801, n40802,
    n40803, n40804, n40805, n40806, n40807, n40808, n40809, n40810, n40811,
    n40812, n40813, n40814, n40815, n40816, n40817, n40818, n40819, n40820,
    n40821, n40822, n40823, n40824, n40825, n40826, n40827, n40828, n40829,
    n40830, n40831, n40832, n40833, n40834, n40835, n40836, n40837, n40838,
    n40839, n40840, n40841, n40842, n40843, n40844, n40845, n40846, n40847,
    n40848, n40849, n40850, n40851, n40852, n40853, n40854, n40855, n40856,
    n40857, n40858, n40859, n40860, n40861, n40862, n40863, n40864, n40865,
    n40866, n40867, n40868, n40869, n40870, n40871, n40872, n40873, n40874,
    n40875, n40876, n40877, n40878, n40879, n40880, n40881, n40882, n40883,
    n40884, n40885, n40886, n40887, n40888, n40889, n40890, n40891, n40892,
    n40893, n40894, n40895, n40896, n40897, n40898, n40899, n40900, n40901,
    n40902, n40903, n40904, n40905, n40906, n40907, n40908, n40909, n40910,
    n40911, n40912, n40913, n40914, n40915, n40916, n40917, n40918, n40919,
    n40920, n40921, n40922, n40923, n40924, n40925, n40926, n40927, n40928,
    n40929, n40930, n40931, n40932, n40933, n40934, n40935, n40936, n40937,
    n40938, n40939, n40940, n40941, n40942, n40943, n40944, n40945, n40946,
    n40947, n40948, n40949, n40950, n40951, n40952, n40953, n40954, n40955,
    n40956, n40957, n40958, n40959, n40960, n40961, n40962, n40963, n40964,
    n40965, n40966, n40967, n40968, n40969, n40970, n40971, n40972, n40973,
    n40974, n40975, n40976, n40977, n40978, n40979, n40980, n40981, n40982,
    n40983, n40984, n40985, n40986, n40987, n40988, n40989, n40990, n40991,
    n40992, n40993, n40994, n40995, n40996, n40997, n40998, n40999, n41000,
    n41001, n41002, n41003, n41004, n41005, n41006, n41007, n41008, n41009,
    n41010, n41011, n41012, n41013, n41014, n41015, n41016, n41017, n41018,
    n41019, n41020, n41021, n41022, n41023, n41024, n41025, n41026, n41027,
    n41028, n41029, n41030, n41031, n41032, n41033, n41034, n41035, n41036,
    n41037, n41038, n41039, n41040, n41041, n41042, n41043, n41044, n41045,
    n41046, n41047, n41048, n41049, n41050, n41051, n41052, n41053, n41054,
    n41055, n41056, n41057, n41058, n41059, n41060, n41061, n41062, n41063,
    n41064, n41065, n41066, n41067, n41068, n41069, n41070, n41071, n41072,
    n41073, n41074, n41075, n41076, n41077, n41078, n41079, n41080, n41081,
    n41082, n41083, n41084, n41085, n41086, n41087, n41088, n41089, n41090,
    n41091, n41092, n41093, n41094, n41095, n41096, n41097, n41098, n41099,
    n41100, n41101, n41102, n41103, n41104, n41105, n41106, n41107, n41108,
    n41109, n41110, n41111, n41112, n41113, n41114, n41115, n41116, n41117,
    n41118, n41119, n41120, n41121, n41122, n41123, n41124, n41125, n41126,
    n41127, n41128, n41129, n41130, n41131, n41132, n41133, n41134, n41135,
    n41136, n41137, n41138, n41139, n41140, n41141, n41142, n41143, n41144,
    n41145, n41146, n41147, n41148, n41149, n41150, n41151, n41152, n41153,
    n41154, n41155, n41156, n41157, n41158, n41159, n41160, n41161, n41162,
    n41163, n41164, n41165, n41166, n41167, n41168, n41169, n41170, n41171,
    n41172, n41173, n41174, n41175, n41176, n41177, n41178, n41179, n41180,
    n41181, n41182, n41183, n41184, n41185, n41186, n41187, n41188, n41189,
    n41190, n41191, n41192, n41193, n41194, n41195, n41196, n41197, n41198,
    n41199, n41200, n41201, n41202, n41203, n41204, n41205, n41206, n41207,
    n41208, n41209, n41210, n41211, n41212, n41213, n41214, n41215, n41216,
    n41217, n41218, n41219, n41220, n41221, n41222, n41223, n41224, n41225,
    n41226, n41227, n41228, n41229, n41230, n41231, n41232, n41233, n41234,
    n41235, n41236, n41237, n41238, n41239, n41240, n41241, n41242, n41243,
    n41244, n41245, n41246, n41247, n41248, n41249, n41250, n41251, n41252,
    n41253, n41254, n41255, n41256, n41257, n41258, n41259, n41260, n41261,
    n41262, n41263, n41264, n41265, n41266, n41267, n41268, n41269, n41270,
    n41271, n41272, n41273, n41274, n41275, n41276, n41277, n41278, n41279,
    n41280, n41281, n41282, n41283, n41284, n41285, n41286, n41287, n41288,
    n41289, n41290, n41291, n41292, n41293, n41294, n41295, n41296, n41297,
    n41298, n41299, n41300, n41301, n41302, n41303, n41304, n41305, n41306,
    n41307, n41308, n41309, n41310, n41311, n41312, n41313, n41314, n41315,
    n41316, n41317, n41318, n41319, n41320, n41321, n41322, n41323, n41324,
    n41325, n41326, n41327, n41328, n41329, n41330, n41331, n41332, n41333,
    n41334, n41335, n41336, n41337, n41338, n41339, n41340, n41341, n41342,
    n41343, n41344, n41345, n41346, n41347, n41348, n41349, n41350, n41351,
    n41352, n41353, n41354, n41355, n41356, n41357, n41358, n41359, n41360,
    n41361, n41362, n41363, n41364, n41365, n41366, n41367, n41368, n41369,
    n41370, n41371, n41372, n41373, n41374, n41375, n41376, n41377, n41378,
    n41379, n41380, n41381, n41382, n41383, n41384, n41385, n41386, n41387,
    n41388, n41389, n41390, n41391, n41392, n41393, n41394, n41395, n41396,
    n41397, n41398, n41399, n41400, n41401, n41402, n41403, n41404, n41405,
    n41406, n41407, n41408, n41409, n41410, n41411, n41412, n41413, n41414,
    n41415, n41416, n41417, n41418, n41419, n41420, n41421, n41422, n41423,
    n41424, n41425, n41426, n41427, n41428, n41429, n41430, n41431, n41432,
    n41433, n41434, n41435, n41436, n41437, n41438, n41439, n41440, n41441,
    n41442, n41443, n41444, n41445, n41446, n41447, n41448, n41449, n41450,
    n41451, n41452, n41453, n41454, n41455, n41456, n41457, n41458, n41459,
    n41460, n41461, n41462, n41463, n41464, n41465, n41466, n41467, n41468,
    n41469, n41470, n41471, n41472, n41473, n41474, n41475, n41476, n41477,
    n41478, n41479, n41480, n41481, n41482, n41483, n41484, n41485, n41486,
    n41487, n41488, n41489, n41490, n41491, n41492, n41493, n41494, n41495,
    n41496, n41497, n41498, n41499, n41500, n41501, n41502, n41503, n41504,
    n41505, n41506, n41507, n41508, n41509, n41510, n41511, n41512, n41513,
    n41514, n41515, n41516, n41517, n41518, n41519, n41520, n41521, n41522,
    n41523, n41524, n41525, n41526, n41527, n41528, n41529, n41530, n41531,
    n41532, n41533, n41534, n41535, n41536, n41537, n41538, n41539, n41540,
    n41541, n41542, n41543, n41544, n41545, n41546, n41547, n41548, n41549,
    n41550, n41551, n41552, n41553, n41554, n41555, n41556, n41557, n41558,
    n41559, n41560, n41561, n41562, n41563, n41564, n41565, n41566, n41567,
    n41568, n41569, n41570, n41571, n41572, n41573, n41574, n41575, n41576,
    n41577, n41578, n41579, n41580, n41581, n41582, n41583, n41584, n41585,
    n41586, n41587, n41588, n41589, n41590, n41591, n41592, n41593, n41594,
    n41595, n41596, n41597, n41598, n41599, n41600, n41601, n41602, n41603,
    n41604, n41605, n41606, n41607, n41608, n41609, n41610, n41611, n41612,
    n41613, n41614, n41615, n41616, n41617, n41618, n41619, n41620, n41621,
    n41622, n41623, n41624, n41625, n41626, n41627, n41628, n41629, n41630,
    n41631, n41632, n41633, n41634, n41635, n41636, n41637, n41638, n41639,
    n41640, n41641, n41642, n41643, n41644, n41645, n41646, n41647, n41648,
    n41649, n41650, n41651, n41652, n41653, n41654, n41655, n41656, n41657,
    n41658, n41659, n41660, n41661, n41662, n41663, n41664, n41665, n41666,
    n41667, n41668, n41669, n41670, n41671, n41672, n41673, n41674, n41675,
    n41676, n41677, n41678, n41679, n41680, n41681, n41682, n41683, n41684,
    n41685, n41686, n41687, n41688, n41689, n41690, n41691, n41692, n41693,
    n41694, n41695, n41696, n41697, n41698, n41699, n41700, n41701, n41702,
    n41703, n41704, n41705, n41706, n41707, n41708, n41709, n41710, n41711,
    n41712, n41713, n41714, n41715, n41716, n41717, n41718, n41719, n41720,
    n41721, n41722, n41723, n41724, n41725, n41726, n41727, n41728, n41729,
    n41730, n41731, n41732, n41733, n41734, n41735, n41736, n41737, n41738,
    n41739, n41740, n41741, n41742, n41743, n41744, n41745, n41746, n41747,
    n41748, n41749, n41750, n41751, n41752, n41753, n41754, n41755, n41756,
    n41757, n41758, n41759, n41760, n41761, n41762, n41763, n41764, n41765,
    n41766, n41767, n41768, n41769, n41770, n41771, n41772, n41773, n41774,
    n41775, n41776, n41777, n41778, n41779, n41780, n41781, n41782, n41783,
    n41784, n41785, n41786, n41787, n41788, n41789, n41790, n41791, n41792,
    n41793, n41794, n41795, n41796, n41797, n41798, n41799, n41800, n41801,
    n41802, n41803, n41804, n41805, n41806, n41807, n41808, n41809, n41810,
    n41811, n41812, n41813, n41814, n41815, n41816, n41817, n41818, n41819,
    n41820, n41821, n41822, n41823, n41824, n41825, n41826, n41827, n41828,
    n41829, n41830, n41831, n41832, n41833, n41834, n41835, n41836, n41837,
    n41838, n41839, n41840, n41841, n41842, n41843, n41844, n41845, n41846,
    n41847, n41848, n41849, n41850, n41851, n41852, n41853, n41854, n41855,
    n41856, n41857, n41858, n41859, n41860, n41861, n41862, n41863, n41864,
    n41865, n41866, n41867, n41868, n41869, n41870, n41871, n41872, n41873,
    n41874, n41875, n41876, n41877, n41878, n41879, n41880, n41881, n41882,
    n41883, n41884, n41885, n41886, n41887, n41888, n41889, n41890, n41891,
    n41892, n41893, n41894, n41895, n41896, n41897, n41898, n41899, n41900,
    n41901, n41902, n41903, n41904, n41905, n41906, n41907, n41908, n41909,
    n41910, n41911, n41912, n41913, n41914, n41915, n41916, n41917, n41918,
    n41919, n41920, n41921, n41922, n41923, n41924, n41925, n41926, n41927,
    n41928, n41929, n41930, n41931, n41932, n41933, n41934, n41935, n41936,
    n41937, n41938, n41939, n41940, n41941, n41942, n41943, n41944, n41945,
    n41946, n41947, n41948, n41949, n41950, n41951, n41952, n41953, n41954,
    n41955, n41956, n41957, n41958, n41959, n41960, n41961, n41962, n41963,
    n41964, n41965, n41966, n41967, n41968, n41969, n41970, n41971, n41972,
    n41973, n41974, n41975, n41976, n41977, n41978, n41979, n41980, n41981,
    n41982, n41983, n41984, n41985, n41986, n41987, n41988, n41989, n41990,
    n41991, n41992, n41993, n41994, n41995, n41996, n41997, n41998, n41999,
    n42000, n42001, n42002, n42003, n42004, n42005, n42006, n42007, n42008,
    n42009, n42010, n42011, n42012, n42013, n42014, n42015, n42016, n42017,
    n42018, n42019, n42020, n42021, n42022, n42023, n42024, n42025, n42026,
    n42027, n42028, n42029, n42030, n42031, n42032, n42033, n42034, n42035,
    n42036, n42037, n42038, n42039, n42040, n42041, n42042, n42043, n42044,
    n42045, n42046, n42047, n42048, n42049, n42050, n42051, n42052, n42053,
    n42054, n42055, n42056, n42057, n42058, n42059, n42060, n42061, n42062,
    n42063, n42064, n42065, n42066, n42067, n42068, n42069, n42070, n42071,
    n42072, n42073, n42074, n42075, n42076, n42077, n42078, n42079, n42080,
    n42081, n42082, n42083, n42084, n42085, n42086, n42087, n42088, n42089,
    n42090, n42091, n42092, n42093, n42094, n42095, n42096, n42097, n42098,
    n42099, n42100, n42101, n42102, n42103, n42104, n42105, n42106, n42107,
    n42108, n42109, n42110, n42111, n42112, n42113, n42114, n42115, n42116,
    n42117, n42118, n42119, n42120, n42121, n42122, n42123, n42124, n42125,
    n42126, n42127, n42128, n42129, n42130, n42131, n42132, n42133, n42134,
    n42135, n42136, n42137, n42138, n42139, n42140, n42141, n42142, n42143,
    n42144, n42145, n42146, n42147, n42148, n42149, n42150, n42151, n42152,
    n42153, n42154, n42155, n42156, n42157, n42158, n42159, n42160, n42161,
    n42162, n42163, n42164, n42165, n42166, n42167, n42168, n42169, n42170,
    n42171, n42172, n42173, n42174, n42175, n42176, n42177, n42178, n42179,
    n42180, n42181, n42182, n42183, n42184, n42185, n42186, n42187, n42188,
    n42189, n42190, n42191, n42192, n42193, n42194, n42195, n42196, n42197,
    n42198, n42199, n42200, n42201, n42202, n42203, n42204, n42205, n42206,
    n42207, n42208, n42209, n42210, n42211, n42212, n42213, n42214, n42215,
    n42216, n42217, n42218, n42219, n42220, n42221, n42222, n42223, n42224,
    n42225, n42226, n42227, n42228, n42229, n42230, n42231, n42232, n42233,
    n42234, n42235, n42236, n42237, n42238, n42239, n42240, n42241, n42242,
    n42243, n42244, n42245, n42246, n42247, n42248, n42249, n42250, n42251,
    n42252, n42253, n42254, n42255, n42256, n42257, n42258, n42259, n42260,
    n42261, n42262, n42263, n42264, n42265, n42266, n42267, n42268, n42269,
    n42270, n42271, n42272, n42273, n42274, n42275, n42276, n42277, n42278,
    n42279, n42280, n42281, n42282, n42283, n42284, n42285, n42286, n42287,
    n42288, n42289, n42290, n42291, n42292, n42293, n42294, n42295, n42296,
    n42297, n42298, n42299, n42300, n42301, n42302, n42303, n42304, n42305,
    n42306, n42307, n42308, n42309, n42310, n42311, n42312, n42313, n42314,
    n42315, n42316, n42317, n42318, n42319, n42320, n42321, n42322, n42323,
    n42324, n42325, n42326, n42327, n42328, n42329, n42330, n42331, n42332,
    n42333, n42334, n42335, n42336, n42337, n42338, n42339, n42340, n42341,
    n42342, n42343, n42344, n42345, n42346, n42347, n42348, n42349, n42350,
    n42351, n42352, n42353, n42354, n42355, n42356, n42357, n42358, n42359,
    n42360, n42361, n42362, n42363, n42364, n42365, n42366, n42367, n42368,
    n42369, n42370, n42371, n42372, n42373, n42374, n42375, n42376, n42377,
    n42378, n42379, n42380, n42381, n42382, n42383, n42384, n42385, n42386,
    n42387, n42388, n42389, n42390, n42391, n42392, n42393, n42394, n42395,
    n42396, n42397, n42398, n42399, n42400, n42401, n42402, n42403, n42404,
    n42405, n42406, n42407, n42408, n42409, n42410, n42411, n42412, n42413,
    n42414, n42415, n42416, n42417, n42418, n42419, n42420, n42421, n42422,
    n42423, n42424, n42425, n42426, n42427, n42428, n42429, n42430, n42431,
    n42432, n42433, n42434, n42435, n42436, n42437, n42438, n42439, n42440,
    n42441, n42442, n42443, n42444, n42445, n42446, n42447, n42448, n42449,
    n42450, n42451, n42452, n42453, n42454, n42455, n42456, n42457, n42458,
    n42459, n42460, n42461, n42462, n42463, n42464, n42465, n42466, n42467,
    n42468, n42469, n42470, n42471, n42472, n42473, n42474, n42475, n42476,
    n42477, n42478, n42479, n42480, n42481, n42482, n42483, n42484, n42485,
    n42486, n42487, n42488, n42489, n42490, n42491, n42492, n42493, n42494,
    n42495, n42496, n42497, n42498, n42499, n42500, n42501, n42502, n42503,
    n42504, n42505, n42506, n42507, n42508, n42509, n42510, n42511, n42512,
    n42513, n42514, n42515, n42516, n42517, n42518, n42519, n42520, n42521,
    n42522, n42523, n42524, n42525, n42526, n42527, n42528, n42529, n42530,
    n42531, n42532, n42533, n42534, n42535, n42536, n42537, n42538, n42539,
    n42540, n42541, n42542, n42543, n42544, n42545, n42546, n42547, n42548,
    n42549, n42550, n42551, n42552, n42553, n42554, n42555, n42556, n42557,
    n42558, n42559, n42560, n42561, n42562, n42563, n42564, n42565, n42566,
    n42567, n42568, n42569, n42570, n42571, n42572, n42573, n42574, n42575,
    n42576, n42577, n42578, n42579, n42580, n42581, n42582, n42583, n42584,
    n42585, n42586, n42587, n42588, n42589, n42590, n42591, n42592, n42593,
    n42594, n42595, n42596, n42597, n42598, n42599, n42600, n42601, n42602,
    n42603, n42604, n42605, n42606, n42607, n42608, n42609, n42610, n42611,
    n42612, n42613, n42614, n42615, n42616, n42617, n42618, n42619, n42620,
    n42621, n42622, n42623, n42624, n42625, n42626, n42627, n42628, n42629,
    n42630, n42631, n42632, n42633, n42634, n42635, n42636, n42637, n42638,
    n42639, n42640, n42641, n42642, n42643, n42644, n42645, n42646, n42647,
    n42648, n42649, n42650, n42651, n42652, n42653, n42654, n42655, n42656,
    n42657, n42658, n42659, n42660, n42661, n42662, n42663, n42664, n42665,
    n42666, n42667, n42668, n42669, n42670, n42671, n42672, n42673, n42674,
    n42675, n42676, n42677, n42678, n42679, n42680, n42681, n42682, n42683,
    n42684, n42685, n42686, n42687, n42688, n42689, n42690, n42691, n42692,
    n42693, n42694, n42695, n42696, n42697, n42698, n42699, n42700, n42701,
    n42702, n42703, n42704, n42705, n42706, n42707, n42708, n42709, n42710,
    n42711, n42712, n42713, n42714, n42715, n42716, n42717, n42718, n42719,
    n42720, n42721, n42722, n42723, n42724, n42725, n42726, n42727, n42728,
    n42729, n42730, n42731, n42732, n42733, n42734, n42735, n42736, n42737,
    n42738, n42739, n42740, n42741, n42742, n42743, n42744, n42745, n42746,
    n42747, n42748, n42749, n42750, n42751, n42752, n42753, n42754, n42755,
    n42756, n42757, n42758, n42759, n42760, n42761, n42762, n42763, n42764,
    n42765, n42766, n42767, n42768, n42769, n42770, n42771, n42772, n42773,
    n42774, n42775, n42776, n42777, n42778, n42779, n42780, n42781, n42782,
    n42783, n42784, n42785, n42786, n42787, n42788, n42789, n42790, n42791,
    n42792, n42793, n42794, n42795, n42796, n42797, n42798, n42799, n42800,
    n42801, n42802, n42803, n42804, n42805, n42806, n42807, n42808, n42809,
    n42810, n42811, n42812, n42813, n42814, n42815, n42816, n42817, n42818,
    n42819, n42820, n42821, n42822, n42823, n42824, n42825, n42826, n42827,
    n42828, n42829, n42830, n42831, n42832, n42833, n42834, n42835, n42836,
    n42837, n42838, n42839, n42840, n42841, n42842, n42843, n42844, n42845,
    n42846, n42847, n42848, n42849, n42850, n42851, n42852, n42853, n42854,
    n42855, n42856, n42857, n42858, n42859, n42860, n42861, n42862, n42863,
    n42864, n42865, n42866, n42867, n42868, n42869, n42870, n42871, n42872,
    n42873, n42874, n42875, n42876, n42877, n42878, n42879, n42880, n42881,
    n42882, n42883, n42884, n42885, n42886, n42887, n42888, n42889, n42890,
    n42891, n42892, n42893, n42894, n42895, n42896, n42897, n42898, n42899,
    n42900, n42901, n42902, n42903, n42904, n42905, n42906, n42907, n42908,
    n42909, n42910, n42911, n42912, n42913, n42914, n42915, n42916, n42917,
    n42918, n42919, n42920, n42921, n42922, n42923, n42924, n42925, n42926,
    n42927, n42928, n42929, n42930, n42931, n42932, n42933, n42934, n42935,
    n42936, n42937, n42938, n42939, n42940, n42941, n42942, n42943, n42944,
    n42945, n42946, n42947, n42948, n42949, n42950, n42951, n42952, n42953,
    n42954, n42955, n42956, n42957, n42958, n42959, n42960, n42961, n42962,
    n42963, n42964, n42965, n42966, n42967, n42968, n42969, n42970, n42971,
    n42972, n42973, n42974, n42975, n42976, n42977, n42978, n42979, n42980,
    n42981, n42982, n42983, n42984, n42985, n42986, n42987, n42988, n42989,
    n42990, n42991, n42992, n42993, n42994, n42995, n42996, n42997, n42998,
    n42999, n43000, n43001, n43002, n43003, n43004, n43005, n43006, n43007,
    n43008, n43009, n43010, n43011, n43012, n43013, n43014, n43015, n43016,
    n43017, n43018, n43019, n43020, n43021, n43022, n43023, n43024, n43025,
    n43026, n43027, n43028, n43029, n43030, n43031, n43032, n43033, n43034,
    n43035, n43036, n43037, n43038, n43039, n43040, n43041, n43042, n43043,
    n43044, n43045, n43046, n43047, n43048, n43049, n43050, n43051, n43052,
    n43053, n43054, n43055, n43056, n43057, n43058, n43059, n43060, n43061,
    n43062, n43063, n43064, n43065, n43066, n43067, n43068, n43069, n43070,
    n43071, n43072, n43073, n43074, n43075, n43076, n43077, n43078, n43079,
    n43080, n43081, n43082, n43083, n43084, n43085, n43086, n43087, n43088,
    n43089, n43090, n43091, n43092, n43093, n43094, n43095, n43096, n43097,
    n43098, n43099, n43100, n43101, n43102, n43103, n43104, n43105, n43106,
    n43107, n43108, n43109, n43110, n43111, n43112, n43113, n43114, n43115,
    n43116, n43117, n43118, n43119, n43120, n43121, n43122, n43123, n43124,
    n43125, n43126, n43127, n43128, n43129, n43130, n43131, n43132, n43133,
    n43134, n43135, n43136, n43137, n43138, n43139, n43140, n43141, n43142,
    n43143, n43144, n43145, n43146, n43147, n43148, n43149, n43150, n43151,
    n43152, n43153, n43154, n43155, n43156, n43157, n43158, n43159, n43160,
    n43161, n43162, n43163, n43164, n43165, n43166, n43167, n43168, n43169,
    n43170, n43171, n43172, n43173, n43174, n43175, n43176, n43177, n43178,
    n43179, n43180, n43181, n43182, n43183, n43184, n43185, n43186, n43187,
    n43188, n43189, n43190, n43191, n43192, n43193, n43194, n43195, n43196,
    n43197, n43198, n43199, n43200, n43201, n43202, n43203, n43204, n43205,
    n43206, n43207, n43208, n43209, n43210, n43211, n43212, n43213, n43214,
    n43215, n43216, n43217, n43218, n43219, n43220, n43221, n43222, n43223,
    n43224, n43225, n43226, n43227, n43228, n43229, n43230, n43231, n43232,
    n43233, n43234, n43235, n43236, n43237, n43238, n43239, n43240, n43241,
    n43242, n43243, n43244, n43245, n43246, n43247, n43248, n43249, n43250,
    n43251, n43252, n43253, n43254, n43255, n43256, n43257, n43258, n43259,
    n43260, n43261, n43262, n43263, n43264, n43265, n43266, n43267, n43268,
    n43269, n43270, n43271, n43272, n43273, n43274, n43275, n43276, n43277,
    n43278, n43279, n43280, n43281, n43282, n43283, n43284, n43285, n43286,
    n43287, n43288, n43289, n43290, n43291, n43292, n43293, n43294, n43295,
    n43296, n43297, n43298, n43299, n43300, n43301, n43302, n43303, n43304,
    n43305, n43306, n43307, n43308, n43309, n43310, n43311, n43312, n43313,
    n43314, n43315, n43316, n43317, n43318, n43319, n43320, n43321, n43322,
    n43323, n43324, n43325, n43326, n43327, n43328, n43329, n43330, n43331,
    n43332, n43333, n43334, n43335, n43336, n43337, n43338, n43339, n43340,
    n43341, n43342, n43343, n43344, n43345, n43346, n43347, n43348, n43349,
    n43350, n43351, n43352, n43353, n43354, n43355, n43356, n43357, n43358,
    n43359, n43360, n43361, n43362, n43363, n43364, n43365, n43366, n43367,
    n43368, n43369, n43370, n43371, n43372, n43373, n43374, n43375, n43376,
    n43377, n43378, n43379, n43380, n43381, n43382, n43383, n43384, n43385,
    n43386, n43387, n43388, n43389, n43390, n43391, n43392, n43393, n43394,
    n43395, n43396, n43397, n43398, n43399, n43400, n43401, n43402, n43403,
    n43404, n43405, n43406, n43407, n43408, n43409, n43410, n43411, n43412,
    n43413, n43414, n43415, n43416, n43417, n43418, n43419, n43420, n43421,
    n43422, n43423, n43424, n43425, n43426, n43427, n43428, n43429, n43430,
    n43431, n43432, n43433, n43434, n43435, n43436, n43437, n43438, n43439,
    n43440, n43441, n43442, n43443, n43444, n43445, n43446, n43447, n43448,
    n43449, n43450, n43451, n43452, n43453, n43454, n43455, n43456, n43457,
    n43458, n43459, n43460, n43461, n43462, n43463, n43464, n43465, n43466,
    n43467, n43468, n43469, n43470, n43471, n43472, n43473, n43474, n43475,
    n43476, n43477, n43478, n43479, n43480, n43481, n43482, n43483, n43484,
    n43485, n43486, n43487, n43488, n43489, n43490, n43491, n43492, n43493,
    n43494, n43495, n43496, n43497, n43498, n43499, n43500, n43501, n43502,
    n43503, n43504, n43505, n43506, n43507, n43508, n43509, n43510, n43511,
    n43512, n43513, n43514, n43515, n43516, n43517, n43518, n43519, n43520,
    n43521, n43522, n43523, n43524, n43525, n43526, n43527, n43528, n43529,
    n43530, n43531, n43532, n43533, n43534, n43535, n43536, n43537, n43538,
    n43539, n43540, n43541, n43542, n43543, n43544, n43545, n43546, n43547,
    n43548, n43549, n43550, n43551, n43552, n43553, n43554, n43555, n43556,
    n43557, n43558, n43559, n43560, n43561, n43562, n43563, n43564, n43565,
    n43566, n43567, n43568, n43569, n43570, n43571, n43572, n43573, n43574,
    n43575, n43576, n43577, n43578, n43579, n43580, n43581, n43582, n43583,
    n43584, n43585, n43586, n43587, n43588, n43589, n43590, n43591, n43592,
    n43593, n43594, n43595, n43596, n43597, n43598, n43599, n43600, n43601,
    n43602, n43603, n43604, n43605, n43606, n43607, n43608, n43609, n43610,
    n43611, n43612, n43613, n43614, n43615, n43616, n43617, n43618, n43619,
    n43620, n43621, n43622, n43623, n43624, n43625, n43626, n43627, n43628,
    n43629, n43630, n43631, n43632, n43633, n43634, n43635, n43636, n43637,
    n43638, n43639, n43640, n43641, n43642, n43643, n43644, n43645, n43646,
    n43647, n43648, n43649, n43650, n43651, n43652, n43653, n43654, n43655,
    n43656, n43657, n43658, n43659, n43660, n43661, n43662, n43663, n43664,
    n43665, n43666, n43667, n43668, n43669, n43670, n43671, n43672, n43673,
    n43674, n43675, n43676, n43677, n43678, n43679, n43680, n43681, n43682,
    n43683, n43684, n43685, n43686, n43687, n43688, n43689, n43690, n43691,
    n43692, n43693, n43694, n43695, n43696, n43697, n43698, n43699, n43700,
    n43701, n43702, n43703, n43704, n43705, n43706, n43707, n43708, n43709,
    n43710, n43711, n43712, n43713, n43714, n43715, n43716, n43717, n43718,
    n43719, n43720, n43721, n43722, n43723, n43724, n43725, n43726, n43727,
    n43728, n43729, n43730, n43731, n43732, n43733, n43734, n43735, n43736,
    n43737, n43738, n43739, n43740, n43741, n43742, n43743, n43744, n43745,
    n43746, n43747, n43748, n43749, n43750, n43751, n43752, n43753, n43754,
    n43755, n43756, n43757, n43758, n43759, n43760, n43761, n43762, n43763,
    n43764, n43765, n43766, n43767, n43768, n43769, n43770, n43771, n43772,
    n43773, n43774, n43775, n43776, n43777, n43778, n43779, n43780, n43781,
    n43782, n43783, n43784, n43785, n43786, n43787, n43788, n43789, n43790,
    n43791, n43792, n43793, n43794, n43795, n43796, n43797, n43798, n43799,
    n43800, n43801, n43802, n43803, n43804, n43805, n43806, n43807, n43808,
    n43809, n43810, n43811, n43812, n43813, n43814, n43815, n43816, n43817,
    n43818, n43819, n43820, n43821, n43822, n43823, n43824, n43825, n43826,
    n43827, n43828, n43829, n43830, n43831, n43832, n43833, n43834, n43835,
    n43836, n43837, n43838, n43839, n43840, n43841, n43842, n43843, n43844,
    n43845, n43846, n43847, n43848, n43849, n43850, n43851, n43852, n43853,
    n43854, n43855, n43856, n43857, n43858, n43859, n43860, n43861, n43862,
    n43863, n43864, n43865, n43866, n43867, n43868, n43869, n43870, n43871,
    n43872, n43873, n43874, n43875, n43876, n43877, n43878, n43879, n43880,
    n43881, n43882, n43883, n43884, n43885, n43886, n43887, n43888, n43889,
    n43890, n43891, n43892, n43893, n43894, n43895, n43896, n43897, n43898,
    n43899, n43900, n43901, n43902, n43903, n43904, n43905, n43906, n43907,
    n43908, n43909, n43910, n43911, n43912, n43913, n43914, n43915, n43916,
    n43917, n43918, n43919, n43920, n43921, n43922, n43923, n43924, n43925,
    n43926, n43927, n43928, n43929, n43930, n43931, n43932, n43933, n43934,
    n43935, n43936, n43937, n43938, n43939, n43940, n43941, n43942, n43943,
    n43944, n43945, n43946, n43947, n43948, n43949, n43950, n43951, n43952,
    n43953, n43954, n43955, n43956, n43957, n43958, n43959, n43960, n43961,
    n43962, n43963, n43964, n43965, n43966, n43967, n43968, n43969, n43970,
    n43971, n43972, n43973, n43974, n43975, n43976, n43977, n43978, n43979,
    n43980, n43981, n43982, n43983, n43984, n43985, n43986, n43987, n43988,
    n43989, n43990, n43991, n43992, n43993, n43994, n43995, n43996, n43997,
    n43998, n43999, n44000, n44001, n44002, n44003, n44004, n44005, n44006,
    n44007, n44008, n44009, n44010, n44011, n44012, n44013, n44014, n44015,
    n44016, n44017, n44018, n44019, n44020, n44021, n44022, n44023, n44024,
    n44025, n44026, n44027, n44028, n44029, n44030, n44031, n44032, n44033,
    n44034, n44035, n44036, n44037, n44038, n44039, n44040, n44041, n44042,
    n44043, n44044, n44045, n44046, n44047, n44048, n44049, n44050, n44051,
    n44052, n44053, n44054, n44055, n44056, n44057, n44058, n44059, n44060,
    n44061, n44062, n44063, n44064, n44065, n44066, n44067, n44068, n44069,
    n44070, n44071, n44072, n44073, n44074, n44075, n44076, n44077, n44078,
    n44079, n44080, n44081, n44082, n44083, n44084, n44085, n44086, n44087,
    n44088, n44089, n44090, n44091, n44092, n44093, n44094, n44095, n44096,
    n44097, n44098, n44099, n44100, n44101, n44102, n44103, n44104, n44105,
    n44106, n44107, n44108, n44109, n44110, n44111, n44112, n44113, n44114,
    n44115, n44116, n44117, n44118, n44119, n44120, n44121, n44122, n44123,
    n44124, n44125, n44126, n44127, n44128, n44129, n44130, n44131, n44132,
    n44133, n44134, n44135, n44136, n44137, n44138, n44139, n44140, n44141,
    n44142, n44143, n44144, n44145, n44146, n44147, n44148, n44149, n44150,
    n44151, n44152, n44153, n44154, n44155, n44156, n44157, n44158, n44159,
    n44160, n44161, n44162, n44163, n44164, n44165, n44166, n44167, n44168,
    n44169, n44170, n44171, n44172, n44173, n44174, n44175, n44176, n44177,
    n44178, n44179, n44180, n44181, n44182, n44183, n44184, n44185, n44186,
    n44187, n44188, n44189, n44190, n44191, n44192, n44193, n44194, n44195,
    n44196, n44197, n44198, n44199, n44200, n44201, n44202, n44203, n44204,
    n44205, n44206, n44207, n44208, n44209, n44210, n44211, n44212, n44213,
    n44214, n44215, n44216, n44217, n44218, n44219, n44220, n44221, n44222,
    n44223, n44224, n44225, n44226, n44227, n44228, n44229, n44230, n44231,
    n44232, n44233, n44234, n44235, n44236, n44237, n44238, n44239, n44240,
    n44241, n44242, n44243, n44244, n44245, n44246, n44247, n44248, n44249,
    n44250, n44251, n44252, n44253, n44254, n44255, n44256, n44257, n44258,
    n44259, n44260, n44261, n44262, n44263, n44264, n44265, n44266, n44267,
    n44268, n44269, n44270, n44271, n44272, n44273, n44274, n44275, n44276,
    n44277, n44278, n44279, n44280, n44281, n44282, n44283, n44284, n44285,
    n44286, n44287, n44288, n44289, n44290, n44291, n44292, n44293, n44294,
    n44295, n44296, n44297, n44298, n44299, n44300, n44301, n44302, n44303,
    n44304, n44305, n44306, n44307, n44308, n44309, n44310, n44311, n44312,
    n44313, n44314, n44315, n44316, n44317, n44318, n44319, n44320, n44321,
    n44322, n44323, n44324, n44325, n44326, n44327, n44328, n44329, n44330,
    n44331, n44332, n44333, n44334, n44335, n44336, n44337, n44338, n44339,
    n44340, n44341, n44342, n44343, n44344, n44345, n44346, n44347, n44348,
    n44349, n44350, n44351, n44352, n44353, n44354, n44355, n44356, n44357,
    n44358, n44359, n44360, n44361, n44362, n44363, n44364, n44365, n44366,
    n44367, n44368, n44369, n44370, n44371, n44372, n44373, n44374, n44375,
    n44376, n44377, n44378, n44379, n44380, n44381, n44382, n44383, n44384,
    n44385, n44386, n44387, n44388, n44389, n44390, n44391, n44392, n44393,
    n44394, n44395, n44396, n44397, n44398, n44399, n44400, n44401, n44402,
    n44403, n44404, n44405, n44406, n44407, n44408, n44409, n44410, n44411,
    n44412, n44413, n44414, n44415, n44416, n44417, n44418, n44419, n44420,
    n44421, n44422, n44423, n44424, n44425, n44426, n44427, n44428, n44429,
    n44430, n44431, n44432, n44433, n44434, n44435, n44436, n44437, n44438,
    n44439, n44440, n44441, n44442, n44443, n44444, n44445, n44446, n44447,
    n44448, n44449, n44450, n44451, n44452, n44453, n44454, n44455, n44456,
    n44457, n44458, n44459, n44460, n44461, n44462, n44463, n44464, n44465,
    n44466, n44467, n44468, n44469, n44470, n44471, n44472, n44473, n44474,
    n44475, n44476, n44477, n44478, n44479, n44480, n44481, n44482, n44483,
    n44484, n44485, n44486, n44487, n44488, n44489, n44490, n44491, n44492,
    n44493, n44494, n44495, n44496, n44497, n44498, n44499, n44500, n44501,
    n44502, n44503, n44504, n44505, n44506, n44507, n44508, n44509, n44510,
    n44511, n44512, n44513, n44514, n44515, n44516, n44517, n44518, n44519,
    n44520, n44521, n44522, n44523, n44524, n44525, n44526, n44527, n44528,
    n44529, n44530, n44531, n44532, n44533, n44534, n44535, n44536, n44537,
    n44538, n44539, n44540, n44541, n44542, n44543, n44544, n44545, n44546,
    n44547, n44548, n44549, n44550, n44551, n44552, n44553, n44554, n44555,
    n44556, n44557, n44558, n44559, n44560, n44561, n44562, n44563, n44564,
    n44565, n44566, n44567, n44568, n44569, n44570, n44571, n44572, n44573,
    n44574, n44575, n44576, n44577, n44578, n44579, n44580, n44581, n44582,
    n44583, n44584, n44585, n44586, n44587, n44588, n44589, n44590, n44591,
    n44592, n44593, n44594, n44595, n44596, n44597, n44598, n44599, n44600,
    n44601, n44602, n44603, n44604, n44605, n44606, n44607, n44608, n44609,
    n44610, n44611, n44612, n44613, n44614, n44615, n44616, n44617, n44618,
    n44619, n44620, n44621, n44622, n44623, n44624, n44625, n44626, n44627,
    n44628, n44629, n44630, n44631, n44632, n44633, n44634, n44635, n44636,
    n44637, n44638, n44639, n44640, n44641, n44642, n44643, n44644, n44645,
    n44646, n44647, n44648, n44649, n44650, n44651, n44652, n44653, n44654,
    n44655, n44656, n44657, n44658, n44659, n44660, n44661, n44662, n44663,
    n44664, n44665, n44666, n44667, n44668, n44669, n44670, n44671, n44672,
    n44673, n44674, n44675, n44676, n44677, n44678, n44679, n44680, n44681,
    n44682, n44683, n44684, n44685, n44686, n44687, n44688, n44689, n44690,
    n44691, n44692, n44693, n44694, n44695, n44696, n44697, n44698, n44699,
    n44700, n44701, n44702, n44703, n44704, n44705, n44706, n44707, n44708,
    n44709, n44710, n44711, n44712, n44713, n44714, n44715, n44716, n44717,
    n44718, n44719, n44720, n44721, n44722, n44723, n44724, n44725, n44726,
    n44727, n44728, n44729, n44730, n44731, n44732, n44733, n44734, n44735,
    n44736, n44737, n44738, n44739, n44740, n44741, n44742, n44743, n44744,
    n44745, n44746, n44747, n44748, n44749, n44750, n44751, n44752, n44753,
    n44754, n44755, n44756, n44757, n44758, n44759, n44760, n44761, n44762,
    n44763, n44764, n44765, n44766, n44767, n44768, n44769, n44770, n44771,
    n44772, n44773, n44774, n44775, n44776, n44777, n44778, n44779, n44780,
    n44781, n44782, n44783, n44784, n44785, n44786, n44787, n44788, n44789,
    n44790, n44791, n44792, n44793, n44794, n44795, n44796, n44797, n44798,
    n44799, n44800, n44801, n44802, n44803, n44804, n44805, n44806, n44807,
    n44808, n44809, n44810, n44811, n44812, n44813, n44814, n44815, n44816,
    n44817, n44818, n44819, n44820, n44821, n44822, n44823, n44824, n44825,
    n44826, n44827, n44828, n44829, n44830, n44831, n44832, n44833, n44834,
    n44835, n44836, n44837, n44838, n44839, n44840, n44841, n44842, n44843,
    n44844, n44845, n44846, n44847, n44848, n44849, n44850, n44851, n44852,
    n44853, n44854, n44855, n44856, n44857, n44858, n44859, n44860, n44861,
    n44862, n44863, n44864, n44865, n44866, n44867, n44868, n44869, n44870,
    n44871, n44872, n44873, n44874, n44875, n44876, n44877, n44878, n44879,
    n44880, n44881, n44882, n44883, n44884, n44885, n44886, n44887, n44888,
    n44889, n44890, n44891, n44892, n44893, n44894, n44895, n44896, n44897,
    n44898, n44899, n44900, n44901, n44902, n44903, n44904, n44905, n44906,
    n44907, n44908, n44909, n44910, n44911, n44912, n44913, n44914, n44915,
    n44916, n44917, n44918, n44919, n44920, n44921, n44922, n44923, n44924,
    n44925, n44926, n44927, n44928, n44929, n44930, n44931, n44932, n44933,
    n44934, n44935, n44936, n44937, n44938, n44939, n44940, n44941, n44942,
    n44943, n44944, n44945, n44946, n44947, n44948, n44949, n44950, n44951,
    n44952, n44953, n44954, n44955, n44956, n44957, n44958, n44959, n44960,
    n44961, n44962, n44963, n44964, n44965, n44966, n44967, n44968, n44969,
    n44970, n44971, n44972, n44973, n44974, n44975, n44976, n44977, n44978,
    n44979, n44980, n44981, n44982, n44983, n44984, n44985, n44986, n44987,
    n44988, n44989, n44990, n44991, n44992, n44993, n44994, n44995, n44996,
    n44997, n44998, n44999, n45000, n45001, n45002, n45003, n45004, n45005,
    n45006, n45007, n45008, n45009, n45010, n45011, n45012, n45013, n45014,
    n45015, n45016, n45017, n45018, n45019, n45020, n45021, n45022, n45023,
    n45024, n45025, n45026, n45027, n45028, n45029, n45030, n45031, n45032,
    n45033, n45034, n45035, n45036, n45037, n45038, n45039, n45040, n45041,
    n45042, n45043, n45044, n45045, n45046, n45047, n45048, n45049, n45050,
    n45051, n45052, n45053, n45054, n45055, n45056, n45057, n45058, n45059,
    n45060, n45061, n45062, n45063, n45064, n45065, n45066, n45067, n45068,
    n45069, n45070, n45071, n45072, n45073, n45074, n45075, n45076, n45077,
    n45078, n45079, n45080, n45081, n45082, n45083, n45084, n45085, n45086,
    n45087, n45088, n45089, n45090, n45091, n45092, n45093, n45094, n45095,
    n45096, n45097, n45098, n45099, n45100, n45101, n45102, n45103, n45104,
    n45105, n45106, n45107, n45108, n45109, n45110, n45111, n45112, n45113,
    n45114, n45115, n45116, n45117, n45118, n45119, n45120, n45121, n45122,
    n45123, n45124, n45125, n45126, n45127, n45128, n45129, n45130, n45131,
    n45132, n45133, n45134, n45135, n45136, n45137, n45138, n45139, n45140,
    n45141, n45142, n45143, n45144, n45145, n45146, n45147, n45148, n45149,
    n45150, n45151, n45152, n45153, n45154, n45155, n45156, n45157, n45158,
    n45159, n45160, n45161, n45162, n45163, n45164, n45165, n45166, n45167,
    n45168, n45169, n45170, n45171, n45172, n45173, n45174, n45175, n45176,
    n45177, n45178, n45179, n45180, n45181, n45182, n45183, n45184, n45185,
    n45186, n45187, n45188, n45189, n45190, n45191, n45192, n45193, n45194,
    n45195, n45196, n45197, n45198, n45199, n45200, n45201, n45202, n45203,
    n45204, n45205, n45206, n45207, n45208, n45209, n45210, n45211, n45212,
    n45213, n45214, n45215, n45216, n45217, n45218, n45219, n45220, n45221,
    n45222, n45223, n45224, n45225, n45226, n45227, n45228, n45229, n45230,
    n45231, n45232, n45233, n45234, n45235, n45236, n45237, n45238, n45239,
    n45240, n45241, n45242, n45243, n45244, n45245, n45246, n45247, n45248,
    n45249, n45250, n45251, n45252, n45253, n45254, n45255, n45256, n45257,
    n45258, n45259, n45260, n45261, n45262, n45263, n45264, n45265, n45266,
    n45267, n45268, n45269, n45270, n45271, n45272, n45273, n45274, n45275,
    n45276, n45277, n45278, n45279, n45280, n45281, n45282, n45283, n45284,
    n45285, n45286, n45287, n45288, n45289, n45290, n45291, n45292, n45293,
    n45294, n45295, n45296, n45297, n45298, n45299, n45300, n45301, n45302,
    n45303, n45304, n45305, n45306, n45307, n45308, n45309, n45310, n45311,
    n45312, n45313, n45314, n45315, n45316, n45317, n45318, n45319, n45320,
    n45321, n45322, n45323, n45324, n45325, n45326, n45327, n45328, n45329,
    n45330, n45331, n45332, n45333, n45334, n45335, n45336, n45337, n45338,
    n45339, n45340, n45341, n45342, n45343, n45344, n45345, n45346, n45347,
    n45348, n45349, n45350, n45351, n45352, n45353, n45354, n45355, n45356,
    n45357, n45358, n45359, n45360, n45361, n45362, n45363, n45364, n45365,
    n45366, n45367, n45368, n45369, n45370, n45371, n45372, n45373, n45374,
    n45375, n45376, n45377, n45378, n45379, n45380, n45381, n45382, n45383,
    n45384, n45385, n45386, n45387, n45388, n45389, n45390, n45391, n45392,
    n45393, n45394, n45395, n45396, n45397, n45398, n45399, n45400, n45401,
    n45402, n45403, n45404, n45405, n45406, n45407, n45408, n45409, n45410,
    n45411, n45412, n45413, n45414, n45415, n45416, n45417, n45418, n45419,
    n45420, n45421, n45422, n45423, n45424, n45425, n45426, n45427, n45428,
    n45429, n45430, n45431, n45432, n45433, n45434, n45435, n45436, n45437,
    n45438, n45439, n45440, n45441, n45442, n45443, n45444, n45445, n45446,
    n45447, n45448, n45449, n45450, n45451, n45452, n45453, n45454, n45455,
    n45456, n45457, n45458, n45459, n45460, n45461, n45462, n45463, n45464,
    n45465, n45466, n45467, n45468, n45469, n45470, n45471, n45472, n45473,
    n45474, n45475, n45476, n45477, n45478, n45479, n45480, n45481, n45482,
    n45483, n45484, n45485, n45486, n45487, n45488, n45489, n45490, n45491,
    n45492, n45493, n45494, n45495, n45496, n45497, n45498, n45499, n45500,
    n45501, n45502, n45503, n45504, n45505, n45506, n45507, n45508, n45509,
    n45510, n45511, n45512, n45513, n45514, n45515, n45516, n45517, n45518,
    n45519, n45520, n45521, n45522, n45523, n45524, n45525, n45526, n45527,
    n45528, n45529, n45530, n45531, n45532, n45533, n45534, n45535, n45536,
    n45537, n45538, n45539, n45540, n45541, n45542, n45543, n45544, n45545,
    n45546, n45547, n45548, n45549, n45550, n45551, n45552, n45553, n45554,
    n45555, n45556, n45557, n45558, n45559, n45560, n45561, n45562, n45563,
    n45564, n45565, n45566, n45567, n45568, n45569, n45570, n45571, n45572,
    n45573, n45574, n45575, n45576, n45577, n45578, n45579, n45580, n45581,
    n45582, n45583, n45584, n45585, n45586, n45587, n45588, n45589, n45590,
    n45591, n45592, n45593, n45594, n45595, n45596, n45597, n45598, n45599,
    n45600, n45601, n45602, n45603, n45604, n45605, n45606, n45607, n45608,
    n45609, n45610, n45611, n45612, n45613, n45614, n45615, n45616, n45617,
    n45618, n45619, n45620, n45621, n45622, n45623, n45624, n45625, n45626,
    n45627, n45628, n45629, n45630, n45631, n45632, n45633, n45634, n45635,
    n45636, n45637, n45638, n45639, n45640, n45641, n45642, n45643, n45644,
    n45645, n45646, n45647, n45648, n45649, n45650, n45651, n45652, n45653,
    n45654, n45655, n45656, n45657, n45658, n45659, n45660, n45661, n45662,
    n45663, n45664, n45665, n45666, n45667, n45668, n45669, n45670, n45671,
    n45672, n45673, n45674, n45675, n45676, n45677, n45678, n45679, n45680,
    n45681, n45682, n45683, n45684, n45685, n45686, n45687, n45688, n45689,
    n45690, n45691, n45692, n45693, n45694, n45695, n45696, n45697, n45698,
    n45699, n45700, n45701, n45702, n45703, n45704, n45705, n45706, n45707,
    n45708, n45709, n45710, n45711, n45712, n45713, n45714, n45715, n45716,
    n45717, n45718, n45719, n45720, n45721, n45722, n45723, n45724, n45725,
    n45726, n45727, n45728, n45729, n45730, n45731, n45732, n45733, n45734,
    n45735, n45736, n45737, n45738, n45739, n45740, n45741, n45742, n45743,
    n45744, n45745, n45746, n45747, n45748, n45749, n45750, n45751, n45752,
    n45753, n45754, n45755, n45756, n45757, n45758, n45759, n45760, n45761,
    n45762, n45763, n45764, n45765, n45766, n45767, n45768, n45769, n45770,
    n45771, n45772, n45773, n45774, n45775, n45776, n45777, n45778, n45779,
    n45780, n45781, n45782, n45783, n45784, n45785, n45786, n45787, n45788,
    n45789, n45790, n45791, n45792, n45793, n45794, n45795, n45796, n45797,
    n45798, n45799, n45800, n45801, n45802, n45803, n45804, n45805, n45806,
    n45807, n45808, n45809, n45810, n45811, n45812, n45813, n45814, n45815,
    n45816, n45817, n45818, n45819, n45820, n45821, n45822, n45823, n45824,
    n45825, n45826, n45827, n45828, n45829, n45830, n45831, n45832, n45833,
    n45834, n45835, n45836, n45837, n45838, n45839, n45840, n45841, n45842,
    n45843, n45844, n45845, n45846, n45847, n45848, n45849, n45850, n45851,
    n45852, n45853, n45854, n45855, n45856, n45857, n45858, n45859, n45860,
    n45861, n45862, n45863, n45864, n45865, n45866, n45867, n45868, n45869,
    n45870, n45871, n45872, n45873, n45874, n45875, n45876, n45877, n45878,
    n45879, n45880, n45881, n45882, n45883, n45884, n45885, n45886, n45887,
    n45888, n45889, n45890, n45891, n45892, n45893, n45894, n45895, n45896,
    n45897, n45898, n45899, n45900, n45901, n45902, n45903, n45904, n45905,
    n45906, n45907, n45908, n45909, n45910, n45911, n45912, n45913, n45914,
    n45915, n45916, n45917, n45918, n45919, n45920, n45921, n45922, n45923,
    n45924, n45925, n45926, n45927, n45928, n45929, n45930, n45931, n45932,
    n45933, n45934, n45935, n45936, n45937, n45938, n45939, n45940, n45941,
    n45942, n45943, n45944, n45945, n45946, n45947, n45948, n45949, n45950,
    n45951, n45952, n45953, n45954, n45955, n45956, n45957, n45958, n45959,
    n45960, n45961, n45962, n45963, n45964, n45965, n45966, n45967, n45968,
    n45969, n45970, n45971, n45972, n45973, n45974, n45975, n45976, n45977,
    n45978, n45979, n45980, n45981, n45982, n45983, n45984, n45985, n45986,
    n45987, n45988, n45989, n45990, n45991, n45992, n45993, n45994, n45995,
    n45996, n45997, n45998, n45999, n46000, n46001, n46002, n46003, n46004,
    n46005, n46006, n46007, n46008, n46009, n46010, n46011, n46012, n46013,
    n46014, n46015, n46016, n46017, n46018, n46019, n46020, n46021, n46022,
    n46023, n46024, n46025, n46026, n46027, n46028, n46029, n46030, n46031,
    n46032, n46033, n46034, n46035, n46036, n46037, n46038, n46039, n46040,
    n46041, n46042, n46043, n46044, n46045, n46046, n46047, n46048, n46049,
    n46050, n46051, n46052, n46053, n46054, n46055, n46056, n46057, n46058,
    n46059, n46060, n46061, n46062, n46063, n46064, n46065, n46066, n46067,
    n46068, n46069, n46070, n46071, n46072, n46073, n46074, n46075, n46076,
    n46077, n46078, n46079, n46080, n46081, n46082, n46083, n46084, n46085,
    n46086, n46087, n46088, n46089, n46090, n46091, n46092, n46093, n46094,
    n46095, n46096, n46097, n46098, n46099, n46100, n46101, n46102, n46103,
    n46104, n46105, n46106, n46107, n46108, n46109, n46110, n46111, n46112,
    n46113, n46114, n46115, n46116, n46117, n46118, n46119, n46120, n46121,
    n46122, n46123, n46124, n46125, n46126, n46127, n46128, n46129, n46130,
    n46131, n46132, n46133, n46134, n46135, n46136, n46137, n46138, n46139,
    n46140, n46141, n46142, n46143, n46144, n46145, n46146, n46147, n46148,
    n46149, n46150, n46151, n46152, n46153, n46154, n46155, n46156, n46157,
    n46158, n46159, n46160, n46161, n46162, n46163, n46164, n46165, n46166,
    n46167, n46168, n46169, n46170, n46171, n46172, n46173, n46174, n46175,
    n46176, n46177, n46178, n46179, n46180, n46181, n46182, n46183, n46184,
    n46185, n46186, n46187, n46188, n46189, n46190, n46191, n46192, n46193,
    n46194, n46195, n46196, n46197, n46198, n46199, n46200, n46201, n46202,
    n46203, n46204, n46205, n46206, n46207, n46208, n46209, n46210, n46211,
    n46212, n46213, n46214, n46215, n46216, n46217, n46218, n46219, n46220,
    n46221, n46222, n46223, n46224, n46225, n46226, n46227, n46228, n46229,
    n46230, n46231, n46232, n46233, n46234, n46235, n46236, n46237, n46238,
    n46239, n46240, n46241, n46242, n46243, n46244, n46245, n46246, n46247,
    n46248, n46249, n46250, n46251, n46252, n46253, n46254, n46255, n46256,
    n46257, n46258, n46259, n46260, n46261, n46262, n46263, n46264, n46265,
    n46266, n46267, n46268, n46269, n46270, n46271, n46272, n46273, n46274,
    n46275, n46276, n46277, n46278, n46279, n46280, n46281, n46282, n46283,
    n46284, n46285, n46286, n46287, n46288, n46289, n46290, n46291, n46292,
    n46293, n46294, n46295, n46296, n46297, n46298, n46299, n46300, n46301,
    n46302, n46303, n46304, n46305, n46306, n46307, n46308, n46309, n46310,
    n46311, n46312, n46313, n46314, n46315, n46316, n46317, n46318, n46319,
    n46320, n46321, n46322, n46323, n46324, n46325, n46326, n46327, n46328,
    n46329, n46330, n46331, n46332, n46333, n46334, n46335, n46336, n46337,
    n46338, n46339, n46340, n46341, n46342, n46343, n46344, n46345, n46346,
    n46347, n46348, n46349, n46350, n46351, n46352, n46353, n46354, n46355,
    n46356, n46357, n46358, n46359, n46360, n46361, n46362, n46363, n46364,
    n46365, n46366, n46367, n46368, n46369, n46370, n46371, n46372, n46373,
    n46374, n46375, n46376, n46377, n46378, n46379, n46380, n46381, n46382,
    n46383, n46384, n46385, n46386, n46387, n46388, n46389, n46390, n46391,
    n46392, n46393, n46394, n46395, n46396, n46397, n46398, n46399, n46400,
    n46401, n46402, n46403, n46404, n46405, n46406, n46407, n46408, n46409,
    n46410, n46411, n46412, n46413, n46414, n46415, n46416, n46417, n46418,
    n46419, n46420, n46421, n46422, n46423, n46424, n46425, n46426, n46427,
    n46428, n46429, n46430, n46431, n46432, n46433, n46434, n46435, n46436,
    n46437, n46438, n46439, n46440, n46441, n46442, n46443, n46444, n46445,
    n46446, n46447, n46448, n46449, n46450, n46451, n46452, n46453, n46454,
    n46455, n46456, n46457, n46458, n46459, n46460, n46461, n46462, n46463,
    n46464, n46465, n46466, n46467, n46468, n46469, n46470, n46471, n46472,
    n46473, n46474, n46475, n46476, n46477, n46478, n46479, n46480, n46481,
    n46482, n46483, n46484, n46485, n46486, n46487, n46488, n46489, n46490,
    n46491, n46492, n46493, n46494, n46495, n46496, n46497, n46498, n46499,
    n46500, n46501, n46502, n46503, n46504, n46505, n46506, n46507, n46508,
    n46509, n46510, n46511, n46512, n46513, n46514, n46515, n46516, n46517,
    n46518, n46519, n46520, n46521, n46522, n46523, n46524, n46525, n46526,
    n46527, n46528, n46529, n46530, n46531, n46532, n46533, n46534, n46535,
    n46536, n46537, n46538, n46539, n46540, n46541, n46542, n46543, n46544,
    n46545, n46546, n46547, n46548, n46549, n46550, n46551, n46552, n46553,
    n46554, n46555, n46556, n46557, n46558, n46559, n46560, n46561, n46562,
    n46563, n46564, n46565, n46566, n46567, n46568, n46569, n46570, n46571,
    n46572, n46573, n46574, n46575, n46576, n46577, n46578, n46579, n46580,
    n46581, n46582, n46583, n46584, n46585, n46586, n46587, n46588, n46589,
    n46590, n46591, n46592, n46593, n46594, n46595, n46596, n46597, n46598,
    n46599, n46600, n46601, n46602, n46603, n46604, n46605, n46606, n46607,
    n46608, n46609, n46610, n46611, n46612, n46613, n46614, n46615, n46616,
    n46617, n46618, n46619, n46620, n46621, n46622, n46623, n46624, n46625,
    n46626, n46627, n46628, n46629, n46630, n46631, n46632, n46633, n46634,
    n46635, n46636, n46637, n46638, n46639, n46640, n46641, n46642, n46643,
    n46644, n46645, n46646, n46647, n46648, n46649, n46650, n46651, n46652,
    n46653, n46654, n46655, n46656, n46657, n46658, n46659, n46660, n46661,
    n46662, n46663, n46664, n46665, n46666, n46667, n46668, n46669, n46670,
    n46671, n46672, n46673, n46674, n46675, n46676, n46677, n46678, n46679,
    n46680, n46681, n46682, n46683, n46684, n46685, n46686, n46687, n46688,
    n46689, n46690, n46691, n46692, n46693, n46694, n46695, n46696, n46697,
    n46698, n46699, n46700, n46701, n46702, n46703, n46704, n46705, n46706,
    n46707, n46708, n46709, n46710, n46711, n46712, n46713, n46714, n46715,
    n46716, n46717, n46718, n46719, n46720, n46721, n46722, n46723, n46724,
    n46725, n46726, n46727, n46728, n46729, n46730, n46731, n46732, n46733,
    n46734, n46735, n46736, n46737, n46738, n46739, n46740, n46741, n46742,
    n46743, n46744, n46745, n46746, n46747, n46748, n46749, n46750, n46751,
    n46752, n46753, n46754, n46755, n46756, n46757, n46758, n46759, n46760,
    n46761, n46762, n46763, n46764, n46765, n46766, n46767, n46768, n46769,
    n46770, n46771, n46772, n46773, n46774, n46775, n46776, n46777, n46778,
    n46779, n46780, n46781, n46782, n46783, n46784, n46785, n46786, n46787,
    n46788, n46789, n46790, n46791, n46792, n46793, n46794, n46795, n46796,
    n46797, n46798, n46799, n46800, n46801, n46802, n46803, n46804, n46805,
    n46806, n46807, n46808, n46809, n46810, n46811, n46812, n46813, n46814,
    n46815, n46816, n46817, n46818, n46819, n46820, n46821, n46822, n46823,
    n46824, n46825, n46826, n46827, n46828, n46829, n46830, n46831, n46832,
    n46833, n46834, n46835, n46836, n46837, n46838, n46839, n46840, n46841,
    n46842, n46843, n46844, n46845, n46846, n46847, n46848, n46849, n46850,
    n46851, n46852, n46853, n46854, n46855, n46856, n46857, n46858, n46859,
    n46860, n46861, n46862, n46863, n46864, n46865, n46866, n46867, n46868,
    n46869, n46870, n46871, n46872, n46873, n46874, n46875, n46876, n46877,
    n46878, n46879, n46880, n46881, n46882, n46883, n46884, n46885, n46886,
    n46887, n46888, n46889, n46890, n46891, n46892, n46893, n46894, n46895,
    n46896, n46897, n46898, n46899, n46900, n46901, n46902, n46903, n46904,
    n46905, n46906, n46907, n46908, n46909, n46910, n46911, n46912, n46913,
    n46914, n46915, n46916, n46917, n46918, n46919, n46920, n46921, n46922,
    n46923, n46924, n46925, n46926, n46927, n46928, n46929, n46930, n46931,
    n46932, n46933, n46934, n46935, n46936, n46937, n46938, n46939, n46940,
    n46941, n46942, n46943, n46944, n46945, n46946, n46947, n46948, n46949,
    n46950, n46951, n46952, n46953, n46954, n46955, n46956, n46957, n46958,
    n46959, n46960, n46961, n46962, n46963, n46964, n46965, n46966, n46967,
    n46968, n46969, n46970, n46971, n46972, n46973, n46974, n46975, n46976,
    n46977, n46978, n46979, n46980, n46981, n46982, n46983, n46984, n46985,
    n46986, n46987, n46988, n46989, n46990, n46991, n46992, n46993, n46994,
    n46995, n46996, n46997, n46998, n46999, n47000, n47001, n47002, n47003,
    n47004, n47005, n47006, n47007, n47008, n47009, n47010, n47011, n47012,
    n47013, n47014, n47015, n47016, n47017, n47018, n47019, n47020, n47021,
    n47022, n47023, n47024, n47025, n47026, n47027, n47028, n47029, n47030,
    n47031, n47032, n47033, n47034, n47035, n47036, n47037, n47038, n47039,
    n47040, n47041, n47042, n47043, n47044, n47045, n47046, n47047, n47048,
    n47049, n47050, n47051, n47052, n47053, n47054, n47055, n47056, n47057,
    n47058, n47059, n47060, n47061, n47062, n47063, n47064, n47065, n47066,
    n47067, n47068, n47069, n47070, n47071, n47072, n47073, n47074, n47075,
    n47076, n47077, n47078, n47079, n47080, n47081, n47082, n47083, n47084,
    n47085, n47086, n47087, n47088, n47089, n47090, n47091, n47092, n47093,
    n47094, n47095, n47096, n47097, n47098, n47099, n47100, n47101, n47102,
    n47103, n47104, n47105, n47106, n47107, n47108, n47109, n47110, n47111,
    n47112, n47113, n47114, n47115, n47116, n47117, n47118, n47119, n47120,
    n47121, n47122, n47123, n47124, n47125, n47126, n47127, n47128, n47129,
    n47130, n47131, n47132, n47133, n47134, n47135, n47136, n47137, n47138,
    n47139, n47140, n47141, n47142, n47143, n47144, n47145, n47146, n47147,
    n47148, n47149, n47150, n47151, n47152, n47153, n47154, n47155, n47156,
    n47157, n47158, n47159, n47160, n47161, n47162, n47163, n47164, n47165,
    n47166, n47167, n47168, n47169, n47170, n47171, n47172, n47173, n47174,
    n47175, n47176, n47177, n47178, n47179, n47180, n47181, n47182, n47183,
    n47184, n47185, n47186, n47187, n47188, n47189, n47190, n47191, n47192,
    n47193, n47194, n47195, n47196, n47197, n47198, n47199, n47200, n47201,
    n47202, n47203, n47204, n47205, n47206, n47207, n47208, n47209, n47210,
    n47211, n47212, n47213, n47214, n47215, n47216, n47217, n47218, n47219,
    n47220, n47221, n47222, n47223, n47224, n47225, n47226, n47227, n47228,
    n47229, n47230, n47231, n47232, n47233, n47234, n47235, n47236, n47237,
    n47238, n47239, n47240, n47241, n47242, n47243, n47244, n47245, n47246,
    n47247, n47248, n47249, n47250, n47251, n47252, n47253, n47254, n47255,
    n47256, n47257, n47258, n47259, n47260, n47261, n47262, n47263, n47264,
    n47265, n47266, n47267, n47268, n47269, n47270, n47271, n47272, n47273,
    n47274, n47275, n47276, n47277, n47278, n47279, n47280, n47281, n47282,
    n47283, n47284, n47285, n47286, n47287, n47288, n47289, n47290, n47291,
    n47292, n47293, n47294, n47295, n47296, n47297, n47298, n47299, n47300,
    n47301, n47302, n47303, n47304, n47305, n47306, n47307, n47308, n47309,
    n47310, n47311, n47312, n47313, n47314, n47315, n47316, n47317, n47318,
    n47319, n47320, n47321, n47322, n47323, n47324, n47325, n47326, n47327,
    n47328, n47329, n47330, n47331, n47332, n47333, n47334, n47335, n47336,
    n47337, n47338, n47339, n47340, n47341, n47342, n47343, n47344, n47345,
    n47346, n47347, n47348, n47349, n47350, n47351, n47352, n47353, n47354,
    n47355, n47356, n47357, n47358, n47359, n47360, n47361, n47362, n47363,
    n47364, n47365, n47366, n47367, n47368, n47369, n47370, n47371, n47372,
    n47373, n47374, n47375, n47376, n47377, n47378, n47379, n47380, n47381,
    n47382, n47383, n47384, n47385, n47386, n47387, n47388, n47389, n47390,
    n47391, n47392, n47393, n47394, n47395, n47396, n47397, n47398, n47399,
    n47400, n47401, n47402, n47403, n47404, n47405, n47406, n47407, n47408,
    n47409, n47410, n47411, n47412, n47413, n47414, n47415, n47416, n47417,
    n47418, n47419, n47420, n47421, n47422, n47423, n47424, n47425, n47426,
    n47427, n47428, n47429, n47430, n47431, n47432, n47433, n47434, n47435,
    n47436, n47437, n47438, n47439, n47440, n47441, n47442, n47443, n47444,
    n47445, n47446, n47447, n47448, n47449, n47450, n47451, n47452, n47453,
    n47454, n47455, n47456, n47457, n47458, n47459, n47460, n47461, n47462,
    n47463, n47464, n47465, n47466, n47467, n47468, n47469, n47470, n47471,
    n47472, n47473, n47474, n47475, n47476, n47477, n47478, n47479, n47480,
    n47481, n47482, n47483, n47484, n47485, n47486, n47487, n47488, n47489,
    n47490, n47491, n47492, n47493, n47494, n47495, n47496, n47497, n47498,
    n47499, n47500, n47501, n47502, n47503, n47504, n47505, n47506, n47507,
    n47508, n47509, n47510, n47511, n47512, n47513, n47514, n47515, n47516,
    n47517, n47518, n47519, n47520, n47521, n47522, n47523, n47524, n47525,
    n47526, n47527, n47528, n47529, n47530, n47531, n47532, n47533, n47534,
    n47535, n47536, n47537, n47538, n47539, n47540, n47541, n47542, n47543,
    n47544, n47545, n47546, n47547, n47548, n47549, n47550, n47551, n47552,
    n47553, n47554, n47555, n47556, n47557, n47558, n47559, n47560, n47561,
    n47562, n47563, n47564, n47565, n47566, n47567, n47568, n47569, n47570,
    n47571, n47572, n47573, n47574, n47575, n47576, n47577, n47578, n47579,
    n47580, n47581, n47582, n47583, n47584, n47585, n47586, n47587, n47588,
    n47589, n47590, n47591, n47592, n47593, n47594, n47595, n47596, n47597,
    n47598, n47599, n47600, n47601, n47602, n47603, n47604, n47605, n47606,
    n47607, n47608, n47609, n47610, n47611, n47612, n47613, n47614, n47615,
    n47616, n47617, n47618, n47619, n47620, n47621, n47622, n47623, n47624,
    n47625, n47626, n47627, n47628, n47629, n47630, n47631, n47632, n47633,
    n47634, n47635, n47636, n47637, n47638, n47639, n47640, n47641, n47642,
    n47643, n47644, n47645, n47646, n47647, n47648, n47649, n47650, n47651,
    n47652, n47653, n47654, n47655, n47656, n47657, n47658, n47659, n47660,
    n47661, n47662, n47663, n47664, n47665, n47666, n47667, n47668, n47669,
    n47670, n47671, n47672, n47673, n47674, n47675, n47676, n47677, n47678,
    n47679, n47680, n47681, n47682, n47683, n47684, n47685, n47686, n47687,
    n47688, n47689, n47690, n47691, n47692, n47693, n47694, n47695, n47696,
    n47697, n47698, n47699, n47700, n47701, n47702, n47703, n47704, n47705,
    n47706, n47707, n47708, n47709, n47710, n47711, n47712, n47713, n47714,
    n47715, n47716, n47717, n47718, n47719, n47720, n47721, n47722, n47723,
    n47724, n47725, n47726, n47727, n47728, n47729, n47730, n47731, n47732,
    n47733, n47734, n47735, n47736, n47737, n47738, n47739, n47740, n47741,
    n47742, n47743, n47744, n47745, n47746, n47747, n47748, n47749, n47750,
    n47751, n47752, n47753, n47754, n47755, n47756, n47757, n47758, n47759,
    n47760, n47761, n47762, n47763, n47764, n47765, n47766, n47767, n47768,
    n47769, n47770, n47771, n47772, n47773, n47774, n47775, n47776, n47777,
    n47778, n47779, n47780, n47781, n47782, n47783, n47784, n47785, n47786,
    n47787, n47788, n47789, n47790, n47791, n47792, n47793, n47794, n47795,
    n47796, n47797, n47798, n47799, n47800, n47801, n47802, n47803, n47804,
    n47805, n47806, n47807, n47808, n47809, n47810, n47811, n47812, n47813,
    n47814, n47815, n47816, n47817, n47818, n47819, n47820, n47821, n47822,
    n47823, n47824, n47825, n47826, n47827, n47828, n47829, n47830, n47831,
    n47832, n47833, n47834, n47835, n47836, n47837, n47838, n47839, n47840,
    n47841, n47842, n47843, n47844, n47845, n47846, n47847, n47848, n47849,
    n47850, n47851, n47852, n47853, n47854, n47855, n47856, n47857, n47858,
    n47859, n47860, n47861, n47862, n47863, n47864, n47865, n47866, n47867,
    n47868, n47869, n47870, n47871, n47872, n47873, n47874, n47875, n47876,
    n47877, n47878, n47879, n47880, n47881, n47882, n47883, n47884, n47885,
    n47886, n47887, n47888, n47889, n47890, n47891, n47892, n47893, n47894,
    n47895, n47896, n47897, n47898, n47899, n47900, n47901, n47902, n47903,
    n47904, n47905, n47906, n47907, n47908, n47909, n47910, n47911, n47912,
    n47913, n47914, n47915, n47916, n47917, n47918, n47919, n47920, n47921,
    n47922, n47923, n47924, n47925, n47926, n47927, n47928, n47929, n47930,
    n47931, n47932, n47933, n47934, n47935, n47936, n47937, n47938, n47939,
    n47940, n47941, n47942, n47943, n47944, n47945, n47946, n47947, n47948,
    n47949, n47950, n47951, n47952, n47953, n47954, n47955, n47956, n47957,
    n47958, n47959, n47960, n47961, n47962, n47963, n47964, n47965, n47966,
    n47967, n47968, n47969, n47970, n47971, n47972, n47973, n47974, n47975,
    n47976, n47977, n47978, n47979, n47980, n47981, n47982, n47983, n47984,
    n47985, n47986, n47987, n47988, n47989, n47990, n47991, n47992, n47993,
    n47994, n47995, n47996, n47997, n47998, n47999, n48000, n48001, n48002,
    n48003, n48004, n48005, n48006, n48007, n48008, n48009, n48010, n48011,
    n48012, n48013, n48014, n48015, n48016, n48017, n48018, n48019, n48020,
    n48021, n48022, n48023, n48024, n48025, n48026, n48027, n48028, n48029,
    n48030, n48031, n48032, n48033, n48034, n48035, n48036, n48037, n48038,
    n48039, n48040, n48041, n48042, n48043, n48044, n48045, n48046, n48047,
    n48048, n48049, n48050, n48051, n48052, n48053, n48054, n48055, n48056,
    n48057, n48058, n48059, n48060, n48061, n48062, n48063, n48064, n48065,
    n48066, n48067, n48068, n48069, n48070, n48071, n48072, n48073, n48074,
    n48075, n48076, n48077, n48078, n48079, n48080, n48081, n48082, n48083,
    n48084, n48085, n48086, n48087, n48088, n48089, n48090, n48091, n48092,
    n48093, n48094, n48095, n48096, n48097, n48098, n48099, n48100, n48101,
    n48102, n48103, n48104, n48105, n48106, n48107, n48108, n48109, n48110,
    n48111, n48112, n48113, n48114, n48115, n48116, n48117, n48118, n48119,
    n48120, n48121, n48122, n48123, n48124, n48125, n48126, n48127, n48128,
    n48129, n48130, n48131, n48132, n48133, n48134, n48135, n48136, n48137,
    n48138, n48139, n48140, n48141, n48142, n48143, n48144, n48145, n48146,
    n48147, n48148, n48149, n48150, n48151, n48152, n48153, n48154, n48155,
    n48156, n48157, n48158, n48159, n48160, n48161, n48162, n48163, n48164,
    n48165, n48166, n48167, n48168, n48169, n48170, n48171, n48172, n48173,
    n48174, n48175, n48176, n48177, n48178, n48179, n48180, n48181, n48182,
    n48183, n48184, n48185, n48186, n48187, n48188, n48189, n48190, n48191,
    n48192, n48193, n48194, n48195, n48196, n48197, n48198, n48199, n48200,
    n48201, n48202, n48203, n48204, n48205, n48206, n48207, n48208, n48209,
    n48210, n48211, n48212, n48213, n48214, n48215, n48216, n48217, n48218,
    n48219, n48220, n48221, n48222, n48223, n48224, n48225, n48226, n48227,
    n48228, n48229, n48230, n48231, n48232, n48233, n48234, n48235, n48236,
    n48237, n48238, n48239, n48240, n48241, n48242, n48243, n48244, n48245,
    n48246, n48247, n48248, n48249, n48250, n48251, n48252, n48253, n48254,
    n48255, n48256, n48257, n48258, n48259, n48260, n48261, n48262, n48263,
    n48264, n48265, n48266, n48267, n48268, n48269, n48270, n48271, n48272,
    n48273, n48274, n48275, n48276, n48277, n48278, n48279, n48280, n48281,
    n48282, n48283, n48284, n48285, n48286, n48287, n48288, n48289, n48290,
    n48291, n48292, n48293, n48294, n48295, n48296, n48297, n48298, n48299,
    n48300, n48301, n48302, n48303, n48304, n48305, n48306, n48307, n48308,
    n48309, n48310, n48311, n48312, n48313, n48314, n48315, n48316, n48317,
    n48318, n48319, n48320, n48321, n48322, n48323, n48324, n48325, n48326,
    n48327, n48328, n48329, n48330, n48331, n48332, n48333, n48334, n48335,
    n48336, n48337, n48338, n48339, n48340, n48341, n48342, n48343, n48344,
    n48345, n48346, n48347, n48348, n48349, n48350, n48351, n48352, n48353,
    n48354, n48355, n48356, n48357, n48358, n48359, n48360, n48361, n48362,
    n48363, n48364, n48365, n48366, n48367, n48368, n48369, n48370, n48371,
    n48372, n48373, n48374, n48375, n48376, n48377, n48378, n48379, n48380,
    n48381, n48382, n48383, n48384, n48385, n48386, n48387, n48388, n48389,
    n48390, n48391, n48392, n48393, n48394, n48395, n48396, n48397, n48398,
    n48399, n48400, n48401, n48402, n48403, n48404, n48405, n48406, n48407,
    n48408, n48409, n48410, n48411, n48412, n48413, n48414, n48415, n48416,
    n48417, n48418, n48419, n48420, n48421, n48422, n48423, n48424, n48425,
    n48426, n48427, n48428, n48429, n48430, n48431, n48432, n48433, n48434,
    n48435, n48436, n48437, n48438, n48439, n48440, n48441, n48442, n48443,
    n48444, n48445, n48446, n48447, n48448, n48449, n48450, n48451, n48452,
    n48453, n48454, n48455, n48456, n48457, n48458, n48459, n48460, n48461,
    n48462, n48463, n48464, n48465, n48466, n48467, n48468, n48469, n48470,
    n48471, n48472, n48473, n48474, n48475, n48476, n48477, n48478, n48479,
    n48480, n48481, n48482, n48483, n48484, n48485, n48486, n48487, n48488,
    n48489, n48490, n48491, n48492, n48493, n48494, n48495, n48496, n48497,
    n48498, n48499, n48500, n48501, n48502, n48503, n48504, n48505, n48506,
    n48507, n48508, n48509, n48510, n48511, n48512, n48513, n48514, n48515,
    n48516, n48517, n48518, n48519, n48520, n48521, n48522, n48523, n48524,
    n48525, n48526, n48527, n48528, n48529, n48530, n48531, n48532, n48533,
    n48534, n48535, n48536, n48537, n48538, n48539, n48540, n48541, n48542,
    n48543, n48544, n48545, n48546, n48547, n48548, n48549, n48550, n48551,
    n48552, n48553, n48554, n48555, n48556, n48557, n48558, n48559, n48560,
    n48561, n48562, n48563, n48564, n48565, n48566, n48567, n48568, n48569,
    n48570, n48571, n48572, n48573, n48574, n48575, n48576, n48577, n48578,
    n48579, n48580, n48581, n48582, n48583, n48584, n48585, n48586, n48587,
    n48588, n48589, n48590, n48591, n48592, n48593, n48594, n48595, n48596,
    n48597, n48598, n48599, n48600, n48601, n48602, n48603, n48604, n48605,
    n48606, n48607, n48608, n48609, n48610, n48611, n48612, n48613, n48614,
    n48615, n48616, n48617, n48618, n48619, n48620, n48621, n48622, n48623,
    n48624, n48625, n48626, n48627, n48628, n48629, n48630, n48631, n48632,
    n48633, n48634, n48635, n48636, n48637, n48638, n48639, n48640, n48641,
    n48642, n48643, n48644, n48645, n48646, n48647, n48648, n48649, n48650,
    n48651, n48652, n48653, n48654, n48655, n48656, n48657, n48658, n48659,
    n48660, n48661, n48662, n48663, n48664, n48665, n48666, n48667, n48668,
    n48669, n48670, n48671, n48672, n48673, n48674, n48675, n48676, n48677,
    n48678, n48679, n48680, n48681, n48682, n48683, n48684, n48685, n48686,
    n48687, n48688, n48689, n48690, n48691, n48692, n48693, n48694, n48695,
    n48696, n48697, n48698, n48699, n48700, n48701, n48702, n48703, n48704,
    n48705, n48706, n48707, n48708, n48709, n48710, n48711, n48712, n48713,
    n48714, n48715, n48716, n48717, n48718, n48719, n48720, n48721, n48722,
    n48723, n48724, n48725, n48726, n48727, n48728, n48729, n48730, n48731,
    n48732, n48733, n48734, n48735, n48736, n48737, n48738, n48739, n48740,
    n48741, n48742, n48743, n48744, n48745, n48746, n48747, n48748, n48749,
    n48750, n48751, n48752, n48753, n48754, n48755, n48756, n48757, n48758,
    n48759, n48760, n48761, n48762, n48763, n48764, n48765, n48766, n48767,
    n48768, n48769, n48770, n48771, n48772, n48773, n48774, n48775, n48776,
    n48777, n48778, n48779, n48780, n48781, n48782, n48783, n48784, n48785,
    n48786, n48787, n48788, n48789, n48790, n48791, n48792, n48793, n48794,
    n48795, n48796, n48797, n48798, n48799, n48800, n48801, n48802, n48803,
    n48804, n48805, n48806, n48807, n48808, n48809, n48810, n48811, n48812,
    n48813, n48814, n48815, n48816, n48817, n48818, n48819, n48820, n48821,
    n48822, n48823, n48824, n48825, n48826, n48827, n48828, n48829, n48830,
    n48831, n48832, n48833, n48834, n48835, n48836, n48837, n48838, n48839,
    n48840, n48841, n48842, n48843, n48844, n48845, n48846, n48847, n48848,
    n48849, n48850, n48851, n48852, n48853, n48854, n48855, n48856, n48857,
    n48858, n48859, n48860, n48861, n48862, n48863, n48864, n48865, n48866,
    n48867, n48868, n48869, n48870, n48871, n48872, n48873, n48874, n48875,
    n48876, n48877, n48878, n48879, n48880, n48881, n48882, n48883, n48884,
    n48885, n48886, n48887, n48888, n48889, n48890, n48891, n48892, n48893,
    n48894, n48895, n48896, n48897, n48898, n48899, n48900, n48901, n48902,
    n48903, n48904, n48905, n48906, n48907, n48908, n48909, n48910, n48911,
    n48912, n48913, n48914, n48915, n48916, n48917, n48918, n48919, n48920,
    n48921, n48922, n48923, n48924, n48925, n48926, n48927, n48928, n48929,
    n48930, n48931, n48932, n48933, n48934, n48935, n48936, n48937, n48938,
    n48939, n48940, n48941, n48942, n48943, n48944, n48945, n48946, n48947,
    n48948, n48949, n48950, n48951, n48952, n48953, n48954, n48955, n48956,
    n48957, n48958, n48959, n48960, n48961, n48962, n48963, n48964, n48965,
    n48966, n48967, n48968, n48969, n48970, n48971, n48972, n48973, n48974,
    n48975, n48976, n48977, n48978, n48979, n48980, n48981, n48982, n48983,
    n48984, n48985, n48986, n48987, n48988, n48989, n48990, n48991, n48992,
    n48993, n48994, n48995, n48996, n48997, n48998, n48999, n49000, n49001,
    n49002, n49003, n49004, n49005, n49006, n49007, n49008, n49009, n49010,
    n49011, n49012, n49013, n49014, n49015, n49016, n49017, n49018, n49019,
    n49020, n49021, n49022, n49023, n49024, n49025, n49026, n49027, n49028,
    n49029, n49030, n49031, n49032, n49033, n49034, n49035, n49036, n49037,
    n49038, n49039, n49040, n49041, n49042, n49043, n49044, n49045, n49046,
    n49047, n49048, n49049, n49050, n49051, n49052, n49053, n49054, n49055,
    n49056, n49057, n49058, n49059, n49060, n49061, n49062, n49063, n49064,
    n49065, n49066, n49067, n49068, n49069, n49070, n49071, n49072, n49073,
    n49074, n49075, n49076, n49077, n49078, n49079, n49080, n49081, n49082,
    n49083, n49084, n49085, n49086, n49087, n49088, n49089, n49090, n49091,
    n49092, n49093, n49094, n49095, n49096, n49097, n49098, n49099, n49100,
    n49101, n49102, n49103, n49104, n49105, n49106, n49107, n49108, n49109,
    n49110, n49111, n49112, n49113, n49114, n49115, n49116, n49117, n49118,
    n49119, n49120, n49121, n49122, n49123, n49124, n49125, n49126, n49127,
    n49128, n49129, n49130, n49131, n49132, n49133, n49134, n49135, n49136,
    n49137, n49138, n49139, n49140, n49141, n49142, n49143, n49144, n49145,
    n49146, n49147, n49148, n49149, n49150, n49151, n49152, n49153, n49154,
    n49155, n49156, n49157, n49158, n49159, n49160, n49161, n49162, n49163,
    n49164, n49165, n49166, n49167, n49168, n49169, n49170, n49171, n49172,
    n49173, n49174, n49175, n49176, n49177, n49178, n49179, n49180, n49181,
    n49182, n49183, n49184, n49185, n49186, n49187, n49188, n49189, n49190,
    n49191, n49192, n49193, n49194, n49195, n49196, n49197, n49198, n49199,
    n49200, n49201, n49202, n49203, n49204, n49205, n49206, n49207, n49208,
    n49209, n49210, n49211, n49212, n49213, n49214, n49215, n49216, n49217,
    n49218, n49219, n49220, n49221, n49222, n49223, n49224, n49225, n49226,
    n49227, n49228, n49229, n49230, n49231, n49232, n49233, n49234, n49235,
    n49236, n49237, n49238, n49239, n49240, n49241, n49242, n49243, n49244,
    n49245, n49246, n49247, n49248, n49249, n49250, n49251, n49252, n49253,
    n49254, n49255, n49256, n49257, n49258, n49259, n49260, n49261, n49262,
    n49263, n49264, n49265, n49266, n49267, n49268, n49269, n49270, n49271,
    n49272, n49273, n49274, n49275, n49276, n49277, n49278, n49279, n49280,
    n49281, n49282, n49283, n49284, n49285, n49286, n49287, n49288, n49289,
    n49290, n49291, n49292, n49293, n49294, n49295, n49296, n49297, n49298,
    n49299, n49300, n49301, n49302, n49303, n49304, n49305, n49306, n49307,
    n49308, n49309, n49310, n49311, n49312, n49313, n49314, n49315, n49316,
    n49317, n49318, n49319, n49320, n49321, n49322, n49323, n49324, n49325,
    n49326, n49327, n49328, n49329, n49330, n49331, n49332, n49333, n49334,
    n49335, n49336, n49337, n49338, n49339, n49340, n49341, n49342, n49343,
    n49344, n49345, n49346, n49347, n49348, n49349, n49350, n49351, n49352,
    n49353, n49354, n49355, n49356, n49357, n49358, n49359, n49360, n49361,
    n49362, n49363, n49364, n49365, n49366, n49367, n49368, n49369, n49370,
    n49371, n49372, n49373, n49374, n49375, n49376, n49377, n49378, n49379,
    n49380, n49381, n49382, n49383, n49384, n49385, n49386, n49387, n49388,
    n49389, n49390, n49391, n49392, n49393, n49394, n49395, n49396, n49397,
    n49398, n49399, n49400, n49401, n49402, n49403, n49404, n49405, n49406,
    n49407, n49408, n49409, n49410, n49411, n49412, n49413, n49414, n49415,
    n49416, n49417, n49418, n49419, n49420, n49421, n49422, n49423, n49424,
    n49425, n49426, n49427, n49428, n49429, n49430, n49431, n49432, n49433,
    n49434, n49435, n49436, n49437, n49438, n49439, n49440, n49441, n49442,
    n49443, n49444, n49445, n49446, n49447, n49448, n49449, n49450, n49451,
    n49452, n49453, n49454, n49455, n49456, n49457, n49458, n49459, n49460,
    n49461, n49462, n49463, n49464, n49465, n49466, n49467, n49468, n49469,
    n49470, n49471, n49472, n49473, n49474, n49475, n49476, n49477, n49478,
    n49479, n49480, n49481, n49482, n49483, n49484, n49485, n49486, n49487,
    n49488, n49489, n49490, n49491, n49492, n49493, n49494, n49495, n49496,
    n49497, n49498, n49499, n49500, n49501, n49502, n49503, n49504, n49505,
    n49506, n49507, n49508, n49509, n49510, n49511, n49512, n49513, n49514,
    n49515, n49516, n49517, n49518, n49519, n49520, n49521, n49522, n49523,
    n49524, n49525, n49526, n49527, n49528, n49529, n49530, n49531, n49532,
    n49533, n49534, n49535, n49536, n49537, n49538, n49539, n49540, n49541,
    n49542, n49543, n49544, n49545, n49546, n49547, n49548, n49549, n49550,
    n49551, n49552, n49553, n49554, n49555, n49556, n49557, n49558, n49559,
    n49560, n49561, n49562, n49563, n49564, n49565, n49566, n49567, n49568,
    n49569, n49570, n49571, n49572, n49573, n49574, n49575, n49576, n49577,
    n49578, n49579, n49580, n49581, n49582, n49583, n49584, n49585, n49586,
    n49587, n49588, n49589, n49590, n49591, n49592, n49593, n49594, n49595,
    n49596, n49597, n49598, n49599, n49600, n49601, n49602, n49603, n49604,
    n49605, n49606, n49607, n49608, n49609, n49610, n49611, n49612, n49613,
    n49614, n49615, n49616, n49617, n49618, n49619, n49620, n49621, n49622,
    n49623, n49624, n49625, n49626, n49627, n49628, n49629, n49630, n49631,
    n49632, n49633, n49634, n49635, n49636, n49637, n49638, n49639, n49640,
    n49641, n49642, n49643, n49644, n49645, n49646, n49647, n49648, n49649,
    n49650, n49651, n49652, n49653, n49654, n49655, n49656, n49657, n49658,
    n49659, n49660, n49661, n49662, n49663, n49664, n49665, n49666, n49667,
    n49668, n49669, n49670, n49671, n49672, n49673, n49674, n49675, n49676,
    n49677, n49678, n49679, n49680, n49681, n49682, n49683, n49684, n49685,
    n49686, n49687, n49688, n49689, n49690, n49691, n49692, n49693, n49694,
    n49695, n49696, n49697, n49698, n49699, n49700, n49701, n49702, n49703,
    n49704, n49705, n49706, n49707, n49708, n49709, n49710, n49711, n49712,
    n49713, n49714, n49715, n49716, n49717, n49718, n49719, n49720, n49721,
    n49722, n49723, n49724, n49725, n49726, n49727, n49728, n49729, n49730,
    n49731, n49732, n49733, n49734, n49735, n49736, n49737, n49738, n49739,
    n49740, n49741, n49742, n49743, n49744, n49745, n49746, n49747, n49748,
    n49749, n49750, n49751, n49752, n49753, n49754, n49755, n49756, n49757,
    n49758, n49759, n49760, n49761, n49762, n49763, n49764, n49765, n49766,
    n49767, n49768, n49769, n49770, n49771, n49772, n49773, n49774, n49775,
    n49776, n49777, n49778, n49779, n49780, n49781, n49782, n49783, n49784,
    n49785, n49786, n49787, n49788, n49789, n49790, n49791, n49792, n49793,
    n49794, n49795, n49796, n49797, n49798, n49799, n49800, n49801, n49802,
    n49803, n49804, n49805, n49806, n49807, n49808, n49809, n49810, n49811,
    n49812, n49813, n49814, n49815, n49816, n49817, n49818, n49819, n49820,
    n49821, n49822, n49823, n49824, n49825, n49826, n49827, n49828, n49829,
    n49830, n49831, n49832, n49833, n49834, n49835, n49836, n49837, n49838,
    n49839, n49840, n49841, n49842, n49843, n49844, n49845, n49846, n49847,
    n49848, n49849, n49850, n49851, n49852, n49853, n49854, n49855, n49856,
    n49857, n49858, n49859, n49860, n49861, n49862, n49863, n49864, n49865,
    n49866, n49867, n49868, n49869, n49870, n49871, n49872, n49873, n49874,
    n49875, n49876, n49877, n49878, n49879, n49880, n49881, n49882, n49883,
    n49884, n49885, n49886, n49887, n49888, n49889, n49890, n49891, n49892,
    n49893, n49894, n49895, n49896, n49897, n49898, n49899, n49900, n49901,
    n49902, n49903, n49904, n49905, n49906, n49907, n49908, n49909, n49910,
    n49911, n49912, n49913, n49914, n49915, n49916, n49917, n49918, n49919,
    n49920, n49921, n49922, n49923, n49924, n49925, n49926, n49927, n49928,
    n49929, n49930, n49931, n49932, n49933, n49934, n49935, n49936, n49937,
    n49938, n49939, n49940, n49941, n49942, n49943, n49944, n49945, n49946,
    n49947, n49948, n49949, n49950, n49951, n49952, n49953, n49954, n49955,
    n49956, n49957, n49958, n49959, n49960, n49961, n49962, n49963, n49964,
    n49965, n49966, n49967, n49968, n49969, n49970, n49971, n49972, n49973,
    n49974, n49975, n49976, n49977, n49978, n49979, n49980, n49981, n49982,
    n49983, n49984, n49985, n49986, n49987, n49988, n49989, n49990, n49991,
    n49992, n49993, n49994, n49995, n49996, n49997, n49998, n49999, n50000,
    n50001, n50002, n50003, n50004, n50005, n50006, n50007, n50008, n50009,
    n50010, n50011, n50012, n50013, n50014, n50015, n50016, n50017, n50018,
    n50019, n50020, n50021, n50022, n50023, n50024, n50025, n50026, n50027,
    n50028, n50029, n50030, n50031, n50032, n50033, n50034, n50035, n50036,
    n50037, n50038, n50039, n50040, n50041, n50042, n50043, n50044, n50045,
    n50046, n50047, n50048, n50049, n50050, n50051, n50052, n50053, n50054,
    n50055, n50056, n50057, n50058, n50059, n50060, n50061, n50062, n50063,
    n50064, n50065, n50066, n50067, n50068, n50069, n50070, n50071, n50072,
    n50073, n50074, n50075, n50076, n50077, n50078, n50079, n50080, n50081,
    n50082, n50083, n50084, n50085, n50086, n50087, n50088, n50089, n50090,
    n50091, n50092, n50093, n50094, n50095, n50096, n50097, n50098, n50099,
    n50100, n50101, n50102, n50103, n50104, n50105, n50106, n50107, n50108,
    n50109, n50110, n50111, n50112, n50113, n50114, n50115, n50116, n50117,
    n50118, n50119, n50120, n50121, n50122, n50123, n50124, n50125, n50126,
    n50127, n50128, n50129, n50130, n50131, n50132, n50133, n50134, n50135,
    n50136, n50137, n50138, n50139, n50140, n50141, n50142, n50143, n50144,
    n50145, n50146, n50147, n50148, n50149, n50150, n50151, n50152, n50153,
    n50154, n50155, n50156, n50157, n50158, n50159, n50160, n50161, n50162,
    n50163, n50164, n50165, n50166, n50167, n50168, n50169, n50170, n50171,
    n50172, n50173, n50174, n50175, n50176, n50177, n50178, n50179, n50180,
    n50181, n50182, n50183, n50184, n50185, n50186, n50187, n50188, n50189,
    n50190, n50191, n50192, n50193, n50194, n50195, n50196, n50197, n50198,
    n50199, n50200, n50201, n50202, n50203, n50204, n50205, n50206, n50207,
    n50208, n50209, n50210, n50211, n50212, n50213, n50214, n50215, n50216,
    n50217, n50218, n50219, n50220, n50221, n50222, n50223, n50224, n50225,
    n50226, n50227, n50228, n50229, n50230, n50231, n50232, n50233, n50234,
    n50235, n50236, n50237, n50238, n50239, n50240, n50241, n50242, n50243,
    n50244, n50245, n50246, n50247, n50248, n50249, n50250, n50251, n50252,
    n50253, n50254, n50255, n50256, n50257, n50258, n50259, n50260, n50261,
    n50262, n50263, n50264, n50265, n50266, n50267, n50268, n50269, n50270,
    n50271, n50272, n50273, n50274, n50275, n50276, n50277, n50278, n50279,
    n50280, n50281, n50282, n50283, n50284, n50285, n50286, n50287, n50288,
    n50289, n50290, n50291, n50292, n50293, n50294, n50295, n50296, n50297,
    n50298, n50299, n50300, n50301, n50302, n50303, n50304, n50305, n50306,
    n50307, n50308, n50309, n50310, n50311, n50312, n50313, n50314, n50315,
    n50316, n50317, n50318, n50319, n50320, n50321, n50322, n50323, n50324,
    n50325, n50326, n50327, n50328, n50329, n50330, n50331, n50332, n50333,
    n50334, n50335, n50336, n50337, n50338, n50339, n50340, n50341, n50342,
    n50343, n50344, n50345, n50346, n50347, n50348, n50349, n50350, n50351,
    n50352, n50353, n50354, n50355, n50356, n50357, n50358, n50359, n50360,
    n50361, n50362, n50363, n50364, n50365, n50366, n50367, n50368, n50369,
    n50370, n50371, n50372, n50373, n50374, n50375, n50376, n50377, n50378,
    n50379, n50380, n50381, n50382, n50383, n50384, n50385, n50386, n50387,
    n50388, n50389, n50390, n50391, n50392, n50393, n50394, n50395, n50396,
    n50397, n50398, n50399, n50400, n50401, n50402, n50403, n50404, n50405,
    n50406, n50407, n50408, n50409, n50410, n50411, n50412, n50413, n50414,
    n50415, n50416, n50417, n50418, n50419, n50420, n50421, n50422, n50423,
    n50424, n50425, n50426, n50427, n50428, n50429, n50430, n50431, n50432,
    n50433, n50434, n50435, n50436, n50437, n50438, n50439, n50440, n50441,
    n50442, n50443, n50444, n50445, n50446, n50447, n50448, n50449, n50450,
    n50451, n50452, n50453, n50454, n50455, n50456, n50457, n50458, n50459,
    n50460, n50461, n50462, n50463, n50464, n50465, n50466, n50467, n50468,
    n50469, n50470, n50471, n50472, n50473, n50474, n50475, n50476, n50477,
    n50478, n50479, n50480, n50481, n50482, n50483, n50484, n50485, n50486,
    n50487, n50488, n50489, n50490, n50491, n50492, n50493, n50494, n50495,
    n50496, n50497, n50498, n50499, n50500, n50501, n50502, n50503, n50504,
    n50505, n50506, n50507, n50508, n50509, n50510, n50511, n50512, n50513,
    n50514, n50515, n50516, n50517, n50518, n50519, n50520, n50521, n50522,
    n50523, n50524, n50525, n50526, n50527, n50528, n50529, n50530, n50531,
    n50532, n50533, n50534, n50535, n50536, n50537, n50538, n50539, n50540,
    n50541, n50542, n50543, n50544, n50545, n50546, n50547, n50548, n50549,
    n50550, n50551, n50552, n50553, n50554, n50555, n50556, n50557, n50558,
    n50559, n50560, n50561, n50562, n50563, n50564, n50565, n50566, n50567,
    n50568, n50569, n50570, n50571, n50572, n50573, n50574, n50575, n50576,
    n50577, n50578, n50579, n50580, n50581, n50582, n50583, n50584, n50585,
    n50586, n50587, n50588, n50589, n50590, n50591, n50592, n50593, n50594,
    n50595, n50596, n50597, n50598, n50599, n50600, n50601, n50602, n50603,
    n50604, n50605, n50606, n50607, n50608, n50609, n50610, n50611, n50612,
    n50613, n50614, n50615, n50616, n50617, n50618, n50619, n50620, n50621,
    n50622, n50623, n50624, n50625, n50626, n50627, n50628, n50629, n50630,
    n50631, n50632, n50633, n50634, n50635, n50636, n50637, n50638, n50639,
    n50640, n50641, n50642, n50643, n50644, n50645, n50646, n50647, n50648,
    n50649, n50650, n50651, n50652, n50653, n50654, n50655, n50656, n50657,
    n50658, n50659, n50660, n50661, n50662, n50663, n50664, n50665, n50666,
    n50667, n50668, n50669, n50670, n50671, n50672, n50673, n50674, n50675,
    n50676, n50677, n50678, n50679, n50680, n50681, n50682, n50683, n50684,
    n50685, n50686, n50687, n50688, n50689, n50690, n50691, n50692, n50693,
    n50694, n50695, n50696, n50697, n50698, n50699, n50700, n50701, n50702,
    n50703, n50704, n50705, n50706, n50707, n50708, n50709, n50710, n50711,
    n50712, n50713, n50714, n50715, n50716, n50717, n50718, n50719, n50720,
    n50721, n50722, n50723, n50724, n50725, n50726, n50727, n50728, n50729,
    n50730, n50731, n50732, n50733, n50734, n50735, n50736, n50737, n50738,
    n50739, n50740, n50741, n50742, n50743, n50744, n50745, n50746, n50747,
    n50748, n50749, n50750, n50751, n50752, n50753, n50754, n50755, n50756,
    n50757, n50758, n50759, n50760, n50761, n50762, n50763, n50764, n50765,
    n50766, n50767, n50768, n50769, n50770, n50771, n50772, n50773, n50774,
    n50775, n50776, n50777, n50778, n50779, n50780, n50781, n50782, n50783,
    n50784, n50785, n50786, n50787, n50788, n50789, n50790, n50791, n50792,
    n50793, n50794, n50795, n50796, n50797, n50798, n50799, n50800, n50801,
    n50802, n50803, n50804, n50805, n50806, n50807, n50808, n50809, n50810,
    n50811, n50812, n50813, n50814, n50815, n50816, n50817, n50818, n50819,
    n50820, n50821, n50822, n50823, n50824, n50825, n50826, n50827, n50828,
    n50829, n50830, n50831, n50832, n50833, n50834, n50835, n50836, n50837,
    n50838, n50839, n50840, n50841, n50842, n50843, n50844, n50845, n50846,
    n50847, n50848, n50849, n50850, n50851, n50852, n50853, n50854, n50855,
    n50856, n50857, n50858, n50859, n50860, n50861, n50862, n50863, n50864,
    n50865, n50866, n50867, n50868, n50869, n50870, n50871, n50872, n50873,
    n50874, n50875, n50876, n50877, n50878, n50879, n50880, n50881, n50882,
    n50883, n50884, n50885, n50886, n50887, n50888, n50889, n50890, n50891,
    n50892, n50893, n50894, n50895, n50896, n50897, n50898, n50899, n50900,
    n50901, n50902, n50903, n50904, n50905, n50906, n50907, n50908, n50909,
    n50910, n50911, n50912, n50913, n50914, n50915, n50916, n50917, n50918,
    n50919, n50920, n50921, n50922, n50923, n50924, n50925, n50926, n50927,
    n50928, n50929, n50930, n50931, n50932, n50933, n50934, n50935, n50936,
    n50937, n50938, n50939, n50940, n50941, n50942, n50943, n50944, n50945,
    n50946, n50947, n50948, n50949, n50950, n50951, n50952, n50953, n50954,
    n50955, n50956, n50957, n50958, n50959, n50960, n50961, n50962, n50963,
    n50964, n50965, n50966, n50967, n50968, n50969, n50970, n50971, n50972,
    n50973, n50974, n50975, n50976, n50977, n50978, n50979, n50980, n50981,
    n50982, n50983, n50984, n50985, n50986, n50987, n50988, n50989, n50990,
    n50991, n50992, n50993, n50994, n50995, n50996, n50997, n50998, n50999,
    n51000, n51001, n51002, n51003, n51004, n51005, n51006, n51007, n51008,
    n51009, n51010, n51011, n51012, n51013, n51014, n51015, n51016, n51017,
    n51018, n51019, n51020, n51021, n51022, n51023, n51024, n51025, n51026,
    n51027, n51028, n51029, n51030, n51031, n51032, n51033, n51034, n51035,
    n51036, n51037, n51038, n51039, n51040, n51041, n51042, n51043, n51044,
    n51045, n51046, n51047, n51048, n51049, n51050, n51051, n51052, n51053,
    n51054, n51055, n51056, n51057, n51058, n51059, n51060, n51061, n51062,
    n51063, n51064, n51065, n51066, n51067, n51068, n51069, n51070, n51071,
    n51072, n51073, n51074, n51075, n51076, n51077, n51078, n51079, n51080,
    n51081, n51082, n51083, n51084, n51085, n51086, n51087, n51088, n51089,
    n51090, n51091, n51092, n51093, n51094, n51095, n51096, n51097, n51098,
    n51099, n51100, n51101, n51102, n51103, n51104, n51105, n51106, n51107,
    n51108, n51109, n51110, n51111, n51112, n51113, n51114, n51115, n51116,
    n51117, n51118, n51119, n51120, n51121, n51122, n51123, n51124, n51125,
    n51126, n51127, n51128, n51129, n51130, n51131, n51132, n51133, n51134,
    n51135, n51136, n51137, n51138, n51139, n51140, n51141, n51142, n51143,
    n51144, n51145, n51146, n51147, n51148, n51149, n51150, n51151, n51152,
    n51153, n51154, n51155, n51156, n51157, n51158, n51159, n51160, n51161,
    n51162, n51163, n51164, n51165, n51166, n51167, n51168, n51169, n51170,
    n51171, n51172, n51173, n51174, n51175, n51176, n51177, n51178, n51179,
    n51180, n51181, n51182, n51183, n51184, n51185, n51186, n51187, n51188,
    n51189, n51190, n51191, n51192, n51193, n51194, n51195, n51196, n51197,
    n51198, n51199, n51200, n51201, n51202, n51203, n51204, n51205, n51206,
    n51207, n51208, n51209, n51210, n51211, n51212, n51213, n51214, n51215,
    n51216, n51217, n51218, n51219, n51220, n51221, n51222, n51223, n51224,
    n51225, n51226, n51227, n51228, n51229, n51230, n51231, n51232, n51233,
    n51234, n51235, n51236, n51237, n51238, n51239, n51240, n51241, n51242,
    n51243, n51244, n51245, n51246, n51247, n51248, n51249, n51250, n51251,
    n51252, n51253, n51254, n51255, n51256, n51257, n51258, n51259, n51260,
    n51261, n51262, n51263, n51264, n51265, n51266, n51267, n51268, n51269,
    n51270, n51271, n51272, n51273, n51274, n51275, n51276, n51277, n51278,
    n51279, n51280, n51281, n51282, n51283, n51284, n51285, n51286, n51287,
    n51288, n51289, n51290, n51291, n51292, n51293, n51294, n51295, n51296,
    n51297, n51298, n51299, n51300, n51301, n51302, n51303, n51304, n51305,
    n51306, n51307, n51308, n51309, n51310, n51311, n51312, n51313, n51314,
    n51315, n51316, n51317, n51318, n51319, n51320, n51321, n51322, n51323,
    n51324, n51325, n51326, n51327, n51328, n51329, n51330, n51331, n51332,
    n51333, n51334, n51335, n51336, n51337, n51338, n51339, n51340, n51341,
    n51342, n51343, n51344, n51345, n51346, n51347, n51348, n51349, n51350,
    n51351, n51352, n51353, n51354, n51355, n51356, n51357, n51358, n51359,
    n51360, n51361, n51362, n51363, n51364, n51365, n51366, n51367, n51368,
    n51369, n51370, n51371, n51372, n51373, n51374, n51375, n51376, n51377,
    n51378, n51379, n51380, n51381, n51382, n51383, n51384, n51385, n51386,
    n51387, n51388, n51389, n51390, n51391, n51392, n51393, n51394, n51395,
    n51396, n51397, n51398, n51399, n51400, n51401, n51402, n51403, n51404,
    n51405, n51406, n51407, n51408, n51409, n51410, n51411, n51412, n51413,
    n51414, n51415, n51416, n51417, n51418, n51419, n51420, n51421, n51422,
    n51423, n51424, n51425, n51426, n51427, n51428, n51429, n51430, n51431,
    n51432, n51433, n51434, n51435, n51436, n51437, n51438, n51439, n51440,
    n51441, n51442, n51443, n51444, n51445, n51446, n51447, n51448, n51449,
    n51450, n51451, n51452, n51453, n51454, n51455, n51456, n51457, n51458,
    n51459, n51460, n51461, n51462, n51463, n51464, n51465, n51466, n51467,
    n51468, n51469, n51470, n51471, n51472, n51473, n51474, n51475, n51476,
    n51477, n51478, n51479, n51480, n51481, n51482, n51483, n51484, n51485,
    n51486, n51487, n51488, n51489, n51490, n51491, n51492, n51493, n51494,
    n51495, n51496, n51497, n51498, n51499, n51500, n51501, n51502, n51503,
    n51504, n51505, n51506, n51507, n51508, n51509, n51510, n51511, n51512,
    n51513, n51514, n51515, n51516, n51517, n51518, n51519, n51520, n51521,
    n51522, n51523, n51524, n51525, n51526, n51527, n51528, n51529, n51530,
    n51531, n51532, n51533, n51534, n51535, n51536, n51537, n51538, n51539,
    n51540, n51541, n51542, n51543, n51544, n51545, n51546, n51547, n51548,
    n51549, n51550, n51551, n51552, n51553, n51554, n51555, n51556, n51557,
    n51558, n51559, n51560, n51561, n51562, n51563, n51564, n51565, n51566,
    n51567, n51568, n51569, n51570, n51571, n51572, n51573, n51574, n51575,
    n51576, n51577, n51578, n51579, n51580, n51581, n51582, n51583, n51584,
    n51585, n51586, n51587, n51588, n51589, n51590, n51591, n51592, n51593,
    n51594, n51595, n51596, n51597, n51598, n51599, n51600, n51601, n51602,
    n51603, n51604, n51605, n51606, n51607, n51608, n51609, n51610, n51611,
    n51612, n51613, n51614, n51615, n51616, n51617, n51618, n51619, n51620,
    n51621, n51622, n51623, n51624, n51625, n51626, n51627, n51628, n51629,
    n51630, n51631, n51632, n51633, n51634, n51635, n51636, n51637, n51638,
    n51639, n51640, n51641, n51642, n51643, n51644, n51645, n51646, n51647,
    n51648, n51649, n51650, n51651, n51652, n51653, n51654, n51655, n51656,
    n51657, n51658, n51659, n51660, n51661, n51662, n51663, n51664, n51665,
    n51666, n51667, n51668, n51669, n51670, n51671, n51672, n51673, n51674,
    n51675, n51676, n51677, n51678, n51679, n51680, n51681, n51682, n51683,
    n51684, n51685, n51686, n51687, n51688, n51689, n51690, n51691, n51692,
    n51693, n51694, n51695, n51696, n51697, n51698, n51699, n51700, n51701,
    n51702, n51703, n51704, n51705, n51706, n51707, n51708, n51709, n51710,
    n51711, n51712, n51713, n51714, n51715, n51716, n51717, n51718, n51719,
    n51720, n51721, n51722, n51723, n51724, n51725, n51726, n51727, n51728,
    n51729, n51730, n51731, n51732, n51733, n51734, n51735, n51736, n51737,
    n51738, n51739, n51740, n51741, n51742, n51743, n51744, n51745, n51746,
    n51747, n51748, n51749, n51750, n51751, n51752, n51753, n51754, n51755,
    n51756, n51757, n51758, n51759, n51760, n51761, n51762, n51763, n51764,
    n51765, n51766, n51767, n51768, n51769, n51770, n51771, n51772, n51773,
    n51774, n51775, n51776, n51777, n51778, n51779, n51780, n51781, n51782,
    n51783, n51784, n51785, n51786, n51787, n51788, n51789, n51790, n51791,
    n51792, n51793, n51794, n51795, n51796, n51797, n51798, n51799, n51800,
    n51801, n51802, n51803, n51804, n51805, n51806, n51807, n51808, n51809,
    n51810, n51811, n51812, n51813, n51814, n51815, n51816, n51817, n51818,
    n51819, n51820, n51821, n51822, n51823, n51824, n51825, n51826, n51827,
    n51828, n51829, n51830, n51831, n51832, n51833, n51834, n51835, n51836,
    n51837, n51838, n51839, n51840, n51841, n51842, n51843, n51844, n51845,
    n51846, n51847, n51848, n51849, n51850, n51851, n51852, n51853, n51854,
    n51855, n51856, n51857, n51858, n51859, n51860, n51861, n51862, n51863,
    n51864, n51865, n51866, n51867, n51868, n51869, n51870, n51871, n51872,
    n51873, n51874, n51875, n51876, n51877, n51878, n51879, n51880, n51881,
    n51882, n51883, n51884, n51885, n51886, n51887, n51888, n51889, n51890,
    n51891, n51892, n51893, n51894, n51895, n51896, n51897, n51898, n51899,
    n51900, n51901, n51902, n51903, n51904, n51905, n51906, n51907, n51908,
    n51909, n51910, n51911, n51912, n51913, n51914, n51915, n51916, n51917,
    n51918, n51919, n51920, n51921, n51922, n51923, n51924, n51925, n51926,
    n51927, n51928, n51929, n51930, n51931, n51932, n51933, n51934, n51935,
    n51936, n51937, n51938, n51939, n51940, n51941, n51942, n51943, n51944,
    n51945, n51946, n51947, n51948, n51949, n51950, n51951, n51952, n51953,
    n51954, n51955, n51956, n51957, n51958, n51959, n51960, n51961, n51962,
    n51963, n51964, n51965, n51966, n51967, n51968, n51969, n51970, n51971,
    n51972, n51973, n51974, n51975, n51976, n51977, n51978, n51979, n51980,
    n51981, n51982, n51983, n51984, n51985, n51986, n51987, n51988, n51989,
    n51990, n51991, n51992, n51993, n51994, n51995, n51996, n51997, n51998,
    n51999, n52000, n52001, n52002, n52003, n52004, n52005, n52006, n52007,
    n52008, n52009, n52010, n52011, n52012, n52013, n52014, n52015, n52016,
    n52017, n52018, n52019, n52020, n52021, n52022, n52023, n52024, n52025,
    n52026, n52027, n52028, n52029, n52030, n52031, n52032, n52033, n52034,
    n52035, n52036, n52037, n52038, n52039, n52040, n52041, n52042, n52043,
    n52044, n52045, n52046, n52047, n52048, n52049, n52050, n52051, n52052,
    n52053, n52054, n52055, n52056, n52057, n52058, n52059, n52060, n52061,
    n52062, n52063, n52064, n52065, n52066, n52067, n52068, n52069, n52070,
    n52071, n52072, n52073, n52074, n52075, n52076, n52077, n52078, n52079,
    n52080, n52081, n52082, n52083, n52084, n52085, n52086, n52087, n52088,
    n52089, n52090, n52091, n52092, n52093, n52094, n52095, n52096, n52097,
    n52098, n52099, n52100, n52101, n52102, n52103, n52104, n52105, n52106,
    n52107, n52108, n52109, n52110, n52111, n52112, n52113, n52114, n52115,
    n52116, n52117, n52118, n52119, n52120, n52121, n52122, n52123, n52124,
    n52125, n52126, n52127, n52128, n52129, n52130, n52131, n52132, n52133,
    n52134, n52135, n52136, n52137, n52138, n52139, n52140, n52141, n52142,
    n52143, n52144, n52145, n52146, n52147, n52148, n52149, n52150, n52151,
    n52152, n52153, n52154, n52155, n52156, n52157, n52158, n52159, n52160,
    n52161, n52162, n52163, n52164, n52165, n52166, n52167, n52168, n52169,
    n52170, n52171, n52172, n52173, n52174, n52175, n52176, n52177, n52178,
    n52179, n52180, n52181, n52182, n52183, n52184, n52185, n52186, n52187,
    n52188, n52189, n52190, n52191, n52192, n52193, n52194, n52195, n52196,
    n52197, n52198, n52199, n52200, n52201, n52202, n52203, n52204, n52205,
    n52206, n52207, n52208, n52209, n52210, n52211, n52212, n52213, n52214,
    n52215, n52216, n52217, n52218, n52219, n52220, n52221, n52222, n52223,
    n52224, n52225, n52226, n52227, n52228, n52229, n52230, n52231, n52232,
    n52233, n52234, n52235, n52236, n52237, n52238, n52239, n52240, n52241,
    n52242, n52243, n52244, n52245, n52246, n52247, n52248, n52249, n52250,
    n52251, n52252, n52253, n52254, n52255, n52256, n52257, n52258, n52259,
    n52260, n52261, n52262, n52263, n52264, n52265, n52266, n52267, n52268,
    n52269, n52270, n52271, n52272, n52273, n52274, n52275, n52276, n52277,
    n52278, n52279, n52280, n52281, n52282, n52283, n52284, n52285, n52286,
    n52287, n52288, n52289, n52290, n52291, n52292, n52293, n52294, n52295,
    n52296, n52297, n52298, n52299, n52300, n52301, n52302, n52303, n52304,
    n52305, n52306, n52307, n52308, n52309, n52310, n52311, n52312, n52313,
    n52314, n52315, n52316, n52317, n52318, n52319, n52320, n52321, n52322,
    n52323, n52324, n52325, n52326, n52327, n52328, n52329, n52330, n52331,
    n52332, n52333, n52334, n52335, n52336, n52337, n52338, n52339, n52340,
    n52341, n52342, n52343, n52344, n52345, n52346, n52347, n52348, n52349,
    n52350, n52351, n52352, n52353, n52354, n52355, n52356, n52357, n52358,
    n52359, n52360, n52361, n52362, n52363, n52364, n52365, n52366, n52367,
    n52368, n52369, n52370, n52371, n52372, n52373, n52374, n52375, n52376,
    n52377, n52378, n52379, n52380, n52381, n52382, n52383, n52384, n52385,
    n52386, n52387, n52388, n52389, n52390, n52391, n52392, n52393, n52394,
    n52395, n52396, n52397, n52398, n52399, n52400, n52401, n52402, n52403,
    n52404, n52405, n52406, n52407, n52408, n52409, n52410, n52411, n52412,
    n52413, n52414, n52415, n52416, n52417, n52418, n52419, n52420, n52421,
    n52422, n52423, n52424, n52425, n52426, n52427, n52428, n52429, n52430,
    n52431, n52432, n52433, n52434, n52435, n52436, n52437, n52438, n52439,
    n52440, n52441, n52442, n52443, n52444, n52445, n52446, n52447, n52448,
    n52449, n52450, n52451, n52452, n52453, n52454, n52455, n52456, n52457,
    n52458, n52459, n52460, n52461, n52462, n52463, n52464, n52465, n52466,
    n52467, n52468, n52469, n52470, n52471, n52472, n52473, n52474, n52475,
    n52476, n52477, n52478, n52479, n52480, n52481, n52482, n52483, n52484,
    n52485, n52486, n52487, n52488, n52489, n52490, n52491, n52492, n52493,
    n52494, n52495, n52496, n52497, n52498, n52499, n52500, n52501, n52502,
    n52503, n52504, n52505, n52506, n52507, n52508, n52509, n52510, n52511,
    n52512, n52513, n52514, n52515, n52516, n52517, n52518, n52519, n52520,
    n52521, n52522, n52523, n52524, n52525, n52526, n52527, n52528, n52529,
    n52530, n52531, n52532, n52533, n52534, n52535, n52536, n52537, n52538,
    n52539, n52540, n52541, n52542, n52543, n52544, n52545, n52546, n52547,
    n52548, n52549, n52550, n52551, n52552, n52553, n52554, n52555, n52556,
    n52557, n52558, n52559, n52560, n52561, n52562, n52563, n52564, n52565,
    n52566, n52567, n52568, n52569, n52570, n52571, n52572, n52573, n52574,
    n52575, n52576, n52577, n52578, n52579, n52580, n52581, n52582, n52583,
    n52584, n52585, n52586, n52587, n52588, n52589, n52590, n52591, n52592,
    n52593, n52594, n52595, n52596, n52597, n52598, n52599, n52600, n52601,
    n52602, n52603, n52604, n52605, n52606, n52607, n52608, n52609, n52610,
    n52611, n52612, n52613, n52614, n52615, n52616, n52617, n52618, n52619,
    n52620, n52621, n52622, n52623, n52624, n52625, n52626, n52627, n52628,
    n52629, n52630, n52631, n52632, n52633, n52634, n52635, n52636, n52637,
    n52638, n52639, n52640, n52641, n52642, n52643, n52644, n52645, n52646,
    n52647, n52648, n52649, n52650, n52651, n52652, n52653, n52654, n52655,
    n52656, n52657, n52658, n52659, n52660, n52661, n52662, n52663, n52664,
    n52665, n52666, n52667, n52668, n52669, n52670, n52671, n52672, n52673,
    n52674, n52675, n52676, n52677, n52678, n52679, n52680, n52681, n52682,
    n52683, n52684, n52685, n52686, n52687, n52688, n52689, n52690, n52691,
    n52692, n52693, n52694, n52695, n52696, n52697, n52698, n52699, n52700,
    n52701, n52702, n52703, n52704, n52705, n52706, n52707, n52708, n52709,
    n52710, n52711, n52712, n52713, n52714, n52715, n52716, n52717, n52718,
    n52719, n52720, n52721, n52722, n52723, n52724, n52725, n52726, n52727,
    n52728, n52729, n52730, n52731, n52732, n52733, n52734, n52735, n52736,
    n52737, n52738, n52739, n52740, n52741, n52742, n52743, n52744, n52745,
    n52746, n52747, n52748, n52749, n52750, n52751, n52752, n52753, n52754,
    n52755, n52756, n52757, n52758, n52759, n52760, n52761, n52762, n52763,
    n52764, n52765, n52766, n52767, n52768, n52769, n52770, n52771, n52772,
    n52773, n52774, n52775, n52776, n52777, n52778, n52779, n52780, n52781,
    n52782, n52783, n52784, n52785, n52786, n52787, n52788, n52789, n52790,
    n52791, n52792, n52793, n52794, n52795, n52796, n52797, n52798, n52799,
    n52800, n52801, n52802, n52803, n52804, n52805, n52806, n52807, n52808,
    n52809, n52810, n52811, n52812, n52813, n52814, n52815, n52816, n52817,
    n52818, n52819, n52820, n52821, n52822, n52823, n52824, n52825, n52826,
    n52827, n52828, n52829, n52830, n52831, n52832, n52833, n52834, n52835,
    n52836, n52837, n52838, n52839, n52840, n52841, n52842, n52843, n52844,
    n52845, n52846, n52847, n52848, n52849, n52850, n52851, n52852, n52853,
    n52854, n52855, n52856, n52857, n52858, n52859, n52860, n52861, n52862,
    n52863, n52864, n52865, n52866, n52867, n52868, n52869, n52870, n52871,
    n52872, n52873, n52874, n52875, n52876, n52877, n52878, n52879, n52880,
    n52881, n52882, n52883, n52884, n52885, n52886, n52887, n52888, n52889,
    n52890, n52891, n52892, n52893, n52894, n52895, n52896, n52897, n52898,
    n52899, n52900, n52901, n52902, n52903, n52904, n52905, n52906, n52907,
    n52908, n52909, n52910, n52911, n52912, n52913, n52914, n52915, n52916,
    n52917, n52918, n52919, n52920, n52921, n52922, n52923, n52924, n52925,
    n52926, n52927, n52928, n52929, n52930, n52931, n52932, n52933, n52934,
    n52935, n52936, n52937, n52938, n52939, n52940, n52941, n52942, n52943,
    n52944, n52945, n52946, n52947, n52948, n52949, n52950, n52951, n52952,
    n52953, n52954, n52955, n52956, n52957, n52958, n52959, n52960, n52961,
    n52962, n52963, n52964, n52965, n52966, n52967, n52968, n52969, n52970,
    n52971, n52972, n52973, n52974, n52975, n52976, n52977, n52978, n52979,
    n52980, n52981, n52982, n52983, n52984, n52985, n52986, n52987, n52988,
    n52989, n52990, n52991, n52992, n52993, n52994, n52995, n52996, n52997,
    n52998, n52999, n53000, n53001, n53002, n53003, n53004, n53005, n53006,
    n53007, n53008, n53009, n53010, n53011, n53012, n53013, n53014, n53015,
    n53016, n53017, n53018, n53019, n53020, n53021, n53022, n53023, n53024,
    n53025, n53026, n53027, n53028, n53029, n53030, n53031, n53032, n53033,
    n53034, n53035, n53036, n53037, n53038, n53039, n53040, n53041, n53042,
    n53043, n53044, n53045, n53046, n53047, n53048, n53049, n53050, n53051,
    n53052, n53053, n53054, n53055, n53056, n53057, n53058, n53059, n53060,
    n53061, n53062, n53063, n53064, n53065, n53066, n53067, n53068, n53069,
    n53070, n53071, n53072, n53073, n53074, n53075, n53076, n53077, n53078,
    n53079, n53080, n53081, n53082, n53083, n53084, n53085, n53086, n53087,
    n53088, n53089, n53090, n53091, n53092, n53093, n53094, n53095, n53096,
    n53097, n53098, n53099, n53100, n53101, n53102, n53103, n53104, n53105,
    n53106, n53107, n53108, n53109, n53110, n53111, n53112, n53113, n53114,
    n53115, n53116, n53117, n53118, n53119, n53120, n53121, n53122, n53123,
    n53124, n53125, n53126, n53127, n53128, n53129, n53130, n53131, n53132,
    n53133, n53134, n53135, n53136, n53137, n53138, n53139, n53140, n53141,
    n53142, n53143, n53144, n53145, n53146, n53147, n53148, n53149, n53150,
    n53151, n53152, n53153, n53154, n53155, n53156, n53157, n53158, n53159,
    n53160, n53161, n53162, n53163, n53164, n53165, n53166, n53167, n53168,
    n53169, n53170, n53171, n53172, n53173, n53174, n53175, n53176, n53177,
    n53178, n53179, n53180, n53181, n53182, n53183, n53184, n53185, n53186,
    n53187, n53188, n53189, n53190, n53191, n53192, n53193, n53194, n53195,
    n53196, n53197, n53198, n53199, n53200, n53201, n53202, n53203, n53204,
    n53205, n53206, n53207, n53208, n53209, n53210, n53211, n53212, n53213,
    n53214, n53215, n53216, n53217, n53218, n53219, n53220, n53221, n53222,
    n53223, n53224, n53225, n53226, n53227, n53228, n53229, n53230, n53231,
    n53232, n53233, n53234, n53235, n53236, n53237, n53238, n53239, n53240,
    n53241, n53242, n53243, n53244, n53245, n53246, n53247, n53248, n53249,
    n53250, n53251, n53252, n53253, n53254, n53255, n53256, n53257, n53258,
    n53259, n53260, n53261, n53262, n53263, n53264, n53265, n53266, n53267,
    n53268, n53269, n53270, n53271, n53272, n53273, n53274, n53275, n53276,
    n53277, n53278, n53279, n53280, n53281, n53282, n53283, n53284, n53285,
    n53286, n53287, n53288, n53289, n53290, n53291, n53292, n53293, n53294,
    n53295, n53296, n53297, n53298, n53299, n53300, n53301, n53302, n53303,
    n53304, n53305, n53306, n53307, n53308, n53309, n53310, n53311, n53312,
    n53313, n53314, n53315, n53316, n53317, n53318, n53319, n53320, n53321,
    n53322, n53323, n53324, n53325, n53326, n53327, n53328, n53329, n53330,
    n53331, n53332, n53333, n53334, n53335, n53336, n53337, n53338, n53339,
    n53340, n53341, n53342, n53343, n53344, n53345, n53346, n53347, n53348,
    n53349, n53350, n53351, n53352, n53353, n53354, n53355, n53356, n53357,
    n53358, n53359, n53360, n53361, n53362, n53363, n53364, n53365, n53366,
    n53367, n53368, n53369, n53370, n53371, n53372, n53373, n53374, n53375,
    n53376, n53377, n53378, n53379, n53380, n53381, n53382, n53383, n53384,
    n53385, n53386, n53387, n53388, n53389, n53390, n53391, n53392, n53393,
    n53394, n53395, n53396, n53397, n53398, n53399, n53400, n53401, n53402,
    n53403, n53404, n53405, n53406, n53407, n53408, n53409, n53410, n53411,
    n53412, n53413, n53414, n53415, n53416, n53417, n53418, n53419, n53420,
    n53421, n53422, n53423, n53424, n53425, n53426, n53427, n53428, n53429,
    n53430, n53431, n53432, n53433, n53434, n53435, n53436, n53437, n53438,
    n53439, n53440, n53441, n53442, n53443, n53444, n53445, n53446, n53447,
    n53448, n53449, n53450, n53451, n53452, n53453, n53454, n53455, n53456,
    n53457, n53458, n53459, n53460, n53461, n53462, n53463, n53464, n53465,
    n53466, n53467, n53468, n53469, n53470, n53471, n53472, n53473, n53474,
    n53475, n53476, n53477, n53478, n53479, n53480, n53481, n53482, n53483,
    n53484, n53485, n53486, n53487, n53488, n53489, n53490, n53491, n53492,
    n53493, n53494, n53495, n53496, n53497, n53498, n53499, n53500, n53501,
    n53502, n53503, n53504, n53505, n53506, n53507, n53508, n53509, n53510,
    n53511, n53512, n53513, n53514, n53515, n53516, n53517, n53518, n53519,
    n53520, n53521, n53522, n53523, n53524, n53525, n53526, n53527, n53528,
    n53529, n53530, n53531, n53532, n53533, n53534, n53535, n53536, n53537,
    n53538, n53539, n53540, n53541, n53542, n53543, n53544, n53545, n53546,
    n53547, n53548, n53549, n53550, n53551, n53552, n53553, n53554, n53555,
    n53556, n53557, n53558, n53559, n53560, n53561, n53562, n53563, n53564,
    n53565, n53566, n53567, n53568, n53569, n53570, n53571, n53572, n53573,
    n53574, n53575, n53576, n53577, n53578, n53579, n53580, n53581, n53582,
    n53583, n53584, n53585, n53586, n53587, n53588, n53589, n53590, n53591,
    n53592, n53593, n53594, n53595, n53596, n53597, n53598, n53599, n53600,
    n53601, n53602, n53603, n53604, n53605, n53606, n53607, n53608, n53609,
    n53610, n53611, n53612, n53613, n53614, n53615, n53616, n53617, n53618,
    n53619, n53620, n53621, n53622, n53623, n53624, n53625, n53626, n53627,
    n53628, n53629, n53630, n53631, n53632, n53633, n53634, n53635, n53636,
    n53637, n53638, n53639, n53640, n53641, n53642, n53643, n53644, n53645,
    n53646, n53647, n53648, n53649, n53650, n53651, n53652, n53653, n53654,
    n53655, n53656, n53657, n53658, n53659, n53660, n53661, n53662, n53663,
    n53664, n53665, n53666, n53667, n53668, n53669, n53670, n53671, n53672,
    n53673, n53674, n53675, n53676, n53677, n53678, n53679, n53680, n53681,
    n53682, n53683, n53684, n53685, n53686, n53687, n53688, n53689, n53690,
    n53691, n53692, n53693, n53694, n53695, n53696, n53697, n53698, n53699,
    n53700, n53701, n53702, n53703, n53704, n53705, n53706, n53707, n53708,
    n53709, n53710, n53711, n53712, n53713, n53714, n53715, n53716, n53717,
    n53718, n53719, n53720, n53721, n53722, n53723, n53724, n53725, n53726,
    n53727, n53728, n53729, n53730, n53731, n53732, n53733, n53734, n53735,
    n53736, n53737, n53738, n53739, n53740, n53741, n53742, n53743, n53744,
    n53745, n53746, n53747, n53748, n53749, n53750, n53751, n53752, n53753,
    n53754, n53755, n53756, n53757, n53758, n53759, n53760, n53761, n53762,
    n53763, n53764, n53765, n53766, n53767, n53768, n53769, n53770, n53771,
    n53772, n53773, n53774, n53775, n53776, n53777, n53778, n53779, n53780,
    n53781, n53782, n53783, n53784, n53785, n53786, n53787, n53788, n53789,
    n53790, n53791, n53792, n53793, n53794, n53795, n53796, n53797, n53798,
    n53799, n53800, n53801, n53802, n53803, n53804, n53805, n53806, n53807,
    n53808, n53809, n53810, n53811, n53812, n53813, n53814, n53815, n53816,
    n53817, n53818, n53819, n53820, n53821, n53822, n53823, n53824, n53825,
    n53826, n53827, n53828, n53829, n53830, n53831, n53832, n53833, n53834,
    n53835, n53836, n53837, n53838, n53839, n53840, n53841, n53842, n53843,
    n53844, n53845, n53846, n53847, n53848, n53849, n53850, n53851, n53852,
    n53853, n53854, n53855, n53856, n53857, n53858, n53859, n53860, n53861,
    n53862, n53863, n53864, n53865, n53866, n53867, n53868, n53869, n53870,
    n53871, n53872, n53873, n53874, n53875, n53876, n53877, n53878, n53879,
    n53880, n53881, n53882, n53883, n53884, n53885, n53886, n53887, n53888,
    n53889, n53890, n53891, n53892, n53893, n53894, n53895, n53896, n53897,
    n53898, n53899, n53900, n53901, n53902, n53903, n53904, n53905, n53906,
    n53907, n53908, n53909, n53910, n53911, n53912, n53913, n53914, n53915,
    n53916, n53917, n53918, n53919, n53920, n53921, n53922, n53923, n53924,
    n53925, n53926, n53927, n53928, n53929, n53930, n53931, n53932, n53933,
    n53934, n53935, n53936, n53937, n53938, n53939, n53940, n53941, n53942,
    n53943, n53944, n53945, n53946, n53947, n53948, n53949, n53950, n53951,
    n53952, n53953, n53954, n53955, n53956, n53957, n53958, n53959, n53960,
    n53961, n53962, n53963, n53964, n53965, n53966, n53967, n53968, n53969,
    n53970, n53971, n53972, n53973, n53974, n53975, n53976, n53977, n53978,
    n53979, n53980, n53981, n53982, n53983, n53984, n53985, n53986, n53987,
    n53988, n53989, n53990, n53991, n53992, n53993, n53994, n53995, n53996,
    n53997, n53998, n53999, n54000, n54001, n54002, n54003, n54004, n54005,
    n54006, n54007, n54008, n54009, n54010, n54011, n54012, n54013, n54014,
    n54015, n54016, n54017, n54018, n54019, n54020, n54021, n54022, n54023,
    n54024, n54025, n54026, n54027, n54028, n54029, n54030, n54031, n54032,
    n54033, n54034, n54035, n54036, n54037, n54038, n54039, n54040, n54041,
    n54042, n54043, n54044, n54045, n54046, n54047, n54048, n54049, n54050,
    n54051, n54052, n54053, n54054, n54055, n54056, n54057, n54058, n54059,
    n54060, n54061, n54062, n54063, n54064, n54065, n54066, n54067, n54068,
    n54069, n54070, n54071, n54072, n54073, n54074, n54075, n54076, n54077,
    n54078, n54079, n54080, n54081, n54082, n54083, n54084, n54085, n54086,
    n54087, n54088, n54089, n54090, n54091, n54092, n54093, n54094, n54095,
    n54096, n54097, n54098, n54099, n54100, n54101, n54102, n54103, n54104,
    n54105, n54106, n54107, n54108, n54109, n54110, n54111, n54112, n54113,
    n54114, n54115, n54116, n54117, n54118, n54119, n54120, n54121, n54122,
    n54123, n54124, n54125, n54126, n54127, n54128, n54129, n54130, n54131,
    n54132, n54133, n54134, n54135, n54136, n54137, n54138, n54139, n54140,
    n54141, n54142, n54143, n54144, n54145, n54146, n54147, n54148, n54149,
    n54150, n54151, n54152, n54153, n54154, n54155, n54156, n54157, n54158,
    n54159, n54160, n54161, n54162, n54163, n54164, n54165, n54166, n54167,
    n54168, n54169, n54170, n54171, n54172, n54173, n54174, n54175, n54176,
    n54177, n54178, n54179, n54180, n54181, n54182, n54183, n54184, n54185,
    n54186, n54187, n54188, n54189, n54190, n54191, n54192, n54193, n54194,
    n54195, n54196, n54197, n54198, n54199, n54200, n54201, n54202, n54203,
    n54204, n54205, n54206, n54207, n54208, n54209, n54210, n54211, n54212,
    n54213, n54214, n54215, n54216, n54217, n54218, n54219, n54220, n54221,
    n54222, n54223, n54224, n54225, n54226, n54227, n54228, n54229, n54230,
    n54231, n54232, n54233, n54234, n54235, n54236, n54237, n54238, n54239,
    n54240, n54241, n54242, n54243, n54244, n54245, n54246, n54247, n54248,
    n54249, n54250, n54251, n54252, n54253, n54254, n54255, n54256, n54257,
    n54258, n54259, n54260, n54261, n54262, n54263, n54264, n54265, n54266,
    n54267, n54268, n54269, n54270, n54271, n54272, n54273, n54274, n54275,
    n54276, n54277, n54278, n54279, n54280, n54281, n54282, n54283, n54284,
    n54285, n54286, n54287, n54288, n54289, n54290, n54291, n54292, n54293,
    n54294, n54295, n54296, n54297, n54298, n54299, n54300, n54301, n54302,
    n54303, n54304, n54305, n54306, n54307, n54308, n54309, n54310, n54311,
    n54312, n54313, n54314, n54315, n54316, n54317, n54318, n54319, n54320,
    n54321, n54322, n54323, n54324, n54325, n54326, n54327, n54328, n54329,
    n54330, n54331, n54332, n54333, n54334, n54335, n54336, n54337, n54338,
    n54339, n54340, n54341, n54342, n54343, n54344, n54345, n54346, n54347,
    n54348, n54349, n54350, n54351, n54352, n54353, n54354, n54355, n54356,
    n54357, n54358, n54359, n54360, n54361, n54362, n54363, n54364, n54365,
    n54366, n54367, n54368, n54369, n54370, n54371, n54372, n54373, n54374,
    n54375, n54376, n54377, n54378, n54379, n54380, n54381, n54382, n54383,
    n54384, n54385, n54386, n54387, n54388, n54389, n54390, n54391, n54392,
    n54393, n54394, n54395, n54396, n54397, n54398, n54399, n54400, n54401,
    n54402, n54403, n54404, n54405, n54406, n54407, n54408, n54409, n54410,
    n54411, n54412, n54413, n54414, n54415, n54416, n54417, n54418, n54419,
    n54420, n54421, n54422, n54423, n54424, n54425, n54426, n54427, n54428,
    n54429, n54430, n54431, n54432, n54433, n54434, n54435, n54436, n54437,
    n54438, n54439, n54440, n54441, n54442, n54443, n54444, n54445, n54446,
    n54447, n54448, n54449, n54450, n54451, n54452, n54453, n54454, n54455,
    n54456, n54457, n54458, n54459, n54460, n54461, n54462, n54463, n54464,
    n54465, n54466, n54467, n54468, n54469, n54470, n54471, n54472, n54473,
    n54474, n54475, n54476, n54477, n54478, n54479, n54480, n54481, n54482,
    n54483, n54484, n54485, n54486, n54487, n54488, n54489, n54490, n54491,
    n54492, n54493, n54494, n54495, n54496, n54497, n54498, n54499, n54500,
    n54501, n54502, n54503, n54504, n54505, n54506, n54507, n54508, n54509,
    n54510, n54511, n54512, n54513, n54514, n54515, n54516, n54517, n54518,
    n54519, n54520, n54521, n54522, n54523, n54524, n54525, n54526, n54527,
    n54528, n54529, n54530, n54531, n54532, n54533, n54534, n54535, n54536,
    n54537, n54538, n54539, n54540, n54541, n54542, n54543, n54544, n54545,
    n54546, n54547, n54548, n54549, n54550, n54551, n54552, n54553, n54554,
    n54555, n54556, n54557, n54558, n54559, n54560, n54561, n54562, n54563,
    n54564, n54565, n54566, n54567, n54568, n54569, n54570, n54571, n54572,
    n54573, n54574, n54575, n54576, n54577, n54578, n54579, n54580, n54581,
    n54582, n54583, n54584, n54585, n54586, n54587, n54588, n54589, n54590,
    n54591, n54592, n54593, n54594, n54595, n54596, n54597, n54598, n54599,
    n54600, n54601, n54602, n54603, n54604, n54605, n54606, n54607, n54608,
    n54609, n54610, n54611, n54612, n54613, n54614, n54615, n54616, n54617,
    n54618, n54619, n54620, n54621, n54622, n54623, n54624, n54625, n54626,
    n54627, n54628, n54629, n54630, n54631, n54632, n54633, n54634, n54635,
    n54636, n54637, n54638, n54639, n54640, n54641, n54642, n54643, n54644,
    n54645, n54646, n54647, n54648, n54649, n54650, n54651, n54652, n54653,
    n54654, n54655, n54656, n54657, n54658, n54659, n54660, n54661, n54662,
    n54663, n54664, n54665, n54666, n54667, n54668, n54669, n54670, n54671,
    n54672, n54673, n54674, n54675, n54676, n54677, n54678, n54679, n54680,
    n54681, n54682, n54683, n54684, n54685, n54686, n54687, n54688, n54689,
    n54690, n54691, n54692, n54693, n54694, n54695, n54696, n54697, n54698,
    n54699, n54700, n54701, n54702, n54703, n54704, n54705, n54706, n54707,
    n54708, n54709, n54710, n54711, n54712, n54713, n54714, n54715, n54716,
    n54717, n54718, n54719, n54720, n54721, n54722, n54723, n54724, n54725,
    n54726, n54727, n54728, n54729, n54730, n54731, n54732, n54733, n54734,
    n54735, n54736, n54737, n54738, n54739, n54740, n54741, n54742, n54743,
    n54744, n54745, n54746, n54747, n54748, n54749, n54750, n54751, n54752,
    n54753, n54754, n54755, n54756, n54757, n54758, n54759, n54760, n54761,
    n54762, n54763, n54764, n54765, n54766, n54767, n54768, n54769, n54770,
    n54771, n54772, n54773, n54774, n54775, n54776, n54777, n54778, n54779,
    n54780, n54781, n54782, n54783, n54784, n54785, n54786, n54787, n54788,
    n54789, n54790, n54791, n54792, n54793, n54794, n54795, n54796, n54797,
    n54798, n54799, n54800, n54801, n54802, n54803, n54804, n54805, n54806,
    n54807, n54808, n54809, n54810, n54811, n54812, n54813, n54814, n54815,
    n54816, n54817, n54818, n54819, n54820, n54821, n54822, n54823, n54824,
    n54825, n54826, n54827, n54828, n54829, n54830, n54831, n54832, n54833,
    n54834, n54835, n54836, n54837, n54838, n54839, n54840, n54841, n54842,
    n54843, n54844, n54845, n54846, n54847, n54848, n54849, n54850, n54851,
    n54852, n54853, n54854, n54855, n54856, n54857, n54858, n54859, n54860,
    n54861, n54862, n54863, n54864, n54865, n54866, n54867, n54868, n54869,
    n54870, n54871, n54872, n54873, n54874, n54875, n54876, n54877, n54878,
    n54879, n54880, n54881, n54882, n54883, n54884, n54885, n54886, n54887,
    n54888, n54889, n54890, n54891, n54892, n54893, n54894, n54895, n54896,
    n54897, n54898, n54899, n54900, n54901, n54902, n54903, n54904, n54905,
    n54906, n54907, n54908, n54909, n54910, n54911, n54912, n54913, n54914,
    n54915, n54916, n54917, n54918, n54919, n54920, n54921, n54922, n54923,
    n54924, n54925, n54926, n54927, n54928, n54929, n54930, n54931, n54932,
    n54933, n54934, n54935, n54936, n54937, n54938, n54939, n54940, n54941,
    n54942, n54943, n54944, n54945, n54946, n54947, n54948, n54949, n54950,
    n54951, n54952, n54953, n54954, n54955, n54956, n54957, n54958, n54959,
    n54960, n54961, n54962, n54963, n54964, n54965, n54966, n54967, n54968,
    n54969, n54970, n54971, n54972, n54973, n54974, n54975, n54976, n54977,
    n54978, n54979, n54980, n54981, n54982, n54983, n54984, n54985, n54986,
    n54987, n54988, n54989, n54990, n54991, n54992, n54993, n54994, n54995,
    n54996, n54997, n54998, n54999, n55000, n55001, n55002, n55003, n55004,
    n55005, n55006, n55007, n55008, n55009, n55010, n55011, n55012, n55013,
    n55014, n55015, n55016, n55017, n55018, n55019, n55020, n55021, n55022,
    n55023, n55024, n55025, n55026, n55027, n55028, n55029, n55030, n55031,
    n55032, n55033, n55034, n55035, n55036, n55037, n55038, n55039, n55040,
    n55041, n55042, n55043, n55044, n55045, n55046, n55047, n55048, n55049,
    n55050, n55051, n55052, n55053, n55054, n55055, n55056, n55057, n55058,
    n55059, n55060, n55061, n55062, n55063, n55064, n55065, n55066, n55067,
    n55068, n55069, n55070, n55071, n55072, n55073, n55074, n55075, n55076,
    n55077, n55078, n55079, n55080, n55081, n55082, n55083, n55084, n55085,
    n55086, n55087, n55088, n55089, n55090, n55091, n55092, n55093, n55094,
    n55095, n55096, n55097, n55098, n55099, n55100, n55101, n55102, n55103,
    n55104, n55105, n55106, n55107, n55108, n55109, n55110, n55111, n55112,
    n55113, n55114, n55115, n55116, n55117, n55118, n55119, n55120, n55121,
    n55122, n55123, n55124, n55125, n55126, n55127, n55128, n55129, n55130,
    n55131, n55132, n55133, n55134, n55135, n55136, n55137, n55138, n55139,
    n55140, n55141, n55142, n55143, n55144, n55145, n55146, n55147, n55148,
    n55149, n55150, n55151, n55152, n55153, n55154, n55155, n55156, n55157,
    n55158, n55159, n55160, n55161, n55162, n55163, n55164, n55165, n55166,
    n55167, n55168, n55169, n55170, n55171, n55172, n55173, n55174, n55175,
    n55176, n55177, n55178, n55179, n55180, n55181, n55182, n55183, n55184,
    n55185, n55186, n55187, n55188, n55189, n55190, n55191, n55192, n55193,
    n55194, n55195, n55196, n55197, n55198, n55199, n55200, n55201, n55202,
    n55203, n55204, n55205, n55206, n55207, n55208, n55209, n55210, n55211,
    n55212, n55213, n55214, n55215, n55216, n55217, n55218, n55219, n55220,
    n55221, n55222, n55223, n55224, n55225, n55226, n55227, n55228, n55229,
    n55230, n55231, n55232, n55233, n55234, n55235, n55236, n55237, n55238,
    n55239, n55240, n55241, n55242, n55243, n55244, n55245, n55246, n55247,
    n55248, n55249, n55250, n55251, n55252, n55253, n55254, n55255, n55256,
    n55257, n55258, n55259, n55260, n55261, n55262, n55263, n55264, n55265,
    n55266, n55267, n55268, n55269, n55270, n55271, n55272, n55273, n55274,
    n55275, n55276, n55277, n55278, n55279, n55280, n55281, n55282, n55283,
    n55284, n55285, n55286, n55287, n55288, n55289, n55290, n55291, n55292,
    n55293, n55294, n55295, n55296, n55297, n55298, n55299, n55300, n55301,
    n55302, n55303, n55304, n55305, n55306, n55307, n55308, n55309, n55310,
    n55311, n55312, n55313, n55314, n55315, n55316, n55317, n55318, n55319,
    n55320, n55321, n55322, n55323, n55324, n55325, n55326, n55327, n55328,
    n55329, n55330, n55331, n55332, n55333, n55334, n55335, n55336, n55337,
    n55338, n55339, n55340, n55341, n55342, n55343, n55344, n55345, n55346,
    n55347, n55348, n55349, n55350, n55351, n55352, n55353, n55354, n55355,
    n55356, n55357, n55358, n55359, n55360, n55361, n55362, n55363, n55364,
    n55365, n55366, n55367, n55368, n55369, n55370, n55371, n55372, n55373,
    n55374, n55375, n55376, n55377, n55378, n55379, n55380, n55381, n55382,
    n55383, n55384, n55385, n55386, n55387, n55388, n55389, n55390, n55391,
    n55392, n55393, n55394, n55395, n55396, n55397, n55398, n55399, n55400,
    n55401, n55402, n55403, n55404, n55405, n55406, n55407, n55408, n55409,
    n55410, n55411, n55412, n55413, n55414, n55415, n55416, n55417, n55418,
    n55419, n55420, n55421, n55422, n55423, n55424, n55425, n55426, n55427,
    n55428, n55429, n55430, n55431, n55432, n55433, n55434, n55435, n55436,
    n55437, n55438, n55439, n55440, n55441, n55442, n55443, n55444, n55445,
    n55446, n55447, n55448, n55449, n55450, n55451, n55452, n55453, n55454,
    n55455, n55456, n55457, n55458, n55459, n55460, n55461, n55462, n55463,
    n55464, n55465, n55466, n55467, n55468, n55469, n55470, n55471, n55472,
    n55473, n55474, n55475, n55476, n55477, n55478, n55479, n55480, n55481,
    n55482, n55483, n55484, n55485, n55486, n55487, n55488, n55489, n55490,
    n55491, n55492, n55493, n55494, n55495, n55496, n55497, n55498, n55499,
    n55500, n55501, n55502, n55503, n55504, n55505, n55506, n55507, n55508,
    n55509, n55510, n55511, n55512, n55513, n55514, n55515, n55516, n55517,
    n55518, n55519, n55520, n55521, n55522, n55523, n55524, n55525, n55526,
    n55527, n55528, n55529, n55530, n55531, n55532, n55533, n55534, n55535,
    n55536, n55537, n55538, n55539, n55540, n55541, n55542, n55543, n55544,
    n55545, n55546, n55547, n55548, n55549, n55550, n55551, n55552, n55553,
    n55554, n55555, n55556, n55557, n55558, n55559, n55560, n55561, n55562,
    n55563, n55564, n55565, n55566, n55567, n55568, n55569, n55570, n55571,
    n55572, n55573, n55574, n55575, n55576, n55577, n55578, n55579, n55580,
    n55581, n55582, n55583, n55584, n55585, n55586, n55587, n55588, n55589,
    n55590, n55591, n55592, n55593, n55594, n55595, n55596, n55597, n55598,
    n55599, n55600, n55601, n55602, n55603, n55604, n55605, n55606, n55607,
    n55608, n55609, n55610, n55611, n55612, n55613, n55614, n55615, n55616,
    n55617, n55618, n55619, n55620, n55621, n55622, n55623, n55624, n55625,
    n55626, n55627, n55628, n55629, n55630, n55631, n55632, n55633, n55634,
    n55635, n55636, n55637, n55638, n55639, n55640, n55641, n55642, n55643,
    n55644, n55645, n55646, n55647, n55648, n55649, n55650, n55651, n55652,
    n55653, n55654, n55655, n55656, n55657, n55658, n55659, n55660, n55661,
    n55662, n55663, n55664, n55665, n55666, n55667, n55668, n55669, n55670,
    n55671, n55672, n55673, n55674, n55675, n55676, n55677, n55678, n55679,
    n55680, n55681, n55682, n55683, n55684, n55685, n55686, n55687, n55688,
    n55689, n55690, n55691, n55692, n55693, n55694, n55695, n55696, n55697,
    n55698, n55699, n55700, n55701, n55702, n55703, n55704, n55705, n55706,
    n55707, n55708, n55709, n55710, n55711, n55712, n55713, n55714, n55715,
    n55716, n55717, n55718, n55719, n55720, n55721, n55722, n55723, n55724,
    n55725, n55726, n55727, n55728, n55729, n55730, n55731, n55732, n55733,
    n55734, n55735, n55736, n55737, n55738, n55739, n55740, n55741, n55742,
    n55743, n55744, n55745, n55746, n55747, n55748, n55749, n55750, n55751,
    n55752, n55753, n55754, n55755, n55756, n55757, n55758, n55759, n55760,
    n55761, n55762, n55763, n55764, n55765, n55766, n55767, n55768, n55769,
    n55770, n55771, n55772, n55773, n55774, n55775, n55776, n55777, n55778,
    n55779, n55780, n55781, n55782, n55783, n55784, n55785, n55786, n55787,
    n55788, n55789, n55790, n55791, n55792, n55793, n55794, n55795, n55796,
    n55797, n55798, n55799, n55800, n55801, n55802, n55803, n55804, n55805,
    n55806, n55807, n55808, n55809, n55810, n55811, n55812, n55813, n55814,
    n55815, n55816, n55817, n55818, n55819, n55820, n55821, n55822, n55823,
    n55824, n55825, n55826, n55827, n55828, n55829, n55830, n55831, n55832,
    n55833, n55834, n55835, n55836, n55837, n55838, n55839, n55840, n55841,
    n55842, n55843, n55844, n55845, n55846, n55847, n55848, n55849, n55850,
    n55851, n55852, n55853, n55854, n55855, n55856, n55857, n55858, n55859,
    n55860, n55861, n55862, n55863, n55864, n55865, n55866, n55867, n55868,
    n55869, n55870, n55871, n55872, n55873, n55874, n55875, n55876, n55877,
    n55878, n55879, n55880, n55881, n55882, n55883, n55884, n55885, n55886,
    n55887, n55888, n55889, n55890, n55891, n55892, n55893, n55894, n55895,
    n55896, n55897, n55898, n55899, n55900, n55901, n55902, n55903, n55904,
    n55905, n55906, n55907, n55908, n55909, n55910, n55911, n55912, n55913,
    n55914, n55915, n55916, n55917, n55918, n55919, n55920, n55921, n55922,
    n55923, n55924, n55925, n55926, n55927, n55928, n55929, n55930, n55931,
    n55932, n55933, n55934, n55935, n55936, n55937, n55938, n55939, n55940,
    n55941, n55942, n55943, n55944, n55945, n55946, n55947, n55948, n55949,
    n55950, n55951, n55952, n55953, n55954, n55955, n55956, n55957, n55958,
    n55959, n55960, n55961, n55962, n55963, n55964, n55965, n55966, n55967,
    n55968, n55969, n55970, n55971, n55972, n55973, n55974, n55975, n55976,
    n55977, n55978, n55979, n55980, n55981, n55982, n55983, n55984, n55985,
    n55986, n55987, n55988, n55989, n55990, n55991, n55992, n55993, n55994,
    n55995, n55996, n55997, n55998, n55999, n56000, n56001, n56002, n56003,
    n56004, n56005, n56006, n56007, n56008, n56009, n56010, n56011, n56012,
    n56013, n56014, n56015, n56016, n56017, n56018, n56019, n56020, n56021,
    n56022, n56023, n56024, n56025, n56026, n56027, n56028, n56029, n56030,
    n56031, n56032, n56033, n56034, n56035, n56036, n56037, n56038, n56039,
    n56040, n56041, n56042, n56043, n56044, n56045, n56046, n56047, n56048,
    n56049, n56050, n56051, n56052, n56053, n56054, n56055, n56056, n56057,
    n56058, n56059, n56060, n56061, n56062, n56063, n56064, n56065, n56066,
    n56067, n56068, n56069, n56070, n56071, n56072, n56073, n56074, n56075,
    n56076, n56077, n56078, n56079, n56080, n56081, n56082, n56083, n56084,
    n56085, n56086, n56087, n56088, n56089, n56090, n56091, n56092, n56093,
    n56094, n56095, n56096, n56097, n56098, n56099, n56100, n56101, n56102,
    n56103, n56104, n56105, n56106, n56107, n56108, n56109, n56110, n56111,
    n56112, n56113, n56114, n56115, n56116, n56117, n56118, n56119, n56120,
    n56121, n56122, n56123, n56124, n56125, n56126, n56127, n56128, n56129,
    n56130, n56131, n56132, n56133, n56134, n56135, n56136, n56137, n56138,
    n56139, n56140, n56141, n56142, n56143, n56144, n56145, n56146, n56147,
    n56148, n56149, n56150, n56151, n56152, n56153, n56154, n56155, n56156,
    n56157, n56158, n56159, n56160, n56161, n56162, n56163, n56164, n56165,
    n56166, n56167, n56168, n56169, n56170, n56171, n56172, n56173, n56174,
    n56175, n56176, n56177, n56178, n56179, n56180, n56181, n56182, n56183,
    n56184, n56185, n56186, n56187, n56188, n56189, n56190, n56191, n56192,
    n56193, n56194, n56195, n56196, n56197, n56198, n56199, n56200, n56201,
    n56202, n56203, n56204, n56205, n56206, n56207, n56208, n56209, n56210,
    n56211, n56212, n56213, n56214, n56215, n56216, n56217, n56218, n56219,
    n56220, n56221, n56222, n56223, n56224, n56225, n56226, n56227, n56228,
    n56229, n56230, n56231, n56232, n56233, n56234, n56235, n56236, n56237,
    n56238, n56239, n56240, n56241, n56242, n56243, n56244, n56245, n56246,
    n56247, n56248, n56249, n56250, n56251, n56252, n56253, n56254, n56255,
    n56256, n56257, n56258, n56259, n56260, n56261, n56262, n56263, n56264,
    n56265, n56266, n56267, n56268, n56269, n56270, n56271, n56272, n56273,
    n56274, n56275, n56276, n56277, n56278, n56279, n56280, n56281, n56282,
    n56283, n56284, n56285, n56286, n56287, n56288, n56289, n56290, n56291,
    n56292, n56293, n56294, n56295, n56296, n56297, n56298, n56299, n56300,
    n56301, n56302, n56303, n56304, n56305, n56306, n56307, n56308, n56309,
    n56310, n56311, n56312, n56313, n56314, n56315, n56316, n56317, n56318,
    n56319, n56320, n56321, n56322, n56323, n56324, n56325, n56326, n56327,
    n56328, n56329, n56330, n56331, n56332, n56333, n56334, n56335, n56336,
    n56337, n56338, n56339, n56340, n56341, n56342, n56343, n56344, n56345,
    n56346, n56347, n56348, n56349, n56350, n56351, n56352, n56353, n56354,
    n56355, n56356, n56357, n56358, n56359, n56360, n56361, n56362, n56363,
    n56364, n56365, n56366, n56367, n56368, n56369, n56370, n56371, n56372,
    n56373, n56374, n56375, n56376, n56377, n56378, n56379, n56380, n56381,
    n56382, n56383, n56384, n56385, n56386, n56387, n56388, n56389, n56390,
    n56391, n56392, n56393, n56394, n56395, n56396, n56397, n56398, n56399,
    n56400, n56401, n56402, n56403, n56404, n56405, n56406, n56407, n56408,
    n56409, n56410, n56411, n56412, n56413, n56414, n56415, n56416, n56417,
    n56418, n56419, n56420, n56421, n56422, n56423, n56424, n56425, n56426,
    n56427, n56428, n56429, n56430, n56431, n56432, n56433, n56434, n56435,
    n56436, n56437, n56438, n56439, n56440, n56441, n56442, n56443, n56444,
    n56445, n56446, n56447, n56448, n56449, n56450, n56451, n56452, n56453,
    n56454, n56455, n56456, n56457, n56458, n56459, n56460, n56461, n56462,
    n56463, n56464, n56465, n56466, n56467, n56468, n56469, n56470, n56471,
    n56472, n56473, n56474, n56475, n56476, n56477, n56478, n56479, n56480,
    n56481, n56482, n56483, n56484, n56485, n56486, n56487, n56488, n56489,
    n56490, n56491, n56492, n56493, n56494, n56495, n56496, n56497, n56498,
    n56499, n56500, n56501, n56502, n56503, n56504, n56505, n56506, n56507,
    n56508, n56509, n56510, n56511, n56512, n56513, n56514, n56515, n56516,
    n56517, n56518, n56519, n56520, n56521, n56522, n56523, n56524, n56525,
    n56526, n56527, n56528, n56529, n56530, n56531, n56532, n56533, n56534,
    n56535, n56536, n56537, n56538, n56539, n56540, n56541, n56542, n56543,
    n56544, n56545, n56546, n56547, n56548, n56549, n56550, n56551, n56552,
    n56553, n56554, n56555, n56556, n56557, n56558, n56559, n56560, n56561,
    n56562, n56563, n56564, n56565, n56566, n56567, n56568, n56569, n56570,
    n56571, n56572, n56573, n56574, n56575, n56576, n56577, n56578, n56579,
    n56580, n56581, n56582, n56583, n56584, n56585, n56586, n56587, n56588,
    n56589, n56590, n56591, n56592, n56593, n56594, n56595, n56596, n56597,
    n56598, n56599, n56600, n56601, n56602, n56603, n56604, n56605, n56606,
    n56607, n56608, n56609, n56610, n56611, n56612, n56613, n56614, n56615,
    n56616, n56617, n56618, n56619, n56620, n56621, n56622, n56623, n56624,
    n56625, n56626, n56627, n56628, n56629, n56630, n56631, n56632, n56633,
    n56634, n56635, n56636, n56637, n56638, n56639, n56640, n56641, n56642,
    n56643, n56644, n56645, n56646, n56647, n56648, n56649, n56650, n56651,
    n56652, n56653, n56654, n56655, n56656, n56657, n56658, n56659, n56660,
    n56661, n56662, n56663, n56664, n56665, n56666, n56667, n56668, n56669,
    n56670, n56671, n56672, n56673, n56674, n56675, n56676, n56677, n56678,
    n56679, n56680, n56681, n56682, n56683, n56684, n56685, n56686, n56687,
    n56688, n56689, n56690, n56691, n56692, n56693, n56694, n56695, n56696,
    n56697, n56698, n56699, n56700, n56701, n56702, n56703, n56704, n56705,
    n56706, n56707, n56708, n56709, n56710, n56711, n56712, n56713, n56714,
    n56715, n56716, n56717, n56718, n56719, n56720, n56721, n56722, n56723,
    n56724, n56725, n56726, n56727, n56728, n56729, n56730, n56731, n56732,
    n56733, n56734, n56735, n56736, n56737, n56738, n56739, n56740, n56741,
    n56742, n56743, n56744, n56745, n56746, n56747, n56748, n56749, n56750,
    n56751, n56752, n56753, n56754, n56755, n56756, n56757, n56758, n56759,
    n56760, n56761, n56762, n56763, n56764, n56765, n56766, n56767, n56768,
    n56769, n56770, n56771, n56772, n56773, n56774, n56775, n56776, n56777,
    n56778, n56779, n56780, n56781, n56782, n56783, n56784, n56785, n56786,
    n56787, n56788, n56789, n56790, n56791, n56792, n56793, n56794, n56795,
    n56796, n56797, n56798, n56799, n56800, n56801, n56802, n56803, n56804,
    n56805, n56806, n56807, n56808, n56809, n56810, n56811, n56812, n56813,
    n56814, n56815, n56816, n56817, n56818, n56819, n56820, n56821, n56822,
    n56823, n56824, n56825, n56826, n56827, n56828, n56829, n56830, n56831,
    n56832, n56833, n56834, n56835, n56836, n56837, n56838, n56839, n56840,
    n56841, n56842, n56843, n56844, n56845, n56846, n56847, n56848, n56849,
    n56850, n56851, n56852, n56853, n56854, n56855, n56856, n56857, n56858,
    n56859, n56860, n56861, n56862, n56863, n56864, n56865, n56866, n56867,
    n56868, n56869, n56870, n56871, n56872, n56873, n56874, n56875, n56876,
    n56877, n56878, n56879, n56880, n56881, n56882, n56883, n56884, n56885,
    n56886, n56887, n56888, n56889, n56890, n56891, n56892, n56893, n56894,
    n56895, n56896, n56897, n56898, n56899, n56900, n56901, n56902, n56903,
    n56904, n56905, n56906, n56907, n56908, n56909, n56910, n56911, n56912,
    n56913, n56914, n56915, n56916, n56917, n56918, n56919, n56920, n56921,
    n56922, n56923, n56924, n56925, n56926, n56927, n56928, n56929, n56930,
    n56931, n56932, n56933, n56934, n56935, n56936, n56937, n56938, n56939,
    n56940, n56941, n56942, n56943, n56944, n56945, n56946, n56947, n56948,
    n56949, n56950, n56951, n56952, n56953, n56954, n56955, n56956, n56957,
    n56958, n56959, n56960, n56961, n56962, n56963, n56964, n56965, n56966,
    n56967, n56968, n56969, n56970, n56971, n56972, n56973, n56974, n56975,
    n56976, n56977, n56978, n56979, n56980, n56981, n56982, n56983, n56984,
    n56985, n56986, n56987, n56988, n56989, n56990, n56991, n56992, n56993,
    n56994, n56995, n56996, n56997, n56998, n56999, n57000, n57001, n57002,
    n57003, n57004, n57005, n57006, n57007, n57008, n57009, n57010, n57011,
    n57012, n57013, n57014, n57015, n57016, n57017, n57018, n57019, n57020,
    n57021, n57022, n57023, n57024, n57025, n57026, n57027, n57028, n57029,
    n57030, n57031, n57032, n57033, n57034, n57035, n57036, n57037, n57038,
    n57039, n57040, n57041, n57042, n57043, n57044, n57045, n57046, n57047,
    n57048, n57049, n57050, n57051, n57052, n57053, n57054, n57055, n57056,
    n57057, n57058, n57059, n57060, n57061, n57062, n57063, n57064, n57065,
    n57066, n57067, n57068, n57069, n57070, n57071, n57072, n57073, n57074,
    n57075, n57076, n57077, n57078, n57079, n57080, n57081, n57082, n57083,
    n57084, n57085, n57086, n57087, n57088, n57089, n57090, n57091, n57092,
    n57093, n57094, n57095, n57096, n57097, n57098, n57099, n57100, n57101,
    n57102, n57103, n57104, n57105, n57106, n57107, n57108, n57109, n57110,
    n57111, n57112, n57113, n57114, n57115, n57116, n57117, n57118, n57119,
    n57120, n57121, n57122, n57123, n57124, n57125, n57126, n57127, n57128,
    n57129, n57130, n57131, n57132, n57133, n57134, n57135, n57136, n57137,
    n57138, n57139, n57140, n57141, n57142, n57143, n57144, n57145, n57146,
    n57147, n57148, n57149, n57150, n57151, n57152, n57153, n57154, n57155,
    n57156, n57157, n57158, n57159, n57160, n57161, n57162, n57163, n57164,
    n57165, n57166, n57167, n57168, n57169, n57170, n57171, n57172, n57173,
    n57174, n57175, n57176, n57177, n57178, n57179, n57180, n57181, n57182,
    n57183, n57184, n57185, n57186, n57187, n57188, n57189, n57190, n57191,
    n57192, n57193, n57194, n57195, n57196, n57197, n57198, n57199, n57200,
    n57201, n57202, n57203, n57204, n57205, n57206, n57207, n57208, n57209,
    n57210, n57211, n57212, n57213, n57214, n57215, n57216, n57217, n57218,
    n57219, n57220, n57221, n57222, n57223, n57224, n57225, n57226, n57227,
    n57228, n57229, n57230, n57231, n57232, n57233, n57234, n57235, n57236,
    n57237, n57238, n57239, n57240, n57241, n57242, n57243, n57244, n57245,
    n57246, n57247, n57248, n57249, n57250, n57251, n57252, n57253, n57254,
    n57255, n57256, n57257, n57258, n57259, n57260, n57261, n57262, n57263,
    n57264, n57265, n57266, n57267, n57268, n57269, n57270, n57271, n57272,
    n57273, n57274, n57275, n57276, n57277, n57278, n57279, n57280, n57281,
    n57282, n57283, n57284, n57285, n57286, n57287, n57288, n57289, n57290,
    n57291, n57292, n57293, n57294, n57295, n57296, n57297, n57298, n57299,
    n57300, n57301, n57302, n57303, n57304, n57305, n57306, n57307, n57308,
    n57309, n57310, n57311, n57312, n57313, n57314, n57315, n57316, n57317,
    n57318, n57319, n57320, n57321, n57322, n57323, n57324, n57325, n57326,
    n57327, n57328, n57329, n57330, n57331, n57332, n57333, n57334, n57335,
    n57336, n57337, n57338, n57339, n57340, n57341, n57342, n57343, n57344,
    n57345, n57346, n57347, n57348, n57349, n57350, n57351, n57352, n57353,
    n57354, n57355, n57356, n57357, n57358, n57359, n57360, n57361, n57362,
    n57363, n57364, n57365, n57366, n57367, n57368, n57369, n57370, n57371,
    n57372, n57373, n57374, n57375, n57376, n57377, n57378, n57379, n57380,
    n57381, n57382, n57383, n57384, n57385, n57386, n57387, n57388, n57389,
    n57390, n57391, n57392, n57393, n57394, n57395, n57396, n57397, n57398,
    n57399, n57400, n57401, n57402, n57403, n57404, n57405, n57406, n57407,
    n57408, n57409, n57410, n57411, n57412, n57413, n57414, n57415, n57416,
    n57417, n57418, n57419, n57420, n57421, n57422, n57423, n57424, n57425,
    n57426, n57427, n57428, n57429, n57430, n57431, n57432, n57433, n57434,
    n57435, n57436, n57437, n57438, n57439, n57440, n57441, n57442, n57443,
    n57444, n57445, n57446, n57447, n57448, n57449, n57450, n57451, n57452,
    n57453, n57454, n57455, n57456, n57457, n57458, n57459, n57460, n57461,
    n57462, n57463, n57464, n57465, n57466, n57467, n57468, n57469, n57470,
    n57471, n57472, n57473, n57474, n57475, n57476, n57477, n57478, n57479,
    n57480, n57481, n57482, n57483, n57484, n57485, n57486, n57487, n57488,
    n57489, n57490, n57491, n57492, n57493, n57494, n57495, n57496, n57497,
    n57498, n57499, n57500, n57501, n57502, n57503, n57504, n57505, n57506,
    n57507, n57508, n57509, n57510, n57511, n57512, n57513, n57514, n57515,
    n57516, n57517, n57518, n57519, n57520, n57521, n57522, n57523, n57524,
    n57525, n57526, n57527, n57528, n57529, n57530, n57531, n57532, n57533,
    n57534, n57535, n57536, n57537, n57538, n57539, n57540, n57541, n57542,
    n57543, n57544, n57545, n57546, n57547, n57548, n57549, n57550, n57551,
    n57552, n57553, n57554, n57555, n57556, n57557, n57558, n57559, n57560,
    n57561, n57562, n57563, n57564, n57565, n57566, n57567, n57568, n57569,
    n57570, n57571, n57572, n57573, n57574, n57575, n57576, n57577, n57578,
    n57579, n57580, n57581, n57582, n57583, n57584, n57585, n57586, n57587,
    n57588, n57589, n57590, n57591, n57592, n57593, n57594, n57595, n57596,
    n57597, n57598, n57599, n57600, n57601, n57602, n57603, n57604, n57605,
    n57606, n57607, n57608, n57609, n57610, n57611, n57612, n57613, n57614,
    n57615, n57616, n57617, n57618, n57619, n57620, n57621, n57622, n57623,
    n57624, n57625, n57626, n57627, n57628, n57629, n57630, n57631, n57632,
    n57633, n57634, n57635, n57636, n57637, n57638, n57639, n57640, n57641,
    n57642, n57643, n57644, n57645, n57646, n57647, n57648, n57649, n57650,
    n57651, n57652, n57653, n57654, n57655, n57656, n57657, n57658, n57659,
    n57660, n57661, n57662, n57663, n57664, n57665, n57666, n57667, n57668,
    n57669, n57670, n57671, n57672, n57673, n57674, n57675, n57676, n57677,
    n57678, n57679, n57680, n57681, n57682, n57683, n57684, n57685, n57686,
    n57687, n57688, n57689, n57690, n57691, n57692, n57693, n57694, n57695,
    n57696, n57697, n57698, n57699, n57700, n57701, n57702, n57703, n57704,
    n57705, n57706, n57707, n57708, n57709, n57710, n57711, n57712, n57713,
    n57714, n57715, n57716, n57717, n57718, n57719, n57720, n57721, n57722,
    n57723, n57724, n57725, n57726, n57727, n57728, n57729, n57730, n57731,
    n57732, n57733, n57734, n57735, n57736, n57737, n57738, n57739, n57740,
    n57741, n57742, n57743, n57744, n57745, n57746, n57747, n57748, n57749,
    n57750, n57751, n57752, n57753, n57754, n57755, n57756, n57757, n57758,
    n57759, n57760, n57761, n57762, n57763, n57764, n57765, n57766, n57767,
    n57768, n57769, n57770, n57771, n57772, n57773, n57774, n57775, n57776,
    n57777, n57778, n57779, n57780, n57781, n57782, n57783, n57784, n57785,
    n57786, n57787, n57788, n57789, n57790, n57791, n57792, n57793, n57794,
    n57795, n57796, n57797, n57798, n57799, n57800, n57801, n57802, n57803,
    n57804, n57805, n57806, n57807, n57808, n57809, n57810, n57811, n57812,
    n57813, n57814, n57815, n57816, n57817, n57818, n57819, n57820, n57821,
    n57822, n57823, n57824, n57825, n57826, n57827, n57828, n57829, n57830,
    n57831, n57832, n57833, n57834, n57835, n57836, n57837, n57838, n57839,
    n57840, n57841, n57842, n57843, n57844, n57845, n57846, n57847, n57848,
    n57849, n57850, n57851, n57852, n57853, n57854, n57855, n57856, n57857,
    n57858, n57859, n57860, n57861, n57862, n57863, n57864, n57865, n57866,
    n57867, n57868, n57869, n57870, n57871, n57872, n57873, n57874, n57875,
    n57876, n57877, n57878, n57879, n57880, n57881, n57882, n57883, n57884,
    n57885, n57886, n57887, n57888, n57889, n57890, n57891, n57892, n57893,
    n57894, n57895, n57896, n57897, n57898, n57899, n57900, n57901, n57902,
    n57903, n57904, n57905, n57906, n57907, n57908, n57909, n57910, n57911,
    n57912, n57913, n57914, n57915, n57916, n57917, n57918, n57919, n57920,
    n57921, n57922, n57923, n57924, n57925, n57926, n57927, n57928, n57929,
    n57930, n57931, n57932, n57933, n57934, n57935, n57936, n57937, n57938,
    n57939, n57940, n57941, n57942, n57943, n57944, n57945, n57946, n57947,
    n57948, n57949, n57950, n57951, n57952, n57953, n57954, n57955, n57956,
    n57957, n57958, n57959, n57960, n57961, n57962, n57963, n57964, n57965,
    n57966, n57967, n57968, n57969, n57970, n57971, n57972, n57973, n57974,
    n57975, n57976, n57977, n57978, n57979, n57980, n57981, n57982, n57983,
    n57984, n57985, n57986, n57987, n57988, n57989, n57990, n57991, n57992,
    n57993, n57994, n57995, n57996, n57997, n57998, n57999, n58000, n58001,
    n58002, n58003, n58004, n58005, n58006, n58007, n58008, n58009, n58010,
    n58011, n58012, n58013, n58014, n58015, n58016, n58017, n58018, n58019,
    n58020, n58021, n58022, n58023, n58024, n58025, n58026, n58027, n58028,
    n58029, n58030, n58031, n58032, n58033, n58034, n58035, n58036, n58037,
    n58038, n58039, n58040, n58041, n58042, n58043, n58044, n58045, n58046,
    n58047, n58048, n58049, n58050, n58051, n58052, n58053, n58054, n58055,
    n58056, n58057, n58058, n58059, n58060, n58061, n58062, n58063, n58064,
    n58065, n58066, n58067, n58068, n58069, n58070, n58071, n58072, n58073,
    n58074, n58075, n58076, n58077, n58078, n58079, n58080, n58081, n58082,
    n58083, n58084, n58085, n58086, n58087, n58088, n58089, n58090, n58091,
    n58092, n58093, n58094, n58095, n58096, n58097, n58098, n58099, n58100,
    n58101, n58102, n58103, n58104, n58105, n58106, n58107, n58108, n58109,
    n58110, n58111, n58112, n58113, n58114, n58115, n58116, n58117, n58118,
    n58119, n58120, n58121, n58122, n58123, n58124, n58125, n58126, n58127,
    n58128, n58129, n58130, n58131, n58132, n58133, n58134, n58135, n58136,
    n58137, n58138, n58139, n58140, n58141, n58142, n58143, n58144, n58145,
    n58146, n58147, n58148, n58149, n58150, n58151, n58152, n58153, n58154,
    n58155, n58156, n58157, n58158, n58159, n58160, n58161, n58162, n58163,
    n58164, n58165, n58166, n58167, n58168, n58169, n58170, n58171, n58172,
    n58173, n58174, n58175, n58176, n58177, n58178, n58179, n58180, n58181,
    n58182, n58183, n58184, n58185, n58186, n58187, n58188, n58189, n58190,
    n58191, n58192, n58193, n58194, n58195, n58196, n58197, n58198, n58199,
    n58200, n58201, n58202, n58203, n58204, n58205, n58206, n58207, n58208,
    n58209, n58210, n58211, n58212, n58213, n58214, n58215, n58216, n58217,
    n58218, n58219, n58220, n58221, n58222, n58223, n58224, n58225, n58226,
    n58227, n58228, n58229, n58230, n58231, n58232, n58233, n58234, n58235,
    n58236, n58237, n58238, n58239, n58240, n58241, n58242, n58243, n58244,
    n58245, n58246, n58247, n58248, n58249, n58250, n58251, n58252, n58253,
    n58254, n58255, n58256, n58257, n58258, n58259, n58260, n58261, n58262,
    n58263, n58264, n58265, n58266, n58267, n58268, n58269, n58270, n58271,
    n58272, n58273, n58274, n58275, n58276, n58277, n58278, n58279, n58280,
    n58281, n58282, n58283, n58284, n58285, n58286, n58287, n58288, n58289,
    n58290, n58291, n58292, n58293, n58294, n58295, n58296, n58297, n58298,
    n58299, n58300, n58301, n58302, n58303, n58304, n58305, n58306, n58307,
    n58308, n58309, n58310, n58311, n58312, n58313, n58314, n58315, n58316,
    n58317, n58318, n58319, n58320, n58321, n58322, n58323, n58324, n58325,
    n58326, n58327, n58328, n58329, n58330, n58331, n58332, n58333, n58334,
    n58335, n58336, n58337, n58338, n58339, n58340, n58341, n58342, n58343,
    n58344, n58345, n58346, n58347, n58348, n58349, n58350, n58351, n58352,
    n58353, n58354, n58355, n58356, n58357, n58358, n58359, n58360, n58361,
    n58362, n58363, n58364, n58365, n58366, n58367, n58368, n58369, n58370,
    n58371, n58372, n58373, n58374, n58375, n58376, n58377, n58378, n58379,
    n58380, n58381, n58382, n58383, n58384, n58385, n58386, n58387, n58388,
    n58389, n58390, n58391, n58392, n58393, n58394, n58395, n58396, n58397,
    n58398, n58399, n58400, n58401, n58402, n58403, n58404, n58405, n58406,
    n58407, n58408, n58409, n58410, n58411, n58412, n58413, n58414, n58415,
    n58416, n58417, n58418, n58419, n58420, n58421, n58422, n58423, n58424,
    n58425, n58426, n58427, n58428, n58429, n58430, n58431, n58432, n58433,
    n58434, n58435, n58436, n58437, n58438, n58439, n58440, n58441, n58442,
    n58443, n58444, n58445, n58446, n58447, n58448, n58449, n58450, n58451,
    n58452, n58453, n58454, n58455, n58456, n58457, n58458, n58459, n58460,
    n58461, n58462, n58463, n58464, n58465, n58466, n58467, n58468, n58469,
    n58470, n58471, n58472, n58473, n58474, n58475, n58476, n58477, n58478,
    n58479, n58480, n58481, n58482, n58483, n58484, n58485, n58486, n58487,
    n58488, n58489, n58490, n58491, n58492, n58493, n58494, n58495, n58496,
    n58497, n58498, n58499, n58500, n58501, n58502, n58503, n58504, n58505,
    n58506, n58507, n58508, n58509, n58510, n58511, n58512, n58513, n58514,
    n58515, n58516, n58517, n58518, n58519, n58520, n58521, n58522, n58523,
    n58524, n58525, n58526, n58527, n58528, n58529, n58530, n58531, n58532,
    n58533, n58534, n58535, n58536, n58537, n58538, n58539, n58540, n58541,
    n58542, n58543, n58544, n58545, n58546, n58547, n58548, n58549, n58550,
    n58551, n58552, n58553, n58554, n58555, n58556, n58557, n58558, n58559,
    n58560, n58561, n58562, n58563, n58564, n58565, n58566, n58567, n58568,
    n58569, n58570, n58571, n58572, n58573, n58574, n58575, n58576, n58577,
    n58578, n58579, n58580, n58581, n58582, n58583, n58584, n58585, n58586,
    n58587, n58588, n58589, n58590, n58591, n58592, n58593, n58594, n58595,
    n58596, n58597, n58598, n58599, n58600, n58601, n58602, n58603, n58604,
    n58605, n58606, n58607, n58608, n58609, n58610, n58611, n58612, n58613,
    n58614, n58615, n58616, n58617, n58618, n58619, n58620, n58621, n58622,
    n58623, n58624, n58625, n58626, n58627, n58628, n58629, n58630, n58631,
    n58632, n58633, n58634, n58635, n58636, n58637, n58638, n58639, n58640,
    n58641, n58642, n58643, n58644, n58645, n58646, n58647, n58648, n58649,
    n58650, n58651, n58652, n58653, n58654, n58655, n58656, n58657, n58658,
    n58659, n58660, n58661, n58662, n58663, n58664, n58665, n58666, n58667,
    n58668, n58669, n58670, n58671, n58672, n58673, n58674, n58675, n58676,
    n58677, n58678, n58679, n58680, n58681, n58682, n58683, n58684, n58685,
    n58686, n58687, n58688, n58689, n58690, n58691, n58692, n58693, n58694,
    n58695, n58696, n58697, n58698, n58699, n58700, n58701, n58702, n58703,
    n58704, n58705, n58706, n58707, n58708, n58709, n58710, n58711, n58712,
    n58713, n58714, n58715, n58716, n58717, n58718, n58719, n58720, n58721,
    n58722, n58723, n58724, n58725, n58726, n58727, n58728, n58729, n58730,
    n58731, n58732, n58733, n58734, n58735, n58736, n58737, n58738, n58739,
    n58740, n58741, n58742, n58743, n58744, n58745, n58746, n58747, n58748,
    n58749, n58750, n58751, n58752, n58753, n58754, n58755, n58756, n58757,
    n58758, n58759, n58760, n58761, n58762, n58763, n58764, n58765, n58766,
    n58767, n58768, n58769, n58770, n58771, n58772, n58773, n58774, n58775,
    n58776, n58777, n58778, n58779, n58780, n58781, n58782, n58783, n58784,
    n58785, n58786, n58787, n58788, n58789, n58790, n58791, n58792, n58793,
    n58794, n58795, n58796, n58797, n58798, n58799, n58800, n58801, n58802,
    n58803, n58804, n58805, n58806, n58807, n58808, n58809, n58810, n58811,
    n58812, n58813, n58814, n58815, n58816, n58817, n58818, n58819, n58820,
    n58821, n58822, n58823, n58824, n58825, n58826, n58827, n58828, n58829,
    n58830, n58831, n58832, n58833, n58834, n58835, n58836, n58837, n58838,
    n58839, n58840, n58841, n58842, n58843, n58844, n58845, n58846, n58847,
    n58848, n58849, n58850, n58851, n58852, n58853, n58854, n58855, n58856,
    n58857, n58858, n58859, n58860, n58861, n58862, n58863, n58864, n58865,
    n58866, n58867, n58868, n58869, n58870, n58871, n58872, n58873, n58874,
    n58875, n58876, n58877, n58878, n58879, n58880, n58881, n58882, n58883,
    n58884, n58885, n58886, n58887, n58888, n58889, n58890, n58891, n58892,
    n58893, n58894, n58895, n58896, n58897, n58898, n58899, n58900, n58901,
    n58902, n58903, n58904, n58905, n58906, n58907, n58908, n58909, n58910,
    n58911, n58912, n58913, n58914, n58915, n58916, n58917, n58918, n58919,
    n58920, n58921, n58922, n58923, n58924, n58925, n58926, n58927, n58928,
    n58929, n58930, n58931, n58932, n58933, n58934, n58935, n58936, n58937,
    n58938, n58939, n58940, n58941, n58942, n58943, n58944, n58945, n58946,
    n58947, n58948, n58949, n58950, n58951, n58952, n58953, n58954, n58955,
    n58956, n58957, n58958, n58959, n58960, n58961, n58962, n58963, n58964,
    n58965, n58966, n58967, n58968, n58969, n58970, n58971, n58972, n58973,
    n58974, n58975, n58976, n58977, n58978, n58979, n58980, n58981, n58982,
    n58983, n58984, n58985, n58986, n58987, n58988, n58989, n58990, n58991,
    n58992, n58993, n58994, n58995, n58996, n58997, n58998, n58999, n59000,
    n59001, n59002, n59003, n59004, n59005, n59006, n59007, n59008, n59009,
    n59010, n59011, n59012, n59013, n59014, n59015, n59016, n59017, n59018,
    n59019, n59020, n59021, n59022, n59023, n59024, n59025, n59026, n59027,
    n59028, n59029, n59030, n59031, n59032, n59033, n59034, n59035, n59036,
    n59037, n59038, n59039, n59040, n59041, n59042, n59043, n59044, n59045,
    n59046, n59047, n59048, n59049, n59050, n59051, n59052, n59053, n59054,
    n59055, n59056, n59057, n59058, n59059, n59060, n59061, n59062, n59063,
    n59064, n59065, n59066, n59067, n59068, n59069, n59070, n59071, n59072,
    n59073, n59074, n59075, n59076, n59077, n59078, n59079, n59080, n59081,
    n59082, n59083, n59084, n59085, n59086, n59087, n59088, n59089, n59090,
    n59091, n59092, n59093, n59094, n59095, n59096, n59097, n59098, n59099,
    n59100, n59101, n59102, n59103, n59104, n59105, n59106, n59107, n59108,
    n59109, n59110, n59111, n59112, n59113, n59114, n59115, n59116, n59117,
    n59118, n59119, n59120, n59121, n59122, n59123, n59124, n59125, n59126,
    n59127, n59128, n59129, n59130, n59131, n59132, n59133, n59134, n59135,
    n59136, n59137, n59138, n59139, n59140, n59141, n59142, n59143, n59144,
    n59145, n59146, n59147, n59148, n59149, n59150, n59151, n59152, n59153,
    n59154, n59155, n59156, n59157, n59158, n59159, n59160, n59161, n59162,
    n59163, n59164, n59165, n59166, n59167, n59168, n59169, n59170, n59171,
    n59172, n59173, n59174, n59175, n59176, n59177, n59178, n59179, n59180,
    n59181, n59182, n59183, n59184, n59185, n59186, n59187, n59188, n59189,
    n59190, n59191, n59192, n59193, n59194, n59195, n59196, n59197, n59198,
    n59199, n59200, n59201, n59202, n59203, n59204, n59205, n59206, n59207,
    n59208, n59209, n59210, n59211, n59212, n59213, n59214, n59215, n59216,
    n59217, n59218, n59219, n59220, n59221, n59222, n59223, n59224, n59225,
    n59226, n59227, n59228, n59229, n59230, n59231, n59232, n59233, n59234,
    n59235, n59236, n59237, n59238, n59239, n59240, n59241, n59242, n59243,
    n59244, n59245, n59246, n59247, n59248, n59249, n59250, n59251, n59252,
    n59253, n59254, n59255, n59256, n59257, n59258, n59259, n59260, n59261,
    n59262, n59263, n59264, n59265, n59266, n59267, n59268, n59269, n59270,
    n59271, n59272, n59273, n59274, n59275, n59276, n59277, n59278, n59279,
    n59280, n59281, n59282, n59283, n59284, n59285, n59286, n59287, n59288,
    n59289, n59290, n59291, n59292, n59293, n59294, n59295, n59296, n59297,
    n59298, n59299, n59300, n59301, n59302, n59303, n59304, n59305, n59306,
    n59307, n59308, n59309, n59310, n59311, n59312, n59313, n59314, n59315,
    n59316, n59317, n59318, n59319, n59320, n59321, n59322, n59323, n59324,
    n59325, n59326, n59327, n59328, n59329, n59330, n59331, n59332, n59333,
    n59334, n59335, n59336, n59337, n59338, n59339, n59340, n59341, n59342,
    n59343, n59344, n59345, n59346, n59347, n59348, n59349, n59350, n59351,
    n59352, n59353, n59354, n59355, n59356, n59357, n59358, n59359, n59360,
    n59361, n59362, n59363, n59364, n59365, n59366, n59367, n59368, n59369,
    n59370, n59371, n59372, n59373, n59374, n59375, n59376, n59377, n59378,
    n59379, n59380, n59381, n59382, n59383, n59384, n59385, n59386, n59387,
    n59388, n59389, n59390, n59391, n59392, n59393, n59394, n59395, n59396,
    n59397, n59398, n59399, n59400, n59401, n59402, n59403, n59404, n59405,
    n59406, n59407, n59408, n59409, n59410, n59411, n59412, n59413, n59414,
    n59415, n59416, n59417, n59418, n59419, n59420, n59421, n59422, n59423,
    n59424, n59425, n59426, n59427, n59428, n59429, n59430, n59431, n59432,
    n59433, n59434, n59435, n59436, n59437, n59438, n59439, n59440, n59441,
    n59442, n59443, n59444, n59445, n59446, n59447, n59448, n59449, n59450,
    n59451, n59452, n59453, n59454, n59455, n59456, n59457, n59458, n59459,
    n59460, n59461, n59462, n59463, n59464, n59465, n59466, n59467, n59468,
    n59469, n59470, n59471, n59472, n59473, n59474, n59475, n59476, n59477,
    n59478, n59479, n59480, n59481, n59482, n59483, n59484, n59485, n59486,
    n59487, n59488, n59489, n59490, n59491, n59492, n59493, n59494, n59495,
    n59496, n59497, n59498, n59499, n59500, n59501, n59502, n59503, n59504,
    n59505, n59506, n59507, n59508, n59509, n59510, n59511, n59512, n59513,
    n59514, n59515, n59516, n59517, n59518, n59519, n59520, n59521, n59522,
    n59523, n59524, n59525, n59526, n59527, n59528, n59529, n59530, n59531,
    n59532, n59533, n59534, n59535, n59536, n59537, n59538, n59539, n59540,
    n59541, n59542, n59543, n59544, n59545, n59546, n59547, n59548, n59549,
    n59550, n59551, n59552, n59553, n59554, n59555, n59556, n59557, n59558,
    n59559, n59560, n59561, n59562, n59563, n59564, n59565, n59566, n59567,
    n59568, n59569, n59570, n59571, n59572, n59573, n59574, n59575, n59576,
    n59577, n59578, n59579, n59580, n59581, n59582, n59583, n59584, n59585,
    n59586, n59587, n59588, n59589, n59590, n59591, n59592, n59593, n59594,
    n59595, n59596, n59597, n59598, n59599, n59600, n59601, n59602, n59603,
    n59604, n59605, n59606, n59607, n59608, n59609, n59610, n59611, n59612,
    n59613, n59614, n59615, n59616, n59617, n59618, n59619, n59620, n59621,
    n59622, n59623, n59624, n59625, n59626, n59627, n59628, n59629, n59630,
    n59631, n59632, n59633, n59634, n59635, n59636, n59637, n59638, n59639,
    n59640, n59641, n59642, n59643, n59644, n59645, n59646, n59647, n59648,
    n59649, n59650, n59651, n59652, n59653, n59654, n59655, n59656, n59657,
    n59658, n59659, n59660, n59661, n59662, n59663, n59664, n59665, n59666,
    n59667, n59668, n59669, n59670, n59671, n59672, n59673, n59674, n59675,
    n59676, n59677, n59678, n59679, n59680, n59681, n59682, n59683, n59684,
    n59685, n59686, n59687, n59688, n59689, n59690, n59691, n59692, n59693,
    n59694, n59695, n59696, n59697, n59698, n59699, n59700, n59701, n59702,
    n59703, n59704, n59705, n59706, n59707, n59708, n59709, n59710, n59711,
    n59712, n59713, n59714, n59715, n59716, n59717, n59718, n59719, n59720,
    n59721, n59722, n59723, n59724, n59725, n59726, n59727, n59728, n59729,
    n59730, n59731, n59732, n59733, n59734, n59735, n59736, n59737, n59738,
    n59739, n59740, n59741, n59742, n59743, n59744, n59745, n59746, n59747,
    n59748, n59749, n59750, n59751, n59752, n59753, n59754, n59755, n59756,
    n59757, n59758, n59759, n59760, n59761, n59762, n59763, n59764, n59765,
    n59766, n59767, n59768, n59769, n59770, n59771, n59772, n59773, n59774,
    n59775, n59776, n59777, n59778, n59779, n59780, n59781, n59782, n59783,
    n59784, n59785, n59786, n59787, n59788, n59789, n59790, n59791, n59792,
    n59793, n59794, n59795, n59796, n59797, n59798, n59799, n59800, n59801,
    n59802, n59803, n59804, n59805, n59806, n59807, n59808, n59809, n59810,
    n59811, n59812, n59813, n59814, n59815, n59816, n59817, n59818, n59819,
    n59820, n59821, n59822, n59823, n59824, n59825, n59826, n59827, n59828,
    n59829, n59830, n59831, n59832, n59833, n59834, n59835, n59836, n59837,
    n59838, n59839, n59840, n59841, n59842, n59843, n59844, n59845, n59846,
    n59847, n59848, n59849, n59850, n59851, n59852, n59853, n59854, n59855,
    n59856, n59857, n59858, n59859, n59860, n59861, n59862, n59863, n59864,
    n59865, n59866, n59867, n59868, n59869, n59870, n59871, n59872, n59873,
    n59874, n59875, n59876, n59877, n59878, n59879, n59880, n59881, n59882,
    n59883, n59884, n59885, n59886, n59887, n59888, n59889, n59890, n59891,
    n59892, n59893, n59894, n59895, n59896, n59897, n59898, n59899, n59900,
    n59901, n59902, n59903, n59904, n59905, n59906, n59907, n59908, n59909,
    n59910, n59911, n59912, n59913, n59914, n59915, n59916, n59917, n59918,
    n59919, n59920, n59921, n59922, n59923, n59924, n59925, n59926, n59927,
    n59928, n59929, n59930, n59931, n59932, n59933, n59934, n59935, n59936,
    n59937, n59938, n59939, n59940, n59941, n59942, n59943, n59944, n59945,
    n59946, n59947, n59948, n59949, n59950, n59951, n59952, n59953, n59954,
    n59955, n59956, n59957, n59958, n59959, n59960, n59961, n59962, n59963,
    n59964, n59965, n59966, n59967, n59968, n59969, n59970, n59971, n59972,
    n59973, n59974, n59975, n59976, n59977, n59978, n59979, n59980, n59981,
    n59982, n59983, n59984, n59985, n59986, n59987, n59988, n59989, n59990,
    n59991, n59992, n59993, n59994, n59995, n59996, n59997, n59998, n59999,
    n60000, n60001, n60002, n60003, n60004, n60005, n60006, n60007, n60008,
    n60009, n60010, n60011, n60012, n60013, n60014, n60015, n60016, n60017,
    n60018, n60019, n60020, n60021, n60022, n60023, n60024, n60025, n60026,
    n60027, n60028, n60029, n60030, n60031, n60032, n60033, n60034, n60035,
    n60036, n60037, n60038, n60039, n60040, n60041, n60042, n60043, n60044,
    n60045, n60046, n60047, n60048, n60049, n60050, n60051, n60052, n60053,
    n60054, n60055, n60056, n60057, n60058, n60059, n60060, n60061, n60062,
    n60063, n60064, n60065, n60066, n60067, n60068, n60069, n60070, n60071,
    n60072, n60073, n60074, n60075, n60076, n60077, n60078, n60079, n60080,
    n60081, n60082, n60083, n60084, n60085, n60086, n60087, n60088, n60089,
    n60090, n60091, n60092, n60093, n60094, n60095, n60096, n60097, n60098,
    n60099, n60100, n60101, n60102, n60103, n60104, n60105, n60106, n60107,
    n60108, n60109, n60110, n60111, n60112, n60113, n60114, n60115, n60116,
    n60117, n60118, n60119, n60120, n60121, n60122, n60123, n60124, n60125,
    n60126, n60127, n60128, n60129, n60130, n60131, n60132, n60133, n60134,
    n60135, n60136, n60137, n60138, n60139, n60140, n60141, n60142, n60143,
    n60144, n60145, n60146, n60147, n60148, n60149, n60150, n60151, n60152,
    n60153, n60154, n60155, n60156, n60157, n60158, n60159, n60160, n60161,
    n60162, n60163, n60164, n60165, n60166, n60167, n60168, n60169, n60170,
    n60171, n60172, n60173, n60174, n60175, n60176, n60177, n60178, n60179,
    n60180, n60181, n60182, n60183, n60184, n60185, n60186, n60187, n60188,
    n60189, n60190, n60191, n60192, n60193, n60194, n60195, n60196, n60197,
    n60198, n60199, n60200, n60201, n60202, n60203, n60204, n60205, n60206,
    n60207, n60208, n60209, n60210, n60211, n60212, n60213, n60214, n60215,
    n60216, n60217, n60218, n60219, n60220, n60221, n60222, n60223, n60224,
    n60225, n60226, n60227, n60228, n60229, n60230, n60231, n60232, n60233,
    n60234, n60235, n60236, n60237, n60238, n60239, n60240, n60241, n60242,
    n60243, n60244, n60245, n60246, n60247, n60248, n60249, n60250, n60251,
    n60252, n60253, n60254, n60255, n60256, n60257, n60258, n60259, n60260,
    n60261, n60262, n60263, n60264, n60265, n60266, n60267, n60268, n60269,
    n60270, n60271, n60272, n60273, n60274, n60275, n60276, n60277, n60278,
    n60279, n60280, n60281, n60282, n60283, n60284, n60285, n60286, n60287,
    n60288, n60289, n60290, n60291, n60292, n60293, n60294, n60295, n60296,
    n60297, n60298, n60299, n60300, n60301, n60302, n60303, n60304, n60305,
    n60306, n60307, n60308, n60309, n60310, n60311, n60312, n60313, n60314,
    n60315, n60316, n60317, n60318, n60319, n60320, n60321, n60322, n60323,
    n60324, n60325, n60326, n60327, n60328, n60329, n60330, n60331, n60332,
    n60333, n60334, n60335, n60336, n60337, n60338, n60339, n60340, n60341,
    n60342, n60343, n60344, n60345, n60346, n60347, n60348, n60349, n60350,
    n60351, n60352, n60353, n60354, n60355, n60356, n60357, n60358, n60359,
    n60360, n60361, n60362, n60363, n60364, n60365, n60366, n60367, n60368,
    n60369, n60370, n60371, n60372, n60373, n60374, n60375, n60376, n60377,
    n60378, n60379, n60380, n60381, n60382, n60383, n60384, n60385, n60386,
    n60387, n60388, n60389, n60390, n60391, n60392, n60393, n60394, n60395,
    n60396, n60397, n60398, n60399, n60400, n60401, n60402, n60403, n60404,
    n60405, n60406, n60407, n60408, n60409, n60410, n60411, n60412, n60413,
    n60414, n60415, n60416, n60417, n60418, n60419, n60420, n60421, n60422,
    n60423, n60424, n60425, n60426, n60427, n60428, n60429, n60430, n60431,
    n60432, n60433, n60434, n60435, n60436, n60437, n60438, n60439, n60440,
    n60441, n60442, n60443, n60444, n60445, n60446, n60447, n60448, n60449,
    n60450, n60451, n60452, n60453, n60454, n60455, n60456, n60457, n60458,
    n60459, n60460, n60461, n60462, n60463, n60464, n60465, n60466, n60467,
    n60468, n60469, n60470, n60471, n60472, n60473, n60474, n60475, n60476,
    n60477, n60478, n60479, n60480, n60481, n60482, n60483, n60484, n60485,
    n60486, n60487, n60488, n60489, n60490, n60491, n60492, n60493, n60494,
    n60495, n60496, n60497, n60498, n60499, n60500, n60501, n60502, n60503,
    n60504, n60505, n60506, n60507, n60508, n60509, n60510, n60511, n60512,
    n60513, n60514, n60515, n60516, n60517, n60518, n60519, n60520, n60521,
    n60522, n60523, n60524, n60525, n60526, n60527, n60528, n60529, n60530,
    n60531, n60532, n60533, n60534, n60535, n60536, n60537, n60538, n60539,
    n60540, n60541, n60542, n60543, n60544, n60545, n60546, n60547, n60548,
    n60549, n60550, n60551, n60552, n60553, n60554, n60555, n60556, n60557,
    n60558, n60559, n60560, n60561, n60562, n60563, n60564, n60565, n60566,
    n60567, n60568, n60569, n60570, n60571, n60572, n60573, n60574, n60575,
    n60576, n60577, n60578, n60579, n60580, n60581, n60582, n60583, n60584,
    n60585, n60586, n60587, n60588, n60589, n60590, n60591, n60592, n60593,
    n60594, n60595, n60596, n60597, n60598, n60599, n60600, n60601, n60602,
    n60603, n60604, n60605, n60606, n60607, n60608, n60609, n60610, n60611,
    n60612, n60613, n60614, n60615, n60616, n60617, n60618, n60619, n60620,
    n60621, n60622, n60623, n60624, n60625, n60626, n60627, n60628, n60629,
    n60630, n60631, n60632, n60633, n60634, n60635, n60636, n60637, n60638,
    n60639, n60640, n60641, n60642, n60643, n60644, n60645, n60646, n60647,
    n60648, n60649, n60650, n60651, n60652, n60653, n60654, n60655, n60656,
    n60657, n60658, n60659, n60660, n60661, n60662, n60663, n60664, n60665,
    n60666, n60667, n60668, n60669, n60670, n60671, n60672, n60673, n60674,
    n60675, n60676, n60677, n60678, n60679, n60680, n60681, n60682, n60683,
    n60684, n60685, n60686, n60687, n60688, n60689, n60690, n60691, n60692,
    n60693, n60694, n60695, n60696, n60697, n60698, n60699, n60700, n60701,
    n60702, n60703, n60704, n60705, n60706, n60707, n60708, n60709, n60710,
    n60711, n60712, n60713, n60714, n60715, n60716, n60717, n60718, n60719,
    n60720, n60721, n60722, n60723, n60724, n60725, n60726, n60727, n60728,
    n60729, n60730, n60731, n60732, n60733, n60734, n60735, n60736, n60737,
    n60738, n60739, n60740, n60741, n60742, n60743, n60744, n60745, n60746,
    n60747, n60748, n60749, n60750, n60751, n60752, n60753, n60754, n60755,
    n60756, n60757, n60758, n60759, n60760, n60761, n60762, n60763, n60764,
    n60765, n60766, n60767, n60768, n60769, n60770, n60771, n60772, n60773,
    n60774, n60775, n60776, n60777, n60778, n60779, n60780, n60781, n60782,
    n60783, n60784, n60785, n60786, n60787, n60788, n60789, n60790, n60791,
    n60792, n60793, n60794, n60795, n60796, n60797, n60798, n60799, n60800,
    n60801, n60802, n60803, n60804, n60805, n60806, n60807, n60808, n60809,
    n60810, n60811, n60812, n60813, n60814, n60815, n60816, n60817, n60818,
    n60819, n60820, n60821, n60822, n60823, n60824, n60825, n60826, n60827,
    n60828, n60829, n60830, n60831, n60832, n60833, n60834, n60835, n60836,
    n60837, n60838, n60839, n60840, n60841, n60842, n60843, n60844, n60845,
    n60846, n60847, n60848, n60849, n60850, n60851, n60852, n60853, n60854,
    n60855, n60856, n60857, n60858, n60859, n60860, n60861, n60862, n60863,
    n60864, n60865, n60866, n60867, n60868, n60869, n60870, n60871, n60872,
    n60873, n60874, n60875, n60876, n60877, n60878, n60879, n60880, n60881,
    n60882, n60883, n60884, n60885, n60886, n60887, n60888, n60889, n60890,
    n60891, n60892, n60893, n60894, n60895, n60896, n60897, n60898, n60899,
    n60900, n60901, n60902, n60903, n60904, n60905, n60906, n60907, n60908,
    n60909, n60910, n60911, n60912, n60913, n60914, n60915, n60916, n60917,
    n60918, n60919, n60920, n60921, n60922, n60923, n60924, n60925, n60926,
    n60927, n60928, n60929, n60930, n60931, n60932, n60933, n60934, n60935,
    n60936, n60937, n60938, n60939, n60940, n60941, n60942, n60943, n60944,
    n60945, n60946, n60947, n60948, n60949, n60950, n60951, n60952, n60953,
    n60954, n60955, n60956, n60957, n60958, n60959, n60960, n60961, n60962,
    n60963, n60964, n60965, n60966, n60967, n60968, n60969, n60970, n60971,
    n60972, n60973, n60974, n60975, n60976, n60977, n60978, n60979, n60980,
    n60981, n60982, n60983, n60984, n60985, n60986, n60987, n60988, n60989,
    n60990, n60991, n60992, n60993, n60994, n60995, n60996, n60997, n60998,
    n60999, n61000, n61001, n61002, n61003, n61004, n61005, n61006, n61007,
    n61008, n61009, n61010, n61011, n61012, n61013, n61014, n61015, n61016,
    n61017, n61018, n61019, n61020, n61021, n61022, n61023, n61024, n61025,
    n61026, n61027, n61028, n61029, n61030, n61031, n61032, n61033, n61034,
    n61035, n61036, n61037, n61038, n61039, n61040, n61041, n61042, n61043,
    n61044, n61045, n61046, n61047, n61048, n61049, n61050, n61051, n61052,
    n61053, n61054, n61055, n61056, n61057, n61058, n61059, n61060, n61061,
    n61062, n61063, n61064, n61065, n61066, n61067, n61068, n61069, n61070,
    n61071, n61072, n61073, n61074, n61075, n61076, n61077, n61078, n61079,
    n61080, n61081, n61082, n61083, n61084, n61085, n61086, n61087, n61088,
    n61089, n61090, n61091, n61092, n61093, n61094, n61095, n61096, n61097,
    n61098, n61099, n61100, n61101, n61102, n61103, n61104, n61105, n61106,
    n61107, n61108, n61109, n61110, n61111, n61112, n61113, n61114, n61115,
    n61116, n61117, n61118, n61119, n61120, n61121, n61122, n61123, n61124,
    n61125, n61126, n61127, n61128, n61129, n61130, n61131, n61132, n61133,
    n61134, n61135, n61136, n61137, n61138, n61139, n61140, n61141, n61142,
    n61143, n61144, n61145, n61146, n61147, n61148, n61149, n61150, n61151,
    n61152, n61153, n61154, n61155, n61156, n61157, n61158, n61159, n61160,
    n61161, n61162, n61163, n61164, n61165, n61166, n61167, n61168, n61169,
    n61170, n61171, n61172, n61173, n61174, n61175, n61176, n61177, n61178,
    n61179, n61180, n61181, n61182, n61183, n61184, n61185, n61186, n61187,
    n61188, n61189, n61190, n61191, n61192, n61193, n61194, n61195, n61196,
    n61197, n61198, n61199, n61200, n61201, n61202, n61203, n61204, n61205,
    n61206, n61207, n61208, n61209, n61210, n61211, n61212, n61213, n61214,
    n61215, n61216, n61217, n61218, n61219, n61220, n61221, n61222, n61223,
    n61224, n61225, n61226, n61227, n61228, n61229, n61230, n61231, n61232,
    n61233, n61234, n61235, n61236, n61237, n61238, n61239, n61240, n61241,
    n61242, n61243, n61244, n61245, n61246, n61247, n61248, n61249, n61250,
    n61251, n61252, n61253, n61254, n61255, n61256, n61257, n61258, n61259,
    n61260, n61261, n61262, n61263, n61264, n61265, n61266, n61267, n61268,
    n61269, n61270, n61271, n61272, n61273, n61274, n61275, n61276, n61277,
    n61278, n61279, n61280, n61281, n61282, n61283, n61284, n61285, n61286,
    n61287, n61288, n61289, n61290, n61291, n61292, n61293, n61294, n61295,
    n61296, n61297, n61298, n61299, n61300, n61301, n61302, n61303, n61304,
    n61305, n61306, n61307, n61308, n61309, n61310, n61311, n61312, n61313,
    n61314, n61315, n61316, n61317, n61318, n61319, n61320, n61321, n61322,
    n61323, n61324, n61325, n61326, n61327, n61328, n61329, n61330, n61331,
    n61332, n61333, n61334, n61335, n61336, n61337, n61338, n61339, n61340,
    n61341, n61342, n61343, n61344, n61345, n61346, n61347, n61348, n61349,
    n61350, n61351, n61352, n61353, n61354, n61355, n61356, n61357, n61358,
    n61359, n61360, n61361, n61362, n61363, n61364, n61365, n61366, n61367,
    n61368, n61369, n61370, n61371, n61372, n61373, n61374, n61375, n61376,
    n61377, n61378, n61379, n61380, n61381, n61382, n61383, n61384, n61385,
    n61386, n61387, n61388, n61389, n61390, n61391, n61392, n61393, n61394,
    n61395, n61396, n61397, n61398, n61399, n61400, n61401, n61402, n61403,
    n61404, n61405, n61406, n61407, n61408, n61409, n61410, n61411, n61412,
    n61413, n61414, n61415, n61416, n61417, n61418, n61419, n61420, n61421,
    n61422, n61423, n61424, n61425, n61426, n61427, n61428, n61429, n61430,
    n61431, n61432, n61433, n61434, n61435, n61436, n61437, n61438, n61439,
    n61440, n61441, n61442, n61443, n61444, n61445, n61446, n61447, n61448,
    n61449, n61450, n61451, n61452, n61453, n61454, n61455, n61456, n61457,
    n61458, n61459, n61460, n61461, n61462, n61463, n61464, n61465, n61466,
    n61467, n61468, n61469, n61470, n61471, n61472, n61473, n61474, n61475,
    n61476, n61477, n61478, n61479, n61480, n61481, n61482, n61483, n61484,
    n61485, n61486, n61487, n61488, n61489, n61490, n61491, n61492, n61493,
    n61494, n61495, n61496, n61497, n61498, n61499, n61500, n61501, n61502,
    n61503, n61504, n61505, n61506, n61507, n61508, n61509, n61510, n61511,
    n61512, n61513, n61514, n61515, n61516, n61517, n61518, n61519, n61520,
    n61521, n61522, n61523, n61524, n61525, n61526, n61527, n61528, n61529,
    n61530, n61531, n61532, n61533, n61534, n61535, n61536, n61537, n61538,
    n61539, n61540, n61541, n61542, n61543, n61544, n61545, n61546, n61547,
    n61548, n61549, n61550, n61551, n61552, n61553, n61554, n61555, n61556,
    n61557, n61558, n61559, n61560, n61561, n61562, n61563, n61564, n61565,
    n61566, n61567, n61568, n61569, n61570, n61571, n61572, n61573, n61574,
    n61575, n61576, n61577, n61578, n61579, n61580, n61581, n61582, n61583,
    n61584, n61585, n61586, n61587, n61588, n61589, n61590, n61591, n61592,
    n61593, n61594, n61595, n61596, n61597, n61598, n61599, n61600, n61601,
    n61602, n61603, n61604, n61605, n61606, n61607, n61608, n61609, n61610,
    n61611, n61612, n61613, n61614, n61615, n61616, n61617, n61618, n61619,
    n61620, n61621, n61622, n61623, n61624, n61625, n61626, n61627, n61628,
    n61629, n61630, n61631, n61632, n61633, n61634, n61635, n61636, n61637,
    n61638, n61639, n61640, n61641, n61642, n61643, n61644, n61645, n61646,
    n61647, n61648, n61649, n61650, n61651, n61652, n61653, n61654, n61655,
    n61656, n61657, n61658, n61659, n61660, n61661, n61662, n61663, n61664,
    n61665, n61666, n61667, n61668, n61669, n61670, n61671, n61672, n61673,
    n61674, n61675, n61676, n61677, n61678, n61679, n61680, n61681, n61682,
    n61683, n61684, n61685, n61686, n61687, n61688, n61689, n61690, n61691,
    n61692, n61693, n61694, n61695, n61696, n61697, n61698, n61699, n61700,
    n61701, n61702, n61703, n61704, n61705, n61706, n61707, n61708, n61709,
    n61710, n61711, n61712, n61713, n61714, n61715, n61716, n61717, n61718,
    n61719, n61720, n61721, n61722, n61723, n61724, n61725, n61726, n61727,
    n61728, n61729, n61730, n61731, n61732, n61733, n61734, n61735, n61736,
    n61737, n61738, n61739, n61740, n61741, n61742, n61743, n61744, n61745,
    n61746, n61747, n61748, n61749, n61750, n61751, n61752, n61753, n61754,
    n61755, n61756, n61757, n61758, n61759, n61760, n61761, n61762, n61763,
    n61764, n61765, n61766, n61767, n61768, n61769, n61770, n61771, n61772,
    n61773, n61774, n61775, n61776, n61777, n61778, n61779, n61780, n61781,
    n61782, n61783, n61784, n61785, n61786, n61787, n61788, n61789, n61790,
    n61791, n61792, n61793, n61794, n61795, n61796, n61797, n61798, n61799,
    n61800, n61801, n61802, n61803, n61804, n61805, n61806, n61807, n61808,
    n61809, n61810, n61811, n61812, n61813, n61814, n61815, n61816, n61817,
    n61818, n61819, n61820, n61821, n61822, n61823, n61824, n61825, n61826,
    n61827, n61828, n61829, n61830, n61831, n61832, n61833, n61834, n61835,
    n61836, n61837, n61838, n61839, n61840, n61841, n61842, n61843, n61844,
    n61845, n61846, n61847, n61848, n61849, n61850, n61851, n61852, n61853,
    n61854, n61855, n61856, n61857, n61858, n61859, n61860, n61861, n61862,
    n61863, n61864, n61865, n61866, n61867, n61868, n61869, n61870, n61871,
    n61872, n61873, n61874, n61875, n61876, n61877, n61878, n61879, n61880,
    n61881, n61882, n61883, n61884, n61885, n61886, n61887, n61888, n61889,
    n61890, n61891, n61892, n61893, n61894, n61895, n61896, n61897, n61898,
    n61899, n61900, n61901, n61902, n61903, n61904, n61905, n61906, n61907,
    n61908, n61909, n61910, n61911, n61912, n61913, n61914, n61915, n61916,
    n61917, n61918, n61919, n61920, n61921, n61922, n61923, n61924, n61925,
    n61926, n61927, n61928, n61929, n61930, n61931, n61932, n61933, n61934,
    n61935, n61936, n61937, n61938, n61939, n61940, n61941, n61942, n61943,
    n61944, n61945, n61946, n61947, n61948, n61949, n61950, n61951, n61952,
    n61953, n61954, n61955, n61956, n61957, n61958, n61959, n61960, n61961,
    n61962, n61963, n61964, n61965, n61966, n61967, n61968, n61969, n61970,
    n61971, n61972, n61973, n61974, n61975, n61976, n61977, n61978, n61979,
    n61980, n61981, n61982, n61983, n61984, n61985, n61986, n61987, n61988,
    n61989, n61990, n61991, n61992, n61993, n61994, n61995, n61996, n61997,
    n61998, n61999, n62000, n62001, n62002, n62003, n62004, n62005, n62006,
    n62007, n62008, n62009, n62010, n62011, n62012, n62013, n62014, n62015,
    n62016, n62017, n62018, n62019, n62020, n62021, n62022, n62023, n62024,
    n62025, n62026, n62027, n62028, n62029, n62030, n62031, n62032, n62033,
    n62034, n62035, n62036, n62037, n62038, n62039, n62040, n62041, n62042,
    n62043, n62044, n62045, n62046, n62047, n62048, n62049, n62050, n62051,
    n62052, n62053, n62054, n62055, n62056, n62057, n62058, n62059, n62060,
    n62061, n62062, n62063, n62064, n62065, n62066, n62067, n62068, n62069,
    n62070, n62071, n62072, n62073, n62074, n62075, n62076, n62077, n62078,
    n62079, n62080, n62081, n62082, n62083, n62084, n62085, n62086, n62087,
    n62088, n62089, n62090, n62091, n62092, n62093, n62094, n62095, n62096,
    n62097, n62098, n62099, n62100, n62101, n62102, n62103, n62104, n62105,
    n62106, n62107, n62108, n62109, n62110, n62111, n62112, n62113, n62114,
    n62115, n62116, n62117, n62118, n62119, n62120, n62121, n62122, n62123,
    n62124, n62125, n62126, n62127, n62128, n62129, n62130, n62131, n62132,
    n62133, n62134, n62135, n62136, n62137, n62138, n62139, n62140, n62141,
    n62142, n62143, n62144, n62145, n62146, n62147, n62148, n62149, n62150,
    n62151, n62152, n62153, n62154, n62155, n62156, n62157, n62158, n62159,
    n62160, n62161, n62162, n62163, n62164, n62165, n62166, n62167, n62168,
    n62169, n62170, n62171, n62172, n62173, n62174, n62175, n62176, n62177,
    n62178, n62179, n62180, n62181, n62182, n62183, n62184, n62185, n62186,
    n62187, n62188, n62189, n62190, n62191, n62192, n62193, n62194, n62195,
    n62196, n62197, n62198, n62199, n62200, n62201, n62202, n62203, n62204,
    n62205, n62206, n62207, n62208, n62209, n62210, n62211, n62212, n62213,
    n62214, n62215, n62216, n62217, n62218, n62219, n62220, n62221, n62222,
    n62223, n62224, n62225, n62226, n62227, n62228, n62229, n62230, n62231,
    n62232, n62233, n62234, n62235, n62236, n62237, n62238, n62239, n62240,
    n62241, n62242, n62243, n62244, n62245, n62246, n62247, n62248, n62249,
    n62250, n62251, n62252, n62253, n62254, n62255, n62256, n62257, n62258,
    n62259, n62260, n62261, n62262, n62263, n62264, n62265, n62266, n62267,
    n62268, n62269, n62270, n62271, n62272, n62273, n62274, n62275, n62276,
    n62277, n62278, n62279, n62280, n62281, n62282, n62283, n62284, n62285,
    n62286, n62287, n62288, n62289, n62290, n62291, n62292, n62293, n62294,
    n62295, n62296, n62297, n62298, n62299, n62300, n62301, n62302, n62303,
    n62304, n62305, n62306, n62307, n62308, n62309, n62310, n62311, n62312,
    n62313, n62314, n62315, n62316, n62317, n62318, n62319, n62320, n62321,
    n62322, n62323, n62324, n62325, n62326, n62327, n62328, n62329, n62330,
    n62331, n62332, n62333, n62334, n62335, n62336, n62337, n62338, n62339,
    n62340, n62341, n62342, n62343, n62344, n62345, n62346, n62347, n62348,
    n62349, n62350, n62351, n62352, n62353, n62354, n62355, n62356, n62357,
    n62358, n62359, n62360, n62361, n62362, n62363, n62364, n62365, n62366,
    n62367, n62368, n62369, n62370, n62371, n62372, n62373, n62374, n62375,
    n62376, n62377, n62378, n62379, n62380, n62381, n62382, n62383, n62384,
    n62385, n62386, n62387, n62388, n62389, n62390, n62391, n62392, n62393,
    n62394, n62395, n62396, n62397, n62398, n62399, n62400, n62401, n62402,
    n62403, n62404, n62405, n62406, n62407, n62408, n62409, n62410, n62411,
    n62412, n62413, n62414, n62415, n62416, n62417, n62418, n62419, n62420,
    n62421, n62422, n62423, n62424, n62425, n62426, n62427, n62428, n62429,
    n62430, n62431, n62432, n62433, n62434, n62435, n62436, n62437, n62438,
    n62439, n62440, n62441, n62442, n62443, n62444, n62445, n62446, n62447,
    n62448, n62449, n62450, n62451, n62452, n62453, n62454, n62455, n62456,
    n62457, n62458, n62459, n62460, n62461, n62462, n62463, n62464, n62465,
    n62466, n62467, n62468, n62469, n62470, n62471, n62472, n62473, n62474,
    n62475, n62476, n62477, n62478, n62479, n62480, n62481, n62482, n62483,
    n62484, n62485, n62486, n62487, n62488, n62489, n62490, n62491, n62492,
    n62493, n62494, n62495, n62496, n62497, n62498, n62499, n62500, n62501,
    n62502, n62503, n62504, n62505, n62506, n62507, n62508, n62509, n62510,
    n62511, n62512, n62513, n62514, n62515, n62516, n62517, n62518, n62519,
    n62520, n62521, n62522, n62523, n62524, n62525, n62526, n62527, n62528,
    n62529, n62530, n62531, n62532, n62533, n62534, n62535, n62536, n62537,
    n62538, n62539, n62540, n62541, n62542, n62543, n62544, n62545, n62546,
    n62547, n62548, n62549, n62550, n62551, n62552, n62553, n62554, n62555,
    n62556, n62557, n62558, n62559, n62560, n62561, n62562, n62563, n62564,
    n62565, n62566, n62567, n62568, n62569, n62570, n62571, n62572, n62573,
    n62574, n62575, n62576, n62577, n62578, n62579, n62580, n62581, n62582,
    n62583, n62584, n62585, n62586, n62587, n62588, n62589, n62590, n62591,
    n62592, n62593, n62594, n62595, n62596, n62597, n62598, n62599, n62600,
    n62601, n62602, n62603, n62604, n62605, n62606, n62607, n62608, n62609,
    n62610, n62611, n62612, n62613, n62614, n62615, n62616, n62617, n62618,
    n62619, n62620, n62621, n62622, n62623, n62624, n62625, n62626, n62627,
    n62628, n62629, n62630, n62631, n62632, n62633, n62634, n62635, n62636,
    n62637, n62638, n62639, n62640, n62641, n62642, n62643, n62644, n62645,
    n62646, n62647, n62648, n62649, n62650, n62651, n62652, n62653, n62654,
    n62655, n62656, n62657, n62658, n62659, n62660, n62661, n62662, n62663,
    n62664, n62665, n62666, n62667, n62668, n62669, n62670, n62671, n62672,
    n62673, n62674, n62675, n62676, n62677, n62678, n62679, n62680, n62681,
    n62682, n62683, n62684, n62685, n62686, n62687, n62688, n62689, n62690,
    n62691, n62692, n62693, n62694, n62695, n62696, n62697, n62698, n62699,
    n62700, n62701, n62702, n62703, n62704, n62705, n62706, n62707, n62708,
    n62709, n62710, n62711, n62712, n62713, n62714, n62715, n62716, n62717,
    n62718, n62719, n62720, n62721, n62722, n62723, n62724, n62725, n62726,
    n62727, n62728, n62729, n62730, n62731, n62732, n62733, n62734, n62735,
    n62736, n62737, n62738, n62739, n62740, n62741, n62742, n62743, n62744,
    n62745, n62746, n62747, n62748, n62749, n62750, n62751, n62752, n62753,
    n62754, n62755, n62756, n62757, n62758, n62759, n62760, n62761, n62762,
    n62763, n62764, n62765, n62766, n62767, n62768, n62769, n62770, n62771,
    n62772, n62773, n62774, n62775, n62776, n62777, n62778, n62779, n62780,
    n62781, n62782, n62783, n62784, n62785, n62786, n62787, n62788, n62789,
    n62790, n62791, n62792, n62793, n62794, n62795, n62796, n62797, n62798,
    n62799, n62800, n62801, n62802, n62803, n62804, n62805, n62806, n62807,
    n62808, n62809, n62810, n62811, n62812, n62813, n62814, n62815, n62816,
    n62817, n62818, n62819, n62820, n62821, n62822, n62823, n62824, n62825,
    n62826, n62827, n62828, n62829, n62830, n62831, n62832, n62833, n62834,
    n62835, n62836, n62837, n62838, n62839, n62840, n62841, n62842, n62843,
    n62844, n62845, n62846, n62847, n62848, n62849, n62850, n62851, n62852,
    n62853, n62854, n62855, n62856, n62857, n62858, n62859, n62860, n62861,
    n62862, n62863, n62864, n62865, n62866, n62867, n62868, n62869, n62870,
    n62871, n62872, n62873, n62874, n62875, n62876, n62877, n62878, n62879,
    n62880, n62881, n62882, n62883, n62884, n62885, n62886, n62887, n62888,
    n62889, n62890, n62891, n62892, n62893, n62894, n62895, n62896, n62897,
    n62898, n62899, n62900, n62901, n62902, n62903, n62904, n62905, n62906,
    n62907, n62908, n62909, n62910, n62911, n62912, n62913, n62914, n62915,
    n62916, n62917, n62918, n62919, n62920, n62921, n62922, n62923, n62924,
    n62925, n62926, n62927, n62928, n62929, n62930, n62931, n62932, n62933,
    n62934, n62935, n62936, n62937, n62938, n62939, n62940, n62941, n62942,
    n62943, n62944, n62945, n62946, n62947, n62948, n62949, n62950, n62951,
    n62952, n62953, n62954, n62955, n62956, n62957, n62958, n62959, n62960,
    n62961, n62962, n62963, n62964, n62965, n62966, n62967, n62968, n62969,
    n62970, n62971, n62972, n62973, n62974, n62975, n62976, n62977, n62978,
    n62979, n62980, n62981, n62982, n62983, n62984, n62985, n62986, n62987,
    n62988, n62989, n62990, n62991, n62992, n62993, n62994, n62995, n62996,
    n62997, n62998, n62999, n63000, n63001, n63002, n63003, n63004, n63005,
    n63006, n63007, n63008, n63009, n63010, n63011, n63012, n63013, n63014,
    n63015, n63016, n63017, n63018, n63019, n63020, n63021, n63022, n63023,
    n63024, n63025, n63026, n63027, n63028, n63029, n63030, n63031, n63032,
    n63033, n63034, n63035, n63036, n63037, n63038, n63039, n63040, n63041,
    n63042, n63043, n63044, n63045, n63046, n63047, n63048, n63049, n63050,
    n63051, n63052, n63053, n63054, n63055, n63056, n63057, n63058, n63059,
    n63060, n63061, n63062, n63063, n63064, n63065, n63066, n63067, n63068,
    n63069, n63070, n63071, n63072, n63073, n63074, n63075, n63076, n63077,
    n63078, n63079, n63080, n63081, n63082, n63083, n63084, n63085, n63086,
    n63087, n63088, n63089, n63090, n63091, n63092, n63093, n63094, n63095,
    n63096, n63097, n63098, n63099, n63100, n63101, n63102, n63103, n63104,
    n63105, n63106, n63107, n63108, n63109, n63110, n63111, n63112, n63113,
    n63114, n63115, n63116, n63117, n63118, n63119, n63120, n63121, n63122,
    n63123, n63124, n63125, n63126, n63127, n63128, n63129, n63130, n63131,
    n63132, n63133, n63134, n63135, n63136, n63137, n63138, n63139, n63140,
    n63141, n63142, n63143, n63144, n63145, n63146, n63147, n63148, n63149,
    n63150, n63151, n63152, n63153, n63154, n63155, n63156, n63157, n63158,
    n63159, n63160, n63161, n63162, n63163, n63164, n63165, n63166, n63167,
    n63168, n63169, n63170, n63171, n63172, n63173, n63174, n63175, n63176,
    n63177, n63178, n63179, n63180, n63181, n63182, n63183, n63184, n63185,
    n63186, n63187, n63188, n63189, n63190, n63191, n63192, n63193, n63194,
    n63195, n63196, n63197, n63198, n63199, n63200, n63201, n63202, n63203,
    n63204, n63205, n63206, n63207, n63208, n63209, n63210, n63211, n63212,
    n63213, n63214, n63215, n63216, n63217, n63218, n63219, n63220, n63221,
    n63222, n63223, n63224, n63225, n63226, n63227, n63228, n63229, n63230,
    n63231, n63232, n63233, n63234, n63235, n63236, n63237, n63238, n63239,
    n63240, n63241, n63242, n63243, n63244, n63245, n63246, n63247, n63248,
    n63249, n63250, n63251, n63252, n63253, n63254, n63255, n63256, n63257,
    n63258, n63259, n63260, n63261, n63262, n63263, n63264, n63265, n63266,
    n63267, n63268, n63269, n63270, n63271, n63272, n63273, n63274, n63275,
    n63276, n63277, n63278, n63279, n63280, n63281, n63282, n63283, n63284,
    n63285, n63286, n63287, n63288, n63289, n63290, n63291, n63292, n63293,
    n63294, n63295, n63296, n63297, n63298, n63299, n63300, n63301, n63302,
    n63303, n63304, n63305, n63306, n63307, n63308, n63309, n63310, n63311,
    n63312, n63313, n63314, n63315, n63316, n63317, n63318, n63319, n63320,
    n63321, n63322, n63323, n63324, n63325, n63326, n63327, n63328, n63329,
    n63330, n63331, n63332, n63333, n63334, n63335, n63336, n63337, n63338,
    n63339, n63340, n63341, n63342, n63343, n63344, n63345, n63346, n63347,
    n63348, n63349, n63350, n63351, n63352, n63353, n63354, n63355, n63356,
    n63357, n63358, n63359, n63360, n63361, n63362, n63363, n63364, n63365,
    n63366, n63367, n63368, n63369, n63370, n63371, n63372, n63373, n63374,
    n63375, n63376, n63377, n63378, n63379, n63380, n63381, n63382, n63383,
    n63384, n63385, n63386, n63387, n63388, n63389, n63390, n63391, n63392,
    n63393, n63394, n63395, n63396, n63397, n63398, n63399, n63400, n63401,
    n63402, n63403, n63404, n63405, n63406, n63407, n63408, n63409, n63410,
    n63411, n63412, n63413, n63414, n63415, n63416, n63417, n63418, n63419,
    n63420, n63421, n63422, n63423, n63424, n63425, n63426, n63427, n63428,
    n63429, n63430, n63431, n63432, n63433, n63434, n63435, n63436, n63437,
    n63438, n63439, n63440, n63441, n63442, n63443, n63444, n63445, n63446,
    n63447, n63448, n63449, n63450, n63451, n63452, n63453, n63454, n63455,
    n63456, n63457, n63458, n63459, n63460, n63461, n63462, n63463, n63464,
    n63465, n63466, n63467, n63468, n63469, n63470, n63471, n63472, n63473,
    n63474, n63475, n63476, n63477, n63478, n63479, n63480, n63481, n63482,
    n63483, n63484, n63485, n63486, n63487, n63488, n63489, n63490, n63491,
    n63492, n63493, n63494, n63495, n63496, n63497, n63498, n63499, n63500,
    n63501, n63502, n63503, n63504, n63505, n63506, n63507, n63508, n63509,
    n63510, n63511, n63512, n63513, n63514, n63515, n63516, n63517, n63518,
    n63519, n63520, n63521, n63522, n63523, n63524, n63525, n63526, n63527,
    n63528, n63529, n63530, n63531, n63532, n63533, n63534, n63535, n63536,
    n63537, n63538, n63539, n63540, n63541, n63542, n63543, n63544, n63545,
    n63546, n63547, n63548, n63549, n63550, n63551, n63552, n63553, n63554,
    n63555, n63556, n63557, n63558, n63559, n63560, n63561, n63562, n63563,
    n63564, n63565, n63566, n63567, n63568, n63569, n63570, n63571, n63572,
    n63573, n63574, n63575, n63576, n63577, n63578, n63579, n63580, n63581,
    n63582, n63583, n63584, n63585, n63586, n63587, n63588, n63589, n63590,
    n63591, n63592, n63593, n63594, n63595, n63596, n63597, n63598, n63599,
    n63600, n63601, n63602, n63603, n63604, n63605, n63606, n63607, n63608,
    n63609, n63610, n63611, n63612, n63613, n63614, n63615, n63616, n63617,
    n63618, n63619, n63620, n63621, n63622, n63623, n63624, n63625, n63626,
    n63627, n63628, n63629, n63630, n63631, n63632, n63633, n63634, n63635,
    n63636, n63637, n63638, n63639, n63640, n63641, n63642, n63643, n63644,
    n63645, n63646, n63647, n63648, n63649, n63650, n63651, n63652, n63653,
    n63654, n63655, n63656, n63657, n63658, n63659, n63660, n63661, n63662,
    n63663, n63664, n63665, n63666, n63667, n63668, n63669, n63670, n63671,
    n63672, n63673, n63674, n63675, n63676, n63677, n63678, n63679, n63680,
    n63681, n63682, n63683, n63684, n63685, n63686, n63687, n63688, n63689,
    n63690, n63691, n63692, n63693, n63694, n63695, n63696, n63697, n63698,
    n63699, n63700, n63701, n63702, n63703, n63704, n63705, n63706, n63707,
    n63708, n63709, n63710, n63711, n63712, n63713, n63714, n63715, n63716,
    n63717, n63718, n63719, n63720, n63721, n63722, n63723, n63724, n63725,
    n63726, n63727, n63728, n63729, n63730, n63731, n63732, n63733, n63734,
    n63735, n63736, n63737, n63738, n63739, n63740, n63741, n63742, n63743,
    n63744, n63745, n63746, n63747, n63748, n63749, n63750, n63751, n63752,
    n63753, n63754, n63755, n63756, n63757, n63758, n63759, n63760, n63761,
    n63762, n63763, n63764, n63765, n63766, n63767, n63768, n63769, n63770,
    n63771, n63772, n63773, n63774, n63775, n63776, n63777, n63778, n63779,
    n63780, n63781, n63782, n63783, n63784, n63785, n63786, n63787, n63788,
    n63789, n63790, n63791, n63792, n63793, n63794, n63795, n63796, n63797,
    n63798, n63799, n63800, n63801, n63802, n63803, n63804, n63805, n63806,
    n63807, n63808, n63809, n63810, n63811, n63812, n63813, n63814, n63815,
    n63816, n63817, n63818, n63819, n63820, n63821, n63822, n63823, n63824,
    n63825, n63826, n63827, n63828, n63829, n63830, n63831, n63832, n63833,
    n63834, n63835, n63836, n63837, n63838, n63839, n63840, n63841, n63842,
    n63843, n63844, n63845, n63846, n63847, n63848, n63849, n63850, n63851,
    n63852, n63853, n63854, n63855, n63856, n63857, n63858, n63859, n63860,
    n63861, n63862, n63863, n63864, n63865, n63866, n63867, n63868, n63869,
    n63870, n63871, n63872, n63873, n63874, n63875, n63876, n63877, n63878,
    n63879, n63880, n63881, n63882, n63883, n63884, n63885, n63886, n63887,
    n63888, n63889, n63890, n63891, n63892, n63893, n63894, n63895, n63896,
    n63897, n63898, n63899, n63900, n63901, n63902, n63903, n63904, n63905,
    n63906, n63907, n63908, n63909, n63910, n63911, n63912, n63913, n63914,
    n63915, n63916, n63917, n63918, n63919, n63920, n63921, n63922, n63923,
    n63924, n63925, n63926, n63927, n63928, n63929, n63930, n63931, n63932,
    n63933, n63934, n63935, n63936, n63937, n63938, n63939, n63940, n63941,
    n63942, n63943, n63944, n63945, n63946, n63947, n63948, n63949, n63950,
    n63951, n63952, n63953, n63954, n63955, n63956, n63957, n63958, n63959,
    n63960, n63961, n63962, n63963, n63964, n63965, n63966, n63967, n63968,
    n63969, n63970, n63971, n63972, n63973, n63974, n63975, n63976, n63977,
    n63978, n63979, n63980, n63981, n63982, n63983, n63984, n63985, n63986,
    n63987, n63988, n63989, n63990, n63991, n63992, n63993, n63994, n63995,
    n63996, n63997, n63998, n63999, n64000, n64001, n64002, n64003, n64004,
    n64005, n64006, n64007, n64008, n64009, n64010, n64011, n64012, n64013,
    n64014, n64015, n64016, n64017, n64018, n64019, n64020, n64021, n64022,
    n64023, n64024, n64025, n64026, n64027, n64028, n64029, n64030, n64031,
    n64032, n64033, n64034, n64035, n64036, n64037, n64038, n64039, n64040,
    n64041, n64042, n64043, n64044, n64045, n64046, n64047, n64048, n64049,
    n64050, n64051, n64052, n64053, n64054, n64055, n64056, n64057, n64058,
    n64059, n64060, n64061, n64062, n64063, n64064, n64065, n64066, n64067,
    n64068, n64069, n64070, n64071, n64072, n64073, n64074, n64075, n64076,
    n64077, n64078, n64079, n64080, n64081, n64082, n64083, n64084, n64085,
    n64086, n64087, n64088, n64089, n64090, n64091, n64092, n64093, n64094,
    n64095, n64096, n64097, n64098, n64099, n64100, n64101, n64102, n64103,
    n64104, n64105, n64106, n64107, n64108, n64109, n64110, n64111, n64112,
    n64113, n64114, n64115, n64116, n64117, n64118, n64119, n64120, n64121,
    n64122, n64123, n64124, n64125, n64126, n64127, n64128, n64129, n64130,
    n64131, n64132, n64133, n64134, n64135, n64136, n64137, n64138, n64139,
    n64140, n64141, n64142, n64143, n64144, n64145, n64146, n64147, n64148,
    n64149, n64150, n64151, n64152, n64153, n64154, n64155, n64156, n64157,
    n64158, n64159, n64160, n64161, n64162, n64163, n64164, n64165, n64166,
    n64167, n64168, n64169, n64170, n64171, n64172, n64173, n64174, n64175,
    n64176, n64177, n64178, n64179, n64180, n64181, n64182, n64183, n64184,
    n64185, n64186, n64187, n64188, n64189, n64190, n64191, n64192, n64193,
    n64194, n64195, n64196, n64197, n64198, n64199, n64200, n64201, n64202,
    n64203, n64204, n64205, n64206, n64207, n64208, n64209, n64210, n64211,
    n64212, n64213, n64214, n64215, n64216, n64217, n64218, n64219, n64220,
    n64221, n64222, n64223, n64224, n64225, n64226, n64227, n64228, n64229,
    n64230, n64231, n64232, n64233, n64234, n64235, n64236, n64237, n64238,
    n64239, n64240, n64241, n64242, n64243, n64244, n64245, n64246, n64247,
    n64248, n64249, n64250, n64251, n64252, n64253, n64254, n64255, n64256,
    n64257, n64258, n64259, n64260, n64261, n64262, n64263, n64264, n64265,
    n64266, n64267, n64268, n64269, n64270, n64271, n64272, n64273, n64274,
    n64275, n64276, n64277, n64278, n64279, n64280, n64281, n64282, n64283,
    n64284, n64285, n64286, n64287, n64288, n64289, n64290, n64291, n64292,
    n64293, n64294, n64295, n64296, n64297, n64298, n64299, n64300, n64301,
    n64302, n64303, n64304, n64305, n64306, n64307, n64308, n64309, n64310,
    n64311, n64312, n64313, n64314, n64315, n64316, n64317, n64318, n64319,
    n64320, n64321, n64322, n64323, n64324, n64325, n64326, n64327, n64328,
    n64329, n64330, n64331, n64332, n64333, n64334, n64335, n64336, n64337,
    n64338, n64339, n64340, n64341, n64342, n64343, n64344, n64345, n64346,
    n64347, n64348, n64349, n64350, n64351, n64352, n64353, n64354, n64355,
    n64356, n64357, n64358, n64359, n64360, n64361, n64362, n64363, n64364,
    n64365, n64366, n64367, n64368, n64369, n64370, n64371, n64372, n64373,
    n64374, n64375, n64376, n64377, n64378, n64379, n64380, n64381, n64382,
    n64383, n64384, n64385, n64386, n64387, n64388, n64389, n64390, n64391,
    n64392, n64393, n64394, n64395, n64396, n64397, n64398, n64399, n64400,
    n64401, n64402, n64403, n64404, n64405, n64406, n64407, n64408, n64409,
    n64410, n64411, n64412, n64413, n64414, n64415, n64416, n64417, n64418,
    n64419, n64420, n64421, n64422, n64423, n64424, n64425, n64426, n64427,
    n64428, n64429, n64430, n64431, n64432, n64433, n64434, n64435, n64436,
    n64437, n64438, n64439, n64440, n64441, n64442, n64443, n64444, n64445,
    n64446, n64447, n64448, n64449, n64450, n64451, n64452, n64453, n64454,
    n64455, n64456, n64457, n64458, n64459, n64460, n64461, n64462, n64463,
    n64464, n64465, n64466, n64467, n64468, n64469, n64470, n64471, n64472,
    n64473, n64474, n64475, n64476, n64477, n64478, n64479, n64480, n64481,
    n64482, n64483, n64484, n64485, n64486, n64487, n64488, n64489, n64490,
    n64491, n64492, n64493, n64494, n64495, n64496, n64497, n64498, n64499,
    n64500, n64501, n64502, n64503, n64504, n64505, n64506, n64507, n64508,
    n64509, n64510, n64511, n64512, n64513, n64514, n64515, n64516, n64517,
    n64518, n64519, n64520, n64521, n64522, n64523, n64524, n64525, n64526,
    n64527, n64528, n64529, n64530, n64531, n64532, n64533, n64534, n64535,
    n64536, n64537, n64538, n64539, n64540, n64541, n64542, n64543, n64544,
    n64545, n64546, n64547, n64548, n64549, n64550, n64551, n64552, n64553,
    n64554, n64555, n64556, n64557, n64558, n64559, n64560, n64561, n64562,
    n64563, n64564, n64565, n64566, n64567, n64568, n64569, n64570, n64571,
    n64572, n64573, n64574, n64575, n64576, n64577, n64578, n64579, n64580,
    n64581, n64582, n64583, n64584, n64585, n64586, n64587, n64588, n64589,
    n64590, n64591, n64592, n64593, n64594, n64595, n64596, n64597, n64598,
    n64599, n64600, n64601, n64602, n64603, n64604, n64605, n64606, n64607,
    n64608, n64609, n64610, n64611, n64612, n64613, n64614, n64615, n64616,
    n64617, n64618, n64619, n64620, n64621, n64622, n64623, n64624, n64625,
    n64626, n64627, n64628, n64629, n64630, n64631, n64632, n64633, n64634,
    n64635, n64636, n64637, n64638, n64639, n64640, n64641, n64642, n64643,
    n64644, n64645, n64646, n64647, n64648, n64649, n64650, n64651, n64652,
    n64653, n64654, n64655, n64656, n64657, n64658, n64659, n64660, n64661,
    n64662, n64663, n64664, n64665, n64666, n64667, n64668, n64669, n64670,
    n64671, n64672, n64673, n64674, n64675, n64676, n64677, n64678, n64679,
    n64680, n64681, n64682, n64683, n64684, n64685, n64686, n64687, n64688,
    n64689, n64690, n64691, n64692, n64693, n64694, n64695, n64696, n64697,
    n64698, n64699, n64700, n64701, n64702, n64703, n64704, n64705, n64706,
    n64707, n64708, n64709, n64710, n64711, n64712, n64713, n64714, n64715,
    n64716, n64717, n64718, n64719, n64720, n64721, n64722, n64723, n64724,
    n64725, n64726, n64727, n64728, n64729, n64730, n64731, n64732, n64733,
    n64734, n64735, n64736, n64737, n64738, n64739, n64740, n64741, n64742,
    n64743, n64744, n64745, n64746, n64747, n64748, n64749, n64750, n64751,
    n64752, n64753, n64754, n64755, n64756, n64757, n64758, n64759, n64760,
    n64761, n64762, n64763, n64764, n64765, n64766, n64767, n64768, n64769,
    n64770, n64771, n64772, n64773, n64774, n64775, n64776, n64777, n64778,
    n64779, n64780, n64781, n64782, n64783, n64784, n64785, n64786, n64787,
    n64788, n64789, n64790, n64791, n64792, n64793, n64794, n64795, n64796,
    n64797, n64798, n64799, n64800, n64801, n64802, n64803, n64804, n64805,
    n64806, n64807, n64808, n64809, n64810, n64811, n64812, n64813, n64814,
    n64815, n64816, n64817, n64818, n64819, n64820, n64821, n64822, n64823,
    n64824, n64825, n64826, n64827, n64828, n64829, n64830, n64831, n64832,
    n64833, n64834, n64835, n64836, n64837, n64838, n64839, n64840, n64841,
    n64842, n64843, n64844, n64845, n64846, n64847, n64848, n64849, n64850,
    n64851, n64852, n64853, n64854, n64855, n64856, n64857, n64858, n64859,
    n64860, n64861, n64862, n64863, n64864, n64865, n64866, n64867, n64868,
    n64869, n64870, n64871, n64872, n64873, n64874, n64875, n64876, n64877,
    n64878, n64879, n64880, n64881, n64882, n64883, n64884, n64885, n64886,
    n64887, n64888, n64889, n64890, n64891, n64892, n64893, n64894, n64895,
    n64896, n64897, n64898, n64899, n64900, n64901, n64902, n64903, n64904,
    n64905, n64906, n64907, n64908, n64909, n64910, n64911, n64912, n64913,
    n64914, n64915, n64916, n64917, n64918, n64919, n64920, n64921, n64922,
    n64923, n64924, n64925, n64926, n64927, n64928, n64929, n64930, n64931,
    n64932, n64933, n64934, n64935, n64936, n64937, n64938, n64939, n64940,
    n64941, n64942, n64943, n64944, n64945, n64946, n64947, n64948, n64949,
    n64950, n64951, n64952, n64953, n64954, n64955, n64956, n64957, n64958,
    n64959, n64960, n64961, n64962, n64963, n64964, n64965, n64966, n64967,
    n64968, n64969, n64970, n64971, n64972, n64973, n64974, n64975, n64976,
    n64977, n64978, n64979, n64980, n64981, n64982, n64983, n64984, n64985,
    n64986, n64987, n64988, n64989, n64990, n64991, n64992, n64993, n64994,
    n64995, n64996, n64997, n64998, n64999, n65000, n65001, n65002, n65003,
    n65004, n65005, n65006, n65007, n65008, n65009, n65010, n65011, n65012,
    n65013, n65014, n65015, n65016, n65017, n65018, n65019, n65020, n65021,
    n65022, n65023, n65024, n65025, n65026, n65027, n65028, n65029, n65030,
    n65031, n65032, n65033, n65034, n65035, n65036, n65037, n65038, n65039,
    n65040, n65041, n65042, n65043, n65044, n65045, n65046, n65047, n65048,
    n65049, n65050, n65051, n65052, n65053, n65054, n65055, n65056, n65057,
    n65058, n65059, n65060, n65061, n65062, n65063, n65064, n65065, n65066,
    n65067, n65068, n65069, n65070, n65071, n65072, n65073, n65074, n65075,
    n65076, n65077, n65078, n65079, n65080, n65081, n65082, n65083, n65084,
    n65085, n65086, n65087, n65088, n65089, n65090, n65091, n65092, n65093,
    n65094, n65095, n65096, n65097, n65098, n65099, n65100, n65101, n65102,
    n65103, n65104, n65105, n65106, n65107, n65108, n65109, n65110, n65111,
    n65112, n65113, n65114, n65115, n65116, n65117, n65118, n65119, n65120,
    n65121, n65122, n65123, n65124, n65125, n65126, n65127, n65128, n65129,
    n65130, n65131, n65132, n65133, n65134, n65135, n65136, n65137, n65138,
    n65139, n65140, n65141, n65142, n65143, n65144, n65145, n65146, n65147,
    n65148, n65149, n65150, n65151, n65152, n65153, n65154, n65155, n65156,
    n65157, n65158, n65159, n65160, n65161, n65162, n65163, n65164, n65165,
    n65166, n65167, n65168, n65169, n65170, n65171, n65172, n65173, n65174,
    n65175, n65176, n65177, n65178, n65179, n65180, n65181, n65182, n65183,
    n65184, n65185, n65186, n65187, n65188, n65189, n65190, n65191, n65192,
    n65193, n65194, n65195, n65196, n65197, n65198, n65199, n65200, n65201,
    n65202, n65203, n65204, n65205, n65206, n65207, n65208, n65209, n65210,
    n65211, n65212, n65213, n65214, n65215, n65216, n65217, n65218, n65219,
    n65220, n65221, n65222, n65223, n65224, n65225, n65226, n65227, n65228,
    n65229, n65230, n65231, n65232, n65233, n65234, n65235, n65236, n65237,
    n65238, n65239, n65240, n65241, n65242, n65243, n65244, n65245, n65246,
    n65247, n65248, n65249, n65250, n65251, n65252, n65253, n65254, n65255,
    n65256, n65257, n65258, n65259, n65260, n65261, n65262, n65263, n65264,
    n65265, n65266, n65267, n65268, n65269, n65270, n65271, n65272, n65273,
    n65274, n65275, n65276, n65277, n65278, n65279, n65280, n65281, n65282,
    n65283, n65284, n65285, n65286, n65287, n65288, n65289, n65290, n65291,
    n65292, n65293, n65294, n65295, n65296, n65297, n65298, n65299, n65300,
    n65301, n65302, n65303, n65304, n65305, n65306, n65307, n65308, n65309,
    n65310, n65311, n65312, n65313, n65314, n65315, n65316, n65317, n65318,
    n65319, n65320, n65321, n65322, n65323, n65324, n65325, n65326, n65327,
    n65328, n65329, n65330, n65331, n65332, n65333, n65334, n65335, n65336,
    n65337, n65338, n65339, n65340, n65341, n65342, n65343, n65344, n65345,
    n65346, n65347, n65348, n65349, n65350, n65351, n65352, n65353, n65354,
    n65355, n65356, n65357, n65358, n65359, n65360, n65361, n65362, n65363,
    n65364, n65365, n65366, n65367, n65368, n65369, n65370, n65371, n65372,
    n65373, n65374, n65375, n65376, n65377, n65378, n65379, n65380, n65381,
    n65382, n65383, n65384, n65385, n65386, n65387, n65388, n65389, n65390,
    n65391, n65392, n65393, n65394, n65395, n65396, n65397, n65398, n65399,
    n65400, n65401, n65402, n65403, n65404, n65405, n65406, n65407, n65408,
    n65409, n65410, n65411, n65412, n65413, n65414, n65415, n65416, n65417,
    n65418, n65419, n65420, n65421, n65422, n65423, n65424, n65425, n65426,
    n65427, n65428, n65429, n65430, n65431, n65432, n65433, n65434, n65435,
    n65436, n65437, n65438, n65439, n65440, n65441, n65442, n65443, n65444,
    n65445, n65446, n65447, n65448, n65449, n65450, n65451, n65452, n65453,
    n65454, n65455, n65456, n65457, n65458, n65459, n65460, n65461, n65462,
    n65463, n65464, n65465, n65466, n65467, n65468, n65469, n65470, n65471,
    n65472, n65473, n65474, n65475, n65476, n65477, n65478, n65479, n65480,
    n65481, n65482, n65483, n65484, n65485, n65486, n65487, n65488, n65489,
    n65490, n65491, n65492, n65493, n65494, n65495, n65496, n65497, n65498,
    n65499, n65500, n65501, n65502, n65503, n65504, n65505, n65506, n65507,
    n65508, n65509, n65510, n65511, n65512, n65513, n65514, n65515, n65516,
    n65517, n65518, n65519, n65520, n65521, n65522, n65523, n65524, n65525,
    n65526, n65527, n65528, n65529, n65530, n65531, n65532, n65533, n65534,
    n65535, n65536, n65537, n65538, n65539, n65540, n65541, n65542, n65543,
    n65544, n65545, n65546, n65547, n65548, n65549, n65550, n65551, n65552,
    n65553, n65554, n65555, n65556, n65557, n65558, n65559, n65560, n65561,
    n65562, n65563, n65564, n65565, n65566, n65567, n65568, n65569, n65570,
    n65571, n65572, n65573, n65574, n65575, n65576, n65577, n65578, n65579,
    n65580, n65581, n65582, n65583, n65584, n65585, n65586, n65587, n65588,
    n65589, n65590, n65591, n65592, n65593, n65594, n65595, n65596, n65597,
    n65598, n65599, n65600, n65601, n65602, n65603, n65604, n65605, n65606,
    n65607, n65608, n65609, n65610, n65611, n65612, n65613, n65614, n65615,
    n65616, n65617, n65618, n65619, n65620, n65621, n65622, n65623, n65624,
    n65625, n65626, n65627, n65628, n65629, n65630, n65631, n65632, n65633,
    n65634, n65635, n65636, n65637, n65638, n65639, n65640, n65641, n65642,
    n65643, n65644, n65645, n65646, n65647, n65648, n65649, n65650, n65651,
    n65652, n65653, n65654, n65655, n65656, n65657, n65658, n65659, n65660,
    n65661, n65662, n65663, n65664, n65665, n65666, n65667, n65668, n65669,
    n65670, n65671, n65672, n65673, n65674, n65675, n65676, n65677, n65678,
    n65679, n65680, n65681, n65682, n65683, n65684, n65685, n65686, n65687,
    n65688, n65689, n65690, n65691, n65692, n65693, n65694, n65695, n65696,
    n65697, n65698, n65699, n65700, n65701, n65702, n65703, n65704, n65705,
    n65706, n65707, n65708, n65709, n65710, n65711, n65712, n65713, n65714,
    n65715, n65716, n65717, n65718, n65719, n65720, n65721, n65722, n65723,
    n65724, n65725, n65726, n65727, n65728, n65729, n65730, n65731, n65732,
    n65733, n65734, n65735, n65736, n65737, n65738, n65739, n65740, n65741,
    n65742, n65743, n65744, n65745, n65746, n65747, n65748, n65749, n65750,
    n65751, n65752, n65753, n65754, n65755, n65756, n65757, n65758, n65759,
    n65760, n65761, n65762, n65763, n65764, n65765, n65766, n65767, n65768,
    n65769, n65770, n65771, n65772, n65773, n65774, n65775, n65776, n65777,
    n65778, n65779, n65780, n65781, n65782, n65783, n65784, n65785, n65786,
    n65787, n65788, n65789, n65790, n65791, n65792, n65793, n65794, n65795,
    n65796, n65797, n65798, n65799, n65800, n65801, n65802, n65803, n65804,
    n65805, n65806, n65807, n65808, n65809, n65810, n65811, n65812, n65813,
    n65814, n65815, n65816, n65817, n65818, n65819, n65820, n65821, n65822,
    n65823, n65824, n65825, n65826, n65827, n65828, n65829, n65830, n65831,
    n65832, n65833, n65834, n65835, n65836, n65837, n65838, n65839, n65840,
    n65841, n65842, n65843, n65844, n65845, n65846, n65847, n65848, n65849,
    n65850, n65851, n65852, n65853, n65854, n65855, n65856, n65857, n65858,
    n65859, n65860, n65861, n65862, n65863, n65864, n65865, n65866, n65867,
    n65868, n65869, n65870, n65871, n65872, n65873, n65874, n65875, n65876,
    n65877, n65878, n65879, n65880, n65881, n65882, n65883, n65884, n65885,
    n65886, n65887, n65888, n65889, n65890, n65891, n65892, n65893, n65894,
    n65895, n65896, n65897, n65898, n65899, n65900, n65901, n65902, n65903,
    n65904, n65905, n65906, n65907, n65908, n65909, n65910, n65911, n65912,
    n65913, n65914, n65915, n65916, n65917, n65918, n65919, n65920, n65921,
    n65922, n65923, n65924, n65925, n65926, n65927, n65928, n65929, n65930,
    n65931, n65932, n65933, n65934, n65935, n65936, n65937, n65938, n65939,
    n65940, n65941, n65942, n65943, n65944, n65945, n65946, n65947, n65948,
    n65949, n65950, n65951, n65952, n65953, n65954, n65955, n65956, n65957,
    n65958, n65959, n65960, n65961, n65962, n65963, n65964, n65965, n65966,
    n65967, n65968, n65969, n65970, n65971, n65972, n65973, n65974, n65975,
    n65976, n65977, n65978, n65979, n65980, n65981, n65982, n65983, n65984,
    n65985, n65986, n65987, n65988, n65989, n65990, n65991, n65992, n65993,
    n65994, n65995, n65996, n65997, n65998, n65999, n66000, n66001, n66002,
    n66003, n66004, n66005, n66006, n66007, n66008, n66009, n66010, n66011,
    n66012, n66013, n66014, n66015, n66016, n66017, n66018, n66019, n66020,
    n66021, n66022, n66023, n66024, n66025, n66026, n66027, n66028, n66029,
    n66030, n66031, n66032, n66033, n66034, n66035, n66036, n66037, n66038,
    n66039, n66040, n66041, n66042, n66043, n66044, n66045, n66046, n66047,
    n66048, n66049, n66050, n66051, n66052, n66053, n66054, n66055, n66056,
    n66057, n66058, n66059, n66060, n66061, n66062, n66063, n66064, n66065,
    n66066, n66067, n66068, n66069, n66070, n66071, n66072, n66073, n66074,
    n66075, n66076, n66077, n66078, n66079, n66080, n66081, n66082, n66083,
    n66084, n66085, n66086, n66087, n66088, n66089, n66090, n66091, n66092,
    n66093, n66094, n66095, n66096, n66097, n66098, n66099, n66100, n66101,
    n66102, n66103, n66104, n66105, n66106, n66107, n66108, n66109, n66110,
    n66111, n66112, n66113, n66114, n66115, n66116, n66117, n66118, n66119,
    n66120, n66121, n66122, n66123, n66124, n66125, n66126, n66127, n66128,
    n66129, n66130, n66131, n66132, n66133, n66134, n66135, n66136, n66137,
    n66138, n66139, n66140, n66141, n66142, n66143, n66144, n66145, n66146,
    n66147, n66148, n66149, n66150, n66151, n66152, n66153, n66154, n66155,
    n66156, n66157, n66158, n66159, n66160, n66161, n66162, n66163, n66164,
    n66165, n66166, n66167, n66168, n66169, n66170, n66171, n66172, n66173,
    n66174, n66175, n66176, n66177, n66178, n66179, n66180, n66181, n66182,
    n66183, n66184, n66185, n66186, n66187, n66188, n66189, n66190, n66191,
    n66192, n66193, n66194, n66195, n66196, n66197, n66198, n66199, n66200,
    n66201, n66202, n66203, n66204, n66205, n66206, n66207, n66208, n66209,
    n66210, n66211, n66212, n66213, n66214, n66215, n66216, n66217, n66218,
    n66219, n66220, n66221, n66222, n66223, n66224, n66225, n66226, n66227,
    n66228, n66229, n66230, n66231, n66232, n66233, n66234, n66235, n66236,
    n66237, n66238, n66239, n66240, n66241, n66242, n66243, n66244, n66245,
    n66246, n66247, n66248, n66249, n66250, n66251, n66252, n66253, n66254,
    n66255, n66256, n66257, n66258, n66259, n66260, n66261, n66262, n66263,
    n66264, n66265, n66266, n66267, n66268, n66269, n66270, n66271, n66272,
    n66273, n66274, n66275, n66276, n66277, n66278, n66279, n66280, n66281,
    n66282, n66283, n66284, n66285, n66286, n66287, n66288, n66289, n66290,
    n66291, n66292, n66293, n66294, n66295, n66296, n66297, n66298, n66299,
    n66300, n66301, n66302, n66303, n66304, n66305, n66306, n66307, n66308,
    n66309, n66310, n66311, n66312, n66313, n66314, n66315, n66316, n66317,
    n66318, n66319, n66320, n66321, n66322, n66323, n66324, n66325, n66326,
    n66327, n66328, n66329, n66330, n66331, n66332, n66333, n66334, n66335,
    n66336, n66337, n66338, n66339, n66340, n66341, n66342, n66343, n66344,
    n66345, n66346, n66347, n66348, n66349, n66350, n66351, n66352, n66353,
    n66354, n66355, n66356, n66357, n66358, n66359, n66360, n66361, n66362,
    n66363, n66364, n66365, n66366, n66367, n66368, n66369, n66370, n66371,
    n66372, n66373, n66374, n66375, n66376, n66377, n66378, n66379, n66380,
    n66381, n66382, n66383, n66384, n66385, n66386, n66387, n66388, n66389,
    n66390, n66391, n66392, n66393, n66394, n66395, n66396, n66397, n66398,
    n66399, n66400, n66401, n66402, n66403, n66404, n66405, n66406, n66407,
    n66408, n66409, n66410, n66411, n66412, n66413, n66414, n66415, n66416,
    n66417, n66418, n66419, n66420, n66421, n66422, n66423, n66424, n66425,
    n66426, n66427, n66428, n66429, n66430, n66431, n66432, n66433, n66434,
    n66435, n66436, n66437, n66438, n66439, n66440, n66441, n66442, n66443,
    n66444, n66445, n66446, n66447, n66448, n66449, n66450, n66451, n66452,
    n66453, n66454, n66455, n66456, n66457, n66458, n66459, n66460, n66461,
    n66462, n66463, n66464, n66465, n66466, n66467, n66468, n66469, n66470,
    n66471, n66472, n66473, n66474, n66475, n66476, n66477, n66478, n66479,
    n66480, n66481, n66482, n66483, n66484, n66485, n66486, n66487, n66488,
    n66489, n66490, n66491, n66492, n66493, n66494, n66495, n66496, n66497,
    n66498, n66499, n66500, n66501, n66502, n66503, n66504, n66505, n66506,
    n66507, n66508, n66509, n66510, n66511, n66512, n66513, n66514, n66515,
    n66516, n66517, n66518, n66519, n66520, n66521, n66522, n66523, n66524,
    n66525, n66526, n66527, n66528, n66529, n66530, n66531, n66532, n66533,
    n66534, n66535, n66536, n66537, n66538, n66539, n66540, n66541, n66542,
    n66543, n66544, n66545, n66546, n66547, n66548, n66549, n66550, n66551,
    n66552, n66553, n66554, n66555, n66556, n66557, n66558, n66559, n66560,
    n66561, n66562, n66563, n66564, n66565, n66566, n66567, n66568, n66569,
    n66570, n66571, n66572, n66573, n66574, n66575, n66576, n66577, n66578,
    n66579, n66580, n66581, n66582, n66583, n66584, n66585, n66586, n66587,
    n66588, n66589, n66590, n66591, n66592, n66593, n66594, n66595, n66596,
    n66597, n66598, n66599, n66600, n66601, n66602, n66603, n66604, n66605,
    n66606, n66607, n66608, n66609, n66610, n66611, n66612, n66613, n66614,
    n66615, n66616, n66617, n66618, n66619, n66620, n66621, n66622, n66623,
    n66624, n66625, n66626, n66627, n66628, n66629, n66630, n66631, n66632,
    n66633, n66634, n66635, n66636, n66637, n66638, n66639, n66640, n66641,
    n66642, n66643, n66644, n66645, n66646, n66647, n66648, n66649, n66650,
    n66651, n66652, n66653, n66654, n66655, n66656, n66657, n66658, n66659,
    n66660, n66661, n66662, n66663, n66664, n66665, n66666, n66667, n66668,
    n66669, n66670, n66671, n66672, n66673, n66674, n66675, n66676, n66677,
    n66678, n66679, n66680, n66681, n66682, n66683, n66684, n66685, n66686,
    n66687, n66688, n66689, n66690, n66691, n66692, n66693, n66694, n66695,
    n66696, n66697, n66698, n66699, n66700, n66701, n66702, n66703, n66704,
    n66705, n66706, n66707, n66708, n66709, n66710, n66711, n66712, n66713,
    n66714, n66715, n66716, n66717, n66718, n66719, n66720, n66721, n66722,
    n66723, n66724, n66725, n66726, n66727, n66728, n66729, n66730, n66731,
    n66732, n66733, n66734, n66735, n66736, n66737, n66738, n66739, n66740,
    n66741, n66742, n66743, n66744, n66745, n66746, n66747, n66748, n66749,
    n66750, n66751, n66752, n66753, n66754, n66755, n66756, n66757, n66758,
    n66759, n66760, n66761, n66762, n66763, n66764, n66765, n66766, n66767,
    n66768, n66769, n66770, n66771, n66772, n66773, n66774, n66775, n66776,
    n66777, n66778, n66779, n66780, n66781, n66782, n66783, n66784, n66785,
    n66786, n66787, n66788, n66789, n66790, n66791, n66792, n66793, n66794,
    n66795, n66796, n66797, n66798, n66799, n66800, n66801, n66802, n66803,
    n66804, n66805, n66806, n66807, n66808, n66809, n66810, n66811, n66812,
    n66813, n66814, n66815, n66816, n66817, n66818, n66819, n66820, n66821,
    n66822, n66823, n66824, n66825, n66826, n66827, n66828, n66829, n66830,
    n66831, n66832, n66833, n66834, n66835, n66836, n66837, n66838, n66839,
    n66840, n66841, n66842, n66843, n66844, n66845, n66846, n66847, n66848,
    n66849, n66850, n66851, n66852, n66853, n66854, n66855, n66856, n66857,
    n66858, n66859, n66860, n66861, n66862, n66863, n66864, n66865, n66866,
    n66867, n66868, n66869, n66870, n66871, n66872, n66873, n66874, n66875,
    n66876, n66877, n66878, n66879, n66880, n66881, n66882, n66883, n66884,
    n66885, n66886, n66887, n66888, n66889, n66890, n66891, n66892, n66893,
    n66894, n66895, n66896, n66897, n66898, n66899, n66900, n66901, n66902,
    n66903, n66904, n66905, n66906, n66907, n66908, n66909, n66910, n66911,
    n66912, n66913, n66914, n66915, n66916, n66917, n66918, n66919, n66920,
    n66921, n66922, n66923, n66924, n66925, n66926, n66927, n66928, n66929,
    n66930, n66931, n66932, n66933, n66934, n66935, n66936, n66937, n66938,
    n66939, n66940, n66941, n66942, n66943, n66944, n66945, n66946, n66947,
    n66948, n66949, n66950, n66951, n66952, n66953, n66954, n66955, n66956,
    n66957, n66958, n66959, n66960, n66961, n66962, n66963, n66964, n66965,
    n66966, n66967, n66968, n66969, n66970, n66971, n66972, n66973, n66974,
    n66975, n66976, n66977, n66978, n66979, n66980, n66981, n66982, n66983,
    n66984, n66985, n66986, n66987, n66988, n66989, n66990, n66991, n66992,
    n66993, n66994, n66995, n66996, n66997, n66998, n66999, n67000, n67001,
    n67002, n67003, n67004, n67005, n67006, n67007, n67008, n67009, n67010,
    n67011, n67012, n67013, n67014, n67015, n67016, n67017, n67018, n67019,
    n67020, n67021, n67022, n67023, n67024, n67025, n67026, n67027, n67028,
    n67029, n67030, n67031, n67032, n67033, n67034, n67035, n67036, n67037,
    n67038, n67039, n67040, n67041, n67042, n67043, n67044, n67045, n67046,
    n67047, n67048, n67049, n67050, n67051, n67052, n67053, n67054, n67055,
    n67056, n67057, n67058, n67059, n67060, n67061, n67062, n67063, n67064,
    n67065, n67066, n67067, n67068, n67069, n67070, n67071, n67072, n67073,
    n67074, n67075, n67076, n67077, n67078, n67079, n67080, n67081, n67082,
    n67083, n67084, n67085, n67086, n67087, n67088, n67089, n67090, n67091,
    n67092, n67093, n67094, n67095, n67096, n67097, n67098, n67099, n67100,
    n67101, n67102, n67103, n67104, n67105, n67106, n67107, n67108, n67109,
    n67110, n67111, n67112, n67113, n67114, n67115, n67116, n67117, n67118,
    n67119, n67120, n67121, n67122, n67123, n67124, n67125, n67126, n67127,
    n67128, n67129, n67130, n67131, n67132, n67133, n67134, n67135, n67136,
    n67137, n67138, n67139, n67140, n67141, n67142, n67143, n67144, n67145,
    n67146, n67147, n67148, n67149, n67150, n67151, n67152, n67153, n67154,
    n67155, n67156, n67157, n67158, n67159, n67160, n67161, n67162, n67163,
    n67164, n67165, n67166, n67167, n67168, n67169, n67170, n67171, n67172,
    n67173, n67174, n67175, n67176, n67177, n67178, n67179, n67180, n67181,
    n67182, n67183, n67184, n67185, n67186, n67187, n67188, n67189, n67190,
    n67191, n67192, n67193, n67194, n67195, n67196, n67197, n67198, n67199,
    n67200, n67201, n67202, n67203, n67204, n67205, n67206, n67207, n67208,
    n67209, n67210, n67211, n67212, n67213, n67214, n67215, n67216, n67217,
    n67218, n67219, n67220, n67221, n67222, n67223, n67224, n67225, n67226,
    n67227, n67228, n67229, n67230, n67231, n67232, n67233, n67234, n67235,
    n67236, n67237, n67238, n67239, n67240, n67241, n67242, n67243, n67244,
    n67245, n67246, n67247, n67248, n67249, n67250, n67251, n67252, n67253,
    n67254, n67255, n67256, n67257, n67258, n67259, n67260, n67261, n67262,
    n67263, n67264, n67265, n67266, n67267, n67268, n67269, n67270, n67271,
    n67272, n67273, n67274, n67275, n67276, n67277, n67278, n67279, n67280,
    n67281, n67282, n67283, n67284, n67285, n67286, n67287, n67288, n67289,
    n67290, n67291, n67292, n67293, n67294, n67295, n67296, n67297, n67298,
    n67299, n67300, n67301, n67302, n67303, n67304, n67305, n67306, n67307,
    n67308, n67309, n67310, n67311, n67312, n67313, n67314, n67315, n67316,
    n67317, n67318, n67319, n67320, n67321, n67322, n67323, n67324, n67325,
    n67326, n67327, n67328, n67329, n67330, n67331, n67332, n67333, n67334,
    n67335, n67336, n67337, n67338, n67339, n67340, n67341, n67342, n67343,
    n67344, n67345, n67346, n67347, n67348, n67349, n67350, n67351, n67352,
    n67353, n67354, n67355, n67356, n67357, n67358, n67359, n67360, n67361,
    n67362, n67363, n67364, n67365, n67366, n67367, n67368, n67369, n67370,
    n67371, n67372, n67373, n67374, n67375, n67376, n67377, n67378, n67379,
    n67380, n67381, n67382, n67383, n67384, n67385, n67386, n67387, n67388,
    n67389, n67390, n67391, n67392, n67393, n67394, n67395, n67396, n67397,
    n67398, n67399, n67400, n67401, n67402, n67403, n67404, n67405, n67406,
    n67407, n67408, n67409, n67410, n67411, n67412, n67413, n67414, n67415,
    n67416, n67417, n67418, n67419, n67420, n67421, n67422, n67423, n67424,
    n67425, n67426, n67427, n67428, n67429, n67430, n67431, n67432, n67433,
    n67434, n67435, n67436, n67437, n67438, n67439, n67440, n67441, n67442,
    n67443, n67444, n67445, n67446, n67447, n67448, n67449, n67450, n67451,
    n67452, n67453, n67454, n67455, n67456, n67457, n67458, n67459, n67460,
    n67461, n67462, n67463, n67464, n67465, n67466, n67467, n67468, n67469,
    n67470, n67471, n67472, n67473, n67474, n67475, n67476, n67477, n67478,
    n67479, n67480, n67481, n67482, n67483, n67484, n67485, n67486, n67487,
    n67488, n67489, n67490, n67491, n67492, n67493, n67494, n67495, n67496,
    n67497, n67498, n67499, n67500, n67501, n67502, n67503, n67504, n67505,
    n67506, n67507, n67508, n67509, n67510, n67511, n67512, n67513, n67514,
    n67515, n67516, n67517, n67518, n67519, n67520, n67521, n67522, n67523,
    n67524, n67525, n67526, n67527, n67528, n67529, n67530, n67531, n67532,
    n67533, n67534, n67535, n67536, n67537, n67538, n67539, n67540, n67541,
    n67542, n67543, n67544, n67545, n67546, n67547, n67548, n67549, n67550,
    n67551, n67552, n67553, n67554, n67555, n67556, n67557, n67558, n67559,
    n67560, n67561, n67562, n67563, n67564, n67565, n67566, n67567, n67568,
    n67569, n67570, n67571, n67572, n67573, n67574, n67575, n67576, n67577,
    n67578, n67579, n67580, n67581, n67582, n67583, n67584, n67585, n67586,
    n67587, n67588, n67589, n67590, n67591, n67592, n67593, n67594, n67595,
    n67596, n67597, n67598, n67599, n67600, n67601, n67602, n67603, n67604,
    n67605, n67606, n67607, n67608, n67609, n67610, n67611, n67612, n67613,
    n67614, n67615, n67616, n67617, n67618, n67619, n67620, n67621, n67622,
    n67623, n67624, n67625, n67626, n67627, n67628, n67629, n67630, n67631,
    n67632, n67633, n67634, n67635, n67636, n67637, n67638, n67639, n67640,
    n67641, n67642, n67643, n67644, n67645, n67646, n67647, n67648, n67649,
    n67650, n67651, n67652, n67653, n67654, n67655, n67656, n67657, n67658,
    n67659, n67660, n67661, n67662, n67663, n67664, n67665, n67666, n67667,
    n67668, n67669, n67670, n67671, n67672, n67673, n67674, n67675, n67676,
    n67677, n67678, n67679, n67680, n67681, n67682, n67683, n67684, n67685,
    n67686, n67687, n67688, n67689, n67690, n67691, n67692, n67693, n67694,
    n67695, n67696, n67697, n67698, n67699, n67700, n67701, n67702, n67703,
    n67704, n67705, n67706, n67707, n67708, n67709, n67710, n67711, n67712,
    n67713, n67714, n67715, n67716, n67717, n67718, n67719, n67720, n67721,
    n67722, n67723, n67724, n67725, n67726, n67727, n67728, n67729, n67730,
    n67731, n67732, n67733, n67734, n67735, n67736, n67737, n67738, n67739,
    n67740, n67741, n67742, n67743, n67744, n67745, n67746, n67747, n67748,
    n67749, n67750, n67751, n67752, n67753, n67754, n67755, n67756, n67757,
    n67758, n67759, n67760, n67761, n67762, n67763, n67764, n67765, n67766,
    n67767, n67768, n67769, n67770, n67771, n67772, n67773, n67774, n67775,
    n67776, n67777, n67778, n67779, n67780, n67781, n67782, n67783, n67784,
    n67785, n67786, n67787, n67788, n67789, n67790, n67791, n67792, n67793,
    n67794, n67795, n67796, n67797, n67798, n67799, n67800, n67801, n67802,
    n67803, n67804, n67805, n67806, n67807, n67808, n67809, n67810, n67811,
    n67812, n67813, n67814, n67815, n67816, n67817, n67818, n67819, n67820,
    n67821, n67822, n67823, n67824, n67825, n67826, n67827, n67828, n67829,
    n67830, n67831, n67832, n67833, n67834, n67835, n67836, n67837, n67838,
    n67839, n67840, n67841, n67842, n67843, n67844, n67845, n67846, n67847,
    n67848, n67849, n67850, n67851, n67852, n67853, n67854, n67855, n67856,
    n67857, n67858, n67859, n67860, n67861, n67862, n67863, n67864, n67865,
    n67866, n67867, n67868, n67869, n67870, n67871, n67872, n67873, n67874,
    n67875, n67876, n67877, n67878, n67879, n67880, n67881, n67882, n67883,
    n67884, n67885, n67886, n67887, n67888, n67889, n67890, n67891, n67892,
    n67893, n67894, n67895, n67896, n67897, n67898, n67899, n67900, n67901,
    n67902, n67903, n67904, n67905, n67906, n67907, n67908, n67909, n67910,
    n67911, n67912, n67913, n67914, n67915, n67916, n67917, n67918, n67919,
    n67920, n67921, n67922, n67923, n67924, n67925, n67926, n67927, n67928,
    n67929, n67930, n67931, n67932, n67933, n67934, n67935, n67936, n67937,
    n67938, n67939, n67940, n67941, n67942, n67943, n67944, n67945, n67946,
    n67947, n67948, n67949, n67950, n67951, n67952, n67953, n67954, n67955,
    n67956, n67957, n67958, n67959, n67960, n67961, n67962, n67963, n67964,
    n67965, n67966, n67967, n67968, n67969, n67970, n67971, n67972, n67973,
    n67974, n67975, n67976, n67977, n67978, n67979, n67980, n67981, n67982,
    n67983, n67984, n67985, n67986, n67987, n67988, n67989, n67990, n67991,
    n67992, n67993, n67994, n67995, n67996, n67997, n67998, n67999, n68000,
    n68001, n68002, n68003, n68004, n68005, n68006, n68007, n68008, n68009,
    n68010, n68011, n68012, n68013, n68014, n68015, n68016, n68017, n68018,
    n68019, n68020, n68021, n68022, n68023, n68024, n68025, n68026, n68027,
    n68028, n68029, n68030, n68031, n68032, n68033, n68034, n68035, n68036,
    n68037, n68038, n68039, n68040, n68041, n68042, n68043, n68044, n68045,
    n68046, n68047, n68048, n68049, n68050, n68051, n68052, n68053, n68054,
    n68055, n68056, n68057, n68058, n68059, n68060, n68061, n68062, n68063,
    n68064, n68065, n68066, n68067, n68068, n68069, n68070, n68071, n68072,
    n68073, n68074, n68075, n68076, n68077, n68078, n68079, n68080, n68081,
    n68082, n68083, n68084, n68085, n68086, n68087, n68088, n68089, n68090,
    n68091, n68092, n68093, n68094, n68095, n68096, n68097, n68098, n68099,
    n68100, n68101, n68102, n68103, n68104, n68105, n68106, n68107, n68108,
    n68109, n68110, n68111, n68112, n68113, n68114, n68115, n68116, n68117,
    n68118, n68119, n68120, n68121, n68122, n68123, n68124, n68125, n68126,
    n68127, n68128, n68129, n68130, n68131, n68132, n68133, n68134, n68135,
    n68136, n68137, n68138, n68139, n68140, n68141, n68142, n68143, n68144,
    n68145, n68146, n68147, n68148, n68149, n68150, n68151, n68152, n68153,
    n68154, n68155, n68156, n68157, n68158, n68159, n68160, n68161, n68162,
    n68163, n68164, n68165, n68166, n68167, n68168, n68169, n68170, n68171,
    n68172, n68173, n68174, n68175, n68176, n68177, n68178, n68179, n68180,
    n68181, n68182, n68183, n68184, n68185, n68186, n68187, n68188, n68189,
    n68190, n68191, n68192, n68193, n68194, n68195, n68196, n68197, n68198,
    n68199, n68200, n68201, n68202, n68203, n68204, n68205, n68206, n68207,
    n68208, n68209, n68210, n68211, n68212, n68213, n68214, n68215, n68216,
    n68217, n68218, n68219, n68220, n68221, n68222, n68223, n68224, n68225,
    n68226, n68227, n68228, n68229, n68230, n68231, n68232, n68233, n68234,
    n68235, n68236, n68237, n68238, n68239, n68240, n68241, n68242, n68243,
    n68244, n68245, n68246, n68247, n68248, n68249, n68250, n68251, n68252,
    n68253, n68254, n68255, n68256, n68257, n68258, n68259, n68260, n68261,
    n68262, n68263, n68264, n68265, n68266, n68267, n68268, n68269, n68270,
    n68271, n68272, n68273, n68274, n68275, n68276, n68277, n68278, n68279,
    n68280, n68281, n68282, n68283, n68284, n68285, n68286, n68287, n68288,
    n68289, n68290, n68291, n68292, n68293, n68294, n68295, n68296, n68297,
    n68298, n68299, n68300, n68301, n68302, n68303, n68304, n68305, n68306,
    n68307, n68308, n68309, n68310, n68311, n68312, n68313, n68314, n68315,
    n68316, n68317, n68318, n68319, n68320, n68321, n68322, n68323, n68324,
    n68325, n68326, n68327, n68328, n68329, n68330, n68331, n68332, n68333,
    n68334, n68335, n68336, n68337, n68338, n68339, n68340, n68341, n68342,
    n68343, n68344, n68345, n68346, n68347, n68348, n68349, n68350, n68351,
    n68352, n68353, n68354, n68355, n68356, n68357, n68358, n68359, n68360,
    n68361, n68362, n68363, n68364, n68365, n68366, n68367, n68368, n68369,
    n68370, n68371, n68372, n68373, n68374, n68375, n68376, n68377, n68378,
    n68379, n68380, n68381, n68382, n68383, n68384, n68385, n68386, n68387,
    n68388, n68389, n68390, n68391, n68392, n68393, n68394, n68395, n68396,
    n68397, n68398, n68399, n68400, n68401, n68402, n68403, n68404, n68405,
    n68406, n68407, n68408, n68409, n68410, n68411, n68412, n68413, n68414,
    n68415, n68416, n68417, n68418, n68419, n68420, n68421, n68422, n68423,
    n68424, n68425, n68426, n68427, n68428, n68429, n68430, n68431, n68432,
    n68433, n68434, n68435, n68436, n68437, n68438, n68439, n68440, n68441,
    n68442, n68443, n68444, n68445, n68446, n68447, n68448, n68449, n68450,
    n68451, n68452, n68453, n68454, n68455, n68456, n68457, n68458, n68459,
    n68460, n68461, n68462, n68463, n68464, n68465, n68466, n68467, n68468,
    n68469, n68470, n68471, n68472, n68473, n68474, n68475, n68476, n68477,
    n68478, n68479, n68480, n68481, n68482, n68483, n68484, n68485, n68486,
    n68487, n68488, n68489, n68490, n68491, n68492, n68493, n68494, n68495,
    n68496, n68497, n68498, n68499, n68500, n68501, n68502, n68503, n68504,
    n68505, n68506, n68507, n68508, n68509, n68510, n68511, n68512, n68513,
    n68514, n68515, n68516, n68517, n68518, n68519, n68520, n68521, n68522,
    n68523, n68524, n68525, n68526, n68527, n68528, n68529, n68530, n68531,
    n68532, n68533, n68534, n68535, n68536, n68537, n68538, n68539, n68540,
    n68541, n68542, n68543, n68544, n68545, n68546, n68547, n68548, n68549,
    n68550, n68551, n68552, n68553, n68554, n68555, n68556, n68557, n68558,
    n68559, n68560, n68561, n68562, n68563, n68564, n68565, n68566, n68567,
    n68568, n68569, n68570, n68571, n68572, n68573, n68574, n68575, n68576,
    n68577, n68578, n68579, n68580, n68581, n68582, n68583, n68584, n68585,
    n68586, n68587, n68588, n68589, n68590, n68591, n68592, n68593, n68594,
    n68595, n68596, n68597, n68598, n68599, n68600, n68601, n68602, n68603,
    n68604, n68605, n68606, n68607, n68608, n68609, n68610, n68611, n68612,
    n68613, n68614, n68615, n68616, n68617, n68618, n68619, n68620, n68621,
    n68622, n68623, n68624, n68625, n68626, n68627, n68628, n68629, n68630,
    n68631, n68632, n68633, n68634, n68635, n68636, n68637, n68638, n68639,
    n68640, n68641, n68642, n68643, n68644, n68645, n68646, n68647, n68648,
    n68649, n68650, n68651, n68652, n68653, n68654, n68655, n68656, n68657,
    n68658, n68659, n68660, n68661, n68662, n68663, n68664, n68665, n68666,
    n68667, n68668, n68669, n68670, n68671, n68672, n68673, n68674, n68675,
    n68676, n68677, n68678, n68679, n68680, n68681, n68682, n68683, n68684,
    n68685, n68686, n68687, n68688, n68689, n68690, n68691, n68692, n68693,
    n68694, n68695, n68696, n68697, n68698, n68699, n68700, n68701, n68702,
    n68703, n68704, n68705, n68706, n68707, n68708, n68709, n68710, n68711,
    n68712, n68713, n68714, n68715, n68716, n68717, n68718, n68719, n68720,
    n68721, n68722, n68723, n68724, n68725, n68726, n68727, n68728, n68729,
    n68730, n68731, n68732, n68733, n68734, n68735, n68736, n68737, n68738,
    n68739, n68740, n68741, n68742, n68743, n68744, n68745, n68746, n68747,
    n68748, n68749, n68750, n68751, n68752, n68753, n68754, n68755, n68756,
    n68757, n68758, n68759, n68760, n68761, n68762, n68763, n68764, n68765,
    n68766, n68767, n68768, n68769, n68770, n68771, n68772, n68773, n68774,
    n68775, n68776, n68777, n68778, n68779, n68780, n68781, n68782, n68783,
    n68784, n68785, n68786, n68787, n68788, n68789, n68790, n68791, n68792,
    n68793, n68794, n68795, n68796, n68797, n68798, n68799, n68800, n68801,
    n68802, n68803, n68804, n68805, n68806, n68807, n68808, n68809, n68810,
    n68811, n68812, n68813, n68814, n68815, n68816, n68817, n68818, n68819,
    n68820, n68821, n68822, n68823, n68824, n68825, n68826, n68827, n68828,
    n68829, n68830, n68831, n68832, n68833, n68834, n68835, n68836, n68837,
    n68838, n68839, n68840, n68841, n68842, n68843, n68844, n68845, n68846,
    n68847, n68848, n68849, n68850, n68851, n68852, n68853, n68854, n68855,
    n68856, n68857, n68858, n68859, n68860, n68861, n68862, n68863, n68864,
    n68865, n68866, n68867, n68868, n68869, n68870, n68871, n68872, n68873,
    n68874, n68875, n68876, n68877, n68878, n68879, n68880, n68881, n68882,
    n68883, n68884, n68885, n68886, n68887, n68888, n68889, n68890, n68891,
    n68892, n68893, n68894, n68895, n68896, n68897, n68898, n68899, n68900,
    n68901, n68902, n68903, n68904, n68905, n68906, n68907, n68908, n68909,
    n68910, n68911, n68912, n68913, n68914, n68915, n68916, n68917, n68918,
    n68919, n68920, n68921, n68922, n68923, n68924, n68925, n68926, n68927,
    n68928, n68929, n68930, n68931, n68932, n68933, n68934, n68935, n68936,
    n68937, n68938, n68939, n68940, n68941, n68942, n68943, n68944, n68945,
    n68946, n68947, n68948, n68949, n68950, n68951, n68952, n68953, n68954,
    n68955, n68956, n68957, n68958, n68959, n68960, n68961, n68962, n68963,
    n68964, n68965, n68966, n68967, n68968, n68969, n68970, n68971, n68972,
    n68973, n68974, n68975, n68976, n68977, n68978, n68979, n68980, n68981,
    n68982, n68983, n68984, n68985, n68986, n68987, n68988, n68989, n68990,
    n68991, n68992, n68993, n68994, n68995, n68996, n68997, n68998, n68999,
    n69000, n69001, n69002, n69003, n69004, n69005, n69006, n69007, n69008,
    n69009, n69010, n69011, n69012, n69013, n69014, n69015, n69016, n69017,
    n69018, n69019, n69020, n69021, n69022, n69023, n69024, n69025, n69026,
    n69027, n69028, n69029, n69030, n69031, n69032, n69033, n69034, n69035,
    n69036, n69037, n69038, n69039, n69040, n69041, n69042, n69043, n69044,
    n69045, n69046, n69047, n69048, n69049, n69050, n69051, n69052, n69053,
    n69054, n69055, n69056, n69057, n69058, n69059, n69060, n69061, n69062,
    n69063, n69064, n69065, n69066, n69067, n69068, n69069, n69070, n69071,
    n69072, n69073, n69074, n69075, n69076, n69077, n69078, n69079, n69080,
    n69081, n69082, n69083, n69084, n69085, n69086, n69087, n69088, n69089,
    n69090, n69091, n69092, n69093, n69094, n69095, n69096, n69097, n69098,
    n69099, n69100, n69101, n69102, n69103, n69104, n69105, n69106, n69107,
    n69108, n69109, n69110, n69111, n69112, n69113, n69114, n69115, n69116,
    n69117, n69118, n69119, n69120, n69121, n69122, n69123, n69124, n69125,
    n69126, n69127, n69128, n69129, n69130, n69131, n69132, n69133, n69134,
    n69135, n69136, n69137, n69138, n69139, n69140, n69141, n69142, n69143,
    n69144, n69145, n69146, n69147, n69148, n69149, n69150, n69151, n69152,
    n69153, n69154, n69155, n69156, n69157, n69158, n69159, n69160, n69161,
    n69162, n69163, n69164, n69165, n69166, n69167, n69168, n69169, n69170,
    n69171, n69172, n69173, n69174, n69175, n69176, n69177, n69178, n69179,
    n69180, n69181, n69182, n69183, n69184, n69185, n69186, n69187, n69188,
    n69189, n69190, n69191, n69192, n69193, n69194, n69195, n69196, n69197,
    n69198, n69199, n69200, n69201, n69202, n69203, n69204, n69205, n69206,
    n69207, n69208, n69209, n69210, n69211, n69212, n69213, n69214, n69215,
    n69216, n69217, n69218, n69219, n69220, n69221, n69222, n69223, n69224,
    n69225, n69226, n69227, n69228, n69229, n69230, n69231, n69232, n69233,
    n69234, n69235, n69236, n69237, n69238, n69239, n69240, n69241, n69242,
    n69243, n69244, n69245, n69246, n69247, n69248, n69249, n69250, n69251,
    n69252, n69253, n69254, n69255, n69256, n69257, n69258, n69259, n69260,
    n69261, n69262, n69263, n69264, n69265, n69266, n69267, n69268, n69269,
    n69270, n69271, n69272, n69273, n69274, n69275, n69276, n69277, n69278,
    n69279, n69280, n69281, n69282, n69283, n69284, n69285, n69286, n69287,
    n69288, n69289, n69290, n69291, n69292, n69293, n69294, n69295, n69296,
    n69297, n69298, n69299, n69300, n69301, n69302, n69303, n69304, n69305,
    n69306, n69307, n69308, n69309, n69310, n69311, n69312, n69313, n69314,
    n69315, n69316, n69317, n69318, n69319, n69320, n69321, n69322, n69323,
    n69324, n69325, n69326, n69327, n69328, n69329, n69330, n69331, n69332,
    n69333, n69334, n69335, n69336, n69337, n69338, n69339, n69340, n69341,
    n69342, n69343, n69344, n69345, n69346, n69347, n69348, n69349, n69350,
    n69351, n69352, n69353, n69354, n69355, n69356, n69357, n69358, n69359,
    n69360, n69361, n69362, n69363, n69364, n69365, n69366, n69367, n69368,
    n69369, n69370, n69371, n69372, n69373, n69374, n69375, n69376, n69377,
    n69378, n69379, n69380, n69381, n69382, n69383, n69384, n69385, n69386,
    n69387, n69388, n69389, n69390, n69391, n69392, n69393, n69394, n69395,
    n69396, n69397, n69398, n69399, n69400, n69401, n69402, n69403, n69404,
    n69405, n69406, n69407, n69408, n69409, n69410, n69411, n69412, n69413,
    n69414, n69415, n69416, n69417, n69418, n69419, n69420, n69421, n69422,
    n69423, n69424, n69425, n69426, n69427, n69428, n69429, n69430, n69431,
    n69432, n69433, n69434, n69435, n69436, n69437, n69438, n69439, n69440,
    n69441, n69442, n69443, n69444, n69445, n69446, n69447, n69448, n69449,
    n69450, n69451, n69452, n69453, n69454, n69455, n69456, n69457, n69458,
    n69459, n69460, n69461, n69462, n69463, n69464, n69465, n69466, n69467,
    n69468, n69469, n69470, n69471, n69472, n69473, n69474, n69475, n69476,
    n69477, n69478, n69479, n69480, n69481, n69482, n69483, n69484, n69485,
    n69486, n69487, n69488, n69489, n69490, n69491, n69492, n69493, n69494,
    n69495, n69496, n69497, n69498, n69499, n69500, n69501, n69502, n69503,
    n69504, n69505, n69506, n69507, n69508, n69509, n69510, n69511, n69512,
    n69513, n69514, n69515, n69516, n69517, n69518, n69519, n69520, n69521,
    n69522, n69523, n69524, n69525, n69526, n69527, n69528, n69529, n69530,
    n69531, n69532, n69533, n69534, n69535, n69536, n69537, n69538, n69539,
    n69540, n69541, n69542, n69543, n69544, n69545, n69546, n69547, n69548,
    n69549, n69550, n69551, n69552, n69553, n69554, n69555, n69556, n69557,
    n69558, n69559, n69560, n69561, n69562, n69563, n69564, n69565, n69566,
    n69567, n69568, n69569, n69570, n69571, n69572, n69573, n69574, n69575,
    n69576, n69577, n69578, n69579, n69580, n69581, n69582, n69583, n69584,
    n69585, n69586, n69587, n69588, n69589, n69590, n69591, n69592, n69593,
    n69594, n69595, n69596, n69597, n69598, n69599, n69600, n69601, n69602,
    n69603, n69604, n69605, n69606, n69607, n69608, n69609, n69610, n69611,
    n69612, n69613, n69614, n69615, n69616, n69617, n69618, n69619, n69620,
    n69621, n69622, n69623, n69624, n69625, n69626, n69627, n69628, n69629,
    n69630, n69631, n69632, n69633, n69634, n69635, n69636, n69637, n69638,
    n69639, n69640, n69641, n69642, n69643, n69644, n69645, n69646, n69647,
    n69648, n69649, n69650, n69651, n69652, n69653, n69654, n69655, n69656,
    n69657, n69658, n69659, n69660, n69661, n69662, n69663, n69664, n69665,
    n69666, n69667, n69668, n69669, n69670, n69671, n69672, n69673, n69674,
    n69675, n69676, n69677, n69678, n69679, n69680, n69681, n69682, n69683,
    n69684, n69685, n69686, n69687, n69688, n69689, n69690, n69691, n69692,
    n69693, n69694, n69695, n69696, n69697, n69698, n69699, n69700, n69701,
    n69702, n69703, n69704, n69705, n69706, n69707, n69708, n69709, n69710,
    n69711, n69712, n69713, n69714, n69715, n69716, n69717, n69718, n69719,
    n69720, n69721, n69722, n69723, n69724, n69725, n69726, n69727, n69728,
    n69729, n69730, n69731, n69732, n69733, n69734, n69735, n69736, n69737,
    n69738, n69739, n69740, n69741, n69742, n69743, n69744, n69745, n69746,
    n69747, n69748, n69749, n69750, n69751, n69752, n69753, n69754, n69755,
    n69756, n69757, n69758, n69759, n69760, n69761, n69762, n69763, n69764,
    n69765, n69766, n69767, n69768, n69769, n69770, n69771, n69772, n69773,
    n69774, n69775, n69776, n69777, n69778, n69779, n69780, n69781, n69782,
    n69783, n69784, n69785, n69786, n69787, n69788, n69789, n69790, n69791,
    n69792, n69793, n69794, n69795, n69796, n69797, n69798, n69799, n69800,
    n69801, n69802, n69803, n69804, n69805, n69806, n69807, n69808, n69809,
    n69810, n69811, n69812, n69813, n69814, n69815, n69816, n69817, n69818,
    n69819, n69820, n69821, n69822, n69823, n69824, n69825, n69826, n69827,
    n69828, n69829, n69830, n69831, n69832, n69833, n69834, n69835, n69836,
    n69837, n69838, n69839, n69840, n69841, n69842, n69843, n69844, n69845,
    n69846, n69847, n69848, n69849, n69850, n69851, n69852, n69853, n69854,
    n69855, n69856, n69857, n69858, n69859, n69860, n69861, n69862, n69863,
    n69864, n69865, n69866, n69867, n69868, n69869, n69870, n69871, n69872,
    n69873, n69874, n69875, n69876, n69877, n69878, n69879, n69880, n69881,
    n69882, n69883, n69884, n69885, n69886, n69887, n69888, n69889, n69890,
    n69891, n69892, n69893, n69894, n69895, n69896, n69897, n69898, n69899,
    n69900, n69901, n69902, n69903, n69904, n69905, n69906, n69907, n69908,
    n69909, n69910, n69911, n69912, n69913, n69914, n69915, n69916, n69917,
    n69918, n69919, n69920, n69921, n69922, n69923, n69924, n69925, n69926,
    n69927, n69928, n69929, n69930, n69931, n69932, n69933, n69934, n69935,
    n69936, n69937, n69938, n69939, n69940, n69941, n69942, n69943, n69944,
    n69945, n69946, n69947, n69948, n69949, n69950, n69951, n69952, n69953,
    n69954, n69955, n69956, n69957, n69958, n69959, n69960, n69961, n69962,
    n69963, n69964, n69965, n69966, n69967, n69968, n69969, n69970, n69971,
    n69972, n69973, n69974, n69975, n69976, n69977, n69978, n69979, n69980,
    n69981, n69982, n69983, n69984, n69985, n69986, n69987, n69988, n69989,
    n69990, n69991, n69992, n69993, n69994, n69995, n69996, n69997, n69998,
    n69999, n70000, n70001, n70002, n70003, n70004, n70005, n70006, n70007,
    n70008, n70009, n70010, n70011, n70012, n70013, n70014, n70015, n70016,
    n70017, n70018, n70019, n70020, n70021, n70022, n70023, n70024, n70025,
    n70026, n70027, n70028, n70029, n70030, n70031, n70032, n70033, n70034,
    n70035, n70036, n70037, n70038, n70039, n70040, n70041, n70042, n70043,
    n70044, n70045, n70046, n70047, n70048, n70049, n70050, n70051, n70052,
    n70053, n70054, n70055, n70056, n70057, n70058, n70059, n70060, n70061,
    n70062, n70063, n70064, n70065, n70066, n70067, n70068, n70069, n70070,
    n70071, n70072, n70073, n70074, n70075, n70076, n70077, n70078, n70079,
    n70080, n70081, n70082, n70083, n70084, n70085, n70086, n70087, n70088,
    n70089, n70090, n70091, n70092, n70093, n70094, n70095, n70096, n70097,
    n70098, n70099, n70100, n70101, n70102, n70103, n70104, n70105, n70106,
    n70107, n70108, n70109, n70110, n70111, n70112, n70113, n70114, n70115,
    n70116, n70117, n70118, n70119, n70120, n70121, n70122, n70123, n70124,
    n70125, n70126, n70127, n70128, n70129, n70130, n70131, n70132, n70133,
    n70134, n70135, n70136, n70137, n70138, n70139, n70140, n70141, n70142,
    n70143, n70144, n70145, n70146, n70147, n70148, n70149, n70150, n70151,
    n70152, n70153, n70154, n70155, n70156, n70157, n70158, n70159, n70160,
    n70161, n70162, n70163, n70164, n70165, n70166, n70167, n70168, n70169,
    n70170, n70171, n70172, n70173, n70174, n70175, n70176, n70177, n70178,
    n70179, n70180, n70181, n70182, n70183, n70184, n70185, n70186, n70187,
    n70188, n70189, n70190, n70191, n70192, n70193, n70194, n70195, n70196,
    n70197, n70198, n70199, n70200, n70201, n70202, n70203, n70204, n70205,
    n70206, n70207, n70208, n70209, n70210, n70211, n70212, n70213, n70214,
    n70215, n70216, n70217, n70218, n70219, n70220, n70221, n70222, n70223,
    n70224, n70225, n70226, n70227, n70228, n70229, n70230, n70231, n70232,
    n70233, n70234, n70235, n70236, n70237, n70238, n70239, n70240, n70241,
    n70242, n70243, n70244, n70245, n70246, n70247, n70248, n70249, n70250,
    n70251, n70252, n70253, n70254, n70255, n70256, n70257, n70258, n70259,
    n70260, n70261, n70262, n70263, n70264, n70265, n70266, n70267, n70268,
    n70269, n70270, n70271, n70272, n70273, n70274, n70275, n70276, n70277,
    n70278, n70279, n70280, n70281, n70282, n70283, n70284, n70285, n70286,
    n70287, n70288, n70289, n70290, n70291, n70292, n70293, n70294, n70295,
    n70296, n70297, n70298, n70299, n70300, n70301, n70302, n70303, n70304,
    n70305, n70306, n70307, n70308, n70309, n70310, n70311, n70312, n70313,
    n70314, n70315, n70316, n70317, n70318, n70319, n70320, n70321, n70322,
    n70323, n70324, n70325, n70326, n70327, n70328, n70329, n70330, n70331,
    n70332, n70333, n70334, n70335, n70336, n70337, n70338, n70339, n70340,
    n70341, n70342, n70343, n70344, n70345, n70346, n70347, n70348, n70349,
    n70350, n70351, n70352, n70353, n70354, n70355, n70356, n70357, n70358,
    n70359, n70360, n70361, n70362, n70363, n70364, n70365, n70366, n70367,
    n70368, n70369, n70370, n70371, n70372, n70373, n70374, n70375, n70376,
    n70377, n70378, n70379, n70380, n70381, n70382, n70383, n70384, n70385,
    n70386, n70387, n70388, n70389, n70390, n70391, n70392, n70393, n70394,
    n70395, n70396, n70397, n70398, n70399, n70400, n70401, n70402, n70403,
    n70404, n70405, n70406, n70407, n70408, n70409, n70410, n70411, n70412,
    n70413, n70414, n70415, n70416, n70417, n70418, n70419, n70420, n70421,
    n70422, n70423, n70424, n70425, n70426, n70427, n70428, n70429, n70430,
    n70431, n70432, n70433, n70434, n70435, n70436, n70437, n70438, n70439,
    n70440, n70441, n70442, n70443, n70444, n70445, n70446, n70447, n70448,
    n70449, n70450, n70451, n70452, n70453, n70454, n70455, n70456, n70457,
    n70458, n70459, n70460, n70461, n70462, n70463, n70464, n70465, n70466,
    n70467, n70468, n70469, n70470, n70471, n70472, n70473, n70474, n70475,
    n70476, n70477, n70478, n70479, n70480, n70481, n70482, n70483, n70484,
    n70485, n70486, n70487, n70488, n70489, n70490, n70491, n70492, n70493,
    n70494, n70495, n70496, n70497, n70498, n70499, n70500, n70501, n70502,
    n70503, n70504, n70505, n70506, n70507, n70508, n70509, n70510, n70511,
    n70512, n70513, n70514, n70515, n70516, n70517, n70518, n70519, n70520,
    n70521, n70522, n70523, n70524, n70525, n70526, n70527, n70528, n70529,
    n70530, n70531, n70532, n70533, n70534, n70535, n70536, n70537, n70538,
    n70539, n70540, n70541, n70542, n70543, n70544, n70545, n70546, n70547,
    n70548, n70549, n70550, n70551, n70552, n70553, n70554, n70555, n70556,
    n70557, n70558, n70559, n70560, n70561, n70562, n70563, n70564, n70565,
    n70566, n70567, n70568, n70569, n70570, n70571, n70572, n70573, n70574,
    n70575, n70576, n70577, n70578, n70579, n70580, n70581, n70582, n70583,
    n70584, n70585, n70586, n70587, n70588, n70589, n70590, n70591, n70592,
    n70593, n70594, n70595, n70596, n70597, n70598, n70599, n70600, n70601,
    n70602, n70603, n70604, n70605, n70606, n70607, n70608, n70609, n70610,
    n70611, n70612, n70613, n70614, n70615, n70616, n70617, n70618, n70619,
    n70620, n70621, n70622, n70623, n70624, n70625, n70626, n70627, n70628,
    n70629, n70630, n70631, n70632, n70633, n70634, n70635, n70636, n70637,
    n70638, n70639, n70640, n70641, n70642, n70643, n70644, n70645, n70646,
    n70647, n70648, n70649, n70650, n70651, n70652, n70653, n70654, n70655,
    n70656, n70657, n70658, n70659, n70660, n70661, n70662, n70663, n70664,
    n70665, n70666, n70667, n70668, n70669, n70670, n70671, n70672, n70673,
    n70674, n70675, n70676, n70677, n70678, n70679, n70680, n70681, n70682,
    n70683, n70684, n70685, n70686, n70687, n70688, n70689, n70690, n70691,
    n70692, n70693, n70694, n70695, n70696, n70697, n70698, n70699, n70700,
    n70701, n70702, n70703, n70704, n70705, n70706, n70707, n70708, n70709,
    n70710, n70711, n70712, n70713, n70714, n70715, n70716, n70717, n70718,
    n70719, n70720, n70721, n70722, n70723, n70724, n70725, n70726, n70727,
    n70728, n70729, n70730, n70731, n70732, n70733, n70734, n70735, n70736,
    n70737, n70738, n70739, n70740, n70741, n70742, n70743, n70744, n70745,
    n70746, n70747, n70748, n70749, n70750, n70751, n70752, n70753, n70754,
    n70755, n70756, n70757, n70758, n70759, n70760, n70761, n70762, n70763,
    n70764, n70765, n70766, n70767, n70768, n70769, n70770, n70771, n70772,
    n70773, n70774, n70775, n70776, n70777, n70778, n70779, n70780, n70781,
    n70782, n70783, n70784, n70785, n70786, n70787, n70788, n70789, n70790,
    n70791, n70792, n70793, n70794, n70795, n70796, n70797, n70798, n70799,
    n70800, n70801, n70802, n70803, n70804, n70805, n70806, n70807, n70808,
    n70809, n70810, n70811, n70812, n70813, n70814, n70815, n70816, n70817,
    n70818, n70819, n70820, n70821, n70822, n70823, n70824, n70825, n70826,
    n70827, n70828, n70829, n70830, n70831, n70832, n70833, n70834, n70835,
    n70836, n70837, n70838, n70839, n70840, n70841, n70842, n70843, n70844,
    n70845, n70846, n70847, n70848, n70849, n70850, n70851, n70852, n70853,
    n70854, n70855, n70856, n70857, n70858, n70859, n70860, n70861, n70862,
    n70863, n70864, n70865, n70866, n70867, n70868, n70869, n70870, n70871,
    n70872, n70873, n70874, n70875, n70876, n70877, n70878, n70879, n70880,
    n70881, n70882, n70883, n70884, n70885, n70886, n70887, n70888, n70889,
    n70890, n70891, n70892, n70893, n70894, n70895, n70896, n70897, n70898,
    n70899, n70900, n70901, n70902, n70903, n70904, n70905, n70906, n70907,
    n70908, n70909, n70910, n70911, n70912, n70913, n70914, n70915, n70916,
    n70917, n70918, n70919, n70920, n70921, n70922, n70923, n70924, n70925,
    n70926, n70927, n70928, n70929, n70930, n70931, n70932, n70933, n70934,
    n70935, n70936, n70937, n70938, n70939, n70940, n70941, n70942, n70943,
    n70944, n70945, n70946, n70947, n70948, n70949, n70950, n70951, n70952,
    n70953, n70954, n70955, n70956, n70957, n70958, n70959, n70960, n70961,
    n70962, n70963, n70964, n70965, n70966, n70967, n70968, n70969, n70970,
    n70971, n70972, n70973, n70974, n70975, n70976, n70977, n70978, n70979,
    n70980, n70981, n70982, n70983, n70984, n70985, n70986, n70987, n70988,
    n70989, n70990, n70991, n70992, n70993, n70994, n70995, n70996, n70997,
    n70998, n70999, n71000, n71001, n71002, n71003, n71004, n71005, n71006,
    n71007, n71008, n71009, n71010, n71011, n71012, n71013, n71014, n71015,
    n71016, n71017, n71018, n71019, n71020, n71021, n71022, n71023, n71024,
    n71025, n71026, n71027, n71028, n71029, n71030, n71031, n71032, n71033,
    n71034, n71035, n71036, n71037, n71038, n71039, n71040, n71041, n71042,
    n71043, n71044, n71045, n71046, n71047, n71048, n71049, n71050, n71051,
    n71052, n71053, n71054, n71055, n71056, n71057, n71058, n71059, n71060,
    n71061, n71062, n71063, n71064, n71065, n71066, n71067, n71068, n71069,
    n71070, n71071, n71072, n71073, n71074, n71075, n71076, n71077, n71078,
    n71079, n71080, n71081, n71082, n71083, n71084, n71085, n71086, n71087,
    n71088, n71089, n71090, n71091, n71092, n71093, n71094, n71095, n71096,
    n71097, n71098, n71099, n71100, n71101, n71102, n71103, n71104, n71105,
    n71106, n71107, n71108, n71109, n71110, n71111, n71112, n71113, n71114,
    n71115, n71116, n71117, n71118, n71119, n71120, n71121, n71122, n71123,
    n71124, n71125, n71126, n71127, n71128, n71129, n71130, n71131, n71132,
    n71133, n71134, n71135, n71136, n71137, n71138, n71139, n71140, n71141,
    n71142, n71143, n71144, n71145, n71146, n71147, n71148, n71149, n71150,
    n71151, n71152, n71153, n71154, n71155, n71156, n71157, n71158, n71159,
    n71160, n71161, n71162, n71163, n71164, n71165, n71166, n71167, n71168,
    n71169, n71170, n71171, n71172, n71173, n71174, n71175, n71176, n71177,
    n71178, n71179, n71180, n71181, n71182, n71183, n71184, n71185, n71186,
    n71187, n71188, n71189, n71190, n71191, n71192, n71193, n71194, n71195,
    n71196, n71197, n71198, n71199, n71200, n71201, n71202, n71203, n71204,
    n71205, n71206, n71207, n71208, n71209, n71210, n71211, n71212, n71213,
    n71214, n71215, n71216, n71217, n71218, n71219, n71220, n71221, n71222,
    n71223, n71224, n71225, n71226, n71227, n71228, n71229, n71230, n71231,
    n71232, n71233, n71234, n71235, n71236, n71237, n71238, n71239, n71240,
    n71241, n71242, n71243, n71244, n71245, n71246, n71247, n71248, n71249,
    n71250, n71251, n71252, n71253, n71254, n71255, n71256, n71257, n71258,
    n71259, n71260, n71261, n71262, n71263, n71264, n71265, n71266, n71267,
    n71268, n71269, n71270, n71271, n71272, n71273, n71274, n71275, n71276,
    n71277, n71278, n71279, n71280, n71281, n71282, n71283, n71284, n71285,
    n71286, n71287, n71288, n71289, n71290, n71291, n71292, n71293, n71294,
    n71295, n71296, n71297, n71298, n71299, n71300, n71301, n71302, n71303,
    n71304, n71305, n71306, n71307, n71308, n71309, n71310, n71311, n71312,
    n71313, n71314, n71315, n71316, n71317, n71318, n71319, n71320, n71321,
    n71322, n71323, n71324, n71325, n71326, n71327, n71328, n71329, n71330,
    n71331, n71332, n71333, n71334, n71335, n71336, n71337, n71338, n71339,
    n71340, n71341, n71342, n71343, n71344, n71345, n71346, n71347, n71348,
    n71349, n71350, n71351, n71352, n71353, n71354, n71355, n71356, n71357,
    n71358, n71359, n71360, n71361, n71362, n71363, n71364, n71365, n71366,
    n71367, n71368, n71369, n71370;
  assign n109 = fair_cnt<0>_out  & ~fair_cnt<1>_out ;
  assign n110 = ~fair_cnt<1>_out  & ~n109;
  assign n111 = fair_cnt<2>_out  & ~n110;
  assign n112 = ~next_sys_fair<4>_out  & n111;
  assign n113 = ~next_sys_fair<4>_out  & ~n112;
  assign n114 = ~reg_stateG3_0_out & ~n113;
  assign n115 = ~reg_stateG3_0_out & ~n114;
  assign n116 = ~reg_stateG3_1_out & ~n115;
  assign n117 = ~reg_stateG3_1_out & ~n116;
  assign n118 = ~reg_stateG3_2_out & ~n117;
  assign n119 = ~reg_stateG3_2_out & ~n118;
  assign n120 = ~reg_stateG2_out & ~n119;
  assign n121 = ~reg_stateG2_out & ~n120;
  assign n122 = ~reg_stateA1_out & ~n121;
  assign n123 = ~reg_stateA1_out & ~n122;
  assign n124 = reg_controllable_locked_out & ~n123;
  assign n125 = ~reg_controllable_locked_out & ~n121;
  assign n126 = ~n124 & ~n125;
  assign n127 = ~reg_controllable_hgrant2_out & ~n126;
  assign n128 = ~reg_controllable_hgrant2_out & ~n127;
  assign n129 = ~reg_controllable_hgrant1_out & ~n128;
  assign n130 = ~reg_controllable_hgrant1_out & ~n129;
  assign n131 = ~reg_controllable_hgrant3_out & ~n130;
  assign n132 = ~reg_controllable_hgrant3_out & ~n131;
  assign n133 = ~next_sys_fair<2>_out  & ~n132;
  assign n134 = ~next_sys_fair<2>_out  & ~n133;
  assign n135 = ~reg_controllable_hgrant4_out & ~n134;
  assign n136 = ~reg_controllable_hgrant4_out & ~n135;
  assign n137 = ~reg_controllable_hgrant5_out & ~n136;
  assign n138 = ~reg_controllable_hgrant5_out & ~n137;
  assign n139 = ~reg_stateG10_9_out & ~n138;
  assign n140 = ~reg_stateG10_9_out & ~n139;
  assign n141 = next_sys_fair<0>_out  & ~n140;
  assign n142 = ~fair_cnt<2>_out  & ~n110;
  assign n143 = ~fair_cnt<2>_out  & ~n142;
  assign n144 = ~next_sys_fair<4>_out  & ~n143;
  assign n145 = ~next_sys_fair<4>_out  & ~n144;
  assign n146 = ~reg_stateG3_0_out & ~n145;
  assign n147 = ~reg_stateG3_0_out & ~n146;
  assign n148 = ~reg_stateG3_1_out & ~n147;
  assign n149 = ~reg_stateG3_1_out & ~n148;
  assign n150 = ~reg_stateG3_2_out & ~n149;
  assign n151 = ~reg_stateG3_2_out & ~n150;
  assign n152 = ~reg_stateG2_out & ~n151;
  assign n153 = ~reg_stateG2_out & ~n152;
  assign n154 = ~reg_stateA1_out & ~n153;
  assign n155 = ~reg_stateA1_out & ~n154;
  assign n156 = reg_controllable_locked_out & ~n155;
  assign n157 = fair_cnt<0>_out  & fair_cnt<1>_out ;
  assign n158 = ~fair_cnt<2>_out  & n157;
  assign n159 = ~fair_cnt<2>_out  & ~n158;
  assign n160 = ~next_sys_fair<4>_out  & ~n159;
  assign n161 = ~next_sys_fair<4>_out  & ~n160;
  assign n162 = ~reg_stateG3_0_out & ~n161;
  assign n163 = ~reg_stateG3_0_out & ~n162;
  assign n164 = ~reg_stateG3_1_out & ~n163;
  assign n165 = ~reg_stateG3_1_out & ~n164;
  assign n166 = ~reg_stateG3_2_out & ~n165;
  assign n167 = ~reg_stateG3_2_out & ~n166;
  assign n168 = next_env_fair_out & ~n167;
  assign n169 = fair_cnt<2>_out  & ~next_sys_fair<4>_out ;
  assign n170 = ~next_sys_fair<4>_out  & ~n169;
  assign n171 = ~reg_stateG3_0_out & ~n170;
  assign n172 = ~reg_stateG3_0_out & ~n171;
  assign n173 = ~reg_stateG3_1_out & ~n172;
  assign n174 = ~reg_stateG3_1_out & ~n173;
  assign n175 = ~reg_stateG3_2_out & ~n174;
  assign n176 = ~reg_stateG3_2_out & ~n175;
  assign n177 = ~next_env_fair_out & ~n176;
  assign n178 = ~n168 & ~n177;
  assign n179 = ~reg_stateG2_out & ~n178;
  assign n180 = ~reg_stateG2_out & ~n179;
  assign n181 = ~reg_controllable_locked_out & ~n180;
  assign n182 = ~n156 & ~n181;
  assign n183 = ~reg_controllable_hgrant2_out & ~n182;
  assign n184 = ~reg_controllable_hgrant2_out & ~n183;
  assign n185 = ~reg_controllable_hgrant1_out & ~n184;
  assign n186 = ~reg_controllable_hgrant1_out & ~n185;
  assign n187 = ~reg_controllable_hgrant3_out & ~n186;
  assign n188 = ~reg_controllable_hgrant3_out & ~n187;
  assign n189 = ~next_sys_fair<2>_out  & ~n188;
  assign n190 = ~next_sys_fair<2>_out  & ~n189;
  assign n191 = ~reg_controllable_hgrant4_out & ~n190;
  assign n192 = ~reg_controllable_hgrant4_out & ~n191;
  assign n193 = ~reg_controllable_hgrant5_out & ~n192;
  assign n194 = ~reg_controllable_hgrant5_out & ~n193;
  assign n195 = ~reg_stateG10_9_out & ~n194;
  assign n196 = ~reg_stateG10_9_out & ~n195;
  assign n197 = ~next_sys_fair<0>_out  & ~n196;
  assign n198 = ~n141 & ~n197;
  assign n199 = next_sys_fair<3>_out  & ~n198;
  assign n200 = ~reg_controllable_hgrant4_out & ~n188;
  assign n201 = ~reg_controllable_hgrant4_out & ~n200;
  assign n202 = ~reg_controllable_hgrant5_out & ~n201;
  assign n203 = ~reg_controllable_hgrant5_out & ~n202;
  assign n204 = ~reg_stateG10_9_out & ~n203;
  assign n205 = ~reg_stateG10_9_out & ~n204;
  assign n206 = ~next_sys_fair<3>_out  & ~n205;
  assign n207 = ~n199 & ~n206;
  assign n208 = reg_controllable_hmaster1_out & ~n207;
  assign n209 = reg_controllable_hmaster2_out & ~n207;
  assign n210 = reg_stateG3_2_out & ~n117;
  assign n211 = ~reg_stateG3_2_out & ~n113;
  assign n212 = ~n210 & ~n211;
  assign n213 = reg_stateA1_out & ~n212;
  assign n214 = ~reg_stateG2_out & ~n212;
  assign n215 = ~reg_stateG2_out & ~n214;
  assign n216 = ~reg_stateA1_out & ~n215;
  assign n217 = ~n213 & ~n216;
  assign n218 = reg_controllable_hmastlock_out & ~n217;
  assign n219 = ~reg_controllable_hmastlock_out & ~n123;
  assign n220 = ~n218 & ~n219;
  assign n221 = reg_controllable_locked_out & ~n220;
  assign n222 = reg_controllable_hmastlock_out & ~n121;
  assign n223 = ~reg_controllable_hmastlock_out & ~n217;
  assign n224 = ~n222 & ~n223;
  assign n225 = ~reg_controllable_locked_out & ~n224;
  assign n226 = ~n221 & ~n225;
  assign n227 = ~reg_controllable_hgrant2_out & ~n226;
  assign n228 = ~reg_controllable_hgrant2_out & ~n227;
  assign n229 = ~reg_controllable_hgrant1_out & ~n228;
  assign n230 = ~reg_controllable_hgrant1_out & ~n229;
  assign n231 = ~reg_controllable_hgrant3_out & ~n230;
  assign n232 = ~reg_controllable_hgrant3_out & ~n231;
  assign n233 = ~next_sys_fair<2>_out  & ~n232;
  assign n234 = ~next_sys_fair<2>_out  & ~n233;
  assign n235 = ~reg_controllable_hgrant4_out & ~n234;
  assign n236 = ~reg_controllable_hgrant4_out & ~n235;
  assign n237 = ~reg_controllable_hgrant5_out & ~n236;
  assign n238 = ~reg_controllable_hgrant5_out & ~n237;
  assign n239 = ~reg_stateG10_9_out & ~n238;
  assign n240 = ~reg_stateG10_9_out & ~n239;
  assign n241 = next_sys_fair<0>_out  & ~n240;
  assign n242 = reg_stateG3_2_out & ~n165;
  assign n243 = reg_stateG3_0_out & ~n161;
  assign n244 = fair_cnt<1>_out  & ~fair_cnt<2>_out ;
  assign n245 = ~fair_cnt<2>_out  & ~n244;
  assign n246 = ~next_sys_fair<4>_out  & ~n245;
  assign n247 = ~next_sys_fair<4>_out  & ~n246;
  assign n248 = ~reg_stateG3_0_out & ~n247;
  assign n249 = ~n243 & ~n248;
  assign n250 = reg_stateG3_1_out & ~n249;
  assign n251 = reg_stateG3_0_out & ~n145;
  assign n252 = ~n162 & ~n251;
  assign n253 = ~reg_stateG3_1_out & ~n252;
  assign n254 = ~n250 & ~n253;
  assign n255 = ~reg_stateG3_2_out & ~n254;
  assign n256 = ~n242 & ~n255;
  assign n257 = next_env_fair_out & ~n256;
  assign n258 = reg_stateG3_2_out & ~n174;
  assign n259 = ~n171 & ~n251;
  assign n260 = ~reg_stateG3_1_out & ~n259;
  assign n261 = ~n250 & ~n260;
  assign n262 = ~reg_stateG3_2_out & ~n261;
  assign n263 = ~n258 & ~n262;
  assign n264 = ~next_env_fair_out & ~n263;
  assign n265 = ~n257 & ~n264;
  assign n266 = reg_stateA1_out & ~n265;
  assign n267 = ~reg_stateG2_out & ~n265;
  assign n268 = ~reg_stateG2_out & ~n267;
  assign n269 = ~reg_stateA1_out & ~n268;
  assign n270 = ~n266 & ~n269;
  assign n271 = reg_controllable_hmastlock_out & ~n270;
  assign n272 = ~reg_controllable_hmastlock_out & ~n155;
  assign n273 = ~n271 & ~n272;
  assign n274 = reg_controllable_locked_out & ~n273;
  assign n275 = reg_controllable_hmastlock_out & ~n180;
  assign n276 = ~reg_controllable_hmastlock_out & ~n270;
  assign n277 = ~n275 & ~n276;
  assign n278 = ~reg_controllable_locked_out & ~n277;
  assign n279 = ~n274 & ~n278;
  assign n280 = ~reg_controllable_hgrant2_out & ~n279;
  assign n281 = ~reg_controllable_hgrant2_out & ~n280;
  assign n282 = ~reg_controllable_hgrant1_out & ~n281;
  assign n283 = ~reg_controllable_hgrant1_out & ~n282;
  assign n284 = ~reg_controllable_hgrant3_out & ~n283;
  assign n285 = ~reg_controllable_hgrant3_out & ~n284;
  assign n286 = ~next_sys_fair<2>_out  & ~n285;
  assign n287 = ~next_sys_fair<2>_out  & ~n286;
  assign n288 = ~reg_controllable_hgrant4_out & ~n287;
  assign n289 = ~reg_controllable_hgrant4_out & ~n288;
  assign n290 = ~reg_controllable_hgrant5_out & ~n289;
  assign n291 = ~reg_controllable_hgrant5_out & ~n290;
  assign n292 = ~reg_stateG10_9_out & ~n291;
  assign n293 = ~reg_stateG10_9_out & ~n292;
  assign n294 = ~next_sys_fair<0>_out  & ~n293;
  assign n295 = ~n241 & ~n294;
  assign n296 = next_sys_fair<3>_out  & ~n295;
  assign n297 = ~reg_controllable_hgrant4_out & ~n285;
  assign n298 = ~reg_controllable_hgrant4_out & ~n297;
  assign n299 = ~reg_controllable_hgrant5_out & ~n298;
  assign n300 = ~reg_controllable_hgrant5_out & ~n299;
  assign n301 = ~reg_stateG10_9_out & ~n300;
  assign n302 = ~reg_stateG10_9_out & ~n301;
  assign n303 = ~next_sys_fair<3>_out  & ~n302;
  assign n304 = ~n296 & ~n303;
  assign n305 = ~reg_controllable_hmaster2_out & ~n304;
  assign n306 = ~n209 & ~n305;
  assign n307 = ~reg_controllable_hmaster1_out & ~n306;
  assign n308 = ~n208 & ~n307;
  assign n309 = next_sys_fair<1>_out  & ~n308;
  assign n310 = next_sys_fair<3>_out  & ~n196;
  assign n311 = next_sys_fair<2>_out  & ~n188;
  assign n312 = ~n133 & ~n311;
  assign n313 = ~reg_controllable_hgrant4_out & ~n312;
  assign n314 = ~reg_controllable_hgrant4_out & ~n313;
  assign n315 = ~reg_controllable_hgrant5_out & ~n314;
  assign n316 = ~reg_controllable_hgrant5_out & ~n315;
  assign n317 = ~reg_stateG10_9_out & ~n316;
  assign n318 = ~reg_stateG10_9_out & ~n317;
  assign n319 = ~next_sys_fair<3>_out  & ~n318;
  assign n320 = ~n310 & ~n319;
  assign n321 = reg_controllable_hmaster1_out & ~n320;
  assign n322 = reg_controllable_hmaster2_out & ~n320;
  assign n323 = next_sys_fair<3>_out  & ~n293;
  assign n324 = next_sys_fair<2>_out  & ~n285;
  assign n325 = ~n114 & ~n251;
  assign n326 = ~reg_stateG3_1_out & ~n325;
  assign n327 = ~n250 & ~n326;
  assign n328 = ~reg_stateG3_2_out & ~n327;
  assign n329 = ~n258 & ~n328;
  assign n330 = reg_stateA1_out & ~n329;
  assign n331 = ~reg_stateG2_out & ~n329;
  assign n332 = ~reg_stateG2_out & ~n331;
  assign n333 = ~reg_stateA1_out & ~n332;
  assign n334 = ~n330 & ~n333;
  assign n335 = reg_controllable_hmastlock_out & ~n334;
  assign n336 = ~n219 & ~n335;
  assign n337 = reg_controllable_locked_out & ~n336;
  assign n338 = ~reg_controllable_hmastlock_out & ~n334;
  assign n339 = ~n222 & ~n338;
  assign n340 = ~reg_controllable_locked_out & ~n339;
  assign n341 = ~n337 & ~n340;
  assign n342 = ~reg_controllable_hgrant2_out & ~n341;
  assign n343 = ~reg_controllable_hgrant2_out & ~n342;
  assign n344 = ~reg_controllable_hgrant1_out & ~n343;
  assign n345 = ~reg_controllable_hgrant1_out & ~n344;
  assign n346 = ~reg_controllable_hgrant3_out & ~n345;
  assign n347 = ~reg_controllable_hgrant3_out & ~n346;
  assign n348 = ~next_sys_fair<2>_out  & ~n347;
  assign n349 = ~n324 & ~n348;
  assign n350 = ~reg_controllable_hgrant4_out & ~n349;
  assign n351 = ~reg_controllable_hgrant4_out & ~n350;
  assign n352 = ~reg_controllable_hgrant5_out & ~n351;
  assign n353 = ~reg_controllable_hgrant5_out & ~n352;
  assign n354 = ~reg_stateG10_9_out & ~n353;
  assign n355 = ~reg_stateG10_9_out & ~n354;
  assign n356 = next_sys_fair<0>_out  & ~n355;
  assign n357 = ~reg_stateG3_2_out & ~n170;
  assign n358 = ~n258 & ~n357;
  assign n359 = next_env_fair_out & ~n358;
  assign n360 = ~next_env_fair_out & ~n212;
  assign n361 = ~n359 & ~n360;
  assign n362 = reg_stateG2_out & ~n361;
  assign n363 = ~n214 & ~n362;
  assign n364 = reg_stateA1_out & ~n363;
  assign n365 = ~n216 & ~n364;
  assign n366 = reg_controllable_hmastlock_out & ~n365;
  assign n367 = ~n219 & ~n366;
  assign n368 = reg_controllable_locked_out & ~n367;
  assign n369 = ~reg_controllable_hmastlock_out & ~n365;
  assign n370 = ~n222 & ~n369;
  assign n371 = ~reg_controllable_locked_out & ~n370;
  assign n372 = ~n368 & ~n371;
  assign n373 = ~reg_controllable_hgrant2_out & ~n372;
  assign n374 = ~reg_controllable_hgrant2_out & ~n373;
  assign n375 = ~reg_controllable_hgrant1_out & ~n374;
  assign n376 = ~reg_controllable_hgrant1_out & ~n375;
  assign n377 = ~reg_controllable_hgrant3_out & ~n376;
  assign n378 = ~reg_controllable_hgrant3_out & ~n377;
  assign n379 = ~next_sys_fair<2>_out  & ~n378;
  assign n380 = ~n324 & ~n379;
  assign n381 = ~reg_controllable_hgrant4_out & ~n380;
  assign n382 = ~reg_controllable_hgrant4_out & ~n381;
  assign n383 = ~reg_controllable_hgrant5_out & ~n382;
  assign n384 = ~reg_controllable_hgrant5_out & ~n383;
  assign n385 = ~reg_stateG10_9_out & ~n384;
  assign n386 = ~reg_stateG10_9_out & ~n385;
  assign n387 = ~next_sys_fair<0>_out  & ~n386;
  assign n388 = ~n356 & ~n387;
  assign n389 = ~next_sys_fair<3>_out  & ~n388;
  assign n390 = ~n323 & ~n389;
  assign n391 = ~reg_controllable_hmaster2_out & ~n390;
  assign n392 = ~n322 & ~n391;
  assign n393 = ~reg_controllable_hmaster1_out & ~n392;
  assign n394 = ~n321 & ~n393;
  assign n395 = ~next_sys_fair<1>_out  & ~n394;
  assign n396 = ~n309 & ~n395;
  assign n397 = reg_controllable_hmaster0_out & ~n396;
  assign n398 = next_sys_fair<1>_out  & ~n207;
  assign n399 = ~next_sys_fair<1>_out  & ~n320;
  assign n400 = ~n398 & ~n399;
  assign n401 = ~reg_controllable_hmaster0_out & ~n400;
  assign n402 = ~n397 & ~n401;
  assign n403 = reg_controllable_hmaster3_out & ~n402;
  assign n404 = ~reg_controllable_hmaster3_out & ~n400;
  assign n405 = ~n403 & ~n404;
  assign n406 = ~reg_controllable_hgrant6_out & ~n405;
  assign n407 = ~reg_controllable_hgrant6_out & ~n406;
  assign n408 = ~reg_controllable_hgrant8_out & ~n407;
  assign n409 = ~reg_controllable_hgrant8_out & ~n408;
  assign n410 = ~reg_controllable_hgrant7_out & ~n409;
  assign n411 = ~reg_controllable_hgrant7_out & ~n410;
  assign n412 = reg_controllable_hgrant9_out & ~n411;
  assign n413 = next_sys_fair<3>_out  & ~n194;
  assign n414 = ~next_sys_fair<3>_out  & ~n203;
  assign n415 = ~n413 & ~n414;
  assign n416 = next_sys_fair<1>_out  & ~n415;
  assign n417 = next_sys_fair<0>_out  & ~n138;
  assign n418 = ~next_sys_fair<0>_out  & ~n194;
  assign n419 = ~n417 & ~n418;
  assign n420 = next_sys_fair<3>_out  & ~n419;
  assign n421 = ~next_sys_fair<3>_out  & ~n316;
  assign n422 = ~n420 & ~n421;
  assign n423 = ~next_sys_fair<1>_out  & ~n422;
  assign n424 = ~n416 & ~n423;
  assign n425 = reg_controllable_hmaster3_out & ~n424;
  assign n426 = next_sys_fair<3>_out  & ~n291;
  assign n427 = ~next_sys_fair<3>_out  & ~n300;
  assign n428 = ~n426 & ~n427;
  assign n429 = reg_controllable_hmaster2_out & ~n428;
  assign n430 = ~reg_controllable_hmaster2_out & ~n415;
  assign n431 = ~n429 & ~n430;
  assign n432 = reg_controllable_hmaster1_out & ~n431;
  assign n433 = ~reg_controllable_hmaster1_out & ~n415;
  assign n434 = ~n432 & ~n433;
  assign n435 = next_sys_fair<1>_out  & ~n434;
  assign n436 = next_sys_fair<0>_out  & ~n238;
  assign n437 = ~next_sys_fair<0>_out  & ~n291;
  assign n438 = ~n436 & ~n437;
  assign n439 = next_sys_fair<3>_out  & ~n438;
  assign n440 = next_sys_fair<0>_out  & ~n353;
  assign n441 = ~next_sys_fair<0>_out  & ~n384;
  assign n442 = ~n440 & ~n441;
  assign n443 = ~next_sys_fair<3>_out  & ~n442;
  assign n444 = ~n439 & ~n443;
  assign n445 = reg_controllable_hmaster2_out & ~n444;
  assign n446 = ~reg_controllable_hmaster2_out & ~n422;
  assign n447 = ~n445 & ~n446;
  assign n448 = reg_controllable_hmaster1_out & ~n447;
  assign n449 = ~reg_controllable_hmaster1_out & ~n422;
  assign n450 = ~n448 & ~n449;
  assign n451 = ~next_sys_fair<1>_out  & ~n450;
  assign n452 = ~n435 & ~n451;
  assign n453 = reg_controllable_hmaster0_out & ~n452;
  assign n454 = ~reg_controllable_hmaster0_out & ~n424;
  assign n455 = ~n453 & ~n454;
  assign n456 = ~reg_controllable_hmaster3_out & ~n455;
  assign n457 = ~n425 & ~n456;
  assign n458 = ~reg_controllable_hgrant6_out & ~n457;
  assign n459 = ~reg_controllable_hgrant6_out & ~n458;
  assign n460 = ~reg_stateG10_7_out & ~n459;
  assign n461 = ~reg_stateG10_7_out & ~n460;
  assign n462 = ~reg_controllable_hgrant8_out & ~n461;
  assign n463 = ~reg_controllable_hgrant8_out & ~n462;
  assign n464 = reg_controllable_hgrant7_out & ~n463;
  assign n465 = next_sys_fair<0>_out  & ~n194;
  assign n466 = ~next_sys_fair<0>_out  & ~n138;
  assign n467 = ~n465 & ~n466;
  assign n468 = next_sys_fair<3>_out  & ~n467;
  assign n469 = ~n414 & ~n468;
  assign n470 = next_sys_fair<1>_out  & ~n469;
  assign n471 = ~n413 & ~n421;
  assign n472 = ~next_sys_fair<1>_out  & ~n471;
  assign n473 = ~n470 & ~n472;
  assign n474 = reg_controllable_hmaster0_out & ~n473;
  assign n475 = reg_controllable_hmaster1_out & ~n469;
  assign n476 = reg_controllable_hmaster2_out & ~n469;
  assign n477 = next_sys_fair<0>_out  & ~n291;
  assign n478 = ~next_sys_fair<0>_out  & ~n238;
  assign n479 = ~n477 & ~n478;
  assign n480 = next_sys_fair<3>_out  & ~n479;
  assign n481 = ~n427 & ~n480;
  assign n482 = ~reg_controllable_hmaster2_out & ~n481;
  assign n483 = ~n476 & ~n482;
  assign n484 = ~reg_controllable_hmaster1_out & ~n483;
  assign n485 = ~n475 & ~n484;
  assign n486 = next_sys_fair<1>_out  & ~n485;
  assign n487 = reg_controllable_hmaster1_out & ~n471;
  assign n488 = reg_controllable_hmaster2_out & ~n471;
  assign n489 = ~n426 & ~n443;
  assign n490 = ~reg_controllable_hmaster2_out & ~n489;
  assign n491 = ~n488 & ~n490;
  assign n492 = ~reg_controllable_hmaster1_out & ~n491;
  assign n493 = ~n487 & ~n492;
  assign n494 = ~next_sys_fair<1>_out  & ~n493;
  assign n495 = ~n486 & ~n494;
  assign n496 = ~reg_controllable_hmaster0_out & ~n495;
  assign n497 = ~n474 & ~n496;
  assign n498 = reg_controllable_hmaster3_out & ~n497;
  assign n499 = ~reg_controllable_hmaster3_out & ~n473;
  assign n500 = ~n498 & ~n499;
  assign n501 = ~reg_stateG10_8_out & ~n500;
  assign n502 = ~reg_stateG10_8_out & ~n501;
  assign n503 = ~reg_controllable_hgrant6_out & ~n502;
  assign n504 = ~reg_controllable_hgrant6_out & ~n503;
  assign n505 = reg_controllable_hgrant8_out & ~n504;
  assign n506 = ~reg_stateG10_6_out & ~n415;
  assign n507 = ~reg_stateG10_6_out & ~n506;
  assign n508 = next_sys_fair<1>_out  & ~n507;
  assign n509 = ~n421 & ~n468;
  assign n510 = ~reg_stateG10_6_out & ~n509;
  assign n511 = ~reg_stateG10_6_out & ~n510;
  assign n512 = ~next_sys_fair<1>_out  & ~n511;
  assign n513 = ~n508 & ~n512;
  assign n514 = reg_controllable_hmaster3_out & ~n513;
  assign n515 = reg_controllable_hmaster0_out & ~n513;
  assign n516 = ~reg_stateG10_6_out & ~n434;
  assign n517 = ~reg_stateG10_6_out & ~n516;
  assign n518 = next_sys_fair<1>_out  & ~n517;
  assign n519 = ~n443 & ~n480;
  assign n520 = reg_controllable_hmaster2_out & ~n519;
  assign n521 = ~reg_controllable_hmaster2_out & ~n509;
  assign n522 = ~n520 & ~n521;
  assign n523 = reg_controllable_hmaster1_out & ~n522;
  assign n524 = ~reg_controllable_hmaster1_out & ~n509;
  assign n525 = ~n523 & ~n524;
  assign n526 = ~reg_stateG10_6_out & ~n525;
  assign n527 = ~reg_stateG10_6_out & ~n526;
  assign n528 = ~next_sys_fair<1>_out  & ~n527;
  assign n529 = ~n518 & ~n528;
  assign n530 = ~reg_controllable_hmaster0_out & ~n529;
  assign n531 = ~n515 & ~n530;
  assign n532 = ~reg_controllable_hmaster3_out & ~n531;
  assign n533 = ~n514 & ~n532;
  assign n534 = reg_controllable_hgrant6_out & ~n533;
  assign n535 = ~reg_stateG10_5_out & ~n192;
  assign n536 = ~reg_stateG10_5_out & ~n535;
  assign n537 = reg_controllable_hgrant5_out & ~n536;
  assign n538 = ~reg_stateG10_4_out & ~n190;
  assign n539 = ~reg_stateG10_4_out & ~n538;
  assign n540 = reg_controllable_hgrant4_out & ~n539;
  assign n541 = fair_cnt<2>_out  & next_env_fair_out;
  assign n542 = ~next_env_fair_out & n111;
  assign n543 = ~n541 & ~n542;
  assign n544 = reg_stateA1_out & ~n543;
  assign n545 = reg_stateA1_out & ~n544;
  assign n546 = reg_controllable_hmastlock_out & ~n545;
  assign n547 = ~reg_stateG3_0_out & fair_cnt<2>_out ;
  assign n548 = ~reg_stateG3_0_out & ~n547;
  assign n549 = ~reg_stateG3_1_out & ~n548;
  assign n550 = ~reg_stateG3_1_out & ~n549;
  assign n551 = ~reg_stateG3_2_out & ~n550;
  assign n552 = ~reg_stateG3_2_out & ~n551;
  assign n553 = next_env_fair_out & ~n552;
  assign n554 = ~reg_stateG3_0_out & n111;
  assign n555 = ~reg_stateG3_0_out & ~n554;
  assign n556 = ~reg_stateG3_1_out & ~n555;
  assign n557 = ~reg_stateG3_1_out & ~n556;
  assign n558 = ~reg_stateG3_2_out & ~n557;
  assign n559 = ~reg_stateG3_2_out & ~n558;
  assign n560 = ~next_env_fair_out & ~n559;
  assign n561 = ~n553 & ~n560;
  assign n562 = ~reg_stateG2_out & ~n561;
  assign n563 = ~reg_stateG2_out & ~n562;
  assign n564 = reg_stateA1_out & ~n563;
  assign n565 = reg_stateA1_out & ~n564;
  assign n566 = ~reg_controllable_hmastlock_out & ~n565;
  assign n567 = ~n546 & ~n566;
  assign n568 = reg_controllable_locked_out & ~n567;
  assign n569 = reg_controllable_hmastlock_out & ~n565;
  assign n570 = ~reg_controllable_hmastlock_out & ~n545;
  assign n571 = ~n569 & ~n570;
  assign n572 = ~reg_controllable_locked_out & ~n571;
  assign n573 = ~n568 & ~n572;
  assign n574 = ~reg_controllable_hgrant2_out & ~n573;
  assign n575 = ~reg_controllable_hgrant2_out & ~n574;
  assign n576 = ~reg_controllable_hgrant1_out & ~n575;
  assign n577 = ~reg_controllable_hgrant1_out & ~n576;
  assign n578 = ~reg_controllable_hgrant3_out & ~n577;
  assign n579 = ~reg_controllable_hgrant3_out & ~n578;
  assign n580 = next_sys_fair<2>_out  & ~n579;
  assign n581 = ~reg_stateG10_3_out & ~n186;
  assign n582 = ~reg_stateG10_3_out & ~n581;
  assign n583 = reg_controllable_hgrant3_out & ~n582;
  assign n584 = ~reg_stateG10_1_out & ~n184;
  assign n585 = ~reg_stateG10_1_out & ~n584;
  assign n586 = reg_controllable_hgrant1_out & ~n585;
  assign n587 = ~reg_stateG10_2_out & ~n182;
  assign n588 = ~reg_stateG10_2_out & ~n587;
  assign n589 = reg_controllable_hgrant2_out & ~n588;
  assign n590 = ~reg_stateA1_out & ~n265;
  assign n591 = ~n544 & ~n590;
  assign n592 = reg_controllable_hmastlock_out & ~n591;
  assign n593 = ~n154 & ~n564;
  assign n594 = ~reg_controllable_hmastlock_out & ~n593;
  assign n595 = ~n592 & ~n594;
  assign n596 = reg_controllable_locked_out & ~n595;
  assign n597 = ~reg_stateA1_out & ~n180;
  assign n598 = ~n564 & ~n597;
  assign n599 = reg_controllable_hmastlock_out & ~n598;
  assign n600 = ~reg_controllable_hmastlock_out & ~n591;
  assign n601 = ~n599 & ~n600;
  assign n602 = ~reg_controllable_locked_out & ~n601;
  assign n603 = ~n596 & ~n602;
  assign n604 = ~reg_controllable_hgrant2_out & ~n603;
  assign n605 = ~n589 & ~n604;
  assign n606 = ~reg_controllable_hgrant1_out & ~n605;
  assign n607 = ~n586 & ~n606;
  assign n608 = ~reg_controllable_hgrant3_out & ~n607;
  assign n609 = ~n583 & ~n608;
  assign n610 = ~next_sys_fair<2>_out  & ~n609;
  assign n611 = ~n580 & ~n610;
  assign n612 = ~reg_controllable_hgrant4_out & ~n611;
  assign n613 = ~n540 & ~n612;
  assign n614 = ~reg_controllable_hgrant5_out & ~n613;
  assign n615 = ~n537 & ~n614;
  assign n616 = next_sys_fair<3>_out  & ~n615;
  assign n617 = next_sys_fair<2>_out  & ~n132;
  assign n618 = ~n189 & ~n617;
  assign n619 = ~reg_controllable_hgrant4_out & ~n618;
  assign n620 = ~reg_controllable_hgrant4_out & ~n619;
  assign n621 = ~reg_stateG10_5_out & ~n620;
  assign n622 = ~reg_stateG10_5_out & ~n621;
  assign n623 = reg_controllable_hgrant5_out & ~n622;
  assign n624 = ~reg_stateG10_4_out & ~n188;
  assign n625 = ~reg_stateG10_4_out & ~n624;
  assign n626 = reg_controllable_hgrant4_out & ~n625;
  assign n627 = next_sys_fair<2>_out  & ~n609;
  assign n628 = ~reg_stateG10_1_out & ~n128;
  assign n629 = ~reg_stateG10_1_out & ~n628;
  assign n630 = reg_controllable_hgrant1_out & ~n629;
  assign n631 = ~n606 & ~n630;
  assign n632 = ~reg_controllable_hgrant3_out & ~n631;
  assign n633 = ~n583 & ~n632;
  assign n634 = ~next_sys_fair<2>_out  & ~n633;
  assign n635 = ~n627 & ~n634;
  assign n636 = ~reg_controllable_hgrant4_out & ~n635;
  assign n637 = ~n626 & ~n636;
  assign n638 = ~reg_controllable_hgrant5_out & ~n637;
  assign n639 = ~n623 & ~n638;
  assign n640 = next_sys_fair<0>_out  & ~n639;
  assign n641 = ~reg_stateG10_5_out & ~n201;
  assign n642 = ~reg_stateG10_5_out & ~n641;
  assign n643 = reg_controllable_hgrant5_out & ~n642;
  assign n644 = ~reg_stateG10_4_out & ~n618;
  assign n645 = ~reg_stateG10_4_out & ~n644;
  assign n646 = reg_controllable_hgrant4_out & ~n645;
  assign n647 = ~reg_controllable_hgrant4_out & ~n609;
  assign n648 = ~n646 & ~n647;
  assign n649 = ~reg_controllable_hgrant5_out & ~n648;
  assign n650 = ~n643 & ~n649;
  assign n651 = ~next_sys_fair<0>_out  & ~n650;
  assign n652 = ~n640 & ~n651;
  assign n653 = ~next_sys_fair<3>_out  & ~n652;
  assign n654 = ~n616 & ~n653;
  assign n655 = reg_controllable_hmaster1_out & ~n654;
  assign n656 = reg_controllable_hmaster2_out & ~n654;
  assign n657 = ~reg_controllable_hgrant2_out & ~n565;
  assign n658 = ~reg_controllable_hgrant2_out & ~n657;
  assign n659 = ~reg_controllable_hgrant1_out & ~n658;
  assign n660 = ~reg_controllable_hgrant1_out & ~n659;
  assign n661 = ~reg_controllable_hgrant3_out & ~n660;
  assign n662 = ~reg_controllable_hgrant3_out & ~n661;
  assign n663 = next_sys_fair<2>_out  & ~n662;
  assign n664 = reg_controllable_locked_out & ~n593;
  assign n665 = ~reg_controllable_locked_out & ~n598;
  assign n666 = ~n664 & ~n665;
  assign n667 = ~reg_controllable_hgrant2_out & ~n666;
  assign n668 = ~n589 & ~n667;
  assign n669 = ~reg_controllable_hgrant1_out & ~n668;
  assign n670 = ~n586 & ~n669;
  assign n671 = ~reg_controllable_hgrant3_out & ~n670;
  assign n672 = ~n583 & ~n671;
  assign n673 = ~next_sys_fair<2>_out  & ~n672;
  assign n674 = ~n663 & ~n673;
  assign n675 = ~reg_controllable_hgrant4_out & ~n674;
  assign n676 = ~n540 & ~n675;
  assign n677 = ~reg_controllable_hgrant5_out & ~n676;
  assign n678 = ~n537 & ~n677;
  assign n679 = next_sys_fair<3>_out  & ~n678;
  assign n680 = next_sys_fair<2>_out  & ~n672;
  assign n681 = ~n630 & ~n669;
  assign n682 = ~reg_controllable_hgrant3_out & ~n681;
  assign n683 = ~n583 & ~n682;
  assign n684 = ~next_sys_fair<2>_out  & ~n683;
  assign n685 = ~n680 & ~n684;
  assign n686 = ~reg_controllable_hgrant4_out & ~n685;
  assign n687 = ~n626 & ~n686;
  assign n688 = ~reg_controllable_hgrant5_out & ~n687;
  assign n689 = ~n623 & ~n688;
  assign n690 = next_sys_fair<0>_out  & ~n689;
  assign n691 = ~reg_controllable_hgrant4_out & ~n672;
  assign n692 = ~n646 & ~n691;
  assign n693 = ~reg_controllable_hgrant5_out & ~n692;
  assign n694 = ~n643 & ~n693;
  assign n695 = ~next_sys_fair<0>_out  & ~n694;
  assign n696 = ~n690 & ~n695;
  assign n697 = ~next_sys_fair<3>_out  & ~n696;
  assign n698 = ~n679 & ~n697;
  assign n699 = ~reg_controllable_hmaster2_out & ~n698;
  assign n700 = ~n656 & ~n699;
  assign n701 = ~reg_controllable_hmaster1_out & ~n700;
  assign n702 = ~n655 & ~n701;
  assign n703 = next_sys_fair<1>_out  & ~n702;
  assign n704 = ~reg_stateG10_5_out & ~n314;
  assign n705 = ~reg_stateG10_5_out & ~n704;
  assign n706 = reg_controllable_hgrant5_out & ~n705;
  assign n707 = ~reg_stateG10_4_out & ~n312;
  assign n708 = ~reg_stateG10_4_out & ~n707;
  assign n709 = reg_controllable_hgrant4_out & ~n708;
  assign n710 = ~reg_stateG10_3_out & ~n130;
  assign n711 = ~reg_stateG10_3_out & ~n710;
  assign n712 = reg_controllable_hgrant3_out & ~n711;
  assign n713 = ~n608 & ~n712;
  assign n714 = next_sys_fair<2>_out  & ~n713;
  assign n715 = ~reg_stateG10_2_out & ~n126;
  assign n716 = ~reg_stateG10_2_out & ~n715;
  assign n717 = reg_controllable_hgrant2_out & ~n716;
  assign n718 = reg_stateG3_2_out & fair_cnt<2>_out ;
  assign n719 = reg_stateG3_1_out & fair_cnt<2>_out ;
  assign n720 = reg_stateG3_0_out & fair_cnt<2>_out ;
  assign n721 = fair_cnt<2>_out  & next_sys_fair<4>_out ;
  assign n722 = ~n112 & ~n721;
  assign n723 = ~reg_stateG3_0_out & ~n722;
  assign n724 = ~n720 & ~n723;
  assign n725 = ~reg_stateG3_1_out & ~n724;
  assign n726 = ~n719 & ~n725;
  assign n727 = ~reg_stateG3_2_out & ~n726;
  assign n728 = ~n718 & ~n727;
  assign n729 = next_env_fair_out & ~n728;
  assign n730 = ~n542 & ~n729;
  assign n731 = reg_stateA1_out & ~n730;
  assign n732 = ~reg_stateA1_out & ~n329;
  assign n733 = ~n731 & ~n732;
  assign n734 = reg_controllable_hmastlock_out & ~n733;
  assign n735 = ~reg_stateG3_0_out & ~n723;
  assign n736 = ~reg_stateG3_1_out & ~n735;
  assign n737 = ~reg_stateG3_1_out & ~n736;
  assign n738 = ~reg_stateG3_2_out & ~n737;
  assign n739 = ~reg_stateG3_2_out & ~n738;
  assign n740 = next_env_fair_out & ~n739;
  assign n741 = ~n560 & ~n740;
  assign n742 = ~reg_stateG2_out & ~n741;
  assign n743 = ~reg_stateG2_out & ~n742;
  assign n744 = reg_stateA1_out & ~n743;
  assign n745 = ~n122 & ~n744;
  assign n746 = ~reg_controllable_hmastlock_out & ~n745;
  assign n747 = ~n734 & ~n746;
  assign n748 = reg_controllable_locked_out & ~n747;
  assign n749 = reg_controllable_hmastlock_out & ~n745;
  assign n750 = ~reg_controllable_hmastlock_out & ~n733;
  assign n751 = ~n749 & ~n750;
  assign n752 = ~reg_controllable_locked_out & ~n751;
  assign n753 = ~n748 & ~n752;
  assign n754 = ~reg_controllable_hgrant2_out & ~n753;
  assign n755 = ~n717 & ~n754;
  assign n756 = ~reg_controllable_hgrant1_out & ~n755;
  assign n757 = ~n630 & ~n756;
  assign n758 = ~reg_controllable_hgrant3_out & ~n757;
  assign n759 = ~n712 & ~n758;
  assign n760 = ~next_sys_fair<2>_out  & ~n759;
  assign n761 = ~n714 & ~n760;
  assign n762 = ~reg_controllable_hgrant4_out & ~n761;
  assign n763 = ~n709 & ~n762;
  assign n764 = ~reg_controllable_hgrant5_out & ~n763;
  assign n765 = ~n706 & ~n764;
  assign n766 = next_sys_fair<0>_out  & ~n765;
  assign n767 = ~n604 & ~n717;
  assign n768 = ~reg_controllable_hgrant1_out & ~n767;
  assign n769 = ~n586 & ~n768;
  assign n770 = ~reg_controllable_hgrant3_out & ~n769;
  assign n771 = ~n583 & ~n770;
  assign n772 = next_sys_fair<2>_out  & ~n771;
  assign n773 = reg_stateG2_out & ~n543;
  assign n774 = next_env_fair_out & ~n722;
  assign n775 = ~n542 & ~n774;
  assign n776 = ~reg_stateG2_out & ~n775;
  assign n777 = ~n773 & ~n776;
  assign n778 = reg_stateA1_out & ~n777;
  assign n779 = ~reg_stateA1_out & ~n363;
  assign n780 = ~n778 & ~n779;
  assign n781 = reg_controllable_hmastlock_out & ~n780;
  assign n782 = ~n746 & ~n781;
  assign n783 = reg_controllable_locked_out & ~n782;
  assign n784 = ~reg_controllable_hmastlock_out & ~n780;
  assign n785 = ~n749 & ~n784;
  assign n786 = ~reg_controllable_locked_out & ~n785;
  assign n787 = ~n783 & ~n786;
  assign n788 = ~reg_controllable_hgrant2_out & ~n787;
  assign n789 = ~n717 & ~n788;
  assign n790 = ~reg_controllable_hgrant1_out & ~n789;
  assign n791 = ~n630 & ~n790;
  assign n792 = ~reg_controllable_hgrant3_out & ~n791;
  assign n793 = ~n712 & ~n792;
  assign n794 = ~next_sys_fair<2>_out  & ~n793;
  assign n795 = ~n772 & ~n794;
  assign n796 = ~reg_controllable_hgrant4_out & ~n795;
  assign n797 = ~n709 & ~n796;
  assign n798 = ~reg_controllable_hgrant5_out & ~n797;
  assign n799 = ~n706 & ~n798;
  assign n800 = ~next_sys_fair<0>_out  & ~n799;
  assign n801 = ~n766 & ~n800;
  assign n802 = ~next_sys_fair<3>_out  & ~n801;
  assign n803 = ~n616 & ~n802;
  assign n804 = reg_controllable_hmaster1_out & ~n803;
  assign n805 = reg_controllable_hmaster2_out & ~n803;
  assign n806 = ~n671 & ~n712;
  assign n807 = next_sys_fair<2>_out  & ~n806;
  assign n808 = ~reg_controllable_hgrant2_out & ~n745;
  assign n809 = ~n717 & ~n808;
  assign n810 = ~reg_controllable_hgrant1_out & ~n809;
  assign n811 = ~n630 & ~n810;
  assign n812 = ~reg_controllable_hgrant3_out & ~n811;
  assign n813 = ~n712 & ~n812;
  assign n814 = ~next_sys_fair<2>_out  & ~n813;
  assign n815 = ~n807 & ~n814;
  assign n816 = ~reg_controllable_hgrant4_out & ~n815;
  assign n817 = ~n709 & ~n816;
  assign n818 = ~reg_controllable_hgrant5_out & ~n817;
  assign n819 = ~n706 & ~n818;
  assign n820 = next_sys_fair<0>_out  & ~n819;
  assign n821 = ~n667 & ~n717;
  assign n822 = ~reg_controllable_hgrant1_out & ~n821;
  assign n823 = ~n586 & ~n822;
  assign n824 = ~reg_controllable_hgrant3_out & ~n823;
  assign n825 = ~n583 & ~n824;
  assign n826 = next_sys_fair<2>_out  & ~n825;
  assign n827 = ~n814 & ~n826;
  assign n828 = ~reg_controllable_hgrant4_out & ~n827;
  assign n829 = ~n709 & ~n828;
  assign n830 = ~reg_controllable_hgrant5_out & ~n829;
  assign n831 = ~n706 & ~n830;
  assign n832 = ~next_sys_fair<0>_out  & ~n831;
  assign n833 = ~n820 & ~n832;
  assign n834 = ~next_sys_fair<3>_out  & ~n833;
  assign n835 = ~n679 & ~n834;
  assign n836 = ~reg_controllable_hmaster2_out & ~n835;
  assign n837 = ~n805 & ~n836;
  assign n838 = ~reg_controllable_hmaster1_out & ~n837;
  assign n839 = ~n804 & ~n838;
  assign n840 = ~next_sys_fair<1>_out  & ~n839;
  assign n841 = ~n703 & ~n840;
  assign n842 = reg_controllable_hmaster3_out & ~n841;
  assign n843 = reg_controllable_hmaster2_out & ~n698;
  assign n844 = ~reg_stateG10_3_out & ~n283;
  assign n845 = ~reg_stateG10_3_out & ~n844;
  assign n846 = reg_controllable_hgrant3_out & ~n845;
  assign n847 = ~n671 & ~n846;
  assign n848 = ~next_sys_fair<2>_out  & ~n847;
  assign n849 = ~n663 & ~n848;
  assign n850 = ~reg_controllable_hgrant4_out & ~n849;
  assign n851 = ~n540 & ~n850;
  assign n852 = ~reg_controllable_hgrant5_out & ~n851;
  assign n853 = ~n537 & ~n852;
  assign n854 = next_sys_fair<3>_out  & ~n853;
  assign n855 = next_sys_fair<2>_out  & ~n847;
  assign n856 = ~n682 & ~n846;
  assign n857 = ~next_sys_fair<2>_out  & ~n856;
  assign n858 = ~n855 & ~n857;
  assign n859 = ~reg_controllable_hgrant4_out & ~n858;
  assign n860 = ~n626 & ~n859;
  assign n861 = ~reg_controllable_hgrant5_out & ~n860;
  assign n862 = ~n623 & ~n861;
  assign n863 = next_sys_fair<0>_out  & ~n862;
  assign n864 = ~reg_controllable_hgrant4_out & ~n847;
  assign n865 = ~n646 & ~n864;
  assign n866 = ~reg_controllable_hgrant5_out & ~n865;
  assign n867 = ~n643 & ~n866;
  assign n868 = ~next_sys_fair<0>_out  & ~n867;
  assign n869 = ~n863 & ~n868;
  assign n870 = ~next_sys_fair<3>_out  & ~n869;
  assign n871 = ~n854 & ~n870;
  assign n872 = ~reg_controllable_hmaster2_out & ~n871;
  assign n873 = ~n843 & ~n872;
  assign n874 = reg_controllable_hmaster1_out & ~n873;
  assign n875 = ~reg_stateG10_5_out & ~n289;
  assign n876 = ~reg_stateG10_5_out & ~n875;
  assign n877 = reg_controllable_hgrant5_out & ~n876;
  assign n878 = ~n677 & ~n877;
  assign n879 = next_sys_fair<3>_out  & ~n878;
  assign n880 = next_sys_fair<2>_out  & ~n232;
  assign n881 = ~n286 & ~n880;
  assign n882 = ~reg_controllable_hgrant4_out & ~n881;
  assign n883 = ~reg_controllable_hgrant4_out & ~n882;
  assign n884 = ~reg_stateG10_5_out & ~n883;
  assign n885 = ~reg_stateG10_5_out & ~n884;
  assign n886 = reg_controllable_hgrant5_out & ~n885;
  assign n887 = ~n688 & ~n886;
  assign n888 = next_sys_fair<0>_out  & ~n887;
  assign n889 = ~reg_stateG10_5_out & ~n298;
  assign n890 = ~reg_stateG10_5_out & ~n889;
  assign n891 = reg_controllable_hgrant5_out & ~n890;
  assign n892 = ~n693 & ~n891;
  assign n893 = ~next_sys_fair<0>_out  & ~n892;
  assign n894 = ~n888 & ~n893;
  assign n895 = ~next_sys_fair<3>_out  & ~n894;
  assign n896 = ~n879 & ~n895;
  assign n897 = reg_controllable_hmaster2_out & ~n896;
  assign n898 = ~reg_stateG10_1_out & ~n281;
  assign n899 = ~reg_stateG10_1_out & ~n898;
  assign n900 = reg_controllable_hgrant1_out & ~n899;
  assign n901 = ~n669 & ~n900;
  assign n902 = ~reg_controllable_hgrant3_out & ~n901;
  assign n903 = ~n583 & ~n902;
  assign n904 = ~next_sys_fair<2>_out  & ~n903;
  assign n905 = ~n663 & ~n904;
  assign n906 = ~reg_controllable_hgrant4_out & ~n905;
  assign n907 = ~n540 & ~n906;
  assign n908 = ~reg_controllable_hgrant5_out & ~n907;
  assign n909 = ~n537 & ~n908;
  assign n910 = next_sys_fair<3>_out  & ~n909;
  assign n911 = next_sys_fair<2>_out  & ~n903;
  assign n912 = ~reg_stateG10_1_out & ~n228;
  assign n913 = ~reg_stateG10_1_out & ~n912;
  assign n914 = reg_controllable_hgrant1_out & ~n913;
  assign n915 = ~n669 & ~n914;
  assign n916 = ~reg_controllable_hgrant3_out & ~n915;
  assign n917 = ~n583 & ~n916;
  assign n918 = ~next_sys_fair<2>_out  & ~n917;
  assign n919 = ~n911 & ~n918;
  assign n920 = ~reg_controllable_hgrant4_out & ~n919;
  assign n921 = ~n626 & ~n920;
  assign n922 = ~reg_controllable_hgrant5_out & ~n921;
  assign n923 = ~n623 & ~n922;
  assign n924 = next_sys_fair<0>_out  & ~n923;
  assign n925 = ~reg_controllable_hgrant4_out & ~n903;
  assign n926 = ~n646 & ~n925;
  assign n927 = ~reg_controllable_hgrant5_out & ~n926;
  assign n928 = ~n643 & ~n927;
  assign n929 = ~next_sys_fair<0>_out  & ~n928;
  assign n930 = ~n924 & ~n929;
  assign n931 = ~next_sys_fair<3>_out  & ~n930;
  assign n932 = ~n910 & ~n931;
  assign n933 = ~reg_controllable_hmaster2_out & ~n932;
  assign n934 = ~n897 & ~n933;
  assign n935 = ~reg_controllable_hmaster1_out & ~n934;
  assign n936 = ~n874 & ~n935;
  assign n937 = next_sys_fair<1>_out  & ~n936;
  assign n938 = reg_controllable_hmaster2_out & ~n835;
  assign n939 = ~reg_stateG10_3_out & ~n230;
  assign n940 = ~reg_stateG10_3_out & ~n939;
  assign n941 = reg_controllable_hgrant3_out & ~n940;
  assign n942 = ~n671 & ~n941;
  assign n943 = next_sys_fair<2>_out  & ~n942;
  assign n944 = ~reg_stateG10_3_out & ~n345;
  assign n945 = ~reg_stateG10_3_out & ~n944;
  assign n946 = reg_controllable_hgrant3_out & ~n945;
  assign n947 = ~n812 & ~n946;
  assign n948 = ~next_sys_fair<2>_out  & ~n947;
  assign n949 = ~n943 & ~n948;
  assign n950 = ~reg_controllable_hgrant4_out & ~n949;
  assign n951 = ~n709 & ~n950;
  assign n952 = ~reg_controllable_hgrant5_out & ~n951;
  assign n953 = ~n706 & ~n952;
  assign n954 = next_sys_fair<0>_out  & ~n953;
  assign n955 = ~n824 & ~n846;
  assign n956 = next_sys_fair<2>_out  & ~n955;
  assign n957 = ~reg_stateG10_3_out & ~n376;
  assign n958 = ~reg_stateG10_3_out & ~n957;
  assign n959 = reg_controllable_hgrant3_out & ~n958;
  assign n960 = ~n812 & ~n959;
  assign n961 = ~next_sys_fair<2>_out  & ~n960;
  assign n962 = ~n956 & ~n961;
  assign n963 = ~reg_controllable_hgrant4_out & ~n962;
  assign n964 = ~n709 & ~n963;
  assign n965 = ~reg_controllable_hgrant5_out & ~n964;
  assign n966 = ~n706 & ~n965;
  assign n967 = ~next_sys_fair<0>_out  & ~n966;
  assign n968 = ~n954 & ~n967;
  assign n969 = ~next_sys_fair<3>_out  & ~n968;
  assign n970 = ~n854 & ~n969;
  assign n971 = ~reg_controllable_hmaster2_out & ~n970;
  assign n972 = ~n938 & ~n971;
  assign n973 = reg_controllable_hmaster1_out & ~n972;
  assign n974 = ~reg_stateG10_5_out & ~n351;
  assign n975 = ~reg_stateG10_5_out & ~n974;
  assign n976 = reg_controllable_hgrant5_out & ~n975;
  assign n977 = ~n818 & ~n976;
  assign n978 = next_sys_fair<0>_out  & ~n977;
  assign n979 = ~reg_stateG10_5_out & ~n382;
  assign n980 = ~reg_stateG10_5_out & ~n979;
  assign n981 = reg_controllable_hgrant5_out & ~n980;
  assign n982 = ~n830 & ~n981;
  assign n983 = ~next_sys_fair<0>_out  & ~n982;
  assign n984 = ~n978 & ~n983;
  assign n985 = ~next_sys_fair<3>_out  & ~n984;
  assign n986 = ~n879 & ~n985;
  assign n987 = reg_controllable_hmaster2_out & ~n986;
  assign n988 = ~n712 & ~n902;
  assign n989 = next_sys_fair<2>_out  & ~n988;
  assign n990 = ~reg_stateG10_1_out & ~n343;
  assign n991 = ~reg_stateG10_1_out & ~n990;
  assign n992 = reg_controllable_hgrant1_out & ~n991;
  assign n993 = ~n810 & ~n992;
  assign n994 = ~reg_controllable_hgrant3_out & ~n993;
  assign n995 = ~n712 & ~n994;
  assign n996 = ~next_sys_fair<2>_out  & ~n995;
  assign n997 = ~n989 & ~n996;
  assign n998 = ~reg_controllable_hgrant4_out & ~n997;
  assign n999 = ~n709 & ~n998;
  assign n1000 = ~reg_controllable_hgrant5_out & ~n999;
  assign n1001 = ~n706 & ~n1000;
  assign n1002 = next_sys_fair<0>_out  & ~n1001;
  assign n1003 = ~n822 & ~n900;
  assign n1004 = ~reg_controllable_hgrant3_out & ~n1003;
  assign n1005 = ~n583 & ~n1004;
  assign n1006 = next_sys_fair<2>_out  & ~n1005;
  assign n1007 = ~reg_stateG10_1_out & ~n374;
  assign n1008 = ~reg_stateG10_1_out & ~n1007;
  assign n1009 = reg_controllable_hgrant1_out & ~n1008;
  assign n1010 = ~n810 & ~n1009;
  assign n1011 = ~reg_controllable_hgrant3_out & ~n1010;
  assign n1012 = ~n712 & ~n1011;
  assign n1013 = ~next_sys_fair<2>_out  & ~n1012;
  assign n1014 = ~n1006 & ~n1013;
  assign n1015 = ~reg_controllable_hgrant4_out & ~n1014;
  assign n1016 = ~n709 & ~n1015;
  assign n1017 = ~reg_controllable_hgrant5_out & ~n1016;
  assign n1018 = ~n706 & ~n1017;
  assign n1019 = ~next_sys_fair<0>_out  & ~n1018;
  assign n1020 = ~n1002 & ~n1019;
  assign n1021 = ~next_sys_fair<3>_out  & ~n1020;
  assign n1022 = ~n910 & ~n1021;
  assign n1023 = ~reg_controllable_hmaster2_out & ~n1022;
  assign n1024 = ~n987 & ~n1023;
  assign n1025 = ~reg_controllable_hmaster1_out & ~n1024;
  assign n1026 = ~n973 & ~n1025;
  assign n1027 = ~next_sys_fair<1>_out  & ~n1026;
  assign n1028 = ~n937 & ~n1027;
  assign n1029 = reg_controllable_hmaster0_out & ~n1028;
  assign n1030 = ~reg_stateG10_2_out & ~n279;
  assign n1031 = ~reg_stateG10_2_out & ~n1030;
  assign n1032 = reg_controllable_hgrant2_out & ~n1031;
  assign n1033 = ~n667 & ~n1032;
  assign n1034 = ~reg_controllable_hgrant1_out & ~n1033;
  assign n1035 = ~n586 & ~n1034;
  assign n1036 = ~reg_controllable_hgrant3_out & ~n1035;
  assign n1037 = ~n583 & ~n1036;
  assign n1038 = ~next_sys_fair<2>_out  & ~n1037;
  assign n1039 = ~n663 & ~n1038;
  assign n1040 = ~reg_controllable_hgrant4_out & ~n1039;
  assign n1041 = ~n540 & ~n1040;
  assign n1042 = ~reg_controllable_hgrant5_out & ~n1041;
  assign n1043 = ~n537 & ~n1042;
  assign n1044 = next_sys_fair<3>_out  & ~n1043;
  assign n1045 = next_sys_fair<2>_out  & ~n1037;
  assign n1046 = ~n630 & ~n1034;
  assign n1047 = ~reg_controllable_hgrant3_out & ~n1046;
  assign n1048 = ~n583 & ~n1047;
  assign n1049 = ~next_sys_fair<2>_out  & ~n1048;
  assign n1050 = ~n1045 & ~n1049;
  assign n1051 = ~reg_controllable_hgrant4_out & ~n1050;
  assign n1052 = ~n626 & ~n1051;
  assign n1053 = ~reg_controllable_hgrant5_out & ~n1052;
  assign n1054 = ~n623 & ~n1053;
  assign n1055 = next_sys_fair<0>_out  & ~n1054;
  assign n1056 = ~reg_controllable_hgrant4_out & ~n1037;
  assign n1057 = ~n646 & ~n1056;
  assign n1058 = ~reg_controllable_hgrant5_out & ~n1057;
  assign n1059 = ~n643 & ~n1058;
  assign n1060 = ~next_sys_fair<0>_out  & ~n1059;
  assign n1061 = ~n1055 & ~n1060;
  assign n1062 = ~next_sys_fair<3>_out  & ~n1061;
  assign n1063 = ~n1044 & ~n1062;
  assign n1064 = ~reg_controllable_hmaster2_out & ~n1063;
  assign n1065 = ~n843 & ~n1064;
  assign n1066 = reg_controllable_hmaster1_out & ~n1065;
  assign n1067 = ~reg_stateG10_4_out & ~n287;
  assign n1068 = ~reg_stateG10_4_out & ~n1067;
  assign n1069 = reg_controllable_hgrant4_out & ~n1068;
  assign n1070 = ~n675 & ~n1069;
  assign n1071 = ~reg_controllable_hgrant5_out & ~n1070;
  assign n1072 = ~n537 & ~n1071;
  assign n1073 = next_sys_fair<3>_out  & ~n1072;
  assign n1074 = ~reg_stateG10_4_out & ~n285;
  assign n1075 = ~reg_stateG10_4_out & ~n1074;
  assign n1076 = reg_controllable_hgrant4_out & ~n1075;
  assign n1077 = ~n686 & ~n1076;
  assign n1078 = ~reg_controllable_hgrant5_out & ~n1077;
  assign n1079 = ~n623 & ~n1078;
  assign n1080 = next_sys_fair<0>_out  & ~n1079;
  assign n1081 = ~reg_stateG10_4_out & ~n881;
  assign n1082 = ~reg_stateG10_4_out & ~n1081;
  assign n1083 = reg_controllable_hgrant4_out & ~n1082;
  assign n1084 = ~n691 & ~n1083;
  assign n1085 = ~reg_controllable_hgrant5_out & ~n1084;
  assign n1086 = ~n643 & ~n1085;
  assign n1087 = ~next_sys_fair<0>_out  & ~n1086;
  assign n1088 = ~n1080 & ~n1087;
  assign n1089 = ~next_sys_fair<3>_out  & ~n1088;
  assign n1090 = ~n1073 & ~n1089;
  assign n1091 = reg_controllable_hmaster2_out & ~n1090;
  assign n1092 = ~n699 & ~n1091;
  assign n1093 = ~reg_controllable_hmaster1_out & ~n1092;
  assign n1094 = ~n1066 & ~n1093;
  assign n1095 = next_sys_fair<1>_out  & ~n1094;
  assign n1096 = ~n712 & ~n1036;
  assign n1097 = next_sys_fair<2>_out  & ~n1096;
  assign n1098 = ~reg_stateG10_2_out & ~n341;
  assign n1099 = ~reg_stateG10_2_out & ~n1098;
  assign n1100 = reg_controllable_hgrant2_out & ~n1099;
  assign n1101 = ~n808 & ~n1100;
  assign n1102 = ~reg_controllable_hgrant1_out & ~n1101;
  assign n1103 = ~n630 & ~n1102;
  assign n1104 = ~reg_controllable_hgrant3_out & ~n1103;
  assign n1105 = ~n712 & ~n1104;
  assign n1106 = ~next_sys_fair<2>_out  & ~n1105;
  assign n1107 = ~n1097 & ~n1106;
  assign n1108 = ~reg_controllable_hgrant4_out & ~n1107;
  assign n1109 = ~n709 & ~n1108;
  assign n1110 = ~reg_controllable_hgrant5_out & ~n1109;
  assign n1111 = ~n706 & ~n1110;
  assign n1112 = next_sys_fair<0>_out  & ~n1111;
  assign n1113 = ~reg_stateG10_2_out & ~n226;
  assign n1114 = ~reg_stateG10_2_out & ~n1113;
  assign n1115 = reg_controllable_hgrant2_out & ~n1114;
  assign n1116 = ~n667 & ~n1115;
  assign n1117 = ~reg_controllable_hgrant1_out & ~n1116;
  assign n1118 = ~n586 & ~n1117;
  assign n1119 = ~reg_controllable_hgrant3_out & ~n1118;
  assign n1120 = ~n583 & ~n1119;
  assign n1121 = next_sys_fair<2>_out  & ~n1120;
  assign n1122 = ~reg_stateG10_2_out & ~n372;
  assign n1123 = ~reg_stateG10_2_out & ~n1122;
  assign n1124 = reg_controllable_hgrant2_out & ~n1123;
  assign n1125 = ~n808 & ~n1124;
  assign n1126 = ~reg_controllable_hgrant1_out & ~n1125;
  assign n1127 = ~n630 & ~n1126;
  assign n1128 = ~reg_controllable_hgrant3_out & ~n1127;
  assign n1129 = ~n712 & ~n1128;
  assign n1130 = ~next_sys_fair<2>_out  & ~n1129;
  assign n1131 = ~n1121 & ~n1130;
  assign n1132 = ~reg_controllable_hgrant4_out & ~n1131;
  assign n1133 = ~n709 & ~n1132;
  assign n1134 = ~reg_controllable_hgrant5_out & ~n1133;
  assign n1135 = ~n706 & ~n1134;
  assign n1136 = ~next_sys_fair<0>_out  & ~n1135;
  assign n1137 = ~n1112 & ~n1136;
  assign n1138 = ~next_sys_fair<3>_out  & ~n1137;
  assign n1139 = ~n1044 & ~n1138;
  assign n1140 = ~reg_controllable_hmaster2_out & ~n1139;
  assign n1141 = ~n938 & ~n1140;
  assign n1142 = reg_controllable_hmaster1_out & ~n1141;
  assign n1143 = ~reg_stateG10_4_out & ~n349;
  assign n1144 = ~reg_stateG10_4_out & ~n1143;
  assign n1145 = reg_controllable_hgrant4_out & ~n1144;
  assign n1146 = ~n816 & ~n1145;
  assign n1147 = ~reg_controllable_hgrant5_out & ~n1146;
  assign n1148 = ~n706 & ~n1147;
  assign n1149 = next_sys_fair<0>_out  & ~n1148;
  assign n1150 = ~reg_stateG10_4_out & ~n380;
  assign n1151 = ~reg_stateG10_4_out & ~n1150;
  assign n1152 = reg_controllable_hgrant4_out & ~n1151;
  assign n1153 = ~n828 & ~n1152;
  assign n1154 = ~reg_controllable_hgrant5_out & ~n1153;
  assign n1155 = ~n706 & ~n1154;
  assign n1156 = ~next_sys_fair<0>_out  & ~n1155;
  assign n1157 = ~n1149 & ~n1156;
  assign n1158 = ~next_sys_fair<3>_out  & ~n1157;
  assign n1159 = ~n1073 & ~n1158;
  assign n1160 = reg_controllable_hmaster2_out & ~n1159;
  assign n1161 = ~n836 & ~n1160;
  assign n1162 = ~reg_controllable_hmaster1_out & ~n1161;
  assign n1163 = ~n1142 & ~n1162;
  assign n1164 = ~next_sys_fair<1>_out  & ~n1163;
  assign n1165 = ~n1095 & ~n1164;
  assign n1166 = ~reg_controllable_hmaster0_out & ~n1165;
  assign n1167 = ~n1029 & ~n1166;
  assign n1168 = ~reg_controllable_hmaster3_out & ~n1167;
  assign n1169 = ~n842 & ~n1168;
  assign n1170 = ~reg_controllable_hgrant6_out & ~n1169;
  assign n1171 = ~n534 & ~n1170;
  assign n1172 = ~reg_controllable_hgrant8_out & ~n1171;
  assign n1173 = ~n505 & ~n1172;
  assign n1174 = ~reg_controllable_hgrant7_out & ~n1173;
  assign n1175 = ~n464 & ~n1174;
  assign n1176 = ~reg_controllable_hgrant9_out & ~n1175;
  assign n1177 = ~n412 & ~n1176;
  assign n1178 = reg_controllable_nhgrant0_out & ~n1177;
  assign n1179 = next_sys_fair<0>_out  & ~n203;
  assign n1180 = ~next_sys_fair<0>_out  & ~n316;
  assign n1181 = ~n1179 & ~n1180;
  assign n1182 = ~next_sys_fair<3>_out  & ~n1181;
  assign n1183 = ~n413 & ~n1182;
  assign n1184 = next_sys_fair<1>_out  & ~n1183;
  assign n1185 = ~n472 & ~n1184;
  assign n1186 = reg_controllable_hmaster3_out & ~n1185;
  assign n1187 = reg_controllable_hmaster0_out & ~n1185;
  assign n1188 = reg_controllable_hmaster1_out & ~n1183;
  assign n1189 = reg_controllable_hmaster2_out & ~n1183;
  assign n1190 = next_sys_fair<0>_out  & ~n300;
  assign n1191 = ~n233 & ~n324;
  assign n1192 = ~reg_controllable_hgrant4_out & ~n1191;
  assign n1193 = ~reg_controllable_hgrant4_out & ~n1192;
  assign n1194 = ~reg_controllable_hgrant5_out & ~n1193;
  assign n1195 = ~reg_controllable_hgrant5_out & ~n1194;
  assign n1196 = ~next_sys_fair<0>_out  & ~n1195;
  assign n1197 = ~n1190 & ~n1196;
  assign n1198 = ~next_sys_fair<3>_out  & ~n1197;
  assign n1199 = ~n426 & ~n1198;
  assign n1200 = ~reg_controllable_hmaster2_out & ~n1199;
  assign n1201 = ~n1189 & ~n1200;
  assign n1202 = ~reg_controllable_hmaster1_out & ~n1201;
  assign n1203 = ~n1188 & ~n1202;
  assign n1204 = next_sys_fair<1>_out  & ~n1203;
  assign n1205 = ~n494 & ~n1204;
  assign n1206 = ~reg_controllable_hmaster0_out & ~n1205;
  assign n1207 = ~n1187 & ~n1206;
  assign n1208 = ~reg_controllable_hmaster3_out & ~n1207;
  assign n1209 = ~n1186 & ~n1208;
  assign n1210 = ~reg_controllable_hgrant6_out & ~n1209;
  assign n1211 = ~reg_controllable_hgrant6_out & ~n1210;
  assign n1212 = ~reg_controllable_hgrant8_out & ~n1211;
  assign n1213 = ~reg_controllable_hgrant8_out & ~n1212;
  assign n1214 = ~reg_controllable_hgrant7_out & ~n1213;
  assign n1215 = ~reg_controllable_hgrant7_out & ~n1214;
  assign n1216 = ~reg_controllable_hgrant9_out & ~n1215;
  assign n1217 = ~reg_controllable_hgrant9_out & ~n1216;
  assign n1218 = ~reg_controllable_nhgrant0_out & ~n1217;
  assign n1219 = ~n1178 & ~n1218;
  assign n1220 = reg_i_hready_out & ~n1219;
  assign n1221 = next_env_fair_out & ~n174;
  assign n1222 = ~next_env_fair_out & ~n117;
  assign n1223 = ~n1221 & ~n1222;
  assign n1224 = reg_stateA1_out & ~n1223;
  assign n1225 = reg_stateA1_out & ~n1224;
  assign n1226 = reg_controllable_hmastlock_out & ~n1225;
  assign n1227 = ~reg_stateA1_out & ~n174;
  assign n1228 = ~n1224 & ~n1227;
  assign n1229 = ~reg_controllable_hmastlock_out & ~n1228;
  assign n1230 = ~n1226 & ~n1229;
  assign n1231 = reg_controllable_locked_out & ~n1230;
  assign n1232 = ~reg_controllable_locked_out & ~n1228;
  assign n1233 = ~n1231 & ~n1232;
  assign n1234 = ~reg_controllable_hgrant2_out & ~n1233;
  assign n1235 = ~reg_controllable_hgrant2_out & ~n1234;
  assign n1236 = ~reg_controllable_hgrant1_out & ~n1235;
  assign n1237 = ~reg_controllable_hgrant1_out & ~n1236;
  assign n1238 = ~reg_controllable_hgrant3_out & ~n1237;
  assign n1239 = ~reg_controllable_hgrant3_out & ~n1238;
  assign n1240 = ~next_sys_fair<2>_out  & ~n1239;
  assign n1241 = ~next_sys_fair<2>_out  & ~n1240;
  assign n1242 = ~reg_controllable_hgrant4_out & ~n1241;
  assign n1243 = ~reg_controllable_hgrant4_out & ~n1242;
  assign n1244 = ~reg_controllable_hgrant5_out & ~n1243;
  assign n1245 = ~reg_controllable_hgrant5_out & ~n1244;
  assign n1246 = ~reg_stateG10_9_out & ~n1245;
  assign n1247 = ~reg_stateG10_9_out & ~n1246;
  assign n1248 = next_sys_fair<0>_out  & ~n1247;
  assign n1249 = ~next_env_fair_out & ~n149;
  assign n1250 = ~next_env_fair_out & ~n1249;
  assign n1251 = reg_stateA1_out & ~n1250;
  assign n1252 = reg_stateA1_out & ~n1251;
  assign n1253 = reg_controllable_hmastlock_out & ~n1252;
  assign n1254 = ~reg_controllable_hmastlock_out & ~n1250;
  assign n1255 = ~n1253 & ~n1254;
  assign n1256 = reg_controllable_locked_out & ~n1255;
  assign n1257 = next_env_fair_out & ~n165;
  assign n1258 = ~next_env_fair_out & ~n174;
  assign n1259 = ~n1257 & ~n1258;
  assign n1260 = ~reg_controllable_locked_out & ~n1259;
  assign n1261 = ~n1256 & ~n1260;
  assign n1262 = ~reg_controllable_hgrant2_out & ~n1261;
  assign n1263 = ~reg_controllable_hgrant2_out & ~n1262;
  assign n1264 = ~reg_controllable_hgrant1_out & ~n1263;
  assign n1265 = ~reg_controllable_hgrant1_out & ~n1264;
  assign n1266 = ~reg_controllable_hgrant3_out & ~n1265;
  assign n1267 = ~reg_controllable_hgrant3_out & ~n1266;
  assign n1268 = ~next_sys_fair<2>_out  & ~n1267;
  assign n1269 = ~next_sys_fair<2>_out  & ~n1268;
  assign n1270 = ~reg_controllable_hgrant4_out & ~n1269;
  assign n1271 = ~reg_controllable_hgrant4_out & ~n1270;
  assign n1272 = ~reg_controllable_hgrant5_out & ~n1271;
  assign n1273 = ~reg_controllable_hgrant5_out & ~n1272;
  assign n1274 = ~reg_stateG10_9_out & ~n1273;
  assign n1275 = ~reg_stateG10_9_out & ~n1274;
  assign n1276 = ~next_sys_fair<0>_out  & ~n1275;
  assign n1277 = ~n1248 & ~n1276;
  assign n1278 = next_sys_fair<3>_out  & ~n1277;
  assign n1279 = ~reg_controllable_hgrant4_out & ~n1267;
  assign n1280 = ~reg_controllable_hgrant4_out & ~n1279;
  assign n1281 = ~reg_controllable_hgrant5_out & ~n1280;
  assign n1282 = ~reg_controllable_hgrant5_out & ~n1281;
  assign n1283 = ~reg_stateG10_9_out & ~n1282;
  assign n1284 = ~reg_stateG10_9_out & ~n1283;
  assign n1285 = ~next_sys_fair<3>_out  & ~n1284;
  assign n1286 = ~n1278 & ~n1285;
  assign n1287 = reg_controllable_hmaster1_out & ~n1286;
  assign n1288 = reg_controllable_hmaster2_out & ~n1286;
  assign n1289 = ~reg_stateG2_out & ~n117;
  assign n1290 = ~reg_stateG2_out & ~n1289;
  assign n1291 = ~reg_stateA1_out & ~n1290;
  assign n1292 = ~reg_stateA1_out & ~n1291;
  assign n1293 = ~reg_controllable_hmastlock_out & ~n1292;
  assign n1294 = ~n218 & ~n1293;
  assign n1295 = reg_controllable_locked_out & ~n1294;
  assign n1296 = reg_controllable_hmastlock_out & ~n1290;
  assign n1297 = ~n223 & ~n1296;
  assign n1298 = ~reg_controllable_locked_out & ~n1297;
  assign n1299 = ~n1295 & ~n1298;
  assign n1300 = ~reg_controllable_hgrant2_out & ~n1299;
  assign n1301 = ~reg_controllable_hgrant2_out & ~n1300;
  assign n1302 = ~reg_controllable_hgrant1_out & ~n1301;
  assign n1303 = ~reg_controllable_hgrant1_out & ~n1302;
  assign n1304 = ~reg_controllable_hgrant3_out & ~n1303;
  assign n1305 = ~reg_controllable_hgrant3_out & ~n1304;
  assign n1306 = ~next_sys_fair<2>_out  & ~n1305;
  assign n1307 = ~next_sys_fair<2>_out  & ~n1306;
  assign n1308 = ~reg_controllable_hgrant4_out & ~n1307;
  assign n1309 = ~reg_controllable_hgrant4_out & ~n1308;
  assign n1310 = ~reg_controllable_hgrant5_out & ~n1309;
  assign n1311 = ~reg_controllable_hgrant5_out & ~n1310;
  assign n1312 = ~reg_stateG10_9_out & ~n1311;
  assign n1313 = ~reg_stateG10_9_out & ~n1312;
  assign n1314 = next_sys_fair<0>_out  & ~n1313;
  assign n1315 = ~reg_stateG2_out & ~n1250;
  assign n1316 = ~reg_stateG2_out & ~n1315;
  assign n1317 = ~reg_stateA1_out & ~n1316;
  assign n1318 = ~reg_stateA1_out & ~n1317;
  assign n1319 = ~reg_controllable_hmastlock_out & ~n1318;
  assign n1320 = ~n271 & ~n1319;
  assign n1321 = reg_controllable_locked_out & ~n1320;
  assign n1322 = ~reg_stateG2_out & ~n1259;
  assign n1323 = ~reg_stateG2_out & ~n1322;
  assign n1324 = reg_controllable_hmastlock_out & ~n1323;
  assign n1325 = ~n276 & ~n1324;
  assign n1326 = ~reg_controllable_locked_out & ~n1325;
  assign n1327 = ~n1321 & ~n1326;
  assign n1328 = ~reg_controllable_hgrant2_out & ~n1327;
  assign n1329 = ~reg_controllable_hgrant2_out & ~n1328;
  assign n1330 = ~reg_controllable_hgrant1_out & ~n1329;
  assign n1331 = ~reg_controllable_hgrant1_out & ~n1330;
  assign n1332 = ~reg_controllable_hgrant3_out & ~n1331;
  assign n1333 = ~reg_controllable_hgrant3_out & ~n1332;
  assign n1334 = ~next_sys_fair<2>_out  & ~n1333;
  assign n1335 = ~next_sys_fair<2>_out  & ~n1334;
  assign n1336 = ~reg_controllable_hgrant4_out & ~n1335;
  assign n1337 = ~reg_controllable_hgrant4_out & ~n1336;
  assign n1338 = ~reg_controllable_hgrant5_out & ~n1337;
  assign n1339 = ~reg_controllable_hgrant5_out & ~n1338;
  assign n1340 = ~reg_stateG10_9_out & ~n1339;
  assign n1341 = ~reg_stateG10_9_out & ~n1340;
  assign n1342 = ~next_sys_fair<0>_out  & ~n1341;
  assign n1343 = ~n1314 & ~n1342;
  assign n1344 = next_sys_fair<3>_out  & ~n1343;
  assign n1345 = ~reg_controllable_hgrant4_out & ~n1333;
  assign n1346 = ~reg_controllable_hgrant4_out & ~n1345;
  assign n1347 = ~reg_controllable_hgrant5_out & ~n1346;
  assign n1348 = ~reg_controllable_hgrant5_out & ~n1347;
  assign n1349 = ~reg_stateG10_9_out & ~n1348;
  assign n1350 = ~reg_stateG10_9_out & ~n1349;
  assign n1351 = ~next_sys_fair<3>_out  & ~n1350;
  assign n1352 = ~n1344 & ~n1351;
  assign n1353 = ~reg_controllable_hmaster2_out & ~n1352;
  assign n1354 = ~n1288 & ~n1353;
  assign n1355 = ~reg_controllable_hmaster1_out & ~n1354;
  assign n1356 = ~n1287 & ~n1355;
  assign n1357 = next_sys_fair<1>_out  & ~n1356;
  assign n1358 = next_sys_fair<3>_out  & ~n1275;
  assign n1359 = next_sys_fair<2>_out  & ~n1267;
  assign n1360 = ~n118 & ~n258;
  assign n1361 = next_env_fair_out & ~n1360;
  assign n1362 = ~n1222 & ~n1361;
  assign n1363 = reg_stateA1_out & ~n1362;
  assign n1364 = reg_stateA1_out & ~n1363;
  assign n1365 = reg_controllable_hmastlock_out & ~n1364;
  assign n1366 = ~reg_stateA1_out & ~n1360;
  assign n1367 = ~n1363 & ~n1366;
  assign n1368 = ~reg_controllable_hmastlock_out & ~n1367;
  assign n1369 = ~n1365 & ~n1368;
  assign n1370 = reg_controllable_locked_out & ~n1369;
  assign n1371 = ~reg_controllable_locked_out & ~n1367;
  assign n1372 = ~n1370 & ~n1371;
  assign n1373 = ~reg_controllable_hgrant2_out & ~n1372;
  assign n1374 = ~reg_controllable_hgrant2_out & ~n1373;
  assign n1375 = ~reg_controllable_hgrant1_out & ~n1374;
  assign n1376 = ~reg_controllable_hgrant1_out & ~n1375;
  assign n1377 = ~reg_controllable_hgrant3_out & ~n1376;
  assign n1378 = ~reg_controllable_hgrant3_out & ~n1377;
  assign n1379 = ~next_sys_fair<2>_out  & ~n1378;
  assign n1380 = ~n1359 & ~n1379;
  assign n1381 = ~reg_controllable_hgrant4_out & ~n1380;
  assign n1382 = ~reg_controllable_hgrant4_out & ~n1381;
  assign n1383 = ~reg_controllable_hgrant5_out & ~n1382;
  assign n1384 = ~reg_controllable_hgrant5_out & ~n1383;
  assign n1385 = ~reg_stateG10_9_out & ~n1384;
  assign n1386 = ~reg_stateG10_9_out & ~n1385;
  assign n1387 = next_sys_fair<0>_out  & ~n1386;
  assign n1388 = reg_stateG2_out & ~n1223;
  assign n1389 = ~n1289 & ~n1388;
  assign n1390 = reg_stateA1_out & ~n1389;
  assign n1391 = reg_stateA1_out & ~n1390;
  assign n1392 = reg_controllable_hmastlock_out & ~n1391;
  assign n1393 = ~reg_controllable_hmastlock_out & ~n1389;
  assign n1394 = ~n1392 & ~n1393;
  assign n1395 = reg_controllable_locked_out & ~n1394;
  assign n1396 = ~reg_controllable_locked_out & ~n1389;
  assign n1397 = ~n1395 & ~n1396;
  assign n1398 = ~reg_controllable_hgrant2_out & ~n1397;
  assign n1399 = ~reg_controllable_hgrant2_out & ~n1398;
  assign n1400 = ~reg_controllable_hgrant1_out & ~n1399;
  assign n1401 = ~reg_controllable_hgrant1_out & ~n1400;
  assign n1402 = ~reg_controllable_hgrant3_out & ~n1401;
  assign n1403 = ~reg_controllable_hgrant3_out & ~n1402;
  assign n1404 = ~next_sys_fair<2>_out  & ~n1403;
  assign n1405 = ~n1359 & ~n1404;
  assign n1406 = ~reg_controllable_hgrant4_out & ~n1405;
  assign n1407 = ~reg_controllable_hgrant4_out & ~n1406;
  assign n1408 = ~reg_controllable_hgrant5_out & ~n1407;
  assign n1409 = ~reg_controllable_hgrant5_out & ~n1408;
  assign n1410 = ~reg_stateG10_9_out & ~n1409;
  assign n1411 = ~reg_stateG10_9_out & ~n1410;
  assign n1412 = ~next_sys_fair<0>_out  & ~n1411;
  assign n1413 = ~n1387 & ~n1412;
  assign n1414 = ~next_sys_fair<3>_out  & ~n1413;
  assign n1415 = ~n1358 & ~n1414;
  assign n1416 = reg_controllable_hmaster1_out & ~n1415;
  assign n1417 = reg_controllable_hmaster2_out & ~n1415;
  assign n1418 = next_sys_fair<3>_out  & ~n1341;
  assign n1419 = next_sys_fair<2>_out  & ~n1333;
  assign n1420 = ~reg_stateG2_out & ~n1360;
  assign n1421 = ~reg_stateG2_out & ~n1420;
  assign n1422 = ~reg_stateA1_out & ~n1421;
  assign n1423 = ~reg_stateA1_out & ~n1422;
  assign n1424 = ~reg_controllable_hmastlock_out & ~n1423;
  assign n1425 = ~n335 & ~n1424;
  assign n1426 = reg_controllable_locked_out & ~n1425;
  assign n1427 = reg_controllable_hmastlock_out & ~n1421;
  assign n1428 = ~n338 & ~n1427;
  assign n1429 = ~reg_controllable_locked_out & ~n1428;
  assign n1430 = ~n1426 & ~n1429;
  assign n1431 = ~reg_controllable_hgrant2_out & ~n1430;
  assign n1432 = ~reg_controllable_hgrant2_out & ~n1431;
  assign n1433 = ~reg_controllable_hgrant1_out & ~n1432;
  assign n1434 = ~reg_controllable_hgrant1_out & ~n1433;
  assign n1435 = ~reg_controllable_hgrant3_out & ~n1434;
  assign n1436 = ~reg_controllable_hgrant3_out & ~n1435;
  assign n1437 = ~next_sys_fair<2>_out  & ~n1436;
  assign n1438 = ~n1419 & ~n1437;
  assign n1439 = ~reg_controllable_hgrant4_out & ~n1438;
  assign n1440 = ~reg_controllable_hgrant4_out & ~n1439;
  assign n1441 = ~reg_controllable_hgrant5_out & ~n1440;
  assign n1442 = ~reg_controllable_hgrant5_out & ~n1441;
  assign n1443 = ~reg_stateG10_9_out & ~n1442;
  assign n1444 = ~reg_stateG10_9_out & ~n1443;
  assign n1445 = next_sys_fair<0>_out  & ~n1444;
  assign n1446 = ~n366 & ~n1293;
  assign n1447 = reg_controllable_locked_out & ~n1446;
  assign n1448 = ~n369 & ~n1296;
  assign n1449 = ~reg_controllable_locked_out & ~n1448;
  assign n1450 = ~n1447 & ~n1449;
  assign n1451 = ~reg_controllable_hgrant2_out & ~n1450;
  assign n1452 = ~reg_controllable_hgrant2_out & ~n1451;
  assign n1453 = ~reg_controllable_hgrant1_out & ~n1452;
  assign n1454 = ~reg_controllable_hgrant1_out & ~n1453;
  assign n1455 = ~reg_controllable_hgrant3_out & ~n1454;
  assign n1456 = ~reg_controllable_hgrant3_out & ~n1455;
  assign n1457 = ~next_sys_fair<2>_out  & ~n1456;
  assign n1458 = ~n1419 & ~n1457;
  assign n1459 = ~reg_controllable_hgrant4_out & ~n1458;
  assign n1460 = ~reg_controllable_hgrant4_out & ~n1459;
  assign n1461 = ~reg_controllable_hgrant5_out & ~n1460;
  assign n1462 = ~reg_controllable_hgrant5_out & ~n1461;
  assign n1463 = ~reg_stateG10_9_out & ~n1462;
  assign n1464 = ~reg_stateG10_9_out & ~n1463;
  assign n1465 = ~next_sys_fair<0>_out  & ~n1464;
  assign n1466 = ~n1445 & ~n1465;
  assign n1467 = ~next_sys_fair<3>_out  & ~n1466;
  assign n1468 = ~n1418 & ~n1467;
  assign n1469 = ~reg_controllable_hmaster2_out & ~n1468;
  assign n1470 = ~n1417 & ~n1469;
  assign n1471 = ~reg_controllable_hmaster1_out & ~n1470;
  assign n1472 = ~n1416 & ~n1471;
  assign n1473 = ~next_sys_fair<1>_out  & ~n1472;
  assign n1474 = ~n1357 & ~n1473;
  assign n1475 = reg_controllable_hmaster0_out & ~n1474;
  assign n1476 = ~reg_stateG2_out & ~n174;
  assign n1477 = ~reg_stateG2_out & ~n1476;
  assign n1478 = ~reg_stateA1_out & ~n1477;
  assign n1479 = ~reg_stateA1_out & ~n1478;
  assign n1480 = ~reg_controllable_hmastlock_out & ~n1479;
  assign n1481 = ~reg_controllable_hmastlock_out & ~n1480;
  assign n1482 = reg_controllable_locked_out & ~n1481;
  assign n1483 = ~reg_controllable_locked_out & ~n1477;
  assign n1484 = ~n1482 & ~n1483;
  assign n1485 = ~reg_controllable_hgrant2_out & ~n1484;
  assign n1486 = ~reg_controllable_hgrant2_out & ~n1485;
  assign n1487 = ~reg_controllable_hgrant1_out & ~n1486;
  assign n1488 = ~reg_controllable_hgrant1_out & ~n1487;
  assign n1489 = ~reg_controllable_hgrant3_out & ~n1488;
  assign n1490 = ~reg_controllable_hgrant3_out & ~n1489;
  assign n1491 = ~next_sys_fair<2>_out  & ~n1490;
  assign n1492 = ~next_sys_fair<2>_out  & ~n1491;
  assign n1493 = ~reg_controllable_hgrant4_out & ~n1492;
  assign n1494 = ~reg_controllable_hgrant4_out & ~n1493;
  assign n1495 = ~reg_controllable_hgrant5_out & ~n1494;
  assign n1496 = ~reg_controllable_hgrant5_out & ~n1495;
  assign n1497 = ~reg_stateG10_9_out & ~n1496;
  assign n1498 = ~reg_stateG10_9_out & ~n1497;
  assign n1499 = next_sys_fair<0>_out  & ~n1498;
  assign n1500 = ~reg_controllable_hmastlock_out & ~n1293;
  assign n1501 = reg_controllable_locked_out & ~n1500;
  assign n1502 = ~reg_controllable_locked_out & ~n1290;
  assign n1503 = ~n1501 & ~n1502;
  assign n1504 = ~reg_controllable_hgrant2_out & ~n1503;
  assign n1505 = ~reg_controllable_hgrant2_out & ~n1504;
  assign n1506 = ~reg_controllable_hgrant1_out & ~n1505;
  assign n1507 = ~reg_controllable_hgrant1_out & ~n1506;
  assign n1508 = ~reg_controllable_hgrant3_out & ~n1507;
  assign n1509 = ~reg_controllable_hgrant3_out & ~n1508;
  assign n1510 = ~next_sys_fair<2>_out  & ~n1509;
  assign n1511 = ~next_sys_fair<2>_out  & ~n1510;
  assign n1512 = ~reg_controllable_hgrant4_out & ~n1511;
  assign n1513 = ~reg_controllable_hgrant4_out & ~n1512;
  assign n1514 = ~reg_controllable_hgrant5_out & ~n1513;
  assign n1515 = ~reg_controllable_hgrant5_out & ~n1514;
  assign n1516 = ~reg_stateG10_9_out & ~n1515;
  assign n1517 = ~reg_stateG10_9_out & ~n1516;
  assign n1518 = ~next_sys_fair<0>_out  & ~n1517;
  assign n1519 = ~n1499 & ~n1518;
  assign n1520 = next_sys_fair<3>_out  & ~n1519;
  assign n1521 = ~reg_controllable_hmastlock_out & ~n1319;
  assign n1522 = reg_controllable_locked_out & ~n1521;
  assign n1523 = ~reg_controllable_locked_out & ~n1323;
  assign n1524 = ~n1522 & ~n1523;
  assign n1525 = ~reg_controllable_hgrant2_out & ~n1524;
  assign n1526 = ~reg_controllable_hgrant2_out & ~n1525;
  assign n1527 = ~reg_controllable_hgrant1_out & ~n1526;
  assign n1528 = ~reg_controllable_hgrant1_out & ~n1527;
  assign n1529 = ~reg_controllable_hgrant3_out & ~n1528;
  assign n1530 = ~reg_controllable_hgrant3_out & ~n1529;
  assign n1531 = ~reg_controllable_hgrant4_out & ~n1530;
  assign n1532 = ~reg_controllable_hgrant4_out & ~n1531;
  assign n1533 = ~reg_controllable_hgrant5_out & ~n1532;
  assign n1534 = ~reg_controllable_hgrant5_out & ~n1533;
  assign n1535 = ~reg_stateG10_9_out & ~n1534;
  assign n1536 = ~reg_stateG10_9_out & ~n1535;
  assign n1537 = ~next_sys_fair<3>_out  & ~n1536;
  assign n1538 = ~n1520 & ~n1537;
  assign n1539 = ~reg_controllable_hmaster2_out & ~n1538;
  assign n1540 = ~n1288 & ~n1539;
  assign n1541 = ~reg_controllable_hmaster1_out & ~n1540;
  assign n1542 = ~n1287 & ~n1541;
  assign n1543 = next_sys_fair<1>_out  & ~n1542;
  assign n1544 = ~next_sys_fair<2>_out  & ~n1530;
  assign n1545 = ~next_sys_fair<2>_out  & ~n1544;
  assign n1546 = ~reg_controllable_hgrant4_out & ~n1545;
  assign n1547 = ~reg_controllable_hgrant4_out & ~n1546;
  assign n1548 = ~reg_controllable_hgrant5_out & ~n1547;
  assign n1549 = ~reg_controllable_hgrant5_out & ~n1548;
  assign n1550 = ~reg_stateG10_9_out & ~n1549;
  assign n1551 = ~reg_stateG10_9_out & ~n1550;
  assign n1552 = next_sys_fair<3>_out  & ~n1551;
  assign n1553 = next_sys_fair<2>_out  & ~n1530;
  assign n1554 = ~reg_controllable_hmastlock_out & ~n1424;
  assign n1555 = reg_controllable_locked_out & ~n1554;
  assign n1556 = ~reg_controllable_locked_out & ~n1421;
  assign n1557 = ~n1555 & ~n1556;
  assign n1558 = ~reg_controllable_hgrant2_out & ~n1557;
  assign n1559 = ~reg_controllable_hgrant2_out & ~n1558;
  assign n1560 = ~reg_controllable_hgrant1_out & ~n1559;
  assign n1561 = ~reg_controllable_hgrant1_out & ~n1560;
  assign n1562 = ~reg_controllable_hgrant3_out & ~n1561;
  assign n1563 = ~reg_controllable_hgrant3_out & ~n1562;
  assign n1564 = ~next_sys_fair<2>_out  & ~n1563;
  assign n1565 = ~n1553 & ~n1564;
  assign n1566 = ~reg_controllable_hgrant4_out & ~n1565;
  assign n1567 = ~reg_controllable_hgrant4_out & ~n1566;
  assign n1568 = ~reg_controllable_hgrant5_out & ~n1567;
  assign n1569 = ~reg_controllable_hgrant5_out & ~n1568;
  assign n1570 = ~reg_stateG10_9_out & ~n1569;
  assign n1571 = ~reg_stateG10_9_out & ~n1570;
  assign n1572 = next_sys_fair<0>_out  & ~n1571;
  assign n1573 = ~n1510 & ~n1553;
  assign n1574 = ~reg_controllable_hgrant4_out & ~n1573;
  assign n1575 = ~reg_controllable_hgrant4_out & ~n1574;
  assign n1576 = ~reg_controllable_hgrant5_out & ~n1575;
  assign n1577 = ~reg_controllable_hgrant5_out & ~n1576;
  assign n1578 = ~reg_stateG10_9_out & ~n1577;
  assign n1579 = ~reg_stateG10_9_out & ~n1578;
  assign n1580 = ~next_sys_fair<0>_out  & ~n1579;
  assign n1581 = ~n1572 & ~n1580;
  assign n1582 = ~next_sys_fair<3>_out  & ~n1581;
  assign n1583 = ~n1552 & ~n1582;
  assign n1584 = ~reg_controllable_hmaster2_out & ~n1583;
  assign n1585 = ~n1417 & ~n1584;
  assign n1586 = ~reg_controllable_hmaster1_out & ~n1585;
  assign n1587 = ~n1416 & ~n1586;
  assign n1588 = ~next_sys_fair<1>_out  & ~n1587;
  assign n1589 = ~n1543 & ~n1588;
  assign n1590 = ~reg_controllable_hmaster0_out & ~n1589;
  assign n1591 = ~n1475 & ~n1590;
  assign n1592 = reg_controllable_hmaster3_out & ~n1591;
  assign n1593 = ~next_sys_fair<0>_out  & ~n1551;
  assign n1594 = ~n1499 & ~n1593;
  assign n1595 = next_sys_fair<3>_out  & ~n1594;
  assign n1596 = ~n1537 & ~n1595;
  assign n1597 = reg_controllable_hmaster1_out & ~n1596;
  assign n1598 = next_sys_fair<2>_out  & ~n1509;
  assign n1599 = ~n1544 & ~n1598;
  assign n1600 = ~reg_controllable_hgrant4_out & ~n1599;
  assign n1601 = ~reg_controllable_hgrant4_out & ~n1600;
  assign n1602 = ~reg_controllable_hgrant5_out & ~n1601;
  assign n1603 = ~reg_controllable_hgrant5_out & ~n1602;
  assign n1604 = ~reg_stateG10_9_out & ~n1603;
  assign n1605 = ~reg_stateG10_9_out & ~n1604;
  assign n1606 = next_sys_fair<0>_out  & ~n1605;
  assign n1607 = ~next_sys_fair<0>_out  & ~n1536;
  assign n1608 = ~n1606 & ~n1607;
  assign n1609 = ~next_sys_fair<3>_out  & ~n1608;
  assign n1610 = ~n1595 & ~n1609;
  assign n1611 = reg_controllable_hmaster2_out & ~n1610;
  assign n1612 = next_sys_fair<0>_out  & ~n1579;
  assign n1613 = ~n1607 & ~n1612;
  assign n1614 = ~next_sys_fair<3>_out  & ~n1613;
  assign n1615 = ~n1595 & ~n1614;
  assign n1616 = ~reg_controllable_hmaster2_out & ~n1615;
  assign n1617 = ~n1611 & ~n1616;
  assign n1618 = ~reg_controllable_hmaster1_out & ~n1617;
  assign n1619 = ~n1597 & ~n1618;
  assign n1620 = next_sys_fair<1>_out  & ~n1619;
  assign n1621 = next_sys_fair<0>_out  & ~n1517;
  assign n1622 = ~n1593 & ~n1621;
  assign n1623 = next_sys_fair<3>_out  & ~n1622;
  assign n1624 = ~n1582 & ~n1623;
  assign n1625 = reg_controllable_hmaster2_out & ~n1624;
  assign n1626 = ~n1564 & ~n1598;
  assign n1627 = ~reg_controllable_hgrant4_out & ~n1626;
  assign n1628 = ~reg_controllable_hgrant4_out & ~n1627;
  assign n1629 = ~reg_controllable_hgrant5_out & ~n1628;
  assign n1630 = ~reg_controllable_hgrant5_out & ~n1629;
  assign n1631 = ~reg_stateG10_9_out & ~n1630;
  assign n1632 = ~reg_stateG10_9_out & ~n1631;
  assign n1633 = next_sys_fair<0>_out  & ~n1632;
  assign n1634 = ~n1580 & ~n1633;
  assign n1635 = ~next_sys_fair<3>_out  & ~n1634;
  assign n1636 = ~n1552 & ~n1635;
  assign n1637 = ~reg_controllable_hmaster2_out & ~n1636;
  assign n1638 = ~n1625 & ~n1637;
  assign n1639 = reg_controllable_hmaster1_out & ~n1638;
  assign n1640 = ~reg_controllable_hmaster1_out & ~n1583;
  assign n1641 = ~n1639 & ~n1640;
  assign n1642 = ~next_sys_fair<1>_out  & ~n1641;
  assign n1643 = ~n1620 & ~n1642;
  assign n1644 = reg_controllable_hmaster0_out & ~n1643;
  assign n1645 = next_sys_fair<0>_out  & ~n1536;
  assign n1646 = ~next_sys_fair<0>_out  & ~n1605;
  assign n1647 = ~n1645 & ~n1646;
  assign n1648 = ~next_sys_fair<3>_out  & ~n1647;
  assign n1649 = ~n1595 & ~n1648;
  assign n1650 = reg_controllable_hmaster2_out & ~n1649;
  assign n1651 = ~n1580 & ~n1645;
  assign n1652 = ~next_sys_fair<3>_out  & ~n1651;
  assign n1653 = ~n1595 & ~n1652;
  assign n1654 = ~reg_controllable_hmaster2_out & ~n1653;
  assign n1655 = ~n1650 & ~n1654;
  assign n1656 = ~reg_controllable_hmaster1_out & ~n1655;
  assign n1657 = ~n1597 & ~n1656;
  assign n1658 = next_sys_fair<1>_out  & ~n1657;
  assign n1659 = next_sys_fair<0>_out  & ~n1551;
  assign n1660 = ~n1518 & ~n1659;
  assign n1661 = next_sys_fair<3>_out  & ~n1660;
  assign n1662 = ~n1582 & ~n1661;
  assign n1663 = reg_controllable_hmaster2_out & ~n1662;
  assign n1664 = ~reg_controllable_hgrant4_out & ~n1509;
  assign n1665 = ~reg_controllable_hgrant4_out & ~n1664;
  assign n1666 = ~reg_controllable_hgrant5_out & ~n1665;
  assign n1667 = ~reg_controllable_hgrant5_out & ~n1666;
  assign n1668 = ~reg_stateG10_9_out & ~n1667;
  assign n1669 = ~reg_stateG10_9_out & ~n1668;
  assign n1670 = ~next_sys_fair<0>_out  & ~n1669;
  assign n1671 = ~n1572 & ~n1670;
  assign n1672 = ~next_sys_fair<3>_out  & ~n1671;
  assign n1673 = ~n1552 & ~n1672;
  assign n1674 = ~reg_controllable_hmaster2_out & ~n1673;
  assign n1675 = ~n1663 & ~n1674;
  assign n1676 = reg_controllable_hmaster1_out & ~n1675;
  assign n1677 = ~n1640 & ~n1676;
  assign n1678 = ~next_sys_fair<1>_out  & ~n1677;
  assign n1679 = ~n1658 & ~n1678;
  assign n1680 = ~reg_controllable_hmaster0_out & ~n1679;
  assign n1681 = ~n1644 & ~n1680;
  assign n1682 = ~reg_controllable_hmaster3_out & ~n1681;
  assign n1683 = ~n1592 & ~n1682;
  assign n1684 = ~reg_controllable_hgrant6_out & ~n1683;
  assign n1685 = ~reg_controllable_hgrant6_out & ~n1684;
  assign n1686 = ~reg_controllable_hgrant8_out & ~n1685;
  assign n1687 = ~reg_controllable_hgrant8_out & ~n1686;
  assign n1688 = ~reg_controllable_hgrant7_out & ~n1687;
  assign n1689 = ~reg_controllable_hgrant7_out & ~n1688;
  assign n1690 = reg_controllable_hgrant9_out & ~n1689;
  assign n1691 = next_sys_fair<3>_out  & ~n1273;
  assign n1692 = ~next_sys_fair<3>_out  & ~n1282;
  assign n1693 = ~n1691 & ~n1692;
  assign n1694 = reg_controllable_hmaster1_out & ~n1693;
  assign n1695 = reg_controllable_hmaster2_out & ~n1693;
  assign n1696 = next_sys_fair<0>_out  & ~n1515;
  assign n1697 = ~next_sys_fair<0>_out  & ~n1549;
  assign n1698 = ~n1696 & ~n1697;
  assign n1699 = next_sys_fair<3>_out  & ~n1698;
  assign n1700 = ~next_sys_fair<3>_out  & ~n1534;
  assign n1701 = ~n1699 & ~n1700;
  assign n1702 = ~reg_controllable_hmaster2_out & ~n1701;
  assign n1703 = ~n1695 & ~n1702;
  assign n1704 = ~reg_controllable_hmaster1_out & ~n1703;
  assign n1705 = ~n1694 & ~n1704;
  assign n1706 = next_sys_fair<1>_out  & ~n1705;
  assign n1707 = next_sys_fair<0>_out  & ~n1245;
  assign n1708 = ~next_sys_fair<0>_out  & ~n1273;
  assign n1709 = ~n1707 & ~n1708;
  assign n1710 = next_sys_fair<3>_out  & ~n1709;
  assign n1711 = next_sys_fair<0>_out  & ~n1384;
  assign n1712 = ~next_sys_fair<0>_out  & ~n1409;
  assign n1713 = ~n1711 & ~n1712;
  assign n1714 = ~next_sys_fair<3>_out  & ~n1713;
  assign n1715 = ~n1710 & ~n1714;
  assign n1716 = reg_controllable_hmaster1_out & ~n1715;
  assign n1717 = reg_controllable_hmaster2_out & ~n1715;
  assign n1718 = next_sys_fair<0>_out  & ~n1496;
  assign n1719 = ~n1697 & ~n1718;
  assign n1720 = next_sys_fair<3>_out  & ~n1719;
  assign n1721 = next_sys_fair<0>_out  & ~n1569;
  assign n1722 = ~next_sys_fair<0>_out  & ~n1577;
  assign n1723 = ~n1721 & ~n1722;
  assign n1724 = ~next_sys_fair<3>_out  & ~n1723;
  assign n1725 = ~n1720 & ~n1724;
  assign n1726 = ~reg_controllable_hmaster2_out & ~n1725;
  assign n1727 = ~n1717 & ~n1726;
  assign n1728 = ~reg_controllable_hmaster1_out & ~n1727;
  assign n1729 = ~n1716 & ~n1728;
  assign n1730 = ~next_sys_fair<1>_out  & ~n1729;
  assign n1731 = ~n1706 & ~n1730;
  assign n1732 = reg_controllable_hmaster0_out & ~n1731;
  assign n1733 = next_sys_fair<0>_out  & ~n1549;
  assign n1734 = ~next_sys_fair<0>_out  & ~n1515;
  assign n1735 = ~n1733 & ~n1734;
  assign n1736 = next_sys_fair<3>_out  & ~n1735;
  assign n1737 = ~n1700 & ~n1736;
  assign n1738 = ~reg_controllable_hmaster2_out & ~n1737;
  assign n1739 = ~n1695 & ~n1738;
  assign n1740 = ~reg_controllable_hmaster1_out & ~n1739;
  assign n1741 = ~n1694 & ~n1740;
  assign n1742 = next_sys_fair<1>_out  & ~n1741;
  assign n1743 = ~n1730 & ~n1742;
  assign n1744 = ~reg_controllable_hmaster0_out & ~n1743;
  assign n1745 = ~n1732 & ~n1744;
  assign n1746 = reg_controllable_hmaster3_out & ~n1745;
  assign n1747 = next_sys_fair<3>_out  & ~n1339;
  assign n1748 = ~next_sys_fair<3>_out  & ~n1348;
  assign n1749 = ~n1747 & ~n1748;
  assign n1750 = reg_controllable_hmaster2_out & ~n1749;
  assign n1751 = next_sys_fair<3>_out  & ~n1549;
  assign n1752 = ~n1700 & ~n1751;
  assign n1753 = ~reg_controllable_hmaster2_out & ~n1752;
  assign n1754 = ~n1750 & ~n1753;
  assign n1755 = reg_controllable_hmaster1_out & ~n1754;
  assign n1756 = next_sys_fair<0>_out  & ~n1603;
  assign n1757 = ~next_sys_fair<0>_out  & ~n1534;
  assign n1758 = ~n1756 & ~n1757;
  assign n1759 = ~next_sys_fair<3>_out  & ~n1758;
  assign n1760 = ~n1751 & ~n1759;
  assign n1761 = reg_controllable_hmaster2_out & ~n1760;
  assign n1762 = next_sys_fair<0>_out  & ~n1577;
  assign n1763 = ~n1757 & ~n1762;
  assign n1764 = ~next_sys_fair<3>_out  & ~n1763;
  assign n1765 = ~n1751 & ~n1764;
  assign n1766 = ~reg_controllable_hmaster2_out & ~n1765;
  assign n1767 = ~n1761 & ~n1766;
  assign n1768 = ~reg_controllable_hmaster1_out & ~n1767;
  assign n1769 = ~n1755 & ~n1768;
  assign n1770 = next_sys_fair<1>_out  & ~n1769;
  assign n1771 = next_sys_fair<0>_out  & ~n1311;
  assign n1772 = ~next_sys_fair<0>_out  & ~n1339;
  assign n1773 = ~n1771 & ~n1772;
  assign n1774 = next_sys_fair<3>_out  & ~n1773;
  assign n1775 = next_sys_fair<0>_out  & ~n1442;
  assign n1776 = ~next_sys_fair<0>_out  & ~n1462;
  assign n1777 = ~n1775 & ~n1776;
  assign n1778 = ~next_sys_fair<3>_out  & ~n1777;
  assign n1779 = ~n1774 & ~n1778;
  assign n1780 = reg_controllable_hmaster2_out & ~n1779;
  assign n1781 = next_sys_fair<0>_out  & ~n1630;
  assign n1782 = ~n1722 & ~n1781;
  assign n1783 = ~next_sys_fair<3>_out  & ~n1782;
  assign n1784 = ~n1720 & ~n1783;
  assign n1785 = ~reg_controllable_hmaster2_out & ~n1784;
  assign n1786 = ~n1780 & ~n1785;
  assign n1787 = reg_controllable_hmaster1_out & ~n1786;
  assign n1788 = ~reg_controllable_hmaster1_out & ~n1725;
  assign n1789 = ~n1787 & ~n1788;
  assign n1790 = ~next_sys_fair<1>_out  & ~n1789;
  assign n1791 = ~n1770 & ~n1790;
  assign n1792 = reg_controllable_hmaster0_out & ~n1791;
  assign n1793 = reg_controllable_hmaster1_out & ~n1752;
  assign n1794 = next_sys_fair<0>_out  & ~n1534;
  assign n1795 = ~next_sys_fair<0>_out  & ~n1603;
  assign n1796 = ~n1794 & ~n1795;
  assign n1797 = ~next_sys_fair<3>_out  & ~n1796;
  assign n1798 = ~n1751 & ~n1797;
  assign n1799 = reg_controllable_hmaster2_out & ~n1798;
  assign n1800 = ~n1722 & ~n1794;
  assign n1801 = ~next_sys_fair<3>_out  & ~n1800;
  assign n1802 = ~n1751 & ~n1801;
  assign n1803 = ~reg_controllable_hmaster2_out & ~n1802;
  assign n1804 = ~n1799 & ~n1803;
  assign n1805 = ~reg_controllable_hmaster1_out & ~n1804;
  assign n1806 = ~n1793 & ~n1805;
  assign n1807 = next_sys_fair<1>_out  & ~n1806;
  assign n1808 = ~n1718 & ~n1734;
  assign n1809 = next_sys_fair<3>_out  & ~n1808;
  assign n1810 = ~n1724 & ~n1809;
  assign n1811 = reg_controllable_hmaster2_out & ~n1810;
  assign n1812 = ~next_sys_fair<0>_out  & ~n1667;
  assign n1813 = ~n1721 & ~n1812;
  assign n1814 = ~next_sys_fair<3>_out  & ~n1813;
  assign n1815 = ~n1720 & ~n1814;
  assign n1816 = ~reg_controllable_hmaster2_out & ~n1815;
  assign n1817 = ~n1811 & ~n1816;
  assign n1818 = reg_controllable_hmaster1_out & ~n1817;
  assign n1819 = ~n1788 & ~n1818;
  assign n1820 = ~next_sys_fair<1>_out  & ~n1819;
  assign n1821 = ~n1807 & ~n1820;
  assign n1822 = ~reg_controllable_hmaster0_out & ~n1821;
  assign n1823 = ~n1792 & ~n1822;
  assign n1824 = ~reg_controllable_hmaster3_out & ~n1823;
  assign n1825 = ~n1746 & ~n1824;
  assign n1826 = ~reg_controllable_hgrant6_out & ~n1825;
  assign n1827 = ~reg_controllable_hgrant6_out & ~n1826;
  assign n1828 = ~reg_stateG10_7_out & ~n1827;
  assign n1829 = ~reg_stateG10_7_out & ~n1828;
  assign n1830 = ~reg_controllable_hgrant8_out & ~n1829;
  assign n1831 = ~reg_controllable_hgrant8_out & ~n1830;
  assign n1832 = reg_controllable_hgrant7_out & ~n1831;
  assign n1833 = next_sys_fair<0>_out  & ~n1273;
  assign n1834 = ~next_sys_fair<0>_out  & ~n1245;
  assign n1835 = ~n1833 & ~n1834;
  assign n1836 = next_sys_fair<3>_out  & ~n1835;
  assign n1837 = ~n1692 & ~n1836;
  assign n1838 = reg_controllable_hmaster1_out & ~n1837;
  assign n1839 = reg_controllable_hmaster2_out & ~n1837;
  assign n1840 = ~next_sys_fair<0>_out  & ~n1496;
  assign n1841 = ~n1696 & ~n1840;
  assign n1842 = next_sys_fair<3>_out  & ~n1841;
  assign n1843 = ~n1700 & ~n1842;
  assign n1844 = ~reg_controllable_hmaster2_out & ~n1843;
  assign n1845 = ~n1839 & ~n1844;
  assign n1846 = ~reg_controllable_hmaster1_out & ~n1845;
  assign n1847 = ~n1838 & ~n1846;
  assign n1848 = next_sys_fair<1>_out  & ~n1847;
  assign n1849 = ~n1691 & ~n1714;
  assign n1850 = reg_controllable_hmaster1_out & ~n1849;
  assign n1851 = reg_controllable_hmaster2_out & ~n1849;
  assign n1852 = ~n1724 & ~n1751;
  assign n1853 = ~reg_controllable_hmaster2_out & ~n1852;
  assign n1854 = ~n1851 & ~n1853;
  assign n1855 = ~reg_controllable_hmaster1_out & ~n1854;
  assign n1856 = ~n1850 & ~n1855;
  assign n1857 = ~next_sys_fair<1>_out  & ~n1856;
  assign n1858 = ~n1848 & ~n1857;
  assign n1859 = reg_controllable_hmaster0_out & ~n1858;
  assign n1860 = next_sys_fair<0>_out  & ~n1339;
  assign n1861 = ~next_sys_fair<0>_out  & ~n1311;
  assign n1862 = ~n1860 & ~n1861;
  assign n1863 = next_sys_fair<3>_out  & ~n1862;
  assign n1864 = ~n1748 & ~n1863;
  assign n1865 = ~reg_controllable_hmaster2_out & ~n1864;
  assign n1866 = ~n1839 & ~n1865;
  assign n1867 = ~reg_controllable_hmaster1_out & ~n1866;
  assign n1868 = ~n1838 & ~n1867;
  assign n1869 = next_sys_fair<1>_out  & ~n1868;
  assign n1870 = ~n1747 & ~n1778;
  assign n1871 = ~reg_controllable_hmaster2_out & ~n1870;
  assign n1872 = ~n1851 & ~n1871;
  assign n1873 = ~reg_controllable_hmaster1_out & ~n1872;
  assign n1874 = ~n1850 & ~n1873;
  assign n1875 = ~next_sys_fair<1>_out  & ~n1874;
  assign n1876 = ~n1869 & ~n1875;
  assign n1877 = ~reg_controllable_hmaster0_out & ~n1876;
  assign n1878 = ~n1859 & ~n1877;
  assign n1879 = reg_controllable_hmaster3_out & ~n1878;
  assign n1880 = ~n1733 & ~n1840;
  assign n1881 = next_sys_fair<3>_out  & ~n1880;
  assign n1882 = ~n1700 & ~n1881;
  assign n1883 = reg_controllable_hmaster1_out & ~n1882;
  assign n1884 = ~n1759 & ~n1881;
  assign n1885 = reg_controllable_hmaster2_out & ~n1884;
  assign n1886 = ~n1764 & ~n1881;
  assign n1887 = ~reg_controllable_hmaster2_out & ~n1886;
  assign n1888 = ~n1885 & ~n1887;
  assign n1889 = ~reg_controllable_hmaster1_out & ~n1888;
  assign n1890 = ~n1883 & ~n1889;
  assign n1891 = next_sys_fair<1>_out  & ~n1890;
  assign n1892 = ~n1699 & ~n1724;
  assign n1893 = reg_controllable_hmaster2_out & ~n1892;
  assign n1894 = ~n1751 & ~n1783;
  assign n1895 = ~reg_controllable_hmaster2_out & ~n1894;
  assign n1896 = ~n1893 & ~n1895;
  assign n1897 = reg_controllable_hmaster1_out & ~n1896;
  assign n1898 = ~reg_controllable_hmaster1_out & ~n1852;
  assign n1899 = ~n1897 & ~n1898;
  assign n1900 = ~next_sys_fair<1>_out  & ~n1899;
  assign n1901 = ~n1891 & ~n1900;
  assign n1902 = reg_controllable_hmaster0_out & ~n1901;
  assign n1903 = ~n1797 & ~n1881;
  assign n1904 = reg_controllable_hmaster2_out & ~n1903;
  assign n1905 = ~n1801 & ~n1881;
  assign n1906 = ~reg_controllable_hmaster2_out & ~n1905;
  assign n1907 = ~n1904 & ~n1906;
  assign n1908 = ~reg_controllable_hmaster1_out & ~n1907;
  assign n1909 = ~n1883 & ~n1908;
  assign n1910 = next_sys_fair<1>_out  & ~n1909;
  assign n1911 = ~n1724 & ~n1736;
  assign n1912 = reg_controllable_hmaster2_out & ~n1911;
  assign n1913 = ~n1751 & ~n1814;
  assign n1914 = ~reg_controllable_hmaster2_out & ~n1913;
  assign n1915 = ~n1912 & ~n1914;
  assign n1916 = reg_controllable_hmaster1_out & ~n1915;
  assign n1917 = ~n1898 & ~n1916;
  assign n1918 = ~next_sys_fair<1>_out  & ~n1917;
  assign n1919 = ~n1910 & ~n1918;
  assign n1920 = ~reg_controllable_hmaster0_out & ~n1919;
  assign n1921 = ~n1902 & ~n1920;
  assign n1922 = ~reg_controllable_hmaster3_out & ~n1921;
  assign n1923 = ~n1879 & ~n1922;
  assign n1924 = ~reg_stateG10_8_out & ~n1923;
  assign n1925 = ~reg_stateG10_8_out & ~n1924;
  assign n1926 = ~reg_controllable_hgrant6_out & ~n1925;
  assign n1927 = ~reg_controllable_hgrant6_out & ~n1926;
  assign n1928 = reg_controllable_hgrant8_out & ~n1927;
  assign n1929 = ~reg_stateG10_6_out & ~n1705;
  assign n1930 = ~reg_stateG10_6_out & ~n1929;
  assign n1931 = next_sys_fair<1>_out  & ~n1930;
  assign n1932 = ~n1714 & ~n1836;
  assign n1933 = reg_controllable_hmaster1_out & ~n1932;
  assign n1934 = reg_controllable_hmaster2_out & ~n1932;
  assign n1935 = ~n1724 & ~n1881;
  assign n1936 = ~reg_controllable_hmaster2_out & ~n1935;
  assign n1937 = ~n1934 & ~n1936;
  assign n1938 = ~reg_controllable_hmaster1_out & ~n1937;
  assign n1939 = ~n1933 & ~n1938;
  assign n1940 = ~reg_stateG10_6_out & ~n1939;
  assign n1941 = ~reg_stateG10_6_out & ~n1940;
  assign n1942 = ~next_sys_fair<1>_out  & ~n1941;
  assign n1943 = ~n1931 & ~n1942;
  assign n1944 = reg_controllable_hmaster0_out & ~n1943;
  assign n1945 = ~reg_stateG10_6_out & ~n1741;
  assign n1946 = ~reg_stateG10_6_out & ~n1945;
  assign n1947 = next_sys_fair<1>_out  & ~n1946;
  assign n1948 = ~n1942 & ~n1947;
  assign n1949 = ~reg_controllable_hmaster0_out & ~n1948;
  assign n1950 = ~n1944 & ~n1949;
  assign n1951 = reg_controllable_hmaster3_out & ~n1950;
  assign n1952 = ~n1768 & ~n1793;
  assign n1953 = ~reg_stateG10_6_out & ~n1952;
  assign n1954 = ~reg_stateG10_6_out & ~n1953;
  assign n1955 = next_sys_fair<1>_out  & ~n1954;
  assign n1956 = ~n1724 & ~n1842;
  assign n1957 = reg_controllable_hmaster2_out & ~n1956;
  assign n1958 = ~n1783 & ~n1881;
  assign n1959 = ~reg_controllable_hmaster2_out & ~n1958;
  assign n1960 = ~n1957 & ~n1959;
  assign n1961 = reg_controllable_hmaster1_out & ~n1960;
  assign n1962 = ~reg_controllable_hmaster1_out & ~n1935;
  assign n1963 = ~n1961 & ~n1962;
  assign n1964 = ~reg_stateG10_6_out & ~n1963;
  assign n1965 = ~reg_stateG10_6_out & ~n1964;
  assign n1966 = ~next_sys_fair<1>_out  & ~n1965;
  assign n1967 = ~n1955 & ~n1966;
  assign n1968 = reg_controllable_hmaster0_out & ~n1967;
  assign n1969 = ~n1755 & ~n1805;
  assign n1970 = ~reg_stateG10_6_out & ~n1969;
  assign n1971 = ~reg_stateG10_6_out & ~n1970;
  assign n1972 = next_sys_fair<1>_out  & ~n1971;
  assign n1973 = ~n1778 & ~n1863;
  assign n1974 = reg_controllable_hmaster2_out & ~n1973;
  assign n1975 = ~n1814 & ~n1881;
  assign n1976 = ~reg_controllable_hmaster2_out & ~n1975;
  assign n1977 = ~n1974 & ~n1976;
  assign n1978 = reg_controllable_hmaster1_out & ~n1977;
  assign n1979 = ~n1962 & ~n1978;
  assign n1980 = ~reg_stateG10_6_out & ~n1979;
  assign n1981 = ~reg_stateG10_6_out & ~n1980;
  assign n1982 = ~next_sys_fair<1>_out  & ~n1981;
  assign n1983 = ~n1972 & ~n1982;
  assign n1984 = ~reg_controllable_hmaster0_out & ~n1983;
  assign n1985 = ~n1968 & ~n1984;
  assign n1986 = ~reg_controllable_hmaster3_out & ~n1985;
  assign n1987 = ~n1951 & ~n1986;
  assign n1988 = reg_controllable_hgrant6_out & ~n1987;
  assign n1989 = ~reg_stateG10_5_out & ~n1271;
  assign n1990 = ~reg_stateG10_5_out & ~n1989;
  assign n1991 = reg_controllable_hgrant5_out & ~n1990;
  assign n1992 = ~reg_stateG10_4_out & ~n1269;
  assign n1993 = ~reg_stateG10_4_out & ~n1992;
  assign n1994 = reg_controllable_hgrant4_out & ~n1993;
  assign n1995 = next_env_fair_out & ~n550;
  assign n1996 = ~next_env_fair_out & ~n557;
  assign n1997 = ~n1995 & ~n1996;
  assign n1998 = ~reg_stateG2_out & ~n1997;
  assign n1999 = ~reg_stateG2_out & ~n1998;
  assign n2000 = reg_stateA1_out & ~n1999;
  assign n2001 = reg_stateA1_out & ~n2000;
  assign n2002 = ~reg_controllable_hmastlock_out & ~n2001;
  assign n2003 = ~n546 & ~n2002;
  assign n2004 = reg_controllable_locked_out & ~n2003;
  assign n2005 = reg_controllable_hmastlock_out & ~n2001;
  assign n2006 = ~n570 & ~n2005;
  assign n2007 = ~reg_controllable_locked_out & ~n2006;
  assign n2008 = ~n2004 & ~n2007;
  assign n2009 = ~reg_controllable_hgrant2_out & ~n2008;
  assign n2010 = ~reg_controllable_hgrant2_out & ~n2009;
  assign n2011 = ~reg_controllable_hgrant1_out & ~n2010;
  assign n2012 = ~reg_controllable_hgrant1_out & ~n2011;
  assign n2013 = ~reg_controllable_hgrant3_out & ~n2012;
  assign n2014 = ~reg_controllable_hgrant3_out & ~n2013;
  assign n2015 = next_sys_fair<2>_out  & ~n2014;
  assign n2016 = ~reg_stateG10_3_out & ~n1265;
  assign n2017 = ~reg_stateG10_3_out & ~n2016;
  assign n2018 = reg_controllable_hgrant3_out & ~n2017;
  assign n2019 = ~reg_stateG10_1_out & ~n1263;
  assign n2020 = ~reg_stateG10_1_out & ~n2019;
  assign n2021 = reg_controllable_hgrant1_out & ~n2020;
  assign n2022 = ~reg_stateG10_2_out & ~n1261;
  assign n2023 = ~reg_stateG10_2_out & ~n2022;
  assign n2024 = reg_controllable_hgrant2_out & ~n2023;
  assign n2025 = reg_stateG2_out & ~n1250;
  assign n2026 = ~n1998 & ~n2025;
  assign n2027 = reg_stateA1_out & ~n2026;
  assign n2028 = ~reg_stateA1_out & ~n1250;
  assign n2029 = ~n2027 & ~n2028;
  assign n2030 = ~reg_controllable_hmastlock_out & ~n2029;
  assign n2031 = ~n592 & ~n2030;
  assign n2032 = reg_controllable_locked_out & ~n2031;
  assign n2033 = reg_stateG2_out & ~n1259;
  assign n2034 = ~n1998 & ~n2033;
  assign n2035 = reg_stateA1_out & ~n2034;
  assign n2036 = ~reg_stateA1_out & ~n1259;
  assign n2037 = ~n2035 & ~n2036;
  assign n2038 = reg_controllable_hmastlock_out & ~n2037;
  assign n2039 = ~n600 & ~n2038;
  assign n2040 = ~reg_controllable_locked_out & ~n2039;
  assign n2041 = ~n2032 & ~n2040;
  assign n2042 = ~reg_controllable_hgrant2_out & ~n2041;
  assign n2043 = ~n2024 & ~n2042;
  assign n2044 = ~reg_controllable_hgrant1_out & ~n2043;
  assign n2045 = ~n2021 & ~n2044;
  assign n2046 = ~reg_controllable_hgrant3_out & ~n2045;
  assign n2047 = ~n2018 & ~n2046;
  assign n2048 = ~next_sys_fair<2>_out  & ~n2047;
  assign n2049 = ~n2015 & ~n2048;
  assign n2050 = ~reg_controllable_hgrant4_out & ~n2049;
  assign n2051 = ~n1994 & ~n2050;
  assign n2052 = ~reg_controllable_hgrant5_out & ~n2051;
  assign n2053 = ~n1991 & ~n2052;
  assign n2054 = next_sys_fair<3>_out  & ~n2053;
  assign n2055 = next_sys_fair<2>_out  & ~n1239;
  assign n2056 = ~n1268 & ~n2055;
  assign n2057 = ~reg_controllable_hgrant4_out & ~n2056;
  assign n2058 = ~reg_controllable_hgrant4_out & ~n2057;
  assign n2059 = ~reg_stateG10_5_out & ~n2058;
  assign n2060 = ~reg_stateG10_5_out & ~n2059;
  assign n2061 = reg_controllable_hgrant5_out & ~n2060;
  assign n2062 = ~reg_stateG10_4_out & ~n1267;
  assign n2063 = ~reg_stateG10_4_out & ~n2062;
  assign n2064 = reg_controllable_hgrant4_out & ~n2063;
  assign n2065 = next_sys_fair<2>_out  & ~n2047;
  assign n2066 = ~reg_stateG10_1_out & ~n1235;
  assign n2067 = ~reg_stateG10_1_out & ~n2066;
  assign n2068 = reg_controllable_hgrant1_out & ~n2067;
  assign n2069 = ~n2044 & ~n2068;
  assign n2070 = ~reg_controllable_hgrant3_out & ~n2069;
  assign n2071 = ~n2018 & ~n2070;
  assign n2072 = ~next_sys_fair<2>_out  & ~n2071;
  assign n2073 = ~n2065 & ~n2072;
  assign n2074 = ~reg_controllable_hgrant4_out & ~n2073;
  assign n2075 = ~n2064 & ~n2074;
  assign n2076 = ~reg_controllable_hgrant5_out & ~n2075;
  assign n2077 = ~n2061 & ~n2076;
  assign n2078 = next_sys_fair<0>_out  & ~n2077;
  assign n2079 = ~reg_stateG10_5_out & ~n1280;
  assign n2080 = ~reg_stateG10_5_out & ~n2079;
  assign n2081 = reg_controllable_hgrant5_out & ~n2080;
  assign n2082 = ~reg_stateG10_4_out & ~n2056;
  assign n2083 = ~reg_stateG10_4_out & ~n2082;
  assign n2084 = reg_controllable_hgrant4_out & ~n2083;
  assign n2085 = ~reg_controllable_hgrant4_out & ~n2047;
  assign n2086 = ~n2084 & ~n2085;
  assign n2087 = ~reg_controllable_hgrant5_out & ~n2086;
  assign n2088 = ~n2081 & ~n2087;
  assign n2089 = ~next_sys_fair<0>_out  & ~n2088;
  assign n2090 = ~n2078 & ~n2089;
  assign n2091 = ~next_sys_fair<3>_out  & ~n2090;
  assign n2092 = ~n2054 & ~n2091;
  assign n2093 = reg_controllable_hmaster1_out & ~n2092;
  assign n2094 = reg_controllable_hmaster2_out & ~n2092;
  assign n2095 = ~reg_stateG10_5_out & ~n1513;
  assign n2096 = ~reg_stateG10_5_out & ~n2095;
  assign n2097 = reg_controllable_hgrant5_out & ~n2096;
  assign n2098 = ~reg_stateG10_4_out & ~n1511;
  assign n2099 = ~reg_stateG10_4_out & ~n2098;
  assign n2100 = reg_controllable_hgrant4_out & ~n2099;
  assign n2101 = ~reg_stateG10_3_out & ~n1507;
  assign n2102 = ~reg_stateG10_3_out & ~n2101;
  assign n2103 = reg_controllable_hgrant3_out & ~n2102;
  assign n2104 = ~reg_stateG10_1_out & ~n1505;
  assign n2105 = ~reg_stateG10_1_out & ~n2104;
  assign n2106 = reg_controllable_hgrant1_out & ~n2105;
  assign n2107 = ~reg_stateG10_2_out & ~n1503;
  assign n2108 = ~reg_stateG10_2_out & ~n2107;
  assign n2109 = reg_controllable_hgrant2_out & ~n2108;
  assign n2110 = ~reg_controllable_hgrant2_out & ~n1290;
  assign n2111 = ~n2109 & ~n2110;
  assign n2112 = ~reg_controllable_hgrant1_out & ~n2111;
  assign n2113 = ~n2106 & ~n2112;
  assign n2114 = ~reg_controllable_hgrant3_out & ~n2113;
  assign n2115 = ~n2103 & ~n2114;
  assign n2116 = ~next_sys_fair<2>_out  & ~n2115;
  assign n2117 = ~next_sys_fair<2>_out  & ~n2116;
  assign n2118 = ~reg_controllable_hgrant4_out & ~n2117;
  assign n2119 = ~n2100 & ~n2118;
  assign n2120 = ~reg_controllable_hgrant5_out & ~n2119;
  assign n2121 = ~n2097 & ~n2120;
  assign n2122 = next_sys_fair<0>_out  & ~n2121;
  assign n2123 = ~reg_stateG10_5_out & ~n1547;
  assign n2124 = ~reg_stateG10_5_out & ~n2123;
  assign n2125 = reg_controllable_hgrant5_out & ~n2124;
  assign n2126 = ~reg_stateG10_4_out & ~n1545;
  assign n2127 = ~reg_stateG10_4_out & ~n2126;
  assign n2128 = reg_controllable_hgrant4_out & ~n2127;
  assign n2129 = ~reg_stateG10_3_out & ~n1528;
  assign n2130 = ~reg_stateG10_3_out & ~n2129;
  assign n2131 = reg_controllable_hgrant3_out & ~n2130;
  assign n2132 = ~reg_stateG10_1_out & ~n1526;
  assign n2133 = ~reg_stateG10_1_out & ~n2132;
  assign n2134 = reg_controllable_hgrant1_out & ~n2133;
  assign n2135 = ~reg_stateG10_2_out & ~n1524;
  assign n2136 = ~reg_stateG10_2_out & ~n2135;
  assign n2137 = reg_controllable_hgrant2_out & ~n2136;
  assign n2138 = reg_controllable_locked_out & ~n1316;
  assign n2139 = ~n1523 & ~n2138;
  assign n2140 = ~reg_controllable_hgrant2_out & ~n2139;
  assign n2141 = ~n2137 & ~n2140;
  assign n2142 = ~reg_controllable_hgrant1_out & ~n2141;
  assign n2143 = ~n2134 & ~n2142;
  assign n2144 = ~reg_controllable_hgrant3_out & ~n2143;
  assign n2145 = ~n2131 & ~n2144;
  assign n2146 = ~next_sys_fair<2>_out  & ~n2145;
  assign n2147 = ~next_sys_fair<2>_out  & ~n2146;
  assign n2148 = ~reg_controllable_hgrant4_out & ~n2147;
  assign n2149 = ~n2128 & ~n2148;
  assign n2150 = ~reg_controllable_hgrant5_out & ~n2149;
  assign n2151 = ~n2125 & ~n2150;
  assign n2152 = ~next_sys_fair<0>_out  & ~n2151;
  assign n2153 = ~n2122 & ~n2152;
  assign n2154 = next_sys_fair<3>_out  & ~n2153;
  assign n2155 = next_sys_fair<2>_out  & ~n1490;
  assign n2156 = ~n1544 & ~n2155;
  assign n2157 = ~reg_controllable_hgrant4_out & ~n2156;
  assign n2158 = ~reg_controllable_hgrant4_out & ~n2157;
  assign n2159 = ~reg_stateG10_5_out & ~n2158;
  assign n2160 = ~reg_stateG10_5_out & ~n2159;
  assign n2161 = reg_controllable_hgrant5_out & ~n2160;
  assign n2162 = ~reg_stateG10_4_out & ~n1530;
  assign n2163 = ~reg_stateG10_4_out & ~n2162;
  assign n2164 = reg_controllable_hgrant4_out & ~n2163;
  assign n2165 = next_sys_fair<2>_out  & ~n2145;
  assign n2166 = ~reg_stateG10_1_out & ~n1486;
  assign n2167 = ~reg_stateG10_1_out & ~n2166;
  assign n2168 = reg_controllable_hgrant1_out & ~n2167;
  assign n2169 = ~n2142 & ~n2168;
  assign n2170 = ~reg_controllable_hgrant3_out & ~n2169;
  assign n2171 = ~n2131 & ~n2170;
  assign n2172 = ~next_sys_fair<2>_out  & ~n2171;
  assign n2173 = ~n2165 & ~n2172;
  assign n2174 = ~reg_controllable_hgrant4_out & ~n2173;
  assign n2175 = ~n2164 & ~n2174;
  assign n2176 = ~reg_controllable_hgrant5_out & ~n2175;
  assign n2177 = ~n2161 & ~n2176;
  assign n2178 = next_sys_fair<0>_out  & ~n2177;
  assign n2179 = ~reg_stateG10_5_out & ~n1532;
  assign n2180 = ~reg_stateG10_5_out & ~n2179;
  assign n2181 = reg_controllable_hgrant5_out & ~n2180;
  assign n2182 = ~reg_stateG10_4_out & ~n2156;
  assign n2183 = ~reg_stateG10_4_out & ~n2182;
  assign n2184 = reg_controllable_hgrant4_out & ~n2183;
  assign n2185 = ~reg_controllable_hgrant4_out & ~n2145;
  assign n2186 = ~n2184 & ~n2185;
  assign n2187 = ~reg_controllable_hgrant5_out & ~n2186;
  assign n2188 = ~n2181 & ~n2187;
  assign n2189 = ~next_sys_fair<0>_out  & ~n2188;
  assign n2190 = ~n2178 & ~n2189;
  assign n2191 = ~next_sys_fair<3>_out  & ~n2190;
  assign n2192 = ~n2154 & ~n2191;
  assign n2193 = ~reg_controllable_hmaster2_out & ~n2192;
  assign n2194 = ~n2094 & ~n2193;
  assign n2195 = ~reg_controllable_hmaster1_out & ~n2194;
  assign n2196 = ~n2093 & ~n2195;
  assign n2197 = next_sys_fair<1>_out  & ~n2196;
  assign n2198 = ~reg_stateG10_5_out & ~n1382;
  assign n2199 = ~reg_stateG10_5_out & ~n2198;
  assign n2200 = reg_controllable_hgrant5_out & ~n2199;
  assign n2201 = ~reg_stateG10_4_out & ~n1380;
  assign n2202 = ~reg_stateG10_4_out & ~n2201;
  assign n2203 = reg_controllable_hgrant4_out & ~n2202;
  assign n2204 = ~reg_stateG10_3_out & ~n1237;
  assign n2205 = ~reg_stateG10_3_out & ~n2204;
  assign n2206 = reg_controllable_hgrant3_out & ~n2205;
  assign n2207 = ~n2046 & ~n2206;
  assign n2208 = next_sys_fair<2>_out  & ~n2207;
  assign n2209 = ~reg_stateG10_3_out & ~n1376;
  assign n2210 = ~reg_stateG10_3_out & ~n2209;
  assign n2211 = reg_controllable_hgrant3_out & ~n2210;
  assign n2212 = ~reg_stateG10_1_out & ~n1374;
  assign n2213 = ~reg_stateG10_1_out & ~n2212;
  assign n2214 = reg_controllable_hgrant1_out & ~n2213;
  assign n2215 = ~reg_stateG10_2_out & ~n1372;
  assign n2216 = ~reg_stateG10_2_out & ~n2215;
  assign n2217 = reg_controllable_hgrant2_out & ~n2216;
  assign n2218 = reg_stateG2_out & ~n1362;
  assign n2219 = reg_stateG3_2_out & ~n550;
  assign n2220 = ~n738 & ~n2219;
  assign n2221 = next_env_fair_out & ~n2220;
  assign n2222 = ~n1996 & ~n2221;
  assign n2223 = ~reg_stateG2_out & ~n2222;
  assign n2224 = ~n2218 & ~n2223;
  assign n2225 = reg_stateA1_out & ~n2224;
  assign n2226 = ~n1366 & ~n2225;
  assign n2227 = ~reg_controllable_hmastlock_out & ~n2226;
  assign n2228 = ~n734 & ~n2227;
  assign n2229 = reg_controllable_locked_out & ~n2228;
  assign n2230 = reg_controllable_hmastlock_out & ~n2226;
  assign n2231 = ~n750 & ~n2230;
  assign n2232 = ~reg_controllable_locked_out & ~n2231;
  assign n2233 = ~n2229 & ~n2232;
  assign n2234 = ~reg_controllable_hgrant2_out & ~n2233;
  assign n2235 = ~n2217 & ~n2234;
  assign n2236 = ~reg_controllable_hgrant1_out & ~n2235;
  assign n2237 = ~n2214 & ~n2236;
  assign n2238 = ~reg_controllable_hgrant3_out & ~n2237;
  assign n2239 = ~n2211 & ~n2238;
  assign n2240 = ~next_sys_fair<2>_out  & ~n2239;
  assign n2241 = ~n2208 & ~n2240;
  assign n2242 = ~reg_controllable_hgrant4_out & ~n2241;
  assign n2243 = ~n2203 & ~n2242;
  assign n2244 = ~reg_controllable_hgrant5_out & ~n2243;
  assign n2245 = ~n2200 & ~n2244;
  assign n2246 = next_sys_fair<0>_out  & ~n2245;
  assign n2247 = ~reg_stateG10_5_out & ~n1407;
  assign n2248 = ~reg_stateG10_5_out & ~n2247;
  assign n2249 = reg_controllable_hgrant5_out & ~n2248;
  assign n2250 = ~reg_stateG10_4_out & ~n1405;
  assign n2251 = ~reg_stateG10_4_out & ~n2250;
  assign n2252 = reg_controllable_hgrant4_out & ~n2251;
  assign n2253 = ~reg_stateG10_2_out & ~n1233;
  assign n2254 = ~reg_stateG10_2_out & ~n2253;
  assign n2255 = reg_controllable_hgrant2_out & ~n2254;
  assign n2256 = ~n2042 & ~n2255;
  assign n2257 = ~reg_controllable_hgrant1_out & ~n2256;
  assign n2258 = ~n2021 & ~n2257;
  assign n2259 = ~reg_controllable_hgrant3_out & ~n2258;
  assign n2260 = ~n2018 & ~n2259;
  assign n2261 = next_sys_fair<2>_out  & ~n2260;
  assign n2262 = ~reg_stateG10_3_out & ~n1401;
  assign n2263 = ~reg_stateG10_3_out & ~n2262;
  assign n2264 = reg_controllable_hgrant3_out & ~n2263;
  assign n2265 = ~reg_stateG10_1_out & ~n1399;
  assign n2266 = ~reg_stateG10_1_out & ~n2265;
  assign n2267 = reg_controllable_hgrant1_out & ~n2266;
  assign n2268 = ~reg_stateG10_2_out & ~n1397;
  assign n2269 = ~reg_stateG10_2_out & ~n2268;
  assign n2270 = reg_controllable_hgrant2_out & ~n2269;
  assign n2271 = next_env_fair_out & ~n737;
  assign n2272 = ~n1996 & ~n2271;
  assign n2273 = ~reg_stateG2_out & ~n2272;
  assign n2274 = ~n1388 & ~n2273;
  assign n2275 = reg_stateA1_out & ~n2274;
  assign n2276 = ~reg_stateA1_out & ~n1389;
  assign n2277 = ~n2275 & ~n2276;
  assign n2278 = ~reg_controllable_hmastlock_out & ~n2277;
  assign n2279 = ~n781 & ~n2278;
  assign n2280 = reg_controllable_locked_out & ~n2279;
  assign n2281 = reg_controllable_hmastlock_out & ~n2277;
  assign n2282 = ~n784 & ~n2281;
  assign n2283 = ~reg_controllable_locked_out & ~n2282;
  assign n2284 = ~n2280 & ~n2283;
  assign n2285 = ~reg_controllable_hgrant2_out & ~n2284;
  assign n2286 = ~n2270 & ~n2285;
  assign n2287 = ~reg_controllable_hgrant1_out & ~n2286;
  assign n2288 = ~n2267 & ~n2287;
  assign n2289 = ~reg_controllable_hgrant3_out & ~n2288;
  assign n2290 = ~n2264 & ~n2289;
  assign n2291 = ~next_sys_fair<2>_out  & ~n2290;
  assign n2292 = ~n2261 & ~n2291;
  assign n2293 = ~reg_controllable_hgrant4_out & ~n2292;
  assign n2294 = ~n2252 & ~n2293;
  assign n2295 = ~reg_controllable_hgrant5_out & ~n2294;
  assign n2296 = ~n2249 & ~n2295;
  assign n2297 = ~next_sys_fair<0>_out  & ~n2296;
  assign n2298 = ~n2246 & ~n2297;
  assign n2299 = ~next_sys_fair<3>_out  & ~n2298;
  assign n2300 = ~n2054 & ~n2299;
  assign n2301 = reg_controllable_hmaster1_out & ~n2300;
  assign n2302 = reg_controllable_hmaster2_out & ~n2300;
  assign n2303 = next_sys_fair<3>_out  & ~n2151;
  assign n2304 = ~reg_stateG10_5_out & ~n1567;
  assign n2305 = ~reg_stateG10_5_out & ~n2304;
  assign n2306 = reg_controllable_hgrant5_out & ~n2305;
  assign n2307 = ~reg_stateG10_4_out & ~n1565;
  assign n2308 = ~reg_stateG10_4_out & ~n2307;
  assign n2309 = reg_controllable_hgrant4_out & ~n2308;
  assign n2310 = ~reg_stateG10_3_out & ~n1488;
  assign n2311 = ~reg_stateG10_3_out & ~n2310;
  assign n2312 = reg_controllable_hgrant3_out & ~n2311;
  assign n2313 = ~n2144 & ~n2312;
  assign n2314 = next_sys_fair<2>_out  & ~n2313;
  assign n2315 = ~reg_stateG10_3_out & ~n1561;
  assign n2316 = ~reg_stateG10_3_out & ~n2315;
  assign n2317 = reg_controllable_hgrant3_out & ~n2316;
  assign n2318 = ~reg_stateG10_1_out & ~n1559;
  assign n2319 = ~reg_stateG10_1_out & ~n2318;
  assign n2320 = reg_controllable_hgrant1_out & ~n2319;
  assign n2321 = ~reg_stateG10_2_out & ~n1557;
  assign n2322 = ~reg_stateG10_2_out & ~n2321;
  assign n2323 = reg_controllable_hgrant2_out & ~n2322;
  assign n2324 = ~reg_controllable_hgrant2_out & ~n1421;
  assign n2325 = ~n2323 & ~n2324;
  assign n2326 = ~reg_controllable_hgrant1_out & ~n2325;
  assign n2327 = ~n2320 & ~n2326;
  assign n2328 = ~reg_controllable_hgrant3_out & ~n2327;
  assign n2329 = ~n2317 & ~n2328;
  assign n2330 = ~next_sys_fair<2>_out  & ~n2329;
  assign n2331 = ~n2314 & ~n2330;
  assign n2332 = ~reg_controllable_hgrant4_out & ~n2331;
  assign n2333 = ~n2309 & ~n2332;
  assign n2334 = ~reg_controllable_hgrant5_out & ~n2333;
  assign n2335 = ~n2306 & ~n2334;
  assign n2336 = next_sys_fair<0>_out  & ~n2335;
  assign n2337 = ~reg_stateG10_5_out & ~n1575;
  assign n2338 = ~reg_stateG10_5_out & ~n2337;
  assign n2339 = reg_controllable_hgrant5_out & ~n2338;
  assign n2340 = ~reg_stateG10_4_out & ~n1573;
  assign n2341 = ~reg_stateG10_4_out & ~n2340;
  assign n2342 = reg_controllable_hgrant4_out & ~n2341;
  assign n2343 = ~reg_stateG10_2_out & ~n1484;
  assign n2344 = ~reg_stateG10_2_out & ~n2343;
  assign n2345 = reg_controllable_hgrant2_out & ~n2344;
  assign n2346 = ~n2140 & ~n2345;
  assign n2347 = ~reg_controllable_hgrant1_out & ~n2346;
  assign n2348 = ~n2134 & ~n2347;
  assign n2349 = ~reg_controllable_hgrant3_out & ~n2348;
  assign n2350 = ~n2131 & ~n2349;
  assign n2351 = next_sys_fair<2>_out  & ~n2350;
  assign n2352 = ~n2116 & ~n2351;
  assign n2353 = ~reg_controllable_hgrant4_out & ~n2352;
  assign n2354 = ~n2342 & ~n2353;
  assign n2355 = ~reg_controllable_hgrant5_out & ~n2354;
  assign n2356 = ~n2339 & ~n2355;
  assign n2357 = ~next_sys_fair<0>_out  & ~n2356;
  assign n2358 = ~n2336 & ~n2357;
  assign n2359 = ~next_sys_fair<3>_out  & ~n2358;
  assign n2360 = ~n2303 & ~n2359;
  assign n2361 = ~reg_controllable_hmaster2_out & ~n2360;
  assign n2362 = ~n2302 & ~n2361;
  assign n2363 = ~reg_controllable_hmaster1_out & ~n2362;
  assign n2364 = ~n2301 & ~n2363;
  assign n2365 = ~next_sys_fair<1>_out  & ~n2364;
  assign n2366 = ~n2197 & ~n2365;
  assign n2367 = reg_controllable_hmaster0_out & ~n2366;
  assign n2368 = next_sys_fair<0>_out  & ~n2151;
  assign n2369 = ~next_sys_fair<0>_out  & ~n2121;
  assign n2370 = ~n2368 & ~n2369;
  assign n2371 = next_sys_fair<3>_out  & ~n2370;
  assign n2372 = ~n2191 & ~n2371;
  assign n2373 = ~reg_controllable_hmaster2_out & ~n2372;
  assign n2374 = ~n2094 & ~n2373;
  assign n2375 = ~reg_controllable_hmaster1_out & ~n2374;
  assign n2376 = ~n2093 & ~n2375;
  assign n2377 = next_sys_fair<1>_out  & ~n2376;
  assign n2378 = ~n2365 & ~n2377;
  assign n2379 = ~reg_controllable_hmaster0_out & ~n2378;
  assign n2380 = ~n2367 & ~n2379;
  assign n2381 = reg_controllable_hmaster3_out & ~n2380;
  assign n2382 = ~n2191 & ~n2303;
  assign n2383 = reg_controllable_hmaster2_out & ~n2382;
  assign n2384 = ~reg_stateG10_3_out & ~n1331;
  assign n2385 = ~reg_stateG10_3_out & ~n2384;
  assign n2386 = reg_controllable_hgrant3_out & ~n2385;
  assign n2387 = ~n2144 & ~n2386;
  assign n2388 = ~next_sys_fair<2>_out  & ~n2387;
  assign n2389 = ~next_sys_fair<2>_out  & ~n2388;
  assign n2390 = ~reg_controllable_hgrant4_out & ~n2389;
  assign n2391 = ~n2128 & ~n2390;
  assign n2392 = ~reg_controllable_hgrant5_out & ~n2391;
  assign n2393 = ~n2125 & ~n2392;
  assign n2394 = next_sys_fair<3>_out  & ~n2393;
  assign n2395 = next_sys_fair<2>_out  & ~n2387;
  assign n2396 = ~n2170 & ~n2386;
  assign n2397 = ~next_sys_fair<2>_out  & ~n2396;
  assign n2398 = ~n2395 & ~n2397;
  assign n2399 = ~reg_controllable_hgrant4_out & ~n2398;
  assign n2400 = ~n2164 & ~n2399;
  assign n2401 = ~reg_controllable_hgrant5_out & ~n2400;
  assign n2402 = ~n2161 & ~n2401;
  assign n2403 = next_sys_fair<0>_out  & ~n2402;
  assign n2404 = ~reg_controllable_hgrant4_out & ~n2387;
  assign n2405 = ~n2184 & ~n2404;
  assign n2406 = ~reg_controllable_hgrant5_out & ~n2405;
  assign n2407 = ~n2181 & ~n2406;
  assign n2408 = ~next_sys_fair<0>_out  & ~n2407;
  assign n2409 = ~n2403 & ~n2408;
  assign n2410 = ~next_sys_fair<3>_out  & ~n2409;
  assign n2411 = ~n2394 & ~n2410;
  assign n2412 = ~reg_controllable_hmaster2_out & ~n2411;
  assign n2413 = ~n2383 & ~n2412;
  assign n2414 = reg_controllable_hmaster1_out & ~n2413;
  assign n2415 = ~reg_stateG10_5_out & ~n1337;
  assign n2416 = ~reg_stateG10_5_out & ~n2415;
  assign n2417 = reg_controllable_hgrant5_out & ~n2416;
  assign n2418 = ~n2150 & ~n2417;
  assign n2419 = next_sys_fair<3>_out  & ~n2418;
  assign n2420 = next_sys_fair<2>_out  & ~n1305;
  assign n2421 = ~n1334 & ~n2420;
  assign n2422 = ~reg_controllable_hgrant4_out & ~n2421;
  assign n2423 = ~reg_controllable_hgrant4_out & ~n2422;
  assign n2424 = ~reg_stateG10_5_out & ~n2423;
  assign n2425 = ~reg_stateG10_5_out & ~n2424;
  assign n2426 = reg_controllable_hgrant5_out & ~n2425;
  assign n2427 = ~reg_stateG10_4_out & ~n1599;
  assign n2428 = ~reg_stateG10_4_out & ~n2427;
  assign n2429 = reg_controllable_hgrant4_out & ~n2428;
  assign n2430 = next_sys_fair<2>_out  & ~n2115;
  assign n2431 = ~n2172 & ~n2430;
  assign n2432 = ~reg_controllable_hgrant4_out & ~n2431;
  assign n2433 = ~n2429 & ~n2432;
  assign n2434 = ~reg_controllable_hgrant5_out & ~n2433;
  assign n2435 = ~n2426 & ~n2434;
  assign n2436 = next_sys_fair<0>_out  & ~n2435;
  assign n2437 = ~reg_stateG10_5_out & ~n1346;
  assign n2438 = ~reg_stateG10_5_out & ~n2437;
  assign n2439 = reg_controllable_hgrant5_out & ~n2438;
  assign n2440 = ~n2187 & ~n2439;
  assign n2441 = ~next_sys_fair<0>_out  & ~n2440;
  assign n2442 = ~n2436 & ~n2441;
  assign n2443 = ~next_sys_fair<3>_out  & ~n2442;
  assign n2444 = ~n2419 & ~n2443;
  assign n2445 = reg_controllable_hmaster2_out & ~n2444;
  assign n2446 = ~reg_stateG10_1_out & ~n1329;
  assign n2447 = ~reg_stateG10_1_out & ~n2446;
  assign n2448 = reg_controllable_hgrant1_out & ~n2447;
  assign n2449 = ~n2142 & ~n2448;
  assign n2450 = ~reg_controllable_hgrant3_out & ~n2449;
  assign n2451 = ~n2131 & ~n2450;
  assign n2452 = ~next_sys_fair<2>_out  & ~n2451;
  assign n2453 = ~next_sys_fair<2>_out  & ~n2452;
  assign n2454 = ~reg_controllable_hgrant4_out & ~n2453;
  assign n2455 = ~n2128 & ~n2454;
  assign n2456 = ~reg_controllable_hgrant5_out & ~n2455;
  assign n2457 = ~n2125 & ~n2456;
  assign n2458 = next_sys_fair<3>_out  & ~n2457;
  assign n2459 = ~n1510 & ~n2155;
  assign n2460 = ~reg_controllable_hgrant4_out & ~n2459;
  assign n2461 = ~reg_controllable_hgrant4_out & ~n2460;
  assign n2462 = ~reg_stateG10_5_out & ~n2461;
  assign n2463 = ~reg_stateG10_5_out & ~n2462;
  assign n2464 = reg_controllable_hgrant5_out & ~n2463;
  assign n2465 = next_sys_fair<2>_out  & ~n2451;
  assign n2466 = ~reg_stateG10_1_out & ~n1301;
  assign n2467 = ~reg_stateG10_1_out & ~n2466;
  assign n2468 = reg_controllable_hgrant1_out & ~n2467;
  assign n2469 = ~n2112 & ~n2468;
  assign n2470 = ~reg_controllable_hgrant3_out & ~n2469;
  assign n2471 = ~n2103 & ~n2470;
  assign n2472 = ~next_sys_fair<2>_out  & ~n2471;
  assign n2473 = ~n2465 & ~n2472;
  assign n2474 = ~reg_controllable_hgrant4_out & ~n2473;
  assign n2475 = ~n2342 & ~n2474;
  assign n2476 = ~reg_controllable_hgrant5_out & ~n2475;
  assign n2477 = ~n2464 & ~n2476;
  assign n2478 = next_sys_fair<0>_out  & ~n2477;
  assign n2479 = ~reg_controllable_hgrant4_out & ~n2451;
  assign n2480 = ~n2184 & ~n2479;
  assign n2481 = ~reg_controllable_hgrant5_out & ~n2480;
  assign n2482 = ~n2181 & ~n2481;
  assign n2483 = ~next_sys_fair<0>_out  & ~n2482;
  assign n2484 = ~n2478 & ~n2483;
  assign n2485 = ~next_sys_fair<3>_out  & ~n2484;
  assign n2486 = ~n2458 & ~n2485;
  assign n2487 = ~reg_controllable_hmaster2_out & ~n2486;
  assign n2488 = ~n2445 & ~n2487;
  assign n2489 = ~reg_controllable_hmaster1_out & ~n2488;
  assign n2490 = ~n2414 & ~n2489;
  assign n2491 = next_sys_fair<1>_out  & ~n2490;
  assign n2492 = ~n2154 & ~n2359;
  assign n2493 = reg_controllable_hmaster2_out & ~n2492;
  assign n2494 = ~reg_stateG10_5_out & ~n1628;
  assign n2495 = ~reg_stateG10_5_out & ~n2494;
  assign n2496 = reg_controllable_hgrant5_out & ~n2495;
  assign n2497 = ~reg_stateG10_4_out & ~n1626;
  assign n2498 = ~reg_stateG10_4_out & ~n2497;
  assign n2499 = reg_controllable_hgrant4_out & ~n2498;
  assign n2500 = ~reg_stateG10_3_out & ~n1303;
  assign n2501 = ~reg_stateG10_3_out & ~n2500;
  assign n2502 = reg_controllable_hgrant3_out & ~n2501;
  assign n2503 = ~n2114 & ~n2502;
  assign n2504 = next_sys_fair<2>_out  & ~n2503;
  assign n2505 = ~reg_stateG10_3_out & ~n1434;
  assign n2506 = ~reg_stateG10_3_out & ~n2505;
  assign n2507 = reg_controllable_hgrant3_out & ~n2506;
  assign n2508 = ~n2328 & ~n2507;
  assign n2509 = ~next_sys_fair<2>_out  & ~n2508;
  assign n2510 = ~n2504 & ~n2509;
  assign n2511 = ~reg_controllable_hgrant4_out & ~n2510;
  assign n2512 = ~n2499 & ~n2511;
  assign n2513 = ~reg_controllable_hgrant5_out & ~n2512;
  assign n2514 = ~n2496 & ~n2513;
  assign n2515 = next_sys_fair<0>_out  & ~n2514;
  assign n2516 = ~n2349 & ~n2386;
  assign n2517 = next_sys_fair<2>_out  & ~n2516;
  assign n2518 = ~reg_stateG10_3_out & ~n1454;
  assign n2519 = ~reg_stateG10_3_out & ~n2518;
  assign n2520 = reg_controllable_hgrant3_out & ~n2519;
  assign n2521 = ~n2114 & ~n2520;
  assign n2522 = ~next_sys_fair<2>_out  & ~n2521;
  assign n2523 = ~n2517 & ~n2522;
  assign n2524 = ~reg_controllable_hgrant4_out & ~n2523;
  assign n2525 = ~n2342 & ~n2524;
  assign n2526 = ~reg_controllable_hgrant5_out & ~n2525;
  assign n2527 = ~n2339 & ~n2526;
  assign n2528 = ~next_sys_fair<0>_out  & ~n2527;
  assign n2529 = ~n2515 & ~n2528;
  assign n2530 = ~next_sys_fair<3>_out  & ~n2529;
  assign n2531 = ~n2394 & ~n2530;
  assign n2532 = ~reg_controllable_hmaster2_out & ~n2531;
  assign n2533 = ~n2493 & ~n2532;
  assign n2534 = reg_controllable_hmaster1_out & ~n2533;
  assign n2535 = ~reg_stateG10_5_out & ~n1440;
  assign n2536 = ~reg_stateG10_5_out & ~n2535;
  assign n2537 = reg_controllable_hgrant5_out & ~n2536;
  assign n2538 = ~n2334 & ~n2537;
  assign n2539 = next_sys_fair<0>_out  & ~n2538;
  assign n2540 = ~reg_stateG10_5_out & ~n1460;
  assign n2541 = ~reg_stateG10_5_out & ~n2540;
  assign n2542 = reg_controllable_hgrant5_out & ~n2541;
  assign n2543 = ~n2355 & ~n2542;
  assign n2544 = ~next_sys_fair<0>_out  & ~n2543;
  assign n2545 = ~n2539 & ~n2544;
  assign n2546 = ~next_sys_fair<3>_out  & ~n2545;
  assign n2547 = ~n2419 & ~n2546;
  assign n2548 = reg_controllable_hmaster2_out & ~n2547;
  assign n2549 = ~n2312 & ~n2450;
  assign n2550 = next_sys_fair<2>_out  & ~n2549;
  assign n2551 = ~reg_stateG10_1_out & ~n1432;
  assign n2552 = ~reg_stateG10_1_out & ~n2551;
  assign n2553 = reg_controllable_hgrant1_out & ~n2552;
  assign n2554 = ~n2326 & ~n2553;
  assign n2555 = ~reg_controllable_hgrant3_out & ~n2554;
  assign n2556 = ~n2317 & ~n2555;
  assign n2557 = ~next_sys_fair<2>_out  & ~n2556;
  assign n2558 = ~n2550 & ~n2557;
  assign n2559 = ~reg_controllable_hgrant4_out & ~n2558;
  assign n2560 = ~n2309 & ~n2559;
  assign n2561 = ~reg_controllable_hgrant5_out & ~n2560;
  assign n2562 = ~n2306 & ~n2561;
  assign n2563 = next_sys_fair<0>_out  & ~n2562;
  assign n2564 = ~n2347 & ~n2448;
  assign n2565 = ~reg_controllable_hgrant3_out & ~n2564;
  assign n2566 = ~n2131 & ~n2565;
  assign n2567 = next_sys_fair<2>_out  & ~n2566;
  assign n2568 = ~reg_stateG10_1_out & ~n1452;
  assign n2569 = ~reg_stateG10_1_out & ~n2568;
  assign n2570 = reg_controllable_hgrant1_out & ~n2569;
  assign n2571 = ~n2112 & ~n2570;
  assign n2572 = ~reg_controllable_hgrant3_out & ~n2571;
  assign n2573 = ~n2103 & ~n2572;
  assign n2574 = ~next_sys_fair<2>_out  & ~n2573;
  assign n2575 = ~n2567 & ~n2574;
  assign n2576 = ~reg_controllable_hgrant4_out & ~n2575;
  assign n2577 = ~n2342 & ~n2576;
  assign n2578 = ~reg_controllable_hgrant5_out & ~n2577;
  assign n2579 = ~n2339 & ~n2578;
  assign n2580 = ~next_sys_fair<0>_out  & ~n2579;
  assign n2581 = ~n2563 & ~n2580;
  assign n2582 = ~next_sys_fair<3>_out  & ~n2581;
  assign n2583 = ~n2458 & ~n2582;
  assign n2584 = ~reg_controllable_hmaster2_out & ~n2583;
  assign n2585 = ~n2548 & ~n2584;
  assign n2586 = ~reg_controllable_hmaster1_out & ~n2585;
  assign n2587 = ~n2534 & ~n2586;
  assign n2588 = ~next_sys_fair<1>_out  & ~n2587;
  assign n2589 = ~n2491 & ~n2588;
  assign n2590 = reg_controllable_hmaster0_out & ~n2589;
  assign n2591 = ~reg_stateG10_2_out & ~n1327;
  assign n2592 = ~reg_stateG10_2_out & ~n2591;
  assign n2593 = reg_controllable_hgrant2_out & ~n2592;
  assign n2594 = ~n2140 & ~n2593;
  assign n2595 = ~reg_controllable_hgrant1_out & ~n2594;
  assign n2596 = ~n2134 & ~n2595;
  assign n2597 = ~reg_controllable_hgrant3_out & ~n2596;
  assign n2598 = ~n2131 & ~n2597;
  assign n2599 = ~next_sys_fair<2>_out  & ~n2598;
  assign n2600 = ~next_sys_fair<2>_out  & ~n2599;
  assign n2601 = ~reg_controllable_hgrant4_out & ~n2600;
  assign n2602 = ~n2128 & ~n2601;
  assign n2603 = ~reg_controllable_hgrant5_out & ~n2602;
  assign n2604 = ~n2125 & ~n2603;
  assign n2605 = next_sys_fair<3>_out  & ~n2604;
  assign n2606 = next_sys_fair<2>_out  & ~n2598;
  assign n2607 = ~n2168 & ~n2595;
  assign n2608 = ~reg_controllable_hgrant3_out & ~n2607;
  assign n2609 = ~n2131 & ~n2608;
  assign n2610 = ~next_sys_fair<2>_out  & ~n2609;
  assign n2611 = ~n2606 & ~n2610;
  assign n2612 = ~reg_controllable_hgrant4_out & ~n2611;
  assign n2613 = ~n2164 & ~n2612;
  assign n2614 = ~reg_controllable_hgrant5_out & ~n2613;
  assign n2615 = ~n2161 & ~n2614;
  assign n2616 = next_sys_fair<0>_out  & ~n2615;
  assign n2617 = ~reg_controllable_hgrant4_out & ~n2598;
  assign n2618 = ~n2184 & ~n2617;
  assign n2619 = ~reg_controllable_hgrant5_out & ~n2618;
  assign n2620 = ~n2181 & ~n2619;
  assign n2621 = ~next_sys_fair<0>_out  & ~n2620;
  assign n2622 = ~n2616 & ~n2621;
  assign n2623 = ~next_sys_fair<3>_out  & ~n2622;
  assign n2624 = ~n2605 & ~n2623;
  assign n2625 = ~reg_controllable_hmaster2_out & ~n2624;
  assign n2626 = ~n2383 & ~n2625;
  assign n2627 = reg_controllable_hmaster1_out & ~n2626;
  assign n2628 = ~reg_stateG10_4_out & ~n1335;
  assign n2629 = ~reg_stateG10_4_out & ~n2628;
  assign n2630 = reg_controllable_hgrant4_out & ~n2629;
  assign n2631 = ~n2148 & ~n2630;
  assign n2632 = ~reg_controllable_hgrant5_out & ~n2631;
  assign n2633 = ~n2125 & ~n2632;
  assign n2634 = next_sys_fair<3>_out  & ~n2633;
  assign n2635 = ~reg_stateG10_4_out & ~n1333;
  assign n2636 = ~reg_stateG10_4_out & ~n2635;
  assign n2637 = reg_controllable_hgrant4_out & ~n2636;
  assign n2638 = ~n2174 & ~n2637;
  assign n2639 = ~reg_controllable_hgrant5_out & ~n2638;
  assign n2640 = ~n2161 & ~n2639;
  assign n2641 = next_sys_fair<0>_out  & ~n2640;
  assign n2642 = ~reg_stateG10_5_out & ~n1601;
  assign n2643 = ~reg_stateG10_5_out & ~n2642;
  assign n2644 = reg_controllable_hgrant5_out & ~n2643;
  assign n2645 = ~reg_stateG10_4_out & ~n2421;
  assign n2646 = ~reg_stateG10_4_out & ~n2645;
  assign n2647 = reg_controllable_hgrant4_out & ~n2646;
  assign n2648 = ~n2146 & ~n2430;
  assign n2649 = ~reg_controllable_hgrant4_out & ~n2648;
  assign n2650 = ~n2647 & ~n2649;
  assign n2651 = ~reg_controllable_hgrant5_out & ~n2650;
  assign n2652 = ~n2644 & ~n2651;
  assign n2653 = ~next_sys_fair<0>_out  & ~n2652;
  assign n2654 = ~n2641 & ~n2653;
  assign n2655 = ~next_sys_fair<3>_out  & ~n2654;
  assign n2656 = ~n2634 & ~n2655;
  assign n2657 = reg_controllable_hmaster2_out & ~n2656;
  assign n2658 = ~reg_stateG10_4_out & ~n2459;
  assign n2659 = ~reg_stateG10_4_out & ~n2658;
  assign n2660 = reg_controllable_hgrant4_out & ~n2659;
  assign n2661 = ~n2116 & ~n2165;
  assign n2662 = ~reg_controllable_hgrant4_out & ~n2661;
  assign n2663 = ~n2660 & ~n2662;
  assign n2664 = ~reg_controllable_hgrant5_out & ~n2663;
  assign n2665 = ~n2339 & ~n2664;
  assign n2666 = ~next_sys_fair<0>_out  & ~n2665;
  assign n2667 = ~n2178 & ~n2666;
  assign n2668 = ~next_sys_fair<3>_out  & ~n2667;
  assign n2669 = ~n2303 & ~n2668;
  assign n2670 = ~reg_controllable_hmaster2_out & ~n2669;
  assign n2671 = ~n2657 & ~n2670;
  assign n2672 = ~reg_controllable_hmaster1_out & ~n2671;
  assign n2673 = ~n2627 & ~n2672;
  assign n2674 = next_sys_fair<1>_out  & ~n2673;
  assign n2675 = ~n2359 & ~n2371;
  assign n2676 = reg_controllable_hmaster2_out & ~n2675;
  assign n2677 = ~n2312 & ~n2597;
  assign n2678 = next_sys_fair<2>_out  & ~n2677;
  assign n2679 = ~reg_stateG10_2_out & ~n1430;
  assign n2680 = ~reg_stateG10_2_out & ~n2679;
  assign n2681 = reg_controllable_hgrant2_out & ~n2680;
  assign n2682 = ~n2324 & ~n2681;
  assign n2683 = ~reg_controllable_hgrant1_out & ~n2682;
  assign n2684 = ~n2320 & ~n2683;
  assign n2685 = ~reg_controllable_hgrant3_out & ~n2684;
  assign n2686 = ~n2317 & ~n2685;
  assign n2687 = ~next_sys_fair<2>_out  & ~n2686;
  assign n2688 = ~n2678 & ~n2687;
  assign n2689 = ~reg_controllable_hgrant4_out & ~n2688;
  assign n2690 = ~n2309 & ~n2689;
  assign n2691 = ~reg_controllable_hgrant5_out & ~n2690;
  assign n2692 = ~n2306 & ~n2691;
  assign n2693 = next_sys_fair<0>_out  & ~n2692;
  assign n2694 = ~reg_stateG10_5_out & ~n1665;
  assign n2695 = ~reg_stateG10_5_out & ~n2694;
  assign n2696 = reg_controllable_hgrant5_out & ~n2695;
  assign n2697 = ~reg_stateG10_4_out & ~n1509;
  assign n2698 = ~reg_stateG10_4_out & ~n2697;
  assign n2699 = reg_controllable_hgrant4_out & ~n2698;
  assign n2700 = ~reg_stateG10_2_out & ~n1299;
  assign n2701 = ~reg_stateG10_2_out & ~n2700;
  assign n2702 = reg_controllable_hgrant2_out & ~n2701;
  assign n2703 = ~n2110 & ~n2702;
  assign n2704 = ~reg_controllable_hgrant1_out & ~n2703;
  assign n2705 = ~n2106 & ~n2704;
  assign n2706 = ~reg_controllable_hgrant3_out & ~n2705;
  assign n2707 = ~n2103 & ~n2706;
  assign n2708 = next_sys_fair<2>_out  & ~n2707;
  assign n2709 = ~reg_stateG10_2_out & ~n1450;
  assign n2710 = ~reg_stateG10_2_out & ~n2709;
  assign n2711 = reg_controllable_hgrant2_out & ~n2710;
  assign n2712 = ~n2110 & ~n2711;
  assign n2713 = ~reg_controllable_hgrant1_out & ~n2712;
  assign n2714 = ~n2106 & ~n2713;
  assign n2715 = ~reg_controllable_hgrant3_out & ~n2714;
  assign n2716 = ~n2103 & ~n2715;
  assign n2717 = ~next_sys_fair<2>_out  & ~n2716;
  assign n2718 = ~n2708 & ~n2717;
  assign n2719 = ~reg_controllable_hgrant4_out & ~n2718;
  assign n2720 = ~n2699 & ~n2719;
  assign n2721 = ~reg_controllable_hgrant5_out & ~n2720;
  assign n2722 = ~n2696 & ~n2721;
  assign n2723 = ~next_sys_fair<0>_out  & ~n2722;
  assign n2724 = ~n2693 & ~n2723;
  assign n2725 = ~next_sys_fair<3>_out  & ~n2724;
  assign n2726 = ~n2605 & ~n2725;
  assign n2727 = ~reg_controllable_hmaster2_out & ~n2726;
  assign n2728 = ~n2676 & ~n2727;
  assign n2729 = reg_controllable_hmaster1_out & ~n2728;
  assign n2730 = ~reg_stateG10_4_out & ~n1438;
  assign n2731 = ~reg_stateG10_4_out & ~n2730;
  assign n2732 = reg_controllable_hgrant4_out & ~n2731;
  assign n2733 = ~n2332 & ~n2732;
  assign n2734 = ~reg_controllable_hgrant5_out & ~n2733;
  assign n2735 = ~n2306 & ~n2734;
  assign n2736 = next_sys_fair<0>_out  & ~n2735;
  assign n2737 = ~reg_stateG10_4_out & ~n1458;
  assign n2738 = ~reg_stateG10_4_out & ~n2737;
  assign n2739 = reg_controllable_hgrant4_out & ~n2738;
  assign n2740 = ~n2353 & ~n2739;
  assign n2741 = ~reg_controllable_hgrant5_out & ~n2740;
  assign n2742 = ~n2339 & ~n2741;
  assign n2743 = ~next_sys_fair<0>_out  & ~n2742;
  assign n2744 = ~n2736 & ~n2743;
  assign n2745 = ~next_sys_fair<3>_out  & ~n2744;
  assign n2746 = ~n2634 & ~n2745;
  assign n2747 = reg_controllable_hmaster2_out & ~n2746;
  assign n2748 = ~n2361 & ~n2747;
  assign n2749 = ~reg_controllable_hmaster1_out & ~n2748;
  assign n2750 = ~n2729 & ~n2749;
  assign n2751 = ~next_sys_fair<1>_out  & ~n2750;
  assign n2752 = ~n2674 & ~n2751;
  assign n2753 = ~reg_controllable_hmaster0_out & ~n2752;
  assign n2754 = ~n2590 & ~n2753;
  assign n2755 = ~reg_controllable_hmaster3_out & ~n2754;
  assign n2756 = ~n2381 & ~n2755;
  assign n2757 = ~reg_controllable_hgrant6_out & ~n2756;
  assign n2758 = ~n1988 & ~n2757;
  assign n2759 = ~reg_controllable_hgrant8_out & ~n2758;
  assign n2760 = ~n1928 & ~n2759;
  assign n2761 = ~reg_controllable_hgrant7_out & ~n2760;
  assign n2762 = ~n1832 & ~n2761;
  assign n2763 = ~reg_controllable_hgrant9_out & ~n2762;
  assign n2764 = ~n1690 & ~n2763;
  assign n2765 = reg_controllable_nhgrant0_out & ~n2764;
  assign n2766 = next_sys_fair<0>_out  & ~n1282;
  assign n2767 = ~n1240 & ~n1359;
  assign n2768 = ~reg_controllable_hgrant4_out & ~n2767;
  assign n2769 = ~reg_controllable_hgrant4_out & ~n2768;
  assign n2770 = ~reg_controllable_hgrant5_out & ~n2769;
  assign n2771 = ~reg_controllable_hgrant5_out & ~n2770;
  assign n2772 = ~next_sys_fair<0>_out  & ~n2771;
  assign n2773 = ~n2766 & ~n2772;
  assign n2774 = ~next_sys_fair<3>_out  & ~n2773;
  assign n2775 = ~n1691 & ~n2774;
  assign n2776 = reg_controllable_hmaster1_out & ~n2775;
  assign n2777 = reg_controllable_hmaster2_out & ~n2775;
  assign n2778 = ~n1491 & ~n1553;
  assign n2779 = ~reg_controllable_hgrant4_out & ~n2778;
  assign n2780 = ~reg_controllable_hgrant4_out & ~n2779;
  assign n2781 = ~reg_controllable_hgrant5_out & ~n2780;
  assign n2782 = ~reg_controllable_hgrant5_out & ~n2781;
  assign n2783 = ~next_sys_fair<0>_out  & ~n2782;
  assign n2784 = ~n1794 & ~n2783;
  assign n2785 = ~next_sys_fair<3>_out  & ~n2784;
  assign n2786 = ~n1699 & ~n2785;
  assign n2787 = ~reg_controllable_hmaster2_out & ~n2786;
  assign n2788 = ~n2777 & ~n2787;
  assign n2789 = ~reg_controllable_hmaster1_out & ~n2788;
  assign n2790 = ~n2776 & ~n2789;
  assign n2791 = next_sys_fair<1>_out  & ~n2790;
  assign n2792 = ~n1857 & ~n2791;
  assign n2793 = reg_controllable_hmaster0_out & ~n2792;
  assign n2794 = ~n1736 & ~n2785;
  assign n2795 = ~reg_controllable_hmaster2_out & ~n2794;
  assign n2796 = ~n2777 & ~n2795;
  assign n2797 = ~reg_controllable_hmaster1_out & ~n2796;
  assign n2798 = ~n2776 & ~n2797;
  assign n2799 = next_sys_fair<1>_out  & ~n2798;
  assign n2800 = ~n1857 & ~n2799;
  assign n2801 = ~reg_controllable_hmaster0_out & ~n2800;
  assign n2802 = ~n2793 & ~n2801;
  assign n2803 = reg_controllable_hmaster3_out & ~n2802;
  assign n2804 = ~n1751 & ~n2785;
  assign n2805 = reg_controllable_hmaster1_out & ~n2804;
  assign n2806 = ~n1756 & ~n2783;
  assign n2807 = ~next_sys_fair<3>_out  & ~n2806;
  assign n2808 = ~n1751 & ~n2807;
  assign n2809 = reg_controllable_hmaster2_out & ~n2808;
  assign n2810 = ~n1762 & ~n2783;
  assign n2811 = ~next_sys_fair<3>_out  & ~n2810;
  assign n2812 = ~n1751 & ~n2811;
  assign n2813 = ~reg_controllable_hmaster2_out & ~n2812;
  assign n2814 = ~n2809 & ~n2813;
  assign n2815 = ~reg_controllable_hmaster1_out & ~n2814;
  assign n2816 = ~n2805 & ~n2815;
  assign n2817 = next_sys_fair<1>_out  & ~n2816;
  assign n2818 = ~n1900 & ~n2817;
  assign n2819 = reg_controllable_hmaster0_out & ~n2818;
  assign n2820 = ~n1491 & ~n1598;
  assign n2821 = ~reg_controllable_hgrant4_out & ~n2820;
  assign n2822 = ~reg_controllable_hgrant4_out & ~n2821;
  assign n2823 = ~reg_controllable_hgrant5_out & ~n2822;
  assign n2824 = ~reg_controllable_hgrant5_out & ~n2823;
  assign n2825 = ~next_sys_fair<0>_out  & ~n2824;
  assign n2826 = ~n1794 & ~n2825;
  assign n2827 = ~next_sys_fair<3>_out  & ~n2826;
  assign n2828 = ~n1751 & ~n2827;
  assign n2829 = reg_controllable_hmaster2_out & ~n2828;
  assign n2830 = next_sys_fair<0>_out  & ~n1348;
  assign n2831 = ~n1306 & ~n1419;
  assign n2832 = ~reg_controllable_hgrant4_out & ~n2831;
  assign n2833 = ~reg_controllable_hgrant4_out & ~n2832;
  assign n2834 = ~reg_controllable_hgrant5_out & ~n2833;
  assign n2835 = ~reg_controllable_hgrant5_out & ~n2834;
  assign n2836 = ~next_sys_fair<0>_out  & ~n2835;
  assign n2837 = ~n2830 & ~n2836;
  assign n2838 = ~next_sys_fair<3>_out  & ~n2837;
  assign n2839 = ~n1747 & ~n2838;
  assign n2840 = ~reg_controllable_hmaster2_out & ~n2839;
  assign n2841 = ~n2829 & ~n2840;
  assign n2842 = ~reg_controllable_hmaster1_out & ~n2841;
  assign n2843 = ~n2805 & ~n2842;
  assign n2844 = next_sys_fair<1>_out  & ~n2843;
  assign n2845 = reg_controllable_hmaster2_out & ~n1852;
  assign n2846 = ~n1871 & ~n2845;
  assign n2847 = ~reg_controllable_hmaster1_out & ~n2846;
  assign n2848 = ~n1916 & ~n2847;
  assign n2849 = ~next_sys_fair<1>_out  & ~n2848;
  assign n2850 = ~n2844 & ~n2849;
  assign n2851 = ~reg_controllable_hmaster0_out & ~n2850;
  assign n2852 = ~n2819 & ~n2851;
  assign n2853 = ~reg_controllable_hmaster3_out & ~n2852;
  assign n2854 = ~n2803 & ~n2853;
  assign n2855 = ~reg_controllable_hgrant6_out & ~n2854;
  assign n2856 = ~reg_controllable_hgrant6_out & ~n2855;
  assign n2857 = ~reg_controllable_hgrant8_out & ~n2856;
  assign n2858 = ~reg_controllable_hgrant8_out & ~n2857;
  assign n2859 = ~reg_controllable_hgrant7_out & ~n2858;
  assign n2860 = ~reg_controllable_hgrant7_out & ~n2859;
  assign n2861 = ~reg_controllable_hgrant9_out & ~n2860;
  assign n2862 = ~reg_controllable_hgrant9_out & ~n2861;
  assign n2863 = ~reg_controllable_nhgrant0_out & ~n2862;
  assign n2864 = ~n2765 & ~n2863;
  assign n2865 = ~reg_i_hready_out & ~n2864;
  assign n2866 = ~n1220 & ~n2865;
  assign n2867 = reg_controllable_ndecide_out & ~n2866;
  assign n2868 = ~reg_controllable_locked_out & ~n125;
  assign n2869 = ~reg_controllable_hgrant2_out & ~n2868;
  assign n2870 = ~reg_controllable_hgrant2_out & ~n2869;
  assign n2871 = ~reg_controllable_hgrant1_out & ~n2870;
  assign n2872 = ~reg_controllable_hgrant1_out & ~n2871;
  assign n2873 = ~reg_controllable_hgrant3_out & ~n2872;
  assign n2874 = ~reg_controllable_hgrant3_out & ~n2873;
  assign n2875 = ~next_sys_fair<2>_out  & ~n2874;
  assign n2876 = ~next_sys_fair<2>_out  & ~n2875;
  assign n2877 = ~reg_controllable_hgrant4_out & ~n2876;
  assign n2878 = ~reg_controllable_hgrant4_out & ~n2877;
  assign n2879 = ~reg_controllable_hgrant5_out & ~n2878;
  assign n2880 = ~reg_controllable_hgrant5_out & ~n2879;
  assign n2881 = reg_stateG10_9_out & ~n2880;
  assign n2882 = ~n139 & ~n2881;
  assign n2883 = next_sys_fair<0>_out  & ~n2882;
  assign n2884 = ~reg_stateG2_out & ~n176;
  assign n2885 = ~reg_stateG2_out & ~n2884;
  assign n2886 = ~reg_controllable_locked_out & ~n2885;
  assign n2887 = ~reg_controllable_locked_out & ~n2886;
  assign n2888 = ~reg_controllable_hgrant2_out & ~n2887;
  assign n2889 = ~reg_controllable_hgrant2_out & ~n2888;
  assign n2890 = ~reg_controllable_hgrant1_out & ~n2889;
  assign n2891 = ~reg_controllable_hgrant1_out & ~n2890;
  assign n2892 = ~reg_controllable_hgrant3_out & ~n2891;
  assign n2893 = ~reg_controllable_hgrant3_out & ~n2892;
  assign n2894 = ~next_sys_fair<2>_out  & ~n2893;
  assign n2895 = ~next_sys_fair<2>_out  & ~n2894;
  assign n2896 = ~reg_controllable_hgrant4_out & ~n2895;
  assign n2897 = ~reg_controllable_hgrant4_out & ~n2896;
  assign n2898 = ~reg_controllable_hgrant5_out & ~n2897;
  assign n2899 = ~reg_controllable_hgrant5_out & ~n2898;
  assign n2900 = reg_stateG10_9_out & ~n2899;
  assign n2901 = ~n156 & ~n2886;
  assign n2902 = ~reg_controllable_hgrant2_out & ~n2901;
  assign n2903 = ~reg_controllable_hgrant2_out & ~n2902;
  assign n2904 = ~reg_controllable_hgrant1_out & ~n2903;
  assign n2905 = ~reg_controllable_hgrant1_out & ~n2904;
  assign n2906 = ~reg_controllable_hgrant3_out & ~n2905;
  assign n2907 = ~reg_controllable_hgrant3_out & ~n2906;
  assign n2908 = ~next_sys_fair<2>_out  & ~n2907;
  assign n2909 = ~next_sys_fair<2>_out  & ~n2908;
  assign n2910 = ~reg_controllable_hgrant4_out & ~n2909;
  assign n2911 = ~reg_controllable_hgrant4_out & ~n2910;
  assign n2912 = ~reg_controllable_hgrant5_out & ~n2911;
  assign n2913 = ~reg_controllable_hgrant5_out & ~n2912;
  assign n2914 = ~reg_stateG10_9_out & ~n2913;
  assign n2915 = ~n2900 & ~n2914;
  assign n2916 = ~next_sys_fair<0>_out  & ~n2915;
  assign n2917 = ~n2883 & ~n2916;
  assign n2918 = next_sys_fair<3>_out  & ~n2917;
  assign n2919 = ~reg_controllable_hgrant4_out & ~n2893;
  assign n2920 = ~reg_controllable_hgrant4_out & ~n2919;
  assign n2921 = ~reg_controllable_hgrant5_out & ~n2920;
  assign n2922 = ~reg_controllable_hgrant5_out & ~n2921;
  assign n2923 = reg_stateG10_9_out & ~n2922;
  assign n2924 = ~reg_controllable_hgrant4_out & ~n2907;
  assign n2925 = ~reg_controllable_hgrant4_out & ~n2924;
  assign n2926 = ~reg_controllable_hgrant5_out & ~n2925;
  assign n2927 = ~reg_controllable_hgrant5_out & ~n2926;
  assign n2928 = ~reg_stateG10_9_out & ~n2927;
  assign n2929 = ~n2923 & ~n2928;
  assign n2930 = ~next_sys_fair<3>_out  & ~n2929;
  assign n2931 = ~n2918 & ~n2930;
  assign n2932 = reg_controllable_hmaster1_out & ~n2931;
  assign n2933 = reg_controllable_hmaster2_out & ~n2931;
  assign n2934 = reg_stateA1_out & ~n117;
  assign n2935 = ~n1291 & ~n2934;
  assign n2936 = reg_controllable_hmastlock_out & ~n2935;
  assign n2937 = reg_controllable_hmastlock_out & ~n2936;
  assign n2938 = reg_controllable_locked_out & ~n2937;
  assign n2939 = ~reg_controllable_hmastlock_out & ~n1290;
  assign n2940 = ~n222 & ~n2939;
  assign n2941 = ~reg_controllable_locked_out & ~n2940;
  assign n2942 = ~n2938 & ~n2941;
  assign n2943 = ~reg_controllable_hgrant2_out & ~n2942;
  assign n2944 = ~reg_controllable_hgrant2_out & ~n2943;
  assign n2945 = ~reg_controllable_hgrant1_out & ~n2944;
  assign n2946 = ~reg_controllable_hgrant1_out & ~n2945;
  assign n2947 = ~reg_controllable_hgrant3_out & ~n2946;
  assign n2948 = ~reg_controllable_hgrant3_out & ~n2947;
  assign n2949 = ~next_sys_fair<2>_out  & ~n2948;
  assign n2950 = ~next_sys_fair<2>_out  & ~n2949;
  assign n2951 = ~reg_controllable_hgrant4_out & ~n2950;
  assign n2952 = ~reg_controllable_hgrant4_out & ~n2951;
  assign n2953 = ~reg_controllable_hgrant5_out & ~n2952;
  assign n2954 = ~reg_controllable_hgrant5_out & ~n2953;
  assign n2955 = reg_stateG10_9_out & ~n2954;
  assign n2956 = ~n221 & ~n2941;
  assign n2957 = ~reg_controllable_hgrant2_out & ~n2956;
  assign n2958 = ~reg_controllable_hgrant2_out & ~n2957;
  assign n2959 = ~reg_controllable_hgrant1_out & ~n2958;
  assign n2960 = ~reg_controllable_hgrant1_out & ~n2959;
  assign n2961 = ~reg_controllable_hgrant3_out & ~n2960;
  assign n2962 = ~reg_controllable_hgrant3_out & ~n2961;
  assign n2963 = ~next_sys_fair<2>_out  & ~n2962;
  assign n2964 = ~next_sys_fair<2>_out  & ~n2963;
  assign n2965 = ~reg_controllable_hgrant4_out & ~n2964;
  assign n2966 = ~reg_controllable_hgrant4_out & ~n2965;
  assign n2967 = ~reg_controllable_hgrant5_out & ~n2966;
  assign n2968 = ~reg_controllable_hgrant5_out & ~n2967;
  assign n2969 = ~reg_stateG10_9_out & ~n2968;
  assign n2970 = ~n2955 & ~n2969;
  assign n2971 = next_sys_fair<0>_out  & ~n2970;
  assign n2972 = ~n1476 & ~n2033;
  assign n2973 = reg_stateA1_out & ~n2972;
  assign n2974 = ~n1478 & ~n2973;
  assign n2975 = reg_controllable_hmastlock_out & ~n2974;
  assign n2976 = reg_controllable_hmastlock_out & ~n2975;
  assign n2977 = reg_controllable_locked_out & ~n2976;
  assign n2978 = reg_controllable_hmastlock_out & ~n2885;
  assign n2979 = ~reg_controllable_hmastlock_out & ~n1477;
  assign n2980 = ~n2978 & ~n2979;
  assign n2981 = ~reg_controllable_locked_out & ~n2980;
  assign n2982 = ~n2977 & ~n2981;
  assign n2983 = ~reg_controllable_hgrant2_out & ~n2982;
  assign n2984 = ~reg_controllable_hgrant2_out & ~n2983;
  assign n2985 = ~reg_controllable_hgrant1_out & ~n2984;
  assign n2986 = ~reg_controllable_hgrant1_out & ~n2985;
  assign n2987 = ~reg_controllable_hgrant3_out & ~n2986;
  assign n2988 = ~reg_controllable_hgrant3_out & ~n2987;
  assign n2989 = ~next_sys_fair<2>_out  & ~n2988;
  assign n2990 = ~next_sys_fair<2>_out  & ~n2989;
  assign n2991 = ~reg_controllable_hgrant4_out & ~n2990;
  assign n2992 = ~reg_controllable_hgrant4_out & ~n2991;
  assign n2993 = ~reg_controllable_hgrant5_out & ~n2992;
  assign n2994 = ~reg_controllable_hgrant5_out & ~n2993;
  assign n2995 = reg_stateG10_9_out & ~n2994;
  assign n2996 = reg_stateG2_out & ~n265;
  assign n2997 = ~reg_stateG2_out & ~n263;
  assign n2998 = ~n2996 & ~n2997;
  assign n2999 = reg_stateA1_out & ~n2998;
  assign n3000 = ~reg_stateG2_out & ~n2997;
  assign n3001 = ~reg_stateA1_out & ~n3000;
  assign n3002 = ~n2999 & ~n3001;
  assign n3003 = reg_controllable_hmastlock_out & ~n3002;
  assign n3004 = ~n272 & ~n3003;
  assign n3005 = reg_controllable_locked_out & ~n3004;
  assign n3006 = ~n2981 & ~n3005;
  assign n3007 = ~reg_controllable_hgrant2_out & ~n3006;
  assign n3008 = ~reg_controllable_hgrant2_out & ~n3007;
  assign n3009 = ~reg_controllable_hgrant1_out & ~n3008;
  assign n3010 = ~reg_controllable_hgrant1_out & ~n3009;
  assign n3011 = ~reg_controllable_hgrant3_out & ~n3010;
  assign n3012 = ~reg_controllable_hgrant3_out & ~n3011;
  assign n3013 = ~next_sys_fair<2>_out  & ~n3012;
  assign n3014 = ~next_sys_fair<2>_out  & ~n3013;
  assign n3015 = ~reg_controllable_hgrant4_out & ~n3014;
  assign n3016 = ~reg_controllable_hgrant4_out & ~n3015;
  assign n3017 = ~reg_controllable_hgrant5_out & ~n3016;
  assign n3018 = ~reg_controllable_hgrant5_out & ~n3017;
  assign n3019 = ~reg_stateG10_9_out & ~n3018;
  assign n3020 = ~n2995 & ~n3019;
  assign n3021 = ~next_sys_fair<0>_out  & ~n3020;
  assign n3022 = ~n2971 & ~n3021;
  assign n3023 = next_sys_fair<3>_out  & ~n3022;
  assign n3024 = ~reg_controllable_hgrant4_out & ~n2988;
  assign n3025 = ~reg_controllable_hgrant4_out & ~n3024;
  assign n3026 = ~reg_controllable_hgrant5_out & ~n3025;
  assign n3027 = ~reg_controllable_hgrant5_out & ~n3026;
  assign n3028 = reg_stateG10_9_out & ~n3027;
  assign n3029 = ~reg_controllable_hgrant4_out & ~n3012;
  assign n3030 = ~reg_controllable_hgrant4_out & ~n3029;
  assign n3031 = ~reg_controllable_hgrant5_out & ~n3030;
  assign n3032 = ~reg_controllable_hgrant5_out & ~n3031;
  assign n3033 = ~reg_stateG10_9_out & ~n3032;
  assign n3034 = ~n3028 & ~n3033;
  assign n3035 = ~next_sys_fair<3>_out  & ~n3034;
  assign n3036 = ~n3023 & ~n3035;
  assign n3037 = ~reg_controllable_hmaster2_out & ~n3036;
  assign n3038 = ~n2933 & ~n3037;
  assign n3039 = ~reg_controllable_hmaster1_out & ~n3038;
  assign n3040 = ~n2932 & ~n3039;
  assign n3041 = reg_i_hlock9_out & ~n3040;
  assign n3042 = next_sys_fair<0>_out  & ~n2880;
  assign n3043 = ~next_sys_fair<0>_out  & ~n2899;
  assign n3044 = ~n3042 & ~n3043;
  assign n3045 = next_sys_fair<3>_out  & ~n3044;
  assign n3046 = ~next_sys_fair<3>_out  & ~n2922;
  assign n3047 = ~n3045 & ~n3046;
  assign n3048 = reg_controllable_hmaster1_out & ~n3047;
  assign n3049 = reg_controllable_hmaster2_out & ~n3047;
  assign n3050 = reg_controllable_hmastlock_out & ~n1296;
  assign n3051 = reg_controllable_locked_out & ~n3050;
  assign n3052 = ~reg_controllable_hmastlock_out & ~n2935;
  assign n3053 = ~n222 & ~n3052;
  assign n3054 = ~reg_controllable_locked_out & ~n3053;
  assign n3055 = ~n3051 & ~n3054;
  assign n3056 = ~reg_controllable_hgrant2_out & ~n3055;
  assign n3057 = ~reg_controllable_hgrant2_out & ~n3056;
  assign n3058 = ~reg_controllable_hgrant1_out & ~n3057;
  assign n3059 = ~reg_controllable_hgrant1_out & ~n3058;
  assign n3060 = ~reg_controllable_hgrant3_out & ~n3059;
  assign n3061 = ~reg_controllable_hgrant3_out & ~n3060;
  assign n3062 = ~next_sys_fair<2>_out  & ~n3061;
  assign n3063 = ~next_sys_fair<2>_out  & ~n3062;
  assign n3064 = ~reg_controllable_hgrant4_out & ~n3063;
  assign n3065 = ~reg_controllable_hgrant4_out & ~n3064;
  assign n3066 = ~reg_controllable_hgrant5_out & ~n3065;
  assign n3067 = ~reg_controllable_hgrant5_out & ~n3066;
  assign n3068 = reg_stateG10_9_out & ~n3067;
  assign n3069 = ~n225 & ~n3051;
  assign n3070 = ~reg_controllable_hgrant2_out & ~n3069;
  assign n3071 = ~reg_controllable_hgrant2_out & ~n3070;
  assign n3072 = ~reg_controllable_hgrant1_out & ~n3071;
  assign n3073 = ~reg_controllable_hgrant1_out & ~n3072;
  assign n3074 = ~reg_controllable_hgrant3_out & ~n3073;
  assign n3075 = ~reg_controllable_hgrant3_out & ~n3074;
  assign n3076 = ~next_sys_fair<2>_out  & ~n3075;
  assign n3077 = ~next_sys_fair<2>_out  & ~n3076;
  assign n3078 = ~reg_controllable_hgrant4_out & ~n3077;
  assign n3079 = ~reg_controllable_hgrant4_out & ~n3078;
  assign n3080 = ~reg_controllable_hgrant5_out & ~n3079;
  assign n3081 = ~reg_controllable_hgrant5_out & ~n3080;
  assign n3082 = ~reg_stateG10_9_out & ~n3081;
  assign n3083 = ~n3068 & ~n3082;
  assign n3084 = next_sys_fair<0>_out  & ~n3083;
  assign n3085 = reg_controllable_hmastlock_out & ~n1477;
  assign n3086 = reg_controllable_hmastlock_out & ~n3085;
  assign n3087 = reg_controllable_locked_out & ~n3086;
  assign n3088 = ~reg_controllable_hmastlock_out & ~n2974;
  assign n3089 = ~n2978 & ~n3088;
  assign n3090 = ~reg_controllable_locked_out & ~n3089;
  assign n3091 = ~n3087 & ~n3090;
  assign n3092 = ~reg_controllable_hgrant2_out & ~n3091;
  assign n3093 = ~reg_controllable_hgrant2_out & ~n3092;
  assign n3094 = ~reg_controllable_hgrant1_out & ~n3093;
  assign n3095 = ~reg_controllable_hgrant1_out & ~n3094;
  assign n3096 = ~reg_controllable_hgrant3_out & ~n3095;
  assign n3097 = ~reg_controllable_hgrant3_out & ~n3096;
  assign n3098 = ~next_sys_fair<2>_out  & ~n3097;
  assign n3099 = ~next_sys_fair<2>_out  & ~n3098;
  assign n3100 = ~reg_controllable_hgrant4_out & ~n3099;
  assign n3101 = ~reg_controllable_hgrant4_out & ~n3100;
  assign n3102 = ~reg_controllable_hgrant5_out & ~n3101;
  assign n3103 = ~reg_controllable_hgrant5_out & ~n3102;
  assign n3104 = reg_stateG10_9_out & ~n3103;
  assign n3105 = ~reg_controllable_hmastlock_out & ~n3002;
  assign n3106 = ~n2978 & ~n3105;
  assign n3107 = ~reg_controllable_locked_out & ~n3106;
  assign n3108 = ~n3087 & ~n3107;
  assign n3109 = ~reg_controllable_hgrant2_out & ~n3108;
  assign n3110 = ~reg_controllable_hgrant2_out & ~n3109;
  assign n3111 = ~reg_controllable_hgrant1_out & ~n3110;
  assign n3112 = ~reg_controllable_hgrant1_out & ~n3111;
  assign n3113 = ~reg_controllable_hgrant3_out & ~n3112;
  assign n3114 = ~reg_controllable_hgrant3_out & ~n3113;
  assign n3115 = ~next_sys_fair<2>_out  & ~n3114;
  assign n3116 = ~next_sys_fair<2>_out  & ~n3115;
  assign n3117 = ~reg_controllable_hgrant4_out & ~n3116;
  assign n3118 = ~reg_controllable_hgrant4_out & ~n3117;
  assign n3119 = ~reg_controllable_hgrant5_out & ~n3118;
  assign n3120 = ~reg_controllable_hgrant5_out & ~n3119;
  assign n3121 = ~reg_stateG10_9_out & ~n3120;
  assign n3122 = ~n3104 & ~n3121;
  assign n3123 = ~next_sys_fair<0>_out  & ~n3122;
  assign n3124 = ~n3084 & ~n3123;
  assign n3125 = next_sys_fair<3>_out  & ~n3124;
  assign n3126 = ~reg_controllable_hgrant4_out & ~n3097;
  assign n3127 = ~reg_controllable_hgrant4_out & ~n3126;
  assign n3128 = ~reg_controllable_hgrant5_out & ~n3127;
  assign n3129 = ~reg_controllable_hgrant5_out & ~n3128;
  assign n3130 = reg_stateG10_9_out & ~n3129;
  assign n3131 = ~reg_controllable_hgrant4_out & ~n3114;
  assign n3132 = ~reg_controllable_hgrant4_out & ~n3131;
  assign n3133 = ~reg_controllable_hgrant5_out & ~n3132;
  assign n3134 = ~reg_controllable_hgrant5_out & ~n3133;
  assign n3135 = ~reg_stateG10_9_out & ~n3134;
  assign n3136 = ~n3130 & ~n3135;
  assign n3137 = ~next_sys_fair<3>_out  & ~n3136;
  assign n3138 = ~n3125 & ~n3137;
  assign n3139 = ~reg_controllable_hmaster2_out & ~n3138;
  assign n3140 = ~n3049 & ~n3139;
  assign n3141 = ~reg_controllable_hmaster1_out & ~n3140;
  assign n3142 = ~n3048 & ~n3141;
  assign n3143 = ~reg_i_hlock9_out & ~n3142;
  assign n3144 = ~n3041 & ~n3143;
  assign n3145 = next_sys_fair<1>_out  & ~n3144;
  assign n3146 = next_sys_fair<3>_out  & ~n2915;
  assign n3147 = next_sys_fair<2>_out  & ~n2893;
  assign n3148 = ~n2875 & ~n3147;
  assign n3149 = ~reg_controllable_hgrant4_out & ~n3148;
  assign n3150 = ~reg_controllable_hgrant4_out & ~n3149;
  assign n3151 = ~reg_controllable_hgrant5_out & ~n3150;
  assign n3152 = ~reg_controllable_hgrant5_out & ~n3151;
  assign n3153 = reg_stateG10_9_out & ~n3152;
  assign n3154 = next_sys_fair<2>_out  & ~n2907;
  assign n3155 = ~n133 & ~n3154;
  assign n3156 = ~reg_controllable_hgrant4_out & ~n3155;
  assign n3157 = ~reg_controllable_hgrant4_out & ~n3156;
  assign n3158 = ~reg_controllable_hgrant5_out & ~n3157;
  assign n3159 = ~reg_controllable_hgrant5_out & ~n3158;
  assign n3160 = ~reg_stateG10_9_out & ~n3159;
  assign n3161 = ~n3153 & ~n3160;
  assign n3162 = ~next_sys_fair<3>_out  & ~n3161;
  assign n3163 = ~n3146 & ~n3162;
  assign n3164 = reg_controllable_hmaster1_out & ~n3163;
  assign n3165 = reg_controllable_hmaster2_out & ~n3163;
  assign n3166 = next_sys_fair<3>_out  & ~n3020;
  assign n3167 = next_sys_fair<2>_out  & ~n2988;
  assign n3168 = reg_stateA1_out & ~n1360;
  assign n3169 = ~n1422 & ~n3168;
  assign n3170 = reg_controllable_hmastlock_out & ~n3169;
  assign n3171 = reg_controllable_hmastlock_out & ~n3170;
  assign n3172 = reg_controllable_locked_out & ~n3171;
  assign n3173 = ~reg_controllable_hmastlock_out & ~n1421;
  assign n3174 = ~n222 & ~n3173;
  assign n3175 = ~reg_controllable_locked_out & ~n3174;
  assign n3176 = ~n3172 & ~n3175;
  assign n3177 = ~reg_controllable_hgrant2_out & ~n3176;
  assign n3178 = ~reg_controllable_hgrant2_out & ~n3177;
  assign n3179 = ~reg_controllable_hgrant1_out & ~n3178;
  assign n3180 = ~reg_controllable_hgrant1_out & ~n3179;
  assign n3181 = ~reg_controllable_hgrant3_out & ~n3180;
  assign n3182 = ~reg_controllable_hgrant3_out & ~n3181;
  assign n3183 = ~next_sys_fair<2>_out  & ~n3182;
  assign n3184 = ~n3167 & ~n3183;
  assign n3185 = ~reg_controllable_hgrant4_out & ~n3184;
  assign n3186 = ~reg_controllable_hgrant4_out & ~n3185;
  assign n3187 = ~reg_controllable_hgrant5_out & ~n3186;
  assign n3188 = ~reg_controllable_hgrant5_out & ~n3187;
  assign n3189 = reg_stateG10_9_out & ~n3188;
  assign n3190 = next_sys_fair<2>_out  & ~n3012;
  assign n3191 = ~n337 & ~n3175;
  assign n3192 = ~reg_controllable_hgrant2_out & ~n3191;
  assign n3193 = ~reg_controllable_hgrant2_out & ~n3192;
  assign n3194 = ~reg_controllable_hgrant1_out & ~n3193;
  assign n3195 = ~reg_controllable_hgrant1_out & ~n3194;
  assign n3196 = ~reg_controllable_hgrant3_out & ~n3195;
  assign n3197 = ~reg_controllable_hgrant3_out & ~n3196;
  assign n3198 = ~next_sys_fair<2>_out  & ~n3197;
  assign n3199 = ~n3190 & ~n3198;
  assign n3200 = ~reg_controllable_hgrant4_out & ~n3199;
  assign n3201 = ~reg_controllable_hgrant4_out & ~n3200;
  assign n3202 = ~reg_controllable_hgrant5_out & ~n3201;
  assign n3203 = ~reg_controllable_hgrant5_out & ~n3202;
  assign n3204 = ~reg_stateG10_9_out & ~n3203;
  assign n3205 = ~n3189 & ~n3204;
  assign n3206 = next_sys_fair<0>_out  & ~n3205;
  assign n3207 = ~n1291 & ~n1390;
  assign n3208 = reg_controllable_hmastlock_out & ~n3207;
  assign n3209 = reg_controllable_hmastlock_out & ~n3208;
  assign n3210 = reg_controllable_locked_out & ~n3209;
  assign n3211 = ~n2941 & ~n3210;
  assign n3212 = ~reg_controllable_hgrant2_out & ~n3211;
  assign n3213 = ~reg_controllable_hgrant2_out & ~n3212;
  assign n3214 = ~reg_controllable_hgrant1_out & ~n3213;
  assign n3215 = ~reg_controllable_hgrant1_out & ~n3214;
  assign n3216 = ~reg_controllable_hgrant3_out & ~n3215;
  assign n3217 = ~reg_controllable_hgrant3_out & ~n3216;
  assign n3218 = ~next_sys_fair<2>_out  & ~n3217;
  assign n3219 = ~n3167 & ~n3218;
  assign n3220 = ~reg_controllable_hgrant4_out & ~n3219;
  assign n3221 = ~reg_controllable_hgrant4_out & ~n3220;
  assign n3222 = ~reg_controllable_hgrant5_out & ~n3221;
  assign n3223 = ~reg_controllable_hgrant5_out & ~n3222;
  assign n3224 = reg_stateG10_9_out & ~n3223;
  assign n3225 = ~n368 & ~n2941;
  assign n3226 = ~reg_controllable_hgrant2_out & ~n3225;
  assign n3227 = ~reg_controllable_hgrant2_out & ~n3226;
  assign n3228 = ~reg_controllable_hgrant1_out & ~n3227;
  assign n3229 = ~reg_controllable_hgrant1_out & ~n3228;
  assign n3230 = ~reg_controllable_hgrant3_out & ~n3229;
  assign n3231 = ~reg_controllable_hgrant3_out & ~n3230;
  assign n3232 = ~next_sys_fair<2>_out  & ~n3231;
  assign n3233 = ~n3190 & ~n3232;
  assign n3234 = ~reg_controllable_hgrant4_out & ~n3233;
  assign n3235 = ~reg_controllable_hgrant4_out & ~n3234;
  assign n3236 = ~reg_controllable_hgrant5_out & ~n3235;
  assign n3237 = ~reg_controllable_hgrant5_out & ~n3236;
  assign n3238 = ~reg_stateG10_9_out & ~n3237;
  assign n3239 = ~n3224 & ~n3238;
  assign n3240 = ~next_sys_fair<0>_out  & ~n3239;
  assign n3241 = ~n3206 & ~n3240;
  assign n3242 = ~next_sys_fair<3>_out  & ~n3241;
  assign n3243 = ~n3166 & ~n3242;
  assign n3244 = ~reg_controllable_hmaster2_out & ~n3243;
  assign n3245 = ~n3165 & ~n3244;
  assign n3246 = ~reg_controllable_hmaster1_out & ~n3245;
  assign n3247 = ~n3164 & ~n3246;
  assign n3248 = reg_i_hlock9_out & ~n3247;
  assign n3249 = next_sys_fair<3>_out  & ~n2899;
  assign n3250 = ~next_sys_fair<3>_out  & ~n3152;
  assign n3251 = ~n3249 & ~n3250;
  assign n3252 = reg_controllable_hmaster1_out & ~n3251;
  assign n3253 = reg_controllable_hmaster2_out & ~n3251;
  assign n3254 = next_sys_fair<3>_out  & ~n3122;
  assign n3255 = next_sys_fair<2>_out  & ~n3097;
  assign n3256 = reg_controllable_hmastlock_out & ~n1427;
  assign n3257 = reg_controllable_locked_out & ~n3256;
  assign n3258 = ~reg_controllable_hmastlock_out & ~n3169;
  assign n3259 = ~n222 & ~n3258;
  assign n3260 = ~reg_controllable_locked_out & ~n3259;
  assign n3261 = ~n3257 & ~n3260;
  assign n3262 = ~reg_controllable_hgrant2_out & ~n3261;
  assign n3263 = ~reg_controllable_hgrant2_out & ~n3262;
  assign n3264 = ~reg_controllable_hgrant1_out & ~n3263;
  assign n3265 = ~reg_controllable_hgrant1_out & ~n3264;
  assign n3266 = ~reg_controllable_hgrant3_out & ~n3265;
  assign n3267 = ~reg_controllable_hgrant3_out & ~n3266;
  assign n3268 = ~next_sys_fair<2>_out  & ~n3267;
  assign n3269 = ~n3255 & ~n3268;
  assign n3270 = ~reg_controllable_hgrant4_out & ~n3269;
  assign n3271 = ~reg_controllable_hgrant4_out & ~n3270;
  assign n3272 = ~reg_controllable_hgrant5_out & ~n3271;
  assign n3273 = ~reg_controllable_hgrant5_out & ~n3272;
  assign n3274 = reg_stateG10_9_out & ~n3273;
  assign n3275 = next_sys_fair<2>_out  & ~n3114;
  assign n3276 = ~n340 & ~n3257;
  assign n3277 = ~reg_controllable_hgrant2_out & ~n3276;
  assign n3278 = ~reg_controllable_hgrant2_out & ~n3277;
  assign n3279 = ~reg_controllable_hgrant1_out & ~n3278;
  assign n3280 = ~reg_controllable_hgrant1_out & ~n3279;
  assign n3281 = ~reg_controllable_hgrant3_out & ~n3280;
  assign n3282 = ~reg_controllable_hgrant3_out & ~n3281;
  assign n3283 = ~next_sys_fair<2>_out  & ~n3282;
  assign n3284 = ~n3275 & ~n3283;
  assign n3285 = ~reg_controllable_hgrant4_out & ~n3284;
  assign n3286 = ~reg_controllable_hgrant4_out & ~n3285;
  assign n3287 = ~reg_controllable_hgrant5_out & ~n3286;
  assign n3288 = ~reg_controllable_hgrant5_out & ~n3287;
  assign n3289 = ~reg_stateG10_9_out & ~n3288;
  assign n3290 = ~n3274 & ~n3289;
  assign n3291 = next_sys_fair<0>_out  & ~n3290;
  assign n3292 = ~reg_controllable_hmastlock_out & ~n3207;
  assign n3293 = ~n222 & ~n3292;
  assign n3294 = ~reg_controllable_locked_out & ~n3293;
  assign n3295 = ~n3051 & ~n3294;
  assign n3296 = ~reg_controllable_hgrant2_out & ~n3295;
  assign n3297 = ~reg_controllable_hgrant2_out & ~n3296;
  assign n3298 = ~reg_controllable_hgrant1_out & ~n3297;
  assign n3299 = ~reg_controllable_hgrant1_out & ~n3298;
  assign n3300 = ~reg_controllable_hgrant3_out & ~n3299;
  assign n3301 = ~reg_controllable_hgrant3_out & ~n3300;
  assign n3302 = ~next_sys_fair<2>_out  & ~n3301;
  assign n3303 = ~n3255 & ~n3302;
  assign n3304 = ~reg_controllable_hgrant4_out & ~n3303;
  assign n3305 = ~reg_controllable_hgrant4_out & ~n3304;
  assign n3306 = ~reg_controllable_hgrant5_out & ~n3305;
  assign n3307 = ~reg_controllable_hgrant5_out & ~n3306;
  assign n3308 = reg_stateG10_9_out & ~n3307;
  assign n3309 = ~n371 & ~n3051;
  assign n3310 = ~reg_controllable_hgrant2_out & ~n3309;
  assign n3311 = ~reg_controllable_hgrant2_out & ~n3310;
  assign n3312 = ~reg_controllable_hgrant1_out & ~n3311;
  assign n3313 = ~reg_controllable_hgrant1_out & ~n3312;
  assign n3314 = ~reg_controllable_hgrant3_out & ~n3313;
  assign n3315 = ~reg_controllable_hgrant3_out & ~n3314;
  assign n3316 = ~next_sys_fair<2>_out  & ~n3315;
  assign n3317 = ~n3275 & ~n3316;
  assign n3318 = ~reg_controllable_hgrant4_out & ~n3317;
  assign n3319 = ~reg_controllable_hgrant4_out & ~n3318;
  assign n3320 = ~reg_controllable_hgrant5_out & ~n3319;
  assign n3321 = ~reg_controllable_hgrant5_out & ~n3320;
  assign n3322 = ~reg_stateG10_9_out & ~n3321;
  assign n3323 = ~n3308 & ~n3322;
  assign n3324 = ~next_sys_fair<0>_out  & ~n3323;
  assign n3325 = ~n3291 & ~n3324;
  assign n3326 = ~next_sys_fair<3>_out  & ~n3325;
  assign n3327 = ~n3254 & ~n3326;
  assign n3328 = ~reg_controllable_hmaster2_out & ~n3327;
  assign n3329 = ~n3253 & ~n3328;
  assign n3330 = ~reg_controllable_hmaster1_out & ~n3329;
  assign n3331 = ~n3252 & ~n3330;
  assign n3332 = ~reg_i_hlock9_out & ~n3331;
  assign n3333 = ~n3248 & ~n3332;
  assign n3334 = ~next_sys_fair<1>_out  & ~n3333;
  assign n3335 = ~n3145 & ~n3334;
  assign n3336 = reg_controllable_hmaster0_out & ~n3335;
  assign n3337 = reg_i_hlock9_out & ~n2931;
  assign n3338 = ~reg_i_hlock9_out & ~n3047;
  assign n3339 = ~n3337 & ~n3338;
  assign n3340 = next_sys_fair<1>_out  & ~n3339;
  assign n3341 = reg_i_hlock9_out & ~n3163;
  assign n3342 = ~reg_i_hlock9_out & ~n3251;
  assign n3343 = ~n3341 & ~n3342;
  assign n3344 = ~next_sys_fair<1>_out  & ~n3343;
  assign n3345 = ~n3340 & ~n3344;
  assign n3346 = ~reg_controllable_hmaster0_out & ~n3345;
  assign n3347 = ~n3336 & ~n3346;
  assign n3348 = reg_controllable_hmaster3_out & ~n3347;
  assign n3349 = ~reg_controllable_hmaster3_out & ~n3345;
  assign n3350 = ~n3348 & ~n3349;
  assign n3351 = ~reg_controllable_hgrant6_out & ~n3350;
  assign n3352 = ~reg_controllable_hgrant6_out & ~n3351;
  assign n3353 = ~reg_controllable_hgrant8_out & ~n3352;
  assign n3354 = ~reg_controllable_hgrant8_out & ~n3353;
  assign n3355 = ~reg_controllable_hgrant7_out & ~n3354;
  assign n3356 = ~reg_controllable_hgrant7_out & ~n3355;
  assign n3357 = reg_controllable_hgrant9_out & ~n3356;
  assign n3358 = ~n3046 & ~n3249;
  assign n3359 = next_sys_fair<1>_out  & ~n3358;
  assign n3360 = ~n3045 & ~n3250;
  assign n3361 = ~next_sys_fair<1>_out  & ~n3360;
  assign n3362 = ~n3359 & ~n3361;
  assign n3363 = reg_controllable_hmaster3_out & ~n3362;
  assign n3364 = next_sys_fair<3>_out  & ~n2994;
  assign n3365 = ~next_sys_fair<3>_out  & ~n3027;
  assign n3366 = ~n3364 & ~n3365;
  assign n3367 = reg_controllable_hmaster2_out & ~n3366;
  assign n3368 = ~reg_controllable_hmaster2_out & ~n3358;
  assign n3369 = ~n3367 & ~n3368;
  assign n3370 = reg_controllable_hmaster1_out & ~n3369;
  assign n3371 = ~reg_controllable_hmaster1_out & ~n3358;
  assign n3372 = ~n3370 & ~n3371;
  assign n3373 = next_sys_fair<1>_out  & ~n3372;
  assign n3374 = next_sys_fair<0>_out  & ~n2954;
  assign n3375 = ~next_sys_fair<0>_out  & ~n2994;
  assign n3376 = ~n3374 & ~n3375;
  assign n3377 = next_sys_fair<3>_out  & ~n3376;
  assign n3378 = next_sys_fair<0>_out  & ~n3188;
  assign n3379 = ~next_sys_fair<0>_out  & ~n3223;
  assign n3380 = ~n3378 & ~n3379;
  assign n3381 = ~next_sys_fair<3>_out  & ~n3380;
  assign n3382 = ~n3377 & ~n3381;
  assign n3383 = reg_controllable_hmaster2_out & ~n3382;
  assign n3384 = ~reg_controllable_hmaster2_out & ~n3360;
  assign n3385 = ~n3383 & ~n3384;
  assign n3386 = reg_controllable_hmaster1_out & ~n3385;
  assign n3387 = ~reg_controllable_hmaster1_out & ~n3360;
  assign n3388 = ~n3386 & ~n3387;
  assign n3389 = ~next_sys_fair<1>_out  & ~n3388;
  assign n3390 = ~n3373 & ~n3389;
  assign n3391 = reg_controllable_hmaster0_out & ~n3390;
  assign n3392 = ~reg_controllable_hmaster0_out & ~n3362;
  assign n3393 = ~n3391 & ~n3392;
  assign n3394 = ~reg_controllable_hmaster3_out & ~n3393;
  assign n3395 = ~n3363 & ~n3394;
  assign n3396 = ~reg_controllable_hgrant6_out & ~n3395;
  assign n3397 = ~reg_controllable_hgrant6_out & ~n3396;
  assign n3398 = reg_stateG10_7_out & ~n3397;
  assign n3399 = next_sys_fair<3>_out  & ~n2913;
  assign n3400 = ~next_sys_fair<3>_out  & ~n2927;
  assign n3401 = ~n3399 & ~n3400;
  assign n3402 = next_sys_fair<1>_out  & ~n3401;
  assign n3403 = ~next_sys_fair<0>_out  & ~n2913;
  assign n3404 = ~n417 & ~n3403;
  assign n3405 = next_sys_fair<3>_out  & ~n3404;
  assign n3406 = ~next_sys_fair<3>_out  & ~n3159;
  assign n3407 = ~n3405 & ~n3406;
  assign n3408 = ~next_sys_fair<1>_out  & ~n3407;
  assign n3409 = ~n3402 & ~n3408;
  assign n3410 = reg_controllable_hmaster3_out & ~n3409;
  assign n3411 = next_sys_fair<3>_out  & ~n3018;
  assign n3412 = ~next_sys_fair<3>_out  & ~n3032;
  assign n3413 = ~n3411 & ~n3412;
  assign n3414 = reg_controllable_hmaster2_out & ~n3413;
  assign n3415 = ~reg_controllable_hmaster2_out & ~n3401;
  assign n3416 = ~n3414 & ~n3415;
  assign n3417 = reg_controllable_hmaster1_out & ~n3416;
  assign n3418 = ~reg_controllable_hmaster1_out & ~n3401;
  assign n3419 = ~n3417 & ~n3418;
  assign n3420 = next_sys_fair<1>_out  & ~n3419;
  assign n3421 = next_sys_fair<0>_out  & ~n2968;
  assign n3422 = ~next_sys_fair<0>_out  & ~n3018;
  assign n3423 = ~n3421 & ~n3422;
  assign n3424 = next_sys_fair<3>_out  & ~n3423;
  assign n3425 = next_sys_fair<0>_out  & ~n3203;
  assign n3426 = ~next_sys_fair<0>_out  & ~n3237;
  assign n3427 = ~n3425 & ~n3426;
  assign n3428 = ~next_sys_fair<3>_out  & ~n3427;
  assign n3429 = ~n3424 & ~n3428;
  assign n3430 = reg_controllable_hmaster2_out & ~n3429;
  assign n3431 = ~reg_controllable_hmaster2_out & ~n3407;
  assign n3432 = ~n3430 & ~n3431;
  assign n3433 = reg_controllable_hmaster1_out & ~n3432;
  assign n3434 = ~reg_controllable_hmaster1_out & ~n3407;
  assign n3435 = ~n3433 & ~n3434;
  assign n3436 = ~next_sys_fair<1>_out  & ~n3435;
  assign n3437 = ~n3420 & ~n3436;
  assign n3438 = reg_controllable_hmaster0_out & ~n3437;
  assign n3439 = ~reg_controllable_hmaster0_out & ~n3409;
  assign n3440 = ~n3438 & ~n3439;
  assign n3441 = ~reg_controllable_hmaster3_out & ~n3440;
  assign n3442 = ~n3410 & ~n3441;
  assign n3443 = ~reg_controllable_hgrant6_out & ~n3442;
  assign n3444 = ~reg_controllable_hgrant6_out & ~n3443;
  assign n3445 = ~reg_stateG10_7_out & ~n3444;
  assign n3446 = ~n3398 & ~n3445;
  assign n3447 = ~reg_controllable_hgrant8_out & ~n3446;
  assign n3448 = ~reg_controllable_hgrant8_out & ~n3447;
  assign n3449 = reg_controllable_hgrant7_out & ~n3448;
  assign n3450 = next_sys_fair<0>_out  & ~n2899;
  assign n3451 = ~next_sys_fair<0>_out  & ~n2880;
  assign n3452 = ~n3450 & ~n3451;
  assign n3453 = next_sys_fair<3>_out  & ~n3452;
  assign n3454 = ~n3046 & ~n3453;
  assign n3455 = next_sys_fair<1>_out  & ~n3454;
  assign n3456 = ~next_sys_fair<1>_out  & ~n3251;
  assign n3457 = ~n3455 & ~n3456;
  assign n3458 = reg_controllable_hmaster0_out & ~n3457;
  assign n3459 = reg_controllable_hmaster1_out & ~n3454;
  assign n3460 = reg_controllable_hmaster2_out & ~n3454;
  assign n3461 = next_sys_fair<0>_out  & ~n2994;
  assign n3462 = ~next_sys_fair<0>_out  & ~n2954;
  assign n3463 = ~n3461 & ~n3462;
  assign n3464 = next_sys_fair<3>_out  & ~n3463;
  assign n3465 = ~n3365 & ~n3464;
  assign n3466 = ~reg_controllable_hmaster2_out & ~n3465;
  assign n3467 = ~n3460 & ~n3466;
  assign n3468 = ~reg_controllable_hmaster1_out & ~n3467;
  assign n3469 = ~n3459 & ~n3468;
  assign n3470 = next_sys_fair<1>_out  & ~n3469;
  assign n3471 = ~n3364 & ~n3381;
  assign n3472 = ~reg_controllable_hmaster2_out & ~n3471;
  assign n3473 = ~n3253 & ~n3472;
  assign n3474 = ~reg_controllable_hmaster1_out & ~n3473;
  assign n3475 = ~n3252 & ~n3474;
  assign n3476 = ~next_sys_fair<1>_out  & ~n3475;
  assign n3477 = ~n3470 & ~n3476;
  assign n3478 = ~reg_controllable_hmaster0_out & ~n3477;
  assign n3479 = ~n3458 & ~n3478;
  assign n3480 = reg_controllable_hmaster3_out & ~n3479;
  assign n3481 = ~reg_controllable_hmaster3_out & ~n3457;
  assign n3482 = ~n3480 & ~n3481;
  assign n3483 = reg_stateG10_8_out & ~n3482;
  assign n3484 = next_sys_fair<0>_out  & ~n2913;
  assign n3485 = ~n466 & ~n3484;
  assign n3486 = next_sys_fair<3>_out  & ~n3485;
  assign n3487 = ~n3400 & ~n3486;
  assign n3488 = next_sys_fair<1>_out  & ~n3487;
  assign n3489 = ~n3399 & ~n3406;
  assign n3490 = ~next_sys_fair<1>_out  & ~n3489;
  assign n3491 = ~n3488 & ~n3490;
  assign n3492 = reg_controllable_hmaster0_out & ~n3491;
  assign n3493 = reg_controllable_hmaster1_out & ~n3487;
  assign n3494 = reg_controllable_hmaster2_out & ~n3487;
  assign n3495 = next_sys_fair<0>_out  & ~n3018;
  assign n3496 = ~next_sys_fair<0>_out  & ~n2968;
  assign n3497 = ~n3495 & ~n3496;
  assign n3498 = next_sys_fair<3>_out  & ~n3497;
  assign n3499 = ~n3412 & ~n3498;
  assign n3500 = ~reg_controllable_hmaster2_out & ~n3499;
  assign n3501 = ~n3494 & ~n3500;
  assign n3502 = ~reg_controllable_hmaster1_out & ~n3501;
  assign n3503 = ~n3493 & ~n3502;
  assign n3504 = next_sys_fair<1>_out  & ~n3503;
  assign n3505 = reg_controllable_hmaster1_out & ~n3489;
  assign n3506 = reg_controllable_hmaster2_out & ~n3489;
  assign n3507 = ~n3411 & ~n3428;
  assign n3508 = ~reg_controllable_hmaster2_out & ~n3507;
  assign n3509 = ~n3506 & ~n3508;
  assign n3510 = ~reg_controllable_hmaster1_out & ~n3509;
  assign n3511 = ~n3505 & ~n3510;
  assign n3512 = ~next_sys_fair<1>_out  & ~n3511;
  assign n3513 = ~n3504 & ~n3512;
  assign n3514 = ~reg_controllable_hmaster0_out & ~n3513;
  assign n3515 = ~n3492 & ~n3514;
  assign n3516 = reg_controllable_hmaster3_out & ~n3515;
  assign n3517 = ~reg_controllable_hmaster3_out & ~n3491;
  assign n3518 = ~n3516 & ~n3517;
  assign n3519 = ~reg_stateG10_8_out & ~n3518;
  assign n3520 = ~n3483 & ~n3519;
  assign n3521 = ~reg_controllable_hgrant6_out & ~n3520;
  assign n3522 = ~reg_controllable_hgrant6_out & ~n3521;
  assign n3523 = reg_controllable_hgrant8_out & ~n3522;
  assign n3524 = reg_stateG10_6_out & ~n3358;
  assign n3525 = ~reg_stateG10_6_out & ~n3401;
  assign n3526 = ~n3524 & ~n3525;
  assign n3527 = reg_i_hlock6_out & ~n3526;
  assign n3528 = ~reg_i_hlock6_out & ~n3358;
  assign n3529 = ~n3527 & ~n3528;
  assign n3530 = next_sys_fair<1>_out  & ~n3529;
  assign n3531 = ~n3250 & ~n3453;
  assign n3532 = reg_stateG10_6_out & ~n3531;
  assign n3533 = ~n3406 & ~n3486;
  assign n3534 = ~reg_stateG10_6_out & ~n3533;
  assign n3535 = ~n3532 & ~n3534;
  assign n3536 = reg_i_hlock6_out & ~n3535;
  assign n3537 = ~reg_i_hlock6_out & ~n3531;
  assign n3538 = ~n3536 & ~n3537;
  assign n3539 = ~next_sys_fair<1>_out  & ~n3538;
  assign n3540 = ~n3530 & ~n3539;
  assign n3541 = reg_controllable_hmaster3_out & ~n3540;
  assign n3542 = reg_controllable_hmaster0_out & ~n3540;
  assign n3543 = reg_stateG10_6_out & ~n3372;
  assign n3544 = ~reg_stateG10_6_out & ~n3419;
  assign n3545 = ~n3543 & ~n3544;
  assign n3546 = reg_i_hlock6_out & ~n3545;
  assign n3547 = next_sys_fair<3>_out  & ~n3103;
  assign n3548 = ~next_sys_fair<3>_out  & ~n3129;
  assign n3549 = ~n3547 & ~n3548;
  assign n3550 = reg_controllable_hmaster2_out & ~n3549;
  assign n3551 = ~n3368 & ~n3550;
  assign n3552 = reg_controllable_hmaster1_out & ~n3551;
  assign n3553 = ~n3371 & ~n3552;
  assign n3554 = reg_stateG10_6_out & ~n3553;
  assign n3555 = next_sys_fair<3>_out  & ~n3120;
  assign n3556 = ~next_sys_fair<3>_out  & ~n3134;
  assign n3557 = ~n3555 & ~n3556;
  assign n3558 = reg_controllable_hmaster2_out & ~n3557;
  assign n3559 = ~n3368 & ~n3558;
  assign n3560 = reg_controllable_hmaster1_out & ~n3559;
  assign n3561 = ~n3371 & ~n3560;
  assign n3562 = ~reg_stateG10_6_out & ~n3561;
  assign n3563 = ~n3554 & ~n3562;
  assign n3564 = ~reg_i_hlock6_out & ~n3563;
  assign n3565 = ~n3546 & ~n3564;
  assign n3566 = next_sys_fair<1>_out  & ~n3565;
  assign n3567 = ~n3381 & ~n3464;
  assign n3568 = reg_controllable_hmaster2_out & ~n3567;
  assign n3569 = ~reg_controllable_hmaster2_out & ~n3531;
  assign n3570 = ~n3568 & ~n3569;
  assign n3571 = reg_controllable_hmaster1_out & ~n3570;
  assign n3572 = ~reg_controllable_hmaster1_out & ~n3531;
  assign n3573 = ~n3571 & ~n3572;
  assign n3574 = reg_stateG10_6_out & ~n3573;
  assign n3575 = ~n3428 & ~n3498;
  assign n3576 = reg_controllable_hmaster2_out & ~n3575;
  assign n3577 = ~reg_controllable_hmaster2_out & ~n3533;
  assign n3578 = ~n3576 & ~n3577;
  assign n3579 = reg_controllable_hmaster1_out & ~n3578;
  assign n3580 = ~reg_controllable_hmaster1_out & ~n3533;
  assign n3581 = ~n3579 & ~n3580;
  assign n3582 = ~reg_stateG10_6_out & ~n3581;
  assign n3583 = ~n3574 & ~n3582;
  assign n3584 = reg_i_hlock6_out & ~n3583;
  assign n3585 = next_sys_fair<0>_out  & ~n3103;
  assign n3586 = ~next_sys_fair<0>_out  & ~n3067;
  assign n3587 = ~n3585 & ~n3586;
  assign n3588 = next_sys_fair<3>_out  & ~n3587;
  assign n3589 = next_sys_fair<0>_out  & ~n3273;
  assign n3590 = ~next_sys_fair<0>_out  & ~n3307;
  assign n3591 = ~n3589 & ~n3590;
  assign n3592 = ~next_sys_fair<3>_out  & ~n3591;
  assign n3593 = ~n3588 & ~n3592;
  assign n3594 = reg_controllable_hmaster2_out & ~n3593;
  assign n3595 = ~n3569 & ~n3594;
  assign n3596 = reg_controllable_hmaster1_out & ~n3595;
  assign n3597 = ~n3572 & ~n3596;
  assign n3598 = reg_stateG10_6_out & ~n3597;
  assign n3599 = next_sys_fair<0>_out  & ~n3120;
  assign n3600 = ~next_sys_fair<0>_out  & ~n3081;
  assign n3601 = ~n3599 & ~n3600;
  assign n3602 = next_sys_fair<3>_out  & ~n3601;
  assign n3603 = next_sys_fair<0>_out  & ~n3288;
  assign n3604 = ~next_sys_fair<0>_out  & ~n3321;
  assign n3605 = ~n3603 & ~n3604;
  assign n3606 = ~next_sys_fair<3>_out  & ~n3605;
  assign n3607 = ~n3602 & ~n3606;
  assign n3608 = reg_controllable_hmaster2_out & ~n3607;
  assign n3609 = ~n3569 & ~n3608;
  assign n3610 = reg_controllable_hmaster1_out & ~n3609;
  assign n3611 = ~n3572 & ~n3610;
  assign n3612 = ~reg_stateG10_6_out & ~n3611;
  assign n3613 = ~n3598 & ~n3612;
  assign n3614 = ~reg_i_hlock6_out & ~n3613;
  assign n3615 = ~n3584 & ~n3614;
  assign n3616 = ~next_sys_fair<1>_out  & ~n3615;
  assign n3617 = ~n3566 & ~n3616;
  assign n3618 = ~reg_controllable_hmaster0_out & ~n3617;
  assign n3619 = ~n3542 & ~n3618;
  assign n3620 = ~reg_controllable_hmaster3_out & ~n3619;
  assign n3621 = ~n3541 & ~n3620;
  assign n3622 = reg_controllable_hgrant6_out & ~n3621;
  assign n3623 = reg_stateG10_5_out & ~n2897;
  assign n3624 = ~reg_stateG10_5_out & ~n2911;
  assign n3625 = ~n3623 & ~n3624;
  assign n3626 = reg_i_hlock5_out & ~n3625;
  assign n3627 = ~reg_i_hlock5_out & ~n2897;
  assign n3628 = ~n3626 & ~n3627;
  assign n3629 = reg_controllable_hgrant5_out & ~n3628;
  assign n3630 = reg_stateG10_4_out & ~n2895;
  assign n3631 = ~reg_stateG10_4_out & ~n2909;
  assign n3632 = ~n3630 & ~n3631;
  assign n3633 = reg_i_hlock4_out & ~n3632;
  assign n3634 = ~reg_i_hlock4_out & ~n2895;
  assign n3635 = ~n3633 & ~n3634;
  assign n3636 = reg_controllable_hgrant4_out & ~n3635;
  assign n3637 = reg_stateG10_3_out & ~n2891;
  assign n3638 = reg_i_hlock3_out & ~n2905;
  assign n3639 = ~reg_i_hlock3_out & ~n2891;
  assign n3640 = ~n3638 & ~n3639;
  assign n3641 = ~reg_stateG10_3_out & ~n3640;
  assign n3642 = ~n3637 & ~n3641;
  assign n3643 = reg_controllable_hgrant3_out & ~n3642;
  assign n3644 = reg_stateG10_1_out & ~n2889;
  assign n3645 = ~reg_stateG10_1_out & ~n2903;
  assign n3646 = ~n3644 & ~n3645;
  assign n3647 = reg_i_hlock1_out & ~n3646;
  assign n3648 = ~reg_i_hlock1_out & ~n2889;
  assign n3649 = ~n3647 & ~n3648;
  assign n3650 = reg_controllable_hgrant1_out & ~n3649;
  assign n3651 = reg_stateG10_2_out & ~n2887;
  assign n3652 = ~reg_stateG10_2_out & ~n2901;
  assign n3653 = ~n3651 & ~n3652;
  assign n3654 = reg_i_hlock2_out & ~n3653;
  assign n3655 = ~reg_i_hlock2_out & ~n2887;
  assign n3656 = ~n3654 & ~n3655;
  assign n3657 = reg_controllable_hgrant2_out & ~n3656;
  assign n3658 = ~reg_stateA1_out & ~n263;
  assign n3659 = ~n544 & ~n3658;
  assign n3660 = reg_controllable_hmastlock_out & ~n3659;
  assign n3661 = ~n594 & ~n3660;
  assign n3662 = reg_controllable_locked_out & ~n3661;
  assign n3663 = ~reg_stateA1_out & ~n2885;
  assign n3664 = ~n564 & ~n3663;
  assign n3665 = reg_controllable_hmastlock_out & ~n3664;
  assign n3666 = ~reg_controllable_hmastlock_out & ~n3659;
  assign n3667 = ~n3665 & ~n3666;
  assign n3668 = ~reg_controllable_locked_out & ~n3667;
  assign n3669 = ~n3662 & ~n3668;
  assign n3670 = ~reg_controllable_hgrant2_out & ~n3669;
  assign n3671 = ~n3657 & ~n3670;
  assign n3672 = ~reg_controllable_hgrant1_out & ~n3671;
  assign n3673 = ~n3650 & ~n3672;
  assign n3674 = ~reg_controllable_hgrant3_out & ~n3673;
  assign n3675 = ~n3643 & ~n3674;
  assign n3676 = ~next_sys_fair<2>_out  & ~n3675;
  assign n3677 = ~n580 & ~n3676;
  assign n3678 = ~reg_controllable_hgrant4_out & ~n3677;
  assign n3679 = ~n3636 & ~n3678;
  assign n3680 = ~reg_controllable_hgrant5_out & ~n3679;
  assign n3681 = ~n3629 & ~n3680;
  assign n3682 = next_sys_fair<3>_out  & ~n3681;
  assign n3683 = next_sys_fair<2>_out  & ~n2874;
  assign n3684 = ~n2894 & ~n3683;
  assign n3685 = ~reg_controllable_hgrant4_out & ~n3684;
  assign n3686 = ~reg_controllable_hgrant4_out & ~n3685;
  assign n3687 = reg_stateG10_5_out & ~n3686;
  assign n3688 = ~n617 & ~n2908;
  assign n3689 = ~reg_controllable_hgrant4_out & ~n3688;
  assign n3690 = ~reg_controllable_hgrant4_out & ~n3689;
  assign n3691 = ~reg_stateG10_5_out & ~n3690;
  assign n3692 = ~n3687 & ~n3691;
  assign n3693 = reg_i_hlock5_out & ~n3692;
  assign n3694 = ~reg_i_hlock5_out & ~n3686;
  assign n3695 = ~n3693 & ~n3694;
  assign n3696 = reg_controllable_hgrant5_out & ~n3695;
  assign n3697 = reg_stateG10_4_out & ~n2893;
  assign n3698 = ~reg_stateG10_4_out & ~n2907;
  assign n3699 = ~n3697 & ~n3698;
  assign n3700 = reg_i_hlock4_out & ~n3699;
  assign n3701 = ~reg_i_hlock4_out & ~n2893;
  assign n3702 = ~n3700 & ~n3701;
  assign n3703 = reg_controllable_hgrant4_out & ~n3702;
  assign n3704 = next_sys_fair<2>_out  & ~n3675;
  assign n3705 = reg_stateG10_1_out & ~n2870;
  assign n3706 = ~n628 & ~n3705;
  assign n3707 = reg_i_hlock1_out & ~n3706;
  assign n3708 = ~reg_i_hlock1_out & ~n2870;
  assign n3709 = ~n3707 & ~n3708;
  assign n3710 = reg_controllable_hgrant1_out & ~n3709;
  assign n3711 = ~n3672 & ~n3710;
  assign n3712 = ~reg_controllable_hgrant3_out & ~n3711;
  assign n3713 = ~n3643 & ~n3712;
  assign n3714 = ~next_sys_fair<2>_out  & ~n3713;
  assign n3715 = ~n3704 & ~n3714;
  assign n3716 = ~reg_controllable_hgrant4_out & ~n3715;
  assign n3717 = ~n3703 & ~n3716;
  assign n3718 = ~reg_controllable_hgrant5_out & ~n3717;
  assign n3719 = ~n3696 & ~n3718;
  assign n3720 = next_sys_fair<0>_out  & ~n3719;
  assign n3721 = reg_stateG10_5_out & ~n2920;
  assign n3722 = ~reg_stateG10_5_out & ~n2925;
  assign n3723 = ~n3721 & ~n3722;
  assign n3724 = reg_i_hlock5_out & ~n3723;
  assign n3725 = ~reg_i_hlock5_out & ~n2920;
  assign n3726 = ~n3724 & ~n3725;
  assign n3727 = reg_controllable_hgrant5_out & ~n3726;
  assign n3728 = reg_stateG10_4_out & ~n3684;
  assign n3729 = ~reg_stateG10_4_out & ~n3688;
  assign n3730 = ~n3728 & ~n3729;
  assign n3731 = reg_i_hlock4_out & ~n3730;
  assign n3732 = ~reg_i_hlock4_out & ~n3684;
  assign n3733 = ~n3731 & ~n3732;
  assign n3734 = reg_controllable_hgrant4_out & ~n3733;
  assign n3735 = ~reg_controllable_hgrant4_out & ~n3675;
  assign n3736 = ~n3734 & ~n3735;
  assign n3737 = ~reg_controllable_hgrant5_out & ~n3736;
  assign n3738 = ~n3727 & ~n3737;
  assign n3739 = ~next_sys_fair<0>_out  & ~n3738;
  assign n3740 = ~n3720 & ~n3739;
  assign n3741 = ~next_sys_fair<3>_out  & ~n3740;
  assign n3742 = ~n3682 & ~n3741;
  assign n3743 = reg_controllable_hmaster1_out & ~n3742;
  assign n3744 = reg_controllable_hmaster2_out & ~n3742;
  assign n3745 = ~reg_controllable_locked_out & ~n3664;
  assign n3746 = ~n664 & ~n3745;
  assign n3747 = ~reg_controllable_hgrant2_out & ~n3746;
  assign n3748 = ~n3657 & ~n3747;
  assign n3749 = ~reg_controllable_hgrant1_out & ~n3748;
  assign n3750 = ~n3650 & ~n3749;
  assign n3751 = ~reg_controllable_hgrant3_out & ~n3750;
  assign n3752 = ~n3643 & ~n3751;
  assign n3753 = ~next_sys_fair<2>_out  & ~n3752;
  assign n3754 = ~n663 & ~n3753;
  assign n3755 = ~reg_controllable_hgrant4_out & ~n3754;
  assign n3756 = ~n3636 & ~n3755;
  assign n3757 = ~reg_controllable_hgrant5_out & ~n3756;
  assign n3758 = ~n3629 & ~n3757;
  assign n3759 = next_sys_fair<3>_out  & ~n3758;
  assign n3760 = next_sys_fair<2>_out  & ~n3752;
  assign n3761 = ~n3710 & ~n3749;
  assign n3762 = ~reg_controllable_hgrant3_out & ~n3761;
  assign n3763 = ~n3643 & ~n3762;
  assign n3764 = ~next_sys_fair<2>_out  & ~n3763;
  assign n3765 = ~n3760 & ~n3764;
  assign n3766 = ~reg_controllable_hgrant4_out & ~n3765;
  assign n3767 = ~n3703 & ~n3766;
  assign n3768 = ~reg_controllable_hgrant5_out & ~n3767;
  assign n3769 = ~n3696 & ~n3768;
  assign n3770 = next_sys_fair<0>_out  & ~n3769;
  assign n3771 = ~reg_controllable_hgrant4_out & ~n3752;
  assign n3772 = ~n3734 & ~n3771;
  assign n3773 = ~reg_controllable_hgrant5_out & ~n3772;
  assign n3774 = ~n3727 & ~n3773;
  assign n3775 = ~next_sys_fair<0>_out  & ~n3774;
  assign n3776 = ~n3770 & ~n3775;
  assign n3777 = ~next_sys_fair<3>_out  & ~n3776;
  assign n3778 = ~n3759 & ~n3777;
  assign n3779 = ~reg_controllable_hmaster2_out & ~n3778;
  assign n3780 = ~n3744 & ~n3779;
  assign n3781 = ~reg_controllable_hmaster1_out & ~n3780;
  assign n3782 = ~n3743 & ~n3781;
  assign n3783 = next_sys_fair<1>_out  & ~n3782;
  assign n3784 = reg_stateG10_5_out & ~n3150;
  assign n3785 = ~reg_stateG10_5_out & ~n3157;
  assign n3786 = ~n3784 & ~n3785;
  assign n3787 = reg_i_hlock5_out & ~n3786;
  assign n3788 = ~reg_i_hlock5_out & ~n3150;
  assign n3789 = ~n3787 & ~n3788;
  assign n3790 = reg_controllable_hgrant5_out & ~n3789;
  assign n3791 = reg_stateG10_4_out & ~n3148;
  assign n3792 = ~reg_stateG10_4_out & ~n3155;
  assign n3793 = ~n3791 & ~n3792;
  assign n3794 = reg_i_hlock4_out & ~n3793;
  assign n3795 = ~reg_i_hlock4_out & ~n3148;
  assign n3796 = ~n3794 & ~n3795;
  assign n3797 = reg_controllable_hgrant4_out & ~n3796;
  assign n3798 = reg_stateG10_3_out & ~n2872;
  assign n3799 = reg_i_hlock3_out & ~n130;
  assign n3800 = ~reg_i_hlock3_out & ~n2872;
  assign n3801 = ~n3799 & ~n3800;
  assign n3802 = ~reg_stateG10_3_out & ~n3801;
  assign n3803 = ~n3798 & ~n3802;
  assign n3804 = reg_controllable_hgrant3_out & ~n3803;
  assign n3805 = ~n3674 & ~n3804;
  assign n3806 = next_sys_fair<2>_out  & ~n3805;
  assign n3807 = reg_stateG10_2_out & ~n2868;
  assign n3808 = ~n715 & ~n3807;
  assign n3809 = reg_i_hlock2_out & ~n3808;
  assign n3810 = ~reg_i_hlock2_out & ~n2868;
  assign n3811 = ~n3809 & ~n3810;
  assign n3812 = reg_controllable_hgrant2_out & ~n3811;
  assign n3813 = ~n754 & ~n3812;
  assign n3814 = ~reg_controllable_hgrant1_out & ~n3813;
  assign n3815 = ~n3710 & ~n3814;
  assign n3816 = ~reg_controllable_hgrant3_out & ~n3815;
  assign n3817 = ~n3804 & ~n3816;
  assign n3818 = ~next_sys_fair<2>_out  & ~n3817;
  assign n3819 = ~n3806 & ~n3818;
  assign n3820 = ~reg_controllable_hgrant4_out & ~n3819;
  assign n3821 = ~n3797 & ~n3820;
  assign n3822 = ~reg_controllable_hgrant5_out & ~n3821;
  assign n3823 = ~n3790 & ~n3822;
  assign n3824 = next_sys_fair<0>_out  & ~n3823;
  assign n3825 = ~n3670 & ~n3812;
  assign n3826 = ~reg_controllable_hgrant1_out & ~n3825;
  assign n3827 = ~n3650 & ~n3826;
  assign n3828 = ~reg_controllable_hgrant3_out & ~n3827;
  assign n3829 = ~n3643 & ~n3828;
  assign n3830 = next_sys_fair<2>_out  & ~n3829;
  assign n3831 = ~n788 & ~n3812;
  assign n3832 = ~reg_controllable_hgrant1_out & ~n3831;
  assign n3833 = ~n3710 & ~n3832;
  assign n3834 = ~reg_controllable_hgrant3_out & ~n3833;
  assign n3835 = ~n3804 & ~n3834;
  assign n3836 = ~next_sys_fair<2>_out  & ~n3835;
  assign n3837 = ~n3830 & ~n3836;
  assign n3838 = ~reg_controllable_hgrant4_out & ~n3837;
  assign n3839 = ~n3797 & ~n3838;
  assign n3840 = ~reg_controllable_hgrant5_out & ~n3839;
  assign n3841 = ~n3790 & ~n3840;
  assign n3842 = ~next_sys_fair<0>_out  & ~n3841;
  assign n3843 = ~n3824 & ~n3842;
  assign n3844 = ~next_sys_fair<3>_out  & ~n3843;
  assign n3845 = ~n3682 & ~n3844;
  assign n3846 = reg_controllable_hmaster1_out & ~n3845;
  assign n3847 = reg_controllable_hmaster2_out & ~n3845;
  assign n3848 = ~n3751 & ~n3804;
  assign n3849 = next_sys_fair<2>_out  & ~n3848;
  assign n3850 = ~n808 & ~n3812;
  assign n3851 = ~reg_controllable_hgrant1_out & ~n3850;
  assign n3852 = ~n3710 & ~n3851;
  assign n3853 = ~reg_controllable_hgrant3_out & ~n3852;
  assign n3854 = ~n3804 & ~n3853;
  assign n3855 = ~next_sys_fair<2>_out  & ~n3854;
  assign n3856 = ~n3849 & ~n3855;
  assign n3857 = ~reg_controllable_hgrant4_out & ~n3856;
  assign n3858 = ~n3797 & ~n3857;
  assign n3859 = ~reg_controllable_hgrant5_out & ~n3858;
  assign n3860 = ~n3790 & ~n3859;
  assign n3861 = next_sys_fair<0>_out  & ~n3860;
  assign n3862 = ~n3747 & ~n3812;
  assign n3863 = ~reg_controllable_hgrant1_out & ~n3862;
  assign n3864 = ~n3650 & ~n3863;
  assign n3865 = ~reg_controllable_hgrant3_out & ~n3864;
  assign n3866 = ~n3643 & ~n3865;
  assign n3867 = next_sys_fair<2>_out  & ~n3866;
  assign n3868 = ~n3855 & ~n3867;
  assign n3869 = ~reg_controllable_hgrant4_out & ~n3868;
  assign n3870 = ~n3797 & ~n3869;
  assign n3871 = ~reg_controllable_hgrant5_out & ~n3870;
  assign n3872 = ~n3790 & ~n3871;
  assign n3873 = ~next_sys_fair<0>_out  & ~n3872;
  assign n3874 = ~n3861 & ~n3873;
  assign n3875 = ~next_sys_fair<3>_out  & ~n3874;
  assign n3876 = ~n3759 & ~n3875;
  assign n3877 = ~reg_controllable_hmaster2_out & ~n3876;
  assign n3878 = ~n3847 & ~n3877;
  assign n3879 = ~reg_controllable_hmaster1_out & ~n3878;
  assign n3880 = ~n3846 & ~n3879;
  assign n3881 = ~next_sys_fair<1>_out  & ~n3880;
  assign n3882 = ~n3783 & ~n3881;
  assign n3883 = reg_controllable_hmaster3_out & ~n3882;
  assign n3884 = reg_controllable_hmaster2_out & ~n3778;
  assign n3885 = reg_i_hlock3_out & ~n2986;
  assign n3886 = ~reg_i_hlock3_out & ~n3095;
  assign n3887 = ~n3885 & ~n3886;
  assign n3888 = reg_stateG10_3_out & ~n3887;
  assign n3889 = reg_i_hlock3_out & ~n3010;
  assign n3890 = ~reg_i_hlock3_out & ~n3112;
  assign n3891 = ~n3889 & ~n3890;
  assign n3892 = ~reg_stateG10_3_out & ~n3891;
  assign n3893 = ~n3888 & ~n3892;
  assign n3894 = reg_controllable_hgrant3_out & ~n3893;
  assign n3895 = ~n3751 & ~n3894;
  assign n3896 = ~next_sys_fair<2>_out  & ~n3895;
  assign n3897 = ~n663 & ~n3896;
  assign n3898 = ~reg_controllable_hgrant4_out & ~n3897;
  assign n3899 = ~n3636 & ~n3898;
  assign n3900 = ~reg_controllable_hgrant5_out & ~n3899;
  assign n3901 = ~n3629 & ~n3900;
  assign n3902 = next_sys_fair<3>_out  & ~n3901;
  assign n3903 = next_sys_fair<2>_out  & ~n3895;
  assign n3904 = ~n3762 & ~n3894;
  assign n3905 = ~next_sys_fair<2>_out  & ~n3904;
  assign n3906 = ~n3903 & ~n3905;
  assign n3907 = ~reg_controllable_hgrant4_out & ~n3906;
  assign n3908 = ~n3703 & ~n3907;
  assign n3909 = ~reg_controllable_hgrant5_out & ~n3908;
  assign n3910 = ~n3696 & ~n3909;
  assign n3911 = next_sys_fair<0>_out  & ~n3910;
  assign n3912 = ~reg_controllable_hgrant4_out & ~n3895;
  assign n3913 = ~n3734 & ~n3912;
  assign n3914 = ~reg_controllable_hgrant5_out & ~n3913;
  assign n3915 = ~n3727 & ~n3914;
  assign n3916 = ~next_sys_fair<0>_out  & ~n3915;
  assign n3917 = ~n3911 & ~n3916;
  assign n3918 = ~next_sys_fair<3>_out  & ~n3917;
  assign n3919 = ~n3902 & ~n3918;
  assign n3920 = ~reg_controllable_hmaster2_out & ~n3919;
  assign n3921 = ~n3884 & ~n3920;
  assign n3922 = reg_controllable_hmaster1_out & ~n3921;
  assign n3923 = reg_stateG10_5_out & ~n2992;
  assign n3924 = ~reg_stateG10_5_out & ~n3016;
  assign n3925 = ~n3923 & ~n3924;
  assign n3926 = reg_i_hlock5_out & ~n3925;
  assign n3927 = reg_stateG10_5_out & ~n3101;
  assign n3928 = ~reg_stateG10_5_out & ~n3118;
  assign n3929 = ~n3927 & ~n3928;
  assign n3930 = ~reg_i_hlock5_out & ~n3929;
  assign n3931 = ~n3926 & ~n3930;
  assign n3932 = reg_controllable_hgrant5_out & ~n3931;
  assign n3933 = ~n3757 & ~n3932;
  assign n3934 = next_sys_fair<3>_out  & ~n3933;
  assign n3935 = next_sys_fair<2>_out  & ~n2948;
  assign n3936 = ~n2989 & ~n3935;
  assign n3937 = ~reg_controllable_hgrant4_out & ~n3936;
  assign n3938 = ~reg_controllable_hgrant4_out & ~n3937;
  assign n3939 = reg_stateG10_5_out & ~n3938;
  assign n3940 = next_sys_fair<2>_out  & ~n2962;
  assign n3941 = ~n3013 & ~n3940;
  assign n3942 = ~reg_controllable_hgrant4_out & ~n3941;
  assign n3943 = ~reg_controllable_hgrant4_out & ~n3942;
  assign n3944 = ~reg_stateG10_5_out & ~n3943;
  assign n3945 = ~n3939 & ~n3944;
  assign n3946 = reg_i_hlock5_out & ~n3945;
  assign n3947 = next_sys_fair<2>_out  & ~n3061;
  assign n3948 = ~n3098 & ~n3947;
  assign n3949 = ~reg_controllable_hgrant4_out & ~n3948;
  assign n3950 = ~reg_controllable_hgrant4_out & ~n3949;
  assign n3951 = reg_stateG10_5_out & ~n3950;
  assign n3952 = next_sys_fair<2>_out  & ~n3075;
  assign n3953 = ~n3115 & ~n3952;
  assign n3954 = ~reg_controllable_hgrant4_out & ~n3953;
  assign n3955 = ~reg_controllable_hgrant4_out & ~n3954;
  assign n3956 = ~reg_stateG10_5_out & ~n3955;
  assign n3957 = ~n3951 & ~n3956;
  assign n3958 = ~reg_i_hlock5_out & ~n3957;
  assign n3959 = ~n3946 & ~n3958;
  assign n3960 = reg_controllable_hgrant5_out & ~n3959;
  assign n3961 = ~n3768 & ~n3960;
  assign n3962 = next_sys_fair<0>_out  & ~n3961;
  assign n3963 = reg_stateG10_5_out & ~n3025;
  assign n3964 = ~reg_stateG10_5_out & ~n3030;
  assign n3965 = ~n3963 & ~n3964;
  assign n3966 = reg_i_hlock5_out & ~n3965;
  assign n3967 = reg_stateG10_5_out & ~n3127;
  assign n3968 = ~reg_stateG10_5_out & ~n3132;
  assign n3969 = ~n3967 & ~n3968;
  assign n3970 = ~reg_i_hlock5_out & ~n3969;
  assign n3971 = ~n3966 & ~n3970;
  assign n3972 = reg_controllable_hgrant5_out & ~n3971;
  assign n3973 = ~n3773 & ~n3972;
  assign n3974 = ~next_sys_fair<0>_out  & ~n3973;
  assign n3975 = ~n3962 & ~n3974;
  assign n3976 = ~next_sys_fair<3>_out  & ~n3975;
  assign n3977 = ~n3934 & ~n3976;
  assign n3978 = reg_controllable_hmaster2_out & ~n3977;
  assign n3979 = reg_stateG10_1_out & ~n2984;
  assign n3980 = ~reg_stateG10_1_out & ~n3008;
  assign n3981 = ~n3979 & ~n3980;
  assign n3982 = reg_i_hlock1_out & ~n3981;
  assign n3983 = reg_stateG10_1_out & ~n3093;
  assign n3984 = ~reg_stateG10_1_out & ~n3110;
  assign n3985 = ~n3983 & ~n3984;
  assign n3986 = ~reg_i_hlock1_out & ~n3985;
  assign n3987 = ~n3982 & ~n3986;
  assign n3988 = reg_controllable_hgrant1_out & ~n3987;
  assign n3989 = ~n3749 & ~n3988;
  assign n3990 = ~reg_controllable_hgrant3_out & ~n3989;
  assign n3991 = ~n3643 & ~n3990;
  assign n3992 = ~next_sys_fair<2>_out  & ~n3991;
  assign n3993 = ~n663 & ~n3992;
  assign n3994 = ~reg_controllable_hgrant4_out & ~n3993;
  assign n3995 = ~n3636 & ~n3994;
  assign n3996 = ~reg_controllable_hgrant5_out & ~n3995;
  assign n3997 = ~n3629 & ~n3996;
  assign n3998 = next_sys_fair<3>_out  & ~n3997;
  assign n3999 = next_sys_fair<2>_out  & ~n3991;
  assign n4000 = reg_stateG10_1_out & ~n2944;
  assign n4001 = ~reg_stateG10_1_out & ~n2958;
  assign n4002 = ~n4000 & ~n4001;
  assign n4003 = reg_i_hlock1_out & ~n4002;
  assign n4004 = reg_stateG10_1_out & ~n3057;
  assign n4005 = ~reg_stateG10_1_out & ~n3071;
  assign n4006 = ~n4004 & ~n4005;
  assign n4007 = ~reg_i_hlock1_out & ~n4006;
  assign n4008 = ~n4003 & ~n4007;
  assign n4009 = reg_controllable_hgrant1_out & ~n4008;
  assign n4010 = ~n3749 & ~n4009;
  assign n4011 = ~reg_controllable_hgrant3_out & ~n4010;
  assign n4012 = ~n3643 & ~n4011;
  assign n4013 = ~next_sys_fair<2>_out  & ~n4012;
  assign n4014 = ~n3999 & ~n4013;
  assign n4015 = ~reg_controllable_hgrant4_out & ~n4014;
  assign n4016 = ~n3703 & ~n4015;
  assign n4017 = ~reg_controllable_hgrant5_out & ~n4016;
  assign n4018 = ~n3696 & ~n4017;
  assign n4019 = next_sys_fair<0>_out  & ~n4018;
  assign n4020 = ~reg_controllable_hgrant4_out & ~n3991;
  assign n4021 = ~n3734 & ~n4020;
  assign n4022 = ~reg_controllable_hgrant5_out & ~n4021;
  assign n4023 = ~n3727 & ~n4022;
  assign n4024 = ~next_sys_fair<0>_out  & ~n4023;
  assign n4025 = ~n4019 & ~n4024;
  assign n4026 = ~next_sys_fair<3>_out  & ~n4025;
  assign n4027 = ~n3998 & ~n4026;
  assign n4028 = ~reg_controllable_hmaster2_out & ~n4027;
  assign n4029 = ~n3978 & ~n4028;
  assign n4030 = ~reg_controllable_hmaster1_out & ~n4029;
  assign n4031 = ~n3922 & ~n4030;
  assign n4032 = next_sys_fair<1>_out  & ~n4031;
  assign n4033 = reg_controllable_hmaster2_out & ~n3876;
  assign n4034 = reg_i_hlock3_out & ~n2946;
  assign n4035 = ~reg_i_hlock3_out & ~n3059;
  assign n4036 = ~n4034 & ~n4035;
  assign n4037 = reg_stateG10_3_out & ~n4036;
  assign n4038 = reg_i_hlock3_out & ~n2960;
  assign n4039 = ~reg_i_hlock3_out & ~n3073;
  assign n4040 = ~n4038 & ~n4039;
  assign n4041 = ~reg_stateG10_3_out & ~n4040;
  assign n4042 = ~n4037 & ~n4041;
  assign n4043 = reg_controllable_hgrant3_out & ~n4042;
  assign n4044 = ~n3751 & ~n4043;
  assign n4045 = next_sys_fair<2>_out  & ~n4044;
  assign n4046 = reg_i_hlock3_out & ~n3180;
  assign n4047 = ~reg_i_hlock3_out & ~n3265;
  assign n4048 = ~n4046 & ~n4047;
  assign n4049 = reg_stateG10_3_out & ~n4048;
  assign n4050 = reg_i_hlock3_out & ~n3195;
  assign n4051 = ~reg_i_hlock3_out & ~n3280;
  assign n4052 = ~n4050 & ~n4051;
  assign n4053 = ~reg_stateG10_3_out & ~n4052;
  assign n4054 = ~n4049 & ~n4053;
  assign n4055 = reg_controllable_hgrant3_out & ~n4054;
  assign n4056 = ~n3853 & ~n4055;
  assign n4057 = ~next_sys_fair<2>_out  & ~n4056;
  assign n4058 = ~n4045 & ~n4057;
  assign n4059 = ~reg_controllable_hgrant4_out & ~n4058;
  assign n4060 = ~n3797 & ~n4059;
  assign n4061 = ~reg_controllable_hgrant5_out & ~n4060;
  assign n4062 = ~n3790 & ~n4061;
  assign n4063 = next_sys_fair<0>_out  & ~n4062;
  assign n4064 = ~n3865 & ~n3894;
  assign n4065 = next_sys_fair<2>_out  & ~n4064;
  assign n4066 = reg_i_hlock3_out & ~n3215;
  assign n4067 = ~reg_i_hlock3_out & ~n3299;
  assign n4068 = ~n4066 & ~n4067;
  assign n4069 = reg_stateG10_3_out & ~n4068;
  assign n4070 = reg_i_hlock3_out & ~n3229;
  assign n4071 = ~reg_i_hlock3_out & ~n3313;
  assign n4072 = ~n4070 & ~n4071;
  assign n4073 = ~reg_stateG10_3_out & ~n4072;
  assign n4074 = ~n4069 & ~n4073;
  assign n4075 = reg_controllable_hgrant3_out & ~n4074;
  assign n4076 = ~n3853 & ~n4075;
  assign n4077 = ~next_sys_fair<2>_out  & ~n4076;
  assign n4078 = ~n4065 & ~n4077;
  assign n4079 = ~reg_controllable_hgrant4_out & ~n4078;
  assign n4080 = ~n3797 & ~n4079;
  assign n4081 = ~reg_controllable_hgrant5_out & ~n4080;
  assign n4082 = ~n3790 & ~n4081;
  assign n4083 = ~next_sys_fair<0>_out  & ~n4082;
  assign n4084 = ~n4063 & ~n4083;
  assign n4085 = ~next_sys_fair<3>_out  & ~n4084;
  assign n4086 = ~n3902 & ~n4085;
  assign n4087 = ~reg_controllable_hmaster2_out & ~n4086;
  assign n4088 = ~n4033 & ~n4087;
  assign n4089 = reg_controllable_hmaster1_out & ~n4088;
  assign n4090 = reg_stateG10_5_out & ~n3186;
  assign n4091 = ~reg_stateG10_5_out & ~n3201;
  assign n4092 = ~n4090 & ~n4091;
  assign n4093 = reg_i_hlock5_out & ~n4092;
  assign n4094 = reg_stateG10_5_out & ~n3271;
  assign n4095 = ~reg_stateG10_5_out & ~n3286;
  assign n4096 = ~n4094 & ~n4095;
  assign n4097 = ~reg_i_hlock5_out & ~n4096;
  assign n4098 = ~n4093 & ~n4097;
  assign n4099 = reg_controllable_hgrant5_out & ~n4098;
  assign n4100 = ~n3859 & ~n4099;
  assign n4101 = next_sys_fair<0>_out  & ~n4100;
  assign n4102 = reg_stateG10_5_out & ~n3221;
  assign n4103 = ~reg_stateG10_5_out & ~n3235;
  assign n4104 = ~n4102 & ~n4103;
  assign n4105 = reg_i_hlock5_out & ~n4104;
  assign n4106 = reg_stateG10_5_out & ~n3305;
  assign n4107 = ~reg_stateG10_5_out & ~n3319;
  assign n4108 = ~n4106 & ~n4107;
  assign n4109 = ~reg_i_hlock5_out & ~n4108;
  assign n4110 = ~n4105 & ~n4109;
  assign n4111 = reg_controllable_hgrant5_out & ~n4110;
  assign n4112 = ~n3871 & ~n4111;
  assign n4113 = ~next_sys_fair<0>_out  & ~n4112;
  assign n4114 = ~n4101 & ~n4113;
  assign n4115 = ~next_sys_fair<3>_out  & ~n4114;
  assign n4116 = ~n3934 & ~n4115;
  assign n4117 = reg_controllable_hmaster2_out & ~n4116;
  assign n4118 = ~n3804 & ~n3990;
  assign n4119 = next_sys_fair<2>_out  & ~n4118;
  assign n4120 = reg_stateG10_1_out & ~n3178;
  assign n4121 = ~reg_stateG10_1_out & ~n3193;
  assign n4122 = ~n4120 & ~n4121;
  assign n4123 = reg_i_hlock1_out & ~n4122;
  assign n4124 = reg_stateG10_1_out & ~n3263;
  assign n4125 = ~reg_stateG10_1_out & ~n3278;
  assign n4126 = ~n4124 & ~n4125;
  assign n4127 = ~reg_i_hlock1_out & ~n4126;
  assign n4128 = ~n4123 & ~n4127;
  assign n4129 = reg_controllable_hgrant1_out & ~n4128;
  assign n4130 = ~n3851 & ~n4129;
  assign n4131 = ~reg_controllable_hgrant3_out & ~n4130;
  assign n4132 = ~n3804 & ~n4131;
  assign n4133 = ~next_sys_fair<2>_out  & ~n4132;
  assign n4134 = ~n4119 & ~n4133;
  assign n4135 = ~reg_controllable_hgrant4_out & ~n4134;
  assign n4136 = ~n3797 & ~n4135;
  assign n4137 = ~reg_controllable_hgrant5_out & ~n4136;
  assign n4138 = ~n3790 & ~n4137;
  assign n4139 = next_sys_fair<0>_out  & ~n4138;
  assign n4140 = ~n3863 & ~n3988;
  assign n4141 = ~reg_controllable_hgrant3_out & ~n4140;
  assign n4142 = ~n3643 & ~n4141;
  assign n4143 = next_sys_fair<2>_out  & ~n4142;
  assign n4144 = reg_stateG10_1_out & ~n3213;
  assign n4145 = ~reg_stateG10_1_out & ~n3227;
  assign n4146 = ~n4144 & ~n4145;
  assign n4147 = reg_i_hlock1_out & ~n4146;
  assign n4148 = reg_stateG10_1_out & ~n3297;
  assign n4149 = ~reg_stateG10_1_out & ~n3311;
  assign n4150 = ~n4148 & ~n4149;
  assign n4151 = ~reg_i_hlock1_out & ~n4150;
  assign n4152 = ~n4147 & ~n4151;
  assign n4153 = reg_controllable_hgrant1_out & ~n4152;
  assign n4154 = ~n3851 & ~n4153;
  assign n4155 = ~reg_controllable_hgrant3_out & ~n4154;
  assign n4156 = ~n3804 & ~n4155;
  assign n4157 = ~next_sys_fair<2>_out  & ~n4156;
  assign n4158 = ~n4143 & ~n4157;
  assign n4159 = ~reg_controllable_hgrant4_out & ~n4158;
  assign n4160 = ~n3797 & ~n4159;
  assign n4161 = ~reg_controllable_hgrant5_out & ~n4160;
  assign n4162 = ~n3790 & ~n4161;
  assign n4163 = ~next_sys_fair<0>_out  & ~n4162;
  assign n4164 = ~n4139 & ~n4163;
  assign n4165 = ~next_sys_fair<3>_out  & ~n4164;
  assign n4166 = ~n3998 & ~n4165;
  assign n4167 = ~reg_controllable_hmaster2_out & ~n4166;
  assign n4168 = ~n4117 & ~n4167;
  assign n4169 = ~reg_controllable_hmaster1_out & ~n4168;
  assign n4170 = ~n4089 & ~n4169;
  assign n4171 = ~next_sys_fair<1>_out  & ~n4170;
  assign n4172 = ~n4032 & ~n4171;
  assign n4173 = reg_controllable_hmaster0_out & ~n4172;
  assign n4174 = reg_stateG10_2_out & ~n2982;
  assign n4175 = ~reg_stateG10_2_out & ~n3006;
  assign n4176 = ~n4174 & ~n4175;
  assign n4177 = reg_i_hlock2_out & ~n4176;
  assign n4178 = reg_stateG10_2_out & ~n3091;
  assign n4179 = ~reg_stateG10_2_out & ~n3108;
  assign n4180 = ~n4178 & ~n4179;
  assign n4181 = ~reg_i_hlock2_out & ~n4180;
  assign n4182 = ~n4177 & ~n4181;
  assign n4183 = reg_controllable_hgrant2_out & ~n4182;
  assign n4184 = ~n3747 & ~n4183;
  assign n4185 = ~reg_controllable_hgrant1_out & ~n4184;
  assign n4186 = ~n3650 & ~n4185;
  assign n4187 = ~reg_controllable_hgrant3_out & ~n4186;
  assign n4188 = ~n3643 & ~n4187;
  assign n4189 = ~next_sys_fair<2>_out  & ~n4188;
  assign n4190 = ~n663 & ~n4189;
  assign n4191 = ~reg_controllable_hgrant4_out & ~n4190;
  assign n4192 = ~n3636 & ~n4191;
  assign n4193 = ~reg_controllable_hgrant5_out & ~n4192;
  assign n4194 = ~n3629 & ~n4193;
  assign n4195 = next_sys_fair<3>_out  & ~n4194;
  assign n4196 = next_sys_fair<2>_out  & ~n4188;
  assign n4197 = ~n3710 & ~n4185;
  assign n4198 = ~reg_controllable_hgrant3_out & ~n4197;
  assign n4199 = ~n3643 & ~n4198;
  assign n4200 = ~next_sys_fair<2>_out  & ~n4199;
  assign n4201 = ~n4196 & ~n4200;
  assign n4202 = ~reg_controllable_hgrant4_out & ~n4201;
  assign n4203 = ~n3703 & ~n4202;
  assign n4204 = ~reg_controllable_hgrant5_out & ~n4203;
  assign n4205 = ~n3696 & ~n4204;
  assign n4206 = next_sys_fair<0>_out  & ~n4205;
  assign n4207 = ~reg_controllable_hgrant4_out & ~n4188;
  assign n4208 = ~n3734 & ~n4207;
  assign n4209 = ~reg_controllable_hgrant5_out & ~n4208;
  assign n4210 = ~n3727 & ~n4209;
  assign n4211 = ~next_sys_fair<0>_out  & ~n4210;
  assign n4212 = ~n4206 & ~n4211;
  assign n4213 = ~next_sys_fair<3>_out  & ~n4212;
  assign n4214 = ~n4195 & ~n4213;
  assign n4215 = ~reg_controllable_hmaster2_out & ~n4214;
  assign n4216 = ~n3884 & ~n4215;
  assign n4217 = reg_controllable_hmaster1_out & ~n4216;
  assign n4218 = reg_stateG10_4_out & ~n2990;
  assign n4219 = ~reg_stateG10_4_out & ~n3014;
  assign n4220 = ~n4218 & ~n4219;
  assign n4221 = reg_i_hlock4_out & ~n4220;
  assign n4222 = reg_stateG10_4_out & ~n3099;
  assign n4223 = ~reg_stateG10_4_out & ~n3116;
  assign n4224 = ~n4222 & ~n4223;
  assign n4225 = ~reg_i_hlock4_out & ~n4224;
  assign n4226 = ~n4221 & ~n4225;
  assign n4227 = reg_controllable_hgrant4_out & ~n4226;
  assign n4228 = ~n3755 & ~n4227;
  assign n4229 = ~reg_controllable_hgrant5_out & ~n4228;
  assign n4230 = ~n3629 & ~n4229;
  assign n4231 = next_sys_fair<3>_out  & ~n4230;
  assign n4232 = reg_stateG10_4_out & ~n2988;
  assign n4233 = ~reg_stateG10_4_out & ~n3012;
  assign n4234 = ~n4232 & ~n4233;
  assign n4235 = reg_i_hlock4_out & ~n4234;
  assign n4236 = reg_stateG10_4_out & ~n3097;
  assign n4237 = ~reg_stateG10_4_out & ~n3114;
  assign n4238 = ~n4236 & ~n4237;
  assign n4239 = ~reg_i_hlock4_out & ~n4238;
  assign n4240 = ~n4235 & ~n4239;
  assign n4241 = reg_controllable_hgrant4_out & ~n4240;
  assign n4242 = ~n3766 & ~n4241;
  assign n4243 = ~reg_controllable_hgrant5_out & ~n4242;
  assign n4244 = ~n3696 & ~n4243;
  assign n4245 = next_sys_fair<0>_out  & ~n4244;
  assign n4246 = reg_stateG10_4_out & ~n3936;
  assign n4247 = ~reg_stateG10_4_out & ~n3941;
  assign n4248 = ~n4246 & ~n4247;
  assign n4249 = reg_i_hlock4_out & ~n4248;
  assign n4250 = reg_stateG10_4_out & ~n3948;
  assign n4251 = ~reg_stateG10_4_out & ~n3953;
  assign n4252 = ~n4250 & ~n4251;
  assign n4253 = ~reg_i_hlock4_out & ~n4252;
  assign n4254 = ~n4249 & ~n4253;
  assign n4255 = reg_controllable_hgrant4_out & ~n4254;
  assign n4256 = ~n3771 & ~n4255;
  assign n4257 = ~reg_controllable_hgrant5_out & ~n4256;
  assign n4258 = ~n3727 & ~n4257;
  assign n4259 = ~next_sys_fair<0>_out  & ~n4258;
  assign n4260 = ~n4245 & ~n4259;
  assign n4261 = ~next_sys_fair<3>_out  & ~n4260;
  assign n4262 = ~n4231 & ~n4261;
  assign n4263 = reg_controllable_hmaster2_out & ~n4262;
  assign n4264 = ~n3779 & ~n4263;
  assign n4265 = ~reg_controllable_hmaster1_out & ~n4264;
  assign n4266 = ~n4217 & ~n4265;
  assign n4267 = next_sys_fair<1>_out  & ~n4266;
  assign n4268 = ~n3804 & ~n4187;
  assign n4269 = next_sys_fair<2>_out  & ~n4268;
  assign n4270 = reg_stateG10_2_out & ~n3176;
  assign n4271 = ~reg_stateG10_2_out & ~n3191;
  assign n4272 = ~n4270 & ~n4271;
  assign n4273 = reg_i_hlock2_out & ~n4272;
  assign n4274 = reg_stateG10_2_out & ~n3261;
  assign n4275 = ~reg_stateG10_2_out & ~n3276;
  assign n4276 = ~n4274 & ~n4275;
  assign n4277 = ~reg_i_hlock2_out & ~n4276;
  assign n4278 = ~n4273 & ~n4277;
  assign n4279 = reg_controllable_hgrant2_out & ~n4278;
  assign n4280 = ~n808 & ~n4279;
  assign n4281 = ~reg_controllable_hgrant1_out & ~n4280;
  assign n4282 = ~n3710 & ~n4281;
  assign n4283 = ~reg_controllable_hgrant3_out & ~n4282;
  assign n4284 = ~n3804 & ~n4283;
  assign n4285 = ~next_sys_fair<2>_out  & ~n4284;
  assign n4286 = ~n4269 & ~n4285;
  assign n4287 = ~reg_controllable_hgrant4_out & ~n4286;
  assign n4288 = ~n3797 & ~n4287;
  assign n4289 = ~reg_controllable_hgrant5_out & ~n4288;
  assign n4290 = ~n3790 & ~n4289;
  assign n4291 = next_sys_fair<0>_out  & ~n4290;
  assign n4292 = reg_stateG10_2_out & ~n2942;
  assign n4293 = ~reg_stateG10_2_out & ~n2956;
  assign n4294 = ~n4292 & ~n4293;
  assign n4295 = reg_i_hlock2_out & ~n4294;
  assign n4296 = reg_stateG10_2_out & ~n3055;
  assign n4297 = ~reg_stateG10_2_out & ~n3069;
  assign n4298 = ~n4296 & ~n4297;
  assign n4299 = ~reg_i_hlock2_out & ~n4298;
  assign n4300 = ~n4295 & ~n4299;
  assign n4301 = reg_controllable_hgrant2_out & ~n4300;
  assign n4302 = ~n3747 & ~n4301;
  assign n4303 = ~reg_controllable_hgrant1_out & ~n4302;
  assign n4304 = ~n3650 & ~n4303;
  assign n4305 = ~reg_controllable_hgrant3_out & ~n4304;
  assign n4306 = ~n3643 & ~n4305;
  assign n4307 = next_sys_fair<2>_out  & ~n4306;
  assign n4308 = reg_stateG10_2_out & ~n3211;
  assign n4309 = ~reg_stateG10_2_out & ~n3225;
  assign n4310 = ~n4308 & ~n4309;
  assign n4311 = reg_i_hlock2_out & ~n4310;
  assign n4312 = reg_stateG10_2_out & ~n3295;
  assign n4313 = ~reg_stateG10_2_out & ~n3309;
  assign n4314 = ~n4312 & ~n4313;
  assign n4315 = ~reg_i_hlock2_out & ~n4314;
  assign n4316 = ~n4311 & ~n4315;
  assign n4317 = reg_controllable_hgrant2_out & ~n4316;
  assign n4318 = ~n808 & ~n4317;
  assign n4319 = ~reg_controllable_hgrant1_out & ~n4318;
  assign n4320 = ~n3710 & ~n4319;
  assign n4321 = ~reg_controllable_hgrant3_out & ~n4320;
  assign n4322 = ~n3804 & ~n4321;
  assign n4323 = ~next_sys_fair<2>_out  & ~n4322;
  assign n4324 = ~n4307 & ~n4323;
  assign n4325 = ~reg_controllable_hgrant4_out & ~n4324;
  assign n4326 = ~n3797 & ~n4325;
  assign n4327 = ~reg_controllable_hgrant5_out & ~n4326;
  assign n4328 = ~n3790 & ~n4327;
  assign n4329 = ~next_sys_fair<0>_out  & ~n4328;
  assign n4330 = ~n4291 & ~n4329;
  assign n4331 = ~next_sys_fair<3>_out  & ~n4330;
  assign n4332 = ~n4195 & ~n4331;
  assign n4333 = ~reg_controllable_hmaster2_out & ~n4332;
  assign n4334 = ~n4033 & ~n4333;
  assign n4335 = reg_controllable_hmaster1_out & ~n4334;
  assign n4336 = reg_stateG10_4_out & ~n3184;
  assign n4337 = ~reg_stateG10_4_out & ~n3199;
  assign n4338 = ~n4336 & ~n4337;
  assign n4339 = reg_i_hlock4_out & ~n4338;
  assign n4340 = reg_stateG10_4_out & ~n3269;
  assign n4341 = ~reg_stateG10_4_out & ~n3284;
  assign n4342 = ~n4340 & ~n4341;
  assign n4343 = ~reg_i_hlock4_out & ~n4342;
  assign n4344 = ~n4339 & ~n4343;
  assign n4345 = reg_controllable_hgrant4_out & ~n4344;
  assign n4346 = ~n3857 & ~n4345;
  assign n4347 = ~reg_controllable_hgrant5_out & ~n4346;
  assign n4348 = ~n3790 & ~n4347;
  assign n4349 = next_sys_fair<0>_out  & ~n4348;
  assign n4350 = reg_stateG10_4_out & ~n3219;
  assign n4351 = ~reg_stateG10_4_out & ~n3233;
  assign n4352 = ~n4350 & ~n4351;
  assign n4353 = reg_i_hlock4_out & ~n4352;
  assign n4354 = reg_stateG10_4_out & ~n3303;
  assign n4355 = ~reg_stateG10_4_out & ~n3317;
  assign n4356 = ~n4354 & ~n4355;
  assign n4357 = ~reg_i_hlock4_out & ~n4356;
  assign n4358 = ~n4353 & ~n4357;
  assign n4359 = reg_controllable_hgrant4_out & ~n4358;
  assign n4360 = ~n3869 & ~n4359;
  assign n4361 = ~reg_controllable_hgrant5_out & ~n4360;
  assign n4362 = ~n3790 & ~n4361;
  assign n4363 = ~next_sys_fair<0>_out  & ~n4362;
  assign n4364 = ~n4349 & ~n4363;
  assign n4365 = ~next_sys_fair<3>_out  & ~n4364;
  assign n4366 = ~n4231 & ~n4365;
  assign n4367 = reg_controllable_hmaster2_out & ~n4366;
  assign n4368 = ~n3877 & ~n4367;
  assign n4369 = ~reg_controllable_hmaster1_out & ~n4368;
  assign n4370 = ~n4335 & ~n4369;
  assign n4371 = ~next_sys_fair<1>_out  & ~n4370;
  assign n4372 = ~n4267 & ~n4371;
  assign n4373 = ~reg_controllable_hmaster0_out & ~n4372;
  assign n4374 = ~n4173 & ~n4373;
  assign n4375 = ~reg_controllable_hmaster3_out & ~n4374;
  assign n4376 = ~n3883 & ~n4375;
  assign n4377 = ~reg_controllable_hgrant6_out & ~n4376;
  assign n4378 = ~n3622 & ~n4377;
  assign n4379 = ~reg_controllable_hgrant8_out & ~n4378;
  assign n4380 = ~n3523 & ~n4379;
  assign n4381 = ~reg_controllable_hgrant7_out & ~n4380;
  assign n4382 = ~n3449 & ~n4381;
  assign n4383 = ~reg_controllable_hgrant9_out & ~n4382;
  assign n4384 = ~n3357 & ~n4383;
  assign n4385 = reg_controllable_nhgrant0_out & ~n4384;
  assign n4386 = next_sys_fair<0>_out  & ~n2927;
  assign n4387 = ~next_sys_fair<0>_out  & ~n3159;
  assign n4388 = ~n4386 & ~n4387;
  assign n4389 = ~next_sys_fair<3>_out  & ~n4388;
  assign n4390 = ~n3399 & ~n4389;
  assign n4391 = next_sys_fair<1>_out  & ~n4390;
  assign n4392 = ~n3490 & ~n4391;
  assign n4393 = reg_controllable_hmaster3_out & ~n4392;
  assign n4394 = reg_controllable_hmaster0_out & ~n4392;
  assign n4395 = reg_controllable_hmaster1_out & ~n4390;
  assign n4396 = reg_controllable_hmaster2_out & ~n4390;
  assign n4397 = next_sys_fair<0>_out  & ~n3032;
  assign n4398 = ~n2963 & ~n3190;
  assign n4399 = ~reg_controllable_hgrant4_out & ~n4398;
  assign n4400 = ~reg_controllable_hgrant4_out & ~n4399;
  assign n4401 = ~reg_controllable_hgrant5_out & ~n4400;
  assign n4402 = ~reg_controllable_hgrant5_out & ~n4401;
  assign n4403 = ~next_sys_fair<0>_out  & ~n4402;
  assign n4404 = ~n4397 & ~n4403;
  assign n4405 = ~next_sys_fair<3>_out  & ~n4404;
  assign n4406 = ~n3411 & ~n4405;
  assign n4407 = ~reg_controllable_hmaster2_out & ~n4406;
  assign n4408 = ~n4396 & ~n4407;
  assign n4409 = ~reg_controllable_hmaster1_out & ~n4408;
  assign n4410 = ~n4395 & ~n4409;
  assign n4411 = next_sys_fair<1>_out  & ~n4410;
  assign n4412 = ~n3512 & ~n4411;
  assign n4413 = ~reg_controllable_hmaster0_out & ~n4412;
  assign n4414 = ~n4394 & ~n4413;
  assign n4415 = ~reg_controllable_hmaster3_out & ~n4414;
  assign n4416 = ~n4393 & ~n4415;
  assign n4417 = ~reg_controllable_hgrant6_out & ~n4416;
  assign n4418 = ~reg_controllable_hgrant6_out & ~n4417;
  assign n4419 = ~reg_controllable_hgrant8_out & ~n4418;
  assign n4420 = ~reg_controllable_hgrant8_out & ~n4419;
  assign n4421 = ~reg_controllable_hgrant7_out & ~n4420;
  assign n4422 = ~reg_controllable_hgrant7_out & ~n4421;
  assign n4423 = ~reg_controllable_hgrant9_out & ~n4422;
  assign n4424 = ~reg_controllable_hgrant9_out & ~n4423;
  assign n4425 = ~reg_controllable_nhgrant0_out & ~n4424;
  assign n4426 = ~n4385 & ~n4425;
  assign n4427 = reg_i_hready_out & ~n4426;
  assign n4428 = next_sys_fair<2>_out  & ~n545;
  assign n4429 = ~next_sys_fair<2>_out  & ~n3659;
  assign n4430 = ~n4428 & ~n4429;
  assign n4431 = next_sys_fair<3>_out  & ~n4430;
  assign n4432 = ~next_sys_fair<3>_out  & ~n3659;
  assign n4433 = ~n4431 & ~n4432;
  assign n4434 = reg_controllable_hmaster1_out & ~n4433;
  assign n4435 = reg_controllable_hmaster2_out & ~n4433;
  assign n4436 = ~n2936 & ~n2939;
  assign n4437 = ~next_sys_fair<2>_out  & ~n4436;
  assign n4438 = ~next_sys_fair<2>_out  & ~n4437;
  assign n4439 = reg_stateG10_9_out & ~n4438;
  assign n4440 = ~n218 & ~n2939;
  assign n4441 = ~next_sys_fair<2>_out  & ~n4440;
  assign n4442 = ~next_sys_fair<2>_out  & ~n4441;
  assign n4443 = ~reg_stateG10_9_out & ~n4442;
  assign n4444 = ~n4439 & ~n4443;
  assign n4445 = next_sys_fair<0>_out  & ~n4444;
  assign n4446 = ~n2975 & ~n2979;
  assign n4447 = ~next_sys_fair<2>_out  & ~n4446;
  assign n4448 = ~next_sys_fair<2>_out  & ~n4447;
  assign n4449 = reg_stateG10_9_out & ~n4448;
  assign n4450 = ~n2979 & ~n3003;
  assign n4451 = ~next_sys_fair<2>_out  & ~n4450;
  assign n4452 = ~next_sys_fair<2>_out  & ~n4451;
  assign n4453 = ~reg_stateG10_9_out & ~n4452;
  assign n4454 = ~n4449 & ~n4453;
  assign n4455 = ~next_sys_fair<0>_out  & ~n4454;
  assign n4456 = ~n4445 & ~n4455;
  assign n4457 = next_sys_fair<3>_out  & ~n4456;
  assign n4458 = reg_stateG10_9_out & ~n4446;
  assign n4459 = ~reg_stateG10_9_out & ~n4450;
  assign n4460 = ~n4458 & ~n4459;
  assign n4461 = ~next_sys_fair<3>_out  & ~n4460;
  assign n4462 = ~n4457 & ~n4461;
  assign n4463 = ~reg_controllable_hmaster2_out & ~n4462;
  assign n4464 = ~n4435 & ~n4463;
  assign n4465 = ~reg_controllable_hmaster1_out & ~n4464;
  assign n4466 = ~n4434 & ~n4465;
  assign n4467 = reg_i_hlock9_out & ~n4466;
  assign n4468 = ~n1296 & ~n3052;
  assign n4469 = ~next_sys_fair<2>_out  & ~n4468;
  assign n4470 = ~next_sys_fair<2>_out  & ~n4469;
  assign n4471 = reg_stateG10_9_out & ~n4470;
  assign n4472 = ~next_sys_fair<2>_out  & ~n1297;
  assign n4473 = ~next_sys_fair<2>_out  & ~n4472;
  assign n4474 = ~reg_stateG10_9_out & ~n4473;
  assign n4475 = ~n4471 & ~n4474;
  assign n4476 = next_sys_fair<0>_out  & ~n4475;
  assign n4477 = ~n3085 & ~n3088;
  assign n4478 = ~next_sys_fair<2>_out  & ~n4477;
  assign n4479 = ~next_sys_fair<2>_out  & ~n4478;
  assign n4480 = reg_stateG10_9_out & ~n4479;
  assign n4481 = ~n3085 & ~n3105;
  assign n4482 = ~next_sys_fair<2>_out  & ~n4481;
  assign n4483 = ~next_sys_fair<2>_out  & ~n4482;
  assign n4484 = ~reg_stateG10_9_out & ~n4483;
  assign n4485 = ~n4480 & ~n4484;
  assign n4486 = ~next_sys_fair<0>_out  & ~n4485;
  assign n4487 = ~n4476 & ~n4486;
  assign n4488 = next_sys_fair<3>_out  & ~n4487;
  assign n4489 = reg_stateG10_9_out & ~n4477;
  assign n4490 = ~reg_stateG10_9_out & ~n4481;
  assign n4491 = ~n4489 & ~n4490;
  assign n4492 = ~next_sys_fair<3>_out  & ~n4491;
  assign n4493 = ~n4488 & ~n4492;
  assign n4494 = ~reg_controllable_hmaster2_out & ~n4493;
  assign n4495 = ~n4435 & ~n4494;
  assign n4496 = ~reg_controllable_hmaster1_out & ~n4495;
  assign n4497 = ~n4434 & ~n4496;
  assign n4498 = ~reg_i_hlock9_out & ~n4497;
  assign n4499 = ~n4467 & ~n4498;
  assign n4500 = next_sys_fair<1>_out  & ~n4499;
  assign n4501 = next_sys_fair<2>_out  & ~n3659;
  assign n4502 = ~next_sys_fair<2>_out  & ~n733;
  assign n4503 = ~n4501 & ~n4502;
  assign n4504 = next_sys_fair<0>_out  & ~n4503;
  assign n4505 = ~next_sys_fair<2>_out  & ~n780;
  assign n4506 = ~n4501 & ~n4505;
  assign n4507 = ~next_sys_fair<0>_out  & ~n4506;
  assign n4508 = ~n4504 & ~n4507;
  assign n4509 = ~next_sys_fair<3>_out  & ~n4508;
  assign n4510 = ~n4431 & ~n4509;
  assign n4511 = reg_controllable_hmaster1_out & ~n4510;
  assign n4512 = reg_controllable_hmaster2_out & ~n4510;
  assign n4513 = next_sys_fair<3>_out  & ~n4454;
  assign n4514 = next_sys_fair<2>_out  & ~n4446;
  assign n4515 = ~n3170 & ~n3173;
  assign n4516 = ~next_sys_fair<2>_out  & ~n4515;
  assign n4517 = ~n4514 & ~n4516;
  assign n4518 = reg_stateG10_9_out & ~n4517;
  assign n4519 = next_sys_fair<2>_out  & ~n4450;
  assign n4520 = ~n335 & ~n3173;
  assign n4521 = ~next_sys_fair<2>_out  & ~n4520;
  assign n4522 = ~n4519 & ~n4521;
  assign n4523 = ~reg_stateG10_9_out & ~n4522;
  assign n4524 = ~n4518 & ~n4523;
  assign n4525 = next_sys_fair<0>_out  & ~n4524;
  assign n4526 = ~n2939 & ~n3208;
  assign n4527 = ~next_sys_fair<2>_out  & ~n4526;
  assign n4528 = ~n4514 & ~n4527;
  assign n4529 = reg_stateG10_9_out & ~n4528;
  assign n4530 = ~n366 & ~n2939;
  assign n4531 = ~next_sys_fair<2>_out  & ~n4530;
  assign n4532 = ~n4519 & ~n4531;
  assign n4533 = ~reg_stateG10_9_out & ~n4532;
  assign n4534 = ~n4529 & ~n4533;
  assign n4535 = ~next_sys_fair<0>_out  & ~n4534;
  assign n4536 = ~n4525 & ~n4535;
  assign n4537 = ~next_sys_fair<3>_out  & ~n4536;
  assign n4538 = ~n4513 & ~n4537;
  assign n4539 = ~reg_controllable_hmaster2_out & ~n4538;
  assign n4540 = ~n4512 & ~n4539;
  assign n4541 = ~reg_controllable_hmaster1_out & ~n4540;
  assign n4542 = ~n4511 & ~n4541;
  assign n4543 = reg_i_hlock9_out & ~n4542;
  assign n4544 = next_sys_fair<3>_out  & ~n4485;
  assign n4545 = next_sys_fair<2>_out  & ~n4477;
  assign n4546 = ~n1427 & ~n3258;
  assign n4547 = ~next_sys_fair<2>_out  & ~n4546;
  assign n4548 = ~n4545 & ~n4547;
  assign n4549 = reg_stateG10_9_out & ~n4548;
  assign n4550 = next_sys_fair<2>_out  & ~n4481;
  assign n4551 = ~next_sys_fair<2>_out  & ~n1428;
  assign n4552 = ~n4550 & ~n4551;
  assign n4553 = ~reg_stateG10_9_out & ~n4552;
  assign n4554 = ~n4549 & ~n4553;
  assign n4555 = next_sys_fair<0>_out  & ~n4554;
  assign n4556 = ~n1296 & ~n3292;
  assign n4557 = ~next_sys_fair<2>_out  & ~n4556;
  assign n4558 = ~n4545 & ~n4557;
  assign n4559 = reg_stateG10_9_out & ~n4558;
  assign n4560 = ~next_sys_fair<2>_out  & ~n1448;
  assign n4561 = ~n4550 & ~n4560;
  assign n4562 = ~reg_stateG10_9_out & ~n4561;
  assign n4563 = ~n4559 & ~n4562;
  assign n4564 = ~next_sys_fair<0>_out  & ~n4563;
  assign n4565 = ~n4555 & ~n4564;
  assign n4566 = ~next_sys_fair<3>_out  & ~n4565;
  assign n4567 = ~n4544 & ~n4566;
  assign n4568 = ~reg_controllable_hmaster2_out & ~n4567;
  assign n4569 = ~n4512 & ~n4568;
  assign n4570 = ~reg_controllable_hmaster1_out & ~n4569;
  assign n4571 = ~n4511 & ~n4570;
  assign n4572 = ~reg_i_hlock9_out & ~n4571;
  assign n4573 = ~n4543 & ~n4572;
  assign n4574 = ~next_sys_fair<1>_out  & ~n4573;
  assign n4575 = ~n4500 & ~n4574;
  assign n4576 = reg_controllable_hmaster0_out & ~n4575;
  assign n4577 = next_sys_fair<0>_out  & ~n4448;
  assign n4578 = ~next_sys_fair<0>_out  & ~n4438;
  assign n4579 = ~n4577 & ~n4578;
  assign n4580 = next_sys_fair<3>_out  & ~n4579;
  assign n4581 = ~next_sys_fair<3>_out  & ~n4446;
  assign n4582 = ~n4580 & ~n4581;
  assign n4583 = ~reg_controllable_hmaster2_out & ~n4582;
  assign n4584 = ~n4435 & ~n4583;
  assign n4585 = ~reg_controllable_hmaster1_out & ~n4584;
  assign n4586 = ~n4434 & ~n4585;
  assign n4587 = next_sys_fair<1>_out  & ~n4586;
  assign n4588 = next_sys_fair<3>_out  & ~n4448;
  assign n4589 = next_sys_fair<0>_out  & ~n4517;
  assign n4590 = ~next_sys_fair<0>_out  & ~n4528;
  assign n4591 = ~n4589 & ~n4590;
  assign n4592 = ~next_sys_fair<3>_out  & ~n4591;
  assign n4593 = ~n4588 & ~n4592;
  assign n4594 = ~reg_controllable_hmaster2_out & ~n4593;
  assign n4595 = ~n4512 & ~n4594;
  assign n4596 = ~reg_controllable_hmaster1_out & ~n4595;
  assign n4597 = ~n4511 & ~n4596;
  assign n4598 = ~next_sys_fair<1>_out  & ~n4597;
  assign n4599 = ~n4587 & ~n4598;
  assign n4600 = ~reg_controllable_hmaster0_out & ~n4599;
  assign n4601 = ~n4576 & ~n4600;
  assign n4602 = reg_controllable_hmaster3_out & ~n4601;
  assign n4603 = ~n4581 & ~n4588;
  assign n4604 = reg_controllable_hmaster2_out & ~n4603;
  assign n4605 = reg_i_hlock3_out & ~n4446;
  assign n4606 = ~reg_i_hlock3_out & ~n4477;
  assign n4607 = ~n4605 & ~n4606;
  assign n4608 = reg_stateG10_3_out & ~n4607;
  assign n4609 = reg_i_hlock3_out & ~n4450;
  assign n4610 = ~reg_i_hlock3_out & ~n4481;
  assign n4611 = ~n4609 & ~n4610;
  assign n4612 = ~reg_stateG10_3_out & ~n4611;
  assign n4613 = ~n4608 & ~n4612;
  assign n4614 = ~next_sys_fair<2>_out  & ~n4613;
  assign n4615 = ~next_sys_fair<2>_out  & ~n4614;
  assign n4616 = next_sys_fair<3>_out  & ~n4615;
  assign n4617 = ~next_sys_fair<3>_out  & ~n4613;
  assign n4618 = ~n4616 & ~n4617;
  assign n4619 = ~reg_controllable_hmaster2_out & ~n4618;
  assign n4620 = ~n4604 & ~n4619;
  assign n4621 = reg_controllable_hmaster1_out & ~n4620;
  assign n4622 = reg_stateG10_5_out & ~n4448;
  assign n4623 = ~reg_stateG10_5_out & ~n4452;
  assign n4624 = ~n4622 & ~n4623;
  assign n4625 = reg_i_hlock5_out & ~n4624;
  assign n4626 = reg_stateG10_5_out & ~n4479;
  assign n4627 = ~reg_stateG10_5_out & ~n4483;
  assign n4628 = ~n4626 & ~n4627;
  assign n4629 = ~reg_i_hlock5_out & ~n4628;
  assign n4630 = ~n4625 & ~n4629;
  assign n4631 = next_sys_fair<3>_out  & ~n4630;
  assign n4632 = next_sys_fair<2>_out  & ~n4436;
  assign n4633 = ~n4447 & ~n4632;
  assign n4634 = reg_stateG10_5_out & ~n4633;
  assign n4635 = next_sys_fair<2>_out  & ~n4440;
  assign n4636 = ~n4451 & ~n4635;
  assign n4637 = ~reg_stateG10_5_out & ~n4636;
  assign n4638 = ~n4634 & ~n4637;
  assign n4639 = reg_i_hlock5_out & ~n4638;
  assign n4640 = next_sys_fair<2>_out  & ~n4468;
  assign n4641 = ~n4478 & ~n4640;
  assign n4642 = reg_stateG10_5_out & ~n4641;
  assign n4643 = next_sys_fair<2>_out  & ~n1297;
  assign n4644 = ~n4482 & ~n4643;
  assign n4645 = ~reg_stateG10_5_out & ~n4644;
  assign n4646 = ~n4642 & ~n4645;
  assign n4647 = ~reg_i_hlock5_out & ~n4646;
  assign n4648 = ~n4639 & ~n4647;
  assign n4649 = next_sys_fair<0>_out  & ~n4648;
  assign n4650 = reg_stateG10_5_out & ~n4446;
  assign n4651 = ~reg_stateG10_5_out & ~n4450;
  assign n4652 = ~n4650 & ~n4651;
  assign n4653 = reg_i_hlock5_out & ~n4652;
  assign n4654 = reg_stateG10_5_out & ~n4477;
  assign n4655 = ~reg_stateG10_5_out & ~n4481;
  assign n4656 = ~n4654 & ~n4655;
  assign n4657 = ~reg_i_hlock5_out & ~n4656;
  assign n4658 = ~n4653 & ~n4657;
  assign n4659 = ~next_sys_fair<0>_out  & ~n4658;
  assign n4660 = ~n4649 & ~n4659;
  assign n4661 = ~next_sys_fair<3>_out  & ~n4660;
  assign n4662 = ~n4631 & ~n4661;
  assign n4663 = reg_controllable_hmaster2_out & ~n4662;
  assign n4664 = reg_stateG10_1_out & ~n4446;
  assign n4665 = ~reg_stateG10_1_out & ~n4450;
  assign n4666 = ~n4664 & ~n4665;
  assign n4667 = reg_i_hlock1_out & ~n4666;
  assign n4668 = reg_stateG10_1_out & ~n4477;
  assign n4669 = ~reg_stateG10_1_out & ~n4481;
  assign n4670 = ~n4668 & ~n4669;
  assign n4671 = ~reg_i_hlock1_out & ~n4670;
  assign n4672 = ~n4667 & ~n4671;
  assign n4673 = ~next_sys_fair<2>_out  & ~n4672;
  assign n4674 = ~next_sys_fair<2>_out  & ~n4673;
  assign n4675 = next_sys_fair<3>_out  & ~n4674;
  assign n4676 = next_sys_fair<2>_out  & ~n4672;
  assign n4677 = reg_stateG10_1_out & ~n4436;
  assign n4678 = ~reg_stateG10_1_out & ~n4440;
  assign n4679 = ~n4677 & ~n4678;
  assign n4680 = reg_i_hlock1_out & ~n4679;
  assign n4681 = reg_stateG10_1_out & ~n4468;
  assign n4682 = ~reg_stateG10_1_out & ~n1297;
  assign n4683 = ~n4681 & ~n4682;
  assign n4684 = ~reg_i_hlock1_out & ~n4683;
  assign n4685 = ~n4680 & ~n4684;
  assign n4686 = ~next_sys_fair<2>_out  & ~n4685;
  assign n4687 = ~n4676 & ~n4686;
  assign n4688 = next_sys_fair<0>_out  & ~n4687;
  assign n4689 = ~next_sys_fair<0>_out  & ~n4672;
  assign n4690 = ~n4688 & ~n4689;
  assign n4691 = ~next_sys_fair<3>_out  & ~n4690;
  assign n4692 = ~n4675 & ~n4691;
  assign n4693 = ~reg_controllable_hmaster2_out & ~n4692;
  assign n4694 = ~n4663 & ~n4693;
  assign n4695 = ~reg_controllable_hmaster1_out & ~n4694;
  assign n4696 = ~n4621 & ~n4695;
  assign n4697 = next_sys_fair<1>_out  & ~n4696;
  assign n4698 = next_sys_fair<0>_out  & ~n4438;
  assign n4699 = ~next_sys_fair<0>_out  & ~n4448;
  assign n4700 = ~n4698 & ~n4699;
  assign n4701 = next_sys_fair<3>_out  & ~n4700;
  assign n4702 = ~n4592 & ~n4701;
  assign n4703 = reg_controllable_hmaster2_out & ~n4702;
  assign n4704 = reg_i_hlock3_out & ~n4436;
  assign n4705 = ~reg_i_hlock3_out & ~n4468;
  assign n4706 = ~n4704 & ~n4705;
  assign n4707 = reg_stateG10_3_out & ~n4706;
  assign n4708 = reg_i_hlock3_out & ~n4440;
  assign n4709 = ~reg_i_hlock3_out & ~n1297;
  assign n4710 = ~n4708 & ~n4709;
  assign n4711 = ~reg_stateG10_3_out & ~n4710;
  assign n4712 = ~n4707 & ~n4711;
  assign n4713 = next_sys_fair<2>_out  & ~n4712;
  assign n4714 = reg_i_hlock3_out & ~n4515;
  assign n4715 = ~reg_i_hlock3_out & ~n4546;
  assign n4716 = ~n4714 & ~n4715;
  assign n4717 = reg_stateG10_3_out & ~n4716;
  assign n4718 = reg_i_hlock3_out & ~n4520;
  assign n4719 = ~reg_i_hlock3_out & ~n1428;
  assign n4720 = ~n4718 & ~n4719;
  assign n4721 = ~reg_stateG10_3_out & ~n4720;
  assign n4722 = ~n4717 & ~n4721;
  assign n4723 = ~next_sys_fair<2>_out  & ~n4722;
  assign n4724 = ~n4713 & ~n4723;
  assign n4725 = next_sys_fair<0>_out  & ~n4724;
  assign n4726 = next_sys_fair<2>_out  & ~n4613;
  assign n4727 = reg_i_hlock3_out & ~n4526;
  assign n4728 = ~reg_i_hlock3_out & ~n4556;
  assign n4729 = ~n4727 & ~n4728;
  assign n4730 = reg_stateG10_3_out & ~n4729;
  assign n4731 = reg_i_hlock3_out & ~n4530;
  assign n4732 = ~reg_i_hlock3_out & ~n1448;
  assign n4733 = ~n4731 & ~n4732;
  assign n4734 = ~reg_stateG10_3_out & ~n4733;
  assign n4735 = ~n4730 & ~n4734;
  assign n4736 = ~next_sys_fair<2>_out  & ~n4735;
  assign n4737 = ~n4726 & ~n4736;
  assign n4738 = ~next_sys_fair<0>_out  & ~n4737;
  assign n4739 = ~n4725 & ~n4738;
  assign n4740 = ~next_sys_fair<3>_out  & ~n4739;
  assign n4741 = ~n4616 & ~n4740;
  assign n4742 = ~reg_controllable_hmaster2_out & ~n4741;
  assign n4743 = ~n4703 & ~n4742;
  assign n4744 = reg_controllable_hmaster1_out & ~n4743;
  assign n4745 = reg_stateG10_5_out & ~n4517;
  assign n4746 = ~reg_stateG10_5_out & ~n4522;
  assign n4747 = ~n4745 & ~n4746;
  assign n4748 = reg_i_hlock5_out & ~n4747;
  assign n4749 = reg_stateG10_5_out & ~n4548;
  assign n4750 = ~reg_stateG10_5_out & ~n4552;
  assign n4751 = ~n4749 & ~n4750;
  assign n4752 = ~reg_i_hlock5_out & ~n4751;
  assign n4753 = ~n4748 & ~n4752;
  assign n4754 = next_sys_fair<0>_out  & ~n4753;
  assign n4755 = reg_stateG10_5_out & ~n4528;
  assign n4756 = ~reg_stateG10_5_out & ~n4532;
  assign n4757 = ~n4755 & ~n4756;
  assign n4758 = reg_i_hlock5_out & ~n4757;
  assign n4759 = reg_stateG10_5_out & ~n4558;
  assign n4760 = ~reg_stateG10_5_out & ~n4561;
  assign n4761 = ~n4759 & ~n4760;
  assign n4762 = ~reg_i_hlock5_out & ~n4761;
  assign n4763 = ~n4758 & ~n4762;
  assign n4764 = ~next_sys_fair<0>_out  & ~n4763;
  assign n4765 = ~n4754 & ~n4764;
  assign n4766 = ~next_sys_fair<3>_out  & ~n4765;
  assign n4767 = ~n4631 & ~n4766;
  assign n4768 = reg_controllable_hmaster2_out & ~n4767;
  assign n4769 = reg_stateG10_1_out & ~n4515;
  assign n4770 = ~reg_stateG10_1_out & ~n4520;
  assign n4771 = ~n4769 & ~n4770;
  assign n4772 = reg_i_hlock1_out & ~n4771;
  assign n4773 = reg_stateG10_1_out & ~n4546;
  assign n4774 = ~reg_stateG10_1_out & ~n1428;
  assign n4775 = ~n4773 & ~n4774;
  assign n4776 = ~reg_i_hlock1_out & ~n4775;
  assign n4777 = ~n4772 & ~n4776;
  assign n4778 = ~next_sys_fair<2>_out  & ~n4777;
  assign n4779 = ~n4676 & ~n4778;
  assign n4780 = next_sys_fair<0>_out  & ~n4779;
  assign n4781 = reg_stateG10_1_out & ~n4526;
  assign n4782 = ~reg_stateG10_1_out & ~n4530;
  assign n4783 = ~n4781 & ~n4782;
  assign n4784 = reg_i_hlock1_out & ~n4783;
  assign n4785 = reg_stateG10_1_out & ~n4556;
  assign n4786 = ~reg_stateG10_1_out & ~n1448;
  assign n4787 = ~n4785 & ~n4786;
  assign n4788 = ~reg_i_hlock1_out & ~n4787;
  assign n4789 = ~n4784 & ~n4788;
  assign n4790 = ~next_sys_fair<2>_out  & ~n4789;
  assign n4791 = ~n4676 & ~n4790;
  assign n4792 = ~next_sys_fair<0>_out  & ~n4791;
  assign n4793 = ~n4780 & ~n4792;
  assign n4794 = ~next_sys_fair<3>_out  & ~n4793;
  assign n4795 = ~n4675 & ~n4794;
  assign n4796 = ~reg_controllable_hmaster2_out & ~n4795;
  assign n4797 = ~n4768 & ~n4796;
  assign n4798 = ~reg_controllable_hmaster1_out & ~n4797;
  assign n4799 = ~n4744 & ~n4798;
  assign n4800 = ~next_sys_fair<1>_out  & ~n4799;
  assign n4801 = ~n4697 & ~n4800;
  assign n4802 = reg_controllable_hmaster0_out & ~n4801;
  assign n4803 = reg_stateG10_2_out & ~n4446;
  assign n4804 = ~reg_stateG10_2_out & ~n4450;
  assign n4805 = ~n4803 & ~n4804;
  assign n4806 = reg_i_hlock2_out & ~n4805;
  assign n4807 = reg_stateG10_2_out & ~n4477;
  assign n4808 = ~reg_stateG10_2_out & ~n4481;
  assign n4809 = ~n4807 & ~n4808;
  assign n4810 = ~reg_i_hlock2_out & ~n4809;
  assign n4811 = ~n4806 & ~n4810;
  assign n4812 = ~next_sys_fair<2>_out  & ~n4811;
  assign n4813 = ~next_sys_fair<2>_out  & ~n4812;
  assign n4814 = next_sys_fair<3>_out  & ~n4813;
  assign n4815 = ~next_sys_fair<3>_out  & ~n4811;
  assign n4816 = ~n4814 & ~n4815;
  assign n4817 = ~reg_controllable_hmaster2_out & ~n4816;
  assign n4818 = ~n4604 & ~n4817;
  assign n4819 = reg_controllable_hmaster1_out & ~n4818;
  assign n4820 = reg_stateG10_4_out & ~n4448;
  assign n4821 = ~reg_stateG10_4_out & ~n4452;
  assign n4822 = ~n4820 & ~n4821;
  assign n4823 = reg_i_hlock4_out & ~n4822;
  assign n4824 = reg_stateG10_4_out & ~n4479;
  assign n4825 = ~reg_stateG10_4_out & ~n4483;
  assign n4826 = ~n4824 & ~n4825;
  assign n4827 = ~reg_i_hlock4_out & ~n4826;
  assign n4828 = ~n4823 & ~n4827;
  assign n4829 = next_sys_fair<3>_out  & ~n4828;
  assign n4830 = reg_stateG10_4_out & ~n4446;
  assign n4831 = ~reg_stateG10_4_out & ~n4450;
  assign n4832 = ~n4830 & ~n4831;
  assign n4833 = reg_i_hlock4_out & ~n4832;
  assign n4834 = reg_stateG10_4_out & ~n4477;
  assign n4835 = ~reg_stateG10_4_out & ~n4481;
  assign n4836 = ~n4834 & ~n4835;
  assign n4837 = ~reg_i_hlock4_out & ~n4836;
  assign n4838 = ~n4833 & ~n4837;
  assign n4839 = next_sys_fair<0>_out  & ~n4838;
  assign n4840 = reg_stateG10_4_out & ~n4633;
  assign n4841 = ~reg_stateG10_4_out & ~n4636;
  assign n4842 = ~n4840 & ~n4841;
  assign n4843 = reg_i_hlock4_out & ~n4842;
  assign n4844 = reg_stateG10_4_out & ~n4641;
  assign n4845 = ~reg_stateG10_4_out & ~n4644;
  assign n4846 = ~n4844 & ~n4845;
  assign n4847 = ~reg_i_hlock4_out & ~n4846;
  assign n4848 = ~n4843 & ~n4847;
  assign n4849 = ~next_sys_fair<0>_out  & ~n4848;
  assign n4850 = ~n4839 & ~n4849;
  assign n4851 = ~next_sys_fair<3>_out  & ~n4850;
  assign n4852 = ~n4829 & ~n4851;
  assign n4853 = reg_controllable_hmaster2_out & ~n4852;
  assign n4854 = next_sys_fair<3>_out  & ~n4452;
  assign n4855 = next_sys_fair<0>_out  & ~n4450;
  assign n4856 = ~n4441 & ~n4519;
  assign n4857 = ~next_sys_fair<0>_out  & ~n4856;
  assign n4858 = ~n4855 & ~n4857;
  assign n4859 = ~next_sys_fair<3>_out  & ~n4858;
  assign n4860 = ~n4854 & ~n4859;
  assign n4861 = ~reg_controllable_hmaster2_out & ~n4860;
  assign n4862 = ~n4853 & ~n4861;
  assign n4863 = ~reg_controllable_hmaster1_out & ~n4862;
  assign n4864 = ~n4819 & ~n4863;
  assign n4865 = reg_stateG10_6_out & ~n4864;
  assign n4866 = ~next_sys_fair<3>_out  & ~n4450;
  assign n4867 = ~n4854 & ~n4866;
  assign n4868 = reg_controllable_hmaster2_out & ~n4867;
  assign n4869 = ~n4817 & ~n4868;
  assign n4870 = reg_controllable_hmaster1_out & ~n4869;
  assign n4871 = ~n4863 & ~n4870;
  assign n4872 = ~reg_stateG10_6_out & ~n4871;
  assign n4873 = ~n4865 & ~n4872;
  assign n4874 = reg_i_hlock6_out & ~n4873;
  assign n4875 = next_sys_fair<3>_out  & ~n4479;
  assign n4876 = ~next_sys_fair<3>_out  & ~n4477;
  assign n4877 = ~n4875 & ~n4876;
  assign n4878 = reg_controllable_hmaster2_out & ~n4877;
  assign n4879 = ~n4817 & ~n4878;
  assign n4880 = reg_controllable_hmaster1_out & ~n4879;
  assign n4881 = ~n4863 & ~n4880;
  assign n4882 = reg_stateG10_6_out & ~n4881;
  assign n4883 = next_sys_fair<3>_out  & ~n4483;
  assign n4884 = ~next_sys_fair<3>_out  & ~n4481;
  assign n4885 = ~n4883 & ~n4884;
  assign n4886 = reg_controllable_hmaster2_out & ~n4885;
  assign n4887 = ~n4817 & ~n4886;
  assign n4888 = reg_controllable_hmaster1_out & ~n4887;
  assign n4889 = ~n4863 & ~n4888;
  assign n4890 = ~reg_stateG10_6_out & ~n4889;
  assign n4891 = ~n4882 & ~n4890;
  assign n4892 = ~reg_i_hlock6_out & ~n4891;
  assign n4893 = ~n4874 & ~n4892;
  assign n4894 = next_sys_fair<1>_out  & ~n4893;
  assign n4895 = ~n4580 & ~n4592;
  assign n4896 = reg_controllable_hmaster2_out & ~n4895;
  assign n4897 = next_sys_fair<2>_out  & ~n4811;
  assign n4898 = reg_stateG10_2_out & ~n4515;
  assign n4899 = ~reg_stateG10_2_out & ~n4520;
  assign n4900 = ~n4898 & ~n4899;
  assign n4901 = reg_i_hlock2_out & ~n4900;
  assign n4902 = reg_stateG10_2_out & ~n4546;
  assign n4903 = ~reg_stateG10_2_out & ~n1428;
  assign n4904 = ~n4902 & ~n4903;
  assign n4905 = ~reg_i_hlock2_out & ~n4904;
  assign n4906 = ~n4901 & ~n4905;
  assign n4907 = ~next_sys_fair<2>_out  & ~n4906;
  assign n4908 = ~n4897 & ~n4907;
  assign n4909 = next_sys_fair<0>_out  & ~n4908;
  assign n4910 = reg_stateG10_2_out & ~n4436;
  assign n4911 = ~reg_stateG10_2_out & ~n4440;
  assign n4912 = ~n4910 & ~n4911;
  assign n4913 = reg_i_hlock2_out & ~n4912;
  assign n4914 = reg_stateG10_2_out & ~n4468;
  assign n4915 = ~reg_stateG10_2_out & ~n1297;
  assign n4916 = ~n4914 & ~n4915;
  assign n4917 = ~reg_i_hlock2_out & ~n4916;
  assign n4918 = ~n4913 & ~n4917;
  assign n4919 = next_sys_fair<2>_out  & ~n4918;
  assign n4920 = reg_stateG10_2_out & ~n4526;
  assign n4921 = ~reg_stateG10_2_out & ~n4530;
  assign n4922 = ~n4920 & ~n4921;
  assign n4923 = reg_i_hlock2_out & ~n4922;
  assign n4924 = reg_stateG10_2_out & ~n4556;
  assign n4925 = ~reg_stateG10_2_out & ~n1448;
  assign n4926 = ~n4924 & ~n4925;
  assign n4927 = ~reg_i_hlock2_out & ~n4926;
  assign n4928 = ~n4923 & ~n4927;
  assign n4929 = ~next_sys_fair<2>_out  & ~n4928;
  assign n4930 = ~n4919 & ~n4929;
  assign n4931 = ~next_sys_fair<0>_out  & ~n4930;
  assign n4932 = ~n4909 & ~n4931;
  assign n4933 = ~next_sys_fair<3>_out  & ~n4932;
  assign n4934 = ~n4814 & ~n4933;
  assign n4935 = ~reg_controllable_hmaster2_out & ~n4934;
  assign n4936 = ~n4896 & ~n4935;
  assign n4937 = reg_controllable_hmaster1_out & ~n4936;
  assign n4938 = reg_stateG10_4_out & ~n4517;
  assign n4939 = ~reg_stateG10_4_out & ~n4522;
  assign n4940 = ~n4938 & ~n4939;
  assign n4941 = reg_i_hlock4_out & ~n4940;
  assign n4942 = reg_stateG10_4_out & ~n4548;
  assign n4943 = ~reg_stateG10_4_out & ~n4552;
  assign n4944 = ~n4942 & ~n4943;
  assign n4945 = ~reg_i_hlock4_out & ~n4944;
  assign n4946 = ~n4941 & ~n4945;
  assign n4947 = next_sys_fair<0>_out  & ~n4946;
  assign n4948 = reg_stateG10_4_out & ~n4528;
  assign n4949 = ~reg_stateG10_4_out & ~n4532;
  assign n4950 = ~n4948 & ~n4949;
  assign n4951 = reg_i_hlock4_out & ~n4950;
  assign n4952 = reg_stateG10_4_out & ~n4558;
  assign n4953 = ~reg_stateG10_4_out & ~n4561;
  assign n4954 = ~n4952 & ~n4953;
  assign n4955 = ~reg_i_hlock4_out & ~n4954;
  assign n4956 = ~n4951 & ~n4955;
  assign n4957 = ~next_sys_fair<0>_out  & ~n4956;
  assign n4958 = ~n4947 & ~n4957;
  assign n4959 = ~next_sys_fair<3>_out  & ~n4958;
  assign n4960 = ~n4829 & ~n4959;
  assign n4961 = reg_controllable_hmaster2_out & ~n4960;
  assign n4962 = next_sys_fair<0>_out  & ~n4522;
  assign n4963 = ~next_sys_fair<0>_out  & ~n4532;
  assign n4964 = ~n4962 & ~n4963;
  assign n4965 = ~next_sys_fair<3>_out  & ~n4964;
  assign n4966 = ~n4854 & ~n4965;
  assign n4967 = ~reg_controllable_hmaster2_out & ~n4966;
  assign n4968 = ~n4961 & ~n4967;
  assign n4969 = ~reg_controllable_hmaster1_out & ~n4968;
  assign n4970 = ~n4937 & ~n4969;
  assign n4971 = reg_stateG10_6_out & ~n4970;
  assign n4972 = next_sys_fair<0>_out  & ~n4452;
  assign n4973 = ~next_sys_fair<0>_out  & ~n4442;
  assign n4974 = ~n4972 & ~n4973;
  assign n4975 = next_sys_fair<3>_out  & ~n4974;
  assign n4976 = ~n4965 & ~n4975;
  assign n4977 = reg_controllable_hmaster2_out & ~n4976;
  assign n4978 = ~n4935 & ~n4977;
  assign n4979 = reg_controllable_hmaster1_out & ~n4978;
  assign n4980 = ~n4969 & ~n4979;
  assign n4981 = ~reg_stateG10_6_out & ~n4980;
  assign n4982 = ~n4971 & ~n4981;
  assign n4983 = reg_i_hlock6_out & ~n4982;
  assign n4984 = next_sys_fair<0>_out  & ~n4479;
  assign n4985 = ~next_sys_fair<0>_out  & ~n4470;
  assign n4986 = ~n4984 & ~n4985;
  assign n4987 = next_sys_fair<3>_out  & ~n4986;
  assign n4988 = next_sys_fair<0>_out  & ~n4548;
  assign n4989 = ~next_sys_fair<0>_out  & ~n4558;
  assign n4990 = ~n4988 & ~n4989;
  assign n4991 = ~next_sys_fair<3>_out  & ~n4990;
  assign n4992 = ~n4987 & ~n4991;
  assign n4993 = reg_controllable_hmaster2_out & ~n4992;
  assign n4994 = ~n4935 & ~n4993;
  assign n4995 = reg_controllable_hmaster1_out & ~n4994;
  assign n4996 = ~n4969 & ~n4995;
  assign n4997 = reg_stateG10_6_out & ~n4996;
  assign n4998 = next_sys_fair<0>_out  & ~n4483;
  assign n4999 = ~next_sys_fair<0>_out  & ~n4473;
  assign n5000 = ~n4998 & ~n4999;
  assign n5001 = next_sys_fair<3>_out  & ~n5000;
  assign n5002 = next_sys_fair<0>_out  & ~n4552;
  assign n5003 = ~next_sys_fair<0>_out  & ~n4561;
  assign n5004 = ~n5002 & ~n5003;
  assign n5005 = ~next_sys_fair<3>_out  & ~n5004;
  assign n5006 = ~n5001 & ~n5005;
  assign n5007 = reg_controllable_hmaster2_out & ~n5006;
  assign n5008 = ~n4935 & ~n5007;
  assign n5009 = reg_controllable_hmaster1_out & ~n5008;
  assign n5010 = ~n4969 & ~n5009;
  assign n5011 = ~reg_stateG10_6_out & ~n5010;
  assign n5012 = ~n4997 & ~n5011;
  assign n5013 = ~reg_i_hlock6_out & ~n5012;
  assign n5014 = ~n4983 & ~n5013;
  assign n5015 = ~next_sys_fair<1>_out  & ~n5014;
  assign n5016 = ~n4894 & ~n5015;
  assign n5017 = ~reg_controllable_hmaster0_out & ~n5016;
  assign n5018 = ~n4802 & ~n5017;
  assign n5019 = ~reg_controllable_hmaster3_out & ~n5018;
  assign n5020 = ~n4602 & ~n5019;
  assign n5021 = reg_stateG10_8_out & ~n5020;
  assign n5022 = ~n4866 & ~n4975;
  assign n5023 = ~reg_controllable_hmaster2_out & ~n5022;
  assign n5024 = ~n4435 & ~n5023;
  assign n5025 = ~reg_controllable_hmaster1_out & ~n5024;
  assign n5026 = ~n4434 & ~n5025;
  assign n5027 = next_sys_fair<1>_out  & ~n5026;
  assign n5028 = ~n4512 & ~n4967;
  assign n5029 = ~reg_controllable_hmaster1_out & ~n5028;
  assign n5030 = ~n4511 & ~n5029;
  assign n5031 = ~next_sys_fair<1>_out  & ~n5030;
  assign n5032 = ~n5027 & ~n5031;
  assign n5033 = ~reg_controllable_hmaster0_out & ~n5032;
  assign n5034 = ~n4576 & ~n5033;
  assign n5035 = reg_controllable_hmaster3_out & ~n5034;
  assign n5036 = ~n5019 & ~n5035;
  assign n5037 = ~reg_stateG10_8_out & ~n5036;
  assign n5038 = ~n5021 & ~n5037;
  assign n5039 = reg_stateG10_7_out & ~n5038;
  assign n5040 = ~n4619 & ~n4868;
  assign n5041 = reg_controllable_hmaster1_out & ~n5040;
  assign n5042 = ~n4695 & ~n5041;
  assign n5043 = next_sys_fair<1>_out  & ~n5042;
  assign n5044 = next_sys_fair<0>_out  & ~n4442;
  assign n5045 = ~next_sys_fair<0>_out  & ~n4452;
  assign n5046 = ~n5044 & ~n5045;
  assign n5047 = next_sys_fair<3>_out  & ~n5046;
  assign n5048 = ~n4965 & ~n5047;
  assign n5049 = reg_controllable_hmaster2_out & ~n5048;
  assign n5050 = ~n4742 & ~n5049;
  assign n5051 = reg_controllable_hmaster1_out & ~n5050;
  assign n5052 = ~n4798 & ~n5051;
  assign n5053 = ~next_sys_fair<1>_out  & ~n5052;
  assign n5054 = ~n5043 & ~n5053;
  assign n5055 = reg_controllable_hmaster0_out & ~n5054;
  assign n5056 = ~n5017 & ~n5055;
  assign n5057 = ~reg_controllable_hmaster3_out & ~n5056;
  assign n5058 = ~n4602 & ~n5057;
  assign n5059 = reg_stateG10_8_out & ~n5058;
  assign n5060 = ~n5035 & ~n5057;
  assign n5061 = ~reg_stateG10_8_out & ~n5060;
  assign n5062 = ~n5059 & ~n5061;
  assign n5063 = ~reg_stateG10_7_out & ~n5062;
  assign n5064 = ~n5039 & ~n5063;
  assign n5065 = ~reg_i_hready_out & ~n5064;
  assign n5066 = ~n4427 & ~n5065;
  assign n5067 = reg_i_hlock7_out & ~n5066;
  assign n5068 = next_sys_fair<1>_out  & ~n3553;
  assign n5069 = next_sys_fair<0>_out  & ~n3067;
  assign n5070 = ~next_sys_fair<0>_out  & ~n3103;
  assign n5071 = ~n5069 & ~n5070;
  assign n5072 = next_sys_fair<3>_out  & ~n5071;
  assign n5073 = ~n3592 & ~n5072;
  assign n5074 = reg_controllable_hmaster2_out & ~n5073;
  assign n5075 = ~n3384 & ~n5074;
  assign n5076 = reg_controllable_hmaster1_out & ~n5075;
  assign n5077 = ~n3387 & ~n5076;
  assign n5078 = ~next_sys_fair<1>_out  & ~n5077;
  assign n5079 = ~n5068 & ~n5078;
  assign n5080 = reg_controllable_hmaster0_out & ~n5079;
  assign n5081 = ~n3392 & ~n5080;
  assign n5082 = ~reg_controllable_hmaster3_out & ~n5081;
  assign n5083 = ~n3363 & ~n5082;
  assign n5084 = ~reg_controllable_hgrant6_out & ~n5083;
  assign n5085 = ~reg_controllable_hgrant6_out & ~n5084;
  assign n5086 = reg_stateG10_7_out & ~n5085;
  assign n5087 = next_sys_fair<1>_out  & ~n3561;
  assign n5088 = next_sys_fair<0>_out  & ~n3081;
  assign n5089 = ~next_sys_fair<0>_out  & ~n3120;
  assign n5090 = ~n5088 & ~n5089;
  assign n5091 = next_sys_fair<3>_out  & ~n5090;
  assign n5092 = ~n3606 & ~n5091;
  assign n5093 = reg_controllable_hmaster2_out & ~n5092;
  assign n5094 = ~n3384 & ~n5093;
  assign n5095 = reg_controllable_hmaster1_out & ~n5094;
  assign n5096 = ~n3387 & ~n5095;
  assign n5097 = ~next_sys_fair<1>_out  & ~n5096;
  assign n5098 = ~n5087 & ~n5097;
  assign n5099 = reg_controllable_hmaster0_out & ~n5098;
  assign n5100 = ~n3392 & ~n5099;
  assign n5101 = ~reg_controllable_hmaster3_out & ~n5100;
  assign n5102 = ~n3363 & ~n5101;
  assign n5103 = ~reg_controllable_hgrant6_out & ~n5102;
  assign n5104 = ~reg_controllable_hgrant6_out & ~n5103;
  assign n5105 = ~reg_stateG10_7_out & ~n5104;
  assign n5106 = ~n5086 & ~n5105;
  assign n5107 = ~reg_controllable_hgrant8_out & ~n5106;
  assign n5108 = ~reg_controllable_hgrant8_out & ~n5107;
  assign n5109 = reg_controllable_hgrant7_out & ~n5108;
  assign n5110 = ~n4381 & ~n5109;
  assign n5111 = ~reg_controllable_hgrant9_out & ~n5110;
  assign n5112 = ~n3357 & ~n5111;
  assign n5113 = reg_controllable_nhgrant0_out & ~n5112;
  assign n5114 = ~n4425 & ~n5113;
  assign n5115 = reg_i_hready_out & ~n5114;
  assign n5116 = ~n4619 & ~n4878;
  assign n5117 = reg_controllable_hmaster1_out & ~n5116;
  assign n5118 = ~n4695 & ~n5117;
  assign n5119 = next_sys_fair<1>_out  & ~n5118;
  assign n5120 = next_sys_fair<0>_out  & ~n4470;
  assign n5121 = ~next_sys_fair<0>_out  & ~n4479;
  assign n5122 = ~n5120 & ~n5121;
  assign n5123 = next_sys_fair<3>_out  & ~n5122;
  assign n5124 = ~n4991 & ~n5123;
  assign n5125 = reg_controllable_hmaster2_out & ~n5124;
  assign n5126 = ~n4742 & ~n5125;
  assign n5127 = reg_controllable_hmaster1_out & ~n5126;
  assign n5128 = ~n4798 & ~n5127;
  assign n5129 = ~next_sys_fair<1>_out  & ~n5128;
  assign n5130 = ~n5119 & ~n5129;
  assign n5131 = reg_controllable_hmaster0_out & ~n5130;
  assign n5132 = ~n5017 & ~n5131;
  assign n5133 = ~reg_controllable_hmaster3_out & ~n5132;
  assign n5134 = ~n4602 & ~n5133;
  assign n5135 = reg_stateG10_8_out & ~n5134;
  assign n5136 = ~n5035 & ~n5133;
  assign n5137 = ~reg_stateG10_8_out & ~n5136;
  assign n5138 = ~n5135 & ~n5137;
  assign n5139 = reg_stateG10_7_out & ~n5138;
  assign n5140 = ~n4619 & ~n4886;
  assign n5141 = reg_controllable_hmaster1_out & ~n5140;
  assign n5142 = ~n4695 & ~n5141;
  assign n5143 = next_sys_fair<1>_out  & ~n5142;
  assign n5144 = next_sys_fair<0>_out  & ~n4473;
  assign n5145 = ~next_sys_fair<0>_out  & ~n4483;
  assign n5146 = ~n5144 & ~n5145;
  assign n5147 = next_sys_fair<3>_out  & ~n5146;
  assign n5148 = ~n5005 & ~n5147;
  assign n5149 = reg_controllable_hmaster2_out & ~n5148;
  assign n5150 = ~n4742 & ~n5149;
  assign n5151 = reg_controllable_hmaster1_out & ~n5150;
  assign n5152 = ~n4798 & ~n5151;
  assign n5153 = ~next_sys_fair<1>_out  & ~n5152;
  assign n5154 = ~n5143 & ~n5153;
  assign n5155 = reg_controllable_hmaster0_out & ~n5154;
  assign n5156 = ~n5017 & ~n5155;
  assign n5157 = ~reg_controllable_hmaster3_out & ~n5156;
  assign n5158 = ~n4602 & ~n5157;
  assign n5159 = reg_stateG10_8_out & ~n5158;
  assign n5160 = ~n5035 & ~n5157;
  assign n5161 = ~reg_stateG10_8_out & ~n5160;
  assign n5162 = ~n5159 & ~n5161;
  assign n5163 = ~reg_stateG10_7_out & ~n5162;
  assign n5164 = ~n5139 & ~n5163;
  assign n5165 = ~reg_i_hready_out & ~n5164;
  assign n5166 = ~n5115 & ~n5165;
  assign n5167 = ~reg_i_hlock7_out & ~n5166;
  assign n5168 = ~n5067 & ~n5167;
  assign n5169 = reg_i_hlock8_out & ~n5168;
  assign n5170 = ~n3548 & ~n3588;
  assign n5171 = ~reg_controllable_hmaster2_out & ~n5170;
  assign n5172 = ~n3460 & ~n5171;
  assign n5173 = ~reg_controllable_hmaster1_out & ~n5172;
  assign n5174 = ~n3459 & ~n5173;
  assign n5175 = next_sys_fair<1>_out  & ~n5174;
  assign n5176 = ~n3547 & ~n3592;
  assign n5177 = ~reg_controllable_hmaster2_out & ~n5176;
  assign n5178 = ~n3253 & ~n5177;
  assign n5179 = ~reg_controllable_hmaster1_out & ~n5178;
  assign n5180 = ~n3252 & ~n5179;
  assign n5181 = ~next_sys_fair<1>_out  & ~n5180;
  assign n5182 = ~n5175 & ~n5181;
  assign n5183 = ~reg_controllable_hmaster0_out & ~n5182;
  assign n5184 = ~n3458 & ~n5183;
  assign n5185 = reg_controllable_hmaster3_out & ~n5184;
  assign n5186 = ~n3481 & ~n5185;
  assign n5187 = reg_stateG10_8_out & ~n5186;
  assign n5188 = ~n3556 & ~n3602;
  assign n5189 = ~reg_controllable_hmaster2_out & ~n5188;
  assign n5190 = ~n3460 & ~n5189;
  assign n5191 = ~reg_controllable_hmaster1_out & ~n5190;
  assign n5192 = ~n3459 & ~n5191;
  assign n5193 = next_sys_fair<1>_out  & ~n5192;
  assign n5194 = ~n3555 & ~n3606;
  assign n5195 = ~reg_controllable_hmaster2_out & ~n5194;
  assign n5196 = ~n3253 & ~n5195;
  assign n5197 = ~reg_controllable_hmaster1_out & ~n5196;
  assign n5198 = ~n3252 & ~n5197;
  assign n5199 = ~next_sys_fair<1>_out  & ~n5198;
  assign n5200 = ~n5193 & ~n5199;
  assign n5201 = ~reg_controllable_hmaster0_out & ~n5200;
  assign n5202 = ~n3458 & ~n5201;
  assign n5203 = reg_controllable_hmaster3_out & ~n5202;
  assign n5204 = ~n3481 & ~n5203;
  assign n5205 = ~reg_stateG10_8_out & ~n5204;
  assign n5206 = ~n5187 & ~n5205;
  assign n5207 = ~reg_controllable_hgrant6_out & ~n5206;
  assign n5208 = ~reg_controllable_hgrant6_out & ~n5207;
  assign n5209 = reg_controllable_hgrant8_out & ~n5208;
  assign n5210 = ~n4379 & ~n5209;
  assign n5211 = ~reg_controllable_hgrant7_out & ~n5210;
  assign n5212 = ~n3449 & ~n5211;
  assign n5213 = ~reg_controllable_hgrant9_out & ~n5212;
  assign n5214 = ~n3357 & ~n5213;
  assign n5215 = reg_controllable_nhgrant0_out & ~n5214;
  assign n5216 = ~n4425 & ~n5215;
  assign n5217 = reg_i_hready_out & ~n5216;
  assign n5218 = ~n4876 & ~n4987;
  assign n5219 = ~reg_controllable_hmaster2_out & ~n5218;
  assign n5220 = ~n4435 & ~n5219;
  assign n5221 = ~reg_controllable_hmaster1_out & ~n5220;
  assign n5222 = ~n4434 & ~n5221;
  assign n5223 = next_sys_fair<1>_out  & ~n5222;
  assign n5224 = ~n4875 & ~n4991;
  assign n5225 = ~reg_controllable_hmaster2_out & ~n5224;
  assign n5226 = ~n4512 & ~n5225;
  assign n5227 = ~reg_controllable_hmaster1_out & ~n5226;
  assign n5228 = ~n4511 & ~n5227;
  assign n5229 = ~next_sys_fair<1>_out  & ~n5228;
  assign n5230 = ~n5223 & ~n5229;
  assign n5231 = ~reg_controllable_hmaster0_out & ~n5230;
  assign n5232 = ~n4576 & ~n5231;
  assign n5233 = reg_controllable_hmaster3_out & ~n5232;
  assign n5234 = ~n5019 & ~n5233;
  assign n5235 = reg_stateG10_8_out & ~n5234;
  assign n5236 = ~n4884 & ~n5001;
  assign n5237 = ~reg_controllable_hmaster2_out & ~n5236;
  assign n5238 = ~n4435 & ~n5237;
  assign n5239 = ~reg_controllable_hmaster1_out & ~n5238;
  assign n5240 = ~n4434 & ~n5239;
  assign n5241 = next_sys_fair<1>_out  & ~n5240;
  assign n5242 = ~n4883 & ~n5005;
  assign n5243 = ~reg_controllable_hmaster2_out & ~n5242;
  assign n5244 = ~n4512 & ~n5243;
  assign n5245 = ~reg_controllable_hmaster1_out & ~n5244;
  assign n5246 = ~n4511 & ~n5245;
  assign n5247 = ~next_sys_fair<1>_out  & ~n5246;
  assign n5248 = ~n5241 & ~n5247;
  assign n5249 = ~reg_controllable_hmaster0_out & ~n5248;
  assign n5250 = ~n4576 & ~n5249;
  assign n5251 = reg_controllable_hmaster3_out & ~n5250;
  assign n5252 = ~n5019 & ~n5251;
  assign n5253 = ~reg_stateG10_8_out & ~n5252;
  assign n5254 = ~n5235 & ~n5253;
  assign n5255 = reg_stateG10_7_out & ~n5254;
  assign n5256 = ~n5057 & ~n5233;
  assign n5257 = reg_stateG10_8_out & ~n5256;
  assign n5258 = ~n5057 & ~n5251;
  assign n5259 = ~reg_stateG10_8_out & ~n5258;
  assign n5260 = ~n5257 & ~n5259;
  assign n5261 = ~reg_stateG10_7_out & ~n5260;
  assign n5262 = ~n5255 & ~n5261;
  assign n5263 = ~reg_i_hready_out & ~n5262;
  assign n5264 = ~n5217 & ~n5263;
  assign n5265 = reg_i_hlock7_out & ~n5264;
  assign n5266 = ~n5109 & ~n5211;
  assign n5267 = ~reg_controllable_hgrant9_out & ~n5266;
  assign n5268 = ~n3357 & ~n5267;
  assign n5269 = reg_controllable_nhgrant0_out & ~n5268;
  assign n5270 = ~n4425 & ~n5269;
  assign n5271 = reg_i_hready_out & ~n5270;
  assign n5272 = ~n5133 & ~n5233;
  assign n5273 = reg_stateG10_8_out & ~n5272;
  assign n5274 = ~n5133 & ~n5251;
  assign n5275 = ~reg_stateG10_8_out & ~n5274;
  assign n5276 = ~n5273 & ~n5275;
  assign n5277 = reg_stateG10_7_out & ~n5276;
  assign n5278 = ~n5157 & ~n5233;
  assign n5279 = reg_stateG10_8_out & ~n5278;
  assign n5280 = ~n5157 & ~n5251;
  assign n5281 = ~reg_stateG10_8_out & ~n5280;
  assign n5282 = ~n5279 & ~n5281;
  assign n5283 = ~reg_stateG10_7_out & ~n5282;
  assign n5284 = ~n5277 & ~n5283;
  assign n5285 = ~reg_i_hready_out & ~n5284;
  assign n5286 = ~n5271 & ~n5285;
  assign n5287 = ~reg_i_hlock7_out & ~n5286;
  assign n5288 = ~n5265 & ~n5287;
  assign n5289 = ~reg_i_hlock8_out & ~n5288;
  assign n5290 = ~n5169 & ~n5289;
  assign n5291 = reg_i_hlock0_out & ~n5290;
  assign n5292 = next_sys_fair<0>_out  & ~n2922;
  assign n5293 = ~next_sys_fair<0>_out  & ~n3152;
  assign n5294 = ~n5292 & ~n5293;
  assign n5295 = ~next_sys_fair<3>_out  & ~n5294;
  assign n5296 = ~n3249 & ~n5295;
  assign n5297 = next_sys_fair<1>_out  & ~n5296;
  assign n5298 = ~n3456 & ~n5297;
  assign n5299 = reg_controllable_hmaster3_out & ~n5298;
  assign n5300 = reg_controllable_hmaster0_out & ~n5298;
  assign n5301 = reg_controllable_hmaster1_out & ~n5296;
  assign n5302 = reg_controllable_hmaster2_out & ~n5296;
  assign n5303 = next_sys_fair<0>_out  & ~n3134;
  assign n5304 = ~n3076 & ~n3275;
  assign n5305 = ~reg_controllable_hgrant4_out & ~n5304;
  assign n5306 = ~reg_controllable_hgrant4_out & ~n5305;
  assign n5307 = ~reg_controllable_hgrant5_out & ~n5306;
  assign n5308 = ~reg_controllable_hgrant5_out & ~n5307;
  assign n5309 = ~next_sys_fair<0>_out  & ~n5308;
  assign n5310 = ~n5303 & ~n5309;
  assign n5311 = ~next_sys_fair<3>_out  & ~n5310;
  assign n5312 = ~n3555 & ~n5311;
  assign n5313 = ~reg_controllable_hmaster2_out & ~n5312;
  assign n5314 = ~n5302 & ~n5313;
  assign n5315 = ~reg_controllable_hmaster1_out & ~n5314;
  assign n5316 = ~n5301 & ~n5315;
  assign n5317 = next_sys_fair<1>_out  & ~n5316;
  assign n5318 = ~n5199 & ~n5317;
  assign n5319 = ~reg_controllable_hmaster0_out & ~n5318;
  assign n5320 = ~n5300 & ~n5319;
  assign n5321 = ~reg_controllable_hmaster3_out & ~n5320;
  assign n5322 = ~n5299 & ~n5321;
  assign n5323 = ~reg_controllable_hgrant6_out & ~n5322;
  assign n5324 = ~reg_controllable_hgrant6_out & ~n5323;
  assign n5325 = ~reg_controllable_hgrant8_out & ~n5324;
  assign n5326 = ~reg_controllable_hgrant8_out & ~n5325;
  assign n5327 = ~reg_controllable_hgrant7_out & ~n5326;
  assign n5328 = ~reg_controllable_hgrant7_out & ~n5327;
  assign n5329 = ~reg_controllable_hgrant9_out & ~n5328;
  assign n5330 = ~reg_controllable_hgrant9_out & ~n5329;
  assign n5331 = ~reg_controllable_nhgrant0_out & ~n5330;
  assign n5332 = ~n4385 & ~n5331;
  assign n5333 = reg_i_hready_out & ~n5332;
  assign n5334 = next_sys_fair<0>_out  & ~n4481;
  assign n5335 = ~n4472 & ~n4550;
  assign n5336 = ~next_sys_fair<0>_out  & ~n5335;
  assign n5337 = ~n5334 & ~n5336;
  assign n5338 = ~next_sys_fair<3>_out  & ~n5337;
  assign n5339 = ~n4883 & ~n5338;
  assign n5340 = ~reg_controllable_hmaster2_out & ~n5339;
  assign n5341 = ~n4853 & ~n5340;
  assign n5342 = ~reg_controllable_hmaster1_out & ~n5341;
  assign n5343 = ~n4819 & ~n5342;
  assign n5344 = reg_stateG10_6_out & ~n5343;
  assign n5345 = ~n4870 & ~n5342;
  assign n5346 = ~reg_stateG10_6_out & ~n5345;
  assign n5347 = ~n5344 & ~n5346;
  assign n5348 = reg_i_hlock6_out & ~n5347;
  assign n5349 = ~n4880 & ~n5342;
  assign n5350 = reg_stateG10_6_out & ~n5349;
  assign n5351 = ~n4888 & ~n5342;
  assign n5352 = ~reg_stateG10_6_out & ~n5351;
  assign n5353 = ~n5350 & ~n5352;
  assign n5354 = ~reg_i_hlock6_out & ~n5353;
  assign n5355 = ~n5348 & ~n5354;
  assign n5356 = next_sys_fair<1>_out  & ~n5355;
  assign n5357 = ~n4961 & ~n5243;
  assign n5358 = ~reg_controllable_hmaster1_out & ~n5357;
  assign n5359 = ~n4937 & ~n5358;
  assign n5360 = reg_stateG10_6_out & ~n5359;
  assign n5361 = ~n4979 & ~n5358;
  assign n5362 = ~reg_stateG10_6_out & ~n5361;
  assign n5363 = ~n5360 & ~n5362;
  assign n5364 = reg_i_hlock6_out & ~n5363;
  assign n5365 = ~n4995 & ~n5358;
  assign n5366 = reg_stateG10_6_out & ~n5365;
  assign n5367 = ~n5009 & ~n5358;
  assign n5368 = ~reg_stateG10_6_out & ~n5367;
  assign n5369 = ~n5366 & ~n5368;
  assign n5370 = ~reg_i_hlock6_out & ~n5369;
  assign n5371 = ~n5364 & ~n5370;
  assign n5372 = ~next_sys_fair<1>_out  & ~n5371;
  assign n5373 = ~n5356 & ~n5372;
  assign n5374 = ~reg_controllable_hmaster0_out & ~n5373;
  assign n5375 = ~n4802 & ~n5374;
  assign n5376 = ~reg_controllable_hmaster3_out & ~n5375;
  assign n5377 = ~n4602 & ~n5376;
  assign n5378 = reg_stateG10_8_out & ~n5377;
  assign n5379 = ~n5035 & ~n5376;
  assign n5380 = ~reg_stateG10_8_out & ~n5379;
  assign n5381 = ~n5378 & ~n5380;
  assign n5382 = reg_stateG10_7_out & ~n5381;
  assign n5383 = ~n5055 & ~n5374;
  assign n5384 = ~reg_controllable_hmaster3_out & ~n5383;
  assign n5385 = ~n4602 & ~n5384;
  assign n5386 = reg_stateG10_8_out & ~n5385;
  assign n5387 = ~n5035 & ~n5384;
  assign n5388 = ~reg_stateG10_8_out & ~n5387;
  assign n5389 = ~n5386 & ~n5388;
  assign n5390 = ~reg_stateG10_7_out & ~n5389;
  assign n5391 = ~n5382 & ~n5390;
  assign n5392 = ~reg_i_hready_out & ~n5391;
  assign n5393 = ~n5333 & ~n5392;
  assign n5394 = reg_i_hlock7_out & ~n5393;
  assign n5395 = ~n5113 & ~n5331;
  assign n5396 = reg_i_hready_out & ~n5395;
  assign n5397 = ~n5131 & ~n5374;
  assign n5398 = ~reg_controllable_hmaster3_out & ~n5397;
  assign n5399 = ~n4602 & ~n5398;
  assign n5400 = reg_stateG10_8_out & ~n5399;
  assign n5401 = ~n5035 & ~n5398;
  assign n5402 = ~reg_stateG10_8_out & ~n5401;
  assign n5403 = ~n5400 & ~n5402;
  assign n5404 = reg_stateG10_7_out & ~n5403;
  assign n5405 = ~n5155 & ~n5374;
  assign n5406 = ~reg_controllable_hmaster3_out & ~n5405;
  assign n5407 = ~n4602 & ~n5406;
  assign n5408 = reg_stateG10_8_out & ~n5407;
  assign n5409 = ~n5035 & ~n5406;
  assign n5410 = ~reg_stateG10_8_out & ~n5409;
  assign n5411 = ~n5408 & ~n5410;
  assign n5412 = ~reg_stateG10_7_out & ~n5411;
  assign n5413 = ~n5404 & ~n5412;
  assign n5414 = ~reg_i_hready_out & ~n5413;
  assign n5415 = ~n5396 & ~n5414;
  assign n5416 = ~reg_i_hlock7_out & ~n5415;
  assign n5417 = ~n5394 & ~n5416;
  assign n5418 = reg_i_hlock8_out & ~n5417;
  assign n5419 = ~n5215 & ~n5331;
  assign n5420 = reg_i_hready_out & ~n5419;
  assign n5421 = ~n5233 & ~n5376;
  assign n5422 = reg_stateG10_8_out & ~n5421;
  assign n5423 = ~n5251 & ~n5376;
  assign n5424 = ~reg_stateG10_8_out & ~n5423;
  assign n5425 = ~n5422 & ~n5424;
  assign n5426 = reg_stateG10_7_out & ~n5425;
  assign n5427 = ~n5233 & ~n5384;
  assign n5428 = reg_stateG10_8_out & ~n5427;
  assign n5429 = ~n5251 & ~n5384;
  assign n5430 = ~reg_stateG10_8_out & ~n5429;
  assign n5431 = ~n5428 & ~n5430;
  assign n5432 = ~reg_stateG10_7_out & ~n5431;
  assign n5433 = ~n5426 & ~n5432;
  assign n5434 = ~reg_i_hready_out & ~n5433;
  assign n5435 = ~n5420 & ~n5434;
  assign n5436 = reg_i_hlock7_out & ~n5435;
  assign n5437 = ~n5269 & ~n5331;
  assign n5438 = reg_i_hready_out & ~n5437;
  assign n5439 = ~n5233 & ~n5398;
  assign n5440 = reg_stateG10_8_out & ~n5439;
  assign n5441 = ~n5251 & ~n5398;
  assign n5442 = ~reg_stateG10_8_out & ~n5441;
  assign n5443 = ~n5440 & ~n5442;
  assign n5444 = reg_stateG10_7_out & ~n5443;
  assign n5445 = ~n5233 & ~n5406;
  assign n5446 = reg_stateG10_8_out & ~n5445;
  assign n5447 = ~n5251 & ~n5406;
  assign n5448 = ~reg_stateG10_8_out & ~n5447;
  assign n5449 = ~n5446 & ~n5448;
  assign n5450 = ~reg_stateG10_7_out & ~n5449;
  assign n5451 = ~n5444 & ~n5450;
  assign n5452 = ~reg_i_hready_out & ~n5451;
  assign n5453 = ~n5438 & ~n5452;
  assign n5454 = ~reg_i_hlock7_out & ~n5453;
  assign n5455 = ~n5436 & ~n5454;
  assign n5456 = ~reg_i_hlock8_out & ~n5455;
  assign n5457 = ~n5418 & ~n5456;
  assign n5458 = ~reg_i_hlock0_out & ~n5457;
  assign n5459 = ~n5291 & ~n5458;
  assign n5460 = reg_i_hbusreq9_out & ~n5459;
  assign n5461 = reg_i_hbusreq0_out & ~n5459;
  assign n5462 = reg_i_hbusreq5_out & ~n5459;
  assign n5463 = reg_i_hbusreq6_out & ~n5459;
  assign n5464 = reg_i_hbusreq7_out & ~n5459;
  assign n5465 = reg_i_hbusreq8_out & ~n5459;
  assign n5466 = reg_i_hbusreq3_out & ~n5459;
  assign n5467 = reg_i_hbusreq4_out & ~n5459;
  assign n5468 = reg_i_hbusreq2_out & ~n5459;
  assign n5469 = reg_i_hbusreq1_out & ~n5459;
  assign n5470 = ~reg_controllable_locked_out & ~n123;
  assign n5471 = ~reg_controllable_locked_out & ~n5470;
  assign n5472 = ~reg_controllable_hgrant2_out & ~n5471;
  assign n5473 = ~reg_controllable_hgrant2_out & ~n5472;
  assign n5474 = ~reg_controllable_hgrant1_out & ~n5473;
  assign n5475 = ~reg_controllable_hgrant1_out & ~n5474;
  assign n5476 = ~reg_controllable_hgrant3_out & ~n5475;
  assign n5477 = ~reg_controllable_hgrant3_out & ~n5476;
  assign n5478 = ~next_sys_fair<2>_out  & ~n5477;
  assign n5479 = ~next_sys_fair<2>_out  & ~n5478;
  assign n5480 = ~reg_controllable_hgrant4_out & ~n5479;
  assign n5481 = ~reg_controllable_hgrant4_out & ~n5480;
  assign n5482 = ~reg_controllable_hgrant5_out & ~n5481;
  assign n5483 = ~reg_controllable_hgrant5_out & ~n5482;
  assign n5484 = next_sys_fair<0>_out  & ~n5483;
  assign n5485 = ~next_env_fair_out & ~n151;
  assign n5486 = ~next_env_fair_out & ~n5485;
  assign n5487 = ~reg_stateG2_out & ~n5486;
  assign n5488 = ~reg_stateG2_out & ~n5487;
  assign n5489 = ~reg_stateA1_out & ~n5488;
  assign n5490 = ~reg_stateA1_out & ~n5489;
  assign n5491 = ~reg_controllable_locked_out & ~n5490;
  assign n5492 = ~reg_controllable_locked_out & ~n5491;
  assign n5493 = ~reg_controllable_hgrant2_out & ~n5492;
  assign n5494 = ~reg_controllable_hgrant2_out & ~n5493;
  assign n5495 = ~reg_controllable_hgrant1_out & ~n5494;
  assign n5496 = ~reg_controllable_hgrant1_out & ~n5495;
  assign n5497 = ~reg_controllable_hgrant3_out & ~n5496;
  assign n5498 = ~reg_controllable_hgrant3_out & ~n5497;
  assign n5499 = ~next_sys_fair<2>_out  & ~n5498;
  assign n5500 = ~next_sys_fair<2>_out  & ~n5499;
  assign n5501 = ~reg_controllable_hgrant4_out & ~n5500;
  assign n5502 = ~reg_controllable_hgrant4_out & ~n5501;
  assign n5503 = ~reg_controllable_hgrant5_out & ~n5502;
  assign n5504 = ~reg_controllable_hgrant5_out & ~n5503;
  assign n5505 = ~next_sys_fair<0>_out  & ~n5504;
  assign n5506 = ~n5484 & ~n5505;
  assign n5507 = next_sys_fair<3>_out  & ~n5506;
  assign n5508 = ~reg_controllable_hgrant4_out & ~n5498;
  assign n5509 = ~reg_controllable_hgrant4_out & ~n5508;
  assign n5510 = ~reg_controllable_hgrant5_out & ~n5509;
  assign n5511 = ~reg_controllable_hgrant5_out & ~n5510;
  assign n5512 = next_sys_fair<0>_out  & ~n5511;
  assign n5513 = next_sys_fair<2>_out  & ~n5498;
  assign n5514 = ~reg_stateA1_out & ~n3663;
  assign n5515 = ~reg_controllable_locked_out & ~n5514;
  assign n5516 = ~reg_controllable_locked_out & ~n5515;
  assign n5517 = ~reg_controllable_hgrant2_out & ~n5516;
  assign n5518 = ~reg_controllable_hgrant2_out & ~n5517;
  assign n5519 = ~reg_controllable_hgrant1_out & ~n5518;
  assign n5520 = ~reg_controllable_hgrant1_out & ~n5519;
  assign n5521 = ~reg_controllable_hgrant3_out & ~n5520;
  assign n5522 = ~reg_controllable_hgrant3_out & ~n5521;
  assign n5523 = ~next_sys_fair<2>_out  & ~n5522;
  assign n5524 = ~n5513 & ~n5523;
  assign n5525 = ~reg_controllable_hgrant4_out & ~n5524;
  assign n5526 = ~reg_controllable_hgrant4_out & ~n5525;
  assign n5527 = ~reg_controllable_hgrant5_out & ~n5526;
  assign n5528 = ~reg_controllable_hgrant5_out & ~n5527;
  assign n5529 = ~next_sys_fair<0>_out  & ~n5528;
  assign n5530 = ~n5512 & ~n5529;
  assign n5531 = ~next_sys_fair<3>_out  & ~n5530;
  assign n5532 = ~n5507 & ~n5531;
  assign n5533 = reg_controllable_hmaster1_out & ~n5532;
  assign n5534 = reg_controllable_hmaster2_out & ~n5532;
  assign n5535 = reg_controllable_hmastlock_out & ~n123;
  assign n5536 = ~n1293 & ~n5535;
  assign n5537 = ~reg_controllable_locked_out & ~n5536;
  assign n5538 = ~reg_controllable_locked_out & ~n5537;
  assign n5539 = ~reg_controllable_hgrant2_out & ~n5538;
  assign n5540 = ~reg_controllable_hgrant2_out & ~n5539;
  assign n5541 = ~reg_controllable_hgrant1_out & ~n5540;
  assign n5542 = ~reg_controllable_hgrant1_out & ~n5541;
  assign n5543 = ~reg_controllable_hgrant3_out & ~n5542;
  assign n5544 = ~reg_controllable_hgrant3_out & ~n5543;
  assign n5545 = ~next_sys_fair<2>_out  & ~n5544;
  assign n5546 = ~next_sys_fair<2>_out  & ~n5545;
  assign n5547 = ~reg_controllable_hgrant4_out & ~n5546;
  assign n5548 = ~reg_controllable_hgrant4_out & ~n5547;
  assign n5549 = ~reg_controllable_hgrant5_out & ~n5548;
  assign n5550 = ~reg_controllable_hgrant5_out & ~n5549;
  assign n5551 = next_sys_fair<0>_out  & ~n5550;
  assign n5552 = reg_controllable_hmastlock_out & ~n5490;
  assign n5553 = ~n1319 & ~n5552;
  assign n5554 = ~reg_controllable_locked_out & ~n5553;
  assign n5555 = ~reg_controllable_locked_out & ~n5554;
  assign n5556 = ~reg_controllable_hgrant2_out & ~n5555;
  assign n5557 = ~reg_controllable_hgrant2_out & ~n5556;
  assign n5558 = ~reg_controllable_hgrant1_out & ~n5557;
  assign n5559 = ~reg_controllable_hgrant1_out & ~n5558;
  assign n5560 = ~reg_controllable_hgrant3_out & ~n5559;
  assign n5561 = ~reg_controllable_hgrant3_out & ~n5560;
  assign n5562 = ~next_sys_fair<2>_out  & ~n5561;
  assign n5563 = ~next_sys_fair<2>_out  & ~n5562;
  assign n5564 = ~reg_controllable_hgrant4_out & ~n5563;
  assign n5565 = ~reg_controllable_hgrant4_out & ~n5564;
  assign n5566 = ~reg_controllable_hgrant5_out & ~n5565;
  assign n5567 = ~reg_controllable_hgrant5_out & ~n5566;
  assign n5568 = ~next_sys_fair<0>_out  & ~n5567;
  assign n5569 = ~n5551 & ~n5568;
  assign n5570 = next_sys_fair<3>_out  & ~n5569;
  assign n5571 = ~reg_controllable_hgrant4_out & ~n5561;
  assign n5572 = ~reg_controllable_hgrant4_out & ~n5571;
  assign n5573 = ~reg_controllable_hgrant5_out & ~n5572;
  assign n5574 = ~reg_controllable_hgrant5_out & ~n5573;
  assign n5575 = next_sys_fair<0>_out  & ~n5574;
  assign n5576 = next_sys_fair<2>_out  & ~n5561;
  assign n5577 = reg_controllable_hmastlock_out & ~n5514;
  assign n5578 = ~n1480 & ~n5577;
  assign n5579 = ~reg_controllable_locked_out & ~n5578;
  assign n5580 = ~reg_controllable_locked_out & ~n5579;
  assign n5581 = ~reg_controllable_hgrant2_out & ~n5580;
  assign n5582 = ~reg_controllable_hgrant2_out & ~n5581;
  assign n5583 = ~reg_controllable_hgrant1_out & ~n5582;
  assign n5584 = ~reg_controllable_hgrant1_out & ~n5583;
  assign n5585 = ~reg_controllable_hgrant3_out & ~n5584;
  assign n5586 = ~reg_controllable_hgrant3_out & ~n5585;
  assign n5587 = ~next_sys_fair<2>_out  & ~n5586;
  assign n5588 = ~n5576 & ~n5587;
  assign n5589 = ~reg_controllable_hgrant4_out & ~n5588;
  assign n5590 = ~reg_controllable_hgrant4_out & ~n5589;
  assign n5591 = ~reg_controllable_hgrant5_out & ~n5590;
  assign n5592 = ~reg_controllable_hgrant5_out & ~n5591;
  assign n5593 = ~next_sys_fair<0>_out  & ~n5592;
  assign n5594 = ~n5575 & ~n5593;
  assign n5595 = ~next_sys_fair<3>_out  & ~n5594;
  assign n5596 = ~n5570 & ~n5595;
  assign n5597 = ~reg_controllable_hmaster2_out & ~n5596;
  assign n5598 = ~n5534 & ~n5597;
  assign n5599 = ~reg_controllable_hmaster1_out & ~n5598;
  assign n5600 = ~n5533 & ~n5599;
  assign n5601 = next_sys_fair<1>_out  & ~n5600;
  assign n5602 = next_sys_fair<3>_out  & ~n5504;
  assign n5603 = ~n5478 & ~n5513;
  assign n5604 = ~reg_controllable_hgrant4_out & ~n5603;
  assign n5605 = ~reg_controllable_hgrant4_out & ~n5604;
  assign n5606 = ~reg_controllable_hgrant5_out & ~n5605;
  assign n5607 = ~reg_controllable_hgrant5_out & ~n5606;
  assign n5608 = ~next_sys_fair<3>_out  & ~n5607;
  assign n5609 = ~n5602 & ~n5608;
  assign n5610 = reg_controllable_hmaster1_out & ~n5609;
  assign n5611 = reg_controllable_hmaster2_out & ~n5609;
  assign n5612 = next_sys_fair<3>_out  & ~n5567;
  assign n5613 = ~n1424 & ~n5535;
  assign n5614 = ~reg_controllable_locked_out & ~n5613;
  assign n5615 = ~reg_controllable_locked_out & ~n5614;
  assign n5616 = ~reg_controllable_hgrant2_out & ~n5615;
  assign n5617 = ~reg_controllable_hgrant2_out & ~n5616;
  assign n5618 = ~reg_controllable_hgrant1_out & ~n5617;
  assign n5619 = ~reg_controllable_hgrant1_out & ~n5618;
  assign n5620 = ~reg_controllable_hgrant3_out & ~n5619;
  assign n5621 = ~reg_controllable_hgrant3_out & ~n5620;
  assign n5622 = ~next_sys_fair<2>_out  & ~n5621;
  assign n5623 = ~n5576 & ~n5622;
  assign n5624 = ~reg_controllable_hgrant4_out & ~n5623;
  assign n5625 = ~reg_controllable_hgrant4_out & ~n5624;
  assign n5626 = ~reg_controllable_hgrant5_out & ~n5625;
  assign n5627 = ~reg_controllable_hgrant5_out & ~n5626;
  assign n5628 = next_sys_fair<0>_out  & ~n5627;
  assign n5629 = ~n5545 & ~n5576;
  assign n5630 = ~reg_controllable_hgrant4_out & ~n5629;
  assign n5631 = ~reg_controllable_hgrant4_out & ~n5630;
  assign n5632 = ~reg_controllable_hgrant5_out & ~n5631;
  assign n5633 = ~reg_controllable_hgrant5_out & ~n5632;
  assign n5634 = ~next_sys_fair<0>_out  & ~n5633;
  assign n5635 = ~n5628 & ~n5634;
  assign n5636 = ~next_sys_fair<3>_out  & ~n5635;
  assign n5637 = ~n5612 & ~n5636;
  assign n5638 = ~reg_controllable_hmaster2_out & ~n5637;
  assign n5639 = ~n5611 & ~n5638;
  assign n5640 = ~reg_controllable_hmaster1_out & ~n5639;
  assign n5641 = ~n5610 & ~n5640;
  assign n5642 = ~next_sys_fair<1>_out  & ~n5641;
  assign n5643 = ~n5601 & ~n5642;
  assign n5644 = reg_controllable_hmaster0_out & ~n5643;
  assign n5645 = next_sys_fair<1>_out  & ~n5532;
  assign n5646 = ~next_sys_fair<1>_out  & ~n5609;
  assign n5647 = ~n5645 & ~n5646;
  assign n5648 = ~reg_controllable_hmaster0_out & ~n5647;
  assign n5649 = ~n5644 & ~n5648;
  assign n5650 = reg_controllable_hmaster3_out & ~n5649;
  assign n5651 = ~reg_controllable_hmaster3_out & ~n5647;
  assign n5652 = ~n5650 & ~n5651;
  assign n5653 = ~reg_controllable_hgrant6_out & ~n5652;
  assign n5654 = ~reg_controllable_hgrant6_out & ~n5653;
  assign n5655 = ~reg_controllable_hgrant8_out & ~n5654;
  assign n5656 = ~reg_controllable_hgrant8_out & ~n5655;
  assign n5657 = ~reg_controllable_hgrant7_out & ~n5656;
  assign n5658 = ~reg_controllable_hgrant7_out & ~n5657;
  assign n5659 = reg_controllable_hgrant9_out & ~n5658;
  assign n5660 = ~n5531 & ~n5602;
  assign n5661 = next_sys_fair<1>_out  & ~n5660;
  assign n5662 = ~n5507 & ~n5608;
  assign n5663 = ~next_sys_fair<1>_out  & ~n5662;
  assign n5664 = ~n5661 & ~n5663;
  assign n5665 = reg_controllable_hmaster3_out & ~n5664;
  assign n5666 = ~n5595 & ~n5612;
  assign n5667 = reg_controllable_hmaster2_out & ~n5666;
  assign n5668 = ~reg_controllable_hmaster2_out & ~n5660;
  assign n5669 = ~n5667 & ~n5668;
  assign n5670 = reg_controllable_hmaster1_out & ~n5669;
  assign n5671 = ~reg_controllable_hmaster1_out & ~n5660;
  assign n5672 = ~n5670 & ~n5671;
  assign n5673 = next_sys_fair<1>_out  & ~n5672;
  assign n5674 = ~n5570 & ~n5636;
  assign n5675 = reg_controllable_hmaster2_out & ~n5674;
  assign n5676 = ~reg_controllable_hmaster2_out & ~n5662;
  assign n5677 = ~n5675 & ~n5676;
  assign n5678 = reg_controllable_hmaster1_out & ~n5677;
  assign n5679 = ~reg_controllable_hmaster1_out & ~n5662;
  assign n5680 = ~n5678 & ~n5679;
  assign n5681 = ~next_sys_fair<1>_out  & ~n5680;
  assign n5682 = ~n5673 & ~n5681;
  assign n5683 = reg_controllable_hmaster0_out & ~n5682;
  assign n5684 = ~reg_controllable_hmaster0_out & ~n5664;
  assign n5685 = ~n5683 & ~n5684;
  assign n5686 = ~reg_controllable_hmaster3_out & ~n5685;
  assign n5687 = ~n5665 & ~n5686;
  assign n5688 = ~reg_controllable_hgrant6_out & ~n5687;
  assign n5689 = ~reg_controllable_hgrant6_out & ~n5688;
  assign n5690 = ~reg_controllable_hgrant8_out & ~n5689;
  assign n5691 = ~reg_controllable_hgrant8_out & ~n5690;
  assign n5692 = reg_controllable_hgrant7_out & ~n5691;
  assign n5693 = next_sys_fair<0>_out  & ~n5504;
  assign n5694 = ~next_sys_fair<0>_out  & ~n5483;
  assign n5695 = ~n5693 & ~n5694;
  assign n5696 = next_sys_fair<3>_out  & ~n5695;
  assign n5697 = ~n5531 & ~n5696;
  assign n5698 = next_sys_fair<1>_out  & ~n5697;
  assign n5699 = ~n5646 & ~n5698;
  assign n5700 = reg_controllable_hmaster0_out & ~n5699;
  assign n5701 = reg_controllable_hmaster1_out & ~n5697;
  assign n5702 = reg_controllable_hmaster2_out & ~n5697;
  assign n5703 = next_sys_fair<0>_out  & ~n5567;
  assign n5704 = ~next_sys_fair<0>_out  & ~n5550;
  assign n5705 = ~n5703 & ~n5704;
  assign n5706 = next_sys_fair<3>_out  & ~n5705;
  assign n5707 = ~n5595 & ~n5706;
  assign n5708 = ~reg_controllable_hmaster2_out & ~n5707;
  assign n5709 = ~n5702 & ~n5708;
  assign n5710 = ~reg_controllable_hmaster1_out & ~n5709;
  assign n5711 = ~n5701 & ~n5710;
  assign n5712 = next_sys_fair<1>_out  & ~n5711;
  assign n5713 = ~n5642 & ~n5712;
  assign n5714 = ~reg_controllable_hmaster0_out & ~n5713;
  assign n5715 = ~n5700 & ~n5714;
  assign n5716 = reg_controllable_hmaster3_out & ~n5715;
  assign n5717 = ~reg_controllable_hmaster3_out & ~n5699;
  assign n5718 = ~n5716 & ~n5717;
  assign n5719 = ~reg_controllable_hgrant6_out & ~n5718;
  assign n5720 = ~reg_controllable_hgrant6_out & ~n5719;
  assign n5721 = reg_controllable_hgrant8_out & ~n5720;
  assign n5722 = ~n5608 & ~n5696;
  assign n5723 = ~next_sys_fair<1>_out  & ~n5722;
  assign n5724 = ~n5661 & ~n5723;
  assign n5725 = reg_controllable_hmaster3_out & ~n5724;
  assign n5726 = reg_controllable_hmaster0_out & ~n5724;
  assign n5727 = ~n5636 & ~n5706;
  assign n5728 = reg_controllable_hmaster2_out & ~n5727;
  assign n5729 = ~reg_controllable_hmaster2_out & ~n5722;
  assign n5730 = ~n5728 & ~n5729;
  assign n5731 = reg_controllable_hmaster1_out & ~n5730;
  assign n5732 = ~reg_controllable_hmaster1_out & ~n5722;
  assign n5733 = ~n5731 & ~n5732;
  assign n5734 = ~next_sys_fair<1>_out  & ~n5733;
  assign n5735 = ~n5673 & ~n5734;
  assign n5736 = ~reg_controllable_hmaster0_out & ~n5735;
  assign n5737 = ~n5726 & ~n5736;
  assign n5738 = ~reg_controllable_hmaster3_out & ~n5737;
  assign n5739 = ~n5725 & ~n5738;
  assign n5740 = reg_controllable_hgrant6_out & ~n5739;
  assign n5741 = reg_controllable_hgrant5_out & ~n5502;
  assign n5742 = reg_controllable_hgrant4_out & ~n5500;
  assign n5743 = reg_controllable_hgrant3_out & ~n5496;
  assign n5744 = reg_controllable_hgrant1_out & ~n5494;
  assign n5745 = reg_controllable_hgrant2_out & ~n5492;
  assign n5746 = reg_controllable_hmastlock_out & ~n1253;
  assign n5747 = reg_controllable_locked_out & ~n5746;
  assign n5748 = reg_controllable_hmastlock_out & ~n5488;
  assign n5749 = ~n1254 & ~n5748;
  assign n5750 = ~reg_controllable_locked_out & ~n5749;
  assign n5751 = ~n5747 & ~n5750;
  assign n5752 = ~reg_controllable_hgrant2_out & ~n5751;
  assign n5753 = ~n5745 & ~n5752;
  assign n5754 = ~reg_controllable_hgrant1_out & ~n5753;
  assign n5755 = ~n5744 & ~n5754;
  assign n5756 = ~reg_controllable_hgrant3_out & ~n5755;
  assign n5757 = ~n5743 & ~n5756;
  assign n5758 = ~next_sys_fair<2>_out  & ~n5757;
  assign n5759 = ~next_sys_fair<2>_out  & ~n5758;
  assign n5760 = ~reg_controllable_hgrant4_out & ~n5759;
  assign n5761 = ~n5742 & ~n5760;
  assign n5762 = ~reg_controllable_hgrant5_out & ~n5761;
  assign n5763 = ~n5741 & ~n5762;
  assign n5764 = next_sys_fair<3>_out  & ~n5763;
  assign n5765 = next_sys_fair<2>_out  & ~n5477;
  assign n5766 = ~n5499 & ~n5765;
  assign n5767 = ~reg_controllable_hgrant4_out & ~n5766;
  assign n5768 = ~reg_controllable_hgrant4_out & ~n5767;
  assign n5769 = reg_controllable_hgrant5_out & ~n5768;
  assign n5770 = reg_controllable_hgrant4_out & ~n5498;
  assign n5771 = next_sys_fair<2>_out  & ~n5757;
  assign n5772 = reg_controllable_hgrant1_out & ~n5473;
  assign n5773 = ~n5754 & ~n5772;
  assign n5774 = ~reg_controllable_hgrant3_out & ~n5773;
  assign n5775 = ~n5743 & ~n5774;
  assign n5776 = ~next_sys_fair<2>_out  & ~n5775;
  assign n5777 = ~n5771 & ~n5776;
  assign n5778 = ~reg_controllable_hgrant4_out & ~n5777;
  assign n5779 = ~n5770 & ~n5778;
  assign n5780 = ~reg_controllable_hgrant5_out & ~n5779;
  assign n5781 = ~n5769 & ~n5780;
  assign n5782 = next_sys_fair<0>_out  & ~n5781;
  assign n5783 = reg_controllable_hgrant5_out & ~n5526;
  assign n5784 = ~n5523 & ~n5765;
  assign n5785 = reg_controllable_hgrant4_out & ~n5784;
  assign n5786 = reg_controllable_hgrant3_out & ~n5520;
  assign n5787 = reg_controllable_hgrant1_out & ~n5518;
  assign n5788 = reg_controllable_hgrant2_out & ~n5516;
  assign n5789 = reg_controllable_hmastlock_out & ~n1226;
  assign n5790 = reg_controllable_locked_out & ~n5789;
  assign n5791 = next_env_fair_out & ~n176;
  assign n5792 = ~next_env_fair_out & ~n119;
  assign n5793 = ~n5791 & ~n5792;
  assign n5794 = ~reg_stateG2_out & ~n5793;
  assign n5795 = ~reg_stateG2_out & ~n5794;
  assign n5796 = reg_stateA1_out & ~n5795;
  assign n5797 = ~n3663 & ~n5796;
  assign n5798 = reg_controllable_hmastlock_out & ~n5797;
  assign n5799 = ~n1229 & ~n5798;
  assign n5800 = ~reg_controllable_locked_out & ~n5799;
  assign n5801 = ~n5790 & ~n5800;
  assign n5802 = ~reg_controllable_hgrant2_out & ~n5801;
  assign n5803 = ~n5788 & ~n5802;
  assign n5804 = ~reg_controllable_hgrant1_out & ~n5803;
  assign n5805 = ~n5787 & ~n5804;
  assign n5806 = ~reg_controllable_hgrant3_out & ~n5805;
  assign n5807 = ~n5786 & ~n5806;
  assign n5808 = ~next_sys_fair<2>_out  & ~n5807;
  assign n5809 = ~n5771 & ~n5808;
  assign n5810 = ~reg_controllable_hgrant4_out & ~n5809;
  assign n5811 = ~n5785 & ~n5810;
  assign n5812 = ~reg_controllable_hgrant5_out & ~n5811;
  assign n5813 = ~n5783 & ~n5812;
  assign n5814 = ~next_sys_fair<0>_out  & ~n5813;
  assign n5815 = ~n5782 & ~n5814;
  assign n5816 = ~next_sys_fair<3>_out  & ~n5815;
  assign n5817 = ~n5764 & ~n5816;
  assign n5818 = reg_controllable_hmaster1_out & ~n5817;
  assign n5819 = reg_controllable_hmaster2_out & ~n5817;
  assign n5820 = ~reg_controllable_locked_out & ~n5488;
  assign n5821 = ~reg_controllable_locked_out & ~n5820;
  assign n5822 = ~reg_controllable_hgrant2_out & ~n5821;
  assign n5823 = ~n5745 & ~n5822;
  assign n5824 = ~reg_controllable_hgrant1_out & ~n5823;
  assign n5825 = ~n5744 & ~n5824;
  assign n5826 = ~reg_controllable_hgrant3_out & ~n5825;
  assign n5827 = ~n5743 & ~n5826;
  assign n5828 = ~next_sys_fair<2>_out  & ~n5827;
  assign n5829 = ~next_sys_fair<2>_out  & ~n5828;
  assign n5830 = ~reg_controllable_hgrant4_out & ~n5829;
  assign n5831 = ~n5742 & ~n5830;
  assign n5832 = ~reg_controllable_hgrant5_out & ~n5831;
  assign n5833 = ~n5741 & ~n5832;
  assign n5834 = next_sys_fair<3>_out  & ~n5833;
  assign n5835 = next_sys_fair<2>_out  & ~n5827;
  assign n5836 = ~n5772 & ~n5824;
  assign n5837 = ~reg_controllable_hgrant3_out & ~n5836;
  assign n5838 = ~n5743 & ~n5837;
  assign n5839 = ~next_sys_fair<2>_out  & ~n5838;
  assign n5840 = ~n5835 & ~n5839;
  assign n5841 = ~reg_controllable_hgrant4_out & ~n5840;
  assign n5842 = ~n5770 & ~n5841;
  assign n5843 = ~reg_controllable_hgrant5_out & ~n5842;
  assign n5844 = ~n5769 & ~n5843;
  assign n5845 = next_sys_fair<0>_out  & ~n5844;
  assign n5846 = ~reg_controllable_locked_out & ~n5797;
  assign n5847 = ~reg_controllable_locked_out & ~n5846;
  assign n5848 = ~reg_controllable_hgrant2_out & ~n5847;
  assign n5849 = ~n5788 & ~n5848;
  assign n5850 = ~reg_controllable_hgrant1_out & ~n5849;
  assign n5851 = ~n5787 & ~n5850;
  assign n5852 = ~reg_controllable_hgrant3_out & ~n5851;
  assign n5853 = ~n5786 & ~n5852;
  assign n5854 = ~next_sys_fair<2>_out  & ~n5853;
  assign n5855 = ~n5835 & ~n5854;
  assign n5856 = ~reg_controllable_hgrant4_out & ~n5855;
  assign n5857 = ~n5785 & ~n5856;
  assign n5858 = ~reg_controllable_hgrant5_out & ~n5857;
  assign n5859 = ~n5783 & ~n5858;
  assign n5860 = ~next_sys_fair<0>_out  & ~n5859;
  assign n5861 = ~n5845 & ~n5860;
  assign n5862 = ~next_sys_fair<3>_out  & ~n5861;
  assign n5863 = ~n5834 & ~n5862;
  assign n5864 = ~reg_controllable_hmaster2_out & ~n5863;
  assign n5865 = ~n5819 & ~n5864;
  assign n5866 = ~reg_controllable_hmaster1_out & ~n5865;
  assign n5867 = ~n5818 & ~n5866;
  assign n5868 = next_sys_fair<1>_out  & ~n5867;
  assign n5869 = reg_controllable_hgrant5_out & ~n5605;
  assign n5870 = reg_controllable_hgrant4_out & ~n5603;
  assign n5871 = reg_controllable_hgrant3_out & ~n5475;
  assign n5872 = ~n5756 & ~n5871;
  assign n5873 = next_sys_fair<2>_out  & ~n5872;
  assign n5874 = reg_controllable_hgrant2_out & ~n5471;
  assign n5875 = reg_controllable_hmastlock_out & ~n1365;
  assign n5876 = reg_controllable_locked_out & ~n5875;
  assign n5877 = ~n222 & ~n1368;
  assign n5878 = ~reg_controllable_locked_out & ~n5877;
  assign n5879 = ~n5876 & ~n5878;
  assign n5880 = ~reg_controllable_hgrant2_out & ~n5879;
  assign n5881 = ~n5874 & ~n5880;
  assign n5882 = ~reg_controllable_hgrant1_out & ~n5881;
  assign n5883 = ~n5772 & ~n5882;
  assign n5884 = ~reg_controllable_hgrant3_out & ~n5883;
  assign n5885 = ~n5871 & ~n5884;
  assign n5886 = ~next_sys_fair<2>_out  & ~n5885;
  assign n5887 = ~n5873 & ~n5886;
  assign n5888 = ~reg_controllable_hgrant4_out & ~n5887;
  assign n5889 = ~n5870 & ~n5888;
  assign n5890 = ~reg_controllable_hgrant5_out & ~n5889;
  assign n5891 = ~n5869 & ~n5890;
  assign n5892 = next_sys_fair<0>_out  & ~n5891;
  assign n5893 = ~n5752 & ~n5874;
  assign n5894 = ~reg_controllable_hgrant1_out & ~n5893;
  assign n5895 = ~n5744 & ~n5894;
  assign n5896 = ~reg_controllable_hgrant3_out & ~n5895;
  assign n5897 = ~n5743 & ~n5896;
  assign n5898 = next_sys_fair<2>_out  & ~n5897;
  assign n5899 = reg_controllable_hmastlock_out & ~n1392;
  assign n5900 = reg_controllable_locked_out & ~n5899;
  assign n5901 = ~n222 & ~n1393;
  assign n5902 = ~reg_controllable_locked_out & ~n5901;
  assign n5903 = ~n5900 & ~n5902;
  assign n5904 = ~reg_controllable_hgrant2_out & ~n5903;
  assign n5905 = ~n5874 & ~n5904;
  assign n5906 = ~reg_controllable_hgrant1_out & ~n5905;
  assign n5907 = ~n5772 & ~n5906;
  assign n5908 = ~reg_controllable_hgrant3_out & ~n5907;
  assign n5909 = ~n5871 & ~n5908;
  assign n5910 = ~next_sys_fair<2>_out  & ~n5909;
  assign n5911 = ~n5898 & ~n5910;
  assign n5912 = ~reg_controllable_hgrant4_out & ~n5911;
  assign n5913 = ~n5870 & ~n5912;
  assign n5914 = ~reg_controllable_hgrant5_out & ~n5913;
  assign n5915 = ~n5869 & ~n5914;
  assign n5916 = ~next_sys_fair<0>_out  & ~n5915;
  assign n5917 = ~n5892 & ~n5916;
  assign n5918 = ~next_sys_fair<3>_out  & ~n5917;
  assign n5919 = ~n5764 & ~n5918;
  assign n5920 = reg_controllable_hmaster1_out & ~n5919;
  assign n5921 = reg_controllable_hmaster2_out & ~n5919;
  assign n5922 = ~n5826 & ~n5871;
  assign n5923 = next_sys_fair<2>_out  & ~n5922;
  assign n5924 = ~n2869 & ~n5874;
  assign n5925 = ~reg_controllable_hgrant1_out & ~n5924;
  assign n5926 = ~n5772 & ~n5925;
  assign n5927 = ~reg_controllable_hgrant3_out & ~n5926;
  assign n5928 = ~n5871 & ~n5927;
  assign n5929 = ~next_sys_fair<2>_out  & ~n5928;
  assign n5930 = ~n5923 & ~n5929;
  assign n5931 = ~reg_controllable_hgrant4_out & ~n5930;
  assign n5932 = ~n5870 & ~n5931;
  assign n5933 = ~reg_controllable_hgrant5_out & ~n5932;
  assign n5934 = ~n5869 & ~n5933;
  assign n5935 = next_sys_fair<0>_out  & ~n5934;
  assign n5936 = ~n5822 & ~n5874;
  assign n5937 = ~reg_controllable_hgrant1_out & ~n5936;
  assign n5938 = ~n5744 & ~n5937;
  assign n5939 = ~reg_controllable_hgrant3_out & ~n5938;
  assign n5940 = ~n5743 & ~n5939;
  assign n5941 = next_sys_fair<2>_out  & ~n5940;
  assign n5942 = ~n5929 & ~n5941;
  assign n5943 = ~reg_controllable_hgrant4_out & ~n5942;
  assign n5944 = ~n5870 & ~n5943;
  assign n5945 = ~reg_controllable_hgrant5_out & ~n5944;
  assign n5946 = ~n5869 & ~n5945;
  assign n5947 = ~next_sys_fair<0>_out  & ~n5946;
  assign n5948 = ~n5935 & ~n5947;
  assign n5949 = ~next_sys_fair<3>_out  & ~n5948;
  assign n5950 = ~n5834 & ~n5949;
  assign n5951 = ~reg_controllable_hmaster2_out & ~n5950;
  assign n5952 = ~n5921 & ~n5951;
  assign n5953 = ~reg_controllable_hmaster1_out & ~n5952;
  assign n5954 = ~n5920 & ~n5953;
  assign n5955 = ~next_sys_fair<1>_out  & ~n5954;
  assign n5956 = ~n5868 & ~n5955;
  assign n5957 = reg_controllable_hmaster3_out & ~n5956;
  assign n5958 = reg_controllable_hmaster2_out & ~n5863;
  assign n5959 = reg_controllable_hgrant3_out & ~n5559;
  assign n5960 = ~n5826 & ~n5959;
  assign n5961 = ~next_sys_fair<2>_out  & ~n5960;
  assign n5962 = ~next_sys_fair<2>_out  & ~n5961;
  assign n5963 = ~reg_controllable_hgrant4_out & ~n5962;
  assign n5964 = ~n5742 & ~n5963;
  assign n5965 = ~reg_controllable_hgrant5_out & ~n5964;
  assign n5966 = ~n5741 & ~n5965;
  assign n5967 = next_sys_fair<3>_out  & ~n5966;
  assign n5968 = next_sys_fair<2>_out  & ~n5960;
  assign n5969 = ~n5837 & ~n5959;
  assign n5970 = ~next_sys_fair<2>_out  & ~n5969;
  assign n5971 = ~n5968 & ~n5970;
  assign n5972 = ~reg_controllable_hgrant4_out & ~n5971;
  assign n5973 = ~n5770 & ~n5972;
  assign n5974 = ~reg_controllable_hgrant5_out & ~n5973;
  assign n5975 = ~n5769 & ~n5974;
  assign n5976 = next_sys_fair<0>_out  & ~n5975;
  assign n5977 = reg_controllable_hgrant3_out & ~n5584;
  assign n5978 = ~n5852 & ~n5977;
  assign n5979 = ~next_sys_fair<2>_out  & ~n5978;
  assign n5980 = ~n5968 & ~n5979;
  assign n5981 = ~reg_controllable_hgrant4_out & ~n5980;
  assign n5982 = ~n5785 & ~n5981;
  assign n5983 = ~reg_controllable_hgrant5_out & ~n5982;
  assign n5984 = ~n5783 & ~n5983;
  assign n5985 = ~next_sys_fair<0>_out  & ~n5984;
  assign n5986 = ~n5976 & ~n5985;
  assign n5987 = ~next_sys_fair<3>_out  & ~n5986;
  assign n5988 = ~n5967 & ~n5987;
  assign n5989 = ~reg_controllable_hmaster2_out & ~n5988;
  assign n5990 = ~n5958 & ~n5989;
  assign n5991 = reg_controllable_hmaster1_out & ~n5990;
  assign n5992 = reg_controllable_hgrant5_out & ~n5565;
  assign n5993 = ~n5832 & ~n5992;
  assign n5994 = next_sys_fair<3>_out  & ~n5993;
  assign n5995 = next_sys_fair<2>_out  & ~n5544;
  assign n5996 = ~n5562 & ~n5995;
  assign n5997 = ~reg_controllable_hgrant4_out & ~n5996;
  assign n5998 = ~reg_controllable_hgrant4_out & ~n5997;
  assign n5999 = reg_controllable_hgrant5_out & ~n5998;
  assign n6000 = ~n5843 & ~n5999;
  assign n6001 = next_sys_fair<0>_out  & ~n6000;
  assign n6002 = reg_controllable_hgrant5_out & ~n5590;
  assign n6003 = ~n5858 & ~n6002;
  assign n6004 = ~next_sys_fair<0>_out  & ~n6003;
  assign n6005 = ~n6001 & ~n6004;
  assign n6006 = ~next_sys_fair<3>_out  & ~n6005;
  assign n6007 = ~n5994 & ~n6006;
  assign n6008 = reg_controllable_hmaster2_out & ~n6007;
  assign n6009 = reg_controllable_hgrant1_out & ~n5557;
  assign n6010 = ~n5824 & ~n6009;
  assign n6011 = ~reg_controllable_hgrant3_out & ~n6010;
  assign n6012 = ~n5743 & ~n6011;
  assign n6013 = ~next_sys_fair<2>_out  & ~n6012;
  assign n6014 = ~next_sys_fair<2>_out  & ~n6013;
  assign n6015 = ~reg_controllable_hgrant4_out & ~n6014;
  assign n6016 = ~n5742 & ~n6015;
  assign n6017 = ~reg_controllable_hgrant5_out & ~n6016;
  assign n6018 = ~n5741 & ~n6017;
  assign n6019 = next_sys_fair<3>_out  & ~n6018;
  assign n6020 = next_sys_fair<2>_out  & ~n6012;
  assign n6021 = reg_controllable_hgrant1_out & ~n5540;
  assign n6022 = ~n5824 & ~n6021;
  assign n6023 = ~reg_controllable_hgrant3_out & ~n6022;
  assign n6024 = ~n5743 & ~n6023;
  assign n6025 = ~next_sys_fair<2>_out  & ~n6024;
  assign n6026 = ~n6020 & ~n6025;
  assign n6027 = ~reg_controllable_hgrant4_out & ~n6026;
  assign n6028 = ~n5770 & ~n6027;
  assign n6029 = ~reg_controllable_hgrant5_out & ~n6028;
  assign n6030 = ~n5769 & ~n6029;
  assign n6031 = next_sys_fair<0>_out  & ~n6030;
  assign n6032 = reg_controllable_hgrant1_out & ~n5582;
  assign n6033 = ~n5850 & ~n6032;
  assign n6034 = ~reg_controllable_hgrant3_out & ~n6033;
  assign n6035 = ~n5786 & ~n6034;
  assign n6036 = ~next_sys_fair<2>_out  & ~n6035;
  assign n6037 = ~n6020 & ~n6036;
  assign n6038 = ~reg_controllable_hgrant4_out & ~n6037;
  assign n6039 = ~n5785 & ~n6038;
  assign n6040 = ~reg_controllable_hgrant5_out & ~n6039;
  assign n6041 = ~n5783 & ~n6040;
  assign n6042 = ~next_sys_fair<0>_out  & ~n6041;
  assign n6043 = ~n6031 & ~n6042;
  assign n6044 = ~next_sys_fair<3>_out  & ~n6043;
  assign n6045 = ~n6019 & ~n6044;
  assign n6046 = ~reg_controllable_hmaster2_out & ~n6045;
  assign n6047 = ~n6008 & ~n6046;
  assign n6048 = ~reg_controllable_hmaster1_out & ~n6047;
  assign n6049 = ~n5991 & ~n6048;
  assign n6050 = next_sys_fair<1>_out  & ~n6049;
  assign n6051 = reg_controllable_hmaster2_out & ~n5950;
  assign n6052 = reg_controllable_hgrant3_out & ~n5542;
  assign n6053 = ~n5826 & ~n6052;
  assign n6054 = next_sys_fair<2>_out  & ~n6053;
  assign n6055 = reg_controllable_hgrant3_out & ~n5619;
  assign n6056 = ~n5927 & ~n6055;
  assign n6057 = ~next_sys_fair<2>_out  & ~n6056;
  assign n6058 = ~n6054 & ~n6057;
  assign n6059 = ~reg_controllable_hgrant4_out & ~n6058;
  assign n6060 = ~n5870 & ~n6059;
  assign n6061 = ~reg_controllable_hgrant5_out & ~n6060;
  assign n6062 = ~n5869 & ~n6061;
  assign n6063 = next_sys_fair<0>_out  & ~n6062;
  assign n6064 = ~n5939 & ~n5959;
  assign n6065 = next_sys_fair<2>_out  & ~n6064;
  assign n6066 = ~n5927 & ~n6052;
  assign n6067 = ~next_sys_fair<2>_out  & ~n6066;
  assign n6068 = ~n6065 & ~n6067;
  assign n6069 = ~reg_controllable_hgrant4_out & ~n6068;
  assign n6070 = ~n5870 & ~n6069;
  assign n6071 = ~reg_controllable_hgrant5_out & ~n6070;
  assign n6072 = ~n5869 & ~n6071;
  assign n6073 = ~next_sys_fair<0>_out  & ~n6072;
  assign n6074 = ~n6063 & ~n6073;
  assign n6075 = ~next_sys_fair<3>_out  & ~n6074;
  assign n6076 = ~n5967 & ~n6075;
  assign n6077 = ~reg_controllable_hmaster2_out & ~n6076;
  assign n6078 = ~n6051 & ~n6077;
  assign n6079 = reg_controllable_hmaster1_out & ~n6078;
  assign n6080 = reg_controllable_hgrant5_out & ~n5625;
  assign n6081 = ~n5933 & ~n6080;
  assign n6082 = next_sys_fair<0>_out  & ~n6081;
  assign n6083 = reg_controllable_hgrant5_out & ~n5631;
  assign n6084 = ~n5945 & ~n6083;
  assign n6085 = ~next_sys_fair<0>_out  & ~n6084;
  assign n6086 = ~n6082 & ~n6085;
  assign n6087 = ~next_sys_fair<3>_out  & ~n6086;
  assign n6088 = ~n5994 & ~n6087;
  assign n6089 = reg_controllable_hmaster2_out & ~n6088;
  assign n6090 = ~n5871 & ~n6011;
  assign n6091 = next_sys_fair<2>_out  & ~n6090;
  assign n6092 = reg_controllable_hgrant1_out & ~n5617;
  assign n6093 = ~n5925 & ~n6092;
  assign n6094 = ~reg_controllable_hgrant3_out & ~n6093;
  assign n6095 = ~n5871 & ~n6094;
  assign n6096 = ~next_sys_fair<2>_out  & ~n6095;
  assign n6097 = ~n6091 & ~n6096;
  assign n6098 = ~reg_controllable_hgrant4_out & ~n6097;
  assign n6099 = ~n5870 & ~n6098;
  assign n6100 = ~reg_controllable_hgrant5_out & ~n6099;
  assign n6101 = ~n5869 & ~n6100;
  assign n6102 = next_sys_fair<0>_out  & ~n6101;
  assign n6103 = ~n5937 & ~n6009;
  assign n6104 = ~reg_controllable_hgrant3_out & ~n6103;
  assign n6105 = ~n5743 & ~n6104;
  assign n6106 = next_sys_fair<2>_out  & ~n6105;
  assign n6107 = ~n5925 & ~n6021;
  assign n6108 = ~reg_controllable_hgrant3_out & ~n6107;
  assign n6109 = ~n5871 & ~n6108;
  assign n6110 = ~next_sys_fair<2>_out  & ~n6109;
  assign n6111 = ~n6106 & ~n6110;
  assign n6112 = ~reg_controllable_hgrant4_out & ~n6111;
  assign n6113 = ~n5870 & ~n6112;
  assign n6114 = ~reg_controllable_hgrant5_out & ~n6113;
  assign n6115 = ~n5869 & ~n6114;
  assign n6116 = ~next_sys_fair<0>_out  & ~n6115;
  assign n6117 = ~n6102 & ~n6116;
  assign n6118 = ~next_sys_fair<3>_out  & ~n6117;
  assign n6119 = ~n6019 & ~n6118;
  assign n6120 = ~reg_controllable_hmaster2_out & ~n6119;
  assign n6121 = ~n6089 & ~n6120;
  assign n6122 = ~reg_controllable_hmaster1_out & ~n6121;
  assign n6123 = ~n6079 & ~n6122;
  assign n6124 = ~next_sys_fair<1>_out  & ~n6123;
  assign n6125 = ~n6050 & ~n6124;
  assign n6126 = reg_controllable_hmaster0_out & ~n6125;
  assign n6127 = reg_controllable_hgrant2_out & ~n5555;
  assign n6128 = ~n5822 & ~n6127;
  assign n6129 = ~reg_controllable_hgrant1_out & ~n6128;
  assign n6130 = ~n5744 & ~n6129;
  assign n6131 = ~reg_controllable_hgrant3_out & ~n6130;
  assign n6132 = ~n5743 & ~n6131;
  assign n6133 = ~next_sys_fair<2>_out  & ~n6132;
  assign n6134 = ~next_sys_fair<2>_out  & ~n6133;
  assign n6135 = ~reg_controllable_hgrant4_out & ~n6134;
  assign n6136 = ~n5742 & ~n6135;
  assign n6137 = ~reg_controllable_hgrant5_out & ~n6136;
  assign n6138 = ~n5741 & ~n6137;
  assign n6139 = next_sys_fair<3>_out  & ~n6138;
  assign n6140 = next_sys_fair<2>_out  & ~n6132;
  assign n6141 = ~n5772 & ~n6129;
  assign n6142 = ~reg_controllable_hgrant3_out & ~n6141;
  assign n6143 = ~n5743 & ~n6142;
  assign n6144 = ~next_sys_fair<2>_out  & ~n6143;
  assign n6145 = ~n6140 & ~n6144;
  assign n6146 = ~reg_controllable_hgrant4_out & ~n6145;
  assign n6147 = ~n5770 & ~n6146;
  assign n6148 = ~reg_controllable_hgrant5_out & ~n6147;
  assign n6149 = ~n5769 & ~n6148;
  assign n6150 = next_sys_fair<0>_out  & ~n6149;
  assign n6151 = reg_controllable_hgrant2_out & ~n5580;
  assign n6152 = ~n5848 & ~n6151;
  assign n6153 = ~reg_controllable_hgrant1_out & ~n6152;
  assign n6154 = ~n5787 & ~n6153;
  assign n6155 = ~reg_controllable_hgrant3_out & ~n6154;
  assign n6156 = ~n5786 & ~n6155;
  assign n6157 = ~next_sys_fair<2>_out  & ~n6156;
  assign n6158 = ~n6140 & ~n6157;
  assign n6159 = ~reg_controllable_hgrant4_out & ~n6158;
  assign n6160 = ~n5785 & ~n6159;
  assign n6161 = ~reg_controllable_hgrant5_out & ~n6160;
  assign n6162 = ~n5783 & ~n6161;
  assign n6163 = ~next_sys_fair<0>_out  & ~n6162;
  assign n6164 = ~n6150 & ~n6163;
  assign n6165 = ~next_sys_fair<3>_out  & ~n6164;
  assign n6166 = ~n6139 & ~n6165;
  assign n6167 = ~reg_controllable_hmaster2_out & ~n6166;
  assign n6168 = ~n5958 & ~n6167;
  assign n6169 = reg_controllable_hmaster1_out & ~n6168;
  assign n6170 = reg_controllable_hgrant4_out & ~n5563;
  assign n6171 = ~n5830 & ~n6170;
  assign n6172 = ~reg_controllable_hgrant5_out & ~n6171;
  assign n6173 = ~n5741 & ~n6172;
  assign n6174 = next_sys_fair<3>_out  & ~n6173;
  assign n6175 = reg_controllable_hgrant4_out & ~n5561;
  assign n6176 = ~n5841 & ~n6175;
  assign n6177 = ~reg_controllable_hgrant5_out & ~n6176;
  assign n6178 = ~n5769 & ~n6177;
  assign n6179 = next_sys_fair<0>_out  & ~n6178;
  assign n6180 = ~n5587 & ~n5995;
  assign n6181 = reg_controllable_hgrant4_out & ~n6180;
  assign n6182 = ~n5856 & ~n6181;
  assign n6183 = ~reg_controllable_hgrant5_out & ~n6182;
  assign n6184 = ~n5783 & ~n6183;
  assign n6185 = ~next_sys_fair<0>_out  & ~n6184;
  assign n6186 = ~n6179 & ~n6185;
  assign n6187 = ~next_sys_fair<3>_out  & ~n6186;
  assign n6188 = ~n6174 & ~n6187;
  assign n6189 = reg_controllable_hmaster2_out & ~n6188;
  assign n6190 = ~n5864 & ~n6189;
  assign n6191 = ~reg_controllable_hmaster1_out & ~n6190;
  assign n6192 = ~n6169 & ~n6191;
  assign n6193 = next_sys_fair<1>_out  & ~n6192;
  assign n6194 = ~n5871 & ~n6131;
  assign n6195 = next_sys_fair<2>_out  & ~n6194;
  assign n6196 = reg_controllable_hgrant2_out & ~n5615;
  assign n6197 = ~n2869 & ~n6196;
  assign n6198 = ~reg_controllable_hgrant1_out & ~n6197;
  assign n6199 = ~n5772 & ~n6198;
  assign n6200 = ~reg_controllable_hgrant3_out & ~n6199;
  assign n6201 = ~n5871 & ~n6200;
  assign n6202 = ~next_sys_fair<2>_out  & ~n6201;
  assign n6203 = ~n6195 & ~n6202;
  assign n6204 = ~reg_controllable_hgrant4_out & ~n6203;
  assign n6205 = ~n5870 & ~n6204;
  assign n6206 = ~reg_controllable_hgrant5_out & ~n6205;
  assign n6207 = ~n5869 & ~n6206;
  assign n6208 = next_sys_fair<0>_out  & ~n6207;
  assign n6209 = reg_controllable_hgrant2_out & ~n5538;
  assign n6210 = ~n5822 & ~n6209;
  assign n6211 = ~reg_controllable_hgrant1_out & ~n6210;
  assign n6212 = ~n5744 & ~n6211;
  assign n6213 = ~reg_controllable_hgrant3_out & ~n6212;
  assign n6214 = ~n5743 & ~n6213;
  assign n6215 = next_sys_fair<2>_out  & ~n6214;
  assign n6216 = ~n2869 & ~n6209;
  assign n6217 = ~reg_controllable_hgrant1_out & ~n6216;
  assign n6218 = ~n5772 & ~n6217;
  assign n6219 = ~reg_controllable_hgrant3_out & ~n6218;
  assign n6220 = ~n5871 & ~n6219;
  assign n6221 = ~next_sys_fair<2>_out  & ~n6220;
  assign n6222 = ~n6215 & ~n6221;
  assign n6223 = ~reg_controllable_hgrant4_out & ~n6222;
  assign n6224 = ~n5870 & ~n6223;
  assign n6225 = ~reg_controllable_hgrant5_out & ~n6224;
  assign n6226 = ~n5869 & ~n6225;
  assign n6227 = ~next_sys_fair<0>_out  & ~n6226;
  assign n6228 = ~n6208 & ~n6227;
  assign n6229 = ~next_sys_fair<3>_out  & ~n6228;
  assign n6230 = ~n6139 & ~n6229;
  assign n6231 = ~reg_controllable_hmaster2_out & ~n6230;
  assign n6232 = ~n6051 & ~n6231;
  assign n6233 = reg_controllable_hmaster1_out & ~n6232;
  assign n6234 = reg_controllable_hgrant4_out & ~n5623;
  assign n6235 = ~n5931 & ~n6234;
  assign n6236 = ~reg_controllable_hgrant5_out & ~n6235;
  assign n6237 = ~n5869 & ~n6236;
  assign n6238 = next_sys_fair<0>_out  & ~n6237;
  assign n6239 = reg_controllable_hgrant4_out & ~n5629;
  assign n6240 = ~n5943 & ~n6239;
  assign n6241 = ~reg_controllable_hgrant5_out & ~n6240;
  assign n6242 = ~n5869 & ~n6241;
  assign n6243 = ~next_sys_fair<0>_out  & ~n6242;
  assign n6244 = ~n6238 & ~n6243;
  assign n6245 = ~next_sys_fair<3>_out  & ~n6244;
  assign n6246 = ~n6174 & ~n6245;
  assign n6247 = reg_controllable_hmaster2_out & ~n6246;
  assign n6248 = ~n5951 & ~n6247;
  assign n6249 = ~reg_controllable_hmaster1_out & ~n6248;
  assign n6250 = ~n6233 & ~n6249;
  assign n6251 = ~next_sys_fair<1>_out  & ~n6250;
  assign n6252 = ~n6193 & ~n6251;
  assign n6253 = ~reg_controllable_hmaster0_out & ~n6252;
  assign n6254 = ~n6126 & ~n6253;
  assign n6255 = ~reg_controllable_hmaster3_out & ~n6254;
  assign n6256 = ~n5957 & ~n6255;
  assign n6257 = ~reg_controllable_hgrant6_out & ~n6256;
  assign n6258 = ~n5740 & ~n6257;
  assign n6259 = ~reg_controllable_hgrant8_out & ~n6258;
  assign n6260 = ~n5721 & ~n6259;
  assign n6261 = ~reg_controllable_hgrant7_out & ~n6260;
  assign n6262 = ~n5692 & ~n6261;
  assign n6263 = ~reg_controllable_hgrant9_out & ~n6262;
  assign n6264 = ~n5659 & ~n6263;
  assign n6265 = reg_controllable_nhgrant0_out & ~n6264;
  assign n6266 = ~n156 & ~n5491;
  assign n6267 = ~reg_controllable_hgrant2_out & ~n6266;
  assign n6268 = ~reg_controllable_hgrant2_out & ~n6267;
  assign n6269 = ~reg_controllable_hgrant1_out & ~n6268;
  assign n6270 = ~reg_controllable_hgrant1_out & ~n6269;
  assign n6271 = ~reg_controllable_hgrant3_out & ~n6270;
  assign n6272 = ~reg_controllable_hgrant3_out & ~n6271;
  assign n6273 = ~next_sys_fair<2>_out  & ~n6272;
  assign n6274 = ~next_sys_fair<2>_out  & ~n6273;
  assign n6275 = ~reg_controllable_hgrant4_out & ~n6274;
  assign n6276 = ~reg_controllable_hgrant4_out & ~n6275;
  assign n6277 = ~reg_controllable_hgrant5_out & ~n6276;
  assign n6278 = ~reg_controllable_hgrant5_out & ~n6277;
  assign n6279 = next_sys_fair<3>_out  & ~n6278;
  assign n6280 = ~reg_controllable_hgrant4_out & ~n6272;
  assign n6281 = ~reg_controllable_hgrant4_out & ~n6280;
  assign n6282 = ~reg_controllable_hgrant5_out & ~n6281;
  assign n6283 = ~reg_controllable_hgrant5_out & ~n6282;
  assign n6284 = next_sys_fair<0>_out  & ~n6283;
  assign n6285 = next_sys_fair<2>_out  & ~n6272;
  assign n6286 = ~reg_controllable_hgrant2_out & ~n123;
  assign n6287 = ~reg_controllable_hgrant2_out & ~n6286;
  assign n6288 = ~reg_controllable_hgrant1_out & ~n6287;
  assign n6289 = ~reg_controllable_hgrant1_out & ~n6288;
  assign n6290 = ~reg_controllable_hgrant3_out & ~n6289;
  assign n6291 = ~reg_controllable_hgrant3_out & ~n6290;
  assign n6292 = ~next_sys_fair<2>_out  & ~n6291;
  assign n6293 = ~n6285 & ~n6292;
  assign n6294 = ~reg_controllable_hgrant4_out & ~n6293;
  assign n6295 = ~reg_controllable_hgrant4_out & ~n6294;
  assign n6296 = ~reg_controllable_hgrant5_out & ~n6295;
  assign n6297 = ~reg_controllable_hgrant5_out & ~n6296;
  assign n6298 = ~next_sys_fair<0>_out  & ~n6297;
  assign n6299 = ~n6284 & ~n6298;
  assign n6300 = ~next_sys_fair<3>_out  & ~n6299;
  assign n6301 = ~n6279 & ~n6300;
  assign n6302 = next_sys_fair<1>_out  & ~n6301;
  assign n6303 = ~next_sys_fair<3>_out  & ~n6297;
  assign n6304 = ~n6279 & ~n6303;
  assign n6305 = ~next_sys_fair<1>_out  & ~n6304;
  assign n6306 = ~n6302 & ~n6305;
  assign n6307 = reg_controllable_hmaster3_out & ~n6306;
  assign n6308 = reg_controllable_hmaster0_out & ~n6306;
  assign n6309 = reg_controllable_hmaster1_out & ~n6301;
  assign n6310 = reg_controllable_hmaster2_out & ~n6301;
  assign n6311 = ~n274 & ~n5554;
  assign n6312 = ~reg_controllable_hgrant2_out & ~n6311;
  assign n6313 = ~reg_controllable_hgrant2_out & ~n6312;
  assign n6314 = ~reg_controllable_hgrant1_out & ~n6313;
  assign n6315 = ~reg_controllable_hgrant1_out & ~n6314;
  assign n6316 = ~reg_controllable_hgrant3_out & ~n6315;
  assign n6317 = ~reg_controllable_hgrant3_out & ~n6316;
  assign n6318 = ~next_sys_fair<2>_out  & ~n6317;
  assign n6319 = ~next_sys_fair<2>_out  & ~n6318;
  assign n6320 = ~reg_controllable_hgrant4_out & ~n6319;
  assign n6321 = ~reg_controllable_hgrant4_out & ~n6320;
  assign n6322 = ~reg_controllable_hgrant5_out & ~n6321;
  assign n6323 = ~reg_controllable_hgrant5_out & ~n6322;
  assign n6324 = next_sys_fair<3>_out  & ~n6323;
  assign n6325 = ~reg_controllable_hgrant4_out & ~n6317;
  assign n6326 = ~reg_controllable_hgrant4_out & ~n6325;
  assign n6327 = ~reg_controllable_hgrant5_out & ~n6326;
  assign n6328 = ~reg_controllable_hgrant5_out & ~n6327;
  assign n6329 = next_sys_fair<0>_out  & ~n6328;
  assign n6330 = next_sys_fair<2>_out  & ~n6317;
  assign n6331 = ~n221 & ~n5537;
  assign n6332 = ~reg_controllable_hgrant2_out & ~n6331;
  assign n6333 = ~reg_controllable_hgrant2_out & ~n6332;
  assign n6334 = ~reg_controllable_hgrant1_out & ~n6333;
  assign n6335 = ~reg_controllable_hgrant1_out & ~n6334;
  assign n6336 = ~reg_controllable_hgrant3_out & ~n6335;
  assign n6337 = ~reg_controllable_hgrant3_out & ~n6336;
  assign n6338 = ~next_sys_fair<2>_out  & ~n6337;
  assign n6339 = ~n6330 & ~n6338;
  assign n6340 = ~reg_controllable_hgrant4_out & ~n6339;
  assign n6341 = ~reg_controllable_hgrant4_out & ~n6340;
  assign n6342 = ~reg_controllable_hgrant5_out & ~n6341;
  assign n6343 = ~reg_controllable_hgrant5_out & ~n6342;
  assign n6344 = ~next_sys_fair<0>_out  & ~n6343;
  assign n6345 = ~n6329 & ~n6344;
  assign n6346 = ~next_sys_fair<3>_out  & ~n6345;
  assign n6347 = ~n6324 & ~n6346;
  assign n6348 = ~reg_controllable_hmaster2_out & ~n6347;
  assign n6349 = ~n6310 & ~n6348;
  assign n6350 = ~reg_controllable_hmaster1_out & ~n6349;
  assign n6351 = ~n6309 & ~n6350;
  assign n6352 = next_sys_fair<1>_out  & ~n6351;
  assign n6353 = reg_controllable_hmaster1_out & ~n6304;
  assign n6354 = reg_controllable_hmaster2_out & ~n6304;
  assign n6355 = ~n337 & ~n5614;
  assign n6356 = ~reg_controllable_hgrant2_out & ~n6355;
  assign n6357 = ~reg_controllable_hgrant2_out & ~n6356;
  assign n6358 = ~reg_controllable_hgrant1_out & ~n6357;
  assign n6359 = ~reg_controllable_hgrant1_out & ~n6358;
  assign n6360 = ~reg_controllable_hgrant3_out & ~n6359;
  assign n6361 = ~reg_controllable_hgrant3_out & ~n6360;
  assign n6362 = ~next_sys_fair<2>_out  & ~n6361;
  assign n6363 = ~n6330 & ~n6362;
  assign n6364 = ~reg_controllable_hgrant4_out & ~n6363;
  assign n6365 = ~reg_controllable_hgrant4_out & ~n6364;
  assign n6366 = ~reg_controllable_hgrant5_out & ~n6365;
  assign n6367 = ~reg_controllable_hgrant5_out & ~n6366;
  assign n6368 = next_sys_fair<0>_out  & ~n6367;
  assign n6369 = ~n368 & ~n5537;
  assign n6370 = ~reg_controllable_hgrant2_out & ~n6369;
  assign n6371 = ~reg_controllable_hgrant2_out & ~n6370;
  assign n6372 = ~reg_controllable_hgrant1_out & ~n6371;
  assign n6373 = ~reg_controllable_hgrant1_out & ~n6372;
  assign n6374 = ~reg_controllable_hgrant3_out & ~n6373;
  assign n6375 = ~reg_controllable_hgrant3_out & ~n6374;
  assign n6376 = ~next_sys_fair<2>_out  & ~n6375;
  assign n6377 = ~n6330 & ~n6376;
  assign n6378 = ~reg_controllable_hgrant4_out & ~n6377;
  assign n6379 = ~reg_controllable_hgrant4_out & ~n6378;
  assign n6380 = ~reg_controllable_hgrant5_out & ~n6379;
  assign n6381 = ~reg_controllable_hgrant5_out & ~n6380;
  assign n6382 = ~next_sys_fair<0>_out  & ~n6381;
  assign n6383 = ~n6368 & ~n6382;
  assign n6384 = ~next_sys_fair<3>_out  & ~n6383;
  assign n6385 = ~n6324 & ~n6384;
  assign n6386 = ~reg_controllable_hmaster2_out & ~n6385;
  assign n6387 = ~n6354 & ~n6386;
  assign n6388 = ~reg_controllable_hmaster1_out & ~n6387;
  assign n6389 = ~n6353 & ~n6388;
  assign n6390 = ~next_sys_fair<1>_out  & ~n6389;
  assign n6391 = ~n6352 & ~n6390;
  assign n6392 = ~reg_controllable_hmaster0_out & ~n6391;
  assign n6393 = ~n6308 & ~n6392;
  assign n6394 = ~reg_controllable_hmaster3_out & ~n6393;
  assign n6395 = ~n6307 & ~n6394;
  assign n6396 = ~reg_controllable_hgrant6_out & ~n6395;
  assign n6397 = ~reg_controllable_hgrant6_out & ~n6396;
  assign n6398 = ~reg_controllable_hgrant8_out & ~n6397;
  assign n6399 = ~reg_controllable_hgrant8_out & ~n6398;
  assign n6400 = ~reg_controllable_hgrant7_out & ~n6399;
  assign n6401 = ~reg_controllable_hgrant7_out & ~n6400;
  assign n6402 = ~reg_controllable_hgrant9_out & ~n6401;
  assign n6403 = ~reg_controllable_hgrant9_out & ~n6402;
  assign n6404 = ~reg_controllable_nhgrant0_out & ~n6403;
  assign n6405 = ~n6265 & ~n6404;
  assign n6406 = reg_i_hready_out & ~n6405;
  assign n6407 = ~next_sys_fair<2>_out  & ~n1255;
  assign n6408 = ~next_sys_fair<2>_out  & ~n6407;
  assign n6409 = next_sys_fair<3>_out  & ~n6408;
  assign n6410 = next_sys_fair<0>_out  & ~n1255;
  assign n6411 = next_sys_fair<2>_out  & ~n1255;
  assign n6412 = ~next_sys_fair<2>_out  & ~n1230;
  assign n6413 = ~n6411 & ~n6412;
  assign n6414 = ~next_sys_fair<0>_out  & ~n6413;
  assign n6415 = ~n6410 & ~n6414;
  assign n6416 = ~next_sys_fair<3>_out  & ~n6415;
  assign n6417 = ~n6409 & ~n6416;
  assign n6418 = reg_controllable_hmaster1_out & ~n6417;
  assign n6419 = reg_controllable_hmaster2_out & ~n6417;
  assign n6420 = ~next_sys_fair<2>_out  & ~n1500;
  assign n6421 = ~next_sys_fair<2>_out  & ~n6420;
  assign n6422 = next_sys_fair<0>_out  & ~n6421;
  assign n6423 = ~next_sys_fair<2>_out  & ~n1521;
  assign n6424 = ~next_sys_fair<2>_out  & ~n6423;
  assign n6425 = ~next_sys_fair<0>_out  & ~n6424;
  assign n6426 = ~n6422 & ~n6425;
  assign n6427 = next_sys_fair<3>_out  & ~n6426;
  assign n6428 = next_sys_fair<0>_out  & ~n1521;
  assign n6429 = next_sys_fair<2>_out  & ~n1521;
  assign n6430 = ~next_sys_fair<2>_out  & ~n1481;
  assign n6431 = ~n6429 & ~n6430;
  assign n6432 = ~next_sys_fair<0>_out  & ~n6431;
  assign n6433 = ~n6428 & ~n6432;
  assign n6434 = ~next_sys_fair<3>_out  & ~n6433;
  assign n6435 = ~n6427 & ~n6434;
  assign n6436 = ~reg_controllable_hmaster2_out & ~n6435;
  assign n6437 = ~n6419 & ~n6436;
  assign n6438 = ~reg_controllable_hmaster1_out & ~n6437;
  assign n6439 = ~n6418 & ~n6438;
  assign n6440 = next_sys_fair<1>_out  & ~n6439;
  assign n6441 = ~next_sys_fair<2>_out  & ~n1369;
  assign n6442 = ~n6411 & ~n6441;
  assign n6443 = next_sys_fair<0>_out  & ~n6442;
  assign n6444 = ~next_sys_fair<2>_out  & ~n1394;
  assign n6445 = ~n6411 & ~n6444;
  assign n6446 = ~next_sys_fair<0>_out  & ~n6445;
  assign n6447 = ~n6443 & ~n6446;
  assign n6448 = ~next_sys_fair<3>_out  & ~n6447;
  assign n6449 = ~n6409 & ~n6448;
  assign n6450 = reg_controllable_hmaster1_out & ~n6449;
  assign n6451 = reg_controllable_hmaster2_out & ~n6449;
  assign n6452 = next_sys_fair<3>_out  & ~n6424;
  assign n6453 = ~next_sys_fair<2>_out  & ~n1554;
  assign n6454 = ~n6429 & ~n6453;
  assign n6455 = next_sys_fair<0>_out  & ~n6454;
  assign n6456 = ~n6420 & ~n6429;
  assign n6457 = ~next_sys_fair<0>_out  & ~n6456;
  assign n6458 = ~n6455 & ~n6457;
  assign n6459 = ~next_sys_fair<3>_out  & ~n6458;
  assign n6460 = ~n6452 & ~n6459;
  assign n6461 = ~reg_controllable_hmaster2_out & ~n6460;
  assign n6462 = ~n6451 & ~n6461;
  assign n6463 = ~reg_controllable_hmaster1_out & ~n6462;
  assign n6464 = ~n6450 & ~n6463;
  assign n6465 = ~next_sys_fair<1>_out  & ~n6464;
  assign n6466 = ~n6440 & ~n6465;
  assign n6467 = reg_controllable_hmaster0_out & ~n6466;
  assign n6468 = next_sys_fair<0>_out  & ~n6424;
  assign n6469 = ~next_sys_fair<0>_out  & ~n6421;
  assign n6470 = ~n6468 & ~n6469;
  assign n6471 = next_sys_fair<3>_out  & ~n6470;
  assign n6472 = ~n6434 & ~n6471;
  assign n6473 = ~reg_controllable_hmaster2_out & ~n6472;
  assign n6474 = ~n6419 & ~n6473;
  assign n6475 = ~reg_controllable_hmaster1_out & ~n6474;
  assign n6476 = ~n6418 & ~n6475;
  assign n6477 = next_sys_fair<1>_out  & ~n6476;
  assign n6478 = ~n6465 & ~n6477;
  assign n6479 = ~reg_controllable_hmaster0_out & ~n6478;
  assign n6480 = ~n6467 & ~n6479;
  assign n6481 = reg_controllable_hmaster3_out & ~n6480;
  assign n6482 = ~n6434 & ~n6452;
  assign n6483 = reg_controllable_hmaster1_out & ~n6482;
  assign n6484 = next_sys_fair<2>_out  & ~n1500;
  assign n6485 = ~n6423 & ~n6484;
  assign n6486 = next_sys_fair<0>_out  & ~n6485;
  assign n6487 = ~n6432 & ~n6486;
  assign n6488 = ~next_sys_fair<3>_out  & ~n6487;
  assign n6489 = ~n6452 & ~n6488;
  assign n6490 = reg_controllable_hmaster2_out & ~n6489;
  assign n6491 = next_sys_fair<0>_out  & ~n6456;
  assign n6492 = ~n6432 & ~n6491;
  assign n6493 = ~next_sys_fair<3>_out  & ~n6492;
  assign n6494 = ~n6452 & ~n6493;
  assign n6495 = ~reg_controllable_hmaster2_out & ~n6494;
  assign n6496 = ~n6490 & ~n6495;
  assign n6497 = ~reg_controllable_hmaster1_out & ~n6496;
  assign n6498 = ~n6483 & ~n6497;
  assign n6499 = next_sys_fair<1>_out  & ~n6498;
  assign n6500 = ~n6427 & ~n6459;
  assign n6501 = reg_controllable_hmaster2_out & ~n6500;
  assign n6502 = ~n6453 & ~n6484;
  assign n6503 = next_sys_fair<0>_out  & ~n6502;
  assign n6504 = ~n6457 & ~n6503;
  assign n6505 = ~next_sys_fair<3>_out  & ~n6504;
  assign n6506 = ~n6452 & ~n6505;
  assign n6507 = ~reg_controllable_hmaster2_out & ~n6506;
  assign n6508 = ~n6501 & ~n6507;
  assign n6509 = reg_controllable_hmaster1_out & ~n6508;
  assign n6510 = ~reg_controllable_hmaster1_out & ~n6460;
  assign n6511 = ~n6509 & ~n6510;
  assign n6512 = ~next_sys_fair<1>_out  & ~n6511;
  assign n6513 = ~n6499 & ~n6512;
  assign n6514 = reg_controllable_hmaster0_out & ~n6513;
  assign n6515 = ~n6430 & ~n6484;
  assign n6516 = ~next_sys_fair<0>_out  & ~n6515;
  assign n6517 = ~n6428 & ~n6516;
  assign n6518 = ~next_sys_fair<3>_out  & ~n6517;
  assign n6519 = ~n6452 & ~n6518;
  assign n6520 = reg_controllable_hmaster2_out & ~n6519;
  assign n6521 = ~next_sys_fair<2>_out  & ~n1320;
  assign n6522 = ~next_sys_fair<2>_out  & ~n6521;
  assign n6523 = next_sys_fair<3>_out  & ~n6522;
  assign n6524 = next_sys_fair<0>_out  & ~n1320;
  assign n6525 = next_sys_fair<2>_out  & ~n1320;
  assign n6526 = ~next_sys_fair<2>_out  & ~n1294;
  assign n6527 = ~n6525 & ~n6526;
  assign n6528 = ~next_sys_fair<0>_out  & ~n6527;
  assign n6529 = ~n6524 & ~n6528;
  assign n6530 = ~next_sys_fair<3>_out  & ~n6529;
  assign n6531 = ~n6523 & ~n6530;
  assign n6532 = ~reg_controllable_hmaster2_out & ~n6531;
  assign n6533 = ~n6520 & ~n6532;
  assign n6534 = ~reg_controllable_hmaster1_out & ~n6533;
  assign n6535 = ~n6483 & ~n6534;
  assign n6536 = next_sys_fair<1>_out  & ~n6535;
  assign n6537 = ~n6459 & ~n6471;
  assign n6538 = reg_controllable_hmaster2_out & ~n6537;
  assign n6539 = ~next_sys_fair<0>_out  & ~n1500;
  assign n6540 = ~n6455 & ~n6539;
  assign n6541 = ~next_sys_fair<3>_out  & ~n6540;
  assign n6542 = ~n6452 & ~n6541;
  assign n6543 = ~reg_controllable_hmaster2_out & ~n6542;
  assign n6544 = ~n6538 & ~n6543;
  assign n6545 = reg_controllable_hmaster1_out & ~n6544;
  assign n6546 = reg_controllable_hmaster2_out & ~n6460;
  assign n6547 = ~next_sys_fair<2>_out  & ~n1425;
  assign n6548 = ~n6525 & ~n6547;
  assign n6549 = next_sys_fair<0>_out  & ~n6548;
  assign n6550 = ~next_sys_fair<2>_out  & ~n1446;
  assign n6551 = ~n6525 & ~n6550;
  assign n6552 = ~next_sys_fair<0>_out  & ~n6551;
  assign n6553 = ~n6549 & ~n6552;
  assign n6554 = ~next_sys_fair<3>_out  & ~n6553;
  assign n6555 = ~n6523 & ~n6554;
  assign n6556 = ~reg_controllable_hmaster2_out & ~n6555;
  assign n6557 = ~n6546 & ~n6556;
  assign n6558 = ~reg_controllable_hmaster1_out & ~n6557;
  assign n6559 = ~n6545 & ~n6558;
  assign n6560 = ~next_sys_fair<1>_out  & ~n6559;
  assign n6561 = ~n6536 & ~n6560;
  assign n6562 = ~reg_controllable_hmaster0_out & ~n6561;
  assign n6563 = ~n6514 & ~n6562;
  assign n6564 = ~reg_controllable_hmaster3_out & ~n6563;
  assign n6565 = ~n6481 & ~n6564;
  assign n6566 = ~reg_i_hready_out & ~n6565;
  assign n6567 = ~n6406 & ~n6566;
  assign n6568 = reg_i_hlock0_out & ~n6567;
  assign n6569 = ~reg_controllable_locked_out & ~n181;
  assign n6570 = ~reg_controllable_hgrant2_out & ~n6569;
  assign n6571 = ~reg_controllable_hgrant2_out & ~n6570;
  assign n6572 = ~reg_controllable_hgrant1_out & ~n6571;
  assign n6573 = ~reg_controllable_hgrant1_out & ~n6572;
  assign n6574 = ~reg_controllable_hgrant3_out & ~n6573;
  assign n6575 = ~reg_controllable_hgrant3_out & ~n6574;
  assign n6576 = ~next_sys_fair<2>_out  & ~n6575;
  assign n6577 = ~next_sys_fair<2>_out  & ~n6576;
  assign n6578 = ~reg_controllable_hgrant4_out & ~n6577;
  assign n6579 = ~reg_controllable_hgrant4_out & ~n6578;
  assign n6580 = ~reg_controllable_hgrant5_out & ~n6579;
  assign n6581 = ~reg_controllable_hgrant5_out & ~n6580;
  assign n6582 = ~next_sys_fair<0>_out  & ~n6581;
  assign n6583 = ~n3042 & ~n6582;
  assign n6584 = next_sys_fair<3>_out  & ~n6583;
  assign n6585 = ~reg_controllable_hgrant4_out & ~n6575;
  assign n6586 = ~reg_controllable_hgrant4_out & ~n6585;
  assign n6587 = ~reg_controllable_hgrant5_out & ~n6586;
  assign n6588 = ~reg_controllable_hgrant5_out & ~n6587;
  assign n6589 = next_sys_fair<0>_out  & ~n6588;
  assign n6590 = next_sys_fair<2>_out  & ~n6575;
  assign n6591 = ~n2894 & ~n6590;
  assign n6592 = ~reg_controllable_hgrant4_out & ~n6591;
  assign n6593 = ~reg_controllable_hgrant4_out & ~n6592;
  assign n6594 = ~reg_controllable_hgrant5_out & ~n6593;
  assign n6595 = ~reg_controllable_hgrant5_out & ~n6594;
  assign n6596 = ~next_sys_fair<0>_out  & ~n6595;
  assign n6597 = ~n6589 & ~n6596;
  assign n6598 = ~next_sys_fair<3>_out  & ~n6597;
  assign n6599 = ~n6584 & ~n6598;
  assign n6600 = reg_controllable_hmaster1_out & ~n6599;
  assign n6601 = reg_controllable_hmaster2_out & ~n6599;
  assign n6602 = ~n2941 & ~n3051;
  assign n6603 = ~reg_controllable_hgrant2_out & ~n6602;
  assign n6604 = ~reg_controllable_hgrant2_out & ~n6603;
  assign n6605 = ~reg_controllable_hgrant1_out & ~n6604;
  assign n6606 = ~reg_controllable_hgrant1_out & ~n6605;
  assign n6607 = ~reg_controllable_hgrant3_out & ~n6606;
  assign n6608 = ~reg_controllable_hgrant3_out & ~n6607;
  assign n6609 = ~next_sys_fair<2>_out  & ~n6608;
  assign n6610 = ~next_sys_fair<2>_out  & ~n6609;
  assign n6611 = ~reg_controllable_hgrant4_out & ~n6610;
  assign n6612 = ~reg_controllable_hgrant4_out & ~n6611;
  assign n6613 = ~reg_controllable_hgrant5_out & ~n6612;
  assign n6614 = ~reg_controllable_hgrant5_out & ~n6613;
  assign n6615 = next_sys_fair<0>_out  & ~n6614;
  assign n6616 = reg_controllable_hmastlock_out & ~n1324;
  assign n6617 = reg_controllable_locked_out & ~n6616;
  assign n6618 = ~reg_controllable_hmastlock_out & ~n1323;
  assign n6619 = ~n275 & ~n6618;
  assign n6620 = ~reg_controllable_locked_out & ~n6619;
  assign n6621 = ~n6617 & ~n6620;
  assign n6622 = ~reg_controllable_hgrant2_out & ~n6621;
  assign n6623 = ~reg_controllable_hgrant2_out & ~n6622;
  assign n6624 = ~reg_controllable_hgrant1_out & ~n6623;
  assign n6625 = ~reg_controllable_hgrant1_out & ~n6624;
  assign n6626 = ~reg_controllable_hgrant3_out & ~n6625;
  assign n6627 = ~reg_controllable_hgrant3_out & ~n6626;
  assign n6628 = ~next_sys_fair<2>_out  & ~n6627;
  assign n6629 = ~next_sys_fair<2>_out  & ~n6628;
  assign n6630 = ~reg_controllable_hgrant4_out & ~n6629;
  assign n6631 = ~reg_controllable_hgrant4_out & ~n6630;
  assign n6632 = ~reg_controllable_hgrant5_out & ~n6631;
  assign n6633 = ~reg_controllable_hgrant5_out & ~n6632;
  assign n6634 = ~next_sys_fair<0>_out  & ~n6633;
  assign n6635 = ~n6615 & ~n6634;
  assign n6636 = next_sys_fair<3>_out  & ~n6635;
  assign n6637 = ~reg_controllable_hgrant4_out & ~n6627;
  assign n6638 = ~reg_controllable_hgrant4_out & ~n6637;
  assign n6639 = ~reg_controllable_hgrant5_out & ~n6638;
  assign n6640 = ~reg_controllable_hgrant5_out & ~n6639;
  assign n6641 = next_sys_fair<0>_out  & ~n6640;
  assign n6642 = next_sys_fair<2>_out  & ~n6627;
  assign n6643 = ~n2981 & ~n3087;
  assign n6644 = ~reg_controllable_hgrant2_out & ~n6643;
  assign n6645 = ~reg_controllable_hgrant2_out & ~n6644;
  assign n6646 = ~reg_controllable_hgrant1_out & ~n6645;
  assign n6647 = ~reg_controllable_hgrant1_out & ~n6646;
  assign n6648 = ~reg_controllable_hgrant3_out & ~n6647;
  assign n6649 = ~reg_controllable_hgrant3_out & ~n6648;
  assign n6650 = ~next_sys_fair<2>_out  & ~n6649;
  assign n6651 = ~n6642 & ~n6650;
  assign n6652 = ~reg_controllable_hgrant4_out & ~n6651;
  assign n6653 = ~reg_controllable_hgrant4_out & ~n6652;
  assign n6654 = ~reg_controllable_hgrant5_out & ~n6653;
  assign n6655 = ~reg_controllable_hgrant5_out & ~n6654;
  assign n6656 = ~next_sys_fair<0>_out  & ~n6655;
  assign n6657 = ~n6641 & ~n6656;
  assign n6658 = ~next_sys_fair<3>_out  & ~n6657;
  assign n6659 = ~n6636 & ~n6658;
  assign n6660 = ~reg_controllable_hmaster2_out & ~n6659;
  assign n6661 = ~n6601 & ~n6660;
  assign n6662 = ~reg_controllable_hmaster1_out & ~n6661;
  assign n6663 = ~n6600 & ~n6662;
  assign n6664 = next_sys_fair<1>_out  & ~n6663;
  assign n6665 = next_sys_fair<3>_out  & ~n6581;
  assign n6666 = ~n2875 & ~n6590;
  assign n6667 = ~reg_controllable_hgrant4_out & ~n6666;
  assign n6668 = ~reg_controllable_hgrant4_out & ~n6667;
  assign n6669 = ~reg_controllable_hgrant5_out & ~n6668;
  assign n6670 = ~reg_controllable_hgrant5_out & ~n6669;
  assign n6671 = ~next_sys_fair<3>_out  & ~n6670;
  assign n6672 = ~n6665 & ~n6671;
  assign n6673 = reg_controllable_hmaster1_out & ~n6672;
  assign n6674 = reg_controllable_hmaster2_out & ~n6672;
  assign n6675 = next_sys_fair<3>_out  & ~n6633;
  assign n6676 = ~n3175 & ~n3257;
  assign n6677 = ~reg_controllable_hgrant2_out & ~n6676;
  assign n6678 = ~reg_controllable_hgrant2_out & ~n6677;
  assign n6679 = ~reg_controllable_hgrant1_out & ~n6678;
  assign n6680 = ~reg_controllable_hgrant1_out & ~n6679;
  assign n6681 = ~reg_controllable_hgrant3_out & ~n6680;
  assign n6682 = ~reg_controllable_hgrant3_out & ~n6681;
  assign n6683 = ~next_sys_fair<2>_out  & ~n6682;
  assign n6684 = ~n6642 & ~n6683;
  assign n6685 = ~reg_controllable_hgrant4_out & ~n6684;
  assign n6686 = ~reg_controllable_hgrant4_out & ~n6685;
  assign n6687 = ~reg_controllable_hgrant5_out & ~n6686;
  assign n6688 = ~reg_controllable_hgrant5_out & ~n6687;
  assign n6689 = next_sys_fair<0>_out  & ~n6688;
  assign n6690 = ~n6609 & ~n6642;
  assign n6691 = ~reg_controllable_hgrant4_out & ~n6690;
  assign n6692 = ~reg_controllable_hgrant4_out & ~n6691;
  assign n6693 = ~reg_controllable_hgrant5_out & ~n6692;
  assign n6694 = ~reg_controllable_hgrant5_out & ~n6693;
  assign n6695 = ~next_sys_fair<0>_out  & ~n6694;
  assign n6696 = ~n6689 & ~n6695;
  assign n6697 = ~next_sys_fair<3>_out  & ~n6696;
  assign n6698 = ~n6675 & ~n6697;
  assign n6699 = ~reg_controllable_hmaster2_out & ~n6698;
  assign n6700 = ~n6674 & ~n6699;
  assign n6701 = ~reg_controllable_hmaster1_out & ~n6700;
  assign n6702 = ~n6673 & ~n6701;
  assign n6703 = ~next_sys_fair<1>_out  & ~n6702;
  assign n6704 = ~n6664 & ~n6703;
  assign n6705 = reg_controllable_hmaster0_out & ~n6704;
  assign n6706 = next_sys_fair<1>_out  & ~n6599;
  assign n6707 = ~next_sys_fair<1>_out  & ~n6672;
  assign n6708 = ~n6706 & ~n6707;
  assign n6709 = ~reg_controllable_hmaster0_out & ~n6708;
  assign n6710 = ~n6705 & ~n6709;
  assign n6711 = reg_controllable_hmaster3_out & ~n6710;
  assign n6712 = ~reg_controllable_hmaster3_out & ~n6708;
  assign n6713 = ~n6711 & ~n6712;
  assign n6714 = ~reg_controllable_hgrant6_out & ~n6713;
  assign n6715 = ~reg_controllable_hgrant6_out & ~n6714;
  assign n6716 = ~reg_controllable_hgrant8_out & ~n6715;
  assign n6717 = ~reg_controllable_hgrant8_out & ~n6716;
  assign n6718 = ~reg_controllable_hgrant7_out & ~n6717;
  assign n6719 = ~reg_controllable_hgrant7_out & ~n6718;
  assign n6720 = reg_controllable_hgrant9_out & ~n6719;
  assign n6721 = ~n6598 & ~n6665;
  assign n6722 = next_sys_fair<1>_out  & ~n6721;
  assign n6723 = ~n6584 & ~n6671;
  assign n6724 = ~next_sys_fair<1>_out  & ~n6723;
  assign n6725 = ~n6722 & ~n6724;
  assign n6726 = reg_controllable_hmaster3_out & ~n6725;
  assign n6727 = ~n6658 & ~n6675;
  assign n6728 = reg_controllable_hmaster2_out & ~n6727;
  assign n6729 = ~reg_controllable_hmaster2_out & ~n6721;
  assign n6730 = ~n6728 & ~n6729;
  assign n6731 = reg_controllable_hmaster1_out & ~n6730;
  assign n6732 = ~reg_controllable_hmaster1_out & ~n6721;
  assign n6733 = ~n6731 & ~n6732;
  assign n6734 = next_sys_fair<1>_out  & ~n6733;
  assign n6735 = ~n6636 & ~n6697;
  assign n6736 = reg_controllable_hmaster2_out & ~n6735;
  assign n6737 = ~reg_controllable_hmaster2_out & ~n6723;
  assign n6738 = ~n6736 & ~n6737;
  assign n6739 = reg_controllable_hmaster1_out & ~n6738;
  assign n6740 = ~reg_controllable_hmaster1_out & ~n6723;
  assign n6741 = ~n6739 & ~n6740;
  assign n6742 = ~next_sys_fair<1>_out  & ~n6741;
  assign n6743 = ~n6734 & ~n6742;
  assign n6744 = reg_controllable_hmaster0_out & ~n6743;
  assign n6745 = ~reg_controllable_hmaster0_out & ~n6725;
  assign n6746 = ~n6744 & ~n6745;
  assign n6747 = ~reg_controllable_hmaster3_out & ~n6746;
  assign n6748 = ~n6726 & ~n6747;
  assign n6749 = ~reg_controllable_hgrant6_out & ~n6748;
  assign n6750 = ~reg_controllable_hgrant6_out & ~n6749;
  assign n6751 = ~reg_controllable_hgrant8_out & ~n6750;
  assign n6752 = ~reg_controllable_hgrant8_out & ~n6751;
  assign n6753 = reg_controllable_hgrant7_out & ~n6752;
  assign n6754 = next_sys_fair<0>_out  & ~n6581;
  assign n6755 = ~n3451 & ~n6754;
  assign n6756 = next_sys_fair<3>_out  & ~n6755;
  assign n6757 = ~n6598 & ~n6756;
  assign n6758 = next_sys_fair<1>_out  & ~n6757;
  assign n6759 = ~n6707 & ~n6758;
  assign n6760 = reg_controllable_hmaster0_out & ~n6759;
  assign n6761 = reg_controllable_hmaster1_out & ~n6757;
  assign n6762 = reg_controllable_hmaster2_out & ~n6757;
  assign n6763 = next_sys_fair<0>_out  & ~n6633;
  assign n6764 = ~next_sys_fair<0>_out  & ~n6614;
  assign n6765 = ~n6763 & ~n6764;
  assign n6766 = next_sys_fair<3>_out  & ~n6765;
  assign n6767 = ~n6658 & ~n6766;
  assign n6768 = ~reg_controllable_hmaster2_out & ~n6767;
  assign n6769 = ~n6762 & ~n6768;
  assign n6770 = ~reg_controllable_hmaster1_out & ~n6769;
  assign n6771 = ~n6761 & ~n6770;
  assign n6772 = next_sys_fair<1>_out  & ~n6771;
  assign n6773 = ~n6703 & ~n6772;
  assign n6774 = ~reg_controllable_hmaster0_out & ~n6773;
  assign n6775 = ~n6760 & ~n6774;
  assign n6776 = reg_controllable_hmaster3_out & ~n6775;
  assign n6777 = ~reg_controllable_hmaster3_out & ~n6759;
  assign n6778 = ~n6776 & ~n6777;
  assign n6779 = ~reg_controllable_hgrant6_out & ~n6778;
  assign n6780 = ~reg_controllable_hgrant6_out & ~n6779;
  assign n6781 = reg_controllable_hgrant8_out & ~n6780;
  assign n6782 = ~n6671 & ~n6756;
  assign n6783 = ~next_sys_fair<1>_out  & ~n6782;
  assign n6784 = ~n6722 & ~n6783;
  assign n6785 = reg_controllable_hmaster3_out & ~n6784;
  assign n6786 = reg_controllable_hmaster0_out & ~n6784;
  assign n6787 = ~n6697 & ~n6766;
  assign n6788 = reg_controllable_hmaster2_out & ~n6787;
  assign n6789 = ~reg_controllable_hmaster2_out & ~n6782;
  assign n6790 = ~n6788 & ~n6789;
  assign n6791 = reg_controllable_hmaster1_out & ~n6790;
  assign n6792 = ~reg_controllable_hmaster1_out & ~n6782;
  assign n6793 = ~n6791 & ~n6792;
  assign n6794 = ~next_sys_fair<1>_out  & ~n6793;
  assign n6795 = ~n6734 & ~n6794;
  assign n6796 = ~reg_controllable_hmaster0_out & ~n6795;
  assign n6797 = ~n6786 & ~n6796;
  assign n6798 = ~reg_controllable_hmaster3_out & ~n6797;
  assign n6799 = ~n6785 & ~n6798;
  assign n6800 = reg_controllable_hgrant6_out & ~n6799;
  assign n6801 = reg_controllable_hgrant5_out & ~n6579;
  assign n6802 = reg_controllable_hgrant4_out & ~n6577;
  assign n6803 = reg_controllable_hgrant3_out & ~n6573;
  assign n6804 = reg_controllable_hgrant1_out & ~n6571;
  assign n6805 = reg_controllable_hgrant2_out & ~n6569;
  assign n6806 = reg_controllable_hmastlock_out & ~n1259;
  assign n6807 = reg_controllable_hmastlock_out & ~n6806;
  assign n6808 = reg_controllable_locked_out & ~n6807;
  assign n6809 = ~reg_controllable_hmastlock_out & ~n1259;
  assign n6810 = ~n275 & ~n6809;
  assign n6811 = ~reg_controllable_locked_out & ~n6810;
  assign n6812 = ~n6808 & ~n6811;
  assign n6813 = ~reg_controllable_hgrant2_out & ~n6812;
  assign n6814 = ~n6805 & ~n6813;
  assign n6815 = ~reg_controllable_hgrant1_out & ~n6814;
  assign n6816 = ~n6804 & ~n6815;
  assign n6817 = ~reg_controllable_hgrant3_out & ~n6816;
  assign n6818 = ~n6803 & ~n6817;
  assign n6819 = ~next_sys_fair<2>_out  & ~n6818;
  assign n6820 = ~next_sys_fair<2>_out  & ~n6819;
  assign n6821 = ~reg_controllable_hgrant4_out & ~n6820;
  assign n6822 = ~n6802 & ~n6821;
  assign n6823 = ~reg_controllable_hgrant5_out & ~n6822;
  assign n6824 = ~n6801 & ~n6823;
  assign n6825 = next_sys_fair<3>_out  & ~n6824;
  assign n6826 = ~n3683 & ~n6576;
  assign n6827 = ~reg_controllable_hgrant4_out & ~n6826;
  assign n6828 = ~reg_controllable_hgrant4_out & ~n6827;
  assign n6829 = reg_controllable_hgrant5_out & ~n6828;
  assign n6830 = reg_controllable_hgrant4_out & ~n6575;
  assign n6831 = next_sys_fair<2>_out  & ~n6818;
  assign n6832 = reg_controllable_hgrant1_out & ~n2870;
  assign n6833 = ~n6815 & ~n6832;
  assign n6834 = ~reg_controllable_hgrant3_out & ~n6833;
  assign n6835 = ~n6803 & ~n6834;
  assign n6836 = ~next_sys_fair<2>_out  & ~n6835;
  assign n6837 = ~n6831 & ~n6836;
  assign n6838 = ~reg_controllable_hgrant4_out & ~n6837;
  assign n6839 = ~n6830 & ~n6838;
  assign n6840 = ~reg_controllable_hgrant5_out & ~n6839;
  assign n6841 = ~n6829 & ~n6840;
  assign n6842 = next_sys_fair<0>_out  & ~n6841;
  assign n6843 = reg_controllable_hgrant5_out & ~n6593;
  assign n6844 = reg_controllable_hgrant4_out & ~n3684;
  assign n6845 = reg_controllable_hgrant3_out & ~n2891;
  assign n6846 = reg_controllable_hgrant1_out & ~n2889;
  assign n6847 = reg_controllable_hgrant2_out & ~n2887;
  assign n6848 = reg_controllable_hmastlock_out & ~n1228;
  assign n6849 = reg_controllable_hmastlock_out & ~n6848;
  assign n6850 = reg_controllable_locked_out & ~n6849;
  assign n6851 = ~n5800 & ~n6850;
  assign n6852 = ~reg_controllable_hgrant2_out & ~n6851;
  assign n6853 = ~n6847 & ~n6852;
  assign n6854 = ~reg_controllable_hgrant1_out & ~n6853;
  assign n6855 = ~n6846 & ~n6854;
  assign n6856 = ~reg_controllable_hgrant3_out & ~n6855;
  assign n6857 = ~n6845 & ~n6856;
  assign n6858 = ~next_sys_fair<2>_out  & ~n6857;
  assign n6859 = ~n6831 & ~n6858;
  assign n6860 = ~reg_controllable_hgrant4_out & ~n6859;
  assign n6861 = ~n6844 & ~n6860;
  assign n6862 = ~reg_controllable_hgrant5_out & ~n6861;
  assign n6863 = ~n6843 & ~n6862;
  assign n6864 = ~next_sys_fair<0>_out  & ~n6863;
  assign n6865 = ~n6842 & ~n6864;
  assign n6866 = ~next_sys_fair<3>_out  & ~n6865;
  assign n6867 = ~n6825 & ~n6866;
  assign n6868 = reg_controllable_hmaster1_out & ~n6867;
  assign n6869 = reg_controllable_hmaster2_out & ~n6867;
  assign n6870 = ~reg_controllable_hgrant1_out & ~n6569;
  assign n6871 = ~n6804 & ~n6870;
  assign n6872 = ~reg_controllable_hgrant3_out & ~n6871;
  assign n6873 = ~n6803 & ~n6872;
  assign n6874 = ~next_sys_fair<2>_out  & ~n6873;
  assign n6875 = ~next_sys_fair<2>_out  & ~n6874;
  assign n6876 = ~reg_controllable_hgrant4_out & ~n6875;
  assign n6877 = ~n6802 & ~n6876;
  assign n6878 = ~reg_controllable_hgrant5_out & ~n6877;
  assign n6879 = ~n6801 & ~n6878;
  assign n6880 = next_sys_fair<3>_out  & ~n6879;
  assign n6881 = next_sys_fair<2>_out  & ~n6873;
  assign n6882 = ~n6832 & ~n6870;
  assign n6883 = ~reg_controllable_hgrant3_out & ~n6882;
  assign n6884 = ~n6803 & ~n6883;
  assign n6885 = ~next_sys_fair<2>_out  & ~n6884;
  assign n6886 = ~n6881 & ~n6885;
  assign n6887 = ~reg_controllable_hgrant4_out & ~n6886;
  assign n6888 = ~n6830 & ~n6887;
  assign n6889 = ~reg_controllable_hgrant5_out & ~n6888;
  assign n6890 = ~n6829 & ~n6889;
  assign n6891 = next_sys_fair<0>_out  & ~n6890;
  assign n6892 = ~n5848 & ~n6847;
  assign n6893 = ~reg_controllable_hgrant1_out & ~n6892;
  assign n6894 = ~n6846 & ~n6893;
  assign n6895 = ~reg_controllable_hgrant3_out & ~n6894;
  assign n6896 = ~n6845 & ~n6895;
  assign n6897 = ~next_sys_fair<2>_out  & ~n6896;
  assign n6898 = ~n6881 & ~n6897;
  assign n6899 = ~reg_controllable_hgrant4_out & ~n6898;
  assign n6900 = ~n6844 & ~n6899;
  assign n6901 = ~reg_controllable_hgrant5_out & ~n6900;
  assign n6902 = ~n6843 & ~n6901;
  assign n6903 = ~next_sys_fair<0>_out  & ~n6902;
  assign n6904 = ~n6891 & ~n6903;
  assign n6905 = ~next_sys_fair<3>_out  & ~n6904;
  assign n6906 = ~n6880 & ~n6905;
  assign n6907 = ~reg_controllable_hmaster2_out & ~n6906;
  assign n6908 = ~n6869 & ~n6907;
  assign n6909 = ~reg_controllable_hmaster1_out & ~n6908;
  assign n6910 = ~n6868 & ~n6909;
  assign n6911 = next_sys_fair<1>_out  & ~n6910;
  assign n6912 = reg_controllable_hgrant5_out & ~n6668;
  assign n6913 = reg_controllable_hgrant4_out & ~n6666;
  assign n6914 = reg_controllable_hgrant3_out & ~n2872;
  assign n6915 = ~n6817 & ~n6914;
  assign n6916 = next_sys_fair<2>_out  & ~n6915;
  assign n6917 = reg_controllable_hgrant2_out & ~n2868;
  assign n6918 = reg_controllable_hmastlock_out & ~n1367;
  assign n6919 = reg_controllable_hmastlock_out & ~n6918;
  assign n6920 = reg_controllable_locked_out & ~n6919;
  assign n6921 = ~n5878 & ~n6920;
  assign n6922 = ~reg_controllable_hgrant2_out & ~n6921;
  assign n6923 = ~n6917 & ~n6922;
  assign n6924 = ~reg_controllable_hgrant1_out & ~n6923;
  assign n6925 = ~n6832 & ~n6924;
  assign n6926 = ~reg_controllable_hgrant3_out & ~n6925;
  assign n6927 = ~n6914 & ~n6926;
  assign n6928 = ~next_sys_fair<2>_out  & ~n6927;
  assign n6929 = ~n6916 & ~n6928;
  assign n6930 = ~reg_controllable_hgrant4_out & ~n6929;
  assign n6931 = ~n6913 & ~n6930;
  assign n6932 = ~reg_controllable_hgrant5_out & ~n6931;
  assign n6933 = ~n6912 & ~n6932;
  assign n6934 = next_sys_fair<0>_out  & ~n6933;
  assign n6935 = ~n6813 & ~n6917;
  assign n6936 = ~reg_controllable_hgrant1_out & ~n6935;
  assign n6937 = ~n6804 & ~n6936;
  assign n6938 = ~reg_controllable_hgrant3_out & ~n6937;
  assign n6939 = ~n6803 & ~n6938;
  assign n6940 = next_sys_fair<2>_out  & ~n6939;
  assign n6941 = reg_controllable_hmastlock_out & ~n1389;
  assign n6942 = reg_controllable_hmastlock_out & ~n6941;
  assign n6943 = reg_controllable_locked_out & ~n6942;
  assign n6944 = ~n5902 & ~n6943;
  assign n6945 = ~reg_controllable_hgrant2_out & ~n6944;
  assign n6946 = ~n6917 & ~n6945;
  assign n6947 = ~reg_controllable_hgrant1_out & ~n6946;
  assign n6948 = ~n6832 & ~n6947;
  assign n6949 = ~reg_controllable_hgrant3_out & ~n6948;
  assign n6950 = ~n6914 & ~n6949;
  assign n6951 = ~next_sys_fair<2>_out  & ~n6950;
  assign n6952 = ~n6940 & ~n6951;
  assign n6953 = ~reg_controllable_hgrant4_out & ~n6952;
  assign n6954 = ~n6913 & ~n6953;
  assign n6955 = ~reg_controllable_hgrant5_out & ~n6954;
  assign n6956 = ~n6912 & ~n6955;
  assign n6957 = ~next_sys_fair<0>_out  & ~n6956;
  assign n6958 = ~n6934 & ~n6957;
  assign n6959 = ~next_sys_fair<3>_out  & ~n6958;
  assign n6960 = ~n6825 & ~n6959;
  assign n6961 = reg_controllable_hmaster1_out & ~n6960;
  assign n6962 = reg_controllable_hmaster2_out & ~n6960;
  assign n6963 = ~n6872 & ~n6914;
  assign n6964 = next_sys_fair<2>_out  & ~n6963;
  assign n6965 = ~reg_controllable_hgrant1_out & ~n2868;
  assign n6966 = ~n6832 & ~n6965;
  assign n6967 = ~reg_controllable_hgrant3_out & ~n6966;
  assign n6968 = ~n6914 & ~n6967;
  assign n6969 = ~next_sys_fair<2>_out  & ~n6968;
  assign n6970 = ~n6964 & ~n6969;
  assign n6971 = ~reg_controllable_hgrant4_out & ~n6970;
  assign n6972 = ~n6913 & ~n6971;
  assign n6973 = ~reg_controllable_hgrant5_out & ~n6972;
  assign n6974 = ~n6912 & ~n6973;
  assign n6975 = next_sys_fair<0>_out  & ~n6974;
  assign n6976 = ~n6570 & ~n6917;
  assign n6977 = ~reg_controllable_hgrant1_out & ~n6976;
  assign n6978 = ~n6804 & ~n6977;
  assign n6979 = ~reg_controllable_hgrant3_out & ~n6978;
  assign n6980 = ~n6803 & ~n6979;
  assign n6981 = next_sys_fair<2>_out  & ~n6980;
  assign n6982 = ~n6969 & ~n6981;
  assign n6983 = ~reg_controllable_hgrant4_out & ~n6982;
  assign n6984 = ~n6913 & ~n6983;
  assign n6985 = ~reg_controllable_hgrant5_out & ~n6984;
  assign n6986 = ~n6912 & ~n6985;
  assign n6987 = ~next_sys_fair<0>_out  & ~n6986;
  assign n6988 = ~n6975 & ~n6987;
  assign n6989 = ~next_sys_fair<3>_out  & ~n6988;
  assign n6990 = ~n6880 & ~n6989;
  assign n6991 = ~reg_controllable_hmaster2_out & ~n6990;
  assign n6992 = ~n6962 & ~n6991;
  assign n6993 = ~reg_controllable_hmaster1_out & ~n6992;
  assign n6994 = ~n6961 & ~n6993;
  assign n6995 = ~next_sys_fair<1>_out  & ~n6994;
  assign n6996 = ~n6911 & ~n6995;
  assign n6997 = reg_controllable_hmaster3_out & ~n6996;
  assign n6998 = reg_controllable_hmaster2_out & ~n6906;
  assign n6999 = reg_controllable_hgrant3_out & ~n6625;
  assign n7000 = ~n6872 & ~n6999;
  assign n7001 = ~next_sys_fair<2>_out  & ~n7000;
  assign n7002 = ~next_sys_fair<2>_out  & ~n7001;
  assign n7003 = ~reg_controllable_hgrant4_out & ~n7002;
  assign n7004 = ~n6802 & ~n7003;
  assign n7005 = ~reg_controllable_hgrant5_out & ~n7004;
  assign n7006 = ~n6801 & ~n7005;
  assign n7007 = next_sys_fair<3>_out  & ~n7006;
  assign n7008 = next_sys_fair<2>_out  & ~n7000;
  assign n7009 = ~n6883 & ~n6999;
  assign n7010 = ~next_sys_fair<2>_out  & ~n7009;
  assign n7011 = ~n7008 & ~n7010;
  assign n7012 = ~reg_controllable_hgrant4_out & ~n7011;
  assign n7013 = ~n6830 & ~n7012;
  assign n7014 = ~reg_controllable_hgrant5_out & ~n7013;
  assign n7015 = ~n6829 & ~n7014;
  assign n7016 = next_sys_fair<0>_out  & ~n7015;
  assign n7017 = reg_controllable_hgrant3_out & ~n6647;
  assign n7018 = ~n6895 & ~n7017;
  assign n7019 = ~next_sys_fair<2>_out  & ~n7018;
  assign n7020 = ~n7008 & ~n7019;
  assign n7021 = ~reg_controllable_hgrant4_out & ~n7020;
  assign n7022 = ~n6844 & ~n7021;
  assign n7023 = ~reg_controllable_hgrant5_out & ~n7022;
  assign n7024 = ~n6843 & ~n7023;
  assign n7025 = ~next_sys_fair<0>_out  & ~n7024;
  assign n7026 = ~n7016 & ~n7025;
  assign n7027 = ~next_sys_fair<3>_out  & ~n7026;
  assign n7028 = ~n7007 & ~n7027;
  assign n7029 = ~reg_controllable_hmaster2_out & ~n7028;
  assign n7030 = ~n6998 & ~n7029;
  assign n7031 = reg_controllable_hmaster1_out & ~n7030;
  assign n7032 = reg_controllable_hgrant5_out & ~n6631;
  assign n7033 = ~n6878 & ~n7032;
  assign n7034 = next_sys_fair<3>_out  & ~n7033;
  assign n7035 = next_sys_fair<2>_out  & ~n6608;
  assign n7036 = ~n6628 & ~n7035;
  assign n7037 = ~reg_controllable_hgrant4_out & ~n7036;
  assign n7038 = ~reg_controllable_hgrant4_out & ~n7037;
  assign n7039 = reg_controllable_hgrant5_out & ~n7038;
  assign n7040 = ~n6889 & ~n7039;
  assign n7041 = next_sys_fair<0>_out  & ~n7040;
  assign n7042 = reg_controllable_hgrant5_out & ~n6653;
  assign n7043 = ~n6901 & ~n7042;
  assign n7044 = ~next_sys_fair<0>_out  & ~n7043;
  assign n7045 = ~n7041 & ~n7044;
  assign n7046 = ~next_sys_fair<3>_out  & ~n7045;
  assign n7047 = ~n7034 & ~n7046;
  assign n7048 = reg_controllable_hmaster2_out & ~n7047;
  assign n7049 = reg_controllable_hgrant1_out & ~n6623;
  assign n7050 = ~n6870 & ~n7049;
  assign n7051 = ~reg_controllable_hgrant3_out & ~n7050;
  assign n7052 = ~n6803 & ~n7051;
  assign n7053 = ~next_sys_fair<2>_out  & ~n7052;
  assign n7054 = ~next_sys_fair<2>_out  & ~n7053;
  assign n7055 = ~reg_controllable_hgrant4_out & ~n7054;
  assign n7056 = ~n6802 & ~n7055;
  assign n7057 = ~reg_controllable_hgrant5_out & ~n7056;
  assign n7058 = ~n6801 & ~n7057;
  assign n7059 = next_sys_fair<3>_out  & ~n7058;
  assign n7060 = next_sys_fair<2>_out  & ~n7052;
  assign n7061 = reg_controllable_hgrant1_out & ~n6604;
  assign n7062 = ~n6870 & ~n7061;
  assign n7063 = ~reg_controllable_hgrant3_out & ~n7062;
  assign n7064 = ~n6803 & ~n7063;
  assign n7065 = ~next_sys_fair<2>_out  & ~n7064;
  assign n7066 = ~n7060 & ~n7065;
  assign n7067 = ~reg_controllable_hgrant4_out & ~n7066;
  assign n7068 = ~n6830 & ~n7067;
  assign n7069 = ~reg_controllable_hgrant5_out & ~n7068;
  assign n7070 = ~n6829 & ~n7069;
  assign n7071 = next_sys_fair<0>_out  & ~n7070;
  assign n7072 = reg_controllable_hgrant1_out & ~n6645;
  assign n7073 = ~n6893 & ~n7072;
  assign n7074 = ~reg_controllable_hgrant3_out & ~n7073;
  assign n7075 = ~n6845 & ~n7074;
  assign n7076 = ~next_sys_fair<2>_out  & ~n7075;
  assign n7077 = ~n7060 & ~n7076;
  assign n7078 = ~reg_controllable_hgrant4_out & ~n7077;
  assign n7079 = ~n6844 & ~n7078;
  assign n7080 = ~reg_controllable_hgrant5_out & ~n7079;
  assign n7081 = ~n6843 & ~n7080;
  assign n7082 = ~next_sys_fair<0>_out  & ~n7081;
  assign n7083 = ~n7071 & ~n7082;
  assign n7084 = ~next_sys_fair<3>_out  & ~n7083;
  assign n7085 = ~n7059 & ~n7084;
  assign n7086 = ~reg_controllable_hmaster2_out & ~n7085;
  assign n7087 = ~n7048 & ~n7086;
  assign n7088 = ~reg_controllable_hmaster1_out & ~n7087;
  assign n7089 = ~n7031 & ~n7088;
  assign n7090 = next_sys_fair<1>_out  & ~n7089;
  assign n7091 = reg_controllable_hmaster2_out & ~n6990;
  assign n7092 = reg_controllable_hgrant3_out & ~n6606;
  assign n7093 = ~n6872 & ~n7092;
  assign n7094 = next_sys_fair<2>_out  & ~n7093;
  assign n7095 = reg_controllable_hgrant3_out & ~n6680;
  assign n7096 = ~n6967 & ~n7095;
  assign n7097 = ~next_sys_fair<2>_out  & ~n7096;
  assign n7098 = ~n7094 & ~n7097;
  assign n7099 = ~reg_controllable_hgrant4_out & ~n7098;
  assign n7100 = ~n6913 & ~n7099;
  assign n7101 = ~reg_controllable_hgrant5_out & ~n7100;
  assign n7102 = ~n6912 & ~n7101;
  assign n7103 = next_sys_fair<0>_out  & ~n7102;
  assign n7104 = ~n6979 & ~n6999;
  assign n7105 = next_sys_fair<2>_out  & ~n7104;
  assign n7106 = ~n6967 & ~n7092;
  assign n7107 = ~next_sys_fair<2>_out  & ~n7106;
  assign n7108 = ~n7105 & ~n7107;
  assign n7109 = ~reg_controllable_hgrant4_out & ~n7108;
  assign n7110 = ~n6913 & ~n7109;
  assign n7111 = ~reg_controllable_hgrant5_out & ~n7110;
  assign n7112 = ~n6912 & ~n7111;
  assign n7113 = ~next_sys_fair<0>_out  & ~n7112;
  assign n7114 = ~n7103 & ~n7113;
  assign n7115 = ~next_sys_fair<3>_out  & ~n7114;
  assign n7116 = ~n7007 & ~n7115;
  assign n7117 = ~reg_controllable_hmaster2_out & ~n7116;
  assign n7118 = ~n7091 & ~n7117;
  assign n7119 = reg_controllable_hmaster1_out & ~n7118;
  assign n7120 = reg_controllable_hgrant5_out & ~n6686;
  assign n7121 = ~n6973 & ~n7120;
  assign n7122 = next_sys_fair<0>_out  & ~n7121;
  assign n7123 = reg_controllable_hgrant5_out & ~n6692;
  assign n7124 = ~n6985 & ~n7123;
  assign n7125 = ~next_sys_fair<0>_out  & ~n7124;
  assign n7126 = ~n7122 & ~n7125;
  assign n7127 = ~next_sys_fair<3>_out  & ~n7126;
  assign n7128 = ~n7034 & ~n7127;
  assign n7129 = reg_controllable_hmaster2_out & ~n7128;
  assign n7130 = ~n6914 & ~n7051;
  assign n7131 = next_sys_fair<2>_out  & ~n7130;
  assign n7132 = reg_controllable_hgrant1_out & ~n6678;
  assign n7133 = ~n6965 & ~n7132;
  assign n7134 = ~reg_controllable_hgrant3_out & ~n7133;
  assign n7135 = ~n6914 & ~n7134;
  assign n7136 = ~next_sys_fair<2>_out  & ~n7135;
  assign n7137 = ~n7131 & ~n7136;
  assign n7138 = ~reg_controllable_hgrant4_out & ~n7137;
  assign n7139 = ~n6913 & ~n7138;
  assign n7140 = ~reg_controllable_hgrant5_out & ~n7139;
  assign n7141 = ~n6912 & ~n7140;
  assign n7142 = next_sys_fair<0>_out  & ~n7141;
  assign n7143 = ~n6977 & ~n7049;
  assign n7144 = ~reg_controllable_hgrant3_out & ~n7143;
  assign n7145 = ~n6803 & ~n7144;
  assign n7146 = next_sys_fair<2>_out  & ~n7145;
  assign n7147 = ~n6965 & ~n7061;
  assign n7148 = ~reg_controllable_hgrant3_out & ~n7147;
  assign n7149 = ~n6914 & ~n7148;
  assign n7150 = ~next_sys_fair<2>_out  & ~n7149;
  assign n7151 = ~n7146 & ~n7150;
  assign n7152 = ~reg_controllable_hgrant4_out & ~n7151;
  assign n7153 = ~n6913 & ~n7152;
  assign n7154 = ~reg_controllable_hgrant5_out & ~n7153;
  assign n7155 = ~n6912 & ~n7154;
  assign n7156 = ~next_sys_fair<0>_out  & ~n7155;
  assign n7157 = ~n7142 & ~n7156;
  assign n7158 = ~next_sys_fair<3>_out  & ~n7157;
  assign n7159 = ~n7059 & ~n7158;
  assign n7160 = ~reg_controllable_hmaster2_out & ~n7159;
  assign n7161 = ~n7129 & ~n7160;
  assign n7162 = ~reg_controllable_hmaster1_out & ~n7161;
  assign n7163 = ~n7119 & ~n7162;
  assign n7164 = ~next_sys_fair<1>_out  & ~n7163;
  assign n7165 = ~n7090 & ~n7164;
  assign n7166 = reg_controllable_hmaster0_out & ~n7165;
  assign n7167 = reg_controllable_hgrant2_out & ~n6621;
  assign n7168 = ~n6570 & ~n7167;
  assign n7169 = ~reg_controllable_hgrant1_out & ~n7168;
  assign n7170 = ~n6804 & ~n7169;
  assign n7171 = ~reg_controllable_hgrant3_out & ~n7170;
  assign n7172 = ~n6803 & ~n7171;
  assign n7173 = ~next_sys_fair<2>_out  & ~n7172;
  assign n7174 = ~next_sys_fair<2>_out  & ~n7173;
  assign n7175 = ~reg_controllable_hgrant4_out & ~n7174;
  assign n7176 = ~n6802 & ~n7175;
  assign n7177 = ~reg_controllable_hgrant5_out & ~n7176;
  assign n7178 = ~n6801 & ~n7177;
  assign n7179 = next_sys_fair<3>_out  & ~n7178;
  assign n7180 = next_sys_fair<2>_out  & ~n7172;
  assign n7181 = ~n6832 & ~n7169;
  assign n7182 = ~reg_controllable_hgrant3_out & ~n7181;
  assign n7183 = ~n6803 & ~n7182;
  assign n7184 = ~next_sys_fair<2>_out  & ~n7183;
  assign n7185 = ~n7180 & ~n7184;
  assign n7186 = ~reg_controllable_hgrant4_out & ~n7185;
  assign n7187 = ~n6830 & ~n7186;
  assign n7188 = ~reg_controllable_hgrant5_out & ~n7187;
  assign n7189 = ~n6829 & ~n7188;
  assign n7190 = next_sys_fair<0>_out  & ~n7189;
  assign n7191 = reg_controllable_hgrant2_out & ~n6643;
  assign n7192 = ~n5848 & ~n7191;
  assign n7193 = ~reg_controllable_hgrant1_out & ~n7192;
  assign n7194 = ~n6846 & ~n7193;
  assign n7195 = ~reg_controllable_hgrant3_out & ~n7194;
  assign n7196 = ~n6845 & ~n7195;
  assign n7197 = ~next_sys_fair<2>_out  & ~n7196;
  assign n7198 = ~n7180 & ~n7197;
  assign n7199 = ~reg_controllable_hgrant4_out & ~n7198;
  assign n7200 = ~n6844 & ~n7199;
  assign n7201 = ~reg_controllable_hgrant5_out & ~n7200;
  assign n7202 = ~n6843 & ~n7201;
  assign n7203 = ~next_sys_fair<0>_out  & ~n7202;
  assign n7204 = ~n7190 & ~n7203;
  assign n7205 = ~next_sys_fair<3>_out  & ~n7204;
  assign n7206 = ~n7179 & ~n7205;
  assign n7207 = ~reg_controllable_hmaster2_out & ~n7206;
  assign n7208 = ~n6998 & ~n7207;
  assign n7209 = reg_controllable_hmaster1_out & ~n7208;
  assign n7210 = reg_controllable_hgrant4_out & ~n6629;
  assign n7211 = ~n6876 & ~n7210;
  assign n7212 = ~reg_controllable_hgrant5_out & ~n7211;
  assign n7213 = ~n6801 & ~n7212;
  assign n7214 = next_sys_fair<3>_out  & ~n7213;
  assign n7215 = reg_controllable_hgrant4_out & ~n6627;
  assign n7216 = ~n6887 & ~n7215;
  assign n7217 = ~reg_controllable_hgrant5_out & ~n7216;
  assign n7218 = ~n6829 & ~n7217;
  assign n7219 = next_sys_fair<0>_out  & ~n7218;
  assign n7220 = ~n6650 & ~n7035;
  assign n7221 = reg_controllable_hgrant4_out & ~n7220;
  assign n7222 = ~n6899 & ~n7221;
  assign n7223 = ~reg_controllable_hgrant5_out & ~n7222;
  assign n7224 = ~n6843 & ~n7223;
  assign n7225 = ~next_sys_fair<0>_out  & ~n7224;
  assign n7226 = ~n7219 & ~n7225;
  assign n7227 = ~next_sys_fair<3>_out  & ~n7226;
  assign n7228 = ~n7214 & ~n7227;
  assign n7229 = reg_controllable_hmaster2_out & ~n7228;
  assign n7230 = ~n6907 & ~n7229;
  assign n7231 = ~reg_controllable_hmaster1_out & ~n7230;
  assign n7232 = ~n7209 & ~n7231;
  assign n7233 = next_sys_fair<1>_out  & ~n7232;
  assign n7234 = ~n6914 & ~n7171;
  assign n7235 = next_sys_fair<2>_out  & ~n7234;
  assign n7236 = reg_controllable_hgrant2_out & ~n6676;
  assign n7237 = ~n2869 & ~n7236;
  assign n7238 = ~reg_controllable_hgrant1_out & ~n7237;
  assign n7239 = ~n6832 & ~n7238;
  assign n7240 = ~reg_controllable_hgrant3_out & ~n7239;
  assign n7241 = ~n6914 & ~n7240;
  assign n7242 = ~next_sys_fair<2>_out  & ~n7241;
  assign n7243 = ~n7235 & ~n7242;
  assign n7244 = ~reg_controllable_hgrant4_out & ~n7243;
  assign n7245 = ~n6913 & ~n7244;
  assign n7246 = ~reg_controllable_hgrant5_out & ~n7245;
  assign n7247 = ~n6912 & ~n7246;
  assign n7248 = next_sys_fair<0>_out  & ~n7247;
  assign n7249 = reg_controllable_hgrant2_out & ~n6602;
  assign n7250 = ~n6570 & ~n7249;
  assign n7251 = ~reg_controllable_hgrant1_out & ~n7250;
  assign n7252 = ~n6804 & ~n7251;
  assign n7253 = ~reg_controllable_hgrant3_out & ~n7252;
  assign n7254 = ~n6803 & ~n7253;
  assign n7255 = next_sys_fair<2>_out  & ~n7254;
  assign n7256 = ~n2869 & ~n7249;
  assign n7257 = ~reg_controllable_hgrant1_out & ~n7256;
  assign n7258 = ~n6832 & ~n7257;
  assign n7259 = ~reg_controllable_hgrant3_out & ~n7258;
  assign n7260 = ~n6914 & ~n7259;
  assign n7261 = ~next_sys_fair<2>_out  & ~n7260;
  assign n7262 = ~n7255 & ~n7261;
  assign n7263 = ~reg_controllable_hgrant4_out & ~n7262;
  assign n7264 = ~n6913 & ~n7263;
  assign n7265 = ~reg_controllable_hgrant5_out & ~n7264;
  assign n7266 = ~n6912 & ~n7265;
  assign n7267 = ~next_sys_fair<0>_out  & ~n7266;
  assign n7268 = ~n7248 & ~n7267;
  assign n7269 = ~next_sys_fair<3>_out  & ~n7268;
  assign n7270 = ~n7179 & ~n7269;
  assign n7271 = ~reg_controllable_hmaster2_out & ~n7270;
  assign n7272 = ~n7091 & ~n7271;
  assign n7273 = reg_controllable_hmaster1_out & ~n7272;
  assign n7274 = reg_controllable_hgrant4_out & ~n6684;
  assign n7275 = ~n6971 & ~n7274;
  assign n7276 = ~reg_controllable_hgrant5_out & ~n7275;
  assign n7277 = ~n6912 & ~n7276;
  assign n7278 = next_sys_fair<0>_out  & ~n7277;
  assign n7279 = reg_controllable_hgrant4_out & ~n6690;
  assign n7280 = ~n6983 & ~n7279;
  assign n7281 = ~reg_controllable_hgrant5_out & ~n7280;
  assign n7282 = ~n6912 & ~n7281;
  assign n7283 = ~next_sys_fair<0>_out  & ~n7282;
  assign n7284 = ~n7278 & ~n7283;
  assign n7285 = ~next_sys_fair<3>_out  & ~n7284;
  assign n7286 = ~n7214 & ~n7285;
  assign n7287 = reg_controllable_hmaster2_out & ~n7286;
  assign n7288 = ~n6991 & ~n7287;
  assign n7289 = ~reg_controllable_hmaster1_out & ~n7288;
  assign n7290 = ~n7273 & ~n7289;
  assign n7291 = ~next_sys_fair<1>_out  & ~n7290;
  assign n7292 = ~n7233 & ~n7291;
  assign n7293 = ~reg_controllable_hmaster0_out & ~n7292;
  assign n7294 = ~n7166 & ~n7293;
  assign n7295 = ~reg_controllable_hmaster3_out & ~n7294;
  assign n7296 = ~n6997 & ~n7295;
  assign n7297 = ~reg_controllable_hgrant6_out & ~n7296;
  assign n7298 = ~n6800 & ~n7297;
  assign n7299 = ~reg_controllable_hgrant8_out & ~n7298;
  assign n7300 = ~n6781 & ~n7299;
  assign n7301 = ~reg_controllable_hgrant7_out & ~n7300;
  assign n7302 = ~n6753 & ~n7301;
  assign n7303 = ~reg_controllable_hgrant9_out & ~n7302;
  assign n7304 = ~n6720 & ~n7303;
  assign n7305 = reg_controllable_nhgrant0_out & ~n7304;
  assign n7306 = ~next_sys_fair<0>_out  & ~n6670;
  assign n7307 = ~n6589 & ~n7306;
  assign n7308 = ~next_sys_fair<3>_out  & ~n7307;
  assign n7309 = ~n6665 & ~n7308;
  assign n7310 = next_sys_fair<1>_out  & ~n7309;
  assign n7311 = ~n6707 & ~n7310;
  assign n7312 = reg_controllable_hmaster3_out & ~n7311;
  assign n7313 = reg_controllable_hmaster0_out & ~n7311;
  assign n7314 = reg_controllable_hmaster1_out & ~n7309;
  assign n7315 = reg_controllable_hmaster2_out & ~n7309;
  assign n7316 = ~n278 & ~n6617;
  assign n7317 = ~reg_controllable_hgrant2_out & ~n7316;
  assign n7318 = ~reg_controllable_hgrant2_out & ~n7317;
  assign n7319 = ~reg_controllable_hgrant1_out & ~n7318;
  assign n7320 = ~reg_controllable_hgrant1_out & ~n7319;
  assign n7321 = ~reg_controllable_hgrant3_out & ~n7320;
  assign n7322 = ~reg_controllable_hgrant3_out & ~n7321;
  assign n7323 = ~next_sys_fair<2>_out  & ~n7322;
  assign n7324 = ~next_sys_fair<2>_out  & ~n7323;
  assign n7325 = ~reg_controllable_hgrant4_out & ~n7324;
  assign n7326 = ~reg_controllable_hgrant4_out & ~n7325;
  assign n7327 = ~reg_controllable_hgrant5_out & ~n7326;
  assign n7328 = ~reg_controllable_hgrant5_out & ~n7327;
  assign n7329 = next_sys_fair<3>_out  & ~n7328;
  assign n7330 = ~reg_controllable_hgrant4_out & ~n7322;
  assign n7331 = ~reg_controllable_hgrant4_out & ~n7330;
  assign n7332 = ~reg_controllable_hgrant5_out & ~n7331;
  assign n7333 = ~reg_controllable_hgrant5_out & ~n7332;
  assign n7334 = next_sys_fair<0>_out  & ~n7333;
  assign n7335 = next_sys_fair<2>_out  & ~n7322;
  assign n7336 = ~n3076 & ~n7335;
  assign n7337 = ~reg_controllable_hgrant4_out & ~n7336;
  assign n7338 = ~reg_controllable_hgrant4_out & ~n7337;
  assign n7339 = ~reg_controllable_hgrant5_out & ~n7338;
  assign n7340 = ~reg_controllable_hgrant5_out & ~n7339;
  assign n7341 = ~next_sys_fair<0>_out  & ~n7340;
  assign n7342 = ~n7334 & ~n7341;
  assign n7343 = ~next_sys_fair<3>_out  & ~n7342;
  assign n7344 = ~n7329 & ~n7343;
  assign n7345 = ~reg_controllable_hmaster2_out & ~n7344;
  assign n7346 = ~n7315 & ~n7345;
  assign n7347 = ~reg_controllable_hmaster1_out & ~n7346;
  assign n7348 = ~n7314 & ~n7347;
  assign n7349 = next_sys_fair<1>_out  & ~n7348;
  assign n7350 = ~n3283 & ~n7335;
  assign n7351 = ~reg_controllable_hgrant4_out & ~n7350;
  assign n7352 = ~reg_controllable_hgrant4_out & ~n7351;
  assign n7353 = ~reg_controllable_hgrant5_out & ~n7352;
  assign n7354 = ~reg_controllable_hgrant5_out & ~n7353;
  assign n7355 = next_sys_fair<0>_out  & ~n7354;
  assign n7356 = ~n3316 & ~n7335;
  assign n7357 = ~reg_controllable_hgrant4_out & ~n7356;
  assign n7358 = ~reg_controllable_hgrant4_out & ~n7357;
  assign n7359 = ~reg_controllable_hgrant5_out & ~n7358;
  assign n7360 = ~reg_controllable_hgrant5_out & ~n7359;
  assign n7361 = ~next_sys_fair<0>_out  & ~n7360;
  assign n7362 = ~n7355 & ~n7361;
  assign n7363 = ~next_sys_fair<3>_out  & ~n7362;
  assign n7364 = ~n7329 & ~n7363;
  assign n7365 = ~reg_controllable_hmaster2_out & ~n7364;
  assign n7366 = ~n6674 & ~n7365;
  assign n7367 = ~reg_controllable_hmaster1_out & ~n7366;
  assign n7368 = ~n6673 & ~n7367;
  assign n7369 = ~next_sys_fair<1>_out  & ~n7368;
  assign n7370 = ~n7349 & ~n7369;
  assign n7371 = ~reg_controllable_hmaster0_out & ~n7370;
  assign n7372 = ~n7313 & ~n7371;
  assign n7373 = ~reg_controllable_hmaster3_out & ~n7372;
  assign n7374 = ~n7312 & ~n7373;
  assign n7375 = ~reg_controllable_hgrant6_out & ~n7374;
  assign n7376 = ~reg_controllable_hgrant6_out & ~n7375;
  assign n7377 = ~reg_controllable_hgrant8_out & ~n7376;
  assign n7378 = ~reg_controllable_hgrant8_out & ~n7377;
  assign n7379 = ~reg_controllable_hgrant7_out & ~n7378;
  assign n7380 = ~reg_controllable_hgrant7_out & ~n7379;
  assign n7381 = ~reg_controllable_hgrant9_out & ~n7380;
  assign n7382 = ~reg_controllable_hgrant9_out & ~n7381;
  assign n7383 = ~reg_controllable_nhgrant0_out & ~n7382;
  assign n7384 = ~n7305 & ~n7383;
  assign n7385 = reg_i_hready_out & ~n7384;
  assign n7386 = ~next_sys_fair<2>_out  & ~n1259;
  assign n7387 = ~next_sys_fair<2>_out  & ~n7386;
  assign n7388 = next_sys_fair<3>_out  & ~n7387;
  assign n7389 = next_sys_fair<0>_out  & ~n1259;
  assign n7390 = next_sys_fair<2>_out  & ~n1259;
  assign n7391 = ~next_sys_fair<2>_out  & ~n1228;
  assign n7392 = ~n7390 & ~n7391;
  assign n7393 = ~next_sys_fair<0>_out  & ~n7392;
  assign n7394 = ~n7389 & ~n7393;
  assign n7395 = ~next_sys_fair<3>_out  & ~n7394;
  assign n7396 = ~n7388 & ~n7395;
  assign n7397 = reg_controllable_hmaster1_out & ~n7396;
  assign n7398 = reg_controllable_hmaster2_out & ~n7396;
  assign n7399 = ~next_sys_fair<2>_out  & ~n1290;
  assign n7400 = ~next_sys_fair<2>_out  & ~n7399;
  assign n7401 = next_sys_fair<0>_out  & ~n7400;
  assign n7402 = ~next_sys_fair<2>_out  & ~n1323;
  assign n7403 = ~next_sys_fair<2>_out  & ~n7402;
  assign n7404 = ~next_sys_fair<0>_out  & ~n7403;
  assign n7405 = ~n7401 & ~n7404;
  assign n7406 = next_sys_fair<3>_out  & ~n7405;
  assign n7407 = next_sys_fair<0>_out  & ~n1323;
  assign n7408 = next_sys_fair<2>_out  & ~n1323;
  assign n7409 = ~next_sys_fair<2>_out  & ~n1477;
  assign n7410 = ~n7408 & ~n7409;
  assign n7411 = ~next_sys_fair<0>_out  & ~n7410;
  assign n7412 = ~n7407 & ~n7411;
  assign n7413 = ~next_sys_fair<3>_out  & ~n7412;
  assign n7414 = ~n7406 & ~n7413;
  assign n7415 = ~reg_controllable_hmaster2_out & ~n7414;
  assign n7416 = ~n7398 & ~n7415;
  assign n7417 = ~reg_controllable_hmaster1_out & ~n7416;
  assign n7418 = ~n7397 & ~n7417;
  assign n7419 = next_sys_fair<1>_out  & ~n7418;
  assign n7420 = ~next_sys_fair<2>_out  & ~n1367;
  assign n7421 = ~n7390 & ~n7420;
  assign n7422 = next_sys_fair<0>_out  & ~n7421;
  assign n7423 = ~next_sys_fair<2>_out  & ~n1389;
  assign n7424 = ~n7390 & ~n7423;
  assign n7425 = ~next_sys_fair<0>_out  & ~n7424;
  assign n7426 = ~n7422 & ~n7425;
  assign n7427 = ~next_sys_fair<3>_out  & ~n7426;
  assign n7428 = ~n7388 & ~n7427;
  assign n7429 = reg_controllable_hmaster1_out & ~n7428;
  assign n7430 = reg_controllable_hmaster2_out & ~n7428;
  assign n7431 = next_sys_fair<3>_out  & ~n7403;
  assign n7432 = ~next_sys_fair<2>_out  & ~n1421;
  assign n7433 = ~n7408 & ~n7432;
  assign n7434 = next_sys_fair<0>_out  & ~n7433;
  assign n7435 = ~n7399 & ~n7408;
  assign n7436 = ~next_sys_fair<0>_out  & ~n7435;
  assign n7437 = ~n7434 & ~n7436;
  assign n7438 = ~next_sys_fair<3>_out  & ~n7437;
  assign n7439 = ~n7431 & ~n7438;
  assign n7440 = ~reg_controllable_hmaster2_out & ~n7439;
  assign n7441 = ~n7430 & ~n7440;
  assign n7442 = ~reg_controllable_hmaster1_out & ~n7441;
  assign n7443 = ~n7429 & ~n7442;
  assign n7444 = ~next_sys_fair<1>_out  & ~n7443;
  assign n7445 = ~n7419 & ~n7444;
  assign n7446 = reg_controllable_hmaster0_out & ~n7445;
  assign n7447 = next_sys_fair<0>_out  & ~n7403;
  assign n7448 = ~next_sys_fair<0>_out  & ~n7400;
  assign n7449 = ~n7447 & ~n7448;
  assign n7450 = next_sys_fair<3>_out  & ~n7449;
  assign n7451 = ~n7413 & ~n7450;
  assign n7452 = ~reg_controllable_hmaster2_out & ~n7451;
  assign n7453 = ~n7398 & ~n7452;
  assign n7454 = ~reg_controllable_hmaster1_out & ~n7453;
  assign n7455 = ~n7397 & ~n7454;
  assign n7456 = next_sys_fair<1>_out  & ~n7455;
  assign n7457 = ~n7444 & ~n7456;
  assign n7458 = ~reg_controllable_hmaster0_out & ~n7457;
  assign n7459 = ~n7446 & ~n7458;
  assign n7460 = reg_controllable_hmaster3_out & ~n7459;
  assign n7461 = ~n7413 & ~n7431;
  assign n7462 = reg_controllable_hmaster1_out & ~n7461;
  assign n7463 = next_sys_fair<2>_out  & ~n1290;
  assign n7464 = ~n7402 & ~n7463;
  assign n7465 = next_sys_fair<0>_out  & ~n7464;
  assign n7466 = ~n7411 & ~n7465;
  assign n7467 = ~next_sys_fair<3>_out  & ~n7466;
  assign n7468 = ~n7431 & ~n7467;
  assign n7469 = reg_controllable_hmaster2_out & ~n7468;
  assign n7470 = next_sys_fair<0>_out  & ~n7435;
  assign n7471 = ~n7411 & ~n7470;
  assign n7472 = ~next_sys_fair<3>_out  & ~n7471;
  assign n7473 = ~n7431 & ~n7472;
  assign n7474 = ~reg_controllable_hmaster2_out & ~n7473;
  assign n7475 = ~n7469 & ~n7474;
  assign n7476 = ~reg_controllable_hmaster1_out & ~n7475;
  assign n7477 = ~n7462 & ~n7476;
  assign n7478 = next_sys_fair<1>_out  & ~n7477;
  assign n7479 = ~n7406 & ~n7438;
  assign n7480 = reg_controllable_hmaster2_out & ~n7479;
  assign n7481 = ~n7432 & ~n7463;
  assign n7482 = next_sys_fair<0>_out  & ~n7481;
  assign n7483 = ~n7436 & ~n7482;
  assign n7484 = ~next_sys_fair<3>_out  & ~n7483;
  assign n7485 = ~n7431 & ~n7484;
  assign n7486 = ~reg_controllable_hmaster2_out & ~n7485;
  assign n7487 = ~n7480 & ~n7486;
  assign n7488 = reg_controllable_hmaster1_out & ~n7487;
  assign n7489 = ~reg_controllable_hmaster1_out & ~n7439;
  assign n7490 = ~n7488 & ~n7489;
  assign n7491 = ~next_sys_fair<1>_out  & ~n7490;
  assign n7492 = ~n7478 & ~n7491;
  assign n7493 = reg_controllable_hmaster0_out & ~n7492;
  assign n7494 = ~n7409 & ~n7463;
  assign n7495 = ~next_sys_fair<0>_out  & ~n7494;
  assign n7496 = ~n7407 & ~n7495;
  assign n7497 = ~next_sys_fair<3>_out  & ~n7496;
  assign n7498 = ~n7431 & ~n7497;
  assign n7499 = reg_controllable_hmaster2_out & ~n7498;
  assign n7500 = ~next_sys_fair<2>_out  & ~n1325;
  assign n7501 = ~next_sys_fair<2>_out  & ~n7500;
  assign n7502 = next_sys_fair<3>_out  & ~n7501;
  assign n7503 = next_sys_fair<0>_out  & ~n1325;
  assign n7504 = next_sys_fair<2>_out  & ~n1325;
  assign n7505 = ~n4472 & ~n7504;
  assign n7506 = ~next_sys_fair<0>_out  & ~n7505;
  assign n7507 = ~n7503 & ~n7506;
  assign n7508 = ~next_sys_fair<3>_out  & ~n7507;
  assign n7509 = ~n7502 & ~n7508;
  assign n7510 = ~reg_controllable_hmaster2_out & ~n7509;
  assign n7511 = ~n7499 & ~n7510;
  assign n7512 = ~reg_controllable_hmaster1_out & ~n7511;
  assign n7513 = ~n7462 & ~n7512;
  assign n7514 = next_sys_fair<1>_out  & ~n7513;
  assign n7515 = ~n7438 & ~n7450;
  assign n7516 = reg_controllable_hmaster2_out & ~n7515;
  assign n7517 = ~next_sys_fair<0>_out  & ~n1290;
  assign n7518 = ~n7434 & ~n7517;
  assign n7519 = ~next_sys_fair<3>_out  & ~n7518;
  assign n7520 = ~n7431 & ~n7519;
  assign n7521 = ~reg_controllable_hmaster2_out & ~n7520;
  assign n7522 = ~n7516 & ~n7521;
  assign n7523 = reg_controllable_hmaster1_out & ~n7522;
  assign n7524 = reg_controllable_hmaster2_out & ~n7439;
  assign n7525 = ~n4551 & ~n7504;
  assign n7526 = next_sys_fair<0>_out  & ~n7525;
  assign n7527 = ~n4560 & ~n7504;
  assign n7528 = ~next_sys_fair<0>_out  & ~n7527;
  assign n7529 = ~n7526 & ~n7528;
  assign n7530 = ~next_sys_fair<3>_out  & ~n7529;
  assign n7531 = ~n7502 & ~n7530;
  assign n7532 = ~reg_controllable_hmaster2_out & ~n7531;
  assign n7533 = ~n7524 & ~n7532;
  assign n7534 = ~reg_controllable_hmaster1_out & ~n7533;
  assign n7535 = ~n7523 & ~n7534;
  assign n7536 = ~next_sys_fair<1>_out  & ~n7535;
  assign n7537 = ~n7514 & ~n7536;
  assign n7538 = ~reg_controllable_hmaster0_out & ~n7537;
  assign n7539 = ~n7493 & ~n7538;
  assign n7540 = ~reg_controllable_hmaster3_out & ~n7539;
  assign n7541 = ~n7460 & ~n7540;
  assign n7542 = ~reg_i_hready_out & ~n7541;
  assign n7543 = ~n7385 & ~n7542;
  assign n7544 = ~reg_i_hlock0_out & ~n7543;
  assign n7545 = ~n6568 & ~n7544;
  assign n7546 = ~reg_i_hbusreq1_out & ~n7545;
  assign n7547 = ~n5469 & ~n7546;
  assign n7548 = ~reg_i_hbusreq2_out & ~n7547;
  assign n7549 = ~n5468 & ~n7548;
  assign n7550 = ~reg_i_hbusreq4_out & ~n7549;
  assign n7551 = ~n5467 & ~n7550;
  assign n7552 = ~reg_i_hbusreq3_out & ~n7551;
  assign n7553 = ~n5466 & ~n7552;
  assign n7554 = ~reg_i_hbusreq8_out & ~n7553;
  assign n7555 = ~n5465 & ~n7554;
  assign n7556 = ~reg_i_hbusreq7_out & ~n7555;
  assign n7557 = ~n5464 & ~n7556;
  assign n7558 = ~reg_i_hbusreq6_out & ~n7557;
  assign n7559 = ~n5463 & ~n7558;
  assign n7560 = ~reg_i_hbusreq5_out & ~n7559;
  assign n7561 = ~n5462 & ~n7560;
  assign n7562 = ~reg_i_hbusreq0_out & ~n7561;
  assign n7563 = ~n5461 & ~n7562;
  assign n7564 = ~reg_i_hbusreq9_out & ~n7563;
  assign n7565 = ~n5460 & ~n7564;
  assign n7566 = ~reg_controllable_ndecide_out & ~n7565;
  assign n7567 = ~n2867 & ~n7566;
  assign n7568 = ~env_safe_err_happened_out & n7567;
  assign n7569 = ~env_safe_err_happened_out & ~n7568;
  assign n7570 = n87 & ~n7569;
  assign n7571 = n87 & ~n7570;
  assign n7572 = i_hlock0 & ~i_hbusreq0;
  assign n7573 = i_hlock1 & ~i_hbusreq1;
  assign n7574 = ~n7572 & ~n7573;
  assign n7575 = i_hlock2 & ~i_hbusreq2;
  assign n7576 = n7574 & ~n7575;
  assign n7577 = i_hlock3 & ~i_hbusreq3;
  assign n7578 = n7576 & ~n7577;
  assign n7579 = i_hlock4 & ~i_hbusreq4;
  assign n7580 = n7578 & ~n7579;
  assign n7581 = i_hlock5 & ~i_hbusreq5;
  assign n7582 = n7580 & ~n7581;
  assign n7583 = i_hlock6 & ~i_hbusreq6;
  assign n7584 = n7582 & ~n7583;
  assign n7585 = i_hlock7 & ~i_hbusreq7;
  assign n7586 = n7584 & ~n7585;
  assign n7587 = i_hlock8 & ~i_hbusreq8;
  assign n7588 = n7586 & ~n7587;
  assign n7589 = i_hlock9 & ~i_hbusreq9;
  assign n7590 = n7588 & ~n7589;
  assign n7591 = n87 & env_safe_err_happened_out;
  assign n7592 = n7590 & ~n7591;
  assign n7593 = n87 & next_sys_fair<4>_out ;
  assign n7594 = n87 & next_sys_fair<3>_out ;
  assign n7595 = n87 & next_sys_fair<2>_out ;
  assign n7596 = n87 & next_sys_fair<0>_out ;
  assign n7597 = n87 & next_sys_fair<1>_out ;
  assign n7598 = n7596 & n7597;
  assign n7599 = ~n7595 & n7598;
  assign n7600 = n7594 & n7599;
  assign n7601 = ~n7593 & n7600;
  assign n7602 = ~controllable_hmaster1 & controllable_hmaster0;
  assign n7603 = ~controllable_hmaster2 & n7602;
  assign n7604 = controllable_hmaster3 & n7603;
  assign n7605 = i_hbusreq9 & ~n7604;
  assign n7606 = n7601 & ~n7605;
  assign n7607 = ~n7596 & n7597;
  assign n7608 = n7595 & n7607;
  assign n7609 = ~n7594 & n7608;
  assign n7610 = ~n7593 & n7609;
  assign n7611 = ~controllable_hmaster1 & ~controllable_hmaster0;
  assign n7612 = controllable_hmaster2 & n7611;
  assign n7613 = ~controllable_hmaster3 & n7612;
  assign n7614 = i_hbusreq4 & ~n7613;
  assign n7615 = n7610 & ~n7614;
  assign n7616 = ~n7595 & n7607;
  assign n7617 = n7594 & n7616;
  assign n7618 = ~n7593 & n7617;
  assign n7619 = ~controllable_hmaster2 & n7611;
  assign n7620 = controllable_hmaster3 & n7619;
  assign n7621 = i_hbusreq8 & ~n7620;
  assign n7622 = n7618 & ~n7621;
  assign n7623 = n7595 & n7598;
  assign n7624 = ~n7594 & n7623;
  assign n7625 = ~n7593 & n7624;
  assign n7626 = controllable_hmaster2 & n7602;
  assign n7627 = ~controllable_hmaster3 & n7626;
  assign n7628 = i_hbusreq5 & ~n7627;
  assign n7629 = n7625 & ~n7628;
  assign n7630 = ~n7622 & ~n7629;
  assign n7631 = ~n7615 & n7630;
  assign n7632 = n7596 & ~n7597;
  assign n7633 = n7595 & n7632;
  assign n7634 = ~n7594 & n7633;
  assign n7635 = ~n7593 & n7634;
  assign n7636 = controllable_hmaster1 & controllable_hmaster0;
  assign n7637 = ~controllable_hmaster2 & n7636;
  assign n7638 = ~controllable_hmaster3 & n7637;
  assign n7639 = i_hbusreq3 & ~n7638;
  assign n7640 = n7635 & ~n7639;
  assign n7641 = n87 & reg_stateG2_out;
  assign n7642 = ~n7596 & ~n7597;
  assign n7643 = ~n7595 & n7642;
  assign n7644 = ~n7594 & n7643;
  assign n7645 = ~n7593 & n7644;
  assign n7646 = ~n7641 & n7645;
  assign n7647 = n87 & reg_stateG3_0_out;
  assign n7648 = n87 & reg_stateG3_1_out;
  assign n7649 = ~n7647 & ~n7648;
  assign n7650 = n87 & reg_stateG3_2_out;
  assign n7651 = n7649 & ~n7650;
  assign n7652 = ~n7595 & n7632;
  assign n7653 = ~n7594 & n7652;
  assign n7654 = ~n7593 & n7653;
  assign n7655 = n7651 & n7654;
  assign n7656 = ~n7646 & ~n7655;
  assign n7657 = ~n7594 & n7616;
  assign n7658 = ~n7593 & n7657;
  assign n7659 = ~controllable_hmaster3 & n7619;
  assign n7660 = i_hbusreq0 & ~n7659;
  assign n7661 = n7658 & ~n7660;
  assign n7662 = n7595 & n7642;
  assign n7663 = ~n7594 & n7662;
  assign n7664 = ~n7593 & n7663;
  assign n7665 = controllable_hmaster1 & ~controllable_hmaster0;
  assign n7666 = ~controllable_hmaster2 & n7665;
  assign n7667 = ~controllable_hmaster3 & n7666;
  assign n7668 = i_hbusreq2 & ~n7667;
  assign n7669 = n7664 & ~n7668;
  assign n7670 = ~n7594 & n7599;
  assign n7671 = ~n7593 & n7670;
  assign n7672 = ~controllable_hmaster3 & n7603;
  assign n7673 = i_hbusreq1 & ~n7672;
  assign n7674 = n7671 & ~n7673;
  assign n7675 = ~n7669 & ~n7674;
  assign n7676 = ~n7661 & n7675;
  assign n7677 = n7656 & n7676;
  assign n7678 = n7594 & n7652;
  assign n7679 = ~n7593 & n7678;
  assign n7680 = controllable_hmaster2 & n7636;
  assign n7681 = ~controllable_hmaster3 & n7680;
  assign n7682 = i_hbusreq7 & ~n7681;
  assign n7683 = n7679 & ~n7682;
  assign n7684 = n7594 & n7643;
  assign n7685 = ~n7593 & n7684;
  assign n7686 = controllable_hmaster2 & n7665;
  assign n7687 = ~controllable_hmaster3 & n7686;
  assign n7688 = i_hbusreq6 & ~n7687;
  assign n7689 = n7685 & ~n7688;
  assign n7690 = ~n7683 & ~n7689;
  assign n7691 = n7677 & n7690;
  assign n7692 = ~n7640 & n7691;
  assign n7693 = n7631 & n7692;
  assign n7694 = ~n7606 & n7693;
  assign n7695 = n87 & fair_cnt<0>_out ;
  assign n7696 = n87 & next_env_fair_out;
  assign n7697 = i_hready & n7696;
  assign n7698 = n7695 & n7697;
  assign n7699 = n87 & fair_cnt<1>_out ;
  assign n7700 = n7698 & n7699;
  assign n7701 = n87 & fair_cnt<2>_out ;
  assign n7702 = ~n7700 & ~n7701;
  assign n7703 = n7700 & n7701;
  assign n7704 = ~n7702 & ~n7703;
  assign n7705 = n7694 & n7704;
  assign n7706 = ~n7640 & n7690;
  assign n7707 = ~n7661 & n7706;
  assign n7708 = n7656 & n7707;
  assign n7709 = ~n7698 & ~n7699;
  assign n7710 = ~n7700 & ~n7709;
  assign n7711 = ~n7606 & n7710;
  assign n7712 = n7675 & n7711;
  assign n7713 = n7631 & n7712;
  assign n7714 = n7708 & n7713;
  assign n7715 = ~n7615 & ~n7640;
  assign n7716 = ~n7695 & ~n7697;
  assign n7717 = ~n7698 & ~n7716;
  assign n7718 = ~n7606 & n7717;
  assign n7719 = ~n7622 & n7718;
  assign n7720 = ~n7629 & n7690;
  assign n7721 = n7719 & n7720;
  assign n7722 = n7715 & n7721;
  assign n7723 = n7677 & n7722;
  assign n7724 = n87 & reg_stateA1_out;
  assign n7725 = ~n7696 & n7724;
  assign n7726 = ~n7697 & ~n7725;
  assign n7727 = ~n7606 & n7726;
  assign n7728 = n7693 & n7727;
  assign n7729 = controllable_busreq & n7724;
  assign n7730 = ~i_hburst1 & ~i_hburst0;
  assign n7731 = controllable_hmastlock & n7730;
  assign n7732 = ~n7724 & n7731;
  assign n7733 = ~n7729 & ~n7732;
  assign n7734 = i_hready & ~controllable_ndecide;
  assign n7735 = ~controllable_ndecide & ~n7734;
  assign n7736 = ~n7733 & ~n7735;
  assign n7737 = ~n7733 & ~n7736;
  assign n7738 = controllable_hmaster1 & ~n7737;
  assign n7739 = controllable_hmaster2 & ~n7737;
  assign n7740 = controllable_hmaster2 & ~n7739;
  assign n7741 = ~controllable_hmaster1 & ~n7740;
  assign n7742 = ~n7738 & ~n7741;
  assign n7743 = controllable_hmaster3 & ~n7742;
  assign n7744 = controllable_hmaster3 & ~n7743;
  assign n7745 = i_hbusreq7 & ~n7744;
  assign n7746 = i_hbusreq8 & ~n7742;
  assign n7747 = i_hbusreq6 & ~n7742;
  assign n7748 = i_hbusreq5 & ~n7737;
  assign n7749 = i_hbusreq4 & ~n7737;
  assign n7750 = i_hbusreq9 & ~n7737;
  assign n7751 = i_hbusreq3 & ~n7737;
  assign n7752 = i_hbusreq1 & ~n7737;
  assign n7753 = i_hbusreq2 & ~n7735;
  assign n7754 = i_hbusreq0 & ~n7735;
  assign n7755 = i_hbusreq0 & ~n7754;
  assign n7756 = ~i_hbusreq2 & ~n7755;
  assign n7757 = ~n7753 & ~n7756;
  assign n7758 = ~n7733 & ~n7757;
  assign n7759 = ~n7733 & ~n7758;
  assign n7760 = ~i_hbusreq1 & ~n7759;
  assign n7761 = ~n7752 & ~n7760;
  assign n7762 = ~i_hbusreq3 & ~n7761;
  assign n7763 = ~n7751 & ~n7762;
  assign n7764 = ~i_hbusreq9 & ~n7763;
  assign n7765 = ~n7750 & ~n7764;
  assign n7766 = ~i_hbusreq4 & ~n7765;
  assign n7767 = ~n7749 & ~n7766;
  assign n7768 = ~i_hbusreq5 & ~n7767;
  assign n7769 = ~n7748 & ~n7768;
  assign n7770 = controllable_hmaster1 & ~n7769;
  assign n7771 = controllable_hmaster2 & ~n7769;
  assign n7772 = controllable_hmaster2 & ~n7771;
  assign n7773 = ~controllable_hmaster1 & ~n7772;
  assign n7774 = ~n7770 & ~n7773;
  assign n7775 = ~i_hbusreq6 & ~n7774;
  assign n7776 = ~n7747 & ~n7775;
  assign n7777 = ~i_hbusreq8 & ~n7776;
  assign n7778 = ~n7746 & ~n7777;
  assign n7779 = controllable_hmaster3 & ~n7778;
  assign n7780 = controllable_hmaster3 & ~n7779;
  assign n7781 = ~i_hbusreq7 & ~n7780;
  assign n7782 = ~n7745 & ~n7781;
  assign n7783 = ~n7728 & ~n7782;
  assign n7784 = ~n7728 & ~n7783;
  assign n7785 = ~n7723 & ~n7784;
  assign n7786 = ~n7723 & ~n7785;
  assign n7787 = ~n7714 & ~n7786;
  assign n7788 = ~n7714 & ~n7787;
  assign n7789 = n7705 & ~n7788;
  assign n7790 = ~n7705 & ~n7782;
  assign n7791 = ~n7789 & ~n7790;
  assign n7792 = controllable_hgrant9 & ~n7791;
  assign n7793 = controllable_hgrant7 & ~n7791;
  assign n7794 = controllable_hgrant8 & ~n7791;
  assign n7795 = controllable_hmastlock & n7651;
  assign n7796 = ~controllable_nstart & n7795;
  assign n7797 = ~i_hburst0 & n7796;
  assign n7798 = i_hburst1 & n7797;
  assign n7799 = i_hready & n7798;
  assign n7800 = n7647 & n7648;
  assign n7801 = ~n7650 & n7800;
  assign n7802 = i_hready & n7801;
  assign n7803 = n7648 & ~n7802;
  assign n7804 = i_hready & ~n7650;
  assign n7805 = n7647 & ~n7648;
  assign n7806 = n7804 & n7805;
  assign n7807 = ~n7803 & ~n7806;
  assign n7808 = ~n7799 & n7807;
  assign n7809 = controllable_hgrant6 & ~n7742;
  assign n7810 = controllable_hgrant5 & ~n7737;
  assign n7811 = controllable_hgrant4 & ~n7737;
  assign n7812 = controllable_hgrant3 & ~n7737;
  assign n7813 = controllable_hgrant1 & ~n7737;
  assign n7814 = controllable_hgrant2 & ~n7735;
  assign n7815 = ~controllable_hmastlock & n7735;
  assign n7816 = ~controllable_hmastlock & ~n7815;
  assign n7817 = controllable_locked & ~n7816;
  assign n7818 = controllable_hmastlock & ~n7735;
  assign n7819 = ~controllable_locked & ~n7818;
  assign n7820 = ~n7817 & ~n7819;
  assign n7821 = ~controllable_hgrant2 & n7820;
  assign n7822 = ~n7814 & ~n7821;
  assign n7823 = ~n7733 & ~n7822;
  assign n7824 = ~n7733 & ~n7823;
  assign n7825 = ~controllable_hgrant1 & ~n7824;
  assign n7826 = ~n7813 & ~n7825;
  assign n7827 = ~controllable_hgrant3 & ~n7826;
  assign n7828 = ~n7812 & ~n7827;
  assign n7829 = ~controllable_hgrant4 & ~n7828;
  assign n7830 = ~n7811 & ~n7829;
  assign n7831 = ~controllable_hgrant5 & ~n7830;
  assign n7832 = ~n7810 & ~n7831;
  assign n7833 = controllable_hmaster1 & ~n7832;
  assign n7834 = controllable_hmaster2 & ~n7832;
  assign n7835 = controllable_hmaster2 & ~n7834;
  assign n7836 = ~controllable_hmaster1 & ~n7835;
  assign n7837 = ~n7833 & ~n7836;
  assign n7838 = ~controllable_hgrant6 & ~n7837;
  assign n7839 = ~n7809 & ~n7838;
  assign n7840 = controllable_hmaster3 & ~n7839;
  assign n7841 = controllable_hmaster3 & ~n7840;
  assign n7842 = i_hbusreq7 & ~n7841;
  assign n7843 = i_hbusreq8 & ~n7839;
  assign n7844 = controllable_hgrant6 & ~n7776;
  assign n7845 = i_hbusreq6 & ~n7837;
  assign n7846 = controllable_hgrant5 & ~n7769;
  assign n7847 = i_hbusreq5 & ~n7830;
  assign n7848 = controllable_hgrant4 & ~n7767;
  assign n7849 = i_hbusreq4 & ~n7828;
  assign n7850 = i_hbusreq9 & ~n7828;
  assign n7851 = controllable_hgrant3 & ~n7763;
  assign n7852 = i_hbusreq3 & ~n7826;
  assign n7853 = controllable_hgrant1 & ~n7761;
  assign n7854 = i_hbusreq1 & ~n7824;
  assign n7855 = controllable_hgrant2 & ~n7757;
  assign n7856 = i_hbusreq2 & ~n7820;
  assign n7857 = i_hbusreq0 & ~n7820;
  assign n7858 = controllable_ndecide & controllable_hmastlock;
  assign n7859 = controllable_locked & n7858;
  assign n7860 = ~controllable_ndecide & ~controllable_hmastlock;
  assign n7861 = ~controllable_hmastlock & ~n7860;
  assign n7862 = ~controllable_locked & n7861;
  assign n7863 = ~n7859 & ~n7862;
  assign n7864 = ~i_hbusreq0 & ~n7863;
  assign n7865 = ~n7857 & ~n7864;
  assign n7866 = ~i_hbusreq2 & ~n7865;
  assign n7867 = ~n7856 & ~n7866;
  assign n7868 = ~controllable_hgrant2 & n7867;
  assign n7869 = ~n7855 & ~n7868;
  assign n7870 = ~n7733 & ~n7869;
  assign n7871 = ~n7733 & ~n7870;
  assign n7872 = ~i_hbusreq1 & ~n7871;
  assign n7873 = ~n7854 & ~n7872;
  assign n7874 = ~controllable_hgrant1 & ~n7873;
  assign n7875 = ~n7853 & ~n7874;
  assign n7876 = ~i_hbusreq3 & ~n7875;
  assign n7877 = ~n7852 & ~n7876;
  assign n7878 = ~controllable_hgrant3 & ~n7877;
  assign n7879 = ~n7851 & ~n7878;
  assign n7880 = ~i_hbusreq9 & ~n7879;
  assign n7881 = ~n7850 & ~n7880;
  assign n7882 = ~i_hbusreq4 & ~n7881;
  assign n7883 = ~n7849 & ~n7882;
  assign n7884 = ~controllable_hgrant4 & ~n7883;
  assign n7885 = ~n7848 & ~n7884;
  assign n7886 = ~i_hbusreq5 & ~n7885;
  assign n7887 = ~n7847 & ~n7886;
  assign n7888 = ~controllable_hgrant5 & ~n7887;
  assign n7889 = ~n7846 & ~n7888;
  assign n7890 = controllable_hmaster1 & ~n7889;
  assign n7891 = controllable_hmaster2 & ~n7889;
  assign n7892 = controllable_hmaster2 & ~n7891;
  assign n7893 = ~controllable_hmaster1 & ~n7892;
  assign n7894 = ~n7890 & ~n7893;
  assign n7895 = ~i_hbusreq6 & ~n7894;
  assign n7896 = ~n7845 & ~n7895;
  assign n7897 = ~controllable_hgrant6 & ~n7896;
  assign n7898 = ~n7844 & ~n7897;
  assign n7899 = ~i_hbusreq8 & ~n7898;
  assign n7900 = ~n7843 & ~n7899;
  assign n7901 = controllable_hmaster3 & ~n7900;
  assign n7902 = controllable_hmaster3 & ~n7901;
  assign n7903 = ~i_hbusreq7 & ~n7902;
  assign n7904 = ~n7842 & ~n7903;
  assign n7905 = ~n7728 & ~n7904;
  assign n7906 = ~n7728 & ~n7905;
  assign n7907 = ~n7723 & ~n7906;
  assign n7908 = ~n7723 & ~n7907;
  assign n7909 = ~n7714 & ~n7908;
  assign n7910 = ~n7714 & ~n7909;
  assign n7911 = n7705 & ~n7910;
  assign n7912 = ~n7705 & ~n7904;
  assign n7913 = ~n7911 & ~n7912;
  assign n7914 = ~n7808 & ~n7913;
  assign n7915 = ~i_hready & n7798;
  assign n7916 = ~n7647 & ~n7804;
  assign n7917 = n7647 & n7804;
  assign n7918 = ~n7916 & ~n7917;
  assign n7919 = ~n7649 & n7918;
  assign n7920 = ~n7915 & ~n7919;
  assign n7921 = ~n7904 & ~n7920;
  assign n7922 = i_hready & n7649;
  assign n7923 = n7650 & ~n7922;
  assign n7924 = ~n7802 & ~n7923;
  assign n7925 = controllable_busreq & n7641;
  assign n7926 = ~controllable_nstart & ~n7641;
  assign n7927 = n7731 & n7926;
  assign n7928 = ~n7925 & ~n7927;
  assign n7929 = ~n7824 & ~n7928;
  assign n7930 = ~i_hready & ~controllable_hmastlock;
  assign n7931 = ~controllable_hmastlock & ~n7930;
  assign n7932 = controllable_locked & ~n7931;
  assign n7933 = i_hready & controllable_hmastlock;
  assign n7934 = ~controllable_locked & ~n7933;
  assign n7935 = ~n7932 & ~n7934;
  assign n7936 = ~controllable_hgrant2 & n7935;
  assign n7937 = ~n7814 & ~n7936;
  assign n7938 = ~n7733 & ~n7937;
  assign n7939 = ~n7733 & ~n7938;
  assign n7940 = n7928 & ~n7939;
  assign n7941 = ~n7929 & ~n7940;
  assign n7942 = ~controllable_hgrant1 & ~n7941;
  assign n7943 = ~n7813 & ~n7942;
  assign n7944 = ~controllable_hgrant3 & ~n7943;
  assign n7945 = ~n7812 & ~n7944;
  assign n7946 = ~controllable_hgrant4 & ~n7945;
  assign n7947 = ~n7811 & ~n7946;
  assign n7948 = ~controllable_hgrant5 & ~n7947;
  assign n7949 = ~n7810 & ~n7948;
  assign n7950 = controllable_hmaster1 & ~n7949;
  assign n7951 = controllable_hmaster2 & ~n7949;
  assign n7952 = controllable_hmaster2 & ~n7951;
  assign n7953 = ~controllable_hmaster1 & ~n7952;
  assign n7954 = ~n7950 & ~n7953;
  assign n7955 = ~controllable_hgrant6 & ~n7954;
  assign n7956 = ~n7809 & ~n7955;
  assign n7957 = controllable_hmaster3 & ~n7956;
  assign n7958 = controllable_hmaster3 & ~n7957;
  assign n7959 = i_hbusreq7 & ~n7958;
  assign n7960 = i_hbusreq8 & ~n7956;
  assign n7961 = i_hbusreq6 & ~n7954;
  assign n7962 = i_hbusreq5 & ~n7947;
  assign n7963 = i_hbusreq4 & ~n7945;
  assign n7964 = i_hbusreq9 & ~n7945;
  assign n7965 = i_hbusreq3 & ~n7943;
  assign n7966 = i_hbusreq1 & ~n7941;
  assign n7967 = ~n7871 & ~n7928;
  assign n7968 = i_hbusreq2 & ~n7935;
  assign n7969 = i_hbusreq0 & ~n7935;
  assign n7970 = i_hready & controllable_ndecide;
  assign n7971 = controllable_ndecide & ~n7970;
  assign n7972 = ~controllable_hmastlock & n7971;
  assign n7973 = ~n7858 & ~n7972;
  assign n7974 = controllable_locked & ~n7973;
  assign n7975 = controllable_hmastlock & ~n7971;
  assign n7976 = ~n7860 & ~n7975;
  assign n7977 = ~controllable_locked & n7976;
  assign n7978 = ~n7974 & ~n7977;
  assign n7979 = ~i_hbusreq0 & ~n7978;
  assign n7980 = ~n7969 & ~n7979;
  assign n7981 = ~i_hbusreq2 & ~n7980;
  assign n7982 = ~n7968 & ~n7981;
  assign n7983 = ~controllable_hgrant2 & n7982;
  assign n7984 = ~n7855 & ~n7983;
  assign n7985 = ~n7733 & ~n7984;
  assign n7986 = ~n7733 & ~n7985;
  assign n7987 = n7928 & ~n7986;
  assign n7988 = ~n7967 & ~n7987;
  assign n7989 = ~i_hbusreq1 & ~n7988;
  assign n7990 = ~n7966 & ~n7989;
  assign n7991 = ~controllable_hgrant1 & ~n7990;
  assign n7992 = ~n7853 & ~n7991;
  assign n7993 = ~i_hbusreq3 & ~n7992;
  assign n7994 = ~n7965 & ~n7993;
  assign n7995 = ~controllable_hgrant3 & ~n7994;
  assign n7996 = ~n7851 & ~n7995;
  assign n7997 = ~i_hbusreq9 & ~n7996;
  assign n7998 = ~n7964 & ~n7997;
  assign n7999 = ~i_hbusreq4 & ~n7998;
  assign n8000 = ~n7963 & ~n7999;
  assign n8001 = ~controllable_hgrant4 & ~n8000;
  assign n8002 = ~n7848 & ~n8001;
  assign n8003 = ~i_hbusreq5 & ~n8002;
  assign n8004 = ~n7962 & ~n8003;
  assign n8005 = ~controllable_hgrant5 & ~n8004;
  assign n8006 = ~n7846 & ~n8005;
  assign n8007 = controllable_hmaster1 & ~n8006;
  assign n8008 = controllable_hmaster2 & ~n8006;
  assign n8009 = controllable_hmaster2 & ~n8008;
  assign n8010 = ~controllable_hmaster1 & ~n8009;
  assign n8011 = ~n8007 & ~n8010;
  assign n8012 = ~i_hbusreq6 & ~n8011;
  assign n8013 = ~n7961 & ~n8012;
  assign n8014 = ~controllable_hgrant6 & ~n8013;
  assign n8015 = ~n7844 & ~n8014;
  assign n8016 = ~i_hbusreq8 & ~n8015;
  assign n8017 = ~n7960 & ~n8016;
  assign n8018 = controllable_hmaster3 & ~n8017;
  assign n8019 = controllable_hmaster3 & ~n8018;
  assign n8020 = ~i_hbusreq7 & ~n8019;
  assign n8021 = ~n7959 & ~n8020;
  assign n8022 = ~n7924 & ~n8021;
  assign n8023 = ~n7733 & n7814;
  assign n8024 = ~n7733 & ~n8023;
  assign n8025 = n7928 & ~n8024;
  assign n8026 = ~n7929 & ~n8025;
  assign n8027 = ~controllable_hgrant1 & ~n8026;
  assign n8028 = ~n7813 & ~n8027;
  assign n8029 = ~controllable_hgrant3 & ~n8028;
  assign n8030 = ~n7812 & ~n8029;
  assign n8031 = ~controllable_hgrant4 & ~n8030;
  assign n8032 = ~n7811 & ~n8031;
  assign n8033 = ~controllable_hgrant5 & ~n8032;
  assign n8034 = ~n7810 & ~n8033;
  assign n8035 = controllable_hmaster1 & ~n8034;
  assign n8036 = controllable_hmaster2 & ~n8034;
  assign n8037 = ~i_hready & ~controllable_hgrant2;
  assign n8038 = ~controllable_hgrant2 & ~n8037;
  assign n8039 = ~n7733 & ~n8038;
  assign n8040 = ~n7733 & ~n8039;
  assign n8041 = n7928 & ~n8040;
  assign n8042 = n7928 & ~n8041;
  assign n8043 = ~controllable_hgrant1 & ~n8042;
  assign n8044 = ~controllable_hgrant1 & ~n8043;
  assign n8045 = ~controllable_hgrant3 & ~n8044;
  assign n8046 = ~controllable_hgrant3 & ~n8045;
  assign n8047 = ~controllable_hgrant4 & ~n8046;
  assign n8048 = ~controllable_hgrant4 & ~n8047;
  assign n8049 = ~controllable_hgrant5 & ~n8048;
  assign n8050 = ~controllable_hgrant5 & ~n8049;
  assign n8051 = ~controllable_hmaster2 & ~n8050;
  assign n8052 = ~n8036 & ~n8051;
  assign n8053 = ~controllable_hmaster1 & ~n8052;
  assign n8054 = ~n8035 & ~n8053;
  assign n8055 = ~controllable_hgrant6 & ~n8054;
  assign n8056 = ~n7809 & ~n8055;
  assign n8057 = controllable_hmaster3 & ~n8056;
  assign n8058 = ~controllable_hgrant6 & ~n8050;
  assign n8059 = ~controllable_hgrant6 & ~n8058;
  assign n8060 = ~controllable_hmaster3 & ~n8059;
  assign n8061 = ~n8057 & ~n8060;
  assign n8062 = i_hbusreq7 & ~n8061;
  assign n8063 = i_hbusreq8 & ~n8056;
  assign n8064 = i_hbusreq6 & ~n8054;
  assign n8065 = i_hbusreq5 & ~n8032;
  assign n8066 = i_hbusreq4 & ~n8030;
  assign n8067 = i_hbusreq9 & ~n8030;
  assign n8068 = i_hbusreq3 & ~n8028;
  assign n8069 = i_hbusreq1 & ~n8026;
  assign n8070 = ~i_hbusreq0 & controllable_ndecide;
  assign n8071 = ~i_hbusreq0 & ~n8070;
  assign n8072 = ~i_hbusreq2 & ~n8071;
  assign n8073 = ~i_hbusreq2 & ~n8072;
  assign n8074 = ~controllable_hgrant2 & n8073;
  assign n8075 = ~n7855 & ~n8074;
  assign n8076 = ~n7733 & ~n8075;
  assign n8077 = ~n7733 & ~n8076;
  assign n8078 = n7928 & ~n8077;
  assign n8079 = ~n7967 & ~n8078;
  assign n8080 = ~i_hbusreq1 & ~n8079;
  assign n8081 = ~n8069 & ~n8080;
  assign n8082 = ~controllable_hgrant1 & ~n8081;
  assign n8083 = ~n7853 & ~n8082;
  assign n8084 = ~i_hbusreq3 & ~n8083;
  assign n8085 = ~n8068 & ~n8084;
  assign n8086 = ~controllable_hgrant3 & ~n8085;
  assign n8087 = ~n7851 & ~n8086;
  assign n8088 = ~i_hbusreq9 & ~n8087;
  assign n8089 = ~n8067 & ~n8088;
  assign n8090 = ~i_hbusreq4 & ~n8089;
  assign n8091 = ~n8066 & ~n8090;
  assign n8092 = ~controllable_hgrant4 & ~n8091;
  assign n8093 = ~n7848 & ~n8092;
  assign n8094 = ~i_hbusreq5 & ~n8093;
  assign n8095 = ~n8065 & ~n8094;
  assign n8096 = ~controllable_hgrant5 & ~n8095;
  assign n8097 = ~n7846 & ~n8096;
  assign n8098 = controllable_hmaster1 & ~n8097;
  assign n8099 = controllable_hmaster2 & ~n8097;
  assign n8100 = i_hbusreq5 & ~n8048;
  assign n8101 = i_hbusreq4 & ~n8046;
  assign n8102 = i_hbusreq9 & ~n8046;
  assign n8103 = i_hbusreq3 & ~n8044;
  assign n8104 = i_hbusreq1 & ~n8042;
  assign n8105 = i_hready & i_hbusreq2;
  assign n8106 = i_hready & i_hbusreq0;
  assign n8107 = ~i_hbusreq0 & n7970;
  assign n8108 = ~n8106 & ~n8107;
  assign n8109 = ~i_hbusreq2 & ~n8108;
  assign n8110 = ~n8105 & ~n8109;
  assign n8111 = ~controllable_hgrant2 & n8110;
  assign n8112 = ~controllable_hgrant2 & ~n8111;
  assign n8113 = ~n7733 & ~n8112;
  assign n8114 = ~n7733 & ~n8113;
  assign n8115 = n7928 & ~n8114;
  assign n8116 = n7928 & ~n8115;
  assign n8117 = ~i_hbusreq1 & ~n8116;
  assign n8118 = ~n8104 & ~n8117;
  assign n8119 = ~controllable_hgrant1 & ~n8118;
  assign n8120 = ~controllable_hgrant1 & ~n8119;
  assign n8121 = ~i_hbusreq3 & ~n8120;
  assign n8122 = ~n8103 & ~n8121;
  assign n8123 = ~controllable_hgrant3 & ~n8122;
  assign n8124 = ~controllable_hgrant3 & ~n8123;
  assign n8125 = ~i_hbusreq9 & ~n8124;
  assign n8126 = ~n8102 & ~n8125;
  assign n8127 = ~i_hbusreq4 & ~n8126;
  assign n8128 = ~n8101 & ~n8127;
  assign n8129 = ~controllable_hgrant4 & ~n8128;
  assign n8130 = ~controllable_hgrant4 & ~n8129;
  assign n8131 = ~i_hbusreq5 & ~n8130;
  assign n8132 = ~n8100 & ~n8131;
  assign n8133 = ~controllable_hgrant5 & ~n8132;
  assign n8134 = ~controllable_hgrant5 & ~n8133;
  assign n8135 = ~controllable_hmaster2 & ~n8134;
  assign n8136 = ~n8099 & ~n8135;
  assign n8137 = ~controllable_hmaster1 & ~n8136;
  assign n8138 = ~n8098 & ~n8137;
  assign n8139 = ~i_hbusreq6 & ~n8138;
  assign n8140 = ~n8064 & ~n8139;
  assign n8141 = ~controllable_hgrant6 & ~n8140;
  assign n8142 = ~n7844 & ~n8141;
  assign n8143 = ~i_hbusreq8 & ~n8142;
  assign n8144 = ~n8063 & ~n8143;
  assign n8145 = controllable_hmaster3 & ~n8144;
  assign n8146 = i_hbusreq8 & ~n8059;
  assign n8147 = i_hbusreq6 & ~n8050;
  assign n8148 = ~i_hbusreq6 & ~n8134;
  assign n8149 = ~n8147 & ~n8148;
  assign n8150 = ~controllable_hgrant6 & ~n8149;
  assign n8151 = ~controllable_hgrant6 & ~n8150;
  assign n8152 = ~i_hbusreq8 & ~n8151;
  assign n8153 = ~n8146 & ~n8152;
  assign n8154 = ~controllable_hmaster3 & ~n8153;
  assign n8155 = ~n8145 & ~n8154;
  assign n8156 = ~i_hbusreq7 & ~n8155;
  assign n8157 = ~n8062 & ~n8156;
  assign n8158 = n7924 & ~n8157;
  assign n8159 = ~n8022 & ~n8158;
  assign n8160 = n7920 & ~n8159;
  assign n8161 = ~n7921 & ~n8160;
  assign n8162 = ~n7728 & ~n8161;
  assign n8163 = ~n7728 & ~n8162;
  assign n8164 = ~n7723 & ~n8163;
  assign n8165 = ~n7723 & ~n8164;
  assign n8166 = ~n7714 & ~n8165;
  assign n8167 = ~n7714 & ~n8166;
  assign n8168 = n7705 & ~n8167;
  assign n8169 = ~n7705 & ~n8161;
  assign n8170 = ~n8168 & ~n8169;
  assign n8171 = n7808 & ~n8170;
  assign n8172 = ~n7914 & ~n8171;
  assign n8173 = ~controllable_hgrant8 & ~n8172;
  assign n8174 = ~n7794 & ~n8173;
  assign n8175 = controllable_nhgrant0 & ~n8174;
  assign n8176 = ~controllable_nhgrant0 & ~n7791;
  assign n8177 = ~n8175 & ~n8176;
  assign n8178 = ~controllable_hgrant7 & ~n8177;
  assign n8179 = ~n7793 & ~n8178;
  assign n8180 = ~controllable_hgrant9 & ~n8179;
  assign n8181 = ~n7792 & ~n8180;
  assign n8182 = n7593 & ~n8181;
  assign n8183 = n87 & reg_stateG10_7_out;
  assign n8184 = controllable_hgrant7 & ~n8183;
  assign n8185 = ~i_hbusreq7 & ~n8184;
  assign n8186 = n87 & reg_stateG10_8_out;
  assign n8187 = controllable_hgrant8 & ~n8186;
  assign n8188 = ~i_hbusreq8 & ~n8187;
  assign n8189 = n87 & reg_stateG10_9_out;
  assign n8190 = controllable_hgrant9 & ~n8189;
  assign n8191 = ~i_hbusreq9 & ~n8190;
  assign n8192 = n7594 & ~n7606;
  assign n8193 = n7630 & ~n8192;
  assign n8194 = n7595 & n7720;
  assign n8195 = n7675 & ~n8194;
  assign n8196 = ~n7791 & ~n8195;
  assign n8197 = n7597 & ~n7606;
  assign n8198 = ~n7683 & ~n8197;
  assign n8199 = ~n7629 & ~n8198;
  assign n8200 = n7715 & ~n8199;
  assign n8201 = n7675 & ~n8200;
  assign n8202 = ~n7655 & ~n8201;
  assign n8203 = n7596 & ~n7606;
  assign n8204 = ~n7622 & ~n8203;
  assign n8205 = ~n7683 & ~n8204;
  assign n8206 = ~n7689 & ~n8205;
  assign n8207 = ~n7629 & ~n8206;
  assign n8208 = ~n7615 & ~n8207;
  assign n8209 = ~n7640 & ~n8208;
  assign n8210 = ~n7669 & ~n8209;
  assign n8211 = ~n7674 & ~n8210;
  assign n8212 = ~n7661 & ~n8211;
  assign n8213 = ~n7655 & ~n8212;
  assign n8214 = ~n7646 & ~n8213;
  assign n8215 = n87 & reg_stateG10_6_out;
  assign n8216 = controllable_hgrant6 & ~n8215;
  assign n8217 = ~i_hbusreq6 & ~n8216;
  assign n8218 = controllable_hmastlock & ~n7818;
  assign n8219 = ~n7733 & ~n8218;
  assign n8220 = ~n7733 & ~n8219;
  assign n8221 = ~n7928 & ~n8220;
  assign n8222 = n7928 & ~n8218;
  assign n8223 = ~n8221 & ~n8222;
  assign n8224 = controllable_hmaster2 & ~n8223;
  assign n8225 = controllable_hmaster2 & ~n8224;
  assign n8226 = controllable_hmaster1 & ~n8225;
  assign n8227 = controllable_hmaster1 & ~n8226;
  assign n8228 = ~n8217 & ~n8227;
  assign n8229 = ~n8217 & ~n8228;
  assign n8230 = i_hlock6 & ~n8229;
  assign n8231 = ~controllable_hmastlock & ~n7735;
  assign n8232 = ~controllable_hmastlock & ~n8231;
  assign n8233 = ~n7733 & ~n8232;
  assign n8234 = ~n7733 & ~n8233;
  assign n8235 = ~n7928 & ~n8234;
  assign n8236 = n7928 & ~n8232;
  assign n8237 = ~n8235 & ~n8236;
  assign n8238 = controllable_hmaster2 & ~n8237;
  assign n8239 = controllable_hmaster2 & ~n8238;
  assign n8240 = controllable_hmaster1 & ~n8239;
  assign n8241 = controllable_hmaster1 & ~n8240;
  assign n8242 = ~n8217 & ~n8241;
  assign n8243 = ~n8217 & ~n8242;
  assign n8244 = ~i_hlock6 & ~n8243;
  assign n8245 = ~n8230 & ~n8244;
  assign n8246 = ~controllable_hmaster0 & ~n8245;
  assign n8247 = ~controllable_hmaster0 & ~n8246;
  assign n8248 = ~controllable_hmaster3 & ~n8247;
  assign n8249 = ~controllable_hmaster3 & ~n8248;
  assign n8250 = i_hbusreq7 & ~n8249;
  assign n8251 = i_hbusreq8 & ~n8247;
  assign n8252 = i_hbusreq6 & ~n8245;
  assign n8253 = i_hbusreq5 & ~n8223;
  assign n8254 = i_hbusreq4 & ~n8223;
  assign n8255 = i_hbusreq9 & ~n8223;
  assign n8256 = i_hbusreq3 & ~n8223;
  assign n8257 = i_hbusreq1 & ~n8223;
  assign n8258 = i_hbusreq2 & ~n8218;
  assign n8259 = i_hbusreq0 & ~n8218;
  assign n8260 = i_hbusreq0 & ~n8259;
  assign n8261 = ~i_hbusreq2 & ~n8260;
  assign n8262 = ~n8258 & ~n8261;
  assign n8263 = ~n7733 & ~n8262;
  assign n8264 = ~n7733 & ~n8263;
  assign n8265 = ~n7928 & ~n8264;
  assign n8266 = n7928 & ~n8262;
  assign n8267 = ~n8265 & ~n8266;
  assign n8268 = ~i_hbusreq1 & ~n8267;
  assign n8269 = ~n8257 & ~n8268;
  assign n8270 = ~i_hbusreq3 & ~n8269;
  assign n8271 = ~n8256 & ~n8270;
  assign n8272 = ~i_hbusreq9 & ~n8271;
  assign n8273 = ~n8255 & ~n8272;
  assign n8274 = ~i_hbusreq4 & ~n8273;
  assign n8275 = ~n8254 & ~n8274;
  assign n8276 = ~i_hbusreq5 & ~n8275;
  assign n8277 = ~n8253 & ~n8276;
  assign n8278 = controllable_hmaster2 & ~n8277;
  assign n8279 = controllable_hmaster2 & ~n8278;
  assign n8280 = controllable_hmaster1 & ~n8279;
  assign n8281 = controllable_hmaster1 & ~n8280;
  assign n8282 = ~n8217 & ~n8281;
  assign n8283 = ~n8217 & ~n8282;
  assign n8284 = i_hlock6 & ~n8283;
  assign n8285 = i_hbusreq5 & ~n8237;
  assign n8286 = i_hbusreq4 & ~n8237;
  assign n8287 = i_hbusreq9 & ~n8237;
  assign n8288 = i_hbusreq3 & ~n8237;
  assign n8289 = i_hbusreq1 & ~n8237;
  assign n8290 = i_hbusreq2 & ~n8232;
  assign n8291 = i_hbusreq0 & ~n8232;
  assign n8292 = i_hbusreq0 & ~n8291;
  assign n8293 = ~i_hbusreq2 & ~n8292;
  assign n8294 = ~n8290 & ~n8293;
  assign n8295 = ~n7733 & ~n8294;
  assign n8296 = ~n7733 & ~n8295;
  assign n8297 = ~n7928 & ~n8296;
  assign n8298 = n7928 & ~n8294;
  assign n8299 = ~n8297 & ~n8298;
  assign n8300 = ~i_hbusreq1 & ~n8299;
  assign n8301 = ~n8289 & ~n8300;
  assign n8302 = ~i_hbusreq3 & ~n8301;
  assign n8303 = ~n8288 & ~n8302;
  assign n8304 = ~i_hbusreq9 & ~n8303;
  assign n8305 = ~n8287 & ~n8304;
  assign n8306 = ~i_hbusreq4 & ~n8305;
  assign n8307 = ~n8286 & ~n8306;
  assign n8308 = ~i_hbusreq5 & ~n8307;
  assign n8309 = ~n8285 & ~n8308;
  assign n8310 = controllable_hmaster2 & ~n8309;
  assign n8311 = controllable_hmaster2 & ~n8310;
  assign n8312 = controllable_hmaster1 & ~n8311;
  assign n8313 = controllable_hmaster1 & ~n8312;
  assign n8314 = ~n8217 & ~n8313;
  assign n8315 = ~n8217 & ~n8314;
  assign n8316 = ~i_hlock6 & ~n8315;
  assign n8317 = ~n8284 & ~n8316;
  assign n8318 = ~i_hbusreq6 & ~n8317;
  assign n8319 = ~n8252 & ~n8318;
  assign n8320 = ~controllable_hmaster0 & ~n8319;
  assign n8321 = ~controllable_hmaster0 & ~n8320;
  assign n8322 = ~i_hbusreq8 & ~n8321;
  assign n8323 = ~n8251 & ~n8322;
  assign n8324 = ~controllable_hmaster3 & ~n8323;
  assign n8325 = ~controllable_hmaster3 & ~n8324;
  assign n8326 = ~i_hbusreq7 & ~n8325;
  assign n8327 = ~n8250 & ~n8326;
  assign n8328 = n7924 & ~n8327;
  assign n8329 = n7924 & ~n8328;
  assign n8330 = n8214 & ~n8329;
  assign n8331 = n8214 & ~n8330;
  assign n8332 = n8202 & ~n8331;
  assign n8333 = n8202 & ~n8332;
  assign n8334 = n7728 & ~n8333;
  assign n8335 = ~n7782 & ~n8202;
  assign n8336 = ~n7782 & ~n8214;
  assign n8337 = ~n7782 & ~n7924;
  assign n8338 = ~n7743 & ~n8248;
  assign n8339 = i_hbusreq7 & ~n8338;
  assign n8340 = ~n7779 & ~n8324;
  assign n8341 = ~i_hbusreq7 & ~n8340;
  assign n8342 = ~n8339 & ~n8341;
  assign n8343 = n7924 & ~n8342;
  assign n8344 = ~n8337 & ~n8343;
  assign n8345 = n8214 & ~n8344;
  assign n8346 = ~n8336 & ~n8345;
  assign n8347 = n8202 & ~n8346;
  assign n8348 = ~n8335 & ~n8347;
  assign n8349 = ~n7728 & ~n8348;
  assign n8350 = ~n8334 & ~n8349;
  assign n8351 = ~n7723 & ~n8350;
  assign n8352 = ~n7723 & ~n8351;
  assign n8353 = ~n7714 & ~n8352;
  assign n8354 = ~n7714 & ~n8353;
  assign n8355 = n7705 & ~n8354;
  assign n8356 = n7723 & ~n8348;
  assign n8357 = controllable_hmaster1 & ~n7735;
  assign n8358 = controllable_hmaster2 & ~n7735;
  assign n8359 = controllable_hmaster2 & ~n8358;
  assign n8360 = ~controllable_hmaster1 & ~n8359;
  assign n8361 = ~n8357 & ~n8360;
  assign n8362 = controllable_hmaster3 & ~n8361;
  assign n8363 = n87 & reg_stateG10_3_out;
  assign n8364 = controllable_hgrant3 & ~n8363;
  assign n8365 = ~i_hbusreq3 & ~n8364;
  assign n8366 = ~n8223 & ~n8365;
  assign n8367 = ~n8365 & ~n8366;
  assign n8368 = i_hlock3 & ~n8367;
  assign n8369 = ~n8237 & ~n8365;
  assign n8370 = ~n8365 & ~n8369;
  assign n8371 = ~i_hlock3 & ~n8370;
  assign n8372 = ~n8368 & ~n8371;
  assign n8373 = ~controllable_hmaster2 & ~n8372;
  assign n8374 = ~controllable_hmaster2 & ~n8373;
  assign n8375 = controllable_hmaster1 & ~n8374;
  assign n8376 = n87 & reg_stateG10_5_out;
  assign n8377 = controllable_hgrant5 & ~n8376;
  assign n8378 = ~i_hbusreq5 & ~n8377;
  assign n8379 = ~n8223 & ~n8378;
  assign n8380 = ~n8378 & ~n8379;
  assign n8381 = i_hlock5 & ~n8380;
  assign n8382 = ~n8237 & ~n8378;
  assign n8383 = ~n8378 & ~n8382;
  assign n8384 = ~i_hlock5 & ~n8383;
  assign n8385 = ~n8381 & ~n8384;
  assign n8386 = controllable_hmaster2 & ~n8385;
  assign n8387 = n87 & reg_stateG10_1_out;
  assign n8388 = controllable_hgrant1 & ~n8387;
  assign n8389 = ~i_hbusreq1 & ~n8388;
  assign n8390 = ~n8223 & ~n8389;
  assign n8391 = ~n8389 & ~n8390;
  assign n8392 = i_hlock1 & ~n8391;
  assign n8393 = ~n8237 & ~n8389;
  assign n8394 = ~n8389 & ~n8393;
  assign n8395 = ~i_hlock1 & ~n8394;
  assign n8396 = ~n8392 & ~n8395;
  assign n8397 = ~controllable_hmaster2 & ~n8396;
  assign n8398 = ~n8386 & ~n8397;
  assign n8399 = ~controllable_hmaster1 & ~n8398;
  assign n8400 = ~n8375 & ~n8399;
  assign n8401 = controllable_hmaster0 & ~n8400;
  assign n8402 = n87 & reg_stateG10_2_out;
  assign n8403 = controllable_hgrant2 & ~n8402;
  assign n8404 = ~i_hbusreq2 & ~n8403;
  assign n8405 = i_hready & ~n8404;
  assign n8406 = ~n8404 & ~n8405;
  assign n8407 = ~controllable_ndecide & ~n8406;
  assign n8408 = ~controllable_ndecide & ~n8407;
  assign n8409 = controllable_hmastlock & ~n8408;
  assign n8410 = controllable_hmastlock & ~n8409;
  assign n8411 = i_hlock2 & ~n8410;
  assign n8412 = ~controllable_hmastlock & ~n8408;
  assign n8413 = ~controllable_hmastlock & ~n8412;
  assign n8414 = ~i_hlock2 & ~n8413;
  assign n8415 = ~n8411 & ~n8414;
  assign n8416 = ~n7733 & ~n8415;
  assign n8417 = ~n7733 & ~n8416;
  assign n8418 = ~n7928 & ~n8417;
  assign n8419 = n7928 & ~n8415;
  assign n8420 = ~n8418 & ~n8419;
  assign n8421 = ~controllable_hmaster2 & ~n8420;
  assign n8422 = ~controllable_hmaster2 & ~n8421;
  assign n8423 = controllable_hmaster1 & ~n8422;
  assign n8424 = n87 & reg_stateG10_4_out;
  assign n8425 = controllable_hgrant4 & ~n8424;
  assign n8426 = ~i_hbusreq4 & ~n8425;
  assign n8427 = ~n8223 & ~n8426;
  assign n8428 = ~n8426 & ~n8427;
  assign n8429 = i_hlock4 & ~n8428;
  assign n8430 = ~n8237 & ~n8426;
  assign n8431 = ~n8426 & ~n8430;
  assign n8432 = ~i_hlock4 & ~n8431;
  assign n8433 = ~n8429 & ~n8432;
  assign n8434 = controllable_hmaster2 & ~n8433;
  assign n8435 = i_hlock0 & ~n8218;
  assign n8436 = ~i_hlock0 & ~n8232;
  assign n8437 = ~n8435 & ~n8436;
  assign n8438 = ~n7733 & ~n8437;
  assign n8439 = ~n7733 & ~n8438;
  assign n8440 = ~n7928 & ~n8439;
  assign n8441 = n7928 & ~n8437;
  assign n8442 = ~n8440 & ~n8441;
  assign n8443 = ~controllable_hmaster2 & ~n8442;
  assign n8444 = ~n8434 & ~n8443;
  assign n8445 = ~controllable_hmaster1 & ~n8444;
  assign n8446 = ~n8423 & ~n8445;
  assign n8447 = n8217 & ~n8446;
  assign n8448 = ~n8224 & ~n8421;
  assign n8449 = controllable_hmaster1 & ~n8448;
  assign n8450 = ~n8445 & ~n8449;
  assign n8451 = ~n8217 & ~n8450;
  assign n8452 = ~n8447 & ~n8451;
  assign n8453 = i_hlock6 & ~n8452;
  assign n8454 = ~n8238 & ~n8421;
  assign n8455 = controllable_hmaster1 & ~n8454;
  assign n8456 = ~n8445 & ~n8455;
  assign n8457 = ~n8217 & ~n8456;
  assign n8458 = ~n8447 & ~n8457;
  assign n8459 = ~i_hlock6 & ~n8458;
  assign n8460 = ~n8453 & ~n8459;
  assign n8461 = ~controllable_hmaster0 & ~n8460;
  assign n8462 = ~n8401 & ~n8461;
  assign n8463 = ~controllable_hmaster3 & ~n8462;
  assign n8464 = ~n8362 & ~n8463;
  assign n8465 = i_hbusreq7 & ~n8464;
  assign n8466 = i_hbusreq8 & ~n8361;
  assign n8467 = i_hbusreq6 & ~n8361;
  assign n8468 = i_hbusreq5 & ~n7735;
  assign n8469 = i_hbusreq4 & ~n7735;
  assign n8470 = i_hbusreq9 & ~n7735;
  assign n8471 = i_hbusreq3 & ~n7735;
  assign n8472 = i_hbusreq1 & ~n7735;
  assign n8473 = ~i_hbusreq1 & ~n7757;
  assign n8474 = ~n8472 & ~n8473;
  assign n8475 = ~i_hbusreq3 & ~n8474;
  assign n8476 = ~n8471 & ~n8475;
  assign n8477 = ~i_hbusreq9 & ~n8476;
  assign n8478 = ~n8470 & ~n8477;
  assign n8479 = ~i_hbusreq4 & ~n8478;
  assign n8480 = ~n8469 & ~n8479;
  assign n8481 = ~i_hbusreq5 & ~n8480;
  assign n8482 = ~n8468 & ~n8481;
  assign n8483 = controllable_hmaster1 & ~n8482;
  assign n8484 = controllable_hmaster2 & ~n8482;
  assign n8485 = controllable_hmaster2 & ~n8484;
  assign n8486 = ~controllable_hmaster1 & ~n8485;
  assign n8487 = ~n8483 & ~n8486;
  assign n8488 = ~i_hbusreq6 & ~n8487;
  assign n8489 = ~n8467 & ~n8488;
  assign n8490 = ~i_hbusreq8 & ~n8489;
  assign n8491 = ~n8466 & ~n8490;
  assign n8492 = controllable_hmaster3 & ~n8491;
  assign n8493 = i_hbusreq8 & ~n8462;
  assign n8494 = i_hbusreq6 & ~n8400;
  assign n8495 = i_hbusreq5 & ~n8372;
  assign n8496 = i_hbusreq4 & ~n8372;
  assign n8497 = i_hbusreq9 & ~n8372;
  assign n8498 = i_hbusreq3 & ~n8372;
  assign n8499 = ~n8269 & ~n8365;
  assign n8500 = ~n8365 & ~n8499;
  assign n8501 = i_hlock3 & ~n8500;
  assign n8502 = ~n8301 & ~n8365;
  assign n8503 = ~n8365 & ~n8502;
  assign n8504 = ~i_hlock3 & ~n8503;
  assign n8505 = ~n8501 & ~n8504;
  assign n8506 = ~i_hbusreq3 & ~n8505;
  assign n8507 = ~n8498 & ~n8506;
  assign n8508 = ~i_hbusreq9 & ~n8507;
  assign n8509 = ~n8497 & ~n8508;
  assign n8510 = ~i_hbusreq4 & ~n8509;
  assign n8511 = ~n8496 & ~n8510;
  assign n8512 = ~i_hbusreq5 & ~n8511;
  assign n8513 = ~n8495 & ~n8512;
  assign n8514 = ~controllable_hmaster2 & ~n8513;
  assign n8515 = ~controllable_hmaster2 & ~n8514;
  assign n8516 = controllable_hmaster1 & ~n8515;
  assign n8517 = i_hbusreq5 & ~n8385;
  assign n8518 = ~n8275 & ~n8378;
  assign n8519 = ~n8378 & ~n8518;
  assign n8520 = i_hlock5 & ~n8519;
  assign n8521 = ~n8307 & ~n8378;
  assign n8522 = ~n8378 & ~n8521;
  assign n8523 = ~i_hlock5 & ~n8522;
  assign n8524 = ~n8520 & ~n8523;
  assign n8525 = ~i_hbusreq5 & ~n8524;
  assign n8526 = ~n8517 & ~n8525;
  assign n8527 = controllable_hmaster2 & ~n8526;
  assign n8528 = i_hbusreq5 & ~n8396;
  assign n8529 = i_hbusreq4 & ~n8396;
  assign n8530 = i_hbusreq9 & ~n8396;
  assign n8531 = i_hbusreq3 & ~n8396;
  assign n8532 = i_hbusreq1 & ~n8396;
  assign n8533 = ~n8267 & ~n8389;
  assign n8534 = ~n8389 & ~n8533;
  assign n8535 = i_hlock1 & ~n8534;
  assign n8536 = ~n8299 & ~n8389;
  assign n8537 = ~n8389 & ~n8536;
  assign n8538 = ~i_hlock1 & ~n8537;
  assign n8539 = ~n8535 & ~n8538;
  assign n8540 = ~i_hbusreq1 & ~n8539;
  assign n8541 = ~n8532 & ~n8540;
  assign n8542 = ~i_hbusreq3 & ~n8541;
  assign n8543 = ~n8531 & ~n8542;
  assign n8544 = ~i_hbusreq9 & ~n8543;
  assign n8545 = ~n8530 & ~n8544;
  assign n8546 = ~i_hbusreq4 & ~n8545;
  assign n8547 = ~n8529 & ~n8546;
  assign n8548 = ~i_hbusreq5 & ~n8547;
  assign n8549 = ~n8528 & ~n8548;
  assign n8550 = ~controllable_hmaster2 & ~n8549;
  assign n8551 = ~n8527 & ~n8550;
  assign n8552 = ~controllable_hmaster1 & ~n8551;
  assign n8553 = ~n8516 & ~n8552;
  assign n8554 = ~i_hbusreq6 & ~n8553;
  assign n8555 = ~n8494 & ~n8554;
  assign n8556 = controllable_hmaster0 & ~n8555;
  assign n8557 = i_hbusreq6 & ~n8460;
  assign n8558 = i_hbusreq5 & ~n8420;
  assign n8559 = i_hbusreq4 & ~n8420;
  assign n8560 = i_hbusreq9 & ~n8420;
  assign n8561 = i_hbusreq3 & ~n8420;
  assign n8562 = i_hbusreq1 & ~n8420;
  assign n8563 = i_hbusreq2 & ~n8415;
  assign n8564 = i_hbusreq0 & ~n8410;
  assign n8565 = i_hbusreq0 & ~n8564;
  assign n8566 = i_hlock2 & ~n8565;
  assign n8567 = i_hbusreq0 & ~n8413;
  assign n8568 = i_hbusreq0 & ~n8567;
  assign n8569 = ~i_hlock2 & ~n8568;
  assign n8570 = ~n8566 & ~n8569;
  assign n8571 = ~i_hbusreq2 & ~n8570;
  assign n8572 = ~n8563 & ~n8571;
  assign n8573 = ~n7733 & ~n8572;
  assign n8574 = ~n7733 & ~n8573;
  assign n8575 = ~n7928 & ~n8574;
  assign n8576 = n7928 & ~n8572;
  assign n8577 = ~n8575 & ~n8576;
  assign n8578 = ~i_hbusreq1 & ~n8577;
  assign n8579 = ~n8562 & ~n8578;
  assign n8580 = ~i_hbusreq3 & ~n8579;
  assign n8581 = ~n8561 & ~n8580;
  assign n8582 = ~i_hbusreq9 & ~n8581;
  assign n8583 = ~n8560 & ~n8582;
  assign n8584 = ~i_hbusreq4 & ~n8583;
  assign n8585 = ~n8559 & ~n8584;
  assign n8586 = ~i_hbusreq5 & ~n8585;
  assign n8587 = ~n8558 & ~n8586;
  assign n8588 = ~controllable_hmaster2 & ~n8587;
  assign n8589 = ~controllable_hmaster2 & ~n8588;
  assign n8590 = controllable_hmaster1 & ~n8589;
  assign n8591 = i_hbusreq5 & ~n8433;
  assign n8592 = i_hbusreq4 & ~n8433;
  assign n8593 = i_hbusreq9 & ~n8428;
  assign n8594 = ~n8271 & ~n8426;
  assign n8595 = ~n8426 & ~n8594;
  assign n8596 = ~i_hbusreq9 & ~n8595;
  assign n8597 = ~n8593 & ~n8596;
  assign n8598 = i_hlock4 & ~n8597;
  assign n8599 = i_hbusreq9 & ~n8431;
  assign n8600 = ~n8303 & ~n8426;
  assign n8601 = ~n8426 & ~n8600;
  assign n8602 = ~i_hbusreq9 & ~n8601;
  assign n8603 = ~n8599 & ~n8602;
  assign n8604 = ~i_hlock4 & ~n8603;
  assign n8605 = ~n8598 & ~n8604;
  assign n8606 = ~i_hbusreq4 & ~n8605;
  assign n8607 = ~n8592 & ~n8606;
  assign n8608 = ~i_hbusreq5 & ~n8607;
  assign n8609 = ~n8591 & ~n8608;
  assign n8610 = controllable_hmaster2 & ~n8609;
  assign n8611 = ~n8443 & ~n8610;
  assign n8612 = ~controllable_hmaster1 & ~n8611;
  assign n8613 = ~n8590 & ~n8612;
  assign n8614 = n8217 & ~n8613;
  assign n8615 = ~n8278 & ~n8588;
  assign n8616 = controllable_hmaster1 & ~n8615;
  assign n8617 = ~n8612 & ~n8616;
  assign n8618 = ~n8217 & ~n8617;
  assign n8619 = ~n8614 & ~n8618;
  assign n8620 = i_hlock6 & ~n8619;
  assign n8621 = ~n8310 & ~n8588;
  assign n8622 = controllable_hmaster1 & ~n8621;
  assign n8623 = ~n8612 & ~n8622;
  assign n8624 = ~n8217 & ~n8623;
  assign n8625 = ~n8614 & ~n8624;
  assign n8626 = ~i_hlock6 & ~n8625;
  assign n8627 = ~n8620 & ~n8626;
  assign n8628 = ~i_hbusreq6 & ~n8627;
  assign n8629 = ~n8557 & ~n8628;
  assign n8630 = ~controllable_hmaster0 & ~n8629;
  assign n8631 = ~n8556 & ~n8630;
  assign n8632 = ~i_hbusreq8 & ~n8631;
  assign n8633 = ~n8493 & ~n8632;
  assign n8634 = ~controllable_hmaster3 & ~n8633;
  assign n8635 = ~n8492 & ~n8634;
  assign n8636 = ~i_hbusreq7 & ~n8635;
  assign n8637 = ~n8465 & ~n8636;
  assign n8638 = n7924 & ~n8637;
  assign n8639 = ~n8337 & ~n8638;
  assign n8640 = ~n7920 & ~n8639;
  assign n8641 = n7920 & ~n8348;
  assign n8642 = ~n8640 & ~n8641;
  assign n8643 = ~n7723 & ~n8642;
  assign n8644 = ~n8356 & ~n8643;
  assign n8645 = n7714 & ~n8644;
  assign n8646 = ~n7714 & ~n8639;
  assign n8647 = ~n8645 & ~n8646;
  assign n8648 = ~n7705 & ~n8647;
  assign n8649 = ~n8355 & ~n8648;
  assign n8650 = ~n7808 & ~n8649;
  assign n8651 = ~n7920 & ~n8333;
  assign n8652 = ~n7735 & n7928;
  assign n8653 = ~n8221 & ~n8652;
  assign n8654 = i_hlock9 & ~n8653;
  assign n8655 = ~n8235 & ~n8652;
  assign n8656 = ~i_hlock9 & ~n8655;
  assign n8657 = ~n8654 & ~n8656;
  assign n8658 = ~controllable_hmaster2 & ~n8657;
  assign n8659 = ~controllable_hmaster2 & ~n8658;
  assign n8660 = ~controllable_hmaster1 & ~n8659;
  assign n8661 = ~controllable_hmaster1 & ~n8660;
  assign n8662 = controllable_hmaster0 & ~n8661;
  assign n8663 = controllable_hmaster0 & ~n8662;
  assign n8664 = controllable_hmaster3 & ~n8663;
  assign n8665 = controllable_hmaster3 & ~n8664;
  assign n8666 = i_hbusreq7 & ~n8665;
  assign n8667 = i_hbusreq8 & ~n8663;
  assign n8668 = i_hbusreq6 & ~n8661;
  assign n8669 = i_hbusreq5 & ~n8657;
  assign n8670 = i_hbusreq4 & ~n8657;
  assign n8671 = i_hbusreq9 & ~n8657;
  assign n8672 = i_hbusreq3 & ~n8653;
  assign n8673 = i_hbusreq1 & ~n8653;
  assign n8674 = ~i_hlock0 & ~n7735;
  assign n8675 = ~i_hlock0 & ~n8674;
  assign n8676 = ~i_hbusreq0 & ~n8675;
  assign n8677 = ~n7754 & ~n8676;
  assign n8678 = ~i_hbusreq2 & ~n8677;
  assign n8679 = ~n7753 & ~n8678;
  assign n8680 = ~n7733 & ~n8679;
  assign n8681 = i_hlock0 & ~n8232;
  assign n8682 = ~n8674 & ~n8681;
  assign n8683 = ~i_hbusreq0 & ~n8682;
  assign n8684 = ~n7754 & ~n8683;
  assign n8685 = ~i_hbusreq2 & ~n8684;
  assign n8686 = ~n7753 & ~n8685;
  assign n8687 = n7733 & ~n8686;
  assign n8688 = ~n8680 & ~n8687;
  assign n8689 = n7928 & ~n8688;
  assign n8690 = ~n8265 & ~n8689;
  assign n8691 = ~i_hbusreq1 & ~n8690;
  assign n8692 = ~n8673 & ~n8691;
  assign n8693 = ~i_hbusreq3 & ~n8692;
  assign n8694 = ~n8672 & ~n8693;
  assign n8695 = i_hlock9 & ~n8694;
  assign n8696 = i_hbusreq3 & ~n8655;
  assign n8697 = i_hbusreq1 & ~n8655;
  assign n8698 = ~n8297 & ~n8689;
  assign n8699 = ~i_hbusreq1 & ~n8698;
  assign n8700 = ~n8697 & ~n8699;
  assign n8701 = ~i_hbusreq3 & ~n8700;
  assign n8702 = ~n8696 & ~n8701;
  assign n8703 = ~i_hlock9 & ~n8702;
  assign n8704 = ~n8695 & ~n8703;
  assign n8705 = ~i_hbusreq9 & ~n8704;
  assign n8706 = ~n8671 & ~n8705;
  assign n8707 = ~i_hbusreq4 & ~n8706;
  assign n8708 = ~n8670 & ~n8707;
  assign n8709 = ~i_hbusreq5 & ~n8708;
  assign n8710 = ~n8669 & ~n8709;
  assign n8711 = ~controllable_hmaster2 & ~n8710;
  assign n8712 = ~controllable_hmaster2 & ~n8711;
  assign n8713 = ~controllable_hmaster1 & ~n8712;
  assign n8714 = ~controllable_hmaster1 & ~n8713;
  assign n8715 = ~i_hbusreq6 & ~n8714;
  assign n8716 = ~n8668 & ~n8715;
  assign n8717 = controllable_hmaster0 & ~n8716;
  assign n8718 = controllable_hmaster0 & ~n8717;
  assign n8719 = ~i_hbusreq8 & ~n8718;
  assign n8720 = ~n8667 & ~n8719;
  assign n8721 = controllable_hmaster3 & ~n8720;
  assign n8722 = controllable_hmaster3 & ~n8721;
  assign n8723 = ~i_hbusreq7 & ~n8722;
  assign n8724 = ~n8666 & ~n8723;
  assign n8725 = ~n8214 & ~n8724;
  assign n8726 = ~controllable_hmaster2 & ~n8653;
  assign n8727 = ~controllable_hmaster2 & ~n8726;
  assign n8728 = ~controllable_hmaster1 & ~n8727;
  assign n8729 = ~controllable_hmaster1 & ~n8728;
  assign n8730 = ~controllable_hmaster0 & ~n8729;
  assign n8731 = ~controllable_hmaster0 & ~n8730;
  assign n8732 = i_hlock8 & ~n8731;
  assign n8733 = ~controllable_hmaster2 & ~n8655;
  assign n8734 = ~controllable_hmaster2 & ~n8733;
  assign n8735 = ~controllable_hmaster1 & ~n8734;
  assign n8736 = ~controllable_hmaster1 & ~n8735;
  assign n8737 = ~controllable_hmaster0 & ~n8736;
  assign n8738 = ~controllable_hmaster0 & ~n8737;
  assign n8739 = ~i_hlock8 & ~n8738;
  assign n8740 = ~n8732 & ~n8739;
  assign n8741 = controllable_hmaster3 & ~n8740;
  assign n8742 = controllable_hmaster3 & ~n8741;
  assign n8743 = i_hbusreq7 & ~n8742;
  assign n8744 = i_hbusreq8 & ~n8740;
  assign n8745 = i_hbusreq6 & ~n8729;
  assign n8746 = i_hbusreq5 & ~n8653;
  assign n8747 = i_hbusreq4 & ~n8653;
  assign n8748 = i_hbusreq9 & ~n8653;
  assign n8749 = ~i_hbusreq9 & ~n8694;
  assign n8750 = ~n8748 & ~n8749;
  assign n8751 = ~i_hbusreq4 & ~n8750;
  assign n8752 = ~n8747 & ~n8751;
  assign n8753 = ~i_hbusreq5 & ~n8752;
  assign n8754 = ~n8746 & ~n8753;
  assign n8755 = ~controllable_hmaster2 & ~n8754;
  assign n8756 = ~controllable_hmaster2 & ~n8755;
  assign n8757 = ~controllable_hmaster1 & ~n8756;
  assign n8758 = ~controllable_hmaster1 & ~n8757;
  assign n8759 = ~i_hbusreq6 & ~n8758;
  assign n8760 = ~n8745 & ~n8759;
  assign n8761 = ~controllable_hmaster0 & ~n8760;
  assign n8762 = ~controllable_hmaster0 & ~n8761;
  assign n8763 = i_hlock8 & ~n8762;
  assign n8764 = i_hbusreq6 & ~n8736;
  assign n8765 = i_hbusreq5 & ~n8655;
  assign n8766 = i_hbusreq4 & ~n8655;
  assign n8767 = i_hbusreq9 & ~n8655;
  assign n8768 = ~i_hbusreq9 & ~n8702;
  assign n8769 = ~n8767 & ~n8768;
  assign n8770 = ~i_hbusreq4 & ~n8769;
  assign n8771 = ~n8766 & ~n8770;
  assign n8772 = ~i_hbusreq5 & ~n8771;
  assign n8773 = ~n8765 & ~n8772;
  assign n8774 = ~controllable_hmaster2 & ~n8773;
  assign n8775 = ~controllable_hmaster2 & ~n8774;
  assign n8776 = ~controllable_hmaster1 & ~n8775;
  assign n8777 = ~controllable_hmaster1 & ~n8776;
  assign n8778 = ~i_hbusreq6 & ~n8777;
  assign n8779 = ~n8764 & ~n8778;
  assign n8780 = ~controllable_hmaster0 & ~n8779;
  assign n8781 = ~controllable_hmaster0 & ~n8780;
  assign n8782 = ~i_hlock8 & ~n8781;
  assign n8783 = ~n8763 & ~n8782;
  assign n8784 = ~i_hbusreq8 & ~n8783;
  assign n8785 = ~n8744 & ~n8784;
  assign n8786 = controllable_hmaster3 & ~n8785;
  assign n8787 = controllable_hmaster3 & ~n8786;
  assign n8788 = ~i_hbusreq7 & ~n8787;
  assign n8789 = ~n8743 & ~n8788;
  assign n8790 = n8214 & ~n8789;
  assign n8791 = ~n8725 & ~n8790;
  assign n8792 = ~n8202 & ~n8791;
  assign n8793 = controllable_hmaster2 & ~n8653;
  assign n8794 = controllable_hmaster2 & ~n8793;
  assign n8795 = controllable_hmaster1 & ~n8794;
  assign n8796 = controllable_hmaster1 & ~n8795;
  assign n8797 = controllable_hmaster0 & ~n8796;
  assign n8798 = controllable_hmaster0 & ~n8797;
  assign n8799 = ~controllable_hmaster3 & ~n8798;
  assign n8800 = ~controllable_hmaster3 & ~n8799;
  assign n8801 = i_hlock7 & ~n8800;
  assign n8802 = controllable_hmaster2 & ~n8655;
  assign n8803 = controllable_hmaster2 & ~n8802;
  assign n8804 = controllable_hmaster1 & ~n8803;
  assign n8805 = controllable_hmaster1 & ~n8804;
  assign n8806 = controllable_hmaster0 & ~n8805;
  assign n8807 = controllable_hmaster0 & ~n8806;
  assign n8808 = ~controllable_hmaster3 & ~n8807;
  assign n8809 = ~controllable_hmaster3 & ~n8808;
  assign n8810 = ~i_hlock7 & ~n8809;
  assign n8811 = ~n8801 & ~n8810;
  assign n8812 = i_hbusreq7 & ~n8811;
  assign n8813 = i_hbusreq8 & ~n8798;
  assign n8814 = i_hbusreq6 & ~n8796;
  assign n8815 = controllable_hmaster2 & ~n8754;
  assign n8816 = controllable_hmaster2 & ~n8815;
  assign n8817 = controllable_hmaster1 & ~n8816;
  assign n8818 = controllable_hmaster1 & ~n8817;
  assign n8819 = ~i_hbusreq6 & ~n8818;
  assign n8820 = ~n8814 & ~n8819;
  assign n8821 = controllable_hmaster0 & ~n8820;
  assign n8822 = controllable_hmaster0 & ~n8821;
  assign n8823 = ~i_hbusreq8 & ~n8822;
  assign n8824 = ~n8813 & ~n8823;
  assign n8825 = ~controllable_hmaster3 & ~n8824;
  assign n8826 = ~controllable_hmaster3 & ~n8825;
  assign n8827 = i_hlock7 & ~n8826;
  assign n8828 = i_hbusreq8 & ~n8807;
  assign n8829 = i_hbusreq6 & ~n8805;
  assign n8830 = controllable_hmaster2 & ~n8773;
  assign n8831 = controllable_hmaster2 & ~n8830;
  assign n8832 = controllable_hmaster1 & ~n8831;
  assign n8833 = controllable_hmaster1 & ~n8832;
  assign n8834 = ~i_hbusreq6 & ~n8833;
  assign n8835 = ~n8829 & ~n8834;
  assign n8836 = controllable_hmaster0 & ~n8835;
  assign n8837 = controllable_hmaster0 & ~n8836;
  assign n8838 = ~i_hbusreq8 & ~n8837;
  assign n8839 = ~n8828 & ~n8838;
  assign n8840 = ~controllable_hmaster3 & ~n8839;
  assign n8841 = ~controllable_hmaster3 & ~n8840;
  assign n8842 = ~i_hlock7 & ~n8841;
  assign n8843 = ~n8827 & ~n8842;
  assign n8844 = ~i_hbusreq7 & ~n8843;
  assign n8845 = ~n8812 & ~n8844;
  assign n8846 = ~n8214 & ~n8845;
  assign n8847 = i_hlock6 & ~n8796;
  assign n8848 = ~i_hlock6 & ~n8805;
  assign n8849 = ~n8847 & ~n8848;
  assign n8850 = ~controllable_hmaster0 & ~n8849;
  assign n8851 = ~controllable_hmaster0 & ~n8850;
  assign n8852 = ~controllable_hmaster3 & ~n8851;
  assign n8853 = ~controllable_hmaster3 & ~n8852;
  assign n8854 = i_hbusreq7 & ~n8853;
  assign n8855 = i_hbusreq8 & ~n8851;
  assign n8856 = i_hbusreq6 & ~n8849;
  assign n8857 = i_hlock6 & ~n8818;
  assign n8858 = ~i_hlock6 & ~n8833;
  assign n8859 = ~n8857 & ~n8858;
  assign n8860 = ~i_hbusreq6 & ~n8859;
  assign n8861 = ~n8856 & ~n8860;
  assign n8862 = ~controllable_hmaster0 & ~n8861;
  assign n8863 = ~controllable_hmaster0 & ~n8862;
  assign n8864 = ~i_hbusreq8 & ~n8863;
  assign n8865 = ~n8855 & ~n8864;
  assign n8866 = ~controllable_hmaster3 & ~n8865;
  assign n8867 = ~controllable_hmaster3 & ~n8866;
  assign n8868 = ~i_hbusreq7 & ~n8867;
  assign n8869 = ~n8854 & ~n8868;
  assign n8870 = n8214 & ~n8869;
  assign n8871 = ~n8846 & ~n8870;
  assign n8872 = n8202 & ~n8871;
  assign n8873 = ~n8792 & ~n8872;
  assign n8874 = n7920 & ~n8873;
  assign n8875 = ~n8651 & ~n8874;
  assign n8876 = n7728 & ~n8875;
  assign n8877 = ~n7920 & ~n8348;
  assign n8878 = ~n7739 & ~n8658;
  assign n8879 = ~controllable_hmaster1 & ~n8878;
  assign n8880 = ~n7738 & ~n8879;
  assign n8881 = controllable_hmaster0 & ~n8880;
  assign n8882 = ~controllable_hmaster0 & ~n7742;
  assign n8883 = ~n8881 & ~n8882;
  assign n8884 = controllable_hmaster3 & ~n8883;
  assign n8885 = controllable_hmaster3 & ~n8884;
  assign n8886 = i_hbusreq7 & ~n8885;
  assign n8887 = i_hbusreq8 & ~n8883;
  assign n8888 = i_hbusreq6 & ~n8880;
  assign n8889 = ~n7771 & ~n8711;
  assign n8890 = ~controllable_hmaster1 & ~n8889;
  assign n8891 = ~n7770 & ~n8890;
  assign n8892 = ~i_hbusreq6 & ~n8891;
  assign n8893 = ~n8888 & ~n8892;
  assign n8894 = controllable_hmaster0 & ~n8893;
  assign n8895 = ~controllable_hmaster0 & ~n7776;
  assign n8896 = ~n8894 & ~n8895;
  assign n8897 = ~i_hbusreq8 & ~n8896;
  assign n8898 = ~n8887 & ~n8897;
  assign n8899 = controllable_hmaster3 & ~n8898;
  assign n8900 = controllable_hmaster3 & ~n8899;
  assign n8901 = ~i_hbusreq7 & ~n8900;
  assign n8902 = ~n8886 & ~n8901;
  assign n8903 = ~n8214 & ~n8902;
  assign n8904 = controllable_hmaster0 & ~n7742;
  assign n8905 = ~n7739 & ~n8726;
  assign n8906 = ~controllable_hmaster1 & ~n8905;
  assign n8907 = ~n7738 & ~n8906;
  assign n8908 = ~controllable_hmaster0 & ~n8907;
  assign n8909 = ~n8904 & ~n8908;
  assign n8910 = i_hlock8 & ~n8909;
  assign n8911 = ~n7739 & ~n8733;
  assign n8912 = ~controllable_hmaster1 & ~n8911;
  assign n8913 = ~n7738 & ~n8912;
  assign n8914 = ~controllable_hmaster0 & ~n8913;
  assign n8915 = ~n8904 & ~n8914;
  assign n8916 = ~i_hlock8 & ~n8915;
  assign n8917 = ~n8910 & ~n8916;
  assign n8918 = controllable_hmaster3 & ~n8917;
  assign n8919 = controllable_hmaster3 & ~n8918;
  assign n8920 = i_hbusreq7 & ~n8919;
  assign n8921 = i_hbusreq8 & ~n8917;
  assign n8922 = controllable_hmaster0 & ~n7776;
  assign n8923 = i_hbusreq6 & ~n8907;
  assign n8924 = ~n7771 & ~n8755;
  assign n8925 = ~controllable_hmaster1 & ~n8924;
  assign n8926 = ~n7770 & ~n8925;
  assign n8927 = ~i_hbusreq6 & ~n8926;
  assign n8928 = ~n8923 & ~n8927;
  assign n8929 = ~controllable_hmaster0 & ~n8928;
  assign n8930 = ~n8922 & ~n8929;
  assign n8931 = i_hlock8 & ~n8930;
  assign n8932 = i_hbusreq6 & ~n8913;
  assign n8933 = ~n7771 & ~n8774;
  assign n8934 = ~controllable_hmaster1 & ~n8933;
  assign n8935 = ~n7770 & ~n8934;
  assign n8936 = ~i_hbusreq6 & ~n8935;
  assign n8937 = ~n8932 & ~n8936;
  assign n8938 = ~controllable_hmaster0 & ~n8937;
  assign n8939 = ~n8922 & ~n8938;
  assign n8940 = ~i_hlock8 & ~n8939;
  assign n8941 = ~n8931 & ~n8940;
  assign n8942 = ~i_hbusreq8 & ~n8941;
  assign n8943 = ~n8921 & ~n8942;
  assign n8944 = controllable_hmaster3 & ~n8943;
  assign n8945 = controllable_hmaster3 & ~n8944;
  assign n8946 = ~i_hbusreq7 & ~n8945;
  assign n8947 = ~n8920 & ~n8946;
  assign n8948 = n8214 & ~n8947;
  assign n8949 = ~n8903 & ~n8948;
  assign n8950 = ~n8202 & ~n8949;
  assign n8951 = ~n7743 & ~n8799;
  assign n8952 = i_hlock7 & ~n8951;
  assign n8953 = ~n7743 & ~n8808;
  assign n8954 = ~i_hlock7 & ~n8953;
  assign n8955 = ~n8952 & ~n8954;
  assign n8956 = i_hbusreq7 & ~n8955;
  assign n8957 = ~n7779 & ~n8825;
  assign n8958 = i_hlock7 & ~n8957;
  assign n8959 = ~n7779 & ~n8840;
  assign n8960 = ~i_hlock7 & ~n8959;
  assign n8961 = ~n8958 & ~n8960;
  assign n8962 = ~i_hbusreq7 & ~n8961;
  assign n8963 = ~n8956 & ~n8962;
  assign n8964 = ~n8214 & ~n8963;
  assign n8965 = ~n7743 & ~n8852;
  assign n8966 = i_hbusreq7 & ~n8965;
  assign n8967 = ~n7779 & ~n8866;
  assign n8968 = ~i_hbusreq7 & ~n8967;
  assign n8969 = ~n8966 & ~n8968;
  assign n8970 = n8214 & ~n8969;
  assign n8971 = ~n8964 & ~n8970;
  assign n8972 = n8202 & ~n8971;
  assign n8973 = ~n8950 & ~n8972;
  assign n8974 = n7920 & ~n8973;
  assign n8975 = ~n8877 & ~n8974;
  assign n8976 = ~n7728 & ~n8975;
  assign n8977 = ~n8876 & ~n8976;
  assign n8978 = ~n7723 & ~n8977;
  assign n8979 = ~n7723 & ~n8978;
  assign n8980 = ~n7714 & ~n8979;
  assign n8981 = ~n7714 & ~n8980;
  assign n8982 = n7705 & ~n8981;
  assign n8983 = ~n8358 & ~n8658;
  assign n8984 = ~controllable_hmaster1 & ~n8983;
  assign n8985 = ~n8357 & ~n8984;
  assign n8986 = controllable_hmaster0 & ~n8985;
  assign n8987 = n7928 & ~n8652;
  assign n8988 = ~controllable_hmaster2 & ~n8987;
  assign n8989 = ~n8358 & ~n8988;
  assign n8990 = ~controllable_hmaster1 & ~n8989;
  assign n8991 = ~n8357 & ~n8990;
  assign n8992 = ~controllable_hmaster0 & ~n8991;
  assign n8993 = ~n8986 & ~n8992;
  assign n8994 = controllable_hmaster3 & ~n8993;
  assign n8995 = ~controllable_hmaster3 & ~n8987;
  assign n8996 = ~n8994 & ~n8995;
  assign n8997 = i_hbusreq7 & ~n8996;
  assign n8998 = i_hbusreq8 & ~n8993;
  assign n8999 = i_hbusreq6 & ~n8985;
  assign n9000 = ~n8484 & ~n8711;
  assign n9001 = ~controllable_hmaster1 & ~n9000;
  assign n9002 = ~n8483 & ~n9001;
  assign n9003 = ~i_hbusreq6 & ~n9002;
  assign n9004 = ~n8999 & ~n9003;
  assign n9005 = controllable_hmaster0 & ~n9004;
  assign n9006 = i_hbusreq6 & ~n8991;
  assign n9007 = i_hbusreq5 & ~n8987;
  assign n9008 = i_hbusreq4 & ~n8987;
  assign n9009 = i_hbusreq9 & ~n8987;
  assign n9010 = i_hbusreq3 & ~n8987;
  assign n9011 = i_hbusreq1 & ~n8987;
  assign n9012 = ~n7757 & n7928;
  assign n9013 = n7928 & ~n9012;
  assign n9014 = ~i_hbusreq1 & ~n9013;
  assign n9015 = ~n9011 & ~n9014;
  assign n9016 = ~i_hbusreq3 & ~n9015;
  assign n9017 = ~n9010 & ~n9016;
  assign n9018 = ~i_hbusreq9 & ~n9017;
  assign n9019 = ~n9009 & ~n9018;
  assign n9020 = ~i_hbusreq4 & ~n9019;
  assign n9021 = ~n9008 & ~n9020;
  assign n9022 = ~i_hbusreq5 & ~n9021;
  assign n9023 = ~n9007 & ~n9022;
  assign n9024 = ~controllable_hmaster2 & ~n9023;
  assign n9025 = ~n8484 & ~n9024;
  assign n9026 = ~controllable_hmaster1 & ~n9025;
  assign n9027 = ~n8483 & ~n9026;
  assign n9028 = ~i_hbusreq6 & ~n9027;
  assign n9029 = ~n9006 & ~n9028;
  assign n9030 = ~controllable_hmaster0 & ~n9029;
  assign n9031 = ~n9005 & ~n9030;
  assign n9032 = ~i_hbusreq8 & ~n9031;
  assign n9033 = ~n8998 & ~n9032;
  assign n9034 = controllable_hmaster3 & ~n9033;
  assign n9035 = i_hbusreq8 & ~n8987;
  assign n9036 = i_hbusreq6 & ~n8987;
  assign n9037 = ~i_hbusreq6 & ~n9023;
  assign n9038 = ~n9036 & ~n9037;
  assign n9039 = ~i_hbusreq8 & ~n9038;
  assign n9040 = ~n9035 & ~n9039;
  assign n9041 = ~controllable_hmaster3 & ~n9040;
  assign n9042 = ~n9034 & ~n9041;
  assign n9043 = ~i_hbusreq7 & ~n9042;
  assign n9044 = ~n8997 & ~n9043;
  assign n9045 = ~n8214 & ~n9044;
  assign n9046 = controllable_hmaster0 & ~n8991;
  assign n9047 = ~n8358 & ~n8726;
  assign n9048 = ~controllable_hmaster1 & ~n9047;
  assign n9049 = ~n8357 & ~n9048;
  assign n9050 = ~controllable_hmaster0 & ~n9049;
  assign n9051 = ~n9046 & ~n9050;
  assign n9052 = i_hlock8 & ~n9051;
  assign n9053 = ~n8358 & ~n8733;
  assign n9054 = ~controllable_hmaster1 & ~n9053;
  assign n9055 = ~n8357 & ~n9054;
  assign n9056 = ~controllable_hmaster0 & ~n9055;
  assign n9057 = ~n9046 & ~n9056;
  assign n9058 = ~i_hlock8 & ~n9057;
  assign n9059 = ~n9052 & ~n9058;
  assign n9060 = controllable_hmaster3 & ~n9059;
  assign n9061 = ~n8995 & ~n9060;
  assign n9062 = i_hbusreq7 & ~n9061;
  assign n9063 = i_hbusreq8 & ~n9059;
  assign n9064 = controllable_hmaster0 & ~n9029;
  assign n9065 = i_hbusreq6 & ~n9049;
  assign n9066 = ~n8484 & ~n8755;
  assign n9067 = ~controllable_hmaster1 & ~n9066;
  assign n9068 = ~n8483 & ~n9067;
  assign n9069 = ~i_hbusreq6 & ~n9068;
  assign n9070 = ~n9065 & ~n9069;
  assign n9071 = ~controllable_hmaster0 & ~n9070;
  assign n9072 = ~n9064 & ~n9071;
  assign n9073 = i_hlock8 & ~n9072;
  assign n9074 = i_hbusreq6 & ~n9055;
  assign n9075 = ~n8484 & ~n8774;
  assign n9076 = ~controllable_hmaster1 & ~n9075;
  assign n9077 = ~n8483 & ~n9076;
  assign n9078 = ~i_hbusreq6 & ~n9077;
  assign n9079 = ~n9074 & ~n9078;
  assign n9080 = ~controllable_hmaster0 & ~n9079;
  assign n9081 = ~n9064 & ~n9080;
  assign n9082 = ~i_hlock8 & ~n9081;
  assign n9083 = ~n9073 & ~n9082;
  assign n9084 = ~i_hbusreq8 & ~n9083;
  assign n9085 = ~n9063 & ~n9084;
  assign n9086 = controllable_hmaster3 & ~n9085;
  assign n9087 = ~n9041 & ~n9086;
  assign n9088 = ~i_hbusreq7 & ~n9087;
  assign n9089 = ~n9062 & ~n9088;
  assign n9090 = n8214 & ~n9089;
  assign n9091 = ~n9045 & ~n9090;
  assign n9092 = ~n8202 & ~n9091;
  assign n9093 = controllable_hmaster3 & ~n8991;
  assign n9094 = ~n8793 & ~n8988;
  assign n9095 = controllable_hmaster1 & ~n9094;
  assign n9096 = ~controllable_hmaster1 & ~n8987;
  assign n9097 = ~n9095 & ~n9096;
  assign n9098 = controllable_hmaster0 & ~n9097;
  assign n9099 = ~controllable_hmaster0 & ~n8987;
  assign n9100 = ~n9098 & ~n9099;
  assign n9101 = ~controllable_hmaster3 & ~n9100;
  assign n9102 = ~n9093 & ~n9101;
  assign n9103 = i_hlock7 & ~n9102;
  assign n9104 = ~n8802 & ~n8988;
  assign n9105 = controllable_hmaster1 & ~n9104;
  assign n9106 = ~n9096 & ~n9105;
  assign n9107 = controllable_hmaster0 & ~n9106;
  assign n9108 = ~n9099 & ~n9107;
  assign n9109 = ~controllable_hmaster3 & ~n9108;
  assign n9110 = ~n9093 & ~n9109;
  assign n9111 = ~i_hlock7 & ~n9110;
  assign n9112 = ~n9103 & ~n9111;
  assign n9113 = i_hbusreq7 & ~n9112;
  assign n9114 = i_hbusreq8 & ~n8991;
  assign n9115 = ~i_hbusreq8 & ~n9029;
  assign n9116 = ~n9114 & ~n9115;
  assign n9117 = controllable_hmaster3 & ~n9116;
  assign n9118 = i_hbusreq8 & ~n9100;
  assign n9119 = i_hbusreq6 & ~n9097;
  assign n9120 = ~n8815 & ~n9024;
  assign n9121 = controllable_hmaster1 & ~n9120;
  assign n9122 = ~controllable_hmaster1 & ~n9023;
  assign n9123 = ~n9121 & ~n9122;
  assign n9124 = ~i_hbusreq6 & ~n9123;
  assign n9125 = ~n9119 & ~n9124;
  assign n9126 = controllable_hmaster0 & ~n9125;
  assign n9127 = ~controllable_hmaster0 & ~n9038;
  assign n9128 = ~n9126 & ~n9127;
  assign n9129 = ~i_hbusreq8 & ~n9128;
  assign n9130 = ~n9118 & ~n9129;
  assign n9131 = ~controllable_hmaster3 & ~n9130;
  assign n9132 = ~n9117 & ~n9131;
  assign n9133 = i_hlock7 & ~n9132;
  assign n9134 = i_hbusreq8 & ~n9108;
  assign n9135 = i_hbusreq6 & ~n9106;
  assign n9136 = ~n8830 & ~n9024;
  assign n9137 = controllable_hmaster1 & ~n9136;
  assign n9138 = ~n9122 & ~n9137;
  assign n9139 = ~i_hbusreq6 & ~n9138;
  assign n9140 = ~n9135 & ~n9139;
  assign n9141 = controllable_hmaster0 & ~n9140;
  assign n9142 = ~n9127 & ~n9141;
  assign n9143 = ~i_hbusreq8 & ~n9142;
  assign n9144 = ~n9134 & ~n9143;
  assign n9145 = ~controllable_hmaster3 & ~n9144;
  assign n9146 = ~n9117 & ~n9145;
  assign n9147 = ~i_hlock7 & ~n9146;
  assign n9148 = ~n9133 & ~n9147;
  assign n9149 = ~i_hbusreq7 & ~n9148;
  assign n9150 = ~n9113 & ~n9149;
  assign n9151 = ~n8214 & ~n9150;
  assign n9152 = controllable_hmaster0 & ~n8987;
  assign n9153 = i_hlock6 & ~n9097;
  assign n9154 = ~i_hlock6 & ~n9106;
  assign n9155 = ~n9153 & ~n9154;
  assign n9156 = ~controllable_hmaster0 & ~n9155;
  assign n9157 = ~n9152 & ~n9156;
  assign n9158 = ~controllable_hmaster3 & ~n9157;
  assign n9159 = ~n9093 & ~n9158;
  assign n9160 = i_hbusreq7 & ~n9159;
  assign n9161 = i_hbusreq8 & ~n9157;
  assign n9162 = controllable_hmaster0 & ~n9038;
  assign n9163 = i_hbusreq6 & ~n9155;
  assign n9164 = i_hlock6 & ~n9123;
  assign n9165 = ~i_hlock6 & ~n9138;
  assign n9166 = ~n9164 & ~n9165;
  assign n9167 = ~i_hbusreq6 & ~n9166;
  assign n9168 = ~n9163 & ~n9167;
  assign n9169 = ~controllable_hmaster0 & ~n9168;
  assign n9170 = ~n9162 & ~n9169;
  assign n9171 = ~i_hbusreq8 & ~n9170;
  assign n9172 = ~n9161 & ~n9171;
  assign n9173 = ~controllable_hmaster3 & ~n9172;
  assign n9174 = ~n9117 & ~n9173;
  assign n9175 = ~i_hbusreq7 & ~n9174;
  assign n9176 = ~n9160 & ~n9175;
  assign n9177 = n8214 & ~n9176;
  assign n9178 = ~n9151 & ~n9177;
  assign n9179 = n8202 & ~n9178;
  assign n9180 = ~n9092 & ~n9179;
  assign n9181 = n7920 & ~n9180;
  assign n9182 = ~n8877 & ~n9181;
  assign n9183 = n7728 & ~n9182;
  assign n9184 = ~n8986 & ~n9050;
  assign n9185 = i_hlock8 & ~n9184;
  assign n9186 = ~n8986 & ~n9056;
  assign n9187 = ~i_hlock8 & ~n9186;
  assign n9188 = ~n9185 & ~n9187;
  assign n9189 = controllable_hmaster3 & ~n9188;
  assign n9190 = i_hlock3 & ~n8653;
  assign n9191 = ~i_hlock3 & ~n8655;
  assign n9192 = ~n9190 & ~n9191;
  assign n9193 = ~controllable_hmaster2 & ~n9192;
  assign n9194 = ~n8793 & ~n9193;
  assign n9195 = controllable_hmaster1 & ~n9194;
  assign n9196 = i_hlock5 & ~n8653;
  assign n9197 = ~i_hlock5 & ~n8655;
  assign n9198 = ~n9196 & ~n9197;
  assign n9199 = controllable_hmaster2 & ~n9198;
  assign n9200 = i_hlock1 & ~n8653;
  assign n9201 = ~i_hlock1 & ~n8655;
  assign n9202 = ~n9200 & ~n9201;
  assign n9203 = ~controllable_hmaster2 & ~n9202;
  assign n9204 = ~n9199 & ~n9203;
  assign n9205 = ~controllable_hmaster1 & ~n9204;
  assign n9206 = ~n9195 & ~n9205;
  assign n9207 = controllable_hmaster0 & ~n9206;
  assign n9208 = i_hlock2 & ~n8218;
  assign n9209 = ~i_hlock2 & ~n8232;
  assign n9210 = ~n9208 & ~n9209;
  assign n9211 = ~n7733 & ~n9210;
  assign n9212 = ~n7733 & ~n9211;
  assign n9213 = ~n7928 & ~n9212;
  assign n9214 = ~n8652 & ~n9213;
  assign n9215 = ~controllable_hmaster2 & ~n9214;
  assign n9216 = ~n8793 & ~n9215;
  assign n9217 = controllable_hmaster1 & ~n9216;
  assign n9218 = i_hlock4 & ~n8653;
  assign n9219 = ~i_hlock4 & ~n8655;
  assign n9220 = ~n9218 & ~n9219;
  assign n9221 = controllable_hmaster2 & ~n9220;
  assign n9222 = ~n8440 & ~n8652;
  assign n9223 = ~controllable_hmaster2 & ~n9222;
  assign n9224 = ~n9221 & ~n9223;
  assign n9225 = ~controllable_hmaster1 & ~n9224;
  assign n9226 = ~n9217 & ~n9225;
  assign n9227 = i_hlock6 & ~n9226;
  assign n9228 = ~n8802 & ~n9215;
  assign n9229 = controllable_hmaster1 & ~n9228;
  assign n9230 = ~n9225 & ~n9229;
  assign n9231 = ~i_hlock6 & ~n9230;
  assign n9232 = ~n9227 & ~n9231;
  assign n9233 = ~controllable_hmaster0 & ~n9232;
  assign n9234 = ~n9207 & ~n9233;
  assign n9235 = ~controllable_hmaster3 & ~n9234;
  assign n9236 = ~n9189 & ~n9235;
  assign n9237 = i_hlock7 & ~n9236;
  assign n9238 = ~n8802 & ~n9193;
  assign n9239 = controllable_hmaster1 & ~n9238;
  assign n9240 = ~n9205 & ~n9239;
  assign n9241 = controllable_hmaster0 & ~n9240;
  assign n9242 = ~n9233 & ~n9241;
  assign n9243 = ~controllable_hmaster3 & ~n9242;
  assign n9244 = ~n9189 & ~n9243;
  assign n9245 = ~i_hlock7 & ~n9244;
  assign n9246 = ~n9237 & ~n9245;
  assign n9247 = i_hbusreq7 & ~n9246;
  assign n9248 = i_hbusreq8 & ~n9188;
  assign n9249 = ~i_hbusreq1 & ~n8679;
  assign n9250 = ~n8472 & ~n9249;
  assign n9251 = ~i_hbusreq3 & ~n9250;
  assign n9252 = ~n8471 & ~n9251;
  assign n9253 = ~i_hbusreq9 & ~n9252;
  assign n9254 = ~n8470 & ~n9253;
  assign n9255 = ~i_hbusreq4 & ~n9254;
  assign n9256 = ~n8469 & ~n9255;
  assign n9257 = ~i_hbusreq5 & ~n9256;
  assign n9258 = ~n8468 & ~n9257;
  assign n9259 = controllable_hmaster1 & ~n9258;
  assign n9260 = controllable_hmaster2 & ~n9258;
  assign n9261 = ~n8711 & ~n9260;
  assign n9262 = ~controllable_hmaster1 & ~n9261;
  assign n9263 = ~n9259 & ~n9262;
  assign n9264 = ~i_hbusreq6 & ~n9263;
  assign n9265 = ~n8999 & ~n9264;
  assign n9266 = controllable_hmaster0 & ~n9265;
  assign n9267 = n7928 & ~n8679;
  assign n9268 = ~n8265 & ~n9267;
  assign n9269 = ~i_hbusreq1 & ~n9268;
  assign n9270 = ~n8673 & ~n9269;
  assign n9271 = ~i_hbusreq3 & ~n9270;
  assign n9272 = ~n8672 & ~n9271;
  assign n9273 = ~i_hbusreq9 & ~n9272;
  assign n9274 = ~n8748 & ~n9273;
  assign n9275 = ~i_hbusreq4 & ~n9274;
  assign n9276 = ~n8747 & ~n9275;
  assign n9277 = ~i_hbusreq5 & ~n9276;
  assign n9278 = ~n8746 & ~n9277;
  assign n9279 = ~controllable_hmaster2 & ~n9278;
  assign n9280 = ~n9260 & ~n9279;
  assign n9281 = ~controllable_hmaster1 & ~n9280;
  assign n9282 = ~n9259 & ~n9281;
  assign n9283 = ~i_hbusreq6 & ~n9282;
  assign n9284 = ~n9065 & ~n9283;
  assign n9285 = ~controllable_hmaster0 & ~n9284;
  assign n9286 = ~n9266 & ~n9285;
  assign n9287 = i_hlock8 & ~n9286;
  assign n9288 = ~n8297 & ~n9267;
  assign n9289 = ~i_hbusreq1 & ~n9288;
  assign n9290 = ~n8697 & ~n9289;
  assign n9291 = ~i_hbusreq3 & ~n9290;
  assign n9292 = ~n8696 & ~n9291;
  assign n9293 = ~i_hbusreq9 & ~n9292;
  assign n9294 = ~n8767 & ~n9293;
  assign n9295 = ~i_hbusreq4 & ~n9294;
  assign n9296 = ~n8766 & ~n9295;
  assign n9297 = ~i_hbusreq5 & ~n9296;
  assign n9298 = ~n8765 & ~n9297;
  assign n9299 = ~controllable_hmaster2 & ~n9298;
  assign n9300 = ~n9260 & ~n9299;
  assign n9301 = ~controllable_hmaster1 & ~n9300;
  assign n9302 = ~n9259 & ~n9301;
  assign n9303 = ~i_hbusreq6 & ~n9302;
  assign n9304 = ~n9074 & ~n9303;
  assign n9305 = ~controllable_hmaster0 & ~n9304;
  assign n9306 = ~n9266 & ~n9305;
  assign n9307 = ~i_hlock8 & ~n9306;
  assign n9308 = ~n9287 & ~n9307;
  assign n9309 = ~i_hbusreq8 & ~n9308;
  assign n9310 = ~n9248 & ~n9309;
  assign n9311 = controllable_hmaster3 & ~n9310;
  assign n9312 = i_hbusreq8 & ~n9234;
  assign n9313 = i_hbusreq6 & ~n9206;
  assign n9314 = controllable_hmaster2 & ~n9278;
  assign n9315 = i_hbusreq5 & ~n9192;
  assign n9316 = i_hbusreq4 & ~n9192;
  assign n9317 = i_hbusreq9 & ~n9192;
  assign n9318 = i_hbusreq3 & ~n9192;
  assign n9319 = i_hlock3 & ~n9270;
  assign n9320 = ~i_hlock3 & ~n9290;
  assign n9321 = ~n9319 & ~n9320;
  assign n9322 = ~i_hbusreq3 & ~n9321;
  assign n9323 = ~n9318 & ~n9322;
  assign n9324 = ~i_hbusreq9 & ~n9323;
  assign n9325 = ~n9317 & ~n9324;
  assign n9326 = ~i_hbusreq4 & ~n9325;
  assign n9327 = ~n9316 & ~n9326;
  assign n9328 = ~i_hbusreq5 & ~n9327;
  assign n9329 = ~n9315 & ~n9328;
  assign n9330 = ~controllable_hmaster2 & ~n9329;
  assign n9331 = ~n9314 & ~n9330;
  assign n9332 = controllable_hmaster1 & ~n9331;
  assign n9333 = i_hbusreq5 & ~n9198;
  assign n9334 = i_hlock5 & ~n9276;
  assign n9335 = ~i_hlock5 & ~n9296;
  assign n9336 = ~n9334 & ~n9335;
  assign n9337 = ~i_hbusreq5 & ~n9336;
  assign n9338 = ~n9333 & ~n9337;
  assign n9339 = controllable_hmaster2 & ~n9338;
  assign n9340 = i_hbusreq5 & ~n9202;
  assign n9341 = i_hbusreq4 & ~n9202;
  assign n9342 = i_hbusreq9 & ~n9202;
  assign n9343 = i_hbusreq3 & ~n9202;
  assign n9344 = i_hbusreq1 & ~n9202;
  assign n9345 = i_hlock1 & ~n9268;
  assign n9346 = ~i_hlock1 & ~n9288;
  assign n9347 = ~n9345 & ~n9346;
  assign n9348 = ~i_hbusreq1 & ~n9347;
  assign n9349 = ~n9344 & ~n9348;
  assign n9350 = ~i_hbusreq3 & ~n9349;
  assign n9351 = ~n9343 & ~n9350;
  assign n9352 = ~i_hbusreq9 & ~n9351;
  assign n9353 = ~n9342 & ~n9352;
  assign n9354 = ~i_hbusreq4 & ~n9353;
  assign n9355 = ~n9341 & ~n9354;
  assign n9356 = ~i_hbusreq5 & ~n9355;
  assign n9357 = ~n9340 & ~n9356;
  assign n9358 = ~controllable_hmaster2 & ~n9357;
  assign n9359 = ~n9339 & ~n9358;
  assign n9360 = ~controllable_hmaster1 & ~n9359;
  assign n9361 = ~n9332 & ~n9360;
  assign n9362 = ~i_hbusreq6 & ~n9361;
  assign n9363 = ~n9313 & ~n9362;
  assign n9364 = controllable_hmaster0 & ~n9363;
  assign n9365 = i_hbusreq6 & ~n9232;
  assign n9366 = i_hbusreq5 & ~n9214;
  assign n9367 = i_hbusreq4 & ~n9214;
  assign n9368 = i_hbusreq9 & ~n9214;
  assign n9369 = i_hbusreq3 & ~n9214;
  assign n9370 = i_hbusreq1 & ~n9214;
  assign n9371 = i_hbusreq2 & ~n9210;
  assign n9372 = i_hlock2 & ~n8260;
  assign n9373 = ~i_hlock2 & ~n8292;
  assign n9374 = ~n9372 & ~n9373;
  assign n9375 = ~i_hbusreq2 & ~n9374;
  assign n9376 = ~n9371 & ~n9375;
  assign n9377 = ~n7733 & ~n9376;
  assign n9378 = ~n7733 & ~n9377;
  assign n9379 = ~n7928 & ~n9378;
  assign n9380 = ~n9267 & ~n9379;
  assign n9381 = ~i_hbusreq1 & ~n9380;
  assign n9382 = ~n9370 & ~n9381;
  assign n9383 = ~i_hbusreq3 & ~n9382;
  assign n9384 = ~n9369 & ~n9383;
  assign n9385 = ~i_hbusreq9 & ~n9384;
  assign n9386 = ~n9368 & ~n9385;
  assign n9387 = ~i_hbusreq4 & ~n9386;
  assign n9388 = ~n9367 & ~n9387;
  assign n9389 = ~i_hbusreq5 & ~n9388;
  assign n9390 = ~n9366 & ~n9389;
  assign n9391 = ~controllable_hmaster2 & ~n9390;
  assign n9392 = ~n9314 & ~n9391;
  assign n9393 = controllable_hmaster1 & ~n9392;
  assign n9394 = i_hbusreq5 & ~n9220;
  assign n9395 = i_hbusreq4 & ~n9220;
  assign n9396 = i_hlock4 & ~n9274;
  assign n9397 = ~i_hlock4 & ~n9294;
  assign n9398 = ~n9396 & ~n9397;
  assign n9399 = ~i_hbusreq4 & ~n9398;
  assign n9400 = ~n9395 & ~n9399;
  assign n9401 = ~i_hbusreq5 & ~n9400;
  assign n9402 = ~n9394 & ~n9401;
  assign n9403 = controllable_hmaster2 & ~n9402;
  assign n9404 = i_hbusreq5 & ~n9222;
  assign n9405 = i_hbusreq4 & ~n9222;
  assign n9406 = i_hbusreq9 & ~n9222;
  assign n9407 = i_hbusreq3 & ~n9222;
  assign n9408 = i_hbusreq1 & ~n9222;
  assign n9409 = ~n8435 & ~n8674;
  assign n9410 = ~i_hbusreq0 & ~n9409;
  assign n9411 = ~n7754 & ~n9410;
  assign n9412 = ~i_hbusreq2 & ~n9411;
  assign n9413 = ~n7753 & ~n9412;
  assign n9414 = n7928 & ~n9413;
  assign n9415 = ~n8440 & ~n9414;
  assign n9416 = ~i_hbusreq1 & ~n9415;
  assign n9417 = ~n9408 & ~n9416;
  assign n9418 = ~i_hbusreq3 & ~n9417;
  assign n9419 = ~n9407 & ~n9418;
  assign n9420 = ~i_hbusreq9 & ~n9419;
  assign n9421 = ~n9406 & ~n9420;
  assign n9422 = ~i_hbusreq4 & ~n9421;
  assign n9423 = ~n9405 & ~n9422;
  assign n9424 = ~i_hbusreq5 & ~n9423;
  assign n9425 = ~n9404 & ~n9424;
  assign n9426 = ~controllable_hmaster2 & ~n9425;
  assign n9427 = ~n9403 & ~n9426;
  assign n9428 = ~controllable_hmaster1 & ~n9427;
  assign n9429 = ~n9393 & ~n9428;
  assign n9430 = i_hlock6 & ~n9429;
  assign n9431 = controllable_hmaster2 & ~n9298;
  assign n9432 = ~n9391 & ~n9431;
  assign n9433 = controllable_hmaster1 & ~n9432;
  assign n9434 = ~n9428 & ~n9433;
  assign n9435 = ~i_hlock6 & ~n9434;
  assign n9436 = ~n9430 & ~n9435;
  assign n9437 = ~i_hbusreq6 & ~n9436;
  assign n9438 = ~n9365 & ~n9437;
  assign n9439 = ~controllable_hmaster0 & ~n9438;
  assign n9440 = ~n9364 & ~n9439;
  assign n9441 = ~i_hbusreq8 & ~n9440;
  assign n9442 = ~n9312 & ~n9441;
  assign n9443 = ~controllable_hmaster3 & ~n9442;
  assign n9444 = ~n9311 & ~n9443;
  assign n9445 = i_hlock7 & ~n9444;
  assign n9446 = i_hbusreq8 & ~n9242;
  assign n9447 = i_hbusreq6 & ~n9240;
  assign n9448 = ~n9330 & ~n9431;
  assign n9449 = controllable_hmaster1 & ~n9448;
  assign n9450 = ~n9360 & ~n9449;
  assign n9451 = ~i_hbusreq6 & ~n9450;
  assign n9452 = ~n9447 & ~n9451;
  assign n9453 = controllable_hmaster0 & ~n9452;
  assign n9454 = ~n9439 & ~n9453;
  assign n9455 = ~i_hbusreq8 & ~n9454;
  assign n9456 = ~n9446 & ~n9455;
  assign n9457 = ~controllable_hmaster3 & ~n9456;
  assign n9458 = ~n9311 & ~n9457;
  assign n9459 = ~i_hlock7 & ~n9458;
  assign n9460 = ~n9445 & ~n9459;
  assign n9461 = ~i_hbusreq7 & ~n9460;
  assign n9462 = ~n9247 & ~n9461;
  assign n9463 = ~n8214 & ~n9462;
  assign n9464 = i_hlock9 & ~n9272;
  assign n9465 = ~i_hlock9 & ~n9292;
  assign n9466 = ~n9464 & ~n9465;
  assign n9467 = ~i_hbusreq9 & ~n9466;
  assign n9468 = ~n8671 & ~n9467;
  assign n9469 = ~i_hbusreq4 & ~n9468;
  assign n9470 = ~n8670 & ~n9469;
  assign n9471 = ~i_hbusreq5 & ~n9470;
  assign n9472 = ~n8669 & ~n9471;
  assign n9473 = ~controllable_hmaster2 & ~n9472;
  assign n9474 = ~n9260 & ~n9473;
  assign n9475 = ~controllable_hmaster1 & ~n9474;
  assign n9476 = ~n9259 & ~n9475;
  assign n9477 = ~i_hbusreq6 & ~n9476;
  assign n9478 = ~n8999 & ~n9477;
  assign n9479 = controllable_hmaster0 & ~n9478;
  assign n9480 = ~n8755 & ~n9260;
  assign n9481 = ~controllable_hmaster1 & ~n9480;
  assign n9482 = ~n9259 & ~n9481;
  assign n9483 = ~i_hbusreq6 & ~n9482;
  assign n9484 = ~n9065 & ~n9483;
  assign n9485 = ~controllable_hmaster0 & ~n9484;
  assign n9486 = ~n9479 & ~n9485;
  assign n9487 = i_hlock8 & ~n9486;
  assign n9488 = ~n8774 & ~n9260;
  assign n9489 = ~controllable_hmaster1 & ~n9488;
  assign n9490 = ~n9259 & ~n9489;
  assign n9491 = ~i_hbusreq6 & ~n9490;
  assign n9492 = ~n9074 & ~n9491;
  assign n9493 = ~controllable_hmaster0 & ~n9492;
  assign n9494 = ~n9479 & ~n9493;
  assign n9495 = ~i_hlock8 & ~n9494;
  assign n9496 = ~n9487 & ~n9495;
  assign n9497 = ~i_hbusreq8 & ~n9496;
  assign n9498 = ~n9248 & ~n9497;
  assign n9499 = controllable_hmaster3 & ~n9498;
  assign n9500 = ~n9443 & ~n9499;
  assign n9501 = i_hlock7 & ~n9500;
  assign n9502 = ~n9457 & ~n9499;
  assign n9503 = ~i_hlock7 & ~n9502;
  assign n9504 = ~n9501 & ~n9503;
  assign n9505 = ~i_hbusreq7 & ~n9504;
  assign n9506 = ~n9247 & ~n9505;
  assign n9507 = n8214 & ~n9506;
  assign n9508 = ~n9463 & ~n9507;
  assign n9509 = ~n8202 & ~n9508;
  assign n9510 = ~n9285 & ~n9479;
  assign n9511 = i_hlock8 & ~n9510;
  assign n9512 = ~n9305 & ~n9479;
  assign n9513 = ~i_hlock8 & ~n9512;
  assign n9514 = ~n9511 & ~n9513;
  assign n9515 = ~i_hbusreq8 & ~n9514;
  assign n9516 = ~n9248 & ~n9515;
  assign n9517 = controllable_hmaster3 & ~n9516;
  assign n9518 = ~n8815 & ~n9330;
  assign n9519 = controllable_hmaster1 & ~n9518;
  assign n9520 = ~n9360 & ~n9519;
  assign n9521 = ~i_hbusreq6 & ~n9520;
  assign n9522 = ~n9313 & ~n9521;
  assign n9523 = controllable_hmaster0 & ~n9522;
  assign n9524 = ~n9439 & ~n9523;
  assign n9525 = ~i_hbusreq8 & ~n9524;
  assign n9526 = ~n9312 & ~n9525;
  assign n9527 = ~controllable_hmaster3 & ~n9526;
  assign n9528 = ~n9517 & ~n9527;
  assign n9529 = i_hlock7 & ~n9528;
  assign n9530 = ~n8830 & ~n9330;
  assign n9531 = controllable_hmaster1 & ~n9530;
  assign n9532 = ~n9360 & ~n9531;
  assign n9533 = ~i_hbusreq6 & ~n9532;
  assign n9534 = ~n9447 & ~n9533;
  assign n9535 = controllable_hmaster0 & ~n9534;
  assign n9536 = ~n9439 & ~n9535;
  assign n9537 = ~i_hbusreq8 & ~n9536;
  assign n9538 = ~n9446 & ~n9537;
  assign n9539 = ~controllable_hmaster3 & ~n9538;
  assign n9540 = ~n9517 & ~n9539;
  assign n9541 = ~i_hlock7 & ~n9540;
  assign n9542 = ~n9529 & ~n9541;
  assign n9543 = ~i_hbusreq7 & ~n9542;
  assign n9544 = ~n9247 & ~n9543;
  assign n9545 = ~n8214 & ~n9544;
  assign n9546 = ~n8815 & ~n9391;
  assign n9547 = controllable_hmaster1 & ~n9546;
  assign n9548 = ~n9428 & ~n9547;
  assign n9549 = i_hlock6 & ~n9548;
  assign n9550 = ~n8830 & ~n9391;
  assign n9551 = controllable_hmaster1 & ~n9550;
  assign n9552 = ~n9428 & ~n9551;
  assign n9553 = ~i_hlock6 & ~n9552;
  assign n9554 = ~n9549 & ~n9553;
  assign n9555 = ~i_hbusreq6 & ~n9554;
  assign n9556 = ~n9365 & ~n9555;
  assign n9557 = ~controllable_hmaster0 & ~n9556;
  assign n9558 = ~n9364 & ~n9557;
  assign n9559 = ~i_hbusreq8 & ~n9558;
  assign n9560 = ~n9312 & ~n9559;
  assign n9561 = ~controllable_hmaster3 & ~n9560;
  assign n9562 = ~n9517 & ~n9561;
  assign n9563 = i_hlock7 & ~n9562;
  assign n9564 = ~n9453 & ~n9557;
  assign n9565 = ~i_hbusreq8 & ~n9564;
  assign n9566 = ~n9446 & ~n9565;
  assign n9567 = ~controllable_hmaster3 & ~n9566;
  assign n9568 = ~n9517 & ~n9567;
  assign n9569 = ~i_hlock7 & ~n9568;
  assign n9570 = ~n9563 & ~n9569;
  assign n9571 = ~i_hbusreq7 & ~n9570;
  assign n9572 = ~n9247 & ~n9571;
  assign n9573 = n8214 & ~n9572;
  assign n9574 = ~n9545 & ~n9573;
  assign n9575 = n8202 & ~n9574;
  assign n9576 = ~n9509 & ~n9575;
  assign n9577 = n7920 & ~n9576;
  assign n9578 = ~n8877 & ~n9577;
  assign n9579 = ~n7728 & ~n9578;
  assign n9580 = ~n9183 & ~n9579;
  assign n9581 = n7723 & ~n9580;
  assign n9582 = ~n7723 & ~n9578;
  assign n9583 = ~n9581 & ~n9582;
  assign n9584 = n7714 & ~n9583;
  assign n9585 = n7723 & ~n9578;
  assign n9586 = ~n8640 & ~n9577;
  assign n9587 = n7728 & ~n9586;
  assign n9588 = ~n7736 & ~n8687;
  assign n9589 = ~i_hbusreq1 & ~n9588;
  assign n9590 = ~n8472 & ~n9589;
  assign n9591 = ~i_hbusreq3 & ~n9590;
  assign n9592 = ~n8471 & ~n9591;
  assign n9593 = ~i_hbusreq9 & ~n9592;
  assign n9594 = ~n8470 & ~n9593;
  assign n9595 = ~i_hbusreq4 & ~n9594;
  assign n9596 = ~n8469 & ~n9595;
  assign n9597 = ~i_hbusreq5 & ~n9596;
  assign n9598 = ~n8468 & ~n9597;
  assign n9599 = controllable_hmaster1 & ~n9598;
  assign n9600 = controllable_hmaster2 & ~n9598;
  assign n9601 = ~n8711 & ~n9600;
  assign n9602 = ~controllable_hmaster1 & ~n9601;
  assign n9603 = ~n9599 & ~n9602;
  assign n9604 = ~i_hbusreq6 & ~n9603;
  assign n9605 = ~n8999 & ~n9604;
  assign n9606 = controllable_hmaster0 & ~n9605;
  assign n9607 = ~n8755 & ~n9600;
  assign n9608 = ~controllable_hmaster1 & ~n9607;
  assign n9609 = ~n9599 & ~n9608;
  assign n9610 = ~i_hbusreq6 & ~n9609;
  assign n9611 = ~n9065 & ~n9610;
  assign n9612 = ~controllable_hmaster0 & ~n9611;
  assign n9613 = ~n9606 & ~n9612;
  assign n9614 = i_hlock8 & ~n9613;
  assign n9615 = ~n8774 & ~n9600;
  assign n9616 = ~controllable_hmaster1 & ~n9615;
  assign n9617 = ~n9599 & ~n9616;
  assign n9618 = ~i_hbusreq6 & ~n9617;
  assign n9619 = ~n9074 & ~n9618;
  assign n9620 = ~controllable_hmaster0 & ~n9619;
  assign n9621 = ~n9606 & ~n9620;
  assign n9622 = ~i_hlock8 & ~n9621;
  assign n9623 = ~n9614 & ~n9622;
  assign n9624 = ~i_hbusreq8 & ~n9623;
  assign n9625 = ~n9248 & ~n9624;
  assign n9626 = controllable_hmaster3 & ~n9625;
  assign n9627 = i_hlock3 & ~n8692;
  assign n9628 = ~i_hlock3 & ~n8700;
  assign n9629 = ~n9627 & ~n9628;
  assign n9630 = ~i_hbusreq3 & ~n9629;
  assign n9631 = ~n9318 & ~n9630;
  assign n9632 = ~i_hbusreq9 & ~n9631;
  assign n9633 = ~n9317 & ~n9632;
  assign n9634 = ~i_hbusreq4 & ~n9633;
  assign n9635 = ~n9316 & ~n9634;
  assign n9636 = ~i_hbusreq5 & ~n9635;
  assign n9637 = ~n9315 & ~n9636;
  assign n9638 = ~controllable_hmaster2 & ~n9637;
  assign n9639 = ~n8815 & ~n9638;
  assign n9640 = controllable_hmaster1 & ~n9639;
  assign n9641 = i_hlock5 & ~n8752;
  assign n9642 = ~i_hlock5 & ~n8771;
  assign n9643 = ~n9641 & ~n9642;
  assign n9644 = ~i_hbusreq5 & ~n9643;
  assign n9645 = ~n9333 & ~n9644;
  assign n9646 = controllable_hmaster2 & ~n9645;
  assign n9647 = i_hlock1 & ~n8690;
  assign n9648 = ~i_hlock1 & ~n8698;
  assign n9649 = ~n9647 & ~n9648;
  assign n9650 = ~i_hbusreq1 & ~n9649;
  assign n9651 = ~n9344 & ~n9650;
  assign n9652 = ~i_hbusreq3 & ~n9651;
  assign n9653 = ~n9343 & ~n9652;
  assign n9654 = ~i_hbusreq9 & ~n9653;
  assign n9655 = ~n9342 & ~n9654;
  assign n9656 = ~i_hbusreq4 & ~n9655;
  assign n9657 = ~n9341 & ~n9656;
  assign n9658 = ~i_hbusreq5 & ~n9657;
  assign n9659 = ~n9340 & ~n9658;
  assign n9660 = ~controllable_hmaster2 & ~n9659;
  assign n9661 = ~n9646 & ~n9660;
  assign n9662 = ~controllable_hmaster1 & ~n9661;
  assign n9663 = ~n9640 & ~n9662;
  assign n9664 = ~i_hbusreq6 & ~n9663;
  assign n9665 = ~n9313 & ~n9664;
  assign n9666 = controllable_hmaster0 & ~n9665;
  assign n9667 = ~n8689 & ~n9379;
  assign n9668 = ~i_hbusreq1 & ~n9667;
  assign n9669 = ~n9370 & ~n9668;
  assign n9670 = ~i_hbusreq3 & ~n9669;
  assign n9671 = ~n9369 & ~n9670;
  assign n9672 = ~i_hbusreq9 & ~n9671;
  assign n9673 = ~n9368 & ~n9672;
  assign n9674 = ~i_hbusreq4 & ~n9673;
  assign n9675 = ~n9367 & ~n9674;
  assign n9676 = ~i_hbusreq5 & ~n9675;
  assign n9677 = ~n9366 & ~n9676;
  assign n9678 = ~controllable_hmaster2 & ~n9677;
  assign n9679 = ~n8815 & ~n9678;
  assign n9680 = controllable_hmaster1 & ~n9679;
  assign n9681 = i_hlock4 & ~n8750;
  assign n9682 = ~i_hlock4 & ~n8769;
  assign n9683 = ~n9681 & ~n9682;
  assign n9684 = ~i_hbusreq4 & ~n9683;
  assign n9685 = ~n9395 & ~n9684;
  assign n9686 = ~i_hbusreq5 & ~n9685;
  assign n9687 = ~n9394 & ~n9686;
  assign n9688 = controllable_hmaster2 & ~n9687;
  assign n9689 = ~n7733 & ~n9413;
  assign n9690 = n7733 & ~n7735;
  assign n9691 = ~n9689 & ~n9690;
  assign n9692 = n7928 & ~n9691;
  assign n9693 = ~n8440 & ~n9692;
  assign n9694 = ~i_hbusreq1 & ~n9693;
  assign n9695 = ~n9408 & ~n9694;
  assign n9696 = ~i_hbusreq3 & ~n9695;
  assign n9697 = ~n9407 & ~n9696;
  assign n9698 = ~i_hbusreq9 & ~n9697;
  assign n9699 = ~n9406 & ~n9698;
  assign n9700 = ~i_hbusreq4 & ~n9699;
  assign n9701 = ~n9405 & ~n9700;
  assign n9702 = ~i_hbusreq5 & ~n9701;
  assign n9703 = ~n9404 & ~n9702;
  assign n9704 = ~controllable_hmaster2 & ~n9703;
  assign n9705 = ~n9688 & ~n9704;
  assign n9706 = ~controllable_hmaster1 & ~n9705;
  assign n9707 = ~n9680 & ~n9706;
  assign n9708 = i_hlock6 & ~n9707;
  assign n9709 = ~n8830 & ~n9678;
  assign n9710 = controllable_hmaster1 & ~n9709;
  assign n9711 = ~n9706 & ~n9710;
  assign n9712 = ~i_hlock6 & ~n9711;
  assign n9713 = ~n9708 & ~n9712;
  assign n9714 = ~i_hbusreq6 & ~n9713;
  assign n9715 = ~n9365 & ~n9714;
  assign n9716 = ~controllable_hmaster0 & ~n9715;
  assign n9717 = ~n9666 & ~n9716;
  assign n9718 = ~i_hbusreq8 & ~n9717;
  assign n9719 = ~n9312 & ~n9718;
  assign n9720 = ~controllable_hmaster3 & ~n9719;
  assign n9721 = ~n9626 & ~n9720;
  assign n9722 = i_hlock7 & ~n9721;
  assign n9723 = ~n8830 & ~n9638;
  assign n9724 = controllable_hmaster1 & ~n9723;
  assign n9725 = ~n9662 & ~n9724;
  assign n9726 = ~i_hbusreq6 & ~n9725;
  assign n9727 = ~n9447 & ~n9726;
  assign n9728 = controllable_hmaster0 & ~n9727;
  assign n9729 = ~n9716 & ~n9728;
  assign n9730 = ~i_hbusreq8 & ~n9729;
  assign n9731 = ~n9446 & ~n9730;
  assign n9732 = ~controllable_hmaster3 & ~n9731;
  assign n9733 = ~n9626 & ~n9732;
  assign n9734 = ~i_hlock7 & ~n9733;
  assign n9735 = ~n9722 & ~n9734;
  assign n9736 = ~i_hbusreq7 & ~n9735;
  assign n9737 = ~n9247 & ~n9736;
  assign n9738 = n7920 & ~n9737;
  assign n9739 = ~n8640 & ~n9738;
  assign n9740 = ~n7728 & ~n9739;
  assign n9741 = ~n9587 & ~n9740;
  assign n9742 = ~n7723 & ~n9741;
  assign n9743 = ~n9585 & ~n9742;
  assign n9744 = ~n7714 & ~n9743;
  assign n9745 = ~n9584 & ~n9744;
  assign n9746 = ~n7705 & ~n9745;
  assign n9747 = ~n8982 & ~n9746;
  assign n9748 = n7808 & ~n9747;
  assign n9749 = ~n8650 & ~n9748;
  assign n9750 = n8195 & ~n9749;
  assign n9751 = ~n8196 & ~n9750;
  assign n9752 = ~n8193 & ~n9751;
  assign n9753 = controllable_hmaster2 & ~n8386;
  assign n9754 = ~controllable_hmaster1 & ~n9753;
  assign n9755 = ~controllable_hmaster1 & ~n9754;
  assign n9756 = controllable_hmaster0 & ~n9755;
  assign n9757 = controllable_hmaster0 & ~n9756;
  assign n9758 = ~controllable_hmaster3 & ~n9757;
  assign n9759 = ~controllable_hmaster3 & ~n9758;
  assign n9760 = i_hbusreq7 & ~n9759;
  assign n9761 = i_hbusreq8 & ~n9757;
  assign n9762 = i_hbusreq6 & ~n9755;
  assign n9763 = controllable_hmaster2 & ~n8527;
  assign n9764 = ~controllable_hmaster1 & ~n9763;
  assign n9765 = ~controllable_hmaster1 & ~n9764;
  assign n9766 = ~i_hbusreq6 & ~n9765;
  assign n9767 = ~n9762 & ~n9766;
  assign n9768 = controllable_hmaster0 & ~n9767;
  assign n9769 = controllable_hmaster0 & ~n9768;
  assign n9770 = ~i_hbusreq8 & ~n9769;
  assign n9771 = ~n9761 & ~n9770;
  assign n9772 = ~controllable_hmaster3 & ~n9771;
  assign n9773 = ~controllable_hmaster3 & ~n9772;
  assign n9774 = ~i_hbusreq7 & ~n9773;
  assign n9775 = ~n9760 & ~n9774;
  assign n9776 = n7924 & ~n9775;
  assign n9777 = n7924 & ~n9776;
  assign n9778 = ~n8214 & ~n9777;
  assign n9779 = controllable_hmaster2 & ~n8434;
  assign n9780 = ~controllable_hmaster1 & ~n9779;
  assign n9781 = ~controllable_hmaster1 & ~n9780;
  assign n9782 = ~controllable_hmaster0 & ~n9781;
  assign n9783 = ~controllable_hmaster0 & ~n9782;
  assign n9784 = ~controllable_hmaster3 & ~n9783;
  assign n9785 = ~controllable_hmaster3 & ~n9784;
  assign n9786 = i_hbusreq7 & ~n9785;
  assign n9787 = i_hbusreq8 & ~n9783;
  assign n9788 = i_hbusreq6 & ~n9781;
  assign n9789 = controllable_hmaster2 & ~n8610;
  assign n9790 = ~controllable_hmaster1 & ~n9789;
  assign n9791 = ~controllable_hmaster1 & ~n9790;
  assign n9792 = ~i_hbusreq6 & ~n9791;
  assign n9793 = ~n9788 & ~n9792;
  assign n9794 = ~controllable_hmaster0 & ~n9793;
  assign n9795 = ~controllable_hmaster0 & ~n9794;
  assign n9796 = ~i_hbusreq8 & ~n9795;
  assign n9797 = ~n9787 & ~n9796;
  assign n9798 = ~controllable_hmaster3 & ~n9797;
  assign n9799 = ~controllable_hmaster3 & ~n9798;
  assign n9800 = ~i_hbusreq7 & ~n9799;
  assign n9801 = ~n9786 & ~n9800;
  assign n9802 = n7924 & ~n9801;
  assign n9803 = n7924 & ~n9802;
  assign n9804 = n8214 & ~n9803;
  assign n9805 = ~n9778 & ~n9804;
  assign n9806 = ~n8202 & ~n9805;
  assign n9807 = controllable_hmaster1 & ~n8375;
  assign n9808 = controllable_hmaster0 & ~n9807;
  assign n9809 = controllable_hmaster0 & ~n9808;
  assign n9810 = ~controllable_hmaster3 & ~n9809;
  assign n9811 = ~controllable_hmaster3 & ~n9810;
  assign n9812 = i_hbusreq7 & ~n9811;
  assign n9813 = i_hbusreq8 & ~n9809;
  assign n9814 = i_hbusreq6 & ~n9807;
  assign n9815 = controllable_hmaster1 & ~n8516;
  assign n9816 = ~i_hbusreq6 & ~n9815;
  assign n9817 = ~n9814 & ~n9816;
  assign n9818 = controllable_hmaster0 & ~n9817;
  assign n9819 = controllable_hmaster0 & ~n9818;
  assign n9820 = ~i_hbusreq8 & ~n9819;
  assign n9821 = ~n9813 & ~n9820;
  assign n9822 = ~controllable_hmaster3 & ~n9821;
  assign n9823 = ~controllable_hmaster3 & ~n9822;
  assign n9824 = ~i_hbusreq7 & ~n9823;
  assign n9825 = ~n9812 & ~n9824;
  assign n9826 = n7924 & ~n9825;
  assign n9827 = n7924 & ~n9826;
  assign n9828 = ~n8214 & ~n9827;
  assign n9829 = controllable_hmaster1 & ~n8423;
  assign n9830 = ~controllable_hmaster0 & ~n9829;
  assign n9831 = ~controllable_hmaster0 & ~n9830;
  assign n9832 = ~controllable_hmaster3 & ~n9831;
  assign n9833 = ~controllable_hmaster3 & ~n9832;
  assign n9834 = i_hbusreq7 & ~n9833;
  assign n9835 = i_hbusreq8 & ~n9831;
  assign n9836 = i_hbusreq6 & ~n9829;
  assign n9837 = controllable_hmaster1 & ~n8590;
  assign n9838 = ~i_hbusreq6 & ~n9837;
  assign n9839 = ~n9836 & ~n9838;
  assign n9840 = ~controllable_hmaster0 & ~n9839;
  assign n9841 = ~controllable_hmaster0 & ~n9840;
  assign n9842 = ~i_hbusreq8 & ~n9841;
  assign n9843 = ~n9835 & ~n9842;
  assign n9844 = ~controllable_hmaster3 & ~n9843;
  assign n9845 = ~controllable_hmaster3 & ~n9844;
  assign n9846 = ~i_hbusreq7 & ~n9845;
  assign n9847 = ~n9834 & ~n9846;
  assign n9848 = n7924 & ~n9847;
  assign n9849 = n7924 & ~n9848;
  assign n9850 = n8214 & ~n9849;
  assign n9851 = ~n9828 & ~n9850;
  assign n9852 = n8202 & ~n9851;
  assign n9853 = ~n9806 & ~n9852;
  assign n9854 = n7728 & ~n9853;
  assign n9855 = ~n7743 & ~n9758;
  assign n9856 = i_hbusreq7 & ~n9855;
  assign n9857 = ~n7779 & ~n9772;
  assign n9858 = ~i_hbusreq7 & ~n9857;
  assign n9859 = ~n9856 & ~n9858;
  assign n9860 = n7924 & ~n9859;
  assign n9861 = ~n8337 & ~n9860;
  assign n9862 = ~n8214 & ~n9861;
  assign n9863 = ~n7743 & ~n9784;
  assign n9864 = i_hbusreq7 & ~n9863;
  assign n9865 = ~n7779 & ~n9798;
  assign n9866 = ~i_hbusreq7 & ~n9865;
  assign n9867 = ~n9864 & ~n9866;
  assign n9868 = n7924 & ~n9867;
  assign n9869 = ~n8337 & ~n9868;
  assign n9870 = n8214 & ~n9869;
  assign n9871 = ~n9862 & ~n9870;
  assign n9872 = ~n8202 & ~n9871;
  assign n9873 = ~n7743 & ~n9810;
  assign n9874 = i_hbusreq7 & ~n9873;
  assign n9875 = ~n7779 & ~n9822;
  assign n9876 = ~i_hbusreq7 & ~n9875;
  assign n9877 = ~n9874 & ~n9876;
  assign n9878 = n7924 & ~n9877;
  assign n9879 = ~n8337 & ~n9878;
  assign n9880 = ~n8214 & ~n9879;
  assign n9881 = ~n7743 & ~n9832;
  assign n9882 = i_hbusreq7 & ~n9881;
  assign n9883 = ~n7779 & ~n9844;
  assign n9884 = ~i_hbusreq7 & ~n9883;
  assign n9885 = ~n9882 & ~n9884;
  assign n9886 = n7924 & ~n9885;
  assign n9887 = ~n8337 & ~n9886;
  assign n9888 = n8214 & ~n9887;
  assign n9889 = ~n9880 & ~n9888;
  assign n9890 = n8202 & ~n9889;
  assign n9891 = ~n9872 & ~n9890;
  assign n9892 = ~n7728 & ~n9891;
  assign n9893 = ~n9854 & ~n9892;
  assign n9894 = ~n7723 & ~n9893;
  assign n9895 = ~n7723 & ~n9894;
  assign n9896 = ~n7714 & ~n9895;
  assign n9897 = ~n7714 & ~n9896;
  assign n9898 = n7705 & ~n9897;
  assign n9899 = n7723 & ~n9891;
  assign n9900 = n7920 & ~n9891;
  assign n9901 = ~n8640 & ~n9900;
  assign n9902 = ~n7723 & ~n9901;
  assign n9903 = ~n9899 & ~n9902;
  assign n9904 = n7714 & ~n9903;
  assign n9905 = ~n8646 & ~n9904;
  assign n9906 = ~n7705 & ~n9905;
  assign n9907 = ~n9898 & ~n9906;
  assign n9908 = ~n7808 & ~n9907;
  assign n9909 = ~n7920 & ~n9853;
  assign n9910 = controllable_hmaster2 & ~n9199;
  assign n9911 = ~controllable_hmaster1 & ~n9910;
  assign n9912 = ~controllable_hmaster1 & ~n9911;
  assign n9913 = controllable_hmaster0 & ~n9912;
  assign n9914 = controllable_hmaster0 & ~n9913;
  assign n9915 = ~controllable_hmaster3 & ~n9914;
  assign n9916 = ~controllable_hmaster3 & ~n9915;
  assign n9917 = i_hbusreq7 & ~n9916;
  assign n9918 = i_hbusreq8 & ~n9914;
  assign n9919 = i_hbusreq6 & ~n9912;
  assign n9920 = controllable_hmaster2 & ~n9646;
  assign n9921 = ~controllable_hmaster1 & ~n9920;
  assign n9922 = ~controllable_hmaster1 & ~n9921;
  assign n9923 = ~i_hbusreq6 & ~n9922;
  assign n9924 = ~n9919 & ~n9923;
  assign n9925 = controllable_hmaster0 & ~n9924;
  assign n9926 = controllable_hmaster0 & ~n9925;
  assign n9927 = ~i_hbusreq8 & ~n9926;
  assign n9928 = ~n9918 & ~n9927;
  assign n9929 = ~controllable_hmaster3 & ~n9928;
  assign n9930 = ~controllable_hmaster3 & ~n9929;
  assign n9931 = ~i_hbusreq7 & ~n9930;
  assign n9932 = ~n9917 & ~n9931;
  assign n9933 = ~n8214 & ~n9932;
  assign n9934 = controllable_hmaster2 & ~n9221;
  assign n9935 = ~controllable_hmaster1 & ~n9934;
  assign n9936 = ~controllable_hmaster1 & ~n9935;
  assign n9937 = ~controllable_hmaster0 & ~n9936;
  assign n9938 = ~controllable_hmaster0 & ~n9937;
  assign n9939 = ~controllable_hmaster3 & ~n9938;
  assign n9940 = ~controllable_hmaster3 & ~n9939;
  assign n9941 = i_hbusreq7 & ~n9940;
  assign n9942 = i_hbusreq8 & ~n9938;
  assign n9943 = i_hbusreq6 & ~n9936;
  assign n9944 = controllable_hmaster2 & ~n9688;
  assign n9945 = ~controllable_hmaster1 & ~n9944;
  assign n9946 = ~controllable_hmaster1 & ~n9945;
  assign n9947 = ~i_hbusreq6 & ~n9946;
  assign n9948 = ~n9943 & ~n9947;
  assign n9949 = ~controllable_hmaster0 & ~n9948;
  assign n9950 = ~controllable_hmaster0 & ~n9949;
  assign n9951 = ~i_hbusreq8 & ~n9950;
  assign n9952 = ~n9942 & ~n9951;
  assign n9953 = ~controllable_hmaster3 & ~n9952;
  assign n9954 = ~controllable_hmaster3 & ~n9953;
  assign n9955 = ~i_hbusreq7 & ~n9954;
  assign n9956 = ~n9941 & ~n9955;
  assign n9957 = n8214 & ~n9956;
  assign n9958 = ~n9933 & ~n9957;
  assign n9959 = ~n8202 & ~n9958;
  assign n9960 = ~controllable_hmaster2 & ~n9193;
  assign n9961 = controllable_hmaster1 & ~n9960;
  assign n9962 = controllable_hmaster1 & ~n9961;
  assign n9963 = controllable_hmaster0 & ~n9962;
  assign n9964 = controllable_hmaster0 & ~n9963;
  assign n9965 = ~controllable_hmaster3 & ~n9964;
  assign n9966 = ~controllable_hmaster3 & ~n9965;
  assign n9967 = i_hbusreq7 & ~n9966;
  assign n9968 = i_hbusreq8 & ~n9964;
  assign n9969 = i_hbusreq6 & ~n9962;
  assign n9970 = ~controllable_hmaster2 & ~n9638;
  assign n9971 = controllable_hmaster1 & ~n9970;
  assign n9972 = controllable_hmaster1 & ~n9971;
  assign n9973 = ~i_hbusreq6 & ~n9972;
  assign n9974 = ~n9969 & ~n9973;
  assign n9975 = controllable_hmaster0 & ~n9974;
  assign n9976 = controllable_hmaster0 & ~n9975;
  assign n9977 = ~i_hbusreq8 & ~n9976;
  assign n9978 = ~n9968 & ~n9977;
  assign n9979 = ~controllable_hmaster3 & ~n9978;
  assign n9980 = ~controllable_hmaster3 & ~n9979;
  assign n9981 = ~i_hbusreq7 & ~n9980;
  assign n9982 = ~n9967 & ~n9981;
  assign n9983 = ~n8214 & ~n9982;
  assign n9984 = ~controllable_hmaster2 & ~n9215;
  assign n9985 = controllable_hmaster1 & ~n9984;
  assign n9986 = controllable_hmaster1 & ~n9985;
  assign n9987 = ~controllable_hmaster0 & ~n9986;
  assign n9988 = ~controllable_hmaster0 & ~n9987;
  assign n9989 = ~controllable_hmaster3 & ~n9988;
  assign n9990 = ~controllable_hmaster3 & ~n9989;
  assign n9991 = i_hbusreq7 & ~n9990;
  assign n9992 = i_hbusreq8 & ~n9988;
  assign n9993 = i_hbusreq6 & ~n9986;
  assign n9994 = ~controllable_hmaster2 & ~n9678;
  assign n9995 = controllable_hmaster1 & ~n9994;
  assign n9996 = controllable_hmaster1 & ~n9995;
  assign n9997 = ~i_hbusreq6 & ~n9996;
  assign n9998 = ~n9993 & ~n9997;
  assign n9999 = ~controllable_hmaster0 & ~n9998;
  assign n10000 = ~controllable_hmaster0 & ~n9999;
  assign n10001 = ~i_hbusreq8 & ~n10000;
  assign n10002 = ~n9992 & ~n10001;
  assign n10003 = ~controllable_hmaster3 & ~n10002;
  assign n10004 = ~controllable_hmaster3 & ~n10003;
  assign n10005 = ~i_hbusreq7 & ~n10004;
  assign n10006 = ~n9991 & ~n10005;
  assign n10007 = n8214 & ~n10006;
  assign n10008 = ~n9983 & ~n10007;
  assign n10009 = n8202 & ~n10008;
  assign n10010 = ~n9959 & ~n10009;
  assign n10011 = n7920 & ~n10010;
  assign n10012 = ~n9909 & ~n10011;
  assign n10013 = n7728 & ~n10012;
  assign n10014 = ~n7920 & ~n9891;
  assign n10015 = ~n7743 & ~n9915;
  assign n10016 = i_hbusreq7 & ~n10015;
  assign n10017 = ~n7779 & ~n9929;
  assign n10018 = ~i_hbusreq7 & ~n10017;
  assign n10019 = ~n10016 & ~n10018;
  assign n10020 = ~n8214 & ~n10019;
  assign n10021 = ~n7743 & ~n9939;
  assign n10022 = i_hbusreq7 & ~n10021;
  assign n10023 = ~n7779 & ~n9953;
  assign n10024 = ~i_hbusreq7 & ~n10023;
  assign n10025 = ~n10022 & ~n10024;
  assign n10026 = n8214 & ~n10025;
  assign n10027 = ~n10020 & ~n10026;
  assign n10028 = ~n8202 & ~n10027;
  assign n10029 = ~n7743 & ~n9965;
  assign n10030 = i_hbusreq7 & ~n10029;
  assign n10031 = ~n7779 & ~n9979;
  assign n10032 = ~i_hbusreq7 & ~n10031;
  assign n10033 = ~n10030 & ~n10032;
  assign n10034 = ~n8214 & ~n10033;
  assign n10035 = ~n7743 & ~n9989;
  assign n10036 = i_hbusreq7 & ~n10035;
  assign n10037 = ~n7779 & ~n10003;
  assign n10038 = ~i_hbusreq7 & ~n10037;
  assign n10039 = ~n10036 & ~n10038;
  assign n10040 = n8214 & ~n10039;
  assign n10041 = ~n10034 & ~n10040;
  assign n10042 = n8202 & ~n10041;
  assign n10043 = ~n10028 & ~n10042;
  assign n10044 = n7920 & ~n10043;
  assign n10045 = ~n10014 & ~n10044;
  assign n10046 = ~n7728 & ~n10045;
  assign n10047 = ~n10013 & ~n10046;
  assign n10048 = ~n7723 & ~n10047;
  assign n10049 = ~n7723 & ~n10048;
  assign n10050 = ~n7714 & ~n10049;
  assign n10051 = ~n7714 & ~n10050;
  assign n10052 = n7705 & ~n10051;
  assign n10053 = controllable_hmaster1 & ~n8987;
  assign n10054 = ~n8988 & ~n9199;
  assign n10055 = ~controllable_hmaster1 & ~n10054;
  assign n10056 = ~n10053 & ~n10055;
  assign n10057 = controllable_hmaster0 & ~n10056;
  assign n10058 = ~n9099 & ~n10057;
  assign n10059 = ~controllable_hmaster3 & ~n10058;
  assign n10060 = ~n9093 & ~n10059;
  assign n10061 = i_hbusreq7 & ~n10060;
  assign n10062 = i_hbusreq8 & ~n10058;
  assign n10063 = i_hbusreq6 & ~n10056;
  assign n10064 = controllable_hmaster1 & ~n9023;
  assign n10065 = ~n9024 & ~n9646;
  assign n10066 = ~controllable_hmaster1 & ~n10065;
  assign n10067 = ~n10064 & ~n10066;
  assign n10068 = ~i_hbusreq6 & ~n10067;
  assign n10069 = ~n10063 & ~n10068;
  assign n10070 = controllable_hmaster0 & ~n10069;
  assign n10071 = ~n9127 & ~n10070;
  assign n10072 = ~i_hbusreq8 & ~n10071;
  assign n10073 = ~n10062 & ~n10072;
  assign n10074 = ~controllable_hmaster3 & ~n10073;
  assign n10075 = ~n9117 & ~n10074;
  assign n10076 = ~i_hbusreq7 & ~n10075;
  assign n10077 = ~n10061 & ~n10076;
  assign n10078 = ~n8214 & ~n10077;
  assign n10079 = ~n8988 & ~n9221;
  assign n10080 = ~controllable_hmaster1 & ~n10079;
  assign n10081 = ~n10053 & ~n10080;
  assign n10082 = ~controllable_hmaster0 & ~n10081;
  assign n10083 = ~n9152 & ~n10082;
  assign n10084 = ~controllable_hmaster3 & ~n10083;
  assign n10085 = ~n9093 & ~n10084;
  assign n10086 = i_hbusreq7 & ~n10085;
  assign n10087 = i_hbusreq8 & ~n10083;
  assign n10088 = i_hbusreq6 & ~n10081;
  assign n10089 = ~n9024 & ~n9688;
  assign n10090 = ~controllable_hmaster1 & ~n10089;
  assign n10091 = ~n10064 & ~n10090;
  assign n10092 = ~i_hbusreq6 & ~n10091;
  assign n10093 = ~n10088 & ~n10092;
  assign n10094 = ~controllable_hmaster0 & ~n10093;
  assign n10095 = ~n9162 & ~n10094;
  assign n10096 = ~i_hbusreq8 & ~n10095;
  assign n10097 = ~n10087 & ~n10096;
  assign n10098 = ~controllable_hmaster3 & ~n10097;
  assign n10099 = ~n9117 & ~n10098;
  assign n10100 = ~i_hbusreq7 & ~n10099;
  assign n10101 = ~n10086 & ~n10100;
  assign n10102 = n8214 & ~n10101;
  assign n10103 = ~n10078 & ~n10102;
  assign n10104 = ~n8202 & ~n10103;
  assign n10105 = controllable_hmaster2 & ~n8987;
  assign n10106 = ~n9193 & ~n10105;
  assign n10107 = controllable_hmaster1 & ~n10106;
  assign n10108 = ~n9096 & ~n10107;
  assign n10109 = controllable_hmaster0 & ~n10108;
  assign n10110 = ~n9099 & ~n10109;
  assign n10111 = ~controllable_hmaster3 & ~n10110;
  assign n10112 = ~n9093 & ~n10111;
  assign n10113 = i_hbusreq7 & ~n10112;
  assign n10114 = i_hbusreq8 & ~n10110;
  assign n10115 = i_hbusreq6 & ~n10108;
  assign n10116 = controllable_hmaster2 & ~n9023;
  assign n10117 = ~n9638 & ~n10116;
  assign n10118 = controllable_hmaster1 & ~n10117;
  assign n10119 = ~n9122 & ~n10118;
  assign n10120 = ~i_hbusreq6 & ~n10119;
  assign n10121 = ~n10115 & ~n10120;
  assign n10122 = controllable_hmaster0 & ~n10121;
  assign n10123 = ~n9127 & ~n10122;
  assign n10124 = ~i_hbusreq8 & ~n10123;
  assign n10125 = ~n10114 & ~n10124;
  assign n10126 = ~controllable_hmaster3 & ~n10125;
  assign n10127 = ~n9117 & ~n10126;
  assign n10128 = ~i_hbusreq7 & ~n10127;
  assign n10129 = ~n10113 & ~n10128;
  assign n10130 = ~n8214 & ~n10129;
  assign n10131 = ~n9215 & ~n10105;
  assign n10132 = controllable_hmaster1 & ~n10131;
  assign n10133 = ~n9096 & ~n10132;
  assign n10134 = ~controllable_hmaster0 & ~n10133;
  assign n10135 = ~n9152 & ~n10134;
  assign n10136 = ~controllable_hmaster3 & ~n10135;
  assign n10137 = ~n9093 & ~n10136;
  assign n10138 = i_hbusreq7 & ~n10137;
  assign n10139 = i_hbusreq8 & ~n10135;
  assign n10140 = i_hbusreq6 & ~n10133;
  assign n10141 = ~n9678 & ~n10116;
  assign n10142 = controllable_hmaster1 & ~n10141;
  assign n10143 = ~n9122 & ~n10142;
  assign n10144 = ~i_hbusreq6 & ~n10143;
  assign n10145 = ~n10140 & ~n10144;
  assign n10146 = ~controllable_hmaster0 & ~n10145;
  assign n10147 = ~n9162 & ~n10146;
  assign n10148 = ~i_hbusreq8 & ~n10147;
  assign n10149 = ~n10139 & ~n10148;
  assign n10150 = ~controllable_hmaster3 & ~n10149;
  assign n10151 = ~n9117 & ~n10150;
  assign n10152 = ~i_hbusreq7 & ~n10151;
  assign n10153 = ~n10138 & ~n10152;
  assign n10154 = n8214 & ~n10153;
  assign n10155 = ~n10130 & ~n10154;
  assign n10156 = n8202 & ~n10155;
  assign n10157 = ~n10104 & ~n10156;
  assign n10158 = n7920 & ~n10157;
  assign n10159 = ~n10014 & ~n10158;
  assign n10160 = n7728 & ~n10159;
  assign n10161 = ~n9358 & ~n9646;
  assign n10162 = ~controllable_hmaster1 & ~n10161;
  assign n10163 = ~n9332 & ~n10162;
  assign n10164 = ~i_hbusreq6 & ~n10163;
  assign n10165 = ~n9313 & ~n10164;
  assign n10166 = controllable_hmaster0 & ~n10165;
  assign n10167 = ~n9439 & ~n10166;
  assign n10168 = ~i_hbusreq8 & ~n10167;
  assign n10169 = ~n9312 & ~n10168;
  assign n10170 = ~controllable_hmaster3 & ~n10169;
  assign n10171 = ~n9517 & ~n10170;
  assign n10172 = i_hlock7 & ~n10171;
  assign n10173 = ~n9449 & ~n10162;
  assign n10174 = ~i_hbusreq6 & ~n10173;
  assign n10175 = ~n9447 & ~n10174;
  assign n10176 = controllable_hmaster0 & ~n10175;
  assign n10177 = ~n9439 & ~n10176;
  assign n10178 = ~i_hbusreq8 & ~n10177;
  assign n10179 = ~n9446 & ~n10178;
  assign n10180 = ~controllable_hmaster3 & ~n10179;
  assign n10181 = ~n9517 & ~n10180;
  assign n10182 = ~i_hlock7 & ~n10181;
  assign n10183 = ~n10172 & ~n10182;
  assign n10184 = ~i_hbusreq7 & ~n10183;
  assign n10185 = ~n9247 & ~n10184;
  assign n10186 = ~n8214 & ~n10185;
  assign n10187 = ~n9426 & ~n9688;
  assign n10188 = ~controllable_hmaster1 & ~n10187;
  assign n10189 = ~n9393 & ~n10188;
  assign n10190 = i_hlock6 & ~n10189;
  assign n10191 = ~n9433 & ~n10188;
  assign n10192 = ~i_hlock6 & ~n10191;
  assign n10193 = ~n10190 & ~n10192;
  assign n10194 = ~i_hbusreq6 & ~n10193;
  assign n10195 = ~n9365 & ~n10194;
  assign n10196 = ~controllable_hmaster0 & ~n10195;
  assign n10197 = ~n9364 & ~n10196;
  assign n10198 = ~i_hbusreq8 & ~n10197;
  assign n10199 = ~n9312 & ~n10198;
  assign n10200 = ~controllable_hmaster3 & ~n10199;
  assign n10201 = ~n9517 & ~n10200;
  assign n10202 = i_hlock7 & ~n10201;
  assign n10203 = ~n9453 & ~n10196;
  assign n10204 = ~i_hbusreq8 & ~n10203;
  assign n10205 = ~n9446 & ~n10204;
  assign n10206 = ~controllable_hmaster3 & ~n10205;
  assign n10207 = ~n9517 & ~n10206;
  assign n10208 = ~i_hlock7 & ~n10207;
  assign n10209 = ~n10202 & ~n10208;
  assign n10210 = ~i_hbusreq7 & ~n10209;
  assign n10211 = ~n9247 & ~n10210;
  assign n10212 = n8214 & ~n10211;
  assign n10213 = ~n10186 & ~n10212;
  assign n10214 = ~n8202 & ~n10213;
  assign n10215 = ~n9314 & ~n9638;
  assign n10216 = controllable_hmaster1 & ~n10215;
  assign n10217 = ~n9360 & ~n10216;
  assign n10218 = ~i_hbusreq6 & ~n10217;
  assign n10219 = ~n9313 & ~n10218;
  assign n10220 = controllable_hmaster0 & ~n10219;
  assign n10221 = ~n9439 & ~n10220;
  assign n10222 = ~i_hbusreq8 & ~n10221;
  assign n10223 = ~n9312 & ~n10222;
  assign n10224 = ~controllable_hmaster3 & ~n10223;
  assign n10225 = ~n9517 & ~n10224;
  assign n10226 = i_hlock7 & ~n10225;
  assign n10227 = ~n9431 & ~n9638;
  assign n10228 = controllable_hmaster1 & ~n10227;
  assign n10229 = ~n9360 & ~n10228;
  assign n10230 = ~i_hbusreq6 & ~n10229;
  assign n10231 = ~n9447 & ~n10230;
  assign n10232 = controllable_hmaster0 & ~n10231;
  assign n10233 = ~n9439 & ~n10232;
  assign n10234 = ~i_hbusreq8 & ~n10233;
  assign n10235 = ~n9446 & ~n10234;
  assign n10236 = ~controllable_hmaster3 & ~n10235;
  assign n10237 = ~n9517 & ~n10236;
  assign n10238 = ~i_hlock7 & ~n10237;
  assign n10239 = ~n10226 & ~n10238;
  assign n10240 = ~i_hbusreq7 & ~n10239;
  assign n10241 = ~n9247 & ~n10240;
  assign n10242 = ~n8214 & ~n10241;
  assign n10243 = ~n9314 & ~n9678;
  assign n10244 = controllable_hmaster1 & ~n10243;
  assign n10245 = ~n9428 & ~n10244;
  assign n10246 = i_hlock6 & ~n10245;
  assign n10247 = ~n9431 & ~n9678;
  assign n10248 = controllable_hmaster1 & ~n10247;
  assign n10249 = ~n9428 & ~n10248;
  assign n10250 = ~i_hlock6 & ~n10249;
  assign n10251 = ~n10246 & ~n10250;
  assign n10252 = ~i_hbusreq6 & ~n10251;
  assign n10253 = ~n9365 & ~n10252;
  assign n10254 = ~controllable_hmaster0 & ~n10253;
  assign n10255 = ~n9364 & ~n10254;
  assign n10256 = ~i_hbusreq8 & ~n10255;
  assign n10257 = ~n9312 & ~n10256;
  assign n10258 = ~controllable_hmaster3 & ~n10257;
  assign n10259 = ~n9517 & ~n10258;
  assign n10260 = i_hlock7 & ~n10259;
  assign n10261 = ~n9453 & ~n10254;
  assign n10262 = ~i_hbusreq8 & ~n10261;
  assign n10263 = ~n9446 & ~n10262;
  assign n10264 = ~controllable_hmaster3 & ~n10263;
  assign n10265 = ~n9517 & ~n10264;
  assign n10266 = ~i_hlock7 & ~n10265;
  assign n10267 = ~n10260 & ~n10266;
  assign n10268 = ~i_hbusreq7 & ~n10267;
  assign n10269 = ~n9247 & ~n10268;
  assign n10270 = n8214 & ~n10269;
  assign n10271 = ~n10242 & ~n10270;
  assign n10272 = n8202 & ~n10271;
  assign n10273 = ~n10214 & ~n10272;
  assign n10274 = n7920 & ~n10273;
  assign n10275 = ~n10014 & ~n10274;
  assign n10276 = ~n7728 & ~n10275;
  assign n10277 = ~n10160 & ~n10276;
  assign n10278 = n7723 & ~n10277;
  assign n10279 = ~n7723 & ~n10275;
  assign n10280 = ~n10278 & ~n10279;
  assign n10281 = n7714 & ~n10280;
  assign n10282 = n7723 & ~n10275;
  assign n10283 = ~n8640 & ~n10274;
  assign n10284 = n7728 & ~n10283;
  assign n10285 = ~n9740 & ~n10284;
  assign n10286 = ~n7723 & ~n10285;
  assign n10287 = ~n10282 & ~n10286;
  assign n10288 = ~n7714 & ~n10287;
  assign n10289 = ~n10281 & ~n10288;
  assign n10290 = ~n7705 & ~n10289;
  assign n10291 = ~n10052 & ~n10290;
  assign n10292 = n7808 & ~n10291;
  assign n10293 = ~n9908 & ~n10292;
  assign n10294 = ~n8195 & ~n10293;
  assign n10295 = ~controllable_hmaster2 & ~n8397;
  assign n10296 = ~controllable_hmaster1 & ~n10295;
  assign n10297 = ~controllable_hmaster1 & ~n10296;
  assign n10298 = controllable_hmaster0 & ~n10297;
  assign n10299 = controllable_hmaster0 & ~n10298;
  assign n10300 = ~controllable_hmaster3 & ~n10299;
  assign n10301 = ~controllable_hmaster3 & ~n10300;
  assign n10302 = i_hbusreq7 & ~n10301;
  assign n10303 = i_hbusreq8 & ~n10299;
  assign n10304 = i_hbusreq6 & ~n10297;
  assign n10305 = ~controllable_hmaster2 & ~n8550;
  assign n10306 = ~controllable_hmaster1 & ~n10305;
  assign n10307 = ~controllable_hmaster1 & ~n10306;
  assign n10308 = ~i_hbusreq6 & ~n10307;
  assign n10309 = ~n10304 & ~n10308;
  assign n10310 = controllable_hmaster0 & ~n10309;
  assign n10311 = controllable_hmaster0 & ~n10310;
  assign n10312 = ~i_hbusreq8 & ~n10311;
  assign n10313 = ~n10303 & ~n10312;
  assign n10314 = ~controllable_hmaster3 & ~n10313;
  assign n10315 = ~controllable_hmaster3 & ~n10314;
  assign n10316 = ~i_hbusreq7 & ~n10315;
  assign n10317 = ~n10302 & ~n10316;
  assign n10318 = n7924 & ~n10317;
  assign n10319 = n7924 & ~n10318;
  assign n10320 = ~n8214 & ~n10319;
  assign n10321 = ~controllable_hmaster2 & ~n8443;
  assign n10322 = ~controllable_hmaster1 & ~n10321;
  assign n10323 = ~controllable_hmaster1 & ~n10322;
  assign n10324 = ~controllable_hmaster0 & ~n10323;
  assign n10325 = ~controllable_hmaster0 & ~n10324;
  assign n10326 = ~controllable_hmaster3 & ~n10325;
  assign n10327 = ~controllable_hmaster3 & ~n10326;
  assign n10328 = n7924 & ~n10327;
  assign n10329 = n7924 & ~n10328;
  assign n10330 = n8214 & ~n10329;
  assign n10331 = ~n10320 & ~n10330;
  assign n10332 = ~n8202 & ~n10331;
  assign n10333 = ~n7737 & n7928;
  assign n10334 = n7928 & ~n10333;
  assign n10335 = controllable_hmaster1 & ~n10334;
  assign n10336 = controllable_hmaster2 & ~n10334;
  assign n10337 = controllable_hmaster2 & ~n10336;
  assign n10338 = ~controllable_hmaster1 & ~n10337;
  assign n10339 = ~n10335 & ~n10338;
  assign n10340 = controllable_hmaster3 & ~n10339;
  assign n10341 = controllable_hmaster3 & ~n10340;
  assign n10342 = i_hbusreq7 & ~n10341;
  assign n10343 = i_hbusreq8 & ~n10339;
  assign n10344 = i_hbusreq6 & ~n10339;
  assign n10345 = i_hbusreq5 & ~n10334;
  assign n10346 = i_hbusreq4 & ~n10334;
  assign n10347 = i_hbusreq9 & ~n10334;
  assign n10348 = i_hbusreq3 & ~n10334;
  assign n10349 = i_hbusreq1 & ~n10334;
  assign n10350 = ~n7759 & n7928;
  assign n10351 = n7928 & ~n10350;
  assign n10352 = ~i_hbusreq1 & ~n10351;
  assign n10353 = ~n10349 & ~n10352;
  assign n10354 = ~i_hbusreq3 & ~n10353;
  assign n10355 = ~n10348 & ~n10354;
  assign n10356 = ~i_hbusreq9 & ~n10355;
  assign n10357 = ~n10347 & ~n10356;
  assign n10358 = ~i_hbusreq4 & ~n10357;
  assign n10359 = ~n10346 & ~n10358;
  assign n10360 = ~i_hbusreq5 & ~n10359;
  assign n10361 = ~n10345 & ~n10360;
  assign n10362 = controllable_hmaster1 & ~n10361;
  assign n10363 = controllable_hmaster2 & ~n10361;
  assign n10364 = controllable_hmaster2 & ~n10363;
  assign n10365 = ~controllable_hmaster1 & ~n10364;
  assign n10366 = ~n10362 & ~n10365;
  assign n10367 = ~i_hbusreq6 & ~n10366;
  assign n10368 = ~n10344 & ~n10367;
  assign n10369 = ~i_hbusreq8 & ~n10368;
  assign n10370 = ~n10343 & ~n10369;
  assign n10371 = controllable_hmaster3 & ~n10370;
  assign n10372 = controllable_hmaster3 & ~n10371;
  assign n10373 = ~i_hbusreq7 & ~n10372;
  assign n10374 = ~n10342 & ~n10373;
  assign n10375 = ~n7924 & ~n10374;
  assign n10376 = controllable_hmaster2 & ~n10105;
  assign n10377 = ~controllable_hmaster1 & ~n10376;
  assign n10378 = ~n10053 & ~n10377;
  assign n10379 = controllable_hmaster3 & ~n10378;
  assign n10380 = n7928 & ~n8222;
  assign n10381 = ~n8365 & ~n10380;
  assign n10382 = ~n8365 & ~n10381;
  assign n10383 = i_hlock3 & ~n10382;
  assign n10384 = n7928 & ~n8236;
  assign n10385 = ~n8365 & ~n10384;
  assign n10386 = ~n8365 & ~n10385;
  assign n10387 = ~i_hlock3 & ~n10386;
  assign n10388 = ~n10383 & ~n10387;
  assign n10389 = ~controllable_hmaster2 & ~n10388;
  assign n10390 = ~controllable_hmaster2 & ~n10389;
  assign n10391 = controllable_hmaster1 & ~n10390;
  assign n10392 = ~n8378 & ~n10380;
  assign n10393 = ~n8378 & ~n10392;
  assign n10394 = i_hlock5 & ~n10393;
  assign n10395 = ~n8378 & ~n10384;
  assign n10396 = ~n8378 & ~n10395;
  assign n10397 = ~i_hlock5 & ~n10396;
  assign n10398 = ~n10394 & ~n10397;
  assign n10399 = controllable_hmaster2 & ~n10398;
  assign n10400 = ~n8389 & ~n10380;
  assign n10401 = ~n8389 & ~n10400;
  assign n10402 = i_hlock1 & ~n10401;
  assign n10403 = ~n8389 & ~n10384;
  assign n10404 = ~n8389 & ~n10403;
  assign n10405 = ~i_hlock1 & ~n10404;
  assign n10406 = ~n10402 & ~n10405;
  assign n10407 = ~controllable_hmaster2 & ~n10406;
  assign n10408 = ~n10399 & ~n10407;
  assign n10409 = ~controllable_hmaster1 & ~n10408;
  assign n10410 = ~n10391 & ~n10409;
  assign n10411 = controllable_hmaster0 & ~n10410;
  assign n10412 = n7928 & ~n8419;
  assign n10413 = ~controllable_hmaster2 & ~n10412;
  assign n10414 = ~controllable_hmaster2 & ~n10413;
  assign n10415 = controllable_hmaster1 & ~n10414;
  assign n10416 = ~n8426 & ~n10380;
  assign n10417 = ~n8426 & ~n10416;
  assign n10418 = i_hlock4 & ~n10417;
  assign n10419 = ~n8426 & ~n10384;
  assign n10420 = ~n8426 & ~n10419;
  assign n10421 = ~i_hlock4 & ~n10420;
  assign n10422 = ~n10418 & ~n10421;
  assign n10423 = controllable_hmaster2 & ~n10422;
  assign n10424 = n7928 & ~n8441;
  assign n10425 = ~controllable_hmaster2 & ~n10424;
  assign n10426 = ~n10423 & ~n10425;
  assign n10427 = ~controllable_hmaster1 & ~n10426;
  assign n10428 = ~n10415 & ~n10427;
  assign n10429 = n8217 & ~n10428;
  assign n10430 = controllable_hmaster2 & ~n10380;
  assign n10431 = ~n10413 & ~n10430;
  assign n10432 = controllable_hmaster1 & ~n10431;
  assign n10433 = ~n10427 & ~n10432;
  assign n10434 = ~n8217 & ~n10433;
  assign n10435 = ~n10429 & ~n10434;
  assign n10436 = i_hlock6 & ~n10435;
  assign n10437 = controllable_hmaster2 & ~n10384;
  assign n10438 = ~n10413 & ~n10437;
  assign n10439 = controllable_hmaster1 & ~n10438;
  assign n10440 = ~n10427 & ~n10439;
  assign n10441 = ~n8217 & ~n10440;
  assign n10442 = ~n10429 & ~n10441;
  assign n10443 = ~i_hlock6 & ~n10442;
  assign n10444 = ~n10436 & ~n10443;
  assign n10445 = ~controllable_hmaster0 & ~n10444;
  assign n10446 = ~n10411 & ~n10445;
  assign n10447 = ~controllable_hmaster3 & ~n10446;
  assign n10448 = ~n10379 & ~n10447;
  assign n10449 = i_hbusreq7 & ~n10448;
  assign n10450 = i_hbusreq8 & ~n10378;
  assign n10451 = i_hbusreq6 & ~n10378;
  assign n10452 = controllable_hmaster2 & ~n10116;
  assign n10453 = ~controllable_hmaster1 & ~n10452;
  assign n10454 = ~n10064 & ~n10453;
  assign n10455 = ~i_hbusreq6 & ~n10454;
  assign n10456 = ~n10451 & ~n10455;
  assign n10457 = ~i_hbusreq8 & ~n10456;
  assign n10458 = ~n10450 & ~n10457;
  assign n10459 = controllable_hmaster3 & ~n10458;
  assign n10460 = i_hbusreq8 & ~n10446;
  assign n10461 = i_hbusreq6 & ~n10410;
  assign n10462 = i_hbusreq5 & ~n10388;
  assign n10463 = i_hbusreq4 & ~n10388;
  assign n10464 = i_hbusreq9 & ~n10388;
  assign n10465 = i_hbusreq3 & ~n10388;
  assign n10466 = i_hbusreq1 & ~n10380;
  assign n10467 = n7928 & ~n8266;
  assign n10468 = ~i_hbusreq1 & ~n10467;
  assign n10469 = ~n10466 & ~n10468;
  assign n10470 = ~n8365 & ~n10469;
  assign n10471 = ~n8365 & ~n10470;
  assign n10472 = i_hlock3 & ~n10471;
  assign n10473 = i_hbusreq1 & ~n10384;
  assign n10474 = n7928 & ~n8298;
  assign n10475 = ~i_hbusreq1 & ~n10474;
  assign n10476 = ~n10473 & ~n10475;
  assign n10477 = ~n8365 & ~n10476;
  assign n10478 = ~n8365 & ~n10477;
  assign n10479 = ~i_hlock3 & ~n10478;
  assign n10480 = ~n10472 & ~n10479;
  assign n10481 = ~i_hbusreq3 & ~n10480;
  assign n10482 = ~n10465 & ~n10481;
  assign n10483 = ~i_hbusreq9 & ~n10482;
  assign n10484 = ~n10464 & ~n10483;
  assign n10485 = ~i_hbusreq4 & ~n10484;
  assign n10486 = ~n10463 & ~n10485;
  assign n10487 = ~i_hbusreq5 & ~n10486;
  assign n10488 = ~n10462 & ~n10487;
  assign n10489 = ~controllable_hmaster2 & ~n10488;
  assign n10490 = ~controllable_hmaster2 & ~n10489;
  assign n10491 = controllable_hmaster1 & ~n10490;
  assign n10492 = i_hbusreq5 & ~n10398;
  assign n10493 = i_hbusreq4 & ~n10380;
  assign n10494 = i_hbusreq9 & ~n10380;
  assign n10495 = i_hbusreq3 & ~n10380;
  assign n10496 = ~i_hbusreq3 & ~n10469;
  assign n10497 = ~n10495 & ~n10496;
  assign n10498 = ~i_hbusreq9 & ~n10497;
  assign n10499 = ~n10494 & ~n10498;
  assign n10500 = ~i_hbusreq4 & ~n10499;
  assign n10501 = ~n10493 & ~n10500;
  assign n10502 = ~n8378 & ~n10501;
  assign n10503 = ~n8378 & ~n10502;
  assign n10504 = i_hlock5 & ~n10503;
  assign n10505 = i_hbusreq4 & ~n10384;
  assign n10506 = i_hbusreq9 & ~n10384;
  assign n10507 = i_hbusreq3 & ~n10384;
  assign n10508 = ~i_hbusreq3 & ~n10476;
  assign n10509 = ~n10507 & ~n10508;
  assign n10510 = ~i_hbusreq9 & ~n10509;
  assign n10511 = ~n10506 & ~n10510;
  assign n10512 = ~i_hbusreq4 & ~n10511;
  assign n10513 = ~n10505 & ~n10512;
  assign n10514 = ~n8378 & ~n10513;
  assign n10515 = ~n8378 & ~n10514;
  assign n10516 = ~i_hlock5 & ~n10515;
  assign n10517 = ~n10504 & ~n10516;
  assign n10518 = ~i_hbusreq5 & ~n10517;
  assign n10519 = ~n10492 & ~n10518;
  assign n10520 = controllable_hmaster2 & ~n10519;
  assign n10521 = i_hbusreq5 & ~n10406;
  assign n10522 = i_hbusreq4 & ~n10406;
  assign n10523 = i_hbusreq9 & ~n10406;
  assign n10524 = i_hbusreq3 & ~n10406;
  assign n10525 = i_hbusreq1 & ~n10406;
  assign n10526 = ~n8389 & ~n10467;
  assign n10527 = ~n8389 & ~n10526;
  assign n10528 = i_hlock1 & ~n10527;
  assign n10529 = ~n8389 & ~n10474;
  assign n10530 = ~n8389 & ~n10529;
  assign n10531 = ~i_hlock1 & ~n10530;
  assign n10532 = ~n10528 & ~n10531;
  assign n10533 = ~i_hbusreq1 & ~n10532;
  assign n10534 = ~n10525 & ~n10533;
  assign n10535 = ~i_hbusreq3 & ~n10534;
  assign n10536 = ~n10524 & ~n10535;
  assign n10537 = ~i_hbusreq9 & ~n10536;
  assign n10538 = ~n10523 & ~n10537;
  assign n10539 = ~i_hbusreq4 & ~n10538;
  assign n10540 = ~n10522 & ~n10539;
  assign n10541 = ~i_hbusreq5 & ~n10540;
  assign n10542 = ~n10521 & ~n10541;
  assign n10543 = ~controllable_hmaster2 & ~n10542;
  assign n10544 = ~n10520 & ~n10543;
  assign n10545 = ~controllable_hmaster1 & ~n10544;
  assign n10546 = ~n10491 & ~n10545;
  assign n10547 = ~i_hbusreq6 & ~n10546;
  assign n10548 = ~n10461 & ~n10547;
  assign n10549 = controllable_hmaster0 & ~n10548;
  assign n10550 = i_hbusreq6 & ~n10444;
  assign n10551 = i_hbusreq5 & ~n10412;
  assign n10552 = i_hbusreq4 & ~n10412;
  assign n10553 = i_hbusreq9 & ~n10412;
  assign n10554 = i_hbusreq3 & ~n10412;
  assign n10555 = i_hbusreq1 & ~n10412;
  assign n10556 = n7928 & ~n8576;
  assign n10557 = ~i_hbusreq1 & ~n10556;
  assign n10558 = ~n10555 & ~n10557;
  assign n10559 = ~i_hbusreq3 & ~n10558;
  assign n10560 = ~n10554 & ~n10559;
  assign n10561 = ~i_hbusreq9 & ~n10560;
  assign n10562 = ~n10553 & ~n10561;
  assign n10563 = ~i_hbusreq4 & ~n10562;
  assign n10564 = ~n10552 & ~n10563;
  assign n10565 = ~i_hbusreq5 & ~n10564;
  assign n10566 = ~n10551 & ~n10565;
  assign n10567 = ~controllable_hmaster2 & ~n10566;
  assign n10568 = ~controllable_hmaster2 & ~n10567;
  assign n10569 = controllable_hmaster1 & ~n10568;
  assign n10570 = i_hbusreq5 & ~n10422;
  assign n10571 = i_hbusreq4 & ~n10422;
  assign n10572 = i_hbusreq9 & ~n10417;
  assign n10573 = ~n8426 & ~n10497;
  assign n10574 = ~n8426 & ~n10573;
  assign n10575 = ~i_hbusreq9 & ~n10574;
  assign n10576 = ~n10572 & ~n10575;
  assign n10577 = i_hlock4 & ~n10576;
  assign n10578 = i_hbusreq9 & ~n10420;
  assign n10579 = ~n8426 & ~n10509;
  assign n10580 = ~n8426 & ~n10579;
  assign n10581 = ~i_hbusreq9 & ~n10580;
  assign n10582 = ~n10578 & ~n10581;
  assign n10583 = ~i_hlock4 & ~n10582;
  assign n10584 = ~n10577 & ~n10583;
  assign n10585 = ~i_hbusreq4 & ~n10584;
  assign n10586 = ~n10571 & ~n10585;
  assign n10587 = ~i_hbusreq5 & ~n10586;
  assign n10588 = ~n10570 & ~n10587;
  assign n10589 = controllable_hmaster2 & ~n10588;
  assign n10590 = ~n10425 & ~n10589;
  assign n10591 = ~controllable_hmaster1 & ~n10590;
  assign n10592 = ~n10569 & ~n10591;
  assign n10593 = n8217 & ~n10592;
  assign n10594 = i_hbusreq5 & ~n10380;
  assign n10595 = ~i_hbusreq5 & ~n10501;
  assign n10596 = ~n10594 & ~n10595;
  assign n10597 = controllable_hmaster2 & ~n10596;
  assign n10598 = ~n10567 & ~n10597;
  assign n10599 = controllable_hmaster1 & ~n10598;
  assign n10600 = ~n10591 & ~n10599;
  assign n10601 = ~n8217 & ~n10600;
  assign n10602 = ~n10593 & ~n10601;
  assign n10603 = i_hlock6 & ~n10602;
  assign n10604 = i_hbusreq5 & ~n10384;
  assign n10605 = ~i_hbusreq5 & ~n10513;
  assign n10606 = ~n10604 & ~n10605;
  assign n10607 = controllable_hmaster2 & ~n10606;
  assign n10608 = ~n10567 & ~n10607;
  assign n10609 = controllable_hmaster1 & ~n10608;
  assign n10610 = ~n10591 & ~n10609;
  assign n10611 = ~n8217 & ~n10610;
  assign n10612 = ~n10593 & ~n10611;
  assign n10613 = ~i_hlock6 & ~n10612;
  assign n10614 = ~n10603 & ~n10613;
  assign n10615 = ~i_hbusreq6 & ~n10614;
  assign n10616 = ~n10550 & ~n10615;
  assign n10617 = ~controllable_hmaster0 & ~n10616;
  assign n10618 = ~n10549 & ~n10617;
  assign n10619 = ~i_hbusreq8 & ~n10618;
  assign n10620 = ~n10460 & ~n10619;
  assign n10621 = ~controllable_hmaster3 & ~n10620;
  assign n10622 = ~n10459 & ~n10621;
  assign n10623 = ~i_hbusreq7 & ~n10622;
  assign n10624 = ~n10449 & ~n10623;
  assign n10625 = n7924 & ~n10624;
  assign n10626 = ~n10375 & ~n10625;
  assign n10627 = n8214 & ~n10626;
  assign n10628 = n8214 & ~n10627;
  assign n10629 = n8202 & ~n10628;
  assign n10630 = ~n10332 & ~n10629;
  assign n10631 = n7728 & ~n10630;
  assign n10632 = ~n7743 & ~n10300;
  assign n10633 = i_hbusreq7 & ~n10632;
  assign n10634 = ~n7779 & ~n10314;
  assign n10635 = ~i_hbusreq7 & ~n10634;
  assign n10636 = ~n10633 & ~n10635;
  assign n10637 = n7924 & ~n10636;
  assign n10638 = ~n8337 & ~n10637;
  assign n10639 = ~n8214 & ~n10638;
  assign n10640 = ~n7743 & ~n10326;
  assign n10641 = i_hbusreq7 & ~n10640;
  assign n10642 = ~n7779 & ~n10326;
  assign n10643 = ~i_hbusreq7 & ~n10642;
  assign n10644 = ~n10641 & ~n10643;
  assign n10645 = n7924 & ~n10644;
  assign n10646 = ~n8337 & ~n10645;
  assign n10647 = n8214 & ~n10646;
  assign n10648 = ~n10639 & ~n10647;
  assign n10649 = ~n8202 & ~n10648;
  assign n10650 = n8214 & ~n8639;
  assign n10651 = ~n8336 & ~n10650;
  assign n10652 = n8202 & ~n10651;
  assign n10653 = ~n10649 & ~n10652;
  assign n10654 = ~n7728 & ~n10653;
  assign n10655 = ~n10631 & ~n10654;
  assign n10656 = ~n7723 & ~n10655;
  assign n10657 = ~n7723 & ~n10656;
  assign n10658 = ~n7714 & ~n10657;
  assign n10659 = ~n7714 & ~n10658;
  assign n10660 = n7705 & ~n10659;
  assign n10661 = n7723 & ~n10653;
  assign n10662 = n7920 & ~n10653;
  assign n10663 = ~n8640 & ~n10662;
  assign n10664 = ~n7723 & ~n10663;
  assign n10665 = ~n10661 & ~n10664;
  assign n10666 = n7714 & ~n10665;
  assign n10667 = ~n8646 & ~n10666;
  assign n10668 = ~n7705 & ~n10667;
  assign n10669 = ~n10660 & ~n10668;
  assign n10670 = ~n7808 & ~n10669;
  assign n10671 = ~n7920 & ~n10630;
  assign n10672 = ~controllable_hmaster2 & ~n9203;
  assign n10673 = ~controllable_hmaster1 & ~n10672;
  assign n10674 = ~controllable_hmaster1 & ~n10673;
  assign n10675 = controllable_hmaster0 & ~n10674;
  assign n10676 = controllable_hmaster0 & ~n10675;
  assign n10677 = ~controllable_hmaster3 & ~n10676;
  assign n10678 = ~controllable_hmaster3 & ~n10677;
  assign n10679 = i_hbusreq7 & ~n10678;
  assign n10680 = i_hbusreq8 & ~n10676;
  assign n10681 = i_hbusreq6 & ~n10674;
  assign n10682 = ~controllable_hmaster2 & ~n9660;
  assign n10683 = ~controllable_hmaster1 & ~n10682;
  assign n10684 = ~controllable_hmaster1 & ~n10683;
  assign n10685 = ~i_hbusreq6 & ~n10684;
  assign n10686 = ~n10681 & ~n10685;
  assign n10687 = controllable_hmaster0 & ~n10686;
  assign n10688 = controllable_hmaster0 & ~n10687;
  assign n10689 = ~i_hbusreq8 & ~n10688;
  assign n10690 = ~n10680 & ~n10689;
  assign n10691 = ~controllable_hmaster3 & ~n10690;
  assign n10692 = ~controllable_hmaster3 & ~n10691;
  assign n10693 = ~i_hbusreq7 & ~n10692;
  assign n10694 = ~n10679 & ~n10693;
  assign n10695 = ~n8214 & ~n10694;
  assign n10696 = ~controllable_hmaster2 & ~n9223;
  assign n10697 = ~controllable_hmaster1 & ~n10696;
  assign n10698 = ~controllable_hmaster1 & ~n10697;
  assign n10699 = ~controllable_hmaster0 & ~n10698;
  assign n10700 = ~controllable_hmaster0 & ~n10699;
  assign n10701 = ~controllable_hmaster3 & ~n10700;
  assign n10702 = ~controllable_hmaster3 & ~n10701;
  assign n10703 = i_hbusreq7 & ~n10702;
  assign n10704 = i_hbusreq8 & ~n10700;
  assign n10705 = i_hbusreq6 & ~n10698;
  assign n10706 = ~controllable_hmaster2 & ~n9704;
  assign n10707 = ~controllable_hmaster1 & ~n10706;
  assign n10708 = ~controllable_hmaster1 & ~n10707;
  assign n10709 = ~i_hbusreq6 & ~n10708;
  assign n10710 = ~n10705 & ~n10709;
  assign n10711 = ~controllable_hmaster0 & ~n10710;
  assign n10712 = ~controllable_hmaster0 & ~n10711;
  assign n10713 = ~i_hbusreq8 & ~n10712;
  assign n10714 = ~n10704 & ~n10713;
  assign n10715 = ~controllable_hmaster3 & ~n10714;
  assign n10716 = ~controllable_hmaster3 & ~n10715;
  assign n10717 = ~i_hbusreq7 & ~n10716;
  assign n10718 = ~n10703 & ~n10717;
  assign n10719 = n8214 & ~n10718;
  assign n10720 = ~n10695 & ~n10719;
  assign n10721 = ~n8202 & ~n10720;
  assign n10722 = n7924 & ~n9737;
  assign n10723 = n7924 & ~n10722;
  assign n10724 = ~n8214 & ~n10723;
  assign n10725 = i_hbusreq7 & ~n8987;
  assign n10726 = n7928 & ~n9588;
  assign n10727 = n7928 & ~n10726;
  assign n10728 = ~i_hbusreq1 & ~n10727;
  assign n10729 = ~n9011 & ~n10728;
  assign n10730 = ~i_hbusreq3 & ~n10729;
  assign n10731 = ~n9010 & ~n10730;
  assign n10732 = ~i_hbusreq9 & ~n10731;
  assign n10733 = ~n9009 & ~n10732;
  assign n10734 = ~i_hbusreq4 & ~n10733;
  assign n10735 = ~n9008 & ~n10734;
  assign n10736 = ~i_hbusreq5 & ~n10735;
  assign n10737 = ~n9007 & ~n10736;
  assign n10738 = controllable_hmaster1 & ~n10737;
  assign n10739 = controllable_hmaster2 & ~n10737;
  assign n10740 = n7928 & ~n8689;
  assign n10741 = ~i_hbusreq1 & ~n10740;
  assign n10742 = ~n9011 & ~n10741;
  assign n10743 = ~i_hbusreq3 & ~n10742;
  assign n10744 = ~n9010 & ~n10743;
  assign n10745 = ~i_hbusreq9 & ~n10744;
  assign n10746 = ~n9009 & ~n10745;
  assign n10747 = ~i_hbusreq4 & ~n10746;
  assign n10748 = ~n9008 & ~n10747;
  assign n10749 = ~i_hbusreq5 & ~n10748;
  assign n10750 = ~n9007 & ~n10749;
  assign n10751 = ~controllable_hmaster2 & ~n10750;
  assign n10752 = ~n10739 & ~n10751;
  assign n10753 = ~controllable_hmaster1 & ~n10752;
  assign n10754 = ~n10738 & ~n10753;
  assign n10755 = ~i_hbusreq6 & ~n10754;
  assign n10756 = ~n9036 & ~n10755;
  assign n10757 = ~i_hbusreq8 & ~n10756;
  assign n10758 = ~n9035 & ~n10757;
  assign n10759 = controllable_hmaster3 & ~n10758;
  assign n10760 = ~i_hbusreq6 & ~n10750;
  assign n10761 = ~n9036 & ~n10760;
  assign n10762 = controllable_hmaster0 & ~n10761;
  assign n10763 = controllable_hmaster1 & ~n10750;
  assign n10764 = controllable_hmaster2 & ~n10750;
  assign n10765 = n7928 & ~n9692;
  assign n10766 = ~i_hbusreq1 & ~n10765;
  assign n10767 = ~n9011 & ~n10766;
  assign n10768 = ~i_hbusreq3 & ~n10767;
  assign n10769 = ~n9010 & ~n10768;
  assign n10770 = ~i_hbusreq9 & ~n10769;
  assign n10771 = ~n9009 & ~n10770;
  assign n10772 = ~i_hbusreq4 & ~n10771;
  assign n10773 = ~n9008 & ~n10772;
  assign n10774 = ~i_hbusreq5 & ~n10773;
  assign n10775 = ~n9007 & ~n10774;
  assign n10776 = ~controllable_hmaster2 & ~n10775;
  assign n10777 = ~n10764 & ~n10776;
  assign n10778 = ~controllable_hmaster1 & ~n10777;
  assign n10779 = ~n10763 & ~n10778;
  assign n10780 = ~i_hbusreq6 & ~n10779;
  assign n10781 = ~n9036 & ~n10780;
  assign n10782 = ~controllable_hmaster0 & ~n10781;
  assign n10783 = ~n10762 & ~n10782;
  assign n10784 = ~i_hbusreq8 & ~n10783;
  assign n10785 = ~n9035 & ~n10784;
  assign n10786 = ~controllable_hmaster3 & ~n10785;
  assign n10787 = ~n10759 & ~n10786;
  assign n10788 = ~i_hbusreq7 & ~n10787;
  assign n10789 = ~n10725 & ~n10788;
  assign n10790 = n8214 & ~n10789;
  assign n10791 = ~n10724 & ~n10790;
  assign n10792 = n8202 & ~n10791;
  assign n10793 = ~n10721 & ~n10792;
  assign n10794 = n7920 & ~n10793;
  assign n10795 = ~n10671 & ~n10794;
  assign n10796 = n7728 & ~n10795;
  assign n10797 = ~n7920 & ~n10653;
  assign n10798 = ~n7743 & ~n10677;
  assign n10799 = i_hbusreq7 & ~n10798;
  assign n10800 = ~n7779 & ~n10691;
  assign n10801 = ~i_hbusreq7 & ~n10800;
  assign n10802 = ~n10799 & ~n10801;
  assign n10803 = ~n8214 & ~n10802;
  assign n10804 = ~n7743 & ~n10701;
  assign n10805 = i_hbusreq7 & ~n10804;
  assign n10806 = ~n7743 & ~n10715;
  assign n10807 = ~i_hbusreq7 & ~n10806;
  assign n10808 = ~n10805 & ~n10807;
  assign n10809 = n8214 & ~n10808;
  assign n10810 = ~n10803 & ~n10809;
  assign n10811 = ~n8202 & ~n10810;
  assign n10812 = ~n7744 & ~n7924;
  assign n10813 = ~n10722 & ~n10812;
  assign n10814 = ~n8214 & ~n10813;
  assign n10815 = n8214 & ~n9737;
  assign n10816 = ~n10814 & ~n10815;
  assign n10817 = n8202 & ~n10816;
  assign n10818 = ~n10811 & ~n10817;
  assign n10819 = n7920 & ~n10818;
  assign n10820 = ~n10797 & ~n10819;
  assign n10821 = ~n7728 & ~n10820;
  assign n10822 = ~n10796 & ~n10821;
  assign n10823 = ~n7723 & ~n10822;
  assign n10824 = ~n7723 & ~n10823;
  assign n10825 = ~n7714 & ~n10824;
  assign n10826 = ~n7714 & ~n10825;
  assign n10827 = n7705 & ~n10826;
  assign n10828 = ~n9203 & ~n10105;
  assign n10829 = ~controllable_hmaster1 & ~n10828;
  assign n10830 = ~n10053 & ~n10829;
  assign n10831 = controllable_hmaster0 & ~n10830;
  assign n10832 = ~n9099 & ~n10831;
  assign n10833 = ~controllable_hmaster3 & ~n10832;
  assign n10834 = ~n9093 & ~n10833;
  assign n10835 = i_hbusreq7 & ~n10834;
  assign n10836 = i_hbusreq8 & ~n10832;
  assign n10837 = i_hbusreq6 & ~n10830;
  assign n10838 = ~n9660 & ~n10116;
  assign n10839 = ~controllable_hmaster1 & ~n10838;
  assign n10840 = ~n10064 & ~n10839;
  assign n10841 = ~i_hbusreq6 & ~n10840;
  assign n10842 = ~n10837 & ~n10841;
  assign n10843 = controllable_hmaster0 & ~n10842;
  assign n10844 = ~n9127 & ~n10843;
  assign n10845 = ~i_hbusreq8 & ~n10844;
  assign n10846 = ~n10836 & ~n10845;
  assign n10847 = ~controllable_hmaster3 & ~n10846;
  assign n10848 = ~n9117 & ~n10847;
  assign n10849 = ~i_hbusreq7 & ~n10848;
  assign n10850 = ~n10835 & ~n10849;
  assign n10851 = ~n8214 & ~n10850;
  assign n10852 = ~n9223 & ~n10105;
  assign n10853 = ~controllable_hmaster1 & ~n10852;
  assign n10854 = ~n10053 & ~n10853;
  assign n10855 = ~controllable_hmaster0 & ~n10854;
  assign n10856 = ~n9152 & ~n10855;
  assign n10857 = ~controllable_hmaster3 & ~n10856;
  assign n10858 = ~n9093 & ~n10857;
  assign n10859 = i_hbusreq7 & ~n10858;
  assign n10860 = ~n9600 & ~n10751;
  assign n10861 = ~controllable_hmaster1 & ~n10860;
  assign n10862 = ~n9599 & ~n10861;
  assign n10863 = ~i_hbusreq6 & ~n10862;
  assign n10864 = ~n9006 & ~n10863;
  assign n10865 = ~i_hbusreq8 & ~n10864;
  assign n10866 = ~n9114 & ~n10865;
  assign n10867 = controllable_hmaster3 & ~n10866;
  assign n10868 = i_hbusreq8 & ~n10856;
  assign n10869 = i_hbusreq6 & ~n10854;
  assign n10870 = ~n9704 & ~n10764;
  assign n10871 = ~controllable_hmaster1 & ~n10870;
  assign n10872 = ~n10763 & ~n10871;
  assign n10873 = ~i_hbusreq6 & ~n10872;
  assign n10874 = ~n10869 & ~n10873;
  assign n10875 = ~controllable_hmaster0 & ~n10874;
  assign n10876 = ~n10762 & ~n10875;
  assign n10877 = ~i_hbusreq8 & ~n10876;
  assign n10878 = ~n10868 & ~n10877;
  assign n10879 = ~controllable_hmaster3 & ~n10878;
  assign n10880 = ~n10867 & ~n10879;
  assign n10881 = ~i_hbusreq7 & ~n10880;
  assign n10882 = ~n10859 & ~n10881;
  assign n10883 = n8214 & ~n10882;
  assign n10884 = ~n10851 & ~n10883;
  assign n10885 = ~n8202 & ~n10884;
  assign n10886 = n8202 & ~n9737;
  assign n10887 = ~n10885 & ~n10886;
  assign n10888 = n7920 & ~n10887;
  assign n10889 = ~n10797 & ~n10888;
  assign n10890 = n7728 & ~n10889;
  assign n10891 = ~n9339 & ~n9660;
  assign n10892 = ~controllable_hmaster1 & ~n10891;
  assign n10893 = ~n9332 & ~n10892;
  assign n10894 = ~i_hbusreq6 & ~n10893;
  assign n10895 = ~n9313 & ~n10894;
  assign n10896 = controllable_hmaster0 & ~n10895;
  assign n10897 = ~n9439 & ~n10896;
  assign n10898 = ~i_hbusreq8 & ~n10897;
  assign n10899 = ~n9312 & ~n10898;
  assign n10900 = ~controllable_hmaster3 & ~n10899;
  assign n10901 = ~n9517 & ~n10900;
  assign n10902 = i_hlock7 & ~n10901;
  assign n10903 = ~n9449 & ~n10892;
  assign n10904 = ~i_hbusreq6 & ~n10903;
  assign n10905 = ~n9447 & ~n10904;
  assign n10906 = controllable_hmaster0 & ~n10905;
  assign n10907 = ~n9439 & ~n10906;
  assign n10908 = ~i_hbusreq8 & ~n10907;
  assign n10909 = ~n9446 & ~n10908;
  assign n10910 = ~controllable_hmaster3 & ~n10909;
  assign n10911 = ~n9517 & ~n10910;
  assign n10912 = ~i_hlock7 & ~n10911;
  assign n10913 = ~n10902 & ~n10912;
  assign n10914 = ~i_hbusreq7 & ~n10913;
  assign n10915 = ~n9247 & ~n10914;
  assign n10916 = ~n8214 & ~n10915;
  assign n10917 = ~n10815 & ~n10916;
  assign n10918 = ~n8202 & ~n10917;
  assign n10919 = ~n10886 & ~n10918;
  assign n10920 = n7920 & ~n10919;
  assign n10921 = ~n10797 & ~n10920;
  assign n10922 = ~n7728 & ~n10921;
  assign n10923 = ~n10890 & ~n10922;
  assign n10924 = n7723 & ~n10923;
  assign n10925 = ~n7723 & ~n10921;
  assign n10926 = ~n10924 & ~n10925;
  assign n10927 = n7714 & ~n10926;
  assign n10928 = n7723 & ~n10921;
  assign n10929 = ~n8640 & ~n10920;
  assign n10930 = n7728 & ~n10929;
  assign n10931 = ~n9740 & ~n10930;
  assign n10932 = ~n7723 & ~n10931;
  assign n10933 = ~n10928 & ~n10932;
  assign n10934 = ~n7714 & ~n10933;
  assign n10935 = ~n10927 & ~n10934;
  assign n10936 = ~n7705 & ~n10935;
  assign n10937 = ~n10827 & ~n10936;
  assign n10938 = n7808 & ~n10937;
  assign n10939 = ~n10670 & ~n10938;
  assign n10940 = n8195 & ~n10939;
  assign n10941 = ~n10294 & ~n10940;
  assign n10942 = n8193 & ~n10941;
  assign n10943 = ~n9752 & ~n10942;
  assign n10944 = n8191 & ~n10943;
  assign n10945 = i_hlock9 & ~n8223;
  assign n10946 = ~i_hlock9 & ~n8237;
  assign n10947 = ~n10945 & ~n10946;
  assign n10948 = ~controllable_hmaster2 & ~n10947;
  assign n10949 = ~controllable_hmaster2 & ~n10948;
  assign n10950 = ~controllable_hmaster1 & ~n10949;
  assign n10951 = ~controllable_hmaster1 & ~n10950;
  assign n10952 = controllable_hmaster0 & ~n10951;
  assign n10953 = controllable_hmaster0 & ~n10952;
  assign n10954 = controllable_hmaster3 & ~n10953;
  assign n10955 = controllable_hmaster3 & ~n10954;
  assign n10956 = i_hbusreq7 & ~n10955;
  assign n10957 = i_hbusreq8 & ~n10953;
  assign n10958 = i_hbusreq6 & ~n10951;
  assign n10959 = i_hbusreq5 & ~n10947;
  assign n10960 = i_hbusreq4 & ~n10947;
  assign n10961 = i_hbusreq9 & ~n10947;
  assign n10962 = i_hlock9 & ~n8271;
  assign n10963 = ~i_hlock9 & ~n8303;
  assign n10964 = ~n10962 & ~n10963;
  assign n10965 = ~i_hbusreq9 & ~n10964;
  assign n10966 = ~n10961 & ~n10965;
  assign n10967 = ~i_hbusreq4 & ~n10966;
  assign n10968 = ~n10960 & ~n10967;
  assign n10969 = ~i_hbusreq5 & ~n10968;
  assign n10970 = ~n10959 & ~n10969;
  assign n10971 = ~controllable_hmaster2 & ~n10970;
  assign n10972 = ~controllable_hmaster2 & ~n10971;
  assign n10973 = ~controllable_hmaster1 & ~n10972;
  assign n10974 = ~controllable_hmaster1 & ~n10973;
  assign n10975 = ~i_hbusreq6 & ~n10974;
  assign n10976 = ~n10958 & ~n10975;
  assign n10977 = controllable_hmaster0 & ~n10976;
  assign n10978 = controllable_hmaster0 & ~n10977;
  assign n10979 = ~i_hbusreq8 & ~n10978;
  assign n10980 = ~n10957 & ~n10979;
  assign n10981 = controllable_hmaster3 & ~n10980;
  assign n10982 = controllable_hmaster3 & ~n10981;
  assign n10983 = ~i_hbusreq7 & ~n10982;
  assign n10984 = ~n10956 & ~n10983;
  assign n10985 = n7924 & ~n10984;
  assign n10986 = n7924 & ~n10985;
  assign n10987 = ~n8214 & ~n10986;
  assign n10988 = ~n8214 & ~n10987;
  assign n10989 = ~n8202 & ~n10988;
  assign n10990 = ~n8332 & ~n10989;
  assign n10991 = n7728 & ~n10990;
  assign n10992 = ~n7739 & ~n10948;
  assign n10993 = ~controllable_hmaster1 & ~n10992;
  assign n10994 = ~n7738 & ~n10993;
  assign n10995 = controllable_hmaster0 & ~n10994;
  assign n10996 = ~n8882 & ~n10995;
  assign n10997 = controllable_hmaster3 & ~n10996;
  assign n10998 = controllable_hmaster3 & ~n10997;
  assign n10999 = i_hbusreq7 & ~n10998;
  assign n11000 = i_hbusreq8 & ~n10996;
  assign n11001 = i_hbusreq6 & ~n10994;
  assign n11002 = ~n7771 & ~n10971;
  assign n11003 = ~controllable_hmaster1 & ~n11002;
  assign n11004 = ~n7770 & ~n11003;
  assign n11005 = ~i_hbusreq6 & ~n11004;
  assign n11006 = ~n11001 & ~n11005;
  assign n11007 = controllable_hmaster0 & ~n11006;
  assign n11008 = ~n8895 & ~n11007;
  assign n11009 = ~i_hbusreq8 & ~n11008;
  assign n11010 = ~n11000 & ~n11009;
  assign n11011 = controllable_hmaster3 & ~n11010;
  assign n11012 = controllable_hmaster3 & ~n11011;
  assign n11013 = ~i_hbusreq7 & ~n11012;
  assign n11014 = ~n10999 & ~n11013;
  assign n11015 = n7924 & ~n11014;
  assign n11016 = ~n8337 & ~n11015;
  assign n11017 = ~n8214 & ~n11016;
  assign n11018 = ~n7782 & n8214;
  assign n11019 = ~n11017 & ~n11018;
  assign n11020 = ~n8202 & ~n11019;
  assign n11021 = ~n8347 & ~n11020;
  assign n11022 = ~n7728 & ~n11021;
  assign n11023 = ~n10991 & ~n11022;
  assign n11024 = ~n7723 & ~n11023;
  assign n11025 = ~n7723 & ~n11024;
  assign n11026 = ~n7714 & ~n11025;
  assign n11027 = ~n7714 & ~n11026;
  assign n11028 = n7705 & ~n11027;
  assign n11029 = n7723 & ~n11021;
  assign n11030 = ~n8358 & ~n10948;
  assign n11031 = ~controllable_hmaster1 & ~n11030;
  assign n11032 = ~n8357 & ~n11031;
  assign n11033 = controllable_hmaster0 & ~n11032;
  assign n11034 = ~controllable_hmaster0 & ~n8361;
  assign n11035 = ~n11033 & ~n11034;
  assign n11036 = controllable_hmaster3 & ~n11035;
  assign n11037 = ~n8463 & ~n11036;
  assign n11038 = i_hbusreq7 & ~n11037;
  assign n11039 = i_hbusreq8 & ~n11035;
  assign n11040 = i_hbusreq6 & ~n11032;
  assign n11041 = ~n8484 & ~n10971;
  assign n11042 = ~controllable_hmaster1 & ~n11041;
  assign n11043 = ~n8483 & ~n11042;
  assign n11044 = ~i_hbusreq6 & ~n11043;
  assign n11045 = ~n11040 & ~n11044;
  assign n11046 = controllable_hmaster0 & ~n11045;
  assign n11047 = ~controllable_hmaster0 & ~n8489;
  assign n11048 = ~n11046 & ~n11047;
  assign n11049 = ~i_hbusreq8 & ~n11048;
  assign n11050 = ~n11039 & ~n11049;
  assign n11051 = controllable_hmaster3 & ~n11050;
  assign n11052 = ~n8634 & ~n11051;
  assign n11053 = ~i_hbusreq7 & ~n11052;
  assign n11054 = ~n11038 & ~n11053;
  assign n11055 = n7924 & ~n11054;
  assign n11056 = ~n8337 & ~n11055;
  assign n11057 = ~n7920 & ~n11056;
  assign n11058 = n7920 & ~n11021;
  assign n11059 = ~n11057 & ~n11058;
  assign n11060 = ~n7723 & ~n11059;
  assign n11061 = ~n11029 & ~n11060;
  assign n11062 = n7714 & ~n11061;
  assign n11063 = ~n7714 & ~n11056;
  assign n11064 = ~n11062 & ~n11063;
  assign n11065 = ~n7705 & ~n11064;
  assign n11066 = ~n11028 & ~n11065;
  assign n11067 = ~n7808 & ~n11066;
  assign n11068 = ~n7920 & ~n10990;
  assign n11069 = ~n8874 & ~n11068;
  assign n11070 = n7728 & ~n11069;
  assign n11071 = ~n7920 & ~n11021;
  assign n11072 = ~n8974 & ~n11071;
  assign n11073 = ~n7728 & ~n11072;
  assign n11074 = ~n11070 & ~n11073;
  assign n11075 = ~n7723 & ~n11074;
  assign n11076 = ~n7723 & ~n11075;
  assign n11077 = ~n7714 & ~n11076;
  assign n11078 = ~n7714 & ~n11077;
  assign n11079 = n7705 & ~n11078;
  assign n11080 = ~n9181 & ~n11071;
  assign n11081 = n7728 & ~n11080;
  assign n11082 = ~n9577 & ~n11071;
  assign n11083 = ~n7728 & ~n11082;
  assign n11084 = ~n11081 & ~n11083;
  assign n11085 = n7723 & ~n11084;
  assign n11086 = ~n7723 & ~n11082;
  assign n11087 = ~n11085 & ~n11086;
  assign n11088 = n7714 & ~n11087;
  assign n11089 = n7723 & ~n11082;
  assign n11090 = ~n9577 & ~n11057;
  assign n11091 = n7728 & ~n11090;
  assign n11092 = ~n9738 & ~n11057;
  assign n11093 = ~n7728 & ~n11092;
  assign n11094 = ~n11091 & ~n11093;
  assign n11095 = ~n7723 & ~n11094;
  assign n11096 = ~n11089 & ~n11095;
  assign n11097 = ~n7714 & ~n11096;
  assign n11098 = ~n11088 & ~n11097;
  assign n11099 = ~n7705 & ~n11098;
  assign n11100 = ~n11079 & ~n11099;
  assign n11101 = n7808 & ~n11100;
  assign n11102 = ~n11067 & ~n11101;
  assign n11103 = n8195 & ~n11102;
  assign n11104 = ~n8196 & ~n11103;
  assign n11105 = ~n8193 & ~n11104;
  assign n11106 = ~n9900 & ~n11057;
  assign n11107 = ~n7723 & ~n11106;
  assign n11108 = ~n9899 & ~n11107;
  assign n11109 = n7714 & ~n11108;
  assign n11110 = ~n11063 & ~n11109;
  assign n11111 = ~n7705 & ~n11110;
  assign n11112 = ~n9898 & ~n11111;
  assign n11113 = ~n7808 & ~n11112;
  assign n11114 = ~n10274 & ~n11057;
  assign n11115 = n7728 & ~n11114;
  assign n11116 = ~n11093 & ~n11115;
  assign n11117 = ~n7723 & ~n11116;
  assign n11118 = ~n10282 & ~n11117;
  assign n11119 = ~n7714 & ~n11118;
  assign n11120 = ~n10281 & ~n11119;
  assign n11121 = ~n7705 & ~n11120;
  assign n11122 = ~n10052 & ~n11121;
  assign n11123 = n7808 & ~n11122;
  assign n11124 = ~n11113 & ~n11123;
  assign n11125 = ~n8195 & ~n11124;
  assign n11126 = i_hlock9 & ~n10380;
  assign n11127 = ~i_hlock9 & ~n10384;
  assign n11128 = ~n11126 & ~n11127;
  assign n11129 = ~controllable_hmaster2 & ~n11128;
  assign n11130 = ~n10105 & ~n11129;
  assign n11131 = ~controllable_hmaster1 & ~n11130;
  assign n11132 = ~n10053 & ~n11131;
  assign n11133 = controllable_hmaster0 & ~n11132;
  assign n11134 = ~controllable_hmaster0 & ~n10378;
  assign n11135 = ~n11133 & ~n11134;
  assign n11136 = controllable_hmaster3 & ~n11135;
  assign n11137 = ~n10447 & ~n11136;
  assign n11138 = i_hbusreq7 & ~n11137;
  assign n11139 = i_hbusreq8 & ~n11135;
  assign n11140 = i_hbusreq6 & ~n11132;
  assign n11141 = i_hbusreq5 & ~n11128;
  assign n11142 = i_hbusreq4 & ~n11128;
  assign n11143 = i_hbusreq9 & ~n11128;
  assign n11144 = i_hlock9 & ~n10497;
  assign n11145 = ~i_hlock9 & ~n10509;
  assign n11146 = ~n11144 & ~n11145;
  assign n11147 = ~i_hbusreq9 & ~n11146;
  assign n11148 = ~n11143 & ~n11147;
  assign n11149 = ~i_hbusreq4 & ~n11148;
  assign n11150 = ~n11142 & ~n11149;
  assign n11151 = ~i_hbusreq5 & ~n11150;
  assign n11152 = ~n11141 & ~n11151;
  assign n11153 = ~controllable_hmaster2 & ~n11152;
  assign n11154 = ~n10116 & ~n11153;
  assign n11155 = ~controllable_hmaster1 & ~n11154;
  assign n11156 = ~n10064 & ~n11155;
  assign n11157 = ~i_hbusreq6 & ~n11156;
  assign n11158 = ~n11140 & ~n11157;
  assign n11159 = controllable_hmaster0 & ~n11158;
  assign n11160 = ~controllable_hmaster0 & ~n10456;
  assign n11161 = ~n11159 & ~n11160;
  assign n11162 = ~i_hbusreq8 & ~n11161;
  assign n11163 = ~n11139 & ~n11162;
  assign n11164 = controllable_hmaster3 & ~n11163;
  assign n11165 = ~n10621 & ~n11164;
  assign n11166 = ~i_hbusreq7 & ~n11165;
  assign n11167 = ~n11138 & ~n11166;
  assign n11168 = n7924 & ~n11167;
  assign n11169 = ~n10375 & ~n11168;
  assign n11170 = n8214 & ~n11169;
  assign n11171 = n8214 & ~n11170;
  assign n11172 = n8202 & ~n11171;
  assign n11173 = ~n10332 & ~n11172;
  assign n11174 = n7728 & ~n11173;
  assign n11175 = n8214 & ~n11056;
  assign n11176 = ~n8336 & ~n11175;
  assign n11177 = n8202 & ~n11176;
  assign n11178 = ~n10649 & ~n11177;
  assign n11179 = ~n7728 & ~n11178;
  assign n11180 = ~n11174 & ~n11179;
  assign n11181 = ~n7723 & ~n11180;
  assign n11182 = ~n7723 & ~n11181;
  assign n11183 = ~n7714 & ~n11182;
  assign n11184 = ~n7714 & ~n11183;
  assign n11185 = n7705 & ~n11184;
  assign n11186 = n7723 & ~n11178;
  assign n11187 = n7920 & ~n11178;
  assign n11188 = ~n11057 & ~n11187;
  assign n11189 = ~n7723 & ~n11188;
  assign n11190 = ~n11186 & ~n11189;
  assign n11191 = n7714 & ~n11190;
  assign n11192 = ~n11063 & ~n11191;
  assign n11193 = ~n7705 & ~n11192;
  assign n11194 = ~n11185 & ~n11193;
  assign n11195 = ~n7808 & ~n11194;
  assign n11196 = ~n7920 & ~n11173;
  assign n11197 = ~n10794 & ~n11196;
  assign n11198 = n7728 & ~n11197;
  assign n11199 = ~n7920 & ~n11178;
  assign n11200 = ~n10819 & ~n11199;
  assign n11201 = ~n7728 & ~n11200;
  assign n11202 = ~n11198 & ~n11201;
  assign n11203 = ~n7723 & ~n11202;
  assign n11204 = ~n7723 & ~n11203;
  assign n11205 = ~n7714 & ~n11204;
  assign n11206 = ~n7714 & ~n11205;
  assign n11207 = n7705 & ~n11206;
  assign n11208 = ~n10888 & ~n11199;
  assign n11209 = n7728 & ~n11208;
  assign n11210 = ~n10920 & ~n11199;
  assign n11211 = ~n7728 & ~n11210;
  assign n11212 = ~n11209 & ~n11211;
  assign n11213 = n7723 & ~n11212;
  assign n11214 = ~n7723 & ~n11210;
  assign n11215 = ~n11213 & ~n11214;
  assign n11216 = n7714 & ~n11215;
  assign n11217 = n7723 & ~n11210;
  assign n11218 = ~n10920 & ~n11057;
  assign n11219 = n7728 & ~n11218;
  assign n11220 = ~n11093 & ~n11219;
  assign n11221 = ~n7723 & ~n11220;
  assign n11222 = ~n11217 & ~n11221;
  assign n11223 = ~n7714 & ~n11222;
  assign n11224 = ~n11216 & ~n11223;
  assign n11225 = ~n7705 & ~n11224;
  assign n11226 = ~n11207 & ~n11225;
  assign n11227 = n7808 & ~n11226;
  assign n11228 = ~n11195 & ~n11227;
  assign n11229 = n8195 & ~n11228;
  assign n11230 = ~n11125 & ~n11229;
  assign n11231 = n8193 & ~n11230;
  assign n11232 = ~n11105 & ~n11231;
  assign n11233 = ~n8191 & ~n11232;
  assign n11234 = ~n10944 & ~n11233;
  assign n11235 = n8188 & ~n11234;
  assign n11236 = ~controllable_hmaster2 & ~n8223;
  assign n11237 = ~controllable_hmaster2 & ~n11236;
  assign n11238 = ~controllable_hmaster1 & ~n11237;
  assign n11239 = ~controllable_hmaster1 & ~n11238;
  assign n11240 = ~controllable_hmaster0 & ~n11239;
  assign n11241 = ~controllable_hmaster0 & ~n11240;
  assign n11242 = i_hlock8 & ~n11241;
  assign n11243 = ~controllable_hmaster2 & ~n8237;
  assign n11244 = ~controllable_hmaster2 & ~n11243;
  assign n11245 = ~controllable_hmaster1 & ~n11244;
  assign n11246 = ~controllable_hmaster1 & ~n11245;
  assign n11247 = ~controllable_hmaster0 & ~n11246;
  assign n11248 = ~controllable_hmaster0 & ~n11247;
  assign n11249 = ~i_hlock8 & ~n11248;
  assign n11250 = ~n11242 & ~n11249;
  assign n11251 = controllable_hmaster3 & ~n11250;
  assign n11252 = controllable_hmaster3 & ~n11251;
  assign n11253 = i_hbusreq7 & ~n11252;
  assign n11254 = i_hbusreq8 & ~n11250;
  assign n11255 = i_hbusreq6 & ~n11239;
  assign n11256 = ~controllable_hmaster2 & ~n8277;
  assign n11257 = ~controllable_hmaster2 & ~n11256;
  assign n11258 = ~controllable_hmaster1 & ~n11257;
  assign n11259 = ~controllable_hmaster1 & ~n11258;
  assign n11260 = ~i_hbusreq6 & ~n11259;
  assign n11261 = ~n11255 & ~n11260;
  assign n11262 = ~controllable_hmaster0 & ~n11261;
  assign n11263 = ~controllable_hmaster0 & ~n11262;
  assign n11264 = i_hlock8 & ~n11263;
  assign n11265 = i_hbusreq6 & ~n11246;
  assign n11266 = ~controllable_hmaster2 & ~n8309;
  assign n11267 = ~controllable_hmaster2 & ~n11266;
  assign n11268 = ~controllable_hmaster1 & ~n11267;
  assign n11269 = ~controllable_hmaster1 & ~n11268;
  assign n11270 = ~i_hbusreq6 & ~n11269;
  assign n11271 = ~n11265 & ~n11270;
  assign n11272 = ~controllable_hmaster0 & ~n11271;
  assign n11273 = ~controllable_hmaster0 & ~n11272;
  assign n11274 = ~i_hlock8 & ~n11273;
  assign n11275 = ~n11264 & ~n11274;
  assign n11276 = ~i_hbusreq8 & ~n11275;
  assign n11277 = ~n11254 & ~n11276;
  assign n11278 = controllable_hmaster3 & ~n11277;
  assign n11279 = controllable_hmaster3 & ~n11278;
  assign n11280 = ~i_hbusreq7 & ~n11279;
  assign n11281 = ~n11253 & ~n11280;
  assign n11282 = n7924 & ~n11281;
  assign n11283 = n7924 & ~n11282;
  assign n11284 = n8214 & ~n11283;
  assign n11285 = n8214 & ~n11284;
  assign n11286 = ~n8202 & ~n11285;
  assign n11287 = ~n8332 & ~n11286;
  assign n11288 = n7728 & ~n11287;
  assign n11289 = ~n7739 & ~n11236;
  assign n11290 = ~controllable_hmaster1 & ~n11289;
  assign n11291 = ~n7738 & ~n11290;
  assign n11292 = ~controllable_hmaster0 & ~n11291;
  assign n11293 = ~n8904 & ~n11292;
  assign n11294 = i_hlock8 & ~n11293;
  assign n11295 = ~n7739 & ~n11243;
  assign n11296 = ~controllable_hmaster1 & ~n11295;
  assign n11297 = ~n7738 & ~n11296;
  assign n11298 = ~controllable_hmaster0 & ~n11297;
  assign n11299 = ~n8904 & ~n11298;
  assign n11300 = ~i_hlock8 & ~n11299;
  assign n11301 = ~n11294 & ~n11300;
  assign n11302 = controllable_hmaster3 & ~n11301;
  assign n11303 = controllable_hmaster3 & ~n11302;
  assign n11304 = i_hbusreq7 & ~n11303;
  assign n11305 = i_hbusreq8 & ~n11301;
  assign n11306 = i_hbusreq6 & ~n11291;
  assign n11307 = ~n7771 & ~n11256;
  assign n11308 = ~controllable_hmaster1 & ~n11307;
  assign n11309 = ~n7770 & ~n11308;
  assign n11310 = ~i_hbusreq6 & ~n11309;
  assign n11311 = ~n11306 & ~n11310;
  assign n11312 = ~controllable_hmaster0 & ~n11311;
  assign n11313 = ~n8922 & ~n11312;
  assign n11314 = i_hlock8 & ~n11313;
  assign n11315 = i_hbusreq6 & ~n11297;
  assign n11316 = ~n7771 & ~n11266;
  assign n11317 = ~controllable_hmaster1 & ~n11316;
  assign n11318 = ~n7770 & ~n11317;
  assign n11319 = ~i_hbusreq6 & ~n11318;
  assign n11320 = ~n11315 & ~n11319;
  assign n11321 = ~controllable_hmaster0 & ~n11320;
  assign n11322 = ~n8922 & ~n11321;
  assign n11323 = ~i_hlock8 & ~n11322;
  assign n11324 = ~n11314 & ~n11323;
  assign n11325 = ~i_hbusreq8 & ~n11324;
  assign n11326 = ~n11305 & ~n11325;
  assign n11327 = controllable_hmaster3 & ~n11326;
  assign n11328 = controllable_hmaster3 & ~n11327;
  assign n11329 = ~i_hbusreq7 & ~n11328;
  assign n11330 = ~n11304 & ~n11329;
  assign n11331 = n7924 & ~n11330;
  assign n11332 = ~n8337 & ~n11331;
  assign n11333 = n8214 & ~n11332;
  assign n11334 = ~n8336 & ~n11333;
  assign n11335 = ~n8202 & ~n11334;
  assign n11336 = ~n8347 & ~n11335;
  assign n11337 = ~n7728 & ~n11336;
  assign n11338 = ~n11288 & ~n11337;
  assign n11339 = ~n7723 & ~n11338;
  assign n11340 = ~n7723 & ~n11339;
  assign n11341 = ~n7714 & ~n11340;
  assign n11342 = ~n7714 & ~n11341;
  assign n11343 = n7705 & ~n11342;
  assign n11344 = n7723 & ~n11336;
  assign n11345 = controllable_hmaster0 & ~n8361;
  assign n11346 = ~n8358 & ~n11236;
  assign n11347 = ~controllable_hmaster1 & ~n11346;
  assign n11348 = ~n8357 & ~n11347;
  assign n11349 = ~controllable_hmaster0 & ~n11348;
  assign n11350 = ~n11345 & ~n11349;
  assign n11351 = i_hlock8 & ~n11350;
  assign n11352 = ~n8358 & ~n11243;
  assign n11353 = ~controllable_hmaster1 & ~n11352;
  assign n11354 = ~n8357 & ~n11353;
  assign n11355 = ~controllable_hmaster0 & ~n11354;
  assign n11356 = ~n11345 & ~n11355;
  assign n11357 = ~i_hlock8 & ~n11356;
  assign n11358 = ~n11351 & ~n11357;
  assign n11359 = controllable_hmaster3 & ~n11358;
  assign n11360 = ~n8463 & ~n11359;
  assign n11361 = i_hbusreq7 & ~n11360;
  assign n11362 = i_hbusreq8 & ~n11358;
  assign n11363 = controllable_hmaster0 & ~n8489;
  assign n11364 = i_hbusreq6 & ~n11348;
  assign n11365 = ~n8484 & ~n11256;
  assign n11366 = ~controllable_hmaster1 & ~n11365;
  assign n11367 = ~n8483 & ~n11366;
  assign n11368 = ~i_hbusreq6 & ~n11367;
  assign n11369 = ~n11364 & ~n11368;
  assign n11370 = ~controllable_hmaster0 & ~n11369;
  assign n11371 = ~n11363 & ~n11370;
  assign n11372 = i_hlock8 & ~n11371;
  assign n11373 = i_hbusreq6 & ~n11354;
  assign n11374 = ~n8484 & ~n11266;
  assign n11375 = ~controllable_hmaster1 & ~n11374;
  assign n11376 = ~n8483 & ~n11375;
  assign n11377 = ~i_hbusreq6 & ~n11376;
  assign n11378 = ~n11373 & ~n11377;
  assign n11379 = ~controllable_hmaster0 & ~n11378;
  assign n11380 = ~n11363 & ~n11379;
  assign n11381 = ~i_hlock8 & ~n11380;
  assign n11382 = ~n11372 & ~n11381;
  assign n11383 = ~i_hbusreq8 & ~n11382;
  assign n11384 = ~n11362 & ~n11383;
  assign n11385 = controllable_hmaster3 & ~n11384;
  assign n11386 = ~n8634 & ~n11385;
  assign n11387 = ~i_hbusreq7 & ~n11386;
  assign n11388 = ~n11361 & ~n11387;
  assign n11389 = n7924 & ~n11388;
  assign n11390 = ~n8337 & ~n11389;
  assign n11391 = ~n7920 & ~n11390;
  assign n11392 = n7920 & ~n11336;
  assign n11393 = ~n11391 & ~n11392;
  assign n11394 = ~n7723 & ~n11393;
  assign n11395 = ~n11344 & ~n11394;
  assign n11396 = n7714 & ~n11395;
  assign n11397 = ~n7714 & ~n11390;
  assign n11398 = ~n11396 & ~n11397;
  assign n11399 = ~n7705 & ~n11398;
  assign n11400 = ~n11343 & ~n11399;
  assign n11401 = ~n7808 & ~n11400;
  assign n11402 = ~n7920 & ~n11287;
  assign n11403 = ~n8874 & ~n11402;
  assign n11404 = n7728 & ~n11403;
  assign n11405 = ~n7920 & ~n11336;
  assign n11406 = ~n8974 & ~n11405;
  assign n11407 = ~n7728 & ~n11406;
  assign n11408 = ~n11404 & ~n11407;
  assign n11409 = ~n7723 & ~n11408;
  assign n11410 = ~n7723 & ~n11409;
  assign n11411 = ~n7714 & ~n11410;
  assign n11412 = ~n7714 & ~n11411;
  assign n11413 = n7705 & ~n11412;
  assign n11414 = ~n9181 & ~n11405;
  assign n11415 = n7728 & ~n11414;
  assign n11416 = ~n9577 & ~n11405;
  assign n11417 = ~n7728 & ~n11416;
  assign n11418 = ~n11415 & ~n11417;
  assign n11419 = n7723 & ~n11418;
  assign n11420 = ~n7723 & ~n11416;
  assign n11421 = ~n11419 & ~n11420;
  assign n11422 = n7714 & ~n11421;
  assign n11423 = n7723 & ~n11416;
  assign n11424 = ~n9577 & ~n11391;
  assign n11425 = n7728 & ~n11424;
  assign n11426 = ~n9738 & ~n11391;
  assign n11427 = ~n7728 & ~n11426;
  assign n11428 = ~n11425 & ~n11427;
  assign n11429 = ~n7723 & ~n11428;
  assign n11430 = ~n11423 & ~n11429;
  assign n11431 = ~n7714 & ~n11430;
  assign n11432 = ~n11422 & ~n11431;
  assign n11433 = ~n7705 & ~n11432;
  assign n11434 = ~n11413 & ~n11433;
  assign n11435 = n7808 & ~n11434;
  assign n11436 = ~n11401 & ~n11435;
  assign n11437 = n8195 & ~n11436;
  assign n11438 = ~n8196 & ~n11437;
  assign n11439 = ~n8193 & ~n11438;
  assign n11440 = ~n9900 & ~n11391;
  assign n11441 = ~n7723 & ~n11440;
  assign n11442 = ~n9899 & ~n11441;
  assign n11443 = n7714 & ~n11442;
  assign n11444 = ~n11397 & ~n11443;
  assign n11445 = ~n7705 & ~n11444;
  assign n11446 = ~n9898 & ~n11445;
  assign n11447 = ~n7808 & ~n11446;
  assign n11448 = ~n10274 & ~n11391;
  assign n11449 = n7728 & ~n11448;
  assign n11450 = ~n11427 & ~n11449;
  assign n11451 = ~n7723 & ~n11450;
  assign n11452 = ~n10282 & ~n11451;
  assign n11453 = ~n7714 & ~n11452;
  assign n11454 = ~n10281 & ~n11453;
  assign n11455 = ~n7705 & ~n11454;
  assign n11456 = ~n10052 & ~n11455;
  assign n11457 = n7808 & ~n11456;
  assign n11458 = ~n11447 & ~n11457;
  assign n11459 = ~n8195 & ~n11458;
  assign n11460 = controllable_hmaster0 & ~n10378;
  assign n11461 = ~controllable_hmaster2 & ~n10380;
  assign n11462 = ~n10105 & ~n11461;
  assign n11463 = ~controllable_hmaster1 & ~n11462;
  assign n11464 = ~n10053 & ~n11463;
  assign n11465 = ~controllable_hmaster0 & ~n11464;
  assign n11466 = ~n11460 & ~n11465;
  assign n11467 = i_hlock8 & ~n11466;
  assign n11468 = ~controllable_hmaster2 & ~n10384;
  assign n11469 = ~n10105 & ~n11468;
  assign n11470 = ~controllable_hmaster1 & ~n11469;
  assign n11471 = ~n10053 & ~n11470;
  assign n11472 = ~controllable_hmaster0 & ~n11471;
  assign n11473 = ~n11460 & ~n11472;
  assign n11474 = ~i_hlock8 & ~n11473;
  assign n11475 = ~n11467 & ~n11474;
  assign n11476 = controllable_hmaster3 & ~n11475;
  assign n11477 = ~n10447 & ~n11476;
  assign n11478 = i_hbusreq7 & ~n11477;
  assign n11479 = i_hbusreq8 & ~n11475;
  assign n11480 = controllable_hmaster0 & ~n10456;
  assign n11481 = i_hbusreq6 & ~n11464;
  assign n11482 = ~controllable_hmaster2 & ~n10596;
  assign n11483 = ~n10116 & ~n11482;
  assign n11484 = ~controllable_hmaster1 & ~n11483;
  assign n11485 = ~n10064 & ~n11484;
  assign n11486 = ~i_hbusreq6 & ~n11485;
  assign n11487 = ~n11481 & ~n11486;
  assign n11488 = ~controllable_hmaster0 & ~n11487;
  assign n11489 = ~n11480 & ~n11488;
  assign n11490 = i_hlock8 & ~n11489;
  assign n11491 = i_hbusreq6 & ~n11471;
  assign n11492 = ~controllable_hmaster2 & ~n10606;
  assign n11493 = ~n10116 & ~n11492;
  assign n11494 = ~controllable_hmaster1 & ~n11493;
  assign n11495 = ~n10064 & ~n11494;
  assign n11496 = ~i_hbusreq6 & ~n11495;
  assign n11497 = ~n11491 & ~n11496;
  assign n11498 = ~controllable_hmaster0 & ~n11497;
  assign n11499 = ~n11480 & ~n11498;
  assign n11500 = ~i_hlock8 & ~n11499;
  assign n11501 = ~n11490 & ~n11500;
  assign n11502 = ~i_hbusreq8 & ~n11501;
  assign n11503 = ~n11479 & ~n11502;
  assign n11504 = controllable_hmaster3 & ~n11503;
  assign n11505 = ~n10621 & ~n11504;
  assign n11506 = ~i_hbusreq7 & ~n11505;
  assign n11507 = ~n11478 & ~n11506;
  assign n11508 = n7924 & ~n11507;
  assign n11509 = ~n10375 & ~n11508;
  assign n11510 = n8214 & ~n11509;
  assign n11511 = n8214 & ~n11510;
  assign n11512 = n8202 & ~n11511;
  assign n11513 = ~n10332 & ~n11512;
  assign n11514 = n7728 & ~n11513;
  assign n11515 = n8214 & ~n11390;
  assign n11516 = ~n8336 & ~n11515;
  assign n11517 = n8202 & ~n11516;
  assign n11518 = ~n10649 & ~n11517;
  assign n11519 = ~n7728 & ~n11518;
  assign n11520 = ~n11514 & ~n11519;
  assign n11521 = ~n7723 & ~n11520;
  assign n11522 = ~n7723 & ~n11521;
  assign n11523 = ~n7714 & ~n11522;
  assign n11524 = ~n7714 & ~n11523;
  assign n11525 = n7705 & ~n11524;
  assign n11526 = n7723 & ~n11518;
  assign n11527 = n7920 & ~n11518;
  assign n11528 = ~n11391 & ~n11527;
  assign n11529 = ~n7723 & ~n11528;
  assign n11530 = ~n11526 & ~n11529;
  assign n11531 = n7714 & ~n11530;
  assign n11532 = ~n11397 & ~n11531;
  assign n11533 = ~n7705 & ~n11532;
  assign n11534 = ~n11525 & ~n11533;
  assign n11535 = ~n7808 & ~n11534;
  assign n11536 = ~n7920 & ~n11513;
  assign n11537 = ~n10794 & ~n11536;
  assign n11538 = n7728 & ~n11537;
  assign n11539 = ~n7920 & ~n11518;
  assign n11540 = ~n10819 & ~n11539;
  assign n11541 = ~n7728 & ~n11540;
  assign n11542 = ~n11538 & ~n11541;
  assign n11543 = ~n7723 & ~n11542;
  assign n11544 = ~n7723 & ~n11543;
  assign n11545 = ~n7714 & ~n11544;
  assign n11546 = ~n7714 & ~n11545;
  assign n11547 = n7705 & ~n11546;
  assign n11548 = ~n10888 & ~n11539;
  assign n11549 = n7728 & ~n11548;
  assign n11550 = ~n10920 & ~n11539;
  assign n11551 = ~n7728 & ~n11550;
  assign n11552 = ~n11549 & ~n11551;
  assign n11553 = n7723 & ~n11552;
  assign n11554 = ~n7723 & ~n11550;
  assign n11555 = ~n11553 & ~n11554;
  assign n11556 = n7714 & ~n11555;
  assign n11557 = n7723 & ~n11550;
  assign n11558 = ~n10920 & ~n11391;
  assign n11559 = n7728 & ~n11558;
  assign n11560 = ~n11427 & ~n11559;
  assign n11561 = ~n7723 & ~n11560;
  assign n11562 = ~n11557 & ~n11561;
  assign n11563 = ~n7714 & ~n11562;
  assign n11564 = ~n11556 & ~n11563;
  assign n11565 = ~n7705 & ~n11564;
  assign n11566 = ~n11547 & ~n11565;
  assign n11567 = n7808 & ~n11566;
  assign n11568 = ~n11535 & ~n11567;
  assign n11569 = n8195 & ~n11568;
  assign n11570 = ~n11459 & ~n11569;
  assign n11571 = n8193 & ~n11570;
  assign n11572 = ~n11439 & ~n11571;
  assign n11573 = n8191 & ~n11572;
  assign n11574 = ~n10987 & ~n11284;
  assign n11575 = ~n8202 & ~n11574;
  assign n11576 = ~n8332 & ~n11575;
  assign n11577 = n7728 & ~n11576;
  assign n11578 = ~n11017 & ~n11333;
  assign n11579 = ~n8202 & ~n11578;
  assign n11580 = ~n8347 & ~n11579;
  assign n11581 = ~n7728 & ~n11580;
  assign n11582 = ~n11577 & ~n11581;
  assign n11583 = ~n7723 & ~n11582;
  assign n11584 = ~n7723 & ~n11583;
  assign n11585 = ~n7714 & ~n11584;
  assign n11586 = ~n7714 & ~n11585;
  assign n11587 = n7705 & ~n11586;
  assign n11588 = n7723 & ~n11580;
  assign n11589 = ~n11033 & ~n11349;
  assign n11590 = i_hlock8 & ~n11589;
  assign n11591 = ~n11033 & ~n11355;
  assign n11592 = ~i_hlock8 & ~n11591;
  assign n11593 = ~n11590 & ~n11592;
  assign n11594 = controllable_hmaster3 & ~n11593;
  assign n11595 = ~n8463 & ~n11594;
  assign n11596 = i_hbusreq7 & ~n11595;
  assign n11597 = i_hbusreq8 & ~n11593;
  assign n11598 = ~n11046 & ~n11370;
  assign n11599 = i_hlock8 & ~n11598;
  assign n11600 = ~n11046 & ~n11379;
  assign n11601 = ~i_hlock8 & ~n11600;
  assign n11602 = ~n11599 & ~n11601;
  assign n11603 = ~i_hbusreq8 & ~n11602;
  assign n11604 = ~n11597 & ~n11603;
  assign n11605 = controllable_hmaster3 & ~n11604;
  assign n11606 = ~n8634 & ~n11605;
  assign n11607 = ~i_hbusreq7 & ~n11606;
  assign n11608 = ~n11596 & ~n11607;
  assign n11609 = n7924 & ~n11608;
  assign n11610 = ~n8337 & ~n11609;
  assign n11611 = ~n7920 & ~n11610;
  assign n11612 = n7920 & ~n11580;
  assign n11613 = ~n11611 & ~n11612;
  assign n11614 = ~n7723 & ~n11613;
  assign n11615 = ~n11588 & ~n11614;
  assign n11616 = n7714 & ~n11615;
  assign n11617 = ~n7714 & ~n11610;
  assign n11618 = ~n11616 & ~n11617;
  assign n11619 = ~n7705 & ~n11618;
  assign n11620 = ~n11587 & ~n11619;
  assign n11621 = ~n7808 & ~n11620;
  assign n11622 = ~n7920 & ~n11576;
  assign n11623 = ~n8874 & ~n11622;
  assign n11624 = n7728 & ~n11623;
  assign n11625 = ~n7920 & ~n11580;
  assign n11626 = ~n8974 & ~n11625;
  assign n11627 = ~n7728 & ~n11626;
  assign n11628 = ~n11624 & ~n11627;
  assign n11629 = ~n7723 & ~n11628;
  assign n11630 = ~n7723 & ~n11629;
  assign n11631 = ~n7714 & ~n11630;
  assign n11632 = ~n7714 & ~n11631;
  assign n11633 = n7705 & ~n11632;
  assign n11634 = ~n9181 & ~n11625;
  assign n11635 = n7728 & ~n11634;
  assign n11636 = ~n9577 & ~n11625;
  assign n11637 = ~n7728 & ~n11636;
  assign n11638 = ~n11635 & ~n11637;
  assign n11639 = n7723 & ~n11638;
  assign n11640 = ~n7723 & ~n11636;
  assign n11641 = ~n11639 & ~n11640;
  assign n11642 = n7714 & ~n11641;
  assign n11643 = n7723 & ~n11636;
  assign n11644 = ~n9577 & ~n11611;
  assign n11645 = n7728 & ~n11644;
  assign n11646 = ~n9738 & ~n11611;
  assign n11647 = ~n7728 & ~n11646;
  assign n11648 = ~n11645 & ~n11647;
  assign n11649 = ~n7723 & ~n11648;
  assign n11650 = ~n11643 & ~n11649;
  assign n11651 = ~n7714 & ~n11650;
  assign n11652 = ~n11642 & ~n11651;
  assign n11653 = ~n7705 & ~n11652;
  assign n11654 = ~n11633 & ~n11653;
  assign n11655 = n7808 & ~n11654;
  assign n11656 = ~n11621 & ~n11655;
  assign n11657 = n8195 & ~n11656;
  assign n11658 = ~n8196 & ~n11657;
  assign n11659 = ~n8193 & ~n11658;
  assign n11660 = ~n9900 & ~n11611;
  assign n11661 = ~n7723 & ~n11660;
  assign n11662 = ~n9899 & ~n11661;
  assign n11663 = n7714 & ~n11662;
  assign n11664 = ~n11617 & ~n11663;
  assign n11665 = ~n7705 & ~n11664;
  assign n11666 = ~n9898 & ~n11665;
  assign n11667 = ~n7808 & ~n11666;
  assign n11668 = ~n10274 & ~n11611;
  assign n11669 = n7728 & ~n11668;
  assign n11670 = ~n11647 & ~n11669;
  assign n11671 = ~n7723 & ~n11670;
  assign n11672 = ~n10282 & ~n11671;
  assign n11673 = ~n7714 & ~n11672;
  assign n11674 = ~n10281 & ~n11673;
  assign n11675 = ~n7705 & ~n11674;
  assign n11676 = ~n10052 & ~n11675;
  assign n11677 = n7808 & ~n11676;
  assign n11678 = ~n11667 & ~n11677;
  assign n11679 = ~n8195 & ~n11678;
  assign n11680 = ~n11133 & ~n11465;
  assign n11681 = i_hlock8 & ~n11680;
  assign n11682 = ~n11133 & ~n11472;
  assign n11683 = ~i_hlock8 & ~n11682;
  assign n11684 = ~n11681 & ~n11683;
  assign n11685 = controllable_hmaster3 & ~n11684;
  assign n11686 = ~n10447 & ~n11685;
  assign n11687 = i_hbusreq7 & ~n11686;
  assign n11688 = i_hbusreq8 & ~n11684;
  assign n11689 = ~n11159 & ~n11488;
  assign n11690 = i_hlock8 & ~n11689;
  assign n11691 = ~n11159 & ~n11498;
  assign n11692 = ~i_hlock8 & ~n11691;
  assign n11693 = ~n11690 & ~n11692;
  assign n11694 = ~i_hbusreq8 & ~n11693;
  assign n11695 = ~n11688 & ~n11694;
  assign n11696 = controllable_hmaster3 & ~n11695;
  assign n11697 = ~n10621 & ~n11696;
  assign n11698 = ~i_hbusreq7 & ~n11697;
  assign n11699 = ~n11687 & ~n11698;
  assign n11700 = n7924 & ~n11699;
  assign n11701 = ~n10375 & ~n11700;
  assign n11702 = n8214 & ~n11701;
  assign n11703 = n8214 & ~n11702;
  assign n11704 = n8202 & ~n11703;
  assign n11705 = ~n10332 & ~n11704;
  assign n11706 = n7728 & ~n11705;
  assign n11707 = n8214 & ~n11610;
  assign n11708 = ~n8336 & ~n11707;
  assign n11709 = n8202 & ~n11708;
  assign n11710 = ~n10649 & ~n11709;
  assign n11711 = ~n7728 & ~n11710;
  assign n11712 = ~n11706 & ~n11711;
  assign n11713 = ~n7723 & ~n11712;
  assign n11714 = ~n7723 & ~n11713;
  assign n11715 = ~n7714 & ~n11714;
  assign n11716 = ~n7714 & ~n11715;
  assign n11717 = n7705 & ~n11716;
  assign n11718 = n7723 & ~n11710;
  assign n11719 = n7920 & ~n11710;
  assign n11720 = ~n11611 & ~n11719;
  assign n11721 = ~n7723 & ~n11720;
  assign n11722 = ~n11718 & ~n11721;
  assign n11723 = n7714 & ~n11722;
  assign n11724 = ~n11617 & ~n11723;
  assign n11725 = ~n7705 & ~n11724;
  assign n11726 = ~n11717 & ~n11725;
  assign n11727 = ~n7808 & ~n11726;
  assign n11728 = ~n7920 & ~n11705;
  assign n11729 = ~n10794 & ~n11728;
  assign n11730 = n7728 & ~n11729;
  assign n11731 = ~n7920 & ~n11710;
  assign n11732 = ~n10819 & ~n11731;
  assign n11733 = ~n7728 & ~n11732;
  assign n11734 = ~n11730 & ~n11733;
  assign n11735 = ~n7723 & ~n11734;
  assign n11736 = ~n7723 & ~n11735;
  assign n11737 = ~n7714 & ~n11736;
  assign n11738 = ~n7714 & ~n11737;
  assign n11739 = n7705 & ~n11738;
  assign n11740 = ~n10888 & ~n11731;
  assign n11741 = n7728 & ~n11740;
  assign n11742 = ~n10920 & ~n11731;
  assign n11743 = ~n7728 & ~n11742;
  assign n11744 = ~n11741 & ~n11743;
  assign n11745 = n7723 & ~n11744;
  assign n11746 = ~n7723 & ~n11742;
  assign n11747 = ~n11745 & ~n11746;
  assign n11748 = n7714 & ~n11747;
  assign n11749 = n7723 & ~n11742;
  assign n11750 = ~n10920 & ~n11611;
  assign n11751 = n7728 & ~n11750;
  assign n11752 = ~n11647 & ~n11751;
  assign n11753 = ~n7723 & ~n11752;
  assign n11754 = ~n11749 & ~n11753;
  assign n11755 = ~n7714 & ~n11754;
  assign n11756 = ~n11748 & ~n11755;
  assign n11757 = ~n7705 & ~n11756;
  assign n11758 = ~n11739 & ~n11757;
  assign n11759 = n7808 & ~n11758;
  assign n11760 = ~n11727 & ~n11759;
  assign n11761 = n8195 & ~n11760;
  assign n11762 = ~n11679 & ~n11761;
  assign n11763 = n8193 & ~n11762;
  assign n11764 = ~n11659 & ~n11763;
  assign n11765 = ~n8191 & ~n11764;
  assign n11766 = ~n11573 & ~n11765;
  assign n11767 = ~n8188 & ~n11766;
  assign n11768 = ~n11235 & ~n11767;
  assign n11769 = n8185 & ~n11768;
  assign n11770 = controllable_hmaster0 & ~n8227;
  assign n11771 = controllable_hmaster0 & ~n11770;
  assign n11772 = ~controllable_hmaster3 & ~n11771;
  assign n11773 = ~controllable_hmaster3 & ~n11772;
  assign n11774 = i_hlock7 & ~n11773;
  assign n11775 = controllable_hmaster0 & ~n8241;
  assign n11776 = controllable_hmaster0 & ~n11775;
  assign n11777 = ~controllable_hmaster3 & ~n11776;
  assign n11778 = ~controllable_hmaster3 & ~n11777;
  assign n11779 = ~i_hlock7 & ~n11778;
  assign n11780 = ~n11774 & ~n11779;
  assign n11781 = i_hbusreq7 & ~n11780;
  assign n11782 = i_hbusreq8 & ~n11771;
  assign n11783 = i_hbusreq6 & ~n8227;
  assign n11784 = ~i_hbusreq6 & ~n8281;
  assign n11785 = ~n11783 & ~n11784;
  assign n11786 = controllable_hmaster0 & ~n11785;
  assign n11787 = controllable_hmaster0 & ~n11786;
  assign n11788 = ~i_hbusreq8 & ~n11787;
  assign n11789 = ~n11782 & ~n11788;
  assign n11790 = ~controllable_hmaster3 & ~n11789;
  assign n11791 = ~controllable_hmaster3 & ~n11790;
  assign n11792 = i_hlock7 & ~n11791;
  assign n11793 = i_hbusreq8 & ~n11776;
  assign n11794 = i_hbusreq6 & ~n8241;
  assign n11795 = ~i_hbusreq6 & ~n8313;
  assign n11796 = ~n11794 & ~n11795;
  assign n11797 = controllable_hmaster0 & ~n11796;
  assign n11798 = controllable_hmaster0 & ~n11797;
  assign n11799 = ~i_hbusreq8 & ~n11798;
  assign n11800 = ~n11793 & ~n11799;
  assign n11801 = ~controllable_hmaster3 & ~n11800;
  assign n11802 = ~controllable_hmaster3 & ~n11801;
  assign n11803 = ~i_hlock7 & ~n11802;
  assign n11804 = ~n11792 & ~n11803;
  assign n11805 = ~i_hbusreq7 & ~n11804;
  assign n11806 = ~n11781 & ~n11805;
  assign n11807 = n7924 & ~n11806;
  assign n11808 = n7924 & ~n11807;
  assign n11809 = ~n8214 & ~n11808;
  assign n11810 = ~n8330 & ~n11809;
  assign n11811 = n8202 & ~n11810;
  assign n11812 = n8202 & ~n11811;
  assign n11813 = n7728 & ~n11812;
  assign n11814 = ~n7743 & ~n11772;
  assign n11815 = i_hlock7 & ~n11814;
  assign n11816 = ~n7743 & ~n11777;
  assign n11817 = ~i_hlock7 & ~n11816;
  assign n11818 = ~n11815 & ~n11817;
  assign n11819 = i_hbusreq7 & ~n11818;
  assign n11820 = ~n7779 & ~n11790;
  assign n11821 = i_hlock7 & ~n11820;
  assign n11822 = ~n7779 & ~n11801;
  assign n11823 = ~i_hlock7 & ~n11822;
  assign n11824 = ~n11821 & ~n11823;
  assign n11825 = ~i_hbusreq7 & ~n11824;
  assign n11826 = ~n11819 & ~n11825;
  assign n11827 = n7924 & ~n11826;
  assign n11828 = ~n8337 & ~n11827;
  assign n11829 = ~n8214 & ~n11828;
  assign n11830 = ~n8345 & ~n11829;
  assign n11831 = n8202 & ~n11830;
  assign n11832 = ~n8335 & ~n11831;
  assign n11833 = ~n7728 & ~n11832;
  assign n11834 = ~n11813 & ~n11833;
  assign n11835 = ~n7723 & ~n11834;
  assign n11836 = ~n7723 & ~n11835;
  assign n11837 = ~n7714 & ~n11836;
  assign n11838 = ~n7714 & ~n11837;
  assign n11839 = n7705 & ~n11838;
  assign n11840 = n7723 & ~n11832;
  assign n11841 = ~n8224 & ~n8373;
  assign n11842 = controllable_hmaster1 & ~n11841;
  assign n11843 = ~n8399 & ~n11842;
  assign n11844 = controllable_hmaster0 & ~n11843;
  assign n11845 = ~n8461 & ~n11844;
  assign n11846 = ~controllable_hmaster3 & ~n11845;
  assign n11847 = ~n8362 & ~n11846;
  assign n11848 = i_hlock7 & ~n11847;
  assign n11849 = ~n8238 & ~n8373;
  assign n11850 = controllable_hmaster1 & ~n11849;
  assign n11851 = ~n8399 & ~n11850;
  assign n11852 = controllable_hmaster0 & ~n11851;
  assign n11853 = ~n8461 & ~n11852;
  assign n11854 = ~controllable_hmaster3 & ~n11853;
  assign n11855 = ~n8362 & ~n11854;
  assign n11856 = ~i_hlock7 & ~n11855;
  assign n11857 = ~n11848 & ~n11856;
  assign n11858 = i_hbusreq7 & ~n11857;
  assign n11859 = i_hbusreq8 & ~n11845;
  assign n11860 = i_hbusreq6 & ~n11843;
  assign n11861 = ~n8278 & ~n8514;
  assign n11862 = controllable_hmaster1 & ~n11861;
  assign n11863 = ~n8552 & ~n11862;
  assign n11864 = ~i_hbusreq6 & ~n11863;
  assign n11865 = ~n11860 & ~n11864;
  assign n11866 = controllable_hmaster0 & ~n11865;
  assign n11867 = ~n8630 & ~n11866;
  assign n11868 = ~i_hbusreq8 & ~n11867;
  assign n11869 = ~n11859 & ~n11868;
  assign n11870 = ~controllable_hmaster3 & ~n11869;
  assign n11871 = ~n8492 & ~n11870;
  assign n11872 = i_hlock7 & ~n11871;
  assign n11873 = i_hbusreq8 & ~n11853;
  assign n11874 = i_hbusreq6 & ~n11851;
  assign n11875 = ~n8310 & ~n8514;
  assign n11876 = controllable_hmaster1 & ~n11875;
  assign n11877 = ~n8552 & ~n11876;
  assign n11878 = ~i_hbusreq6 & ~n11877;
  assign n11879 = ~n11874 & ~n11878;
  assign n11880 = controllable_hmaster0 & ~n11879;
  assign n11881 = ~n8630 & ~n11880;
  assign n11882 = ~i_hbusreq8 & ~n11881;
  assign n11883 = ~n11873 & ~n11882;
  assign n11884 = ~controllable_hmaster3 & ~n11883;
  assign n11885 = ~n8492 & ~n11884;
  assign n11886 = ~i_hlock7 & ~n11885;
  assign n11887 = ~n11872 & ~n11886;
  assign n11888 = ~i_hbusreq7 & ~n11887;
  assign n11889 = ~n11858 & ~n11888;
  assign n11890 = n7924 & ~n11889;
  assign n11891 = ~n8337 & ~n11890;
  assign n11892 = ~n7920 & ~n11891;
  assign n11893 = n7920 & ~n11832;
  assign n11894 = ~n11892 & ~n11893;
  assign n11895 = ~n7723 & ~n11894;
  assign n11896 = ~n11840 & ~n11895;
  assign n11897 = n7714 & ~n11896;
  assign n11898 = ~n7714 & ~n11891;
  assign n11899 = ~n11897 & ~n11898;
  assign n11900 = ~n7705 & ~n11899;
  assign n11901 = ~n11839 & ~n11900;
  assign n11902 = ~n7808 & ~n11901;
  assign n11903 = ~n7920 & ~n11812;
  assign n11904 = ~n8874 & ~n11903;
  assign n11905 = n7728 & ~n11904;
  assign n11906 = ~n7920 & ~n11832;
  assign n11907 = ~n8974 & ~n11906;
  assign n11908 = ~n7728 & ~n11907;
  assign n11909 = ~n11905 & ~n11908;
  assign n11910 = ~n7723 & ~n11909;
  assign n11911 = ~n7723 & ~n11910;
  assign n11912 = ~n7714 & ~n11911;
  assign n11913 = ~n7714 & ~n11912;
  assign n11914 = n7705 & ~n11913;
  assign n11915 = ~n9181 & ~n11906;
  assign n11916 = n7728 & ~n11915;
  assign n11917 = ~n9577 & ~n11906;
  assign n11918 = ~n7728 & ~n11917;
  assign n11919 = ~n11916 & ~n11918;
  assign n11920 = n7723 & ~n11919;
  assign n11921 = ~n7723 & ~n11917;
  assign n11922 = ~n11920 & ~n11921;
  assign n11923 = n7714 & ~n11922;
  assign n11924 = n7723 & ~n11917;
  assign n11925 = ~n9577 & ~n11892;
  assign n11926 = n7728 & ~n11925;
  assign n11927 = ~n9738 & ~n11892;
  assign n11928 = ~n7728 & ~n11927;
  assign n11929 = ~n11926 & ~n11928;
  assign n11930 = ~n7723 & ~n11929;
  assign n11931 = ~n11924 & ~n11930;
  assign n11932 = ~n7714 & ~n11931;
  assign n11933 = ~n11923 & ~n11932;
  assign n11934 = ~n7705 & ~n11933;
  assign n11935 = ~n11914 & ~n11934;
  assign n11936 = n7808 & ~n11935;
  assign n11937 = ~n11902 & ~n11936;
  assign n11938 = n8195 & ~n11937;
  assign n11939 = ~n8196 & ~n11938;
  assign n11940 = ~n8193 & ~n11939;
  assign n11941 = ~n9900 & ~n11892;
  assign n11942 = ~n7723 & ~n11941;
  assign n11943 = ~n9899 & ~n11942;
  assign n11944 = n7714 & ~n11943;
  assign n11945 = ~n11898 & ~n11944;
  assign n11946 = ~n7705 & ~n11945;
  assign n11947 = ~n9898 & ~n11946;
  assign n11948 = ~n7808 & ~n11947;
  assign n11949 = ~n10274 & ~n11892;
  assign n11950 = n7728 & ~n11949;
  assign n11951 = ~n11928 & ~n11950;
  assign n11952 = ~n7723 & ~n11951;
  assign n11953 = ~n10282 & ~n11952;
  assign n11954 = ~n7714 & ~n11953;
  assign n11955 = ~n10281 & ~n11954;
  assign n11956 = ~n7705 & ~n11955;
  assign n11957 = ~n10052 & ~n11956;
  assign n11958 = n7808 & ~n11957;
  assign n11959 = ~n11948 & ~n11958;
  assign n11960 = ~n8195 & ~n11959;
  assign n11961 = ~n10389 & ~n10430;
  assign n11962 = controllable_hmaster1 & ~n11961;
  assign n11963 = ~n10409 & ~n11962;
  assign n11964 = controllable_hmaster0 & ~n11963;
  assign n11965 = ~n10445 & ~n11964;
  assign n11966 = ~controllable_hmaster3 & ~n11965;
  assign n11967 = ~n10379 & ~n11966;
  assign n11968 = i_hlock7 & ~n11967;
  assign n11969 = ~n10389 & ~n10437;
  assign n11970 = controllable_hmaster1 & ~n11969;
  assign n11971 = ~n10409 & ~n11970;
  assign n11972 = controllable_hmaster0 & ~n11971;
  assign n11973 = ~n10445 & ~n11972;
  assign n11974 = ~controllable_hmaster3 & ~n11973;
  assign n11975 = ~n10379 & ~n11974;
  assign n11976 = ~i_hlock7 & ~n11975;
  assign n11977 = ~n11968 & ~n11976;
  assign n11978 = i_hbusreq7 & ~n11977;
  assign n11979 = i_hbusreq8 & ~n11965;
  assign n11980 = i_hbusreq6 & ~n11963;
  assign n11981 = ~n10489 & ~n10597;
  assign n11982 = controllable_hmaster1 & ~n11981;
  assign n11983 = ~n10545 & ~n11982;
  assign n11984 = ~i_hbusreq6 & ~n11983;
  assign n11985 = ~n11980 & ~n11984;
  assign n11986 = controllable_hmaster0 & ~n11985;
  assign n11987 = ~n10617 & ~n11986;
  assign n11988 = ~i_hbusreq8 & ~n11987;
  assign n11989 = ~n11979 & ~n11988;
  assign n11990 = ~controllable_hmaster3 & ~n11989;
  assign n11991 = ~n10459 & ~n11990;
  assign n11992 = i_hlock7 & ~n11991;
  assign n11993 = i_hbusreq8 & ~n11973;
  assign n11994 = i_hbusreq6 & ~n11971;
  assign n11995 = ~n10489 & ~n10607;
  assign n11996 = controllable_hmaster1 & ~n11995;
  assign n11997 = ~n10545 & ~n11996;
  assign n11998 = ~i_hbusreq6 & ~n11997;
  assign n11999 = ~n11994 & ~n11998;
  assign n12000 = controllable_hmaster0 & ~n11999;
  assign n12001 = ~n10617 & ~n12000;
  assign n12002 = ~i_hbusreq8 & ~n12001;
  assign n12003 = ~n11993 & ~n12002;
  assign n12004 = ~controllable_hmaster3 & ~n12003;
  assign n12005 = ~n10459 & ~n12004;
  assign n12006 = ~i_hlock7 & ~n12005;
  assign n12007 = ~n11992 & ~n12006;
  assign n12008 = ~i_hbusreq7 & ~n12007;
  assign n12009 = ~n11978 & ~n12008;
  assign n12010 = n7924 & ~n12009;
  assign n12011 = ~n10375 & ~n12010;
  assign n12012 = n8214 & ~n12011;
  assign n12013 = n8214 & ~n12012;
  assign n12014 = n8202 & ~n12013;
  assign n12015 = ~n10332 & ~n12014;
  assign n12016 = n7728 & ~n12015;
  assign n12017 = n8214 & ~n11891;
  assign n12018 = ~n8336 & ~n12017;
  assign n12019 = n8202 & ~n12018;
  assign n12020 = ~n10649 & ~n12019;
  assign n12021 = ~n7728 & ~n12020;
  assign n12022 = ~n12016 & ~n12021;
  assign n12023 = ~n7723 & ~n12022;
  assign n12024 = ~n7723 & ~n12023;
  assign n12025 = ~n7714 & ~n12024;
  assign n12026 = ~n7714 & ~n12025;
  assign n12027 = n7705 & ~n12026;
  assign n12028 = n7723 & ~n12020;
  assign n12029 = n7920 & ~n12020;
  assign n12030 = ~n11892 & ~n12029;
  assign n12031 = ~n7723 & ~n12030;
  assign n12032 = ~n12028 & ~n12031;
  assign n12033 = n7714 & ~n12032;
  assign n12034 = ~n11898 & ~n12033;
  assign n12035 = ~n7705 & ~n12034;
  assign n12036 = ~n12027 & ~n12035;
  assign n12037 = ~n7808 & ~n12036;
  assign n12038 = ~n7920 & ~n12015;
  assign n12039 = ~n10794 & ~n12038;
  assign n12040 = n7728 & ~n12039;
  assign n12041 = ~n7920 & ~n12020;
  assign n12042 = ~n10819 & ~n12041;
  assign n12043 = ~n7728 & ~n12042;
  assign n12044 = ~n12040 & ~n12043;
  assign n12045 = ~n7723 & ~n12044;
  assign n12046 = ~n7723 & ~n12045;
  assign n12047 = ~n7714 & ~n12046;
  assign n12048 = ~n7714 & ~n12047;
  assign n12049 = n7705 & ~n12048;
  assign n12050 = ~n10888 & ~n12041;
  assign n12051 = n7728 & ~n12050;
  assign n12052 = ~n10920 & ~n12041;
  assign n12053 = ~n7728 & ~n12052;
  assign n12054 = ~n12051 & ~n12053;
  assign n12055 = n7723 & ~n12054;
  assign n12056 = ~n7723 & ~n12052;
  assign n12057 = ~n12055 & ~n12056;
  assign n12058 = n7714 & ~n12057;
  assign n12059 = n7723 & ~n12052;
  assign n12060 = ~n10920 & ~n11892;
  assign n12061 = n7728 & ~n12060;
  assign n12062 = ~n11928 & ~n12061;
  assign n12063 = ~n7723 & ~n12062;
  assign n12064 = ~n12059 & ~n12063;
  assign n12065 = ~n7714 & ~n12064;
  assign n12066 = ~n12058 & ~n12065;
  assign n12067 = ~n7705 & ~n12066;
  assign n12068 = ~n12049 & ~n12067;
  assign n12069 = n7808 & ~n12068;
  assign n12070 = ~n12037 & ~n12069;
  assign n12071 = n8195 & ~n12070;
  assign n12072 = ~n11960 & ~n12071;
  assign n12073 = n8193 & ~n12072;
  assign n12074 = ~n11940 & ~n12073;
  assign n12075 = n8191 & ~n12074;
  assign n12076 = ~n10989 & ~n11811;
  assign n12077 = n7728 & ~n12076;
  assign n12078 = ~n11020 & ~n11831;
  assign n12079 = ~n7728 & ~n12078;
  assign n12080 = ~n12077 & ~n12079;
  assign n12081 = ~n7723 & ~n12080;
  assign n12082 = ~n7723 & ~n12081;
  assign n12083 = ~n7714 & ~n12082;
  assign n12084 = ~n7714 & ~n12083;
  assign n12085 = n7705 & ~n12084;
  assign n12086 = n7723 & ~n12078;
  assign n12087 = ~n11036 & ~n11846;
  assign n12088 = i_hlock7 & ~n12087;
  assign n12089 = ~n11036 & ~n11854;
  assign n12090 = ~i_hlock7 & ~n12089;
  assign n12091 = ~n12088 & ~n12090;
  assign n12092 = i_hbusreq7 & ~n12091;
  assign n12093 = ~n11051 & ~n11870;
  assign n12094 = i_hlock7 & ~n12093;
  assign n12095 = ~n11051 & ~n11884;
  assign n12096 = ~i_hlock7 & ~n12095;
  assign n12097 = ~n12094 & ~n12096;
  assign n12098 = ~i_hbusreq7 & ~n12097;
  assign n12099 = ~n12092 & ~n12098;
  assign n12100 = n7924 & ~n12099;
  assign n12101 = ~n8337 & ~n12100;
  assign n12102 = ~n7920 & ~n12101;
  assign n12103 = n7920 & ~n12078;
  assign n12104 = ~n12102 & ~n12103;
  assign n12105 = ~n7723 & ~n12104;
  assign n12106 = ~n12086 & ~n12105;
  assign n12107 = n7714 & ~n12106;
  assign n12108 = ~n7714 & ~n12101;
  assign n12109 = ~n12107 & ~n12108;
  assign n12110 = ~n7705 & ~n12109;
  assign n12111 = ~n12085 & ~n12110;
  assign n12112 = ~n7808 & ~n12111;
  assign n12113 = ~n7920 & ~n12076;
  assign n12114 = ~n8874 & ~n12113;
  assign n12115 = n7728 & ~n12114;
  assign n12116 = ~n7920 & ~n12078;
  assign n12117 = ~n8974 & ~n12116;
  assign n12118 = ~n7728 & ~n12117;
  assign n12119 = ~n12115 & ~n12118;
  assign n12120 = ~n7723 & ~n12119;
  assign n12121 = ~n7723 & ~n12120;
  assign n12122 = ~n7714 & ~n12121;
  assign n12123 = ~n7714 & ~n12122;
  assign n12124 = n7705 & ~n12123;
  assign n12125 = ~n9181 & ~n12116;
  assign n12126 = n7728 & ~n12125;
  assign n12127 = ~n9577 & ~n12116;
  assign n12128 = ~n7728 & ~n12127;
  assign n12129 = ~n12126 & ~n12128;
  assign n12130 = n7723 & ~n12129;
  assign n12131 = ~n7723 & ~n12127;
  assign n12132 = ~n12130 & ~n12131;
  assign n12133 = n7714 & ~n12132;
  assign n12134 = n7723 & ~n12127;
  assign n12135 = ~n9577 & ~n12102;
  assign n12136 = n7728 & ~n12135;
  assign n12137 = ~n9738 & ~n12102;
  assign n12138 = ~n7728 & ~n12137;
  assign n12139 = ~n12136 & ~n12138;
  assign n12140 = ~n7723 & ~n12139;
  assign n12141 = ~n12134 & ~n12140;
  assign n12142 = ~n7714 & ~n12141;
  assign n12143 = ~n12133 & ~n12142;
  assign n12144 = ~n7705 & ~n12143;
  assign n12145 = ~n12124 & ~n12144;
  assign n12146 = n7808 & ~n12145;
  assign n12147 = ~n12112 & ~n12146;
  assign n12148 = n8195 & ~n12147;
  assign n12149 = ~n8196 & ~n12148;
  assign n12150 = ~n8193 & ~n12149;
  assign n12151 = ~n9900 & ~n12102;
  assign n12152 = ~n7723 & ~n12151;
  assign n12153 = ~n9899 & ~n12152;
  assign n12154 = n7714 & ~n12153;
  assign n12155 = ~n12108 & ~n12154;
  assign n12156 = ~n7705 & ~n12155;
  assign n12157 = ~n9898 & ~n12156;
  assign n12158 = ~n7808 & ~n12157;
  assign n12159 = ~n10274 & ~n12102;
  assign n12160 = n7728 & ~n12159;
  assign n12161 = ~n12138 & ~n12160;
  assign n12162 = ~n7723 & ~n12161;
  assign n12163 = ~n10282 & ~n12162;
  assign n12164 = ~n7714 & ~n12163;
  assign n12165 = ~n10281 & ~n12164;
  assign n12166 = ~n7705 & ~n12165;
  assign n12167 = ~n10052 & ~n12166;
  assign n12168 = n7808 & ~n12167;
  assign n12169 = ~n12158 & ~n12168;
  assign n12170 = ~n8195 & ~n12169;
  assign n12171 = ~n11136 & ~n11966;
  assign n12172 = i_hlock7 & ~n12171;
  assign n12173 = ~n11136 & ~n11974;
  assign n12174 = ~i_hlock7 & ~n12173;
  assign n12175 = ~n12172 & ~n12174;
  assign n12176 = i_hbusreq7 & ~n12175;
  assign n12177 = ~n11164 & ~n11990;
  assign n12178 = i_hlock7 & ~n12177;
  assign n12179 = ~n11164 & ~n12004;
  assign n12180 = ~i_hlock7 & ~n12179;
  assign n12181 = ~n12178 & ~n12180;
  assign n12182 = ~i_hbusreq7 & ~n12181;
  assign n12183 = ~n12176 & ~n12182;
  assign n12184 = n7924 & ~n12183;
  assign n12185 = ~n10375 & ~n12184;
  assign n12186 = n8214 & ~n12185;
  assign n12187 = n8214 & ~n12186;
  assign n12188 = n8202 & ~n12187;
  assign n12189 = ~n10332 & ~n12188;
  assign n12190 = n7728 & ~n12189;
  assign n12191 = n8214 & ~n12101;
  assign n12192 = ~n8336 & ~n12191;
  assign n12193 = n8202 & ~n12192;
  assign n12194 = ~n10649 & ~n12193;
  assign n12195 = ~n7728 & ~n12194;
  assign n12196 = ~n12190 & ~n12195;
  assign n12197 = ~n7723 & ~n12196;
  assign n12198 = ~n7723 & ~n12197;
  assign n12199 = ~n7714 & ~n12198;
  assign n12200 = ~n7714 & ~n12199;
  assign n12201 = n7705 & ~n12200;
  assign n12202 = n7723 & ~n12194;
  assign n12203 = n7920 & ~n12194;
  assign n12204 = ~n12102 & ~n12203;
  assign n12205 = ~n7723 & ~n12204;
  assign n12206 = ~n12202 & ~n12205;
  assign n12207 = n7714 & ~n12206;
  assign n12208 = ~n12108 & ~n12207;
  assign n12209 = ~n7705 & ~n12208;
  assign n12210 = ~n12201 & ~n12209;
  assign n12211 = ~n7808 & ~n12210;
  assign n12212 = ~n7920 & ~n12189;
  assign n12213 = ~n10794 & ~n12212;
  assign n12214 = n7728 & ~n12213;
  assign n12215 = ~n7920 & ~n12194;
  assign n12216 = ~n10819 & ~n12215;
  assign n12217 = ~n7728 & ~n12216;
  assign n12218 = ~n12214 & ~n12217;
  assign n12219 = ~n7723 & ~n12218;
  assign n12220 = ~n7723 & ~n12219;
  assign n12221 = ~n7714 & ~n12220;
  assign n12222 = ~n7714 & ~n12221;
  assign n12223 = n7705 & ~n12222;
  assign n12224 = ~n10888 & ~n12215;
  assign n12225 = n7728 & ~n12224;
  assign n12226 = ~n10920 & ~n12215;
  assign n12227 = ~n7728 & ~n12226;
  assign n12228 = ~n12225 & ~n12227;
  assign n12229 = n7723 & ~n12228;
  assign n12230 = ~n7723 & ~n12226;
  assign n12231 = ~n12229 & ~n12230;
  assign n12232 = n7714 & ~n12231;
  assign n12233 = n7723 & ~n12226;
  assign n12234 = ~n10920 & ~n12102;
  assign n12235 = n7728 & ~n12234;
  assign n12236 = ~n12138 & ~n12235;
  assign n12237 = ~n7723 & ~n12236;
  assign n12238 = ~n12233 & ~n12237;
  assign n12239 = ~n7714 & ~n12238;
  assign n12240 = ~n12232 & ~n12239;
  assign n12241 = ~n7705 & ~n12240;
  assign n12242 = ~n12223 & ~n12241;
  assign n12243 = n7808 & ~n12242;
  assign n12244 = ~n12211 & ~n12243;
  assign n12245 = n8195 & ~n12244;
  assign n12246 = ~n12170 & ~n12245;
  assign n12247 = n8193 & ~n12246;
  assign n12248 = ~n12150 & ~n12247;
  assign n12249 = ~n8191 & ~n12248;
  assign n12250 = ~n12075 & ~n12249;
  assign n12251 = n8188 & ~n12250;
  assign n12252 = ~n11286 & ~n11811;
  assign n12253 = n7728 & ~n12252;
  assign n12254 = ~n11335 & ~n11831;
  assign n12255 = ~n7728 & ~n12254;
  assign n12256 = ~n12253 & ~n12255;
  assign n12257 = ~n7723 & ~n12256;
  assign n12258 = ~n7723 & ~n12257;
  assign n12259 = ~n7714 & ~n12258;
  assign n12260 = ~n7714 & ~n12259;
  assign n12261 = n7705 & ~n12260;
  assign n12262 = n7723 & ~n12254;
  assign n12263 = ~n11359 & ~n11846;
  assign n12264 = i_hlock7 & ~n12263;
  assign n12265 = ~n11359 & ~n11854;
  assign n12266 = ~i_hlock7 & ~n12265;
  assign n12267 = ~n12264 & ~n12266;
  assign n12268 = i_hbusreq7 & ~n12267;
  assign n12269 = ~n11385 & ~n11870;
  assign n12270 = i_hlock7 & ~n12269;
  assign n12271 = ~n11385 & ~n11884;
  assign n12272 = ~i_hlock7 & ~n12271;
  assign n12273 = ~n12270 & ~n12272;
  assign n12274 = ~i_hbusreq7 & ~n12273;
  assign n12275 = ~n12268 & ~n12274;
  assign n12276 = n7924 & ~n12275;
  assign n12277 = ~n8337 & ~n12276;
  assign n12278 = ~n7920 & ~n12277;
  assign n12279 = n7920 & ~n12254;
  assign n12280 = ~n12278 & ~n12279;
  assign n12281 = ~n7723 & ~n12280;
  assign n12282 = ~n12262 & ~n12281;
  assign n12283 = n7714 & ~n12282;
  assign n12284 = ~n7714 & ~n12277;
  assign n12285 = ~n12283 & ~n12284;
  assign n12286 = ~n7705 & ~n12285;
  assign n12287 = ~n12261 & ~n12286;
  assign n12288 = ~n7808 & ~n12287;
  assign n12289 = ~n7920 & ~n12252;
  assign n12290 = ~n8874 & ~n12289;
  assign n12291 = n7728 & ~n12290;
  assign n12292 = ~n7920 & ~n12254;
  assign n12293 = ~n8974 & ~n12292;
  assign n12294 = ~n7728 & ~n12293;
  assign n12295 = ~n12291 & ~n12294;
  assign n12296 = ~n7723 & ~n12295;
  assign n12297 = ~n7723 & ~n12296;
  assign n12298 = ~n7714 & ~n12297;
  assign n12299 = ~n7714 & ~n12298;
  assign n12300 = n7705 & ~n12299;
  assign n12301 = ~n9181 & ~n12292;
  assign n12302 = n7728 & ~n12301;
  assign n12303 = ~n9577 & ~n12292;
  assign n12304 = ~n7728 & ~n12303;
  assign n12305 = ~n12302 & ~n12304;
  assign n12306 = n7723 & ~n12305;
  assign n12307 = ~n7723 & ~n12303;
  assign n12308 = ~n12306 & ~n12307;
  assign n12309 = n7714 & ~n12308;
  assign n12310 = n7723 & ~n12303;
  assign n12311 = ~n9577 & ~n12278;
  assign n12312 = n7728 & ~n12311;
  assign n12313 = ~n9738 & ~n12278;
  assign n12314 = ~n7728 & ~n12313;
  assign n12315 = ~n12312 & ~n12314;
  assign n12316 = ~n7723 & ~n12315;
  assign n12317 = ~n12310 & ~n12316;
  assign n12318 = ~n7714 & ~n12317;
  assign n12319 = ~n12309 & ~n12318;
  assign n12320 = ~n7705 & ~n12319;
  assign n12321 = ~n12300 & ~n12320;
  assign n12322 = n7808 & ~n12321;
  assign n12323 = ~n12288 & ~n12322;
  assign n12324 = n8195 & ~n12323;
  assign n12325 = ~n8196 & ~n12324;
  assign n12326 = ~n8193 & ~n12325;
  assign n12327 = ~n9900 & ~n12278;
  assign n12328 = ~n7723 & ~n12327;
  assign n12329 = ~n9899 & ~n12328;
  assign n12330 = n7714 & ~n12329;
  assign n12331 = ~n12284 & ~n12330;
  assign n12332 = ~n7705 & ~n12331;
  assign n12333 = ~n9898 & ~n12332;
  assign n12334 = ~n7808 & ~n12333;
  assign n12335 = ~n10274 & ~n12278;
  assign n12336 = n7728 & ~n12335;
  assign n12337 = ~n12314 & ~n12336;
  assign n12338 = ~n7723 & ~n12337;
  assign n12339 = ~n10282 & ~n12338;
  assign n12340 = ~n7714 & ~n12339;
  assign n12341 = ~n10281 & ~n12340;
  assign n12342 = ~n7705 & ~n12341;
  assign n12343 = ~n10052 & ~n12342;
  assign n12344 = n7808 & ~n12343;
  assign n12345 = ~n12334 & ~n12344;
  assign n12346 = ~n8195 & ~n12345;
  assign n12347 = ~n11476 & ~n11966;
  assign n12348 = i_hlock7 & ~n12347;
  assign n12349 = ~n11476 & ~n11974;
  assign n12350 = ~i_hlock7 & ~n12349;
  assign n12351 = ~n12348 & ~n12350;
  assign n12352 = i_hbusreq7 & ~n12351;
  assign n12353 = ~n11504 & ~n11990;
  assign n12354 = i_hlock7 & ~n12353;
  assign n12355 = ~n11504 & ~n12004;
  assign n12356 = ~i_hlock7 & ~n12355;
  assign n12357 = ~n12354 & ~n12356;
  assign n12358 = ~i_hbusreq7 & ~n12357;
  assign n12359 = ~n12352 & ~n12358;
  assign n12360 = n7924 & ~n12359;
  assign n12361 = ~n10375 & ~n12360;
  assign n12362 = n8214 & ~n12361;
  assign n12363 = n8214 & ~n12362;
  assign n12364 = n8202 & ~n12363;
  assign n12365 = ~n10332 & ~n12364;
  assign n12366 = n7728 & ~n12365;
  assign n12367 = n8214 & ~n12277;
  assign n12368 = ~n8336 & ~n12367;
  assign n12369 = n8202 & ~n12368;
  assign n12370 = ~n10649 & ~n12369;
  assign n12371 = ~n7728 & ~n12370;
  assign n12372 = ~n12366 & ~n12371;
  assign n12373 = ~n7723 & ~n12372;
  assign n12374 = ~n7723 & ~n12373;
  assign n12375 = ~n7714 & ~n12374;
  assign n12376 = ~n7714 & ~n12375;
  assign n12377 = n7705 & ~n12376;
  assign n12378 = n7723 & ~n12370;
  assign n12379 = n7920 & ~n12370;
  assign n12380 = ~n12278 & ~n12379;
  assign n12381 = ~n7723 & ~n12380;
  assign n12382 = ~n12378 & ~n12381;
  assign n12383 = n7714 & ~n12382;
  assign n12384 = ~n12284 & ~n12383;
  assign n12385 = ~n7705 & ~n12384;
  assign n12386 = ~n12377 & ~n12385;
  assign n12387 = ~n7808 & ~n12386;
  assign n12388 = ~n7920 & ~n12365;
  assign n12389 = ~n10794 & ~n12388;
  assign n12390 = n7728 & ~n12389;
  assign n12391 = ~n7920 & ~n12370;
  assign n12392 = ~n10819 & ~n12391;
  assign n12393 = ~n7728 & ~n12392;
  assign n12394 = ~n12390 & ~n12393;
  assign n12395 = ~n7723 & ~n12394;
  assign n12396 = ~n7723 & ~n12395;
  assign n12397 = ~n7714 & ~n12396;
  assign n12398 = ~n7714 & ~n12397;
  assign n12399 = n7705 & ~n12398;
  assign n12400 = ~n10888 & ~n12391;
  assign n12401 = n7728 & ~n12400;
  assign n12402 = ~n10920 & ~n12391;
  assign n12403 = ~n7728 & ~n12402;
  assign n12404 = ~n12401 & ~n12403;
  assign n12405 = n7723 & ~n12404;
  assign n12406 = ~n7723 & ~n12402;
  assign n12407 = ~n12405 & ~n12406;
  assign n12408 = n7714 & ~n12407;
  assign n12409 = n7723 & ~n12402;
  assign n12410 = ~n10920 & ~n12278;
  assign n12411 = n7728 & ~n12410;
  assign n12412 = ~n12314 & ~n12411;
  assign n12413 = ~n7723 & ~n12412;
  assign n12414 = ~n12409 & ~n12413;
  assign n12415 = ~n7714 & ~n12414;
  assign n12416 = ~n12408 & ~n12415;
  assign n12417 = ~n7705 & ~n12416;
  assign n12418 = ~n12399 & ~n12417;
  assign n12419 = n7808 & ~n12418;
  assign n12420 = ~n12387 & ~n12419;
  assign n12421 = n8195 & ~n12420;
  assign n12422 = ~n12346 & ~n12421;
  assign n12423 = n8193 & ~n12422;
  assign n12424 = ~n12326 & ~n12423;
  assign n12425 = n8191 & ~n12424;
  assign n12426 = ~n11575 & ~n11811;
  assign n12427 = n7728 & ~n12426;
  assign n12428 = ~n11579 & ~n11831;
  assign n12429 = ~n7728 & ~n12428;
  assign n12430 = ~n12427 & ~n12429;
  assign n12431 = ~n7723 & ~n12430;
  assign n12432 = ~n7723 & ~n12431;
  assign n12433 = ~n7714 & ~n12432;
  assign n12434 = ~n7714 & ~n12433;
  assign n12435 = n7705 & ~n12434;
  assign n12436 = n7723 & ~n12428;
  assign n12437 = ~n11594 & ~n11846;
  assign n12438 = i_hlock7 & ~n12437;
  assign n12439 = ~n11594 & ~n11854;
  assign n12440 = ~i_hlock7 & ~n12439;
  assign n12441 = ~n12438 & ~n12440;
  assign n12442 = i_hbusreq7 & ~n12441;
  assign n12443 = ~n11605 & ~n11870;
  assign n12444 = i_hlock7 & ~n12443;
  assign n12445 = ~n11605 & ~n11884;
  assign n12446 = ~i_hlock7 & ~n12445;
  assign n12447 = ~n12444 & ~n12446;
  assign n12448 = ~i_hbusreq7 & ~n12447;
  assign n12449 = ~n12442 & ~n12448;
  assign n12450 = n7924 & ~n12449;
  assign n12451 = ~n8337 & ~n12450;
  assign n12452 = ~n7920 & ~n12451;
  assign n12453 = n7920 & ~n12428;
  assign n12454 = ~n12452 & ~n12453;
  assign n12455 = ~n7723 & ~n12454;
  assign n12456 = ~n12436 & ~n12455;
  assign n12457 = n7714 & ~n12456;
  assign n12458 = ~n7714 & ~n12451;
  assign n12459 = ~n12457 & ~n12458;
  assign n12460 = ~n7705 & ~n12459;
  assign n12461 = ~n12435 & ~n12460;
  assign n12462 = ~n7808 & ~n12461;
  assign n12463 = ~n7920 & ~n12426;
  assign n12464 = ~n8874 & ~n12463;
  assign n12465 = n7728 & ~n12464;
  assign n12466 = ~n7920 & ~n12428;
  assign n12467 = ~n8974 & ~n12466;
  assign n12468 = ~n7728 & ~n12467;
  assign n12469 = ~n12465 & ~n12468;
  assign n12470 = ~n7723 & ~n12469;
  assign n12471 = ~n7723 & ~n12470;
  assign n12472 = ~n7714 & ~n12471;
  assign n12473 = ~n7714 & ~n12472;
  assign n12474 = n7705 & ~n12473;
  assign n12475 = ~n9181 & ~n12466;
  assign n12476 = n7728 & ~n12475;
  assign n12477 = ~n9577 & ~n12466;
  assign n12478 = ~n7728 & ~n12477;
  assign n12479 = ~n12476 & ~n12478;
  assign n12480 = n7723 & ~n12479;
  assign n12481 = ~n7723 & ~n12477;
  assign n12482 = ~n12480 & ~n12481;
  assign n12483 = n7714 & ~n12482;
  assign n12484 = n7723 & ~n12477;
  assign n12485 = ~n9577 & ~n12452;
  assign n12486 = n7728 & ~n12485;
  assign n12487 = ~n9738 & ~n12452;
  assign n12488 = ~n7728 & ~n12487;
  assign n12489 = ~n12486 & ~n12488;
  assign n12490 = ~n7723 & ~n12489;
  assign n12491 = ~n12484 & ~n12490;
  assign n12492 = ~n7714 & ~n12491;
  assign n12493 = ~n12483 & ~n12492;
  assign n12494 = ~n7705 & ~n12493;
  assign n12495 = ~n12474 & ~n12494;
  assign n12496 = n7808 & ~n12495;
  assign n12497 = ~n12462 & ~n12496;
  assign n12498 = n8195 & ~n12497;
  assign n12499 = ~n8196 & ~n12498;
  assign n12500 = ~n8193 & ~n12499;
  assign n12501 = ~n9900 & ~n12452;
  assign n12502 = ~n7723 & ~n12501;
  assign n12503 = ~n9899 & ~n12502;
  assign n12504 = n7714 & ~n12503;
  assign n12505 = ~n12458 & ~n12504;
  assign n12506 = ~n7705 & ~n12505;
  assign n12507 = ~n9898 & ~n12506;
  assign n12508 = ~n7808 & ~n12507;
  assign n12509 = ~n10274 & ~n12452;
  assign n12510 = n7728 & ~n12509;
  assign n12511 = ~n12488 & ~n12510;
  assign n12512 = ~n7723 & ~n12511;
  assign n12513 = ~n10282 & ~n12512;
  assign n12514 = ~n7714 & ~n12513;
  assign n12515 = ~n10281 & ~n12514;
  assign n12516 = ~n7705 & ~n12515;
  assign n12517 = ~n10052 & ~n12516;
  assign n12518 = n7808 & ~n12517;
  assign n12519 = ~n12508 & ~n12518;
  assign n12520 = ~n8195 & ~n12519;
  assign n12521 = ~n11685 & ~n11966;
  assign n12522 = i_hlock7 & ~n12521;
  assign n12523 = ~n11685 & ~n11974;
  assign n12524 = ~i_hlock7 & ~n12523;
  assign n12525 = ~n12522 & ~n12524;
  assign n12526 = i_hbusreq7 & ~n12525;
  assign n12527 = ~n11696 & ~n11990;
  assign n12528 = i_hlock7 & ~n12527;
  assign n12529 = ~n11696 & ~n12004;
  assign n12530 = ~i_hlock7 & ~n12529;
  assign n12531 = ~n12528 & ~n12530;
  assign n12532 = ~i_hbusreq7 & ~n12531;
  assign n12533 = ~n12526 & ~n12532;
  assign n12534 = n7924 & ~n12533;
  assign n12535 = ~n10375 & ~n12534;
  assign n12536 = n8214 & ~n12535;
  assign n12537 = n8214 & ~n12536;
  assign n12538 = n8202 & ~n12537;
  assign n12539 = ~n10332 & ~n12538;
  assign n12540 = n7728 & ~n12539;
  assign n12541 = n8214 & ~n12451;
  assign n12542 = ~n8336 & ~n12541;
  assign n12543 = n8202 & ~n12542;
  assign n12544 = ~n10649 & ~n12543;
  assign n12545 = ~n7728 & ~n12544;
  assign n12546 = ~n12540 & ~n12545;
  assign n12547 = ~n7723 & ~n12546;
  assign n12548 = ~n7723 & ~n12547;
  assign n12549 = ~n7714 & ~n12548;
  assign n12550 = ~n7714 & ~n12549;
  assign n12551 = n7705 & ~n12550;
  assign n12552 = n7723 & ~n12544;
  assign n12553 = n7920 & ~n12544;
  assign n12554 = ~n12452 & ~n12553;
  assign n12555 = ~n7723 & ~n12554;
  assign n12556 = ~n12552 & ~n12555;
  assign n12557 = n7714 & ~n12556;
  assign n12558 = ~n12458 & ~n12557;
  assign n12559 = ~n7705 & ~n12558;
  assign n12560 = ~n12551 & ~n12559;
  assign n12561 = ~n7808 & ~n12560;
  assign n12562 = ~n7920 & ~n12539;
  assign n12563 = ~n10794 & ~n12562;
  assign n12564 = n7728 & ~n12563;
  assign n12565 = ~n7920 & ~n12544;
  assign n12566 = ~n10819 & ~n12565;
  assign n12567 = ~n7728 & ~n12566;
  assign n12568 = ~n12564 & ~n12567;
  assign n12569 = ~n7723 & ~n12568;
  assign n12570 = ~n7723 & ~n12569;
  assign n12571 = ~n7714 & ~n12570;
  assign n12572 = ~n7714 & ~n12571;
  assign n12573 = n7705 & ~n12572;
  assign n12574 = ~n10888 & ~n12565;
  assign n12575 = n7728 & ~n12574;
  assign n12576 = ~n10920 & ~n12565;
  assign n12577 = ~n7728 & ~n12576;
  assign n12578 = ~n12575 & ~n12577;
  assign n12579 = n7723 & ~n12578;
  assign n12580 = ~n7723 & ~n12576;
  assign n12581 = ~n12579 & ~n12580;
  assign n12582 = n7714 & ~n12581;
  assign n12583 = n7723 & ~n12576;
  assign n12584 = ~n10920 & ~n12452;
  assign n12585 = n7728 & ~n12584;
  assign n12586 = ~n12488 & ~n12585;
  assign n12587 = ~n7723 & ~n12586;
  assign n12588 = ~n12583 & ~n12587;
  assign n12589 = ~n7714 & ~n12588;
  assign n12590 = ~n12582 & ~n12589;
  assign n12591 = ~n7705 & ~n12590;
  assign n12592 = ~n12573 & ~n12591;
  assign n12593 = n7808 & ~n12592;
  assign n12594 = ~n12561 & ~n12593;
  assign n12595 = n8195 & ~n12594;
  assign n12596 = ~n12520 & ~n12595;
  assign n12597 = n8193 & ~n12596;
  assign n12598 = ~n12500 & ~n12597;
  assign n12599 = ~n8191 & ~n12598;
  assign n12600 = ~n12425 & ~n12599;
  assign n12601 = ~n8188 & ~n12600;
  assign n12602 = ~n12251 & ~n12601;
  assign n12603 = ~n8185 & ~n12602;
  assign n12604 = ~n11769 & ~n12603;
  assign n12605 = controllable_hgrant7 & ~n12604;
  assign n12606 = controllable_hgrant8 & ~n12604;
  assign n12607 = controllable_hgrant6 & ~n8661;
  assign n12608 = controllable_hgrant5 & ~n8657;
  assign n12609 = controllable_hgrant4 & ~n8657;
  assign n12610 = controllable_hgrant3 & ~n8653;
  assign n12611 = controllable_hgrant1 & ~n8653;
  assign n12612 = controllable_hgrant2 & ~n8218;
  assign n12613 = controllable_hmastlock & ~n7858;
  assign n12614 = controllable_locked & ~n12613;
  assign n12615 = ~controllable_locked & ~n8218;
  assign n12616 = ~n12614 & ~n12615;
  assign n12617 = ~controllable_hgrant2 & ~n12616;
  assign n12618 = ~n12612 & ~n12617;
  assign n12619 = ~n7733 & ~n12618;
  assign n12620 = ~n7733 & ~n12619;
  assign n12621 = ~n7928 & ~n12620;
  assign n12622 = ~n7858 & ~n8231;
  assign n12623 = controllable_locked & ~n12622;
  assign n12624 = controllable_ndecide & ~controllable_hmastlock;
  assign n12625 = ~n7818 & ~n12624;
  assign n12626 = ~controllable_locked & ~n12625;
  assign n12627 = ~n12623 & ~n12626;
  assign n12628 = ~controllable_hgrant2 & ~n12627;
  assign n12629 = ~n7814 & ~n12628;
  assign n12630 = n7928 & ~n12629;
  assign n12631 = ~n12621 & ~n12630;
  assign n12632 = ~controllable_hgrant1 & ~n12631;
  assign n12633 = ~n12611 & ~n12632;
  assign n12634 = ~controllable_hgrant3 & ~n12633;
  assign n12635 = ~n12610 & ~n12634;
  assign n12636 = i_hlock9 & ~n12635;
  assign n12637 = controllable_hgrant3 & ~n8655;
  assign n12638 = controllable_hgrant1 & ~n8655;
  assign n12639 = controllable_hgrant2 & ~n8232;
  assign n12640 = controllable_locked & ~n8232;
  assign n12641 = ~controllable_hmastlock & ~n12624;
  assign n12642 = ~controllable_locked & ~n12641;
  assign n12643 = ~n12640 & ~n12642;
  assign n12644 = ~controllable_hgrant2 & ~n12643;
  assign n12645 = ~n12639 & ~n12644;
  assign n12646 = ~n7733 & ~n12645;
  assign n12647 = ~n7733 & ~n12646;
  assign n12648 = ~n7928 & ~n12647;
  assign n12649 = ~n12630 & ~n12648;
  assign n12650 = ~controllable_hgrant1 & ~n12649;
  assign n12651 = ~n12638 & ~n12650;
  assign n12652 = ~controllable_hgrant3 & ~n12651;
  assign n12653 = ~n12637 & ~n12652;
  assign n12654 = ~i_hlock9 & ~n12653;
  assign n12655 = ~n12636 & ~n12654;
  assign n12656 = ~controllable_hgrant4 & ~n12655;
  assign n12657 = ~n12609 & ~n12656;
  assign n12658 = ~controllable_hgrant5 & ~n12657;
  assign n12659 = ~n12608 & ~n12658;
  assign n12660 = ~controllable_hmaster2 & ~n12659;
  assign n12661 = ~controllable_hmaster2 & ~n12660;
  assign n12662 = ~controllable_hmaster1 & ~n12661;
  assign n12663 = ~controllable_hmaster1 & ~n12662;
  assign n12664 = ~controllable_hgrant6 & ~n12663;
  assign n12665 = ~n12607 & ~n12664;
  assign n12666 = controllable_hmaster0 & ~n12665;
  assign n12667 = controllable_hmaster0 & ~n12666;
  assign n12668 = controllable_hmaster3 & ~n12667;
  assign n12669 = controllable_hmaster3 & ~n12668;
  assign n12670 = i_hbusreq7 & ~n12669;
  assign n12671 = i_hbusreq8 & ~n12667;
  assign n12672 = controllable_hgrant6 & ~n8716;
  assign n12673 = i_hbusreq6 & ~n12663;
  assign n12674 = controllable_hgrant5 & ~n8710;
  assign n12675 = i_hbusreq5 & ~n12657;
  assign n12676 = controllable_hgrant4 & ~n8708;
  assign n12677 = i_hbusreq4 & ~n12655;
  assign n12678 = i_hbusreq9 & ~n12655;
  assign n12679 = controllable_hgrant3 & ~n8694;
  assign n12680 = i_hbusreq3 & ~n12633;
  assign n12681 = controllable_hgrant1 & ~n8692;
  assign n12682 = i_hbusreq1 & ~n12631;
  assign n12683 = controllable_hgrant2 & ~n8262;
  assign n12684 = i_hbusreq2 & ~n12616;
  assign n12685 = i_hbusreq0 & ~n12616;
  assign n12686 = i_hbusreq0 & ~n12685;
  assign n12687 = ~i_hbusreq2 & ~n12686;
  assign n12688 = ~n12684 & ~n12687;
  assign n12689 = ~controllable_hgrant2 & ~n12688;
  assign n12690 = ~n12683 & ~n12689;
  assign n12691 = ~n7733 & ~n12690;
  assign n12692 = ~n7733 & ~n12691;
  assign n12693 = ~n7928 & ~n12692;
  assign n12694 = controllable_hgrant2 & ~n8679;
  assign n12695 = i_hbusreq2 & ~n12627;
  assign n12696 = i_hbusreq0 & ~n12627;
  assign n12697 = ~i_hlock0 & ~n12627;
  assign n12698 = ~i_hlock0 & ~n12697;
  assign n12699 = ~i_hbusreq0 & ~n12698;
  assign n12700 = ~n12696 & ~n12699;
  assign n12701 = ~i_hbusreq2 & ~n12700;
  assign n12702 = ~n12695 & ~n12701;
  assign n12703 = ~controllable_hgrant2 & ~n12702;
  assign n12704 = ~n12694 & ~n12703;
  assign n12705 = ~n7733 & ~n12704;
  assign n12706 = controllable_hgrant2 & ~n8686;
  assign n12707 = i_hlock0 & ~n12643;
  assign n12708 = ~n12697 & ~n12707;
  assign n12709 = ~i_hbusreq0 & ~n12708;
  assign n12710 = ~n12696 & ~n12709;
  assign n12711 = ~i_hbusreq2 & ~n12710;
  assign n12712 = ~n12695 & ~n12711;
  assign n12713 = ~controllable_hgrant2 & ~n12712;
  assign n12714 = ~n12706 & ~n12713;
  assign n12715 = n7733 & ~n12714;
  assign n12716 = ~n12705 & ~n12715;
  assign n12717 = n7928 & ~n12716;
  assign n12718 = ~n12693 & ~n12717;
  assign n12719 = ~i_hbusreq1 & ~n12718;
  assign n12720 = ~n12682 & ~n12719;
  assign n12721 = ~controllable_hgrant1 & ~n12720;
  assign n12722 = ~n12681 & ~n12721;
  assign n12723 = ~i_hbusreq3 & ~n12722;
  assign n12724 = ~n12680 & ~n12723;
  assign n12725 = ~controllable_hgrant3 & ~n12724;
  assign n12726 = ~n12679 & ~n12725;
  assign n12727 = i_hlock9 & ~n12726;
  assign n12728 = controllable_hgrant3 & ~n8702;
  assign n12729 = i_hbusreq3 & ~n12651;
  assign n12730 = controllable_hgrant1 & ~n8700;
  assign n12731 = i_hbusreq1 & ~n12649;
  assign n12732 = controllable_hgrant2 & ~n8294;
  assign n12733 = i_hbusreq2 & ~n12643;
  assign n12734 = i_hbusreq0 & ~n12643;
  assign n12735 = i_hbusreq0 & ~n12734;
  assign n12736 = ~i_hbusreq2 & ~n12735;
  assign n12737 = ~n12733 & ~n12736;
  assign n12738 = ~controllable_hgrant2 & ~n12737;
  assign n12739 = ~n12732 & ~n12738;
  assign n12740 = ~n7733 & ~n12739;
  assign n12741 = ~n7733 & ~n12740;
  assign n12742 = ~n7928 & ~n12741;
  assign n12743 = ~n12717 & ~n12742;
  assign n12744 = ~i_hbusreq1 & ~n12743;
  assign n12745 = ~n12731 & ~n12744;
  assign n12746 = ~controllable_hgrant1 & ~n12745;
  assign n12747 = ~n12730 & ~n12746;
  assign n12748 = ~i_hbusreq3 & ~n12747;
  assign n12749 = ~n12729 & ~n12748;
  assign n12750 = ~controllable_hgrant3 & ~n12749;
  assign n12751 = ~n12728 & ~n12750;
  assign n12752 = ~i_hlock9 & ~n12751;
  assign n12753 = ~n12727 & ~n12752;
  assign n12754 = ~i_hbusreq9 & ~n12753;
  assign n12755 = ~n12678 & ~n12754;
  assign n12756 = ~i_hbusreq4 & ~n12755;
  assign n12757 = ~n12677 & ~n12756;
  assign n12758 = ~controllable_hgrant4 & ~n12757;
  assign n12759 = ~n12676 & ~n12758;
  assign n12760 = ~i_hbusreq5 & ~n12759;
  assign n12761 = ~n12675 & ~n12760;
  assign n12762 = ~controllable_hgrant5 & ~n12761;
  assign n12763 = ~n12674 & ~n12762;
  assign n12764 = ~controllable_hmaster2 & ~n12763;
  assign n12765 = ~controllable_hmaster2 & ~n12764;
  assign n12766 = ~controllable_hmaster1 & ~n12765;
  assign n12767 = ~controllable_hmaster1 & ~n12766;
  assign n12768 = ~i_hbusreq6 & ~n12767;
  assign n12769 = ~n12673 & ~n12768;
  assign n12770 = ~controllable_hgrant6 & ~n12769;
  assign n12771 = ~n12672 & ~n12770;
  assign n12772 = controllable_hmaster0 & ~n12771;
  assign n12773 = controllable_hmaster0 & ~n12772;
  assign n12774 = ~i_hbusreq8 & ~n12773;
  assign n12775 = ~n12671 & ~n12774;
  assign n12776 = controllable_hmaster3 & ~n12775;
  assign n12777 = controllable_hmaster3 & ~n12776;
  assign n12778 = ~i_hbusreq7 & ~n12777;
  assign n12779 = ~n12670 & ~n12778;
  assign n12780 = ~n7924 & ~n12779;
  assign n12781 = ~i_hready & ~controllable_ndecide;
  assign n12782 = ~controllable_ndecide & ~n12781;
  assign n12783 = ~controllable_locked & ~n12782;
  assign n12784 = ~controllable_locked & ~n12783;
  assign n12785 = ~controllable_hgrant2 & ~n12784;
  assign n12786 = ~controllable_hgrant2 & ~n12785;
  assign n12787 = n7928 & ~n12786;
  assign n12788 = n7928 & ~n12787;
  assign n12789 = ~controllable_hgrant1 & ~n12788;
  assign n12790 = ~controllable_hgrant1 & ~n12789;
  assign n12791 = ~controllable_hgrant3 & ~n12790;
  assign n12792 = ~controllable_hgrant3 & ~n12791;
  assign n12793 = ~controllable_hgrant4 & ~n12792;
  assign n12794 = ~controllable_hgrant4 & ~n12793;
  assign n12795 = ~controllable_hgrant5 & ~n12794;
  assign n12796 = ~controllable_hgrant5 & ~n12795;
  assign n12797 = controllable_hmaster1 & ~n12796;
  assign n12798 = controllable_hmaster2 & ~n12796;
  assign n12799 = ~controllable_locked & controllable_ndecide;
  assign n12800 = ~n12623 & ~n12799;
  assign n12801 = ~controllable_hgrant2 & ~n12800;
  assign n12802 = ~n7814 & ~n12801;
  assign n12803 = n7928 & ~n12802;
  assign n12804 = ~n12621 & ~n12803;
  assign n12805 = ~controllable_hgrant1 & ~n12804;
  assign n12806 = ~n12611 & ~n12805;
  assign n12807 = ~controllable_hgrant3 & ~n12806;
  assign n12808 = ~n12610 & ~n12807;
  assign n12809 = i_hlock9 & ~n12808;
  assign n12810 = ~n12648 & ~n12803;
  assign n12811 = ~controllable_hgrant1 & ~n12810;
  assign n12812 = ~n12638 & ~n12811;
  assign n12813 = ~controllable_hgrant3 & ~n12812;
  assign n12814 = ~n12637 & ~n12813;
  assign n12815 = ~i_hlock9 & ~n12814;
  assign n12816 = ~n12809 & ~n12815;
  assign n12817 = ~controllable_hgrant4 & ~n12816;
  assign n12818 = ~n12609 & ~n12817;
  assign n12819 = ~controllable_hgrant5 & ~n12818;
  assign n12820 = ~n12608 & ~n12819;
  assign n12821 = ~controllable_hmaster2 & ~n12820;
  assign n12822 = ~n12798 & ~n12821;
  assign n12823 = ~controllable_hmaster1 & ~n12822;
  assign n12824 = ~n12797 & ~n12823;
  assign n12825 = ~controllable_hgrant6 & ~n12824;
  assign n12826 = ~n12607 & ~n12825;
  assign n12827 = controllable_hmaster0 & ~n12826;
  assign n12828 = ~controllable_hgrant6 & ~n12796;
  assign n12829 = ~controllable_hgrant6 & ~n12828;
  assign n12830 = ~controllable_hmaster0 & ~n12829;
  assign n12831 = ~n12827 & ~n12830;
  assign n12832 = controllable_hmaster3 & ~n12831;
  assign n12833 = ~controllable_hmaster3 & ~n12829;
  assign n12834 = ~n12832 & ~n12833;
  assign n12835 = i_hbusreq7 & ~n12834;
  assign n12836 = i_hbusreq8 & ~n12831;
  assign n12837 = i_hbusreq6 & ~n12824;
  assign n12838 = i_hbusreq5 & ~n12794;
  assign n12839 = i_hbusreq4 & ~n12792;
  assign n12840 = i_hbusreq9 & ~n12792;
  assign n12841 = i_hbusreq3 & ~n12790;
  assign n12842 = i_hbusreq1 & ~n12788;
  assign n12843 = i_hbusreq2 & ~n12784;
  assign n12844 = i_hbusreq0 & ~n12784;
  assign n12845 = ~i_hlock0 & ~n12784;
  assign n12846 = ~i_hlock0 & ~n12845;
  assign n12847 = ~i_hbusreq0 & ~n12846;
  assign n12848 = ~n12844 & ~n12847;
  assign n12849 = ~i_hbusreq2 & ~n12848;
  assign n12850 = ~n12843 & ~n12849;
  assign n12851 = ~controllable_hgrant2 & ~n12850;
  assign n12852 = ~controllable_hgrant2 & ~n12851;
  assign n12853 = ~n7733 & ~n12852;
  assign n12854 = n7733 & ~n12786;
  assign n12855 = ~n12853 & ~n12854;
  assign n12856 = n7928 & ~n12855;
  assign n12857 = n7928 & ~n12856;
  assign n12858 = ~i_hbusreq1 & ~n12857;
  assign n12859 = ~n12842 & ~n12858;
  assign n12860 = ~controllable_hgrant1 & ~n12859;
  assign n12861 = ~controllable_hgrant1 & ~n12860;
  assign n12862 = ~i_hbusreq3 & ~n12861;
  assign n12863 = ~n12841 & ~n12862;
  assign n12864 = ~controllable_hgrant3 & ~n12863;
  assign n12865 = ~controllable_hgrant3 & ~n12864;
  assign n12866 = ~i_hbusreq9 & ~n12865;
  assign n12867 = ~n12840 & ~n12866;
  assign n12868 = ~i_hbusreq4 & ~n12867;
  assign n12869 = ~n12839 & ~n12868;
  assign n12870 = ~controllable_hgrant4 & ~n12869;
  assign n12871 = ~controllable_hgrant4 & ~n12870;
  assign n12872 = ~i_hbusreq5 & ~n12871;
  assign n12873 = ~n12838 & ~n12872;
  assign n12874 = ~controllable_hgrant5 & ~n12873;
  assign n12875 = ~controllable_hgrant5 & ~n12874;
  assign n12876 = controllable_hmaster1 & ~n12875;
  assign n12877 = controllable_hmaster2 & ~n12875;
  assign n12878 = i_hbusreq5 & ~n12818;
  assign n12879 = i_hbusreq4 & ~n12816;
  assign n12880 = i_hbusreq9 & ~n12816;
  assign n12881 = i_hbusreq3 & ~n12806;
  assign n12882 = i_hbusreq1 & ~n12804;
  assign n12883 = i_hbusreq2 & ~n12800;
  assign n12884 = i_hbusreq0 & ~n12800;
  assign n12885 = ~i_hlock0 & ~n12800;
  assign n12886 = ~i_hlock0 & ~n12885;
  assign n12887 = ~i_hbusreq0 & ~n12886;
  assign n12888 = ~n12884 & ~n12887;
  assign n12889 = ~i_hbusreq2 & ~n12888;
  assign n12890 = ~n12883 & ~n12889;
  assign n12891 = ~controllable_hgrant2 & ~n12890;
  assign n12892 = ~n12694 & ~n12891;
  assign n12893 = ~n7733 & ~n12892;
  assign n12894 = controllable_hmastlock & ~n12782;
  assign n12895 = ~n12624 & ~n12894;
  assign n12896 = ~controllable_locked & ~n12895;
  assign n12897 = ~n12640 & ~n12896;
  assign n12898 = i_hlock0 & ~n12897;
  assign n12899 = ~n12885 & ~n12898;
  assign n12900 = ~i_hbusreq0 & ~n12899;
  assign n12901 = ~n12884 & ~n12900;
  assign n12902 = ~i_hbusreq2 & ~n12901;
  assign n12903 = ~n12883 & ~n12902;
  assign n12904 = ~controllable_hgrant2 & ~n12903;
  assign n12905 = ~n12706 & ~n12904;
  assign n12906 = n7733 & ~n12905;
  assign n12907 = ~n12893 & ~n12906;
  assign n12908 = n7928 & ~n12907;
  assign n12909 = ~n12693 & ~n12908;
  assign n12910 = ~i_hbusreq1 & ~n12909;
  assign n12911 = ~n12882 & ~n12910;
  assign n12912 = ~controllable_hgrant1 & ~n12911;
  assign n12913 = ~n12681 & ~n12912;
  assign n12914 = ~i_hbusreq3 & ~n12913;
  assign n12915 = ~n12881 & ~n12914;
  assign n12916 = ~controllable_hgrant3 & ~n12915;
  assign n12917 = ~n12679 & ~n12916;
  assign n12918 = i_hlock9 & ~n12917;
  assign n12919 = i_hbusreq3 & ~n12812;
  assign n12920 = i_hbusreq1 & ~n12810;
  assign n12921 = ~n12742 & ~n12908;
  assign n12922 = ~i_hbusreq1 & ~n12921;
  assign n12923 = ~n12920 & ~n12922;
  assign n12924 = ~controllable_hgrant1 & ~n12923;
  assign n12925 = ~n12730 & ~n12924;
  assign n12926 = ~i_hbusreq3 & ~n12925;
  assign n12927 = ~n12919 & ~n12926;
  assign n12928 = ~controllable_hgrant3 & ~n12927;
  assign n12929 = ~n12728 & ~n12928;
  assign n12930 = ~i_hlock9 & ~n12929;
  assign n12931 = ~n12918 & ~n12930;
  assign n12932 = ~i_hbusreq9 & ~n12931;
  assign n12933 = ~n12880 & ~n12932;
  assign n12934 = ~i_hbusreq4 & ~n12933;
  assign n12935 = ~n12879 & ~n12934;
  assign n12936 = ~controllable_hgrant4 & ~n12935;
  assign n12937 = ~n12676 & ~n12936;
  assign n12938 = ~i_hbusreq5 & ~n12937;
  assign n12939 = ~n12878 & ~n12938;
  assign n12940 = ~controllable_hgrant5 & ~n12939;
  assign n12941 = ~n12674 & ~n12940;
  assign n12942 = ~controllable_hmaster2 & ~n12941;
  assign n12943 = ~n12877 & ~n12942;
  assign n12944 = ~controllable_hmaster1 & ~n12943;
  assign n12945 = ~n12876 & ~n12944;
  assign n12946 = ~i_hbusreq6 & ~n12945;
  assign n12947 = ~n12837 & ~n12946;
  assign n12948 = ~controllable_hgrant6 & ~n12947;
  assign n12949 = ~n12672 & ~n12948;
  assign n12950 = controllable_hmaster0 & ~n12949;
  assign n12951 = i_hbusreq6 & ~n12796;
  assign n12952 = ~i_hbusreq6 & ~n12875;
  assign n12953 = ~n12951 & ~n12952;
  assign n12954 = ~controllable_hgrant6 & ~n12953;
  assign n12955 = ~controllable_hgrant6 & ~n12954;
  assign n12956 = ~controllable_hmaster0 & ~n12955;
  assign n12957 = ~n12950 & ~n12956;
  assign n12958 = ~i_hbusreq8 & ~n12957;
  assign n12959 = ~n12836 & ~n12958;
  assign n12960 = controllable_hmaster3 & ~n12959;
  assign n12961 = i_hbusreq8 & ~n12829;
  assign n12962 = ~i_hbusreq8 & ~n12955;
  assign n12963 = ~n12961 & ~n12962;
  assign n12964 = ~controllable_hmaster3 & ~n12963;
  assign n12965 = ~n12960 & ~n12964;
  assign n12966 = ~i_hbusreq7 & ~n12965;
  assign n12967 = ~n12835 & ~n12966;
  assign n12968 = n7924 & ~n12967;
  assign n12969 = ~n12780 & ~n12968;
  assign n12970 = ~n8214 & ~n12969;
  assign n12971 = ~n8790 & ~n12970;
  assign n12972 = ~n8202 & ~n12971;
  assign n12973 = ~n8872 & ~n12972;
  assign n12974 = n7920 & ~n12973;
  assign n12975 = ~n8651 & ~n12974;
  assign n12976 = n7728 & ~n12975;
  assign n12977 = controllable_hgrant6 & ~n8880;
  assign n12978 = ~n7739 & ~n12660;
  assign n12979 = ~controllable_hmaster1 & ~n12978;
  assign n12980 = ~n7738 & ~n12979;
  assign n12981 = ~controllable_hgrant6 & ~n12980;
  assign n12982 = ~n12977 & ~n12981;
  assign n12983 = controllable_hmaster0 & ~n12982;
  assign n12984 = ~n8882 & ~n12983;
  assign n12985 = controllable_hmaster3 & ~n12984;
  assign n12986 = controllable_hmaster3 & ~n12985;
  assign n12987 = i_hbusreq7 & ~n12986;
  assign n12988 = i_hbusreq8 & ~n12984;
  assign n12989 = controllable_hgrant6 & ~n8893;
  assign n12990 = i_hbusreq6 & ~n12980;
  assign n12991 = ~n7771 & ~n12764;
  assign n12992 = ~controllable_hmaster1 & ~n12991;
  assign n12993 = ~n7770 & ~n12992;
  assign n12994 = ~i_hbusreq6 & ~n12993;
  assign n12995 = ~n12990 & ~n12994;
  assign n12996 = ~controllable_hgrant6 & ~n12995;
  assign n12997 = ~n12989 & ~n12996;
  assign n12998 = controllable_hmaster0 & ~n12997;
  assign n12999 = ~n8895 & ~n12998;
  assign n13000 = ~i_hbusreq8 & ~n12999;
  assign n13001 = ~n12988 & ~n13000;
  assign n13002 = controllable_hmaster3 & ~n13001;
  assign n13003 = controllable_hmaster3 & ~n13002;
  assign n13004 = ~i_hbusreq7 & ~n13003;
  assign n13005 = ~n12987 & ~n13004;
  assign n13006 = ~n7924 & ~n13005;
  assign n13007 = ~n7737 & ~n7928;
  assign n13008 = controllable_locked & ~n7735;
  assign n13009 = ~n12799 & ~n13008;
  assign n13010 = ~controllable_hgrant2 & ~n13009;
  assign n13011 = ~n7814 & ~n13010;
  assign n13012 = ~n7733 & ~n13011;
  assign n13013 = ~n12854 & ~n13012;
  assign n13014 = n7928 & ~n13013;
  assign n13015 = ~n13007 & ~n13014;
  assign n13016 = ~controllable_hgrant1 & ~n13015;
  assign n13017 = ~n7813 & ~n13016;
  assign n13018 = ~controllable_hgrant3 & ~n13017;
  assign n13019 = ~n7812 & ~n13018;
  assign n13020 = ~controllable_hgrant4 & ~n13019;
  assign n13021 = ~n7811 & ~n13020;
  assign n13022 = ~controllable_hgrant5 & ~n13021;
  assign n13023 = ~n7810 & ~n13022;
  assign n13024 = controllable_hmaster1 & ~n13023;
  assign n13025 = controllable_hmaster2 & ~n13023;
  assign n13026 = ~n12821 & ~n13025;
  assign n13027 = ~controllable_hmaster1 & ~n13026;
  assign n13028 = ~n13024 & ~n13027;
  assign n13029 = ~controllable_hgrant6 & ~n13028;
  assign n13030 = ~n12977 & ~n13029;
  assign n13031 = controllable_hmaster0 & ~n13030;
  assign n13032 = ~controllable_hmaster2 & ~n12796;
  assign n13033 = ~n13025 & ~n13032;
  assign n13034 = ~controllable_hmaster1 & ~n13033;
  assign n13035 = ~n13024 & ~n13034;
  assign n13036 = ~controllable_hgrant6 & ~n13035;
  assign n13037 = ~n7809 & ~n13036;
  assign n13038 = ~controllable_hmaster0 & ~n13037;
  assign n13039 = ~n13031 & ~n13038;
  assign n13040 = controllable_hmaster3 & ~n13039;
  assign n13041 = ~n12833 & ~n13040;
  assign n13042 = i_hbusreq7 & ~n13041;
  assign n13043 = i_hbusreq8 & ~n13039;
  assign n13044 = i_hbusreq6 & ~n13028;
  assign n13045 = i_hbusreq5 & ~n13021;
  assign n13046 = i_hbusreq4 & ~n13019;
  assign n13047 = i_hbusreq9 & ~n13019;
  assign n13048 = i_hbusreq3 & ~n13017;
  assign n13049 = i_hbusreq1 & ~n13015;
  assign n13050 = ~n7759 & ~n7928;
  assign n13051 = i_hbusreq2 & ~n13009;
  assign n13052 = i_hbusreq0 & ~n13009;
  assign n13053 = ~n12847 & ~n13052;
  assign n13054 = ~i_hbusreq2 & ~n13053;
  assign n13055 = ~n13051 & ~n13054;
  assign n13056 = ~controllable_hgrant2 & ~n13055;
  assign n13057 = ~n7855 & ~n13056;
  assign n13058 = ~n7733 & ~n13057;
  assign n13059 = ~n12854 & ~n13058;
  assign n13060 = n7928 & ~n13059;
  assign n13061 = ~n13050 & ~n13060;
  assign n13062 = ~i_hbusreq1 & ~n13061;
  assign n13063 = ~n13049 & ~n13062;
  assign n13064 = ~controllable_hgrant1 & ~n13063;
  assign n13065 = ~n7853 & ~n13064;
  assign n13066 = ~i_hbusreq3 & ~n13065;
  assign n13067 = ~n13048 & ~n13066;
  assign n13068 = ~controllable_hgrant3 & ~n13067;
  assign n13069 = ~n7851 & ~n13068;
  assign n13070 = ~i_hbusreq9 & ~n13069;
  assign n13071 = ~n13047 & ~n13070;
  assign n13072 = ~i_hbusreq4 & ~n13071;
  assign n13073 = ~n13046 & ~n13072;
  assign n13074 = ~controllable_hgrant4 & ~n13073;
  assign n13075 = ~n7848 & ~n13074;
  assign n13076 = ~i_hbusreq5 & ~n13075;
  assign n13077 = ~n13045 & ~n13076;
  assign n13078 = ~controllable_hgrant5 & ~n13077;
  assign n13079 = ~n7846 & ~n13078;
  assign n13080 = controllable_hmaster1 & ~n13079;
  assign n13081 = controllable_hmaster2 & ~n13079;
  assign n13082 = ~n12942 & ~n13081;
  assign n13083 = ~controllable_hmaster1 & ~n13082;
  assign n13084 = ~n13080 & ~n13083;
  assign n13085 = ~i_hbusreq6 & ~n13084;
  assign n13086 = ~n13044 & ~n13085;
  assign n13087 = ~controllable_hgrant6 & ~n13086;
  assign n13088 = ~n12989 & ~n13087;
  assign n13089 = controllable_hmaster0 & ~n13088;
  assign n13090 = i_hbusreq6 & ~n13035;
  assign n13091 = ~controllable_hmaster2 & ~n12875;
  assign n13092 = ~n13081 & ~n13091;
  assign n13093 = ~controllable_hmaster1 & ~n13092;
  assign n13094 = ~n13080 & ~n13093;
  assign n13095 = ~i_hbusreq6 & ~n13094;
  assign n13096 = ~n13090 & ~n13095;
  assign n13097 = ~controllable_hgrant6 & ~n13096;
  assign n13098 = ~n7844 & ~n13097;
  assign n13099 = ~controllable_hmaster0 & ~n13098;
  assign n13100 = ~n13089 & ~n13099;
  assign n13101 = ~i_hbusreq8 & ~n13100;
  assign n13102 = ~n13043 & ~n13101;
  assign n13103 = controllable_hmaster3 & ~n13102;
  assign n13104 = ~n12964 & ~n13103;
  assign n13105 = ~i_hbusreq7 & ~n13104;
  assign n13106 = ~n13042 & ~n13105;
  assign n13107 = n7924 & ~n13106;
  assign n13108 = ~n13006 & ~n13107;
  assign n13109 = ~n8214 & ~n13108;
  assign n13110 = ~n8948 & ~n13109;
  assign n13111 = ~n8202 & ~n13110;
  assign n13112 = ~n8972 & ~n13111;
  assign n13113 = n7920 & ~n13112;
  assign n13114 = ~n8877 & ~n13113;
  assign n13115 = ~n7728 & ~n13114;
  assign n13116 = ~n12976 & ~n13115;
  assign n13117 = ~n7723 & ~n13116;
  assign n13118 = ~n7723 & ~n13117;
  assign n13119 = ~n7714 & ~n13118;
  assign n13120 = ~n7714 & ~n13119;
  assign n13121 = n7705 & ~n13120;
  assign n13122 = controllable_hgrant6 & ~n8985;
  assign n13123 = ~n8358 & ~n12660;
  assign n13124 = ~controllable_hmaster1 & ~n13123;
  assign n13125 = ~n8357 & ~n13124;
  assign n13126 = ~controllable_hgrant6 & ~n13125;
  assign n13127 = ~n13122 & ~n13126;
  assign n13128 = controllable_hmaster0 & ~n13127;
  assign n13129 = ~n8992 & ~n13128;
  assign n13130 = controllable_hmaster3 & ~n13129;
  assign n13131 = ~n8995 & ~n13130;
  assign n13132 = i_hbusreq7 & ~n13131;
  assign n13133 = i_hbusreq8 & ~n13129;
  assign n13134 = controllable_hgrant6 & ~n9004;
  assign n13135 = i_hbusreq6 & ~n13125;
  assign n13136 = ~n8484 & ~n12764;
  assign n13137 = ~controllable_hmaster1 & ~n13136;
  assign n13138 = ~n8483 & ~n13137;
  assign n13139 = ~i_hbusreq6 & ~n13138;
  assign n13140 = ~n13135 & ~n13139;
  assign n13141 = ~controllable_hgrant6 & ~n13140;
  assign n13142 = ~n13134 & ~n13141;
  assign n13143 = controllable_hmaster0 & ~n13142;
  assign n13144 = ~n9030 & ~n13143;
  assign n13145 = ~i_hbusreq8 & ~n13144;
  assign n13146 = ~n13133 & ~n13145;
  assign n13147 = controllable_hmaster3 & ~n13146;
  assign n13148 = ~n9041 & ~n13147;
  assign n13149 = ~i_hbusreq7 & ~n13148;
  assign n13150 = ~n13132 & ~n13149;
  assign n13151 = ~n7924 & ~n13150;
  assign n13152 = controllable_hgrant5 & ~n7735;
  assign n13153 = controllable_hgrant4 & ~n7735;
  assign n13154 = controllable_hgrant3 & ~n7735;
  assign n13155 = controllable_hgrant1 & ~n7735;
  assign n13156 = ~n7735 & ~n7928;
  assign n13157 = n7928 & ~n13011;
  assign n13158 = ~n13156 & ~n13157;
  assign n13159 = ~controllable_hgrant1 & ~n13158;
  assign n13160 = ~n13155 & ~n13159;
  assign n13161 = ~controllable_hgrant3 & ~n13160;
  assign n13162 = ~n13154 & ~n13161;
  assign n13163 = ~controllable_hgrant4 & ~n13162;
  assign n13164 = ~n13153 & ~n13163;
  assign n13165 = ~controllable_hgrant5 & ~n13164;
  assign n13166 = ~n13152 & ~n13165;
  assign n13167 = controllable_hmaster1 & ~n13166;
  assign n13168 = controllable_hmaster2 & ~n13166;
  assign n13169 = ~n12821 & ~n13168;
  assign n13170 = ~controllable_hmaster1 & ~n13169;
  assign n13171 = ~n13167 & ~n13170;
  assign n13172 = ~controllable_hgrant6 & ~n13171;
  assign n13173 = ~n13122 & ~n13172;
  assign n13174 = controllable_hmaster0 & ~n13173;
  assign n13175 = controllable_hgrant6 & ~n8991;
  assign n13176 = controllable_hgrant5 & ~n8987;
  assign n13177 = controllable_hgrant4 & ~n8987;
  assign n13178 = controllable_hgrant3 & ~n8987;
  assign n13179 = controllable_hgrant1 & ~n8987;
  assign n13180 = n7928 & ~n13157;
  assign n13181 = ~controllable_hgrant1 & ~n13180;
  assign n13182 = ~n13179 & ~n13181;
  assign n13183 = ~controllable_hgrant3 & ~n13182;
  assign n13184 = ~n13178 & ~n13183;
  assign n13185 = ~controllable_hgrant4 & ~n13184;
  assign n13186 = ~n13177 & ~n13185;
  assign n13187 = ~controllable_hgrant5 & ~n13186;
  assign n13188 = ~n13176 & ~n13187;
  assign n13189 = ~controllable_hmaster2 & ~n13188;
  assign n13190 = ~n13168 & ~n13189;
  assign n13191 = ~controllable_hmaster1 & ~n13190;
  assign n13192 = ~n13167 & ~n13191;
  assign n13193 = ~controllable_hgrant6 & ~n13192;
  assign n13194 = ~n13175 & ~n13193;
  assign n13195 = ~controllable_hmaster0 & ~n13194;
  assign n13196 = ~n13174 & ~n13195;
  assign n13197 = controllable_hmaster3 & ~n13196;
  assign n13198 = controllable_hgrant6 & ~n8987;
  assign n13199 = ~controllable_hgrant6 & ~n13188;
  assign n13200 = ~n13198 & ~n13199;
  assign n13201 = ~controllable_hmaster3 & ~n13200;
  assign n13202 = ~n13197 & ~n13201;
  assign n13203 = i_hbusreq7 & ~n13202;
  assign n13204 = i_hbusreq8 & ~n13196;
  assign n13205 = i_hbusreq6 & ~n13171;
  assign n13206 = controllable_hgrant5 & ~n8482;
  assign n13207 = i_hbusreq5 & ~n13164;
  assign n13208 = controllable_hgrant4 & ~n8480;
  assign n13209 = i_hbusreq4 & ~n13162;
  assign n13210 = i_hbusreq9 & ~n13162;
  assign n13211 = controllable_hgrant3 & ~n8476;
  assign n13212 = i_hbusreq3 & ~n13160;
  assign n13213 = controllable_hgrant1 & ~n8474;
  assign n13214 = i_hbusreq1 & ~n13158;
  assign n13215 = ~n7757 & ~n7928;
  assign n13216 = ~i_hbusreq0 & ~n12784;
  assign n13217 = ~n13052 & ~n13216;
  assign n13218 = ~i_hbusreq2 & ~n13217;
  assign n13219 = ~n13051 & ~n13218;
  assign n13220 = ~controllable_hgrant2 & ~n13219;
  assign n13221 = ~n7855 & ~n13220;
  assign n13222 = n7733 & ~n13221;
  assign n13223 = ~n13058 & ~n13222;
  assign n13224 = n7928 & ~n13223;
  assign n13225 = ~n13215 & ~n13224;
  assign n13226 = ~i_hbusreq1 & ~n13225;
  assign n13227 = ~n13214 & ~n13226;
  assign n13228 = ~controllable_hgrant1 & ~n13227;
  assign n13229 = ~n13213 & ~n13228;
  assign n13230 = ~i_hbusreq3 & ~n13229;
  assign n13231 = ~n13212 & ~n13230;
  assign n13232 = ~controllable_hgrant3 & ~n13231;
  assign n13233 = ~n13211 & ~n13232;
  assign n13234 = ~i_hbusreq9 & ~n13233;
  assign n13235 = ~n13210 & ~n13234;
  assign n13236 = ~i_hbusreq4 & ~n13235;
  assign n13237 = ~n13209 & ~n13236;
  assign n13238 = ~controllable_hgrant4 & ~n13237;
  assign n13239 = ~n13208 & ~n13238;
  assign n13240 = ~i_hbusreq5 & ~n13239;
  assign n13241 = ~n13207 & ~n13240;
  assign n13242 = ~controllable_hgrant5 & ~n13241;
  assign n13243 = ~n13206 & ~n13242;
  assign n13244 = controllable_hmaster1 & ~n13243;
  assign n13245 = controllable_hmaster2 & ~n13243;
  assign n13246 = ~n12942 & ~n13245;
  assign n13247 = ~controllable_hmaster1 & ~n13246;
  assign n13248 = ~n13244 & ~n13247;
  assign n13249 = ~i_hbusreq6 & ~n13248;
  assign n13250 = ~n13205 & ~n13249;
  assign n13251 = ~controllable_hgrant6 & ~n13250;
  assign n13252 = ~n13134 & ~n13251;
  assign n13253 = controllable_hmaster0 & ~n13252;
  assign n13254 = controllable_hgrant6 & ~n9029;
  assign n13255 = i_hbusreq6 & ~n13192;
  assign n13256 = controllable_hgrant5 & ~n9023;
  assign n13257 = i_hbusreq5 & ~n13186;
  assign n13258 = controllable_hgrant4 & ~n9021;
  assign n13259 = i_hbusreq4 & ~n13184;
  assign n13260 = i_hbusreq9 & ~n13184;
  assign n13261 = controllable_hgrant3 & ~n9017;
  assign n13262 = i_hbusreq3 & ~n13182;
  assign n13263 = controllable_hgrant1 & ~n9015;
  assign n13264 = i_hbusreq1 & ~n13180;
  assign n13265 = n7928 & ~n13224;
  assign n13266 = ~i_hbusreq1 & ~n13265;
  assign n13267 = ~n13264 & ~n13266;
  assign n13268 = ~controllable_hgrant1 & ~n13267;
  assign n13269 = ~n13263 & ~n13268;
  assign n13270 = ~i_hbusreq3 & ~n13269;
  assign n13271 = ~n13262 & ~n13270;
  assign n13272 = ~controllable_hgrant3 & ~n13271;
  assign n13273 = ~n13261 & ~n13272;
  assign n13274 = ~i_hbusreq9 & ~n13273;
  assign n13275 = ~n13260 & ~n13274;
  assign n13276 = ~i_hbusreq4 & ~n13275;
  assign n13277 = ~n13259 & ~n13276;
  assign n13278 = ~controllable_hgrant4 & ~n13277;
  assign n13279 = ~n13258 & ~n13278;
  assign n13280 = ~i_hbusreq5 & ~n13279;
  assign n13281 = ~n13257 & ~n13280;
  assign n13282 = ~controllable_hgrant5 & ~n13281;
  assign n13283 = ~n13256 & ~n13282;
  assign n13284 = ~controllable_hmaster2 & ~n13283;
  assign n13285 = ~n13245 & ~n13284;
  assign n13286 = ~controllable_hmaster1 & ~n13285;
  assign n13287 = ~n13244 & ~n13286;
  assign n13288 = ~i_hbusreq6 & ~n13287;
  assign n13289 = ~n13255 & ~n13288;
  assign n13290 = ~controllable_hgrant6 & ~n13289;
  assign n13291 = ~n13254 & ~n13290;
  assign n13292 = ~controllable_hmaster0 & ~n13291;
  assign n13293 = ~n13253 & ~n13292;
  assign n13294 = ~i_hbusreq8 & ~n13293;
  assign n13295 = ~n13204 & ~n13294;
  assign n13296 = controllable_hmaster3 & ~n13295;
  assign n13297 = i_hbusreq8 & ~n13200;
  assign n13298 = controllable_hgrant6 & ~n9038;
  assign n13299 = i_hbusreq6 & ~n13188;
  assign n13300 = ~i_hbusreq6 & ~n13283;
  assign n13301 = ~n13299 & ~n13300;
  assign n13302 = ~controllable_hgrant6 & ~n13301;
  assign n13303 = ~n13298 & ~n13302;
  assign n13304 = ~i_hbusreq8 & ~n13303;
  assign n13305 = ~n13297 & ~n13304;
  assign n13306 = ~controllable_hmaster3 & ~n13305;
  assign n13307 = ~n13296 & ~n13306;
  assign n13308 = ~i_hbusreq7 & ~n13307;
  assign n13309 = ~n13203 & ~n13308;
  assign n13310 = n7924 & ~n13309;
  assign n13311 = ~n13151 & ~n13310;
  assign n13312 = ~n8214 & ~n13311;
  assign n13313 = n7928 & ~n12630;
  assign n13314 = ~controllable_hgrant1 & ~n13313;
  assign n13315 = ~n13179 & ~n13314;
  assign n13316 = ~controllable_hgrant3 & ~n13315;
  assign n13317 = ~n13178 & ~n13316;
  assign n13318 = ~controllable_hgrant4 & ~n13317;
  assign n13319 = ~n13177 & ~n13318;
  assign n13320 = ~controllable_hgrant5 & ~n13319;
  assign n13321 = ~n13176 & ~n13320;
  assign n13322 = ~controllable_hmaster2 & ~n13321;
  assign n13323 = ~n8358 & ~n13322;
  assign n13324 = ~controllable_hmaster1 & ~n13323;
  assign n13325 = ~n8357 & ~n13324;
  assign n13326 = ~controllable_hgrant6 & ~n13325;
  assign n13327 = ~n13175 & ~n13326;
  assign n13328 = controllable_hmaster0 & ~n13327;
  assign n13329 = ~n9050 & ~n13328;
  assign n13330 = i_hlock8 & ~n13329;
  assign n13331 = ~n9056 & ~n13328;
  assign n13332 = ~i_hlock8 & ~n13331;
  assign n13333 = ~n13330 & ~n13332;
  assign n13334 = controllable_hmaster3 & ~n13333;
  assign n13335 = ~n8995 & ~n13334;
  assign n13336 = i_hbusreq7 & ~n13335;
  assign n13337 = i_hbusreq8 & ~n13333;
  assign n13338 = i_hbusreq6 & ~n13325;
  assign n13339 = i_hbusreq5 & ~n13319;
  assign n13340 = i_hbusreq4 & ~n13317;
  assign n13341 = i_hbusreq9 & ~n13317;
  assign n13342 = i_hbusreq3 & ~n13315;
  assign n13343 = i_hbusreq1 & ~n13313;
  assign n13344 = i_hbusreq0 & ~n12696;
  assign n13345 = ~i_hbusreq2 & ~n13344;
  assign n13346 = ~n12695 & ~n13345;
  assign n13347 = ~controllable_hgrant2 & ~n13346;
  assign n13348 = ~n7855 & ~n13347;
  assign n13349 = n7928 & ~n13348;
  assign n13350 = n7928 & ~n13349;
  assign n13351 = ~i_hbusreq1 & ~n13350;
  assign n13352 = ~n13343 & ~n13351;
  assign n13353 = ~controllable_hgrant1 & ~n13352;
  assign n13354 = ~n13263 & ~n13353;
  assign n13355 = ~i_hbusreq3 & ~n13354;
  assign n13356 = ~n13342 & ~n13355;
  assign n13357 = ~controllable_hgrant3 & ~n13356;
  assign n13358 = ~n13261 & ~n13357;
  assign n13359 = ~i_hbusreq9 & ~n13358;
  assign n13360 = ~n13341 & ~n13359;
  assign n13361 = ~i_hbusreq4 & ~n13360;
  assign n13362 = ~n13340 & ~n13361;
  assign n13363 = ~controllable_hgrant4 & ~n13362;
  assign n13364 = ~n13258 & ~n13363;
  assign n13365 = ~i_hbusreq5 & ~n13364;
  assign n13366 = ~n13339 & ~n13365;
  assign n13367 = ~controllable_hgrant5 & ~n13366;
  assign n13368 = ~n13256 & ~n13367;
  assign n13369 = ~controllable_hmaster2 & ~n13368;
  assign n13370 = ~n8484 & ~n13369;
  assign n13371 = ~controllable_hmaster1 & ~n13370;
  assign n13372 = ~n8483 & ~n13371;
  assign n13373 = ~i_hbusreq6 & ~n13372;
  assign n13374 = ~n13338 & ~n13373;
  assign n13375 = ~controllable_hgrant6 & ~n13374;
  assign n13376 = ~n13254 & ~n13375;
  assign n13377 = controllable_hmaster0 & ~n13376;
  assign n13378 = ~n9071 & ~n13377;
  assign n13379 = i_hlock8 & ~n13378;
  assign n13380 = ~n9080 & ~n13377;
  assign n13381 = ~i_hlock8 & ~n13380;
  assign n13382 = ~n13379 & ~n13381;
  assign n13383 = ~i_hbusreq8 & ~n13382;
  assign n13384 = ~n13337 & ~n13383;
  assign n13385 = controllable_hmaster3 & ~n13384;
  assign n13386 = ~n9041 & ~n13385;
  assign n13387 = ~i_hbusreq7 & ~n13386;
  assign n13388 = ~n13336 & ~n13387;
  assign n13389 = ~n7924 & ~n13388;
  assign n13390 = n7928 & ~n12803;
  assign n13391 = ~controllable_hgrant1 & ~n13390;
  assign n13392 = ~n13179 & ~n13391;
  assign n13393 = ~controllable_hgrant3 & ~n13392;
  assign n13394 = ~n13178 & ~n13393;
  assign n13395 = ~controllable_hgrant4 & ~n13394;
  assign n13396 = ~n13177 & ~n13395;
  assign n13397 = ~controllable_hgrant5 & ~n13396;
  assign n13398 = ~n13176 & ~n13397;
  assign n13399 = ~controllable_hmaster2 & ~n13398;
  assign n13400 = ~n13168 & ~n13399;
  assign n13401 = ~controllable_hmaster1 & ~n13400;
  assign n13402 = ~n13167 & ~n13401;
  assign n13403 = ~controllable_hgrant6 & ~n13402;
  assign n13404 = ~n13175 & ~n13403;
  assign n13405 = controllable_hmaster0 & ~n13404;
  assign n13406 = controllable_hgrant6 & ~n9049;
  assign n13407 = controllable_hgrant5 & ~n8653;
  assign n13408 = controllable_hgrant4 & ~n8653;
  assign n13409 = ~n8221 & ~n13157;
  assign n13410 = ~controllable_hgrant1 & ~n13409;
  assign n13411 = ~n12611 & ~n13410;
  assign n13412 = ~controllable_hgrant3 & ~n13411;
  assign n13413 = ~n12610 & ~n13412;
  assign n13414 = ~controllable_hgrant4 & ~n13413;
  assign n13415 = ~n13408 & ~n13414;
  assign n13416 = ~controllable_hgrant5 & ~n13415;
  assign n13417 = ~n13407 & ~n13416;
  assign n13418 = ~controllable_hmaster2 & ~n13417;
  assign n13419 = ~n13168 & ~n13418;
  assign n13420 = ~controllable_hmaster1 & ~n13419;
  assign n13421 = ~n13167 & ~n13420;
  assign n13422 = ~controllable_hgrant6 & ~n13421;
  assign n13423 = ~n13406 & ~n13422;
  assign n13424 = ~controllable_hmaster0 & ~n13423;
  assign n13425 = ~n13405 & ~n13424;
  assign n13426 = i_hlock8 & ~n13425;
  assign n13427 = controllable_hgrant6 & ~n9055;
  assign n13428 = controllable_hgrant5 & ~n8655;
  assign n13429 = controllable_hgrant4 & ~n8655;
  assign n13430 = ~n8235 & ~n13157;
  assign n13431 = ~controllable_hgrant1 & ~n13430;
  assign n13432 = ~n12638 & ~n13431;
  assign n13433 = ~controllable_hgrant3 & ~n13432;
  assign n13434 = ~n12637 & ~n13433;
  assign n13435 = ~controllable_hgrant4 & ~n13434;
  assign n13436 = ~n13429 & ~n13435;
  assign n13437 = ~controllable_hgrant5 & ~n13436;
  assign n13438 = ~n13428 & ~n13437;
  assign n13439 = ~controllable_hmaster2 & ~n13438;
  assign n13440 = ~n13168 & ~n13439;
  assign n13441 = ~controllable_hmaster1 & ~n13440;
  assign n13442 = ~n13167 & ~n13441;
  assign n13443 = ~controllable_hgrant6 & ~n13442;
  assign n13444 = ~n13427 & ~n13443;
  assign n13445 = ~controllable_hmaster0 & ~n13444;
  assign n13446 = ~n13405 & ~n13445;
  assign n13447 = ~i_hlock8 & ~n13446;
  assign n13448 = ~n13426 & ~n13447;
  assign n13449 = controllable_hmaster3 & ~n13448;
  assign n13450 = ~n13201 & ~n13449;
  assign n13451 = i_hbusreq7 & ~n13450;
  assign n13452 = i_hbusreq8 & ~n13448;
  assign n13453 = i_hbusreq6 & ~n13402;
  assign n13454 = i_hbusreq0 & ~n13052;
  assign n13455 = ~i_hbusreq2 & ~n13454;
  assign n13456 = ~n13051 & ~n13455;
  assign n13457 = ~controllable_hgrant2 & ~n13456;
  assign n13458 = ~n7855 & ~n13457;
  assign n13459 = n7928 & ~n13458;
  assign n13460 = ~n13215 & ~n13459;
  assign n13461 = ~i_hbusreq1 & ~n13460;
  assign n13462 = ~n13214 & ~n13461;
  assign n13463 = ~controllable_hgrant1 & ~n13462;
  assign n13464 = ~n13213 & ~n13463;
  assign n13465 = ~i_hbusreq3 & ~n13464;
  assign n13466 = ~n13212 & ~n13465;
  assign n13467 = ~controllable_hgrant3 & ~n13466;
  assign n13468 = ~n13211 & ~n13467;
  assign n13469 = ~i_hbusreq9 & ~n13468;
  assign n13470 = ~n13210 & ~n13469;
  assign n13471 = ~i_hbusreq4 & ~n13470;
  assign n13472 = ~n13209 & ~n13471;
  assign n13473 = ~controllable_hgrant4 & ~n13472;
  assign n13474 = ~n13208 & ~n13473;
  assign n13475 = ~i_hbusreq5 & ~n13474;
  assign n13476 = ~n13207 & ~n13475;
  assign n13477 = ~controllable_hgrant5 & ~n13476;
  assign n13478 = ~n13206 & ~n13477;
  assign n13479 = controllable_hmaster1 & ~n13478;
  assign n13480 = controllable_hmaster2 & ~n13478;
  assign n13481 = i_hbusreq5 & ~n13396;
  assign n13482 = i_hbusreq4 & ~n13394;
  assign n13483 = i_hbusreq9 & ~n13394;
  assign n13484 = i_hbusreq3 & ~n13392;
  assign n13485 = i_hbusreq1 & ~n13390;
  assign n13486 = i_hbusreq0 & ~n12884;
  assign n13487 = ~i_hbusreq2 & ~n13486;
  assign n13488 = ~n12883 & ~n13487;
  assign n13489 = ~controllable_hgrant2 & ~n13488;
  assign n13490 = ~n7855 & ~n13489;
  assign n13491 = n7928 & ~n13490;
  assign n13492 = n7928 & ~n13491;
  assign n13493 = ~i_hbusreq1 & ~n13492;
  assign n13494 = ~n13485 & ~n13493;
  assign n13495 = ~controllable_hgrant1 & ~n13494;
  assign n13496 = ~n13263 & ~n13495;
  assign n13497 = ~i_hbusreq3 & ~n13496;
  assign n13498 = ~n13484 & ~n13497;
  assign n13499 = ~controllable_hgrant3 & ~n13498;
  assign n13500 = ~n13261 & ~n13499;
  assign n13501 = ~i_hbusreq9 & ~n13500;
  assign n13502 = ~n13483 & ~n13501;
  assign n13503 = ~i_hbusreq4 & ~n13502;
  assign n13504 = ~n13482 & ~n13503;
  assign n13505 = ~controllable_hgrant4 & ~n13504;
  assign n13506 = ~n13258 & ~n13505;
  assign n13507 = ~i_hbusreq5 & ~n13506;
  assign n13508 = ~n13481 & ~n13507;
  assign n13509 = ~controllable_hgrant5 & ~n13508;
  assign n13510 = ~n13256 & ~n13509;
  assign n13511 = ~controllable_hmaster2 & ~n13510;
  assign n13512 = ~n13480 & ~n13511;
  assign n13513 = ~controllable_hmaster1 & ~n13512;
  assign n13514 = ~n13479 & ~n13513;
  assign n13515 = ~i_hbusreq6 & ~n13514;
  assign n13516 = ~n13453 & ~n13515;
  assign n13517 = ~controllable_hgrant6 & ~n13516;
  assign n13518 = ~n13254 & ~n13517;
  assign n13519 = controllable_hmaster0 & ~n13518;
  assign n13520 = controllable_hgrant6 & ~n9070;
  assign n13521 = i_hbusreq6 & ~n13421;
  assign n13522 = controllable_hgrant5 & ~n8754;
  assign n13523 = i_hbusreq5 & ~n13415;
  assign n13524 = controllable_hgrant4 & ~n8752;
  assign n13525 = i_hbusreq4 & ~n13413;
  assign n13526 = i_hbusreq9 & ~n13413;
  assign n13527 = i_hbusreq3 & ~n13411;
  assign n13528 = i_hbusreq1 & ~n13409;
  assign n13529 = ~n8676 & ~n13052;
  assign n13530 = ~i_hbusreq2 & ~n13529;
  assign n13531 = ~n13051 & ~n13530;
  assign n13532 = ~controllable_hgrant2 & ~n13531;
  assign n13533 = ~n12694 & ~n13532;
  assign n13534 = ~n7733 & ~n13533;
  assign n13535 = ~n8683 & ~n13052;
  assign n13536 = ~i_hbusreq2 & ~n13535;
  assign n13537 = ~n13051 & ~n13536;
  assign n13538 = ~controllable_hgrant2 & ~n13537;
  assign n13539 = ~n12706 & ~n13538;
  assign n13540 = n7733 & ~n13539;
  assign n13541 = ~n13534 & ~n13540;
  assign n13542 = n7928 & ~n13541;
  assign n13543 = ~n8265 & ~n13542;
  assign n13544 = ~i_hbusreq1 & ~n13543;
  assign n13545 = ~n13528 & ~n13544;
  assign n13546 = ~controllable_hgrant1 & ~n13545;
  assign n13547 = ~n12681 & ~n13546;
  assign n13548 = ~i_hbusreq3 & ~n13547;
  assign n13549 = ~n13527 & ~n13548;
  assign n13550 = ~controllable_hgrant3 & ~n13549;
  assign n13551 = ~n12679 & ~n13550;
  assign n13552 = ~i_hbusreq9 & ~n13551;
  assign n13553 = ~n13526 & ~n13552;
  assign n13554 = ~i_hbusreq4 & ~n13553;
  assign n13555 = ~n13525 & ~n13554;
  assign n13556 = ~controllable_hgrant4 & ~n13555;
  assign n13557 = ~n13524 & ~n13556;
  assign n13558 = ~i_hbusreq5 & ~n13557;
  assign n13559 = ~n13523 & ~n13558;
  assign n13560 = ~controllable_hgrant5 & ~n13559;
  assign n13561 = ~n13522 & ~n13560;
  assign n13562 = ~controllable_hmaster2 & ~n13561;
  assign n13563 = ~n13480 & ~n13562;
  assign n13564 = ~controllable_hmaster1 & ~n13563;
  assign n13565 = ~n13479 & ~n13564;
  assign n13566 = ~i_hbusreq6 & ~n13565;
  assign n13567 = ~n13521 & ~n13566;
  assign n13568 = ~controllable_hgrant6 & ~n13567;
  assign n13569 = ~n13520 & ~n13568;
  assign n13570 = ~controllable_hmaster0 & ~n13569;
  assign n13571 = ~n13519 & ~n13570;
  assign n13572 = i_hlock8 & ~n13571;
  assign n13573 = controllable_hgrant6 & ~n9079;
  assign n13574 = i_hbusreq6 & ~n13442;
  assign n13575 = controllable_hgrant5 & ~n8773;
  assign n13576 = i_hbusreq5 & ~n13436;
  assign n13577 = controllable_hgrant4 & ~n8771;
  assign n13578 = i_hbusreq4 & ~n13434;
  assign n13579 = i_hbusreq9 & ~n13434;
  assign n13580 = i_hbusreq3 & ~n13432;
  assign n13581 = i_hbusreq1 & ~n13430;
  assign n13582 = ~n8297 & ~n13542;
  assign n13583 = ~i_hbusreq1 & ~n13582;
  assign n13584 = ~n13581 & ~n13583;
  assign n13585 = ~controllable_hgrant1 & ~n13584;
  assign n13586 = ~n12730 & ~n13585;
  assign n13587 = ~i_hbusreq3 & ~n13586;
  assign n13588 = ~n13580 & ~n13587;
  assign n13589 = ~controllable_hgrant3 & ~n13588;
  assign n13590 = ~n12728 & ~n13589;
  assign n13591 = ~i_hbusreq9 & ~n13590;
  assign n13592 = ~n13579 & ~n13591;
  assign n13593 = ~i_hbusreq4 & ~n13592;
  assign n13594 = ~n13578 & ~n13593;
  assign n13595 = ~controllable_hgrant4 & ~n13594;
  assign n13596 = ~n13577 & ~n13595;
  assign n13597 = ~i_hbusreq5 & ~n13596;
  assign n13598 = ~n13576 & ~n13597;
  assign n13599 = ~controllable_hgrant5 & ~n13598;
  assign n13600 = ~n13575 & ~n13599;
  assign n13601 = ~controllable_hmaster2 & ~n13600;
  assign n13602 = ~n13480 & ~n13601;
  assign n13603 = ~controllable_hmaster1 & ~n13602;
  assign n13604 = ~n13479 & ~n13603;
  assign n13605 = ~i_hbusreq6 & ~n13604;
  assign n13606 = ~n13574 & ~n13605;
  assign n13607 = ~controllable_hgrant6 & ~n13606;
  assign n13608 = ~n13573 & ~n13607;
  assign n13609 = ~controllable_hmaster0 & ~n13608;
  assign n13610 = ~n13519 & ~n13609;
  assign n13611 = ~i_hlock8 & ~n13610;
  assign n13612 = ~n13572 & ~n13611;
  assign n13613 = ~i_hbusreq8 & ~n13612;
  assign n13614 = ~n13452 & ~n13613;
  assign n13615 = controllable_hmaster3 & ~n13614;
  assign n13616 = n7928 & ~n13459;
  assign n13617 = ~i_hbusreq1 & ~n13616;
  assign n13618 = ~n13264 & ~n13617;
  assign n13619 = ~controllable_hgrant1 & ~n13618;
  assign n13620 = ~n13263 & ~n13619;
  assign n13621 = ~i_hbusreq3 & ~n13620;
  assign n13622 = ~n13262 & ~n13621;
  assign n13623 = ~controllable_hgrant3 & ~n13622;
  assign n13624 = ~n13261 & ~n13623;
  assign n13625 = ~i_hbusreq9 & ~n13624;
  assign n13626 = ~n13260 & ~n13625;
  assign n13627 = ~i_hbusreq4 & ~n13626;
  assign n13628 = ~n13259 & ~n13627;
  assign n13629 = ~controllable_hgrant4 & ~n13628;
  assign n13630 = ~n13258 & ~n13629;
  assign n13631 = ~i_hbusreq5 & ~n13630;
  assign n13632 = ~n13257 & ~n13631;
  assign n13633 = ~controllable_hgrant5 & ~n13632;
  assign n13634 = ~n13256 & ~n13633;
  assign n13635 = ~i_hbusreq6 & ~n13634;
  assign n13636 = ~n13299 & ~n13635;
  assign n13637 = ~controllable_hgrant6 & ~n13636;
  assign n13638 = ~n13298 & ~n13637;
  assign n13639 = ~i_hbusreq8 & ~n13638;
  assign n13640 = ~n13297 & ~n13639;
  assign n13641 = ~controllable_hmaster3 & ~n13640;
  assign n13642 = ~n13615 & ~n13641;
  assign n13643 = ~i_hbusreq7 & ~n13642;
  assign n13644 = ~n13451 & ~n13643;
  assign n13645 = n7924 & ~n13644;
  assign n13646 = ~n13389 & ~n13645;
  assign n13647 = n8214 & ~n13646;
  assign n13648 = ~n13312 & ~n13647;
  assign n13649 = ~n8202 & ~n13648;
  assign n13650 = ~n8992 & ~n13328;
  assign n13651 = controllable_hmaster3 & ~n13650;
  assign n13652 = ~n9101 & ~n13651;
  assign n13653 = i_hlock7 & ~n13652;
  assign n13654 = ~n9109 & ~n13651;
  assign n13655 = ~i_hlock7 & ~n13654;
  assign n13656 = ~n13653 & ~n13655;
  assign n13657 = i_hbusreq7 & ~n13656;
  assign n13658 = i_hbusreq8 & ~n13650;
  assign n13659 = ~n9030 & ~n13377;
  assign n13660 = ~i_hbusreq8 & ~n13659;
  assign n13661 = ~n13658 & ~n13660;
  assign n13662 = controllable_hmaster3 & ~n13661;
  assign n13663 = ~n9131 & ~n13662;
  assign n13664 = i_hlock7 & ~n13663;
  assign n13665 = ~n9145 & ~n13662;
  assign n13666 = ~i_hlock7 & ~n13665;
  assign n13667 = ~n13664 & ~n13666;
  assign n13668 = ~i_hbusreq7 & ~n13667;
  assign n13669 = ~n13657 & ~n13668;
  assign n13670 = ~n7924 & ~n13669;
  assign n13671 = ~n13195 & ~n13405;
  assign n13672 = controllable_hmaster3 & ~n13671;
  assign n13673 = controllable_hgrant6 & ~n9097;
  assign n13674 = controllable_hmaster2 & ~n13417;
  assign n13675 = ~n13189 & ~n13674;
  assign n13676 = controllable_hmaster1 & ~n13675;
  assign n13677 = ~controllable_hmaster1 & ~n13188;
  assign n13678 = ~n13676 & ~n13677;
  assign n13679 = ~controllable_hgrant6 & ~n13678;
  assign n13680 = ~n13673 & ~n13679;
  assign n13681 = controllable_hmaster0 & ~n13680;
  assign n13682 = ~controllable_hmaster0 & ~n13200;
  assign n13683 = ~n13681 & ~n13682;
  assign n13684 = ~controllable_hmaster3 & ~n13683;
  assign n13685 = ~n13672 & ~n13684;
  assign n13686 = i_hlock7 & ~n13685;
  assign n13687 = controllable_hgrant6 & ~n9106;
  assign n13688 = controllable_hmaster2 & ~n13438;
  assign n13689 = ~n13189 & ~n13688;
  assign n13690 = controllable_hmaster1 & ~n13689;
  assign n13691 = ~n13677 & ~n13690;
  assign n13692 = ~controllable_hgrant6 & ~n13691;
  assign n13693 = ~n13687 & ~n13692;
  assign n13694 = controllable_hmaster0 & ~n13693;
  assign n13695 = ~n13682 & ~n13694;
  assign n13696 = ~controllable_hmaster3 & ~n13695;
  assign n13697 = ~n13672 & ~n13696;
  assign n13698 = ~i_hlock7 & ~n13697;
  assign n13699 = ~n13686 & ~n13698;
  assign n13700 = i_hbusreq7 & ~n13699;
  assign n13701 = i_hbusreq8 & ~n13671;
  assign n13702 = ~controllable_hmaster2 & ~n13634;
  assign n13703 = ~n13480 & ~n13702;
  assign n13704 = ~controllable_hmaster1 & ~n13703;
  assign n13705 = ~n13479 & ~n13704;
  assign n13706 = ~i_hbusreq6 & ~n13705;
  assign n13707 = ~n13255 & ~n13706;
  assign n13708 = ~controllable_hgrant6 & ~n13707;
  assign n13709 = ~n13254 & ~n13708;
  assign n13710 = ~controllable_hmaster0 & ~n13709;
  assign n13711 = ~n13519 & ~n13710;
  assign n13712 = ~i_hbusreq8 & ~n13711;
  assign n13713 = ~n13701 & ~n13712;
  assign n13714 = controllable_hmaster3 & ~n13713;
  assign n13715 = i_hbusreq8 & ~n13683;
  assign n13716 = controllable_hgrant6 & ~n9125;
  assign n13717 = i_hbusreq6 & ~n13678;
  assign n13718 = controllable_hmaster2 & ~n13561;
  assign n13719 = ~n13702 & ~n13718;
  assign n13720 = controllable_hmaster1 & ~n13719;
  assign n13721 = ~controllable_hmaster1 & ~n13634;
  assign n13722 = ~n13720 & ~n13721;
  assign n13723 = ~i_hbusreq6 & ~n13722;
  assign n13724 = ~n13717 & ~n13723;
  assign n13725 = ~controllable_hgrant6 & ~n13724;
  assign n13726 = ~n13716 & ~n13725;
  assign n13727 = controllable_hmaster0 & ~n13726;
  assign n13728 = ~controllable_hmaster0 & ~n13638;
  assign n13729 = ~n13727 & ~n13728;
  assign n13730 = ~i_hbusreq8 & ~n13729;
  assign n13731 = ~n13715 & ~n13730;
  assign n13732 = ~controllable_hmaster3 & ~n13731;
  assign n13733 = ~n13714 & ~n13732;
  assign n13734 = i_hlock7 & ~n13733;
  assign n13735 = i_hbusreq8 & ~n13695;
  assign n13736 = controllable_hgrant6 & ~n9140;
  assign n13737 = i_hbusreq6 & ~n13691;
  assign n13738 = controllable_hmaster2 & ~n13600;
  assign n13739 = ~n13702 & ~n13738;
  assign n13740 = controllable_hmaster1 & ~n13739;
  assign n13741 = ~n13721 & ~n13740;
  assign n13742 = ~i_hbusreq6 & ~n13741;
  assign n13743 = ~n13737 & ~n13742;
  assign n13744 = ~controllable_hgrant6 & ~n13743;
  assign n13745 = ~n13736 & ~n13744;
  assign n13746 = controllable_hmaster0 & ~n13745;
  assign n13747 = ~n13728 & ~n13746;
  assign n13748 = ~i_hbusreq8 & ~n13747;
  assign n13749 = ~n13735 & ~n13748;
  assign n13750 = ~controllable_hmaster3 & ~n13749;
  assign n13751 = ~n13714 & ~n13750;
  assign n13752 = ~i_hlock7 & ~n13751;
  assign n13753 = ~n13734 & ~n13752;
  assign n13754 = ~i_hbusreq7 & ~n13753;
  assign n13755 = ~n13700 & ~n13754;
  assign n13756 = n7924 & ~n13755;
  assign n13757 = ~n13670 & ~n13756;
  assign n13758 = ~n8214 & ~n13757;
  assign n13759 = ~n9158 & ~n13651;
  assign n13760 = i_hbusreq7 & ~n13759;
  assign n13761 = ~n9173 & ~n13662;
  assign n13762 = ~i_hbusreq7 & ~n13761;
  assign n13763 = ~n13760 & ~n13762;
  assign n13764 = ~n7924 & ~n13763;
  assign n13765 = controllable_hmaster0 & ~n13200;
  assign n13766 = controllable_hgrant6 & ~n9155;
  assign n13767 = i_hlock6 & ~n13678;
  assign n13768 = ~i_hlock6 & ~n13691;
  assign n13769 = ~n13767 & ~n13768;
  assign n13770 = ~controllable_hgrant6 & ~n13769;
  assign n13771 = ~n13766 & ~n13770;
  assign n13772 = ~controllable_hmaster0 & ~n13771;
  assign n13773 = ~n13765 & ~n13772;
  assign n13774 = ~controllable_hmaster3 & ~n13773;
  assign n13775 = ~n13672 & ~n13774;
  assign n13776 = i_hbusreq7 & ~n13775;
  assign n13777 = i_hbusreq8 & ~n13773;
  assign n13778 = controllable_hmaster0 & ~n13638;
  assign n13779 = controllable_hgrant6 & ~n9168;
  assign n13780 = i_hbusreq6 & ~n13769;
  assign n13781 = i_hlock6 & ~n13722;
  assign n13782 = ~i_hlock6 & ~n13741;
  assign n13783 = ~n13781 & ~n13782;
  assign n13784 = ~i_hbusreq6 & ~n13783;
  assign n13785 = ~n13780 & ~n13784;
  assign n13786 = ~controllable_hgrant6 & ~n13785;
  assign n13787 = ~n13779 & ~n13786;
  assign n13788 = ~controllable_hmaster0 & ~n13787;
  assign n13789 = ~n13778 & ~n13788;
  assign n13790 = ~i_hbusreq8 & ~n13789;
  assign n13791 = ~n13777 & ~n13790;
  assign n13792 = ~controllable_hmaster3 & ~n13791;
  assign n13793 = ~n13714 & ~n13792;
  assign n13794 = ~i_hbusreq7 & ~n13793;
  assign n13795 = ~n13776 & ~n13794;
  assign n13796 = n7924 & ~n13795;
  assign n13797 = ~n13764 & ~n13796;
  assign n13798 = n8214 & ~n13797;
  assign n13799 = ~n13758 & ~n13798;
  assign n13800 = n8202 & ~n13799;
  assign n13801 = ~n13649 & ~n13800;
  assign n13802 = n7920 & ~n13801;
  assign n13803 = ~n8877 & ~n13802;
  assign n13804 = n7728 & ~n13803;
  assign n13805 = ~n9050 & ~n13128;
  assign n13806 = i_hlock8 & ~n13805;
  assign n13807 = ~n9056 & ~n13128;
  assign n13808 = ~i_hlock8 & ~n13807;
  assign n13809 = ~n13806 & ~n13808;
  assign n13810 = controllable_hmaster3 & ~n13809;
  assign n13811 = ~n9235 & ~n13810;
  assign n13812 = i_hlock7 & ~n13811;
  assign n13813 = ~n9243 & ~n13810;
  assign n13814 = ~i_hlock7 & ~n13813;
  assign n13815 = ~n13812 & ~n13814;
  assign n13816 = i_hbusreq7 & ~n13815;
  assign n13817 = i_hbusreq8 & ~n13809;
  assign n13818 = controllable_hgrant6 & ~n9265;
  assign n13819 = ~n9260 & ~n12764;
  assign n13820 = ~controllable_hmaster1 & ~n13819;
  assign n13821 = ~n9259 & ~n13820;
  assign n13822 = ~i_hbusreq6 & ~n13821;
  assign n13823 = ~n13135 & ~n13822;
  assign n13824 = ~controllable_hgrant6 & ~n13823;
  assign n13825 = ~n13818 & ~n13824;
  assign n13826 = controllable_hmaster0 & ~n13825;
  assign n13827 = ~n9285 & ~n13826;
  assign n13828 = i_hlock8 & ~n13827;
  assign n13829 = ~n9305 & ~n13826;
  assign n13830 = ~i_hlock8 & ~n13829;
  assign n13831 = ~n13828 & ~n13830;
  assign n13832 = ~i_hbusreq8 & ~n13831;
  assign n13833 = ~n13817 & ~n13832;
  assign n13834 = controllable_hmaster3 & ~n13833;
  assign n13835 = ~n9443 & ~n13834;
  assign n13836 = i_hlock7 & ~n13835;
  assign n13837 = ~n9457 & ~n13834;
  assign n13838 = ~i_hlock7 & ~n13837;
  assign n13839 = ~n13836 & ~n13838;
  assign n13840 = ~i_hbusreq7 & ~n13839;
  assign n13841 = ~n13816 & ~n13840;
  assign n13842 = ~n7924 & ~n13841;
  assign n13843 = ~n13174 & ~n13424;
  assign n13844 = i_hlock8 & ~n13843;
  assign n13845 = ~n13174 & ~n13445;
  assign n13846 = ~i_hlock8 & ~n13845;
  assign n13847 = ~n13844 & ~n13846;
  assign n13848 = controllable_hmaster3 & ~n13847;
  assign n13849 = controllable_hgrant6 & ~n9206;
  assign n13850 = controllable_hgrant5 & ~n9192;
  assign n13851 = controllable_hgrant4 & ~n9192;
  assign n13852 = controllable_hgrant3 & ~n9192;
  assign n13853 = i_hlock3 & ~n13411;
  assign n13854 = ~i_hlock3 & ~n13432;
  assign n13855 = ~n13853 & ~n13854;
  assign n13856 = ~controllable_hgrant3 & ~n13855;
  assign n13857 = ~n13852 & ~n13856;
  assign n13858 = ~controllable_hgrant4 & ~n13857;
  assign n13859 = ~n13851 & ~n13858;
  assign n13860 = ~controllable_hgrant5 & ~n13859;
  assign n13861 = ~n13850 & ~n13860;
  assign n13862 = ~controllable_hmaster2 & ~n13861;
  assign n13863 = ~n13674 & ~n13862;
  assign n13864 = controllable_hmaster1 & ~n13863;
  assign n13865 = controllable_hgrant5 & ~n9198;
  assign n13866 = i_hlock5 & ~n13415;
  assign n13867 = ~i_hlock5 & ~n13436;
  assign n13868 = ~n13866 & ~n13867;
  assign n13869 = ~controllable_hgrant5 & ~n13868;
  assign n13870 = ~n13865 & ~n13869;
  assign n13871 = controllable_hmaster2 & ~n13870;
  assign n13872 = controllable_hgrant5 & ~n9202;
  assign n13873 = controllable_hgrant4 & ~n9202;
  assign n13874 = controllable_hgrant3 & ~n9202;
  assign n13875 = controllable_hgrant1 & ~n9202;
  assign n13876 = i_hlock1 & ~n13409;
  assign n13877 = ~i_hlock1 & ~n13430;
  assign n13878 = ~n13876 & ~n13877;
  assign n13879 = ~controllable_hgrant1 & ~n13878;
  assign n13880 = ~n13875 & ~n13879;
  assign n13881 = ~controllable_hgrant3 & ~n13880;
  assign n13882 = ~n13874 & ~n13881;
  assign n13883 = ~controllable_hgrant4 & ~n13882;
  assign n13884 = ~n13873 & ~n13883;
  assign n13885 = ~controllable_hgrant5 & ~n13884;
  assign n13886 = ~n13872 & ~n13885;
  assign n13887 = ~controllable_hmaster2 & ~n13886;
  assign n13888 = ~n13871 & ~n13887;
  assign n13889 = ~controllable_hmaster1 & ~n13888;
  assign n13890 = ~n13864 & ~n13889;
  assign n13891 = ~controllable_hgrant6 & ~n13890;
  assign n13892 = ~n13849 & ~n13891;
  assign n13893 = controllable_hmaster0 & ~n13892;
  assign n13894 = controllable_hgrant6 & ~n9232;
  assign n13895 = controllable_hgrant5 & ~n9214;
  assign n13896 = controllable_hgrant4 & ~n9214;
  assign n13897 = controllable_hgrant3 & ~n9214;
  assign n13898 = controllable_hgrant1 & ~n9214;
  assign n13899 = ~n9213 & ~n13157;
  assign n13900 = ~controllable_hgrant1 & ~n13899;
  assign n13901 = ~n13898 & ~n13900;
  assign n13902 = ~controllable_hgrant3 & ~n13901;
  assign n13903 = ~n13897 & ~n13902;
  assign n13904 = ~controllable_hgrant4 & ~n13903;
  assign n13905 = ~n13896 & ~n13904;
  assign n13906 = ~controllable_hgrant5 & ~n13905;
  assign n13907 = ~n13895 & ~n13906;
  assign n13908 = ~controllable_hmaster2 & ~n13907;
  assign n13909 = ~n13674 & ~n13908;
  assign n13910 = controllable_hmaster1 & ~n13909;
  assign n13911 = controllable_hgrant5 & ~n9220;
  assign n13912 = controllable_hgrant4 & ~n9220;
  assign n13913 = i_hlock4 & ~n13413;
  assign n13914 = ~i_hlock4 & ~n13434;
  assign n13915 = ~n13913 & ~n13914;
  assign n13916 = ~controllable_hgrant4 & ~n13915;
  assign n13917 = ~n13912 & ~n13916;
  assign n13918 = ~controllable_hgrant5 & ~n13917;
  assign n13919 = ~n13911 & ~n13918;
  assign n13920 = controllable_hmaster2 & ~n13919;
  assign n13921 = controllable_hgrant5 & ~n9222;
  assign n13922 = controllable_hgrant4 & ~n9222;
  assign n13923 = controllable_hgrant3 & ~n9222;
  assign n13924 = controllable_hgrant1 & ~n9222;
  assign n13925 = ~n8440 & ~n13157;
  assign n13926 = ~controllable_hgrant1 & ~n13925;
  assign n13927 = ~n13924 & ~n13926;
  assign n13928 = ~controllable_hgrant3 & ~n13927;
  assign n13929 = ~n13923 & ~n13928;
  assign n13930 = ~controllable_hgrant4 & ~n13929;
  assign n13931 = ~n13922 & ~n13930;
  assign n13932 = ~controllable_hgrant5 & ~n13931;
  assign n13933 = ~n13921 & ~n13932;
  assign n13934 = ~controllable_hmaster2 & ~n13933;
  assign n13935 = ~n13920 & ~n13934;
  assign n13936 = ~controllable_hmaster1 & ~n13935;
  assign n13937 = ~n13910 & ~n13936;
  assign n13938 = i_hlock6 & ~n13937;
  assign n13939 = ~n13688 & ~n13908;
  assign n13940 = controllable_hmaster1 & ~n13939;
  assign n13941 = ~n13936 & ~n13940;
  assign n13942 = ~i_hlock6 & ~n13941;
  assign n13943 = ~n13938 & ~n13942;
  assign n13944 = ~controllable_hgrant6 & ~n13943;
  assign n13945 = ~n13894 & ~n13944;
  assign n13946 = ~controllable_hmaster0 & ~n13945;
  assign n13947 = ~n13893 & ~n13946;
  assign n13948 = ~controllable_hmaster3 & ~n13947;
  assign n13949 = ~n13848 & ~n13948;
  assign n13950 = i_hlock7 & ~n13949;
  assign n13951 = controllable_hgrant6 & ~n9240;
  assign n13952 = ~n13688 & ~n13862;
  assign n13953 = controllable_hmaster1 & ~n13952;
  assign n13954 = ~n13889 & ~n13953;
  assign n13955 = ~controllable_hgrant6 & ~n13954;
  assign n13956 = ~n13951 & ~n13955;
  assign n13957 = controllable_hmaster0 & ~n13956;
  assign n13958 = ~n13946 & ~n13957;
  assign n13959 = ~controllable_hmaster3 & ~n13958;
  assign n13960 = ~n13848 & ~n13959;
  assign n13961 = ~i_hlock7 & ~n13960;
  assign n13962 = ~n13950 & ~n13961;
  assign n13963 = i_hbusreq7 & ~n13962;
  assign n13964 = i_hbusreq8 & ~n13847;
  assign n13965 = controllable_hgrant5 & ~n9258;
  assign n13966 = controllable_hgrant4 & ~n9256;
  assign n13967 = controllable_hgrant3 & ~n9252;
  assign n13968 = controllable_hgrant1 & ~n9250;
  assign n13969 = ~n7928 & ~n8679;
  assign n13970 = ~i_hlock0 & ~n13009;
  assign n13971 = ~i_hlock0 & ~n13970;
  assign n13972 = ~i_hbusreq0 & ~n13971;
  assign n13973 = ~n13052 & ~n13972;
  assign n13974 = ~i_hbusreq2 & ~n13973;
  assign n13975 = ~n13051 & ~n13974;
  assign n13976 = ~controllable_hgrant2 & ~n13975;
  assign n13977 = ~n12694 & ~n13976;
  assign n13978 = ~n7733 & ~n13977;
  assign n13979 = i_hlock0 & ~n12784;
  assign n13980 = ~n13970 & ~n13979;
  assign n13981 = ~i_hbusreq0 & ~n13980;
  assign n13982 = ~n13052 & ~n13981;
  assign n13983 = ~i_hbusreq2 & ~n13982;
  assign n13984 = ~n13051 & ~n13983;
  assign n13985 = ~controllable_hgrant2 & ~n13984;
  assign n13986 = ~n12694 & ~n13985;
  assign n13987 = n7733 & ~n13986;
  assign n13988 = ~n13978 & ~n13987;
  assign n13989 = n7928 & ~n13988;
  assign n13990 = ~n13969 & ~n13989;
  assign n13991 = ~i_hbusreq1 & ~n13990;
  assign n13992 = ~n13214 & ~n13991;
  assign n13993 = ~controllable_hgrant1 & ~n13992;
  assign n13994 = ~n13968 & ~n13993;
  assign n13995 = ~i_hbusreq3 & ~n13994;
  assign n13996 = ~n13212 & ~n13995;
  assign n13997 = ~controllable_hgrant3 & ~n13996;
  assign n13998 = ~n13967 & ~n13997;
  assign n13999 = ~i_hbusreq9 & ~n13998;
  assign n14000 = ~n13210 & ~n13999;
  assign n14001 = ~i_hbusreq4 & ~n14000;
  assign n14002 = ~n13209 & ~n14001;
  assign n14003 = ~controllable_hgrant4 & ~n14002;
  assign n14004 = ~n13966 & ~n14003;
  assign n14005 = ~i_hbusreq5 & ~n14004;
  assign n14006 = ~n13207 & ~n14005;
  assign n14007 = ~controllable_hgrant5 & ~n14006;
  assign n14008 = ~n13965 & ~n14007;
  assign n14009 = controllable_hmaster1 & ~n14008;
  assign n14010 = controllable_hmaster2 & ~n14008;
  assign n14011 = ~n12942 & ~n14010;
  assign n14012 = ~controllable_hmaster1 & ~n14011;
  assign n14013 = ~n14009 & ~n14012;
  assign n14014 = ~i_hbusreq6 & ~n14013;
  assign n14015 = ~n13205 & ~n14014;
  assign n14016 = ~controllable_hgrant6 & ~n14015;
  assign n14017 = ~n13818 & ~n14016;
  assign n14018 = controllable_hmaster0 & ~n14017;
  assign n14019 = controllable_hgrant6 & ~n9284;
  assign n14020 = controllable_hgrant5 & ~n9278;
  assign n14021 = controllable_hgrant4 & ~n9276;
  assign n14022 = controllable_hgrant3 & ~n9272;
  assign n14023 = controllable_hgrant1 & ~n9270;
  assign n14024 = ~n8265 & ~n13989;
  assign n14025 = ~i_hbusreq1 & ~n14024;
  assign n14026 = ~n13528 & ~n14025;
  assign n14027 = ~controllable_hgrant1 & ~n14026;
  assign n14028 = ~n14023 & ~n14027;
  assign n14029 = ~i_hbusreq3 & ~n14028;
  assign n14030 = ~n13527 & ~n14029;
  assign n14031 = ~controllable_hgrant3 & ~n14030;
  assign n14032 = ~n14022 & ~n14031;
  assign n14033 = ~i_hbusreq9 & ~n14032;
  assign n14034 = ~n13526 & ~n14033;
  assign n14035 = ~i_hbusreq4 & ~n14034;
  assign n14036 = ~n13525 & ~n14035;
  assign n14037 = ~controllable_hgrant4 & ~n14036;
  assign n14038 = ~n14021 & ~n14037;
  assign n14039 = ~i_hbusreq5 & ~n14038;
  assign n14040 = ~n13523 & ~n14039;
  assign n14041 = ~controllable_hgrant5 & ~n14040;
  assign n14042 = ~n14020 & ~n14041;
  assign n14043 = ~controllable_hmaster2 & ~n14042;
  assign n14044 = ~n14010 & ~n14043;
  assign n14045 = ~controllable_hmaster1 & ~n14044;
  assign n14046 = ~n14009 & ~n14045;
  assign n14047 = ~i_hbusreq6 & ~n14046;
  assign n14048 = ~n13521 & ~n14047;
  assign n14049 = ~controllable_hgrant6 & ~n14048;
  assign n14050 = ~n14019 & ~n14049;
  assign n14051 = ~controllable_hmaster0 & ~n14050;
  assign n14052 = ~n14018 & ~n14051;
  assign n14053 = i_hlock8 & ~n14052;
  assign n14054 = controllable_hgrant6 & ~n9304;
  assign n14055 = controllable_hgrant5 & ~n9298;
  assign n14056 = controllable_hgrant4 & ~n9296;
  assign n14057 = controllable_hgrant3 & ~n9292;
  assign n14058 = controllable_hgrant1 & ~n9290;
  assign n14059 = ~n8297 & ~n13989;
  assign n14060 = ~i_hbusreq1 & ~n14059;
  assign n14061 = ~n13581 & ~n14060;
  assign n14062 = ~controllable_hgrant1 & ~n14061;
  assign n14063 = ~n14058 & ~n14062;
  assign n14064 = ~i_hbusreq3 & ~n14063;
  assign n14065 = ~n13580 & ~n14064;
  assign n14066 = ~controllable_hgrant3 & ~n14065;
  assign n14067 = ~n14057 & ~n14066;
  assign n14068 = ~i_hbusreq9 & ~n14067;
  assign n14069 = ~n13579 & ~n14068;
  assign n14070 = ~i_hbusreq4 & ~n14069;
  assign n14071 = ~n13578 & ~n14070;
  assign n14072 = ~controllable_hgrant4 & ~n14071;
  assign n14073 = ~n14056 & ~n14072;
  assign n14074 = ~i_hbusreq5 & ~n14073;
  assign n14075 = ~n13576 & ~n14074;
  assign n14076 = ~controllable_hgrant5 & ~n14075;
  assign n14077 = ~n14055 & ~n14076;
  assign n14078 = ~controllable_hmaster2 & ~n14077;
  assign n14079 = ~n14010 & ~n14078;
  assign n14080 = ~controllable_hmaster1 & ~n14079;
  assign n14081 = ~n14009 & ~n14080;
  assign n14082 = ~i_hbusreq6 & ~n14081;
  assign n14083 = ~n13574 & ~n14082;
  assign n14084 = ~controllable_hgrant6 & ~n14083;
  assign n14085 = ~n14054 & ~n14084;
  assign n14086 = ~controllable_hmaster0 & ~n14085;
  assign n14087 = ~n14018 & ~n14086;
  assign n14088 = ~i_hlock8 & ~n14087;
  assign n14089 = ~n14053 & ~n14088;
  assign n14090 = ~i_hbusreq8 & ~n14089;
  assign n14091 = ~n13964 & ~n14090;
  assign n14092 = controllable_hmaster3 & ~n14091;
  assign n14093 = i_hbusreq8 & ~n13947;
  assign n14094 = controllable_hgrant6 & ~n9363;
  assign n14095 = i_hbusreq6 & ~n13890;
  assign n14096 = controllable_hmaster2 & ~n14042;
  assign n14097 = controllable_hgrant5 & ~n9329;
  assign n14098 = i_hbusreq5 & ~n13859;
  assign n14099 = controllable_hgrant4 & ~n9327;
  assign n14100 = i_hbusreq4 & ~n13857;
  assign n14101 = i_hbusreq9 & ~n13857;
  assign n14102 = controllable_hgrant3 & ~n9323;
  assign n14103 = i_hbusreq3 & ~n13855;
  assign n14104 = i_hlock3 & ~n14028;
  assign n14105 = ~i_hlock3 & ~n14063;
  assign n14106 = ~n14104 & ~n14105;
  assign n14107 = ~i_hbusreq3 & ~n14106;
  assign n14108 = ~n14103 & ~n14107;
  assign n14109 = ~controllable_hgrant3 & ~n14108;
  assign n14110 = ~n14102 & ~n14109;
  assign n14111 = ~i_hbusreq9 & ~n14110;
  assign n14112 = ~n14101 & ~n14111;
  assign n14113 = ~i_hbusreq4 & ~n14112;
  assign n14114 = ~n14100 & ~n14113;
  assign n14115 = ~controllable_hgrant4 & ~n14114;
  assign n14116 = ~n14099 & ~n14115;
  assign n14117 = ~i_hbusreq5 & ~n14116;
  assign n14118 = ~n14098 & ~n14117;
  assign n14119 = ~controllable_hgrant5 & ~n14118;
  assign n14120 = ~n14097 & ~n14119;
  assign n14121 = ~controllable_hmaster2 & ~n14120;
  assign n14122 = ~n14096 & ~n14121;
  assign n14123 = controllable_hmaster1 & ~n14122;
  assign n14124 = controllable_hgrant5 & ~n9338;
  assign n14125 = i_hbusreq5 & ~n13868;
  assign n14126 = i_hlock5 & ~n14038;
  assign n14127 = ~i_hlock5 & ~n14073;
  assign n14128 = ~n14126 & ~n14127;
  assign n14129 = ~i_hbusreq5 & ~n14128;
  assign n14130 = ~n14125 & ~n14129;
  assign n14131 = ~controllable_hgrant5 & ~n14130;
  assign n14132 = ~n14124 & ~n14131;
  assign n14133 = controllable_hmaster2 & ~n14132;
  assign n14134 = controllable_hgrant5 & ~n9357;
  assign n14135 = i_hbusreq5 & ~n13884;
  assign n14136 = controllable_hgrant4 & ~n9355;
  assign n14137 = i_hbusreq4 & ~n13882;
  assign n14138 = i_hbusreq9 & ~n13882;
  assign n14139 = controllable_hgrant3 & ~n9351;
  assign n14140 = i_hbusreq3 & ~n13880;
  assign n14141 = controllable_hgrant1 & ~n9349;
  assign n14142 = i_hbusreq1 & ~n13878;
  assign n14143 = i_hlock1 & ~n14024;
  assign n14144 = ~i_hlock1 & ~n14059;
  assign n14145 = ~n14143 & ~n14144;
  assign n14146 = ~i_hbusreq1 & ~n14145;
  assign n14147 = ~n14142 & ~n14146;
  assign n14148 = ~controllable_hgrant1 & ~n14147;
  assign n14149 = ~n14141 & ~n14148;
  assign n14150 = ~i_hbusreq3 & ~n14149;
  assign n14151 = ~n14140 & ~n14150;
  assign n14152 = ~controllable_hgrant3 & ~n14151;
  assign n14153 = ~n14139 & ~n14152;
  assign n14154 = ~i_hbusreq9 & ~n14153;
  assign n14155 = ~n14138 & ~n14154;
  assign n14156 = ~i_hbusreq4 & ~n14155;
  assign n14157 = ~n14137 & ~n14156;
  assign n14158 = ~controllable_hgrant4 & ~n14157;
  assign n14159 = ~n14136 & ~n14158;
  assign n14160 = ~i_hbusreq5 & ~n14159;
  assign n14161 = ~n14135 & ~n14160;
  assign n14162 = ~controllable_hgrant5 & ~n14161;
  assign n14163 = ~n14134 & ~n14162;
  assign n14164 = ~controllable_hmaster2 & ~n14163;
  assign n14165 = ~n14133 & ~n14164;
  assign n14166 = ~controllable_hmaster1 & ~n14165;
  assign n14167 = ~n14123 & ~n14166;
  assign n14168 = ~i_hbusreq6 & ~n14167;
  assign n14169 = ~n14095 & ~n14168;
  assign n14170 = ~controllable_hgrant6 & ~n14169;
  assign n14171 = ~n14094 & ~n14170;
  assign n14172 = controllable_hmaster0 & ~n14171;
  assign n14173 = controllable_hgrant6 & ~n9438;
  assign n14174 = i_hbusreq6 & ~n13943;
  assign n14175 = controllable_hgrant5 & ~n9390;
  assign n14176 = i_hbusreq5 & ~n13905;
  assign n14177 = controllable_hgrant4 & ~n9388;
  assign n14178 = i_hbusreq4 & ~n13903;
  assign n14179 = i_hbusreq9 & ~n13903;
  assign n14180 = controllable_hgrant3 & ~n9384;
  assign n14181 = i_hbusreq3 & ~n13901;
  assign n14182 = controllable_hgrant1 & ~n9382;
  assign n14183 = i_hbusreq1 & ~n13899;
  assign n14184 = ~n9379 & ~n13989;
  assign n14185 = ~i_hbusreq1 & ~n14184;
  assign n14186 = ~n14183 & ~n14185;
  assign n14187 = ~controllable_hgrant1 & ~n14186;
  assign n14188 = ~n14182 & ~n14187;
  assign n14189 = ~i_hbusreq3 & ~n14188;
  assign n14190 = ~n14181 & ~n14189;
  assign n14191 = ~controllable_hgrant3 & ~n14190;
  assign n14192 = ~n14180 & ~n14191;
  assign n14193 = ~i_hbusreq9 & ~n14192;
  assign n14194 = ~n14179 & ~n14193;
  assign n14195 = ~i_hbusreq4 & ~n14194;
  assign n14196 = ~n14178 & ~n14195;
  assign n14197 = ~controllable_hgrant4 & ~n14196;
  assign n14198 = ~n14177 & ~n14197;
  assign n14199 = ~i_hbusreq5 & ~n14198;
  assign n14200 = ~n14176 & ~n14199;
  assign n14201 = ~controllable_hgrant5 & ~n14200;
  assign n14202 = ~n14175 & ~n14201;
  assign n14203 = ~controllable_hmaster2 & ~n14202;
  assign n14204 = ~n14096 & ~n14203;
  assign n14205 = controllable_hmaster1 & ~n14204;
  assign n14206 = controllable_hgrant5 & ~n9402;
  assign n14207 = i_hbusreq5 & ~n13917;
  assign n14208 = controllable_hgrant4 & ~n9400;
  assign n14209 = i_hbusreq4 & ~n13915;
  assign n14210 = i_hlock4 & ~n14034;
  assign n14211 = ~i_hlock4 & ~n14069;
  assign n14212 = ~n14210 & ~n14211;
  assign n14213 = ~i_hbusreq4 & ~n14212;
  assign n14214 = ~n14209 & ~n14213;
  assign n14215 = ~controllable_hgrant4 & ~n14214;
  assign n14216 = ~n14208 & ~n14215;
  assign n14217 = ~i_hbusreq5 & ~n14216;
  assign n14218 = ~n14207 & ~n14217;
  assign n14219 = ~controllable_hgrant5 & ~n14218;
  assign n14220 = ~n14206 & ~n14219;
  assign n14221 = controllable_hmaster2 & ~n14220;
  assign n14222 = controllable_hgrant5 & ~n9425;
  assign n14223 = i_hbusreq5 & ~n13931;
  assign n14224 = controllable_hgrant4 & ~n9423;
  assign n14225 = i_hbusreq4 & ~n13929;
  assign n14226 = i_hbusreq9 & ~n13929;
  assign n14227 = controllable_hgrant3 & ~n9419;
  assign n14228 = i_hbusreq3 & ~n13927;
  assign n14229 = controllable_hgrant1 & ~n9417;
  assign n14230 = i_hbusreq1 & ~n13925;
  assign n14231 = controllable_hgrant2 & ~n9413;
  assign n14232 = ~n8435 & ~n13970;
  assign n14233 = ~i_hbusreq0 & ~n14232;
  assign n14234 = ~n13052 & ~n14233;
  assign n14235 = ~i_hbusreq2 & ~n14234;
  assign n14236 = ~n13051 & ~n14235;
  assign n14237 = ~controllable_hgrant2 & ~n14236;
  assign n14238 = ~n14231 & ~n14237;
  assign n14239 = ~n7733 & ~n14238;
  assign n14240 = controllable_locked & ~n8218;
  assign n14241 = ~controllable_hmastlock & ~n12782;
  assign n14242 = ~n7858 & ~n14241;
  assign n14243 = ~controllable_locked & ~n14242;
  assign n14244 = ~n14240 & ~n14243;
  assign n14245 = i_hlock0 & ~n14244;
  assign n14246 = ~n13970 & ~n14245;
  assign n14247 = ~i_hbusreq0 & ~n14246;
  assign n14248 = ~n13052 & ~n14247;
  assign n14249 = ~i_hbusreq2 & ~n14248;
  assign n14250 = ~n13051 & ~n14249;
  assign n14251 = ~controllable_hgrant2 & ~n14250;
  assign n14252 = ~n14231 & ~n14251;
  assign n14253 = n7733 & ~n14252;
  assign n14254 = ~n14239 & ~n14253;
  assign n14255 = n7928 & ~n14254;
  assign n14256 = ~n8440 & ~n14255;
  assign n14257 = ~i_hbusreq1 & ~n14256;
  assign n14258 = ~n14230 & ~n14257;
  assign n14259 = ~controllable_hgrant1 & ~n14258;
  assign n14260 = ~n14229 & ~n14259;
  assign n14261 = ~i_hbusreq3 & ~n14260;
  assign n14262 = ~n14228 & ~n14261;
  assign n14263 = ~controllable_hgrant3 & ~n14262;
  assign n14264 = ~n14227 & ~n14263;
  assign n14265 = ~i_hbusreq9 & ~n14264;
  assign n14266 = ~n14226 & ~n14265;
  assign n14267 = ~i_hbusreq4 & ~n14266;
  assign n14268 = ~n14225 & ~n14267;
  assign n14269 = ~controllable_hgrant4 & ~n14268;
  assign n14270 = ~n14224 & ~n14269;
  assign n14271 = ~i_hbusreq5 & ~n14270;
  assign n14272 = ~n14223 & ~n14271;
  assign n14273 = ~controllable_hgrant5 & ~n14272;
  assign n14274 = ~n14222 & ~n14273;
  assign n14275 = ~controllable_hmaster2 & ~n14274;
  assign n14276 = ~n14221 & ~n14275;
  assign n14277 = ~controllable_hmaster1 & ~n14276;
  assign n14278 = ~n14205 & ~n14277;
  assign n14279 = i_hlock6 & ~n14278;
  assign n14280 = controllable_hmaster2 & ~n14077;
  assign n14281 = ~n14203 & ~n14280;
  assign n14282 = controllable_hmaster1 & ~n14281;
  assign n14283 = ~n14277 & ~n14282;
  assign n14284 = ~i_hlock6 & ~n14283;
  assign n14285 = ~n14279 & ~n14284;
  assign n14286 = ~i_hbusreq6 & ~n14285;
  assign n14287 = ~n14174 & ~n14286;
  assign n14288 = ~controllable_hgrant6 & ~n14287;
  assign n14289 = ~n14173 & ~n14288;
  assign n14290 = ~controllable_hmaster0 & ~n14289;
  assign n14291 = ~n14172 & ~n14290;
  assign n14292 = ~i_hbusreq8 & ~n14291;
  assign n14293 = ~n14093 & ~n14292;
  assign n14294 = ~controllable_hmaster3 & ~n14293;
  assign n14295 = ~n14092 & ~n14294;
  assign n14296 = i_hlock7 & ~n14295;
  assign n14297 = i_hbusreq8 & ~n13958;
  assign n14298 = controllable_hgrant6 & ~n9452;
  assign n14299 = i_hbusreq6 & ~n13954;
  assign n14300 = ~n14121 & ~n14280;
  assign n14301 = controllable_hmaster1 & ~n14300;
  assign n14302 = ~n14166 & ~n14301;
  assign n14303 = ~i_hbusreq6 & ~n14302;
  assign n14304 = ~n14299 & ~n14303;
  assign n14305 = ~controllable_hgrant6 & ~n14304;
  assign n14306 = ~n14298 & ~n14305;
  assign n14307 = controllable_hmaster0 & ~n14306;
  assign n14308 = ~n14290 & ~n14307;
  assign n14309 = ~i_hbusreq8 & ~n14308;
  assign n14310 = ~n14297 & ~n14309;
  assign n14311 = ~controllable_hmaster3 & ~n14310;
  assign n14312 = ~n14092 & ~n14311;
  assign n14313 = ~i_hlock7 & ~n14312;
  assign n14314 = ~n14296 & ~n14313;
  assign n14315 = ~i_hbusreq7 & ~n14314;
  assign n14316 = ~n13963 & ~n14315;
  assign n14317 = n7924 & ~n14316;
  assign n14318 = ~n13842 & ~n14317;
  assign n14319 = ~n8214 & ~n14318;
  assign n14320 = controllable_hgrant6 & ~n9478;
  assign n14321 = controllable_hgrant5 & ~n9472;
  assign n14322 = controllable_hgrant4 & ~n9470;
  assign n14323 = n7928 & ~n12704;
  assign n14324 = ~n12693 & ~n14323;
  assign n14325 = ~i_hbusreq1 & ~n14324;
  assign n14326 = ~n12682 & ~n14325;
  assign n14327 = ~controllable_hgrant1 & ~n14326;
  assign n14328 = ~n14023 & ~n14327;
  assign n14329 = ~i_hbusreq3 & ~n14328;
  assign n14330 = ~n12680 & ~n14329;
  assign n14331 = ~controllable_hgrant3 & ~n14330;
  assign n14332 = ~n14022 & ~n14331;
  assign n14333 = i_hlock9 & ~n14332;
  assign n14334 = ~n12742 & ~n14323;
  assign n14335 = ~i_hbusreq1 & ~n14334;
  assign n14336 = ~n12731 & ~n14335;
  assign n14337 = ~controllable_hgrant1 & ~n14336;
  assign n14338 = ~n14058 & ~n14337;
  assign n14339 = ~i_hbusreq3 & ~n14338;
  assign n14340 = ~n12729 & ~n14339;
  assign n14341 = ~controllable_hgrant3 & ~n14340;
  assign n14342 = ~n14057 & ~n14341;
  assign n14343 = ~i_hlock9 & ~n14342;
  assign n14344 = ~n14333 & ~n14343;
  assign n14345 = ~i_hbusreq9 & ~n14344;
  assign n14346 = ~n12678 & ~n14345;
  assign n14347 = ~i_hbusreq4 & ~n14346;
  assign n14348 = ~n12677 & ~n14347;
  assign n14349 = ~controllable_hgrant4 & ~n14348;
  assign n14350 = ~n14322 & ~n14349;
  assign n14351 = ~i_hbusreq5 & ~n14350;
  assign n14352 = ~n12675 & ~n14351;
  assign n14353 = ~controllable_hgrant5 & ~n14352;
  assign n14354 = ~n14321 & ~n14353;
  assign n14355 = ~controllable_hmaster2 & ~n14354;
  assign n14356 = ~n9260 & ~n14355;
  assign n14357 = ~controllable_hmaster1 & ~n14356;
  assign n14358 = ~n9259 & ~n14357;
  assign n14359 = ~i_hbusreq6 & ~n14358;
  assign n14360 = ~n13135 & ~n14359;
  assign n14361 = ~controllable_hgrant6 & ~n14360;
  assign n14362 = ~n14320 & ~n14361;
  assign n14363 = controllable_hmaster0 & ~n14362;
  assign n14364 = ~n9485 & ~n14363;
  assign n14365 = i_hlock8 & ~n14364;
  assign n14366 = ~n9493 & ~n14363;
  assign n14367 = ~i_hlock8 & ~n14366;
  assign n14368 = ~n14365 & ~n14367;
  assign n14369 = ~i_hbusreq8 & ~n14368;
  assign n14370 = ~n13817 & ~n14369;
  assign n14371 = controllable_hmaster3 & ~n14370;
  assign n14372 = ~n9443 & ~n14371;
  assign n14373 = i_hlock7 & ~n14372;
  assign n14374 = ~n9457 & ~n14371;
  assign n14375 = ~i_hlock7 & ~n14374;
  assign n14376 = ~n14373 & ~n14375;
  assign n14377 = ~i_hbusreq7 & ~n14376;
  assign n14378 = ~n13816 & ~n14377;
  assign n14379 = ~n7924 & ~n14378;
  assign n14380 = n7928 & ~n13977;
  assign n14381 = ~n13969 & ~n14380;
  assign n14382 = ~i_hbusreq1 & ~n14381;
  assign n14383 = ~n13214 & ~n14382;
  assign n14384 = ~controllable_hgrant1 & ~n14383;
  assign n14385 = ~n13968 & ~n14384;
  assign n14386 = ~i_hbusreq3 & ~n14385;
  assign n14387 = ~n13212 & ~n14386;
  assign n14388 = ~controllable_hgrant3 & ~n14387;
  assign n14389 = ~n13967 & ~n14388;
  assign n14390 = ~i_hbusreq9 & ~n14389;
  assign n14391 = ~n13210 & ~n14390;
  assign n14392 = ~i_hbusreq4 & ~n14391;
  assign n14393 = ~n13209 & ~n14392;
  assign n14394 = ~controllable_hgrant4 & ~n14393;
  assign n14395 = ~n13966 & ~n14394;
  assign n14396 = ~i_hbusreq5 & ~n14395;
  assign n14397 = ~n13207 & ~n14396;
  assign n14398 = ~controllable_hgrant5 & ~n14397;
  assign n14399 = ~n13965 & ~n14398;
  assign n14400 = controllable_hmaster1 & ~n14399;
  assign n14401 = controllable_hmaster2 & ~n14399;
  assign n14402 = n7928 & ~n12892;
  assign n14403 = ~n12693 & ~n14402;
  assign n14404 = ~i_hbusreq1 & ~n14403;
  assign n14405 = ~n12882 & ~n14404;
  assign n14406 = ~controllable_hgrant1 & ~n14405;
  assign n14407 = ~n14023 & ~n14406;
  assign n14408 = ~i_hbusreq3 & ~n14407;
  assign n14409 = ~n12881 & ~n14408;
  assign n14410 = ~controllable_hgrant3 & ~n14409;
  assign n14411 = ~n14022 & ~n14410;
  assign n14412 = i_hlock9 & ~n14411;
  assign n14413 = ~n12742 & ~n14402;
  assign n14414 = ~i_hbusreq1 & ~n14413;
  assign n14415 = ~n12920 & ~n14414;
  assign n14416 = ~controllable_hgrant1 & ~n14415;
  assign n14417 = ~n14058 & ~n14416;
  assign n14418 = ~i_hbusreq3 & ~n14417;
  assign n14419 = ~n12919 & ~n14418;
  assign n14420 = ~controllable_hgrant3 & ~n14419;
  assign n14421 = ~n14057 & ~n14420;
  assign n14422 = ~i_hlock9 & ~n14421;
  assign n14423 = ~n14412 & ~n14422;
  assign n14424 = ~i_hbusreq9 & ~n14423;
  assign n14425 = ~n12880 & ~n14424;
  assign n14426 = ~i_hbusreq4 & ~n14425;
  assign n14427 = ~n12879 & ~n14426;
  assign n14428 = ~controllable_hgrant4 & ~n14427;
  assign n14429 = ~n14322 & ~n14428;
  assign n14430 = ~i_hbusreq5 & ~n14429;
  assign n14431 = ~n12878 & ~n14430;
  assign n14432 = ~controllable_hgrant5 & ~n14431;
  assign n14433 = ~n14321 & ~n14432;
  assign n14434 = ~controllable_hmaster2 & ~n14433;
  assign n14435 = ~n14401 & ~n14434;
  assign n14436 = ~controllable_hmaster1 & ~n14435;
  assign n14437 = ~n14400 & ~n14436;
  assign n14438 = ~i_hbusreq6 & ~n14437;
  assign n14439 = ~n13205 & ~n14438;
  assign n14440 = ~controllable_hgrant6 & ~n14439;
  assign n14441 = ~n14320 & ~n14440;
  assign n14442 = controllable_hmaster0 & ~n14441;
  assign n14443 = controllable_hgrant6 & ~n9484;
  assign n14444 = ~n8681 & ~n13970;
  assign n14445 = ~i_hbusreq0 & ~n14444;
  assign n14446 = ~n13052 & ~n14445;
  assign n14447 = ~i_hbusreq2 & ~n14446;
  assign n14448 = ~n13051 & ~n14447;
  assign n14449 = ~controllable_hgrant2 & ~n14448;
  assign n14450 = ~n12706 & ~n14449;
  assign n14451 = n7733 & ~n14450;
  assign n14452 = ~n13978 & ~n14451;
  assign n14453 = n7928 & ~n14452;
  assign n14454 = ~n8265 & ~n14453;
  assign n14455 = ~i_hbusreq1 & ~n14454;
  assign n14456 = ~n13528 & ~n14455;
  assign n14457 = ~controllable_hgrant1 & ~n14456;
  assign n14458 = ~n12681 & ~n14457;
  assign n14459 = ~i_hbusreq3 & ~n14458;
  assign n14460 = ~n13527 & ~n14459;
  assign n14461 = ~controllable_hgrant3 & ~n14460;
  assign n14462 = ~n12679 & ~n14461;
  assign n14463 = ~i_hbusreq9 & ~n14462;
  assign n14464 = ~n13526 & ~n14463;
  assign n14465 = ~i_hbusreq4 & ~n14464;
  assign n14466 = ~n13525 & ~n14465;
  assign n14467 = ~controllable_hgrant4 & ~n14466;
  assign n14468 = ~n13524 & ~n14467;
  assign n14469 = ~i_hbusreq5 & ~n14468;
  assign n14470 = ~n13523 & ~n14469;
  assign n14471 = ~controllable_hgrant5 & ~n14470;
  assign n14472 = ~n13522 & ~n14471;
  assign n14473 = ~controllable_hmaster2 & ~n14472;
  assign n14474 = ~n14401 & ~n14473;
  assign n14475 = ~controllable_hmaster1 & ~n14474;
  assign n14476 = ~n14400 & ~n14475;
  assign n14477 = ~i_hbusreq6 & ~n14476;
  assign n14478 = ~n13521 & ~n14477;
  assign n14479 = ~controllable_hgrant6 & ~n14478;
  assign n14480 = ~n14443 & ~n14479;
  assign n14481 = ~controllable_hmaster0 & ~n14480;
  assign n14482 = ~n14442 & ~n14481;
  assign n14483 = i_hlock8 & ~n14482;
  assign n14484 = controllable_hgrant6 & ~n9492;
  assign n14485 = ~n8297 & ~n14453;
  assign n14486 = ~i_hbusreq1 & ~n14485;
  assign n14487 = ~n13581 & ~n14486;
  assign n14488 = ~controllable_hgrant1 & ~n14487;
  assign n14489 = ~n12730 & ~n14488;
  assign n14490 = ~i_hbusreq3 & ~n14489;
  assign n14491 = ~n13580 & ~n14490;
  assign n14492 = ~controllable_hgrant3 & ~n14491;
  assign n14493 = ~n12728 & ~n14492;
  assign n14494 = ~i_hbusreq9 & ~n14493;
  assign n14495 = ~n13579 & ~n14494;
  assign n14496 = ~i_hbusreq4 & ~n14495;
  assign n14497 = ~n13578 & ~n14496;
  assign n14498 = ~controllable_hgrant4 & ~n14497;
  assign n14499 = ~n13577 & ~n14498;
  assign n14500 = ~i_hbusreq5 & ~n14499;
  assign n14501 = ~n13576 & ~n14500;
  assign n14502 = ~controllable_hgrant5 & ~n14501;
  assign n14503 = ~n13575 & ~n14502;
  assign n14504 = ~controllable_hmaster2 & ~n14503;
  assign n14505 = ~n14401 & ~n14504;
  assign n14506 = ~controllable_hmaster1 & ~n14505;
  assign n14507 = ~n14400 & ~n14506;
  assign n14508 = ~i_hbusreq6 & ~n14507;
  assign n14509 = ~n13574 & ~n14508;
  assign n14510 = ~controllable_hgrant6 & ~n14509;
  assign n14511 = ~n14484 & ~n14510;
  assign n14512 = ~controllable_hmaster0 & ~n14511;
  assign n14513 = ~n14442 & ~n14512;
  assign n14514 = ~i_hlock8 & ~n14513;
  assign n14515 = ~n14483 & ~n14514;
  assign n14516 = ~i_hbusreq8 & ~n14515;
  assign n14517 = ~n13964 & ~n14516;
  assign n14518 = controllable_hmaster3 & ~n14517;
  assign n14519 = ~n8265 & ~n14380;
  assign n14520 = ~i_hbusreq1 & ~n14519;
  assign n14521 = ~n13528 & ~n14520;
  assign n14522 = ~controllable_hgrant1 & ~n14521;
  assign n14523 = ~n14023 & ~n14522;
  assign n14524 = ~i_hbusreq3 & ~n14523;
  assign n14525 = ~n13527 & ~n14524;
  assign n14526 = ~controllable_hgrant3 & ~n14525;
  assign n14527 = ~n14022 & ~n14526;
  assign n14528 = ~i_hbusreq9 & ~n14527;
  assign n14529 = ~n13526 & ~n14528;
  assign n14530 = ~i_hbusreq4 & ~n14529;
  assign n14531 = ~n13525 & ~n14530;
  assign n14532 = ~controllable_hgrant4 & ~n14531;
  assign n14533 = ~n14021 & ~n14532;
  assign n14534 = ~i_hbusreq5 & ~n14533;
  assign n14535 = ~n13523 & ~n14534;
  assign n14536 = ~controllable_hgrant5 & ~n14535;
  assign n14537 = ~n14020 & ~n14536;
  assign n14538 = controllable_hmaster2 & ~n14537;
  assign n14539 = i_hlock3 & ~n14523;
  assign n14540 = ~n8297 & ~n14380;
  assign n14541 = ~i_hbusreq1 & ~n14540;
  assign n14542 = ~n13581 & ~n14541;
  assign n14543 = ~controllable_hgrant1 & ~n14542;
  assign n14544 = ~n14058 & ~n14543;
  assign n14545 = ~i_hlock3 & ~n14544;
  assign n14546 = ~n14539 & ~n14545;
  assign n14547 = ~i_hbusreq3 & ~n14546;
  assign n14548 = ~n14103 & ~n14547;
  assign n14549 = ~controllable_hgrant3 & ~n14548;
  assign n14550 = ~n14102 & ~n14549;
  assign n14551 = ~i_hbusreq9 & ~n14550;
  assign n14552 = ~n14101 & ~n14551;
  assign n14553 = ~i_hbusreq4 & ~n14552;
  assign n14554 = ~n14100 & ~n14553;
  assign n14555 = ~controllable_hgrant4 & ~n14554;
  assign n14556 = ~n14099 & ~n14555;
  assign n14557 = ~i_hbusreq5 & ~n14556;
  assign n14558 = ~n14098 & ~n14557;
  assign n14559 = ~controllable_hgrant5 & ~n14558;
  assign n14560 = ~n14097 & ~n14559;
  assign n14561 = ~controllable_hmaster2 & ~n14560;
  assign n14562 = ~n14538 & ~n14561;
  assign n14563 = controllable_hmaster1 & ~n14562;
  assign n14564 = i_hlock5 & ~n14533;
  assign n14565 = ~i_hbusreq3 & ~n14544;
  assign n14566 = ~n13580 & ~n14565;
  assign n14567 = ~controllable_hgrant3 & ~n14566;
  assign n14568 = ~n14057 & ~n14567;
  assign n14569 = ~i_hbusreq9 & ~n14568;
  assign n14570 = ~n13579 & ~n14569;
  assign n14571 = ~i_hbusreq4 & ~n14570;
  assign n14572 = ~n13578 & ~n14571;
  assign n14573 = ~controllable_hgrant4 & ~n14572;
  assign n14574 = ~n14056 & ~n14573;
  assign n14575 = ~i_hlock5 & ~n14574;
  assign n14576 = ~n14564 & ~n14575;
  assign n14577 = ~i_hbusreq5 & ~n14576;
  assign n14578 = ~n14125 & ~n14577;
  assign n14579 = ~controllable_hgrant5 & ~n14578;
  assign n14580 = ~n14124 & ~n14579;
  assign n14581 = controllable_hmaster2 & ~n14580;
  assign n14582 = i_hlock1 & ~n14519;
  assign n14583 = ~i_hlock1 & ~n14540;
  assign n14584 = ~n14582 & ~n14583;
  assign n14585 = ~i_hbusreq1 & ~n14584;
  assign n14586 = ~n14142 & ~n14585;
  assign n14587 = ~controllable_hgrant1 & ~n14586;
  assign n14588 = ~n14141 & ~n14587;
  assign n14589 = ~i_hbusreq3 & ~n14588;
  assign n14590 = ~n14140 & ~n14589;
  assign n14591 = ~controllable_hgrant3 & ~n14590;
  assign n14592 = ~n14139 & ~n14591;
  assign n14593 = ~i_hbusreq9 & ~n14592;
  assign n14594 = ~n14138 & ~n14593;
  assign n14595 = ~i_hbusreq4 & ~n14594;
  assign n14596 = ~n14137 & ~n14595;
  assign n14597 = ~controllable_hgrant4 & ~n14596;
  assign n14598 = ~n14136 & ~n14597;
  assign n14599 = ~i_hbusreq5 & ~n14598;
  assign n14600 = ~n14135 & ~n14599;
  assign n14601 = ~controllable_hgrant5 & ~n14600;
  assign n14602 = ~n14134 & ~n14601;
  assign n14603 = ~controllable_hmaster2 & ~n14602;
  assign n14604 = ~n14581 & ~n14603;
  assign n14605 = ~controllable_hmaster1 & ~n14604;
  assign n14606 = ~n14563 & ~n14605;
  assign n14607 = ~i_hbusreq6 & ~n14606;
  assign n14608 = ~n14095 & ~n14607;
  assign n14609 = ~controllable_hgrant6 & ~n14608;
  assign n14610 = ~n14094 & ~n14609;
  assign n14611 = controllable_hmaster0 & ~n14610;
  assign n14612 = ~n9379 & ~n14380;
  assign n14613 = ~i_hbusreq1 & ~n14612;
  assign n14614 = ~n14183 & ~n14613;
  assign n14615 = ~controllable_hgrant1 & ~n14614;
  assign n14616 = ~n14182 & ~n14615;
  assign n14617 = ~i_hbusreq3 & ~n14616;
  assign n14618 = ~n14181 & ~n14617;
  assign n14619 = ~controllable_hgrant3 & ~n14618;
  assign n14620 = ~n14180 & ~n14619;
  assign n14621 = ~i_hbusreq9 & ~n14620;
  assign n14622 = ~n14179 & ~n14621;
  assign n14623 = ~i_hbusreq4 & ~n14622;
  assign n14624 = ~n14178 & ~n14623;
  assign n14625 = ~controllable_hgrant4 & ~n14624;
  assign n14626 = ~n14177 & ~n14625;
  assign n14627 = ~i_hbusreq5 & ~n14626;
  assign n14628 = ~n14176 & ~n14627;
  assign n14629 = ~controllable_hgrant5 & ~n14628;
  assign n14630 = ~n14175 & ~n14629;
  assign n14631 = ~controllable_hmaster2 & ~n14630;
  assign n14632 = ~n14538 & ~n14631;
  assign n14633 = controllable_hmaster1 & ~n14632;
  assign n14634 = i_hlock4 & ~n14529;
  assign n14635 = ~i_hlock4 & ~n14570;
  assign n14636 = ~n14634 & ~n14635;
  assign n14637 = ~i_hbusreq4 & ~n14636;
  assign n14638 = ~n14209 & ~n14637;
  assign n14639 = ~controllable_hgrant4 & ~n14638;
  assign n14640 = ~n14208 & ~n14639;
  assign n14641 = ~i_hbusreq5 & ~n14640;
  assign n14642 = ~n14207 & ~n14641;
  assign n14643 = ~controllable_hgrant5 & ~n14642;
  assign n14644 = ~n14206 & ~n14643;
  assign n14645 = controllable_hmaster2 & ~n14644;
  assign n14646 = n7928 & ~n14238;
  assign n14647 = ~n8440 & ~n14646;
  assign n14648 = ~i_hbusreq1 & ~n14647;
  assign n14649 = ~n14230 & ~n14648;
  assign n14650 = ~controllable_hgrant1 & ~n14649;
  assign n14651 = ~n14229 & ~n14650;
  assign n14652 = ~i_hbusreq3 & ~n14651;
  assign n14653 = ~n14228 & ~n14652;
  assign n14654 = ~controllable_hgrant3 & ~n14653;
  assign n14655 = ~n14227 & ~n14654;
  assign n14656 = ~i_hbusreq9 & ~n14655;
  assign n14657 = ~n14226 & ~n14656;
  assign n14658 = ~i_hbusreq4 & ~n14657;
  assign n14659 = ~n14225 & ~n14658;
  assign n14660 = ~controllable_hgrant4 & ~n14659;
  assign n14661 = ~n14224 & ~n14660;
  assign n14662 = ~i_hbusreq5 & ~n14661;
  assign n14663 = ~n14223 & ~n14662;
  assign n14664 = ~controllable_hgrant5 & ~n14663;
  assign n14665 = ~n14222 & ~n14664;
  assign n14666 = ~controllable_hmaster2 & ~n14665;
  assign n14667 = ~n14645 & ~n14666;
  assign n14668 = ~controllable_hmaster1 & ~n14667;
  assign n14669 = ~n14633 & ~n14668;
  assign n14670 = i_hlock6 & ~n14669;
  assign n14671 = ~i_hbusreq5 & ~n14574;
  assign n14672 = ~n13576 & ~n14671;
  assign n14673 = ~controllable_hgrant5 & ~n14672;
  assign n14674 = ~n14055 & ~n14673;
  assign n14675 = controllable_hmaster2 & ~n14674;
  assign n14676 = ~n14631 & ~n14675;
  assign n14677 = controllable_hmaster1 & ~n14676;
  assign n14678 = ~n14668 & ~n14677;
  assign n14679 = ~i_hlock6 & ~n14678;
  assign n14680 = ~n14670 & ~n14679;
  assign n14681 = ~i_hbusreq6 & ~n14680;
  assign n14682 = ~n14174 & ~n14681;
  assign n14683 = ~controllable_hgrant6 & ~n14682;
  assign n14684 = ~n14173 & ~n14683;
  assign n14685 = ~controllable_hmaster0 & ~n14684;
  assign n14686 = ~n14611 & ~n14685;
  assign n14687 = ~i_hbusreq8 & ~n14686;
  assign n14688 = ~n14093 & ~n14687;
  assign n14689 = ~controllable_hmaster3 & ~n14688;
  assign n14690 = ~n14518 & ~n14689;
  assign n14691 = i_hlock7 & ~n14690;
  assign n14692 = ~n14561 & ~n14675;
  assign n14693 = controllable_hmaster1 & ~n14692;
  assign n14694 = ~n14605 & ~n14693;
  assign n14695 = ~i_hbusreq6 & ~n14694;
  assign n14696 = ~n14299 & ~n14695;
  assign n14697 = ~controllable_hgrant6 & ~n14696;
  assign n14698 = ~n14298 & ~n14697;
  assign n14699 = controllable_hmaster0 & ~n14698;
  assign n14700 = ~n14685 & ~n14699;
  assign n14701 = ~i_hbusreq8 & ~n14700;
  assign n14702 = ~n14297 & ~n14701;
  assign n14703 = ~controllable_hmaster3 & ~n14702;
  assign n14704 = ~n14518 & ~n14703;
  assign n14705 = ~i_hlock7 & ~n14704;
  assign n14706 = ~n14691 & ~n14705;
  assign n14707 = ~i_hbusreq7 & ~n14706;
  assign n14708 = ~n13963 & ~n14707;
  assign n14709 = n7924 & ~n14708;
  assign n14710 = ~n14379 & ~n14709;
  assign n14711 = n8214 & ~n14710;
  assign n14712 = ~n14319 & ~n14711;
  assign n14713 = ~n8202 & ~n14712;
  assign n14714 = ~n9285 & ~n14363;
  assign n14715 = i_hlock8 & ~n14714;
  assign n14716 = ~n9305 & ~n14363;
  assign n14717 = ~i_hlock8 & ~n14716;
  assign n14718 = ~n14715 & ~n14717;
  assign n14719 = ~i_hbusreq8 & ~n14718;
  assign n14720 = ~n13817 & ~n14719;
  assign n14721 = controllable_hmaster3 & ~n14720;
  assign n14722 = ~n9527 & ~n14721;
  assign n14723 = i_hlock7 & ~n14722;
  assign n14724 = ~n9539 & ~n14721;
  assign n14725 = ~i_hlock7 & ~n14724;
  assign n14726 = ~n14723 & ~n14725;
  assign n14727 = ~i_hbusreq7 & ~n14726;
  assign n14728 = ~n13816 & ~n14727;
  assign n14729 = ~n7924 & ~n14728;
  assign n14730 = ~controllable_hmaster2 & ~n14537;
  assign n14731 = ~n14401 & ~n14730;
  assign n14732 = ~controllable_hmaster1 & ~n14731;
  assign n14733 = ~n14400 & ~n14732;
  assign n14734 = ~i_hbusreq6 & ~n14733;
  assign n14735 = ~n13521 & ~n14734;
  assign n14736 = ~controllable_hgrant6 & ~n14735;
  assign n14737 = ~n14019 & ~n14736;
  assign n14738 = ~controllable_hmaster0 & ~n14737;
  assign n14739 = ~n14442 & ~n14738;
  assign n14740 = i_hlock8 & ~n14739;
  assign n14741 = ~controllable_hmaster2 & ~n14674;
  assign n14742 = ~n14401 & ~n14741;
  assign n14743 = ~controllable_hmaster1 & ~n14742;
  assign n14744 = ~n14400 & ~n14743;
  assign n14745 = ~i_hbusreq6 & ~n14744;
  assign n14746 = ~n13574 & ~n14745;
  assign n14747 = ~controllable_hgrant6 & ~n14746;
  assign n14748 = ~n14054 & ~n14747;
  assign n14749 = ~controllable_hmaster0 & ~n14748;
  assign n14750 = ~n14442 & ~n14749;
  assign n14751 = ~i_hlock8 & ~n14750;
  assign n14752 = ~n14740 & ~n14751;
  assign n14753 = ~i_hbusreq8 & ~n14752;
  assign n14754 = ~n13964 & ~n14753;
  assign n14755 = controllable_hmaster3 & ~n14754;
  assign n14756 = controllable_hgrant6 & ~n9522;
  assign n14757 = controllable_hmaster2 & ~n14472;
  assign n14758 = ~n14561 & ~n14757;
  assign n14759 = controllable_hmaster1 & ~n14758;
  assign n14760 = ~n14605 & ~n14759;
  assign n14761 = ~i_hbusreq6 & ~n14760;
  assign n14762 = ~n14095 & ~n14761;
  assign n14763 = ~controllable_hgrant6 & ~n14762;
  assign n14764 = ~n14756 & ~n14763;
  assign n14765 = controllable_hmaster0 & ~n14764;
  assign n14766 = ~n14685 & ~n14765;
  assign n14767 = ~i_hbusreq8 & ~n14766;
  assign n14768 = ~n14093 & ~n14767;
  assign n14769 = ~controllable_hmaster3 & ~n14768;
  assign n14770 = ~n14755 & ~n14769;
  assign n14771 = i_hlock7 & ~n14770;
  assign n14772 = controllable_hgrant6 & ~n9534;
  assign n14773 = controllable_hmaster2 & ~n14503;
  assign n14774 = ~n14561 & ~n14773;
  assign n14775 = controllable_hmaster1 & ~n14774;
  assign n14776 = ~n14605 & ~n14775;
  assign n14777 = ~i_hbusreq6 & ~n14776;
  assign n14778 = ~n14299 & ~n14777;
  assign n14779 = ~controllable_hgrant6 & ~n14778;
  assign n14780 = ~n14772 & ~n14779;
  assign n14781 = controllable_hmaster0 & ~n14780;
  assign n14782 = ~n14685 & ~n14781;
  assign n14783 = ~i_hbusreq8 & ~n14782;
  assign n14784 = ~n14297 & ~n14783;
  assign n14785 = ~controllable_hmaster3 & ~n14784;
  assign n14786 = ~n14755 & ~n14785;
  assign n14787 = ~i_hlock7 & ~n14786;
  assign n14788 = ~n14771 & ~n14787;
  assign n14789 = ~i_hbusreq7 & ~n14788;
  assign n14790 = ~n13963 & ~n14789;
  assign n14791 = n7924 & ~n14790;
  assign n14792 = ~n14729 & ~n14791;
  assign n14793 = ~n8214 & ~n14792;
  assign n14794 = ~n9561 & ~n14721;
  assign n14795 = i_hlock7 & ~n14794;
  assign n14796 = ~n9567 & ~n14721;
  assign n14797 = ~i_hlock7 & ~n14796;
  assign n14798 = ~n14795 & ~n14797;
  assign n14799 = ~i_hbusreq7 & ~n14798;
  assign n14800 = ~n13816 & ~n14799;
  assign n14801 = ~n7924 & ~n14800;
  assign n14802 = controllable_hgrant6 & ~n9556;
  assign n14803 = ~n14631 & ~n14757;
  assign n14804 = controllable_hmaster1 & ~n14803;
  assign n14805 = ~n14668 & ~n14804;
  assign n14806 = i_hlock6 & ~n14805;
  assign n14807 = ~n14631 & ~n14773;
  assign n14808 = controllable_hmaster1 & ~n14807;
  assign n14809 = ~n14668 & ~n14808;
  assign n14810 = ~i_hlock6 & ~n14809;
  assign n14811 = ~n14806 & ~n14810;
  assign n14812 = ~i_hbusreq6 & ~n14811;
  assign n14813 = ~n14174 & ~n14812;
  assign n14814 = ~controllable_hgrant6 & ~n14813;
  assign n14815 = ~n14802 & ~n14814;
  assign n14816 = ~controllable_hmaster0 & ~n14815;
  assign n14817 = ~n14611 & ~n14816;
  assign n14818 = ~i_hbusreq8 & ~n14817;
  assign n14819 = ~n14093 & ~n14818;
  assign n14820 = ~controllable_hmaster3 & ~n14819;
  assign n14821 = ~n14755 & ~n14820;
  assign n14822 = i_hlock7 & ~n14821;
  assign n14823 = ~n14699 & ~n14816;
  assign n14824 = ~i_hbusreq8 & ~n14823;
  assign n14825 = ~n14297 & ~n14824;
  assign n14826 = ~controllable_hmaster3 & ~n14825;
  assign n14827 = ~n14755 & ~n14826;
  assign n14828 = ~i_hlock7 & ~n14827;
  assign n14829 = ~n14822 & ~n14828;
  assign n14830 = ~i_hbusreq7 & ~n14829;
  assign n14831 = ~n13963 & ~n14830;
  assign n14832 = n7924 & ~n14831;
  assign n14833 = ~n14801 & ~n14832;
  assign n14834 = n8214 & ~n14833;
  assign n14835 = ~n14793 & ~n14834;
  assign n14836 = n8202 & ~n14835;
  assign n14837 = ~n14713 & ~n14836;
  assign n14838 = n7920 & ~n14837;
  assign n14839 = ~n8877 & ~n14838;
  assign n14840 = ~n7728 & ~n14839;
  assign n14841 = ~n13804 & ~n14840;
  assign n14842 = n7723 & ~n14841;
  assign n14843 = ~n7723 & ~n14839;
  assign n14844 = ~n14842 & ~n14843;
  assign n14845 = n7714 & ~n14844;
  assign n14846 = n7723 & ~n14839;
  assign n14847 = ~n8640 & ~n14838;
  assign n14848 = n7728 & ~n14847;
  assign n14849 = controllable_hgrant6 & ~n9605;
  assign n14850 = ~n9600 & ~n12764;
  assign n14851 = ~controllable_hmaster1 & ~n14850;
  assign n14852 = ~n9599 & ~n14851;
  assign n14853 = ~i_hbusreq6 & ~n14852;
  assign n14854 = ~n13135 & ~n14853;
  assign n14855 = ~controllable_hgrant6 & ~n14854;
  assign n14856 = ~n14849 & ~n14855;
  assign n14857 = controllable_hmaster0 & ~n14856;
  assign n14858 = ~n9612 & ~n14857;
  assign n14859 = i_hlock8 & ~n14858;
  assign n14860 = ~n9620 & ~n14857;
  assign n14861 = ~i_hlock8 & ~n14860;
  assign n14862 = ~n14859 & ~n14861;
  assign n14863 = ~i_hbusreq8 & ~n14862;
  assign n14864 = ~n13817 & ~n14863;
  assign n14865 = controllable_hmaster3 & ~n14864;
  assign n14866 = ~n9720 & ~n14865;
  assign n14867 = i_hlock7 & ~n14866;
  assign n14868 = ~n9732 & ~n14865;
  assign n14869 = ~i_hlock7 & ~n14868;
  assign n14870 = ~n14867 & ~n14869;
  assign n14871 = ~i_hbusreq7 & ~n14870;
  assign n14872 = ~n13816 & ~n14871;
  assign n14873 = ~n7924 & ~n14872;
  assign n14874 = controllable_hgrant5 & ~n9598;
  assign n14875 = controllable_hgrant4 & ~n9596;
  assign n14876 = controllable_hgrant3 & ~n9592;
  assign n14877 = controllable_hgrant1 & ~n9590;
  assign n14878 = ~n7928 & ~n9588;
  assign n14879 = i_hlock0 & ~n7735;
  assign n14880 = ~n13970 & ~n14879;
  assign n14881 = ~i_hbusreq0 & ~n14880;
  assign n14882 = ~n13052 & ~n14881;
  assign n14883 = ~i_hbusreq2 & ~n14882;
  assign n14884 = ~n13051 & ~n14883;
  assign n14885 = ~controllable_hgrant2 & ~n14884;
  assign n14886 = ~n7814 & ~n14885;
  assign n14887 = ~n7733 & ~n14886;
  assign n14888 = ~n12898 & ~n13970;
  assign n14889 = ~i_hbusreq0 & ~n14888;
  assign n14890 = ~n13052 & ~n14889;
  assign n14891 = ~i_hbusreq2 & ~n14890;
  assign n14892 = ~n13051 & ~n14891;
  assign n14893 = ~controllable_hgrant2 & ~n14892;
  assign n14894 = ~n12706 & ~n14893;
  assign n14895 = n7733 & ~n14894;
  assign n14896 = ~n14887 & ~n14895;
  assign n14897 = n7928 & ~n14896;
  assign n14898 = ~n14878 & ~n14897;
  assign n14899 = ~i_hbusreq1 & ~n14898;
  assign n14900 = ~n13214 & ~n14899;
  assign n14901 = ~controllable_hgrant1 & ~n14900;
  assign n14902 = ~n14877 & ~n14901;
  assign n14903 = ~i_hbusreq3 & ~n14902;
  assign n14904 = ~n13212 & ~n14903;
  assign n14905 = ~controllable_hgrant3 & ~n14904;
  assign n14906 = ~n14876 & ~n14905;
  assign n14907 = ~i_hbusreq9 & ~n14906;
  assign n14908 = ~n13210 & ~n14907;
  assign n14909 = ~i_hbusreq4 & ~n14908;
  assign n14910 = ~n13209 & ~n14909;
  assign n14911 = ~controllable_hgrant4 & ~n14910;
  assign n14912 = ~n14875 & ~n14911;
  assign n14913 = ~i_hbusreq5 & ~n14912;
  assign n14914 = ~n13207 & ~n14913;
  assign n14915 = ~controllable_hgrant5 & ~n14914;
  assign n14916 = ~n14874 & ~n14915;
  assign n14917 = controllable_hmaster1 & ~n14916;
  assign n14918 = controllable_hmaster2 & ~n14916;
  assign n14919 = ~n12942 & ~n14918;
  assign n14920 = ~controllable_hmaster1 & ~n14919;
  assign n14921 = ~n14917 & ~n14920;
  assign n14922 = ~i_hbusreq6 & ~n14921;
  assign n14923 = ~n13205 & ~n14922;
  assign n14924 = ~controllable_hgrant6 & ~n14923;
  assign n14925 = ~n14849 & ~n14924;
  assign n14926 = controllable_hmaster0 & ~n14925;
  assign n14927 = controllable_hgrant6 & ~n9611;
  assign n14928 = ~n13978 & ~n14895;
  assign n14929 = n7928 & ~n14928;
  assign n14930 = ~n8265 & ~n14929;
  assign n14931 = ~i_hbusreq1 & ~n14930;
  assign n14932 = ~n13528 & ~n14931;
  assign n14933 = ~controllable_hgrant1 & ~n14932;
  assign n14934 = ~n12681 & ~n14933;
  assign n14935 = ~i_hbusreq3 & ~n14934;
  assign n14936 = ~n13527 & ~n14935;
  assign n14937 = ~controllable_hgrant3 & ~n14936;
  assign n14938 = ~n12679 & ~n14937;
  assign n14939 = ~i_hbusreq9 & ~n14938;
  assign n14940 = ~n13526 & ~n14939;
  assign n14941 = ~i_hbusreq4 & ~n14940;
  assign n14942 = ~n13525 & ~n14941;
  assign n14943 = ~controllable_hgrant4 & ~n14942;
  assign n14944 = ~n13524 & ~n14943;
  assign n14945 = ~i_hbusreq5 & ~n14944;
  assign n14946 = ~n13523 & ~n14945;
  assign n14947 = ~controllable_hgrant5 & ~n14946;
  assign n14948 = ~n13522 & ~n14947;
  assign n14949 = ~controllable_hmaster2 & ~n14948;
  assign n14950 = ~n14918 & ~n14949;
  assign n14951 = ~controllable_hmaster1 & ~n14950;
  assign n14952 = ~n14917 & ~n14951;
  assign n14953 = ~i_hbusreq6 & ~n14952;
  assign n14954 = ~n13521 & ~n14953;
  assign n14955 = ~controllable_hgrant6 & ~n14954;
  assign n14956 = ~n14927 & ~n14955;
  assign n14957 = ~controllable_hmaster0 & ~n14956;
  assign n14958 = ~n14926 & ~n14957;
  assign n14959 = i_hlock8 & ~n14958;
  assign n14960 = controllable_hgrant6 & ~n9619;
  assign n14961 = ~n8297 & ~n14929;
  assign n14962 = ~i_hbusreq1 & ~n14961;
  assign n14963 = ~n13581 & ~n14962;
  assign n14964 = ~controllable_hgrant1 & ~n14963;
  assign n14965 = ~n12730 & ~n14964;
  assign n14966 = ~i_hbusreq3 & ~n14965;
  assign n14967 = ~n13580 & ~n14966;
  assign n14968 = ~controllable_hgrant3 & ~n14967;
  assign n14969 = ~n12728 & ~n14968;
  assign n14970 = ~i_hbusreq9 & ~n14969;
  assign n14971 = ~n13579 & ~n14970;
  assign n14972 = ~i_hbusreq4 & ~n14971;
  assign n14973 = ~n13578 & ~n14972;
  assign n14974 = ~controllable_hgrant4 & ~n14973;
  assign n14975 = ~n13577 & ~n14974;
  assign n14976 = ~i_hbusreq5 & ~n14975;
  assign n14977 = ~n13576 & ~n14976;
  assign n14978 = ~controllable_hgrant5 & ~n14977;
  assign n14979 = ~n13575 & ~n14978;
  assign n14980 = ~controllable_hmaster2 & ~n14979;
  assign n14981 = ~n14918 & ~n14980;
  assign n14982 = ~controllable_hmaster1 & ~n14981;
  assign n14983 = ~n14917 & ~n14982;
  assign n14984 = ~i_hbusreq6 & ~n14983;
  assign n14985 = ~n13574 & ~n14984;
  assign n14986 = ~controllable_hgrant6 & ~n14985;
  assign n14987 = ~n14960 & ~n14986;
  assign n14988 = ~controllable_hmaster0 & ~n14987;
  assign n14989 = ~n14926 & ~n14988;
  assign n14990 = ~i_hlock8 & ~n14989;
  assign n14991 = ~n14959 & ~n14990;
  assign n14992 = ~i_hbusreq8 & ~n14991;
  assign n14993 = ~n13964 & ~n14992;
  assign n14994 = controllable_hmaster3 & ~n14993;
  assign n14995 = controllable_hgrant6 & ~n9665;
  assign n14996 = controllable_hmaster2 & ~n14948;
  assign n14997 = controllable_hgrant5 & ~n9637;
  assign n14998 = controllable_hgrant4 & ~n9635;
  assign n14999 = controllable_hgrant3 & ~n9631;
  assign n15000 = i_hlock3 & ~n14934;
  assign n15001 = ~i_hlock3 & ~n14965;
  assign n15002 = ~n15000 & ~n15001;
  assign n15003 = ~i_hbusreq3 & ~n15002;
  assign n15004 = ~n14103 & ~n15003;
  assign n15005 = ~controllable_hgrant3 & ~n15004;
  assign n15006 = ~n14999 & ~n15005;
  assign n15007 = ~i_hbusreq9 & ~n15006;
  assign n15008 = ~n14101 & ~n15007;
  assign n15009 = ~i_hbusreq4 & ~n15008;
  assign n15010 = ~n14100 & ~n15009;
  assign n15011 = ~controllable_hgrant4 & ~n15010;
  assign n15012 = ~n14998 & ~n15011;
  assign n15013 = ~i_hbusreq5 & ~n15012;
  assign n15014 = ~n14098 & ~n15013;
  assign n15015 = ~controllable_hgrant5 & ~n15014;
  assign n15016 = ~n14997 & ~n15015;
  assign n15017 = ~controllable_hmaster2 & ~n15016;
  assign n15018 = ~n14996 & ~n15017;
  assign n15019 = controllable_hmaster1 & ~n15018;
  assign n15020 = controllable_hgrant5 & ~n9645;
  assign n15021 = i_hlock5 & ~n14944;
  assign n15022 = ~i_hlock5 & ~n14975;
  assign n15023 = ~n15021 & ~n15022;
  assign n15024 = ~i_hbusreq5 & ~n15023;
  assign n15025 = ~n14125 & ~n15024;
  assign n15026 = ~controllable_hgrant5 & ~n15025;
  assign n15027 = ~n15020 & ~n15026;
  assign n15028 = controllable_hmaster2 & ~n15027;
  assign n15029 = controllable_hgrant5 & ~n9659;
  assign n15030 = controllable_hgrant4 & ~n9657;
  assign n15031 = controllable_hgrant3 & ~n9653;
  assign n15032 = controllable_hgrant1 & ~n9651;
  assign n15033 = i_hlock1 & ~n14930;
  assign n15034 = ~i_hlock1 & ~n14961;
  assign n15035 = ~n15033 & ~n15034;
  assign n15036 = ~i_hbusreq1 & ~n15035;
  assign n15037 = ~n14142 & ~n15036;
  assign n15038 = ~controllable_hgrant1 & ~n15037;
  assign n15039 = ~n15032 & ~n15038;
  assign n15040 = ~i_hbusreq3 & ~n15039;
  assign n15041 = ~n14140 & ~n15040;
  assign n15042 = ~controllable_hgrant3 & ~n15041;
  assign n15043 = ~n15031 & ~n15042;
  assign n15044 = ~i_hbusreq9 & ~n15043;
  assign n15045 = ~n14138 & ~n15044;
  assign n15046 = ~i_hbusreq4 & ~n15045;
  assign n15047 = ~n14137 & ~n15046;
  assign n15048 = ~controllable_hgrant4 & ~n15047;
  assign n15049 = ~n15030 & ~n15048;
  assign n15050 = ~i_hbusreq5 & ~n15049;
  assign n15051 = ~n14135 & ~n15050;
  assign n15052 = ~controllable_hgrant5 & ~n15051;
  assign n15053 = ~n15029 & ~n15052;
  assign n15054 = ~controllable_hmaster2 & ~n15053;
  assign n15055 = ~n15028 & ~n15054;
  assign n15056 = ~controllable_hmaster1 & ~n15055;
  assign n15057 = ~n15019 & ~n15056;
  assign n15058 = ~i_hbusreq6 & ~n15057;
  assign n15059 = ~n14095 & ~n15058;
  assign n15060 = ~controllable_hgrant6 & ~n15059;
  assign n15061 = ~n14995 & ~n15060;
  assign n15062 = controllable_hmaster0 & ~n15061;
  assign n15063 = controllable_hgrant6 & ~n9715;
  assign n15064 = controllable_hgrant5 & ~n9677;
  assign n15065 = controllable_hgrant4 & ~n9675;
  assign n15066 = controllable_hgrant3 & ~n9671;
  assign n15067 = controllable_hgrant1 & ~n9669;
  assign n15068 = ~n9379 & ~n14929;
  assign n15069 = ~i_hbusreq1 & ~n15068;
  assign n15070 = ~n14183 & ~n15069;
  assign n15071 = ~controllable_hgrant1 & ~n15070;
  assign n15072 = ~n15067 & ~n15071;
  assign n15073 = ~i_hbusreq3 & ~n15072;
  assign n15074 = ~n14181 & ~n15073;
  assign n15075 = ~controllable_hgrant3 & ~n15074;
  assign n15076 = ~n15066 & ~n15075;
  assign n15077 = ~i_hbusreq9 & ~n15076;
  assign n15078 = ~n14179 & ~n15077;
  assign n15079 = ~i_hbusreq4 & ~n15078;
  assign n15080 = ~n14178 & ~n15079;
  assign n15081 = ~controllable_hgrant4 & ~n15080;
  assign n15082 = ~n15065 & ~n15081;
  assign n15083 = ~i_hbusreq5 & ~n15082;
  assign n15084 = ~n14176 & ~n15083;
  assign n15085 = ~controllable_hgrant5 & ~n15084;
  assign n15086 = ~n15064 & ~n15085;
  assign n15087 = ~controllable_hmaster2 & ~n15086;
  assign n15088 = ~n14996 & ~n15087;
  assign n15089 = controllable_hmaster1 & ~n15088;
  assign n15090 = controllable_hgrant5 & ~n9687;
  assign n15091 = controllable_hgrant4 & ~n9685;
  assign n15092 = i_hlock4 & ~n14940;
  assign n15093 = ~i_hlock4 & ~n14971;
  assign n15094 = ~n15092 & ~n15093;
  assign n15095 = ~i_hbusreq4 & ~n15094;
  assign n15096 = ~n14209 & ~n15095;
  assign n15097 = ~controllable_hgrant4 & ~n15096;
  assign n15098 = ~n15091 & ~n15097;
  assign n15099 = ~i_hbusreq5 & ~n15098;
  assign n15100 = ~n14207 & ~n15099;
  assign n15101 = ~controllable_hgrant5 & ~n15100;
  assign n15102 = ~n15090 & ~n15101;
  assign n15103 = controllable_hmaster2 & ~n15102;
  assign n15104 = controllable_hgrant5 & ~n9703;
  assign n15105 = controllable_hgrant4 & ~n9701;
  assign n15106 = controllable_hgrant3 & ~n9697;
  assign n15107 = controllable_hgrant1 & ~n9695;
  assign n15108 = n7733 & ~n13011;
  assign n15109 = ~n14239 & ~n15108;
  assign n15110 = n7928 & ~n15109;
  assign n15111 = ~n8440 & ~n15110;
  assign n15112 = ~i_hbusreq1 & ~n15111;
  assign n15113 = ~n14230 & ~n15112;
  assign n15114 = ~controllable_hgrant1 & ~n15113;
  assign n15115 = ~n15107 & ~n15114;
  assign n15116 = ~i_hbusreq3 & ~n15115;
  assign n15117 = ~n14228 & ~n15116;
  assign n15118 = ~controllable_hgrant3 & ~n15117;
  assign n15119 = ~n15106 & ~n15118;
  assign n15120 = ~i_hbusreq9 & ~n15119;
  assign n15121 = ~n14226 & ~n15120;
  assign n15122 = ~i_hbusreq4 & ~n15121;
  assign n15123 = ~n14225 & ~n15122;
  assign n15124 = ~controllable_hgrant4 & ~n15123;
  assign n15125 = ~n15105 & ~n15124;
  assign n15126 = ~i_hbusreq5 & ~n15125;
  assign n15127 = ~n14223 & ~n15126;
  assign n15128 = ~controllable_hgrant5 & ~n15127;
  assign n15129 = ~n15104 & ~n15128;
  assign n15130 = ~controllable_hmaster2 & ~n15129;
  assign n15131 = ~n15103 & ~n15130;
  assign n15132 = ~controllable_hmaster1 & ~n15131;
  assign n15133 = ~n15089 & ~n15132;
  assign n15134 = i_hlock6 & ~n15133;
  assign n15135 = controllable_hmaster2 & ~n14979;
  assign n15136 = ~n15087 & ~n15135;
  assign n15137 = controllable_hmaster1 & ~n15136;
  assign n15138 = ~n15132 & ~n15137;
  assign n15139 = ~i_hlock6 & ~n15138;
  assign n15140 = ~n15134 & ~n15139;
  assign n15141 = ~i_hbusreq6 & ~n15140;
  assign n15142 = ~n14174 & ~n15141;
  assign n15143 = ~controllable_hgrant6 & ~n15142;
  assign n15144 = ~n15063 & ~n15143;
  assign n15145 = ~controllable_hmaster0 & ~n15144;
  assign n15146 = ~n15062 & ~n15145;
  assign n15147 = ~i_hbusreq8 & ~n15146;
  assign n15148 = ~n14093 & ~n15147;
  assign n15149 = ~controllable_hmaster3 & ~n15148;
  assign n15150 = ~n14994 & ~n15149;
  assign n15151 = i_hlock7 & ~n15150;
  assign n15152 = controllable_hgrant6 & ~n9727;
  assign n15153 = ~n15017 & ~n15135;
  assign n15154 = controllable_hmaster1 & ~n15153;
  assign n15155 = ~n15056 & ~n15154;
  assign n15156 = ~i_hbusreq6 & ~n15155;
  assign n15157 = ~n14299 & ~n15156;
  assign n15158 = ~controllable_hgrant6 & ~n15157;
  assign n15159 = ~n15152 & ~n15158;
  assign n15160 = controllable_hmaster0 & ~n15159;
  assign n15161 = ~n15145 & ~n15160;
  assign n15162 = ~i_hbusreq8 & ~n15161;
  assign n15163 = ~n14297 & ~n15162;
  assign n15164 = ~controllable_hmaster3 & ~n15163;
  assign n15165 = ~n14994 & ~n15164;
  assign n15166 = ~i_hlock7 & ~n15165;
  assign n15167 = ~n15151 & ~n15166;
  assign n15168 = ~i_hbusreq7 & ~n15167;
  assign n15169 = ~n13963 & ~n15168;
  assign n15170 = n7924 & ~n15169;
  assign n15171 = ~n14873 & ~n15170;
  assign n15172 = n7920 & ~n15171;
  assign n15173 = ~n8640 & ~n15172;
  assign n15174 = ~n7728 & ~n15173;
  assign n15175 = ~n14848 & ~n15174;
  assign n15176 = ~n7723 & ~n15175;
  assign n15177 = ~n14846 & ~n15176;
  assign n15178 = ~n7714 & ~n15177;
  assign n15179 = ~n14845 & ~n15178;
  assign n15180 = ~n7705 & ~n15179;
  assign n15181 = ~n13121 & ~n15180;
  assign n15182 = n7808 & ~n15181;
  assign n15183 = ~n8650 & ~n15182;
  assign n15184 = n8195 & ~n15183;
  assign n15185 = ~n8196 & ~n15184;
  assign n15186 = ~n8193 & ~n15185;
  assign n15187 = ~n10059 & ~n13651;
  assign n15188 = i_hbusreq7 & ~n15187;
  assign n15189 = ~n10074 & ~n13662;
  assign n15190 = ~i_hbusreq7 & ~n15189;
  assign n15191 = ~n15188 & ~n15190;
  assign n15192 = ~n7924 & ~n15191;
  assign n15193 = controllable_hgrant6 & ~n10056;
  assign n15194 = controllable_hmaster1 & ~n13188;
  assign n15195 = ~n13189 & ~n13871;
  assign n15196 = ~controllable_hmaster1 & ~n15195;
  assign n15197 = ~n15194 & ~n15196;
  assign n15198 = ~controllable_hgrant6 & ~n15197;
  assign n15199 = ~n15193 & ~n15198;
  assign n15200 = controllable_hmaster0 & ~n15199;
  assign n15201 = ~n13682 & ~n15200;
  assign n15202 = ~controllable_hmaster3 & ~n15201;
  assign n15203 = ~n13672 & ~n15202;
  assign n15204 = i_hbusreq7 & ~n15203;
  assign n15205 = i_hbusreq8 & ~n15201;
  assign n15206 = controllable_hgrant6 & ~n10069;
  assign n15207 = i_hbusreq6 & ~n15197;
  assign n15208 = controllable_hmaster1 & ~n13634;
  assign n15209 = i_hlock5 & ~n13557;
  assign n15210 = ~i_hlock5 & ~n13596;
  assign n15211 = ~n15209 & ~n15210;
  assign n15212 = ~i_hbusreq5 & ~n15211;
  assign n15213 = ~n14125 & ~n15212;
  assign n15214 = ~controllable_hgrant5 & ~n15213;
  assign n15215 = ~n15020 & ~n15214;
  assign n15216 = controllable_hmaster2 & ~n15215;
  assign n15217 = ~n13702 & ~n15216;
  assign n15218 = ~controllable_hmaster1 & ~n15217;
  assign n15219 = ~n15208 & ~n15218;
  assign n15220 = ~i_hbusreq6 & ~n15219;
  assign n15221 = ~n15207 & ~n15220;
  assign n15222 = ~controllable_hgrant6 & ~n15221;
  assign n15223 = ~n15206 & ~n15222;
  assign n15224 = controllable_hmaster0 & ~n15223;
  assign n15225 = ~n13728 & ~n15224;
  assign n15226 = ~i_hbusreq8 & ~n15225;
  assign n15227 = ~n15205 & ~n15226;
  assign n15228 = ~controllable_hmaster3 & ~n15227;
  assign n15229 = ~n13714 & ~n15228;
  assign n15230 = ~i_hbusreq7 & ~n15229;
  assign n15231 = ~n15204 & ~n15230;
  assign n15232 = n7924 & ~n15231;
  assign n15233 = ~n15192 & ~n15232;
  assign n15234 = ~n8214 & ~n15233;
  assign n15235 = ~n10084 & ~n13651;
  assign n15236 = i_hbusreq7 & ~n15235;
  assign n15237 = ~n10098 & ~n13662;
  assign n15238 = ~i_hbusreq7 & ~n15237;
  assign n15239 = ~n15236 & ~n15238;
  assign n15240 = ~n7924 & ~n15239;
  assign n15241 = controllable_hgrant6 & ~n10081;
  assign n15242 = ~n13189 & ~n13920;
  assign n15243 = ~controllable_hmaster1 & ~n15242;
  assign n15244 = ~n15194 & ~n15243;
  assign n15245 = ~controllable_hgrant6 & ~n15244;
  assign n15246 = ~n15241 & ~n15245;
  assign n15247 = ~controllable_hmaster0 & ~n15246;
  assign n15248 = ~n13765 & ~n15247;
  assign n15249 = ~controllable_hmaster3 & ~n15248;
  assign n15250 = ~n13672 & ~n15249;
  assign n15251 = i_hbusreq7 & ~n15250;
  assign n15252 = i_hbusreq8 & ~n15248;
  assign n15253 = controllable_hgrant6 & ~n10093;
  assign n15254 = i_hbusreq6 & ~n15244;
  assign n15255 = i_hlock4 & ~n13553;
  assign n15256 = ~i_hlock4 & ~n13592;
  assign n15257 = ~n15255 & ~n15256;
  assign n15258 = ~i_hbusreq4 & ~n15257;
  assign n15259 = ~n14209 & ~n15258;
  assign n15260 = ~controllable_hgrant4 & ~n15259;
  assign n15261 = ~n15091 & ~n15260;
  assign n15262 = ~i_hbusreq5 & ~n15261;
  assign n15263 = ~n14207 & ~n15262;
  assign n15264 = ~controllable_hgrant5 & ~n15263;
  assign n15265 = ~n15090 & ~n15264;
  assign n15266 = controllable_hmaster2 & ~n15265;
  assign n15267 = ~n13702 & ~n15266;
  assign n15268 = ~controllable_hmaster1 & ~n15267;
  assign n15269 = ~n15208 & ~n15268;
  assign n15270 = ~i_hbusreq6 & ~n15269;
  assign n15271 = ~n15254 & ~n15270;
  assign n15272 = ~controllable_hgrant6 & ~n15271;
  assign n15273 = ~n15253 & ~n15272;
  assign n15274 = ~controllable_hmaster0 & ~n15273;
  assign n15275 = ~n13778 & ~n15274;
  assign n15276 = ~i_hbusreq8 & ~n15275;
  assign n15277 = ~n15252 & ~n15276;
  assign n15278 = ~controllable_hmaster3 & ~n15277;
  assign n15279 = ~n13714 & ~n15278;
  assign n15280 = ~i_hbusreq7 & ~n15279;
  assign n15281 = ~n15251 & ~n15280;
  assign n15282 = n7924 & ~n15281;
  assign n15283 = ~n15240 & ~n15282;
  assign n15284 = n8214 & ~n15283;
  assign n15285 = ~n15234 & ~n15284;
  assign n15286 = ~n8202 & ~n15285;
  assign n15287 = ~n10111 & ~n13651;
  assign n15288 = i_hbusreq7 & ~n15287;
  assign n15289 = ~n10126 & ~n13662;
  assign n15290 = ~i_hbusreq7 & ~n15289;
  assign n15291 = ~n15288 & ~n15290;
  assign n15292 = ~n7924 & ~n15291;
  assign n15293 = controllable_hgrant6 & ~n10108;
  assign n15294 = controllable_hmaster2 & ~n13188;
  assign n15295 = ~n13862 & ~n15294;
  assign n15296 = controllable_hmaster1 & ~n15295;
  assign n15297 = ~n13677 & ~n15296;
  assign n15298 = ~controllable_hgrant6 & ~n15297;
  assign n15299 = ~n15293 & ~n15298;
  assign n15300 = controllable_hmaster0 & ~n15299;
  assign n15301 = ~n13682 & ~n15300;
  assign n15302 = ~controllable_hmaster3 & ~n15301;
  assign n15303 = ~n13672 & ~n15302;
  assign n15304 = i_hbusreq7 & ~n15303;
  assign n15305 = i_hbusreq8 & ~n15301;
  assign n15306 = controllable_hgrant6 & ~n10121;
  assign n15307 = i_hbusreq6 & ~n15297;
  assign n15308 = controllable_hmaster2 & ~n13634;
  assign n15309 = i_hlock3 & ~n13547;
  assign n15310 = ~i_hlock3 & ~n13586;
  assign n15311 = ~n15309 & ~n15310;
  assign n15312 = ~i_hbusreq3 & ~n15311;
  assign n15313 = ~n14103 & ~n15312;
  assign n15314 = ~controllable_hgrant3 & ~n15313;
  assign n15315 = ~n14999 & ~n15314;
  assign n15316 = ~i_hbusreq9 & ~n15315;
  assign n15317 = ~n14101 & ~n15316;
  assign n15318 = ~i_hbusreq4 & ~n15317;
  assign n15319 = ~n14100 & ~n15318;
  assign n15320 = ~controllable_hgrant4 & ~n15319;
  assign n15321 = ~n14998 & ~n15320;
  assign n15322 = ~i_hbusreq5 & ~n15321;
  assign n15323 = ~n14098 & ~n15322;
  assign n15324 = ~controllable_hgrant5 & ~n15323;
  assign n15325 = ~n14997 & ~n15324;
  assign n15326 = ~controllable_hmaster2 & ~n15325;
  assign n15327 = ~n15308 & ~n15326;
  assign n15328 = controllable_hmaster1 & ~n15327;
  assign n15329 = ~n13721 & ~n15328;
  assign n15330 = ~i_hbusreq6 & ~n15329;
  assign n15331 = ~n15307 & ~n15330;
  assign n15332 = ~controllable_hgrant6 & ~n15331;
  assign n15333 = ~n15306 & ~n15332;
  assign n15334 = controllable_hmaster0 & ~n15333;
  assign n15335 = ~n13728 & ~n15334;
  assign n15336 = ~i_hbusreq8 & ~n15335;
  assign n15337 = ~n15305 & ~n15336;
  assign n15338 = ~controllable_hmaster3 & ~n15337;
  assign n15339 = ~n13714 & ~n15338;
  assign n15340 = ~i_hbusreq7 & ~n15339;
  assign n15341 = ~n15304 & ~n15340;
  assign n15342 = n7924 & ~n15341;
  assign n15343 = ~n15292 & ~n15342;
  assign n15344 = ~n8214 & ~n15343;
  assign n15345 = ~n10136 & ~n13651;
  assign n15346 = i_hbusreq7 & ~n15345;
  assign n15347 = ~n10150 & ~n13662;
  assign n15348 = ~i_hbusreq7 & ~n15347;
  assign n15349 = ~n15346 & ~n15348;
  assign n15350 = ~n7924 & ~n15349;
  assign n15351 = controllable_hgrant6 & ~n10133;
  assign n15352 = ~n13908 & ~n15294;
  assign n15353 = controllable_hmaster1 & ~n15352;
  assign n15354 = ~n13677 & ~n15353;
  assign n15355 = ~controllable_hgrant6 & ~n15354;
  assign n15356 = ~n15351 & ~n15355;
  assign n15357 = ~controllable_hmaster0 & ~n15356;
  assign n15358 = ~n13765 & ~n15357;
  assign n15359 = ~controllable_hmaster3 & ~n15358;
  assign n15360 = ~n13672 & ~n15359;
  assign n15361 = i_hbusreq7 & ~n15360;
  assign n15362 = i_hbusreq8 & ~n15358;
  assign n15363 = controllable_hgrant6 & ~n10145;
  assign n15364 = i_hbusreq6 & ~n15354;
  assign n15365 = ~n9379 & ~n13542;
  assign n15366 = ~i_hbusreq1 & ~n15365;
  assign n15367 = ~n14183 & ~n15366;
  assign n15368 = ~controllable_hgrant1 & ~n15367;
  assign n15369 = ~n15067 & ~n15368;
  assign n15370 = ~i_hbusreq3 & ~n15369;
  assign n15371 = ~n14181 & ~n15370;
  assign n15372 = ~controllable_hgrant3 & ~n15371;
  assign n15373 = ~n15066 & ~n15372;
  assign n15374 = ~i_hbusreq9 & ~n15373;
  assign n15375 = ~n14179 & ~n15374;
  assign n15376 = ~i_hbusreq4 & ~n15375;
  assign n15377 = ~n14178 & ~n15376;
  assign n15378 = ~controllable_hgrant4 & ~n15377;
  assign n15379 = ~n15065 & ~n15378;
  assign n15380 = ~i_hbusreq5 & ~n15379;
  assign n15381 = ~n14176 & ~n15380;
  assign n15382 = ~controllable_hgrant5 & ~n15381;
  assign n15383 = ~n15064 & ~n15382;
  assign n15384 = ~controllable_hmaster2 & ~n15383;
  assign n15385 = ~n15308 & ~n15384;
  assign n15386 = controllable_hmaster1 & ~n15385;
  assign n15387 = ~n13721 & ~n15386;
  assign n15388 = ~i_hbusreq6 & ~n15387;
  assign n15389 = ~n15364 & ~n15388;
  assign n15390 = ~controllable_hgrant6 & ~n15389;
  assign n15391 = ~n15363 & ~n15390;
  assign n15392 = ~controllable_hmaster0 & ~n15391;
  assign n15393 = ~n13778 & ~n15392;
  assign n15394 = ~i_hbusreq8 & ~n15393;
  assign n15395 = ~n15362 & ~n15394;
  assign n15396 = ~controllable_hmaster3 & ~n15395;
  assign n15397 = ~n13714 & ~n15396;
  assign n15398 = ~i_hbusreq7 & ~n15397;
  assign n15399 = ~n15361 & ~n15398;
  assign n15400 = n7924 & ~n15399;
  assign n15401 = ~n15350 & ~n15400;
  assign n15402 = n8214 & ~n15401;
  assign n15403 = ~n15344 & ~n15402;
  assign n15404 = n8202 & ~n15403;
  assign n15405 = ~n15286 & ~n15404;
  assign n15406 = n7920 & ~n15405;
  assign n15407 = ~n10014 & ~n15406;
  assign n15408 = n7728 & ~n15407;
  assign n15409 = ~n10170 & ~n14721;
  assign n15410 = i_hlock7 & ~n15409;
  assign n15411 = ~n10180 & ~n14721;
  assign n15412 = ~i_hlock7 & ~n15411;
  assign n15413 = ~n15410 & ~n15412;
  assign n15414 = ~i_hbusreq7 & ~n15413;
  assign n15415 = ~n13816 & ~n15414;
  assign n15416 = ~n7924 & ~n15415;
  assign n15417 = controllable_hgrant6 & ~n10165;
  assign n15418 = i_hlock5 & ~n14468;
  assign n15419 = ~i_hlock5 & ~n14499;
  assign n15420 = ~n15418 & ~n15419;
  assign n15421 = ~i_hbusreq5 & ~n15420;
  assign n15422 = ~n14125 & ~n15421;
  assign n15423 = ~controllable_hgrant5 & ~n15422;
  assign n15424 = ~n15020 & ~n15423;
  assign n15425 = controllable_hmaster2 & ~n15424;
  assign n15426 = ~n14603 & ~n15425;
  assign n15427 = ~controllable_hmaster1 & ~n15426;
  assign n15428 = ~n14563 & ~n15427;
  assign n15429 = ~i_hbusreq6 & ~n15428;
  assign n15430 = ~n14095 & ~n15429;
  assign n15431 = ~controllable_hgrant6 & ~n15430;
  assign n15432 = ~n15417 & ~n15431;
  assign n15433 = controllable_hmaster0 & ~n15432;
  assign n15434 = ~n14685 & ~n15433;
  assign n15435 = ~i_hbusreq8 & ~n15434;
  assign n15436 = ~n14093 & ~n15435;
  assign n15437 = ~controllable_hmaster3 & ~n15436;
  assign n15438 = ~n14755 & ~n15437;
  assign n15439 = i_hlock7 & ~n15438;
  assign n15440 = controllable_hgrant6 & ~n10175;
  assign n15441 = ~n14693 & ~n15427;
  assign n15442 = ~i_hbusreq6 & ~n15441;
  assign n15443 = ~n14299 & ~n15442;
  assign n15444 = ~controllable_hgrant6 & ~n15443;
  assign n15445 = ~n15440 & ~n15444;
  assign n15446 = controllable_hmaster0 & ~n15445;
  assign n15447 = ~n14685 & ~n15446;
  assign n15448 = ~i_hbusreq8 & ~n15447;
  assign n15449 = ~n14297 & ~n15448;
  assign n15450 = ~controllable_hmaster3 & ~n15449;
  assign n15451 = ~n14755 & ~n15450;
  assign n15452 = ~i_hlock7 & ~n15451;
  assign n15453 = ~n15439 & ~n15452;
  assign n15454 = ~i_hbusreq7 & ~n15453;
  assign n15455 = ~n13963 & ~n15454;
  assign n15456 = n7924 & ~n15455;
  assign n15457 = ~n15416 & ~n15456;
  assign n15458 = ~n8214 & ~n15457;
  assign n15459 = ~n10200 & ~n14721;
  assign n15460 = i_hlock7 & ~n15459;
  assign n15461 = ~n10206 & ~n14721;
  assign n15462 = ~i_hlock7 & ~n15461;
  assign n15463 = ~n15460 & ~n15462;
  assign n15464 = ~i_hbusreq7 & ~n15463;
  assign n15465 = ~n13816 & ~n15464;
  assign n15466 = ~n7924 & ~n15465;
  assign n15467 = controllable_hgrant6 & ~n10195;
  assign n15468 = i_hlock4 & ~n14464;
  assign n15469 = ~i_hlock4 & ~n14495;
  assign n15470 = ~n15468 & ~n15469;
  assign n15471 = ~i_hbusreq4 & ~n15470;
  assign n15472 = ~n14209 & ~n15471;
  assign n15473 = ~controllable_hgrant4 & ~n15472;
  assign n15474 = ~n15091 & ~n15473;
  assign n15475 = ~i_hbusreq5 & ~n15474;
  assign n15476 = ~n14207 & ~n15475;
  assign n15477 = ~controllable_hgrant5 & ~n15476;
  assign n15478 = ~n15090 & ~n15477;
  assign n15479 = controllable_hmaster2 & ~n15478;
  assign n15480 = ~n14666 & ~n15479;
  assign n15481 = ~controllable_hmaster1 & ~n15480;
  assign n15482 = ~n14633 & ~n15481;
  assign n15483 = i_hlock6 & ~n15482;
  assign n15484 = ~n14677 & ~n15481;
  assign n15485 = ~i_hlock6 & ~n15484;
  assign n15486 = ~n15483 & ~n15485;
  assign n15487 = ~i_hbusreq6 & ~n15486;
  assign n15488 = ~n14174 & ~n15487;
  assign n15489 = ~controllable_hgrant6 & ~n15488;
  assign n15490 = ~n15467 & ~n15489;
  assign n15491 = ~controllable_hmaster0 & ~n15490;
  assign n15492 = ~n14611 & ~n15491;
  assign n15493 = ~i_hbusreq8 & ~n15492;
  assign n15494 = ~n14093 & ~n15493;
  assign n15495 = ~controllable_hmaster3 & ~n15494;
  assign n15496 = ~n14755 & ~n15495;
  assign n15497 = i_hlock7 & ~n15496;
  assign n15498 = ~n14699 & ~n15491;
  assign n15499 = ~i_hbusreq8 & ~n15498;
  assign n15500 = ~n14297 & ~n15499;
  assign n15501 = ~controllable_hmaster3 & ~n15500;
  assign n15502 = ~n14755 & ~n15501;
  assign n15503 = ~i_hlock7 & ~n15502;
  assign n15504 = ~n15497 & ~n15503;
  assign n15505 = ~i_hbusreq7 & ~n15504;
  assign n15506 = ~n13963 & ~n15505;
  assign n15507 = n7924 & ~n15506;
  assign n15508 = ~n15466 & ~n15507;
  assign n15509 = n8214 & ~n15508;
  assign n15510 = ~n15458 & ~n15509;
  assign n15511 = ~n8202 & ~n15510;
  assign n15512 = ~n10224 & ~n14721;
  assign n15513 = i_hlock7 & ~n15512;
  assign n15514 = ~n10236 & ~n14721;
  assign n15515 = ~i_hlock7 & ~n15514;
  assign n15516 = ~n15513 & ~n15515;
  assign n15517 = ~i_hbusreq7 & ~n15516;
  assign n15518 = ~n13816 & ~n15517;
  assign n15519 = ~n7924 & ~n15518;
  assign n15520 = controllable_hgrant6 & ~n10219;
  assign n15521 = i_hlock3 & ~n14458;
  assign n15522 = ~i_hlock3 & ~n14489;
  assign n15523 = ~n15521 & ~n15522;
  assign n15524 = ~i_hbusreq3 & ~n15523;
  assign n15525 = ~n14103 & ~n15524;
  assign n15526 = ~controllable_hgrant3 & ~n15525;
  assign n15527 = ~n14999 & ~n15526;
  assign n15528 = ~i_hbusreq9 & ~n15527;
  assign n15529 = ~n14101 & ~n15528;
  assign n15530 = ~i_hbusreq4 & ~n15529;
  assign n15531 = ~n14100 & ~n15530;
  assign n15532 = ~controllable_hgrant4 & ~n15531;
  assign n15533 = ~n14998 & ~n15532;
  assign n15534 = ~i_hbusreq5 & ~n15533;
  assign n15535 = ~n14098 & ~n15534;
  assign n15536 = ~controllable_hgrant5 & ~n15535;
  assign n15537 = ~n14997 & ~n15536;
  assign n15538 = ~controllable_hmaster2 & ~n15537;
  assign n15539 = ~n14538 & ~n15538;
  assign n15540 = controllable_hmaster1 & ~n15539;
  assign n15541 = ~n14605 & ~n15540;
  assign n15542 = ~i_hbusreq6 & ~n15541;
  assign n15543 = ~n14095 & ~n15542;
  assign n15544 = ~controllable_hgrant6 & ~n15543;
  assign n15545 = ~n15520 & ~n15544;
  assign n15546 = controllable_hmaster0 & ~n15545;
  assign n15547 = ~n14685 & ~n15546;
  assign n15548 = ~i_hbusreq8 & ~n15547;
  assign n15549 = ~n14093 & ~n15548;
  assign n15550 = ~controllable_hmaster3 & ~n15549;
  assign n15551 = ~n14755 & ~n15550;
  assign n15552 = i_hlock7 & ~n15551;
  assign n15553 = controllable_hgrant6 & ~n10231;
  assign n15554 = ~n14675 & ~n15538;
  assign n15555 = controllable_hmaster1 & ~n15554;
  assign n15556 = ~n14605 & ~n15555;
  assign n15557 = ~i_hbusreq6 & ~n15556;
  assign n15558 = ~n14299 & ~n15557;
  assign n15559 = ~controllable_hgrant6 & ~n15558;
  assign n15560 = ~n15553 & ~n15559;
  assign n15561 = controllable_hmaster0 & ~n15560;
  assign n15562 = ~n14685 & ~n15561;
  assign n15563 = ~i_hbusreq8 & ~n15562;
  assign n15564 = ~n14297 & ~n15563;
  assign n15565 = ~controllable_hmaster3 & ~n15564;
  assign n15566 = ~n14755 & ~n15565;
  assign n15567 = ~i_hlock7 & ~n15566;
  assign n15568 = ~n15552 & ~n15567;
  assign n15569 = ~i_hbusreq7 & ~n15568;
  assign n15570 = ~n13963 & ~n15569;
  assign n15571 = n7924 & ~n15570;
  assign n15572 = ~n15519 & ~n15571;
  assign n15573 = ~n8214 & ~n15572;
  assign n15574 = ~n10258 & ~n14721;
  assign n15575 = i_hlock7 & ~n15574;
  assign n15576 = ~n10264 & ~n14721;
  assign n15577 = ~i_hlock7 & ~n15576;
  assign n15578 = ~n15575 & ~n15577;
  assign n15579 = ~i_hbusreq7 & ~n15578;
  assign n15580 = ~n13816 & ~n15579;
  assign n15581 = ~n7924 & ~n15580;
  assign n15582 = controllable_hgrant6 & ~n10253;
  assign n15583 = ~n9379 & ~n14453;
  assign n15584 = ~i_hbusreq1 & ~n15583;
  assign n15585 = ~n14183 & ~n15584;
  assign n15586 = ~controllable_hgrant1 & ~n15585;
  assign n15587 = ~n15067 & ~n15586;
  assign n15588 = ~i_hbusreq3 & ~n15587;
  assign n15589 = ~n14181 & ~n15588;
  assign n15590 = ~controllable_hgrant3 & ~n15589;
  assign n15591 = ~n15066 & ~n15590;
  assign n15592 = ~i_hbusreq9 & ~n15591;
  assign n15593 = ~n14179 & ~n15592;
  assign n15594 = ~i_hbusreq4 & ~n15593;
  assign n15595 = ~n14178 & ~n15594;
  assign n15596 = ~controllable_hgrant4 & ~n15595;
  assign n15597 = ~n15065 & ~n15596;
  assign n15598 = ~i_hbusreq5 & ~n15597;
  assign n15599 = ~n14176 & ~n15598;
  assign n15600 = ~controllable_hgrant5 & ~n15599;
  assign n15601 = ~n15064 & ~n15600;
  assign n15602 = ~controllable_hmaster2 & ~n15601;
  assign n15603 = ~n14538 & ~n15602;
  assign n15604 = controllable_hmaster1 & ~n15603;
  assign n15605 = ~n14668 & ~n15604;
  assign n15606 = i_hlock6 & ~n15605;
  assign n15607 = ~n14675 & ~n15602;
  assign n15608 = controllable_hmaster1 & ~n15607;
  assign n15609 = ~n14668 & ~n15608;
  assign n15610 = ~i_hlock6 & ~n15609;
  assign n15611 = ~n15606 & ~n15610;
  assign n15612 = ~i_hbusreq6 & ~n15611;
  assign n15613 = ~n14174 & ~n15612;
  assign n15614 = ~controllable_hgrant6 & ~n15613;
  assign n15615 = ~n15582 & ~n15614;
  assign n15616 = ~controllable_hmaster0 & ~n15615;
  assign n15617 = ~n14611 & ~n15616;
  assign n15618 = ~i_hbusreq8 & ~n15617;
  assign n15619 = ~n14093 & ~n15618;
  assign n15620 = ~controllable_hmaster3 & ~n15619;
  assign n15621 = ~n14755 & ~n15620;
  assign n15622 = i_hlock7 & ~n15621;
  assign n15623 = ~n14699 & ~n15616;
  assign n15624 = ~i_hbusreq8 & ~n15623;
  assign n15625 = ~n14297 & ~n15624;
  assign n15626 = ~controllable_hmaster3 & ~n15625;
  assign n15627 = ~n14755 & ~n15626;
  assign n15628 = ~i_hlock7 & ~n15627;
  assign n15629 = ~n15622 & ~n15628;
  assign n15630 = ~i_hbusreq7 & ~n15629;
  assign n15631 = ~n13963 & ~n15630;
  assign n15632 = n7924 & ~n15631;
  assign n15633 = ~n15581 & ~n15632;
  assign n15634 = n8214 & ~n15633;
  assign n15635 = ~n15573 & ~n15634;
  assign n15636 = n8202 & ~n15635;
  assign n15637 = ~n15511 & ~n15636;
  assign n15638 = n7920 & ~n15637;
  assign n15639 = ~n10014 & ~n15638;
  assign n15640 = ~n7728 & ~n15639;
  assign n15641 = ~n15408 & ~n15640;
  assign n15642 = n7723 & ~n15641;
  assign n15643 = ~n7723 & ~n15639;
  assign n15644 = ~n15642 & ~n15643;
  assign n15645 = n7714 & ~n15644;
  assign n15646 = n7723 & ~n15639;
  assign n15647 = ~n8640 & ~n15638;
  assign n15648 = n7728 & ~n15647;
  assign n15649 = ~n15174 & ~n15648;
  assign n15650 = ~n7723 & ~n15649;
  assign n15651 = ~n15646 & ~n15650;
  assign n15652 = ~n7714 & ~n15651;
  assign n15653 = ~n15645 & ~n15652;
  assign n15654 = ~n7705 & ~n15653;
  assign n15655 = ~n10052 & ~n15654;
  assign n15656 = n7808 & ~n15655;
  assign n15657 = ~n9908 & ~n15656;
  assign n15658 = ~n8195 & ~n15657;
  assign n15659 = n7924 & ~n15170;
  assign n15660 = ~n8214 & ~n15659;
  assign n15661 = ~n10105 & ~n13322;
  assign n15662 = ~controllable_hmaster1 & ~n15661;
  assign n15663 = ~n10053 & ~n15662;
  assign n15664 = ~controllable_hgrant6 & ~n15663;
  assign n15665 = ~n13198 & ~n15664;
  assign n15666 = controllable_hmaster0 & ~n15665;
  assign n15667 = ~n9099 & ~n15666;
  assign n15668 = controllable_hmaster3 & ~n15667;
  assign n15669 = ~n8995 & ~n15668;
  assign n15670 = i_hbusreq7 & ~n15669;
  assign n15671 = i_hbusreq8 & ~n15667;
  assign n15672 = controllable_hgrant6 & ~n10756;
  assign n15673 = i_hbusreq6 & ~n15663;
  assign n15674 = controllable_hgrant5 & ~n10750;
  assign n15675 = controllable_hgrant4 & ~n10748;
  assign n15676 = controllable_hgrant3 & ~n10744;
  assign n15677 = controllable_hgrant1 & ~n10742;
  assign n15678 = n7928 & ~n12717;
  assign n15679 = ~i_hbusreq1 & ~n15678;
  assign n15680 = ~n13343 & ~n15679;
  assign n15681 = ~controllable_hgrant1 & ~n15680;
  assign n15682 = ~n15677 & ~n15681;
  assign n15683 = ~i_hbusreq3 & ~n15682;
  assign n15684 = ~n13342 & ~n15683;
  assign n15685 = ~controllable_hgrant3 & ~n15684;
  assign n15686 = ~n15676 & ~n15685;
  assign n15687 = ~i_hbusreq9 & ~n15686;
  assign n15688 = ~n13341 & ~n15687;
  assign n15689 = ~i_hbusreq4 & ~n15688;
  assign n15690 = ~n13340 & ~n15689;
  assign n15691 = ~controllable_hgrant4 & ~n15690;
  assign n15692 = ~n15675 & ~n15691;
  assign n15693 = ~i_hbusreq5 & ~n15692;
  assign n15694 = ~n13339 & ~n15693;
  assign n15695 = ~controllable_hgrant5 & ~n15694;
  assign n15696 = ~n15674 & ~n15695;
  assign n15697 = ~controllable_hmaster2 & ~n15696;
  assign n15698 = ~n10739 & ~n15697;
  assign n15699 = ~controllable_hmaster1 & ~n15698;
  assign n15700 = ~n10738 & ~n15699;
  assign n15701 = ~i_hbusreq6 & ~n15700;
  assign n15702 = ~n15673 & ~n15701;
  assign n15703 = ~controllable_hgrant6 & ~n15702;
  assign n15704 = ~n15672 & ~n15703;
  assign n15705 = controllable_hmaster0 & ~n15704;
  assign n15706 = ~controllable_hmaster0 & ~n10756;
  assign n15707 = ~n15705 & ~n15706;
  assign n15708 = ~i_hbusreq8 & ~n15707;
  assign n15709 = ~n15671 & ~n15708;
  assign n15710 = controllable_hmaster3 & ~n15709;
  assign n15711 = ~n10786 & ~n15710;
  assign n15712 = ~i_hbusreq7 & ~n15711;
  assign n15713 = ~n15670 & ~n15712;
  assign n15714 = ~n7924 & ~n15713;
  assign n15715 = ~n13399 & ~n15294;
  assign n15716 = ~controllable_hmaster1 & ~n15715;
  assign n15717 = ~n15194 & ~n15716;
  assign n15718 = ~controllable_hgrant6 & ~n15717;
  assign n15719 = ~n13198 & ~n15718;
  assign n15720 = controllable_hmaster0 & ~n15719;
  assign n15721 = ~n13682 & ~n15720;
  assign n15722 = controllable_hmaster3 & ~n15721;
  assign n15723 = ~n13201 & ~n15722;
  assign n15724 = i_hbusreq7 & ~n15723;
  assign n15725 = i_hbusreq8 & ~n15721;
  assign n15726 = i_hbusreq6 & ~n15717;
  assign n15727 = controllable_hgrant5 & ~n10737;
  assign n15728 = controllable_hgrant4 & ~n10735;
  assign n15729 = controllable_hgrant3 & ~n10731;
  assign n15730 = controllable_hgrant1 & ~n10729;
  assign n15731 = n7928 & ~n14897;
  assign n15732 = ~i_hbusreq1 & ~n15731;
  assign n15733 = ~n13264 & ~n15732;
  assign n15734 = ~controllable_hgrant1 & ~n15733;
  assign n15735 = ~n15730 & ~n15734;
  assign n15736 = ~i_hbusreq3 & ~n15735;
  assign n15737 = ~n13262 & ~n15736;
  assign n15738 = ~controllable_hgrant3 & ~n15737;
  assign n15739 = ~n15729 & ~n15738;
  assign n15740 = ~i_hbusreq9 & ~n15739;
  assign n15741 = ~n13260 & ~n15740;
  assign n15742 = ~i_hbusreq4 & ~n15741;
  assign n15743 = ~n13259 & ~n15742;
  assign n15744 = ~controllable_hgrant4 & ~n15743;
  assign n15745 = ~n15728 & ~n15744;
  assign n15746 = ~i_hbusreq5 & ~n15745;
  assign n15747 = ~n13257 & ~n15746;
  assign n15748 = ~controllable_hgrant5 & ~n15747;
  assign n15749 = ~n15727 & ~n15748;
  assign n15750 = controllable_hmaster1 & ~n15749;
  assign n15751 = controllable_hmaster2 & ~n15749;
  assign n15752 = n7928 & ~n12908;
  assign n15753 = ~i_hbusreq1 & ~n15752;
  assign n15754 = ~n13485 & ~n15753;
  assign n15755 = ~controllable_hgrant1 & ~n15754;
  assign n15756 = ~n15677 & ~n15755;
  assign n15757 = ~i_hbusreq3 & ~n15756;
  assign n15758 = ~n13484 & ~n15757;
  assign n15759 = ~controllable_hgrant3 & ~n15758;
  assign n15760 = ~n15676 & ~n15759;
  assign n15761 = ~i_hbusreq9 & ~n15760;
  assign n15762 = ~n13483 & ~n15761;
  assign n15763 = ~i_hbusreq4 & ~n15762;
  assign n15764 = ~n13482 & ~n15763;
  assign n15765 = ~controllable_hgrant4 & ~n15764;
  assign n15766 = ~n15675 & ~n15765;
  assign n15767 = ~i_hbusreq5 & ~n15766;
  assign n15768 = ~n13481 & ~n15767;
  assign n15769 = ~controllable_hgrant5 & ~n15768;
  assign n15770 = ~n15674 & ~n15769;
  assign n15771 = ~controllable_hmaster2 & ~n15770;
  assign n15772 = ~n15751 & ~n15771;
  assign n15773 = ~controllable_hmaster1 & ~n15772;
  assign n15774 = ~n15750 & ~n15773;
  assign n15775 = ~i_hbusreq6 & ~n15774;
  assign n15776 = ~n15726 & ~n15775;
  assign n15777 = ~controllable_hgrant6 & ~n15776;
  assign n15778 = ~n15672 & ~n15777;
  assign n15779 = controllable_hmaster0 & ~n15778;
  assign n15780 = n7928 & ~n14929;
  assign n15781 = ~i_hbusreq1 & ~n15780;
  assign n15782 = ~n13264 & ~n15781;
  assign n15783 = ~controllable_hgrant1 & ~n15782;
  assign n15784 = ~n15677 & ~n15783;
  assign n15785 = ~i_hbusreq3 & ~n15784;
  assign n15786 = ~n13262 & ~n15785;
  assign n15787 = ~controllable_hgrant3 & ~n15786;
  assign n15788 = ~n15676 & ~n15787;
  assign n15789 = ~i_hbusreq9 & ~n15788;
  assign n15790 = ~n13260 & ~n15789;
  assign n15791 = ~i_hbusreq4 & ~n15790;
  assign n15792 = ~n13259 & ~n15791;
  assign n15793 = ~controllable_hgrant4 & ~n15792;
  assign n15794 = ~n15675 & ~n15793;
  assign n15795 = ~i_hbusreq5 & ~n15794;
  assign n15796 = ~n13257 & ~n15795;
  assign n15797 = ~controllable_hgrant5 & ~n15796;
  assign n15798 = ~n15674 & ~n15797;
  assign n15799 = ~controllable_hmaster2 & ~n15798;
  assign n15800 = ~n15751 & ~n15799;
  assign n15801 = ~controllable_hmaster1 & ~n15800;
  assign n15802 = ~n15750 & ~n15801;
  assign n15803 = ~i_hbusreq6 & ~n15802;
  assign n15804 = ~n13299 & ~n15803;
  assign n15805 = ~controllable_hgrant6 & ~n15804;
  assign n15806 = ~n15672 & ~n15805;
  assign n15807 = ~controllable_hmaster0 & ~n15806;
  assign n15808 = ~n15779 & ~n15807;
  assign n15809 = ~i_hbusreq8 & ~n15808;
  assign n15810 = ~n15725 & ~n15809;
  assign n15811 = controllable_hmaster3 & ~n15810;
  assign n15812 = controllable_hgrant6 & ~n10761;
  assign n15813 = ~i_hbusreq6 & ~n15798;
  assign n15814 = ~n13299 & ~n15813;
  assign n15815 = ~controllable_hgrant6 & ~n15814;
  assign n15816 = ~n15812 & ~n15815;
  assign n15817 = controllable_hmaster0 & ~n15816;
  assign n15818 = controllable_hgrant6 & ~n10781;
  assign n15819 = controllable_hmaster1 & ~n15798;
  assign n15820 = controllable_hmaster2 & ~n15798;
  assign n15821 = controllable_hgrant5 & ~n10775;
  assign n15822 = controllable_hgrant4 & ~n10773;
  assign n15823 = controllable_hgrant3 & ~n10769;
  assign n15824 = controllable_hgrant1 & ~n10767;
  assign n15825 = n7928 & ~n15110;
  assign n15826 = ~i_hbusreq1 & ~n15825;
  assign n15827 = ~n13264 & ~n15826;
  assign n15828 = ~controllable_hgrant1 & ~n15827;
  assign n15829 = ~n15824 & ~n15828;
  assign n15830 = ~i_hbusreq3 & ~n15829;
  assign n15831 = ~n13262 & ~n15830;
  assign n15832 = ~controllable_hgrant3 & ~n15831;
  assign n15833 = ~n15823 & ~n15832;
  assign n15834 = ~i_hbusreq9 & ~n15833;
  assign n15835 = ~n13260 & ~n15834;
  assign n15836 = ~i_hbusreq4 & ~n15835;
  assign n15837 = ~n13259 & ~n15836;
  assign n15838 = ~controllable_hgrant4 & ~n15837;
  assign n15839 = ~n15822 & ~n15838;
  assign n15840 = ~i_hbusreq5 & ~n15839;
  assign n15841 = ~n13257 & ~n15840;
  assign n15842 = ~controllable_hgrant5 & ~n15841;
  assign n15843 = ~n15821 & ~n15842;
  assign n15844 = ~controllable_hmaster2 & ~n15843;
  assign n15845 = ~n15820 & ~n15844;
  assign n15846 = ~controllable_hmaster1 & ~n15845;
  assign n15847 = ~n15819 & ~n15846;
  assign n15848 = ~i_hbusreq6 & ~n15847;
  assign n15849 = ~n13299 & ~n15848;
  assign n15850 = ~controllable_hgrant6 & ~n15849;
  assign n15851 = ~n15818 & ~n15850;
  assign n15852 = ~controllable_hmaster0 & ~n15851;
  assign n15853 = ~n15817 & ~n15852;
  assign n15854 = ~i_hbusreq8 & ~n15853;
  assign n15855 = ~n13297 & ~n15854;
  assign n15856 = ~controllable_hmaster3 & ~n15855;
  assign n15857 = ~n15811 & ~n15856;
  assign n15858 = ~i_hbusreq7 & ~n15857;
  assign n15859 = ~n15724 & ~n15858;
  assign n15860 = n7924 & ~n15859;
  assign n15861 = ~n15714 & ~n15860;
  assign n15862 = n8214 & ~n15861;
  assign n15863 = ~n15660 & ~n15862;
  assign n15864 = n8202 & ~n15863;
  assign n15865 = ~n10721 & ~n15864;
  assign n15866 = n7920 & ~n15865;
  assign n15867 = ~n10671 & ~n15866;
  assign n15868 = n7728 & ~n15867;
  assign n15869 = ~n10812 & ~n15170;
  assign n15870 = ~n8214 & ~n15869;
  assign n15871 = n8214 & ~n15171;
  assign n15872 = ~n15870 & ~n15871;
  assign n15873 = n8202 & ~n15872;
  assign n15874 = ~n10811 & ~n15873;
  assign n15875 = n7920 & ~n15874;
  assign n15876 = ~n10797 & ~n15875;
  assign n15877 = ~n7728 & ~n15876;
  assign n15878 = ~n15868 & ~n15877;
  assign n15879 = ~n7723 & ~n15878;
  assign n15880 = ~n7723 & ~n15879;
  assign n15881 = ~n7714 & ~n15880;
  assign n15882 = ~n7714 & ~n15881;
  assign n15883 = n7705 & ~n15882;
  assign n15884 = ~n10833 & ~n13651;
  assign n15885 = i_hbusreq7 & ~n15884;
  assign n15886 = ~n10847 & ~n13662;
  assign n15887 = ~i_hbusreq7 & ~n15886;
  assign n15888 = ~n15885 & ~n15887;
  assign n15889 = ~n7924 & ~n15888;
  assign n15890 = controllable_hgrant6 & ~n10830;
  assign n15891 = ~n13887 & ~n15294;
  assign n15892 = ~controllable_hmaster1 & ~n15891;
  assign n15893 = ~n15194 & ~n15892;
  assign n15894 = ~controllable_hgrant6 & ~n15893;
  assign n15895 = ~n15890 & ~n15894;
  assign n15896 = controllable_hmaster0 & ~n15895;
  assign n15897 = ~n13682 & ~n15896;
  assign n15898 = ~controllable_hmaster3 & ~n15897;
  assign n15899 = ~n13672 & ~n15898;
  assign n15900 = i_hbusreq7 & ~n15899;
  assign n15901 = i_hbusreq8 & ~n15897;
  assign n15902 = controllable_hgrant6 & ~n10842;
  assign n15903 = i_hbusreq6 & ~n15893;
  assign n15904 = i_hlock1 & ~n13543;
  assign n15905 = ~i_hlock1 & ~n13582;
  assign n15906 = ~n15904 & ~n15905;
  assign n15907 = ~i_hbusreq1 & ~n15906;
  assign n15908 = ~n14142 & ~n15907;
  assign n15909 = ~controllable_hgrant1 & ~n15908;
  assign n15910 = ~n15032 & ~n15909;
  assign n15911 = ~i_hbusreq3 & ~n15910;
  assign n15912 = ~n14140 & ~n15911;
  assign n15913 = ~controllable_hgrant3 & ~n15912;
  assign n15914 = ~n15031 & ~n15913;
  assign n15915 = ~i_hbusreq9 & ~n15914;
  assign n15916 = ~n14138 & ~n15915;
  assign n15917 = ~i_hbusreq4 & ~n15916;
  assign n15918 = ~n14137 & ~n15917;
  assign n15919 = ~controllable_hgrant4 & ~n15918;
  assign n15920 = ~n15030 & ~n15919;
  assign n15921 = ~i_hbusreq5 & ~n15920;
  assign n15922 = ~n14135 & ~n15921;
  assign n15923 = ~controllable_hgrant5 & ~n15922;
  assign n15924 = ~n15029 & ~n15923;
  assign n15925 = ~controllable_hmaster2 & ~n15924;
  assign n15926 = ~n15308 & ~n15925;
  assign n15927 = ~controllable_hmaster1 & ~n15926;
  assign n15928 = ~n15208 & ~n15927;
  assign n15929 = ~i_hbusreq6 & ~n15928;
  assign n15930 = ~n15903 & ~n15929;
  assign n15931 = ~controllable_hgrant6 & ~n15930;
  assign n15932 = ~n15902 & ~n15931;
  assign n15933 = controllable_hmaster0 & ~n15932;
  assign n15934 = ~n13728 & ~n15933;
  assign n15935 = ~i_hbusreq8 & ~n15934;
  assign n15936 = ~n15901 & ~n15935;
  assign n15937 = ~controllable_hmaster3 & ~n15936;
  assign n15938 = ~n13714 & ~n15937;
  assign n15939 = ~i_hbusreq7 & ~n15938;
  assign n15940 = ~n15900 & ~n15939;
  assign n15941 = n7924 & ~n15940;
  assign n15942 = ~n15889 & ~n15941;
  assign n15943 = ~n8214 & ~n15942;
  assign n15944 = ~n10857 & ~n13651;
  assign n15945 = i_hbusreq7 & ~n15944;
  assign n15946 = controllable_hgrant6 & ~n10864;
  assign n15947 = ~n9600 & ~n15697;
  assign n15948 = ~controllable_hmaster1 & ~n15947;
  assign n15949 = ~n9599 & ~n15948;
  assign n15950 = ~i_hbusreq6 & ~n15949;
  assign n15951 = ~n13338 & ~n15950;
  assign n15952 = ~controllable_hgrant6 & ~n15951;
  assign n15953 = ~n15946 & ~n15952;
  assign n15954 = controllable_hmaster0 & ~n15953;
  assign n15955 = ~controllable_hmaster0 & ~n10864;
  assign n15956 = ~n15954 & ~n15955;
  assign n15957 = ~i_hbusreq8 & ~n15956;
  assign n15958 = ~n13658 & ~n15957;
  assign n15959 = controllable_hmaster3 & ~n15958;
  assign n15960 = ~n10879 & ~n15959;
  assign n15961 = ~i_hbusreq7 & ~n15960;
  assign n15962 = ~n15945 & ~n15961;
  assign n15963 = ~n7924 & ~n15962;
  assign n15964 = controllable_hgrant6 & ~n10854;
  assign n15965 = ~n13934 & ~n15294;
  assign n15966 = ~controllable_hmaster1 & ~n15965;
  assign n15967 = ~n15194 & ~n15966;
  assign n15968 = ~controllable_hgrant6 & ~n15967;
  assign n15969 = ~n15964 & ~n15968;
  assign n15970 = ~controllable_hmaster0 & ~n15969;
  assign n15971 = ~n13765 & ~n15970;
  assign n15972 = ~controllable_hmaster3 & ~n15971;
  assign n15973 = ~n13672 & ~n15972;
  assign n15974 = i_hbusreq7 & ~n15973;
  assign n15975 = ~n14918 & ~n15771;
  assign n15976 = ~controllable_hmaster1 & ~n15975;
  assign n15977 = ~n14917 & ~n15976;
  assign n15978 = ~i_hbusreq6 & ~n15977;
  assign n15979 = ~n13453 & ~n15978;
  assign n15980 = ~controllable_hgrant6 & ~n15979;
  assign n15981 = ~n15946 & ~n15980;
  assign n15982 = controllable_hmaster0 & ~n15981;
  assign n15983 = ~n14918 & ~n15799;
  assign n15984 = ~controllable_hmaster1 & ~n15983;
  assign n15985 = ~n14917 & ~n15984;
  assign n15986 = ~i_hbusreq6 & ~n15985;
  assign n15987 = ~n13255 & ~n15986;
  assign n15988 = ~controllable_hgrant6 & ~n15987;
  assign n15989 = ~n15946 & ~n15988;
  assign n15990 = ~controllable_hmaster0 & ~n15989;
  assign n15991 = ~n15982 & ~n15990;
  assign n15992 = ~i_hbusreq8 & ~n15991;
  assign n15993 = ~n13701 & ~n15992;
  assign n15994 = controllable_hmaster3 & ~n15993;
  assign n15995 = i_hbusreq8 & ~n15971;
  assign n15996 = controllable_hgrant6 & ~n10874;
  assign n15997 = i_hbusreq6 & ~n15967;
  assign n15998 = ~n15130 & ~n15820;
  assign n15999 = ~controllable_hmaster1 & ~n15998;
  assign n16000 = ~n15819 & ~n15999;
  assign n16001 = ~i_hbusreq6 & ~n16000;
  assign n16002 = ~n15997 & ~n16001;
  assign n16003 = ~controllable_hgrant6 & ~n16002;
  assign n16004 = ~n15996 & ~n16003;
  assign n16005 = ~controllable_hmaster0 & ~n16004;
  assign n16006 = ~n15817 & ~n16005;
  assign n16007 = ~i_hbusreq8 & ~n16006;
  assign n16008 = ~n15995 & ~n16007;
  assign n16009 = ~controllable_hmaster3 & ~n16008;
  assign n16010 = ~n15994 & ~n16009;
  assign n16011 = ~i_hbusreq7 & ~n16010;
  assign n16012 = ~n15974 & ~n16011;
  assign n16013 = n7924 & ~n16012;
  assign n16014 = ~n15963 & ~n16013;
  assign n16015 = n8214 & ~n16014;
  assign n16016 = ~n15943 & ~n16015;
  assign n16017 = ~n8202 & ~n16016;
  assign n16018 = n8202 & ~n15171;
  assign n16019 = ~n16017 & ~n16018;
  assign n16020 = n7920 & ~n16019;
  assign n16021 = ~n10797 & ~n16020;
  assign n16022 = n7728 & ~n16021;
  assign n16023 = ~n10900 & ~n14721;
  assign n16024 = i_hlock7 & ~n16023;
  assign n16025 = ~n10910 & ~n14721;
  assign n16026 = ~i_hlock7 & ~n16025;
  assign n16027 = ~n16024 & ~n16026;
  assign n16028 = ~i_hbusreq7 & ~n16027;
  assign n16029 = ~n13816 & ~n16028;
  assign n16030 = ~n7924 & ~n16029;
  assign n16031 = controllable_hgrant6 & ~n10895;
  assign n16032 = i_hlock1 & ~n14454;
  assign n16033 = ~i_hlock1 & ~n14485;
  assign n16034 = ~n16032 & ~n16033;
  assign n16035 = ~i_hbusreq1 & ~n16034;
  assign n16036 = ~n14142 & ~n16035;
  assign n16037 = ~controllable_hgrant1 & ~n16036;
  assign n16038 = ~n15032 & ~n16037;
  assign n16039 = ~i_hbusreq3 & ~n16038;
  assign n16040 = ~n14140 & ~n16039;
  assign n16041 = ~controllable_hgrant3 & ~n16040;
  assign n16042 = ~n15031 & ~n16041;
  assign n16043 = ~i_hbusreq9 & ~n16042;
  assign n16044 = ~n14138 & ~n16043;
  assign n16045 = ~i_hbusreq4 & ~n16044;
  assign n16046 = ~n14137 & ~n16045;
  assign n16047 = ~controllable_hgrant4 & ~n16046;
  assign n16048 = ~n15030 & ~n16047;
  assign n16049 = ~i_hbusreq5 & ~n16048;
  assign n16050 = ~n14135 & ~n16049;
  assign n16051 = ~controllable_hgrant5 & ~n16050;
  assign n16052 = ~n15029 & ~n16051;
  assign n16053 = ~controllable_hmaster2 & ~n16052;
  assign n16054 = ~n14581 & ~n16053;
  assign n16055 = ~controllable_hmaster1 & ~n16054;
  assign n16056 = ~n14563 & ~n16055;
  assign n16057 = ~i_hbusreq6 & ~n16056;
  assign n16058 = ~n14095 & ~n16057;
  assign n16059 = ~controllable_hgrant6 & ~n16058;
  assign n16060 = ~n16031 & ~n16059;
  assign n16061 = controllable_hmaster0 & ~n16060;
  assign n16062 = ~n14685 & ~n16061;
  assign n16063 = ~i_hbusreq8 & ~n16062;
  assign n16064 = ~n14093 & ~n16063;
  assign n16065 = ~controllable_hmaster3 & ~n16064;
  assign n16066 = ~n14755 & ~n16065;
  assign n16067 = i_hlock7 & ~n16066;
  assign n16068 = controllable_hgrant6 & ~n10905;
  assign n16069 = ~n14693 & ~n16055;
  assign n16070 = ~i_hbusreq6 & ~n16069;
  assign n16071 = ~n14299 & ~n16070;
  assign n16072 = ~controllable_hgrant6 & ~n16071;
  assign n16073 = ~n16068 & ~n16072;
  assign n16074 = controllable_hmaster0 & ~n16073;
  assign n16075 = ~n14685 & ~n16074;
  assign n16076 = ~i_hbusreq8 & ~n16075;
  assign n16077 = ~n14297 & ~n16076;
  assign n16078 = ~controllable_hmaster3 & ~n16077;
  assign n16079 = ~n14755 & ~n16078;
  assign n16080 = ~i_hlock7 & ~n16079;
  assign n16081 = ~n16067 & ~n16080;
  assign n16082 = ~i_hbusreq7 & ~n16081;
  assign n16083 = ~n13963 & ~n16082;
  assign n16084 = n7924 & ~n16083;
  assign n16085 = ~n16030 & ~n16084;
  assign n16086 = ~n8214 & ~n16085;
  assign n16087 = ~n15871 & ~n16086;
  assign n16088 = ~n8202 & ~n16087;
  assign n16089 = ~n16018 & ~n16088;
  assign n16090 = n7920 & ~n16089;
  assign n16091 = ~n10797 & ~n16090;
  assign n16092 = ~n7728 & ~n16091;
  assign n16093 = ~n16022 & ~n16092;
  assign n16094 = n7723 & ~n16093;
  assign n16095 = ~n7723 & ~n16091;
  assign n16096 = ~n16094 & ~n16095;
  assign n16097 = n7714 & ~n16096;
  assign n16098 = n7723 & ~n16091;
  assign n16099 = ~n8640 & ~n16090;
  assign n16100 = n7728 & ~n16099;
  assign n16101 = ~n15174 & ~n16100;
  assign n16102 = ~n7723 & ~n16101;
  assign n16103 = ~n16098 & ~n16102;
  assign n16104 = ~n7714 & ~n16103;
  assign n16105 = ~n16097 & ~n16104;
  assign n16106 = ~n7705 & ~n16105;
  assign n16107 = ~n15883 & ~n16106;
  assign n16108 = n7808 & ~n16107;
  assign n16109 = ~n10670 & ~n16108;
  assign n16110 = n8195 & ~n16109;
  assign n16111 = ~n15658 & ~n16110;
  assign n16112 = n8193 & ~n16111;
  assign n16113 = ~n15186 & ~n16112;
  assign n16114 = n8191 & ~n16113;
  assign n16115 = controllable_hgrant6 & ~n10951;
  assign n16116 = controllable_hgrant5 & ~n10947;
  assign n16117 = controllable_hgrant4 & ~n10947;
  assign n16118 = controllable_hgrant3 & ~n8223;
  assign n16119 = controllable_hgrant1 & ~n8223;
  assign n16120 = controllable_locked & controllable_hmastlock;
  assign n16121 = ~n7818 & ~n7860;
  assign n16122 = ~controllable_locked & n16121;
  assign n16123 = ~n16120 & ~n16122;
  assign n16124 = ~controllable_hgrant2 & n16123;
  assign n16125 = ~n12612 & ~n16124;
  assign n16126 = ~n7733 & ~n16125;
  assign n16127 = ~n7733 & ~n16126;
  assign n16128 = ~n7928 & ~n16127;
  assign n16129 = n7928 & ~n16125;
  assign n16130 = ~n16128 & ~n16129;
  assign n16131 = ~controllable_hgrant1 & ~n16130;
  assign n16132 = ~n16119 & ~n16131;
  assign n16133 = ~controllable_hgrant3 & ~n16132;
  assign n16134 = ~n16118 & ~n16133;
  assign n16135 = i_hlock9 & ~n16134;
  assign n16136 = controllable_hgrant3 & ~n8237;
  assign n16137 = controllable_hgrant1 & ~n8237;
  assign n16138 = ~n7815 & ~n7858;
  assign n16139 = controllable_locked & ~n16138;
  assign n16140 = ~controllable_locked & ~controllable_hmastlock;
  assign n16141 = ~n16139 & ~n16140;
  assign n16142 = ~controllable_hgrant2 & n16141;
  assign n16143 = ~n12639 & ~n16142;
  assign n16144 = ~n7733 & ~n16143;
  assign n16145 = ~n7733 & ~n16144;
  assign n16146 = ~n7928 & ~n16145;
  assign n16147 = n7928 & ~n16143;
  assign n16148 = ~n16146 & ~n16147;
  assign n16149 = ~controllable_hgrant1 & ~n16148;
  assign n16150 = ~n16137 & ~n16149;
  assign n16151 = ~controllable_hgrant3 & ~n16150;
  assign n16152 = ~n16136 & ~n16151;
  assign n16153 = ~i_hlock9 & ~n16152;
  assign n16154 = ~n16135 & ~n16153;
  assign n16155 = ~controllable_hgrant4 & ~n16154;
  assign n16156 = ~n16117 & ~n16155;
  assign n16157 = ~controllable_hgrant5 & ~n16156;
  assign n16158 = ~n16116 & ~n16157;
  assign n16159 = ~controllable_hmaster2 & ~n16158;
  assign n16160 = ~controllable_hmaster2 & ~n16159;
  assign n16161 = ~controllable_hmaster1 & ~n16160;
  assign n16162 = ~controllable_hmaster1 & ~n16161;
  assign n16163 = ~controllable_hgrant6 & ~n16162;
  assign n16164 = ~n16115 & ~n16163;
  assign n16165 = controllable_hmaster0 & ~n16164;
  assign n16166 = controllable_hmaster0 & ~n16165;
  assign n16167 = controllable_hmaster3 & ~n16166;
  assign n16168 = controllable_hmaster3 & ~n16167;
  assign n16169 = i_hbusreq7 & ~n16168;
  assign n16170 = i_hbusreq8 & ~n16166;
  assign n16171 = controllable_hgrant6 & ~n10976;
  assign n16172 = i_hbusreq6 & ~n16162;
  assign n16173 = controllable_hgrant5 & ~n10970;
  assign n16174 = i_hbusreq5 & ~n16156;
  assign n16175 = controllable_hgrant4 & ~n10968;
  assign n16176 = i_hbusreq4 & ~n16154;
  assign n16177 = i_hbusreq9 & ~n16154;
  assign n16178 = controllable_hgrant3 & ~n8271;
  assign n16179 = i_hbusreq3 & ~n16132;
  assign n16180 = controllable_hgrant1 & ~n8269;
  assign n16181 = i_hbusreq1 & ~n16130;
  assign n16182 = i_hbusreq2 & ~n16123;
  assign n16183 = i_hbusreq0 & ~n16123;
  assign n16184 = ~n7864 & ~n16183;
  assign n16185 = ~i_hbusreq2 & ~n16184;
  assign n16186 = ~n16182 & ~n16185;
  assign n16187 = ~controllable_hgrant2 & n16186;
  assign n16188 = ~n12683 & ~n16187;
  assign n16189 = ~n7733 & ~n16188;
  assign n16190 = ~n7733 & ~n16189;
  assign n16191 = ~n7928 & ~n16190;
  assign n16192 = n7928 & ~n16188;
  assign n16193 = ~n16191 & ~n16192;
  assign n16194 = ~i_hbusreq1 & ~n16193;
  assign n16195 = ~n16181 & ~n16194;
  assign n16196 = ~controllable_hgrant1 & ~n16195;
  assign n16197 = ~n16180 & ~n16196;
  assign n16198 = ~i_hbusreq3 & ~n16197;
  assign n16199 = ~n16179 & ~n16198;
  assign n16200 = ~controllable_hgrant3 & ~n16199;
  assign n16201 = ~n16178 & ~n16200;
  assign n16202 = i_hlock9 & ~n16201;
  assign n16203 = controllable_hgrant3 & ~n8303;
  assign n16204 = i_hbusreq3 & ~n16150;
  assign n16205 = controllable_hgrant1 & ~n8301;
  assign n16206 = i_hbusreq1 & ~n16148;
  assign n16207 = i_hbusreq2 & ~n16141;
  assign n16208 = i_hbusreq0 & ~n16141;
  assign n16209 = ~n7864 & ~n16208;
  assign n16210 = ~i_hbusreq2 & ~n16209;
  assign n16211 = ~n16207 & ~n16210;
  assign n16212 = ~controllable_hgrant2 & n16211;
  assign n16213 = ~n12732 & ~n16212;
  assign n16214 = ~n7733 & ~n16213;
  assign n16215 = ~n7733 & ~n16214;
  assign n16216 = ~n7928 & ~n16215;
  assign n16217 = n7928 & ~n16213;
  assign n16218 = ~n16216 & ~n16217;
  assign n16219 = ~i_hbusreq1 & ~n16218;
  assign n16220 = ~n16206 & ~n16219;
  assign n16221 = ~controllable_hgrant1 & ~n16220;
  assign n16222 = ~n16205 & ~n16221;
  assign n16223 = ~i_hbusreq3 & ~n16222;
  assign n16224 = ~n16204 & ~n16223;
  assign n16225 = ~controllable_hgrant3 & ~n16224;
  assign n16226 = ~n16203 & ~n16225;
  assign n16227 = ~i_hlock9 & ~n16226;
  assign n16228 = ~n16202 & ~n16227;
  assign n16229 = ~i_hbusreq9 & ~n16228;
  assign n16230 = ~n16177 & ~n16229;
  assign n16231 = ~i_hbusreq4 & ~n16230;
  assign n16232 = ~n16176 & ~n16231;
  assign n16233 = ~controllable_hgrant4 & ~n16232;
  assign n16234 = ~n16175 & ~n16233;
  assign n16235 = ~i_hbusreq5 & ~n16234;
  assign n16236 = ~n16174 & ~n16235;
  assign n16237 = ~controllable_hgrant5 & ~n16236;
  assign n16238 = ~n16173 & ~n16237;
  assign n16239 = ~controllable_hmaster2 & ~n16238;
  assign n16240 = ~controllable_hmaster2 & ~n16239;
  assign n16241 = ~controllable_hmaster1 & ~n16240;
  assign n16242 = ~controllable_hmaster1 & ~n16241;
  assign n16243 = ~i_hbusreq6 & ~n16242;
  assign n16244 = ~n16172 & ~n16243;
  assign n16245 = ~controllable_hgrant6 & ~n16244;
  assign n16246 = ~n16171 & ~n16245;
  assign n16247 = controllable_hmaster0 & ~n16246;
  assign n16248 = controllable_hmaster0 & ~n16247;
  assign n16249 = ~i_hbusreq8 & ~n16248;
  assign n16250 = ~n16170 & ~n16249;
  assign n16251 = controllable_hmaster3 & ~n16250;
  assign n16252 = controllable_hmaster3 & ~n16251;
  assign n16253 = ~i_hbusreq7 & ~n16252;
  assign n16254 = ~n16169 & ~n16253;
  assign n16255 = n7924 & ~n16254;
  assign n16256 = n7924 & ~n16255;
  assign n16257 = ~n8214 & ~n16256;
  assign n16258 = ~n8214 & ~n16257;
  assign n16259 = ~n8202 & ~n16258;
  assign n16260 = ~n8332 & ~n16259;
  assign n16261 = n7728 & ~n16260;
  assign n16262 = controllable_hgrant6 & ~n10994;
  assign n16263 = ~n7739 & ~n16159;
  assign n16264 = ~controllable_hmaster1 & ~n16263;
  assign n16265 = ~n7738 & ~n16264;
  assign n16266 = ~controllable_hgrant6 & ~n16265;
  assign n16267 = ~n16262 & ~n16266;
  assign n16268 = controllable_hmaster0 & ~n16267;
  assign n16269 = ~n8882 & ~n16268;
  assign n16270 = controllable_hmaster3 & ~n16269;
  assign n16271 = controllable_hmaster3 & ~n16270;
  assign n16272 = i_hbusreq7 & ~n16271;
  assign n16273 = i_hbusreq8 & ~n16269;
  assign n16274 = controllable_hgrant6 & ~n11006;
  assign n16275 = i_hbusreq6 & ~n16265;
  assign n16276 = ~n7771 & ~n16239;
  assign n16277 = ~controllable_hmaster1 & ~n16276;
  assign n16278 = ~n7770 & ~n16277;
  assign n16279 = ~i_hbusreq6 & ~n16278;
  assign n16280 = ~n16275 & ~n16279;
  assign n16281 = ~controllable_hgrant6 & ~n16280;
  assign n16282 = ~n16274 & ~n16281;
  assign n16283 = controllable_hmaster0 & ~n16282;
  assign n16284 = ~n8895 & ~n16283;
  assign n16285 = ~i_hbusreq8 & ~n16284;
  assign n16286 = ~n16273 & ~n16285;
  assign n16287 = controllable_hmaster3 & ~n16286;
  assign n16288 = controllable_hmaster3 & ~n16287;
  assign n16289 = ~i_hbusreq7 & ~n16288;
  assign n16290 = ~n16272 & ~n16289;
  assign n16291 = n7924 & ~n16290;
  assign n16292 = ~n8337 & ~n16291;
  assign n16293 = ~n8214 & ~n16292;
  assign n16294 = ~n11018 & ~n16293;
  assign n16295 = ~n8202 & ~n16294;
  assign n16296 = ~n8347 & ~n16295;
  assign n16297 = ~n7728 & ~n16296;
  assign n16298 = ~n16261 & ~n16297;
  assign n16299 = ~n7723 & ~n16298;
  assign n16300 = ~n7723 & ~n16299;
  assign n16301 = ~n7714 & ~n16300;
  assign n16302 = ~n7714 & ~n16301;
  assign n16303 = n7705 & ~n16302;
  assign n16304 = n7723 & ~n16296;
  assign n16305 = controllable_hgrant6 & ~n11032;
  assign n16306 = ~n8358 & ~n16159;
  assign n16307 = ~controllable_hmaster1 & ~n16306;
  assign n16308 = ~n8357 & ~n16307;
  assign n16309 = ~controllable_hgrant6 & ~n16308;
  assign n16310 = ~n16305 & ~n16309;
  assign n16311 = controllable_hmaster0 & ~n16310;
  assign n16312 = ~n11034 & ~n16311;
  assign n16313 = controllable_hmaster3 & ~n16312;
  assign n16314 = ~n8463 & ~n16313;
  assign n16315 = i_hbusreq7 & ~n16314;
  assign n16316 = i_hbusreq8 & ~n16312;
  assign n16317 = controllable_hgrant6 & ~n11045;
  assign n16318 = i_hbusreq6 & ~n16308;
  assign n16319 = ~n8484 & ~n16239;
  assign n16320 = ~controllable_hmaster1 & ~n16319;
  assign n16321 = ~n8483 & ~n16320;
  assign n16322 = ~i_hbusreq6 & ~n16321;
  assign n16323 = ~n16318 & ~n16322;
  assign n16324 = ~controllable_hgrant6 & ~n16323;
  assign n16325 = ~n16317 & ~n16324;
  assign n16326 = controllable_hmaster0 & ~n16325;
  assign n16327 = ~n11047 & ~n16326;
  assign n16328 = ~i_hbusreq8 & ~n16327;
  assign n16329 = ~n16316 & ~n16328;
  assign n16330 = controllable_hmaster3 & ~n16329;
  assign n16331 = ~n8634 & ~n16330;
  assign n16332 = ~i_hbusreq7 & ~n16331;
  assign n16333 = ~n16315 & ~n16332;
  assign n16334 = n7924 & ~n16333;
  assign n16335 = ~n8337 & ~n16334;
  assign n16336 = ~n7920 & ~n16335;
  assign n16337 = n7920 & ~n16296;
  assign n16338 = ~n16336 & ~n16337;
  assign n16339 = ~n7723 & ~n16338;
  assign n16340 = ~n16304 & ~n16339;
  assign n16341 = n7714 & ~n16340;
  assign n16342 = ~n7714 & ~n16335;
  assign n16343 = ~n16341 & ~n16342;
  assign n16344 = ~n7705 & ~n16343;
  assign n16345 = ~n16303 & ~n16344;
  assign n16346 = ~n7808 & ~n16345;
  assign n16347 = ~n7920 & ~n16260;
  assign n16348 = ~n7817 & ~n7934;
  assign n16349 = ~controllable_hgrant2 & n16348;
  assign n16350 = ~n7814 & ~n16349;
  assign n16351 = ~n7733 & ~n16350;
  assign n16352 = n7733 & ~n7937;
  assign n16353 = ~n16351 & ~n16352;
  assign n16354 = n7928 & ~n16353;
  assign n16355 = ~n16128 & ~n16354;
  assign n16356 = ~controllable_hgrant1 & ~n16355;
  assign n16357 = ~n12611 & ~n16356;
  assign n16358 = ~controllable_hgrant3 & ~n16357;
  assign n16359 = ~n12610 & ~n16358;
  assign n16360 = i_hlock9 & ~n16359;
  assign n16361 = ~n16146 & ~n16354;
  assign n16362 = ~controllable_hgrant1 & ~n16361;
  assign n16363 = ~n12638 & ~n16362;
  assign n16364 = ~controllable_hgrant3 & ~n16363;
  assign n16365 = ~n12637 & ~n16364;
  assign n16366 = ~i_hlock9 & ~n16365;
  assign n16367 = ~n16360 & ~n16366;
  assign n16368 = ~controllable_hgrant4 & ~n16367;
  assign n16369 = ~n12609 & ~n16368;
  assign n16370 = ~controllable_hgrant5 & ~n16369;
  assign n16371 = ~n12608 & ~n16370;
  assign n16372 = ~controllable_hmaster2 & ~n16371;
  assign n16373 = ~controllable_hmaster2 & ~n16372;
  assign n16374 = ~controllable_hmaster1 & ~n16373;
  assign n16375 = ~controllable_hmaster1 & ~n16374;
  assign n16376 = ~controllable_hgrant6 & ~n16375;
  assign n16377 = ~n12607 & ~n16376;
  assign n16378 = controllable_hmaster0 & ~n16377;
  assign n16379 = controllable_hmaster0 & ~n16378;
  assign n16380 = controllable_hmaster3 & ~n16379;
  assign n16381 = controllable_hmaster3 & ~n16380;
  assign n16382 = i_hbusreq7 & ~n16381;
  assign n16383 = i_hbusreq8 & ~n16379;
  assign n16384 = i_hbusreq6 & ~n16375;
  assign n16385 = i_hbusreq5 & ~n16369;
  assign n16386 = i_hbusreq4 & ~n16367;
  assign n16387 = i_hbusreq9 & ~n16367;
  assign n16388 = i_hbusreq3 & ~n16357;
  assign n16389 = i_hbusreq1 & ~n16355;
  assign n16390 = i_hbusreq2 & ~n16348;
  assign n16391 = i_hbusreq0 & ~n16348;
  assign n16392 = ~n7859 & ~n7977;
  assign n16393 = i_hlock0 & ~n16392;
  assign n16394 = ~i_hlock0 & ~n16348;
  assign n16395 = ~n16393 & ~n16394;
  assign n16396 = ~i_hbusreq0 & ~n16395;
  assign n16397 = ~n16391 & ~n16396;
  assign n16398 = ~i_hbusreq2 & ~n16397;
  assign n16399 = ~n16390 & ~n16398;
  assign n16400 = ~controllable_hgrant2 & n16399;
  assign n16401 = ~n12694 & ~n16400;
  assign n16402 = ~n7733 & ~n16401;
  assign n16403 = ~n7858 & ~n7930;
  assign n16404 = controllable_locked & ~n16403;
  assign n16405 = ~controllable_locked & ~n7975;
  assign n16406 = ~n16404 & ~n16405;
  assign n16407 = i_hlock0 & ~n16406;
  assign n16408 = ~i_hlock0 & ~n7935;
  assign n16409 = ~n16407 & ~n16408;
  assign n16410 = ~i_hbusreq0 & ~n16409;
  assign n16411 = ~n7969 & ~n16410;
  assign n16412 = ~i_hbusreq2 & ~n16411;
  assign n16413 = ~n7968 & ~n16412;
  assign n16414 = ~controllable_hgrant2 & n16413;
  assign n16415 = ~n12706 & ~n16414;
  assign n16416 = n7733 & ~n16415;
  assign n16417 = ~n16402 & ~n16416;
  assign n16418 = n7928 & ~n16417;
  assign n16419 = ~n16191 & ~n16418;
  assign n16420 = ~i_hbusreq1 & ~n16419;
  assign n16421 = ~n16389 & ~n16420;
  assign n16422 = ~controllable_hgrant1 & ~n16421;
  assign n16423 = ~n12681 & ~n16422;
  assign n16424 = ~i_hbusreq3 & ~n16423;
  assign n16425 = ~n16388 & ~n16424;
  assign n16426 = ~controllable_hgrant3 & ~n16425;
  assign n16427 = ~n12679 & ~n16426;
  assign n16428 = i_hlock9 & ~n16427;
  assign n16429 = i_hbusreq3 & ~n16363;
  assign n16430 = i_hbusreq1 & ~n16361;
  assign n16431 = ~n16216 & ~n16418;
  assign n16432 = ~i_hbusreq1 & ~n16431;
  assign n16433 = ~n16430 & ~n16432;
  assign n16434 = ~controllable_hgrant1 & ~n16433;
  assign n16435 = ~n12730 & ~n16434;
  assign n16436 = ~i_hbusreq3 & ~n16435;
  assign n16437 = ~n16429 & ~n16436;
  assign n16438 = ~controllable_hgrant3 & ~n16437;
  assign n16439 = ~n12728 & ~n16438;
  assign n16440 = ~i_hlock9 & ~n16439;
  assign n16441 = ~n16428 & ~n16440;
  assign n16442 = ~i_hbusreq9 & ~n16441;
  assign n16443 = ~n16387 & ~n16442;
  assign n16444 = ~i_hbusreq4 & ~n16443;
  assign n16445 = ~n16386 & ~n16444;
  assign n16446 = ~controllable_hgrant4 & ~n16445;
  assign n16447 = ~n12676 & ~n16446;
  assign n16448 = ~i_hbusreq5 & ~n16447;
  assign n16449 = ~n16385 & ~n16448;
  assign n16450 = ~controllable_hgrant5 & ~n16449;
  assign n16451 = ~n12674 & ~n16450;
  assign n16452 = ~controllable_hmaster2 & ~n16451;
  assign n16453 = ~controllable_hmaster2 & ~n16452;
  assign n16454 = ~controllable_hmaster1 & ~n16453;
  assign n16455 = ~controllable_hmaster1 & ~n16454;
  assign n16456 = ~i_hbusreq6 & ~n16455;
  assign n16457 = ~n16384 & ~n16456;
  assign n16458 = ~controllable_hgrant6 & ~n16457;
  assign n16459 = ~n12672 & ~n16458;
  assign n16460 = controllable_hmaster0 & ~n16459;
  assign n16461 = controllable_hmaster0 & ~n16460;
  assign n16462 = ~i_hbusreq8 & ~n16461;
  assign n16463 = ~n16383 & ~n16462;
  assign n16464 = controllable_hmaster3 & ~n16463;
  assign n16465 = controllable_hmaster3 & ~n16464;
  assign n16466 = ~i_hbusreq7 & ~n16465;
  assign n16467 = ~n16382 & ~n16466;
  assign n16468 = ~n7924 & ~n16467;
  assign n16469 = ~i_hready & ~controllable_locked;
  assign n16470 = ~controllable_locked & ~n16469;
  assign n16471 = ~controllable_hgrant2 & ~n16470;
  assign n16472 = ~controllable_hgrant2 & ~n16471;
  assign n16473 = ~n7733 & ~n16472;
  assign n16474 = n7733 & ~n8038;
  assign n16475 = ~n16473 & ~n16474;
  assign n16476 = n7928 & ~n16475;
  assign n16477 = n7928 & ~n16476;
  assign n16478 = ~controllable_hgrant1 & ~n16477;
  assign n16479 = ~controllable_hgrant1 & ~n16478;
  assign n16480 = ~controllable_hgrant3 & ~n16479;
  assign n16481 = ~controllable_hgrant3 & ~n16480;
  assign n16482 = i_hlock9 & ~n16481;
  assign n16483 = controllable_locked & n7970;
  assign n16484 = i_hready & ~controllable_locked;
  assign n16485 = ~n16483 & ~n16484;
  assign n16486 = ~controllable_hgrant2 & n16485;
  assign n16487 = ~controllable_hgrant2 & ~n16486;
  assign n16488 = n7733 & ~n16487;
  assign n16489 = ~n16473 & ~n16488;
  assign n16490 = n7928 & ~n16489;
  assign n16491 = n7928 & ~n16490;
  assign n16492 = ~controllable_hgrant1 & ~n16491;
  assign n16493 = ~controllable_hgrant1 & ~n16492;
  assign n16494 = ~controllable_hgrant3 & ~n16493;
  assign n16495 = ~controllable_hgrant3 & ~n16494;
  assign n16496 = ~i_hlock9 & ~n16495;
  assign n16497 = ~n16482 & ~n16496;
  assign n16498 = ~controllable_hgrant4 & ~n16497;
  assign n16499 = ~controllable_hgrant4 & ~n16498;
  assign n16500 = ~controllable_hgrant5 & ~n16499;
  assign n16501 = ~controllable_hgrant5 & ~n16500;
  assign n16502 = controllable_hmaster1 & ~n16501;
  assign n16503 = controllable_hmaster2 & ~n16501;
  assign n16504 = controllable_locked & ~n7817;
  assign n16505 = ~controllable_hgrant2 & n16504;
  assign n16506 = ~n7814 & ~n16505;
  assign n16507 = ~n7733 & ~n16506;
  assign n16508 = n7733 & n7814;
  assign n16509 = ~n16507 & ~n16508;
  assign n16510 = n7928 & ~n16509;
  assign n16511 = ~n16128 & ~n16510;
  assign n16512 = ~controllable_hgrant1 & ~n16511;
  assign n16513 = ~n12611 & ~n16512;
  assign n16514 = ~controllable_hgrant3 & ~n16513;
  assign n16515 = ~n12610 & ~n16514;
  assign n16516 = i_hlock9 & ~n16515;
  assign n16517 = ~controllable_hmastlock & ~n14241;
  assign n16518 = controllable_locked & ~n16517;
  assign n16519 = controllable_locked & ~n16518;
  assign n16520 = ~controllable_hgrant2 & n16519;
  assign n16521 = ~n7814 & ~n16520;
  assign n16522 = n7733 & ~n16521;
  assign n16523 = ~n16507 & ~n16522;
  assign n16524 = n7928 & ~n16523;
  assign n16525 = ~n16146 & ~n16524;
  assign n16526 = ~controllable_hgrant1 & ~n16525;
  assign n16527 = ~n12638 & ~n16526;
  assign n16528 = ~controllable_hgrant3 & ~n16527;
  assign n16529 = ~n12637 & ~n16528;
  assign n16530 = ~i_hlock9 & ~n16529;
  assign n16531 = ~n16516 & ~n16530;
  assign n16532 = ~controllable_hgrant4 & ~n16531;
  assign n16533 = ~n12609 & ~n16532;
  assign n16534 = ~controllable_hgrant5 & ~n16533;
  assign n16535 = ~n12608 & ~n16534;
  assign n16536 = ~controllable_hmaster2 & ~n16535;
  assign n16537 = ~n16503 & ~n16536;
  assign n16538 = ~controllable_hmaster1 & ~n16537;
  assign n16539 = ~n16502 & ~n16538;
  assign n16540 = ~controllable_hgrant6 & ~n16539;
  assign n16541 = ~n12607 & ~n16540;
  assign n16542 = controllable_hmaster0 & ~n16541;
  assign n16543 = ~controllable_hgrant6 & ~n16501;
  assign n16544 = ~controllable_hgrant6 & ~n16543;
  assign n16545 = ~controllable_hmaster0 & ~n16544;
  assign n16546 = ~n16542 & ~n16545;
  assign n16547 = controllable_hmaster3 & ~n16546;
  assign n16548 = ~controllable_hmaster3 & ~n16544;
  assign n16549 = ~n16547 & ~n16548;
  assign n16550 = i_hbusreq7 & ~n16549;
  assign n16551 = i_hbusreq8 & ~n16546;
  assign n16552 = i_hbusreq6 & ~n16539;
  assign n16553 = i_hbusreq5 & ~n16499;
  assign n16554 = i_hbusreq4 & ~n16497;
  assign n16555 = i_hbusreq9 & ~n16497;
  assign n16556 = i_hbusreq3 & ~n16479;
  assign n16557 = i_hbusreq1 & ~n16477;
  assign n16558 = i_hbusreq2 & ~n16470;
  assign n16559 = i_hbusreq0 & ~n16470;
  assign n16560 = ~controllable_locked & ~n7970;
  assign n16561 = ~controllable_locked & ~n16560;
  assign n16562 = i_hlock0 & ~n16561;
  assign n16563 = ~i_hlock0 & ~n16470;
  assign n16564 = ~n16562 & ~n16563;
  assign n16565 = ~i_hbusreq0 & ~n16564;
  assign n16566 = ~n16559 & ~n16565;
  assign n16567 = ~i_hbusreq2 & ~n16566;
  assign n16568 = ~n16558 & ~n16567;
  assign n16569 = ~controllable_hgrant2 & ~n16568;
  assign n16570 = ~controllable_hgrant2 & ~n16569;
  assign n16571 = ~n7733 & ~n16570;
  assign n16572 = ~i_hbusreq0 & ~n16485;
  assign n16573 = ~n8106 & ~n16572;
  assign n16574 = ~i_hbusreq2 & ~n16573;
  assign n16575 = ~n8105 & ~n16574;
  assign n16576 = ~controllable_hgrant2 & n16575;
  assign n16577 = ~controllable_hgrant2 & ~n16576;
  assign n16578 = n7733 & ~n16577;
  assign n16579 = ~n16571 & ~n16578;
  assign n16580 = n7928 & ~n16579;
  assign n16581 = n7928 & ~n16580;
  assign n16582 = ~i_hbusreq1 & ~n16581;
  assign n16583 = ~n16557 & ~n16582;
  assign n16584 = ~controllable_hgrant1 & ~n16583;
  assign n16585 = ~controllable_hgrant1 & ~n16584;
  assign n16586 = ~i_hbusreq3 & ~n16585;
  assign n16587 = ~n16556 & ~n16586;
  assign n16588 = ~controllable_hgrant3 & ~n16587;
  assign n16589 = ~controllable_hgrant3 & ~n16588;
  assign n16590 = i_hlock9 & ~n16589;
  assign n16591 = i_hbusreq3 & ~n16493;
  assign n16592 = i_hbusreq1 & ~n16491;
  assign n16593 = ~n16488 & ~n16571;
  assign n16594 = n7928 & ~n16593;
  assign n16595 = n7928 & ~n16594;
  assign n16596 = ~i_hbusreq1 & ~n16595;
  assign n16597 = ~n16592 & ~n16596;
  assign n16598 = ~controllable_hgrant1 & ~n16597;
  assign n16599 = ~controllable_hgrant1 & ~n16598;
  assign n16600 = ~i_hbusreq3 & ~n16599;
  assign n16601 = ~n16591 & ~n16600;
  assign n16602 = ~controllable_hgrant3 & ~n16601;
  assign n16603 = ~controllable_hgrant3 & ~n16602;
  assign n16604 = ~i_hlock9 & ~n16603;
  assign n16605 = ~n16590 & ~n16604;
  assign n16606 = ~i_hbusreq9 & ~n16605;
  assign n16607 = ~n16555 & ~n16606;
  assign n16608 = ~i_hbusreq4 & ~n16607;
  assign n16609 = ~n16554 & ~n16608;
  assign n16610 = ~controllable_hgrant4 & ~n16609;
  assign n16611 = ~controllable_hgrant4 & ~n16610;
  assign n16612 = ~i_hbusreq5 & ~n16611;
  assign n16613 = ~n16553 & ~n16612;
  assign n16614 = ~controllable_hgrant5 & ~n16613;
  assign n16615 = ~controllable_hgrant5 & ~n16614;
  assign n16616 = controllable_hmaster1 & ~n16615;
  assign n16617 = controllable_hmaster2 & ~n16615;
  assign n16618 = i_hbusreq5 & ~n16533;
  assign n16619 = i_hbusreq4 & ~n16531;
  assign n16620 = i_hbusreq9 & ~n16531;
  assign n16621 = i_hbusreq3 & ~n16513;
  assign n16622 = i_hbusreq1 & ~n16511;
  assign n16623 = i_hbusreq2 & ~n16504;
  assign n16624 = i_hbusreq0 & ~n16504;
  assign n16625 = ~n7859 & ~n12799;
  assign n16626 = i_hlock0 & ~n16625;
  assign n16627 = ~i_hlock0 & ~n16504;
  assign n16628 = ~n16626 & ~n16627;
  assign n16629 = ~i_hbusreq0 & ~n16628;
  assign n16630 = ~n16624 & ~n16629;
  assign n16631 = ~i_hbusreq2 & ~n16630;
  assign n16632 = ~n16623 & ~n16631;
  assign n16633 = ~controllable_hgrant2 & n16632;
  assign n16634 = ~n12694 & ~n16633;
  assign n16635 = ~n7733 & ~n16634;
  assign n16636 = controllable_locked & ~n14242;
  assign n16637 = ~n12615 & ~n16636;
  assign n16638 = i_hlock0 & ~n16637;
  assign n16639 = ~i_hlock0 & ~n16519;
  assign n16640 = ~n16638 & ~n16639;
  assign n16641 = ~i_hbusreq0 & ~n16640;
  assign n16642 = ~i_hbusreq0 & ~n16641;
  assign n16643 = ~i_hbusreq2 & ~n16642;
  assign n16644 = ~i_hbusreq2 & ~n16643;
  assign n16645 = ~controllable_hgrant2 & n16644;
  assign n16646 = ~n12706 & ~n16645;
  assign n16647 = n7733 & ~n16646;
  assign n16648 = ~n16635 & ~n16647;
  assign n16649 = n7928 & ~n16648;
  assign n16650 = ~n16191 & ~n16649;
  assign n16651 = ~i_hbusreq1 & ~n16650;
  assign n16652 = ~n16622 & ~n16651;
  assign n16653 = ~controllable_hgrant1 & ~n16652;
  assign n16654 = ~n12681 & ~n16653;
  assign n16655 = ~i_hbusreq3 & ~n16654;
  assign n16656 = ~n16621 & ~n16655;
  assign n16657 = ~controllable_hgrant3 & ~n16656;
  assign n16658 = ~n12679 & ~n16657;
  assign n16659 = i_hlock9 & ~n16658;
  assign n16660 = i_hbusreq3 & ~n16527;
  assign n16661 = i_hbusreq1 & ~n16525;
  assign n16662 = i_hbusreq2 & ~n16519;
  assign n16663 = i_hbusreq0 & ~n16519;
  assign n16664 = ~n16641 & ~n16663;
  assign n16665 = ~i_hbusreq2 & ~n16664;
  assign n16666 = ~n16662 & ~n16665;
  assign n16667 = ~controllable_hgrant2 & n16666;
  assign n16668 = ~n12706 & ~n16667;
  assign n16669 = n7733 & ~n16668;
  assign n16670 = ~n16635 & ~n16669;
  assign n16671 = n7928 & ~n16670;
  assign n16672 = ~n16216 & ~n16671;
  assign n16673 = ~i_hbusreq1 & ~n16672;
  assign n16674 = ~n16661 & ~n16673;
  assign n16675 = ~controllable_hgrant1 & ~n16674;
  assign n16676 = ~n12730 & ~n16675;
  assign n16677 = ~i_hbusreq3 & ~n16676;
  assign n16678 = ~n16660 & ~n16677;
  assign n16679 = ~controllable_hgrant3 & ~n16678;
  assign n16680 = ~n12728 & ~n16679;
  assign n16681 = ~i_hlock9 & ~n16680;
  assign n16682 = ~n16659 & ~n16681;
  assign n16683 = ~i_hbusreq9 & ~n16682;
  assign n16684 = ~n16620 & ~n16683;
  assign n16685 = ~i_hbusreq4 & ~n16684;
  assign n16686 = ~n16619 & ~n16685;
  assign n16687 = ~controllable_hgrant4 & ~n16686;
  assign n16688 = ~n12676 & ~n16687;
  assign n16689 = ~i_hbusreq5 & ~n16688;
  assign n16690 = ~n16618 & ~n16689;
  assign n16691 = ~controllable_hgrant5 & ~n16690;
  assign n16692 = ~n12674 & ~n16691;
  assign n16693 = ~controllable_hmaster2 & ~n16692;
  assign n16694 = ~n16617 & ~n16693;
  assign n16695 = ~controllable_hmaster1 & ~n16694;
  assign n16696 = ~n16616 & ~n16695;
  assign n16697 = ~i_hbusreq6 & ~n16696;
  assign n16698 = ~n16552 & ~n16697;
  assign n16699 = ~controllable_hgrant6 & ~n16698;
  assign n16700 = ~n12672 & ~n16699;
  assign n16701 = controllable_hmaster0 & ~n16700;
  assign n16702 = i_hbusreq6 & ~n16501;
  assign n16703 = ~i_hbusreq6 & ~n16615;
  assign n16704 = ~n16702 & ~n16703;
  assign n16705 = ~controllable_hgrant6 & ~n16704;
  assign n16706 = ~controllable_hgrant6 & ~n16705;
  assign n16707 = ~controllable_hmaster0 & ~n16706;
  assign n16708 = ~n16701 & ~n16707;
  assign n16709 = ~i_hbusreq8 & ~n16708;
  assign n16710 = ~n16551 & ~n16709;
  assign n16711 = controllable_hmaster3 & ~n16710;
  assign n16712 = i_hbusreq8 & ~n16544;
  assign n16713 = ~i_hbusreq8 & ~n16706;
  assign n16714 = ~n16712 & ~n16713;
  assign n16715 = ~controllable_hmaster3 & ~n16714;
  assign n16716 = ~n16711 & ~n16715;
  assign n16717 = ~i_hbusreq7 & ~n16716;
  assign n16718 = ~n16550 & ~n16717;
  assign n16719 = n7924 & ~n16718;
  assign n16720 = ~n16468 & ~n16719;
  assign n16721 = ~n8214 & ~n16720;
  assign n16722 = controllable_hgrant6 & ~n8729;
  assign n16723 = ~n13008 & ~n16484;
  assign n16724 = ~controllable_hgrant2 & ~n16723;
  assign n16725 = ~n7814 & ~n16724;
  assign n16726 = ~n7733 & ~n16725;
  assign n16727 = i_hready & ~controllable_hmastlock;
  assign n16728 = ~n7818 & ~n16727;
  assign n16729 = controllable_locked & ~n16728;
  assign n16730 = ~n16484 & ~n16729;
  assign n16731 = ~controllable_hgrant2 & ~n16730;
  assign n16732 = ~n7814 & ~n16731;
  assign n16733 = n7733 & ~n16732;
  assign n16734 = ~n16726 & ~n16733;
  assign n16735 = n7928 & ~n16734;
  assign n16736 = ~n8221 & ~n16735;
  assign n16737 = ~controllable_hgrant1 & ~n16736;
  assign n16738 = ~n12611 & ~n16737;
  assign n16739 = ~controllable_hgrant3 & ~n16738;
  assign n16740 = ~n12610 & ~n16739;
  assign n16741 = ~controllable_hgrant4 & ~n16740;
  assign n16742 = ~n13408 & ~n16741;
  assign n16743 = ~controllable_hgrant5 & ~n16742;
  assign n16744 = ~n13407 & ~n16743;
  assign n16745 = ~controllable_hmaster2 & ~n16744;
  assign n16746 = ~controllable_hmaster2 & ~n16745;
  assign n16747 = ~controllable_hmaster1 & ~n16746;
  assign n16748 = ~controllable_hmaster1 & ~n16747;
  assign n16749 = ~controllable_hgrant6 & ~n16748;
  assign n16750 = ~n16722 & ~n16749;
  assign n16751 = ~controllable_hmaster0 & ~n16750;
  assign n16752 = ~controllable_hmaster0 & ~n16751;
  assign n16753 = i_hlock8 & ~n16752;
  assign n16754 = controllable_hgrant6 & ~n8736;
  assign n16755 = ~n8235 & ~n16735;
  assign n16756 = ~controllable_hgrant1 & ~n16755;
  assign n16757 = ~n12638 & ~n16756;
  assign n16758 = ~controllable_hgrant3 & ~n16757;
  assign n16759 = ~n12637 & ~n16758;
  assign n16760 = ~controllable_hgrant4 & ~n16759;
  assign n16761 = ~n13429 & ~n16760;
  assign n16762 = ~controllable_hgrant5 & ~n16761;
  assign n16763 = ~n13428 & ~n16762;
  assign n16764 = ~controllable_hmaster2 & ~n16763;
  assign n16765 = ~controllable_hmaster2 & ~n16764;
  assign n16766 = ~controllable_hmaster1 & ~n16765;
  assign n16767 = ~controllable_hmaster1 & ~n16766;
  assign n16768 = ~controllable_hgrant6 & ~n16767;
  assign n16769 = ~n16754 & ~n16768;
  assign n16770 = ~controllable_hmaster0 & ~n16769;
  assign n16771 = ~controllable_hmaster0 & ~n16770;
  assign n16772 = ~i_hlock8 & ~n16771;
  assign n16773 = ~n16753 & ~n16772;
  assign n16774 = controllable_hmaster3 & ~n16773;
  assign n16775 = controllable_hmaster3 & ~n16774;
  assign n16776 = i_hbusreq7 & ~n16775;
  assign n16777 = i_hbusreq8 & ~n16773;
  assign n16778 = controllable_hgrant6 & ~n8760;
  assign n16779 = i_hbusreq6 & ~n16748;
  assign n16780 = i_hbusreq5 & ~n16742;
  assign n16781 = i_hbusreq4 & ~n16740;
  assign n16782 = i_hbusreq9 & ~n16740;
  assign n16783 = i_hbusreq3 & ~n16738;
  assign n16784 = i_hbusreq1 & ~n16736;
  assign n16785 = i_hbusreq2 & ~n16723;
  assign n16786 = i_hbusreq0 & ~n16723;
  assign n16787 = ~controllable_locked & ~n7971;
  assign n16788 = ~controllable_locked & ~n16787;
  assign n16789 = i_hlock0 & ~n16788;
  assign n16790 = ~i_hlock0 & ~n16723;
  assign n16791 = ~n16789 & ~n16790;
  assign n16792 = ~i_hbusreq0 & ~n16791;
  assign n16793 = ~n16786 & ~n16792;
  assign n16794 = ~i_hbusreq2 & ~n16793;
  assign n16795 = ~n16785 & ~n16794;
  assign n16796 = ~controllable_hgrant2 & ~n16795;
  assign n16797 = ~n12694 & ~n16796;
  assign n16798 = ~n7733 & ~n16797;
  assign n16799 = i_hbusreq2 & ~n16730;
  assign n16800 = i_hbusreq0 & ~n16730;
  assign n16801 = ~controllable_hmastlock & ~n16727;
  assign n16802 = controllable_locked & ~n16801;
  assign n16803 = ~n7975 & ~n16727;
  assign n16804 = ~controllable_locked & ~n16803;
  assign n16805 = ~n16802 & ~n16804;
  assign n16806 = i_hlock0 & ~n16805;
  assign n16807 = ~i_hlock0 & ~n16730;
  assign n16808 = ~n16806 & ~n16807;
  assign n16809 = ~i_hbusreq0 & ~n16808;
  assign n16810 = ~n16800 & ~n16809;
  assign n16811 = ~i_hbusreq2 & ~n16810;
  assign n16812 = ~n16799 & ~n16811;
  assign n16813 = ~controllable_hgrant2 & ~n16812;
  assign n16814 = ~n12706 & ~n16813;
  assign n16815 = n7733 & ~n16814;
  assign n16816 = ~n16798 & ~n16815;
  assign n16817 = n7928 & ~n16816;
  assign n16818 = ~n8265 & ~n16817;
  assign n16819 = ~i_hbusreq1 & ~n16818;
  assign n16820 = ~n16784 & ~n16819;
  assign n16821 = ~controllable_hgrant1 & ~n16820;
  assign n16822 = ~n12681 & ~n16821;
  assign n16823 = ~i_hbusreq3 & ~n16822;
  assign n16824 = ~n16783 & ~n16823;
  assign n16825 = ~controllable_hgrant3 & ~n16824;
  assign n16826 = ~n12679 & ~n16825;
  assign n16827 = ~i_hbusreq9 & ~n16826;
  assign n16828 = ~n16782 & ~n16827;
  assign n16829 = ~i_hbusreq4 & ~n16828;
  assign n16830 = ~n16781 & ~n16829;
  assign n16831 = ~controllable_hgrant4 & ~n16830;
  assign n16832 = ~n13524 & ~n16831;
  assign n16833 = ~i_hbusreq5 & ~n16832;
  assign n16834 = ~n16780 & ~n16833;
  assign n16835 = ~controllable_hgrant5 & ~n16834;
  assign n16836 = ~n13522 & ~n16835;
  assign n16837 = ~controllable_hmaster2 & ~n16836;
  assign n16838 = ~controllable_hmaster2 & ~n16837;
  assign n16839 = ~controllable_hmaster1 & ~n16838;
  assign n16840 = ~controllable_hmaster1 & ~n16839;
  assign n16841 = ~i_hbusreq6 & ~n16840;
  assign n16842 = ~n16779 & ~n16841;
  assign n16843 = ~controllable_hgrant6 & ~n16842;
  assign n16844 = ~n16778 & ~n16843;
  assign n16845 = ~controllable_hmaster0 & ~n16844;
  assign n16846 = ~controllable_hmaster0 & ~n16845;
  assign n16847 = i_hlock8 & ~n16846;
  assign n16848 = controllable_hgrant6 & ~n8779;
  assign n16849 = i_hbusreq6 & ~n16767;
  assign n16850 = i_hbusreq5 & ~n16761;
  assign n16851 = i_hbusreq4 & ~n16759;
  assign n16852 = i_hbusreq9 & ~n16759;
  assign n16853 = i_hbusreq3 & ~n16757;
  assign n16854 = i_hbusreq1 & ~n16755;
  assign n16855 = ~n8297 & ~n16817;
  assign n16856 = ~i_hbusreq1 & ~n16855;
  assign n16857 = ~n16854 & ~n16856;
  assign n16858 = ~controllable_hgrant1 & ~n16857;
  assign n16859 = ~n12730 & ~n16858;
  assign n16860 = ~i_hbusreq3 & ~n16859;
  assign n16861 = ~n16853 & ~n16860;
  assign n16862 = ~controllable_hgrant3 & ~n16861;
  assign n16863 = ~n12728 & ~n16862;
  assign n16864 = ~i_hbusreq9 & ~n16863;
  assign n16865 = ~n16852 & ~n16864;
  assign n16866 = ~i_hbusreq4 & ~n16865;
  assign n16867 = ~n16851 & ~n16866;
  assign n16868 = ~controllable_hgrant4 & ~n16867;
  assign n16869 = ~n13577 & ~n16868;
  assign n16870 = ~i_hbusreq5 & ~n16869;
  assign n16871 = ~n16850 & ~n16870;
  assign n16872 = ~controllable_hgrant5 & ~n16871;
  assign n16873 = ~n13575 & ~n16872;
  assign n16874 = ~controllable_hmaster2 & ~n16873;
  assign n16875 = ~controllable_hmaster2 & ~n16874;
  assign n16876 = ~controllable_hmaster1 & ~n16875;
  assign n16877 = ~controllable_hmaster1 & ~n16876;
  assign n16878 = ~i_hbusreq6 & ~n16877;
  assign n16879 = ~n16849 & ~n16878;
  assign n16880 = ~controllable_hgrant6 & ~n16879;
  assign n16881 = ~n16848 & ~n16880;
  assign n16882 = ~controllable_hmaster0 & ~n16881;
  assign n16883 = ~controllable_hmaster0 & ~n16882;
  assign n16884 = ~i_hlock8 & ~n16883;
  assign n16885 = ~n16847 & ~n16884;
  assign n16886 = ~i_hbusreq8 & ~n16885;
  assign n16887 = ~n16777 & ~n16886;
  assign n16888 = controllable_hmaster3 & ~n16887;
  assign n16889 = controllable_hmaster3 & ~n16888;
  assign n16890 = ~i_hbusreq7 & ~n16889;
  assign n16891 = ~n16776 & ~n16890;
  assign n16892 = n8214 & ~n16891;
  assign n16893 = ~n16721 & ~n16892;
  assign n16894 = ~n8202 & ~n16893;
  assign n16895 = controllable_hgrant6 & ~n8796;
  assign n16896 = controllable_hmaster2 & ~n16744;
  assign n16897 = controllable_hmaster2 & ~n16896;
  assign n16898 = controllable_hmaster1 & ~n16897;
  assign n16899 = controllable_hmaster1 & ~n16898;
  assign n16900 = ~controllable_hgrant6 & ~n16899;
  assign n16901 = ~n16895 & ~n16900;
  assign n16902 = controllable_hmaster0 & ~n16901;
  assign n16903 = controllable_hmaster0 & ~n16902;
  assign n16904 = ~controllable_hmaster3 & ~n16903;
  assign n16905 = ~controllable_hmaster3 & ~n16904;
  assign n16906 = i_hlock7 & ~n16905;
  assign n16907 = controllable_hgrant6 & ~n8805;
  assign n16908 = controllable_hmaster2 & ~n16763;
  assign n16909 = controllable_hmaster2 & ~n16908;
  assign n16910 = controllable_hmaster1 & ~n16909;
  assign n16911 = controllable_hmaster1 & ~n16910;
  assign n16912 = ~controllable_hgrant6 & ~n16911;
  assign n16913 = ~n16907 & ~n16912;
  assign n16914 = controllable_hmaster0 & ~n16913;
  assign n16915 = controllable_hmaster0 & ~n16914;
  assign n16916 = ~controllable_hmaster3 & ~n16915;
  assign n16917 = ~controllable_hmaster3 & ~n16916;
  assign n16918 = ~i_hlock7 & ~n16917;
  assign n16919 = ~n16906 & ~n16918;
  assign n16920 = i_hbusreq7 & ~n16919;
  assign n16921 = i_hbusreq8 & ~n16903;
  assign n16922 = controllable_hgrant6 & ~n8820;
  assign n16923 = i_hbusreq6 & ~n16899;
  assign n16924 = controllable_hmaster2 & ~n16836;
  assign n16925 = controllable_hmaster2 & ~n16924;
  assign n16926 = controllable_hmaster1 & ~n16925;
  assign n16927 = controllable_hmaster1 & ~n16926;
  assign n16928 = ~i_hbusreq6 & ~n16927;
  assign n16929 = ~n16923 & ~n16928;
  assign n16930 = ~controllable_hgrant6 & ~n16929;
  assign n16931 = ~n16922 & ~n16930;
  assign n16932 = controllable_hmaster0 & ~n16931;
  assign n16933 = controllable_hmaster0 & ~n16932;
  assign n16934 = ~i_hbusreq8 & ~n16933;
  assign n16935 = ~n16921 & ~n16934;
  assign n16936 = ~controllable_hmaster3 & ~n16935;
  assign n16937 = ~controllable_hmaster3 & ~n16936;
  assign n16938 = i_hlock7 & ~n16937;
  assign n16939 = i_hbusreq8 & ~n16915;
  assign n16940 = controllable_hgrant6 & ~n8835;
  assign n16941 = i_hbusreq6 & ~n16911;
  assign n16942 = controllable_hmaster2 & ~n16873;
  assign n16943 = controllable_hmaster2 & ~n16942;
  assign n16944 = controllable_hmaster1 & ~n16943;
  assign n16945 = controllable_hmaster1 & ~n16944;
  assign n16946 = ~i_hbusreq6 & ~n16945;
  assign n16947 = ~n16941 & ~n16946;
  assign n16948 = ~controllable_hgrant6 & ~n16947;
  assign n16949 = ~n16940 & ~n16948;
  assign n16950 = controllable_hmaster0 & ~n16949;
  assign n16951 = controllable_hmaster0 & ~n16950;
  assign n16952 = ~i_hbusreq8 & ~n16951;
  assign n16953 = ~n16939 & ~n16952;
  assign n16954 = ~controllable_hmaster3 & ~n16953;
  assign n16955 = ~controllable_hmaster3 & ~n16954;
  assign n16956 = ~i_hlock7 & ~n16955;
  assign n16957 = ~n16938 & ~n16956;
  assign n16958 = ~i_hbusreq7 & ~n16957;
  assign n16959 = ~n16920 & ~n16958;
  assign n16960 = ~n8214 & ~n16959;
  assign n16961 = controllable_hgrant6 & ~n8849;
  assign n16962 = i_hlock6 & ~n16899;
  assign n16963 = ~i_hlock6 & ~n16911;
  assign n16964 = ~n16962 & ~n16963;
  assign n16965 = ~controllable_hgrant6 & ~n16964;
  assign n16966 = ~n16961 & ~n16965;
  assign n16967 = ~controllable_hmaster0 & ~n16966;
  assign n16968 = ~controllable_hmaster0 & ~n16967;
  assign n16969 = ~controllable_hmaster3 & ~n16968;
  assign n16970 = ~controllable_hmaster3 & ~n16969;
  assign n16971 = i_hbusreq7 & ~n16970;
  assign n16972 = i_hbusreq8 & ~n16968;
  assign n16973 = controllable_hgrant6 & ~n8861;
  assign n16974 = i_hbusreq6 & ~n16964;
  assign n16975 = i_hlock6 & ~n16927;
  assign n16976 = ~i_hlock6 & ~n16945;
  assign n16977 = ~n16975 & ~n16976;
  assign n16978 = ~i_hbusreq6 & ~n16977;
  assign n16979 = ~n16974 & ~n16978;
  assign n16980 = ~controllable_hgrant6 & ~n16979;
  assign n16981 = ~n16973 & ~n16980;
  assign n16982 = ~controllable_hmaster0 & ~n16981;
  assign n16983 = ~controllable_hmaster0 & ~n16982;
  assign n16984 = ~i_hbusreq8 & ~n16983;
  assign n16985 = ~n16972 & ~n16984;
  assign n16986 = ~controllable_hmaster3 & ~n16985;
  assign n16987 = ~controllable_hmaster3 & ~n16986;
  assign n16988 = ~i_hbusreq7 & ~n16987;
  assign n16989 = ~n16971 & ~n16988;
  assign n16990 = n8214 & ~n16989;
  assign n16991 = ~n16960 & ~n16990;
  assign n16992 = n8202 & ~n16991;
  assign n16993 = ~n16894 & ~n16992;
  assign n16994 = n7920 & ~n16993;
  assign n16995 = ~n16347 & ~n16994;
  assign n16996 = n7728 & ~n16995;
  assign n16997 = ~n7920 & ~n16296;
  assign n16998 = i_hready & ~controllable_hgrant2;
  assign n16999 = ~n7814 & ~n16998;
  assign n17000 = ~n7733 & ~n16999;
  assign n17001 = ~n7733 & ~n17000;
  assign n17002 = ~controllable_hgrant1 & ~n17001;
  assign n17003 = ~n7813 & ~n17002;
  assign n17004 = ~controllable_hgrant3 & ~n17003;
  assign n17005 = ~n7812 & ~n17004;
  assign n17006 = ~controllable_hgrant4 & ~n17005;
  assign n17007 = ~n7811 & ~n17006;
  assign n17008 = ~controllable_hgrant5 & ~n17007;
  assign n17009 = ~n7810 & ~n17008;
  assign n17010 = controllable_hmaster1 & ~n17009;
  assign n17011 = controllable_hmaster2 & ~n17009;
  assign n17012 = ~n16372 & ~n17011;
  assign n17013 = ~controllable_hmaster1 & ~n17012;
  assign n17014 = ~n17010 & ~n17013;
  assign n17015 = ~controllable_hgrant6 & ~n17014;
  assign n17016 = ~n12977 & ~n17015;
  assign n17017 = controllable_hmaster0 & ~n17016;
  assign n17018 = controllable_hmaster2 & ~n17011;
  assign n17019 = ~controllable_hmaster1 & ~n17018;
  assign n17020 = ~n17010 & ~n17019;
  assign n17021 = ~controllable_hgrant6 & ~n17020;
  assign n17022 = ~n7809 & ~n17021;
  assign n17023 = ~controllable_hmaster0 & ~n17022;
  assign n17024 = ~n17017 & ~n17023;
  assign n17025 = controllable_hmaster3 & ~n17024;
  assign n17026 = controllable_hmaster3 & ~n17025;
  assign n17027 = i_hbusreq7 & ~n17026;
  assign n17028 = i_hbusreq8 & ~n17024;
  assign n17029 = i_hbusreq6 & ~n17014;
  assign n17030 = i_hbusreq5 & ~n17007;
  assign n17031 = i_hbusreq4 & ~n17005;
  assign n17032 = i_hbusreq9 & ~n17005;
  assign n17033 = i_hbusreq3 & ~n17003;
  assign n17034 = i_hbusreq1 & ~n17001;
  assign n17035 = ~i_hbusreq0 & ~n7971;
  assign n17036 = ~n8106 & ~n17035;
  assign n17037 = ~i_hbusreq2 & ~n17036;
  assign n17038 = ~n8105 & ~n17037;
  assign n17039 = ~controllable_hgrant2 & ~n17038;
  assign n17040 = ~n7855 & ~n17039;
  assign n17041 = ~n7733 & ~n17040;
  assign n17042 = ~n7733 & ~n17041;
  assign n17043 = ~i_hbusreq1 & ~n17042;
  assign n17044 = ~n17034 & ~n17043;
  assign n17045 = ~controllable_hgrant1 & ~n17044;
  assign n17046 = ~n7853 & ~n17045;
  assign n17047 = ~i_hbusreq3 & ~n17046;
  assign n17048 = ~n17033 & ~n17047;
  assign n17049 = ~controllable_hgrant3 & ~n17048;
  assign n17050 = ~n7851 & ~n17049;
  assign n17051 = ~i_hbusreq9 & ~n17050;
  assign n17052 = ~n17032 & ~n17051;
  assign n17053 = ~i_hbusreq4 & ~n17052;
  assign n17054 = ~n17031 & ~n17053;
  assign n17055 = ~controllable_hgrant4 & ~n17054;
  assign n17056 = ~n7848 & ~n17055;
  assign n17057 = ~i_hbusreq5 & ~n17056;
  assign n17058 = ~n17030 & ~n17057;
  assign n17059 = ~controllable_hgrant5 & ~n17058;
  assign n17060 = ~n7846 & ~n17059;
  assign n17061 = controllable_hmaster1 & ~n17060;
  assign n17062 = controllable_hmaster2 & ~n17060;
  assign n17063 = ~n16452 & ~n17062;
  assign n17064 = ~controllable_hmaster1 & ~n17063;
  assign n17065 = ~n17061 & ~n17064;
  assign n17066 = ~i_hbusreq6 & ~n17065;
  assign n17067 = ~n17029 & ~n17066;
  assign n17068 = ~controllable_hgrant6 & ~n17067;
  assign n17069 = ~n12989 & ~n17068;
  assign n17070 = controllable_hmaster0 & ~n17069;
  assign n17071 = i_hbusreq6 & ~n17020;
  assign n17072 = controllable_hmaster2 & ~n17062;
  assign n17073 = ~controllable_hmaster1 & ~n17072;
  assign n17074 = ~n17061 & ~n17073;
  assign n17075 = ~i_hbusreq6 & ~n17074;
  assign n17076 = ~n17071 & ~n17075;
  assign n17077 = ~controllable_hgrant6 & ~n17076;
  assign n17078 = ~n7844 & ~n17077;
  assign n17079 = ~controllable_hmaster0 & ~n17078;
  assign n17080 = ~n17070 & ~n17079;
  assign n17081 = ~i_hbusreq8 & ~n17080;
  assign n17082 = ~n17028 & ~n17081;
  assign n17083 = controllable_hmaster3 & ~n17082;
  assign n17084 = controllable_hmaster3 & ~n17083;
  assign n17085 = ~i_hbusreq7 & ~n17084;
  assign n17086 = ~n17027 & ~n17085;
  assign n17087 = ~n7924 & ~n17086;
  assign n17088 = ~n7928 & ~n17001;
  assign n17089 = i_hready & controllable_locked;
  assign n17090 = ~controllable_hgrant2 & n17089;
  assign n17091 = ~n7814 & ~n17090;
  assign n17092 = ~n7733 & ~n17091;
  assign n17093 = ~n16474 & ~n17092;
  assign n17094 = n7928 & ~n17093;
  assign n17095 = ~n17088 & ~n17094;
  assign n17096 = ~controllable_hgrant1 & ~n17095;
  assign n17097 = ~n7813 & ~n17096;
  assign n17098 = ~controllable_hgrant3 & ~n17097;
  assign n17099 = ~n7812 & ~n17098;
  assign n17100 = i_hlock9 & ~n17099;
  assign n17101 = ~n16488 & ~n17092;
  assign n17102 = n7928 & ~n17101;
  assign n17103 = ~n17088 & ~n17102;
  assign n17104 = ~controllable_hgrant1 & ~n17103;
  assign n17105 = ~n7813 & ~n17104;
  assign n17106 = ~controllable_hgrant3 & ~n17105;
  assign n17107 = ~n7812 & ~n17106;
  assign n17108 = ~i_hlock9 & ~n17107;
  assign n17109 = ~n17100 & ~n17108;
  assign n17110 = ~controllable_hgrant4 & ~n17109;
  assign n17111 = ~n7811 & ~n17110;
  assign n17112 = ~controllable_hgrant5 & ~n17111;
  assign n17113 = ~n7810 & ~n17112;
  assign n17114 = controllable_hmaster1 & ~n17113;
  assign n17115 = controllable_hmaster2 & ~n17113;
  assign n17116 = ~n16536 & ~n17115;
  assign n17117 = ~controllable_hmaster1 & ~n17116;
  assign n17118 = ~n17114 & ~n17117;
  assign n17119 = ~controllable_hgrant6 & ~n17118;
  assign n17120 = ~n12977 & ~n17119;
  assign n17121 = controllable_hmaster0 & ~n17120;
  assign n17122 = ~controllable_hmaster2 & ~n16501;
  assign n17123 = ~n17115 & ~n17122;
  assign n17124 = ~controllable_hmaster1 & ~n17123;
  assign n17125 = ~n17114 & ~n17124;
  assign n17126 = ~controllable_hgrant6 & ~n17125;
  assign n17127 = ~n7809 & ~n17126;
  assign n17128 = ~controllable_hmaster0 & ~n17127;
  assign n17129 = ~n17121 & ~n17128;
  assign n17130 = controllable_hmaster3 & ~n17129;
  assign n17131 = ~n16548 & ~n17130;
  assign n17132 = i_hbusreq7 & ~n17131;
  assign n17133 = i_hbusreq8 & ~n17129;
  assign n17134 = i_hbusreq6 & ~n17118;
  assign n17135 = i_hbusreq5 & ~n17111;
  assign n17136 = i_hbusreq4 & ~n17109;
  assign n17137 = i_hbusreq9 & ~n17109;
  assign n17138 = i_hbusreq3 & ~n17097;
  assign n17139 = i_hbusreq1 & ~n17095;
  assign n17140 = ~n7928 & ~n17042;
  assign n17141 = i_hbusreq2 & n17089;
  assign n17142 = i_hbusreq0 & n17089;
  assign n17143 = controllable_locked & ~n7971;
  assign n17144 = ~controllable_locked & ~controllable_ndecide;
  assign n17145 = ~n17143 & ~n17144;
  assign n17146 = i_hlock0 & ~n17145;
  assign n17147 = ~controllable_locked & n7735;
  assign n17148 = ~n17143 & ~n17147;
  assign n17149 = ~i_hlock0 & ~n17148;
  assign n17150 = ~n17146 & ~n17149;
  assign n17151 = ~i_hbusreq0 & ~n17150;
  assign n17152 = ~n17142 & ~n17151;
  assign n17153 = ~i_hbusreq2 & ~n17152;
  assign n17154 = ~n17141 & ~n17153;
  assign n17155 = ~controllable_hgrant2 & ~n17154;
  assign n17156 = ~n7855 & ~n17155;
  assign n17157 = ~n7733 & ~n17156;
  assign n17158 = ~n16578 & ~n17157;
  assign n17159 = n7928 & ~n17158;
  assign n17160 = ~n17140 & ~n17159;
  assign n17161 = ~i_hbusreq1 & ~n17160;
  assign n17162 = ~n17139 & ~n17161;
  assign n17163 = ~controllable_hgrant1 & ~n17162;
  assign n17164 = ~n7853 & ~n17163;
  assign n17165 = ~i_hbusreq3 & ~n17164;
  assign n17166 = ~n17138 & ~n17165;
  assign n17167 = ~controllable_hgrant3 & ~n17166;
  assign n17168 = ~n7851 & ~n17167;
  assign n17169 = i_hlock9 & ~n17168;
  assign n17170 = i_hbusreq3 & ~n17105;
  assign n17171 = i_hbusreq1 & ~n17103;
  assign n17172 = ~n16488 & ~n17157;
  assign n17173 = n7928 & ~n17172;
  assign n17174 = ~n17140 & ~n17173;
  assign n17175 = ~i_hbusreq1 & ~n17174;
  assign n17176 = ~n17171 & ~n17175;
  assign n17177 = ~controllable_hgrant1 & ~n17176;
  assign n17178 = ~n7853 & ~n17177;
  assign n17179 = ~i_hbusreq3 & ~n17178;
  assign n17180 = ~n17170 & ~n17179;
  assign n17181 = ~controllable_hgrant3 & ~n17180;
  assign n17182 = ~n7851 & ~n17181;
  assign n17183 = ~i_hlock9 & ~n17182;
  assign n17184 = ~n17169 & ~n17183;
  assign n17185 = ~i_hbusreq9 & ~n17184;
  assign n17186 = ~n17137 & ~n17185;
  assign n17187 = ~i_hbusreq4 & ~n17186;
  assign n17188 = ~n17136 & ~n17187;
  assign n17189 = ~controllable_hgrant4 & ~n17188;
  assign n17190 = ~n7848 & ~n17189;
  assign n17191 = ~i_hbusreq5 & ~n17190;
  assign n17192 = ~n17135 & ~n17191;
  assign n17193 = ~controllable_hgrant5 & ~n17192;
  assign n17194 = ~n7846 & ~n17193;
  assign n17195 = controllable_hmaster1 & ~n17194;
  assign n17196 = controllable_hmaster2 & ~n17194;
  assign n17197 = ~n16693 & ~n17196;
  assign n17198 = ~controllable_hmaster1 & ~n17197;
  assign n17199 = ~n17195 & ~n17198;
  assign n17200 = ~i_hbusreq6 & ~n17199;
  assign n17201 = ~n17134 & ~n17200;
  assign n17202 = ~controllable_hgrant6 & ~n17201;
  assign n17203 = ~n12989 & ~n17202;
  assign n17204 = controllable_hmaster0 & ~n17203;
  assign n17205 = i_hbusreq6 & ~n17125;
  assign n17206 = ~controllable_hmaster2 & ~n16615;
  assign n17207 = ~n17196 & ~n17206;
  assign n17208 = ~controllable_hmaster1 & ~n17207;
  assign n17209 = ~n17195 & ~n17208;
  assign n17210 = ~i_hbusreq6 & ~n17209;
  assign n17211 = ~n17205 & ~n17210;
  assign n17212 = ~controllable_hgrant6 & ~n17211;
  assign n17213 = ~n7844 & ~n17212;
  assign n17214 = ~controllable_hmaster0 & ~n17213;
  assign n17215 = ~n17204 & ~n17214;
  assign n17216 = ~i_hbusreq8 & ~n17215;
  assign n17217 = ~n17133 & ~n17216;
  assign n17218 = controllable_hmaster3 & ~n17217;
  assign n17219 = ~n16715 & ~n17218;
  assign n17220 = ~i_hbusreq7 & ~n17219;
  assign n17221 = ~n17132 & ~n17220;
  assign n17222 = n7924 & ~n17221;
  assign n17223 = ~n17087 & ~n17222;
  assign n17224 = ~n8214 & ~n17223;
  assign n17225 = controllable_hgrant6 & ~n8907;
  assign n17226 = ~n7739 & ~n16745;
  assign n17227 = ~controllable_hmaster1 & ~n17226;
  assign n17228 = ~n7738 & ~n17227;
  assign n17229 = ~controllable_hgrant6 & ~n17228;
  assign n17230 = ~n17225 & ~n17229;
  assign n17231 = ~controllable_hmaster0 & ~n17230;
  assign n17232 = ~n8904 & ~n17231;
  assign n17233 = i_hlock8 & ~n17232;
  assign n17234 = controllable_hgrant6 & ~n8913;
  assign n17235 = ~n7739 & ~n16764;
  assign n17236 = ~controllable_hmaster1 & ~n17235;
  assign n17237 = ~n7738 & ~n17236;
  assign n17238 = ~controllable_hgrant6 & ~n17237;
  assign n17239 = ~n17234 & ~n17238;
  assign n17240 = ~controllable_hmaster0 & ~n17239;
  assign n17241 = ~n8904 & ~n17240;
  assign n17242 = ~i_hlock8 & ~n17241;
  assign n17243 = ~n17233 & ~n17242;
  assign n17244 = controllable_hmaster3 & ~n17243;
  assign n17245 = controllable_hmaster3 & ~n17244;
  assign n17246 = i_hbusreq7 & ~n17245;
  assign n17247 = i_hbusreq8 & ~n17243;
  assign n17248 = controllable_hgrant6 & ~n8928;
  assign n17249 = i_hbusreq6 & ~n17228;
  assign n17250 = ~n7771 & ~n16837;
  assign n17251 = ~controllable_hmaster1 & ~n17250;
  assign n17252 = ~n7770 & ~n17251;
  assign n17253 = ~i_hbusreq6 & ~n17252;
  assign n17254 = ~n17249 & ~n17253;
  assign n17255 = ~controllable_hgrant6 & ~n17254;
  assign n17256 = ~n17248 & ~n17255;
  assign n17257 = ~controllable_hmaster0 & ~n17256;
  assign n17258 = ~n8922 & ~n17257;
  assign n17259 = i_hlock8 & ~n17258;
  assign n17260 = controllable_hgrant6 & ~n8937;
  assign n17261 = i_hbusreq6 & ~n17237;
  assign n17262 = ~n7771 & ~n16874;
  assign n17263 = ~controllable_hmaster1 & ~n17262;
  assign n17264 = ~n7770 & ~n17263;
  assign n17265 = ~i_hbusreq6 & ~n17264;
  assign n17266 = ~n17261 & ~n17265;
  assign n17267 = ~controllable_hgrant6 & ~n17266;
  assign n17268 = ~n17260 & ~n17267;
  assign n17269 = ~controllable_hmaster0 & ~n17268;
  assign n17270 = ~n8922 & ~n17269;
  assign n17271 = ~i_hlock8 & ~n17270;
  assign n17272 = ~n17259 & ~n17271;
  assign n17273 = ~i_hbusreq8 & ~n17272;
  assign n17274 = ~n17247 & ~n17273;
  assign n17275 = controllable_hmaster3 & ~n17274;
  assign n17276 = controllable_hmaster3 & ~n17275;
  assign n17277 = ~i_hbusreq7 & ~n17276;
  assign n17278 = ~n17246 & ~n17277;
  assign n17279 = n8214 & ~n17278;
  assign n17280 = ~n17224 & ~n17279;
  assign n17281 = ~n8202 & ~n17280;
  assign n17282 = ~n7743 & ~n16904;
  assign n17283 = i_hlock7 & ~n17282;
  assign n17284 = ~n7743 & ~n16916;
  assign n17285 = ~i_hlock7 & ~n17284;
  assign n17286 = ~n17283 & ~n17285;
  assign n17287 = i_hbusreq7 & ~n17286;
  assign n17288 = ~n7779 & ~n16936;
  assign n17289 = i_hlock7 & ~n17288;
  assign n17290 = ~n7779 & ~n16954;
  assign n17291 = ~i_hlock7 & ~n17290;
  assign n17292 = ~n17289 & ~n17291;
  assign n17293 = ~i_hbusreq7 & ~n17292;
  assign n17294 = ~n17287 & ~n17293;
  assign n17295 = ~n8214 & ~n17294;
  assign n17296 = ~n7743 & ~n16969;
  assign n17297 = i_hbusreq7 & ~n17296;
  assign n17298 = ~n7779 & ~n16986;
  assign n17299 = ~i_hbusreq7 & ~n17298;
  assign n17300 = ~n17297 & ~n17299;
  assign n17301 = n8214 & ~n17300;
  assign n17302 = ~n17295 & ~n17301;
  assign n17303 = n8202 & ~n17302;
  assign n17304 = ~n17281 & ~n17303;
  assign n17305 = n7920 & ~n17304;
  assign n17306 = ~n16997 & ~n17305;
  assign n17307 = ~n7728 & ~n17306;
  assign n17308 = ~n16996 & ~n17307;
  assign n17309 = ~n7723 & ~n17308;
  assign n17310 = ~n7723 & ~n17309;
  assign n17311 = ~n7714 & ~n17310;
  assign n17312 = ~n7714 & ~n17311;
  assign n17313 = n7705 & ~n17312;
  assign n17314 = ~n16733 & ~n17000;
  assign n17315 = ~controllable_hgrant1 & ~n17314;
  assign n17316 = ~n13155 & ~n17315;
  assign n17317 = ~controllable_hgrant3 & ~n17316;
  assign n17318 = ~n13154 & ~n17317;
  assign n17319 = ~controllable_hgrant4 & ~n17318;
  assign n17320 = ~n13153 & ~n17319;
  assign n17321 = ~controllable_hgrant5 & ~n17320;
  assign n17322 = ~n13152 & ~n17321;
  assign n17323 = controllable_hmaster1 & ~n17322;
  assign n17324 = controllable_hmaster2 & ~n17322;
  assign n17325 = ~n16372 & ~n17324;
  assign n17326 = ~controllable_hmaster1 & ~n17325;
  assign n17327 = ~n17323 & ~n17326;
  assign n17328 = ~controllable_hgrant6 & ~n17327;
  assign n17329 = ~n13122 & ~n17328;
  assign n17330 = controllable_hmaster0 & ~n17329;
  assign n17331 = n7928 & ~n16735;
  assign n17332 = ~controllable_hgrant1 & ~n17331;
  assign n17333 = ~n13179 & ~n17332;
  assign n17334 = ~controllable_hgrant3 & ~n17333;
  assign n17335 = ~n13178 & ~n17334;
  assign n17336 = ~controllable_hgrant4 & ~n17335;
  assign n17337 = ~n13177 & ~n17336;
  assign n17338 = ~controllable_hgrant5 & ~n17337;
  assign n17339 = ~n13176 & ~n17338;
  assign n17340 = ~controllable_hmaster2 & ~n17339;
  assign n17341 = ~n17324 & ~n17340;
  assign n17342 = ~controllable_hmaster1 & ~n17341;
  assign n17343 = ~n17323 & ~n17342;
  assign n17344 = ~controllable_hgrant6 & ~n17343;
  assign n17345 = ~n13175 & ~n17344;
  assign n17346 = ~controllable_hmaster0 & ~n17345;
  assign n17347 = ~n17330 & ~n17346;
  assign n17348 = controllable_hmaster3 & ~n17347;
  assign n17349 = ~controllable_hgrant6 & ~n17339;
  assign n17350 = ~n13198 & ~n17349;
  assign n17351 = ~controllable_hmaster3 & ~n17350;
  assign n17352 = ~n17348 & ~n17351;
  assign n17353 = i_hbusreq7 & ~n17352;
  assign n17354 = i_hbusreq8 & ~n17347;
  assign n17355 = i_hbusreq6 & ~n17327;
  assign n17356 = i_hbusreq5 & ~n17320;
  assign n17357 = i_hbusreq4 & ~n17318;
  assign n17358 = i_hbusreq9 & ~n17318;
  assign n17359 = i_hbusreq3 & ~n17316;
  assign n17360 = i_hbusreq1 & ~n17314;
  assign n17361 = ~controllable_hmastlock & ~n7971;
  assign n17362 = ~controllable_hmastlock & ~n17361;
  assign n17363 = controllable_locked & ~n17362;
  assign n17364 = ~n16787 & ~n17363;
  assign n17365 = ~i_hbusreq0 & ~n17364;
  assign n17366 = ~n16800 & ~n17365;
  assign n17367 = ~i_hbusreq2 & ~n17366;
  assign n17368 = ~n16799 & ~n17367;
  assign n17369 = ~controllable_hgrant2 & ~n17368;
  assign n17370 = ~n7855 & ~n17369;
  assign n17371 = n7733 & ~n17370;
  assign n17372 = ~n17041 & ~n17371;
  assign n17373 = ~i_hbusreq1 & ~n17372;
  assign n17374 = ~n17360 & ~n17373;
  assign n17375 = ~controllable_hgrant1 & ~n17374;
  assign n17376 = ~n13213 & ~n17375;
  assign n17377 = ~i_hbusreq3 & ~n17376;
  assign n17378 = ~n17359 & ~n17377;
  assign n17379 = ~controllable_hgrant3 & ~n17378;
  assign n17380 = ~n13211 & ~n17379;
  assign n17381 = ~i_hbusreq9 & ~n17380;
  assign n17382 = ~n17358 & ~n17381;
  assign n17383 = ~i_hbusreq4 & ~n17382;
  assign n17384 = ~n17357 & ~n17383;
  assign n17385 = ~controllable_hgrant4 & ~n17384;
  assign n17386 = ~n13208 & ~n17385;
  assign n17387 = ~i_hbusreq5 & ~n17386;
  assign n17388 = ~n17356 & ~n17387;
  assign n17389 = ~controllable_hgrant5 & ~n17388;
  assign n17390 = ~n13206 & ~n17389;
  assign n17391 = controllable_hmaster1 & ~n17390;
  assign n17392 = controllable_hmaster2 & ~n17390;
  assign n17393 = ~n16452 & ~n17392;
  assign n17394 = ~controllable_hmaster1 & ~n17393;
  assign n17395 = ~n17391 & ~n17394;
  assign n17396 = ~i_hbusreq6 & ~n17395;
  assign n17397 = ~n17355 & ~n17396;
  assign n17398 = ~controllable_hgrant6 & ~n17397;
  assign n17399 = ~n13134 & ~n17398;
  assign n17400 = controllable_hmaster0 & ~n17399;
  assign n17401 = i_hbusreq6 & ~n17343;
  assign n17402 = i_hbusreq5 & ~n17337;
  assign n17403 = i_hbusreq4 & ~n17335;
  assign n17404 = i_hbusreq9 & ~n17335;
  assign n17405 = i_hbusreq3 & ~n17333;
  assign n17406 = i_hbusreq1 & ~n17331;
  assign n17407 = ~i_hbusreq0 & ~n16788;
  assign n17408 = ~n16786 & ~n17407;
  assign n17409 = ~i_hbusreq2 & ~n17408;
  assign n17410 = ~n16785 & ~n17409;
  assign n17411 = ~controllable_hgrant2 & ~n17410;
  assign n17412 = ~n7855 & ~n17411;
  assign n17413 = ~n7733 & ~n17412;
  assign n17414 = ~n17371 & ~n17413;
  assign n17415 = n7928 & ~n17414;
  assign n17416 = n7928 & ~n17415;
  assign n17417 = ~i_hbusreq1 & ~n17416;
  assign n17418 = ~n17406 & ~n17417;
  assign n17419 = ~controllable_hgrant1 & ~n17418;
  assign n17420 = ~n13263 & ~n17419;
  assign n17421 = ~i_hbusreq3 & ~n17420;
  assign n17422 = ~n17405 & ~n17421;
  assign n17423 = ~controllable_hgrant3 & ~n17422;
  assign n17424 = ~n13261 & ~n17423;
  assign n17425 = ~i_hbusreq9 & ~n17424;
  assign n17426 = ~n17404 & ~n17425;
  assign n17427 = ~i_hbusreq4 & ~n17426;
  assign n17428 = ~n17403 & ~n17427;
  assign n17429 = ~controllable_hgrant4 & ~n17428;
  assign n17430 = ~n13258 & ~n17429;
  assign n17431 = ~i_hbusreq5 & ~n17430;
  assign n17432 = ~n17402 & ~n17431;
  assign n17433 = ~controllable_hgrant5 & ~n17432;
  assign n17434 = ~n13256 & ~n17433;
  assign n17435 = ~controllable_hmaster2 & ~n17434;
  assign n17436 = ~n17392 & ~n17435;
  assign n17437 = ~controllable_hmaster1 & ~n17436;
  assign n17438 = ~n17391 & ~n17437;
  assign n17439 = ~i_hbusreq6 & ~n17438;
  assign n17440 = ~n17401 & ~n17439;
  assign n17441 = ~controllable_hgrant6 & ~n17440;
  assign n17442 = ~n13254 & ~n17441;
  assign n17443 = ~controllable_hmaster0 & ~n17442;
  assign n17444 = ~n17400 & ~n17443;
  assign n17445 = ~i_hbusreq8 & ~n17444;
  assign n17446 = ~n17354 & ~n17445;
  assign n17447 = controllable_hmaster3 & ~n17446;
  assign n17448 = i_hbusreq8 & ~n17350;
  assign n17449 = i_hbusreq6 & ~n17339;
  assign n17450 = ~i_hbusreq6 & ~n17434;
  assign n17451 = ~n17449 & ~n17450;
  assign n17452 = ~controllable_hgrant6 & ~n17451;
  assign n17453 = ~n13298 & ~n17452;
  assign n17454 = ~i_hbusreq8 & ~n17453;
  assign n17455 = ~n17448 & ~n17454;
  assign n17456 = ~controllable_hmaster3 & ~n17455;
  assign n17457 = ~n17447 & ~n17456;
  assign n17458 = ~i_hbusreq7 & ~n17457;
  assign n17459 = ~n17353 & ~n17458;
  assign n17460 = ~n7924 & ~n17459;
  assign n17461 = ~n7928 & ~n17314;
  assign n17462 = controllable_hmastlock & ~n7975;
  assign n17463 = controllable_locked & ~n17462;
  assign n17464 = controllable_locked & ~n17463;
  assign n17465 = ~controllable_hgrant2 & n17464;
  assign n17466 = ~n7814 & ~n17465;
  assign n17467 = n7733 & ~n17466;
  assign n17468 = ~n17092 & ~n17467;
  assign n17469 = n7928 & ~n17468;
  assign n17470 = ~n17461 & ~n17469;
  assign n17471 = ~controllable_hgrant1 & ~n17470;
  assign n17472 = ~n13155 & ~n17471;
  assign n17473 = ~controllable_hgrant3 & ~n17472;
  assign n17474 = ~n13154 & ~n17473;
  assign n17475 = i_hlock9 & ~n17474;
  assign n17476 = ~n7970 & ~n12781;
  assign n17477 = controllable_hmastlock & ~n17476;
  assign n17478 = ~n14241 & ~n17477;
  assign n17479 = controllable_locked & ~n17478;
  assign n17480 = controllable_locked & ~n17479;
  assign n17481 = ~controllable_hgrant2 & n17480;
  assign n17482 = ~n7814 & ~n17481;
  assign n17483 = n7733 & ~n17482;
  assign n17484 = ~n17092 & ~n17483;
  assign n17485 = n7928 & ~n17484;
  assign n17486 = ~n17461 & ~n17485;
  assign n17487 = ~controllable_hgrant1 & ~n17486;
  assign n17488 = ~n13155 & ~n17487;
  assign n17489 = ~controllable_hgrant3 & ~n17488;
  assign n17490 = ~n13154 & ~n17489;
  assign n17491 = ~i_hlock9 & ~n17490;
  assign n17492 = ~n17475 & ~n17491;
  assign n17493 = ~controllable_hgrant4 & ~n17492;
  assign n17494 = ~n13153 & ~n17493;
  assign n17495 = ~controllable_hgrant5 & ~n17494;
  assign n17496 = ~n13152 & ~n17495;
  assign n17497 = controllable_hmaster1 & ~n17496;
  assign n17498 = controllable_hmaster2 & ~n17496;
  assign n17499 = ~n16536 & ~n17498;
  assign n17500 = ~controllable_hmaster1 & ~n17499;
  assign n17501 = ~n17497 & ~n17500;
  assign n17502 = ~controllable_hgrant6 & ~n17501;
  assign n17503 = ~n13122 & ~n17502;
  assign n17504 = controllable_hmaster0 & ~n17503;
  assign n17505 = ~controllable_hgrant2 & n13008;
  assign n17506 = ~n7814 & ~n17505;
  assign n17507 = ~n7733 & ~n17506;
  assign n17508 = ~n17467 & ~n17507;
  assign n17509 = n7928 & ~n17508;
  assign n17510 = n7928 & ~n17509;
  assign n17511 = ~controllable_hgrant1 & ~n17510;
  assign n17512 = ~n13179 & ~n17511;
  assign n17513 = ~controllable_hgrant3 & ~n17512;
  assign n17514 = ~n13178 & ~n17513;
  assign n17515 = i_hlock9 & ~n17514;
  assign n17516 = ~n17483 & ~n17507;
  assign n17517 = n7928 & ~n17516;
  assign n17518 = n7928 & ~n17517;
  assign n17519 = ~controllable_hgrant1 & ~n17518;
  assign n17520 = ~n13179 & ~n17519;
  assign n17521 = ~controllable_hgrant3 & ~n17520;
  assign n17522 = ~n13178 & ~n17521;
  assign n17523 = ~i_hlock9 & ~n17522;
  assign n17524 = ~n17515 & ~n17523;
  assign n17525 = ~controllable_hgrant4 & ~n17524;
  assign n17526 = ~n13177 & ~n17525;
  assign n17527 = ~controllable_hgrant5 & ~n17526;
  assign n17528 = ~n13176 & ~n17527;
  assign n17529 = ~controllable_hmaster2 & ~n17528;
  assign n17530 = ~n17498 & ~n17529;
  assign n17531 = ~controllable_hmaster1 & ~n17530;
  assign n17532 = ~n17497 & ~n17531;
  assign n17533 = ~controllable_hgrant6 & ~n17532;
  assign n17534 = ~n13175 & ~n17533;
  assign n17535 = ~controllable_hmaster0 & ~n17534;
  assign n17536 = ~n17504 & ~n17535;
  assign n17537 = controllable_hmaster3 & ~n17536;
  assign n17538 = ~controllable_hgrant6 & ~n17528;
  assign n17539 = ~n13198 & ~n17538;
  assign n17540 = ~controllable_hmaster3 & ~n17539;
  assign n17541 = ~n17537 & ~n17540;
  assign n17542 = i_hbusreq7 & ~n17541;
  assign n17543 = i_hbusreq8 & ~n17536;
  assign n17544 = i_hbusreq6 & ~n17501;
  assign n17545 = i_hbusreq5 & ~n17494;
  assign n17546 = i_hbusreq4 & ~n17492;
  assign n17547 = i_hbusreq9 & ~n17492;
  assign n17548 = i_hbusreq3 & ~n17472;
  assign n17549 = i_hbusreq1 & ~n17470;
  assign n17550 = ~n7928 & ~n17372;
  assign n17551 = i_hbusreq2 & ~n17464;
  assign n17552 = i_hbusreq0 & ~n17464;
  assign n17553 = controllable_hmastlock & n7970;
  assign n17554 = ~n12624 & ~n17553;
  assign n17555 = controllable_locked & ~n17554;
  assign n17556 = ~controllable_locked & ~n7735;
  assign n17557 = ~n17555 & ~n17556;
  assign n17558 = ~i_hbusreq0 & ~n17557;
  assign n17559 = ~n17552 & ~n17558;
  assign n17560 = ~i_hbusreq2 & ~n17559;
  assign n17561 = ~n17551 & ~n17560;
  assign n17562 = ~controllable_hgrant2 & n17561;
  assign n17563 = ~n7855 & ~n17562;
  assign n17564 = n7733 & ~n17563;
  assign n17565 = ~n17157 & ~n17564;
  assign n17566 = n7928 & ~n17565;
  assign n17567 = ~n17550 & ~n17566;
  assign n17568 = ~i_hbusreq1 & ~n17567;
  assign n17569 = ~n17549 & ~n17568;
  assign n17570 = ~controllable_hgrant1 & ~n17569;
  assign n17571 = ~n13213 & ~n17570;
  assign n17572 = ~i_hbusreq3 & ~n17571;
  assign n17573 = ~n17548 & ~n17572;
  assign n17574 = ~controllable_hgrant3 & ~n17573;
  assign n17575 = ~n13211 & ~n17574;
  assign n17576 = i_hlock9 & ~n17575;
  assign n17577 = i_hbusreq3 & ~n17488;
  assign n17578 = i_hbusreq1 & ~n17486;
  assign n17579 = i_hbusreq2 & ~n17480;
  assign n17580 = i_hbusreq0 & ~n17480;
  assign n17581 = ~n17558 & ~n17580;
  assign n17582 = ~i_hbusreq2 & ~n17581;
  assign n17583 = ~n17579 & ~n17582;
  assign n17584 = ~controllable_hgrant2 & n17583;
  assign n17585 = ~n7855 & ~n17584;
  assign n17586 = n7733 & ~n17585;
  assign n17587 = ~n17157 & ~n17586;
  assign n17588 = n7928 & ~n17587;
  assign n17589 = ~n17550 & ~n17588;
  assign n17590 = ~i_hbusreq1 & ~n17589;
  assign n17591 = ~n17578 & ~n17590;
  assign n17592 = ~controllable_hgrant1 & ~n17591;
  assign n17593 = ~n13213 & ~n17592;
  assign n17594 = ~i_hbusreq3 & ~n17593;
  assign n17595 = ~n17577 & ~n17594;
  assign n17596 = ~controllable_hgrant3 & ~n17595;
  assign n17597 = ~n13211 & ~n17596;
  assign n17598 = ~i_hlock9 & ~n17597;
  assign n17599 = ~n17576 & ~n17598;
  assign n17600 = ~i_hbusreq9 & ~n17599;
  assign n17601 = ~n17547 & ~n17600;
  assign n17602 = ~i_hbusreq4 & ~n17601;
  assign n17603 = ~n17546 & ~n17602;
  assign n17604 = ~controllable_hgrant4 & ~n17603;
  assign n17605 = ~n13208 & ~n17604;
  assign n17606 = ~i_hbusreq5 & ~n17605;
  assign n17607 = ~n17545 & ~n17606;
  assign n17608 = ~controllable_hgrant5 & ~n17607;
  assign n17609 = ~n13206 & ~n17608;
  assign n17610 = controllable_hmaster1 & ~n17609;
  assign n17611 = controllable_hmaster2 & ~n17609;
  assign n17612 = ~n16693 & ~n17611;
  assign n17613 = ~controllable_hmaster1 & ~n17612;
  assign n17614 = ~n17610 & ~n17613;
  assign n17615 = ~i_hbusreq6 & ~n17614;
  assign n17616 = ~n17544 & ~n17615;
  assign n17617 = ~controllable_hgrant6 & ~n17616;
  assign n17618 = ~n13134 & ~n17617;
  assign n17619 = controllable_hmaster0 & ~n17618;
  assign n17620 = i_hbusreq6 & ~n17532;
  assign n17621 = i_hbusreq5 & ~n17526;
  assign n17622 = i_hbusreq4 & ~n17524;
  assign n17623 = i_hbusreq9 & ~n17524;
  assign n17624 = i_hbusreq3 & ~n17512;
  assign n17625 = i_hbusreq1 & ~n17510;
  assign n17626 = i_hbusreq2 & n13008;
  assign n17627 = i_hbusreq0 & n13008;
  assign n17628 = ~controllable_locked & ~n17144;
  assign n17629 = i_hlock0 & ~n17628;
  assign n17630 = ~controllable_locked & ~n17147;
  assign n17631 = ~i_hlock0 & ~n17630;
  assign n17632 = ~n17629 & ~n17631;
  assign n17633 = ~i_hbusreq0 & ~n17632;
  assign n17634 = ~n17627 & ~n17633;
  assign n17635 = ~i_hbusreq2 & ~n17634;
  assign n17636 = ~n17626 & ~n17635;
  assign n17637 = ~controllable_hgrant2 & ~n17636;
  assign n17638 = ~n7855 & ~n17637;
  assign n17639 = ~n7733 & ~n17638;
  assign n17640 = ~n17564 & ~n17639;
  assign n17641 = n7928 & ~n17640;
  assign n17642 = n7928 & ~n17641;
  assign n17643 = ~i_hbusreq1 & ~n17642;
  assign n17644 = ~n17625 & ~n17643;
  assign n17645 = ~controllable_hgrant1 & ~n17644;
  assign n17646 = ~n13263 & ~n17645;
  assign n17647 = ~i_hbusreq3 & ~n17646;
  assign n17648 = ~n17624 & ~n17647;
  assign n17649 = ~controllable_hgrant3 & ~n17648;
  assign n17650 = ~n13261 & ~n17649;
  assign n17651 = i_hlock9 & ~n17650;
  assign n17652 = i_hbusreq3 & ~n17520;
  assign n17653 = i_hbusreq1 & ~n17518;
  assign n17654 = ~n17586 & ~n17639;
  assign n17655 = n7928 & ~n17654;
  assign n17656 = n7928 & ~n17655;
  assign n17657 = ~i_hbusreq1 & ~n17656;
  assign n17658 = ~n17653 & ~n17657;
  assign n17659 = ~controllable_hgrant1 & ~n17658;
  assign n17660 = ~n13263 & ~n17659;
  assign n17661 = ~i_hbusreq3 & ~n17660;
  assign n17662 = ~n17652 & ~n17661;
  assign n17663 = ~controllable_hgrant3 & ~n17662;
  assign n17664 = ~n13261 & ~n17663;
  assign n17665 = ~i_hlock9 & ~n17664;
  assign n17666 = ~n17651 & ~n17665;
  assign n17667 = ~i_hbusreq9 & ~n17666;
  assign n17668 = ~n17623 & ~n17667;
  assign n17669 = ~i_hbusreq4 & ~n17668;
  assign n17670 = ~n17622 & ~n17669;
  assign n17671 = ~controllable_hgrant4 & ~n17670;
  assign n17672 = ~n13258 & ~n17671;
  assign n17673 = ~i_hbusreq5 & ~n17672;
  assign n17674 = ~n17621 & ~n17673;
  assign n17675 = ~controllable_hgrant5 & ~n17674;
  assign n17676 = ~n13256 & ~n17675;
  assign n17677 = ~controllable_hmaster2 & ~n17676;
  assign n17678 = ~n17611 & ~n17677;
  assign n17679 = ~controllable_hmaster1 & ~n17678;
  assign n17680 = ~n17610 & ~n17679;
  assign n17681 = ~i_hbusreq6 & ~n17680;
  assign n17682 = ~n17620 & ~n17681;
  assign n17683 = ~controllable_hgrant6 & ~n17682;
  assign n17684 = ~n13254 & ~n17683;
  assign n17685 = ~controllable_hmaster0 & ~n17684;
  assign n17686 = ~n17619 & ~n17685;
  assign n17687 = ~i_hbusreq8 & ~n17686;
  assign n17688 = ~n17543 & ~n17687;
  assign n17689 = controllable_hmaster3 & ~n17688;
  assign n17690 = i_hbusreq8 & ~n17539;
  assign n17691 = i_hbusreq6 & ~n17528;
  assign n17692 = ~i_hbusreq6 & ~n17676;
  assign n17693 = ~n17691 & ~n17692;
  assign n17694 = ~controllable_hgrant6 & ~n17693;
  assign n17695 = ~n13298 & ~n17694;
  assign n17696 = ~i_hbusreq8 & ~n17695;
  assign n17697 = ~n17690 & ~n17696;
  assign n17698 = ~controllable_hmaster3 & ~n17697;
  assign n17699 = ~n17689 & ~n17698;
  assign n17700 = ~i_hbusreq7 & ~n17699;
  assign n17701 = ~n17542 & ~n17700;
  assign n17702 = n7924 & ~n17701;
  assign n17703 = ~n17460 & ~n17702;
  assign n17704 = ~n8214 & ~n17703;
  assign n17705 = ~n8358 & ~n16745;
  assign n17706 = ~controllable_hmaster1 & ~n17705;
  assign n17707 = ~n8357 & ~n17706;
  assign n17708 = ~controllable_hgrant6 & ~n17707;
  assign n17709 = ~n13406 & ~n17708;
  assign n17710 = ~controllable_hmaster0 & ~n17709;
  assign n17711 = ~n13328 & ~n17710;
  assign n17712 = i_hlock8 & ~n17711;
  assign n17713 = ~n8358 & ~n16764;
  assign n17714 = ~controllable_hmaster1 & ~n17713;
  assign n17715 = ~n8357 & ~n17714;
  assign n17716 = ~controllable_hgrant6 & ~n17715;
  assign n17717 = ~n13427 & ~n17716;
  assign n17718 = ~controllable_hmaster0 & ~n17717;
  assign n17719 = ~n13328 & ~n17718;
  assign n17720 = ~i_hlock8 & ~n17719;
  assign n17721 = ~n17712 & ~n17720;
  assign n17722 = controllable_hmaster3 & ~n17721;
  assign n17723 = ~n8995 & ~n17722;
  assign n17724 = i_hbusreq7 & ~n17723;
  assign n17725 = i_hbusreq8 & ~n17721;
  assign n17726 = i_hbusreq6 & ~n17707;
  assign n17727 = ~n8484 & ~n16837;
  assign n17728 = ~controllable_hmaster1 & ~n17727;
  assign n17729 = ~n8483 & ~n17728;
  assign n17730 = ~i_hbusreq6 & ~n17729;
  assign n17731 = ~n17726 & ~n17730;
  assign n17732 = ~controllable_hgrant6 & ~n17731;
  assign n17733 = ~n13520 & ~n17732;
  assign n17734 = ~controllable_hmaster0 & ~n17733;
  assign n17735 = ~n13377 & ~n17734;
  assign n17736 = i_hlock8 & ~n17735;
  assign n17737 = i_hbusreq6 & ~n17715;
  assign n17738 = ~n8484 & ~n16874;
  assign n17739 = ~controllable_hmaster1 & ~n17738;
  assign n17740 = ~n8483 & ~n17739;
  assign n17741 = ~i_hbusreq6 & ~n17740;
  assign n17742 = ~n17737 & ~n17741;
  assign n17743 = ~controllable_hgrant6 & ~n17742;
  assign n17744 = ~n13573 & ~n17743;
  assign n17745 = ~controllable_hmaster0 & ~n17744;
  assign n17746 = ~n13377 & ~n17745;
  assign n17747 = ~i_hlock8 & ~n17746;
  assign n17748 = ~n17736 & ~n17747;
  assign n17749 = ~i_hbusreq8 & ~n17748;
  assign n17750 = ~n17725 & ~n17749;
  assign n17751 = controllable_hmaster3 & ~n17750;
  assign n17752 = ~n9041 & ~n17751;
  assign n17753 = ~i_hbusreq7 & ~n17752;
  assign n17754 = ~n17724 & ~n17753;
  assign n17755 = ~n7924 & ~n17754;
  assign n17756 = ~controllable_locked & n7970;
  assign n17757 = ~n13008 & ~n17756;
  assign n17758 = ~controllable_hgrant2 & ~n17757;
  assign n17759 = ~n7814 & ~n17758;
  assign n17760 = ~n7733 & ~n17759;
  assign n17761 = ~n16729 & ~n17756;
  assign n17762 = ~controllable_hgrant2 & ~n17761;
  assign n17763 = ~n7814 & ~n17762;
  assign n17764 = n7733 & ~n17763;
  assign n17765 = ~n17760 & ~n17764;
  assign n17766 = n7928 & ~n17765;
  assign n17767 = ~n8221 & ~n17766;
  assign n17768 = ~controllable_hgrant1 & ~n17767;
  assign n17769 = ~n12611 & ~n17768;
  assign n17770 = ~controllable_hgrant3 & ~n17769;
  assign n17771 = ~n12610 & ~n17770;
  assign n17772 = ~controllable_hgrant4 & ~n17771;
  assign n17773 = ~n13408 & ~n17772;
  assign n17774 = ~controllable_hgrant5 & ~n17773;
  assign n17775 = ~n13407 & ~n17774;
  assign n17776 = ~controllable_hmaster2 & ~n17775;
  assign n17777 = ~n13168 & ~n17776;
  assign n17778 = ~controllable_hmaster1 & ~n17777;
  assign n17779 = ~n13167 & ~n17778;
  assign n17780 = ~controllable_hgrant6 & ~n17779;
  assign n17781 = ~n13406 & ~n17780;
  assign n17782 = ~controllable_hmaster0 & ~n17781;
  assign n17783 = ~n13405 & ~n17782;
  assign n17784 = i_hlock8 & ~n17783;
  assign n17785 = ~n8235 & ~n17766;
  assign n17786 = ~controllable_hgrant1 & ~n17785;
  assign n17787 = ~n12638 & ~n17786;
  assign n17788 = ~controllable_hgrant3 & ~n17787;
  assign n17789 = ~n12637 & ~n17788;
  assign n17790 = ~controllable_hgrant4 & ~n17789;
  assign n17791 = ~n13429 & ~n17790;
  assign n17792 = ~controllable_hgrant5 & ~n17791;
  assign n17793 = ~n13428 & ~n17792;
  assign n17794 = ~controllable_hmaster2 & ~n17793;
  assign n17795 = ~n13168 & ~n17794;
  assign n17796 = ~controllable_hmaster1 & ~n17795;
  assign n17797 = ~n13167 & ~n17796;
  assign n17798 = ~controllable_hgrant6 & ~n17797;
  assign n17799 = ~n13427 & ~n17798;
  assign n17800 = ~controllable_hmaster0 & ~n17799;
  assign n17801 = ~n13405 & ~n17800;
  assign n17802 = ~i_hlock8 & ~n17801;
  assign n17803 = ~n17784 & ~n17802;
  assign n17804 = controllable_hmaster3 & ~n17803;
  assign n17805 = ~n13201 & ~n17804;
  assign n17806 = i_hbusreq7 & ~n17805;
  assign n17807 = i_hbusreq8 & ~n17803;
  assign n17808 = i_hbusreq6 & ~n17779;
  assign n17809 = i_hbusreq5 & ~n17773;
  assign n17810 = i_hbusreq4 & ~n17771;
  assign n17811 = i_hbusreq9 & ~n17771;
  assign n17812 = i_hbusreq3 & ~n17769;
  assign n17813 = i_hbusreq1 & ~n17767;
  assign n17814 = i_hbusreq2 & ~n17757;
  assign n17815 = i_hbusreq0 & ~n17757;
  assign n17816 = ~n16792 & ~n17815;
  assign n17817 = ~i_hbusreq2 & ~n17816;
  assign n17818 = ~n17814 & ~n17817;
  assign n17819 = ~controllable_hgrant2 & ~n17818;
  assign n17820 = ~n12694 & ~n17819;
  assign n17821 = ~n7733 & ~n17820;
  assign n17822 = i_hbusreq2 & ~n17761;
  assign n17823 = i_hbusreq0 & ~n17761;
  assign n17824 = ~n16809 & ~n17823;
  assign n17825 = ~i_hbusreq2 & ~n17824;
  assign n17826 = ~n17822 & ~n17825;
  assign n17827 = ~controllable_hgrant2 & ~n17826;
  assign n17828 = ~n12706 & ~n17827;
  assign n17829 = n7733 & ~n17828;
  assign n17830 = ~n17821 & ~n17829;
  assign n17831 = n7928 & ~n17830;
  assign n17832 = ~n8265 & ~n17831;
  assign n17833 = ~i_hbusreq1 & ~n17832;
  assign n17834 = ~n17813 & ~n17833;
  assign n17835 = ~controllable_hgrant1 & ~n17834;
  assign n17836 = ~n12681 & ~n17835;
  assign n17837 = ~i_hbusreq3 & ~n17836;
  assign n17838 = ~n17812 & ~n17837;
  assign n17839 = ~controllable_hgrant3 & ~n17838;
  assign n17840 = ~n12679 & ~n17839;
  assign n17841 = ~i_hbusreq9 & ~n17840;
  assign n17842 = ~n17811 & ~n17841;
  assign n17843 = ~i_hbusreq4 & ~n17842;
  assign n17844 = ~n17810 & ~n17843;
  assign n17845 = ~controllable_hgrant4 & ~n17844;
  assign n17846 = ~n13524 & ~n17845;
  assign n17847 = ~i_hbusreq5 & ~n17846;
  assign n17848 = ~n17809 & ~n17847;
  assign n17849 = ~controllable_hgrant5 & ~n17848;
  assign n17850 = ~n13522 & ~n17849;
  assign n17851 = ~controllable_hmaster2 & ~n17850;
  assign n17852 = ~n13480 & ~n17851;
  assign n17853 = ~controllable_hmaster1 & ~n17852;
  assign n17854 = ~n13479 & ~n17853;
  assign n17855 = ~i_hbusreq6 & ~n17854;
  assign n17856 = ~n17808 & ~n17855;
  assign n17857 = ~controllable_hgrant6 & ~n17856;
  assign n17858 = ~n13520 & ~n17857;
  assign n17859 = ~controllable_hmaster0 & ~n17858;
  assign n17860 = ~n13519 & ~n17859;
  assign n17861 = i_hlock8 & ~n17860;
  assign n17862 = i_hbusreq6 & ~n17797;
  assign n17863 = i_hbusreq5 & ~n17791;
  assign n17864 = i_hbusreq4 & ~n17789;
  assign n17865 = i_hbusreq9 & ~n17789;
  assign n17866 = i_hbusreq3 & ~n17787;
  assign n17867 = i_hbusreq1 & ~n17785;
  assign n17868 = ~n8297 & ~n17831;
  assign n17869 = ~i_hbusreq1 & ~n17868;
  assign n17870 = ~n17867 & ~n17869;
  assign n17871 = ~controllable_hgrant1 & ~n17870;
  assign n17872 = ~n12730 & ~n17871;
  assign n17873 = ~i_hbusreq3 & ~n17872;
  assign n17874 = ~n17866 & ~n17873;
  assign n17875 = ~controllable_hgrant3 & ~n17874;
  assign n17876 = ~n12728 & ~n17875;
  assign n17877 = ~i_hbusreq9 & ~n17876;
  assign n17878 = ~n17865 & ~n17877;
  assign n17879 = ~i_hbusreq4 & ~n17878;
  assign n17880 = ~n17864 & ~n17879;
  assign n17881 = ~controllable_hgrant4 & ~n17880;
  assign n17882 = ~n13577 & ~n17881;
  assign n17883 = ~i_hbusreq5 & ~n17882;
  assign n17884 = ~n17863 & ~n17883;
  assign n17885 = ~controllable_hgrant5 & ~n17884;
  assign n17886 = ~n13575 & ~n17885;
  assign n17887 = ~controllable_hmaster2 & ~n17886;
  assign n17888 = ~n13480 & ~n17887;
  assign n17889 = ~controllable_hmaster1 & ~n17888;
  assign n17890 = ~n13479 & ~n17889;
  assign n17891 = ~i_hbusreq6 & ~n17890;
  assign n17892 = ~n17862 & ~n17891;
  assign n17893 = ~controllable_hgrant6 & ~n17892;
  assign n17894 = ~n13573 & ~n17893;
  assign n17895 = ~controllable_hmaster0 & ~n17894;
  assign n17896 = ~n13519 & ~n17895;
  assign n17897 = ~i_hlock8 & ~n17896;
  assign n17898 = ~n17861 & ~n17897;
  assign n17899 = ~i_hbusreq8 & ~n17898;
  assign n17900 = ~n17807 & ~n17899;
  assign n17901 = controllable_hmaster3 & ~n17900;
  assign n17902 = ~n13641 & ~n17901;
  assign n17903 = ~i_hbusreq7 & ~n17902;
  assign n17904 = ~n17806 & ~n17903;
  assign n17905 = n7924 & ~n17904;
  assign n17906 = ~n17755 & ~n17905;
  assign n17907 = n8214 & ~n17906;
  assign n17908 = ~n17704 & ~n17907;
  assign n17909 = ~n8202 & ~n17908;
  assign n17910 = ~n8988 & ~n16896;
  assign n17911 = controllable_hmaster1 & ~n17910;
  assign n17912 = ~n9096 & ~n17911;
  assign n17913 = ~controllable_hgrant6 & ~n17912;
  assign n17914 = ~n13673 & ~n17913;
  assign n17915 = controllable_hmaster0 & ~n17914;
  assign n17916 = ~n9099 & ~n17915;
  assign n17917 = ~controllable_hmaster3 & ~n17916;
  assign n17918 = ~n13651 & ~n17917;
  assign n17919 = i_hlock7 & ~n17918;
  assign n17920 = ~n8988 & ~n16908;
  assign n17921 = controllable_hmaster1 & ~n17920;
  assign n17922 = ~n9096 & ~n17921;
  assign n17923 = ~controllable_hgrant6 & ~n17922;
  assign n17924 = ~n13687 & ~n17923;
  assign n17925 = controllable_hmaster0 & ~n17924;
  assign n17926 = ~n9099 & ~n17925;
  assign n17927 = ~controllable_hmaster3 & ~n17926;
  assign n17928 = ~n13651 & ~n17927;
  assign n17929 = ~i_hlock7 & ~n17928;
  assign n17930 = ~n17919 & ~n17929;
  assign n17931 = i_hbusreq7 & ~n17930;
  assign n17932 = i_hbusreq8 & ~n17916;
  assign n17933 = i_hbusreq6 & ~n17912;
  assign n17934 = ~n9024 & ~n16924;
  assign n17935 = controllable_hmaster1 & ~n17934;
  assign n17936 = ~n9122 & ~n17935;
  assign n17937 = ~i_hbusreq6 & ~n17936;
  assign n17938 = ~n17933 & ~n17937;
  assign n17939 = ~controllable_hgrant6 & ~n17938;
  assign n17940 = ~n13716 & ~n17939;
  assign n17941 = controllable_hmaster0 & ~n17940;
  assign n17942 = ~n9127 & ~n17941;
  assign n17943 = ~i_hbusreq8 & ~n17942;
  assign n17944 = ~n17932 & ~n17943;
  assign n17945 = ~controllable_hmaster3 & ~n17944;
  assign n17946 = ~n13662 & ~n17945;
  assign n17947 = i_hlock7 & ~n17946;
  assign n17948 = i_hbusreq8 & ~n17926;
  assign n17949 = i_hbusreq6 & ~n17922;
  assign n17950 = ~n9024 & ~n16942;
  assign n17951 = controllable_hmaster1 & ~n17950;
  assign n17952 = ~n9122 & ~n17951;
  assign n17953 = ~i_hbusreq6 & ~n17952;
  assign n17954 = ~n17949 & ~n17953;
  assign n17955 = ~controllable_hgrant6 & ~n17954;
  assign n17956 = ~n13736 & ~n17955;
  assign n17957 = controllable_hmaster0 & ~n17956;
  assign n17958 = ~n9127 & ~n17957;
  assign n17959 = ~i_hbusreq8 & ~n17958;
  assign n17960 = ~n17948 & ~n17959;
  assign n17961 = ~controllable_hmaster3 & ~n17960;
  assign n17962 = ~n13662 & ~n17961;
  assign n17963 = ~i_hlock7 & ~n17962;
  assign n17964 = ~n17947 & ~n17963;
  assign n17965 = ~i_hbusreq7 & ~n17964;
  assign n17966 = ~n17931 & ~n17965;
  assign n17967 = ~n7924 & ~n17966;
  assign n17968 = controllable_hmaster2 & ~n17775;
  assign n17969 = ~n13189 & ~n17968;
  assign n17970 = controllable_hmaster1 & ~n17969;
  assign n17971 = ~n13677 & ~n17970;
  assign n17972 = ~controllable_hgrant6 & ~n17971;
  assign n17973 = ~n13673 & ~n17972;
  assign n17974 = controllable_hmaster0 & ~n17973;
  assign n17975 = ~n13682 & ~n17974;
  assign n17976 = ~controllable_hmaster3 & ~n17975;
  assign n17977 = ~n13672 & ~n17976;
  assign n17978 = i_hlock7 & ~n17977;
  assign n17979 = controllable_hmaster2 & ~n17793;
  assign n17980 = ~n13189 & ~n17979;
  assign n17981 = controllable_hmaster1 & ~n17980;
  assign n17982 = ~n13677 & ~n17981;
  assign n17983 = ~controllable_hgrant6 & ~n17982;
  assign n17984 = ~n13687 & ~n17983;
  assign n17985 = controllable_hmaster0 & ~n17984;
  assign n17986 = ~n13682 & ~n17985;
  assign n17987 = ~controllable_hmaster3 & ~n17986;
  assign n17988 = ~n13672 & ~n17987;
  assign n17989 = ~i_hlock7 & ~n17988;
  assign n17990 = ~n17978 & ~n17989;
  assign n17991 = i_hbusreq7 & ~n17990;
  assign n17992 = i_hbusreq8 & ~n17975;
  assign n17993 = i_hbusreq6 & ~n17971;
  assign n17994 = controllable_hmaster2 & ~n17850;
  assign n17995 = ~n13702 & ~n17994;
  assign n17996 = controllable_hmaster1 & ~n17995;
  assign n17997 = ~n13721 & ~n17996;
  assign n17998 = ~i_hbusreq6 & ~n17997;
  assign n17999 = ~n17993 & ~n17998;
  assign n18000 = ~controllable_hgrant6 & ~n17999;
  assign n18001 = ~n13716 & ~n18000;
  assign n18002 = controllable_hmaster0 & ~n18001;
  assign n18003 = ~n13728 & ~n18002;
  assign n18004 = ~i_hbusreq8 & ~n18003;
  assign n18005 = ~n17992 & ~n18004;
  assign n18006 = ~controllable_hmaster3 & ~n18005;
  assign n18007 = ~n13714 & ~n18006;
  assign n18008 = i_hlock7 & ~n18007;
  assign n18009 = i_hbusreq8 & ~n17986;
  assign n18010 = i_hbusreq6 & ~n17982;
  assign n18011 = controllable_hmaster2 & ~n17886;
  assign n18012 = ~n13702 & ~n18011;
  assign n18013 = controllable_hmaster1 & ~n18012;
  assign n18014 = ~n13721 & ~n18013;
  assign n18015 = ~i_hbusreq6 & ~n18014;
  assign n18016 = ~n18010 & ~n18015;
  assign n18017 = ~controllable_hgrant6 & ~n18016;
  assign n18018 = ~n13736 & ~n18017;
  assign n18019 = controllable_hmaster0 & ~n18018;
  assign n18020 = ~n13728 & ~n18019;
  assign n18021 = ~i_hbusreq8 & ~n18020;
  assign n18022 = ~n18009 & ~n18021;
  assign n18023 = ~controllable_hmaster3 & ~n18022;
  assign n18024 = ~n13714 & ~n18023;
  assign n18025 = ~i_hlock7 & ~n18024;
  assign n18026 = ~n18008 & ~n18025;
  assign n18027 = ~i_hbusreq7 & ~n18026;
  assign n18028 = ~n17991 & ~n18027;
  assign n18029 = n7924 & ~n18028;
  assign n18030 = ~n17967 & ~n18029;
  assign n18031 = ~n8214 & ~n18030;
  assign n18032 = i_hlock6 & ~n17912;
  assign n18033 = ~i_hlock6 & ~n17922;
  assign n18034 = ~n18032 & ~n18033;
  assign n18035 = ~controllable_hgrant6 & ~n18034;
  assign n18036 = ~n13766 & ~n18035;
  assign n18037 = ~controllable_hmaster0 & ~n18036;
  assign n18038 = ~n9152 & ~n18037;
  assign n18039 = ~controllable_hmaster3 & ~n18038;
  assign n18040 = ~n13651 & ~n18039;
  assign n18041 = i_hbusreq7 & ~n18040;
  assign n18042 = i_hbusreq8 & ~n18038;
  assign n18043 = i_hbusreq6 & ~n18034;
  assign n18044 = i_hlock6 & ~n17936;
  assign n18045 = ~i_hlock6 & ~n17952;
  assign n18046 = ~n18044 & ~n18045;
  assign n18047 = ~i_hbusreq6 & ~n18046;
  assign n18048 = ~n18043 & ~n18047;
  assign n18049 = ~controllable_hgrant6 & ~n18048;
  assign n18050 = ~n13779 & ~n18049;
  assign n18051 = ~controllable_hmaster0 & ~n18050;
  assign n18052 = ~n9162 & ~n18051;
  assign n18053 = ~i_hbusreq8 & ~n18052;
  assign n18054 = ~n18042 & ~n18053;
  assign n18055 = ~controllable_hmaster3 & ~n18054;
  assign n18056 = ~n13662 & ~n18055;
  assign n18057 = ~i_hbusreq7 & ~n18056;
  assign n18058 = ~n18041 & ~n18057;
  assign n18059 = ~n7924 & ~n18058;
  assign n18060 = i_hlock6 & ~n17971;
  assign n18061 = ~i_hlock6 & ~n17982;
  assign n18062 = ~n18060 & ~n18061;
  assign n18063 = ~controllable_hgrant6 & ~n18062;
  assign n18064 = ~n13766 & ~n18063;
  assign n18065 = ~controllable_hmaster0 & ~n18064;
  assign n18066 = ~n13765 & ~n18065;
  assign n18067 = ~controllable_hmaster3 & ~n18066;
  assign n18068 = ~n13672 & ~n18067;
  assign n18069 = i_hbusreq7 & ~n18068;
  assign n18070 = i_hbusreq8 & ~n18066;
  assign n18071 = i_hbusreq6 & ~n18062;
  assign n18072 = i_hlock6 & ~n17997;
  assign n18073 = ~i_hlock6 & ~n18014;
  assign n18074 = ~n18072 & ~n18073;
  assign n18075 = ~i_hbusreq6 & ~n18074;
  assign n18076 = ~n18071 & ~n18075;
  assign n18077 = ~controllable_hgrant6 & ~n18076;
  assign n18078 = ~n13779 & ~n18077;
  assign n18079 = ~controllable_hmaster0 & ~n18078;
  assign n18080 = ~n13778 & ~n18079;
  assign n18081 = ~i_hbusreq8 & ~n18080;
  assign n18082 = ~n18070 & ~n18081;
  assign n18083 = ~controllable_hmaster3 & ~n18082;
  assign n18084 = ~n13714 & ~n18083;
  assign n18085 = ~i_hbusreq7 & ~n18084;
  assign n18086 = ~n18069 & ~n18085;
  assign n18087 = n7924 & ~n18086;
  assign n18088 = ~n18059 & ~n18087;
  assign n18089 = n8214 & ~n18088;
  assign n18090 = ~n18031 & ~n18089;
  assign n18091 = n8202 & ~n18090;
  assign n18092 = ~n17909 & ~n18091;
  assign n18093 = n7920 & ~n18092;
  assign n18094 = ~n16997 & ~n18093;
  assign n18095 = n7728 & ~n18094;
  assign n18096 = ~n16745 & ~n17324;
  assign n18097 = ~controllable_hmaster1 & ~n18096;
  assign n18098 = ~n17323 & ~n18097;
  assign n18099 = ~controllable_hgrant6 & ~n18098;
  assign n18100 = ~n13406 & ~n18099;
  assign n18101 = ~controllable_hmaster0 & ~n18100;
  assign n18102 = ~n17330 & ~n18101;
  assign n18103 = i_hlock8 & ~n18102;
  assign n18104 = ~n16764 & ~n17324;
  assign n18105 = ~controllable_hmaster1 & ~n18104;
  assign n18106 = ~n17323 & ~n18105;
  assign n18107 = ~controllable_hgrant6 & ~n18106;
  assign n18108 = ~n13427 & ~n18107;
  assign n18109 = ~controllable_hmaster0 & ~n18108;
  assign n18110 = ~n17330 & ~n18109;
  assign n18111 = ~i_hlock8 & ~n18110;
  assign n18112 = ~n18103 & ~n18111;
  assign n18113 = controllable_hmaster3 & ~n18112;
  assign n18114 = i_hlock3 & ~n16738;
  assign n18115 = ~i_hlock3 & ~n16757;
  assign n18116 = ~n18114 & ~n18115;
  assign n18117 = ~controllable_hgrant3 & ~n18116;
  assign n18118 = ~n13852 & ~n18117;
  assign n18119 = ~controllable_hgrant4 & ~n18118;
  assign n18120 = ~n13851 & ~n18119;
  assign n18121 = ~controllable_hgrant5 & ~n18120;
  assign n18122 = ~n13850 & ~n18121;
  assign n18123 = ~controllable_hmaster2 & ~n18122;
  assign n18124 = ~n16896 & ~n18123;
  assign n18125 = controllable_hmaster1 & ~n18124;
  assign n18126 = i_hlock5 & ~n16742;
  assign n18127 = ~i_hlock5 & ~n16761;
  assign n18128 = ~n18126 & ~n18127;
  assign n18129 = ~controllable_hgrant5 & ~n18128;
  assign n18130 = ~n13865 & ~n18129;
  assign n18131 = controllable_hmaster2 & ~n18130;
  assign n18132 = i_hlock1 & ~n16736;
  assign n18133 = ~i_hlock1 & ~n16755;
  assign n18134 = ~n18132 & ~n18133;
  assign n18135 = ~controllable_hgrant1 & ~n18134;
  assign n18136 = ~n13875 & ~n18135;
  assign n18137 = ~controllable_hgrant3 & ~n18136;
  assign n18138 = ~n13874 & ~n18137;
  assign n18139 = ~controllable_hgrant4 & ~n18138;
  assign n18140 = ~n13873 & ~n18139;
  assign n18141 = ~controllable_hgrant5 & ~n18140;
  assign n18142 = ~n13872 & ~n18141;
  assign n18143 = ~controllable_hmaster2 & ~n18142;
  assign n18144 = ~n18131 & ~n18143;
  assign n18145 = ~controllable_hmaster1 & ~n18144;
  assign n18146 = ~n18125 & ~n18145;
  assign n18147 = ~controllable_hgrant6 & ~n18146;
  assign n18148 = ~n13849 & ~n18147;
  assign n18149 = controllable_hmaster0 & ~n18148;
  assign n18150 = ~n9213 & ~n16735;
  assign n18151 = ~controllable_hgrant1 & ~n18150;
  assign n18152 = ~n13898 & ~n18151;
  assign n18153 = ~controllable_hgrant3 & ~n18152;
  assign n18154 = ~n13897 & ~n18153;
  assign n18155 = ~controllable_hgrant4 & ~n18154;
  assign n18156 = ~n13896 & ~n18155;
  assign n18157 = ~controllable_hgrant5 & ~n18156;
  assign n18158 = ~n13895 & ~n18157;
  assign n18159 = ~controllable_hmaster2 & ~n18158;
  assign n18160 = ~n16896 & ~n18159;
  assign n18161 = controllable_hmaster1 & ~n18160;
  assign n18162 = i_hlock4 & ~n16740;
  assign n18163 = ~i_hlock4 & ~n16759;
  assign n18164 = ~n18162 & ~n18163;
  assign n18165 = ~controllable_hgrant4 & ~n18164;
  assign n18166 = ~n13912 & ~n18165;
  assign n18167 = ~controllable_hgrant5 & ~n18166;
  assign n18168 = ~n13911 & ~n18167;
  assign n18169 = controllable_hmaster2 & ~n18168;
  assign n18170 = ~n8440 & ~n16735;
  assign n18171 = ~controllable_hgrant1 & ~n18170;
  assign n18172 = ~n13924 & ~n18171;
  assign n18173 = ~controllable_hgrant3 & ~n18172;
  assign n18174 = ~n13923 & ~n18173;
  assign n18175 = ~controllable_hgrant4 & ~n18174;
  assign n18176 = ~n13922 & ~n18175;
  assign n18177 = ~controllable_hgrant5 & ~n18176;
  assign n18178 = ~n13921 & ~n18177;
  assign n18179 = ~controllable_hmaster2 & ~n18178;
  assign n18180 = ~n18169 & ~n18179;
  assign n18181 = ~controllable_hmaster1 & ~n18180;
  assign n18182 = ~n18161 & ~n18181;
  assign n18183 = i_hlock6 & ~n18182;
  assign n18184 = ~n16908 & ~n18159;
  assign n18185 = controllable_hmaster1 & ~n18184;
  assign n18186 = ~n18181 & ~n18185;
  assign n18187 = ~i_hlock6 & ~n18186;
  assign n18188 = ~n18183 & ~n18187;
  assign n18189 = ~controllable_hgrant6 & ~n18188;
  assign n18190 = ~n13894 & ~n18189;
  assign n18191 = ~controllable_hmaster0 & ~n18190;
  assign n18192 = ~n18149 & ~n18191;
  assign n18193 = ~controllable_hmaster3 & ~n18192;
  assign n18194 = ~n18113 & ~n18193;
  assign n18195 = i_hlock7 & ~n18194;
  assign n18196 = ~n16908 & ~n18123;
  assign n18197 = controllable_hmaster1 & ~n18196;
  assign n18198 = ~n18145 & ~n18197;
  assign n18199 = ~controllable_hgrant6 & ~n18198;
  assign n18200 = ~n13951 & ~n18199;
  assign n18201 = controllable_hmaster0 & ~n18200;
  assign n18202 = ~n18191 & ~n18201;
  assign n18203 = ~controllable_hmaster3 & ~n18202;
  assign n18204 = ~n18113 & ~n18203;
  assign n18205 = ~i_hlock7 & ~n18204;
  assign n18206 = ~n18195 & ~n18205;
  assign n18207 = i_hbusreq7 & ~n18206;
  assign n18208 = i_hbusreq8 & ~n18112;
  assign n18209 = i_hlock0 & ~n7971;
  assign n18210 = ~i_hlock0 & i_hready;
  assign n18211 = ~n18209 & ~n18210;
  assign n18212 = ~i_hbusreq0 & ~n18211;
  assign n18213 = ~n8106 & ~n18212;
  assign n18214 = ~i_hbusreq2 & ~n18213;
  assign n18215 = ~n8105 & ~n18214;
  assign n18216 = ~controllable_hgrant2 & ~n18215;
  assign n18217 = ~n12694 & ~n18216;
  assign n18218 = ~n7733 & ~n18217;
  assign n18219 = i_hlock0 & ~n17364;
  assign n18220 = ~n16807 & ~n18219;
  assign n18221 = ~i_hbusreq0 & ~n18220;
  assign n18222 = ~n16800 & ~n18221;
  assign n18223 = ~i_hbusreq2 & ~n18222;
  assign n18224 = ~n16799 & ~n18223;
  assign n18225 = ~controllable_hgrant2 & ~n18224;
  assign n18226 = ~n12694 & ~n18225;
  assign n18227 = n7733 & ~n18226;
  assign n18228 = ~n18218 & ~n18227;
  assign n18229 = ~i_hbusreq1 & ~n18228;
  assign n18230 = ~n17360 & ~n18229;
  assign n18231 = ~controllable_hgrant1 & ~n18230;
  assign n18232 = ~n13968 & ~n18231;
  assign n18233 = ~i_hbusreq3 & ~n18232;
  assign n18234 = ~n17359 & ~n18233;
  assign n18235 = ~controllable_hgrant3 & ~n18234;
  assign n18236 = ~n13967 & ~n18235;
  assign n18237 = ~i_hbusreq9 & ~n18236;
  assign n18238 = ~n17358 & ~n18237;
  assign n18239 = ~i_hbusreq4 & ~n18238;
  assign n18240 = ~n17357 & ~n18239;
  assign n18241 = ~controllable_hgrant4 & ~n18240;
  assign n18242 = ~n13966 & ~n18241;
  assign n18243 = ~i_hbusreq5 & ~n18242;
  assign n18244 = ~n17356 & ~n18243;
  assign n18245 = ~controllable_hgrant5 & ~n18244;
  assign n18246 = ~n13965 & ~n18245;
  assign n18247 = controllable_hmaster1 & ~n18246;
  assign n18248 = controllable_hmaster2 & ~n18246;
  assign n18249 = ~n16452 & ~n18248;
  assign n18250 = ~controllable_hmaster1 & ~n18249;
  assign n18251 = ~n18247 & ~n18250;
  assign n18252 = ~i_hbusreq6 & ~n18251;
  assign n18253 = ~n17355 & ~n18252;
  assign n18254 = ~controllable_hgrant6 & ~n18253;
  assign n18255 = ~n13818 & ~n18254;
  assign n18256 = controllable_hmaster0 & ~n18255;
  assign n18257 = i_hbusreq6 & ~n18098;
  assign n18258 = ~n16798 & ~n18227;
  assign n18259 = n7928 & ~n18258;
  assign n18260 = ~n8265 & ~n18259;
  assign n18261 = ~i_hbusreq1 & ~n18260;
  assign n18262 = ~n16784 & ~n18261;
  assign n18263 = ~controllable_hgrant1 & ~n18262;
  assign n18264 = ~n14023 & ~n18263;
  assign n18265 = ~i_hbusreq3 & ~n18264;
  assign n18266 = ~n16783 & ~n18265;
  assign n18267 = ~controllable_hgrant3 & ~n18266;
  assign n18268 = ~n14022 & ~n18267;
  assign n18269 = ~i_hbusreq9 & ~n18268;
  assign n18270 = ~n16782 & ~n18269;
  assign n18271 = ~i_hbusreq4 & ~n18270;
  assign n18272 = ~n16781 & ~n18271;
  assign n18273 = ~controllable_hgrant4 & ~n18272;
  assign n18274 = ~n14021 & ~n18273;
  assign n18275 = ~i_hbusreq5 & ~n18274;
  assign n18276 = ~n16780 & ~n18275;
  assign n18277 = ~controllable_hgrant5 & ~n18276;
  assign n18278 = ~n14020 & ~n18277;
  assign n18279 = ~controllable_hmaster2 & ~n18278;
  assign n18280 = ~n18248 & ~n18279;
  assign n18281 = ~controllable_hmaster1 & ~n18280;
  assign n18282 = ~n18247 & ~n18281;
  assign n18283 = ~i_hbusreq6 & ~n18282;
  assign n18284 = ~n18257 & ~n18283;
  assign n18285 = ~controllable_hgrant6 & ~n18284;
  assign n18286 = ~n14019 & ~n18285;
  assign n18287 = ~controllable_hmaster0 & ~n18286;
  assign n18288 = ~n18256 & ~n18287;
  assign n18289 = i_hlock8 & ~n18288;
  assign n18290 = i_hbusreq6 & ~n18106;
  assign n18291 = ~n8297 & ~n18259;
  assign n18292 = ~i_hbusreq1 & ~n18291;
  assign n18293 = ~n16854 & ~n18292;
  assign n18294 = ~controllable_hgrant1 & ~n18293;
  assign n18295 = ~n14058 & ~n18294;
  assign n18296 = ~i_hbusreq3 & ~n18295;
  assign n18297 = ~n16853 & ~n18296;
  assign n18298 = ~controllable_hgrant3 & ~n18297;
  assign n18299 = ~n14057 & ~n18298;
  assign n18300 = ~i_hbusreq9 & ~n18299;
  assign n18301 = ~n16852 & ~n18300;
  assign n18302 = ~i_hbusreq4 & ~n18301;
  assign n18303 = ~n16851 & ~n18302;
  assign n18304 = ~controllable_hgrant4 & ~n18303;
  assign n18305 = ~n14056 & ~n18304;
  assign n18306 = ~i_hbusreq5 & ~n18305;
  assign n18307 = ~n16850 & ~n18306;
  assign n18308 = ~controllable_hgrant5 & ~n18307;
  assign n18309 = ~n14055 & ~n18308;
  assign n18310 = ~controllable_hmaster2 & ~n18309;
  assign n18311 = ~n18248 & ~n18310;
  assign n18312 = ~controllable_hmaster1 & ~n18311;
  assign n18313 = ~n18247 & ~n18312;
  assign n18314 = ~i_hbusreq6 & ~n18313;
  assign n18315 = ~n18290 & ~n18314;
  assign n18316 = ~controllable_hgrant6 & ~n18315;
  assign n18317 = ~n14054 & ~n18316;
  assign n18318 = ~controllable_hmaster0 & ~n18317;
  assign n18319 = ~n18256 & ~n18318;
  assign n18320 = ~i_hlock8 & ~n18319;
  assign n18321 = ~n18289 & ~n18320;
  assign n18322 = ~i_hbusreq8 & ~n18321;
  assign n18323 = ~n18208 & ~n18322;
  assign n18324 = controllable_hmaster3 & ~n18323;
  assign n18325 = i_hbusreq8 & ~n18192;
  assign n18326 = i_hbusreq6 & ~n18146;
  assign n18327 = controllable_hmaster2 & ~n18278;
  assign n18328 = i_hbusreq5 & ~n18120;
  assign n18329 = i_hbusreq4 & ~n18118;
  assign n18330 = i_hbusreq9 & ~n18118;
  assign n18331 = i_hbusreq3 & ~n18116;
  assign n18332 = i_hlock3 & ~n18264;
  assign n18333 = ~i_hlock3 & ~n18295;
  assign n18334 = ~n18332 & ~n18333;
  assign n18335 = ~i_hbusreq3 & ~n18334;
  assign n18336 = ~n18331 & ~n18335;
  assign n18337 = ~controllable_hgrant3 & ~n18336;
  assign n18338 = ~n14102 & ~n18337;
  assign n18339 = ~i_hbusreq9 & ~n18338;
  assign n18340 = ~n18330 & ~n18339;
  assign n18341 = ~i_hbusreq4 & ~n18340;
  assign n18342 = ~n18329 & ~n18341;
  assign n18343 = ~controllable_hgrant4 & ~n18342;
  assign n18344 = ~n14099 & ~n18343;
  assign n18345 = ~i_hbusreq5 & ~n18344;
  assign n18346 = ~n18328 & ~n18345;
  assign n18347 = ~controllable_hgrant5 & ~n18346;
  assign n18348 = ~n14097 & ~n18347;
  assign n18349 = ~controllable_hmaster2 & ~n18348;
  assign n18350 = ~n18327 & ~n18349;
  assign n18351 = controllable_hmaster1 & ~n18350;
  assign n18352 = i_hbusreq5 & ~n18128;
  assign n18353 = i_hlock5 & ~n18274;
  assign n18354 = ~i_hlock5 & ~n18305;
  assign n18355 = ~n18353 & ~n18354;
  assign n18356 = ~i_hbusreq5 & ~n18355;
  assign n18357 = ~n18352 & ~n18356;
  assign n18358 = ~controllable_hgrant5 & ~n18357;
  assign n18359 = ~n14124 & ~n18358;
  assign n18360 = controllable_hmaster2 & ~n18359;
  assign n18361 = i_hbusreq5 & ~n18140;
  assign n18362 = i_hbusreq4 & ~n18138;
  assign n18363 = i_hbusreq9 & ~n18138;
  assign n18364 = i_hbusreq3 & ~n18136;
  assign n18365 = i_hbusreq1 & ~n18134;
  assign n18366 = i_hlock1 & ~n18260;
  assign n18367 = ~i_hlock1 & ~n18291;
  assign n18368 = ~n18366 & ~n18367;
  assign n18369 = ~i_hbusreq1 & ~n18368;
  assign n18370 = ~n18365 & ~n18369;
  assign n18371 = ~controllable_hgrant1 & ~n18370;
  assign n18372 = ~n14141 & ~n18371;
  assign n18373 = ~i_hbusreq3 & ~n18372;
  assign n18374 = ~n18364 & ~n18373;
  assign n18375 = ~controllable_hgrant3 & ~n18374;
  assign n18376 = ~n14139 & ~n18375;
  assign n18377 = ~i_hbusreq9 & ~n18376;
  assign n18378 = ~n18363 & ~n18377;
  assign n18379 = ~i_hbusreq4 & ~n18378;
  assign n18380 = ~n18362 & ~n18379;
  assign n18381 = ~controllable_hgrant4 & ~n18380;
  assign n18382 = ~n14136 & ~n18381;
  assign n18383 = ~i_hbusreq5 & ~n18382;
  assign n18384 = ~n18361 & ~n18383;
  assign n18385 = ~controllable_hgrant5 & ~n18384;
  assign n18386 = ~n14134 & ~n18385;
  assign n18387 = ~controllable_hmaster2 & ~n18386;
  assign n18388 = ~n18360 & ~n18387;
  assign n18389 = ~controllable_hmaster1 & ~n18388;
  assign n18390 = ~n18351 & ~n18389;
  assign n18391 = ~i_hbusreq6 & ~n18390;
  assign n18392 = ~n18326 & ~n18391;
  assign n18393 = ~controllable_hgrant6 & ~n18392;
  assign n18394 = ~n14094 & ~n18393;
  assign n18395 = controllable_hmaster0 & ~n18394;
  assign n18396 = i_hbusreq6 & ~n18188;
  assign n18397 = i_hbusreq5 & ~n18156;
  assign n18398 = i_hbusreq4 & ~n18154;
  assign n18399 = i_hbusreq9 & ~n18154;
  assign n18400 = i_hbusreq3 & ~n18152;
  assign n18401 = i_hbusreq1 & ~n18150;
  assign n18402 = ~n9379 & ~n18259;
  assign n18403 = ~i_hbusreq1 & ~n18402;
  assign n18404 = ~n18401 & ~n18403;
  assign n18405 = ~controllable_hgrant1 & ~n18404;
  assign n18406 = ~n14182 & ~n18405;
  assign n18407 = ~i_hbusreq3 & ~n18406;
  assign n18408 = ~n18400 & ~n18407;
  assign n18409 = ~controllable_hgrant3 & ~n18408;
  assign n18410 = ~n14180 & ~n18409;
  assign n18411 = ~i_hbusreq9 & ~n18410;
  assign n18412 = ~n18399 & ~n18411;
  assign n18413 = ~i_hbusreq4 & ~n18412;
  assign n18414 = ~n18398 & ~n18413;
  assign n18415 = ~controllable_hgrant4 & ~n18414;
  assign n18416 = ~n14177 & ~n18415;
  assign n18417 = ~i_hbusreq5 & ~n18416;
  assign n18418 = ~n18397 & ~n18417;
  assign n18419 = ~controllable_hgrant5 & ~n18418;
  assign n18420 = ~n14175 & ~n18419;
  assign n18421 = ~controllable_hmaster2 & ~n18420;
  assign n18422 = ~n18327 & ~n18421;
  assign n18423 = controllable_hmaster1 & ~n18422;
  assign n18424 = i_hbusreq5 & ~n18166;
  assign n18425 = i_hbusreq4 & ~n18164;
  assign n18426 = i_hlock4 & ~n18270;
  assign n18427 = ~i_hlock4 & ~n18301;
  assign n18428 = ~n18426 & ~n18427;
  assign n18429 = ~i_hbusreq4 & ~n18428;
  assign n18430 = ~n18425 & ~n18429;
  assign n18431 = ~controllable_hgrant4 & ~n18430;
  assign n18432 = ~n14208 & ~n18431;
  assign n18433 = ~i_hbusreq5 & ~n18432;
  assign n18434 = ~n18424 & ~n18433;
  assign n18435 = ~controllable_hgrant5 & ~n18434;
  assign n18436 = ~n14206 & ~n18435;
  assign n18437 = controllable_hmaster2 & ~n18436;
  assign n18438 = i_hbusreq5 & ~n18176;
  assign n18439 = i_hbusreq4 & ~n18174;
  assign n18440 = i_hbusreq9 & ~n18174;
  assign n18441 = i_hbusreq3 & ~n18172;
  assign n18442 = i_hbusreq1 & ~n18170;
  assign n18443 = ~n7933 & ~n17361;
  assign n18444 = ~controllable_locked & ~n18443;
  assign n18445 = ~n14240 & ~n18444;
  assign n18446 = i_hlock0 & ~n18445;
  assign n18447 = ~n16790 & ~n18446;
  assign n18448 = ~i_hbusreq0 & ~n18447;
  assign n18449 = ~n16786 & ~n18448;
  assign n18450 = ~i_hbusreq2 & ~n18449;
  assign n18451 = ~n16785 & ~n18450;
  assign n18452 = ~controllable_hgrant2 & ~n18451;
  assign n18453 = ~n14231 & ~n18452;
  assign n18454 = ~n7733 & ~n18453;
  assign n18455 = ~n7818 & ~n17361;
  assign n18456 = controllable_locked & ~n18455;
  assign n18457 = ~n18444 & ~n18456;
  assign n18458 = i_hlock0 & ~n18457;
  assign n18459 = ~n16807 & ~n18458;
  assign n18460 = ~i_hbusreq0 & ~n18459;
  assign n18461 = ~n16800 & ~n18460;
  assign n18462 = ~i_hbusreq2 & ~n18461;
  assign n18463 = ~n16799 & ~n18462;
  assign n18464 = ~controllable_hgrant2 & ~n18463;
  assign n18465 = ~n14231 & ~n18464;
  assign n18466 = n7733 & ~n18465;
  assign n18467 = ~n18454 & ~n18466;
  assign n18468 = n7928 & ~n18467;
  assign n18469 = ~n8440 & ~n18468;
  assign n18470 = ~i_hbusreq1 & ~n18469;
  assign n18471 = ~n18442 & ~n18470;
  assign n18472 = ~controllable_hgrant1 & ~n18471;
  assign n18473 = ~n14229 & ~n18472;
  assign n18474 = ~i_hbusreq3 & ~n18473;
  assign n18475 = ~n18441 & ~n18474;
  assign n18476 = ~controllable_hgrant3 & ~n18475;
  assign n18477 = ~n14227 & ~n18476;
  assign n18478 = ~i_hbusreq9 & ~n18477;
  assign n18479 = ~n18440 & ~n18478;
  assign n18480 = ~i_hbusreq4 & ~n18479;
  assign n18481 = ~n18439 & ~n18480;
  assign n18482 = ~controllable_hgrant4 & ~n18481;
  assign n18483 = ~n14224 & ~n18482;
  assign n18484 = ~i_hbusreq5 & ~n18483;
  assign n18485 = ~n18438 & ~n18484;
  assign n18486 = ~controllable_hgrant5 & ~n18485;
  assign n18487 = ~n14222 & ~n18486;
  assign n18488 = ~controllable_hmaster2 & ~n18487;
  assign n18489 = ~n18437 & ~n18488;
  assign n18490 = ~controllable_hmaster1 & ~n18489;
  assign n18491 = ~n18423 & ~n18490;
  assign n18492 = i_hlock6 & ~n18491;
  assign n18493 = controllable_hmaster2 & ~n18309;
  assign n18494 = ~n18421 & ~n18493;
  assign n18495 = controllable_hmaster1 & ~n18494;
  assign n18496 = ~n18490 & ~n18495;
  assign n18497 = ~i_hlock6 & ~n18496;
  assign n18498 = ~n18492 & ~n18497;
  assign n18499 = ~i_hbusreq6 & ~n18498;
  assign n18500 = ~n18396 & ~n18499;
  assign n18501 = ~controllable_hgrant6 & ~n18500;
  assign n18502 = ~n14173 & ~n18501;
  assign n18503 = ~controllable_hmaster0 & ~n18502;
  assign n18504 = ~n18395 & ~n18503;
  assign n18505 = ~i_hbusreq8 & ~n18504;
  assign n18506 = ~n18325 & ~n18505;
  assign n18507 = ~controllable_hmaster3 & ~n18506;
  assign n18508 = ~n18324 & ~n18507;
  assign n18509 = i_hlock7 & ~n18508;
  assign n18510 = i_hbusreq8 & ~n18202;
  assign n18511 = i_hbusreq6 & ~n18198;
  assign n18512 = ~n18349 & ~n18493;
  assign n18513 = controllable_hmaster1 & ~n18512;
  assign n18514 = ~n18389 & ~n18513;
  assign n18515 = ~i_hbusreq6 & ~n18514;
  assign n18516 = ~n18511 & ~n18515;
  assign n18517 = ~controllable_hgrant6 & ~n18516;
  assign n18518 = ~n14298 & ~n18517;
  assign n18519 = controllable_hmaster0 & ~n18518;
  assign n18520 = ~n18503 & ~n18519;
  assign n18521 = ~i_hbusreq8 & ~n18520;
  assign n18522 = ~n18510 & ~n18521;
  assign n18523 = ~controllable_hmaster3 & ~n18522;
  assign n18524 = ~n18324 & ~n18523;
  assign n18525 = ~i_hlock7 & ~n18524;
  assign n18526 = ~n18509 & ~n18525;
  assign n18527 = ~i_hbusreq7 & ~n18526;
  assign n18528 = ~n18207 & ~n18527;
  assign n18529 = ~n7924 & ~n18528;
  assign n18530 = ~n8221 & ~n17509;
  assign n18531 = ~controllable_hgrant1 & ~n18530;
  assign n18532 = ~n12611 & ~n18531;
  assign n18533 = ~controllable_hgrant3 & ~n18532;
  assign n18534 = ~n12610 & ~n18533;
  assign n18535 = i_hlock9 & ~n18534;
  assign n18536 = ~n8221 & ~n17517;
  assign n18537 = ~controllable_hgrant1 & ~n18536;
  assign n18538 = ~n12611 & ~n18537;
  assign n18539 = ~controllable_hgrant3 & ~n18538;
  assign n18540 = ~n12610 & ~n18539;
  assign n18541 = ~i_hlock9 & ~n18540;
  assign n18542 = ~n18535 & ~n18541;
  assign n18543 = ~controllable_hgrant4 & ~n18542;
  assign n18544 = ~n13408 & ~n18543;
  assign n18545 = ~controllable_hgrant5 & ~n18544;
  assign n18546 = ~n13407 & ~n18545;
  assign n18547 = ~controllable_hmaster2 & ~n18546;
  assign n18548 = ~n17498 & ~n18547;
  assign n18549 = ~controllable_hmaster1 & ~n18548;
  assign n18550 = ~n17497 & ~n18549;
  assign n18551 = ~controllable_hgrant6 & ~n18550;
  assign n18552 = ~n13406 & ~n18551;
  assign n18553 = ~controllable_hmaster0 & ~n18552;
  assign n18554 = ~n17504 & ~n18553;
  assign n18555 = i_hlock8 & ~n18554;
  assign n18556 = ~n8235 & ~n17509;
  assign n18557 = ~controllable_hgrant1 & ~n18556;
  assign n18558 = ~n12638 & ~n18557;
  assign n18559 = ~controllable_hgrant3 & ~n18558;
  assign n18560 = ~n12637 & ~n18559;
  assign n18561 = i_hlock9 & ~n18560;
  assign n18562 = ~n8235 & ~n17517;
  assign n18563 = ~controllable_hgrant1 & ~n18562;
  assign n18564 = ~n12638 & ~n18563;
  assign n18565 = ~controllable_hgrant3 & ~n18564;
  assign n18566 = ~n12637 & ~n18565;
  assign n18567 = ~i_hlock9 & ~n18566;
  assign n18568 = ~n18561 & ~n18567;
  assign n18569 = ~controllable_hgrant4 & ~n18568;
  assign n18570 = ~n13429 & ~n18569;
  assign n18571 = ~controllable_hgrant5 & ~n18570;
  assign n18572 = ~n13428 & ~n18571;
  assign n18573 = ~controllable_hmaster2 & ~n18572;
  assign n18574 = ~n17498 & ~n18573;
  assign n18575 = ~controllable_hmaster1 & ~n18574;
  assign n18576 = ~n17497 & ~n18575;
  assign n18577 = ~controllable_hgrant6 & ~n18576;
  assign n18578 = ~n13427 & ~n18577;
  assign n18579 = ~controllable_hmaster0 & ~n18578;
  assign n18580 = ~n17504 & ~n18579;
  assign n18581 = ~i_hlock8 & ~n18580;
  assign n18582 = ~n18555 & ~n18581;
  assign n18583 = controllable_hmaster3 & ~n18582;
  assign n18584 = controllable_hmaster2 & ~n18546;
  assign n18585 = i_hlock3 & ~n18532;
  assign n18586 = ~i_hlock3 & ~n18558;
  assign n18587 = ~n18585 & ~n18586;
  assign n18588 = ~controllable_hgrant3 & ~n18587;
  assign n18589 = ~n13852 & ~n18588;
  assign n18590 = i_hlock9 & ~n18589;
  assign n18591 = i_hlock3 & ~n18538;
  assign n18592 = ~i_hlock3 & ~n18564;
  assign n18593 = ~n18591 & ~n18592;
  assign n18594 = ~controllable_hgrant3 & ~n18593;
  assign n18595 = ~n13852 & ~n18594;
  assign n18596 = ~i_hlock9 & ~n18595;
  assign n18597 = ~n18590 & ~n18596;
  assign n18598 = ~controllable_hgrant4 & ~n18597;
  assign n18599 = ~n13851 & ~n18598;
  assign n18600 = ~controllable_hgrant5 & ~n18599;
  assign n18601 = ~n13850 & ~n18600;
  assign n18602 = ~controllable_hmaster2 & ~n18601;
  assign n18603 = ~n18584 & ~n18602;
  assign n18604 = controllable_hmaster1 & ~n18603;
  assign n18605 = i_hlock5 & ~n18544;
  assign n18606 = ~i_hlock5 & ~n18570;
  assign n18607 = ~n18605 & ~n18606;
  assign n18608 = ~controllable_hgrant5 & ~n18607;
  assign n18609 = ~n13865 & ~n18608;
  assign n18610 = controllable_hmaster2 & ~n18609;
  assign n18611 = i_hlock1 & ~n18530;
  assign n18612 = ~i_hlock1 & ~n18556;
  assign n18613 = ~n18611 & ~n18612;
  assign n18614 = ~controllable_hgrant1 & ~n18613;
  assign n18615 = ~n13875 & ~n18614;
  assign n18616 = ~controllable_hgrant3 & ~n18615;
  assign n18617 = ~n13874 & ~n18616;
  assign n18618 = i_hlock9 & ~n18617;
  assign n18619 = i_hlock1 & ~n18536;
  assign n18620 = ~i_hlock1 & ~n18562;
  assign n18621 = ~n18619 & ~n18620;
  assign n18622 = ~controllable_hgrant1 & ~n18621;
  assign n18623 = ~n13875 & ~n18622;
  assign n18624 = ~controllable_hgrant3 & ~n18623;
  assign n18625 = ~n13874 & ~n18624;
  assign n18626 = ~i_hlock9 & ~n18625;
  assign n18627 = ~n18618 & ~n18626;
  assign n18628 = ~controllable_hgrant4 & ~n18627;
  assign n18629 = ~n13873 & ~n18628;
  assign n18630 = ~controllable_hgrant5 & ~n18629;
  assign n18631 = ~n13872 & ~n18630;
  assign n18632 = ~controllable_hmaster2 & ~n18631;
  assign n18633 = ~n18610 & ~n18632;
  assign n18634 = ~controllable_hmaster1 & ~n18633;
  assign n18635 = ~n18604 & ~n18634;
  assign n18636 = ~controllable_hgrant6 & ~n18635;
  assign n18637 = ~n13849 & ~n18636;
  assign n18638 = controllable_hmaster0 & ~n18637;
  assign n18639 = ~n9213 & ~n17509;
  assign n18640 = ~controllable_hgrant1 & ~n18639;
  assign n18641 = ~n13898 & ~n18640;
  assign n18642 = ~controllable_hgrant3 & ~n18641;
  assign n18643 = ~n13897 & ~n18642;
  assign n18644 = i_hlock9 & ~n18643;
  assign n18645 = ~n9213 & ~n17517;
  assign n18646 = ~controllable_hgrant1 & ~n18645;
  assign n18647 = ~n13898 & ~n18646;
  assign n18648 = ~controllable_hgrant3 & ~n18647;
  assign n18649 = ~n13897 & ~n18648;
  assign n18650 = ~i_hlock9 & ~n18649;
  assign n18651 = ~n18644 & ~n18650;
  assign n18652 = ~controllable_hgrant4 & ~n18651;
  assign n18653 = ~n13896 & ~n18652;
  assign n18654 = ~controllable_hgrant5 & ~n18653;
  assign n18655 = ~n13895 & ~n18654;
  assign n18656 = ~controllable_hmaster2 & ~n18655;
  assign n18657 = ~n18584 & ~n18656;
  assign n18658 = controllable_hmaster1 & ~n18657;
  assign n18659 = i_hlock4 & ~n18542;
  assign n18660 = ~i_hlock4 & ~n18568;
  assign n18661 = ~n18659 & ~n18660;
  assign n18662 = ~controllable_hgrant4 & ~n18661;
  assign n18663 = ~n13912 & ~n18662;
  assign n18664 = ~controllable_hgrant5 & ~n18663;
  assign n18665 = ~n13911 & ~n18664;
  assign n18666 = controllable_hmaster2 & ~n18665;
  assign n18667 = ~n8440 & ~n17509;
  assign n18668 = ~controllable_hgrant1 & ~n18667;
  assign n18669 = ~n13924 & ~n18668;
  assign n18670 = ~controllable_hgrant3 & ~n18669;
  assign n18671 = ~n13923 & ~n18670;
  assign n18672 = i_hlock9 & ~n18671;
  assign n18673 = ~n8440 & ~n17517;
  assign n18674 = ~controllable_hgrant1 & ~n18673;
  assign n18675 = ~n13924 & ~n18674;
  assign n18676 = ~controllable_hgrant3 & ~n18675;
  assign n18677 = ~n13923 & ~n18676;
  assign n18678 = ~i_hlock9 & ~n18677;
  assign n18679 = ~n18672 & ~n18678;
  assign n18680 = ~controllable_hgrant4 & ~n18679;
  assign n18681 = ~n13922 & ~n18680;
  assign n18682 = ~controllable_hgrant5 & ~n18681;
  assign n18683 = ~n13921 & ~n18682;
  assign n18684 = ~controllable_hmaster2 & ~n18683;
  assign n18685 = ~n18666 & ~n18684;
  assign n18686 = ~controllable_hmaster1 & ~n18685;
  assign n18687 = ~n18658 & ~n18686;
  assign n18688 = i_hlock6 & ~n18687;
  assign n18689 = controllable_hmaster2 & ~n18572;
  assign n18690 = ~n18656 & ~n18689;
  assign n18691 = controllable_hmaster1 & ~n18690;
  assign n18692 = ~n18686 & ~n18691;
  assign n18693 = ~i_hlock6 & ~n18692;
  assign n18694 = ~n18688 & ~n18693;
  assign n18695 = ~controllable_hgrant6 & ~n18694;
  assign n18696 = ~n13894 & ~n18695;
  assign n18697 = ~controllable_hmaster0 & ~n18696;
  assign n18698 = ~n18638 & ~n18697;
  assign n18699 = ~controllable_hmaster3 & ~n18698;
  assign n18700 = ~n18583 & ~n18699;
  assign n18701 = i_hlock7 & ~n18700;
  assign n18702 = ~n18602 & ~n18689;
  assign n18703 = controllable_hmaster1 & ~n18702;
  assign n18704 = ~n18634 & ~n18703;
  assign n18705 = ~controllable_hgrant6 & ~n18704;
  assign n18706 = ~n13951 & ~n18705;
  assign n18707 = controllable_hmaster0 & ~n18706;
  assign n18708 = ~n18697 & ~n18707;
  assign n18709 = ~controllable_hmaster3 & ~n18708;
  assign n18710 = ~n18583 & ~n18709;
  assign n18711 = ~i_hlock7 & ~n18710;
  assign n18712 = ~n18701 & ~n18711;
  assign n18713 = i_hbusreq7 & ~n18712;
  assign n18714 = i_hbusreq8 & ~n18582;
  assign n18715 = ~n7928 & ~n18228;
  assign n18716 = ~i_hlock0 & n17089;
  assign n18717 = ~n17146 & ~n18716;
  assign n18718 = ~i_hbusreq0 & ~n18717;
  assign n18719 = ~n17142 & ~n18718;
  assign n18720 = ~i_hbusreq2 & ~n18719;
  assign n18721 = ~n17141 & ~n18720;
  assign n18722 = ~controllable_hgrant2 & ~n18721;
  assign n18723 = ~n12694 & ~n18722;
  assign n18724 = ~n7733 & ~n18723;
  assign n18725 = i_hlock0 & ~n17557;
  assign n18726 = ~i_hlock0 & ~n17480;
  assign n18727 = ~n18725 & ~n18726;
  assign n18728 = ~i_hbusreq0 & ~n18727;
  assign n18729 = ~n17552 & ~n18728;
  assign n18730 = ~i_hbusreq2 & ~n18729;
  assign n18731 = ~n17551 & ~n18730;
  assign n18732 = ~controllable_hgrant2 & n18731;
  assign n18733 = ~n12694 & ~n18732;
  assign n18734 = n7733 & ~n18733;
  assign n18735 = ~n18724 & ~n18734;
  assign n18736 = n7928 & ~n18735;
  assign n18737 = ~n18715 & ~n18736;
  assign n18738 = ~i_hbusreq1 & ~n18737;
  assign n18739 = ~n17549 & ~n18738;
  assign n18740 = ~controllable_hgrant1 & ~n18739;
  assign n18741 = ~n13968 & ~n18740;
  assign n18742 = ~i_hbusreq3 & ~n18741;
  assign n18743 = ~n17548 & ~n18742;
  assign n18744 = ~controllable_hgrant3 & ~n18743;
  assign n18745 = ~n13967 & ~n18744;
  assign n18746 = i_hlock9 & ~n18745;
  assign n18747 = ~n17580 & ~n18728;
  assign n18748 = ~i_hbusreq2 & ~n18747;
  assign n18749 = ~n17579 & ~n18748;
  assign n18750 = ~controllable_hgrant2 & n18749;
  assign n18751 = ~n12694 & ~n18750;
  assign n18752 = n7733 & ~n18751;
  assign n18753 = ~n18724 & ~n18752;
  assign n18754 = n7928 & ~n18753;
  assign n18755 = ~n18715 & ~n18754;
  assign n18756 = ~i_hbusreq1 & ~n18755;
  assign n18757 = ~n17578 & ~n18756;
  assign n18758 = ~controllable_hgrant1 & ~n18757;
  assign n18759 = ~n13968 & ~n18758;
  assign n18760 = ~i_hbusreq3 & ~n18759;
  assign n18761 = ~n17577 & ~n18760;
  assign n18762 = ~controllable_hgrant3 & ~n18761;
  assign n18763 = ~n13967 & ~n18762;
  assign n18764 = ~i_hlock9 & ~n18763;
  assign n18765 = ~n18746 & ~n18764;
  assign n18766 = ~i_hbusreq9 & ~n18765;
  assign n18767 = ~n17547 & ~n18766;
  assign n18768 = ~i_hbusreq4 & ~n18767;
  assign n18769 = ~n17546 & ~n18768;
  assign n18770 = ~controllable_hgrant4 & ~n18769;
  assign n18771 = ~n13966 & ~n18770;
  assign n18772 = ~i_hbusreq5 & ~n18771;
  assign n18773 = ~n17545 & ~n18772;
  assign n18774 = ~controllable_hgrant5 & ~n18773;
  assign n18775 = ~n13965 & ~n18774;
  assign n18776 = controllable_hmaster1 & ~n18775;
  assign n18777 = controllable_hmaster2 & ~n18775;
  assign n18778 = ~n16693 & ~n18777;
  assign n18779 = ~controllable_hmaster1 & ~n18778;
  assign n18780 = ~n18776 & ~n18779;
  assign n18781 = ~i_hbusreq6 & ~n18780;
  assign n18782 = ~n17544 & ~n18781;
  assign n18783 = ~controllable_hgrant6 & ~n18782;
  assign n18784 = ~n13818 & ~n18783;
  assign n18785 = controllable_hmaster0 & ~n18784;
  assign n18786 = i_hbusreq6 & ~n18550;
  assign n18787 = i_hbusreq5 & ~n18544;
  assign n18788 = i_hbusreq4 & ~n18542;
  assign n18789 = i_hbusreq9 & ~n18542;
  assign n18790 = i_hbusreq3 & ~n18532;
  assign n18791 = i_hbusreq1 & ~n18530;
  assign n18792 = ~i_hlock0 & n13008;
  assign n18793 = ~n17629 & ~n18792;
  assign n18794 = ~i_hbusreq0 & ~n18793;
  assign n18795 = ~n17627 & ~n18794;
  assign n18796 = ~i_hbusreq2 & ~n18795;
  assign n18797 = ~n17626 & ~n18796;
  assign n18798 = ~controllable_hgrant2 & ~n18797;
  assign n18799 = ~n12694 & ~n18798;
  assign n18800 = ~n7733 & ~n18799;
  assign n18801 = ~n18734 & ~n18800;
  assign n18802 = n7928 & ~n18801;
  assign n18803 = ~n8265 & ~n18802;
  assign n18804 = ~i_hbusreq1 & ~n18803;
  assign n18805 = ~n18791 & ~n18804;
  assign n18806 = ~controllable_hgrant1 & ~n18805;
  assign n18807 = ~n14023 & ~n18806;
  assign n18808 = ~i_hbusreq3 & ~n18807;
  assign n18809 = ~n18790 & ~n18808;
  assign n18810 = ~controllable_hgrant3 & ~n18809;
  assign n18811 = ~n14022 & ~n18810;
  assign n18812 = i_hlock9 & ~n18811;
  assign n18813 = i_hbusreq3 & ~n18538;
  assign n18814 = i_hbusreq1 & ~n18536;
  assign n18815 = ~n18752 & ~n18800;
  assign n18816 = n7928 & ~n18815;
  assign n18817 = ~n8265 & ~n18816;
  assign n18818 = ~i_hbusreq1 & ~n18817;
  assign n18819 = ~n18814 & ~n18818;
  assign n18820 = ~controllable_hgrant1 & ~n18819;
  assign n18821 = ~n14023 & ~n18820;
  assign n18822 = ~i_hbusreq3 & ~n18821;
  assign n18823 = ~n18813 & ~n18822;
  assign n18824 = ~controllable_hgrant3 & ~n18823;
  assign n18825 = ~n14022 & ~n18824;
  assign n18826 = ~i_hlock9 & ~n18825;
  assign n18827 = ~n18812 & ~n18826;
  assign n18828 = ~i_hbusreq9 & ~n18827;
  assign n18829 = ~n18789 & ~n18828;
  assign n18830 = ~i_hbusreq4 & ~n18829;
  assign n18831 = ~n18788 & ~n18830;
  assign n18832 = ~controllable_hgrant4 & ~n18831;
  assign n18833 = ~n14021 & ~n18832;
  assign n18834 = ~i_hbusreq5 & ~n18833;
  assign n18835 = ~n18787 & ~n18834;
  assign n18836 = ~controllable_hgrant5 & ~n18835;
  assign n18837 = ~n14020 & ~n18836;
  assign n18838 = ~controllable_hmaster2 & ~n18837;
  assign n18839 = ~n18777 & ~n18838;
  assign n18840 = ~controllable_hmaster1 & ~n18839;
  assign n18841 = ~n18776 & ~n18840;
  assign n18842 = ~i_hbusreq6 & ~n18841;
  assign n18843 = ~n18786 & ~n18842;
  assign n18844 = ~controllable_hgrant6 & ~n18843;
  assign n18845 = ~n14019 & ~n18844;
  assign n18846 = ~controllable_hmaster0 & ~n18845;
  assign n18847 = ~n18785 & ~n18846;
  assign n18848 = i_hlock8 & ~n18847;
  assign n18849 = i_hbusreq6 & ~n18576;
  assign n18850 = i_hbusreq5 & ~n18570;
  assign n18851 = i_hbusreq4 & ~n18568;
  assign n18852 = i_hbusreq9 & ~n18568;
  assign n18853 = i_hbusreq3 & ~n18558;
  assign n18854 = i_hbusreq1 & ~n18556;
  assign n18855 = ~n8297 & ~n18802;
  assign n18856 = ~i_hbusreq1 & ~n18855;
  assign n18857 = ~n18854 & ~n18856;
  assign n18858 = ~controllable_hgrant1 & ~n18857;
  assign n18859 = ~n14058 & ~n18858;
  assign n18860 = ~i_hbusreq3 & ~n18859;
  assign n18861 = ~n18853 & ~n18860;
  assign n18862 = ~controllable_hgrant3 & ~n18861;
  assign n18863 = ~n14057 & ~n18862;
  assign n18864 = i_hlock9 & ~n18863;
  assign n18865 = i_hbusreq3 & ~n18564;
  assign n18866 = i_hbusreq1 & ~n18562;
  assign n18867 = ~n8297 & ~n18816;
  assign n18868 = ~i_hbusreq1 & ~n18867;
  assign n18869 = ~n18866 & ~n18868;
  assign n18870 = ~controllable_hgrant1 & ~n18869;
  assign n18871 = ~n14058 & ~n18870;
  assign n18872 = ~i_hbusreq3 & ~n18871;
  assign n18873 = ~n18865 & ~n18872;
  assign n18874 = ~controllable_hgrant3 & ~n18873;
  assign n18875 = ~n14057 & ~n18874;
  assign n18876 = ~i_hlock9 & ~n18875;
  assign n18877 = ~n18864 & ~n18876;
  assign n18878 = ~i_hbusreq9 & ~n18877;
  assign n18879 = ~n18852 & ~n18878;
  assign n18880 = ~i_hbusreq4 & ~n18879;
  assign n18881 = ~n18851 & ~n18880;
  assign n18882 = ~controllable_hgrant4 & ~n18881;
  assign n18883 = ~n14056 & ~n18882;
  assign n18884 = ~i_hbusreq5 & ~n18883;
  assign n18885 = ~n18850 & ~n18884;
  assign n18886 = ~controllable_hgrant5 & ~n18885;
  assign n18887 = ~n14055 & ~n18886;
  assign n18888 = ~controllable_hmaster2 & ~n18887;
  assign n18889 = ~n18777 & ~n18888;
  assign n18890 = ~controllable_hmaster1 & ~n18889;
  assign n18891 = ~n18776 & ~n18890;
  assign n18892 = ~i_hbusreq6 & ~n18891;
  assign n18893 = ~n18849 & ~n18892;
  assign n18894 = ~controllable_hgrant6 & ~n18893;
  assign n18895 = ~n14054 & ~n18894;
  assign n18896 = ~controllable_hmaster0 & ~n18895;
  assign n18897 = ~n18785 & ~n18896;
  assign n18898 = ~i_hlock8 & ~n18897;
  assign n18899 = ~n18848 & ~n18898;
  assign n18900 = ~i_hbusreq8 & ~n18899;
  assign n18901 = ~n18714 & ~n18900;
  assign n18902 = controllable_hmaster3 & ~n18901;
  assign n18903 = i_hbusreq8 & ~n18698;
  assign n18904 = i_hbusreq6 & ~n18635;
  assign n18905 = controllable_hmaster2 & ~n18837;
  assign n18906 = i_hbusreq5 & ~n18599;
  assign n18907 = i_hbusreq4 & ~n18597;
  assign n18908 = i_hbusreq9 & ~n18597;
  assign n18909 = i_hbusreq3 & ~n18587;
  assign n18910 = i_hlock3 & ~n18807;
  assign n18911 = ~i_hlock3 & ~n18859;
  assign n18912 = ~n18910 & ~n18911;
  assign n18913 = ~i_hbusreq3 & ~n18912;
  assign n18914 = ~n18909 & ~n18913;
  assign n18915 = ~controllable_hgrant3 & ~n18914;
  assign n18916 = ~n14102 & ~n18915;
  assign n18917 = i_hlock9 & ~n18916;
  assign n18918 = i_hbusreq3 & ~n18593;
  assign n18919 = i_hlock3 & ~n18821;
  assign n18920 = ~i_hlock3 & ~n18871;
  assign n18921 = ~n18919 & ~n18920;
  assign n18922 = ~i_hbusreq3 & ~n18921;
  assign n18923 = ~n18918 & ~n18922;
  assign n18924 = ~controllable_hgrant3 & ~n18923;
  assign n18925 = ~n14102 & ~n18924;
  assign n18926 = ~i_hlock9 & ~n18925;
  assign n18927 = ~n18917 & ~n18926;
  assign n18928 = ~i_hbusreq9 & ~n18927;
  assign n18929 = ~n18908 & ~n18928;
  assign n18930 = ~i_hbusreq4 & ~n18929;
  assign n18931 = ~n18907 & ~n18930;
  assign n18932 = ~controllable_hgrant4 & ~n18931;
  assign n18933 = ~n14099 & ~n18932;
  assign n18934 = ~i_hbusreq5 & ~n18933;
  assign n18935 = ~n18906 & ~n18934;
  assign n18936 = ~controllable_hgrant5 & ~n18935;
  assign n18937 = ~n14097 & ~n18936;
  assign n18938 = ~controllable_hmaster2 & ~n18937;
  assign n18939 = ~n18905 & ~n18938;
  assign n18940 = controllable_hmaster1 & ~n18939;
  assign n18941 = i_hbusreq5 & ~n18607;
  assign n18942 = i_hlock5 & ~n18833;
  assign n18943 = ~i_hlock5 & ~n18883;
  assign n18944 = ~n18942 & ~n18943;
  assign n18945 = ~i_hbusreq5 & ~n18944;
  assign n18946 = ~n18941 & ~n18945;
  assign n18947 = ~controllable_hgrant5 & ~n18946;
  assign n18948 = ~n14124 & ~n18947;
  assign n18949 = controllable_hmaster2 & ~n18948;
  assign n18950 = i_hbusreq5 & ~n18629;
  assign n18951 = i_hbusreq4 & ~n18627;
  assign n18952 = i_hbusreq9 & ~n18627;
  assign n18953 = i_hbusreq3 & ~n18615;
  assign n18954 = i_hbusreq1 & ~n18613;
  assign n18955 = i_hlock1 & ~n18803;
  assign n18956 = ~i_hlock1 & ~n18855;
  assign n18957 = ~n18955 & ~n18956;
  assign n18958 = ~i_hbusreq1 & ~n18957;
  assign n18959 = ~n18954 & ~n18958;
  assign n18960 = ~controllable_hgrant1 & ~n18959;
  assign n18961 = ~n14141 & ~n18960;
  assign n18962 = ~i_hbusreq3 & ~n18961;
  assign n18963 = ~n18953 & ~n18962;
  assign n18964 = ~controllable_hgrant3 & ~n18963;
  assign n18965 = ~n14139 & ~n18964;
  assign n18966 = i_hlock9 & ~n18965;
  assign n18967 = i_hbusreq3 & ~n18623;
  assign n18968 = i_hbusreq1 & ~n18621;
  assign n18969 = i_hlock1 & ~n18817;
  assign n18970 = ~i_hlock1 & ~n18867;
  assign n18971 = ~n18969 & ~n18970;
  assign n18972 = ~i_hbusreq1 & ~n18971;
  assign n18973 = ~n18968 & ~n18972;
  assign n18974 = ~controllable_hgrant1 & ~n18973;
  assign n18975 = ~n14141 & ~n18974;
  assign n18976 = ~i_hbusreq3 & ~n18975;
  assign n18977 = ~n18967 & ~n18976;
  assign n18978 = ~controllable_hgrant3 & ~n18977;
  assign n18979 = ~n14139 & ~n18978;
  assign n18980 = ~i_hlock9 & ~n18979;
  assign n18981 = ~n18966 & ~n18980;
  assign n18982 = ~i_hbusreq9 & ~n18981;
  assign n18983 = ~n18952 & ~n18982;
  assign n18984 = ~i_hbusreq4 & ~n18983;
  assign n18985 = ~n18951 & ~n18984;
  assign n18986 = ~controllable_hgrant4 & ~n18985;
  assign n18987 = ~n14136 & ~n18986;
  assign n18988 = ~i_hbusreq5 & ~n18987;
  assign n18989 = ~n18950 & ~n18988;
  assign n18990 = ~controllable_hgrant5 & ~n18989;
  assign n18991 = ~n14134 & ~n18990;
  assign n18992 = ~controllable_hmaster2 & ~n18991;
  assign n18993 = ~n18949 & ~n18992;
  assign n18994 = ~controllable_hmaster1 & ~n18993;
  assign n18995 = ~n18940 & ~n18994;
  assign n18996 = ~i_hbusreq6 & ~n18995;
  assign n18997 = ~n18904 & ~n18996;
  assign n18998 = ~controllable_hgrant6 & ~n18997;
  assign n18999 = ~n14094 & ~n18998;
  assign n19000 = controllable_hmaster0 & ~n18999;
  assign n19001 = i_hbusreq6 & ~n18694;
  assign n19002 = i_hbusreq5 & ~n18653;
  assign n19003 = i_hbusreq4 & ~n18651;
  assign n19004 = i_hbusreq9 & ~n18651;
  assign n19005 = i_hbusreq3 & ~n18641;
  assign n19006 = i_hbusreq1 & ~n18639;
  assign n19007 = ~n9379 & ~n18802;
  assign n19008 = ~i_hbusreq1 & ~n19007;
  assign n19009 = ~n19006 & ~n19008;
  assign n19010 = ~controllable_hgrant1 & ~n19009;
  assign n19011 = ~n14182 & ~n19010;
  assign n19012 = ~i_hbusreq3 & ~n19011;
  assign n19013 = ~n19005 & ~n19012;
  assign n19014 = ~controllable_hgrant3 & ~n19013;
  assign n19015 = ~n14180 & ~n19014;
  assign n19016 = i_hlock9 & ~n19015;
  assign n19017 = i_hbusreq3 & ~n18647;
  assign n19018 = i_hbusreq1 & ~n18645;
  assign n19019 = ~n9379 & ~n18816;
  assign n19020 = ~i_hbusreq1 & ~n19019;
  assign n19021 = ~n19018 & ~n19020;
  assign n19022 = ~controllable_hgrant1 & ~n19021;
  assign n19023 = ~n14182 & ~n19022;
  assign n19024 = ~i_hbusreq3 & ~n19023;
  assign n19025 = ~n19017 & ~n19024;
  assign n19026 = ~controllable_hgrant3 & ~n19025;
  assign n19027 = ~n14180 & ~n19026;
  assign n19028 = ~i_hlock9 & ~n19027;
  assign n19029 = ~n19016 & ~n19028;
  assign n19030 = ~i_hbusreq9 & ~n19029;
  assign n19031 = ~n19004 & ~n19030;
  assign n19032 = ~i_hbusreq4 & ~n19031;
  assign n19033 = ~n19003 & ~n19032;
  assign n19034 = ~controllable_hgrant4 & ~n19033;
  assign n19035 = ~n14177 & ~n19034;
  assign n19036 = ~i_hbusreq5 & ~n19035;
  assign n19037 = ~n19002 & ~n19036;
  assign n19038 = ~controllable_hgrant5 & ~n19037;
  assign n19039 = ~n14175 & ~n19038;
  assign n19040 = ~controllable_hmaster2 & ~n19039;
  assign n19041 = ~n18905 & ~n19040;
  assign n19042 = controllable_hmaster1 & ~n19041;
  assign n19043 = i_hbusreq5 & ~n18663;
  assign n19044 = i_hbusreq4 & ~n18661;
  assign n19045 = i_hlock4 & ~n18829;
  assign n19046 = ~i_hlock4 & ~n18879;
  assign n19047 = ~n19045 & ~n19046;
  assign n19048 = ~i_hbusreq4 & ~n19047;
  assign n19049 = ~n19044 & ~n19048;
  assign n19050 = ~controllable_hgrant4 & ~n19049;
  assign n19051 = ~n14208 & ~n19050;
  assign n19052 = ~i_hbusreq5 & ~n19051;
  assign n19053 = ~n19043 & ~n19052;
  assign n19054 = ~controllable_hgrant5 & ~n19053;
  assign n19055 = ~n14206 & ~n19054;
  assign n19056 = controllable_hmaster2 & ~n19055;
  assign n19057 = i_hbusreq5 & ~n18681;
  assign n19058 = i_hbusreq4 & ~n18679;
  assign n19059 = i_hbusreq9 & ~n18679;
  assign n19060 = i_hbusreq3 & ~n18669;
  assign n19061 = i_hbusreq1 & ~n18667;
  assign n19062 = ~controllable_locked & n12895;
  assign n19063 = ~n14240 & ~n19062;
  assign n19064 = i_hlock0 & ~n19063;
  assign n19065 = ~n18792 & ~n19064;
  assign n19066 = ~i_hbusreq0 & ~n19065;
  assign n19067 = ~n17627 & ~n19066;
  assign n19068 = ~i_hbusreq2 & ~n19067;
  assign n19069 = ~n17626 & ~n19068;
  assign n19070 = ~controllable_hgrant2 & ~n19069;
  assign n19071 = ~n14231 & ~n19070;
  assign n19072 = ~n7733 & ~n19071;
  assign n19073 = ~n12624 & ~n17477;
  assign n19074 = controllable_locked & ~n19073;
  assign n19075 = ~controllable_locked & ~n8232;
  assign n19076 = ~n19074 & ~n19075;
  assign n19077 = i_hlock0 & ~n19076;
  assign n19078 = ~n18726 & ~n19077;
  assign n19079 = ~i_hbusreq0 & ~n19078;
  assign n19080 = ~n17552 & ~n19079;
  assign n19081 = ~i_hbusreq2 & ~n19080;
  assign n19082 = ~n17551 & ~n19081;
  assign n19083 = ~controllable_hgrant2 & n19082;
  assign n19084 = ~n14231 & ~n19083;
  assign n19085 = n7733 & ~n19084;
  assign n19086 = ~n19072 & ~n19085;
  assign n19087 = n7928 & ~n19086;
  assign n19088 = ~n8440 & ~n19087;
  assign n19089 = ~i_hbusreq1 & ~n19088;
  assign n19090 = ~n19061 & ~n19089;
  assign n19091 = ~controllable_hgrant1 & ~n19090;
  assign n19092 = ~n14229 & ~n19091;
  assign n19093 = ~i_hbusreq3 & ~n19092;
  assign n19094 = ~n19060 & ~n19093;
  assign n19095 = ~controllable_hgrant3 & ~n19094;
  assign n19096 = ~n14227 & ~n19095;
  assign n19097 = i_hlock9 & ~n19096;
  assign n19098 = i_hbusreq3 & ~n18675;
  assign n19099 = i_hbusreq1 & ~n18673;
  assign n19100 = ~n17580 & ~n19079;
  assign n19101 = ~i_hbusreq2 & ~n19100;
  assign n19102 = ~n17579 & ~n19101;
  assign n19103 = ~controllable_hgrant2 & n19102;
  assign n19104 = ~n14231 & ~n19103;
  assign n19105 = n7733 & ~n19104;
  assign n19106 = ~n19072 & ~n19105;
  assign n19107 = n7928 & ~n19106;
  assign n19108 = ~n8440 & ~n19107;
  assign n19109 = ~i_hbusreq1 & ~n19108;
  assign n19110 = ~n19099 & ~n19109;
  assign n19111 = ~controllable_hgrant1 & ~n19110;
  assign n19112 = ~n14229 & ~n19111;
  assign n19113 = ~i_hbusreq3 & ~n19112;
  assign n19114 = ~n19098 & ~n19113;
  assign n19115 = ~controllable_hgrant3 & ~n19114;
  assign n19116 = ~n14227 & ~n19115;
  assign n19117 = ~i_hlock9 & ~n19116;
  assign n19118 = ~n19097 & ~n19117;
  assign n19119 = ~i_hbusreq9 & ~n19118;
  assign n19120 = ~n19059 & ~n19119;
  assign n19121 = ~i_hbusreq4 & ~n19120;
  assign n19122 = ~n19058 & ~n19121;
  assign n19123 = ~controllable_hgrant4 & ~n19122;
  assign n19124 = ~n14224 & ~n19123;
  assign n19125 = ~i_hbusreq5 & ~n19124;
  assign n19126 = ~n19057 & ~n19125;
  assign n19127 = ~controllable_hgrant5 & ~n19126;
  assign n19128 = ~n14222 & ~n19127;
  assign n19129 = ~controllable_hmaster2 & ~n19128;
  assign n19130 = ~n19056 & ~n19129;
  assign n19131 = ~controllable_hmaster1 & ~n19130;
  assign n19132 = ~n19042 & ~n19131;
  assign n19133 = i_hlock6 & ~n19132;
  assign n19134 = controllable_hmaster2 & ~n18887;
  assign n19135 = ~n19040 & ~n19134;
  assign n19136 = controllable_hmaster1 & ~n19135;
  assign n19137 = ~n19131 & ~n19136;
  assign n19138 = ~i_hlock6 & ~n19137;
  assign n19139 = ~n19133 & ~n19138;
  assign n19140 = ~i_hbusreq6 & ~n19139;
  assign n19141 = ~n19001 & ~n19140;
  assign n19142 = ~controllable_hgrant6 & ~n19141;
  assign n19143 = ~n14173 & ~n19142;
  assign n19144 = ~controllable_hmaster0 & ~n19143;
  assign n19145 = ~n19000 & ~n19144;
  assign n19146 = ~i_hbusreq8 & ~n19145;
  assign n19147 = ~n18903 & ~n19146;
  assign n19148 = ~controllable_hmaster3 & ~n19147;
  assign n19149 = ~n18902 & ~n19148;
  assign n19150 = i_hlock7 & ~n19149;
  assign n19151 = i_hbusreq8 & ~n18708;
  assign n19152 = i_hbusreq6 & ~n18704;
  assign n19153 = ~n18938 & ~n19134;
  assign n19154 = controllable_hmaster1 & ~n19153;
  assign n19155 = ~n18994 & ~n19154;
  assign n19156 = ~i_hbusreq6 & ~n19155;
  assign n19157 = ~n19152 & ~n19156;
  assign n19158 = ~controllable_hgrant6 & ~n19157;
  assign n19159 = ~n14298 & ~n19158;
  assign n19160 = controllable_hmaster0 & ~n19159;
  assign n19161 = ~n19144 & ~n19160;
  assign n19162 = ~i_hbusreq8 & ~n19161;
  assign n19163 = ~n19151 & ~n19162;
  assign n19164 = ~controllable_hmaster3 & ~n19163;
  assign n19165 = ~n18902 & ~n19164;
  assign n19166 = ~i_hlock7 & ~n19165;
  assign n19167 = ~n19150 & ~n19166;
  assign n19168 = ~i_hbusreq7 & ~n19167;
  assign n19169 = ~n18713 & ~n19168;
  assign n19170 = n7924 & ~n19169;
  assign n19171 = ~n18529 & ~n19170;
  assign n19172 = ~n8214 & ~n19171;
  assign n19173 = ~controllable_hgrant1 & ~n16725;
  assign n19174 = ~n13155 & ~n19173;
  assign n19175 = ~controllable_hgrant3 & ~n19174;
  assign n19176 = ~n13154 & ~n19175;
  assign n19177 = ~controllable_hgrant4 & ~n19176;
  assign n19178 = ~n13153 & ~n19177;
  assign n19179 = ~controllable_hgrant5 & ~n19178;
  assign n19180 = ~n13152 & ~n19179;
  assign n19181 = controllable_hmaster1 & ~n19180;
  assign n19182 = controllable_hmaster2 & ~n19180;
  assign n19183 = n7928 & ~n16350;
  assign n19184 = ~n16128 & ~n19183;
  assign n19185 = ~controllable_hgrant1 & ~n19184;
  assign n19186 = ~n12611 & ~n19185;
  assign n19187 = ~controllable_hgrant3 & ~n19186;
  assign n19188 = ~n12610 & ~n19187;
  assign n19189 = i_hlock9 & ~n19188;
  assign n19190 = ~n16146 & ~n19183;
  assign n19191 = ~controllable_hgrant1 & ~n19190;
  assign n19192 = ~n12638 & ~n19191;
  assign n19193 = ~controllable_hgrant3 & ~n19192;
  assign n19194 = ~n12637 & ~n19193;
  assign n19195 = ~i_hlock9 & ~n19194;
  assign n19196 = ~n19189 & ~n19195;
  assign n19197 = ~controllable_hgrant4 & ~n19196;
  assign n19198 = ~n12609 & ~n19197;
  assign n19199 = ~controllable_hgrant5 & ~n19198;
  assign n19200 = ~n12608 & ~n19199;
  assign n19201 = ~controllable_hmaster2 & ~n19200;
  assign n19202 = ~n19182 & ~n19201;
  assign n19203 = ~controllable_hmaster1 & ~n19202;
  assign n19204 = ~n19181 & ~n19203;
  assign n19205 = ~controllable_hgrant6 & ~n19204;
  assign n19206 = ~n13122 & ~n19205;
  assign n19207 = controllable_hmaster0 & ~n19206;
  assign n19208 = ~n16745 & ~n19182;
  assign n19209 = ~controllable_hmaster1 & ~n19208;
  assign n19210 = ~n19181 & ~n19209;
  assign n19211 = ~controllable_hgrant6 & ~n19210;
  assign n19212 = ~n13406 & ~n19211;
  assign n19213 = ~controllable_hmaster0 & ~n19212;
  assign n19214 = ~n19207 & ~n19213;
  assign n19215 = i_hlock8 & ~n19214;
  assign n19216 = ~n16764 & ~n19182;
  assign n19217 = ~controllable_hmaster1 & ~n19216;
  assign n19218 = ~n19181 & ~n19217;
  assign n19219 = ~controllable_hgrant6 & ~n19218;
  assign n19220 = ~n13427 & ~n19219;
  assign n19221 = ~controllable_hmaster0 & ~n19220;
  assign n19222 = ~n19207 & ~n19221;
  assign n19223 = ~i_hlock8 & ~n19222;
  assign n19224 = ~n19215 & ~n19223;
  assign n19225 = controllable_hmaster3 & ~n19224;
  assign n19226 = n7928 & ~n16725;
  assign n19227 = ~n8221 & ~n19226;
  assign n19228 = ~controllable_hgrant1 & ~n19227;
  assign n19229 = ~n12611 & ~n19228;
  assign n19230 = ~controllable_hgrant3 & ~n19229;
  assign n19231 = ~n12610 & ~n19230;
  assign n19232 = ~controllable_hgrant4 & ~n19231;
  assign n19233 = ~n13408 & ~n19232;
  assign n19234 = ~controllable_hgrant5 & ~n19233;
  assign n19235 = ~n13407 & ~n19234;
  assign n19236 = controllable_hmaster2 & ~n19235;
  assign n19237 = i_hlock3 & ~n19229;
  assign n19238 = ~n8235 & ~n19226;
  assign n19239 = ~controllable_hgrant1 & ~n19238;
  assign n19240 = ~n12638 & ~n19239;
  assign n19241 = ~i_hlock3 & ~n19240;
  assign n19242 = ~n19237 & ~n19241;
  assign n19243 = ~controllable_hgrant3 & ~n19242;
  assign n19244 = ~n13852 & ~n19243;
  assign n19245 = ~controllable_hgrant4 & ~n19244;
  assign n19246 = ~n13851 & ~n19245;
  assign n19247 = ~controllable_hgrant5 & ~n19246;
  assign n19248 = ~n13850 & ~n19247;
  assign n19249 = ~controllable_hmaster2 & ~n19248;
  assign n19250 = ~n19236 & ~n19249;
  assign n19251 = controllable_hmaster1 & ~n19250;
  assign n19252 = i_hlock5 & ~n19233;
  assign n19253 = ~controllable_hgrant3 & ~n19240;
  assign n19254 = ~n12637 & ~n19253;
  assign n19255 = ~controllable_hgrant4 & ~n19254;
  assign n19256 = ~n13429 & ~n19255;
  assign n19257 = ~i_hlock5 & ~n19256;
  assign n19258 = ~n19252 & ~n19257;
  assign n19259 = ~controllable_hgrant5 & ~n19258;
  assign n19260 = ~n13865 & ~n19259;
  assign n19261 = controllable_hmaster2 & ~n19260;
  assign n19262 = i_hlock1 & ~n19227;
  assign n19263 = ~i_hlock1 & ~n19238;
  assign n19264 = ~n19262 & ~n19263;
  assign n19265 = ~controllable_hgrant1 & ~n19264;
  assign n19266 = ~n13875 & ~n19265;
  assign n19267 = ~controllable_hgrant3 & ~n19266;
  assign n19268 = ~n13874 & ~n19267;
  assign n19269 = ~controllable_hgrant4 & ~n19268;
  assign n19270 = ~n13873 & ~n19269;
  assign n19271 = ~controllable_hgrant5 & ~n19270;
  assign n19272 = ~n13872 & ~n19271;
  assign n19273 = ~controllable_hmaster2 & ~n19272;
  assign n19274 = ~n19261 & ~n19273;
  assign n19275 = ~controllable_hmaster1 & ~n19274;
  assign n19276 = ~n19251 & ~n19275;
  assign n19277 = ~controllable_hgrant6 & ~n19276;
  assign n19278 = ~n13849 & ~n19277;
  assign n19279 = controllable_hmaster0 & ~n19278;
  assign n19280 = ~n9213 & ~n19226;
  assign n19281 = ~controllable_hgrant1 & ~n19280;
  assign n19282 = ~n13898 & ~n19281;
  assign n19283 = ~controllable_hgrant3 & ~n19282;
  assign n19284 = ~n13897 & ~n19283;
  assign n19285 = ~controllable_hgrant4 & ~n19284;
  assign n19286 = ~n13896 & ~n19285;
  assign n19287 = ~controllable_hgrant5 & ~n19286;
  assign n19288 = ~n13895 & ~n19287;
  assign n19289 = ~controllable_hmaster2 & ~n19288;
  assign n19290 = ~n19236 & ~n19289;
  assign n19291 = controllable_hmaster1 & ~n19290;
  assign n19292 = i_hlock4 & ~n19231;
  assign n19293 = ~i_hlock4 & ~n19254;
  assign n19294 = ~n19292 & ~n19293;
  assign n19295 = ~controllable_hgrant4 & ~n19294;
  assign n19296 = ~n13912 & ~n19295;
  assign n19297 = ~controllable_hgrant5 & ~n19296;
  assign n19298 = ~n13911 & ~n19297;
  assign n19299 = controllable_hmaster2 & ~n19298;
  assign n19300 = ~n8440 & ~n19226;
  assign n19301 = ~controllable_hgrant1 & ~n19300;
  assign n19302 = ~n13924 & ~n19301;
  assign n19303 = ~controllable_hgrant3 & ~n19302;
  assign n19304 = ~n13923 & ~n19303;
  assign n19305 = ~controllable_hgrant4 & ~n19304;
  assign n19306 = ~n13922 & ~n19305;
  assign n19307 = ~controllable_hgrant5 & ~n19306;
  assign n19308 = ~n13921 & ~n19307;
  assign n19309 = ~controllable_hmaster2 & ~n19308;
  assign n19310 = ~n19299 & ~n19309;
  assign n19311 = ~controllable_hmaster1 & ~n19310;
  assign n19312 = ~n19291 & ~n19311;
  assign n19313 = i_hlock6 & ~n19312;
  assign n19314 = ~controllable_hgrant5 & ~n19256;
  assign n19315 = ~n13428 & ~n19314;
  assign n19316 = controllable_hmaster2 & ~n19315;
  assign n19317 = ~n19289 & ~n19316;
  assign n19318 = controllable_hmaster1 & ~n19317;
  assign n19319 = ~n19311 & ~n19318;
  assign n19320 = ~i_hlock6 & ~n19319;
  assign n19321 = ~n19313 & ~n19320;
  assign n19322 = ~controllable_hgrant6 & ~n19321;
  assign n19323 = ~n13894 & ~n19322;
  assign n19324 = ~controllable_hmaster0 & ~n19323;
  assign n19325 = ~n19279 & ~n19324;
  assign n19326 = ~controllable_hmaster3 & ~n19325;
  assign n19327 = ~n19225 & ~n19326;
  assign n19328 = i_hlock7 & ~n19327;
  assign n19329 = ~n19249 & ~n19316;
  assign n19330 = controllable_hmaster1 & ~n19329;
  assign n19331 = ~n19275 & ~n19330;
  assign n19332 = ~controllable_hgrant6 & ~n19331;
  assign n19333 = ~n13951 & ~n19332;
  assign n19334 = controllable_hmaster0 & ~n19333;
  assign n19335 = ~n19324 & ~n19334;
  assign n19336 = ~controllable_hmaster3 & ~n19335;
  assign n19337 = ~n19225 & ~n19336;
  assign n19338 = ~i_hlock7 & ~n19337;
  assign n19339 = ~n19328 & ~n19338;
  assign n19340 = i_hbusreq7 & ~n19339;
  assign n19341 = i_hbusreq8 & ~n19224;
  assign n19342 = i_hbusreq6 & ~n19204;
  assign n19343 = i_hbusreq5 & ~n19178;
  assign n19344 = i_hbusreq4 & ~n19176;
  assign n19345 = i_hbusreq9 & ~n19176;
  assign n19346 = i_hbusreq3 & ~n19174;
  assign n19347 = i_hbusreq1 & ~n16725;
  assign n19348 = ~i_hbusreq1 & ~n16797;
  assign n19349 = ~n19347 & ~n19348;
  assign n19350 = ~controllable_hgrant1 & ~n19349;
  assign n19351 = ~n13968 & ~n19350;
  assign n19352 = ~i_hbusreq3 & ~n19351;
  assign n19353 = ~n19346 & ~n19352;
  assign n19354 = ~controllable_hgrant3 & ~n19353;
  assign n19355 = ~n13967 & ~n19354;
  assign n19356 = ~i_hbusreq9 & ~n19355;
  assign n19357 = ~n19345 & ~n19356;
  assign n19358 = ~i_hbusreq4 & ~n19357;
  assign n19359 = ~n19344 & ~n19358;
  assign n19360 = ~controllable_hgrant4 & ~n19359;
  assign n19361 = ~n13966 & ~n19360;
  assign n19362 = ~i_hbusreq5 & ~n19361;
  assign n19363 = ~n19343 & ~n19362;
  assign n19364 = ~controllable_hgrant5 & ~n19363;
  assign n19365 = ~n13965 & ~n19364;
  assign n19366 = controllable_hmaster1 & ~n19365;
  assign n19367 = controllable_hmaster2 & ~n19365;
  assign n19368 = i_hbusreq5 & ~n19198;
  assign n19369 = i_hbusreq4 & ~n19196;
  assign n19370 = i_hbusreq9 & ~n19196;
  assign n19371 = i_hbusreq3 & ~n19186;
  assign n19372 = i_hbusreq1 & ~n19184;
  assign n19373 = n7928 & ~n16401;
  assign n19374 = ~n16191 & ~n19373;
  assign n19375 = ~i_hbusreq1 & ~n19374;
  assign n19376 = ~n19372 & ~n19375;
  assign n19377 = ~controllable_hgrant1 & ~n19376;
  assign n19378 = ~n14023 & ~n19377;
  assign n19379 = ~i_hbusreq3 & ~n19378;
  assign n19380 = ~n19371 & ~n19379;
  assign n19381 = ~controllable_hgrant3 & ~n19380;
  assign n19382 = ~n14022 & ~n19381;
  assign n19383 = i_hlock9 & ~n19382;
  assign n19384 = i_hbusreq3 & ~n19192;
  assign n19385 = i_hbusreq1 & ~n19190;
  assign n19386 = ~n16216 & ~n19373;
  assign n19387 = ~i_hbusreq1 & ~n19386;
  assign n19388 = ~n19385 & ~n19387;
  assign n19389 = ~controllable_hgrant1 & ~n19388;
  assign n19390 = ~n14058 & ~n19389;
  assign n19391 = ~i_hbusreq3 & ~n19390;
  assign n19392 = ~n19384 & ~n19391;
  assign n19393 = ~controllable_hgrant3 & ~n19392;
  assign n19394 = ~n14057 & ~n19393;
  assign n19395 = ~i_hlock9 & ~n19394;
  assign n19396 = ~n19383 & ~n19395;
  assign n19397 = ~i_hbusreq9 & ~n19396;
  assign n19398 = ~n19370 & ~n19397;
  assign n19399 = ~i_hbusreq4 & ~n19398;
  assign n19400 = ~n19369 & ~n19399;
  assign n19401 = ~controllable_hgrant4 & ~n19400;
  assign n19402 = ~n14322 & ~n19401;
  assign n19403 = ~i_hbusreq5 & ~n19402;
  assign n19404 = ~n19368 & ~n19403;
  assign n19405 = ~controllable_hgrant5 & ~n19404;
  assign n19406 = ~n14321 & ~n19405;
  assign n19407 = ~controllable_hmaster2 & ~n19406;
  assign n19408 = ~n19367 & ~n19407;
  assign n19409 = ~controllable_hmaster1 & ~n19408;
  assign n19410 = ~n19366 & ~n19409;
  assign n19411 = ~i_hbusreq6 & ~n19410;
  assign n19412 = ~n19342 & ~n19411;
  assign n19413 = ~controllable_hgrant6 & ~n19412;
  assign n19414 = ~n14320 & ~n19413;
  assign n19415 = controllable_hmaster0 & ~n19414;
  assign n19416 = i_hbusreq6 & ~n19210;
  assign n19417 = ~n16837 & ~n19367;
  assign n19418 = ~controllable_hmaster1 & ~n19417;
  assign n19419 = ~n19366 & ~n19418;
  assign n19420 = ~i_hbusreq6 & ~n19419;
  assign n19421 = ~n19416 & ~n19420;
  assign n19422 = ~controllable_hgrant6 & ~n19421;
  assign n19423 = ~n14443 & ~n19422;
  assign n19424 = ~controllable_hmaster0 & ~n19423;
  assign n19425 = ~n19415 & ~n19424;
  assign n19426 = i_hlock8 & ~n19425;
  assign n19427 = i_hbusreq6 & ~n19218;
  assign n19428 = ~n16874 & ~n19367;
  assign n19429 = ~controllable_hmaster1 & ~n19428;
  assign n19430 = ~n19366 & ~n19429;
  assign n19431 = ~i_hbusreq6 & ~n19430;
  assign n19432 = ~n19427 & ~n19431;
  assign n19433 = ~controllable_hgrant6 & ~n19432;
  assign n19434 = ~n14484 & ~n19433;
  assign n19435 = ~controllable_hmaster0 & ~n19434;
  assign n19436 = ~n19415 & ~n19435;
  assign n19437 = ~i_hlock8 & ~n19436;
  assign n19438 = ~n19426 & ~n19437;
  assign n19439 = ~i_hbusreq8 & ~n19438;
  assign n19440 = ~n19341 & ~n19439;
  assign n19441 = controllable_hmaster3 & ~n19440;
  assign n19442 = i_hbusreq8 & ~n19325;
  assign n19443 = i_hbusreq6 & ~n19276;
  assign n19444 = i_hbusreq5 & ~n19233;
  assign n19445 = i_hbusreq4 & ~n19231;
  assign n19446 = i_hbusreq9 & ~n19231;
  assign n19447 = i_hbusreq3 & ~n19229;
  assign n19448 = i_hbusreq1 & ~n19227;
  assign n19449 = n7928 & ~n16797;
  assign n19450 = ~n8265 & ~n19449;
  assign n19451 = ~i_hbusreq1 & ~n19450;
  assign n19452 = ~n19448 & ~n19451;
  assign n19453 = ~controllable_hgrant1 & ~n19452;
  assign n19454 = ~n14023 & ~n19453;
  assign n19455 = ~i_hbusreq3 & ~n19454;
  assign n19456 = ~n19447 & ~n19455;
  assign n19457 = ~controllable_hgrant3 & ~n19456;
  assign n19458 = ~n14022 & ~n19457;
  assign n19459 = ~i_hbusreq9 & ~n19458;
  assign n19460 = ~n19446 & ~n19459;
  assign n19461 = ~i_hbusreq4 & ~n19460;
  assign n19462 = ~n19445 & ~n19461;
  assign n19463 = ~controllable_hgrant4 & ~n19462;
  assign n19464 = ~n14021 & ~n19463;
  assign n19465 = ~i_hbusreq5 & ~n19464;
  assign n19466 = ~n19444 & ~n19465;
  assign n19467 = ~controllable_hgrant5 & ~n19466;
  assign n19468 = ~n14020 & ~n19467;
  assign n19469 = controllable_hmaster2 & ~n19468;
  assign n19470 = i_hbusreq5 & ~n19246;
  assign n19471 = i_hbusreq4 & ~n19244;
  assign n19472 = i_hbusreq9 & ~n19244;
  assign n19473 = i_hbusreq3 & ~n19242;
  assign n19474 = i_hlock3 & ~n19454;
  assign n19475 = i_hbusreq1 & ~n19238;
  assign n19476 = ~n8297 & ~n19449;
  assign n19477 = ~i_hbusreq1 & ~n19476;
  assign n19478 = ~n19475 & ~n19477;
  assign n19479 = ~controllable_hgrant1 & ~n19478;
  assign n19480 = ~n14058 & ~n19479;
  assign n19481 = ~i_hlock3 & ~n19480;
  assign n19482 = ~n19474 & ~n19481;
  assign n19483 = ~i_hbusreq3 & ~n19482;
  assign n19484 = ~n19473 & ~n19483;
  assign n19485 = ~controllable_hgrant3 & ~n19484;
  assign n19486 = ~n14102 & ~n19485;
  assign n19487 = ~i_hbusreq9 & ~n19486;
  assign n19488 = ~n19472 & ~n19487;
  assign n19489 = ~i_hbusreq4 & ~n19488;
  assign n19490 = ~n19471 & ~n19489;
  assign n19491 = ~controllable_hgrant4 & ~n19490;
  assign n19492 = ~n14099 & ~n19491;
  assign n19493 = ~i_hbusreq5 & ~n19492;
  assign n19494 = ~n19470 & ~n19493;
  assign n19495 = ~controllable_hgrant5 & ~n19494;
  assign n19496 = ~n14097 & ~n19495;
  assign n19497 = ~controllable_hmaster2 & ~n19496;
  assign n19498 = ~n19469 & ~n19497;
  assign n19499 = controllable_hmaster1 & ~n19498;
  assign n19500 = i_hbusreq5 & ~n19258;
  assign n19501 = i_hlock5 & ~n19464;
  assign n19502 = i_hbusreq4 & ~n19254;
  assign n19503 = i_hbusreq9 & ~n19254;
  assign n19504 = i_hbusreq3 & ~n19240;
  assign n19505 = ~i_hbusreq3 & ~n19480;
  assign n19506 = ~n19504 & ~n19505;
  assign n19507 = ~controllable_hgrant3 & ~n19506;
  assign n19508 = ~n14057 & ~n19507;
  assign n19509 = ~i_hbusreq9 & ~n19508;
  assign n19510 = ~n19503 & ~n19509;
  assign n19511 = ~i_hbusreq4 & ~n19510;
  assign n19512 = ~n19502 & ~n19511;
  assign n19513 = ~controllable_hgrant4 & ~n19512;
  assign n19514 = ~n14056 & ~n19513;
  assign n19515 = ~i_hlock5 & ~n19514;
  assign n19516 = ~n19501 & ~n19515;
  assign n19517 = ~i_hbusreq5 & ~n19516;
  assign n19518 = ~n19500 & ~n19517;
  assign n19519 = ~controllable_hgrant5 & ~n19518;
  assign n19520 = ~n14124 & ~n19519;
  assign n19521 = controllable_hmaster2 & ~n19520;
  assign n19522 = i_hbusreq5 & ~n19270;
  assign n19523 = i_hbusreq4 & ~n19268;
  assign n19524 = i_hbusreq9 & ~n19268;
  assign n19525 = i_hbusreq3 & ~n19266;
  assign n19526 = i_hbusreq1 & ~n19264;
  assign n19527 = i_hlock1 & ~n19450;
  assign n19528 = ~i_hlock1 & ~n19476;
  assign n19529 = ~n19527 & ~n19528;
  assign n19530 = ~i_hbusreq1 & ~n19529;
  assign n19531 = ~n19526 & ~n19530;
  assign n19532 = ~controllable_hgrant1 & ~n19531;
  assign n19533 = ~n14141 & ~n19532;
  assign n19534 = ~i_hbusreq3 & ~n19533;
  assign n19535 = ~n19525 & ~n19534;
  assign n19536 = ~controllable_hgrant3 & ~n19535;
  assign n19537 = ~n14139 & ~n19536;
  assign n19538 = ~i_hbusreq9 & ~n19537;
  assign n19539 = ~n19524 & ~n19538;
  assign n19540 = ~i_hbusreq4 & ~n19539;
  assign n19541 = ~n19523 & ~n19540;
  assign n19542 = ~controllable_hgrant4 & ~n19541;
  assign n19543 = ~n14136 & ~n19542;
  assign n19544 = ~i_hbusreq5 & ~n19543;
  assign n19545 = ~n19522 & ~n19544;
  assign n19546 = ~controllable_hgrant5 & ~n19545;
  assign n19547 = ~n14134 & ~n19546;
  assign n19548 = ~controllable_hmaster2 & ~n19547;
  assign n19549 = ~n19521 & ~n19548;
  assign n19550 = ~controllable_hmaster1 & ~n19549;
  assign n19551 = ~n19499 & ~n19550;
  assign n19552 = ~i_hbusreq6 & ~n19551;
  assign n19553 = ~n19443 & ~n19552;
  assign n19554 = ~controllable_hgrant6 & ~n19553;
  assign n19555 = ~n14094 & ~n19554;
  assign n19556 = controllable_hmaster0 & ~n19555;
  assign n19557 = i_hbusreq6 & ~n19321;
  assign n19558 = i_hbusreq5 & ~n19286;
  assign n19559 = i_hbusreq4 & ~n19284;
  assign n19560 = i_hbusreq9 & ~n19284;
  assign n19561 = i_hbusreq3 & ~n19282;
  assign n19562 = i_hbusreq1 & ~n19280;
  assign n19563 = ~n9379 & ~n19449;
  assign n19564 = ~i_hbusreq1 & ~n19563;
  assign n19565 = ~n19562 & ~n19564;
  assign n19566 = ~controllable_hgrant1 & ~n19565;
  assign n19567 = ~n14182 & ~n19566;
  assign n19568 = ~i_hbusreq3 & ~n19567;
  assign n19569 = ~n19561 & ~n19568;
  assign n19570 = ~controllable_hgrant3 & ~n19569;
  assign n19571 = ~n14180 & ~n19570;
  assign n19572 = ~i_hbusreq9 & ~n19571;
  assign n19573 = ~n19560 & ~n19572;
  assign n19574 = ~i_hbusreq4 & ~n19573;
  assign n19575 = ~n19559 & ~n19574;
  assign n19576 = ~controllable_hgrant4 & ~n19575;
  assign n19577 = ~n14177 & ~n19576;
  assign n19578 = ~i_hbusreq5 & ~n19577;
  assign n19579 = ~n19558 & ~n19578;
  assign n19580 = ~controllable_hgrant5 & ~n19579;
  assign n19581 = ~n14175 & ~n19580;
  assign n19582 = ~controllable_hmaster2 & ~n19581;
  assign n19583 = ~n19469 & ~n19582;
  assign n19584 = controllable_hmaster1 & ~n19583;
  assign n19585 = i_hbusreq5 & ~n19296;
  assign n19586 = i_hbusreq4 & ~n19294;
  assign n19587 = i_hlock4 & ~n19460;
  assign n19588 = ~i_hlock4 & ~n19510;
  assign n19589 = ~n19587 & ~n19588;
  assign n19590 = ~i_hbusreq4 & ~n19589;
  assign n19591 = ~n19586 & ~n19590;
  assign n19592 = ~controllable_hgrant4 & ~n19591;
  assign n19593 = ~n14208 & ~n19592;
  assign n19594 = ~i_hbusreq5 & ~n19593;
  assign n19595 = ~n19585 & ~n19594;
  assign n19596 = ~controllable_hgrant5 & ~n19595;
  assign n19597 = ~n14206 & ~n19596;
  assign n19598 = controllable_hmaster2 & ~n19597;
  assign n19599 = i_hbusreq5 & ~n19306;
  assign n19600 = i_hbusreq4 & ~n19304;
  assign n19601 = i_hbusreq9 & ~n19304;
  assign n19602 = i_hbusreq3 & ~n19302;
  assign n19603 = i_hbusreq1 & ~n19300;
  assign n19604 = n7928 & ~n18453;
  assign n19605 = ~n8440 & ~n19604;
  assign n19606 = ~i_hbusreq1 & ~n19605;
  assign n19607 = ~n19603 & ~n19606;
  assign n19608 = ~controllable_hgrant1 & ~n19607;
  assign n19609 = ~n14229 & ~n19608;
  assign n19610 = ~i_hbusreq3 & ~n19609;
  assign n19611 = ~n19602 & ~n19610;
  assign n19612 = ~controllable_hgrant3 & ~n19611;
  assign n19613 = ~n14227 & ~n19612;
  assign n19614 = ~i_hbusreq9 & ~n19613;
  assign n19615 = ~n19601 & ~n19614;
  assign n19616 = ~i_hbusreq4 & ~n19615;
  assign n19617 = ~n19600 & ~n19616;
  assign n19618 = ~controllable_hgrant4 & ~n19617;
  assign n19619 = ~n14224 & ~n19618;
  assign n19620 = ~i_hbusreq5 & ~n19619;
  assign n19621 = ~n19599 & ~n19620;
  assign n19622 = ~controllable_hgrant5 & ~n19621;
  assign n19623 = ~n14222 & ~n19622;
  assign n19624 = ~controllable_hmaster2 & ~n19623;
  assign n19625 = ~n19598 & ~n19624;
  assign n19626 = ~controllable_hmaster1 & ~n19625;
  assign n19627 = ~n19584 & ~n19626;
  assign n19628 = i_hlock6 & ~n19627;
  assign n19629 = i_hbusreq5 & ~n19256;
  assign n19630 = ~i_hbusreq5 & ~n19514;
  assign n19631 = ~n19629 & ~n19630;
  assign n19632 = ~controllable_hgrant5 & ~n19631;
  assign n19633 = ~n14055 & ~n19632;
  assign n19634 = controllable_hmaster2 & ~n19633;
  assign n19635 = ~n19582 & ~n19634;
  assign n19636 = controllable_hmaster1 & ~n19635;
  assign n19637 = ~n19626 & ~n19636;
  assign n19638 = ~i_hlock6 & ~n19637;
  assign n19639 = ~n19628 & ~n19638;
  assign n19640 = ~i_hbusreq6 & ~n19639;
  assign n19641 = ~n19557 & ~n19640;
  assign n19642 = ~controllable_hgrant6 & ~n19641;
  assign n19643 = ~n14173 & ~n19642;
  assign n19644 = ~controllable_hmaster0 & ~n19643;
  assign n19645 = ~n19556 & ~n19644;
  assign n19646 = ~i_hbusreq8 & ~n19645;
  assign n19647 = ~n19442 & ~n19646;
  assign n19648 = ~controllable_hmaster3 & ~n19647;
  assign n19649 = ~n19441 & ~n19648;
  assign n19650 = i_hlock7 & ~n19649;
  assign n19651 = i_hbusreq8 & ~n19335;
  assign n19652 = i_hbusreq6 & ~n19331;
  assign n19653 = ~n19497 & ~n19634;
  assign n19654 = controllable_hmaster1 & ~n19653;
  assign n19655 = ~n19550 & ~n19654;
  assign n19656 = ~i_hbusreq6 & ~n19655;
  assign n19657 = ~n19652 & ~n19656;
  assign n19658 = ~controllable_hgrant6 & ~n19657;
  assign n19659 = ~n14298 & ~n19658;
  assign n19660 = controllable_hmaster0 & ~n19659;
  assign n19661 = ~n19644 & ~n19660;
  assign n19662 = ~i_hbusreq8 & ~n19661;
  assign n19663 = ~n19651 & ~n19662;
  assign n19664 = ~controllable_hmaster3 & ~n19663;
  assign n19665 = ~n19441 & ~n19664;
  assign n19666 = ~i_hlock7 & ~n19665;
  assign n19667 = ~n19650 & ~n19666;
  assign n19668 = ~i_hbusreq7 & ~n19667;
  assign n19669 = ~n19340 & ~n19668;
  assign n19670 = ~n7924 & ~n19669;
  assign n19671 = ~n7928 & ~n16725;
  assign n19672 = n7928 & ~n17506;
  assign n19673 = ~n19671 & ~n19672;
  assign n19674 = ~controllable_hgrant1 & ~n19673;
  assign n19675 = ~n13155 & ~n19674;
  assign n19676 = ~controllable_hgrant3 & ~n19675;
  assign n19677 = ~n13154 & ~n19676;
  assign n19678 = ~controllable_hgrant4 & ~n19677;
  assign n19679 = ~n13153 & ~n19678;
  assign n19680 = ~controllable_hgrant5 & ~n19679;
  assign n19681 = ~n13152 & ~n19680;
  assign n19682 = controllable_hmaster1 & ~n19681;
  assign n19683 = controllable_hmaster2 & ~n19681;
  assign n19684 = n7928 & ~n16506;
  assign n19685 = ~n16128 & ~n19684;
  assign n19686 = ~controllable_hgrant1 & ~n19685;
  assign n19687 = ~n12611 & ~n19686;
  assign n19688 = ~controllable_hgrant3 & ~n19687;
  assign n19689 = ~n12610 & ~n19688;
  assign n19690 = i_hlock9 & ~n19689;
  assign n19691 = ~n16146 & ~n19684;
  assign n19692 = ~controllable_hgrant1 & ~n19691;
  assign n19693 = ~n12638 & ~n19692;
  assign n19694 = ~controllable_hgrant3 & ~n19693;
  assign n19695 = ~n12637 & ~n19694;
  assign n19696 = ~i_hlock9 & ~n19695;
  assign n19697 = ~n19690 & ~n19696;
  assign n19698 = ~controllable_hgrant4 & ~n19697;
  assign n19699 = ~n12609 & ~n19698;
  assign n19700 = ~controllable_hgrant5 & ~n19699;
  assign n19701 = ~n12608 & ~n19700;
  assign n19702 = ~controllable_hmaster2 & ~n19701;
  assign n19703 = ~n19683 & ~n19702;
  assign n19704 = ~controllable_hmaster1 & ~n19703;
  assign n19705 = ~n19682 & ~n19704;
  assign n19706 = ~controllable_hgrant6 & ~n19705;
  assign n19707 = ~n13122 & ~n19706;
  assign n19708 = controllable_hmaster0 & ~n19707;
  assign n19709 = ~controllable_hgrant2 & n16729;
  assign n19710 = ~n7814 & ~n19709;
  assign n19711 = n7733 & ~n19710;
  assign n19712 = ~n17507 & ~n19711;
  assign n19713 = n7928 & ~n19712;
  assign n19714 = ~n8221 & ~n19713;
  assign n19715 = ~controllable_hgrant1 & ~n19714;
  assign n19716 = ~n12611 & ~n19715;
  assign n19717 = ~controllable_hgrant3 & ~n19716;
  assign n19718 = ~n12610 & ~n19717;
  assign n19719 = ~controllable_hgrant4 & ~n19718;
  assign n19720 = ~n13408 & ~n19719;
  assign n19721 = ~controllable_hgrant5 & ~n19720;
  assign n19722 = ~n13407 & ~n19721;
  assign n19723 = ~controllable_hmaster2 & ~n19722;
  assign n19724 = ~n19683 & ~n19723;
  assign n19725 = ~controllable_hmaster1 & ~n19724;
  assign n19726 = ~n19682 & ~n19725;
  assign n19727 = ~controllable_hgrant6 & ~n19726;
  assign n19728 = ~n13406 & ~n19727;
  assign n19729 = ~controllable_hmaster0 & ~n19728;
  assign n19730 = ~n19708 & ~n19729;
  assign n19731 = i_hlock8 & ~n19730;
  assign n19732 = ~n8235 & ~n19713;
  assign n19733 = ~controllable_hgrant1 & ~n19732;
  assign n19734 = ~n12638 & ~n19733;
  assign n19735 = ~controllable_hgrant3 & ~n19734;
  assign n19736 = ~n12637 & ~n19735;
  assign n19737 = ~controllable_hgrant4 & ~n19736;
  assign n19738 = ~n13429 & ~n19737;
  assign n19739 = ~controllable_hgrant5 & ~n19738;
  assign n19740 = ~n13428 & ~n19739;
  assign n19741 = ~controllable_hmaster2 & ~n19740;
  assign n19742 = ~n19683 & ~n19741;
  assign n19743 = ~controllable_hmaster1 & ~n19742;
  assign n19744 = ~n19682 & ~n19743;
  assign n19745 = ~controllable_hgrant6 & ~n19744;
  assign n19746 = ~n13427 & ~n19745;
  assign n19747 = ~controllable_hmaster0 & ~n19746;
  assign n19748 = ~n19708 & ~n19747;
  assign n19749 = ~i_hlock8 & ~n19748;
  assign n19750 = ~n19731 & ~n19749;
  assign n19751 = controllable_hmaster3 & ~n19750;
  assign n19752 = ~n8221 & ~n19672;
  assign n19753 = ~controllable_hgrant1 & ~n19752;
  assign n19754 = ~n12611 & ~n19753;
  assign n19755 = ~controllable_hgrant3 & ~n19754;
  assign n19756 = ~n12610 & ~n19755;
  assign n19757 = ~controllable_hgrant4 & ~n19756;
  assign n19758 = ~n13408 & ~n19757;
  assign n19759 = ~controllable_hgrant5 & ~n19758;
  assign n19760 = ~n13407 & ~n19759;
  assign n19761 = controllable_hmaster2 & ~n19760;
  assign n19762 = i_hlock3 & ~n19754;
  assign n19763 = ~n8235 & ~n19672;
  assign n19764 = ~controllable_hgrant1 & ~n19763;
  assign n19765 = ~n12638 & ~n19764;
  assign n19766 = ~i_hlock3 & ~n19765;
  assign n19767 = ~n19762 & ~n19766;
  assign n19768 = ~controllable_hgrant3 & ~n19767;
  assign n19769 = ~n13852 & ~n19768;
  assign n19770 = ~controllable_hgrant4 & ~n19769;
  assign n19771 = ~n13851 & ~n19770;
  assign n19772 = ~controllable_hgrant5 & ~n19771;
  assign n19773 = ~n13850 & ~n19772;
  assign n19774 = ~controllable_hmaster2 & ~n19773;
  assign n19775 = ~n19761 & ~n19774;
  assign n19776 = controllable_hmaster1 & ~n19775;
  assign n19777 = i_hlock5 & ~n19758;
  assign n19778 = ~controllable_hgrant3 & ~n19765;
  assign n19779 = ~n12637 & ~n19778;
  assign n19780 = ~controllable_hgrant4 & ~n19779;
  assign n19781 = ~n13429 & ~n19780;
  assign n19782 = ~i_hlock5 & ~n19781;
  assign n19783 = ~n19777 & ~n19782;
  assign n19784 = ~controllable_hgrant5 & ~n19783;
  assign n19785 = ~n13865 & ~n19784;
  assign n19786 = controllable_hmaster2 & ~n19785;
  assign n19787 = i_hlock1 & ~n19752;
  assign n19788 = ~i_hlock1 & ~n19763;
  assign n19789 = ~n19787 & ~n19788;
  assign n19790 = ~controllable_hgrant1 & ~n19789;
  assign n19791 = ~n13875 & ~n19790;
  assign n19792 = ~controllable_hgrant3 & ~n19791;
  assign n19793 = ~n13874 & ~n19792;
  assign n19794 = ~controllable_hgrant4 & ~n19793;
  assign n19795 = ~n13873 & ~n19794;
  assign n19796 = ~controllable_hgrant5 & ~n19795;
  assign n19797 = ~n13872 & ~n19796;
  assign n19798 = ~controllable_hmaster2 & ~n19797;
  assign n19799 = ~n19786 & ~n19798;
  assign n19800 = ~controllable_hmaster1 & ~n19799;
  assign n19801 = ~n19776 & ~n19800;
  assign n19802 = ~controllable_hgrant6 & ~n19801;
  assign n19803 = ~n13849 & ~n19802;
  assign n19804 = controllable_hmaster0 & ~n19803;
  assign n19805 = ~n9213 & ~n19672;
  assign n19806 = ~controllable_hgrant1 & ~n19805;
  assign n19807 = ~n13898 & ~n19806;
  assign n19808 = ~controllable_hgrant3 & ~n19807;
  assign n19809 = ~n13897 & ~n19808;
  assign n19810 = ~controllable_hgrant4 & ~n19809;
  assign n19811 = ~n13896 & ~n19810;
  assign n19812 = ~controllable_hgrant5 & ~n19811;
  assign n19813 = ~n13895 & ~n19812;
  assign n19814 = ~controllable_hmaster2 & ~n19813;
  assign n19815 = ~n19761 & ~n19814;
  assign n19816 = controllable_hmaster1 & ~n19815;
  assign n19817 = i_hlock4 & ~n19756;
  assign n19818 = ~i_hlock4 & ~n19779;
  assign n19819 = ~n19817 & ~n19818;
  assign n19820 = ~controllable_hgrant4 & ~n19819;
  assign n19821 = ~n13912 & ~n19820;
  assign n19822 = ~controllable_hgrant5 & ~n19821;
  assign n19823 = ~n13911 & ~n19822;
  assign n19824 = controllable_hmaster2 & ~n19823;
  assign n19825 = ~n8440 & ~n19672;
  assign n19826 = ~controllable_hgrant1 & ~n19825;
  assign n19827 = ~n13924 & ~n19826;
  assign n19828 = ~controllable_hgrant3 & ~n19827;
  assign n19829 = ~n13923 & ~n19828;
  assign n19830 = ~controllable_hgrant4 & ~n19829;
  assign n19831 = ~n13922 & ~n19830;
  assign n19832 = ~controllable_hgrant5 & ~n19831;
  assign n19833 = ~n13921 & ~n19832;
  assign n19834 = ~controllable_hmaster2 & ~n19833;
  assign n19835 = ~n19824 & ~n19834;
  assign n19836 = ~controllable_hmaster1 & ~n19835;
  assign n19837 = ~n19816 & ~n19836;
  assign n19838 = i_hlock6 & ~n19837;
  assign n19839 = ~controllable_hgrant5 & ~n19781;
  assign n19840 = ~n13428 & ~n19839;
  assign n19841 = controllable_hmaster2 & ~n19840;
  assign n19842 = ~n19814 & ~n19841;
  assign n19843 = controllable_hmaster1 & ~n19842;
  assign n19844 = ~n19836 & ~n19843;
  assign n19845 = ~i_hlock6 & ~n19844;
  assign n19846 = ~n19838 & ~n19845;
  assign n19847 = ~controllable_hgrant6 & ~n19846;
  assign n19848 = ~n13894 & ~n19847;
  assign n19849 = ~controllable_hmaster0 & ~n19848;
  assign n19850 = ~n19804 & ~n19849;
  assign n19851 = ~controllable_hmaster3 & ~n19850;
  assign n19852 = ~n19751 & ~n19851;
  assign n19853 = i_hlock7 & ~n19852;
  assign n19854 = ~n19774 & ~n19841;
  assign n19855 = controllable_hmaster1 & ~n19854;
  assign n19856 = ~n19800 & ~n19855;
  assign n19857 = ~controllable_hgrant6 & ~n19856;
  assign n19858 = ~n13951 & ~n19857;
  assign n19859 = controllable_hmaster0 & ~n19858;
  assign n19860 = ~n19849 & ~n19859;
  assign n19861 = ~controllable_hmaster3 & ~n19860;
  assign n19862 = ~n19751 & ~n19861;
  assign n19863 = ~i_hlock7 & ~n19862;
  assign n19864 = ~n19853 & ~n19863;
  assign n19865 = i_hbusreq7 & ~n19864;
  assign n19866 = i_hbusreq8 & ~n19750;
  assign n19867 = i_hbusreq6 & ~n19705;
  assign n19868 = i_hbusreq5 & ~n19679;
  assign n19869 = i_hbusreq4 & ~n19677;
  assign n19870 = i_hbusreq9 & ~n19677;
  assign n19871 = i_hbusreq3 & ~n19675;
  assign n19872 = i_hbusreq1 & ~n19673;
  assign n19873 = ~n7928 & ~n16797;
  assign n19874 = n7928 & ~n18799;
  assign n19875 = ~n19873 & ~n19874;
  assign n19876 = ~i_hbusreq1 & ~n19875;
  assign n19877 = ~n19872 & ~n19876;
  assign n19878 = ~controllable_hgrant1 & ~n19877;
  assign n19879 = ~n13968 & ~n19878;
  assign n19880 = ~i_hbusreq3 & ~n19879;
  assign n19881 = ~n19871 & ~n19880;
  assign n19882 = ~controllable_hgrant3 & ~n19881;
  assign n19883 = ~n13967 & ~n19882;
  assign n19884 = ~i_hbusreq9 & ~n19883;
  assign n19885 = ~n19870 & ~n19884;
  assign n19886 = ~i_hbusreq4 & ~n19885;
  assign n19887 = ~n19869 & ~n19886;
  assign n19888 = ~controllable_hgrant4 & ~n19887;
  assign n19889 = ~n13966 & ~n19888;
  assign n19890 = ~i_hbusreq5 & ~n19889;
  assign n19891 = ~n19868 & ~n19890;
  assign n19892 = ~controllable_hgrant5 & ~n19891;
  assign n19893 = ~n13965 & ~n19892;
  assign n19894 = controllable_hmaster1 & ~n19893;
  assign n19895 = controllable_hmaster2 & ~n19893;
  assign n19896 = i_hbusreq5 & ~n19699;
  assign n19897 = i_hbusreq4 & ~n19697;
  assign n19898 = i_hbusreq9 & ~n19697;
  assign n19899 = i_hbusreq3 & ~n19687;
  assign n19900 = i_hbusreq1 & ~n19685;
  assign n19901 = n7928 & ~n16634;
  assign n19902 = ~n16191 & ~n19901;
  assign n19903 = ~i_hbusreq1 & ~n19902;
  assign n19904 = ~n19900 & ~n19903;
  assign n19905 = ~controllable_hgrant1 & ~n19904;
  assign n19906 = ~n14023 & ~n19905;
  assign n19907 = ~i_hbusreq3 & ~n19906;
  assign n19908 = ~n19899 & ~n19907;
  assign n19909 = ~controllable_hgrant3 & ~n19908;
  assign n19910 = ~n14022 & ~n19909;
  assign n19911 = i_hlock9 & ~n19910;
  assign n19912 = i_hbusreq3 & ~n19693;
  assign n19913 = i_hbusreq1 & ~n19691;
  assign n19914 = ~n16216 & ~n19901;
  assign n19915 = ~i_hbusreq1 & ~n19914;
  assign n19916 = ~n19913 & ~n19915;
  assign n19917 = ~controllable_hgrant1 & ~n19916;
  assign n19918 = ~n14058 & ~n19917;
  assign n19919 = ~i_hbusreq3 & ~n19918;
  assign n19920 = ~n19912 & ~n19919;
  assign n19921 = ~controllable_hgrant3 & ~n19920;
  assign n19922 = ~n14057 & ~n19921;
  assign n19923 = ~i_hlock9 & ~n19922;
  assign n19924 = ~n19911 & ~n19923;
  assign n19925 = ~i_hbusreq9 & ~n19924;
  assign n19926 = ~n19898 & ~n19925;
  assign n19927 = ~i_hbusreq4 & ~n19926;
  assign n19928 = ~n19897 & ~n19927;
  assign n19929 = ~controllable_hgrant4 & ~n19928;
  assign n19930 = ~n14322 & ~n19929;
  assign n19931 = ~i_hbusreq5 & ~n19930;
  assign n19932 = ~n19896 & ~n19931;
  assign n19933 = ~controllable_hgrant5 & ~n19932;
  assign n19934 = ~n14321 & ~n19933;
  assign n19935 = ~controllable_hmaster2 & ~n19934;
  assign n19936 = ~n19895 & ~n19935;
  assign n19937 = ~controllable_hmaster1 & ~n19936;
  assign n19938 = ~n19894 & ~n19937;
  assign n19939 = ~i_hbusreq6 & ~n19938;
  assign n19940 = ~n19867 & ~n19939;
  assign n19941 = ~controllable_hgrant6 & ~n19940;
  assign n19942 = ~n14320 & ~n19941;
  assign n19943 = controllable_hmaster0 & ~n19942;
  assign n19944 = i_hbusreq6 & ~n19726;
  assign n19945 = i_hbusreq5 & ~n19720;
  assign n19946 = i_hbusreq4 & ~n19718;
  assign n19947 = i_hbusreq9 & ~n19718;
  assign n19948 = i_hbusreq3 & ~n19716;
  assign n19949 = i_hbusreq1 & ~n19714;
  assign n19950 = i_hbusreq2 & n16729;
  assign n19951 = i_hbusreq0 & n16729;
  assign n19952 = ~controllable_locked & n14242;
  assign n19953 = ~n16802 & ~n19952;
  assign n19954 = i_hlock0 & ~n19953;
  assign n19955 = ~i_hlock0 & n16729;
  assign n19956 = ~n19954 & ~n19955;
  assign n19957 = ~i_hbusreq0 & ~n19956;
  assign n19958 = ~n19951 & ~n19957;
  assign n19959 = ~i_hbusreq2 & ~n19958;
  assign n19960 = ~n19950 & ~n19959;
  assign n19961 = ~controllable_hgrant2 & ~n19960;
  assign n19962 = ~n12706 & ~n19961;
  assign n19963 = n7733 & ~n19962;
  assign n19964 = ~n18800 & ~n19963;
  assign n19965 = n7928 & ~n19964;
  assign n19966 = ~n8265 & ~n19965;
  assign n19967 = ~i_hbusreq1 & ~n19966;
  assign n19968 = ~n19949 & ~n19967;
  assign n19969 = ~controllable_hgrant1 & ~n19968;
  assign n19970 = ~n12681 & ~n19969;
  assign n19971 = ~i_hbusreq3 & ~n19970;
  assign n19972 = ~n19948 & ~n19971;
  assign n19973 = ~controllable_hgrant3 & ~n19972;
  assign n19974 = ~n12679 & ~n19973;
  assign n19975 = ~i_hbusreq9 & ~n19974;
  assign n19976 = ~n19947 & ~n19975;
  assign n19977 = ~i_hbusreq4 & ~n19976;
  assign n19978 = ~n19946 & ~n19977;
  assign n19979 = ~controllable_hgrant4 & ~n19978;
  assign n19980 = ~n13524 & ~n19979;
  assign n19981 = ~i_hbusreq5 & ~n19980;
  assign n19982 = ~n19945 & ~n19981;
  assign n19983 = ~controllable_hgrant5 & ~n19982;
  assign n19984 = ~n13522 & ~n19983;
  assign n19985 = ~controllable_hmaster2 & ~n19984;
  assign n19986 = ~n19895 & ~n19985;
  assign n19987 = ~controllable_hmaster1 & ~n19986;
  assign n19988 = ~n19894 & ~n19987;
  assign n19989 = ~i_hbusreq6 & ~n19988;
  assign n19990 = ~n19944 & ~n19989;
  assign n19991 = ~controllable_hgrant6 & ~n19990;
  assign n19992 = ~n14443 & ~n19991;
  assign n19993 = ~controllable_hmaster0 & ~n19992;
  assign n19994 = ~n19943 & ~n19993;
  assign n19995 = i_hlock8 & ~n19994;
  assign n19996 = i_hbusreq6 & ~n19744;
  assign n19997 = i_hbusreq5 & ~n19738;
  assign n19998 = i_hbusreq4 & ~n19736;
  assign n19999 = i_hbusreq9 & ~n19736;
  assign n20000 = i_hbusreq3 & ~n19734;
  assign n20001 = i_hbusreq1 & ~n19732;
  assign n20002 = ~n8297 & ~n19965;
  assign n20003 = ~i_hbusreq1 & ~n20002;
  assign n20004 = ~n20001 & ~n20003;
  assign n20005 = ~controllable_hgrant1 & ~n20004;
  assign n20006 = ~n12730 & ~n20005;
  assign n20007 = ~i_hbusreq3 & ~n20006;
  assign n20008 = ~n20000 & ~n20007;
  assign n20009 = ~controllable_hgrant3 & ~n20008;
  assign n20010 = ~n12728 & ~n20009;
  assign n20011 = ~i_hbusreq9 & ~n20010;
  assign n20012 = ~n19999 & ~n20011;
  assign n20013 = ~i_hbusreq4 & ~n20012;
  assign n20014 = ~n19998 & ~n20013;
  assign n20015 = ~controllable_hgrant4 & ~n20014;
  assign n20016 = ~n13577 & ~n20015;
  assign n20017 = ~i_hbusreq5 & ~n20016;
  assign n20018 = ~n19997 & ~n20017;
  assign n20019 = ~controllable_hgrant5 & ~n20018;
  assign n20020 = ~n13575 & ~n20019;
  assign n20021 = ~controllable_hmaster2 & ~n20020;
  assign n20022 = ~n19895 & ~n20021;
  assign n20023 = ~controllable_hmaster1 & ~n20022;
  assign n20024 = ~n19894 & ~n20023;
  assign n20025 = ~i_hbusreq6 & ~n20024;
  assign n20026 = ~n19996 & ~n20025;
  assign n20027 = ~controllable_hgrant6 & ~n20026;
  assign n20028 = ~n14484 & ~n20027;
  assign n20029 = ~controllable_hmaster0 & ~n20028;
  assign n20030 = ~n19943 & ~n20029;
  assign n20031 = ~i_hlock8 & ~n20030;
  assign n20032 = ~n19995 & ~n20031;
  assign n20033 = ~i_hbusreq8 & ~n20032;
  assign n20034 = ~n19866 & ~n20033;
  assign n20035 = controllable_hmaster3 & ~n20034;
  assign n20036 = i_hbusreq8 & ~n19850;
  assign n20037 = i_hbusreq6 & ~n19801;
  assign n20038 = i_hbusreq5 & ~n19758;
  assign n20039 = i_hbusreq4 & ~n19756;
  assign n20040 = i_hbusreq9 & ~n19756;
  assign n20041 = i_hbusreq3 & ~n19754;
  assign n20042 = i_hbusreq1 & ~n19752;
  assign n20043 = ~n8265 & ~n19874;
  assign n20044 = ~i_hbusreq1 & ~n20043;
  assign n20045 = ~n20042 & ~n20044;
  assign n20046 = ~controllable_hgrant1 & ~n20045;
  assign n20047 = ~n14023 & ~n20046;
  assign n20048 = ~i_hbusreq3 & ~n20047;
  assign n20049 = ~n20041 & ~n20048;
  assign n20050 = ~controllable_hgrant3 & ~n20049;
  assign n20051 = ~n14022 & ~n20050;
  assign n20052 = ~i_hbusreq9 & ~n20051;
  assign n20053 = ~n20040 & ~n20052;
  assign n20054 = ~i_hbusreq4 & ~n20053;
  assign n20055 = ~n20039 & ~n20054;
  assign n20056 = ~controllable_hgrant4 & ~n20055;
  assign n20057 = ~n14021 & ~n20056;
  assign n20058 = ~i_hbusreq5 & ~n20057;
  assign n20059 = ~n20038 & ~n20058;
  assign n20060 = ~controllable_hgrant5 & ~n20059;
  assign n20061 = ~n14020 & ~n20060;
  assign n20062 = controllable_hmaster2 & ~n20061;
  assign n20063 = i_hbusreq5 & ~n19771;
  assign n20064 = i_hbusreq4 & ~n19769;
  assign n20065 = i_hbusreq9 & ~n19769;
  assign n20066 = i_hbusreq3 & ~n19767;
  assign n20067 = i_hlock3 & ~n20047;
  assign n20068 = i_hbusreq1 & ~n19763;
  assign n20069 = ~n8297 & ~n19874;
  assign n20070 = ~i_hbusreq1 & ~n20069;
  assign n20071 = ~n20068 & ~n20070;
  assign n20072 = ~controllable_hgrant1 & ~n20071;
  assign n20073 = ~n14058 & ~n20072;
  assign n20074 = ~i_hlock3 & ~n20073;
  assign n20075 = ~n20067 & ~n20074;
  assign n20076 = ~i_hbusreq3 & ~n20075;
  assign n20077 = ~n20066 & ~n20076;
  assign n20078 = ~controllable_hgrant3 & ~n20077;
  assign n20079 = ~n14102 & ~n20078;
  assign n20080 = ~i_hbusreq9 & ~n20079;
  assign n20081 = ~n20065 & ~n20080;
  assign n20082 = ~i_hbusreq4 & ~n20081;
  assign n20083 = ~n20064 & ~n20082;
  assign n20084 = ~controllable_hgrant4 & ~n20083;
  assign n20085 = ~n14099 & ~n20084;
  assign n20086 = ~i_hbusreq5 & ~n20085;
  assign n20087 = ~n20063 & ~n20086;
  assign n20088 = ~controllable_hgrant5 & ~n20087;
  assign n20089 = ~n14097 & ~n20088;
  assign n20090 = ~controllable_hmaster2 & ~n20089;
  assign n20091 = ~n20062 & ~n20090;
  assign n20092 = controllable_hmaster1 & ~n20091;
  assign n20093 = i_hbusreq5 & ~n19783;
  assign n20094 = i_hlock5 & ~n20057;
  assign n20095 = i_hbusreq4 & ~n19779;
  assign n20096 = i_hbusreq9 & ~n19779;
  assign n20097 = i_hbusreq3 & ~n19765;
  assign n20098 = ~i_hbusreq3 & ~n20073;
  assign n20099 = ~n20097 & ~n20098;
  assign n20100 = ~controllable_hgrant3 & ~n20099;
  assign n20101 = ~n14057 & ~n20100;
  assign n20102 = ~i_hbusreq9 & ~n20101;
  assign n20103 = ~n20096 & ~n20102;
  assign n20104 = ~i_hbusreq4 & ~n20103;
  assign n20105 = ~n20095 & ~n20104;
  assign n20106 = ~controllable_hgrant4 & ~n20105;
  assign n20107 = ~n14056 & ~n20106;
  assign n20108 = ~i_hlock5 & ~n20107;
  assign n20109 = ~n20094 & ~n20108;
  assign n20110 = ~i_hbusreq5 & ~n20109;
  assign n20111 = ~n20093 & ~n20110;
  assign n20112 = ~controllable_hgrant5 & ~n20111;
  assign n20113 = ~n14124 & ~n20112;
  assign n20114 = controllable_hmaster2 & ~n20113;
  assign n20115 = i_hbusreq5 & ~n19795;
  assign n20116 = i_hbusreq4 & ~n19793;
  assign n20117 = i_hbusreq9 & ~n19793;
  assign n20118 = i_hbusreq3 & ~n19791;
  assign n20119 = i_hbusreq1 & ~n19789;
  assign n20120 = i_hlock1 & ~n20043;
  assign n20121 = ~i_hlock1 & ~n20069;
  assign n20122 = ~n20120 & ~n20121;
  assign n20123 = ~i_hbusreq1 & ~n20122;
  assign n20124 = ~n20119 & ~n20123;
  assign n20125 = ~controllable_hgrant1 & ~n20124;
  assign n20126 = ~n14141 & ~n20125;
  assign n20127 = ~i_hbusreq3 & ~n20126;
  assign n20128 = ~n20118 & ~n20127;
  assign n20129 = ~controllable_hgrant3 & ~n20128;
  assign n20130 = ~n14139 & ~n20129;
  assign n20131 = ~i_hbusreq9 & ~n20130;
  assign n20132 = ~n20117 & ~n20131;
  assign n20133 = ~i_hbusreq4 & ~n20132;
  assign n20134 = ~n20116 & ~n20133;
  assign n20135 = ~controllable_hgrant4 & ~n20134;
  assign n20136 = ~n14136 & ~n20135;
  assign n20137 = ~i_hbusreq5 & ~n20136;
  assign n20138 = ~n20115 & ~n20137;
  assign n20139 = ~controllable_hgrant5 & ~n20138;
  assign n20140 = ~n14134 & ~n20139;
  assign n20141 = ~controllable_hmaster2 & ~n20140;
  assign n20142 = ~n20114 & ~n20141;
  assign n20143 = ~controllable_hmaster1 & ~n20142;
  assign n20144 = ~n20092 & ~n20143;
  assign n20145 = ~i_hbusreq6 & ~n20144;
  assign n20146 = ~n20037 & ~n20145;
  assign n20147 = ~controllable_hgrant6 & ~n20146;
  assign n20148 = ~n14094 & ~n20147;
  assign n20149 = controllable_hmaster0 & ~n20148;
  assign n20150 = i_hbusreq6 & ~n19846;
  assign n20151 = i_hbusreq5 & ~n19811;
  assign n20152 = i_hbusreq4 & ~n19809;
  assign n20153 = i_hbusreq9 & ~n19809;
  assign n20154 = i_hbusreq3 & ~n19807;
  assign n20155 = i_hbusreq1 & ~n19805;
  assign n20156 = ~n9379 & ~n19874;
  assign n20157 = ~i_hbusreq1 & ~n20156;
  assign n20158 = ~n20155 & ~n20157;
  assign n20159 = ~controllable_hgrant1 & ~n20158;
  assign n20160 = ~n14182 & ~n20159;
  assign n20161 = ~i_hbusreq3 & ~n20160;
  assign n20162 = ~n20154 & ~n20161;
  assign n20163 = ~controllable_hgrant3 & ~n20162;
  assign n20164 = ~n14180 & ~n20163;
  assign n20165 = ~i_hbusreq9 & ~n20164;
  assign n20166 = ~n20153 & ~n20165;
  assign n20167 = ~i_hbusreq4 & ~n20166;
  assign n20168 = ~n20152 & ~n20167;
  assign n20169 = ~controllable_hgrant4 & ~n20168;
  assign n20170 = ~n14177 & ~n20169;
  assign n20171 = ~i_hbusreq5 & ~n20170;
  assign n20172 = ~n20151 & ~n20171;
  assign n20173 = ~controllable_hgrant5 & ~n20172;
  assign n20174 = ~n14175 & ~n20173;
  assign n20175 = ~controllable_hmaster2 & ~n20174;
  assign n20176 = ~n20062 & ~n20175;
  assign n20177 = controllable_hmaster1 & ~n20176;
  assign n20178 = i_hbusreq5 & ~n19821;
  assign n20179 = i_hbusreq4 & ~n19819;
  assign n20180 = i_hlock4 & ~n20053;
  assign n20181 = ~i_hlock4 & ~n20103;
  assign n20182 = ~n20180 & ~n20181;
  assign n20183 = ~i_hbusreq4 & ~n20182;
  assign n20184 = ~n20179 & ~n20183;
  assign n20185 = ~controllable_hgrant4 & ~n20184;
  assign n20186 = ~n14208 & ~n20185;
  assign n20187 = ~i_hbusreq5 & ~n20186;
  assign n20188 = ~n20178 & ~n20187;
  assign n20189 = ~controllable_hgrant5 & ~n20188;
  assign n20190 = ~n14206 & ~n20189;
  assign n20191 = controllable_hmaster2 & ~n20190;
  assign n20192 = i_hbusreq5 & ~n19831;
  assign n20193 = i_hbusreq4 & ~n19829;
  assign n20194 = i_hbusreq9 & ~n19829;
  assign n20195 = i_hbusreq3 & ~n19827;
  assign n20196 = i_hbusreq1 & ~n19825;
  assign n20197 = n7928 & ~n19071;
  assign n20198 = ~n8440 & ~n20197;
  assign n20199 = ~i_hbusreq1 & ~n20198;
  assign n20200 = ~n20196 & ~n20199;
  assign n20201 = ~controllable_hgrant1 & ~n20200;
  assign n20202 = ~n14229 & ~n20201;
  assign n20203 = ~i_hbusreq3 & ~n20202;
  assign n20204 = ~n20195 & ~n20203;
  assign n20205 = ~controllable_hgrant3 & ~n20204;
  assign n20206 = ~n14227 & ~n20205;
  assign n20207 = ~i_hbusreq9 & ~n20206;
  assign n20208 = ~n20194 & ~n20207;
  assign n20209 = ~i_hbusreq4 & ~n20208;
  assign n20210 = ~n20193 & ~n20209;
  assign n20211 = ~controllable_hgrant4 & ~n20210;
  assign n20212 = ~n14224 & ~n20211;
  assign n20213 = ~i_hbusreq5 & ~n20212;
  assign n20214 = ~n20192 & ~n20213;
  assign n20215 = ~controllable_hgrant5 & ~n20214;
  assign n20216 = ~n14222 & ~n20215;
  assign n20217 = ~controllable_hmaster2 & ~n20216;
  assign n20218 = ~n20191 & ~n20217;
  assign n20219 = ~controllable_hmaster1 & ~n20218;
  assign n20220 = ~n20177 & ~n20219;
  assign n20221 = i_hlock6 & ~n20220;
  assign n20222 = i_hbusreq5 & ~n19781;
  assign n20223 = ~i_hbusreq5 & ~n20107;
  assign n20224 = ~n20222 & ~n20223;
  assign n20225 = ~controllable_hgrant5 & ~n20224;
  assign n20226 = ~n14055 & ~n20225;
  assign n20227 = controllable_hmaster2 & ~n20226;
  assign n20228 = ~n20175 & ~n20227;
  assign n20229 = controllable_hmaster1 & ~n20228;
  assign n20230 = ~n20219 & ~n20229;
  assign n20231 = ~i_hlock6 & ~n20230;
  assign n20232 = ~n20221 & ~n20231;
  assign n20233 = ~i_hbusreq6 & ~n20232;
  assign n20234 = ~n20150 & ~n20233;
  assign n20235 = ~controllable_hgrant6 & ~n20234;
  assign n20236 = ~n14173 & ~n20235;
  assign n20237 = ~controllable_hmaster0 & ~n20236;
  assign n20238 = ~n20149 & ~n20237;
  assign n20239 = ~i_hbusreq8 & ~n20238;
  assign n20240 = ~n20036 & ~n20239;
  assign n20241 = ~controllable_hmaster3 & ~n20240;
  assign n20242 = ~n20035 & ~n20241;
  assign n20243 = i_hlock7 & ~n20242;
  assign n20244 = i_hbusreq8 & ~n19860;
  assign n20245 = i_hbusreq6 & ~n19856;
  assign n20246 = ~n20090 & ~n20227;
  assign n20247 = controllable_hmaster1 & ~n20246;
  assign n20248 = ~n20143 & ~n20247;
  assign n20249 = ~i_hbusreq6 & ~n20248;
  assign n20250 = ~n20245 & ~n20249;
  assign n20251 = ~controllable_hgrant6 & ~n20250;
  assign n20252 = ~n14298 & ~n20251;
  assign n20253 = controllable_hmaster0 & ~n20252;
  assign n20254 = ~n20237 & ~n20253;
  assign n20255 = ~i_hbusreq8 & ~n20254;
  assign n20256 = ~n20244 & ~n20255;
  assign n20257 = ~controllable_hmaster3 & ~n20256;
  assign n20258 = ~n20035 & ~n20257;
  assign n20259 = ~i_hlock7 & ~n20258;
  assign n20260 = ~n20243 & ~n20259;
  assign n20261 = ~i_hbusreq7 & ~n20260;
  assign n20262 = ~n19865 & ~n20261;
  assign n20263 = n7924 & ~n20262;
  assign n20264 = ~n19670 & ~n20263;
  assign n20265 = n8214 & ~n20264;
  assign n20266 = ~n19172 & ~n20265;
  assign n20267 = ~n8202 & ~n20266;
  assign n20268 = ~controllable_hmaster2 & ~n19235;
  assign n20269 = ~n19182 & ~n20268;
  assign n20270 = ~controllable_hmaster1 & ~n20269;
  assign n20271 = ~n19181 & ~n20270;
  assign n20272 = ~controllable_hgrant6 & ~n20271;
  assign n20273 = ~n13406 & ~n20272;
  assign n20274 = ~controllable_hmaster0 & ~n20273;
  assign n20275 = ~n19207 & ~n20274;
  assign n20276 = i_hlock8 & ~n20275;
  assign n20277 = ~controllable_hmaster2 & ~n19315;
  assign n20278 = ~n19182 & ~n20277;
  assign n20279 = ~controllable_hmaster1 & ~n20278;
  assign n20280 = ~n19181 & ~n20279;
  assign n20281 = ~controllable_hgrant6 & ~n20280;
  assign n20282 = ~n13427 & ~n20281;
  assign n20283 = ~controllable_hmaster0 & ~n20282;
  assign n20284 = ~n19207 & ~n20283;
  assign n20285 = ~i_hlock8 & ~n20284;
  assign n20286 = ~n20276 & ~n20285;
  assign n20287 = controllable_hmaster3 & ~n20286;
  assign n20288 = ~n16896 & ~n19249;
  assign n20289 = controllable_hmaster1 & ~n20288;
  assign n20290 = ~n19275 & ~n20289;
  assign n20291 = ~controllable_hgrant6 & ~n20290;
  assign n20292 = ~n13849 & ~n20291;
  assign n20293 = controllable_hmaster0 & ~n20292;
  assign n20294 = ~n19324 & ~n20293;
  assign n20295 = ~controllable_hmaster3 & ~n20294;
  assign n20296 = ~n20287 & ~n20295;
  assign n20297 = i_hlock7 & ~n20296;
  assign n20298 = ~n16908 & ~n19249;
  assign n20299 = controllable_hmaster1 & ~n20298;
  assign n20300 = ~n19275 & ~n20299;
  assign n20301 = ~controllable_hgrant6 & ~n20300;
  assign n20302 = ~n13951 & ~n20301;
  assign n20303 = controllable_hmaster0 & ~n20302;
  assign n20304 = ~n19324 & ~n20303;
  assign n20305 = ~controllable_hmaster3 & ~n20304;
  assign n20306 = ~n20287 & ~n20305;
  assign n20307 = ~i_hlock7 & ~n20306;
  assign n20308 = ~n20297 & ~n20307;
  assign n20309 = i_hbusreq7 & ~n20308;
  assign n20310 = i_hbusreq8 & ~n20286;
  assign n20311 = i_hbusreq6 & ~n20271;
  assign n20312 = ~controllable_hmaster2 & ~n19468;
  assign n20313 = ~n19367 & ~n20312;
  assign n20314 = ~controllable_hmaster1 & ~n20313;
  assign n20315 = ~n19366 & ~n20314;
  assign n20316 = ~i_hbusreq6 & ~n20315;
  assign n20317 = ~n20311 & ~n20316;
  assign n20318 = ~controllable_hgrant6 & ~n20317;
  assign n20319 = ~n14019 & ~n20318;
  assign n20320 = ~controllable_hmaster0 & ~n20319;
  assign n20321 = ~n19415 & ~n20320;
  assign n20322 = i_hlock8 & ~n20321;
  assign n20323 = i_hbusreq6 & ~n20280;
  assign n20324 = ~controllable_hmaster2 & ~n19633;
  assign n20325 = ~n19367 & ~n20324;
  assign n20326 = ~controllable_hmaster1 & ~n20325;
  assign n20327 = ~n19366 & ~n20326;
  assign n20328 = ~i_hbusreq6 & ~n20327;
  assign n20329 = ~n20323 & ~n20328;
  assign n20330 = ~controllable_hgrant6 & ~n20329;
  assign n20331 = ~n14054 & ~n20330;
  assign n20332 = ~controllable_hmaster0 & ~n20331;
  assign n20333 = ~n19415 & ~n20332;
  assign n20334 = ~i_hlock8 & ~n20333;
  assign n20335 = ~n20322 & ~n20334;
  assign n20336 = ~i_hbusreq8 & ~n20335;
  assign n20337 = ~n20310 & ~n20336;
  assign n20338 = controllable_hmaster3 & ~n20337;
  assign n20339 = i_hbusreq8 & ~n20294;
  assign n20340 = i_hbusreq6 & ~n20290;
  assign n20341 = ~n16924 & ~n19497;
  assign n20342 = controllable_hmaster1 & ~n20341;
  assign n20343 = ~n19550 & ~n20342;
  assign n20344 = ~i_hbusreq6 & ~n20343;
  assign n20345 = ~n20340 & ~n20344;
  assign n20346 = ~controllable_hgrant6 & ~n20345;
  assign n20347 = ~n14756 & ~n20346;
  assign n20348 = controllable_hmaster0 & ~n20347;
  assign n20349 = ~n19644 & ~n20348;
  assign n20350 = ~i_hbusreq8 & ~n20349;
  assign n20351 = ~n20339 & ~n20350;
  assign n20352 = ~controllable_hmaster3 & ~n20351;
  assign n20353 = ~n20338 & ~n20352;
  assign n20354 = i_hlock7 & ~n20353;
  assign n20355 = i_hbusreq8 & ~n20304;
  assign n20356 = i_hbusreq6 & ~n20300;
  assign n20357 = ~n16942 & ~n19497;
  assign n20358 = controllable_hmaster1 & ~n20357;
  assign n20359 = ~n19550 & ~n20358;
  assign n20360 = ~i_hbusreq6 & ~n20359;
  assign n20361 = ~n20356 & ~n20360;
  assign n20362 = ~controllable_hgrant6 & ~n20361;
  assign n20363 = ~n14772 & ~n20362;
  assign n20364 = controllable_hmaster0 & ~n20363;
  assign n20365 = ~n19644 & ~n20364;
  assign n20366 = ~i_hbusreq8 & ~n20365;
  assign n20367 = ~n20355 & ~n20366;
  assign n20368 = ~controllable_hmaster3 & ~n20367;
  assign n20369 = ~n20338 & ~n20368;
  assign n20370 = ~i_hlock7 & ~n20369;
  assign n20371 = ~n20354 & ~n20370;
  assign n20372 = ~i_hbusreq7 & ~n20371;
  assign n20373 = ~n20309 & ~n20372;
  assign n20374 = ~n7924 & ~n20373;
  assign n20375 = ~controllable_hmaster2 & ~n19760;
  assign n20376 = ~n19683 & ~n20375;
  assign n20377 = ~controllable_hmaster1 & ~n20376;
  assign n20378 = ~n19682 & ~n20377;
  assign n20379 = ~controllable_hgrant6 & ~n20378;
  assign n20380 = ~n13406 & ~n20379;
  assign n20381 = ~controllable_hmaster0 & ~n20380;
  assign n20382 = ~n19708 & ~n20381;
  assign n20383 = i_hlock8 & ~n20382;
  assign n20384 = ~controllable_hmaster2 & ~n19840;
  assign n20385 = ~n19683 & ~n20384;
  assign n20386 = ~controllable_hmaster1 & ~n20385;
  assign n20387 = ~n19682 & ~n20386;
  assign n20388 = ~controllable_hgrant6 & ~n20387;
  assign n20389 = ~n13427 & ~n20388;
  assign n20390 = ~controllable_hmaster0 & ~n20389;
  assign n20391 = ~n19708 & ~n20390;
  assign n20392 = ~i_hlock8 & ~n20391;
  assign n20393 = ~n20383 & ~n20392;
  assign n20394 = controllable_hmaster3 & ~n20393;
  assign n20395 = controllable_hmaster2 & ~n19722;
  assign n20396 = ~n19774 & ~n20395;
  assign n20397 = controllable_hmaster1 & ~n20396;
  assign n20398 = ~n19800 & ~n20397;
  assign n20399 = ~controllable_hgrant6 & ~n20398;
  assign n20400 = ~n13849 & ~n20399;
  assign n20401 = controllable_hmaster0 & ~n20400;
  assign n20402 = ~n19849 & ~n20401;
  assign n20403 = ~controllable_hmaster3 & ~n20402;
  assign n20404 = ~n20394 & ~n20403;
  assign n20405 = i_hlock7 & ~n20404;
  assign n20406 = controllable_hmaster2 & ~n19740;
  assign n20407 = ~n19774 & ~n20406;
  assign n20408 = controllable_hmaster1 & ~n20407;
  assign n20409 = ~n19800 & ~n20408;
  assign n20410 = ~controllable_hgrant6 & ~n20409;
  assign n20411 = ~n13951 & ~n20410;
  assign n20412 = controllable_hmaster0 & ~n20411;
  assign n20413 = ~n19849 & ~n20412;
  assign n20414 = ~controllable_hmaster3 & ~n20413;
  assign n20415 = ~n20394 & ~n20414;
  assign n20416 = ~i_hlock7 & ~n20415;
  assign n20417 = ~n20405 & ~n20416;
  assign n20418 = i_hbusreq7 & ~n20417;
  assign n20419 = i_hbusreq8 & ~n20393;
  assign n20420 = i_hbusreq6 & ~n20378;
  assign n20421 = ~controllable_hmaster2 & ~n20061;
  assign n20422 = ~n19895 & ~n20421;
  assign n20423 = ~controllable_hmaster1 & ~n20422;
  assign n20424 = ~n19894 & ~n20423;
  assign n20425 = ~i_hbusreq6 & ~n20424;
  assign n20426 = ~n20420 & ~n20425;
  assign n20427 = ~controllable_hgrant6 & ~n20426;
  assign n20428 = ~n14019 & ~n20427;
  assign n20429 = ~controllable_hmaster0 & ~n20428;
  assign n20430 = ~n19943 & ~n20429;
  assign n20431 = i_hlock8 & ~n20430;
  assign n20432 = i_hbusreq6 & ~n20387;
  assign n20433 = ~controllable_hmaster2 & ~n20226;
  assign n20434 = ~n19895 & ~n20433;
  assign n20435 = ~controllable_hmaster1 & ~n20434;
  assign n20436 = ~n19894 & ~n20435;
  assign n20437 = ~i_hbusreq6 & ~n20436;
  assign n20438 = ~n20432 & ~n20437;
  assign n20439 = ~controllable_hgrant6 & ~n20438;
  assign n20440 = ~n14054 & ~n20439;
  assign n20441 = ~controllable_hmaster0 & ~n20440;
  assign n20442 = ~n19943 & ~n20441;
  assign n20443 = ~i_hlock8 & ~n20442;
  assign n20444 = ~n20431 & ~n20443;
  assign n20445 = ~i_hbusreq8 & ~n20444;
  assign n20446 = ~n20419 & ~n20445;
  assign n20447 = controllable_hmaster3 & ~n20446;
  assign n20448 = i_hbusreq8 & ~n20402;
  assign n20449 = i_hbusreq6 & ~n20398;
  assign n20450 = controllable_hmaster2 & ~n19984;
  assign n20451 = ~n20090 & ~n20450;
  assign n20452 = controllable_hmaster1 & ~n20451;
  assign n20453 = ~n20143 & ~n20452;
  assign n20454 = ~i_hbusreq6 & ~n20453;
  assign n20455 = ~n20449 & ~n20454;
  assign n20456 = ~controllable_hgrant6 & ~n20455;
  assign n20457 = ~n14756 & ~n20456;
  assign n20458 = controllable_hmaster0 & ~n20457;
  assign n20459 = ~n20237 & ~n20458;
  assign n20460 = ~i_hbusreq8 & ~n20459;
  assign n20461 = ~n20448 & ~n20460;
  assign n20462 = ~controllable_hmaster3 & ~n20461;
  assign n20463 = ~n20447 & ~n20462;
  assign n20464 = i_hlock7 & ~n20463;
  assign n20465 = i_hbusreq8 & ~n20413;
  assign n20466 = i_hbusreq6 & ~n20409;
  assign n20467 = controllable_hmaster2 & ~n20020;
  assign n20468 = ~n20090 & ~n20467;
  assign n20469 = controllable_hmaster1 & ~n20468;
  assign n20470 = ~n20143 & ~n20469;
  assign n20471 = ~i_hbusreq6 & ~n20470;
  assign n20472 = ~n20466 & ~n20471;
  assign n20473 = ~controllable_hgrant6 & ~n20472;
  assign n20474 = ~n14772 & ~n20473;
  assign n20475 = controllable_hmaster0 & ~n20474;
  assign n20476 = ~n20237 & ~n20475;
  assign n20477 = ~i_hbusreq8 & ~n20476;
  assign n20478 = ~n20465 & ~n20477;
  assign n20479 = ~controllable_hmaster3 & ~n20478;
  assign n20480 = ~n20447 & ~n20479;
  assign n20481 = ~i_hlock7 & ~n20480;
  assign n20482 = ~n20464 & ~n20481;
  assign n20483 = ~i_hbusreq7 & ~n20482;
  assign n20484 = ~n20418 & ~n20483;
  assign n20485 = n7924 & ~n20484;
  assign n20486 = ~n20374 & ~n20485;
  assign n20487 = ~n8214 & ~n20486;
  assign n20488 = ~n16896 & ~n19289;
  assign n20489 = controllable_hmaster1 & ~n20488;
  assign n20490 = ~n19311 & ~n20489;
  assign n20491 = i_hlock6 & ~n20490;
  assign n20492 = ~n16908 & ~n19289;
  assign n20493 = controllable_hmaster1 & ~n20492;
  assign n20494 = ~n19311 & ~n20493;
  assign n20495 = ~i_hlock6 & ~n20494;
  assign n20496 = ~n20491 & ~n20495;
  assign n20497 = ~controllable_hgrant6 & ~n20496;
  assign n20498 = ~n13894 & ~n20497;
  assign n20499 = ~controllable_hmaster0 & ~n20498;
  assign n20500 = ~n19279 & ~n20499;
  assign n20501 = ~controllable_hmaster3 & ~n20500;
  assign n20502 = ~n20287 & ~n20501;
  assign n20503 = i_hlock7 & ~n20502;
  assign n20504 = ~n19334 & ~n20499;
  assign n20505 = ~controllable_hmaster3 & ~n20504;
  assign n20506 = ~n20287 & ~n20505;
  assign n20507 = ~i_hlock7 & ~n20506;
  assign n20508 = ~n20503 & ~n20507;
  assign n20509 = i_hbusreq7 & ~n20508;
  assign n20510 = i_hbusreq8 & ~n20500;
  assign n20511 = i_hbusreq6 & ~n20496;
  assign n20512 = ~n16924 & ~n19582;
  assign n20513 = controllable_hmaster1 & ~n20512;
  assign n20514 = ~n19626 & ~n20513;
  assign n20515 = i_hlock6 & ~n20514;
  assign n20516 = ~n16942 & ~n19582;
  assign n20517 = controllable_hmaster1 & ~n20516;
  assign n20518 = ~n19626 & ~n20517;
  assign n20519 = ~i_hlock6 & ~n20518;
  assign n20520 = ~n20515 & ~n20519;
  assign n20521 = ~i_hbusreq6 & ~n20520;
  assign n20522 = ~n20511 & ~n20521;
  assign n20523 = ~controllable_hgrant6 & ~n20522;
  assign n20524 = ~n14802 & ~n20523;
  assign n20525 = ~controllable_hmaster0 & ~n20524;
  assign n20526 = ~n19556 & ~n20525;
  assign n20527 = ~i_hbusreq8 & ~n20526;
  assign n20528 = ~n20510 & ~n20527;
  assign n20529 = ~controllable_hmaster3 & ~n20528;
  assign n20530 = ~n20338 & ~n20529;
  assign n20531 = i_hlock7 & ~n20530;
  assign n20532 = i_hbusreq8 & ~n20504;
  assign n20533 = ~n19660 & ~n20525;
  assign n20534 = ~i_hbusreq8 & ~n20533;
  assign n20535 = ~n20532 & ~n20534;
  assign n20536 = ~controllable_hmaster3 & ~n20535;
  assign n20537 = ~n20338 & ~n20536;
  assign n20538 = ~i_hlock7 & ~n20537;
  assign n20539 = ~n20531 & ~n20538;
  assign n20540 = ~i_hbusreq7 & ~n20539;
  assign n20541 = ~n20509 & ~n20540;
  assign n20542 = ~n7924 & ~n20541;
  assign n20543 = ~n19814 & ~n20395;
  assign n20544 = controllable_hmaster1 & ~n20543;
  assign n20545 = ~n19836 & ~n20544;
  assign n20546 = i_hlock6 & ~n20545;
  assign n20547 = ~n19814 & ~n20406;
  assign n20548 = controllable_hmaster1 & ~n20547;
  assign n20549 = ~n19836 & ~n20548;
  assign n20550 = ~i_hlock6 & ~n20549;
  assign n20551 = ~n20546 & ~n20550;
  assign n20552 = ~controllable_hgrant6 & ~n20551;
  assign n20553 = ~n13894 & ~n20552;
  assign n20554 = ~controllable_hmaster0 & ~n20553;
  assign n20555 = ~n19804 & ~n20554;
  assign n20556 = ~controllable_hmaster3 & ~n20555;
  assign n20557 = ~n20394 & ~n20556;
  assign n20558 = i_hlock7 & ~n20557;
  assign n20559 = ~n19859 & ~n20554;
  assign n20560 = ~controllable_hmaster3 & ~n20559;
  assign n20561 = ~n20394 & ~n20560;
  assign n20562 = ~i_hlock7 & ~n20561;
  assign n20563 = ~n20558 & ~n20562;
  assign n20564 = i_hbusreq7 & ~n20563;
  assign n20565 = i_hbusreq8 & ~n20555;
  assign n20566 = i_hbusreq6 & ~n20551;
  assign n20567 = ~n20175 & ~n20450;
  assign n20568 = controllable_hmaster1 & ~n20567;
  assign n20569 = ~n20219 & ~n20568;
  assign n20570 = i_hlock6 & ~n20569;
  assign n20571 = ~n20175 & ~n20467;
  assign n20572 = controllable_hmaster1 & ~n20571;
  assign n20573 = ~n20219 & ~n20572;
  assign n20574 = ~i_hlock6 & ~n20573;
  assign n20575 = ~n20570 & ~n20574;
  assign n20576 = ~i_hbusreq6 & ~n20575;
  assign n20577 = ~n20566 & ~n20576;
  assign n20578 = ~controllable_hgrant6 & ~n20577;
  assign n20579 = ~n14802 & ~n20578;
  assign n20580 = ~controllable_hmaster0 & ~n20579;
  assign n20581 = ~n20149 & ~n20580;
  assign n20582 = ~i_hbusreq8 & ~n20581;
  assign n20583 = ~n20565 & ~n20582;
  assign n20584 = ~controllable_hmaster3 & ~n20583;
  assign n20585 = ~n20447 & ~n20584;
  assign n20586 = i_hlock7 & ~n20585;
  assign n20587 = i_hbusreq8 & ~n20559;
  assign n20588 = ~n20253 & ~n20580;
  assign n20589 = ~i_hbusreq8 & ~n20588;
  assign n20590 = ~n20587 & ~n20589;
  assign n20591 = ~controllable_hmaster3 & ~n20590;
  assign n20592 = ~n20447 & ~n20591;
  assign n20593 = ~i_hlock7 & ~n20592;
  assign n20594 = ~n20586 & ~n20593;
  assign n20595 = ~i_hbusreq7 & ~n20594;
  assign n20596 = ~n20564 & ~n20595;
  assign n20597 = n7924 & ~n20596;
  assign n20598 = ~n20542 & ~n20597;
  assign n20599 = n8214 & ~n20598;
  assign n20600 = ~n20487 & ~n20599;
  assign n20601 = n8202 & ~n20600;
  assign n20602 = ~n20267 & ~n20601;
  assign n20603 = n7920 & ~n20602;
  assign n20604 = ~n16997 & ~n20603;
  assign n20605 = ~n7728 & ~n20604;
  assign n20606 = ~n18095 & ~n20605;
  assign n20607 = n7723 & ~n20606;
  assign n20608 = ~n7723 & ~n20604;
  assign n20609 = ~n20607 & ~n20608;
  assign n20610 = n7714 & ~n20609;
  assign n20611 = n7723 & ~n20604;
  assign n20612 = controllable_locked & ~n17143;
  assign n20613 = ~controllable_hgrant2 & n20612;
  assign n20614 = ~n7814 & ~n20613;
  assign n20615 = n7733 & ~n20614;
  assign n20616 = ~n17507 & ~n20615;
  assign n20617 = n7928 & ~n20616;
  assign n20618 = ~n19671 & ~n20617;
  assign n20619 = ~controllable_hgrant1 & ~n20618;
  assign n20620 = ~n13155 & ~n20619;
  assign n20621 = ~controllable_hgrant3 & ~n20620;
  assign n20622 = ~n13154 & ~n20621;
  assign n20623 = i_hlock9 & ~n20622;
  assign n20624 = controllable_locked & ~n17476;
  assign n20625 = controllable_locked & ~n20624;
  assign n20626 = ~controllable_hgrant2 & n20625;
  assign n20627 = ~n7814 & ~n20626;
  assign n20628 = n7733 & ~n20627;
  assign n20629 = ~n17507 & ~n20628;
  assign n20630 = n7928 & ~n20629;
  assign n20631 = ~n19671 & ~n20630;
  assign n20632 = ~controllable_hgrant1 & ~n20631;
  assign n20633 = ~n13155 & ~n20632;
  assign n20634 = ~controllable_hgrant3 & ~n20633;
  assign n20635 = ~n13154 & ~n20634;
  assign n20636 = ~i_hlock9 & ~n20635;
  assign n20637 = ~n20623 & ~n20636;
  assign n20638 = ~controllable_hgrant4 & ~n20637;
  assign n20639 = ~n13153 & ~n20638;
  assign n20640 = ~controllable_hgrant5 & ~n20639;
  assign n20641 = ~n13152 & ~n20640;
  assign n20642 = controllable_hmaster1 & ~n20641;
  assign n20643 = controllable_hmaster2 & ~n20641;
  assign n20644 = controllable_locked & ~n17363;
  assign n20645 = ~controllable_hgrant2 & n20644;
  assign n20646 = ~n7814 & ~n20645;
  assign n20647 = n7733 & ~n20646;
  assign n20648 = ~n16507 & ~n20647;
  assign n20649 = n7928 & ~n20648;
  assign n20650 = ~n16128 & ~n20649;
  assign n20651 = ~controllable_hgrant1 & ~n20650;
  assign n20652 = ~n12611 & ~n20651;
  assign n20653 = ~controllable_hgrant3 & ~n20652;
  assign n20654 = ~n12610 & ~n20653;
  assign n20655 = i_hlock9 & ~n20654;
  assign n20656 = ~controllable_hmastlock & ~n17476;
  assign n20657 = ~controllable_hmastlock & ~n20656;
  assign n20658 = controllable_locked & ~n20657;
  assign n20659 = controllable_locked & ~n20658;
  assign n20660 = ~controllable_hgrant2 & n20659;
  assign n20661 = ~n7814 & ~n20660;
  assign n20662 = n7733 & ~n20661;
  assign n20663 = ~n16507 & ~n20662;
  assign n20664 = n7928 & ~n20663;
  assign n20665 = ~n16146 & ~n20664;
  assign n20666 = ~controllable_hgrant1 & ~n20665;
  assign n20667 = ~n12638 & ~n20666;
  assign n20668 = ~controllable_hgrant3 & ~n20667;
  assign n20669 = ~n12637 & ~n20668;
  assign n20670 = ~i_hlock9 & ~n20669;
  assign n20671 = ~n20655 & ~n20670;
  assign n20672 = ~controllable_hgrant4 & ~n20671;
  assign n20673 = ~n12609 & ~n20672;
  assign n20674 = ~controllable_hgrant5 & ~n20673;
  assign n20675 = ~n12608 & ~n20674;
  assign n20676 = ~controllable_hmaster2 & ~n20675;
  assign n20677 = ~n20643 & ~n20676;
  assign n20678 = ~controllable_hmaster1 & ~n20677;
  assign n20679 = ~n20642 & ~n20678;
  assign n20680 = ~controllable_hgrant6 & ~n20679;
  assign n20681 = ~n13122 & ~n20680;
  assign n20682 = controllable_hmaster0 & ~n20681;
  assign n20683 = ~n18547 & ~n20643;
  assign n20684 = ~controllable_hmaster1 & ~n20683;
  assign n20685 = ~n20642 & ~n20684;
  assign n20686 = ~controllable_hgrant6 & ~n20685;
  assign n20687 = ~n13406 & ~n20686;
  assign n20688 = ~controllable_hmaster0 & ~n20687;
  assign n20689 = ~n20682 & ~n20688;
  assign n20690 = i_hlock8 & ~n20689;
  assign n20691 = ~n18573 & ~n20643;
  assign n20692 = ~controllable_hmaster1 & ~n20691;
  assign n20693 = ~n20642 & ~n20692;
  assign n20694 = ~controllable_hgrant6 & ~n20693;
  assign n20695 = ~n13427 & ~n20694;
  assign n20696 = ~controllable_hmaster0 & ~n20695;
  assign n20697 = ~n20682 & ~n20696;
  assign n20698 = ~i_hlock8 & ~n20697;
  assign n20699 = ~n20690 & ~n20698;
  assign n20700 = controllable_hmaster3 & ~n20699;
  assign n20701 = ~n8221 & ~n20617;
  assign n20702 = ~controllable_hgrant1 & ~n20701;
  assign n20703 = ~n12611 & ~n20702;
  assign n20704 = ~controllable_hgrant3 & ~n20703;
  assign n20705 = ~n12610 & ~n20704;
  assign n20706 = i_hlock9 & ~n20705;
  assign n20707 = ~n8221 & ~n20630;
  assign n20708 = ~controllable_hgrant1 & ~n20707;
  assign n20709 = ~n12611 & ~n20708;
  assign n20710 = ~controllable_hgrant3 & ~n20709;
  assign n20711 = ~n12610 & ~n20710;
  assign n20712 = ~i_hlock9 & ~n20711;
  assign n20713 = ~n20706 & ~n20712;
  assign n20714 = ~controllable_hgrant4 & ~n20713;
  assign n20715 = ~n13408 & ~n20714;
  assign n20716 = ~controllable_hgrant5 & ~n20715;
  assign n20717 = ~n13407 & ~n20716;
  assign n20718 = controllable_hmaster2 & ~n20717;
  assign n20719 = i_hlock3 & ~n20703;
  assign n20720 = ~n8235 & ~n20617;
  assign n20721 = ~controllable_hgrant1 & ~n20720;
  assign n20722 = ~n12638 & ~n20721;
  assign n20723 = ~i_hlock3 & ~n20722;
  assign n20724 = ~n20719 & ~n20723;
  assign n20725 = ~controllable_hgrant3 & ~n20724;
  assign n20726 = ~n13852 & ~n20725;
  assign n20727 = i_hlock9 & ~n20726;
  assign n20728 = i_hlock3 & ~n20709;
  assign n20729 = ~n8235 & ~n20630;
  assign n20730 = ~controllable_hgrant1 & ~n20729;
  assign n20731 = ~n12638 & ~n20730;
  assign n20732 = ~i_hlock3 & ~n20731;
  assign n20733 = ~n20728 & ~n20732;
  assign n20734 = ~controllable_hgrant3 & ~n20733;
  assign n20735 = ~n13852 & ~n20734;
  assign n20736 = ~i_hlock9 & ~n20735;
  assign n20737 = ~n20727 & ~n20736;
  assign n20738 = ~controllable_hgrant4 & ~n20737;
  assign n20739 = ~n13851 & ~n20738;
  assign n20740 = ~controllable_hgrant5 & ~n20739;
  assign n20741 = ~n13850 & ~n20740;
  assign n20742 = ~controllable_hmaster2 & ~n20741;
  assign n20743 = ~n20718 & ~n20742;
  assign n20744 = controllable_hmaster1 & ~n20743;
  assign n20745 = i_hlock5 & ~n20715;
  assign n20746 = ~controllable_hgrant3 & ~n20722;
  assign n20747 = ~n12637 & ~n20746;
  assign n20748 = i_hlock9 & ~n20747;
  assign n20749 = ~controllable_hgrant3 & ~n20731;
  assign n20750 = ~n12637 & ~n20749;
  assign n20751 = ~i_hlock9 & ~n20750;
  assign n20752 = ~n20748 & ~n20751;
  assign n20753 = ~controllable_hgrant4 & ~n20752;
  assign n20754 = ~n13429 & ~n20753;
  assign n20755 = ~i_hlock5 & ~n20754;
  assign n20756 = ~n20745 & ~n20755;
  assign n20757 = ~controllable_hgrant5 & ~n20756;
  assign n20758 = ~n13865 & ~n20757;
  assign n20759 = controllable_hmaster2 & ~n20758;
  assign n20760 = i_hlock1 & ~n20701;
  assign n20761 = ~i_hlock1 & ~n20720;
  assign n20762 = ~n20760 & ~n20761;
  assign n20763 = ~controllable_hgrant1 & ~n20762;
  assign n20764 = ~n13875 & ~n20763;
  assign n20765 = ~controllable_hgrant3 & ~n20764;
  assign n20766 = ~n13874 & ~n20765;
  assign n20767 = i_hlock9 & ~n20766;
  assign n20768 = i_hlock1 & ~n20707;
  assign n20769 = ~i_hlock1 & ~n20729;
  assign n20770 = ~n20768 & ~n20769;
  assign n20771 = ~controllable_hgrant1 & ~n20770;
  assign n20772 = ~n13875 & ~n20771;
  assign n20773 = ~controllable_hgrant3 & ~n20772;
  assign n20774 = ~n13874 & ~n20773;
  assign n20775 = ~i_hlock9 & ~n20774;
  assign n20776 = ~n20767 & ~n20775;
  assign n20777 = ~controllable_hgrant4 & ~n20776;
  assign n20778 = ~n13873 & ~n20777;
  assign n20779 = ~controllable_hgrant5 & ~n20778;
  assign n20780 = ~n13872 & ~n20779;
  assign n20781 = ~controllable_hmaster2 & ~n20780;
  assign n20782 = ~n20759 & ~n20781;
  assign n20783 = ~controllable_hmaster1 & ~n20782;
  assign n20784 = ~n20744 & ~n20783;
  assign n20785 = ~controllable_hgrant6 & ~n20784;
  assign n20786 = ~n13849 & ~n20785;
  assign n20787 = controllable_hmaster0 & ~n20786;
  assign n20788 = ~n9213 & ~n20617;
  assign n20789 = ~controllable_hgrant1 & ~n20788;
  assign n20790 = ~n13898 & ~n20789;
  assign n20791 = ~controllable_hgrant3 & ~n20790;
  assign n20792 = ~n13897 & ~n20791;
  assign n20793 = i_hlock9 & ~n20792;
  assign n20794 = ~n9213 & ~n20630;
  assign n20795 = ~controllable_hgrant1 & ~n20794;
  assign n20796 = ~n13898 & ~n20795;
  assign n20797 = ~controllable_hgrant3 & ~n20796;
  assign n20798 = ~n13897 & ~n20797;
  assign n20799 = ~i_hlock9 & ~n20798;
  assign n20800 = ~n20793 & ~n20799;
  assign n20801 = ~controllable_hgrant4 & ~n20800;
  assign n20802 = ~n13896 & ~n20801;
  assign n20803 = ~controllable_hgrant5 & ~n20802;
  assign n20804 = ~n13895 & ~n20803;
  assign n20805 = ~controllable_hmaster2 & ~n20804;
  assign n20806 = ~n20718 & ~n20805;
  assign n20807 = controllable_hmaster1 & ~n20806;
  assign n20808 = i_hlock4 & ~n20713;
  assign n20809 = ~i_hlock4 & ~n20752;
  assign n20810 = ~n20808 & ~n20809;
  assign n20811 = ~controllable_hgrant4 & ~n20810;
  assign n20812 = ~n13912 & ~n20811;
  assign n20813 = ~controllable_hgrant5 & ~n20812;
  assign n20814 = ~n13911 & ~n20813;
  assign n20815 = controllable_hmaster2 & ~n20814;
  assign n20816 = ~n8440 & ~n20617;
  assign n20817 = ~controllable_hgrant1 & ~n20816;
  assign n20818 = ~n13924 & ~n20817;
  assign n20819 = ~controllable_hgrant3 & ~n20818;
  assign n20820 = ~n13923 & ~n20819;
  assign n20821 = i_hlock9 & ~n20820;
  assign n20822 = ~n8440 & ~n20630;
  assign n20823 = ~controllable_hgrant1 & ~n20822;
  assign n20824 = ~n13924 & ~n20823;
  assign n20825 = ~controllable_hgrant3 & ~n20824;
  assign n20826 = ~n13923 & ~n20825;
  assign n20827 = ~i_hlock9 & ~n20826;
  assign n20828 = ~n20821 & ~n20827;
  assign n20829 = ~controllable_hgrant4 & ~n20828;
  assign n20830 = ~n13922 & ~n20829;
  assign n20831 = ~controllable_hgrant5 & ~n20830;
  assign n20832 = ~n13921 & ~n20831;
  assign n20833 = ~controllable_hmaster2 & ~n20832;
  assign n20834 = ~n20815 & ~n20833;
  assign n20835 = ~controllable_hmaster1 & ~n20834;
  assign n20836 = ~n20807 & ~n20835;
  assign n20837 = i_hlock6 & ~n20836;
  assign n20838 = ~controllable_hgrant5 & ~n20754;
  assign n20839 = ~n13428 & ~n20838;
  assign n20840 = controllable_hmaster2 & ~n20839;
  assign n20841 = ~n20805 & ~n20840;
  assign n20842 = controllable_hmaster1 & ~n20841;
  assign n20843 = ~n20835 & ~n20842;
  assign n20844 = ~i_hlock6 & ~n20843;
  assign n20845 = ~n20837 & ~n20844;
  assign n20846 = ~controllable_hgrant6 & ~n20845;
  assign n20847 = ~n13894 & ~n20846;
  assign n20848 = ~controllable_hmaster0 & ~n20847;
  assign n20849 = ~n20787 & ~n20848;
  assign n20850 = ~controllable_hmaster3 & ~n20849;
  assign n20851 = ~n20700 & ~n20850;
  assign n20852 = i_hlock7 & ~n20851;
  assign n20853 = ~n20742 & ~n20840;
  assign n20854 = controllable_hmaster1 & ~n20853;
  assign n20855 = ~n20783 & ~n20854;
  assign n20856 = ~controllable_hgrant6 & ~n20855;
  assign n20857 = ~n13951 & ~n20856;
  assign n20858 = controllable_hmaster0 & ~n20857;
  assign n20859 = ~n20848 & ~n20858;
  assign n20860 = ~controllable_hmaster3 & ~n20859;
  assign n20861 = ~n20700 & ~n20860;
  assign n20862 = ~i_hlock7 & ~n20861;
  assign n20863 = ~n20852 & ~n20862;
  assign n20864 = i_hbusreq7 & ~n20863;
  assign n20865 = i_hbusreq8 & ~n20699;
  assign n20866 = i_hbusreq6 & ~n20679;
  assign n20867 = i_hbusreq5 & ~n20639;
  assign n20868 = i_hbusreq4 & ~n20637;
  assign n20869 = i_hbusreq9 & ~n20637;
  assign n20870 = i_hbusreq3 & ~n20620;
  assign n20871 = i_hbusreq1 & ~n20618;
  assign n20872 = i_hbusreq2 & ~n20612;
  assign n20873 = i_hbusreq0 & ~n20612;
  assign n20874 = ~n12799 & ~n16483;
  assign n20875 = i_hlock0 & ~n20874;
  assign n20876 = ~i_hlock0 & ~n20625;
  assign n20877 = ~n20875 & ~n20876;
  assign n20878 = ~i_hbusreq0 & ~n20877;
  assign n20879 = ~n20873 & ~n20878;
  assign n20880 = ~i_hbusreq2 & ~n20879;
  assign n20881 = ~n20872 & ~n20880;
  assign n20882 = ~controllable_hgrant2 & n20881;
  assign n20883 = ~n12694 & ~n20882;
  assign n20884 = n7733 & ~n20883;
  assign n20885 = ~n18800 & ~n20884;
  assign n20886 = n7928 & ~n20885;
  assign n20887 = ~n19873 & ~n20886;
  assign n20888 = ~i_hbusreq1 & ~n20887;
  assign n20889 = ~n20871 & ~n20888;
  assign n20890 = ~controllable_hgrant1 & ~n20889;
  assign n20891 = ~n13968 & ~n20890;
  assign n20892 = ~i_hbusreq3 & ~n20891;
  assign n20893 = ~n20870 & ~n20892;
  assign n20894 = ~controllable_hgrant3 & ~n20893;
  assign n20895 = ~n13967 & ~n20894;
  assign n20896 = i_hlock9 & ~n20895;
  assign n20897 = i_hbusreq3 & ~n20633;
  assign n20898 = i_hbusreq1 & ~n20631;
  assign n20899 = i_hbusreq2 & ~n20625;
  assign n20900 = i_hbusreq0 & ~n20625;
  assign n20901 = ~n20878 & ~n20900;
  assign n20902 = ~i_hbusreq2 & ~n20901;
  assign n20903 = ~n20899 & ~n20902;
  assign n20904 = ~controllable_hgrant2 & n20903;
  assign n20905 = ~n12694 & ~n20904;
  assign n20906 = n7733 & ~n20905;
  assign n20907 = ~n18800 & ~n20906;
  assign n20908 = n7928 & ~n20907;
  assign n20909 = ~n19873 & ~n20908;
  assign n20910 = ~i_hbusreq1 & ~n20909;
  assign n20911 = ~n20898 & ~n20910;
  assign n20912 = ~controllable_hgrant1 & ~n20911;
  assign n20913 = ~n13968 & ~n20912;
  assign n20914 = ~i_hbusreq3 & ~n20913;
  assign n20915 = ~n20897 & ~n20914;
  assign n20916 = ~controllable_hgrant3 & ~n20915;
  assign n20917 = ~n13967 & ~n20916;
  assign n20918 = ~i_hlock9 & ~n20917;
  assign n20919 = ~n20896 & ~n20918;
  assign n20920 = ~i_hbusreq9 & ~n20919;
  assign n20921 = ~n20869 & ~n20920;
  assign n20922 = ~i_hbusreq4 & ~n20921;
  assign n20923 = ~n20868 & ~n20922;
  assign n20924 = ~controllable_hgrant4 & ~n20923;
  assign n20925 = ~n13966 & ~n20924;
  assign n20926 = ~i_hbusreq5 & ~n20925;
  assign n20927 = ~n20867 & ~n20926;
  assign n20928 = ~controllable_hgrant5 & ~n20927;
  assign n20929 = ~n13965 & ~n20928;
  assign n20930 = controllable_hmaster1 & ~n20929;
  assign n20931 = controllable_hmaster2 & ~n20929;
  assign n20932 = i_hbusreq5 & ~n20673;
  assign n20933 = i_hbusreq4 & ~n20671;
  assign n20934 = i_hbusreq9 & ~n20671;
  assign n20935 = i_hbusreq3 & ~n20652;
  assign n20936 = i_hbusreq1 & ~n20650;
  assign n20937 = i_hbusreq2 & ~n20644;
  assign n20938 = i_hbusreq0 & ~n20644;
  assign n20939 = ~controllable_hmastlock & n7970;
  assign n20940 = ~n7858 & ~n20939;
  assign n20941 = controllable_locked & ~n20940;
  assign n20942 = ~n12799 & ~n20941;
  assign n20943 = i_hlock0 & ~n20942;
  assign n20944 = ~i_hlock0 & ~n20659;
  assign n20945 = ~n20943 & ~n20944;
  assign n20946 = ~i_hbusreq0 & ~n20945;
  assign n20947 = ~n20938 & ~n20946;
  assign n20948 = ~i_hbusreq2 & ~n20947;
  assign n20949 = ~n20937 & ~n20948;
  assign n20950 = ~controllable_hgrant2 & n20949;
  assign n20951 = ~n12694 & ~n20950;
  assign n20952 = n7733 & ~n20951;
  assign n20953 = ~n16635 & ~n20952;
  assign n20954 = n7928 & ~n20953;
  assign n20955 = ~n16191 & ~n20954;
  assign n20956 = ~i_hbusreq1 & ~n20955;
  assign n20957 = ~n20936 & ~n20956;
  assign n20958 = ~controllable_hgrant1 & ~n20957;
  assign n20959 = ~n14023 & ~n20958;
  assign n20960 = ~i_hbusreq3 & ~n20959;
  assign n20961 = ~n20935 & ~n20960;
  assign n20962 = ~controllable_hgrant3 & ~n20961;
  assign n20963 = ~n14022 & ~n20962;
  assign n20964 = i_hlock9 & ~n20963;
  assign n20965 = i_hbusreq3 & ~n20667;
  assign n20966 = i_hbusreq1 & ~n20665;
  assign n20967 = i_hbusreq2 & ~n20659;
  assign n20968 = i_hbusreq0 & ~n20659;
  assign n20969 = ~n20946 & ~n20968;
  assign n20970 = ~i_hbusreq2 & ~n20969;
  assign n20971 = ~n20967 & ~n20970;
  assign n20972 = ~controllable_hgrant2 & n20971;
  assign n20973 = ~n12694 & ~n20972;
  assign n20974 = n7733 & ~n20973;
  assign n20975 = ~n16635 & ~n20974;
  assign n20976 = n7928 & ~n20975;
  assign n20977 = ~n16216 & ~n20976;
  assign n20978 = ~i_hbusreq1 & ~n20977;
  assign n20979 = ~n20966 & ~n20978;
  assign n20980 = ~controllable_hgrant1 & ~n20979;
  assign n20981 = ~n14058 & ~n20980;
  assign n20982 = ~i_hbusreq3 & ~n20981;
  assign n20983 = ~n20965 & ~n20982;
  assign n20984 = ~controllable_hgrant3 & ~n20983;
  assign n20985 = ~n14057 & ~n20984;
  assign n20986 = ~i_hlock9 & ~n20985;
  assign n20987 = ~n20964 & ~n20986;
  assign n20988 = ~i_hbusreq9 & ~n20987;
  assign n20989 = ~n20934 & ~n20988;
  assign n20990 = ~i_hbusreq4 & ~n20989;
  assign n20991 = ~n20933 & ~n20990;
  assign n20992 = ~controllable_hgrant4 & ~n20991;
  assign n20993 = ~n14322 & ~n20992;
  assign n20994 = ~i_hbusreq5 & ~n20993;
  assign n20995 = ~n20932 & ~n20994;
  assign n20996 = ~controllable_hgrant5 & ~n20995;
  assign n20997 = ~n14321 & ~n20996;
  assign n20998 = ~controllable_hmaster2 & ~n20997;
  assign n20999 = ~n20931 & ~n20998;
  assign n21000 = ~controllable_hmaster1 & ~n20999;
  assign n21001 = ~n20930 & ~n21000;
  assign n21002 = ~i_hbusreq6 & ~n21001;
  assign n21003 = ~n20866 & ~n21002;
  assign n21004 = ~controllable_hgrant6 & ~n21003;
  assign n21005 = ~n14320 & ~n21004;
  assign n21006 = controllable_hmaster0 & ~n21005;
  assign n21007 = i_hbusreq6 & ~n20685;
  assign n21008 = ~n14241 & ~n17553;
  assign n21009 = controllable_locked & ~n21008;
  assign n21010 = ~n14243 & ~n21009;
  assign n21011 = i_hlock0 & ~n21010;
  assign n21012 = ~n18726 & ~n21011;
  assign n21013 = ~i_hbusreq0 & ~n21012;
  assign n21014 = ~n17552 & ~n21013;
  assign n21015 = ~i_hbusreq2 & ~n21014;
  assign n21016 = ~n17551 & ~n21015;
  assign n21017 = ~controllable_hgrant2 & n21016;
  assign n21018 = ~n12706 & ~n21017;
  assign n21019 = n7733 & ~n21018;
  assign n21020 = ~n18800 & ~n21019;
  assign n21021 = n7928 & ~n21020;
  assign n21022 = ~n8265 & ~n21021;
  assign n21023 = ~i_hbusreq1 & ~n21022;
  assign n21024 = ~n18791 & ~n21023;
  assign n21025 = ~controllable_hgrant1 & ~n21024;
  assign n21026 = ~n12681 & ~n21025;
  assign n21027 = ~i_hbusreq3 & ~n21026;
  assign n21028 = ~n18790 & ~n21027;
  assign n21029 = ~controllable_hgrant3 & ~n21028;
  assign n21030 = ~n12679 & ~n21029;
  assign n21031 = i_hlock9 & ~n21030;
  assign n21032 = ~n17580 & ~n21013;
  assign n21033 = ~i_hbusreq2 & ~n21032;
  assign n21034 = ~n17579 & ~n21033;
  assign n21035 = ~controllable_hgrant2 & n21034;
  assign n21036 = ~n12706 & ~n21035;
  assign n21037 = n7733 & ~n21036;
  assign n21038 = ~n18800 & ~n21037;
  assign n21039 = n7928 & ~n21038;
  assign n21040 = ~n8265 & ~n21039;
  assign n21041 = ~i_hbusreq1 & ~n21040;
  assign n21042 = ~n18814 & ~n21041;
  assign n21043 = ~controllable_hgrant1 & ~n21042;
  assign n21044 = ~n12681 & ~n21043;
  assign n21045 = ~i_hbusreq3 & ~n21044;
  assign n21046 = ~n18813 & ~n21045;
  assign n21047 = ~controllable_hgrant3 & ~n21046;
  assign n21048 = ~n12679 & ~n21047;
  assign n21049 = ~i_hlock9 & ~n21048;
  assign n21050 = ~n21031 & ~n21049;
  assign n21051 = ~i_hbusreq9 & ~n21050;
  assign n21052 = ~n18789 & ~n21051;
  assign n21053 = ~i_hbusreq4 & ~n21052;
  assign n21054 = ~n18788 & ~n21053;
  assign n21055 = ~controllable_hgrant4 & ~n21054;
  assign n21056 = ~n13524 & ~n21055;
  assign n21057 = ~i_hbusreq5 & ~n21056;
  assign n21058 = ~n18787 & ~n21057;
  assign n21059 = ~controllable_hgrant5 & ~n21058;
  assign n21060 = ~n13522 & ~n21059;
  assign n21061 = ~controllable_hmaster2 & ~n21060;
  assign n21062 = ~n20931 & ~n21061;
  assign n21063 = ~controllable_hmaster1 & ~n21062;
  assign n21064 = ~n20930 & ~n21063;
  assign n21065 = ~i_hbusreq6 & ~n21064;
  assign n21066 = ~n21007 & ~n21065;
  assign n21067 = ~controllable_hgrant6 & ~n21066;
  assign n21068 = ~n14443 & ~n21067;
  assign n21069 = ~controllable_hmaster0 & ~n21068;
  assign n21070 = ~n21006 & ~n21069;
  assign n21071 = i_hlock8 & ~n21070;
  assign n21072 = i_hbusreq6 & ~n20693;
  assign n21073 = ~n8297 & ~n21021;
  assign n21074 = ~i_hbusreq1 & ~n21073;
  assign n21075 = ~n18854 & ~n21074;
  assign n21076 = ~controllable_hgrant1 & ~n21075;
  assign n21077 = ~n12730 & ~n21076;
  assign n21078 = ~i_hbusreq3 & ~n21077;
  assign n21079 = ~n18853 & ~n21078;
  assign n21080 = ~controllable_hgrant3 & ~n21079;
  assign n21081 = ~n12728 & ~n21080;
  assign n21082 = i_hlock9 & ~n21081;
  assign n21083 = ~n8297 & ~n21039;
  assign n21084 = ~i_hbusreq1 & ~n21083;
  assign n21085 = ~n18866 & ~n21084;
  assign n21086 = ~controllable_hgrant1 & ~n21085;
  assign n21087 = ~n12730 & ~n21086;
  assign n21088 = ~i_hbusreq3 & ~n21087;
  assign n21089 = ~n18865 & ~n21088;
  assign n21090 = ~controllable_hgrant3 & ~n21089;
  assign n21091 = ~n12728 & ~n21090;
  assign n21092 = ~i_hlock9 & ~n21091;
  assign n21093 = ~n21082 & ~n21092;
  assign n21094 = ~i_hbusreq9 & ~n21093;
  assign n21095 = ~n18852 & ~n21094;
  assign n21096 = ~i_hbusreq4 & ~n21095;
  assign n21097 = ~n18851 & ~n21096;
  assign n21098 = ~controllable_hgrant4 & ~n21097;
  assign n21099 = ~n13577 & ~n21098;
  assign n21100 = ~i_hbusreq5 & ~n21099;
  assign n21101 = ~n18850 & ~n21100;
  assign n21102 = ~controllable_hgrant5 & ~n21101;
  assign n21103 = ~n13575 & ~n21102;
  assign n21104 = ~controllable_hmaster2 & ~n21103;
  assign n21105 = ~n20931 & ~n21104;
  assign n21106 = ~controllable_hmaster1 & ~n21105;
  assign n21107 = ~n20930 & ~n21106;
  assign n21108 = ~i_hbusreq6 & ~n21107;
  assign n21109 = ~n21072 & ~n21108;
  assign n21110 = ~controllable_hgrant6 & ~n21109;
  assign n21111 = ~n14484 & ~n21110;
  assign n21112 = ~controllable_hmaster0 & ~n21111;
  assign n21113 = ~n21006 & ~n21112;
  assign n21114 = ~i_hlock8 & ~n21113;
  assign n21115 = ~n21071 & ~n21114;
  assign n21116 = ~i_hbusreq8 & ~n21115;
  assign n21117 = ~n20865 & ~n21116;
  assign n21118 = controllable_hmaster3 & ~n21117;
  assign n21119 = i_hbusreq8 & ~n20849;
  assign n21120 = i_hbusreq6 & ~n20784;
  assign n21121 = i_hbusreq5 & ~n20715;
  assign n21122 = i_hbusreq4 & ~n20713;
  assign n21123 = i_hbusreq9 & ~n20713;
  assign n21124 = i_hbusreq3 & ~n20703;
  assign n21125 = i_hbusreq1 & ~n20701;
  assign n21126 = ~n8265 & ~n20886;
  assign n21127 = ~i_hbusreq1 & ~n21126;
  assign n21128 = ~n21125 & ~n21127;
  assign n21129 = ~controllable_hgrant1 & ~n21128;
  assign n21130 = ~n14023 & ~n21129;
  assign n21131 = ~i_hbusreq3 & ~n21130;
  assign n21132 = ~n21124 & ~n21131;
  assign n21133 = ~controllable_hgrant3 & ~n21132;
  assign n21134 = ~n14022 & ~n21133;
  assign n21135 = i_hlock9 & ~n21134;
  assign n21136 = i_hbusreq3 & ~n20709;
  assign n21137 = i_hbusreq1 & ~n20707;
  assign n21138 = ~n8265 & ~n20908;
  assign n21139 = ~i_hbusreq1 & ~n21138;
  assign n21140 = ~n21137 & ~n21139;
  assign n21141 = ~controllable_hgrant1 & ~n21140;
  assign n21142 = ~n14023 & ~n21141;
  assign n21143 = ~i_hbusreq3 & ~n21142;
  assign n21144 = ~n21136 & ~n21143;
  assign n21145 = ~controllable_hgrant3 & ~n21144;
  assign n21146 = ~n14022 & ~n21145;
  assign n21147 = ~i_hlock9 & ~n21146;
  assign n21148 = ~n21135 & ~n21147;
  assign n21149 = ~i_hbusreq9 & ~n21148;
  assign n21150 = ~n21123 & ~n21149;
  assign n21151 = ~i_hbusreq4 & ~n21150;
  assign n21152 = ~n21122 & ~n21151;
  assign n21153 = ~controllable_hgrant4 & ~n21152;
  assign n21154 = ~n14021 & ~n21153;
  assign n21155 = ~i_hbusreq5 & ~n21154;
  assign n21156 = ~n21121 & ~n21155;
  assign n21157 = ~controllable_hgrant5 & ~n21156;
  assign n21158 = ~n14020 & ~n21157;
  assign n21159 = controllable_hmaster2 & ~n21158;
  assign n21160 = i_hbusreq5 & ~n20739;
  assign n21161 = i_hbusreq4 & ~n20737;
  assign n21162 = i_hbusreq9 & ~n20737;
  assign n21163 = i_hbusreq3 & ~n20724;
  assign n21164 = i_hlock3 & ~n21130;
  assign n21165 = i_hbusreq1 & ~n20720;
  assign n21166 = ~n8297 & ~n20886;
  assign n21167 = ~i_hbusreq1 & ~n21166;
  assign n21168 = ~n21165 & ~n21167;
  assign n21169 = ~controllable_hgrant1 & ~n21168;
  assign n21170 = ~n14058 & ~n21169;
  assign n21171 = ~i_hlock3 & ~n21170;
  assign n21172 = ~n21164 & ~n21171;
  assign n21173 = ~i_hbusreq3 & ~n21172;
  assign n21174 = ~n21163 & ~n21173;
  assign n21175 = ~controllable_hgrant3 & ~n21174;
  assign n21176 = ~n14102 & ~n21175;
  assign n21177 = i_hlock9 & ~n21176;
  assign n21178 = i_hbusreq3 & ~n20733;
  assign n21179 = i_hlock3 & ~n21142;
  assign n21180 = i_hbusreq1 & ~n20729;
  assign n21181 = ~n8297 & ~n20908;
  assign n21182 = ~i_hbusreq1 & ~n21181;
  assign n21183 = ~n21180 & ~n21182;
  assign n21184 = ~controllable_hgrant1 & ~n21183;
  assign n21185 = ~n14058 & ~n21184;
  assign n21186 = ~i_hlock3 & ~n21185;
  assign n21187 = ~n21179 & ~n21186;
  assign n21188 = ~i_hbusreq3 & ~n21187;
  assign n21189 = ~n21178 & ~n21188;
  assign n21190 = ~controllable_hgrant3 & ~n21189;
  assign n21191 = ~n14102 & ~n21190;
  assign n21192 = ~i_hlock9 & ~n21191;
  assign n21193 = ~n21177 & ~n21192;
  assign n21194 = ~i_hbusreq9 & ~n21193;
  assign n21195 = ~n21162 & ~n21194;
  assign n21196 = ~i_hbusreq4 & ~n21195;
  assign n21197 = ~n21161 & ~n21196;
  assign n21198 = ~controllable_hgrant4 & ~n21197;
  assign n21199 = ~n14099 & ~n21198;
  assign n21200 = ~i_hbusreq5 & ~n21199;
  assign n21201 = ~n21160 & ~n21200;
  assign n21202 = ~controllable_hgrant5 & ~n21201;
  assign n21203 = ~n14097 & ~n21202;
  assign n21204 = ~controllable_hmaster2 & ~n21203;
  assign n21205 = ~n21159 & ~n21204;
  assign n21206 = controllable_hmaster1 & ~n21205;
  assign n21207 = i_hbusreq5 & ~n20756;
  assign n21208 = i_hlock5 & ~n21154;
  assign n21209 = i_hbusreq4 & ~n20752;
  assign n21210 = i_hbusreq9 & ~n20752;
  assign n21211 = i_hbusreq3 & ~n20722;
  assign n21212 = ~i_hbusreq3 & ~n21170;
  assign n21213 = ~n21211 & ~n21212;
  assign n21214 = ~controllable_hgrant3 & ~n21213;
  assign n21215 = ~n14057 & ~n21214;
  assign n21216 = i_hlock9 & ~n21215;
  assign n21217 = i_hbusreq3 & ~n20731;
  assign n21218 = ~i_hbusreq3 & ~n21185;
  assign n21219 = ~n21217 & ~n21218;
  assign n21220 = ~controllable_hgrant3 & ~n21219;
  assign n21221 = ~n14057 & ~n21220;
  assign n21222 = ~i_hlock9 & ~n21221;
  assign n21223 = ~n21216 & ~n21222;
  assign n21224 = ~i_hbusreq9 & ~n21223;
  assign n21225 = ~n21210 & ~n21224;
  assign n21226 = ~i_hbusreq4 & ~n21225;
  assign n21227 = ~n21209 & ~n21226;
  assign n21228 = ~controllable_hgrant4 & ~n21227;
  assign n21229 = ~n14056 & ~n21228;
  assign n21230 = ~i_hlock5 & ~n21229;
  assign n21231 = ~n21208 & ~n21230;
  assign n21232 = ~i_hbusreq5 & ~n21231;
  assign n21233 = ~n21207 & ~n21232;
  assign n21234 = ~controllable_hgrant5 & ~n21233;
  assign n21235 = ~n14124 & ~n21234;
  assign n21236 = controllable_hmaster2 & ~n21235;
  assign n21237 = i_hbusreq5 & ~n20778;
  assign n21238 = i_hbusreq4 & ~n20776;
  assign n21239 = i_hbusreq9 & ~n20776;
  assign n21240 = i_hbusreq3 & ~n20764;
  assign n21241 = i_hbusreq1 & ~n20762;
  assign n21242 = i_hlock1 & ~n21126;
  assign n21243 = ~i_hlock1 & ~n21166;
  assign n21244 = ~n21242 & ~n21243;
  assign n21245 = ~i_hbusreq1 & ~n21244;
  assign n21246 = ~n21241 & ~n21245;
  assign n21247 = ~controllable_hgrant1 & ~n21246;
  assign n21248 = ~n14141 & ~n21247;
  assign n21249 = ~i_hbusreq3 & ~n21248;
  assign n21250 = ~n21240 & ~n21249;
  assign n21251 = ~controllable_hgrant3 & ~n21250;
  assign n21252 = ~n14139 & ~n21251;
  assign n21253 = i_hlock9 & ~n21252;
  assign n21254 = i_hbusreq3 & ~n20772;
  assign n21255 = i_hbusreq1 & ~n20770;
  assign n21256 = i_hlock1 & ~n21138;
  assign n21257 = ~i_hlock1 & ~n21181;
  assign n21258 = ~n21256 & ~n21257;
  assign n21259 = ~i_hbusreq1 & ~n21258;
  assign n21260 = ~n21255 & ~n21259;
  assign n21261 = ~controllable_hgrant1 & ~n21260;
  assign n21262 = ~n14141 & ~n21261;
  assign n21263 = ~i_hbusreq3 & ~n21262;
  assign n21264 = ~n21254 & ~n21263;
  assign n21265 = ~controllable_hgrant3 & ~n21264;
  assign n21266 = ~n14139 & ~n21265;
  assign n21267 = ~i_hlock9 & ~n21266;
  assign n21268 = ~n21253 & ~n21267;
  assign n21269 = ~i_hbusreq9 & ~n21268;
  assign n21270 = ~n21239 & ~n21269;
  assign n21271 = ~i_hbusreq4 & ~n21270;
  assign n21272 = ~n21238 & ~n21271;
  assign n21273 = ~controllable_hgrant4 & ~n21272;
  assign n21274 = ~n14136 & ~n21273;
  assign n21275 = ~i_hbusreq5 & ~n21274;
  assign n21276 = ~n21237 & ~n21275;
  assign n21277 = ~controllable_hgrant5 & ~n21276;
  assign n21278 = ~n14134 & ~n21277;
  assign n21279 = ~controllable_hmaster2 & ~n21278;
  assign n21280 = ~n21236 & ~n21279;
  assign n21281 = ~controllable_hmaster1 & ~n21280;
  assign n21282 = ~n21206 & ~n21281;
  assign n21283 = ~i_hbusreq6 & ~n21282;
  assign n21284 = ~n21120 & ~n21283;
  assign n21285 = ~controllable_hgrant6 & ~n21284;
  assign n21286 = ~n14094 & ~n21285;
  assign n21287 = controllable_hmaster0 & ~n21286;
  assign n21288 = i_hbusreq6 & ~n20845;
  assign n21289 = i_hbusreq5 & ~n20802;
  assign n21290 = i_hbusreq4 & ~n20800;
  assign n21291 = i_hbusreq9 & ~n20800;
  assign n21292 = i_hbusreq3 & ~n20790;
  assign n21293 = i_hbusreq1 & ~n20788;
  assign n21294 = ~n9379 & ~n20886;
  assign n21295 = ~i_hbusreq1 & ~n21294;
  assign n21296 = ~n21293 & ~n21295;
  assign n21297 = ~controllable_hgrant1 & ~n21296;
  assign n21298 = ~n14182 & ~n21297;
  assign n21299 = ~i_hbusreq3 & ~n21298;
  assign n21300 = ~n21292 & ~n21299;
  assign n21301 = ~controllable_hgrant3 & ~n21300;
  assign n21302 = ~n14180 & ~n21301;
  assign n21303 = i_hlock9 & ~n21302;
  assign n21304 = i_hbusreq3 & ~n20796;
  assign n21305 = i_hbusreq1 & ~n20794;
  assign n21306 = ~n9379 & ~n20908;
  assign n21307 = ~i_hbusreq1 & ~n21306;
  assign n21308 = ~n21305 & ~n21307;
  assign n21309 = ~controllable_hgrant1 & ~n21308;
  assign n21310 = ~n14182 & ~n21309;
  assign n21311 = ~i_hbusreq3 & ~n21310;
  assign n21312 = ~n21304 & ~n21311;
  assign n21313 = ~controllable_hgrant3 & ~n21312;
  assign n21314 = ~n14180 & ~n21313;
  assign n21315 = ~i_hlock9 & ~n21314;
  assign n21316 = ~n21303 & ~n21315;
  assign n21317 = ~i_hbusreq9 & ~n21316;
  assign n21318 = ~n21291 & ~n21317;
  assign n21319 = ~i_hbusreq4 & ~n21318;
  assign n21320 = ~n21290 & ~n21319;
  assign n21321 = ~controllable_hgrant4 & ~n21320;
  assign n21322 = ~n14177 & ~n21321;
  assign n21323 = ~i_hbusreq5 & ~n21322;
  assign n21324 = ~n21289 & ~n21323;
  assign n21325 = ~controllable_hgrant5 & ~n21324;
  assign n21326 = ~n14175 & ~n21325;
  assign n21327 = ~controllable_hmaster2 & ~n21326;
  assign n21328 = ~n21159 & ~n21327;
  assign n21329 = controllable_hmaster1 & ~n21328;
  assign n21330 = i_hbusreq5 & ~n20812;
  assign n21331 = i_hbusreq4 & ~n20810;
  assign n21332 = i_hlock4 & ~n21150;
  assign n21333 = ~i_hlock4 & ~n21225;
  assign n21334 = ~n21332 & ~n21333;
  assign n21335 = ~i_hbusreq4 & ~n21334;
  assign n21336 = ~n21331 & ~n21335;
  assign n21337 = ~controllable_hgrant4 & ~n21336;
  assign n21338 = ~n14208 & ~n21337;
  assign n21339 = ~i_hbusreq5 & ~n21338;
  assign n21340 = ~n21330 & ~n21339;
  assign n21341 = ~controllable_hgrant5 & ~n21340;
  assign n21342 = ~n14206 & ~n21341;
  assign n21343 = controllable_hmaster2 & ~n21342;
  assign n21344 = i_hbusreq5 & ~n20830;
  assign n21345 = i_hbusreq4 & ~n20828;
  assign n21346 = i_hbusreq9 & ~n20828;
  assign n21347 = i_hbusreq3 & ~n20818;
  assign n21348 = i_hbusreq1 & ~n20816;
  assign n21349 = ~n17477 & ~n20939;
  assign n21350 = controllable_locked & ~n21349;
  assign n21351 = ~n12896 & ~n21350;
  assign n21352 = i_hlock0 & ~n21351;
  assign n21353 = ~n20876 & ~n21352;
  assign n21354 = ~i_hbusreq0 & ~n21353;
  assign n21355 = ~n20873 & ~n21354;
  assign n21356 = ~i_hbusreq2 & ~n21355;
  assign n21357 = ~n20872 & ~n21356;
  assign n21358 = ~controllable_hgrant2 & n21357;
  assign n21359 = ~n14231 & ~n21358;
  assign n21360 = n7733 & ~n21359;
  assign n21361 = ~n19072 & ~n21360;
  assign n21362 = n7928 & ~n21361;
  assign n21363 = ~n8440 & ~n21362;
  assign n21364 = ~i_hbusreq1 & ~n21363;
  assign n21365 = ~n21348 & ~n21364;
  assign n21366 = ~controllable_hgrant1 & ~n21365;
  assign n21367 = ~n14229 & ~n21366;
  assign n21368 = ~i_hbusreq3 & ~n21367;
  assign n21369 = ~n21347 & ~n21368;
  assign n21370 = ~controllable_hgrant3 & ~n21369;
  assign n21371 = ~n14227 & ~n21370;
  assign n21372 = i_hlock9 & ~n21371;
  assign n21373 = i_hbusreq3 & ~n20824;
  assign n21374 = i_hbusreq1 & ~n20822;
  assign n21375 = ~n20900 & ~n21354;
  assign n21376 = ~i_hbusreq2 & ~n21375;
  assign n21377 = ~n20899 & ~n21376;
  assign n21378 = ~controllable_hgrant2 & n21377;
  assign n21379 = ~n14231 & ~n21378;
  assign n21380 = n7733 & ~n21379;
  assign n21381 = ~n19072 & ~n21380;
  assign n21382 = n7928 & ~n21381;
  assign n21383 = ~n8440 & ~n21382;
  assign n21384 = ~i_hbusreq1 & ~n21383;
  assign n21385 = ~n21374 & ~n21384;
  assign n21386 = ~controllable_hgrant1 & ~n21385;
  assign n21387 = ~n14229 & ~n21386;
  assign n21388 = ~i_hbusreq3 & ~n21387;
  assign n21389 = ~n21373 & ~n21388;
  assign n21390 = ~controllable_hgrant3 & ~n21389;
  assign n21391 = ~n14227 & ~n21390;
  assign n21392 = ~i_hlock9 & ~n21391;
  assign n21393 = ~n21372 & ~n21392;
  assign n21394 = ~i_hbusreq9 & ~n21393;
  assign n21395 = ~n21346 & ~n21394;
  assign n21396 = ~i_hbusreq4 & ~n21395;
  assign n21397 = ~n21345 & ~n21396;
  assign n21398 = ~controllable_hgrant4 & ~n21397;
  assign n21399 = ~n14224 & ~n21398;
  assign n21400 = ~i_hbusreq5 & ~n21399;
  assign n21401 = ~n21344 & ~n21400;
  assign n21402 = ~controllable_hgrant5 & ~n21401;
  assign n21403 = ~n14222 & ~n21402;
  assign n21404 = ~controllable_hmaster2 & ~n21403;
  assign n21405 = ~n21343 & ~n21404;
  assign n21406 = ~controllable_hmaster1 & ~n21405;
  assign n21407 = ~n21329 & ~n21406;
  assign n21408 = i_hlock6 & ~n21407;
  assign n21409 = i_hbusreq5 & ~n20754;
  assign n21410 = ~i_hbusreq5 & ~n21229;
  assign n21411 = ~n21409 & ~n21410;
  assign n21412 = ~controllable_hgrant5 & ~n21411;
  assign n21413 = ~n14055 & ~n21412;
  assign n21414 = controllable_hmaster2 & ~n21413;
  assign n21415 = ~n21327 & ~n21414;
  assign n21416 = controllable_hmaster1 & ~n21415;
  assign n21417 = ~n21406 & ~n21416;
  assign n21418 = ~i_hlock6 & ~n21417;
  assign n21419 = ~n21408 & ~n21418;
  assign n21420 = ~i_hbusreq6 & ~n21419;
  assign n21421 = ~n21288 & ~n21420;
  assign n21422 = ~controllable_hgrant6 & ~n21421;
  assign n21423 = ~n14173 & ~n21422;
  assign n21424 = ~controllable_hmaster0 & ~n21423;
  assign n21425 = ~n21287 & ~n21424;
  assign n21426 = ~i_hbusreq8 & ~n21425;
  assign n21427 = ~n21119 & ~n21426;
  assign n21428 = ~controllable_hmaster3 & ~n21427;
  assign n21429 = ~n21118 & ~n21428;
  assign n21430 = i_hlock7 & ~n21429;
  assign n21431 = i_hbusreq8 & ~n20859;
  assign n21432 = i_hbusreq6 & ~n20855;
  assign n21433 = ~n21204 & ~n21414;
  assign n21434 = controllable_hmaster1 & ~n21433;
  assign n21435 = ~n21281 & ~n21434;
  assign n21436 = ~i_hbusreq6 & ~n21435;
  assign n21437 = ~n21432 & ~n21436;
  assign n21438 = ~controllable_hgrant6 & ~n21437;
  assign n21439 = ~n14298 & ~n21438;
  assign n21440 = controllable_hmaster0 & ~n21439;
  assign n21441 = ~n21424 & ~n21440;
  assign n21442 = ~i_hbusreq8 & ~n21441;
  assign n21443 = ~n21431 & ~n21442;
  assign n21444 = ~controllable_hmaster3 & ~n21443;
  assign n21445 = ~n21118 & ~n21444;
  assign n21446 = ~i_hlock7 & ~n21445;
  assign n21447 = ~n21430 & ~n21446;
  assign n21448 = ~i_hbusreq7 & ~n21447;
  assign n21449 = ~n20864 & ~n21448;
  assign n21450 = n7924 & ~n21449;
  assign n21451 = ~n19670 & ~n21450;
  assign n21452 = n8214 & ~n21451;
  assign n21453 = ~n19172 & ~n21452;
  assign n21454 = ~n8202 & ~n21453;
  assign n21455 = ~controllable_hmaster2 & ~n20717;
  assign n21456 = ~n20643 & ~n21455;
  assign n21457 = ~controllable_hmaster1 & ~n21456;
  assign n21458 = ~n20642 & ~n21457;
  assign n21459 = ~controllable_hgrant6 & ~n21458;
  assign n21460 = ~n13406 & ~n21459;
  assign n21461 = ~controllable_hmaster0 & ~n21460;
  assign n21462 = ~n20682 & ~n21461;
  assign n21463 = i_hlock8 & ~n21462;
  assign n21464 = ~controllable_hmaster2 & ~n20839;
  assign n21465 = ~n20643 & ~n21464;
  assign n21466 = ~controllable_hmaster1 & ~n21465;
  assign n21467 = ~n20642 & ~n21466;
  assign n21468 = ~controllable_hgrant6 & ~n21467;
  assign n21469 = ~n13427 & ~n21468;
  assign n21470 = ~controllable_hmaster0 & ~n21469;
  assign n21471 = ~n20682 & ~n21470;
  assign n21472 = ~i_hlock8 & ~n21471;
  assign n21473 = ~n21463 & ~n21472;
  assign n21474 = controllable_hmaster3 & ~n21473;
  assign n21475 = ~n18584 & ~n20742;
  assign n21476 = controllable_hmaster1 & ~n21475;
  assign n21477 = ~n20783 & ~n21476;
  assign n21478 = ~controllable_hgrant6 & ~n21477;
  assign n21479 = ~n13849 & ~n21478;
  assign n21480 = controllable_hmaster0 & ~n21479;
  assign n21481 = ~n20848 & ~n21480;
  assign n21482 = ~controllable_hmaster3 & ~n21481;
  assign n21483 = ~n21474 & ~n21482;
  assign n21484 = i_hlock7 & ~n21483;
  assign n21485 = ~n18689 & ~n20742;
  assign n21486 = controllable_hmaster1 & ~n21485;
  assign n21487 = ~n20783 & ~n21486;
  assign n21488 = ~controllable_hgrant6 & ~n21487;
  assign n21489 = ~n13951 & ~n21488;
  assign n21490 = controllable_hmaster0 & ~n21489;
  assign n21491 = ~n20848 & ~n21490;
  assign n21492 = ~controllable_hmaster3 & ~n21491;
  assign n21493 = ~n21474 & ~n21492;
  assign n21494 = ~i_hlock7 & ~n21493;
  assign n21495 = ~n21484 & ~n21494;
  assign n21496 = i_hbusreq7 & ~n21495;
  assign n21497 = i_hbusreq8 & ~n21473;
  assign n21498 = i_hbusreq6 & ~n21458;
  assign n21499 = ~controllable_hmaster2 & ~n21158;
  assign n21500 = ~n20931 & ~n21499;
  assign n21501 = ~controllable_hmaster1 & ~n21500;
  assign n21502 = ~n20930 & ~n21501;
  assign n21503 = ~i_hbusreq6 & ~n21502;
  assign n21504 = ~n21498 & ~n21503;
  assign n21505 = ~controllable_hgrant6 & ~n21504;
  assign n21506 = ~n14019 & ~n21505;
  assign n21507 = ~controllable_hmaster0 & ~n21506;
  assign n21508 = ~n21006 & ~n21507;
  assign n21509 = i_hlock8 & ~n21508;
  assign n21510 = i_hbusreq6 & ~n21467;
  assign n21511 = ~controllable_hmaster2 & ~n21413;
  assign n21512 = ~n20931 & ~n21511;
  assign n21513 = ~controllable_hmaster1 & ~n21512;
  assign n21514 = ~n20930 & ~n21513;
  assign n21515 = ~i_hbusreq6 & ~n21514;
  assign n21516 = ~n21510 & ~n21515;
  assign n21517 = ~controllable_hgrant6 & ~n21516;
  assign n21518 = ~n14054 & ~n21517;
  assign n21519 = ~controllable_hmaster0 & ~n21518;
  assign n21520 = ~n21006 & ~n21519;
  assign n21521 = ~i_hlock8 & ~n21520;
  assign n21522 = ~n21509 & ~n21521;
  assign n21523 = ~i_hbusreq8 & ~n21522;
  assign n21524 = ~n21497 & ~n21523;
  assign n21525 = controllable_hmaster3 & ~n21524;
  assign n21526 = i_hbusreq8 & ~n21481;
  assign n21527 = i_hbusreq6 & ~n21477;
  assign n21528 = controllable_hmaster2 & ~n21060;
  assign n21529 = ~n21204 & ~n21528;
  assign n21530 = controllable_hmaster1 & ~n21529;
  assign n21531 = ~n21281 & ~n21530;
  assign n21532 = ~i_hbusreq6 & ~n21531;
  assign n21533 = ~n21527 & ~n21532;
  assign n21534 = ~controllable_hgrant6 & ~n21533;
  assign n21535 = ~n14756 & ~n21534;
  assign n21536 = controllable_hmaster0 & ~n21535;
  assign n21537 = ~n21424 & ~n21536;
  assign n21538 = ~i_hbusreq8 & ~n21537;
  assign n21539 = ~n21526 & ~n21538;
  assign n21540 = ~controllable_hmaster3 & ~n21539;
  assign n21541 = ~n21525 & ~n21540;
  assign n21542 = i_hlock7 & ~n21541;
  assign n21543 = i_hbusreq8 & ~n21491;
  assign n21544 = i_hbusreq6 & ~n21487;
  assign n21545 = controllable_hmaster2 & ~n21103;
  assign n21546 = ~n21204 & ~n21545;
  assign n21547 = controllable_hmaster1 & ~n21546;
  assign n21548 = ~n21281 & ~n21547;
  assign n21549 = ~i_hbusreq6 & ~n21548;
  assign n21550 = ~n21544 & ~n21549;
  assign n21551 = ~controllable_hgrant6 & ~n21550;
  assign n21552 = ~n14772 & ~n21551;
  assign n21553 = controllable_hmaster0 & ~n21552;
  assign n21554 = ~n21424 & ~n21553;
  assign n21555 = ~i_hbusreq8 & ~n21554;
  assign n21556 = ~n21543 & ~n21555;
  assign n21557 = ~controllable_hmaster3 & ~n21556;
  assign n21558 = ~n21525 & ~n21557;
  assign n21559 = ~i_hlock7 & ~n21558;
  assign n21560 = ~n21542 & ~n21559;
  assign n21561 = ~i_hbusreq7 & ~n21560;
  assign n21562 = ~n21496 & ~n21561;
  assign n21563 = n7924 & ~n21562;
  assign n21564 = ~n20374 & ~n21563;
  assign n21565 = ~n8214 & ~n21564;
  assign n21566 = ~n18584 & ~n20805;
  assign n21567 = controllable_hmaster1 & ~n21566;
  assign n21568 = ~n20835 & ~n21567;
  assign n21569 = i_hlock6 & ~n21568;
  assign n21570 = ~n18689 & ~n20805;
  assign n21571 = controllable_hmaster1 & ~n21570;
  assign n21572 = ~n20835 & ~n21571;
  assign n21573 = ~i_hlock6 & ~n21572;
  assign n21574 = ~n21569 & ~n21573;
  assign n21575 = ~controllable_hgrant6 & ~n21574;
  assign n21576 = ~n13894 & ~n21575;
  assign n21577 = ~controllable_hmaster0 & ~n21576;
  assign n21578 = ~n20787 & ~n21577;
  assign n21579 = ~controllable_hmaster3 & ~n21578;
  assign n21580 = ~n21474 & ~n21579;
  assign n21581 = i_hlock7 & ~n21580;
  assign n21582 = ~n20858 & ~n21577;
  assign n21583 = ~controllable_hmaster3 & ~n21582;
  assign n21584 = ~n21474 & ~n21583;
  assign n21585 = ~i_hlock7 & ~n21584;
  assign n21586 = ~n21581 & ~n21585;
  assign n21587 = i_hbusreq7 & ~n21586;
  assign n21588 = i_hbusreq8 & ~n21578;
  assign n21589 = i_hbusreq6 & ~n21574;
  assign n21590 = ~n21327 & ~n21528;
  assign n21591 = controllable_hmaster1 & ~n21590;
  assign n21592 = ~n21406 & ~n21591;
  assign n21593 = i_hlock6 & ~n21592;
  assign n21594 = ~n21327 & ~n21545;
  assign n21595 = controllable_hmaster1 & ~n21594;
  assign n21596 = ~n21406 & ~n21595;
  assign n21597 = ~i_hlock6 & ~n21596;
  assign n21598 = ~n21593 & ~n21597;
  assign n21599 = ~i_hbusreq6 & ~n21598;
  assign n21600 = ~n21589 & ~n21599;
  assign n21601 = ~controllable_hgrant6 & ~n21600;
  assign n21602 = ~n14802 & ~n21601;
  assign n21603 = ~controllable_hmaster0 & ~n21602;
  assign n21604 = ~n21287 & ~n21603;
  assign n21605 = ~i_hbusreq8 & ~n21604;
  assign n21606 = ~n21588 & ~n21605;
  assign n21607 = ~controllable_hmaster3 & ~n21606;
  assign n21608 = ~n21525 & ~n21607;
  assign n21609 = i_hlock7 & ~n21608;
  assign n21610 = i_hbusreq8 & ~n21582;
  assign n21611 = ~n21440 & ~n21603;
  assign n21612 = ~i_hbusreq8 & ~n21611;
  assign n21613 = ~n21610 & ~n21612;
  assign n21614 = ~controllable_hmaster3 & ~n21613;
  assign n21615 = ~n21525 & ~n21614;
  assign n21616 = ~i_hlock7 & ~n21615;
  assign n21617 = ~n21609 & ~n21616;
  assign n21618 = ~i_hbusreq7 & ~n21617;
  assign n21619 = ~n21587 & ~n21618;
  assign n21620 = n7924 & ~n21619;
  assign n21621 = ~n20542 & ~n21620;
  assign n21622 = n8214 & ~n21621;
  assign n21623 = ~n21565 & ~n21622;
  assign n21624 = n8202 & ~n21623;
  assign n21625 = ~n21454 & ~n21624;
  assign n21626 = n7920 & ~n21625;
  assign n21627 = ~n16336 & ~n21626;
  assign n21628 = n7728 & ~n21627;
  assign n21629 = ~n16815 & ~n17000;
  assign n21630 = ~i_hbusreq1 & ~n21629;
  assign n21631 = ~n17360 & ~n21630;
  assign n21632 = ~controllable_hgrant1 & ~n21631;
  assign n21633 = ~n14877 & ~n21632;
  assign n21634 = ~i_hbusreq3 & ~n21633;
  assign n21635 = ~n17359 & ~n21634;
  assign n21636 = ~controllable_hgrant3 & ~n21635;
  assign n21637 = ~n14876 & ~n21636;
  assign n21638 = ~i_hbusreq9 & ~n21637;
  assign n21639 = ~n17358 & ~n21638;
  assign n21640 = ~i_hbusreq4 & ~n21639;
  assign n21641 = ~n17357 & ~n21640;
  assign n21642 = ~controllable_hgrant4 & ~n21641;
  assign n21643 = ~n14875 & ~n21642;
  assign n21644 = ~i_hbusreq5 & ~n21643;
  assign n21645 = ~n17356 & ~n21644;
  assign n21646 = ~controllable_hgrant5 & ~n21645;
  assign n21647 = ~n14874 & ~n21646;
  assign n21648 = controllable_hmaster1 & ~n21647;
  assign n21649 = controllable_hmaster2 & ~n21647;
  assign n21650 = ~n16452 & ~n21649;
  assign n21651 = ~controllable_hmaster1 & ~n21650;
  assign n21652 = ~n21648 & ~n21651;
  assign n21653 = ~i_hbusreq6 & ~n21652;
  assign n21654 = ~n17355 & ~n21653;
  assign n21655 = ~controllable_hgrant6 & ~n21654;
  assign n21656 = ~n14849 & ~n21655;
  assign n21657 = controllable_hmaster0 & ~n21656;
  assign n21658 = ~n16837 & ~n21649;
  assign n21659 = ~controllable_hmaster1 & ~n21658;
  assign n21660 = ~n21648 & ~n21659;
  assign n21661 = ~i_hbusreq6 & ~n21660;
  assign n21662 = ~n18257 & ~n21661;
  assign n21663 = ~controllable_hgrant6 & ~n21662;
  assign n21664 = ~n14927 & ~n21663;
  assign n21665 = ~controllable_hmaster0 & ~n21664;
  assign n21666 = ~n21657 & ~n21665;
  assign n21667 = i_hlock8 & ~n21666;
  assign n21668 = ~n16874 & ~n21649;
  assign n21669 = ~controllable_hmaster1 & ~n21668;
  assign n21670 = ~n21648 & ~n21669;
  assign n21671 = ~i_hbusreq6 & ~n21670;
  assign n21672 = ~n18290 & ~n21671;
  assign n21673 = ~controllable_hgrant6 & ~n21672;
  assign n21674 = ~n14960 & ~n21673;
  assign n21675 = ~controllable_hmaster0 & ~n21674;
  assign n21676 = ~n21657 & ~n21675;
  assign n21677 = ~i_hlock8 & ~n21676;
  assign n21678 = ~n21667 & ~n21677;
  assign n21679 = ~i_hbusreq8 & ~n21678;
  assign n21680 = ~n18208 & ~n21679;
  assign n21681 = controllable_hmaster3 & ~n21680;
  assign n21682 = i_hlock3 & ~n16822;
  assign n21683 = ~i_hlock3 & ~n16859;
  assign n21684 = ~n21682 & ~n21683;
  assign n21685 = ~i_hbusreq3 & ~n21684;
  assign n21686 = ~n18331 & ~n21685;
  assign n21687 = ~controllable_hgrant3 & ~n21686;
  assign n21688 = ~n14999 & ~n21687;
  assign n21689 = ~i_hbusreq9 & ~n21688;
  assign n21690 = ~n18330 & ~n21689;
  assign n21691 = ~i_hbusreq4 & ~n21690;
  assign n21692 = ~n18329 & ~n21691;
  assign n21693 = ~controllable_hgrant4 & ~n21692;
  assign n21694 = ~n14998 & ~n21693;
  assign n21695 = ~i_hbusreq5 & ~n21694;
  assign n21696 = ~n18328 & ~n21695;
  assign n21697 = ~controllable_hgrant5 & ~n21696;
  assign n21698 = ~n14997 & ~n21697;
  assign n21699 = ~controllable_hmaster2 & ~n21698;
  assign n21700 = ~n16924 & ~n21699;
  assign n21701 = controllable_hmaster1 & ~n21700;
  assign n21702 = i_hlock5 & ~n16832;
  assign n21703 = ~i_hlock5 & ~n16869;
  assign n21704 = ~n21702 & ~n21703;
  assign n21705 = ~i_hbusreq5 & ~n21704;
  assign n21706 = ~n18352 & ~n21705;
  assign n21707 = ~controllable_hgrant5 & ~n21706;
  assign n21708 = ~n15020 & ~n21707;
  assign n21709 = controllable_hmaster2 & ~n21708;
  assign n21710 = i_hlock1 & ~n16818;
  assign n21711 = ~i_hlock1 & ~n16855;
  assign n21712 = ~n21710 & ~n21711;
  assign n21713 = ~i_hbusreq1 & ~n21712;
  assign n21714 = ~n18365 & ~n21713;
  assign n21715 = ~controllable_hgrant1 & ~n21714;
  assign n21716 = ~n15032 & ~n21715;
  assign n21717 = ~i_hbusreq3 & ~n21716;
  assign n21718 = ~n18364 & ~n21717;
  assign n21719 = ~controllable_hgrant3 & ~n21718;
  assign n21720 = ~n15031 & ~n21719;
  assign n21721 = ~i_hbusreq9 & ~n21720;
  assign n21722 = ~n18363 & ~n21721;
  assign n21723 = ~i_hbusreq4 & ~n21722;
  assign n21724 = ~n18362 & ~n21723;
  assign n21725 = ~controllable_hgrant4 & ~n21724;
  assign n21726 = ~n15030 & ~n21725;
  assign n21727 = ~i_hbusreq5 & ~n21726;
  assign n21728 = ~n18361 & ~n21727;
  assign n21729 = ~controllable_hgrant5 & ~n21728;
  assign n21730 = ~n15029 & ~n21729;
  assign n21731 = ~controllable_hmaster2 & ~n21730;
  assign n21732 = ~n21709 & ~n21731;
  assign n21733 = ~controllable_hmaster1 & ~n21732;
  assign n21734 = ~n21701 & ~n21733;
  assign n21735 = ~i_hbusreq6 & ~n21734;
  assign n21736 = ~n18326 & ~n21735;
  assign n21737 = ~controllable_hgrant6 & ~n21736;
  assign n21738 = ~n14995 & ~n21737;
  assign n21739 = controllable_hmaster0 & ~n21738;
  assign n21740 = ~n9379 & ~n16817;
  assign n21741 = ~i_hbusreq1 & ~n21740;
  assign n21742 = ~n18401 & ~n21741;
  assign n21743 = ~controllable_hgrant1 & ~n21742;
  assign n21744 = ~n15067 & ~n21743;
  assign n21745 = ~i_hbusreq3 & ~n21744;
  assign n21746 = ~n18400 & ~n21745;
  assign n21747 = ~controllable_hgrant3 & ~n21746;
  assign n21748 = ~n15066 & ~n21747;
  assign n21749 = ~i_hbusreq9 & ~n21748;
  assign n21750 = ~n18399 & ~n21749;
  assign n21751 = ~i_hbusreq4 & ~n21750;
  assign n21752 = ~n18398 & ~n21751;
  assign n21753 = ~controllable_hgrant4 & ~n21752;
  assign n21754 = ~n15065 & ~n21753;
  assign n21755 = ~i_hbusreq5 & ~n21754;
  assign n21756 = ~n18397 & ~n21755;
  assign n21757 = ~controllable_hgrant5 & ~n21756;
  assign n21758 = ~n15064 & ~n21757;
  assign n21759 = ~controllable_hmaster2 & ~n21758;
  assign n21760 = ~n16924 & ~n21759;
  assign n21761 = controllable_hmaster1 & ~n21760;
  assign n21762 = i_hlock4 & ~n16828;
  assign n21763 = ~i_hlock4 & ~n16865;
  assign n21764 = ~n21762 & ~n21763;
  assign n21765 = ~i_hbusreq4 & ~n21764;
  assign n21766 = ~n18425 & ~n21765;
  assign n21767 = ~controllable_hgrant4 & ~n21766;
  assign n21768 = ~n15091 & ~n21767;
  assign n21769 = ~i_hbusreq5 & ~n21768;
  assign n21770 = ~n18424 & ~n21769;
  assign n21771 = ~controllable_hgrant5 & ~n21770;
  assign n21772 = ~n15090 & ~n21771;
  assign n21773 = controllable_hmaster2 & ~n21772;
  assign n21774 = ~n16733 & ~n18454;
  assign n21775 = n7928 & ~n21774;
  assign n21776 = ~n8440 & ~n21775;
  assign n21777 = ~i_hbusreq1 & ~n21776;
  assign n21778 = ~n18442 & ~n21777;
  assign n21779 = ~controllable_hgrant1 & ~n21778;
  assign n21780 = ~n15107 & ~n21779;
  assign n21781 = ~i_hbusreq3 & ~n21780;
  assign n21782 = ~n18441 & ~n21781;
  assign n21783 = ~controllable_hgrant3 & ~n21782;
  assign n21784 = ~n15106 & ~n21783;
  assign n21785 = ~i_hbusreq9 & ~n21784;
  assign n21786 = ~n18440 & ~n21785;
  assign n21787 = ~i_hbusreq4 & ~n21786;
  assign n21788 = ~n18439 & ~n21787;
  assign n21789 = ~controllable_hgrant4 & ~n21788;
  assign n21790 = ~n15105 & ~n21789;
  assign n21791 = ~i_hbusreq5 & ~n21790;
  assign n21792 = ~n18438 & ~n21791;
  assign n21793 = ~controllable_hgrant5 & ~n21792;
  assign n21794 = ~n15104 & ~n21793;
  assign n21795 = ~controllable_hmaster2 & ~n21794;
  assign n21796 = ~n21773 & ~n21795;
  assign n21797 = ~controllable_hmaster1 & ~n21796;
  assign n21798 = ~n21761 & ~n21797;
  assign n21799 = i_hlock6 & ~n21798;
  assign n21800 = ~n16942 & ~n21759;
  assign n21801 = controllable_hmaster1 & ~n21800;
  assign n21802 = ~n21797 & ~n21801;
  assign n21803 = ~i_hlock6 & ~n21802;
  assign n21804 = ~n21799 & ~n21803;
  assign n21805 = ~i_hbusreq6 & ~n21804;
  assign n21806 = ~n18396 & ~n21805;
  assign n21807 = ~controllable_hgrant6 & ~n21806;
  assign n21808 = ~n15063 & ~n21807;
  assign n21809 = ~controllable_hmaster0 & ~n21808;
  assign n21810 = ~n21739 & ~n21809;
  assign n21811 = ~i_hbusreq8 & ~n21810;
  assign n21812 = ~n18325 & ~n21811;
  assign n21813 = ~controllable_hmaster3 & ~n21812;
  assign n21814 = ~n21681 & ~n21813;
  assign n21815 = i_hlock7 & ~n21814;
  assign n21816 = ~n16942 & ~n21699;
  assign n21817 = controllable_hmaster1 & ~n21816;
  assign n21818 = ~n21733 & ~n21817;
  assign n21819 = ~i_hbusreq6 & ~n21818;
  assign n21820 = ~n18511 & ~n21819;
  assign n21821 = ~controllable_hgrant6 & ~n21820;
  assign n21822 = ~n15152 & ~n21821;
  assign n21823 = controllable_hmaster0 & ~n21822;
  assign n21824 = ~n21809 & ~n21823;
  assign n21825 = ~i_hbusreq8 & ~n21824;
  assign n21826 = ~n18510 & ~n21825;
  assign n21827 = ~controllable_hmaster3 & ~n21826;
  assign n21828 = ~n21681 & ~n21827;
  assign n21829 = ~i_hlock7 & ~n21828;
  assign n21830 = ~n21815 & ~n21829;
  assign n21831 = ~i_hbusreq7 & ~n21830;
  assign n21832 = ~n18207 & ~n21831;
  assign n21833 = ~n7924 & ~n21832;
  assign n21834 = ~n7928 & ~n21629;
  assign n21835 = ~controllable_locked & n12782;
  assign n21836 = ~n17089 & ~n21835;
  assign n21837 = i_hlock0 & ~n21836;
  assign n21838 = ~n18716 & ~n21837;
  assign n21839 = ~i_hbusreq0 & ~n21838;
  assign n21840 = ~n17142 & ~n21839;
  assign n21841 = ~i_hbusreq2 & ~n21840;
  assign n21842 = ~n17141 & ~n21841;
  assign n21843 = ~controllable_hgrant2 & ~n21842;
  assign n21844 = ~n7814 & ~n21843;
  assign n21845 = ~n7733 & ~n21844;
  assign n21846 = ~n12615 & ~n21009;
  assign n21847 = i_hlock0 & ~n21846;
  assign n21848 = ~n18726 & ~n21847;
  assign n21849 = ~i_hbusreq0 & ~n21848;
  assign n21850 = ~n17552 & ~n21849;
  assign n21851 = ~i_hbusreq2 & ~n21850;
  assign n21852 = ~n17551 & ~n21851;
  assign n21853 = ~controllable_hgrant2 & n21852;
  assign n21854 = ~n12706 & ~n21853;
  assign n21855 = n7733 & ~n21854;
  assign n21856 = ~n21845 & ~n21855;
  assign n21857 = n7928 & ~n21856;
  assign n21858 = ~n21834 & ~n21857;
  assign n21859 = ~i_hbusreq1 & ~n21858;
  assign n21860 = ~n17549 & ~n21859;
  assign n21861 = ~controllable_hgrant1 & ~n21860;
  assign n21862 = ~n14877 & ~n21861;
  assign n21863 = ~i_hbusreq3 & ~n21862;
  assign n21864 = ~n17548 & ~n21863;
  assign n21865 = ~controllable_hgrant3 & ~n21864;
  assign n21866 = ~n14876 & ~n21865;
  assign n21867 = i_hlock9 & ~n21866;
  assign n21868 = ~n17580 & ~n21849;
  assign n21869 = ~i_hbusreq2 & ~n21868;
  assign n21870 = ~n17579 & ~n21869;
  assign n21871 = ~controllable_hgrant2 & n21870;
  assign n21872 = ~n12706 & ~n21871;
  assign n21873 = n7733 & ~n21872;
  assign n21874 = ~n21845 & ~n21873;
  assign n21875 = n7928 & ~n21874;
  assign n21876 = ~n21834 & ~n21875;
  assign n21877 = ~i_hbusreq1 & ~n21876;
  assign n21878 = ~n17578 & ~n21877;
  assign n21879 = ~controllable_hgrant1 & ~n21878;
  assign n21880 = ~n14877 & ~n21879;
  assign n21881 = ~i_hbusreq3 & ~n21880;
  assign n21882 = ~n17577 & ~n21881;
  assign n21883 = ~controllable_hgrant3 & ~n21882;
  assign n21884 = ~n14876 & ~n21883;
  assign n21885 = ~i_hlock9 & ~n21884;
  assign n21886 = ~n21867 & ~n21885;
  assign n21887 = ~i_hbusreq9 & ~n21886;
  assign n21888 = ~n17547 & ~n21887;
  assign n21889 = ~i_hbusreq4 & ~n21888;
  assign n21890 = ~n17546 & ~n21889;
  assign n21891 = ~controllable_hgrant4 & ~n21890;
  assign n21892 = ~n14875 & ~n21891;
  assign n21893 = ~i_hbusreq5 & ~n21892;
  assign n21894 = ~n17545 & ~n21893;
  assign n21895 = ~controllable_hgrant5 & ~n21894;
  assign n21896 = ~n14874 & ~n21895;
  assign n21897 = controllable_hmaster1 & ~n21896;
  assign n21898 = controllable_hmaster2 & ~n21896;
  assign n21899 = ~n16693 & ~n21898;
  assign n21900 = ~controllable_hmaster1 & ~n21899;
  assign n21901 = ~n21897 & ~n21900;
  assign n21902 = ~i_hbusreq6 & ~n21901;
  assign n21903 = ~n17544 & ~n21902;
  assign n21904 = ~controllable_hgrant6 & ~n21903;
  assign n21905 = ~n14849 & ~n21904;
  assign n21906 = controllable_hmaster0 & ~n21905;
  assign n21907 = ~n18800 & ~n21855;
  assign n21908 = n7928 & ~n21907;
  assign n21909 = ~n8265 & ~n21908;
  assign n21910 = ~i_hbusreq1 & ~n21909;
  assign n21911 = ~n18791 & ~n21910;
  assign n21912 = ~controllable_hgrant1 & ~n21911;
  assign n21913 = ~n12681 & ~n21912;
  assign n21914 = ~i_hbusreq3 & ~n21913;
  assign n21915 = ~n18790 & ~n21914;
  assign n21916 = ~controllable_hgrant3 & ~n21915;
  assign n21917 = ~n12679 & ~n21916;
  assign n21918 = i_hlock9 & ~n21917;
  assign n21919 = ~n18800 & ~n21873;
  assign n21920 = n7928 & ~n21919;
  assign n21921 = ~n8265 & ~n21920;
  assign n21922 = ~i_hbusreq1 & ~n21921;
  assign n21923 = ~n18814 & ~n21922;
  assign n21924 = ~controllable_hgrant1 & ~n21923;
  assign n21925 = ~n12681 & ~n21924;
  assign n21926 = ~i_hbusreq3 & ~n21925;
  assign n21927 = ~n18813 & ~n21926;
  assign n21928 = ~controllable_hgrant3 & ~n21927;
  assign n21929 = ~n12679 & ~n21928;
  assign n21930 = ~i_hlock9 & ~n21929;
  assign n21931 = ~n21918 & ~n21930;
  assign n21932 = ~i_hbusreq9 & ~n21931;
  assign n21933 = ~n18789 & ~n21932;
  assign n21934 = ~i_hbusreq4 & ~n21933;
  assign n21935 = ~n18788 & ~n21934;
  assign n21936 = ~controllable_hgrant4 & ~n21935;
  assign n21937 = ~n13524 & ~n21936;
  assign n21938 = ~i_hbusreq5 & ~n21937;
  assign n21939 = ~n18787 & ~n21938;
  assign n21940 = ~controllable_hgrant5 & ~n21939;
  assign n21941 = ~n13522 & ~n21940;
  assign n21942 = ~controllable_hmaster2 & ~n21941;
  assign n21943 = ~n21898 & ~n21942;
  assign n21944 = ~controllable_hmaster1 & ~n21943;
  assign n21945 = ~n21897 & ~n21944;
  assign n21946 = ~i_hbusreq6 & ~n21945;
  assign n21947 = ~n18786 & ~n21946;
  assign n21948 = ~controllable_hgrant6 & ~n21947;
  assign n21949 = ~n14927 & ~n21948;
  assign n21950 = ~controllable_hmaster0 & ~n21949;
  assign n21951 = ~n21906 & ~n21950;
  assign n21952 = i_hlock8 & ~n21951;
  assign n21953 = ~n8297 & ~n21908;
  assign n21954 = ~i_hbusreq1 & ~n21953;
  assign n21955 = ~n18854 & ~n21954;
  assign n21956 = ~controllable_hgrant1 & ~n21955;
  assign n21957 = ~n12730 & ~n21956;
  assign n21958 = ~i_hbusreq3 & ~n21957;
  assign n21959 = ~n18853 & ~n21958;
  assign n21960 = ~controllable_hgrant3 & ~n21959;
  assign n21961 = ~n12728 & ~n21960;
  assign n21962 = i_hlock9 & ~n21961;
  assign n21963 = ~n8297 & ~n21920;
  assign n21964 = ~i_hbusreq1 & ~n21963;
  assign n21965 = ~n18866 & ~n21964;
  assign n21966 = ~controllable_hgrant1 & ~n21965;
  assign n21967 = ~n12730 & ~n21966;
  assign n21968 = ~i_hbusreq3 & ~n21967;
  assign n21969 = ~n18865 & ~n21968;
  assign n21970 = ~controllable_hgrant3 & ~n21969;
  assign n21971 = ~n12728 & ~n21970;
  assign n21972 = ~i_hlock9 & ~n21971;
  assign n21973 = ~n21962 & ~n21972;
  assign n21974 = ~i_hbusreq9 & ~n21973;
  assign n21975 = ~n18852 & ~n21974;
  assign n21976 = ~i_hbusreq4 & ~n21975;
  assign n21977 = ~n18851 & ~n21976;
  assign n21978 = ~controllable_hgrant4 & ~n21977;
  assign n21979 = ~n13577 & ~n21978;
  assign n21980 = ~i_hbusreq5 & ~n21979;
  assign n21981 = ~n18850 & ~n21980;
  assign n21982 = ~controllable_hgrant5 & ~n21981;
  assign n21983 = ~n13575 & ~n21982;
  assign n21984 = ~controllable_hmaster2 & ~n21983;
  assign n21985 = ~n21898 & ~n21984;
  assign n21986 = ~controllable_hmaster1 & ~n21985;
  assign n21987 = ~n21897 & ~n21986;
  assign n21988 = ~i_hbusreq6 & ~n21987;
  assign n21989 = ~n18849 & ~n21988;
  assign n21990 = ~controllable_hgrant6 & ~n21989;
  assign n21991 = ~n14960 & ~n21990;
  assign n21992 = ~controllable_hmaster0 & ~n21991;
  assign n21993 = ~n21906 & ~n21992;
  assign n21994 = ~i_hlock8 & ~n21993;
  assign n21995 = ~n21952 & ~n21994;
  assign n21996 = ~i_hbusreq8 & ~n21995;
  assign n21997 = ~n18714 & ~n21996;
  assign n21998 = controllable_hmaster3 & ~n21997;
  assign n21999 = controllable_hmaster2 & ~n21941;
  assign n22000 = i_hlock3 & ~n21913;
  assign n22001 = ~i_hlock3 & ~n21957;
  assign n22002 = ~n22000 & ~n22001;
  assign n22003 = ~i_hbusreq3 & ~n22002;
  assign n22004 = ~n18909 & ~n22003;
  assign n22005 = ~controllable_hgrant3 & ~n22004;
  assign n22006 = ~n14999 & ~n22005;
  assign n22007 = i_hlock9 & ~n22006;
  assign n22008 = i_hlock3 & ~n21925;
  assign n22009 = ~i_hlock3 & ~n21967;
  assign n22010 = ~n22008 & ~n22009;
  assign n22011 = ~i_hbusreq3 & ~n22010;
  assign n22012 = ~n18918 & ~n22011;
  assign n22013 = ~controllable_hgrant3 & ~n22012;
  assign n22014 = ~n14999 & ~n22013;
  assign n22015 = ~i_hlock9 & ~n22014;
  assign n22016 = ~n22007 & ~n22015;
  assign n22017 = ~i_hbusreq9 & ~n22016;
  assign n22018 = ~n18908 & ~n22017;
  assign n22019 = ~i_hbusreq4 & ~n22018;
  assign n22020 = ~n18907 & ~n22019;
  assign n22021 = ~controllable_hgrant4 & ~n22020;
  assign n22022 = ~n14998 & ~n22021;
  assign n22023 = ~i_hbusreq5 & ~n22022;
  assign n22024 = ~n18906 & ~n22023;
  assign n22025 = ~controllable_hgrant5 & ~n22024;
  assign n22026 = ~n14997 & ~n22025;
  assign n22027 = ~controllable_hmaster2 & ~n22026;
  assign n22028 = ~n21999 & ~n22027;
  assign n22029 = controllable_hmaster1 & ~n22028;
  assign n22030 = i_hlock5 & ~n21937;
  assign n22031 = ~i_hlock5 & ~n21979;
  assign n22032 = ~n22030 & ~n22031;
  assign n22033 = ~i_hbusreq5 & ~n22032;
  assign n22034 = ~n18941 & ~n22033;
  assign n22035 = ~controllable_hgrant5 & ~n22034;
  assign n22036 = ~n15020 & ~n22035;
  assign n22037 = controllable_hmaster2 & ~n22036;
  assign n22038 = i_hlock1 & ~n21909;
  assign n22039 = ~i_hlock1 & ~n21953;
  assign n22040 = ~n22038 & ~n22039;
  assign n22041 = ~i_hbusreq1 & ~n22040;
  assign n22042 = ~n18954 & ~n22041;
  assign n22043 = ~controllable_hgrant1 & ~n22042;
  assign n22044 = ~n15032 & ~n22043;
  assign n22045 = ~i_hbusreq3 & ~n22044;
  assign n22046 = ~n18953 & ~n22045;
  assign n22047 = ~controllable_hgrant3 & ~n22046;
  assign n22048 = ~n15031 & ~n22047;
  assign n22049 = i_hlock9 & ~n22048;
  assign n22050 = i_hlock1 & ~n21921;
  assign n22051 = ~i_hlock1 & ~n21963;
  assign n22052 = ~n22050 & ~n22051;
  assign n22053 = ~i_hbusreq1 & ~n22052;
  assign n22054 = ~n18968 & ~n22053;
  assign n22055 = ~controllable_hgrant1 & ~n22054;
  assign n22056 = ~n15032 & ~n22055;
  assign n22057 = ~i_hbusreq3 & ~n22056;
  assign n22058 = ~n18967 & ~n22057;
  assign n22059 = ~controllable_hgrant3 & ~n22058;
  assign n22060 = ~n15031 & ~n22059;
  assign n22061 = ~i_hlock9 & ~n22060;
  assign n22062 = ~n22049 & ~n22061;
  assign n22063 = ~i_hbusreq9 & ~n22062;
  assign n22064 = ~n18952 & ~n22063;
  assign n22065 = ~i_hbusreq4 & ~n22064;
  assign n22066 = ~n18951 & ~n22065;
  assign n22067 = ~controllable_hgrant4 & ~n22066;
  assign n22068 = ~n15030 & ~n22067;
  assign n22069 = ~i_hbusreq5 & ~n22068;
  assign n22070 = ~n18950 & ~n22069;
  assign n22071 = ~controllable_hgrant5 & ~n22070;
  assign n22072 = ~n15029 & ~n22071;
  assign n22073 = ~controllable_hmaster2 & ~n22072;
  assign n22074 = ~n22037 & ~n22073;
  assign n22075 = ~controllable_hmaster1 & ~n22074;
  assign n22076 = ~n22029 & ~n22075;
  assign n22077 = ~i_hbusreq6 & ~n22076;
  assign n22078 = ~n18904 & ~n22077;
  assign n22079 = ~controllable_hgrant6 & ~n22078;
  assign n22080 = ~n14995 & ~n22079;
  assign n22081 = controllable_hmaster0 & ~n22080;
  assign n22082 = ~n9379 & ~n21908;
  assign n22083 = ~i_hbusreq1 & ~n22082;
  assign n22084 = ~n19006 & ~n22083;
  assign n22085 = ~controllable_hgrant1 & ~n22084;
  assign n22086 = ~n15067 & ~n22085;
  assign n22087 = ~i_hbusreq3 & ~n22086;
  assign n22088 = ~n19005 & ~n22087;
  assign n22089 = ~controllable_hgrant3 & ~n22088;
  assign n22090 = ~n15066 & ~n22089;
  assign n22091 = i_hlock9 & ~n22090;
  assign n22092 = ~n9379 & ~n21920;
  assign n22093 = ~i_hbusreq1 & ~n22092;
  assign n22094 = ~n19018 & ~n22093;
  assign n22095 = ~controllable_hgrant1 & ~n22094;
  assign n22096 = ~n15067 & ~n22095;
  assign n22097 = ~i_hbusreq3 & ~n22096;
  assign n22098 = ~n19017 & ~n22097;
  assign n22099 = ~controllable_hgrant3 & ~n22098;
  assign n22100 = ~n15066 & ~n22099;
  assign n22101 = ~i_hlock9 & ~n22100;
  assign n22102 = ~n22091 & ~n22101;
  assign n22103 = ~i_hbusreq9 & ~n22102;
  assign n22104 = ~n19004 & ~n22103;
  assign n22105 = ~i_hbusreq4 & ~n22104;
  assign n22106 = ~n19003 & ~n22105;
  assign n22107 = ~controllable_hgrant4 & ~n22106;
  assign n22108 = ~n15065 & ~n22107;
  assign n22109 = ~i_hbusreq5 & ~n22108;
  assign n22110 = ~n19002 & ~n22109;
  assign n22111 = ~controllable_hgrant5 & ~n22110;
  assign n22112 = ~n15064 & ~n22111;
  assign n22113 = ~controllable_hmaster2 & ~n22112;
  assign n22114 = ~n21999 & ~n22113;
  assign n22115 = controllable_hmaster1 & ~n22114;
  assign n22116 = i_hlock4 & ~n21933;
  assign n22117 = ~i_hlock4 & ~n21975;
  assign n22118 = ~n22116 & ~n22117;
  assign n22119 = ~i_hbusreq4 & ~n22118;
  assign n22120 = ~n19044 & ~n22119;
  assign n22121 = ~controllable_hgrant4 & ~n22120;
  assign n22122 = ~n15091 & ~n22121;
  assign n22123 = ~i_hbusreq5 & ~n22122;
  assign n22124 = ~n19043 & ~n22123;
  assign n22125 = ~controllable_hgrant5 & ~n22124;
  assign n22126 = ~n15090 & ~n22125;
  assign n22127 = controllable_hmaster2 & ~n22126;
  assign n22128 = ~i_hbusreq0 & ~n17480;
  assign n22129 = ~n17552 & ~n22128;
  assign n22130 = ~i_hbusreq2 & ~n22129;
  assign n22131 = ~n17551 & ~n22130;
  assign n22132 = ~controllable_hgrant2 & n22131;
  assign n22133 = ~n7814 & ~n22132;
  assign n22134 = n7733 & ~n22133;
  assign n22135 = ~n19072 & ~n22134;
  assign n22136 = n7928 & ~n22135;
  assign n22137 = ~n8440 & ~n22136;
  assign n22138 = ~i_hbusreq1 & ~n22137;
  assign n22139 = ~n19061 & ~n22138;
  assign n22140 = ~controllable_hgrant1 & ~n22139;
  assign n22141 = ~n15107 & ~n22140;
  assign n22142 = ~i_hbusreq3 & ~n22141;
  assign n22143 = ~n19060 & ~n22142;
  assign n22144 = ~controllable_hgrant3 & ~n22143;
  assign n22145 = ~n15106 & ~n22144;
  assign n22146 = i_hlock9 & ~n22145;
  assign n22147 = ~n17483 & ~n19072;
  assign n22148 = n7928 & ~n22147;
  assign n22149 = ~n8440 & ~n22148;
  assign n22150 = ~i_hbusreq1 & ~n22149;
  assign n22151 = ~n19099 & ~n22150;
  assign n22152 = ~controllable_hgrant1 & ~n22151;
  assign n22153 = ~n15107 & ~n22152;
  assign n22154 = ~i_hbusreq3 & ~n22153;
  assign n22155 = ~n19098 & ~n22154;
  assign n22156 = ~controllable_hgrant3 & ~n22155;
  assign n22157 = ~n15106 & ~n22156;
  assign n22158 = ~i_hlock9 & ~n22157;
  assign n22159 = ~n22146 & ~n22158;
  assign n22160 = ~i_hbusreq9 & ~n22159;
  assign n22161 = ~n19059 & ~n22160;
  assign n22162 = ~i_hbusreq4 & ~n22161;
  assign n22163 = ~n19058 & ~n22162;
  assign n22164 = ~controllable_hgrant4 & ~n22163;
  assign n22165 = ~n15105 & ~n22164;
  assign n22166 = ~i_hbusreq5 & ~n22165;
  assign n22167 = ~n19057 & ~n22166;
  assign n22168 = ~controllable_hgrant5 & ~n22167;
  assign n22169 = ~n15104 & ~n22168;
  assign n22170 = ~controllable_hmaster2 & ~n22169;
  assign n22171 = ~n22127 & ~n22170;
  assign n22172 = ~controllable_hmaster1 & ~n22171;
  assign n22173 = ~n22115 & ~n22172;
  assign n22174 = i_hlock6 & ~n22173;
  assign n22175 = controllable_hmaster2 & ~n21983;
  assign n22176 = ~n22113 & ~n22175;
  assign n22177 = controllable_hmaster1 & ~n22176;
  assign n22178 = ~n22172 & ~n22177;
  assign n22179 = ~i_hlock6 & ~n22178;
  assign n22180 = ~n22174 & ~n22179;
  assign n22181 = ~i_hbusreq6 & ~n22180;
  assign n22182 = ~n19001 & ~n22181;
  assign n22183 = ~controllable_hgrant6 & ~n22182;
  assign n22184 = ~n15063 & ~n22183;
  assign n22185 = ~controllable_hmaster0 & ~n22184;
  assign n22186 = ~n22081 & ~n22185;
  assign n22187 = ~i_hbusreq8 & ~n22186;
  assign n22188 = ~n18903 & ~n22187;
  assign n22189 = ~controllable_hmaster3 & ~n22188;
  assign n22190 = ~n21998 & ~n22189;
  assign n22191 = i_hlock7 & ~n22190;
  assign n22192 = ~n22027 & ~n22175;
  assign n22193 = controllable_hmaster1 & ~n22192;
  assign n22194 = ~n22075 & ~n22193;
  assign n22195 = ~i_hbusreq6 & ~n22194;
  assign n22196 = ~n19152 & ~n22195;
  assign n22197 = ~controllable_hgrant6 & ~n22196;
  assign n22198 = ~n15152 & ~n22197;
  assign n22199 = controllable_hmaster0 & ~n22198;
  assign n22200 = ~n22185 & ~n22199;
  assign n22201 = ~i_hbusreq8 & ~n22200;
  assign n22202 = ~n19151 & ~n22201;
  assign n22203 = ~controllable_hmaster3 & ~n22202;
  assign n22204 = ~n21998 & ~n22203;
  assign n22205 = ~i_hlock7 & ~n22204;
  assign n22206 = ~n22191 & ~n22205;
  assign n22207 = ~i_hbusreq7 & ~n22206;
  assign n22208 = ~n18713 & ~n22207;
  assign n22209 = n7924 & ~n22208;
  assign n22210 = ~n21833 & ~n22209;
  assign n22211 = n7920 & ~n22210;
  assign n22212 = ~n16336 & ~n22211;
  assign n22213 = ~n7728 & ~n22212;
  assign n22214 = ~n21628 & ~n22213;
  assign n22215 = ~n7723 & ~n22214;
  assign n22216 = ~n20611 & ~n22215;
  assign n22217 = ~n7714 & ~n22216;
  assign n22218 = ~n20610 & ~n22217;
  assign n22219 = ~n7705 & ~n22218;
  assign n22220 = ~n17313 & ~n22219;
  assign n22221 = n7808 & ~n22220;
  assign n22222 = ~n16346 & ~n22221;
  assign n22223 = n8195 & ~n22222;
  assign n22224 = ~n8196 & ~n22223;
  assign n22225 = ~n8193 & ~n22224;
  assign n22226 = ~n9900 & ~n16336;
  assign n22227 = ~n7723 & ~n22226;
  assign n22228 = ~n9899 & ~n22227;
  assign n22229 = n7714 & ~n22228;
  assign n22230 = ~n16342 & ~n22229;
  assign n22231 = ~n7705 & ~n22230;
  assign n22232 = ~n9898 & ~n22231;
  assign n22233 = ~n7808 & ~n22232;
  assign n22234 = controllable_hgrant6 & ~n9912;
  assign n22235 = controllable_hmaster2 & ~n18131;
  assign n22236 = ~controllable_hmaster1 & ~n22235;
  assign n22237 = ~controllable_hmaster1 & ~n22236;
  assign n22238 = ~controllable_hgrant6 & ~n22237;
  assign n22239 = ~n22234 & ~n22238;
  assign n22240 = controllable_hmaster0 & ~n22239;
  assign n22241 = controllable_hmaster0 & ~n22240;
  assign n22242 = ~controllable_hmaster3 & ~n22241;
  assign n22243 = ~controllable_hmaster3 & ~n22242;
  assign n22244 = i_hbusreq7 & ~n22243;
  assign n22245 = i_hbusreq8 & ~n22241;
  assign n22246 = controllable_hgrant6 & ~n9924;
  assign n22247 = i_hbusreq6 & ~n22237;
  assign n22248 = controllable_hmaster2 & ~n21709;
  assign n22249 = ~controllable_hmaster1 & ~n22248;
  assign n22250 = ~controllable_hmaster1 & ~n22249;
  assign n22251 = ~i_hbusreq6 & ~n22250;
  assign n22252 = ~n22247 & ~n22251;
  assign n22253 = ~controllable_hgrant6 & ~n22252;
  assign n22254 = ~n22246 & ~n22253;
  assign n22255 = controllable_hmaster0 & ~n22254;
  assign n22256 = controllable_hmaster0 & ~n22255;
  assign n22257 = ~i_hbusreq8 & ~n22256;
  assign n22258 = ~n22245 & ~n22257;
  assign n22259 = ~controllable_hmaster3 & ~n22258;
  assign n22260 = ~controllable_hmaster3 & ~n22259;
  assign n22261 = ~i_hbusreq7 & ~n22260;
  assign n22262 = ~n22244 & ~n22261;
  assign n22263 = ~n8214 & ~n22262;
  assign n22264 = controllable_hgrant6 & ~n9936;
  assign n22265 = controllable_hmaster2 & ~n18169;
  assign n22266 = ~controllable_hmaster1 & ~n22265;
  assign n22267 = ~controllable_hmaster1 & ~n22266;
  assign n22268 = ~controllable_hgrant6 & ~n22267;
  assign n22269 = ~n22264 & ~n22268;
  assign n22270 = ~controllable_hmaster0 & ~n22269;
  assign n22271 = ~controllable_hmaster0 & ~n22270;
  assign n22272 = ~controllable_hmaster3 & ~n22271;
  assign n22273 = ~controllable_hmaster3 & ~n22272;
  assign n22274 = i_hbusreq7 & ~n22273;
  assign n22275 = i_hbusreq8 & ~n22271;
  assign n22276 = controllable_hgrant6 & ~n9948;
  assign n22277 = i_hbusreq6 & ~n22267;
  assign n22278 = controllable_hmaster2 & ~n21773;
  assign n22279 = ~controllable_hmaster1 & ~n22278;
  assign n22280 = ~controllable_hmaster1 & ~n22279;
  assign n22281 = ~i_hbusreq6 & ~n22280;
  assign n22282 = ~n22277 & ~n22281;
  assign n22283 = ~controllable_hgrant6 & ~n22282;
  assign n22284 = ~n22276 & ~n22283;
  assign n22285 = ~controllable_hmaster0 & ~n22284;
  assign n22286 = ~controllable_hmaster0 & ~n22285;
  assign n22287 = ~i_hbusreq8 & ~n22286;
  assign n22288 = ~n22275 & ~n22287;
  assign n22289 = ~controllable_hmaster3 & ~n22288;
  assign n22290 = ~controllable_hmaster3 & ~n22289;
  assign n22291 = ~i_hbusreq7 & ~n22290;
  assign n22292 = ~n22274 & ~n22291;
  assign n22293 = n8214 & ~n22292;
  assign n22294 = ~n22263 & ~n22293;
  assign n22295 = ~n8202 & ~n22294;
  assign n22296 = controllable_hgrant6 & ~n9962;
  assign n22297 = ~controllable_hmaster2 & ~n18123;
  assign n22298 = controllable_hmaster1 & ~n22297;
  assign n22299 = controllable_hmaster1 & ~n22298;
  assign n22300 = ~controllable_hgrant6 & ~n22299;
  assign n22301 = ~n22296 & ~n22300;
  assign n22302 = controllable_hmaster0 & ~n22301;
  assign n22303 = controllable_hmaster0 & ~n22302;
  assign n22304 = ~controllable_hmaster3 & ~n22303;
  assign n22305 = ~controllable_hmaster3 & ~n22304;
  assign n22306 = i_hbusreq7 & ~n22305;
  assign n22307 = i_hbusreq8 & ~n22303;
  assign n22308 = controllable_hgrant6 & ~n9974;
  assign n22309 = i_hbusreq6 & ~n22299;
  assign n22310 = ~controllable_hmaster2 & ~n21699;
  assign n22311 = controllable_hmaster1 & ~n22310;
  assign n22312 = controllable_hmaster1 & ~n22311;
  assign n22313 = ~i_hbusreq6 & ~n22312;
  assign n22314 = ~n22309 & ~n22313;
  assign n22315 = ~controllable_hgrant6 & ~n22314;
  assign n22316 = ~n22308 & ~n22315;
  assign n22317 = controllable_hmaster0 & ~n22316;
  assign n22318 = controllable_hmaster0 & ~n22317;
  assign n22319 = ~i_hbusreq8 & ~n22318;
  assign n22320 = ~n22307 & ~n22319;
  assign n22321 = ~controllable_hmaster3 & ~n22320;
  assign n22322 = ~controllable_hmaster3 & ~n22321;
  assign n22323 = ~i_hbusreq7 & ~n22322;
  assign n22324 = ~n22306 & ~n22323;
  assign n22325 = ~n8214 & ~n22324;
  assign n22326 = controllable_hgrant6 & ~n9986;
  assign n22327 = ~controllable_hmaster2 & ~n18159;
  assign n22328 = controllable_hmaster1 & ~n22327;
  assign n22329 = controllable_hmaster1 & ~n22328;
  assign n22330 = ~controllable_hgrant6 & ~n22329;
  assign n22331 = ~n22326 & ~n22330;
  assign n22332 = ~controllable_hmaster0 & ~n22331;
  assign n22333 = ~controllable_hmaster0 & ~n22332;
  assign n22334 = ~controllable_hmaster3 & ~n22333;
  assign n22335 = ~controllable_hmaster3 & ~n22334;
  assign n22336 = i_hbusreq7 & ~n22335;
  assign n22337 = i_hbusreq8 & ~n22333;
  assign n22338 = controllable_hgrant6 & ~n9998;
  assign n22339 = i_hbusreq6 & ~n22329;
  assign n22340 = ~controllable_hmaster2 & ~n21759;
  assign n22341 = controllable_hmaster1 & ~n22340;
  assign n22342 = controllable_hmaster1 & ~n22341;
  assign n22343 = ~i_hbusreq6 & ~n22342;
  assign n22344 = ~n22339 & ~n22343;
  assign n22345 = ~controllable_hgrant6 & ~n22344;
  assign n22346 = ~n22338 & ~n22345;
  assign n22347 = ~controllable_hmaster0 & ~n22346;
  assign n22348 = ~controllable_hmaster0 & ~n22347;
  assign n22349 = ~i_hbusreq8 & ~n22348;
  assign n22350 = ~n22337 & ~n22349;
  assign n22351 = ~controllable_hmaster3 & ~n22350;
  assign n22352 = ~controllable_hmaster3 & ~n22351;
  assign n22353 = ~i_hbusreq7 & ~n22352;
  assign n22354 = ~n22336 & ~n22353;
  assign n22355 = n8214 & ~n22354;
  assign n22356 = ~n22325 & ~n22355;
  assign n22357 = n8202 & ~n22356;
  assign n22358 = ~n22295 & ~n22357;
  assign n22359 = n7920 & ~n22358;
  assign n22360 = ~n9909 & ~n22359;
  assign n22361 = n7728 & ~n22360;
  assign n22362 = ~n7743 & ~n22242;
  assign n22363 = i_hbusreq7 & ~n22362;
  assign n22364 = ~n7779 & ~n22259;
  assign n22365 = ~i_hbusreq7 & ~n22364;
  assign n22366 = ~n22363 & ~n22365;
  assign n22367 = ~n8214 & ~n22366;
  assign n22368 = ~n7743 & ~n22272;
  assign n22369 = i_hbusreq7 & ~n22368;
  assign n22370 = ~n7779 & ~n22289;
  assign n22371 = ~i_hbusreq7 & ~n22370;
  assign n22372 = ~n22369 & ~n22371;
  assign n22373 = n8214 & ~n22372;
  assign n22374 = ~n22367 & ~n22373;
  assign n22375 = ~n8202 & ~n22374;
  assign n22376 = ~n7743 & ~n22304;
  assign n22377 = i_hbusreq7 & ~n22376;
  assign n22378 = ~n7779 & ~n22321;
  assign n22379 = ~i_hbusreq7 & ~n22378;
  assign n22380 = ~n22377 & ~n22379;
  assign n22381 = ~n8214 & ~n22380;
  assign n22382 = ~n7743 & ~n22334;
  assign n22383 = i_hbusreq7 & ~n22382;
  assign n22384 = ~n7779 & ~n22351;
  assign n22385 = ~i_hbusreq7 & ~n22384;
  assign n22386 = ~n22383 & ~n22385;
  assign n22387 = n8214 & ~n22386;
  assign n22388 = ~n22381 & ~n22387;
  assign n22389 = n8202 & ~n22388;
  assign n22390 = ~n22375 & ~n22389;
  assign n22391 = n7920 & ~n22390;
  assign n22392 = ~n10014 & ~n22391;
  assign n22393 = ~n7728 & ~n22392;
  assign n22394 = ~n22361 & ~n22393;
  assign n22395 = ~n7723 & ~n22394;
  assign n22396 = ~n7723 & ~n22395;
  assign n22397 = ~n7714 & ~n22396;
  assign n22398 = ~n7714 & ~n22397;
  assign n22399 = n7705 & ~n22398;
  assign n22400 = ~n8988 & ~n18131;
  assign n22401 = ~controllable_hmaster1 & ~n22400;
  assign n22402 = ~n10053 & ~n22401;
  assign n22403 = ~controllable_hgrant6 & ~n22402;
  assign n22404 = ~n15193 & ~n22403;
  assign n22405 = controllable_hmaster0 & ~n22404;
  assign n22406 = ~n9099 & ~n22405;
  assign n22407 = ~controllable_hmaster3 & ~n22406;
  assign n22408 = ~n13651 & ~n22407;
  assign n22409 = i_hbusreq7 & ~n22408;
  assign n22410 = i_hbusreq8 & ~n22406;
  assign n22411 = i_hbusreq6 & ~n22402;
  assign n22412 = ~n9024 & ~n21709;
  assign n22413 = ~controllable_hmaster1 & ~n22412;
  assign n22414 = ~n10064 & ~n22413;
  assign n22415 = ~i_hbusreq6 & ~n22414;
  assign n22416 = ~n22411 & ~n22415;
  assign n22417 = ~controllable_hgrant6 & ~n22416;
  assign n22418 = ~n15206 & ~n22417;
  assign n22419 = controllable_hmaster0 & ~n22418;
  assign n22420 = ~n9127 & ~n22419;
  assign n22421 = ~i_hbusreq8 & ~n22420;
  assign n22422 = ~n22410 & ~n22421;
  assign n22423 = ~controllable_hmaster3 & ~n22422;
  assign n22424 = ~n13662 & ~n22423;
  assign n22425 = ~i_hbusreq7 & ~n22424;
  assign n22426 = ~n22409 & ~n22425;
  assign n22427 = ~n7924 & ~n22426;
  assign n22428 = i_hlock5 & ~n17773;
  assign n22429 = ~i_hlock5 & ~n17791;
  assign n22430 = ~n22428 & ~n22429;
  assign n22431 = ~controllable_hgrant5 & ~n22430;
  assign n22432 = ~n13865 & ~n22431;
  assign n22433 = controllable_hmaster2 & ~n22432;
  assign n22434 = ~n13189 & ~n22433;
  assign n22435 = ~controllable_hmaster1 & ~n22434;
  assign n22436 = ~n15194 & ~n22435;
  assign n22437 = ~controllable_hgrant6 & ~n22436;
  assign n22438 = ~n15193 & ~n22437;
  assign n22439 = controllable_hmaster0 & ~n22438;
  assign n22440 = ~n13682 & ~n22439;
  assign n22441 = ~controllable_hmaster3 & ~n22440;
  assign n22442 = ~n13672 & ~n22441;
  assign n22443 = i_hbusreq7 & ~n22442;
  assign n22444 = i_hbusreq8 & ~n22440;
  assign n22445 = i_hbusreq6 & ~n22436;
  assign n22446 = i_hbusreq5 & ~n22430;
  assign n22447 = i_hlock5 & ~n17846;
  assign n22448 = ~i_hlock5 & ~n17882;
  assign n22449 = ~n22447 & ~n22448;
  assign n22450 = ~i_hbusreq5 & ~n22449;
  assign n22451 = ~n22446 & ~n22450;
  assign n22452 = ~controllable_hgrant5 & ~n22451;
  assign n22453 = ~n15020 & ~n22452;
  assign n22454 = controllable_hmaster2 & ~n22453;
  assign n22455 = ~n13702 & ~n22454;
  assign n22456 = ~controllable_hmaster1 & ~n22455;
  assign n22457 = ~n15208 & ~n22456;
  assign n22458 = ~i_hbusreq6 & ~n22457;
  assign n22459 = ~n22445 & ~n22458;
  assign n22460 = ~controllable_hgrant6 & ~n22459;
  assign n22461 = ~n15206 & ~n22460;
  assign n22462 = controllable_hmaster0 & ~n22461;
  assign n22463 = ~n13728 & ~n22462;
  assign n22464 = ~i_hbusreq8 & ~n22463;
  assign n22465 = ~n22444 & ~n22464;
  assign n22466 = ~controllable_hmaster3 & ~n22465;
  assign n22467 = ~n13714 & ~n22466;
  assign n22468 = ~i_hbusreq7 & ~n22467;
  assign n22469 = ~n22443 & ~n22468;
  assign n22470 = n7924 & ~n22469;
  assign n22471 = ~n22427 & ~n22470;
  assign n22472 = ~n8214 & ~n22471;
  assign n22473 = ~n8988 & ~n18169;
  assign n22474 = ~controllable_hmaster1 & ~n22473;
  assign n22475 = ~n10053 & ~n22474;
  assign n22476 = ~controllable_hgrant6 & ~n22475;
  assign n22477 = ~n15241 & ~n22476;
  assign n22478 = ~controllable_hmaster0 & ~n22477;
  assign n22479 = ~n9152 & ~n22478;
  assign n22480 = ~controllable_hmaster3 & ~n22479;
  assign n22481 = ~n13651 & ~n22480;
  assign n22482 = i_hbusreq7 & ~n22481;
  assign n22483 = i_hbusreq8 & ~n22479;
  assign n22484 = i_hbusreq6 & ~n22475;
  assign n22485 = ~n9024 & ~n21773;
  assign n22486 = ~controllable_hmaster1 & ~n22485;
  assign n22487 = ~n10064 & ~n22486;
  assign n22488 = ~i_hbusreq6 & ~n22487;
  assign n22489 = ~n22484 & ~n22488;
  assign n22490 = ~controllable_hgrant6 & ~n22489;
  assign n22491 = ~n15253 & ~n22490;
  assign n22492 = ~controllable_hmaster0 & ~n22491;
  assign n22493 = ~n9162 & ~n22492;
  assign n22494 = ~i_hbusreq8 & ~n22493;
  assign n22495 = ~n22483 & ~n22494;
  assign n22496 = ~controllable_hmaster3 & ~n22495;
  assign n22497 = ~n13662 & ~n22496;
  assign n22498 = ~i_hbusreq7 & ~n22497;
  assign n22499 = ~n22482 & ~n22498;
  assign n22500 = ~n7924 & ~n22499;
  assign n22501 = i_hlock4 & ~n17771;
  assign n22502 = ~i_hlock4 & ~n17789;
  assign n22503 = ~n22501 & ~n22502;
  assign n22504 = ~controllable_hgrant4 & ~n22503;
  assign n22505 = ~n13912 & ~n22504;
  assign n22506 = ~controllable_hgrant5 & ~n22505;
  assign n22507 = ~n13911 & ~n22506;
  assign n22508 = controllable_hmaster2 & ~n22507;
  assign n22509 = ~n13189 & ~n22508;
  assign n22510 = ~controllable_hmaster1 & ~n22509;
  assign n22511 = ~n15194 & ~n22510;
  assign n22512 = ~controllable_hgrant6 & ~n22511;
  assign n22513 = ~n15241 & ~n22512;
  assign n22514 = ~controllable_hmaster0 & ~n22513;
  assign n22515 = ~n13765 & ~n22514;
  assign n22516 = ~controllable_hmaster3 & ~n22515;
  assign n22517 = ~n13672 & ~n22516;
  assign n22518 = i_hbusreq7 & ~n22517;
  assign n22519 = i_hbusreq8 & ~n22515;
  assign n22520 = i_hbusreq6 & ~n22511;
  assign n22521 = i_hbusreq5 & ~n22505;
  assign n22522 = i_hbusreq4 & ~n22503;
  assign n22523 = i_hlock4 & ~n17842;
  assign n22524 = ~i_hlock4 & ~n17878;
  assign n22525 = ~n22523 & ~n22524;
  assign n22526 = ~i_hbusreq4 & ~n22525;
  assign n22527 = ~n22522 & ~n22526;
  assign n22528 = ~controllable_hgrant4 & ~n22527;
  assign n22529 = ~n15091 & ~n22528;
  assign n22530 = ~i_hbusreq5 & ~n22529;
  assign n22531 = ~n22521 & ~n22530;
  assign n22532 = ~controllable_hgrant5 & ~n22531;
  assign n22533 = ~n15090 & ~n22532;
  assign n22534 = controllable_hmaster2 & ~n22533;
  assign n22535 = ~n13702 & ~n22534;
  assign n22536 = ~controllable_hmaster1 & ~n22535;
  assign n22537 = ~n15208 & ~n22536;
  assign n22538 = ~i_hbusreq6 & ~n22537;
  assign n22539 = ~n22520 & ~n22538;
  assign n22540 = ~controllable_hgrant6 & ~n22539;
  assign n22541 = ~n15253 & ~n22540;
  assign n22542 = ~controllable_hmaster0 & ~n22541;
  assign n22543 = ~n13778 & ~n22542;
  assign n22544 = ~i_hbusreq8 & ~n22543;
  assign n22545 = ~n22519 & ~n22544;
  assign n22546 = ~controllable_hmaster3 & ~n22545;
  assign n22547 = ~n13714 & ~n22546;
  assign n22548 = ~i_hbusreq7 & ~n22547;
  assign n22549 = ~n22518 & ~n22548;
  assign n22550 = n7924 & ~n22549;
  assign n22551 = ~n22500 & ~n22550;
  assign n22552 = n8214 & ~n22551;
  assign n22553 = ~n22472 & ~n22552;
  assign n22554 = ~n8202 & ~n22553;
  assign n22555 = ~n10105 & ~n18123;
  assign n22556 = controllable_hmaster1 & ~n22555;
  assign n22557 = ~n9096 & ~n22556;
  assign n22558 = ~controllable_hgrant6 & ~n22557;
  assign n22559 = ~n15293 & ~n22558;
  assign n22560 = controllable_hmaster0 & ~n22559;
  assign n22561 = ~n9099 & ~n22560;
  assign n22562 = ~controllable_hmaster3 & ~n22561;
  assign n22563 = ~n13651 & ~n22562;
  assign n22564 = i_hbusreq7 & ~n22563;
  assign n22565 = i_hbusreq8 & ~n22561;
  assign n22566 = i_hbusreq6 & ~n22557;
  assign n22567 = ~n10116 & ~n21699;
  assign n22568 = controllable_hmaster1 & ~n22567;
  assign n22569 = ~n9122 & ~n22568;
  assign n22570 = ~i_hbusreq6 & ~n22569;
  assign n22571 = ~n22566 & ~n22570;
  assign n22572 = ~controllable_hgrant6 & ~n22571;
  assign n22573 = ~n15306 & ~n22572;
  assign n22574 = controllable_hmaster0 & ~n22573;
  assign n22575 = ~n9127 & ~n22574;
  assign n22576 = ~i_hbusreq8 & ~n22575;
  assign n22577 = ~n22565 & ~n22576;
  assign n22578 = ~controllable_hmaster3 & ~n22577;
  assign n22579 = ~n13662 & ~n22578;
  assign n22580 = ~i_hbusreq7 & ~n22579;
  assign n22581 = ~n22564 & ~n22580;
  assign n22582 = ~n7924 & ~n22581;
  assign n22583 = i_hlock3 & ~n17769;
  assign n22584 = ~i_hlock3 & ~n17787;
  assign n22585 = ~n22583 & ~n22584;
  assign n22586 = ~controllable_hgrant3 & ~n22585;
  assign n22587 = ~n13852 & ~n22586;
  assign n22588 = ~controllable_hgrant4 & ~n22587;
  assign n22589 = ~n13851 & ~n22588;
  assign n22590 = ~controllable_hgrant5 & ~n22589;
  assign n22591 = ~n13850 & ~n22590;
  assign n22592 = ~controllable_hmaster2 & ~n22591;
  assign n22593 = ~n15294 & ~n22592;
  assign n22594 = controllable_hmaster1 & ~n22593;
  assign n22595 = ~n13677 & ~n22594;
  assign n22596 = ~controllable_hgrant6 & ~n22595;
  assign n22597 = ~n15293 & ~n22596;
  assign n22598 = controllable_hmaster0 & ~n22597;
  assign n22599 = ~n13682 & ~n22598;
  assign n22600 = ~controllable_hmaster3 & ~n22599;
  assign n22601 = ~n13672 & ~n22600;
  assign n22602 = i_hbusreq7 & ~n22601;
  assign n22603 = i_hbusreq8 & ~n22599;
  assign n22604 = i_hbusreq6 & ~n22595;
  assign n22605 = i_hbusreq5 & ~n22589;
  assign n22606 = i_hbusreq4 & ~n22587;
  assign n22607 = i_hbusreq9 & ~n22587;
  assign n22608 = i_hbusreq3 & ~n22585;
  assign n22609 = i_hlock3 & ~n17836;
  assign n22610 = ~i_hlock3 & ~n17872;
  assign n22611 = ~n22609 & ~n22610;
  assign n22612 = ~i_hbusreq3 & ~n22611;
  assign n22613 = ~n22608 & ~n22612;
  assign n22614 = ~controllable_hgrant3 & ~n22613;
  assign n22615 = ~n14999 & ~n22614;
  assign n22616 = ~i_hbusreq9 & ~n22615;
  assign n22617 = ~n22607 & ~n22616;
  assign n22618 = ~i_hbusreq4 & ~n22617;
  assign n22619 = ~n22606 & ~n22618;
  assign n22620 = ~controllable_hgrant4 & ~n22619;
  assign n22621 = ~n14998 & ~n22620;
  assign n22622 = ~i_hbusreq5 & ~n22621;
  assign n22623 = ~n22605 & ~n22622;
  assign n22624 = ~controllable_hgrant5 & ~n22623;
  assign n22625 = ~n14997 & ~n22624;
  assign n22626 = ~controllable_hmaster2 & ~n22625;
  assign n22627 = ~n15308 & ~n22626;
  assign n22628 = controllable_hmaster1 & ~n22627;
  assign n22629 = ~n13721 & ~n22628;
  assign n22630 = ~i_hbusreq6 & ~n22629;
  assign n22631 = ~n22604 & ~n22630;
  assign n22632 = ~controllable_hgrant6 & ~n22631;
  assign n22633 = ~n15306 & ~n22632;
  assign n22634 = controllable_hmaster0 & ~n22633;
  assign n22635 = ~n13728 & ~n22634;
  assign n22636 = ~i_hbusreq8 & ~n22635;
  assign n22637 = ~n22603 & ~n22636;
  assign n22638 = ~controllable_hmaster3 & ~n22637;
  assign n22639 = ~n13714 & ~n22638;
  assign n22640 = ~i_hbusreq7 & ~n22639;
  assign n22641 = ~n22602 & ~n22640;
  assign n22642 = n7924 & ~n22641;
  assign n22643 = ~n22582 & ~n22642;
  assign n22644 = ~n8214 & ~n22643;
  assign n22645 = ~n10105 & ~n18159;
  assign n22646 = controllable_hmaster1 & ~n22645;
  assign n22647 = ~n9096 & ~n22646;
  assign n22648 = ~controllable_hgrant6 & ~n22647;
  assign n22649 = ~n15351 & ~n22648;
  assign n22650 = ~controllable_hmaster0 & ~n22649;
  assign n22651 = ~n9152 & ~n22650;
  assign n22652 = ~controllable_hmaster3 & ~n22651;
  assign n22653 = ~n13651 & ~n22652;
  assign n22654 = i_hbusreq7 & ~n22653;
  assign n22655 = i_hbusreq8 & ~n22651;
  assign n22656 = i_hbusreq6 & ~n22647;
  assign n22657 = ~n10116 & ~n21759;
  assign n22658 = controllable_hmaster1 & ~n22657;
  assign n22659 = ~n9122 & ~n22658;
  assign n22660 = ~i_hbusreq6 & ~n22659;
  assign n22661 = ~n22656 & ~n22660;
  assign n22662 = ~controllable_hgrant6 & ~n22661;
  assign n22663 = ~n15363 & ~n22662;
  assign n22664 = ~controllable_hmaster0 & ~n22663;
  assign n22665 = ~n9162 & ~n22664;
  assign n22666 = ~i_hbusreq8 & ~n22665;
  assign n22667 = ~n22655 & ~n22666;
  assign n22668 = ~controllable_hmaster3 & ~n22667;
  assign n22669 = ~n13662 & ~n22668;
  assign n22670 = ~i_hbusreq7 & ~n22669;
  assign n22671 = ~n22654 & ~n22670;
  assign n22672 = ~n7924 & ~n22671;
  assign n22673 = ~n9213 & ~n17766;
  assign n22674 = ~controllable_hgrant1 & ~n22673;
  assign n22675 = ~n13898 & ~n22674;
  assign n22676 = ~controllable_hgrant3 & ~n22675;
  assign n22677 = ~n13897 & ~n22676;
  assign n22678 = ~controllable_hgrant4 & ~n22677;
  assign n22679 = ~n13896 & ~n22678;
  assign n22680 = ~controllable_hgrant5 & ~n22679;
  assign n22681 = ~n13895 & ~n22680;
  assign n22682 = ~controllable_hmaster2 & ~n22681;
  assign n22683 = ~n15294 & ~n22682;
  assign n22684 = controllable_hmaster1 & ~n22683;
  assign n22685 = ~n13677 & ~n22684;
  assign n22686 = ~controllable_hgrant6 & ~n22685;
  assign n22687 = ~n15351 & ~n22686;
  assign n22688 = ~controllable_hmaster0 & ~n22687;
  assign n22689 = ~n13765 & ~n22688;
  assign n22690 = ~controllable_hmaster3 & ~n22689;
  assign n22691 = ~n13672 & ~n22690;
  assign n22692 = i_hbusreq7 & ~n22691;
  assign n22693 = i_hbusreq8 & ~n22689;
  assign n22694 = i_hbusreq6 & ~n22685;
  assign n22695 = i_hbusreq5 & ~n22679;
  assign n22696 = i_hbusreq4 & ~n22677;
  assign n22697 = i_hbusreq9 & ~n22677;
  assign n22698 = i_hbusreq3 & ~n22675;
  assign n22699 = i_hbusreq1 & ~n22673;
  assign n22700 = ~n9379 & ~n17831;
  assign n22701 = ~i_hbusreq1 & ~n22700;
  assign n22702 = ~n22699 & ~n22701;
  assign n22703 = ~controllable_hgrant1 & ~n22702;
  assign n22704 = ~n15067 & ~n22703;
  assign n22705 = ~i_hbusreq3 & ~n22704;
  assign n22706 = ~n22698 & ~n22705;
  assign n22707 = ~controllable_hgrant3 & ~n22706;
  assign n22708 = ~n15066 & ~n22707;
  assign n22709 = ~i_hbusreq9 & ~n22708;
  assign n22710 = ~n22697 & ~n22709;
  assign n22711 = ~i_hbusreq4 & ~n22710;
  assign n22712 = ~n22696 & ~n22711;
  assign n22713 = ~controllable_hgrant4 & ~n22712;
  assign n22714 = ~n15065 & ~n22713;
  assign n22715 = ~i_hbusreq5 & ~n22714;
  assign n22716 = ~n22695 & ~n22715;
  assign n22717 = ~controllable_hgrant5 & ~n22716;
  assign n22718 = ~n15064 & ~n22717;
  assign n22719 = ~controllable_hmaster2 & ~n22718;
  assign n22720 = ~n15308 & ~n22719;
  assign n22721 = controllable_hmaster1 & ~n22720;
  assign n22722 = ~n13721 & ~n22721;
  assign n22723 = ~i_hbusreq6 & ~n22722;
  assign n22724 = ~n22694 & ~n22723;
  assign n22725 = ~controllable_hgrant6 & ~n22724;
  assign n22726 = ~n15363 & ~n22725;
  assign n22727 = ~controllable_hmaster0 & ~n22726;
  assign n22728 = ~n13778 & ~n22727;
  assign n22729 = ~i_hbusreq8 & ~n22728;
  assign n22730 = ~n22693 & ~n22729;
  assign n22731 = ~controllable_hmaster3 & ~n22730;
  assign n22732 = ~n13714 & ~n22731;
  assign n22733 = ~i_hbusreq7 & ~n22732;
  assign n22734 = ~n22692 & ~n22733;
  assign n22735 = n7924 & ~n22734;
  assign n22736 = ~n22672 & ~n22735;
  assign n22737 = n8214 & ~n22736;
  assign n22738 = ~n22644 & ~n22737;
  assign n22739 = n8202 & ~n22738;
  assign n22740 = ~n22554 & ~n22739;
  assign n22741 = n7920 & ~n22740;
  assign n22742 = ~n10014 & ~n22741;
  assign n22743 = n7728 & ~n22742;
  assign n22744 = ~n18131 & ~n19273;
  assign n22745 = ~controllable_hmaster1 & ~n22744;
  assign n22746 = ~n19251 & ~n22745;
  assign n22747 = ~controllable_hgrant6 & ~n22746;
  assign n22748 = ~n13849 & ~n22747;
  assign n22749 = controllable_hmaster0 & ~n22748;
  assign n22750 = ~n19324 & ~n22749;
  assign n22751 = ~controllable_hmaster3 & ~n22750;
  assign n22752 = ~n20287 & ~n22751;
  assign n22753 = i_hlock7 & ~n22752;
  assign n22754 = ~n19330 & ~n22745;
  assign n22755 = ~controllable_hgrant6 & ~n22754;
  assign n22756 = ~n13951 & ~n22755;
  assign n22757 = controllable_hmaster0 & ~n22756;
  assign n22758 = ~n19324 & ~n22757;
  assign n22759 = ~controllable_hmaster3 & ~n22758;
  assign n22760 = ~n20287 & ~n22759;
  assign n22761 = ~i_hlock7 & ~n22760;
  assign n22762 = ~n22753 & ~n22761;
  assign n22763 = i_hbusreq7 & ~n22762;
  assign n22764 = i_hbusreq8 & ~n22750;
  assign n22765 = i_hbusreq6 & ~n22746;
  assign n22766 = ~n19548 & ~n21709;
  assign n22767 = ~controllable_hmaster1 & ~n22766;
  assign n22768 = ~n19499 & ~n22767;
  assign n22769 = ~i_hbusreq6 & ~n22768;
  assign n22770 = ~n22765 & ~n22769;
  assign n22771 = ~controllable_hgrant6 & ~n22770;
  assign n22772 = ~n15417 & ~n22771;
  assign n22773 = controllable_hmaster0 & ~n22772;
  assign n22774 = ~n19644 & ~n22773;
  assign n22775 = ~i_hbusreq8 & ~n22774;
  assign n22776 = ~n22764 & ~n22775;
  assign n22777 = ~controllable_hmaster3 & ~n22776;
  assign n22778 = ~n20338 & ~n22777;
  assign n22779 = i_hlock7 & ~n22778;
  assign n22780 = i_hbusreq8 & ~n22758;
  assign n22781 = i_hbusreq6 & ~n22754;
  assign n22782 = ~n19654 & ~n22767;
  assign n22783 = ~i_hbusreq6 & ~n22782;
  assign n22784 = ~n22781 & ~n22783;
  assign n22785 = ~controllable_hgrant6 & ~n22784;
  assign n22786 = ~n15440 & ~n22785;
  assign n22787 = controllable_hmaster0 & ~n22786;
  assign n22788 = ~n19644 & ~n22787;
  assign n22789 = ~i_hbusreq8 & ~n22788;
  assign n22790 = ~n22780 & ~n22789;
  assign n22791 = ~controllable_hmaster3 & ~n22790;
  assign n22792 = ~n20338 & ~n22791;
  assign n22793 = ~i_hlock7 & ~n22792;
  assign n22794 = ~n22779 & ~n22793;
  assign n22795 = ~i_hbusreq7 & ~n22794;
  assign n22796 = ~n22763 & ~n22795;
  assign n22797 = ~n7924 & ~n22796;
  assign n22798 = i_hlock5 & ~n19720;
  assign n22799 = ~i_hlock5 & ~n19738;
  assign n22800 = ~n22798 & ~n22799;
  assign n22801 = ~controllable_hgrant5 & ~n22800;
  assign n22802 = ~n13865 & ~n22801;
  assign n22803 = controllable_hmaster2 & ~n22802;
  assign n22804 = ~n19798 & ~n22803;
  assign n22805 = ~controllable_hmaster1 & ~n22804;
  assign n22806 = ~n19776 & ~n22805;
  assign n22807 = ~controllable_hgrant6 & ~n22806;
  assign n22808 = ~n13849 & ~n22807;
  assign n22809 = controllable_hmaster0 & ~n22808;
  assign n22810 = ~n19849 & ~n22809;
  assign n22811 = ~controllable_hmaster3 & ~n22810;
  assign n22812 = ~n20394 & ~n22811;
  assign n22813 = i_hlock7 & ~n22812;
  assign n22814 = ~n19855 & ~n22805;
  assign n22815 = ~controllable_hgrant6 & ~n22814;
  assign n22816 = ~n13951 & ~n22815;
  assign n22817 = controllable_hmaster0 & ~n22816;
  assign n22818 = ~n19849 & ~n22817;
  assign n22819 = ~controllable_hmaster3 & ~n22818;
  assign n22820 = ~n20394 & ~n22819;
  assign n22821 = ~i_hlock7 & ~n22820;
  assign n22822 = ~n22813 & ~n22821;
  assign n22823 = i_hbusreq7 & ~n22822;
  assign n22824 = i_hbusreq8 & ~n22810;
  assign n22825 = i_hbusreq6 & ~n22806;
  assign n22826 = i_hbusreq5 & ~n22800;
  assign n22827 = i_hlock5 & ~n19980;
  assign n22828 = ~i_hlock5 & ~n20016;
  assign n22829 = ~n22827 & ~n22828;
  assign n22830 = ~i_hbusreq5 & ~n22829;
  assign n22831 = ~n22826 & ~n22830;
  assign n22832 = ~controllable_hgrant5 & ~n22831;
  assign n22833 = ~n15020 & ~n22832;
  assign n22834 = controllable_hmaster2 & ~n22833;
  assign n22835 = ~n20141 & ~n22834;
  assign n22836 = ~controllable_hmaster1 & ~n22835;
  assign n22837 = ~n20092 & ~n22836;
  assign n22838 = ~i_hbusreq6 & ~n22837;
  assign n22839 = ~n22825 & ~n22838;
  assign n22840 = ~controllable_hgrant6 & ~n22839;
  assign n22841 = ~n15417 & ~n22840;
  assign n22842 = controllable_hmaster0 & ~n22841;
  assign n22843 = ~n20237 & ~n22842;
  assign n22844 = ~i_hbusreq8 & ~n22843;
  assign n22845 = ~n22824 & ~n22844;
  assign n22846 = ~controllable_hmaster3 & ~n22845;
  assign n22847 = ~n20447 & ~n22846;
  assign n22848 = i_hlock7 & ~n22847;
  assign n22849 = i_hbusreq8 & ~n22818;
  assign n22850 = i_hbusreq6 & ~n22814;
  assign n22851 = ~n20247 & ~n22836;
  assign n22852 = ~i_hbusreq6 & ~n22851;
  assign n22853 = ~n22850 & ~n22852;
  assign n22854 = ~controllable_hgrant6 & ~n22853;
  assign n22855 = ~n15440 & ~n22854;
  assign n22856 = controllable_hmaster0 & ~n22855;
  assign n22857 = ~n20237 & ~n22856;
  assign n22858 = ~i_hbusreq8 & ~n22857;
  assign n22859 = ~n22849 & ~n22858;
  assign n22860 = ~controllable_hmaster3 & ~n22859;
  assign n22861 = ~n20447 & ~n22860;
  assign n22862 = ~i_hlock7 & ~n22861;
  assign n22863 = ~n22848 & ~n22862;
  assign n22864 = ~i_hbusreq7 & ~n22863;
  assign n22865 = ~n22823 & ~n22864;
  assign n22866 = n7924 & ~n22865;
  assign n22867 = ~n22797 & ~n22866;
  assign n22868 = ~n8214 & ~n22867;
  assign n22869 = ~n18169 & ~n19309;
  assign n22870 = ~controllable_hmaster1 & ~n22869;
  assign n22871 = ~n19291 & ~n22870;
  assign n22872 = i_hlock6 & ~n22871;
  assign n22873 = ~n19318 & ~n22870;
  assign n22874 = ~i_hlock6 & ~n22873;
  assign n22875 = ~n22872 & ~n22874;
  assign n22876 = ~controllable_hgrant6 & ~n22875;
  assign n22877 = ~n13894 & ~n22876;
  assign n22878 = ~controllable_hmaster0 & ~n22877;
  assign n22879 = ~n19279 & ~n22878;
  assign n22880 = ~controllable_hmaster3 & ~n22879;
  assign n22881 = ~n20287 & ~n22880;
  assign n22882 = i_hlock7 & ~n22881;
  assign n22883 = ~n19334 & ~n22878;
  assign n22884 = ~controllable_hmaster3 & ~n22883;
  assign n22885 = ~n20287 & ~n22884;
  assign n22886 = ~i_hlock7 & ~n22885;
  assign n22887 = ~n22882 & ~n22886;
  assign n22888 = i_hbusreq7 & ~n22887;
  assign n22889 = i_hbusreq8 & ~n22879;
  assign n22890 = i_hbusreq6 & ~n22875;
  assign n22891 = ~n19624 & ~n21773;
  assign n22892 = ~controllable_hmaster1 & ~n22891;
  assign n22893 = ~n19584 & ~n22892;
  assign n22894 = i_hlock6 & ~n22893;
  assign n22895 = ~n19636 & ~n22892;
  assign n22896 = ~i_hlock6 & ~n22895;
  assign n22897 = ~n22894 & ~n22896;
  assign n22898 = ~i_hbusreq6 & ~n22897;
  assign n22899 = ~n22890 & ~n22898;
  assign n22900 = ~controllable_hgrant6 & ~n22899;
  assign n22901 = ~n15467 & ~n22900;
  assign n22902 = ~controllable_hmaster0 & ~n22901;
  assign n22903 = ~n19556 & ~n22902;
  assign n22904 = ~i_hbusreq8 & ~n22903;
  assign n22905 = ~n22889 & ~n22904;
  assign n22906 = ~controllable_hmaster3 & ~n22905;
  assign n22907 = ~n20338 & ~n22906;
  assign n22908 = i_hlock7 & ~n22907;
  assign n22909 = i_hbusreq8 & ~n22883;
  assign n22910 = ~n19660 & ~n22902;
  assign n22911 = ~i_hbusreq8 & ~n22910;
  assign n22912 = ~n22909 & ~n22911;
  assign n22913 = ~controllable_hmaster3 & ~n22912;
  assign n22914 = ~n20338 & ~n22913;
  assign n22915 = ~i_hlock7 & ~n22914;
  assign n22916 = ~n22908 & ~n22915;
  assign n22917 = ~i_hbusreq7 & ~n22916;
  assign n22918 = ~n22888 & ~n22917;
  assign n22919 = ~n7924 & ~n22918;
  assign n22920 = i_hlock4 & ~n19718;
  assign n22921 = ~i_hlock4 & ~n19736;
  assign n22922 = ~n22920 & ~n22921;
  assign n22923 = ~controllable_hgrant4 & ~n22922;
  assign n22924 = ~n13912 & ~n22923;
  assign n22925 = ~controllable_hgrant5 & ~n22924;
  assign n22926 = ~n13911 & ~n22925;
  assign n22927 = controllable_hmaster2 & ~n22926;
  assign n22928 = ~n19834 & ~n22927;
  assign n22929 = ~controllable_hmaster1 & ~n22928;
  assign n22930 = ~n19816 & ~n22929;
  assign n22931 = i_hlock6 & ~n22930;
  assign n22932 = ~n19843 & ~n22929;
  assign n22933 = ~i_hlock6 & ~n22932;
  assign n22934 = ~n22931 & ~n22933;
  assign n22935 = ~controllable_hgrant6 & ~n22934;
  assign n22936 = ~n13894 & ~n22935;
  assign n22937 = ~controllable_hmaster0 & ~n22936;
  assign n22938 = ~n19804 & ~n22937;
  assign n22939 = ~controllable_hmaster3 & ~n22938;
  assign n22940 = ~n20394 & ~n22939;
  assign n22941 = i_hlock7 & ~n22940;
  assign n22942 = ~n19859 & ~n22937;
  assign n22943 = ~controllable_hmaster3 & ~n22942;
  assign n22944 = ~n20394 & ~n22943;
  assign n22945 = ~i_hlock7 & ~n22944;
  assign n22946 = ~n22941 & ~n22945;
  assign n22947 = i_hbusreq7 & ~n22946;
  assign n22948 = i_hbusreq8 & ~n22938;
  assign n22949 = i_hbusreq6 & ~n22934;
  assign n22950 = i_hbusreq5 & ~n22924;
  assign n22951 = i_hbusreq4 & ~n22922;
  assign n22952 = i_hlock4 & ~n19976;
  assign n22953 = ~i_hlock4 & ~n20012;
  assign n22954 = ~n22952 & ~n22953;
  assign n22955 = ~i_hbusreq4 & ~n22954;
  assign n22956 = ~n22951 & ~n22955;
  assign n22957 = ~controllable_hgrant4 & ~n22956;
  assign n22958 = ~n15091 & ~n22957;
  assign n22959 = ~i_hbusreq5 & ~n22958;
  assign n22960 = ~n22950 & ~n22959;
  assign n22961 = ~controllable_hgrant5 & ~n22960;
  assign n22962 = ~n15090 & ~n22961;
  assign n22963 = controllable_hmaster2 & ~n22962;
  assign n22964 = ~n20217 & ~n22963;
  assign n22965 = ~controllable_hmaster1 & ~n22964;
  assign n22966 = ~n20177 & ~n22965;
  assign n22967 = i_hlock6 & ~n22966;
  assign n22968 = ~n20229 & ~n22965;
  assign n22969 = ~i_hlock6 & ~n22968;
  assign n22970 = ~n22967 & ~n22969;
  assign n22971 = ~i_hbusreq6 & ~n22970;
  assign n22972 = ~n22949 & ~n22971;
  assign n22973 = ~controllable_hgrant6 & ~n22972;
  assign n22974 = ~n15467 & ~n22973;
  assign n22975 = ~controllable_hmaster0 & ~n22974;
  assign n22976 = ~n20149 & ~n22975;
  assign n22977 = ~i_hbusreq8 & ~n22976;
  assign n22978 = ~n22948 & ~n22977;
  assign n22979 = ~controllable_hmaster3 & ~n22978;
  assign n22980 = ~n20447 & ~n22979;
  assign n22981 = i_hlock7 & ~n22980;
  assign n22982 = i_hbusreq8 & ~n22942;
  assign n22983 = ~n20253 & ~n22975;
  assign n22984 = ~i_hbusreq8 & ~n22983;
  assign n22985 = ~n22982 & ~n22984;
  assign n22986 = ~controllable_hmaster3 & ~n22985;
  assign n22987 = ~n20447 & ~n22986;
  assign n22988 = ~i_hlock7 & ~n22987;
  assign n22989 = ~n22981 & ~n22988;
  assign n22990 = ~i_hbusreq7 & ~n22989;
  assign n22991 = ~n22947 & ~n22990;
  assign n22992 = n7924 & ~n22991;
  assign n22993 = ~n22919 & ~n22992;
  assign n22994 = n8214 & ~n22993;
  assign n22995 = ~n22868 & ~n22994;
  assign n22996 = ~n8202 & ~n22995;
  assign n22997 = ~n18123 & ~n19236;
  assign n22998 = controllable_hmaster1 & ~n22997;
  assign n22999 = ~n19275 & ~n22998;
  assign n23000 = ~controllable_hgrant6 & ~n22999;
  assign n23001 = ~n13849 & ~n23000;
  assign n23002 = controllable_hmaster0 & ~n23001;
  assign n23003 = ~n19324 & ~n23002;
  assign n23004 = ~controllable_hmaster3 & ~n23003;
  assign n23005 = ~n20287 & ~n23004;
  assign n23006 = i_hlock7 & ~n23005;
  assign n23007 = ~n18123 & ~n19316;
  assign n23008 = controllable_hmaster1 & ~n23007;
  assign n23009 = ~n19275 & ~n23008;
  assign n23010 = ~controllable_hgrant6 & ~n23009;
  assign n23011 = ~n13951 & ~n23010;
  assign n23012 = controllable_hmaster0 & ~n23011;
  assign n23013 = ~n19324 & ~n23012;
  assign n23014 = ~controllable_hmaster3 & ~n23013;
  assign n23015 = ~n20287 & ~n23014;
  assign n23016 = ~i_hlock7 & ~n23015;
  assign n23017 = ~n23006 & ~n23016;
  assign n23018 = i_hbusreq7 & ~n23017;
  assign n23019 = i_hbusreq8 & ~n23003;
  assign n23020 = i_hbusreq6 & ~n22999;
  assign n23021 = ~n19469 & ~n21699;
  assign n23022 = controllable_hmaster1 & ~n23021;
  assign n23023 = ~n19550 & ~n23022;
  assign n23024 = ~i_hbusreq6 & ~n23023;
  assign n23025 = ~n23020 & ~n23024;
  assign n23026 = ~controllable_hgrant6 & ~n23025;
  assign n23027 = ~n15520 & ~n23026;
  assign n23028 = controllable_hmaster0 & ~n23027;
  assign n23029 = ~n19644 & ~n23028;
  assign n23030 = ~i_hbusreq8 & ~n23029;
  assign n23031 = ~n23019 & ~n23030;
  assign n23032 = ~controllable_hmaster3 & ~n23031;
  assign n23033 = ~n20338 & ~n23032;
  assign n23034 = i_hlock7 & ~n23033;
  assign n23035 = i_hbusreq8 & ~n23013;
  assign n23036 = i_hbusreq6 & ~n23009;
  assign n23037 = ~n19634 & ~n21699;
  assign n23038 = controllable_hmaster1 & ~n23037;
  assign n23039 = ~n19550 & ~n23038;
  assign n23040 = ~i_hbusreq6 & ~n23039;
  assign n23041 = ~n23036 & ~n23040;
  assign n23042 = ~controllable_hgrant6 & ~n23041;
  assign n23043 = ~n15553 & ~n23042;
  assign n23044 = controllable_hmaster0 & ~n23043;
  assign n23045 = ~n19644 & ~n23044;
  assign n23046 = ~i_hbusreq8 & ~n23045;
  assign n23047 = ~n23035 & ~n23046;
  assign n23048 = ~controllable_hmaster3 & ~n23047;
  assign n23049 = ~n20338 & ~n23048;
  assign n23050 = ~i_hlock7 & ~n23049;
  assign n23051 = ~n23034 & ~n23050;
  assign n23052 = ~i_hbusreq7 & ~n23051;
  assign n23053 = ~n23018 & ~n23052;
  assign n23054 = ~n7924 & ~n23053;
  assign n23055 = i_hlock3 & ~n19716;
  assign n23056 = ~i_hlock3 & ~n19734;
  assign n23057 = ~n23055 & ~n23056;
  assign n23058 = ~controllable_hgrant3 & ~n23057;
  assign n23059 = ~n13852 & ~n23058;
  assign n23060 = ~controllable_hgrant4 & ~n23059;
  assign n23061 = ~n13851 & ~n23060;
  assign n23062 = ~controllable_hgrant5 & ~n23061;
  assign n23063 = ~n13850 & ~n23062;
  assign n23064 = ~controllable_hmaster2 & ~n23063;
  assign n23065 = ~n19761 & ~n23064;
  assign n23066 = controllable_hmaster1 & ~n23065;
  assign n23067 = ~n19800 & ~n23066;
  assign n23068 = ~controllable_hgrant6 & ~n23067;
  assign n23069 = ~n13849 & ~n23068;
  assign n23070 = controllable_hmaster0 & ~n23069;
  assign n23071 = ~n19849 & ~n23070;
  assign n23072 = ~controllable_hmaster3 & ~n23071;
  assign n23073 = ~n20394 & ~n23072;
  assign n23074 = i_hlock7 & ~n23073;
  assign n23075 = ~n19841 & ~n23064;
  assign n23076 = controllable_hmaster1 & ~n23075;
  assign n23077 = ~n19800 & ~n23076;
  assign n23078 = ~controllable_hgrant6 & ~n23077;
  assign n23079 = ~n13951 & ~n23078;
  assign n23080 = controllable_hmaster0 & ~n23079;
  assign n23081 = ~n19849 & ~n23080;
  assign n23082 = ~controllable_hmaster3 & ~n23081;
  assign n23083 = ~n20394 & ~n23082;
  assign n23084 = ~i_hlock7 & ~n23083;
  assign n23085 = ~n23074 & ~n23084;
  assign n23086 = i_hbusreq7 & ~n23085;
  assign n23087 = i_hbusreq8 & ~n23071;
  assign n23088 = i_hbusreq6 & ~n23067;
  assign n23089 = i_hbusreq5 & ~n23061;
  assign n23090 = i_hbusreq4 & ~n23059;
  assign n23091 = i_hbusreq9 & ~n23059;
  assign n23092 = i_hbusreq3 & ~n23057;
  assign n23093 = i_hlock3 & ~n19970;
  assign n23094 = ~i_hlock3 & ~n20006;
  assign n23095 = ~n23093 & ~n23094;
  assign n23096 = ~i_hbusreq3 & ~n23095;
  assign n23097 = ~n23092 & ~n23096;
  assign n23098 = ~controllable_hgrant3 & ~n23097;
  assign n23099 = ~n14999 & ~n23098;
  assign n23100 = ~i_hbusreq9 & ~n23099;
  assign n23101 = ~n23091 & ~n23100;
  assign n23102 = ~i_hbusreq4 & ~n23101;
  assign n23103 = ~n23090 & ~n23102;
  assign n23104 = ~controllable_hgrant4 & ~n23103;
  assign n23105 = ~n14998 & ~n23104;
  assign n23106 = ~i_hbusreq5 & ~n23105;
  assign n23107 = ~n23089 & ~n23106;
  assign n23108 = ~controllable_hgrant5 & ~n23107;
  assign n23109 = ~n14997 & ~n23108;
  assign n23110 = ~controllable_hmaster2 & ~n23109;
  assign n23111 = ~n20062 & ~n23110;
  assign n23112 = controllable_hmaster1 & ~n23111;
  assign n23113 = ~n20143 & ~n23112;
  assign n23114 = ~i_hbusreq6 & ~n23113;
  assign n23115 = ~n23088 & ~n23114;
  assign n23116 = ~controllable_hgrant6 & ~n23115;
  assign n23117 = ~n15520 & ~n23116;
  assign n23118 = controllable_hmaster0 & ~n23117;
  assign n23119 = ~n20237 & ~n23118;
  assign n23120 = ~i_hbusreq8 & ~n23119;
  assign n23121 = ~n23087 & ~n23120;
  assign n23122 = ~controllable_hmaster3 & ~n23121;
  assign n23123 = ~n20447 & ~n23122;
  assign n23124 = i_hlock7 & ~n23123;
  assign n23125 = i_hbusreq8 & ~n23081;
  assign n23126 = i_hbusreq6 & ~n23077;
  assign n23127 = ~n20227 & ~n23110;
  assign n23128 = controllable_hmaster1 & ~n23127;
  assign n23129 = ~n20143 & ~n23128;
  assign n23130 = ~i_hbusreq6 & ~n23129;
  assign n23131 = ~n23126 & ~n23130;
  assign n23132 = ~controllable_hgrant6 & ~n23131;
  assign n23133 = ~n15553 & ~n23132;
  assign n23134 = controllable_hmaster0 & ~n23133;
  assign n23135 = ~n20237 & ~n23134;
  assign n23136 = ~i_hbusreq8 & ~n23135;
  assign n23137 = ~n23125 & ~n23136;
  assign n23138 = ~controllable_hmaster3 & ~n23137;
  assign n23139 = ~n20447 & ~n23138;
  assign n23140 = ~i_hlock7 & ~n23139;
  assign n23141 = ~n23124 & ~n23140;
  assign n23142 = ~i_hbusreq7 & ~n23141;
  assign n23143 = ~n23086 & ~n23142;
  assign n23144 = n7924 & ~n23143;
  assign n23145 = ~n23054 & ~n23144;
  assign n23146 = ~n8214 & ~n23145;
  assign n23147 = ~n18159 & ~n19236;
  assign n23148 = controllable_hmaster1 & ~n23147;
  assign n23149 = ~n19311 & ~n23148;
  assign n23150 = i_hlock6 & ~n23149;
  assign n23151 = ~n18159 & ~n19316;
  assign n23152 = controllable_hmaster1 & ~n23151;
  assign n23153 = ~n19311 & ~n23152;
  assign n23154 = ~i_hlock6 & ~n23153;
  assign n23155 = ~n23150 & ~n23154;
  assign n23156 = ~controllable_hgrant6 & ~n23155;
  assign n23157 = ~n13894 & ~n23156;
  assign n23158 = ~controllable_hmaster0 & ~n23157;
  assign n23159 = ~n19279 & ~n23158;
  assign n23160 = ~controllable_hmaster3 & ~n23159;
  assign n23161 = ~n20287 & ~n23160;
  assign n23162 = i_hlock7 & ~n23161;
  assign n23163 = ~n19334 & ~n23158;
  assign n23164 = ~controllable_hmaster3 & ~n23163;
  assign n23165 = ~n20287 & ~n23164;
  assign n23166 = ~i_hlock7 & ~n23165;
  assign n23167 = ~n23162 & ~n23166;
  assign n23168 = i_hbusreq7 & ~n23167;
  assign n23169 = i_hbusreq8 & ~n23159;
  assign n23170 = i_hbusreq6 & ~n23155;
  assign n23171 = ~n19469 & ~n21759;
  assign n23172 = controllable_hmaster1 & ~n23171;
  assign n23173 = ~n19626 & ~n23172;
  assign n23174 = i_hlock6 & ~n23173;
  assign n23175 = ~n19634 & ~n21759;
  assign n23176 = controllable_hmaster1 & ~n23175;
  assign n23177 = ~n19626 & ~n23176;
  assign n23178 = ~i_hlock6 & ~n23177;
  assign n23179 = ~n23174 & ~n23178;
  assign n23180 = ~i_hbusreq6 & ~n23179;
  assign n23181 = ~n23170 & ~n23180;
  assign n23182 = ~controllable_hgrant6 & ~n23181;
  assign n23183 = ~n15582 & ~n23182;
  assign n23184 = ~controllable_hmaster0 & ~n23183;
  assign n23185 = ~n19556 & ~n23184;
  assign n23186 = ~i_hbusreq8 & ~n23185;
  assign n23187 = ~n23169 & ~n23186;
  assign n23188 = ~controllable_hmaster3 & ~n23187;
  assign n23189 = ~n20338 & ~n23188;
  assign n23190 = i_hlock7 & ~n23189;
  assign n23191 = i_hbusreq8 & ~n23163;
  assign n23192 = ~n19660 & ~n23184;
  assign n23193 = ~i_hbusreq8 & ~n23192;
  assign n23194 = ~n23191 & ~n23193;
  assign n23195 = ~controllable_hmaster3 & ~n23194;
  assign n23196 = ~n20338 & ~n23195;
  assign n23197 = ~i_hlock7 & ~n23196;
  assign n23198 = ~n23190 & ~n23197;
  assign n23199 = ~i_hbusreq7 & ~n23198;
  assign n23200 = ~n23168 & ~n23199;
  assign n23201 = ~n7924 & ~n23200;
  assign n23202 = ~n9213 & ~n19713;
  assign n23203 = ~controllable_hgrant1 & ~n23202;
  assign n23204 = ~n13898 & ~n23203;
  assign n23205 = ~controllable_hgrant3 & ~n23204;
  assign n23206 = ~n13897 & ~n23205;
  assign n23207 = ~controllable_hgrant4 & ~n23206;
  assign n23208 = ~n13896 & ~n23207;
  assign n23209 = ~controllable_hgrant5 & ~n23208;
  assign n23210 = ~n13895 & ~n23209;
  assign n23211 = ~controllable_hmaster2 & ~n23210;
  assign n23212 = ~n19761 & ~n23211;
  assign n23213 = controllable_hmaster1 & ~n23212;
  assign n23214 = ~n19836 & ~n23213;
  assign n23215 = i_hlock6 & ~n23214;
  assign n23216 = ~n19841 & ~n23211;
  assign n23217 = controllable_hmaster1 & ~n23216;
  assign n23218 = ~n19836 & ~n23217;
  assign n23219 = ~i_hlock6 & ~n23218;
  assign n23220 = ~n23215 & ~n23219;
  assign n23221 = ~controllable_hgrant6 & ~n23220;
  assign n23222 = ~n13894 & ~n23221;
  assign n23223 = ~controllable_hmaster0 & ~n23222;
  assign n23224 = ~n19804 & ~n23223;
  assign n23225 = ~controllable_hmaster3 & ~n23224;
  assign n23226 = ~n20394 & ~n23225;
  assign n23227 = i_hlock7 & ~n23226;
  assign n23228 = ~n19859 & ~n23223;
  assign n23229 = ~controllable_hmaster3 & ~n23228;
  assign n23230 = ~n20394 & ~n23229;
  assign n23231 = ~i_hlock7 & ~n23230;
  assign n23232 = ~n23227 & ~n23231;
  assign n23233 = i_hbusreq7 & ~n23232;
  assign n23234 = i_hbusreq8 & ~n23224;
  assign n23235 = i_hbusreq6 & ~n23220;
  assign n23236 = i_hbusreq5 & ~n23208;
  assign n23237 = i_hbusreq4 & ~n23206;
  assign n23238 = i_hbusreq9 & ~n23206;
  assign n23239 = i_hbusreq3 & ~n23204;
  assign n23240 = i_hbusreq1 & ~n23202;
  assign n23241 = ~n9379 & ~n19965;
  assign n23242 = ~i_hbusreq1 & ~n23241;
  assign n23243 = ~n23240 & ~n23242;
  assign n23244 = ~controllable_hgrant1 & ~n23243;
  assign n23245 = ~n15067 & ~n23244;
  assign n23246 = ~i_hbusreq3 & ~n23245;
  assign n23247 = ~n23239 & ~n23246;
  assign n23248 = ~controllable_hgrant3 & ~n23247;
  assign n23249 = ~n15066 & ~n23248;
  assign n23250 = ~i_hbusreq9 & ~n23249;
  assign n23251 = ~n23238 & ~n23250;
  assign n23252 = ~i_hbusreq4 & ~n23251;
  assign n23253 = ~n23237 & ~n23252;
  assign n23254 = ~controllable_hgrant4 & ~n23253;
  assign n23255 = ~n15065 & ~n23254;
  assign n23256 = ~i_hbusreq5 & ~n23255;
  assign n23257 = ~n23236 & ~n23256;
  assign n23258 = ~controllable_hgrant5 & ~n23257;
  assign n23259 = ~n15064 & ~n23258;
  assign n23260 = ~controllable_hmaster2 & ~n23259;
  assign n23261 = ~n20062 & ~n23260;
  assign n23262 = controllable_hmaster1 & ~n23261;
  assign n23263 = ~n20219 & ~n23262;
  assign n23264 = i_hlock6 & ~n23263;
  assign n23265 = ~n20227 & ~n23260;
  assign n23266 = controllable_hmaster1 & ~n23265;
  assign n23267 = ~n20219 & ~n23266;
  assign n23268 = ~i_hlock6 & ~n23267;
  assign n23269 = ~n23264 & ~n23268;
  assign n23270 = ~i_hbusreq6 & ~n23269;
  assign n23271 = ~n23235 & ~n23270;
  assign n23272 = ~controllable_hgrant6 & ~n23271;
  assign n23273 = ~n15582 & ~n23272;
  assign n23274 = ~controllable_hmaster0 & ~n23273;
  assign n23275 = ~n20149 & ~n23274;
  assign n23276 = ~i_hbusreq8 & ~n23275;
  assign n23277 = ~n23234 & ~n23276;
  assign n23278 = ~controllable_hmaster3 & ~n23277;
  assign n23279 = ~n20447 & ~n23278;
  assign n23280 = i_hlock7 & ~n23279;
  assign n23281 = i_hbusreq8 & ~n23228;
  assign n23282 = ~n20253 & ~n23274;
  assign n23283 = ~i_hbusreq8 & ~n23282;
  assign n23284 = ~n23281 & ~n23283;
  assign n23285 = ~controllable_hmaster3 & ~n23284;
  assign n23286 = ~n20447 & ~n23285;
  assign n23287 = ~i_hlock7 & ~n23286;
  assign n23288 = ~n23280 & ~n23287;
  assign n23289 = ~i_hbusreq7 & ~n23288;
  assign n23290 = ~n23233 & ~n23289;
  assign n23291 = n7924 & ~n23290;
  assign n23292 = ~n23201 & ~n23291;
  assign n23293 = n8214 & ~n23292;
  assign n23294 = ~n23146 & ~n23293;
  assign n23295 = n8202 & ~n23294;
  assign n23296 = ~n22996 & ~n23295;
  assign n23297 = n7920 & ~n23296;
  assign n23298 = ~n10014 & ~n23297;
  assign n23299 = ~n7728 & ~n23298;
  assign n23300 = ~n22743 & ~n23299;
  assign n23301 = n7723 & ~n23300;
  assign n23302 = ~n7723 & ~n23298;
  assign n23303 = ~n23301 & ~n23302;
  assign n23304 = n7714 & ~n23303;
  assign n23305 = n7723 & ~n23298;
  assign n23306 = ~n18610 & ~n20781;
  assign n23307 = ~controllable_hmaster1 & ~n23306;
  assign n23308 = ~n20744 & ~n23307;
  assign n23309 = ~controllable_hgrant6 & ~n23308;
  assign n23310 = ~n13849 & ~n23309;
  assign n23311 = controllable_hmaster0 & ~n23310;
  assign n23312 = ~n20848 & ~n23311;
  assign n23313 = ~controllable_hmaster3 & ~n23312;
  assign n23314 = ~n21474 & ~n23313;
  assign n23315 = i_hlock7 & ~n23314;
  assign n23316 = ~n20854 & ~n23307;
  assign n23317 = ~controllable_hgrant6 & ~n23316;
  assign n23318 = ~n13951 & ~n23317;
  assign n23319 = controllable_hmaster0 & ~n23318;
  assign n23320 = ~n20848 & ~n23319;
  assign n23321 = ~controllable_hmaster3 & ~n23320;
  assign n23322 = ~n21474 & ~n23321;
  assign n23323 = ~i_hlock7 & ~n23322;
  assign n23324 = ~n23315 & ~n23323;
  assign n23325 = i_hbusreq7 & ~n23324;
  assign n23326 = i_hbusreq8 & ~n23312;
  assign n23327 = i_hbusreq6 & ~n23308;
  assign n23328 = i_hlock5 & ~n21056;
  assign n23329 = ~i_hlock5 & ~n21099;
  assign n23330 = ~n23328 & ~n23329;
  assign n23331 = ~i_hbusreq5 & ~n23330;
  assign n23332 = ~n18941 & ~n23331;
  assign n23333 = ~controllable_hgrant5 & ~n23332;
  assign n23334 = ~n15020 & ~n23333;
  assign n23335 = controllable_hmaster2 & ~n23334;
  assign n23336 = ~n21279 & ~n23335;
  assign n23337 = ~controllable_hmaster1 & ~n23336;
  assign n23338 = ~n21206 & ~n23337;
  assign n23339 = ~i_hbusreq6 & ~n23338;
  assign n23340 = ~n23327 & ~n23339;
  assign n23341 = ~controllable_hgrant6 & ~n23340;
  assign n23342 = ~n15417 & ~n23341;
  assign n23343 = controllable_hmaster0 & ~n23342;
  assign n23344 = ~n21424 & ~n23343;
  assign n23345 = ~i_hbusreq8 & ~n23344;
  assign n23346 = ~n23326 & ~n23345;
  assign n23347 = ~controllable_hmaster3 & ~n23346;
  assign n23348 = ~n21525 & ~n23347;
  assign n23349 = i_hlock7 & ~n23348;
  assign n23350 = i_hbusreq8 & ~n23320;
  assign n23351 = i_hbusreq6 & ~n23316;
  assign n23352 = ~n21434 & ~n23337;
  assign n23353 = ~i_hbusreq6 & ~n23352;
  assign n23354 = ~n23351 & ~n23353;
  assign n23355 = ~controllable_hgrant6 & ~n23354;
  assign n23356 = ~n15440 & ~n23355;
  assign n23357 = controllable_hmaster0 & ~n23356;
  assign n23358 = ~n21424 & ~n23357;
  assign n23359 = ~i_hbusreq8 & ~n23358;
  assign n23360 = ~n23350 & ~n23359;
  assign n23361 = ~controllable_hmaster3 & ~n23360;
  assign n23362 = ~n21525 & ~n23361;
  assign n23363 = ~i_hlock7 & ~n23362;
  assign n23364 = ~n23349 & ~n23363;
  assign n23365 = ~i_hbusreq7 & ~n23364;
  assign n23366 = ~n23325 & ~n23365;
  assign n23367 = n7924 & ~n23366;
  assign n23368 = ~n22797 & ~n23367;
  assign n23369 = ~n8214 & ~n23368;
  assign n23370 = ~n18666 & ~n20833;
  assign n23371 = ~controllable_hmaster1 & ~n23370;
  assign n23372 = ~n20807 & ~n23371;
  assign n23373 = i_hlock6 & ~n23372;
  assign n23374 = ~n20842 & ~n23371;
  assign n23375 = ~i_hlock6 & ~n23374;
  assign n23376 = ~n23373 & ~n23375;
  assign n23377 = ~controllable_hgrant6 & ~n23376;
  assign n23378 = ~n13894 & ~n23377;
  assign n23379 = ~controllable_hmaster0 & ~n23378;
  assign n23380 = ~n20787 & ~n23379;
  assign n23381 = ~controllable_hmaster3 & ~n23380;
  assign n23382 = ~n21474 & ~n23381;
  assign n23383 = i_hlock7 & ~n23382;
  assign n23384 = ~n20858 & ~n23379;
  assign n23385 = ~controllable_hmaster3 & ~n23384;
  assign n23386 = ~n21474 & ~n23385;
  assign n23387 = ~i_hlock7 & ~n23386;
  assign n23388 = ~n23383 & ~n23387;
  assign n23389 = i_hbusreq7 & ~n23388;
  assign n23390 = i_hbusreq8 & ~n23380;
  assign n23391 = i_hbusreq6 & ~n23376;
  assign n23392 = i_hlock4 & ~n21052;
  assign n23393 = ~i_hlock4 & ~n21095;
  assign n23394 = ~n23392 & ~n23393;
  assign n23395 = ~i_hbusreq4 & ~n23394;
  assign n23396 = ~n19044 & ~n23395;
  assign n23397 = ~controllable_hgrant4 & ~n23396;
  assign n23398 = ~n15091 & ~n23397;
  assign n23399 = ~i_hbusreq5 & ~n23398;
  assign n23400 = ~n19043 & ~n23399;
  assign n23401 = ~controllable_hgrant5 & ~n23400;
  assign n23402 = ~n15090 & ~n23401;
  assign n23403 = controllable_hmaster2 & ~n23402;
  assign n23404 = ~n21404 & ~n23403;
  assign n23405 = ~controllable_hmaster1 & ~n23404;
  assign n23406 = ~n21329 & ~n23405;
  assign n23407 = i_hlock6 & ~n23406;
  assign n23408 = ~n21416 & ~n23405;
  assign n23409 = ~i_hlock6 & ~n23408;
  assign n23410 = ~n23407 & ~n23409;
  assign n23411 = ~i_hbusreq6 & ~n23410;
  assign n23412 = ~n23391 & ~n23411;
  assign n23413 = ~controllable_hgrant6 & ~n23412;
  assign n23414 = ~n15467 & ~n23413;
  assign n23415 = ~controllable_hmaster0 & ~n23414;
  assign n23416 = ~n21287 & ~n23415;
  assign n23417 = ~i_hbusreq8 & ~n23416;
  assign n23418 = ~n23390 & ~n23417;
  assign n23419 = ~controllable_hmaster3 & ~n23418;
  assign n23420 = ~n21525 & ~n23419;
  assign n23421 = i_hlock7 & ~n23420;
  assign n23422 = i_hbusreq8 & ~n23384;
  assign n23423 = ~n21440 & ~n23415;
  assign n23424 = ~i_hbusreq8 & ~n23423;
  assign n23425 = ~n23422 & ~n23424;
  assign n23426 = ~controllable_hmaster3 & ~n23425;
  assign n23427 = ~n21525 & ~n23426;
  assign n23428 = ~i_hlock7 & ~n23427;
  assign n23429 = ~n23421 & ~n23428;
  assign n23430 = ~i_hbusreq7 & ~n23429;
  assign n23431 = ~n23389 & ~n23430;
  assign n23432 = n7924 & ~n23431;
  assign n23433 = ~n22919 & ~n23432;
  assign n23434 = n8214 & ~n23433;
  assign n23435 = ~n23369 & ~n23434;
  assign n23436 = ~n8202 & ~n23435;
  assign n23437 = ~n18602 & ~n20718;
  assign n23438 = controllable_hmaster1 & ~n23437;
  assign n23439 = ~n20783 & ~n23438;
  assign n23440 = ~controllable_hgrant6 & ~n23439;
  assign n23441 = ~n13849 & ~n23440;
  assign n23442 = controllable_hmaster0 & ~n23441;
  assign n23443 = ~n20848 & ~n23442;
  assign n23444 = ~controllable_hmaster3 & ~n23443;
  assign n23445 = ~n21474 & ~n23444;
  assign n23446 = i_hlock7 & ~n23445;
  assign n23447 = ~n18602 & ~n20840;
  assign n23448 = controllable_hmaster1 & ~n23447;
  assign n23449 = ~n20783 & ~n23448;
  assign n23450 = ~controllable_hgrant6 & ~n23449;
  assign n23451 = ~n13951 & ~n23450;
  assign n23452 = controllable_hmaster0 & ~n23451;
  assign n23453 = ~n20848 & ~n23452;
  assign n23454 = ~controllable_hmaster3 & ~n23453;
  assign n23455 = ~n21474 & ~n23454;
  assign n23456 = ~i_hlock7 & ~n23455;
  assign n23457 = ~n23446 & ~n23456;
  assign n23458 = i_hbusreq7 & ~n23457;
  assign n23459 = i_hbusreq8 & ~n23443;
  assign n23460 = i_hbusreq6 & ~n23439;
  assign n23461 = i_hlock3 & ~n21026;
  assign n23462 = ~i_hlock3 & ~n21077;
  assign n23463 = ~n23461 & ~n23462;
  assign n23464 = ~i_hbusreq3 & ~n23463;
  assign n23465 = ~n18909 & ~n23464;
  assign n23466 = ~controllable_hgrant3 & ~n23465;
  assign n23467 = ~n14999 & ~n23466;
  assign n23468 = i_hlock9 & ~n23467;
  assign n23469 = i_hlock3 & ~n21044;
  assign n23470 = ~i_hlock3 & ~n21087;
  assign n23471 = ~n23469 & ~n23470;
  assign n23472 = ~i_hbusreq3 & ~n23471;
  assign n23473 = ~n18918 & ~n23472;
  assign n23474 = ~controllable_hgrant3 & ~n23473;
  assign n23475 = ~n14999 & ~n23474;
  assign n23476 = ~i_hlock9 & ~n23475;
  assign n23477 = ~n23468 & ~n23476;
  assign n23478 = ~i_hbusreq9 & ~n23477;
  assign n23479 = ~n18908 & ~n23478;
  assign n23480 = ~i_hbusreq4 & ~n23479;
  assign n23481 = ~n18907 & ~n23480;
  assign n23482 = ~controllable_hgrant4 & ~n23481;
  assign n23483 = ~n14998 & ~n23482;
  assign n23484 = ~i_hbusreq5 & ~n23483;
  assign n23485 = ~n18906 & ~n23484;
  assign n23486 = ~controllable_hgrant5 & ~n23485;
  assign n23487 = ~n14997 & ~n23486;
  assign n23488 = ~controllable_hmaster2 & ~n23487;
  assign n23489 = ~n21159 & ~n23488;
  assign n23490 = controllable_hmaster1 & ~n23489;
  assign n23491 = ~n21281 & ~n23490;
  assign n23492 = ~i_hbusreq6 & ~n23491;
  assign n23493 = ~n23460 & ~n23492;
  assign n23494 = ~controllable_hgrant6 & ~n23493;
  assign n23495 = ~n15520 & ~n23494;
  assign n23496 = controllable_hmaster0 & ~n23495;
  assign n23497 = ~n21424 & ~n23496;
  assign n23498 = ~i_hbusreq8 & ~n23497;
  assign n23499 = ~n23459 & ~n23498;
  assign n23500 = ~controllable_hmaster3 & ~n23499;
  assign n23501 = ~n21525 & ~n23500;
  assign n23502 = i_hlock7 & ~n23501;
  assign n23503 = i_hbusreq8 & ~n23453;
  assign n23504 = i_hbusreq6 & ~n23449;
  assign n23505 = ~n21414 & ~n23488;
  assign n23506 = controllable_hmaster1 & ~n23505;
  assign n23507 = ~n21281 & ~n23506;
  assign n23508 = ~i_hbusreq6 & ~n23507;
  assign n23509 = ~n23504 & ~n23508;
  assign n23510 = ~controllable_hgrant6 & ~n23509;
  assign n23511 = ~n15553 & ~n23510;
  assign n23512 = controllable_hmaster0 & ~n23511;
  assign n23513 = ~n21424 & ~n23512;
  assign n23514 = ~i_hbusreq8 & ~n23513;
  assign n23515 = ~n23503 & ~n23514;
  assign n23516 = ~controllable_hmaster3 & ~n23515;
  assign n23517 = ~n21525 & ~n23516;
  assign n23518 = ~i_hlock7 & ~n23517;
  assign n23519 = ~n23502 & ~n23518;
  assign n23520 = ~i_hbusreq7 & ~n23519;
  assign n23521 = ~n23458 & ~n23520;
  assign n23522 = n7924 & ~n23521;
  assign n23523 = ~n23054 & ~n23522;
  assign n23524 = ~n8214 & ~n23523;
  assign n23525 = ~n18656 & ~n20718;
  assign n23526 = controllable_hmaster1 & ~n23525;
  assign n23527 = ~n20835 & ~n23526;
  assign n23528 = i_hlock6 & ~n23527;
  assign n23529 = ~n18656 & ~n20840;
  assign n23530 = controllable_hmaster1 & ~n23529;
  assign n23531 = ~n20835 & ~n23530;
  assign n23532 = ~i_hlock6 & ~n23531;
  assign n23533 = ~n23528 & ~n23532;
  assign n23534 = ~controllable_hgrant6 & ~n23533;
  assign n23535 = ~n13894 & ~n23534;
  assign n23536 = ~controllable_hmaster0 & ~n23535;
  assign n23537 = ~n20787 & ~n23536;
  assign n23538 = ~controllable_hmaster3 & ~n23537;
  assign n23539 = ~n21474 & ~n23538;
  assign n23540 = i_hlock7 & ~n23539;
  assign n23541 = ~n20858 & ~n23536;
  assign n23542 = ~controllable_hmaster3 & ~n23541;
  assign n23543 = ~n21474 & ~n23542;
  assign n23544 = ~i_hlock7 & ~n23543;
  assign n23545 = ~n23540 & ~n23544;
  assign n23546 = i_hbusreq7 & ~n23545;
  assign n23547 = i_hbusreq8 & ~n23537;
  assign n23548 = i_hbusreq6 & ~n23533;
  assign n23549 = ~n9379 & ~n21021;
  assign n23550 = ~i_hbusreq1 & ~n23549;
  assign n23551 = ~n19006 & ~n23550;
  assign n23552 = ~controllable_hgrant1 & ~n23551;
  assign n23553 = ~n15067 & ~n23552;
  assign n23554 = ~i_hbusreq3 & ~n23553;
  assign n23555 = ~n19005 & ~n23554;
  assign n23556 = ~controllable_hgrant3 & ~n23555;
  assign n23557 = ~n15066 & ~n23556;
  assign n23558 = i_hlock9 & ~n23557;
  assign n23559 = ~n9379 & ~n21039;
  assign n23560 = ~i_hbusreq1 & ~n23559;
  assign n23561 = ~n19018 & ~n23560;
  assign n23562 = ~controllable_hgrant1 & ~n23561;
  assign n23563 = ~n15067 & ~n23562;
  assign n23564 = ~i_hbusreq3 & ~n23563;
  assign n23565 = ~n19017 & ~n23564;
  assign n23566 = ~controllable_hgrant3 & ~n23565;
  assign n23567 = ~n15066 & ~n23566;
  assign n23568 = ~i_hlock9 & ~n23567;
  assign n23569 = ~n23558 & ~n23568;
  assign n23570 = ~i_hbusreq9 & ~n23569;
  assign n23571 = ~n19004 & ~n23570;
  assign n23572 = ~i_hbusreq4 & ~n23571;
  assign n23573 = ~n19003 & ~n23572;
  assign n23574 = ~controllable_hgrant4 & ~n23573;
  assign n23575 = ~n15065 & ~n23574;
  assign n23576 = ~i_hbusreq5 & ~n23575;
  assign n23577 = ~n19002 & ~n23576;
  assign n23578 = ~controllable_hgrant5 & ~n23577;
  assign n23579 = ~n15064 & ~n23578;
  assign n23580 = ~controllable_hmaster2 & ~n23579;
  assign n23581 = ~n21159 & ~n23580;
  assign n23582 = controllable_hmaster1 & ~n23581;
  assign n23583 = ~n21406 & ~n23582;
  assign n23584 = i_hlock6 & ~n23583;
  assign n23585 = ~n21414 & ~n23580;
  assign n23586 = controllable_hmaster1 & ~n23585;
  assign n23587 = ~n21406 & ~n23586;
  assign n23588 = ~i_hlock6 & ~n23587;
  assign n23589 = ~n23584 & ~n23588;
  assign n23590 = ~i_hbusreq6 & ~n23589;
  assign n23591 = ~n23548 & ~n23590;
  assign n23592 = ~controllable_hgrant6 & ~n23591;
  assign n23593 = ~n15582 & ~n23592;
  assign n23594 = ~controllable_hmaster0 & ~n23593;
  assign n23595 = ~n21287 & ~n23594;
  assign n23596 = ~i_hbusreq8 & ~n23595;
  assign n23597 = ~n23547 & ~n23596;
  assign n23598 = ~controllable_hmaster3 & ~n23597;
  assign n23599 = ~n21525 & ~n23598;
  assign n23600 = i_hlock7 & ~n23599;
  assign n23601 = i_hbusreq8 & ~n23541;
  assign n23602 = ~n21440 & ~n23594;
  assign n23603 = ~i_hbusreq8 & ~n23602;
  assign n23604 = ~n23601 & ~n23603;
  assign n23605 = ~controllable_hmaster3 & ~n23604;
  assign n23606 = ~n21525 & ~n23605;
  assign n23607 = ~i_hlock7 & ~n23606;
  assign n23608 = ~n23600 & ~n23607;
  assign n23609 = ~i_hbusreq7 & ~n23608;
  assign n23610 = ~n23546 & ~n23609;
  assign n23611 = n7924 & ~n23610;
  assign n23612 = ~n23201 & ~n23611;
  assign n23613 = n8214 & ~n23612;
  assign n23614 = ~n23524 & ~n23613;
  assign n23615 = n8202 & ~n23614;
  assign n23616 = ~n23436 & ~n23615;
  assign n23617 = n7920 & ~n23616;
  assign n23618 = ~n16336 & ~n23617;
  assign n23619 = n7728 & ~n23618;
  assign n23620 = ~n22213 & ~n23619;
  assign n23621 = ~n7723 & ~n23620;
  assign n23622 = ~n23305 & ~n23621;
  assign n23623 = ~n7714 & ~n23622;
  assign n23624 = ~n23304 & ~n23623;
  assign n23625 = ~n7705 & ~n23624;
  assign n23626 = ~n22399 & ~n23625;
  assign n23627 = n7808 & ~n23626;
  assign n23628 = ~n22233 & ~n23627;
  assign n23629 = ~n8195 & ~n23628;
  assign n23630 = controllable_hgrant6 & ~n11132;
  assign n23631 = controllable_hgrant5 & ~n11128;
  assign n23632 = controllable_hgrant4 & ~n11128;
  assign n23633 = controllable_hgrant3 & ~n10380;
  assign n23634 = controllable_hgrant1 & ~n10380;
  assign n23635 = n7928 & ~n16129;
  assign n23636 = ~controllable_hgrant1 & ~n23635;
  assign n23637 = ~n23634 & ~n23636;
  assign n23638 = ~controllable_hgrant3 & ~n23637;
  assign n23639 = ~n23633 & ~n23638;
  assign n23640 = i_hlock9 & ~n23639;
  assign n23641 = controllable_hgrant3 & ~n10384;
  assign n23642 = controllable_hgrant1 & ~n10384;
  assign n23643 = n7928 & ~n16147;
  assign n23644 = ~controllable_hgrant1 & ~n23643;
  assign n23645 = ~n23642 & ~n23644;
  assign n23646 = ~controllable_hgrant3 & ~n23645;
  assign n23647 = ~n23641 & ~n23646;
  assign n23648 = ~i_hlock9 & ~n23647;
  assign n23649 = ~n23640 & ~n23648;
  assign n23650 = ~controllable_hgrant4 & ~n23649;
  assign n23651 = ~n23632 & ~n23650;
  assign n23652 = ~controllable_hgrant5 & ~n23651;
  assign n23653 = ~n23631 & ~n23652;
  assign n23654 = ~controllable_hmaster2 & ~n23653;
  assign n23655 = ~n10105 & ~n23654;
  assign n23656 = ~controllable_hmaster1 & ~n23655;
  assign n23657 = ~n10053 & ~n23656;
  assign n23658 = ~controllable_hgrant6 & ~n23657;
  assign n23659 = ~n23630 & ~n23658;
  assign n23660 = controllable_hmaster0 & ~n23659;
  assign n23661 = ~n11134 & ~n23660;
  assign n23662 = controllable_hmaster3 & ~n23661;
  assign n23663 = ~n10447 & ~n23662;
  assign n23664 = i_hbusreq7 & ~n23663;
  assign n23665 = i_hbusreq8 & ~n23661;
  assign n23666 = controllable_hgrant6 & ~n11158;
  assign n23667 = i_hbusreq6 & ~n23657;
  assign n23668 = controllable_hgrant5 & ~n11152;
  assign n23669 = i_hbusreq5 & ~n23651;
  assign n23670 = controllable_hgrant4 & ~n11150;
  assign n23671 = i_hbusreq4 & ~n23649;
  assign n23672 = i_hbusreq9 & ~n23649;
  assign n23673 = controllable_hgrant3 & ~n10497;
  assign n23674 = i_hbusreq3 & ~n23637;
  assign n23675 = controllable_hgrant1 & ~n10469;
  assign n23676 = i_hbusreq1 & ~n23635;
  assign n23677 = n7928 & ~n16192;
  assign n23678 = ~i_hbusreq1 & ~n23677;
  assign n23679 = ~n23676 & ~n23678;
  assign n23680 = ~controllable_hgrant1 & ~n23679;
  assign n23681 = ~n23675 & ~n23680;
  assign n23682 = ~i_hbusreq3 & ~n23681;
  assign n23683 = ~n23674 & ~n23682;
  assign n23684 = ~controllable_hgrant3 & ~n23683;
  assign n23685 = ~n23673 & ~n23684;
  assign n23686 = i_hlock9 & ~n23685;
  assign n23687 = controllable_hgrant3 & ~n10509;
  assign n23688 = i_hbusreq3 & ~n23645;
  assign n23689 = controllable_hgrant1 & ~n10476;
  assign n23690 = i_hbusreq1 & ~n23643;
  assign n23691 = n7928 & ~n16217;
  assign n23692 = ~i_hbusreq1 & ~n23691;
  assign n23693 = ~n23690 & ~n23692;
  assign n23694 = ~controllable_hgrant1 & ~n23693;
  assign n23695 = ~n23689 & ~n23694;
  assign n23696 = ~i_hbusreq3 & ~n23695;
  assign n23697 = ~n23688 & ~n23696;
  assign n23698 = ~controllable_hgrant3 & ~n23697;
  assign n23699 = ~n23687 & ~n23698;
  assign n23700 = ~i_hlock9 & ~n23699;
  assign n23701 = ~n23686 & ~n23700;
  assign n23702 = ~i_hbusreq9 & ~n23701;
  assign n23703 = ~n23672 & ~n23702;
  assign n23704 = ~i_hbusreq4 & ~n23703;
  assign n23705 = ~n23671 & ~n23704;
  assign n23706 = ~controllable_hgrant4 & ~n23705;
  assign n23707 = ~n23670 & ~n23706;
  assign n23708 = ~i_hbusreq5 & ~n23707;
  assign n23709 = ~n23669 & ~n23708;
  assign n23710 = ~controllable_hgrant5 & ~n23709;
  assign n23711 = ~n23668 & ~n23710;
  assign n23712 = ~controllable_hmaster2 & ~n23711;
  assign n23713 = ~n10116 & ~n23712;
  assign n23714 = ~controllable_hmaster1 & ~n23713;
  assign n23715 = ~n10064 & ~n23714;
  assign n23716 = ~i_hbusreq6 & ~n23715;
  assign n23717 = ~n23667 & ~n23716;
  assign n23718 = ~controllable_hgrant6 & ~n23717;
  assign n23719 = ~n23666 & ~n23718;
  assign n23720 = controllable_hmaster0 & ~n23719;
  assign n23721 = ~n11160 & ~n23720;
  assign n23722 = ~i_hbusreq8 & ~n23721;
  assign n23723 = ~n23665 & ~n23722;
  assign n23724 = controllable_hmaster3 & ~n23723;
  assign n23725 = ~n10621 & ~n23724;
  assign n23726 = ~i_hbusreq7 & ~n23725;
  assign n23727 = ~n23664 & ~n23726;
  assign n23728 = n7924 & ~n23727;
  assign n23729 = ~n10375 & ~n23728;
  assign n23730 = n8214 & ~n23729;
  assign n23731 = n8214 & ~n23730;
  assign n23732 = n8202 & ~n23731;
  assign n23733 = ~n10332 & ~n23732;
  assign n23734 = n7728 & ~n23733;
  assign n23735 = n8214 & ~n16335;
  assign n23736 = ~n8336 & ~n23735;
  assign n23737 = n8202 & ~n23736;
  assign n23738 = ~n10649 & ~n23737;
  assign n23739 = ~n7728 & ~n23738;
  assign n23740 = ~n23734 & ~n23739;
  assign n23741 = ~n7723 & ~n23740;
  assign n23742 = ~n7723 & ~n23741;
  assign n23743 = ~n7714 & ~n23742;
  assign n23744 = ~n7714 & ~n23743;
  assign n23745 = n7705 & ~n23744;
  assign n23746 = n7723 & ~n23738;
  assign n23747 = n7920 & ~n23738;
  assign n23748 = ~n16336 & ~n23747;
  assign n23749 = ~n7723 & ~n23748;
  assign n23750 = ~n23746 & ~n23749;
  assign n23751 = n7714 & ~n23750;
  assign n23752 = ~n16342 & ~n23751;
  assign n23753 = ~n7705 & ~n23752;
  assign n23754 = ~n23745 & ~n23753;
  assign n23755 = ~n7808 & ~n23754;
  assign n23756 = ~n7920 & ~n23733;
  assign n23757 = controllable_hgrant6 & ~n10674;
  assign n23758 = ~controllable_hmaster2 & ~n18143;
  assign n23759 = ~controllable_hmaster1 & ~n23758;
  assign n23760 = ~controllable_hmaster1 & ~n23759;
  assign n23761 = ~controllable_hgrant6 & ~n23760;
  assign n23762 = ~n23757 & ~n23761;
  assign n23763 = controllable_hmaster0 & ~n23762;
  assign n23764 = controllable_hmaster0 & ~n23763;
  assign n23765 = ~controllable_hmaster3 & ~n23764;
  assign n23766 = ~controllable_hmaster3 & ~n23765;
  assign n23767 = i_hbusreq7 & ~n23766;
  assign n23768 = i_hbusreq8 & ~n23764;
  assign n23769 = controllable_hgrant6 & ~n10686;
  assign n23770 = i_hbusreq6 & ~n23760;
  assign n23771 = ~controllable_hmaster2 & ~n21731;
  assign n23772 = ~controllable_hmaster1 & ~n23771;
  assign n23773 = ~controllable_hmaster1 & ~n23772;
  assign n23774 = ~i_hbusreq6 & ~n23773;
  assign n23775 = ~n23770 & ~n23774;
  assign n23776 = ~controllable_hgrant6 & ~n23775;
  assign n23777 = ~n23769 & ~n23776;
  assign n23778 = controllable_hmaster0 & ~n23777;
  assign n23779 = controllable_hmaster0 & ~n23778;
  assign n23780 = ~i_hbusreq8 & ~n23779;
  assign n23781 = ~n23768 & ~n23780;
  assign n23782 = ~controllable_hmaster3 & ~n23781;
  assign n23783 = ~controllable_hmaster3 & ~n23782;
  assign n23784 = ~i_hbusreq7 & ~n23783;
  assign n23785 = ~n23767 & ~n23784;
  assign n23786 = ~n8214 & ~n23785;
  assign n23787 = controllable_hgrant6 & ~n10698;
  assign n23788 = ~controllable_hmaster2 & ~n18179;
  assign n23789 = ~controllable_hmaster1 & ~n23788;
  assign n23790 = ~controllable_hmaster1 & ~n23789;
  assign n23791 = ~controllable_hgrant6 & ~n23790;
  assign n23792 = ~n23787 & ~n23791;
  assign n23793 = ~controllable_hmaster0 & ~n23792;
  assign n23794 = ~controllable_hmaster0 & ~n23793;
  assign n23795 = ~controllable_hmaster3 & ~n23794;
  assign n23796 = ~controllable_hmaster3 & ~n23795;
  assign n23797 = i_hbusreq7 & ~n23796;
  assign n23798 = i_hbusreq8 & ~n23794;
  assign n23799 = controllable_hgrant6 & ~n10710;
  assign n23800 = i_hbusreq6 & ~n23790;
  assign n23801 = ~controllable_hmaster2 & ~n21795;
  assign n23802 = ~controllable_hmaster1 & ~n23801;
  assign n23803 = ~controllable_hmaster1 & ~n23802;
  assign n23804 = ~i_hbusreq6 & ~n23803;
  assign n23805 = ~n23800 & ~n23804;
  assign n23806 = ~controllable_hgrant6 & ~n23805;
  assign n23807 = ~n23799 & ~n23806;
  assign n23808 = ~controllable_hmaster0 & ~n23807;
  assign n23809 = ~controllable_hmaster0 & ~n23808;
  assign n23810 = ~i_hbusreq8 & ~n23809;
  assign n23811 = ~n23798 & ~n23810;
  assign n23812 = ~controllable_hmaster3 & ~n23811;
  assign n23813 = ~controllable_hmaster3 & ~n23812;
  assign n23814 = ~i_hbusreq7 & ~n23813;
  assign n23815 = ~n23797 & ~n23814;
  assign n23816 = n8214 & ~n23815;
  assign n23817 = ~n23786 & ~n23816;
  assign n23818 = ~n8202 & ~n23817;
  assign n23819 = n7924 & ~n22209;
  assign n23820 = ~n8214 & ~n23819;
  assign n23821 = n7928 & ~n17314;
  assign n23822 = n7928 & ~n23821;
  assign n23823 = ~controllable_hgrant1 & ~n23822;
  assign n23824 = ~n13179 & ~n23823;
  assign n23825 = ~controllable_hgrant3 & ~n23824;
  assign n23826 = ~n13178 & ~n23825;
  assign n23827 = ~controllable_hgrant4 & ~n23826;
  assign n23828 = ~n13177 & ~n23827;
  assign n23829 = ~controllable_hgrant5 & ~n23828;
  assign n23830 = ~n13176 & ~n23829;
  assign n23831 = controllable_hmaster1 & ~n23830;
  assign n23832 = controllable_hmaster2 & ~n23830;
  assign n23833 = n7928 & ~n16354;
  assign n23834 = ~controllable_hgrant1 & ~n23833;
  assign n23835 = ~n13179 & ~n23834;
  assign n23836 = ~controllable_hgrant3 & ~n23835;
  assign n23837 = ~n13178 & ~n23836;
  assign n23838 = ~controllable_hgrant4 & ~n23837;
  assign n23839 = ~n13177 & ~n23838;
  assign n23840 = ~controllable_hgrant5 & ~n23839;
  assign n23841 = ~n13176 & ~n23840;
  assign n23842 = ~controllable_hmaster2 & ~n23841;
  assign n23843 = ~n23832 & ~n23842;
  assign n23844 = ~controllable_hmaster1 & ~n23843;
  assign n23845 = ~n23831 & ~n23844;
  assign n23846 = ~controllable_hgrant6 & ~n23845;
  assign n23847 = ~n13198 & ~n23846;
  assign n23848 = controllable_hmaster0 & ~n23847;
  assign n23849 = ~n17340 & ~n23832;
  assign n23850 = ~controllable_hmaster1 & ~n23849;
  assign n23851 = ~n23831 & ~n23850;
  assign n23852 = ~controllable_hgrant6 & ~n23851;
  assign n23853 = ~n13198 & ~n23852;
  assign n23854 = ~controllable_hmaster0 & ~n23853;
  assign n23855 = ~n23848 & ~n23854;
  assign n23856 = controllable_hmaster3 & ~n23855;
  assign n23857 = ~n17351 & ~n23856;
  assign n23858 = i_hbusreq7 & ~n23857;
  assign n23859 = i_hbusreq8 & ~n23855;
  assign n23860 = i_hbusreq6 & ~n23845;
  assign n23861 = i_hbusreq5 & ~n23828;
  assign n23862 = i_hbusreq4 & ~n23826;
  assign n23863 = i_hbusreq9 & ~n23826;
  assign n23864 = i_hbusreq3 & ~n23824;
  assign n23865 = i_hbusreq1 & ~n23822;
  assign n23866 = n7928 & ~n21629;
  assign n23867 = n7928 & ~n23866;
  assign n23868 = ~i_hbusreq1 & ~n23867;
  assign n23869 = ~n23865 & ~n23868;
  assign n23870 = ~controllable_hgrant1 & ~n23869;
  assign n23871 = ~n15730 & ~n23870;
  assign n23872 = ~i_hbusreq3 & ~n23871;
  assign n23873 = ~n23864 & ~n23872;
  assign n23874 = ~controllable_hgrant3 & ~n23873;
  assign n23875 = ~n15729 & ~n23874;
  assign n23876 = ~i_hbusreq9 & ~n23875;
  assign n23877 = ~n23863 & ~n23876;
  assign n23878 = ~i_hbusreq4 & ~n23877;
  assign n23879 = ~n23862 & ~n23878;
  assign n23880 = ~controllable_hgrant4 & ~n23879;
  assign n23881 = ~n15728 & ~n23880;
  assign n23882 = ~i_hbusreq5 & ~n23881;
  assign n23883 = ~n23861 & ~n23882;
  assign n23884 = ~controllable_hgrant5 & ~n23883;
  assign n23885 = ~n15727 & ~n23884;
  assign n23886 = controllable_hmaster1 & ~n23885;
  assign n23887 = controllable_hmaster2 & ~n23885;
  assign n23888 = i_hbusreq5 & ~n23839;
  assign n23889 = i_hbusreq4 & ~n23837;
  assign n23890 = i_hbusreq9 & ~n23837;
  assign n23891 = i_hbusreq3 & ~n23835;
  assign n23892 = i_hbusreq1 & ~n23833;
  assign n23893 = n7928 & ~n16418;
  assign n23894 = ~i_hbusreq1 & ~n23893;
  assign n23895 = ~n23892 & ~n23894;
  assign n23896 = ~controllable_hgrant1 & ~n23895;
  assign n23897 = ~n15677 & ~n23896;
  assign n23898 = ~i_hbusreq3 & ~n23897;
  assign n23899 = ~n23891 & ~n23898;
  assign n23900 = ~controllable_hgrant3 & ~n23899;
  assign n23901 = ~n15676 & ~n23900;
  assign n23902 = ~i_hbusreq9 & ~n23901;
  assign n23903 = ~n23890 & ~n23902;
  assign n23904 = ~i_hbusreq4 & ~n23903;
  assign n23905 = ~n23889 & ~n23904;
  assign n23906 = ~controllable_hgrant4 & ~n23905;
  assign n23907 = ~n15675 & ~n23906;
  assign n23908 = ~i_hbusreq5 & ~n23907;
  assign n23909 = ~n23888 & ~n23908;
  assign n23910 = ~controllable_hgrant5 & ~n23909;
  assign n23911 = ~n15674 & ~n23910;
  assign n23912 = ~controllable_hmaster2 & ~n23911;
  assign n23913 = ~n23887 & ~n23912;
  assign n23914 = ~controllable_hmaster1 & ~n23913;
  assign n23915 = ~n23886 & ~n23914;
  assign n23916 = ~i_hbusreq6 & ~n23915;
  assign n23917 = ~n23860 & ~n23916;
  assign n23918 = ~controllable_hgrant6 & ~n23917;
  assign n23919 = ~n15672 & ~n23918;
  assign n23920 = controllable_hmaster0 & ~n23919;
  assign n23921 = i_hbusreq6 & ~n23851;
  assign n23922 = n7928 & ~n16817;
  assign n23923 = ~i_hbusreq1 & ~n23922;
  assign n23924 = ~n17406 & ~n23923;
  assign n23925 = ~controllable_hgrant1 & ~n23924;
  assign n23926 = ~n15677 & ~n23925;
  assign n23927 = ~i_hbusreq3 & ~n23926;
  assign n23928 = ~n17405 & ~n23927;
  assign n23929 = ~controllable_hgrant3 & ~n23928;
  assign n23930 = ~n15676 & ~n23929;
  assign n23931 = ~i_hbusreq9 & ~n23930;
  assign n23932 = ~n17404 & ~n23931;
  assign n23933 = ~i_hbusreq4 & ~n23932;
  assign n23934 = ~n17403 & ~n23933;
  assign n23935 = ~controllable_hgrant4 & ~n23934;
  assign n23936 = ~n15675 & ~n23935;
  assign n23937 = ~i_hbusreq5 & ~n23936;
  assign n23938 = ~n17402 & ~n23937;
  assign n23939 = ~controllable_hgrant5 & ~n23938;
  assign n23940 = ~n15674 & ~n23939;
  assign n23941 = ~controllable_hmaster2 & ~n23940;
  assign n23942 = ~n23887 & ~n23941;
  assign n23943 = ~controllable_hmaster1 & ~n23942;
  assign n23944 = ~n23886 & ~n23943;
  assign n23945 = ~i_hbusreq6 & ~n23944;
  assign n23946 = ~n23921 & ~n23945;
  assign n23947 = ~controllable_hgrant6 & ~n23946;
  assign n23948 = ~n15672 & ~n23947;
  assign n23949 = ~controllable_hmaster0 & ~n23948;
  assign n23950 = ~n23920 & ~n23949;
  assign n23951 = ~i_hbusreq8 & ~n23950;
  assign n23952 = ~n23859 & ~n23951;
  assign n23953 = controllable_hmaster3 & ~n23952;
  assign n23954 = ~i_hbusreq6 & ~n23940;
  assign n23955 = ~n17449 & ~n23954;
  assign n23956 = ~controllable_hgrant6 & ~n23955;
  assign n23957 = ~n15812 & ~n23956;
  assign n23958 = controllable_hmaster0 & ~n23957;
  assign n23959 = controllable_hmaster1 & ~n23940;
  assign n23960 = controllable_hmaster2 & ~n23940;
  assign n23961 = n7928 & ~n21775;
  assign n23962 = ~i_hbusreq1 & ~n23961;
  assign n23963 = ~n17406 & ~n23962;
  assign n23964 = ~controllable_hgrant1 & ~n23963;
  assign n23965 = ~n15824 & ~n23964;
  assign n23966 = ~i_hbusreq3 & ~n23965;
  assign n23967 = ~n17405 & ~n23966;
  assign n23968 = ~controllable_hgrant3 & ~n23967;
  assign n23969 = ~n15823 & ~n23968;
  assign n23970 = ~i_hbusreq9 & ~n23969;
  assign n23971 = ~n17404 & ~n23970;
  assign n23972 = ~i_hbusreq4 & ~n23971;
  assign n23973 = ~n17403 & ~n23972;
  assign n23974 = ~controllable_hgrant4 & ~n23973;
  assign n23975 = ~n15822 & ~n23974;
  assign n23976 = ~i_hbusreq5 & ~n23975;
  assign n23977 = ~n17402 & ~n23976;
  assign n23978 = ~controllable_hgrant5 & ~n23977;
  assign n23979 = ~n15821 & ~n23978;
  assign n23980 = ~controllable_hmaster2 & ~n23979;
  assign n23981 = ~n23960 & ~n23980;
  assign n23982 = ~controllable_hmaster1 & ~n23981;
  assign n23983 = ~n23959 & ~n23982;
  assign n23984 = ~i_hbusreq6 & ~n23983;
  assign n23985 = ~n17449 & ~n23984;
  assign n23986 = ~controllable_hgrant6 & ~n23985;
  assign n23987 = ~n15818 & ~n23986;
  assign n23988 = ~controllable_hmaster0 & ~n23987;
  assign n23989 = ~n23958 & ~n23988;
  assign n23990 = ~i_hbusreq8 & ~n23989;
  assign n23991 = ~n17448 & ~n23990;
  assign n23992 = ~controllable_hmaster3 & ~n23991;
  assign n23993 = ~n23953 & ~n23992;
  assign n23994 = ~i_hbusreq7 & ~n23993;
  assign n23995 = ~n23858 & ~n23994;
  assign n23996 = ~n7924 & ~n23995;
  assign n23997 = n7928 & ~n17469;
  assign n23998 = ~controllable_hgrant1 & ~n23997;
  assign n23999 = ~n13179 & ~n23998;
  assign n24000 = ~controllable_hgrant3 & ~n23999;
  assign n24001 = ~n13178 & ~n24000;
  assign n24002 = i_hlock9 & ~n24001;
  assign n24003 = n7928 & ~n17485;
  assign n24004 = ~controllable_hgrant1 & ~n24003;
  assign n24005 = ~n13179 & ~n24004;
  assign n24006 = ~controllable_hgrant3 & ~n24005;
  assign n24007 = ~n13178 & ~n24006;
  assign n24008 = ~i_hlock9 & ~n24007;
  assign n24009 = ~n24002 & ~n24008;
  assign n24010 = ~controllable_hgrant4 & ~n24009;
  assign n24011 = ~n13177 & ~n24010;
  assign n24012 = ~controllable_hgrant5 & ~n24011;
  assign n24013 = ~n13176 & ~n24012;
  assign n24014 = controllable_hmaster1 & ~n24013;
  assign n24015 = controllable_hmaster2 & ~n24013;
  assign n24016 = n7928 & ~n16510;
  assign n24017 = ~controllable_hgrant1 & ~n24016;
  assign n24018 = ~n13179 & ~n24017;
  assign n24019 = ~controllable_hgrant3 & ~n24018;
  assign n24020 = ~n13178 & ~n24019;
  assign n24021 = i_hlock9 & ~n24020;
  assign n24022 = n7928 & ~n16524;
  assign n24023 = ~controllable_hgrant1 & ~n24022;
  assign n24024 = ~n13179 & ~n24023;
  assign n24025 = ~controllable_hgrant3 & ~n24024;
  assign n24026 = ~n13178 & ~n24025;
  assign n24027 = ~i_hlock9 & ~n24026;
  assign n24028 = ~n24021 & ~n24027;
  assign n24029 = ~controllable_hgrant4 & ~n24028;
  assign n24030 = ~n13177 & ~n24029;
  assign n24031 = ~controllable_hgrant5 & ~n24030;
  assign n24032 = ~n13176 & ~n24031;
  assign n24033 = ~controllable_hmaster2 & ~n24032;
  assign n24034 = ~n24015 & ~n24033;
  assign n24035 = ~controllable_hmaster1 & ~n24034;
  assign n24036 = ~n24014 & ~n24035;
  assign n24037 = ~controllable_hgrant6 & ~n24036;
  assign n24038 = ~n13198 & ~n24037;
  assign n24039 = controllable_hmaster0 & ~n24038;
  assign n24040 = ~n17529 & ~n24015;
  assign n24041 = ~controllable_hmaster1 & ~n24040;
  assign n24042 = ~n24014 & ~n24041;
  assign n24043 = ~controllable_hgrant6 & ~n24042;
  assign n24044 = ~n13198 & ~n24043;
  assign n24045 = ~controllable_hmaster0 & ~n24044;
  assign n24046 = ~n24039 & ~n24045;
  assign n24047 = controllable_hmaster3 & ~n24046;
  assign n24048 = ~n17540 & ~n24047;
  assign n24049 = i_hbusreq7 & ~n24048;
  assign n24050 = i_hbusreq8 & ~n24046;
  assign n24051 = i_hbusreq6 & ~n24036;
  assign n24052 = i_hbusreq5 & ~n24011;
  assign n24053 = i_hbusreq4 & ~n24009;
  assign n24054 = i_hbusreq9 & ~n24009;
  assign n24055 = i_hbusreq3 & ~n23999;
  assign n24056 = i_hbusreq1 & ~n23997;
  assign n24057 = n7928 & ~n21857;
  assign n24058 = ~i_hbusreq1 & ~n24057;
  assign n24059 = ~n24056 & ~n24058;
  assign n24060 = ~controllable_hgrant1 & ~n24059;
  assign n24061 = ~n15730 & ~n24060;
  assign n24062 = ~i_hbusreq3 & ~n24061;
  assign n24063 = ~n24055 & ~n24062;
  assign n24064 = ~controllable_hgrant3 & ~n24063;
  assign n24065 = ~n15729 & ~n24064;
  assign n24066 = i_hlock9 & ~n24065;
  assign n24067 = i_hbusreq3 & ~n24005;
  assign n24068 = i_hbusreq1 & ~n24003;
  assign n24069 = n7928 & ~n21875;
  assign n24070 = ~i_hbusreq1 & ~n24069;
  assign n24071 = ~n24068 & ~n24070;
  assign n24072 = ~controllable_hgrant1 & ~n24071;
  assign n24073 = ~n15730 & ~n24072;
  assign n24074 = ~i_hbusreq3 & ~n24073;
  assign n24075 = ~n24067 & ~n24074;
  assign n24076 = ~controllable_hgrant3 & ~n24075;
  assign n24077 = ~n15729 & ~n24076;
  assign n24078 = ~i_hlock9 & ~n24077;
  assign n24079 = ~n24066 & ~n24078;
  assign n24080 = ~i_hbusreq9 & ~n24079;
  assign n24081 = ~n24054 & ~n24080;
  assign n24082 = ~i_hbusreq4 & ~n24081;
  assign n24083 = ~n24053 & ~n24082;
  assign n24084 = ~controllable_hgrant4 & ~n24083;
  assign n24085 = ~n15728 & ~n24084;
  assign n24086 = ~i_hbusreq5 & ~n24085;
  assign n24087 = ~n24052 & ~n24086;
  assign n24088 = ~controllable_hgrant5 & ~n24087;
  assign n24089 = ~n15727 & ~n24088;
  assign n24090 = controllable_hmaster1 & ~n24089;
  assign n24091 = controllable_hmaster2 & ~n24089;
  assign n24092 = i_hbusreq5 & ~n24030;
  assign n24093 = i_hbusreq4 & ~n24028;
  assign n24094 = i_hbusreq9 & ~n24028;
  assign n24095 = i_hbusreq3 & ~n24018;
  assign n24096 = i_hbusreq1 & ~n24016;
  assign n24097 = n7928 & ~n16649;
  assign n24098 = ~i_hbusreq1 & ~n24097;
  assign n24099 = ~n24096 & ~n24098;
  assign n24100 = ~controllable_hgrant1 & ~n24099;
  assign n24101 = ~n15677 & ~n24100;
  assign n24102 = ~i_hbusreq3 & ~n24101;
  assign n24103 = ~n24095 & ~n24102;
  assign n24104 = ~controllable_hgrant3 & ~n24103;
  assign n24105 = ~n15676 & ~n24104;
  assign n24106 = i_hlock9 & ~n24105;
  assign n24107 = i_hbusreq3 & ~n24024;
  assign n24108 = i_hbusreq1 & ~n24022;
  assign n24109 = n7928 & ~n16671;
  assign n24110 = ~i_hbusreq1 & ~n24109;
  assign n24111 = ~n24108 & ~n24110;
  assign n24112 = ~controllable_hgrant1 & ~n24111;
  assign n24113 = ~n15677 & ~n24112;
  assign n24114 = ~i_hbusreq3 & ~n24113;
  assign n24115 = ~n24107 & ~n24114;
  assign n24116 = ~controllable_hgrant3 & ~n24115;
  assign n24117 = ~n15676 & ~n24116;
  assign n24118 = ~i_hlock9 & ~n24117;
  assign n24119 = ~n24106 & ~n24118;
  assign n24120 = ~i_hbusreq9 & ~n24119;
  assign n24121 = ~n24094 & ~n24120;
  assign n24122 = ~i_hbusreq4 & ~n24121;
  assign n24123 = ~n24093 & ~n24122;
  assign n24124 = ~controllable_hgrant4 & ~n24123;
  assign n24125 = ~n15675 & ~n24124;
  assign n24126 = ~i_hbusreq5 & ~n24125;
  assign n24127 = ~n24092 & ~n24126;
  assign n24128 = ~controllable_hgrant5 & ~n24127;
  assign n24129 = ~n15674 & ~n24128;
  assign n24130 = ~controllable_hmaster2 & ~n24129;
  assign n24131 = ~n24091 & ~n24130;
  assign n24132 = ~controllable_hmaster1 & ~n24131;
  assign n24133 = ~n24090 & ~n24132;
  assign n24134 = ~i_hbusreq6 & ~n24133;
  assign n24135 = ~n24051 & ~n24134;
  assign n24136 = ~controllable_hgrant6 & ~n24135;
  assign n24137 = ~n15672 & ~n24136;
  assign n24138 = controllable_hmaster0 & ~n24137;
  assign n24139 = i_hbusreq6 & ~n24042;
  assign n24140 = n7928 & ~n21908;
  assign n24141 = ~i_hbusreq1 & ~n24140;
  assign n24142 = ~n17625 & ~n24141;
  assign n24143 = ~controllable_hgrant1 & ~n24142;
  assign n24144 = ~n15677 & ~n24143;
  assign n24145 = ~i_hbusreq3 & ~n24144;
  assign n24146 = ~n17624 & ~n24145;
  assign n24147 = ~controllable_hgrant3 & ~n24146;
  assign n24148 = ~n15676 & ~n24147;
  assign n24149 = i_hlock9 & ~n24148;
  assign n24150 = n7928 & ~n21920;
  assign n24151 = ~i_hbusreq1 & ~n24150;
  assign n24152 = ~n17653 & ~n24151;
  assign n24153 = ~controllable_hgrant1 & ~n24152;
  assign n24154 = ~n15677 & ~n24153;
  assign n24155 = ~i_hbusreq3 & ~n24154;
  assign n24156 = ~n17652 & ~n24155;
  assign n24157 = ~controllable_hgrant3 & ~n24156;
  assign n24158 = ~n15676 & ~n24157;
  assign n24159 = ~i_hlock9 & ~n24158;
  assign n24160 = ~n24149 & ~n24159;
  assign n24161 = ~i_hbusreq9 & ~n24160;
  assign n24162 = ~n17623 & ~n24161;
  assign n24163 = ~i_hbusreq4 & ~n24162;
  assign n24164 = ~n17622 & ~n24163;
  assign n24165 = ~controllable_hgrant4 & ~n24164;
  assign n24166 = ~n15675 & ~n24165;
  assign n24167 = ~i_hbusreq5 & ~n24166;
  assign n24168 = ~n17621 & ~n24167;
  assign n24169 = ~controllable_hgrant5 & ~n24168;
  assign n24170 = ~n15674 & ~n24169;
  assign n24171 = ~controllable_hmaster2 & ~n24170;
  assign n24172 = ~n24091 & ~n24171;
  assign n24173 = ~controllable_hmaster1 & ~n24172;
  assign n24174 = ~n24090 & ~n24173;
  assign n24175 = ~i_hbusreq6 & ~n24174;
  assign n24176 = ~n24139 & ~n24175;
  assign n24177 = ~controllable_hgrant6 & ~n24176;
  assign n24178 = ~n15672 & ~n24177;
  assign n24179 = ~controllable_hmaster0 & ~n24178;
  assign n24180 = ~n24138 & ~n24179;
  assign n24181 = ~i_hbusreq8 & ~n24180;
  assign n24182 = ~n24050 & ~n24181;
  assign n24183 = controllable_hmaster3 & ~n24182;
  assign n24184 = ~i_hbusreq6 & ~n24170;
  assign n24185 = ~n17691 & ~n24184;
  assign n24186 = ~controllable_hgrant6 & ~n24185;
  assign n24187 = ~n15812 & ~n24186;
  assign n24188 = controllable_hmaster0 & ~n24187;
  assign n24189 = controllable_hmaster1 & ~n24170;
  assign n24190 = controllable_hmaster2 & ~n24170;
  assign n24191 = n7928 & ~n22136;
  assign n24192 = ~i_hbusreq1 & ~n24191;
  assign n24193 = ~n17625 & ~n24192;
  assign n24194 = ~controllable_hgrant1 & ~n24193;
  assign n24195 = ~n15824 & ~n24194;
  assign n24196 = ~i_hbusreq3 & ~n24195;
  assign n24197 = ~n17624 & ~n24196;
  assign n24198 = ~controllable_hgrant3 & ~n24197;
  assign n24199 = ~n15823 & ~n24198;
  assign n24200 = i_hlock9 & ~n24199;
  assign n24201 = n7928 & ~n22148;
  assign n24202 = ~i_hbusreq1 & ~n24201;
  assign n24203 = ~n17653 & ~n24202;
  assign n24204 = ~controllable_hgrant1 & ~n24203;
  assign n24205 = ~n15824 & ~n24204;
  assign n24206 = ~i_hbusreq3 & ~n24205;
  assign n24207 = ~n17652 & ~n24206;
  assign n24208 = ~controllable_hgrant3 & ~n24207;
  assign n24209 = ~n15823 & ~n24208;
  assign n24210 = ~i_hlock9 & ~n24209;
  assign n24211 = ~n24200 & ~n24210;
  assign n24212 = ~i_hbusreq9 & ~n24211;
  assign n24213 = ~n17623 & ~n24212;
  assign n24214 = ~i_hbusreq4 & ~n24213;
  assign n24215 = ~n17622 & ~n24214;
  assign n24216 = ~controllable_hgrant4 & ~n24215;
  assign n24217 = ~n15822 & ~n24216;
  assign n24218 = ~i_hbusreq5 & ~n24217;
  assign n24219 = ~n17621 & ~n24218;
  assign n24220 = ~controllable_hgrant5 & ~n24219;
  assign n24221 = ~n15821 & ~n24220;
  assign n24222 = ~controllable_hmaster2 & ~n24221;
  assign n24223 = ~n24190 & ~n24222;
  assign n24224 = ~controllable_hmaster1 & ~n24223;
  assign n24225 = ~n24189 & ~n24224;
  assign n24226 = ~i_hbusreq6 & ~n24225;
  assign n24227 = ~n17691 & ~n24226;
  assign n24228 = ~controllable_hgrant6 & ~n24227;
  assign n24229 = ~n15818 & ~n24228;
  assign n24230 = ~controllable_hmaster0 & ~n24229;
  assign n24231 = ~n24188 & ~n24230;
  assign n24232 = ~i_hbusreq8 & ~n24231;
  assign n24233 = ~n17690 & ~n24232;
  assign n24234 = ~controllable_hmaster3 & ~n24233;
  assign n24235 = ~n24183 & ~n24234;
  assign n24236 = ~i_hbusreq7 & ~n24235;
  assign n24237 = ~n24049 & ~n24236;
  assign n24238 = n7924 & ~n24237;
  assign n24239 = ~n23996 & ~n24238;
  assign n24240 = n8214 & ~n24239;
  assign n24241 = ~n23820 & ~n24240;
  assign n24242 = n8202 & ~n24241;
  assign n24243 = ~n23818 & ~n24242;
  assign n24244 = n7920 & ~n24243;
  assign n24245 = ~n23756 & ~n24244;
  assign n24246 = n7728 & ~n24245;
  assign n24247 = ~n7920 & ~n23738;
  assign n24248 = ~n7743 & ~n23765;
  assign n24249 = i_hbusreq7 & ~n24248;
  assign n24250 = ~n7779 & ~n23782;
  assign n24251 = ~i_hbusreq7 & ~n24250;
  assign n24252 = ~n24249 & ~n24251;
  assign n24253 = ~n8214 & ~n24252;
  assign n24254 = ~n7743 & ~n23795;
  assign n24255 = i_hbusreq7 & ~n24254;
  assign n24256 = ~n7743 & ~n23812;
  assign n24257 = ~i_hbusreq7 & ~n24256;
  assign n24258 = ~n24255 & ~n24257;
  assign n24259 = n8214 & ~n24258;
  assign n24260 = ~n24253 & ~n24259;
  assign n24261 = ~n8202 & ~n24260;
  assign n24262 = controllable_hmaster3 & ~n17022;
  assign n24263 = controllable_hmaster3 & ~n24262;
  assign n24264 = ~n7924 & ~n24263;
  assign n24265 = ~n22209 & ~n24264;
  assign n24266 = ~n8214 & ~n24265;
  assign n24267 = n8214 & ~n22210;
  assign n24268 = ~n24266 & ~n24267;
  assign n24269 = n8202 & ~n24268;
  assign n24270 = ~n24261 & ~n24269;
  assign n24271 = n7920 & ~n24270;
  assign n24272 = ~n24247 & ~n24271;
  assign n24273 = ~n7728 & ~n24272;
  assign n24274 = ~n24246 & ~n24273;
  assign n24275 = ~n7723 & ~n24274;
  assign n24276 = ~n7723 & ~n24275;
  assign n24277 = ~n7714 & ~n24276;
  assign n24278 = ~n7714 & ~n24277;
  assign n24279 = n7705 & ~n24278;
  assign n24280 = ~n10105 & ~n18143;
  assign n24281 = ~controllable_hmaster1 & ~n24280;
  assign n24282 = ~n10053 & ~n24281;
  assign n24283 = ~controllable_hgrant6 & ~n24282;
  assign n24284 = ~n15890 & ~n24283;
  assign n24285 = controllable_hmaster0 & ~n24284;
  assign n24286 = ~n9099 & ~n24285;
  assign n24287 = ~controllable_hmaster3 & ~n24286;
  assign n24288 = ~n13651 & ~n24287;
  assign n24289 = i_hbusreq7 & ~n24288;
  assign n24290 = i_hbusreq8 & ~n24286;
  assign n24291 = i_hbusreq6 & ~n24282;
  assign n24292 = ~n10116 & ~n21731;
  assign n24293 = ~controllable_hmaster1 & ~n24292;
  assign n24294 = ~n10064 & ~n24293;
  assign n24295 = ~i_hbusreq6 & ~n24294;
  assign n24296 = ~n24291 & ~n24295;
  assign n24297 = ~controllable_hgrant6 & ~n24296;
  assign n24298 = ~n15902 & ~n24297;
  assign n24299 = controllable_hmaster0 & ~n24298;
  assign n24300 = ~n9127 & ~n24299;
  assign n24301 = ~i_hbusreq8 & ~n24300;
  assign n24302 = ~n24290 & ~n24301;
  assign n24303 = ~controllable_hmaster3 & ~n24302;
  assign n24304 = ~n13662 & ~n24303;
  assign n24305 = ~i_hbusreq7 & ~n24304;
  assign n24306 = ~n24289 & ~n24305;
  assign n24307 = ~n7924 & ~n24306;
  assign n24308 = i_hlock1 & ~n17767;
  assign n24309 = ~i_hlock1 & ~n17785;
  assign n24310 = ~n24308 & ~n24309;
  assign n24311 = ~controllable_hgrant1 & ~n24310;
  assign n24312 = ~n13875 & ~n24311;
  assign n24313 = ~controllable_hgrant3 & ~n24312;
  assign n24314 = ~n13874 & ~n24313;
  assign n24315 = ~controllable_hgrant4 & ~n24314;
  assign n24316 = ~n13873 & ~n24315;
  assign n24317 = ~controllable_hgrant5 & ~n24316;
  assign n24318 = ~n13872 & ~n24317;
  assign n24319 = ~controllable_hmaster2 & ~n24318;
  assign n24320 = ~n15294 & ~n24319;
  assign n24321 = ~controllable_hmaster1 & ~n24320;
  assign n24322 = ~n15194 & ~n24321;
  assign n24323 = ~controllable_hgrant6 & ~n24322;
  assign n24324 = ~n15890 & ~n24323;
  assign n24325 = controllable_hmaster0 & ~n24324;
  assign n24326 = ~n13682 & ~n24325;
  assign n24327 = ~controllable_hmaster3 & ~n24326;
  assign n24328 = ~n13672 & ~n24327;
  assign n24329 = i_hbusreq7 & ~n24328;
  assign n24330 = i_hbusreq8 & ~n24326;
  assign n24331 = i_hbusreq6 & ~n24322;
  assign n24332 = i_hbusreq5 & ~n24316;
  assign n24333 = i_hbusreq4 & ~n24314;
  assign n24334 = i_hbusreq9 & ~n24314;
  assign n24335 = i_hbusreq3 & ~n24312;
  assign n24336 = i_hbusreq1 & ~n24310;
  assign n24337 = i_hlock1 & ~n17832;
  assign n24338 = ~i_hlock1 & ~n17868;
  assign n24339 = ~n24337 & ~n24338;
  assign n24340 = ~i_hbusreq1 & ~n24339;
  assign n24341 = ~n24336 & ~n24340;
  assign n24342 = ~controllable_hgrant1 & ~n24341;
  assign n24343 = ~n15032 & ~n24342;
  assign n24344 = ~i_hbusreq3 & ~n24343;
  assign n24345 = ~n24335 & ~n24344;
  assign n24346 = ~controllable_hgrant3 & ~n24345;
  assign n24347 = ~n15031 & ~n24346;
  assign n24348 = ~i_hbusreq9 & ~n24347;
  assign n24349 = ~n24334 & ~n24348;
  assign n24350 = ~i_hbusreq4 & ~n24349;
  assign n24351 = ~n24333 & ~n24350;
  assign n24352 = ~controllable_hgrant4 & ~n24351;
  assign n24353 = ~n15030 & ~n24352;
  assign n24354 = ~i_hbusreq5 & ~n24353;
  assign n24355 = ~n24332 & ~n24354;
  assign n24356 = ~controllable_hgrant5 & ~n24355;
  assign n24357 = ~n15029 & ~n24356;
  assign n24358 = ~controllable_hmaster2 & ~n24357;
  assign n24359 = ~n15308 & ~n24358;
  assign n24360 = ~controllable_hmaster1 & ~n24359;
  assign n24361 = ~n15208 & ~n24360;
  assign n24362 = ~i_hbusreq6 & ~n24361;
  assign n24363 = ~n24331 & ~n24362;
  assign n24364 = ~controllable_hgrant6 & ~n24363;
  assign n24365 = ~n15902 & ~n24364;
  assign n24366 = controllable_hmaster0 & ~n24365;
  assign n24367 = ~n13728 & ~n24366;
  assign n24368 = ~i_hbusreq8 & ~n24367;
  assign n24369 = ~n24330 & ~n24368;
  assign n24370 = ~controllable_hmaster3 & ~n24369;
  assign n24371 = ~n13714 & ~n24370;
  assign n24372 = ~i_hbusreq7 & ~n24371;
  assign n24373 = ~n24329 & ~n24372;
  assign n24374 = n7924 & ~n24373;
  assign n24375 = ~n24307 & ~n24374;
  assign n24376 = ~n8214 & ~n24375;
  assign n24377 = ~n10105 & ~n18179;
  assign n24378 = ~controllable_hmaster1 & ~n24377;
  assign n24379 = ~n10053 & ~n24378;
  assign n24380 = ~controllable_hgrant6 & ~n24379;
  assign n24381 = ~n15964 & ~n24380;
  assign n24382 = ~controllable_hmaster0 & ~n24381;
  assign n24383 = ~n9152 & ~n24382;
  assign n24384 = ~controllable_hmaster3 & ~n24383;
  assign n24385 = ~n13651 & ~n24384;
  assign n24386 = i_hbusreq7 & ~n24385;
  assign n24387 = i_hbusreq8 & ~n24383;
  assign n24388 = i_hbusreq6 & ~n24379;
  assign n24389 = ~n10764 & ~n21795;
  assign n24390 = ~controllable_hmaster1 & ~n24389;
  assign n24391 = ~n10763 & ~n24390;
  assign n24392 = ~i_hbusreq6 & ~n24391;
  assign n24393 = ~n24388 & ~n24392;
  assign n24394 = ~controllable_hgrant6 & ~n24393;
  assign n24395 = ~n15996 & ~n24394;
  assign n24396 = ~controllable_hmaster0 & ~n24395;
  assign n24397 = ~n10762 & ~n24396;
  assign n24398 = ~i_hbusreq8 & ~n24397;
  assign n24399 = ~n24387 & ~n24398;
  assign n24400 = ~controllable_hmaster3 & ~n24399;
  assign n24401 = ~n15959 & ~n24400;
  assign n24402 = ~i_hbusreq7 & ~n24401;
  assign n24403 = ~n24386 & ~n24402;
  assign n24404 = ~n7924 & ~n24403;
  assign n24405 = ~n8440 & ~n17766;
  assign n24406 = ~controllable_hgrant1 & ~n24405;
  assign n24407 = ~n13924 & ~n24406;
  assign n24408 = ~controllable_hgrant3 & ~n24407;
  assign n24409 = ~n13923 & ~n24408;
  assign n24410 = ~controllable_hgrant4 & ~n24409;
  assign n24411 = ~n13922 & ~n24410;
  assign n24412 = ~controllable_hgrant5 & ~n24411;
  assign n24413 = ~n13921 & ~n24412;
  assign n24414 = ~controllable_hmaster2 & ~n24413;
  assign n24415 = ~n15294 & ~n24414;
  assign n24416 = ~controllable_hmaster1 & ~n24415;
  assign n24417 = ~n15194 & ~n24416;
  assign n24418 = ~controllable_hgrant6 & ~n24417;
  assign n24419 = ~n15964 & ~n24418;
  assign n24420 = ~controllable_hmaster0 & ~n24419;
  assign n24421 = ~n13765 & ~n24420;
  assign n24422 = ~controllable_hmaster3 & ~n24421;
  assign n24423 = ~n13672 & ~n24422;
  assign n24424 = i_hbusreq7 & ~n24423;
  assign n24425 = i_hbusreq8 & ~n24421;
  assign n24426 = i_hbusreq6 & ~n24417;
  assign n24427 = i_hbusreq5 & ~n24411;
  assign n24428 = i_hbusreq4 & ~n24409;
  assign n24429 = i_hbusreq9 & ~n24409;
  assign n24430 = i_hbusreq3 & ~n24407;
  assign n24431 = i_hbusreq1 & ~n24405;
  assign n24432 = ~i_hlock0 & ~n17757;
  assign n24433 = ~n18446 & ~n24432;
  assign n24434 = ~i_hbusreq0 & ~n24433;
  assign n24435 = ~n17815 & ~n24434;
  assign n24436 = ~i_hbusreq2 & ~n24435;
  assign n24437 = ~n17814 & ~n24436;
  assign n24438 = ~controllable_hgrant2 & ~n24437;
  assign n24439 = ~n14231 & ~n24438;
  assign n24440 = ~n7733 & ~n24439;
  assign n24441 = ~n17764 & ~n24440;
  assign n24442 = n7928 & ~n24441;
  assign n24443 = ~n8440 & ~n24442;
  assign n24444 = ~i_hbusreq1 & ~n24443;
  assign n24445 = ~n24431 & ~n24444;
  assign n24446 = ~controllable_hgrant1 & ~n24445;
  assign n24447 = ~n15107 & ~n24446;
  assign n24448 = ~i_hbusreq3 & ~n24447;
  assign n24449 = ~n24430 & ~n24448;
  assign n24450 = ~controllable_hgrant3 & ~n24449;
  assign n24451 = ~n15106 & ~n24450;
  assign n24452 = ~i_hbusreq9 & ~n24451;
  assign n24453 = ~n24429 & ~n24452;
  assign n24454 = ~i_hbusreq4 & ~n24453;
  assign n24455 = ~n24428 & ~n24454;
  assign n24456 = ~controllable_hgrant4 & ~n24455;
  assign n24457 = ~n15105 & ~n24456;
  assign n24458 = ~i_hbusreq5 & ~n24457;
  assign n24459 = ~n24427 & ~n24458;
  assign n24460 = ~controllable_hgrant5 & ~n24459;
  assign n24461 = ~n15104 & ~n24460;
  assign n24462 = ~controllable_hmaster2 & ~n24461;
  assign n24463 = ~n15820 & ~n24462;
  assign n24464 = ~controllable_hmaster1 & ~n24463;
  assign n24465 = ~n15819 & ~n24464;
  assign n24466 = ~i_hbusreq6 & ~n24465;
  assign n24467 = ~n24426 & ~n24466;
  assign n24468 = ~controllable_hgrant6 & ~n24467;
  assign n24469 = ~n15996 & ~n24468;
  assign n24470 = ~controllable_hmaster0 & ~n24469;
  assign n24471 = ~n15817 & ~n24470;
  assign n24472 = ~i_hbusreq8 & ~n24471;
  assign n24473 = ~n24425 & ~n24472;
  assign n24474 = ~controllable_hmaster3 & ~n24473;
  assign n24475 = ~n15994 & ~n24474;
  assign n24476 = ~i_hbusreq7 & ~n24475;
  assign n24477 = ~n24424 & ~n24476;
  assign n24478 = n7924 & ~n24477;
  assign n24479 = ~n24404 & ~n24478;
  assign n24480 = n8214 & ~n24479;
  assign n24481 = ~n24376 & ~n24480;
  assign n24482 = ~n8202 & ~n24481;
  assign n24483 = n8202 & ~n22210;
  assign n24484 = ~n24482 & ~n24483;
  assign n24485 = n7920 & ~n24484;
  assign n24486 = ~n24247 & ~n24485;
  assign n24487 = n7728 & ~n24486;
  assign n24488 = ~n18143 & ~n19261;
  assign n24489 = ~controllable_hmaster1 & ~n24488;
  assign n24490 = ~n19251 & ~n24489;
  assign n24491 = ~controllable_hgrant6 & ~n24490;
  assign n24492 = ~n13849 & ~n24491;
  assign n24493 = controllable_hmaster0 & ~n24492;
  assign n24494 = ~n19324 & ~n24493;
  assign n24495 = ~controllable_hmaster3 & ~n24494;
  assign n24496 = ~n20287 & ~n24495;
  assign n24497 = i_hlock7 & ~n24496;
  assign n24498 = ~n19330 & ~n24489;
  assign n24499 = ~controllable_hgrant6 & ~n24498;
  assign n24500 = ~n13951 & ~n24499;
  assign n24501 = controllable_hmaster0 & ~n24500;
  assign n24502 = ~n19324 & ~n24501;
  assign n24503 = ~controllable_hmaster3 & ~n24502;
  assign n24504 = ~n20287 & ~n24503;
  assign n24505 = ~i_hlock7 & ~n24504;
  assign n24506 = ~n24497 & ~n24505;
  assign n24507 = i_hbusreq7 & ~n24506;
  assign n24508 = i_hbusreq8 & ~n24494;
  assign n24509 = i_hbusreq6 & ~n24490;
  assign n24510 = ~n19521 & ~n21731;
  assign n24511 = ~controllable_hmaster1 & ~n24510;
  assign n24512 = ~n19499 & ~n24511;
  assign n24513 = ~i_hbusreq6 & ~n24512;
  assign n24514 = ~n24509 & ~n24513;
  assign n24515 = ~controllable_hgrant6 & ~n24514;
  assign n24516 = ~n16031 & ~n24515;
  assign n24517 = controllable_hmaster0 & ~n24516;
  assign n24518 = ~n19644 & ~n24517;
  assign n24519 = ~i_hbusreq8 & ~n24518;
  assign n24520 = ~n24508 & ~n24519;
  assign n24521 = ~controllable_hmaster3 & ~n24520;
  assign n24522 = ~n20338 & ~n24521;
  assign n24523 = i_hlock7 & ~n24522;
  assign n24524 = i_hbusreq8 & ~n24502;
  assign n24525 = i_hbusreq6 & ~n24498;
  assign n24526 = ~n19654 & ~n24511;
  assign n24527 = ~i_hbusreq6 & ~n24526;
  assign n24528 = ~n24525 & ~n24527;
  assign n24529 = ~controllable_hgrant6 & ~n24528;
  assign n24530 = ~n16068 & ~n24529;
  assign n24531 = controllable_hmaster0 & ~n24530;
  assign n24532 = ~n19644 & ~n24531;
  assign n24533 = ~i_hbusreq8 & ~n24532;
  assign n24534 = ~n24524 & ~n24533;
  assign n24535 = ~controllable_hmaster3 & ~n24534;
  assign n24536 = ~n20338 & ~n24535;
  assign n24537 = ~i_hlock7 & ~n24536;
  assign n24538 = ~n24523 & ~n24537;
  assign n24539 = ~i_hbusreq7 & ~n24538;
  assign n24540 = ~n24507 & ~n24539;
  assign n24541 = ~n7924 & ~n24540;
  assign n24542 = i_hlock1 & ~n19714;
  assign n24543 = ~i_hlock1 & ~n19732;
  assign n24544 = ~n24542 & ~n24543;
  assign n24545 = ~controllable_hgrant1 & ~n24544;
  assign n24546 = ~n13875 & ~n24545;
  assign n24547 = ~controllable_hgrant3 & ~n24546;
  assign n24548 = ~n13874 & ~n24547;
  assign n24549 = ~controllable_hgrant4 & ~n24548;
  assign n24550 = ~n13873 & ~n24549;
  assign n24551 = ~controllable_hgrant5 & ~n24550;
  assign n24552 = ~n13872 & ~n24551;
  assign n24553 = ~controllable_hmaster2 & ~n24552;
  assign n24554 = ~n19786 & ~n24553;
  assign n24555 = ~controllable_hmaster1 & ~n24554;
  assign n24556 = ~n19776 & ~n24555;
  assign n24557 = ~controllable_hgrant6 & ~n24556;
  assign n24558 = ~n13849 & ~n24557;
  assign n24559 = controllable_hmaster0 & ~n24558;
  assign n24560 = ~n19849 & ~n24559;
  assign n24561 = ~controllable_hmaster3 & ~n24560;
  assign n24562 = ~n20394 & ~n24561;
  assign n24563 = i_hlock7 & ~n24562;
  assign n24564 = ~n19855 & ~n24555;
  assign n24565 = ~controllable_hgrant6 & ~n24564;
  assign n24566 = ~n13951 & ~n24565;
  assign n24567 = controllable_hmaster0 & ~n24566;
  assign n24568 = ~n19849 & ~n24567;
  assign n24569 = ~controllable_hmaster3 & ~n24568;
  assign n24570 = ~n20394 & ~n24569;
  assign n24571 = ~i_hlock7 & ~n24570;
  assign n24572 = ~n24563 & ~n24571;
  assign n24573 = i_hbusreq7 & ~n24572;
  assign n24574 = i_hbusreq8 & ~n24560;
  assign n24575 = i_hbusreq6 & ~n24556;
  assign n24576 = i_hbusreq5 & ~n24550;
  assign n24577 = i_hbusreq4 & ~n24548;
  assign n24578 = i_hbusreq9 & ~n24548;
  assign n24579 = i_hbusreq3 & ~n24546;
  assign n24580 = i_hbusreq1 & ~n24544;
  assign n24581 = i_hlock1 & ~n19966;
  assign n24582 = ~i_hlock1 & ~n20002;
  assign n24583 = ~n24581 & ~n24582;
  assign n24584 = ~i_hbusreq1 & ~n24583;
  assign n24585 = ~n24580 & ~n24584;
  assign n24586 = ~controllable_hgrant1 & ~n24585;
  assign n24587 = ~n15032 & ~n24586;
  assign n24588 = ~i_hbusreq3 & ~n24587;
  assign n24589 = ~n24579 & ~n24588;
  assign n24590 = ~controllable_hgrant3 & ~n24589;
  assign n24591 = ~n15031 & ~n24590;
  assign n24592 = ~i_hbusreq9 & ~n24591;
  assign n24593 = ~n24578 & ~n24592;
  assign n24594 = ~i_hbusreq4 & ~n24593;
  assign n24595 = ~n24577 & ~n24594;
  assign n24596 = ~controllable_hgrant4 & ~n24595;
  assign n24597 = ~n15030 & ~n24596;
  assign n24598 = ~i_hbusreq5 & ~n24597;
  assign n24599 = ~n24576 & ~n24598;
  assign n24600 = ~controllable_hgrant5 & ~n24599;
  assign n24601 = ~n15029 & ~n24600;
  assign n24602 = ~controllable_hmaster2 & ~n24601;
  assign n24603 = ~n20114 & ~n24602;
  assign n24604 = ~controllable_hmaster1 & ~n24603;
  assign n24605 = ~n20092 & ~n24604;
  assign n24606 = ~i_hbusreq6 & ~n24605;
  assign n24607 = ~n24575 & ~n24606;
  assign n24608 = ~controllable_hgrant6 & ~n24607;
  assign n24609 = ~n16031 & ~n24608;
  assign n24610 = controllable_hmaster0 & ~n24609;
  assign n24611 = ~n20237 & ~n24610;
  assign n24612 = ~i_hbusreq8 & ~n24611;
  assign n24613 = ~n24574 & ~n24612;
  assign n24614 = ~controllable_hmaster3 & ~n24613;
  assign n24615 = ~n20447 & ~n24614;
  assign n24616 = i_hlock7 & ~n24615;
  assign n24617 = i_hbusreq8 & ~n24568;
  assign n24618 = i_hbusreq6 & ~n24564;
  assign n24619 = ~n20247 & ~n24604;
  assign n24620 = ~i_hbusreq6 & ~n24619;
  assign n24621 = ~n24618 & ~n24620;
  assign n24622 = ~controllable_hgrant6 & ~n24621;
  assign n24623 = ~n16068 & ~n24622;
  assign n24624 = controllable_hmaster0 & ~n24623;
  assign n24625 = ~n20237 & ~n24624;
  assign n24626 = ~i_hbusreq8 & ~n24625;
  assign n24627 = ~n24617 & ~n24626;
  assign n24628 = ~controllable_hmaster3 & ~n24627;
  assign n24629 = ~n20447 & ~n24628;
  assign n24630 = ~i_hlock7 & ~n24629;
  assign n24631 = ~n24616 & ~n24630;
  assign n24632 = ~i_hbusreq7 & ~n24631;
  assign n24633 = ~n24573 & ~n24632;
  assign n24634 = n7924 & ~n24633;
  assign n24635 = ~n24541 & ~n24634;
  assign n24636 = ~n8214 & ~n24635;
  assign n24637 = ~n18179 & ~n19299;
  assign n24638 = ~controllable_hmaster1 & ~n24637;
  assign n24639 = ~n19291 & ~n24638;
  assign n24640 = i_hlock6 & ~n24639;
  assign n24641 = ~n19318 & ~n24638;
  assign n24642 = ~i_hlock6 & ~n24641;
  assign n24643 = ~n24640 & ~n24642;
  assign n24644 = ~controllable_hgrant6 & ~n24643;
  assign n24645 = ~n13894 & ~n24644;
  assign n24646 = ~controllable_hmaster0 & ~n24645;
  assign n24647 = ~n19279 & ~n24646;
  assign n24648 = ~controllable_hmaster3 & ~n24647;
  assign n24649 = ~n20287 & ~n24648;
  assign n24650 = i_hlock7 & ~n24649;
  assign n24651 = ~n19334 & ~n24646;
  assign n24652 = ~controllable_hmaster3 & ~n24651;
  assign n24653 = ~n20287 & ~n24652;
  assign n24654 = ~i_hlock7 & ~n24653;
  assign n24655 = ~n24650 & ~n24654;
  assign n24656 = i_hbusreq7 & ~n24655;
  assign n24657 = ~n12640 & ~n16804;
  assign n24658 = i_hlock0 & ~n24657;
  assign n24659 = ~n16790 & ~n24658;
  assign n24660 = ~i_hbusreq0 & ~n24659;
  assign n24661 = ~n16786 & ~n24660;
  assign n24662 = ~i_hbusreq2 & ~n24661;
  assign n24663 = ~n16785 & ~n24662;
  assign n24664 = ~controllable_hgrant2 & ~n24663;
  assign n24665 = ~n12706 & ~n24664;
  assign n24666 = n7733 & ~n24665;
  assign n24667 = ~n16726 & ~n24666;
  assign n24668 = ~i_hbusreq1 & ~n24667;
  assign n24669 = ~n19347 & ~n24668;
  assign n24670 = ~controllable_hgrant1 & ~n24669;
  assign n24671 = ~n14877 & ~n24670;
  assign n24672 = ~i_hbusreq3 & ~n24671;
  assign n24673 = ~n19346 & ~n24672;
  assign n24674 = ~controllable_hgrant3 & ~n24673;
  assign n24675 = ~n14876 & ~n24674;
  assign n24676 = ~i_hbusreq9 & ~n24675;
  assign n24677 = ~n19345 & ~n24676;
  assign n24678 = ~i_hbusreq4 & ~n24677;
  assign n24679 = ~n19344 & ~n24678;
  assign n24680 = ~controllable_hgrant4 & ~n24679;
  assign n24681 = ~n14875 & ~n24680;
  assign n24682 = ~i_hbusreq5 & ~n24681;
  assign n24683 = ~n19343 & ~n24682;
  assign n24684 = ~controllable_hgrant5 & ~n24683;
  assign n24685 = ~n14874 & ~n24684;
  assign n24686 = controllable_hmaster1 & ~n24685;
  assign n24687 = controllable_hmaster2 & ~n24685;
  assign n24688 = ~n16139 & ~n16405;
  assign n24689 = i_hlock0 & ~n24688;
  assign n24690 = ~n16394 & ~n24689;
  assign n24691 = ~i_hbusreq0 & ~n24690;
  assign n24692 = ~n16391 & ~n24691;
  assign n24693 = ~i_hbusreq2 & ~n24692;
  assign n24694 = ~n16390 & ~n24693;
  assign n24695 = ~controllable_hgrant2 & n24694;
  assign n24696 = ~n12706 & ~n24695;
  assign n24697 = n7733 & ~n24696;
  assign n24698 = ~n16402 & ~n24697;
  assign n24699 = n7928 & ~n24698;
  assign n24700 = ~n16191 & ~n24699;
  assign n24701 = ~i_hbusreq1 & ~n24700;
  assign n24702 = ~n19372 & ~n24701;
  assign n24703 = ~controllable_hgrant1 & ~n24702;
  assign n24704 = ~n12681 & ~n24703;
  assign n24705 = ~i_hbusreq3 & ~n24704;
  assign n24706 = ~n19371 & ~n24705;
  assign n24707 = ~controllable_hgrant3 & ~n24706;
  assign n24708 = ~n12679 & ~n24707;
  assign n24709 = i_hlock9 & ~n24708;
  assign n24710 = ~n16216 & ~n24699;
  assign n24711 = ~i_hbusreq1 & ~n24710;
  assign n24712 = ~n19385 & ~n24711;
  assign n24713 = ~controllable_hgrant1 & ~n24712;
  assign n24714 = ~n12730 & ~n24713;
  assign n24715 = ~i_hbusreq3 & ~n24714;
  assign n24716 = ~n19384 & ~n24715;
  assign n24717 = ~controllable_hgrant3 & ~n24716;
  assign n24718 = ~n12728 & ~n24717;
  assign n24719 = ~i_hlock9 & ~n24718;
  assign n24720 = ~n24709 & ~n24719;
  assign n24721 = ~i_hbusreq9 & ~n24720;
  assign n24722 = ~n19370 & ~n24721;
  assign n24723 = ~i_hbusreq4 & ~n24722;
  assign n24724 = ~n19369 & ~n24723;
  assign n24725 = ~controllable_hgrant4 & ~n24724;
  assign n24726 = ~n12676 & ~n24725;
  assign n24727 = ~i_hbusreq5 & ~n24726;
  assign n24728 = ~n19368 & ~n24727;
  assign n24729 = ~controllable_hgrant5 & ~n24728;
  assign n24730 = ~n12674 & ~n24729;
  assign n24731 = ~controllable_hmaster2 & ~n24730;
  assign n24732 = ~n24687 & ~n24731;
  assign n24733 = ~controllable_hmaster1 & ~n24732;
  assign n24734 = ~n24686 & ~n24733;
  assign n24735 = ~i_hbusreq6 & ~n24734;
  assign n24736 = ~n19342 & ~n24735;
  assign n24737 = ~controllable_hgrant6 & ~n24736;
  assign n24738 = ~n14849 & ~n24737;
  assign n24739 = controllable_hmaster0 & ~n24738;
  assign n24740 = ~n16798 & ~n24666;
  assign n24741 = n7928 & ~n24740;
  assign n24742 = ~n8265 & ~n24741;
  assign n24743 = ~i_hbusreq1 & ~n24742;
  assign n24744 = ~n19448 & ~n24743;
  assign n24745 = ~controllable_hgrant1 & ~n24744;
  assign n24746 = ~n12681 & ~n24745;
  assign n24747 = ~i_hbusreq3 & ~n24746;
  assign n24748 = ~n19447 & ~n24747;
  assign n24749 = ~controllable_hgrant3 & ~n24748;
  assign n24750 = ~n12679 & ~n24749;
  assign n24751 = ~i_hbusreq9 & ~n24750;
  assign n24752 = ~n19446 & ~n24751;
  assign n24753 = ~i_hbusreq4 & ~n24752;
  assign n24754 = ~n19445 & ~n24753;
  assign n24755 = ~controllable_hgrant4 & ~n24754;
  assign n24756 = ~n13524 & ~n24755;
  assign n24757 = ~i_hbusreq5 & ~n24756;
  assign n24758 = ~n19444 & ~n24757;
  assign n24759 = ~controllable_hgrant5 & ~n24758;
  assign n24760 = ~n13522 & ~n24759;
  assign n24761 = ~controllable_hmaster2 & ~n24760;
  assign n24762 = ~n24687 & ~n24761;
  assign n24763 = ~controllable_hmaster1 & ~n24762;
  assign n24764 = ~n24686 & ~n24763;
  assign n24765 = ~i_hbusreq6 & ~n24764;
  assign n24766 = ~n20311 & ~n24765;
  assign n24767 = ~controllable_hgrant6 & ~n24766;
  assign n24768 = ~n14927 & ~n24767;
  assign n24769 = ~controllable_hmaster0 & ~n24768;
  assign n24770 = ~n24739 & ~n24769;
  assign n24771 = i_hlock8 & ~n24770;
  assign n24772 = ~n8297 & ~n24741;
  assign n24773 = ~i_hbusreq1 & ~n24772;
  assign n24774 = ~n19475 & ~n24773;
  assign n24775 = ~controllable_hgrant1 & ~n24774;
  assign n24776 = ~n12730 & ~n24775;
  assign n24777 = ~i_hbusreq3 & ~n24776;
  assign n24778 = ~n19504 & ~n24777;
  assign n24779 = ~controllable_hgrant3 & ~n24778;
  assign n24780 = ~n12728 & ~n24779;
  assign n24781 = ~i_hbusreq9 & ~n24780;
  assign n24782 = ~n19503 & ~n24781;
  assign n24783 = ~i_hbusreq4 & ~n24782;
  assign n24784 = ~n19502 & ~n24783;
  assign n24785 = ~controllable_hgrant4 & ~n24784;
  assign n24786 = ~n13577 & ~n24785;
  assign n24787 = ~i_hbusreq5 & ~n24786;
  assign n24788 = ~n19629 & ~n24787;
  assign n24789 = ~controllable_hgrant5 & ~n24788;
  assign n24790 = ~n13575 & ~n24789;
  assign n24791 = ~controllable_hmaster2 & ~n24790;
  assign n24792 = ~n24687 & ~n24791;
  assign n24793 = ~controllable_hmaster1 & ~n24792;
  assign n24794 = ~n24686 & ~n24793;
  assign n24795 = ~i_hbusreq6 & ~n24794;
  assign n24796 = ~n20323 & ~n24795;
  assign n24797 = ~controllable_hgrant6 & ~n24796;
  assign n24798 = ~n14960 & ~n24797;
  assign n24799 = ~controllable_hmaster0 & ~n24798;
  assign n24800 = ~n24739 & ~n24799;
  assign n24801 = ~i_hlock8 & ~n24800;
  assign n24802 = ~n24771 & ~n24801;
  assign n24803 = ~i_hbusreq8 & ~n24802;
  assign n24804 = ~n20310 & ~n24803;
  assign n24805 = controllable_hmaster3 & ~n24804;
  assign n24806 = i_hbusreq8 & ~n24647;
  assign n24807 = controllable_hmaster2 & ~n24760;
  assign n24808 = i_hlock3 & ~n24746;
  assign n24809 = ~i_hlock3 & ~n24776;
  assign n24810 = ~n24808 & ~n24809;
  assign n24811 = ~i_hbusreq3 & ~n24810;
  assign n24812 = ~n19473 & ~n24811;
  assign n24813 = ~controllable_hgrant3 & ~n24812;
  assign n24814 = ~n14999 & ~n24813;
  assign n24815 = ~i_hbusreq9 & ~n24814;
  assign n24816 = ~n19472 & ~n24815;
  assign n24817 = ~i_hbusreq4 & ~n24816;
  assign n24818 = ~n19471 & ~n24817;
  assign n24819 = ~controllable_hgrant4 & ~n24818;
  assign n24820 = ~n14998 & ~n24819;
  assign n24821 = ~i_hbusreq5 & ~n24820;
  assign n24822 = ~n19470 & ~n24821;
  assign n24823 = ~controllable_hgrant5 & ~n24822;
  assign n24824 = ~n14997 & ~n24823;
  assign n24825 = ~controllable_hmaster2 & ~n24824;
  assign n24826 = ~n24807 & ~n24825;
  assign n24827 = controllable_hmaster1 & ~n24826;
  assign n24828 = i_hlock5 & ~n24756;
  assign n24829 = ~i_hlock5 & ~n24786;
  assign n24830 = ~n24828 & ~n24829;
  assign n24831 = ~i_hbusreq5 & ~n24830;
  assign n24832 = ~n19500 & ~n24831;
  assign n24833 = ~controllable_hgrant5 & ~n24832;
  assign n24834 = ~n15020 & ~n24833;
  assign n24835 = controllable_hmaster2 & ~n24834;
  assign n24836 = i_hlock1 & ~n24742;
  assign n24837 = ~i_hlock1 & ~n24772;
  assign n24838 = ~n24836 & ~n24837;
  assign n24839 = ~i_hbusreq1 & ~n24838;
  assign n24840 = ~n19526 & ~n24839;
  assign n24841 = ~controllable_hgrant1 & ~n24840;
  assign n24842 = ~n15032 & ~n24841;
  assign n24843 = ~i_hbusreq3 & ~n24842;
  assign n24844 = ~n19525 & ~n24843;
  assign n24845 = ~controllable_hgrant3 & ~n24844;
  assign n24846 = ~n15031 & ~n24845;
  assign n24847 = ~i_hbusreq9 & ~n24846;
  assign n24848 = ~n19524 & ~n24847;
  assign n24849 = ~i_hbusreq4 & ~n24848;
  assign n24850 = ~n19523 & ~n24849;
  assign n24851 = ~controllable_hgrant4 & ~n24850;
  assign n24852 = ~n15030 & ~n24851;
  assign n24853 = ~i_hbusreq5 & ~n24852;
  assign n24854 = ~n19522 & ~n24853;
  assign n24855 = ~controllable_hgrant5 & ~n24854;
  assign n24856 = ~n15029 & ~n24855;
  assign n24857 = ~controllable_hmaster2 & ~n24856;
  assign n24858 = ~n24835 & ~n24857;
  assign n24859 = ~controllable_hmaster1 & ~n24858;
  assign n24860 = ~n24827 & ~n24859;
  assign n24861 = ~i_hbusreq6 & ~n24860;
  assign n24862 = ~n19443 & ~n24861;
  assign n24863 = ~controllable_hgrant6 & ~n24862;
  assign n24864 = ~n14995 & ~n24863;
  assign n24865 = controllable_hmaster0 & ~n24864;
  assign n24866 = i_hbusreq6 & ~n24643;
  assign n24867 = ~n9379 & ~n24741;
  assign n24868 = ~i_hbusreq1 & ~n24867;
  assign n24869 = ~n19562 & ~n24868;
  assign n24870 = ~controllable_hgrant1 & ~n24869;
  assign n24871 = ~n15067 & ~n24870;
  assign n24872 = ~i_hbusreq3 & ~n24871;
  assign n24873 = ~n19561 & ~n24872;
  assign n24874 = ~controllable_hgrant3 & ~n24873;
  assign n24875 = ~n15066 & ~n24874;
  assign n24876 = ~i_hbusreq9 & ~n24875;
  assign n24877 = ~n19560 & ~n24876;
  assign n24878 = ~i_hbusreq4 & ~n24877;
  assign n24879 = ~n19559 & ~n24878;
  assign n24880 = ~controllable_hgrant4 & ~n24879;
  assign n24881 = ~n15065 & ~n24880;
  assign n24882 = ~i_hbusreq5 & ~n24881;
  assign n24883 = ~n19558 & ~n24882;
  assign n24884 = ~controllable_hgrant5 & ~n24883;
  assign n24885 = ~n15064 & ~n24884;
  assign n24886 = ~controllable_hmaster2 & ~n24885;
  assign n24887 = ~n24807 & ~n24886;
  assign n24888 = controllable_hmaster1 & ~n24887;
  assign n24889 = i_hlock4 & ~n24752;
  assign n24890 = ~i_hlock4 & ~n24782;
  assign n24891 = ~n24889 & ~n24890;
  assign n24892 = ~i_hbusreq4 & ~n24891;
  assign n24893 = ~n19586 & ~n24892;
  assign n24894 = ~controllable_hgrant4 & ~n24893;
  assign n24895 = ~n15091 & ~n24894;
  assign n24896 = ~i_hbusreq5 & ~n24895;
  assign n24897 = ~n19585 & ~n24896;
  assign n24898 = ~controllable_hgrant5 & ~n24897;
  assign n24899 = ~n15090 & ~n24898;
  assign n24900 = controllable_hmaster2 & ~n24899;
  assign n24901 = ~n21795 & ~n24900;
  assign n24902 = ~controllable_hmaster1 & ~n24901;
  assign n24903 = ~n24888 & ~n24902;
  assign n24904 = i_hlock6 & ~n24903;
  assign n24905 = controllable_hmaster2 & ~n24790;
  assign n24906 = ~n24886 & ~n24905;
  assign n24907 = controllable_hmaster1 & ~n24906;
  assign n24908 = ~n24902 & ~n24907;
  assign n24909 = ~i_hlock6 & ~n24908;
  assign n24910 = ~n24904 & ~n24909;
  assign n24911 = ~i_hbusreq6 & ~n24910;
  assign n24912 = ~n24866 & ~n24911;
  assign n24913 = ~controllable_hgrant6 & ~n24912;
  assign n24914 = ~n15063 & ~n24913;
  assign n24915 = ~controllable_hmaster0 & ~n24914;
  assign n24916 = ~n24865 & ~n24915;
  assign n24917 = ~i_hbusreq8 & ~n24916;
  assign n24918 = ~n24806 & ~n24917;
  assign n24919 = ~controllable_hmaster3 & ~n24918;
  assign n24920 = ~n24805 & ~n24919;
  assign n24921 = i_hlock7 & ~n24920;
  assign n24922 = i_hbusreq8 & ~n24651;
  assign n24923 = ~n24825 & ~n24905;
  assign n24924 = controllable_hmaster1 & ~n24923;
  assign n24925 = ~n24859 & ~n24924;
  assign n24926 = ~i_hbusreq6 & ~n24925;
  assign n24927 = ~n19652 & ~n24926;
  assign n24928 = ~controllable_hgrant6 & ~n24927;
  assign n24929 = ~n15152 & ~n24928;
  assign n24930 = controllable_hmaster0 & ~n24929;
  assign n24931 = ~n24915 & ~n24930;
  assign n24932 = ~i_hbusreq8 & ~n24931;
  assign n24933 = ~n24922 & ~n24932;
  assign n24934 = ~controllable_hmaster3 & ~n24933;
  assign n24935 = ~n24805 & ~n24934;
  assign n24936 = ~i_hlock7 & ~n24935;
  assign n24937 = ~n24921 & ~n24936;
  assign n24938 = ~i_hbusreq7 & ~n24937;
  assign n24939 = ~n24656 & ~n24938;
  assign n24940 = ~n7924 & ~n24939;
  assign n24941 = ~n8440 & ~n19713;
  assign n24942 = ~controllable_hgrant1 & ~n24941;
  assign n24943 = ~n13924 & ~n24942;
  assign n24944 = ~controllable_hgrant3 & ~n24943;
  assign n24945 = ~n13923 & ~n24944;
  assign n24946 = ~controllable_hgrant4 & ~n24945;
  assign n24947 = ~n13922 & ~n24946;
  assign n24948 = ~controllable_hgrant5 & ~n24947;
  assign n24949 = ~n13921 & ~n24948;
  assign n24950 = ~controllable_hmaster2 & ~n24949;
  assign n24951 = ~n19824 & ~n24950;
  assign n24952 = ~controllable_hmaster1 & ~n24951;
  assign n24953 = ~n19816 & ~n24952;
  assign n24954 = i_hlock6 & ~n24953;
  assign n24955 = ~n19843 & ~n24952;
  assign n24956 = ~i_hlock6 & ~n24955;
  assign n24957 = ~n24954 & ~n24956;
  assign n24958 = ~controllable_hgrant6 & ~n24957;
  assign n24959 = ~n13894 & ~n24958;
  assign n24960 = ~controllable_hmaster0 & ~n24959;
  assign n24961 = ~n19804 & ~n24960;
  assign n24962 = ~controllable_hmaster3 & ~n24961;
  assign n24963 = ~n20394 & ~n24962;
  assign n24964 = i_hlock7 & ~n24963;
  assign n24965 = ~n19859 & ~n24960;
  assign n24966 = ~controllable_hmaster3 & ~n24965;
  assign n24967 = ~n20394 & ~n24966;
  assign n24968 = ~i_hlock7 & ~n24967;
  assign n24969 = ~n24964 & ~n24968;
  assign n24970 = i_hbusreq7 & ~n24969;
  assign n24971 = ~n7928 & ~n24667;
  assign n24972 = ~n13008 & ~n21835;
  assign n24973 = i_hlock0 & ~n24972;
  assign n24974 = ~n18792 & ~n24973;
  assign n24975 = ~i_hbusreq0 & ~n24974;
  assign n24976 = ~n17627 & ~n24975;
  assign n24977 = ~i_hbusreq2 & ~n24976;
  assign n24978 = ~n17626 & ~n24977;
  assign n24979 = ~controllable_hgrant2 & ~n24978;
  assign n24980 = ~n7814 & ~n24979;
  assign n24981 = ~n7733 & ~n24980;
  assign n24982 = ~controllable_locked & n8218;
  assign n24983 = ~n12640 & ~n24982;
  assign n24984 = i_hlock0 & ~n24983;
  assign n24985 = ~n18792 & ~n24984;
  assign n24986 = ~i_hbusreq0 & ~n24985;
  assign n24987 = ~n17627 & ~n24986;
  assign n24988 = ~i_hbusreq2 & ~n24987;
  assign n24989 = ~n17626 & ~n24988;
  assign n24990 = ~controllable_hgrant2 & ~n24989;
  assign n24991 = ~n12706 & ~n24990;
  assign n24992 = n7733 & ~n24991;
  assign n24993 = ~n24981 & ~n24992;
  assign n24994 = n7928 & ~n24993;
  assign n24995 = ~n24971 & ~n24994;
  assign n24996 = ~i_hbusreq1 & ~n24995;
  assign n24997 = ~n19872 & ~n24996;
  assign n24998 = ~controllable_hgrant1 & ~n24997;
  assign n24999 = ~n14877 & ~n24998;
  assign n25000 = ~i_hbusreq3 & ~n24999;
  assign n25001 = ~n19871 & ~n25000;
  assign n25002 = ~controllable_hgrant3 & ~n25001;
  assign n25003 = ~n14876 & ~n25002;
  assign n25004 = ~i_hbusreq9 & ~n25003;
  assign n25005 = ~n19870 & ~n25004;
  assign n25006 = ~i_hbusreq4 & ~n25005;
  assign n25007 = ~n19869 & ~n25006;
  assign n25008 = ~controllable_hgrant4 & ~n25007;
  assign n25009 = ~n14875 & ~n25008;
  assign n25010 = ~i_hbusreq5 & ~n25009;
  assign n25011 = ~n19868 & ~n25010;
  assign n25012 = ~controllable_hgrant5 & ~n25011;
  assign n25013 = ~n14874 & ~n25012;
  assign n25014 = controllable_hmaster1 & ~n25013;
  assign n25015 = controllable_hmaster2 & ~n25013;
  assign n25016 = ~n12615 & ~n16139;
  assign n25017 = i_hlock0 & ~n25016;
  assign n25018 = ~n16627 & ~n25017;
  assign n25019 = ~i_hbusreq0 & ~n25018;
  assign n25020 = ~n16624 & ~n25019;
  assign n25021 = ~i_hbusreq2 & ~n25020;
  assign n25022 = ~n16623 & ~n25021;
  assign n25023 = ~controllable_hgrant2 & n25022;
  assign n25024 = ~n12706 & ~n25023;
  assign n25025 = n7733 & ~n25024;
  assign n25026 = ~n16635 & ~n25025;
  assign n25027 = n7928 & ~n25026;
  assign n25028 = ~n16191 & ~n25027;
  assign n25029 = ~i_hbusreq1 & ~n25028;
  assign n25030 = ~n19900 & ~n25029;
  assign n25031 = ~controllable_hgrant1 & ~n25030;
  assign n25032 = ~n12681 & ~n25031;
  assign n25033 = ~i_hbusreq3 & ~n25032;
  assign n25034 = ~n19899 & ~n25033;
  assign n25035 = ~controllable_hgrant3 & ~n25034;
  assign n25036 = ~n12679 & ~n25035;
  assign n25037 = i_hlock9 & ~n25036;
  assign n25038 = ~n16216 & ~n25027;
  assign n25039 = ~i_hbusreq1 & ~n25038;
  assign n25040 = ~n19913 & ~n25039;
  assign n25041 = ~controllable_hgrant1 & ~n25040;
  assign n25042 = ~n12730 & ~n25041;
  assign n25043 = ~i_hbusreq3 & ~n25042;
  assign n25044 = ~n19912 & ~n25043;
  assign n25045 = ~controllable_hgrant3 & ~n25044;
  assign n25046 = ~n12728 & ~n25045;
  assign n25047 = ~i_hlock9 & ~n25046;
  assign n25048 = ~n25037 & ~n25047;
  assign n25049 = ~i_hbusreq9 & ~n25048;
  assign n25050 = ~n19898 & ~n25049;
  assign n25051 = ~i_hbusreq4 & ~n25050;
  assign n25052 = ~n19897 & ~n25051;
  assign n25053 = ~controllable_hgrant4 & ~n25052;
  assign n25054 = ~n12676 & ~n25053;
  assign n25055 = ~i_hbusreq5 & ~n25054;
  assign n25056 = ~n19896 & ~n25055;
  assign n25057 = ~controllable_hgrant5 & ~n25056;
  assign n25058 = ~n12674 & ~n25057;
  assign n25059 = ~controllable_hmaster2 & ~n25058;
  assign n25060 = ~n25015 & ~n25059;
  assign n25061 = ~controllable_hmaster1 & ~n25060;
  assign n25062 = ~n25014 & ~n25061;
  assign n25063 = ~i_hbusreq6 & ~n25062;
  assign n25064 = ~n19867 & ~n25063;
  assign n25065 = ~controllable_hgrant6 & ~n25064;
  assign n25066 = ~n14849 & ~n25065;
  assign n25067 = controllable_hmaster0 & ~n25066;
  assign n25068 = ~n18800 & ~n24992;
  assign n25069 = n7928 & ~n25068;
  assign n25070 = ~n8265 & ~n25069;
  assign n25071 = ~i_hbusreq1 & ~n25070;
  assign n25072 = ~n20042 & ~n25071;
  assign n25073 = ~controllable_hgrant1 & ~n25072;
  assign n25074 = ~n12681 & ~n25073;
  assign n25075 = ~i_hbusreq3 & ~n25074;
  assign n25076 = ~n20041 & ~n25075;
  assign n25077 = ~controllable_hgrant3 & ~n25076;
  assign n25078 = ~n12679 & ~n25077;
  assign n25079 = ~i_hbusreq9 & ~n25078;
  assign n25080 = ~n20040 & ~n25079;
  assign n25081 = ~i_hbusreq4 & ~n25080;
  assign n25082 = ~n20039 & ~n25081;
  assign n25083 = ~controllable_hgrant4 & ~n25082;
  assign n25084 = ~n13524 & ~n25083;
  assign n25085 = ~i_hbusreq5 & ~n25084;
  assign n25086 = ~n20038 & ~n25085;
  assign n25087 = ~controllable_hgrant5 & ~n25086;
  assign n25088 = ~n13522 & ~n25087;
  assign n25089 = ~controllable_hmaster2 & ~n25088;
  assign n25090 = ~n25015 & ~n25089;
  assign n25091 = ~controllable_hmaster1 & ~n25090;
  assign n25092 = ~n25014 & ~n25091;
  assign n25093 = ~i_hbusreq6 & ~n25092;
  assign n25094 = ~n20420 & ~n25093;
  assign n25095 = ~controllable_hgrant6 & ~n25094;
  assign n25096 = ~n14927 & ~n25095;
  assign n25097 = ~controllable_hmaster0 & ~n25096;
  assign n25098 = ~n25067 & ~n25097;
  assign n25099 = i_hlock8 & ~n25098;
  assign n25100 = ~n8297 & ~n25069;
  assign n25101 = ~i_hbusreq1 & ~n25100;
  assign n25102 = ~n20068 & ~n25101;
  assign n25103 = ~controllable_hgrant1 & ~n25102;
  assign n25104 = ~n12730 & ~n25103;
  assign n25105 = ~i_hbusreq3 & ~n25104;
  assign n25106 = ~n20097 & ~n25105;
  assign n25107 = ~controllable_hgrant3 & ~n25106;
  assign n25108 = ~n12728 & ~n25107;
  assign n25109 = ~i_hbusreq9 & ~n25108;
  assign n25110 = ~n20096 & ~n25109;
  assign n25111 = ~i_hbusreq4 & ~n25110;
  assign n25112 = ~n20095 & ~n25111;
  assign n25113 = ~controllable_hgrant4 & ~n25112;
  assign n25114 = ~n13577 & ~n25113;
  assign n25115 = ~i_hbusreq5 & ~n25114;
  assign n25116 = ~n20222 & ~n25115;
  assign n25117 = ~controllable_hgrant5 & ~n25116;
  assign n25118 = ~n13575 & ~n25117;
  assign n25119 = ~controllable_hmaster2 & ~n25118;
  assign n25120 = ~n25015 & ~n25119;
  assign n25121 = ~controllable_hmaster1 & ~n25120;
  assign n25122 = ~n25014 & ~n25121;
  assign n25123 = ~i_hbusreq6 & ~n25122;
  assign n25124 = ~n20432 & ~n25123;
  assign n25125 = ~controllable_hgrant6 & ~n25124;
  assign n25126 = ~n14960 & ~n25125;
  assign n25127 = ~controllable_hmaster0 & ~n25126;
  assign n25128 = ~n25067 & ~n25127;
  assign n25129 = ~i_hlock8 & ~n25128;
  assign n25130 = ~n25099 & ~n25129;
  assign n25131 = ~i_hbusreq8 & ~n25130;
  assign n25132 = ~n20419 & ~n25131;
  assign n25133 = controllable_hmaster3 & ~n25132;
  assign n25134 = i_hbusreq8 & ~n24961;
  assign n25135 = controllable_hmaster2 & ~n25088;
  assign n25136 = i_hlock3 & ~n25074;
  assign n25137 = ~i_hlock3 & ~n25104;
  assign n25138 = ~n25136 & ~n25137;
  assign n25139 = ~i_hbusreq3 & ~n25138;
  assign n25140 = ~n20066 & ~n25139;
  assign n25141 = ~controllable_hgrant3 & ~n25140;
  assign n25142 = ~n14999 & ~n25141;
  assign n25143 = ~i_hbusreq9 & ~n25142;
  assign n25144 = ~n20065 & ~n25143;
  assign n25145 = ~i_hbusreq4 & ~n25144;
  assign n25146 = ~n20064 & ~n25145;
  assign n25147 = ~controllable_hgrant4 & ~n25146;
  assign n25148 = ~n14998 & ~n25147;
  assign n25149 = ~i_hbusreq5 & ~n25148;
  assign n25150 = ~n20063 & ~n25149;
  assign n25151 = ~controllable_hgrant5 & ~n25150;
  assign n25152 = ~n14997 & ~n25151;
  assign n25153 = ~controllable_hmaster2 & ~n25152;
  assign n25154 = ~n25135 & ~n25153;
  assign n25155 = controllable_hmaster1 & ~n25154;
  assign n25156 = i_hlock5 & ~n25084;
  assign n25157 = ~i_hlock5 & ~n25114;
  assign n25158 = ~n25156 & ~n25157;
  assign n25159 = ~i_hbusreq5 & ~n25158;
  assign n25160 = ~n20093 & ~n25159;
  assign n25161 = ~controllable_hgrant5 & ~n25160;
  assign n25162 = ~n15020 & ~n25161;
  assign n25163 = controllable_hmaster2 & ~n25162;
  assign n25164 = i_hlock1 & ~n25070;
  assign n25165 = ~i_hlock1 & ~n25100;
  assign n25166 = ~n25164 & ~n25165;
  assign n25167 = ~i_hbusreq1 & ~n25166;
  assign n25168 = ~n20119 & ~n25167;
  assign n25169 = ~controllable_hgrant1 & ~n25168;
  assign n25170 = ~n15032 & ~n25169;
  assign n25171 = ~i_hbusreq3 & ~n25170;
  assign n25172 = ~n20118 & ~n25171;
  assign n25173 = ~controllable_hgrant3 & ~n25172;
  assign n25174 = ~n15031 & ~n25173;
  assign n25175 = ~i_hbusreq9 & ~n25174;
  assign n25176 = ~n20117 & ~n25175;
  assign n25177 = ~i_hbusreq4 & ~n25176;
  assign n25178 = ~n20116 & ~n25177;
  assign n25179 = ~controllable_hgrant4 & ~n25178;
  assign n25180 = ~n15030 & ~n25179;
  assign n25181 = ~i_hbusreq5 & ~n25180;
  assign n25182 = ~n20115 & ~n25181;
  assign n25183 = ~controllable_hgrant5 & ~n25182;
  assign n25184 = ~n15029 & ~n25183;
  assign n25185 = ~controllable_hmaster2 & ~n25184;
  assign n25186 = ~n25163 & ~n25185;
  assign n25187 = ~controllable_hmaster1 & ~n25186;
  assign n25188 = ~n25155 & ~n25187;
  assign n25189 = ~i_hbusreq6 & ~n25188;
  assign n25190 = ~n20037 & ~n25189;
  assign n25191 = ~controllable_hgrant6 & ~n25190;
  assign n25192 = ~n14995 & ~n25191;
  assign n25193 = controllable_hmaster0 & ~n25192;
  assign n25194 = i_hbusreq6 & ~n24957;
  assign n25195 = ~n9379 & ~n25069;
  assign n25196 = ~i_hbusreq1 & ~n25195;
  assign n25197 = ~n20155 & ~n25196;
  assign n25198 = ~controllable_hgrant1 & ~n25197;
  assign n25199 = ~n15067 & ~n25198;
  assign n25200 = ~i_hbusreq3 & ~n25199;
  assign n25201 = ~n20154 & ~n25200;
  assign n25202 = ~controllable_hgrant3 & ~n25201;
  assign n25203 = ~n15066 & ~n25202;
  assign n25204 = ~i_hbusreq9 & ~n25203;
  assign n25205 = ~n20153 & ~n25204;
  assign n25206 = ~i_hbusreq4 & ~n25205;
  assign n25207 = ~n20152 & ~n25206;
  assign n25208 = ~controllable_hgrant4 & ~n25207;
  assign n25209 = ~n15065 & ~n25208;
  assign n25210 = ~i_hbusreq5 & ~n25209;
  assign n25211 = ~n20151 & ~n25210;
  assign n25212 = ~controllable_hgrant5 & ~n25211;
  assign n25213 = ~n15064 & ~n25212;
  assign n25214 = ~controllable_hmaster2 & ~n25213;
  assign n25215 = ~n25135 & ~n25214;
  assign n25216 = controllable_hmaster1 & ~n25215;
  assign n25217 = i_hlock4 & ~n25080;
  assign n25218 = ~i_hlock4 & ~n25110;
  assign n25219 = ~n25217 & ~n25218;
  assign n25220 = ~i_hbusreq4 & ~n25219;
  assign n25221 = ~n20179 & ~n25220;
  assign n25222 = ~controllable_hgrant4 & ~n25221;
  assign n25223 = ~n15091 & ~n25222;
  assign n25224 = ~i_hbusreq5 & ~n25223;
  assign n25225 = ~n20178 & ~n25224;
  assign n25226 = ~controllable_hgrant5 & ~n25225;
  assign n25227 = ~n15090 & ~n25226;
  assign n25228 = controllable_hmaster2 & ~n25227;
  assign n25229 = i_hbusreq5 & ~n24947;
  assign n25230 = i_hbusreq4 & ~n24945;
  assign n25231 = i_hbusreq9 & ~n24945;
  assign n25232 = i_hbusreq3 & ~n24943;
  assign n25233 = i_hbusreq1 & ~n24941;
  assign n25234 = ~n19072 & ~n19711;
  assign n25235 = n7928 & ~n25234;
  assign n25236 = ~n8440 & ~n25235;
  assign n25237 = ~i_hbusreq1 & ~n25236;
  assign n25238 = ~n25233 & ~n25237;
  assign n25239 = ~controllable_hgrant1 & ~n25238;
  assign n25240 = ~n15107 & ~n25239;
  assign n25241 = ~i_hbusreq3 & ~n25240;
  assign n25242 = ~n25232 & ~n25241;
  assign n25243 = ~controllable_hgrant3 & ~n25242;
  assign n25244 = ~n15106 & ~n25243;
  assign n25245 = ~i_hbusreq9 & ~n25244;
  assign n25246 = ~n25231 & ~n25245;
  assign n25247 = ~i_hbusreq4 & ~n25246;
  assign n25248 = ~n25230 & ~n25247;
  assign n25249 = ~controllable_hgrant4 & ~n25248;
  assign n25250 = ~n15105 & ~n25249;
  assign n25251 = ~i_hbusreq5 & ~n25250;
  assign n25252 = ~n25229 & ~n25251;
  assign n25253 = ~controllable_hgrant5 & ~n25252;
  assign n25254 = ~n15104 & ~n25253;
  assign n25255 = ~controllable_hmaster2 & ~n25254;
  assign n25256 = ~n25228 & ~n25255;
  assign n25257 = ~controllable_hmaster1 & ~n25256;
  assign n25258 = ~n25216 & ~n25257;
  assign n25259 = i_hlock6 & ~n25258;
  assign n25260 = controllable_hmaster2 & ~n25118;
  assign n25261 = ~n25214 & ~n25260;
  assign n25262 = controllable_hmaster1 & ~n25261;
  assign n25263 = ~n25257 & ~n25262;
  assign n25264 = ~i_hlock6 & ~n25263;
  assign n25265 = ~n25259 & ~n25264;
  assign n25266 = ~i_hbusreq6 & ~n25265;
  assign n25267 = ~n25194 & ~n25266;
  assign n25268 = ~controllable_hgrant6 & ~n25267;
  assign n25269 = ~n15063 & ~n25268;
  assign n25270 = ~controllable_hmaster0 & ~n25269;
  assign n25271 = ~n25193 & ~n25270;
  assign n25272 = ~i_hbusreq8 & ~n25271;
  assign n25273 = ~n25134 & ~n25272;
  assign n25274 = ~controllable_hmaster3 & ~n25273;
  assign n25275 = ~n25133 & ~n25274;
  assign n25276 = i_hlock7 & ~n25275;
  assign n25277 = i_hbusreq8 & ~n24965;
  assign n25278 = ~n25153 & ~n25260;
  assign n25279 = controllable_hmaster1 & ~n25278;
  assign n25280 = ~n25187 & ~n25279;
  assign n25281 = ~i_hbusreq6 & ~n25280;
  assign n25282 = ~n20245 & ~n25281;
  assign n25283 = ~controllable_hgrant6 & ~n25282;
  assign n25284 = ~n15152 & ~n25283;
  assign n25285 = controllable_hmaster0 & ~n25284;
  assign n25286 = ~n25270 & ~n25285;
  assign n25287 = ~i_hbusreq8 & ~n25286;
  assign n25288 = ~n25277 & ~n25287;
  assign n25289 = ~controllable_hmaster3 & ~n25288;
  assign n25290 = ~n25133 & ~n25289;
  assign n25291 = ~i_hlock7 & ~n25290;
  assign n25292 = ~n25276 & ~n25291;
  assign n25293 = ~i_hbusreq7 & ~n25292;
  assign n25294 = ~n24970 & ~n25293;
  assign n25295 = n7924 & ~n25294;
  assign n25296 = ~n24940 & ~n25295;
  assign n25297 = n8214 & ~n25296;
  assign n25298 = ~n24636 & ~n25297;
  assign n25299 = ~n8202 & ~n25298;
  assign n25300 = ~n24483 & ~n25299;
  assign n25301 = n7920 & ~n25300;
  assign n25302 = ~n24247 & ~n25301;
  assign n25303 = ~n7728 & ~n25302;
  assign n25304 = ~n24487 & ~n25303;
  assign n25305 = n7723 & ~n25304;
  assign n25306 = ~n7723 & ~n25302;
  assign n25307 = ~n25305 & ~n25306;
  assign n25308 = n7714 & ~n25307;
  assign n25309 = n7723 & ~n25302;
  assign n25310 = ~n18632 & ~n20759;
  assign n25311 = ~controllable_hmaster1 & ~n25310;
  assign n25312 = ~n20744 & ~n25311;
  assign n25313 = ~controllable_hgrant6 & ~n25312;
  assign n25314 = ~n13849 & ~n25313;
  assign n25315 = controllable_hmaster0 & ~n25314;
  assign n25316 = ~n20848 & ~n25315;
  assign n25317 = ~controllable_hmaster3 & ~n25316;
  assign n25318 = ~n21474 & ~n25317;
  assign n25319 = i_hlock7 & ~n25318;
  assign n25320 = ~n20854 & ~n25311;
  assign n25321 = ~controllable_hgrant6 & ~n25320;
  assign n25322 = ~n13951 & ~n25321;
  assign n25323 = controllable_hmaster0 & ~n25322;
  assign n25324 = ~n20848 & ~n25323;
  assign n25325 = ~controllable_hmaster3 & ~n25324;
  assign n25326 = ~n21474 & ~n25325;
  assign n25327 = ~i_hlock7 & ~n25326;
  assign n25328 = ~n25319 & ~n25327;
  assign n25329 = i_hbusreq7 & ~n25328;
  assign n25330 = i_hbusreq8 & ~n25316;
  assign n25331 = i_hbusreq6 & ~n25312;
  assign n25332 = i_hlock1 & ~n21022;
  assign n25333 = ~i_hlock1 & ~n21073;
  assign n25334 = ~n25332 & ~n25333;
  assign n25335 = ~i_hbusreq1 & ~n25334;
  assign n25336 = ~n18954 & ~n25335;
  assign n25337 = ~controllable_hgrant1 & ~n25336;
  assign n25338 = ~n15032 & ~n25337;
  assign n25339 = ~i_hbusreq3 & ~n25338;
  assign n25340 = ~n18953 & ~n25339;
  assign n25341 = ~controllable_hgrant3 & ~n25340;
  assign n25342 = ~n15031 & ~n25341;
  assign n25343 = i_hlock9 & ~n25342;
  assign n25344 = i_hlock1 & ~n21040;
  assign n25345 = ~i_hlock1 & ~n21083;
  assign n25346 = ~n25344 & ~n25345;
  assign n25347 = ~i_hbusreq1 & ~n25346;
  assign n25348 = ~n18968 & ~n25347;
  assign n25349 = ~controllable_hgrant1 & ~n25348;
  assign n25350 = ~n15032 & ~n25349;
  assign n25351 = ~i_hbusreq3 & ~n25350;
  assign n25352 = ~n18967 & ~n25351;
  assign n25353 = ~controllable_hgrant3 & ~n25352;
  assign n25354 = ~n15031 & ~n25353;
  assign n25355 = ~i_hlock9 & ~n25354;
  assign n25356 = ~n25343 & ~n25355;
  assign n25357 = ~i_hbusreq9 & ~n25356;
  assign n25358 = ~n18952 & ~n25357;
  assign n25359 = ~i_hbusreq4 & ~n25358;
  assign n25360 = ~n18951 & ~n25359;
  assign n25361 = ~controllable_hgrant4 & ~n25360;
  assign n25362 = ~n15030 & ~n25361;
  assign n25363 = ~i_hbusreq5 & ~n25362;
  assign n25364 = ~n18950 & ~n25363;
  assign n25365 = ~controllable_hgrant5 & ~n25364;
  assign n25366 = ~n15029 & ~n25365;
  assign n25367 = ~controllable_hmaster2 & ~n25366;
  assign n25368 = ~n21236 & ~n25367;
  assign n25369 = ~controllable_hmaster1 & ~n25368;
  assign n25370 = ~n21206 & ~n25369;
  assign n25371 = ~i_hbusreq6 & ~n25370;
  assign n25372 = ~n25331 & ~n25371;
  assign n25373 = ~controllable_hgrant6 & ~n25372;
  assign n25374 = ~n16031 & ~n25373;
  assign n25375 = controllable_hmaster0 & ~n25374;
  assign n25376 = ~n21424 & ~n25375;
  assign n25377 = ~i_hbusreq8 & ~n25376;
  assign n25378 = ~n25330 & ~n25377;
  assign n25379 = ~controllable_hmaster3 & ~n25378;
  assign n25380 = ~n21525 & ~n25379;
  assign n25381 = i_hlock7 & ~n25380;
  assign n25382 = i_hbusreq8 & ~n25324;
  assign n25383 = i_hbusreq6 & ~n25320;
  assign n25384 = ~n21434 & ~n25369;
  assign n25385 = ~i_hbusreq6 & ~n25384;
  assign n25386 = ~n25383 & ~n25385;
  assign n25387 = ~controllable_hgrant6 & ~n25386;
  assign n25388 = ~n16068 & ~n25387;
  assign n25389 = controllable_hmaster0 & ~n25388;
  assign n25390 = ~n21424 & ~n25389;
  assign n25391 = ~i_hbusreq8 & ~n25390;
  assign n25392 = ~n25382 & ~n25391;
  assign n25393 = ~controllable_hmaster3 & ~n25392;
  assign n25394 = ~n21525 & ~n25393;
  assign n25395 = ~i_hlock7 & ~n25394;
  assign n25396 = ~n25381 & ~n25395;
  assign n25397 = ~i_hbusreq7 & ~n25396;
  assign n25398 = ~n25329 & ~n25397;
  assign n25399 = n7924 & ~n25398;
  assign n25400 = ~n24541 & ~n25399;
  assign n25401 = ~n8214 & ~n25400;
  assign n25402 = ~n18684 & ~n20815;
  assign n25403 = ~controllable_hmaster1 & ~n25402;
  assign n25404 = ~n20807 & ~n25403;
  assign n25405 = i_hlock6 & ~n25404;
  assign n25406 = ~n20842 & ~n25403;
  assign n25407 = ~i_hlock6 & ~n25406;
  assign n25408 = ~n25405 & ~n25407;
  assign n25409 = ~controllable_hgrant6 & ~n25408;
  assign n25410 = ~n13894 & ~n25409;
  assign n25411 = ~controllable_hmaster0 & ~n25410;
  assign n25412 = ~n20787 & ~n25411;
  assign n25413 = ~controllable_hmaster3 & ~n25412;
  assign n25414 = ~n21474 & ~n25413;
  assign n25415 = i_hlock7 & ~n25414;
  assign n25416 = ~n20858 & ~n25411;
  assign n25417 = ~controllable_hmaster3 & ~n25416;
  assign n25418 = ~n21474 & ~n25417;
  assign n25419 = ~i_hlock7 & ~n25418;
  assign n25420 = ~n25415 & ~n25419;
  assign n25421 = i_hbusreq7 & ~n25420;
  assign n25422 = ~n17553 & ~n20656;
  assign n25423 = controllable_locked & ~n25422;
  assign n25424 = ~n12615 & ~n25423;
  assign n25425 = i_hlock0 & ~n25424;
  assign n25426 = ~n20876 & ~n25425;
  assign n25427 = ~i_hbusreq0 & ~n25426;
  assign n25428 = ~n20873 & ~n25427;
  assign n25429 = ~i_hbusreq2 & ~n25428;
  assign n25430 = ~n20872 & ~n25429;
  assign n25431 = ~controllable_hgrant2 & n25430;
  assign n25432 = ~n12706 & ~n25431;
  assign n25433 = n7733 & ~n25432;
  assign n25434 = ~n24981 & ~n25433;
  assign n25435 = n7928 & ~n25434;
  assign n25436 = ~n24971 & ~n25435;
  assign n25437 = ~i_hbusreq1 & ~n25436;
  assign n25438 = ~n20871 & ~n25437;
  assign n25439 = ~controllable_hgrant1 & ~n25438;
  assign n25440 = ~n14877 & ~n25439;
  assign n25441 = ~i_hbusreq3 & ~n25440;
  assign n25442 = ~n20870 & ~n25441;
  assign n25443 = ~controllable_hgrant3 & ~n25442;
  assign n25444 = ~n14876 & ~n25443;
  assign n25445 = i_hlock9 & ~n25444;
  assign n25446 = ~n20900 & ~n25427;
  assign n25447 = ~i_hbusreq2 & ~n25446;
  assign n25448 = ~n20899 & ~n25447;
  assign n25449 = ~controllable_hgrant2 & n25448;
  assign n25450 = ~n12706 & ~n25449;
  assign n25451 = n7733 & ~n25450;
  assign n25452 = ~n24981 & ~n25451;
  assign n25453 = n7928 & ~n25452;
  assign n25454 = ~n24971 & ~n25453;
  assign n25455 = ~i_hbusreq1 & ~n25454;
  assign n25456 = ~n20898 & ~n25455;
  assign n25457 = ~controllable_hgrant1 & ~n25456;
  assign n25458 = ~n14877 & ~n25457;
  assign n25459 = ~i_hbusreq3 & ~n25458;
  assign n25460 = ~n20897 & ~n25459;
  assign n25461 = ~controllable_hgrant3 & ~n25460;
  assign n25462 = ~n14876 & ~n25461;
  assign n25463 = ~i_hlock9 & ~n25462;
  assign n25464 = ~n25445 & ~n25463;
  assign n25465 = ~i_hbusreq9 & ~n25464;
  assign n25466 = ~n20869 & ~n25465;
  assign n25467 = ~i_hbusreq4 & ~n25466;
  assign n25468 = ~n20868 & ~n25467;
  assign n25469 = ~controllable_hgrant4 & ~n25468;
  assign n25470 = ~n14875 & ~n25469;
  assign n25471 = ~i_hbusreq5 & ~n25470;
  assign n25472 = ~n20867 & ~n25471;
  assign n25473 = ~controllable_hgrant5 & ~n25472;
  assign n25474 = ~n14874 & ~n25473;
  assign n25475 = controllable_hmaster1 & ~n25474;
  assign n25476 = controllable_hmaster2 & ~n25474;
  assign n25477 = ~n7858 & ~n20656;
  assign n25478 = controllable_locked & ~n25477;
  assign n25479 = ~n12615 & ~n25478;
  assign n25480 = i_hlock0 & ~n25479;
  assign n25481 = ~n20944 & ~n25480;
  assign n25482 = ~i_hbusreq0 & ~n25481;
  assign n25483 = ~n20938 & ~n25482;
  assign n25484 = ~i_hbusreq2 & ~n25483;
  assign n25485 = ~n20937 & ~n25484;
  assign n25486 = ~controllable_hgrant2 & n25485;
  assign n25487 = ~n12706 & ~n25486;
  assign n25488 = n7733 & ~n25487;
  assign n25489 = ~n16635 & ~n25488;
  assign n25490 = n7928 & ~n25489;
  assign n25491 = ~n16191 & ~n25490;
  assign n25492 = ~i_hbusreq1 & ~n25491;
  assign n25493 = ~n20936 & ~n25492;
  assign n25494 = ~controllable_hgrant1 & ~n25493;
  assign n25495 = ~n12681 & ~n25494;
  assign n25496 = ~i_hbusreq3 & ~n25495;
  assign n25497 = ~n20935 & ~n25496;
  assign n25498 = ~controllable_hgrant3 & ~n25497;
  assign n25499 = ~n12679 & ~n25498;
  assign n25500 = i_hlock9 & ~n25499;
  assign n25501 = ~n20968 & ~n25482;
  assign n25502 = ~i_hbusreq2 & ~n25501;
  assign n25503 = ~n20967 & ~n25502;
  assign n25504 = ~controllable_hgrant2 & n25503;
  assign n25505 = ~n12706 & ~n25504;
  assign n25506 = n7733 & ~n25505;
  assign n25507 = ~n16635 & ~n25506;
  assign n25508 = n7928 & ~n25507;
  assign n25509 = ~n16216 & ~n25508;
  assign n25510 = ~i_hbusreq1 & ~n25509;
  assign n25511 = ~n20966 & ~n25510;
  assign n25512 = ~controllable_hgrant1 & ~n25511;
  assign n25513 = ~n12730 & ~n25512;
  assign n25514 = ~i_hbusreq3 & ~n25513;
  assign n25515 = ~n20965 & ~n25514;
  assign n25516 = ~controllable_hgrant3 & ~n25515;
  assign n25517 = ~n12728 & ~n25516;
  assign n25518 = ~i_hlock9 & ~n25517;
  assign n25519 = ~n25500 & ~n25518;
  assign n25520 = ~i_hbusreq9 & ~n25519;
  assign n25521 = ~n20934 & ~n25520;
  assign n25522 = ~i_hbusreq4 & ~n25521;
  assign n25523 = ~n20933 & ~n25522;
  assign n25524 = ~controllable_hgrant4 & ~n25523;
  assign n25525 = ~n12676 & ~n25524;
  assign n25526 = ~i_hbusreq5 & ~n25525;
  assign n25527 = ~n20932 & ~n25526;
  assign n25528 = ~controllable_hgrant5 & ~n25527;
  assign n25529 = ~n12674 & ~n25528;
  assign n25530 = ~controllable_hmaster2 & ~n25529;
  assign n25531 = ~n25476 & ~n25530;
  assign n25532 = ~controllable_hmaster1 & ~n25531;
  assign n25533 = ~n25475 & ~n25532;
  assign n25534 = ~i_hbusreq6 & ~n25533;
  assign n25535 = ~n20866 & ~n25534;
  assign n25536 = ~controllable_hgrant6 & ~n25535;
  assign n25537 = ~n14849 & ~n25536;
  assign n25538 = controllable_hmaster0 & ~n25537;
  assign n25539 = ~n18800 & ~n25433;
  assign n25540 = n7928 & ~n25539;
  assign n25541 = ~n8265 & ~n25540;
  assign n25542 = ~i_hbusreq1 & ~n25541;
  assign n25543 = ~n21125 & ~n25542;
  assign n25544 = ~controllable_hgrant1 & ~n25543;
  assign n25545 = ~n12681 & ~n25544;
  assign n25546 = ~i_hbusreq3 & ~n25545;
  assign n25547 = ~n21124 & ~n25546;
  assign n25548 = ~controllable_hgrant3 & ~n25547;
  assign n25549 = ~n12679 & ~n25548;
  assign n25550 = i_hlock9 & ~n25549;
  assign n25551 = ~n18800 & ~n25451;
  assign n25552 = n7928 & ~n25551;
  assign n25553 = ~n8265 & ~n25552;
  assign n25554 = ~i_hbusreq1 & ~n25553;
  assign n25555 = ~n21137 & ~n25554;
  assign n25556 = ~controllable_hgrant1 & ~n25555;
  assign n25557 = ~n12681 & ~n25556;
  assign n25558 = ~i_hbusreq3 & ~n25557;
  assign n25559 = ~n21136 & ~n25558;
  assign n25560 = ~controllable_hgrant3 & ~n25559;
  assign n25561 = ~n12679 & ~n25560;
  assign n25562 = ~i_hlock9 & ~n25561;
  assign n25563 = ~n25550 & ~n25562;
  assign n25564 = ~i_hbusreq9 & ~n25563;
  assign n25565 = ~n21123 & ~n25564;
  assign n25566 = ~i_hbusreq4 & ~n25565;
  assign n25567 = ~n21122 & ~n25566;
  assign n25568 = ~controllable_hgrant4 & ~n25567;
  assign n25569 = ~n13524 & ~n25568;
  assign n25570 = ~i_hbusreq5 & ~n25569;
  assign n25571 = ~n21121 & ~n25570;
  assign n25572 = ~controllable_hgrant5 & ~n25571;
  assign n25573 = ~n13522 & ~n25572;
  assign n25574 = ~controllable_hmaster2 & ~n25573;
  assign n25575 = ~n25476 & ~n25574;
  assign n25576 = ~controllable_hmaster1 & ~n25575;
  assign n25577 = ~n25475 & ~n25576;
  assign n25578 = ~i_hbusreq6 & ~n25577;
  assign n25579 = ~n21498 & ~n25578;
  assign n25580 = ~controllable_hgrant6 & ~n25579;
  assign n25581 = ~n14927 & ~n25580;
  assign n25582 = ~controllable_hmaster0 & ~n25581;
  assign n25583 = ~n25538 & ~n25582;
  assign n25584 = i_hlock8 & ~n25583;
  assign n25585 = ~n8297 & ~n25540;
  assign n25586 = ~i_hbusreq1 & ~n25585;
  assign n25587 = ~n21165 & ~n25586;
  assign n25588 = ~controllable_hgrant1 & ~n25587;
  assign n25589 = ~n12730 & ~n25588;
  assign n25590 = ~i_hbusreq3 & ~n25589;
  assign n25591 = ~n21211 & ~n25590;
  assign n25592 = ~controllable_hgrant3 & ~n25591;
  assign n25593 = ~n12728 & ~n25592;
  assign n25594 = i_hlock9 & ~n25593;
  assign n25595 = ~n8297 & ~n25552;
  assign n25596 = ~i_hbusreq1 & ~n25595;
  assign n25597 = ~n21180 & ~n25596;
  assign n25598 = ~controllable_hgrant1 & ~n25597;
  assign n25599 = ~n12730 & ~n25598;
  assign n25600 = ~i_hbusreq3 & ~n25599;
  assign n25601 = ~n21217 & ~n25600;
  assign n25602 = ~controllable_hgrant3 & ~n25601;
  assign n25603 = ~n12728 & ~n25602;
  assign n25604 = ~i_hlock9 & ~n25603;
  assign n25605 = ~n25594 & ~n25604;
  assign n25606 = ~i_hbusreq9 & ~n25605;
  assign n25607 = ~n21210 & ~n25606;
  assign n25608 = ~i_hbusreq4 & ~n25607;
  assign n25609 = ~n21209 & ~n25608;
  assign n25610 = ~controllable_hgrant4 & ~n25609;
  assign n25611 = ~n13577 & ~n25610;
  assign n25612 = ~i_hbusreq5 & ~n25611;
  assign n25613 = ~n21409 & ~n25612;
  assign n25614 = ~controllable_hgrant5 & ~n25613;
  assign n25615 = ~n13575 & ~n25614;
  assign n25616 = ~controllable_hmaster2 & ~n25615;
  assign n25617 = ~n25476 & ~n25616;
  assign n25618 = ~controllable_hmaster1 & ~n25617;
  assign n25619 = ~n25475 & ~n25618;
  assign n25620 = ~i_hbusreq6 & ~n25619;
  assign n25621 = ~n21510 & ~n25620;
  assign n25622 = ~controllable_hgrant6 & ~n25621;
  assign n25623 = ~n14960 & ~n25622;
  assign n25624 = ~controllable_hmaster0 & ~n25623;
  assign n25625 = ~n25538 & ~n25624;
  assign n25626 = ~i_hlock8 & ~n25625;
  assign n25627 = ~n25584 & ~n25626;
  assign n25628 = ~i_hbusreq8 & ~n25627;
  assign n25629 = ~n21497 & ~n25628;
  assign n25630 = controllable_hmaster3 & ~n25629;
  assign n25631 = i_hbusreq8 & ~n25412;
  assign n25632 = controllable_hmaster2 & ~n25573;
  assign n25633 = i_hlock3 & ~n25545;
  assign n25634 = ~i_hlock3 & ~n25589;
  assign n25635 = ~n25633 & ~n25634;
  assign n25636 = ~i_hbusreq3 & ~n25635;
  assign n25637 = ~n21163 & ~n25636;
  assign n25638 = ~controllable_hgrant3 & ~n25637;
  assign n25639 = ~n14999 & ~n25638;
  assign n25640 = i_hlock9 & ~n25639;
  assign n25641 = i_hlock3 & ~n25557;
  assign n25642 = ~i_hlock3 & ~n25599;
  assign n25643 = ~n25641 & ~n25642;
  assign n25644 = ~i_hbusreq3 & ~n25643;
  assign n25645 = ~n21178 & ~n25644;
  assign n25646 = ~controllable_hgrant3 & ~n25645;
  assign n25647 = ~n14999 & ~n25646;
  assign n25648 = ~i_hlock9 & ~n25647;
  assign n25649 = ~n25640 & ~n25648;
  assign n25650 = ~i_hbusreq9 & ~n25649;
  assign n25651 = ~n21162 & ~n25650;
  assign n25652 = ~i_hbusreq4 & ~n25651;
  assign n25653 = ~n21161 & ~n25652;
  assign n25654 = ~controllable_hgrant4 & ~n25653;
  assign n25655 = ~n14998 & ~n25654;
  assign n25656 = ~i_hbusreq5 & ~n25655;
  assign n25657 = ~n21160 & ~n25656;
  assign n25658 = ~controllable_hgrant5 & ~n25657;
  assign n25659 = ~n14997 & ~n25658;
  assign n25660 = ~controllable_hmaster2 & ~n25659;
  assign n25661 = ~n25632 & ~n25660;
  assign n25662 = controllable_hmaster1 & ~n25661;
  assign n25663 = i_hlock5 & ~n25569;
  assign n25664 = ~i_hlock5 & ~n25611;
  assign n25665 = ~n25663 & ~n25664;
  assign n25666 = ~i_hbusreq5 & ~n25665;
  assign n25667 = ~n21207 & ~n25666;
  assign n25668 = ~controllable_hgrant5 & ~n25667;
  assign n25669 = ~n15020 & ~n25668;
  assign n25670 = controllable_hmaster2 & ~n25669;
  assign n25671 = i_hlock1 & ~n25541;
  assign n25672 = ~i_hlock1 & ~n25585;
  assign n25673 = ~n25671 & ~n25672;
  assign n25674 = ~i_hbusreq1 & ~n25673;
  assign n25675 = ~n21241 & ~n25674;
  assign n25676 = ~controllable_hgrant1 & ~n25675;
  assign n25677 = ~n15032 & ~n25676;
  assign n25678 = ~i_hbusreq3 & ~n25677;
  assign n25679 = ~n21240 & ~n25678;
  assign n25680 = ~controllable_hgrant3 & ~n25679;
  assign n25681 = ~n15031 & ~n25680;
  assign n25682 = i_hlock9 & ~n25681;
  assign n25683 = i_hlock1 & ~n25553;
  assign n25684 = ~i_hlock1 & ~n25595;
  assign n25685 = ~n25683 & ~n25684;
  assign n25686 = ~i_hbusreq1 & ~n25685;
  assign n25687 = ~n21255 & ~n25686;
  assign n25688 = ~controllable_hgrant1 & ~n25687;
  assign n25689 = ~n15032 & ~n25688;
  assign n25690 = ~i_hbusreq3 & ~n25689;
  assign n25691 = ~n21254 & ~n25690;
  assign n25692 = ~controllable_hgrant3 & ~n25691;
  assign n25693 = ~n15031 & ~n25692;
  assign n25694 = ~i_hlock9 & ~n25693;
  assign n25695 = ~n25682 & ~n25694;
  assign n25696 = ~i_hbusreq9 & ~n25695;
  assign n25697 = ~n21239 & ~n25696;
  assign n25698 = ~i_hbusreq4 & ~n25697;
  assign n25699 = ~n21238 & ~n25698;
  assign n25700 = ~controllable_hgrant4 & ~n25699;
  assign n25701 = ~n15030 & ~n25700;
  assign n25702 = ~i_hbusreq5 & ~n25701;
  assign n25703 = ~n21237 & ~n25702;
  assign n25704 = ~controllable_hgrant5 & ~n25703;
  assign n25705 = ~n15029 & ~n25704;
  assign n25706 = ~controllable_hmaster2 & ~n25705;
  assign n25707 = ~n25670 & ~n25706;
  assign n25708 = ~controllable_hmaster1 & ~n25707;
  assign n25709 = ~n25662 & ~n25708;
  assign n25710 = ~i_hbusreq6 & ~n25709;
  assign n25711 = ~n21120 & ~n25710;
  assign n25712 = ~controllable_hgrant6 & ~n25711;
  assign n25713 = ~n14995 & ~n25712;
  assign n25714 = controllable_hmaster0 & ~n25713;
  assign n25715 = i_hbusreq6 & ~n25408;
  assign n25716 = ~n9379 & ~n25540;
  assign n25717 = ~i_hbusreq1 & ~n25716;
  assign n25718 = ~n21293 & ~n25717;
  assign n25719 = ~controllable_hgrant1 & ~n25718;
  assign n25720 = ~n15067 & ~n25719;
  assign n25721 = ~i_hbusreq3 & ~n25720;
  assign n25722 = ~n21292 & ~n25721;
  assign n25723 = ~controllable_hgrant3 & ~n25722;
  assign n25724 = ~n15066 & ~n25723;
  assign n25725 = i_hlock9 & ~n25724;
  assign n25726 = ~n9379 & ~n25552;
  assign n25727 = ~i_hbusreq1 & ~n25726;
  assign n25728 = ~n21305 & ~n25727;
  assign n25729 = ~controllable_hgrant1 & ~n25728;
  assign n25730 = ~n15067 & ~n25729;
  assign n25731 = ~i_hbusreq3 & ~n25730;
  assign n25732 = ~n21304 & ~n25731;
  assign n25733 = ~controllable_hgrant3 & ~n25732;
  assign n25734 = ~n15066 & ~n25733;
  assign n25735 = ~i_hlock9 & ~n25734;
  assign n25736 = ~n25725 & ~n25735;
  assign n25737 = ~i_hbusreq9 & ~n25736;
  assign n25738 = ~n21291 & ~n25737;
  assign n25739 = ~i_hbusreq4 & ~n25738;
  assign n25740 = ~n21290 & ~n25739;
  assign n25741 = ~controllable_hgrant4 & ~n25740;
  assign n25742 = ~n15065 & ~n25741;
  assign n25743 = ~i_hbusreq5 & ~n25742;
  assign n25744 = ~n21289 & ~n25743;
  assign n25745 = ~controllable_hgrant5 & ~n25744;
  assign n25746 = ~n15064 & ~n25745;
  assign n25747 = ~controllable_hmaster2 & ~n25746;
  assign n25748 = ~n25632 & ~n25747;
  assign n25749 = controllable_hmaster1 & ~n25748;
  assign n25750 = i_hlock4 & ~n25565;
  assign n25751 = ~i_hlock4 & ~n25607;
  assign n25752 = ~n25750 & ~n25751;
  assign n25753 = ~i_hbusreq4 & ~n25752;
  assign n25754 = ~n21331 & ~n25753;
  assign n25755 = ~controllable_hgrant4 & ~n25754;
  assign n25756 = ~n15091 & ~n25755;
  assign n25757 = ~i_hbusreq5 & ~n25756;
  assign n25758 = ~n21330 & ~n25757;
  assign n25759 = ~controllable_hgrant5 & ~n25758;
  assign n25760 = ~n15090 & ~n25759;
  assign n25761 = controllable_hmaster2 & ~n25760;
  assign n25762 = ~n22170 & ~n25761;
  assign n25763 = ~controllable_hmaster1 & ~n25762;
  assign n25764 = ~n25749 & ~n25763;
  assign n25765 = i_hlock6 & ~n25764;
  assign n25766 = controllable_hmaster2 & ~n25615;
  assign n25767 = ~n25747 & ~n25766;
  assign n25768 = controllable_hmaster1 & ~n25767;
  assign n25769 = ~n25763 & ~n25768;
  assign n25770 = ~i_hlock6 & ~n25769;
  assign n25771 = ~n25765 & ~n25770;
  assign n25772 = ~i_hbusreq6 & ~n25771;
  assign n25773 = ~n25715 & ~n25772;
  assign n25774 = ~controllable_hgrant6 & ~n25773;
  assign n25775 = ~n15063 & ~n25774;
  assign n25776 = ~controllable_hmaster0 & ~n25775;
  assign n25777 = ~n25714 & ~n25776;
  assign n25778 = ~i_hbusreq8 & ~n25777;
  assign n25779 = ~n25631 & ~n25778;
  assign n25780 = ~controllable_hmaster3 & ~n25779;
  assign n25781 = ~n25630 & ~n25780;
  assign n25782 = i_hlock7 & ~n25781;
  assign n25783 = i_hbusreq8 & ~n25416;
  assign n25784 = ~n25660 & ~n25766;
  assign n25785 = controllable_hmaster1 & ~n25784;
  assign n25786 = ~n25708 & ~n25785;
  assign n25787 = ~i_hbusreq6 & ~n25786;
  assign n25788 = ~n21432 & ~n25787;
  assign n25789 = ~controllable_hgrant6 & ~n25788;
  assign n25790 = ~n15152 & ~n25789;
  assign n25791 = controllable_hmaster0 & ~n25790;
  assign n25792 = ~n25776 & ~n25791;
  assign n25793 = ~i_hbusreq8 & ~n25792;
  assign n25794 = ~n25783 & ~n25793;
  assign n25795 = ~controllable_hmaster3 & ~n25794;
  assign n25796 = ~n25630 & ~n25795;
  assign n25797 = ~i_hlock7 & ~n25796;
  assign n25798 = ~n25782 & ~n25797;
  assign n25799 = ~i_hbusreq7 & ~n25798;
  assign n25800 = ~n25421 & ~n25799;
  assign n25801 = n7924 & ~n25800;
  assign n25802 = ~n24940 & ~n25801;
  assign n25803 = n8214 & ~n25802;
  assign n25804 = ~n25401 & ~n25803;
  assign n25805 = ~n8202 & ~n25804;
  assign n25806 = ~n24483 & ~n25805;
  assign n25807 = n7920 & ~n25806;
  assign n25808 = ~n16336 & ~n25807;
  assign n25809 = n7728 & ~n25808;
  assign n25810 = ~n22213 & ~n25809;
  assign n25811 = ~n7723 & ~n25810;
  assign n25812 = ~n25309 & ~n25811;
  assign n25813 = ~n7714 & ~n25812;
  assign n25814 = ~n25308 & ~n25813;
  assign n25815 = ~n7705 & ~n25814;
  assign n25816 = ~n24279 & ~n25815;
  assign n25817 = n7808 & ~n25816;
  assign n25818 = ~n23755 & ~n25817;
  assign n25819 = n8195 & ~n25818;
  assign n25820 = ~n23629 & ~n25819;
  assign n25821 = n8193 & ~n25820;
  assign n25822 = ~n22225 & ~n25821;
  assign n25823 = ~n8191 & ~n25822;
  assign n25824 = ~n16114 & ~n25823;
  assign n25825 = n8188 & ~n25824;
  assign n25826 = ~n11402 & ~n12974;
  assign n25827 = n7728 & ~n25826;
  assign n25828 = ~n11405 & ~n13113;
  assign n25829 = ~n7728 & ~n25828;
  assign n25830 = ~n25827 & ~n25829;
  assign n25831 = ~n7723 & ~n25830;
  assign n25832 = ~n7723 & ~n25831;
  assign n25833 = ~n7714 & ~n25832;
  assign n25834 = ~n7714 & ~n25833;
  assign n25835 = n7705 & ~n25834;
  assign n25836 = ~n11405 & ~n13802;
  assign n25837 = n7728 & ~n25836;
  assign n25838 = ~n11405 & ~n14838;
  assign n25839 = ~n7728 & ~n25838;
  assign n25840 = ~n25837 & ~n25839;
  assign n25841 = n7723 & ~n25840;
  assign n25842 = ~n7723 & ~n25838;
  assign n25843 = ~n25841 & ~n25842;
  assign n25844 = n7714 & ~n25843;
  assign n25845 = n7723 & ~n25838;
  assign n25846 = ~n11391 & ~n14838;
  assign n25847 = n7728 & ~n25846;
  assign n25848 = ~n11391 & ~n15172;
  assign n25849 = ~n7728 & ~n25848;
  assign n25850 = ~n25847 & ~n25849;
  assign n25851 = ~n7723 & ~n25850;
  assign n25852 = ~n25845 & ~n25851;
  assign n25853 = ~n7714 & ~n25852;
  assign n25854 = ~n25844 & ~n25853;
  assign n25855 = ~n7705 & ~n25854;
  assign n25856 = ~n25835 & ~n25855;
  assign n25857 = n7808 & ~n25856;
  assign n25858 = ~n11401 & ~n25857;
  assign n25859 = n8195 & ~n25858;
  assign n25860 = ~n8196 & ~n25859;
  assign n25861 = ~n8193 & ~n25860;
  assign n25862 = ~n11391 & ~n15638;
  assign n25863 = n7728 & ~n25862;
  assign n25864 = ~n25849 & ~n25863;
  assign n25865 = ~n7723 & ~n25864;
  assign n25866 = ~n15646 & ~n25865;
  assign n25867 = ~n7714 & ~n25866;
  assign n25868 = ~n15645 & ~n25867;
  assign n25869 = ~n7705 & ~n25868;
  assign n25870 = ~n10052 & ~n25869;
  assign n25871 = n7808 & ~n25870;
  assign n25872 = ~n11447 & ~n25871;
  assign n25873 = ~n8195 & ~n25872;
  assign n25874 = ~n11536 & ~n15866;
  assign n25875 = n7728 & ~n25874;
  assign n25876 = ~n11539 & ~n15875;
  assign n25877 = ~n7728 & ~n25876;
  assign n25878 = ~n25875 & ~n25877;
  assign n25879 = ~n7723 & ~n25878;
  assign n25880 = ~n7723 & ~n25879;
  assign n25881 = ~n7714 & ~n25880;
  assign n25882 = ~n7714 & ~n25881;
  assign n25883 = n7705 & ~n25882;
  assign n25884 = ~n11539 & ~n16020;
  assign n25885 = n7728 & ~n25884;
  assign n25886 = ~n11539 & ~n16090;
  assign n25887 = ~n7728 & ~n25886;
  assign n25888 = ~n25885 & ~n25887;
  assign n25889 = n7723 & ~n25888;
  assign n25890 = ~n7723 & ~n25886;
  assign n25891 = ~n25889 & ~n25890;
  assign n25892 = n7714 & ~n25891;
  assign n25893 = n7723 & ~n25886;
  assign n25894 = ~n11391 & ~n16090;
  assign n25895 = n7728 & ~n25894;
  assign n25896 = ~n25849 & ~n25895;
  assign n25897 = ~n7723 & ~n25896;
  assign n25898 = ~n25893 & ~n25897;
  assign n25899 = ~n7714 & ~n25898;
  assign n25900 = ~n25892 & ~n25899;
  assign n25901 = ~n7705 & ~n25900;
  assign n25902 = ~n25883 & ~n25901;
  assign n25903 = n7808 & ~n25902;
  assign n25904 = ~n11535 & ~n25903;
  assign n25905 = n8195 & ~n25904;
  assign n25906 = ~n25873 & ~n25905;
  assign n25907 = n8193 & ~n25906;
  assign n25908 = ~n25861 & ~n25907;
  assign n25909 = n8191 & ~n25908;
  assign n25910 = ~n11284 & ~n16257;
  assign n25911 = ~n8202 & ~n25910;
  assign n25912 = ~n8332 & ~n25911;
  assign n25913 = n7728 & ~n25912;
  assign n25914 = ~n11333 & ~n16293;
  assign n25915 = ~n8202 & ~n25914;
  assign n25916 = ~n8347 & ~n25915;
  assign n25917 = ~n7728 & ~n25916;
  assign n25918 = ~n25913 & ~n25917;
  assign n25919 = ~n7723 & ~n25918;
  assign n25920 = ~n7723 & ~n25919;
  assign n25921 = ~n7714 & ~n25920;
  assign n25922 = ~n7714 & ~n25921;
  assign n25923 = n7705 & ~n25922;
  assign n25924 = n7723 & ~n25916;
  assign n25925 = ~n11349 & ~n16311;
  assign n25926 = i_hlock8 & ~n25925;
  assign n25927 = ~n11355 & ~n16311;
  assign n25928 = ~i_hlock8 & ~n25927;
  assign n25929 = ~n25926 & ~n25928;
  assign n25930 = controllable_hmaster3 & ~n25929;
  assign n25931 = ~n8463 & ~n25930;
  assign n25932 = i_hbusreq7 & ~n25931;
  assign n25933 = i_hbusreq8 & ~n25929;
  assign n25934 = ~n11370 & ~n16326;
  assign n25935 = i_hlock8 & ~n25934;
  assign n25936 = ~n11379 & ~n16326;
  assign n25937 = ~i_hlock8 & ~n25936;
  assign n25938 = ~n25935 & ~n25937;
  assign n25939 = ~i_hbusreq8 & ~n25938;
  assign n25940 = ~n25933 & ~n25939;
  assign n25941 = controllable_hmaster3 & ~n25940;
  assign n25942 = ~n8634 & ~n25941;
  assign n25943 = ~i_hbusreq7 & ~n25942;
  assign n25944 = ~n25932 & ~n25943;
  assign n25945 = n7924 & ~n25944;
  assign n25946 = ~n8337 & ~n25945;
  assign n25947 = ~n7920 & ~n25946;
  assign n25948 = n7920 & ~n25916;
  assign n25949 = ~n25947 & ~n25948;
  assign n25950 = ~n7723 & ~n25949;
  assign n25951 = ~n25924 & ~n25950;
  assign n25952 = n7714 & ~n25951;
  assign n25953 = ~n7714 & ~n25946;
  assign n25954 = ~n25952 & ~n25953;
  assign n25955 = ~n7705 & ~n25954;
  assign n25956 = ~n25923 & ~n25955;
  assign n25957 = ~n7808 & ~n25956;
  assign n25958 = ~n7920 & ~n25912;
  assign n25959 = ~n16994 & ~n25958;
  assign n25960 = n7728 & ~n25959;
  assign n25961 = ~n7920 & ~n25916;
  assign n25962 = ~n17305 & ~n25961;
  assign n25963 = ~n7728 & ~n25962;
  assign n25964 = ~n25960 & ~n25963;
  assign n25965 = ~n7723 & ~n25964;
  assign n25966 = ~n7723 & ~n25965;
  assign n25967 = ~n7714 & ~n25966;
  assign n25968 = ~n7714 & ~n25967;
  assign n25969 = n7705 & ~n25968;
  assign n25970 = ~n18093 & ~n25961;
  assign n25971 = n7728 & ~n25970;
  assign n25972 = ~n20603 & ~n25961;
  assign n25973 = ~n7728 & ~n25972;
  assign n25974 = ~n25971 & ~n25973;
  assign n25975 = n7723 & ~n25974;
  assign n25976 = ~n7723 & ~n25972;
  assign n25977 = ~n25975 & ~n25976;
  assign n25978 = n7714 & ~n25977;
  assign n25979 = n7723 & ~n25972;
  assign n25980 = ~n21626 & ~n25947;
  assign n25981 = n7728 & ~n25980;
  assign n25982 = ~n22211 & ~n25947;
  assign n25983 = ~n7728 & ~n25982;
  assign n25984 = ~n25981 & ~n25983;
  assign n25985 = ~n7723 & ~n25984;
  assign n25986 = ~n25979 & ~n25985;
  assign n25987 = ~n7714 & ~n25986;
  assign n25988 = ~n25978 & ~n25987;
  assign n25989 = ~n7705 & ~n25988;
  assign n25990 = ~n25969 & ~n25989;
  assign n25991 = n7808 & ~n25990;
  assign n25992 = ~n25957 & ~n25991;
  assign n25993 = n8195 & ~n25992;
  assign n25994 = ~n8196 & ~n25993;
  assign n25995 = ~n8193 & ~n25994;
  assign n25996 = ~n9900 & ~n25947;
  assign n25997 = ~n7723 & ~n25996;
  assign n25998 = ~n9899 & ~n25997;
  assign n25999 = n7714 & ~n25998;
  assign n26000 = ~n25953 & ~n25999;
  assign n26001 = ~n7705 & ~n26000;
  assign n26002 = ~n9898 & ~n26001;
  assign n26003 = ~n7808 & ~n26002;
  assign n26004 = ~n23617 & ~n25947;
  assign n26005 = n7728 & ~n26004;
  assign n26006 = ~n25983 & ~n26005;
  assign n26007 = ~n7723 & ~n26006;
  assign n26008 = ~n23305 & ~n26007;
  assign n26009 = ~n7714 & ~n26008;
  assign n26010 = ~n23304 & ~n26009;
  assign n26011 = ~n7705 & ~n26010;
  assign n26012 = ~n22399 & ~n26011;
  assign n26013 = n7808 & ~n26012;
  assign n26014 = ~n26003 & ~n26013;
  assign n26015 = ~n8195 & ~n26014;
  assign n26016 = ~n11465 & ~n23660;
  assign n26017 = i_hlock8 & ~n26016;
  assign n26018 = ~n11472 & ~n23660;
  assign n26019 = ~i_hlock8 & ~n26018;
  assign n26020 = ~n26017 & ~n26019;
  assign n26021 = controllable_hmaster3 & ~n26020;
  assign n26022 = ~n10447 & ~n26021;
  assign n26023 = i_hbusreq7 & ~n26022;
  assign n26024 = i_hbusreq8 & ~n26020;
  assign n26025 = ~n11488 & ~n23720;
  assign n26026 = i_hlock8 & ~n26025;
  assign n26027 = ~n11498 & ~n23720;
  assign n26028 = ~i_hlock8 & ~n26027;
  assign n26029 = ~n26026 & ~n26028;
  assign n26030 = ~i_hbusreq8 & ~n26029;
  assign n26031 = ~n26024 & ~n26030;
  assign n26032 = controllable_hmaster3 & ~n26031;
  assign n26033 = ~n10621 & ~n26032;
  assign n26034 = ~i_hbusreq7 & ~n26033;
  assign n26035 = ~n26023 & ~n26034;
  assign n26036 = n7924 & ~n26035;
  assign n26037 = ~n10375 & ~n26036;
  assign n26038 = n8214 & ~n26037;
  assign n26039 = n8214 & ~n26038;
  assign n26040 = n8202 & ~n26039;
  assign n26041 = ~n10332 & ~n26040;
  assign n26042 = n7728 & ~n26041;
  assign n26043 = n8214 & ~n25946;
  assign n26044 = ~n8336 & ~n26043;
  assign n26045 = n8202 & ~n26044;
  assign n26046 = ~n10649 & ~n26045;
  assign n26047 = ~n7728 & ~n26046;
  assign n26048 = ~n26042 & ~n26047;
  assign n26049 = ~n7723 & ~n26048;
  assign n26050 = ~n7723 & ~n26049;
  assign n26051 = ~n7714 & ~n26050;
  assign n26052 = ~n7714 & ~n26051;
  assign n26053 = n7705 & ~n26052;
  assign n26054 = n7723 & ~n26046;
  assign n26055 = n7920 & ~n26046;
  assign n26056 = ~n25947 & ~n26055;
  assign n26057 = ~n7723 & ~n26056;
  assign n26058 = ~n26054 & ~n26057;
  assign n26059 = n7714 & ~n26058;
  assign n26060 = ~n25953 & ~n26059;
  assign n26061 = ~n7705 & ~n26060;
  assign n26062 = ~n26053 & ~n26061;
  assign n26063 = ~n7808 & ~n26062;
  assign n26064 = ~n7920 & ~n26041;
  assign n26065 = ~n24244 & ~n26064;
  assign n26066 = n7728 & ~n26065;
  assign n26067 = ~n7920 & ~n26046;
  assign n26068 = ~n24271 & ~n26067;
  assign n26069 = ~n7728 & ~n26068;
  assign n26070 = ~n26066 & ~n26069;
  assign n26071 = ~n7723 & ~n26070;
  assign n26072 = ~n7723 & ~n26071;
  assign n26073 = ~n7714 & ~n26072;
  assign n26074 = ~n7714 & ~n26073;
  assign n26075 = n7705 & ~n26074;
  assign n26076 = ~n24485 & ~n26067;
  assign n26077 = n7728 & ~n26076;
  assign n26078 = ~n25301 & ~n26067;
  assign n26079 = ~n7728 & ~n26078;
  assign n26080 = ~n26077 & ~n26079;
  assign n26081 = n7723 & ~n26080;
  assign n26082 = ~n7723 & ~n26078;
  assign n26083 = ~n26081 & ~n26082;
  assign n26084 = n7714 & ~n26083;
  assign n26085 = n7723 & ~n26078;
  assign n26086 = ~n25807 & ~n25947;
  assign n26087 = n7728 & ~n26086;
  assign n26088 = ~n25983 & ~n26087;
  assign n26089 = ~n7723 & ~n26088;
  assign n26090 = ~n26085 & ~n26089;
  assign n26091 = ~n7714 & ~n26090;
  assign n26092 = ~n26084 & ~n26091;
  assign n26093 = ~n7705 & ~n26092;
  assign n26094 = ~n26075 & ~n26093;
  assign n26095 = n7808 & ~n26094;
  assign n26096 = ~n26063 & ~n26095;
  assign n26097 = n8195 & ~n26096;
  assign n26098 = ~n26015 & ~n26097;
  assign n26099 = n8193 & ~n26098;
  assign n26100 = ~n25995 & ~n26099;
  assign n26101 = ~n8191 & ~n26100;
  assign n26102 = ~n25909 & ~n26101;
  assign n26103 = ~n8188 & ~n26102;
  assign n26104 = ~n25825 & ~n26103;
  assign n26105 = n8185 & ~n26104;
  assign n26106 = ~n11903 & ~n12974;
  assign n26107 = n7728 & ~n26106;
  assign n26108 = ~n11906 & ~n13113;
  assign n26109 = ~n7728 & ~n26108;
  assign n26110 = ~n26107 & ~n26109;
  assign n26111 = ~n7723 & ~n26110;
  assign n26112 = ~n7723 & ~n26111;
  assign n26113 = ~n7714 & ~n26112;
  assign n26114 = ~n7714 & ~n26113;
  assign n26115 = n7705 & ~n26114;
  assign n26116 = ~n11906 & ~n13802;
  assign n26117 = n7728 & ~n26116;
  assign n26118 = ~n11906 & ~n14838;
  assign n26119 = ~n7728 & ~n26118;
  assign n26120 = ~n26117 & ~n26119;
  assign n26121 = n7723 & ~n26120;
  assign n26122 = ~n7723 & ~n26118;
  assign n26123 = ~n26121 & ~n26122;
  assign n26124 = n7714 & ~n26123;
  assign n26125 = n7723 & ~n26118;
  assign n26126 = ~n11892 & ~n14838;
  assign n26127 = n7728 & ~n26126;
  assign n26128 = ~n11892 & ~n15172;
  assign n26129 = ~n7728 & ~n26128;
  assign n26130 = ~n26127 & ~n26129;
  assign n26131 = ~n7723 & ~n26130;
  assign n26132 = ~n26125 & ~n26131;
  assign n26133 = ~n7714 & ~n26132;
  assign n26134 = ~n26124 & ~n26133;
  assign n26135 = ~n7705 & ~n26134;
  assign n26136 = ~n26115 & ~n26135;
  assign n26137 = n7808 & ~n26136;
  assign n26138 = ~n11902 & ~n26137;
  assign n26139 = n8195 & ~n26138;
  assign n26140 = ~n8196 & ~n26139;
  assign n26141 = ~n8193 & ~n26140;
  assign n26142 = ~n11892 & ~n15638;
  assign n26143 = n7728 & ~n26142;
  assign n26144 = ~n26129 & ~n26143;
  assign n26145 = ~n7723 & ~n26144;
  assign n26146 = ~n15646 & ~n26145;
  assign n26147 = ~n7714 & ~n26146;
  assign n26148 = ~n15645 & ~n26147;
  assign n26149 = ~n7705 & ~n26148;
  assign n26150 = ~n10052 & ~n26149;
  assign n26151 = n7808 & ~n26150;
  assign n26152 = ~n11948 & ~n26151;
  assign n26153 = ~n8195 & ~n26152;
  assign n26154 = ~n12038 & ~n15866;
  assign n26155 = n7728 & ~n26154;
  assign n26156 = ~n12041 & ~n15875;
  assign n26157 = ~n7728 & ~n26156;
  assign n26158 = ~n26155 & ~n26157;
  assign n26159 = ~n7723 & ~n26158;
  assign n26160 = ~n7723 & ~n26159;
  assign n26161 = ~n7714 & ~n26160;
  assign n26162 = ~n7714 & ~n26161;
  assign n26163 = n7705 & ~n26162;
  assign n26164 = ~n12041 & ~n16020;
  assign n26165 = n7728 & ~n26164;
  assign n26166 = ~n12041 & ~n16090;
  assign n26167 = ~n7728 & ~n26166;
  assign n26168 = ~n26165 & ~n26167;
  assign n26169 = n7723 & ~n26168;
  assign n26170 = ~n7723 & ~n26166;
  assign n26171 = ~n26169 & ~n26170;
  assign n26172 = n7714 & ~n26171;
  assign n26173 = n7723 & ~n26166;
  assign n26174 = ~n11892 & ~n16090;
  assign n26175 = n7728 & ~n26174;
  assign n26176 = ~n26129 & ~n26175;
  assign n26177 = ~n7723 & ~n26176;
  assign n26178 = ~n26173 & ~n26177;
  assign n26179 = ~n7714 & ~n26178;
  assign n26180 = ~n26172 & ~n26179;
  assign n26181 = ~n7705 & ~n26180;
  assign n26182 = ~n26163 & ~n26181;
  assign n26183 = n7808 & ~n26182;
  assign n26184 = ~n12037 & ~n26183;
  assign n26185 = n8195 & ~n26184;
  assign n26186 = ~n26153 & ~n26185;
  assign n26187 = n8193 & ~n26186;
  assign n26188 = ~n26141 & ~n26187;
  assign n26189 = n8191 & ~n26188;
  assign n26190 = ~n11811 & ~n16259;
  assign n26191 = n7728 & ~n26190;
  assign n26192 = ~n11831 & ~n16295;
  assign n26193 = ~n7728 & ~n26192;
  assign n26194 = ~n26191 & ~n26193;
  assign n26195 = ~n7723 & ~n26194;
  assign n26196 = ~n7723 & ~n26195;
  assign n26197 = ~n7714 & ~n26196;
  assign n26198 = ~n7714 & ~n26197;
  assign n26199 = n7705 & ~n26198;
  assign n26200 = n7723 & ~n26192;
  assign n26201 = ~n11846 & ~n16313;
  assign n26202 = i_hlock7 & ~n26201;
  assign n26203 = ~n11854 & ~n16313;
  assign n26204 = ~i_hlock7 & ~n26203;
  assign n26205 = ~n26202 & ~n26204;
  assign n26206 = i_hbusreq7 & ~n26205;
  assign n26207 = ~n11870 & ~n16330;
  assign n26208 = i_hlock7 & ~n26207;
  assign n26209 = ~n11884 & ~n16330;
  assign n26210 = ~i_hlock7 & ~n26209;
  assign n26211 = ~n26208 & ~n26210;
  assign n26212 = ~i_hbusreq7 & ~n26211;
  assign n26213 = ~n26206 & ~n26212;
  assign n26214 = n7924 & ~n26213;
  assign n26215 = ~n8337 & ~n26214;
  assign n26216 = ~n7920 & ~n26215;
  assign n26217 = n7920 & ~n26192;
  assign n26218 = ~n26216 & ~n26217;
  assign n26219 = ~n7723 & ~n26218;
  assign n26220 = ~n26200 & ~n26219;
  assign n26221 = n7714 & ~n26220;
  assign n26222 = ~n7714 & ~n26215;
  assign n26223 = ~n26221 & ~n26222;
  assign n26224 = ~n7705 & ~n26223;
  assign n26225 = ~n26199 & ~n26224;
  assign n26226 = ~n7808 & ~n26225;
  assign n26227 = ~n7920 & ~n26190;
  assign n26228 = ~n16994 & ~n26227;
  assign n26229 = n7728 & ~n26228;
  assign n26230 = ~n7920 & ~n26192;
  assign n26231 = ~n17305 & ~n26230;
  assign n26232 = ~n7728 & ~n26231;
  assign n26233 = ~n26229 & ~n26232;
  assign n26234 = ~n7723 & ~n26233;
  assign n26235 = ~n7723 & ~n26234;
  assign n26236 = ~n7714 & ~n26235;
  assign n26237 = ~n7714 & ~n26236;
  assign n26238 = n7705 & ~n26237;
  assign n26239 = ~n18093 & ~n26230;
  assign n26240 = n7728 & ~n26239;
  assign n26241 = ~n20603 & ~n26230;
  assign n26242 = ~n7728 & ~n26241;
  assign n26243 = ~n26240 & ~n26242;
  assign n26244 = n7723 & ~n26243;
  assign n26245 = ~n7723 & ~n26241;
  assign n26246 = ~n26244 & ~n26245;
  assign n26247 = n7714 & ~n26246;
  assign n26248 = n7723 & ~n26241;
  assign n26249 = ~n21626 & ~n26216;
  assign n26250 = n7728 & ~n26249;
  assign n26251 = ~n22211 & ~n26216;
  assign n26252 = ~n7728 & ~n26251;
  assign n26253 = ~n26250 & ~n26252;
  assign n26254 = ~n7723 & ~n26253;
  assign n26255 = ~n26248 & ~n26254;
  assign n26256 = ~n7714 & ~n26255;
  assign n26257 = ~n26247 & ~n26256;
  assign n26258 = ~n7705 & ~n26257;
  assign n26259 = ~n26238 & ~n26258;
  assign n26260 = n7808 & ~n26259;
  assign n26261 = ~n26226 & ~n26260;
  assign n26262 = n8195 & ~n26261;
  assign n26263 = ~n8196 & ~n26262;
  assign n26264 = ~n8193 & ~n26263;
  assign n26265 = ~n9900 & ~n26216;
  assign n26266 = ~n7723 & ~n26265;
  assign n26267 = ~n9899 & ~n26266;
  assign n26268 = n7714 & ~n26267;
  assign n26269 = ~n26222 & ~n26268;
  assign n26270 = ~n7705 & ~n26269;
  assign n26271 = ~n9898 & ~n26270;
  assign n26272 = ~n7808 & ~n26271;
  assign n26273 = ~n23617 & ~n26216;
  assign n26274 = n7728 & ~n26273;
  assign n26275 = ~n26252 & ~n26274;
  assign n26276 = ~n7723 & ~n26275;
  assign n26277 = ~n23305 & ~n26276;
  assign n26278 = ~n7714 & ~n26277;
  assign n26279 = ~n23304 & ~n26278;
  assign n26280 = ~n7705 & ~n26279;
  assign n26281 = ~n22399 & ~n26280;
  assign n26282 = n7808 & ~n26281;
  assign n26283 = ~n26272 & ~n26282;
  assign n26284 = ~n8195 & ~n26283;
  assign n26285 = ~n11966 & ~n23662;
  assign n26286 = i_hlock7 & ~n26285;
  assign n26287 = ~n11974 & ~n23662;
  assign n26288 = ~i_hlock7 & ~n26287;
  assign n26289 = ~n26286 & ~n26288;
  assign n26290 = i_hbusreq7 & ~n26289;
  assign n26291 = ~n11990 & ~n23724;
  assign n26292 = i_hlock7 & ~n26291;
  assign n26293 = ~n12004 & ~n23724;
  assign n26294 = ~i_hlock7 & ~n26293;
  assign n26295 = ~n26292 & ~n26294;
  assign n26296 = ~i_hbusreq7 & ~n26295;
  assign n26297 = ~n26290 & ~n26296;
  assign n26298 = n7924 & ~n26297;
  assign n26299 = ~n10375 & ~n26298;
  assign n26300 = n8214 & ~n26299;
  assign n26301 = n8214 & ~n26300;
  assign n26302 = n8202 & ~n26301;
  assign n26303 = ~n10332 & ~n26302;
  assign n26304 = n7728 & ~n26303;
  assign n26305 = n8214 & ~n26215;
  assign n26306 = ~n8336 & ~n26305;
  assign n26307 = n8202 & ~n26306;
  assign n26308 = ~n10649 & ~n26307;
  assign n26309 = ~n7728 & ~n26308;
  assign n26310 = ~n26304 & ~n26309;
  assign n26311 = ~n7723 & ~n26310;
  assign n26312 = ~n7723 & ~n26311;
  assign n26313 = ~n7714 & ~n26312;
  assign n26314 = ~n7714 & ~n26313;
  assign n26315 = n7705 & ~n26314;
  assign n26316 = n7723 & ~n26308;
  assign n26317 = n7920 & ~n26308;
  assign n26318 = ~n26216 & ~n26317;
  assign n26319 = ~n7723 & ~n26318;
  assign n26320 = ~n26316 & ~n26319;
  assign n26321 = n7714 & ~n26320;
  assign n26322 = ~n26222 & ~n26321;
  assign n26323 = ~n7705 & ~n26322;
  assign n26324 = ~n26315 & ~n26323;
  assign n26325 = ~n7808 & ~n26324;
  assign n26326 = ~n7920 & ~n26303;
  assign n26327 = ~n24244 & ~n26326;
  assign n26328 = n7728 & ~n26327;
  assign n26329 = ~n7920 & ~n26308;
  assign n26330 = ~n24271 & ~n26329;
  assign n26331 = ~n7728 & ~n26330;
  assign n26332 = ~n26328 & ~n26331;
  assign n26333 = ~n7723 & ~n26332;
  assign n26334 = ~n7723 & ~n26333;
  assign n26335 = ~n7714 & ~n26334;
  assign n26336 = ~n7714 & ~n26335;
  assign n26337 = n7705 & ~n26336;
  assign n26338 = ~n24485 & ~n26329;
  assign n26339 = n7728 & ~n26338;
  assign n26340 = ~n25301 & ~n26329;
  assign n26341 = ~n7728 & ~n26340;
  assign n26342 = ~n26339 & ~n26341;
  assign n26343 = n7723 & ~n26342;
  assign n26344 = ~n7723 & ~n26340;
  assign n26345 = ~n26343 & ~n26344;
  assign n26346 = n7714 & ~n26345;
  assign n26347 = n7723 & ~n26340;
  assign n26348 = ~n25807 & ~n26216;
  assign n26349 = n7728 & ~n26348;
  assign n26350 = ~n26252 & ~n26349;
  assign n26351 = ~n7723 & ~n26350;
  assign n26352 = ~n26347 & ~n26351;
  assign n26353 = ~n7714 & ~n26352;
  assign n26354 = ~n26346 & ~n26353;
  assign n26355 = ~n7705 & ~n26354;
  assign n26356 = ~n26337 & ~n26355;
  assign n26357 = n7808 & ~n26356;
  assign n26358 = ~n26325 & ~n26357;
  assign n26359 = n8195 & ~n26358;
  assign n26360 = ~n26284 & ~n26359;
  assign n26361 = n8193 & ~n26360;
  assign n26362 = ~n26264 & ~n26361;
  assign n26363 = ~n8191 & ~n26362;
  assign n26364 = ~n26189 & ~n26363;
  assign n26365 = n8188 & ~n26364;
  assign n26366 = ~n12289 & ~n12974;
  assign n26367 = n7728 & ~n26366;
  assign n26368 = ~n12292 & ~n13113;
  assign n26369 = ~n7728 & ~n26368;
  assign n26370 = ~n26367 & ~n26369;
  assign n26371 = ~n7723 & ~n26370;
  assign n26372 = ~n7723 & ~n26371;
  assign n26373 = ~n7714 & ~n26372;
  assign n26374 = ~n7714 & ~n26373;
  assign n26375 = n7705 & ~n26374;
  assign n26376 = ~n12292 & ~n13802;
  assign n26377 = n7728 & ~n26376;
  assign n26378 = ~n12292 & ~n14838;
  assign n26379 = ~n7728 & ~n26378;
  assign n26380 = ~n26377 & ~n26379;
  assign n26381 = n7723 & ~n26380;
  assign n26382 = ~n7723 & ~n26378;
  assign n26383 = ~n26381 & ~n26382;
  assign n26384 = n7714 & ~n26383;
  assign n26385 = n7723 & ~n26378;
  assign n26386 = ~n12278 & ~n14838;
  assign n26387 = n7728 & ~n26386;
  assign n26388 = ~n12278 & ~n15172;
  assign n26389 = ~n7728 & ~n26388;
  assign n26390 = ~n26387 & ~n26389;
  assign n26391 = ~n7723 & ~n26390;
  assign n26392 = ~n26385 & ~n26391;
  assign n26393 = ~n7714 & ~n26392;
  assign n26394 = ~n26384 & ~n26393;
  assign n26395 = ~n7705 & ~n26394;
  assign n26396 = ~n26375 & ~n26395;
  assign n26397 = n7808 & ~n26396;
  assign n26398 = ~n12288 & ~n26397;
  assign n26399 = n8195 & ~n26398;
  assign n26400 = ~n8196 & ~n26399;
  assign n26401 = ~n8193 & ~n26400;
  assign n26402 = ~n12278 & ~n15638;
  assign n26403 = n7728 & ~n26402;
  assign n26404 = ~n26389 & ~n26403;
  assign n26405 = ~n7723 & ~n26404;
  assign n26406 = ~n15646 & ~n26405;
  assign n26407 = ~n7714 & ~n26406;
  assign n26408 = ~n15645 & ~n26407;
  assign n26409 = ~n7705 & ~n26408;
  assign n26410 = ~n10052 & ~n26409;
  assign n26411 = n7808 & ~n26410;
  assign n26412 = ~n12334 & ~n26411;
  assign n26413 = ~n8195 & ~n26412;
  assign n26414 = ~n12388 & ~n15866;
  assign n26415 = n7728 & ~n26414;
  assign n26416 = ~n12391 & ~n15875;
  assign n26417 = ~n7728 & ~n26416;
  assign n26418 = ~n26415 & ~n26417;
  assign n26419 = ~n7723 & ~n26418;
  assign n26420 = ~n7723 & ~n26419;
  assign n26421 = ~n7714 & ~n26420;
  assign n26422 = ~n7714 & ~n26421;
  assign n26423 = n7705 & ~n26422;
  assign n26424 = ~n12391 & ~n16020;
  assign n26425 = n7728 & ~n26424;
  assign n26426 = ~n12391 & ~n16090;
  assign n26427 = ~n7728 & ~n26426;
  assign n26428 = ~n26425 & ~n26427;
  assign n26429 = n7723 & ~n26428;
  assign n26430 = ~n7723 & ~n26426;
  assign n26431 = ~n26429 & ~n26430;
  assign n26432 = n7714 & ~n26431;
  assign n26433 = n7723 & ~n26426;
  assign n26434 = ~n12278 & ~n16090;
  assign n26435 = n7728 & ~n26434;
  assign n26436 = ~n26389 & ~n26435;
  assign n26437 = ~n7723 & ~n26436;
  assign n26438 = ~n26433 & ~n26437;
  assign n26439 = ~n7714 & ~n26438;
  assign n26440 = ~n26432 & ~n26439;
  assign n26441 = ~n7705 & ~n26440;
  assign n26442 = ~n26423 & ~n26441;
  assign n26443 = n7808 & ~n26442;
  assign n26444 = ~n12387 & ~n26443;
  assign n26445 = n8195 & ~n26444;
  assign n26446 = ~n26413 & ~n26445;
  assign n26447 = n8193 & ~n26446;
  assign n26448 = ~n26401 & ~n26447;
  assign n26449 = n8191 & ~n26448;
  assign n26450 = ~n11811 & ~n25911;
  assign n26451 = n7728 & ~n26450;
  assign n26452 = ~n11831 & ~n25915;
  assign n26453 = ~n7728 & ~n26452;
  assign n26454 = ~n26451 & ~n26453;
  assign n26455 = ~n7723 & ~n26454;
  assign n26456 = ~n7723 & ~n26455;
  assign n26457 = ~n7714 & ~n26456;
  assign n26458 = ~n7714 & ~n26457;
  assign n26459 = n7705 & ~n26458;
  assign n26460 = n7723 & ~n26452;
  assign n26461 = ~n11846 & ~n25930;
  assign n26462 = i_hlock7 & ~n26461;
  assign n26463 = ~n11854 & ~n25930;
  assign n26464 = ~i_hlock7 & ~n26463;
  assign n26465 = ~n26462 & ~n26464;
  assign n26466 = i_hbusreq7 & ~n26465;
  assign n26467 = ~n11870 & ~n25941;
  assign n26468 = i_hlock7 & ~n26467;
  assign n26469 = ~n11884 & ~n25941;
  assign n26470 = ~i_hlock7 & ~n26469;
  assign n26471 = ~n26468 & ~n26470;
  assign n26472 = ~i_hbusreq7 & ~n26471;
  assign n26473 = ~n26466 & ~n26472;
  assign n26474 = n7924 & ~n26473;
  assign n26475 = ~n8337 & ~n26474;
  assign n26476 = ~n7920 & ~n26475;
  assign n26477 = n7920 & ~n26452;
  assign n26478 = ~n26476 & ~n26477;
  assign n26479 = ~n7723 & ~n26478;
  assign n26480 = ~n26460 & ~n26479;
  assign n26481 = n7714 & ~n26480;
  assign n26482 = ~n7714 & ~n26475;
  assign n26483 = ~n26481 & ~n26482;
  assign n26484 = ~n7705 & ~n26483;
  assign n26485 = ~n26459 & ~n26484;
  assign n26486 = ~n7808 & ~n26485;
  assign n26487 = ~n7920 & ~n26450;
  assign n26488 = ~n16994 & ~n26487;
  assign n26489 = n7728 & ~n26488;
  assign n26490 = ~n7920 & ~n26452;
  assign n26491 = ~n17305 & ~n26490;
  assign n26492 = ~n7728 & ~n26491;
  assign n26493 = ~n26489 & ~n26492;
  assign n26494 = ~n7723 & ~n26493;
  assign n26495 = ~n7723 & ~n26494;
  assign n26496 = ~n7714 & ~n26495;
  assign n26497 = ~n7714 & ~n26496;
  assign n26498 = n7705 & ~n26497;
  assign n26499 = ~n18093 & ~n26490;
  assign n26500 = n7728 & ~n26499;
  assign n26501 = ~n20603 & ~n26490;
  assign n26502 = ~n7728 & ~n26501;
  assign n26503 = ~n26500 & ~n26502;
  assign n26504 = n7723 & ~n26503;
  assign n26505 = ~n7723 & ~n26501;
  assign n26506 = ~n26504 & ~n26505;
  assign n26507 = n7714 & ~n26506;
  assign n26508 = n7723 & ~n26501;
  assign n26509 = ~n21626 & ~n26476;
  assign n26510 = n7728 & ~n26509;
  assign n26511 = ~n22211 & ~n26476;
  assign n26512 = ~n7728 & ~n26511;
  assign n26513 = ~n26510 & ~n26512;
  assign n26514 = ~n7723 & ~n26513;
  assign n26515 = ~n26508 & ~n26514;
  assign n26516 = ~n7714 & ~n26515;
  assign n26517 = ~n26507 & ~n26516;
  assign n26518 = ~n7705 & ~n26517;
  assign n26519 = ~n26498 & ~n26518;
  assign n26520 = n7808 & ~n26519;
  assign n26521 = ~n26486 & ~n26520;
  assign n26522 = n8195 & ~n26521;
  assign n26523 = ~n8196 & ~n26522;
  assign n26524 = ~n8193 & ~n26523;
  assign n26525 = ~n9900 & ~n26476;
  assign n26526 = ~n7723 & ~n26525;
  assign n26527 = ~n9899 & ~n26526;
  assign n26528 = n7714 & ~n26527;
  assign n26529 = ~n26482 & ~n26528;
  assign n26530 = ~n7705 & ~n26529;
  assign n26531 = ~n9898 & ~n26530;
  assign n26532 = ~n7808 & ~n26531;
  assign n26533 = ~n23617 & ~n26476;
  assign n26534 = n7728 & ~n26533;
  assign n26535 = ~n26512 & ~n26534;
  assign n26536 = ~n7723 & ~n26535;
  assign n26537 = ~n23305 & ~n26536;
  assign n26538 = ~n7714 & ~n26537;
  assign n26539 = ~n23304 & ~n26538;
  assign n26540 = ~n7705 & ~n26539;
  assign n26541 = ~n22399 & ~n26540;
  assign n26542 = n7808 & ~n26541;
  assign n26543 = ~n26532 & ~n26542;
  assign n26544 = ~n8195 & ~n26543;
  assign n26545 = ~n11966 & ~n26021;
  assign n26546 = i_hlock7 & ~n26545;
  assign n26547 = ~n11974 & ~n26021;
  assign n26548 = ~i_hlock7 & ~n26547;
  assign n26549 = ~n26546 & ~n26548;
  assign n26550 = i_hbusreq7 & ~n26549;
  assign n26551 = ~n11990 & ~n26032;
  assign n26552 = i_hlock7 & ~n26551;
  assign n26553 = ~n12004 & ~n26032;
  assign n26554 = ~i_hlock7 & ~n26553;
  assign n26555 = ~n26552 & ~n26554;
  assign n26556 = ~i_hbusreq7 & ~n26555;
  assign n26557 = ~n26550 & ~n26556;
  assign n26558 = n7924 & ~n26557;
  assign n26559 = ~n10375 & ~n26558;
  assign n26560 = n8214 & ~n26559;
  assign n26561 = n8214 & ~n26560;
  assign n26562 = n8202 & ~n26561;
  assign n26563 = ~n10332 & ~n26562;
  assign n26564 = n7728 & ~n26563;
  assign n26565 = n8214 & ~n26475;
  assign n26566 = ~n8336 & ~n26565;
  assign n26567 = n8202 & ~n26566;
  assign n26568 = ~n10649 & ~n26567;
  assign n26569 = ~n7728 & ~n26568;
  assign n26570 = ~n26564 & ~n26569;
  assign n26571 = ~n7723 & ~n26570;
  assign n26572 = ~n7723 & ~n26571;
  assign n26573 = ~n7714 & ~n26572;
  assign n26574 = ~n7714 & ~n26573;
  assign n26575 = n7705 & ~n26574;
  assign n26576 = n7723 & ~n26568;
  assign n26577 = n7920 & ~n26568;
  assign n26578 = ~n26476 & ~n26577;
  assign n26579 = ~n7723 & ~n26578;
  assign n26580 = ~n26576 & ~n26579;
  assign n26581 = n7714 & ~n26580;
  assign n26582 = ~n26482 & ~n26581;
  assign n26583 = ~n7705 & ~n26582;
  assign n26584 = ~n26575 & ~n26583;
  assign n26585 = ~n7808 & ~n26584;
  assign n26586 = ~n7920 & ~n26563;
  assign n26587 = ~n24244 & ~n26586;
  assign n26588 = n7728 & ~n26587;
  assign n26589 = ~n7920 & ~n26568;
  assign n26590 = ~n24271 & ~n26589;
  assign n26591 = ~n7728 & ~n26590;
  assign n26592 = ~n26588 & ~n26591;
  assign n26593 = ~n7723 & ~n26592;
  assign n26594 = ~n7723 & ~n26593;
  assign n26595 = ~n7714 & ~n26594;
  assign n26596 = ~n7714 & ~n26595;
  assign n26597 = n7705 & ~n26596;
  assign n26598 = ~n24485 & ~n26589;
  assign n26599 = n7728 & ~n26598;
  assign n26600 = ~n25301 & ~n26589;
  assign n26601 = ~n7728 & ~n26600;
  assign n26602 = ~n26599 & ~n26601;
  assign n26603 = n7723 & ~n26602;
  assign n26604 = ~n7723 & ~n26600;
  assign n26605 = ~n26603 & ~n26604;
  assign n26606 = n7714 & ~n26605;
  assign n26607 = n7723 & ~n26600;
  assign n26608 = ~n25807 & ~n26476;
  assign n26609 = n7728 & ~n26608;
  assign n26610 = ~n26512 & ~n26609;
  assign n26611 = ~n7723 & ~n26610;
  assign n26612 = ~n26607 & ~n26611;
  assign n26613 = ~n7714 & ~n26612;
  assign n26614 = ~n26606 & ~n26613;
  assign n26615 = ~n7705 & ~n26614;
  assign n26616 = ~n26597 & ~n26615;
  assign n26617 = n7808 & ~n26616;
  assign n26618 = ~n26585 & ~n26617;
  assign n26619 = n8195 & ~n26618;
  assign n26620 = ~n26544 & ~n26619;
  assign n26621 = n8193 & ~n26620;
  assign n26622 = ~n26524 & ~n26621;
  assign n26623 = ~n8191 & ~n26622;
  assign n26624 = ~n26449 & ~n26623;
  assign n26625 = ~n8188 & ~n26624;
  assign n26626 = ~n26365 & ~n26625;
  assign n26627 = ~n8185 & ~n26626;
  assign n26628 = ~n26105 & ~n26627;
  assign n26629 = ~controllable_hgrant8 & ~n26628;
  assign n26630 = ~n12606 & ~n26629;
  assign n26631 = controllable_nhgrant0 & ~n26630;
  assign n26632 = ~controllable_nhgrant0 & ~n12604;
  assign n26633 = ~n26631 & ~n26632;
  assign n26634 = ~controllable_hgrant7 & ~n26633;
  assign n26635 = ~n12605 & ~n26634;
  assign n26636 = controllable_hgrant9 & ~n26635;
  assign n26637 = ~controllable_hgrant4 & ~n12635;
  assign n26638 = ~n13408 & ~n26637;
  assign n26639 = ~controllable_hgrant5 & ~n26638;
  assign n26640 = ~n13407 & ~n26639;
  assign n26641 = controllable_hmaster2 & ~n26640;
  assign n26642 = controllable_hmaster2 & ~n26641;
  assign n26643 = controllable_hmaster1 & ~n26642;
  assign n26644 = controllable_hmaster1 & ~n26643;
  assign n26645 = ~controllable_hgrant6 & ~n26644;
  assign n26646 = ~n16895 & ~n26645;
  assign n26647 = controllable_hmaster0 & ~n26646;
  assign n26648 = controllable_hmaster0 & ~n26647;
  assign n26649 = ~controllable_hmaster3 & ~n26648;
  assign n26650 = ~controllable_hmaster3 & ~n26649;
  assign n26651 = i_hlock7 & ~n26650;
  assign n26652 = ~controllable_hgrant4 & ~n12653;
  assign n26653 = ~n13429 & ~n26652;
  assign n26654 = ~controllable_hgrant5 & ~n26653;
  assign n26655 = ~n13428 & ~n26654;
  assign n26656 = controllable_hmaster2 & ~n26655;
  assign n26657 = controllable_hmaster2 & ~n26656;
  assign n26658 = controllable_hmaster1 & ~n26657;
  assign n26659 = controllable_hmaster1 & ~n26658;
  assign n26660 = ~controllable_hgrant6 & ~n26659;
  assign n26661 = ~n16907 & ~n26660;
  assign n26662 = controllable_hmaster0 & ~n26661;
  assign n26663 = controllable_hmaster0 & ~n26662;
  assign n26664 = ~controllable_hmaster3 & ~n26663;
  assign n26665 = ~controllable_hmaster3 & ~n26664;
  assign n26666 = ~i_hlock7 & ~n26665;
  assign n26667 = ~n26651 & ~n26666;
  assign n26668 = i_hbusreq7 & ~n26667;
  assign n26669 = i_hbusreq8 & ~n26648;
  assign n26670 = i_hbusreq6 & ~n26644;
  assign n26671 = i_hbusreq5 & ~n26638;
  assign n26672 = i_hbusreq4 & ~n12635;
  assign n26673 = i_hbusreq9 & ~n12635;
  assign n26674 = ~i_hbusreq9 & ~n12726;
  assign n26675 = ~n26673 & ~n26674;
  assign n26676 = ~i_hbusreq4 & ~n26675;
  assign n26677 = ~n26672 & ~n26676;
  assign n26678 = ~controllable_hgrant4 & ~n26677;
  assign n26679 = ~n13524 & ~n26678;
  assign n26680 = ~i_hbusreq5 & ~n26679;
  assign n26681 = ~n26671 & ~n26680;
  assign n26682 = ~controllable_hgrant5 & ~n26681;
  assign n26683 = ~n13522 & ~n26682;
  assign n26684 = controllable_hmaster2 & ~n26683;
  assign n26685 = controllable_hmaster2 & ~n26684;
  assign n26686 = controllable_hmaster1 & ~n26685;
  assign n26687 = controllable_hmaster1 & ~n26686;
  assign n26688 = ~i_hbusreq6 & ~n26687;
  assign n26689 = ~n26670 & ~n26688;
  assign n26690 = ~controllable_hgrant6 & ~n26689;
  assign n26691 = ~n16922 & ~n26690;
  assign n26692 = controllable_hmaster0 & ~n26691;
  assign n26693 = controllable_hmaster0 & ~n26692;
  assign n26694 = ~i_hbusreq8 & ~n26693;
  assign n26695 = ~n26669 & ~n26694;
  assign n26696 = ~controllable_hmaster3 & ~n26695;
  assign n26697 = ~controllable_hmaster3 & ~n26696;
  assign n26698 = i_hlock7 & ~n26697;
  assign n26699 = i_hbusreq8 & ~n26663;
  assign n26700 = i_hbusreq6 & ~n26659;
  assign n26701 = i_hbusreq5 & ~n26653;
  assign n26702 = i_hbusreq4 & ~n12653;
  assign n26703 = i_hbusreq9 & ~n12653;
  assign n26704 = ~i_hbusreq9 & ~n12751;
  assign n26705 = ~n26703 & ~n26704;
  assign n26706 = ~i_hbusreq4 & ~n26705;
  assign n26707 = ~n26702 & ~n26706;
  assign n26708 = ~controllable_hgrant4 & ~n26707;
  assign n26709 = ~n13577 & ~n26708;
  assign n26710 = ~i_hbusreq5 & ~n26709;
  assign n26711 = ~n26701 & ~n26710;
  assign n26712 = ~controllable_hgrant5 & ~n26711;
  assign n26713 = ~n13575 & ~n26712;
  assign n26714 = controllable_hmaster2 & ~n26713;
  assign n26715 = controllable_hmaster2 & ~n26714;
  assign n26716 = controllable_hmaster1 & ~n26715;
  assign n26717 = controllable_hmaster1 & ~n26716;
  assign n26718 = ~i_hbusreq6 & ~n26717;
  assign n26719 = ~n26700 & ~n26718;
  assign n26720 = ~controllable_hgrant6 & ~n26719;
  assign n26721 = ~n16940 & ~n26720;
  assign n26722 = controllable_hmaster0 & ~n26721;
  assign n26723 = controllable_hmaster0 & ~n26722;
  assign n26724 = ~i_hbusreq8 & ~n26723;
  assign n26725 = ~n26699 & ~n26724;
  assign n26726 = ~controllable_hmaster3 & ~n26725;
  assign n26727 = ~controllable_hmaster3 & ~n26726;
  assign n26728 = ~i_hlock7 & ~n26727;
  assign n26729 = ~n26698 & ~n26728;
  assign n26730 = ~i_hbusreq7 & ~n26729;
  assign n26731 = ~n26668 & ~n26730;
  assign n26732 = ~n7924 & ~n26731;
  assign n26733 = controllable_hmaster3 & ~n12829;
  assign n26734 = ~controllable_hgrant4 & ~n12808;
  assign n26735 = ~n13408 & ~n26734;
  assign n26736 = ~controllable_hgrant5 & ~n26735;
  assign n26737 = ~n13407 & ~n26736;
  assign n26738 = controllable_hmaster2 & ~n26737;
  assign n26739 = ~n13032 & ~n26738;
  assign n26740 = controllable_hmaster1 & ~n26739;
  assign n26741 = ~controllable_hmaster1 & ~n12796;
  assign n26742 = ~n26740 & ~n26741;
  assign n26743 = ~controllable_hgrant6 & ~n26742;
  assign n26744 = ~n16895 & ~n26743;
  assign n26745 = controllable_hmaster0 & ~n26744;
  assign n26746 = ~n12830 & ~n26745;
  assign n26747 = ~controllable_hmaster3 & ~n26746;
  assign n26748 = ~n26733 & ~n26747;
  assign n26749 = i_hlock7 & ~n26748;
  assign n26750 = ~controllable_hgrant4 & ~n12814;
  assign n26751 = ~n13429 & ~n26750;
  assign n26752 = ~controllable_hgrant5 & ~n26751;
  assign n26753 = ~n13428 & ~n26752;
  assign n26754 = controllable_hmaster2 & ~n26753;
  assign n26755 = ~n13032 & ~n26754;
  assign n26756 = controllable_hmaster1 & ~n26755;
  assign n26757 = ~n26741 & ~n26756;
  assign n26758 = ~controllable_hgrant6 & ~n26757;
  assign n26759 = ~n16907 & ~n26758;
  assign n26760 = controllable_hmaster0 & ~n26759;
  assign n26761 = ~n12830 & ~n26760;
  assign n26762 = ~controllable_hmaster3 & ~n26761;
  assign n26763 = ~n26733 & ~n26762;
  assign n26764 = ~i_hlock7 & ~n26763;
  assign n26765 = ~n26749 & ~n26764;
  assign n26766 = i_hbusreq7 & ~n26765;
  assign n26767 = controllable_hmaster3 & ~n12963;
  assign n26768 = i_hbusreq8 & ~n26746;
  assign n26769 = i_hbusreq6 & ~n26742;
  assign n26770 = i_hbusreq5 & ~n26735;
  assign n26771 = i_hbusreq4 & ~n12808;
  assign n26772 = i_hbusreq9 & ~n12808;
  assign n26773 = ~i_hbusreq9 & ~n12917;
  assign n26774 = ~n26772 & ~n26773;
  assign n26775 = ~i_hbusreq4 & ~n26774;
  assign n26776 = ~n26771 & ~n26775;
  assign n26777 = ~controllable_hgrant4 & ~n26776;
  assign n26778 = ~n13524 & ~n26777;
  assign n26779 = ~i_hbusreq5 & ~n26778;
  assign n26780 = ~n26770 & ~n26779;
  assign n26781 = ~controllable_hgrant5 & ~n26780;
  assign n26782 = ~n13522 & ~n26781;
  assign n26783 = controllable_hmaster2 & ~n26782;
  assign n26784 = ~n13091 & ~n26783;
  assign n26785 = controllable_hmaster1 & ~n26784;
  assign n26786 = ~controllable_hmaster1 & ~n12875;
  assign n26787 = ~n26785 & ~n26786;
  assign n26788 = ~i_hbusreq6 & ~n26787;
  assign n26789 = ~n26769 & ~n26788;
  assign n26790 = ~controllable_hgrant6 & ~n26789;
  assign n26791 = ~n16922 & ~n26790;
  assign n26792 = controllable_hmaster0 & ~n26791;
  assign n26793 = ~n12956 & ~n26792;
  assign n26794 = ~i_hbusreq8 & ~n26793;
  assign n26795 = ~n26768 & ~n26794;
  assign n26796 = ~controllable_hmaster3 & ~n26795;
  assign n26797 = ~n26767 & ~n26796;
  assign n26798 = i_hlock7 & ~n26797;
  assign n26799 = i_hbusreq8 & ~n26761;
  assign n26800 = i_hbusreq6 & ~n26757;
  assign n26801 = i_hbusreq5 & ~n26751;
  assign n26802 = i_hbusreq4 & ~n12814;
  assign n26803 = i_hbusreq9 & ~n12814;
  assign n26804 = ~i_hbusreq9 & ~n12929;
  assign n26805 = ~n26803 & ~n26804;
  assign n26806 = ~i_hbusreq4 & ~n26805;
  assign n26807 = ~n26802 & ~n26806;
  assign n26808 = ~controllable_hgrant4 & ~n26807;
  assign n26809 = ~n13577 & ~n26808;
  assign n26810 = ~i_hbusreq5 & ~n26809;
  assign n26811 = ~n26801 & ~n26810;
  assign n26812 = ~controllable_hgrant5 & ~n26811;
  assign n26813 = ~n13575 & ~n26812;
  assign n26814 = controllable_hmaster2 & ~n26813;
  assign n26815 = ~n13091 & ~n26814;
  assign n26816 = controllable_hmaster1 & ~n26815;
  assign n26817 = ~n26786 & ~n26816;
  assign n26818 = ~i_hbusreq6 & ~n26817;
  assign n26819 = ~n26800 & ~n26818;
  assign n26820 = ~controllable_hgrant6 & ~n26819;
  assign n26821 = ~n16940 & ~n26820;
  assign n26822 = controllable_hmaster0 & ~n26821;
  assign n26823 = ~n12956 & ~n26822;
  assign n26824 = ~i_hbusreq8 & ~n26823;
  assign n26825 = ~n26799 & ~n26824;
  assign n26826 = ~controllable_hmaster3 & ~n26825;
  assign n26827 = ~n26767 & ~n26826;
  assign n26828 = ~i_hlock7 & ~n26827;
  assign n26829 = ~n26798 & ~n26828;
  assign n26830 = ~i_hbusreq7 & ~n26829;
  assign n26831 = ~n26766 & ~n26830;
  assign n26832 = n7924 & ~n26831;
  assign n26833 = ~n26732 & ~n26832;
  assign n26834 = ~n8214 & ~n26833;
  assign n26835 = ~n8870 & ~n26834;
  assign n26836 = n8202 & ~n26835;
  assign n26837 = ~n8792 & ~n26836;
  assign n26838 = n7920 & ~n26837;
  assign n26839 = ~n8651 & ~n26838;
  assign n26840 = n7728 & ~n26839;
  assign n26841 = ~n7743 & ~n26649;
  assign n26842 = i_hlock7 & ~n26841;
  assign n26843 = ~n7743 & ~n26664;
  assign n26844 = ~i_hlock7 & ~n26843;
  assign n26845 = ~n26842 & ~n26844;
  assign n26846 = i_hbusreq7 & ~n26845;
  assign n26847 = ~n7779 & ~n26696;
  assign n26848 = i_hlock7 & ~n26847;
  assign n26849 = ~n7779 & ~n26726;
  assign n26850 = ~i_hlock7 & ~n26849;
  assign n26851 = ~n26848 & ~n26850;
  assign n26852 = ~i_hbusreq7 & ~n26851;
  assign n26853 = ~n26846 & ~n26852;
  assign n26854 = ~n7924 & ~n26853;
  assign n26855 = controllable_hmaster3 & ~n13037;
  assign n26856 = ~n26747 & ~n26855;
  assign n26857 = i_hlock7 & ~n26856;
  assign n26858 = ~n26762 & ~n26855;
  assign n26859 = ~i_hlock7 & ~n26858;
  assign n26860 = ~n26857 & ~n26859;
  assign n26861 = i_hbusreq7 & ~n26860;
  assign n26862 = i_hbusreq8 & ~n13037;
  assign n26863 = ~i_hbusreq8 & ~n13098;
  assign n26864 = ~n26862 & ~n26863;
  assign n26865 = controllable_hmaster3 & ~n26864;
  assign n26866 = ~n26796 & ~n26865;
  assign n26867 = i_hlock7 & ~n26866;
  assign n26868 = ~n26826 & ~n26865;
  assign n26869 = ~i_hlock7 & ~n26868;
  assign n26870 = ~n26867 & ~n26869;
  assign n26871 = ~i_hbusreq7 & ~n26870;
  assign n26872 = ~n26861 & ~n26871;
  assign n26873 = n7924 & ~n26872;
  assign n26874 = ~n26854 & ~n26873;
  assign n26875 = ~n8214 & ~n26874;
  assign n26876 = ~n8970 & ~n26875;
  assign n26877 = n8202 & ~n26876;
  assign n26878 = ~n8950 & ~n26877;
  assign n26879 = n7920 & ~n26878;
  assign n26880 = ~n8877 & ~n26879;
  assign n26881 = ~n7728 & ~n26880;
  assign n26882 = ~n26840 & ~n26881;
  assign n26883 = ~n7723 & ~n26882;
  assign n26884 = ~n7723 & ~n26883;
  assign n26885 = ~n7714 & ~n26884;
  assign n26886 = ~n7714 & ~n26885;
  assign n26887 = n7705 & ~n26886;
  assign n26888 = controllable_hmaster2 & ~n13321;
  assign n26889 = ~n8988 & ~n26888;
  assign n26890 = controllable_hmaster1 & ~n26889;
  assign n26891 = ~n9096 & ~n26890;
  assign n26892 = ~controllable_hgrant6 & ~n26891;
  assign n26893 = ~n13198 & ~n26892;
  assign n26894 = controllable_hmaster0 & ~n26893;
  assign n26895 = ~n9099 & ~n26894;
  assign n26896 = ~controllable_hmaster3 & ~n26895;
  assign n26897 = ~n8994 & ~n26896;
  assign n26898 = i_hbusreq7 & ~n26897;
  assign n26899 = i_hbusreq8 & ~n26895;
  assign n26900 = i_hbusreq6 & ~n26891;
  assign n26901 = controllable_hmaster2 & ~n13368;
  assign n26902 = ~n9024 & ~n26901;
  assign n26903 = controllable_hmaster1 & ~n26902;
  assign n26904 = ~n9122 & ~n26903;
  assign n26905 = ~i_hbusreq6 & ~n26904;
  assign n26906 = ~n26900 & ~n26905;
  assign n26907 = ~controllable_hgrant6 & ~n26906;
  assign n26908 = ~n13298 & ~n26907;
  assign n26909 = controllable_hmaster0 & ~n26908;
  assign n26910 = ~n9127 & ~n26909;
  assign n26911 = ~i_hbusreq8 & ~n26910;
  assign n26912 = ~n26899 & ~n26911;
  assign n26913 = ~controllable_hmaster3 & ~n26912;
  assign n26914 = ~n9034 & ~n26913;
  assign n26915 = ~i_hbusreq7 & ~n26914;
  assign n26916 = ~n26898 & ~n26915;
  assign n26917 = ~n7924 & ~n26916;
  assign n26918 = i_hlock9 & ~n13413;
  assign n26919 = ~i_hlock9 & ~n13434;
  assign n26920 = ~n26918 & ~n26919;
  assign n26921 = ~controllable_hgrant4 & ~n26920;
  assign n26922 = ~n12609 & ~n26921;
  assign n26923 = ~controllable_hgrant5 & ~n26922;
  assign n26924 = ~n12608 & ~n26923;
  assign n26925 = ~controllable_hmaster2 & ~n26924;
  assign n26926 = ~n13168 & ~n26925;
  assign n26927 = ~controllable_hmaster1 & ~n26926;
  assign n26928 = ~n13167 & ~n26927;
  assign n26929 = ~controllable_hgrant6 & ~n26928;
  assign n26930 = ~n13122 & ~n26929;
  assign n26931 = controllable_hmaster0 & ~n26930;
  assign n26932 = ~n13195 & ~n26931;
  assign n26933 = controllable_hmaster3 & ~n26932;
  assign n26934 = controllable_hmaster2 & ~n13398;
  assign n26935 = ~n13189 & ~n26934;
  assign n26936 = controllable_hmaster1 & ~n26935;
  assign n26937 = ~n13677 & ~n26936;
  assign n26938 = ~controllable_hgrant6 & ~n26937;
  assign n26939 = ~n13198 & ~n26938;
  assign n26940 = controllable_hmaster0 & ~n26939;
  assign n26941 = ~n13682 & ~n26940;
  assign n26942 = ~controllable_hmaster3 & ~n26941;
  assign n26943 = ~n26933 & ~n26942;
  assign n26944 = i_hbusreq7 & ~n26943;
  assign n26945 = i_hbusreq8 & ~n26932;
  assign n26946 = i_hbusreq6 & ~n26928;
  assign n26947 = i_hbusreq5 & ~n26922;
  assign n26948 = i_hbusreq4 & ~n26920;
  assign n26949 = i_hbusreq9 & ~n26920;
  assign n26950 = i_hlock9 & ~n13551;
  assign n26951 = ~i_hlock9 & ~n13590;
  assign n26952 = ~n26950 & ~n26951;
  assign n26953 = ~i_hbusreq9 & ~n26952;
  assign n26954 = ~n26949 & ~n26953;
  assign n26955 = ~i_hbusreq4 & ~n26954;
  assign n26956 = ~n26948 & ~n26955;
  assign n26957 = ~controllable_hgrant4 & ~n26956;
  assign n26958 = ~n12676 & ~n26957;
  assign n26959 = ~i_hbusreq5 & ~n26958;
  assign n26960 = ~n26947 & ~n26959;
  assign n26961 = ~controllable_hgrant5 & ~n26960;
  assign n26962 = ~n12674 & ~n26961;
  assign n26963 = ~controllable_hmaster2 & ~n26962;
  assign n26964 = ~n13480 & ~n26963;
  assign n26965 = ~controllable_hmaster1 & ~n26964;
  assign n26966 = ~n13479 & ~n26965;
  assign n26967 = ~i_hbusreq6 & ~n26966;
  assign n26968 = ~n26946 & ~n26967;
  assign n26969 = ~controllable_hgrant6 & ~n26968;
  assign n26970 = ~n13134 & ~n26969;
  assign n26971 = controllable_hmaster0 & ~n26970;
  assign n26972 = ~n13710 & ~n26971;
  assign n26973 = ~i_hbusreq8 & ~n26972;
  assign n26974 = ~n26945 & ~n26973;
  assign n26975 = controllable_hmaster3 & ~n26974;
  assign n26976 = i_hbusreq8 & ~n26941;
  assign n26977 = i_hbusreq6 & ~n26937;
  assign n26978 = controllable_hmaster2 & ~n13510;
  assign n26979 = ~n13702 & ~n26978;
  assign n26980 = controllable_hmaster1 & ~n26979;
  assign n26981 = ~n13721 & ~n26980;
  assign n26982 = ~i_hbusreq6 & ~n26981;
  assign n26983 = ~n26977 & ~n26982;
  assign n26984 = ~controllable_hgrant6 & ~n26983;
  assign n26985 = ~n13298 & ~n26984;
  assign n26986 = controllable_hmaster0 & ~n26985;
  assign n26987 = ~n13728 & ~n26986;
  assign n26988 = ~i_hbusreq8 & ~n26987;
  assign n26989 = ~n26976 & ~n26988;
  assign n26990 = ~controllable_hmaster3 & ~n26989;
  assign n26991 = ~n26975 & ~n26990;
  assign n26992 = ~i_hbusreq7 & ~n26991;
  assign n26993 = ~n26944 & ~n26992;
  assign n26994 = n7924 & ~n26993;
  assign n26995 = ~n26917 & ~n26994;
  assign n26996 = ~n8214 & ~n26995;
  assign n26997 = ~n9060 & ~n26896;
  assign n26998 = i_hbusreq7 & ~n26997;
  assign n26999 = ~n9086 & ~n26913;
  assign n27000 = ~i_hbusreq7 & ~n26999;
  assign n27001 = ~n26998 & ~n27000;
  assign n27002 = ~n7924 & ~n27001;
  assign n27003 = controllable_hmaster0 & ~n13194;
  assign n27004 = ~n13424 & ~n27003;
  assign n27005 = i_hlock8 & ~n27004;
  assign n27006 = ~n13445 & ~n27003;
  assign n27007 = ~i_hlock8 & ~n27006;
  assign n27008 = ~n27005 & ~n27007;
  assign n27009 = controllable_hmaster3 & ~n27008;
  assign n27010 = ~n26942 & ~n27009;
  assign n27011 = i_hbusreq7 & ~n27010;
  assign n27012 = i_hbusreq8 & ~n27008;
  assign n27013 = controllable_hmaster0 & ~n13709;
  assign n27014 = ~n13570 & ~n27013;
  assign n27015 = i_hlock8 & ~n27014;
  assign n27016 = ~n13609 & ~n27013;
  assign n27017 = ~i_hlock8 & ~n27016;
  assign n27018 = ~n27015 & ~n27017;
  assign n27019 = ~i_hbusreq8 & ~n27018;
  assign n27020 = ~n27012 & ~n27019;
  assign n27021 = controllable_hmaster3 & ~n27020;
  assign n27022 = ~n26990 & ~n27021;
  assign n27023 = ~i_hbusreq7 & ~n27022;
  assign n27024 = ~n27011 & ~n27023;
  assign n27025 = n7924 & ~n27024;
  assign n27026 = ~n27002 & ~n27025;
  assign n27027 = n8214 & ~n27026;
  assign n27028 = ~n26996 & ~n27027;
  assign n27029 = ~n8202 & ~n27028;
  assign n27030 = ~n8988 & ~n26641;
  assign n27031 = controllable_hmaster1 & ~n27030;
  assign n27032 = ~n9096 & ~n27031;
  assign n27033 = ~controllable_hgrant6 & ~n27032;
  assign n27034 = ~n13673 & ~n27033;
  assign n27035 = controllable_hmaster0 & ~n27034;
  assign n27036 = ~n9099 & ~n27035;
  assign n27037 = ~controllable_hmaster3 & ~n27036;
  assign n27038 = ~n9093 & ~n27037;
  assign n27039 = i_hlock7 & ~n27038;
  assign n27040 = ~n8988 & ~n26656;
  assign n27041 = controllable_hmaster1 & ~n27040;
  assign n27042 = ~n9096 & ~n27041;
  assign n27043 = ~controllable_hgrant6 & ~n27042;
  assign n27044 = ~n13687 & ~n27043;
  assign n27045 = controllable_hmaster0 & ~n27044;
  assign n27046 = ~n9099 & ~n27045;
  assign n27047 = ~controllable_hmaster3 & ~n27046;
  assign n27048 = ~n9093 & ~n27047;
  assign n27049 = ~i_hlock7 & ~n27048;
  assign n27050 = ~n27039 & ~n27049;
  assign n27051 = i_hbusreq7 & ~n27050;
  assign n27052 = i_hbusreq8 & ~n27036;
  assign n27053 = i_hbusreq6 & ~n27032;
  assign n27054 = ~n9024 & ~n26684;
  assign n27055 = controllable_hmaster1 & ~n27054;
  assign n27056 = ~n9122 & ~n27055;
  assign n27057 = ~i_hbusreq6 & ~n27056;
  assign n27058 = ~n27053 & ~n27057;
  assign n27059 = ~controllable_hgrant6 & ~n27058;
  assign n27060 = ~n13716 & ~n27059;
  assign n27061 = controllable_hmaster0 & ~n27060;
  assign n27062 = ~n9127 & ~n27061;
  assign n27063 = ~i_hbusreq8 & ~n27062;
  assign n27064 = ~n27052 & ~n27063;
  assign n27065 = ~controllable_hmaster3 & ~n27064;
  assign n27066 = ~n9117 & ~n27065;
  assign n27067 = i_hlock7 & ~n27066;
  assign n27068 = i_hbusreq8 & ~n27046;
  assign n27069 = i_hbusreq6 & ~n27042;
  assign n27070 = ~n9024 & ~n26714;
  assign n27071 = controllable_hmaster1 & ~n27070;
  assign n27072 = ~n9122 & ~n27071;
  assign n27073 = ~i_hbusreq6 & ~n27072;
  assign n27074 = ~n27069 & ~n27073;
  assign n27075 = ~controllable_hgrant6 & ~n27074;
  assign n27076 = ~n13736 & ~n27075;
  assign n27077 = controllable_hmaster0 & ~n27076;
  assign n27078 = ~n9127 & ~n27077;
  assign n27079 = ~i_hbusreq8 & ~n27078;
  assign n27080 = ~n27068 & ~n27079;
  assign n27081 = ~controllable_hmaster3 & ~n27080;
  assign n27082 = ~n9117 & ~n27081;
  assign n27083 = ~i_hlock7 & ~n27082;
  assign n27084 = ~n27067 & ~n27083;
  assign n27085 = ~i_hbusreq7 & ~n27084;
  assign n27086 = ~n27051 & ~n27085;
  assign n27087 = ~n7924 & ~n27086;
  assign n27088 = controllable_hmaster3 & ~n13194;
  assign n27089 = ~n13189 & ~n26738;
  assign n27090 = controllable_hmaster1 & ~n27089;
  assign n27091 = ~n13677 & ~n27090;
  assign n27092 = ~controllable_hgrant6 & ~n27091;
  assign n27093 = ~n13673 & ~n27092;
  assign n27094 = controllable_hmaster0 & ~n27093;
  assign n27095 = ~n13682 & ~n27094;
  assign n27096 = ~controllable_hmaster3 & ~n27095;
  assign n27097 = ~n27088 & ~n27096;
  assign n27098 = i_hlock7 & ~n27097;
  assign n27099 = ~n13189 & ~n26754;
  assign n27100 = controllable_hmaster1 & ~n27099;
  assign n27101 = ~n13677 & ~n27100;
  assign n27102 = ~controllable_hgrant6 & ~n27101;
  assign n27103 = ~n13687 & ~n27102;
  assign n27104 = controllable_hmaster0 & ~n27103;
  assign n27105 = ~n13682 & ~n27104;
  assign n27106 = ~controllable_hmaster3 & ~n27105;
  assign n27107 = ~n27088 & ~n27106;
  assign n27108 = ~i_hlock7 & ~n27107;
  assign n27109 = ~n27098 & ~n27108;
  assign n27110 = i_hbusreq7 & ~n27109;
  assign n27111 = i_hbusreq8 & ~n13194;
  assign n27112 = ~i_hbusreq8 & ~n13291;
  assign n27113 = ~n27111 & ~n27112;
  assign n27114 = controllable_hmaster3 & ~n27113;
  assign n27115 = i_hbusreq8 & ~n27095;
  assign n27116 = i_hbusreq6 & ~n27091;
  assign n27117 = ~n13284 & ~n26783;
  assign n27118 = controllable_hmaster1 & ~n27117;
  assign n27119 = ~controllable_hmaster1 & ~n13283;
  assign n27120 = ~n27118 & ~n27119;
  assign n27121 = ~i_hbusreq6 & ~n27120;
  assign n27122 = ~n27116 & ~n27121;
  assign n27123 = ~controllable_hgrant6 & ~n27122;
  assign n27124 = ~n13716 & ~n27123;
  assign n27125 = controllable_hmaster0 & ~n27124;
  assign n27126 = ~controllable_hmaster0 & ~n13303;
  assign n27127 = ~n27125 & ~n27126;
  assign n27128 = ~i_hbusreq8 & ~n27127;
  assign n27129 = ~n27115 & ~n27128;
  assign n27130 = ~controllable_hmaster3 & ~n27129;
  assign n27131 = ~n27114 & ~n27130;
  assign n27132 = i_hlock7 & ~n27131;
  assign n27133 = i_hbusreq8 & ~n27105;
  assign n27134 = i_hbusreq6 & ~n27101;
  assign n27135 = ~n13284 & ~n26814;
  assign n27136 = controllable_hmaster1 & ~n27135;
  assign n27137 = ~n27119 & ~n27136;
  assign n27138 = ~i_hbusreq6 & ~n27137;
  assign n27139 = ~n27134 & ~n27138;
  assign n27140 = ~controllable_hgrant6 & ~n27139;
  assign n27141 = ~n13736 & ~n27140;
  assign n27142 = controllable_hmaster0 & ~n27141;
  assign n27143 = ~n27126 & ~n27142;
  assign n27144 = ~i_hbusreq8 & ~n27143;
  assign n27145 = ~n27133 & ~n27144;
  assign n27146 = ~controllable_hmaster3 & ~n27145;
  assign n27147 = ~n27114 & ~n27146;
  assign n27148 = ~i_hlock7 & ~n27147;
  assign n27149 = ~n27132 & ~n27148;
  assign n27150 = ~i_hbusreq7 & ~n27149;
  assign n27151 = ~n27110 & ~n27150;
  assign n27152 = n7924 & ~n27151;
  assign n27153 = ~n27087 & ~n27152;
  assign n27154 = ~n8214 & ~n27153;
  assign n27155 = ~n9156 & ~n26894;
  assign n27156 = ~controllable_hmaster3 & ~n27155;
  assign n27157 = ~n9093 & ~n27156;
  assign n27158 = i_hbusreq7 & ~n27157;
  assign n27159 = i_hbusreq8 & ~n27155;
  assign n27160 = ~n9169 & ~n26909;
  assign n27161 = ~i_hbusreq8 & ~n27160;
  assign n27162 = ~n27159 & ~n27161;
  assign n27163 = ~controllable_hmaster3 & ~n27162;
  assign n27164 = ~n9117 & ~n27163;
  assign n27165 = ~i_hbusreq7 & ~n27164;
  assign n27166 = ~n27158 & ~n27165;
  assign n27167 = ~n7924 & ~n27166;
  assign n27168 = ~n13772 & ~n26940;
  assign n27169 = ~controllable_hmaster3 & ~n27168;
  assign n27170 = ~n27088 & ~n27169;
  assign n27171 = i_hbusreq7 & ~n27170;
  assign n27172 = ~i_hbusreq8 & ~n13709;
  assign n27173 = ~n27111 & ~n27172;
  assign n27174 = controllable_hmaster3 & ~n27173;
  assign n27175 = i_hbusreq8 & ~n27168;
  assign n27176 = ~n13788 & ~n26986;
  assign n27177 = ~i_hbusreq8 & ~n27176;
  assign n27178 = ~n27175 & ~n27177;
  assign n27179 = ~controllable_hmaster3 & ~n27178;
  assign n27180 = ~n27174 & ~n27179;
  assign n27181 = ~i_hbusreq7 & ~n27180;
  assign n27182 = ~n27171 & ~n27181;
  assign n27183 = n7924 & ~n27182;
  assign n27184 = ~n27167 & ~n27183;
  assign n27185 = n8214 & ~n27184;
  assign n27186 = ~n27154 & ~n27185;
  assign n27187 = n8202 & ~n27186;
  assign n27188 = ~n27029 & ~n27187;
  assign n27189 = n7920 & ~n27188;
  assign n27190 = ~n8877 & ~n27189;
  assign n27191 = n7728 & ~n27190;
  assign n27192 = ~n9193 & ~n26641;
  assign n27193 = controllable_hmaster1 & ~n27192;
  assign n27194 = ~n9205 & ~n27193;
  assign n27195 = ~controllable_hgrant6 & ~n27194;
  assign n27196 = ~n13849 & ~n27195;
  assign n27197 = controllable_hmaster0 & ~n27196;
  assign n27198 = ~n9233 & ~n27197;
  assign n27199 = ~controllable_hmaster3 & ~n27198;
  assign n27200 = ~n9189 & ~n27199;
  assign n27201 = i_hlock7 & ~n27200;
  assign n27202 = ~n9193 & ~n26656;
  assign n27203 = controllable_hmaster1 & ~n27202;
  assign n27204 = ~n9205 & ~n27203;
  assign n27205 = ~controllable_hgrant6 & ~n27204;
  assign n27206 = ~n13951 & ~n27205;
  assign n27207 = controllable_hmaster0 & ~n27206;
  assign n27208 = ~n9233 & ~n27207;
  assign n27209 = ~controllable_hmaster3 & ~n27208;
  assign n27210 = ~n9189 & ~n27209;
  assign n27211 = ~i_hlock7 & ~n27210;
  assign n27212 = ~n27201 & ~n27211;
  assign n27213 = i_hbusreq7 & ~n27212;
  assign n27214 = i_hbusreq8 & ~n27198;
  assign n27215 = i_hbusreq6 & ~n27194;
  assign n27216 = ~i_hbusreq9 & ~n14332;
  assign n27217 = ~n26673 & ~n27216;
  assign n27218 = ~i_hbusreq4 & ~n27217;
  assign n27219 = ~n26672 & ~n27218;
  assign n27220 = ~controllable_hgrant4 & ~n27219;
  assign n27221 = ~n14021 & ~n27220;
  assign n27222 = ~i_hbusreq5 & ~n27221;
  assign n27223 = ~n26671 & ~n27222;
  assign n27224 = ~controllable_hgrant5 & ~n27223;
  assign n27225 = ~n14020 & ~n27224;
  assign n27226 = controllable_hmaster2 & ~n27225;
  assign n27227 = ~n9330 & ~n27226;
  assign n27228 = controllable_hmaster1 & ~n27227;
  assign n27229 = ~n9360 & ~n27228;
  assign n27230 = ~i_hbusreq6 & ~n27229;
  assign n27231 = ~n27215 & ~n27230;
  assign n27232 = ~controllable_hgrant6 & ~n27231;
  assign n27233 = ~n14094 & ~n27232;
  assign n27234 = controllable_hmaster0 & ~n27233;
  assign n27235 = ~n9439 & ~n27234;
  assign n27236 = ~i_hbusreq8 & ~n27235;
  assign n27237 = ~n27214 & ~n27236;
  assign n27238 = ~controllable_hmaster3 & ~n27237;
  assign n27239 = ~n9311 & ~n27238;
  assign n27240 = i_hlock7 & ~n27239;
  assign n27241 = i_hbusreq8 & ~n27208;
  assign n27242 = i_hbusreq6 & ~n27204;
  assign n27243 = ~i_hbusreq9 & ~n14342;
  assign n27244 = ~n26703 & ~n27243;
  assign n27245 = ~i_hbusreq4 & ~n27244;
  assign n27246 = ~n26702 & ~n27245;
  assign n27247 = ~controllable_hgrant4 & ~n27246;
  assign n27248 = ~n14056 & ~n27247;
  assign n27249 = ~i_hbusreq5 & ~n27248;
  assign n27250 = ~n26701 & ~n27249;
  assign n27251 = ~controllable_hgrant5 & ~n27250;
  assign n27252 = ~n14055 & ~n27251;
  assign n27253 = controllable_hmaster2 & ~n27252;
  assign n27254 = ~n9330 & ~n27253;
  assign n27255 = controllable_hmaster1 & ~n27254;
  assign n27256 = ~n9360 & ~n27255;
  assign n27257 = ~i_hbusreq6 & ~n27256;
  assign n27258 = ~n27242 & ~n27257;
  assign n27259 = ~controllable_hgrant6 & ~n27258;
  assign n27260 = ~n14298 & ~n27259;
  assign n27261 = controllable_hmaster0 & ~n27260;
  assign n27262 = ~n9439 & ~n27261;
  assign n27263 = ~i_hbusreq8 & ~n27262;
  assign n27264 = ~n27241 & ~n27263;
  assign n27265 = ~controllable_hmaster3 & ~n27264;
  assign n27266 = ~n9311 & ~n27265;
  assign n27267 = ~i_hlock7 & ~n27266;
  assign n27268 = ~n27240 & ~n27267;
  assign n27269 = ~i_hbusreq7 & ~n27268;
  assign n27270 = ~n27213 & ~n27269;
  assign n27271 = ~n7924 & ~n27270;
  assign n27272 = ~n13424 & ~n26931;
  assign n27273 = i_hlock8 & ~n27272;
  assign n27274 = ~n13445 & ~n26931;
  assign n27275 = ~i_hlock8 & ~n27274;
  assign n27276 = ~n27273 & ~n27275;
  assign n27277 = controllable_hmaster3 & ~n27276;
  assign n27278 = ~n13862 & ~n26738;
  assign n27279 = controllable_hmaster1 & ~n27278;
  assign n27280 = ~n13889 & ~n27279;
  assign n27281 = ~controllable_hgrant6 & ~n27280;
  assign n27282 = ~n13849 & ~n27281;
  assign n27283 = controllable_hmaster0 & ~n27282;
  assign n27284 = ~n13946 & ~n27283;
  assign n27285 = ~controllable_hmaster3 & ~n27284;
  assign n27286 = ~n27277 & ~n27285;
  assign n27287 = i_hlock7 & ~n27286;
  assign n27288 = ~n13862 & ~n26754;
  assign n27289 = controllable_hmaster1 & ~n27288;
  assign n27290 = ~n13889 & ~n27289;
  assign n27291 = ~controllable_hgrant6 & ~n27290;
  assign n27292 = ~n13951 & ~n27291;
  assign n27293 = controllable_hmaster0 & ~n27292;
  assign n27294 = ~n13946 & ~n27293;
  assign n27295 = ~controllable_hmaster3 & ~n27294;
  assign n27296 = ~n27277 & ~n27295;
  assign n27297 = ~i_hlock7 & ~n27296;
  assign n27298 = ~n27287 & ~n27297;
  assign n27299 = i_hbusreq7 & ~n27298;
  assign n27300 = i_hbusreq8 & ~n27276;
  assign n27301 = i_hlock9 & ~n14462;
  assign n27302 = ~i_hlock9 & ~n14493;
  assign n27303 = ~n27301 & ~n27302;
  assign n27304 = ~i_hbusreq9 & ~n27303;
  assign n27305 = ~n26949 & ~n27304;
  assign n27306 = ~i_hbusreq4 & ~n27305;
  assign n27307 = ~n26948 & ~n27306;
  assign n27308 = ~controllable_hgrant4 & ~n27307;
  assign n27309 = ~n12676 & ~n27308;
  assign n27310 = ~i_hbusreq5 & ~n27309;
  assign n27311 = ~n26947 & ~n27310;
  assign n27312 = ~controllable_hgrant5 & ~n27311;
  assign n27313 = ~n12674 & ~n27312;
  assign n27314 = ~controllable_hmaster2 & ~n27313;
  assign n27315 = ~n14401 & ~n27314;
  assign n27316 = ~controllable_hmaster1 & ~n27315;
  assign n27317 = ~n14400 & ~n27316;
  assign n27318 = ~i_hbusreq6 & ~n27317;
  assign n27319 = ~n26946 & ~n27318;
  assign n27320 = ~controllable_hgrant6 & ~n27319;
  assign n27321 = ~n13818 & ~n27320;
  assign n27322 = controllable_hmaster0 & ~n27321;
  assign n27323 = ~n14738 & ~n27322;
  assign n27324 = i_hlock8 & ~n27323;
  assign n27325 = ~n14749 & ~n27322;
  assign n27326 = ~i_hlock8 & ~n27325;
  assign n27327 = ~n27324 & ~n27326;
  assign n27328 = ~i_hbusreq8 & ~n27327;
  assign n27329 = ~n27300 & ~n27328;
  assign n27330 = controllable_hmaster3 & ~n27329;
  assign n27331 = i_hbusreq8 & ~n27284;
  assign n27332 = i_hbusreq6 & ~n27280;
  assign n27333 = ~i_hbusreq9 & ~n14411;
  assign n27334 = ~n26772 & ~n27333;
  assign n27335 = ~i_hbusreq4 & ~n27334;
  assign n27336 = ~n26771 & ~n27335;
  assign n27337 = ~controllable_hgrant4 & ~n27336;
  assign n27338 = ~n14021 & ~n27337;
  assign n27339 = ~i_hbusreq5 & ~n27338;
  assign n27340 = ~n26770 & ~n27339;
  assign n27341 = ~controllable_hgrant5 & ~n27340;
  assign n27342 = ~n14020 & ~n27341;
  assign n27343 = controllable_hmaster2 & ~n27342;
  assign n27344 = ~n14561 & ~n27343;
  assign n27345 = controllable_hmaster1 & ~n27344;
  assign n27346 = ~n14605 & ~n27345;
  assign n27347 = ~i_hbusreq6 & ~n27346;
  assign n27348 = ~n27332 & ~n27347;
  assign n27349 = ~controllable_hgrant6 & ~n27348;
  assign n27350 = ~n14094 & ~n27349;
  assign n27351 = controllable_hmaster0 & ~n27350;
  assign n27352 = ~n14685 & ~n27351;
  assign n27353 = ~i_hbusreq8 & ~n27352;
  assign n27354 = ~n27331 & ~n27353;
  assign n27355 = ~controllable_hmaster3 & ~n27354;
  assign n27356 = ~n27330 & ~n27355;
  assign n27357 = i_hlock7 & ~n27356;
  assign n27358 = i_hbusreq8 & ~n27294;
  assign n27359 = i_hbusreq6 & ~n27290;
  assign n27360 = ~i_hbusreq9 & ~n14421;
  assign n27361 = ~n26803 & ~n27360;
  assign n27362 = ~i_hbusreq4 & ~n27361;
  assign n27363 = ~n26802 & ~n27362;
  assign n27364 = ~controllable_hgrant4 & ~n27363;
  assign n27365 = ~n14056 & ~n27364;
  assign n27366 = ~i_hbusreq5 & ~n27365;
  assign n27367 = ~n26801 & ~n27366;
  assign n27368 = ~controllable_hgrant5 & ~n27367;
  assign n27369 = ~n14055 & ~n27368;
  assign n27370 = controllable_hmaster2 & ~n27369;
  assign n27371 = ~n14561 & ~n27370;
  assign n27372 = controllable_hmaster1 & ~n27371;
  assign n27373 = ~n14605 & ~n27372;
  assign n27374 = ~i_hbusreq6 & ~n27373;
  assign n27375 = ~n27359 & ~n27374;
  assign n27376 = ~controllable_hgrant6 & ~n27375;
  assign n27377 = ~n14298 & ~n27376;
  assign n27378 = controllable_hmaster0 & ~n27377;
  assign n27379 = ~n14685 & ~n27378;
  assign n27380 = ~i_hbusreq8 & ~n27379;
  assign n27381 = ~n27358 & ~n27380;
  assign n27382 = ~controllable_hmaster3 & ~n27381;
  assign n27383 = ~n27330 & ~n27382;
  assign n27384 = ~i_hlock7 & ~n27383;
  assign n27385 = ~n27357 & ~n27384;
  assign n27386 = ~i_hbusreq7 & ~n27385;
  assign n27387 = ~n27299 & ~n27386;
  assign n27388 = n7924 & ~n27387;
  assign n27389 = ~n27271 & ~n27388;
  assign n27390 = ~n8214 & ~n27389;
  assign n27391 = ~n9499 & ~n27238;
  assign n27392 = i_hlock7 & ~n27391;
  assign n27393 = ~n9499 & ~n27265;
  assign n27394 = ~i_hlock7 & ~n27393;
  assign n27395 = ~n27392 & ~n27394;
  assign n27396 = ~i_hbusreq7 & ~n27395;
  assign n27397 = ~n27213 & ~n27396;
  assign n27398 = ~n7924 & ~n27397;
  assign n27399 = i_hlock9 & ~n14527;
  assign n27400 = ~i_hlock9 & ~n14568;
  assign n27401 = ~n27399 & ~n27400;
  assign n27402 = ~i_hbusreq9 & ~n27401;
  assign n27403 = ~n26949 & ~n27402;
  assign n27404 = ~i_hbusreq4 & ~n27403;
  assign n27405 = ~n26948 & ~n27404;
  assign n27406 = ~controllable_hgrant4 & ~n27405;
  assign n27407 = ~n14322 & ~n27406;
  assign n27408 = ~i_hbusreq5 & ~n27407;
  assign n27409 = ~n26947 & ~n27408;
  assign n27410 = ~controllable_hgrant5 & ~n27409;
  assign n27411 = ~n14321 & ~n27410;
  assign n27412 = ~controllable_hmaster2 & ~n27411;
  assign n27413 = ~n14401 & ~n27412;
  assign n27414 = ~controllable_hmaster1 & ~n27413;
  assign n27415 = ~n14400 & ~n27414;
  assign n27416 = ~i_hbusreq6 & ~n27415;
  assign n27417 = ~n26946 & ~n27416;
  assign n27418 = ~controllable_hgrant6 & ~n27417;
  assign n27419 = ~n14320 & ~n27418;
  assign n27420 = controllable_hmaster0 & ~n27419;
  assign n27421 = ~n14481 & ~n27420;
  assign n27422 = i_hlock8 & ~n27421;
  assign n27423 = ~n14512 & ~n27420;
  assign n27424 = ~i_hlock8 & ~n27423;
  assign n27425 = ~n27422 & ~n27424;
  assign n27426 = ~i_hbusreq8 & ~n27425;
  assign n27427 = ~n27300 & ~n27426;
  assign n27428 = controllable_hmaster3 & ~n27427;
  assign n27429 = ~n27355 & ~n27428;
  assign n27430 = i_hlock7 & ~n27429;
  assign n27431 = ~n27382 & ~n27428;
  assign n27432 = ~i_hlock7 & ~n27431;
  assign n27433 = ~n27430 & ~n27432;
  assign n27434 = ~i_hbusreq7 & ~n27433;
  assign n27435 = ~n27299 & ~n27434;
  assign n27436 = n7924 & ~n27435;
  assign n27437 = ~n27398 & ~n27436;
  assign n27438 = n8214 & ~n27437;
  assign n27439 = ~n27390 & ~n27438;
  assign n27440 = ~n8202 & ~n27439;
  assign n27441 = ~n9330 & ~n26684;
  assign n27442 = controllable_hmaster1 & ~n27441;
  assign n27443 = ~n9360 & ~n27442;
  assign n27444 = ~i_hbusreq6 & ~n27443;
  assign n27445 = ~n27215 & ~n27444;
  assign n27446 = ~controllable_hgrant6 & ~n27445;
  assign n27447 = ~n14756 & ~n27446;
  assign n27448 = controllable_hmaster0 & ~n27447;
  assign n27449 = ~n9439 & ~n27448;
  assign n27450 = ~i_hbusreq8 & ~n27449;
  assign n27451 = ~n27214 & ~n27450;
  assign n27452 = ~controllable_hmaster3 & ~n27451;
  assign n27453 = ~n9517 & ~n27452;
  assign n27454 = i_hlock7 & ~n27453;
  assign n27455 = ~n9330 & ~n26714;
  assign n27456 = controllable_hmaster1 & ~n27455;
  assign n27457 = ~n9360 & ~n27456;
  assign n27458 = ~i_hbusreq6 & ~n27457;
  assign n27459 = ~n27242 & ~n27458;
  assign n27460 = ~controllable_hgrant6 & ~n27459;
  assign n27461 = ~n14772 & ~n27460;
  assign n27462 = controllable_hmaster0 & ~n27461;
  assign n27463 = ~n9439 & ~n27462;
  assign n27464 = ~i_hbusreq8 & ~n27463;
  assign n27465 = ~n27241 & ~n27464;
  assign n27466 = ~controllable_hmaster3 & ~n27465;
  assign n27467 = ~n9517 & ~n27466;
  assign n27468 = ~i_hlock7 & ~n27467;
  assign n27469 = ~n27454 & ~n27468;
  assign n27470 = ~i_hbusreq7 & ~n27469;
  assign n27471 = ~n27213 & ~n27470;
  assign n27472 = ~n7924 & ~n27471;
  assign n27473 = i_hlock9 & ~n14032;
  assign n27474 = ~i_hlock9 & ~n14067;
  assign n27475 = ~n27473 & ~n27474;
  assign n27476 = ~i_hbusreq9 & ~n27475;
  assign n27477 = ~n26949 & ~n27476;
  assign n27478 = ~i_hbusreq4 & ~n27477;
  assign n27479 = ~n26948 & ~n27478;
  assign n27480 = ~controllable_hgrant4 & ~n27479;
  assign n27481 = ~n14322 & ~n27480;
  assign n27482 = ~i_hbusreq5 & ~n27481;
  assign n27483 = ~n26947 & ~n27482;
  assign n27484 = ~controllable_hgrant5 & ~n27483;
  assign n27485 = ~n14321 & ~n27484;
  assign n27486 = ~controllable_hmaster2 & ~n27485;
  assign n27487 = ~n14010 & ~n27486;
  assign n27488 = ~controllable_hmaster1 & ~n27487;
  assign n27489 = ~n14009 & ~n27488;
  assign n27490 = ~i_hbusreq6 & ~n27489;
  assign n27491 = ~n26946 & ~n27490;
  assign n27492 = ~controllable_hgrant6 & ~n27491;
  assign n27493 = ~n14320 & ~n27492;
  assign n27494 = controllable_hmaster0 & ~n27493;
  assign n27495 = ~n14051 & ~n27494;
  assign n27496 = i_hlock8 & ~n27495;
  assign n27497 = ~n14086 & ~n27494;
  assign n27498 = ~i_hlock8 & ~n27497;
  assign n27499 = ~n27496 & ~n27498;
  assign n27500 = ~i_hbusreq8 & ~n27499;
  assign n27501 = ~n27300 & ~n27500;
  assign n27502 = controllable_hmaster3 & ~n27501;
  assign n27503 = ~n14121 & ~n26783;
  assign n27504 = controllable_hmaster1 & ~n27503;
  assign n27505 = ~n14166 & ~n27504;
  assign n27506 = ~i_hbusreq6 & ~n27505;
  assign n27507 = ~n27332 & ~n27506;
  assign n27508 = ~controllable_hgrant6 & ~n27507;
  assign n27509 = ~n14756 & ~n27508;
  assign n27510 = controllable_hmaster0 & ~n27509;
  assign n27511 = ~n14290 & ~n27510;
  assign n27512 = ~i_hbusreq8 & ~n27511;
  assign n27513 = ~n27331 & ~n27512;
  assign n27514 = ~controllable_hmaster3 & ~n27513;
  assign n27515 = ~n27502 & ~n27514;
  assign n27516 = i_hlock7 & ~n27515;
  assign n27517 = ~n14121 & ~n26814;
  assign n27518 = controllable_hmaster1 & ~n27517;
  assign n27519 = ~n14166 & ~n27518;
  assign n27520 = ~i_hbusreq6 & ~n27519;
  assign n27521 = ~n27359 & ~n27520;
  assign n27522 = ~controllable_hgrant6 & ~n27521;
  assign n27523 = ~n14772 & ~n27522;
  assign n27524 = controllable_hmaster0 & ~n27523;
  assign n27525 = ~n14290 & ~n27524;
  assign n27526 = ~i_hbusreq8 & ~n27525;
  assign n27527 = ~n27358 & ~n27526;
  assign n27528 = ~controllable_hmaster3 & ~n27527;
  assign n27529 = ~n27502 & ~n27528;
  assign n27530 = ~i_hlock7 & ~n27529;
  assign n27531 = ~n27516 & ~n27530;
  assign n27532 = ~i_hbusreq7 & ~n27531;
  assign n27533 = ~n27299 & ~n27532;
  assign n27534 = n7924 & ~n27533;
  assign n27535 = ~n27472 & ~n27534;
  assign n27536 = ~n8214 & ~n27535;
  assign n27537 = ~n9557 & ~n27234;
  assign n27538 = ~i_hbusreq8 & ~n27537;
  assign n27539 = ~n27214 & ~n27538;
  assign n27540 = ~controllable_hmaster3 & ~n27539;
  assign n27541 = ~n9517 & ~n27540;
  assign n27542 = i_hlock7 & ~n27541;
  assign n27543 = ~n9557 & ~n27261;
  assign n27544 = ~i_hbusreq8 & ~n27543;
  assign n27545 = ~n27241 & ~n27544;
  assign n27546 = ~controllable_hmaster3 & ~n27545;
  assign n27547 = ~n9517 & ~n27546;
  assign n27548 = ~i_hlock7 & ~n27547;
  assign n27549 = ~n27542 & ~n27548;
  assign n27550 = ~i_hbusreq7 & ~n27549;
  assign n27551 = ~n27213 & ~n27550;
  assign n27552 = ~n7924 & ~n27551;
  assign n27553 = ~n14738 & ~n27420;
  assign n27554 = i_hlock8 & ~n27553;
  assign n27555 = ~n14749 & ~n27420;
  assign n27556 = ~i_hlock8 & ~n27555;
  assign n27557 = ~n27554 & ~n27556;
  assign n27558 = ~i_hbusreq8 & ~n27557;
  assign n27559 = ~n27300 & ~n27558;
  assign n27560 = controllable_hmaster3 & ~n27559;
  assign n27561 = ~n14816 & ~n27351;
  assign n27562 = ~i_hbusreq8 & ~n27561;
  assign n27563 = ~n27331 & ~n27562;
  assign n27564 = ~controllable_hmaster3 & ~n27563;
  assign n27565 = ~n27560 & ~n27564;
  assign n27566 = i_hlock7 & ~n27565;
  assign n27567 = ~n14816 & ~n27378;
  assign n27568 = ~i_hbusreq8 & ~n27567;
  assign n27569 = ~n27358 & ~n27568;
  assign n27570 = ~controllable_hmaster3 & ~n27569;
  assign n27571 = ~n27560 & ~n27570;
  assign n27572 = ~i_hlock7 & ~n27571;
  assign n27573 = ~n27566 & ~n27572;
  assign n27574 = ~i_hbusreq7 & ~n27573;
  assign n27575 = ~n27299 & ~n27574;
  assign n27576 = n7924 & ~n27575;
  assign n27577 = ~n27552 & ~n27576;
  assign n27578 = n8214 & ~n27577;
  assign n27579 = ~n27536 & ~n27578;
  assign n27580 = n8202 & ~n27579;
  assign n27581 = ~n27440 & ~n27580;
  assign n27582 = n7920 & ~n27581;
  assign n27583 = ~n8877 & ~n27582;
  assign n27584 = ~n7728 & ~n27583;
  assign n27585 = ~n27191 & ~n27584;
  assign n27586 = n7723 & ~n27585;
  assign n27587 = ~n7723 & ~n27583;
  assign n27588 = ~n27586 & ~n27587;
  assign n27589 = n7714 & ~n27588;
  assign n27590 = n7723 & ~n27583;
  assign n27591 = ~n8640 & ~n27582;
  assign n27592 = n7728 & ~n27591;
  assign n27593 = ~n9638 & ~n26684;
  assign n27594 = controllable_hmaster1 & ~n27593;
  assign n27595 = ~n9662 & ~n27594;
  assign n27596 = ~i_hbusreq6 & ~n27595;
  assign n27597 = ~n27215 & ~n27596;
  assign n27598 = ~controllable_hgrant6 & ~n27597;
  assign n27599 = ~n14995 & ~n27598;
  assign n27600 = controllable_hmaster0 & ~n27599;
  assign n27601 = ~n9716 & ~n27600;
  assign n27602 = ~i_hbusreq8 & ~n27601;
  assign n27603 = ~n27214 & ~n27602;
  assign n27604 = ~controllable_hmaster3 & ~n27603;
  assign n27605 = ~n9626 & ~n27604;
  assign n27606 = i_hlock7 & ~n27605;
  assign n27607 = ~n9638 & ~n26714;
  assign n27608 = controllable_hmaster1 & ~n27607;
  assign n27609 = ~n9662 & ~n27608;
  assign n27610 = ~i_hbusreq6 & ~n27609;
  assign n27611 = ~n27242 & ~n27610;
  assign n27612 = ~controllable_hgrant6 & ~n27611;
  assign n27613 = ~n15152 & ~n27612;
  assign n27614 = controllable_hmaster0 & ~n27613;
  assign n27615 = ~n9716 & ~n27614;
  assign n27616 = ~i_hbusreq8 & ~n27615;
  assign n27617 = ~n27241 & ~n27616;
  assign n27618 = ~controllable_hmaster3 & ~n27617;
  assign n27619 = ~n9626 & ~n27618;
  assign n27620 = ~i_hlock7 & ~n27619;
  assign n27621 = ~n27606 & ~n27620;
  assign n27622 = ~i_hbusreq7 & ~n27621;
  assign n27623 = ~n27213 & ~n27622;
  assign n27624 = ~n7924 & ~n27623;
  assign n27625 = i_hlock9 & ~n14938;
  assign n27626 = ~i_hlock9 & ~n14969;
  assign n27627 = ~n27625 & ~n27626;
  assign n27628 = ~i_hbusreq9 & ~n27627;
  assign n27629 = ~n26949 & ~n27628;
  assign n27630 = ~i_hbusreq4 & ~n27629;
  assign n27631 = ~n26948 & ~n27630;
  assign n27632 = ~controllable_hgrant4 & ~n27631;
  assign n27633 = ~n12676 & ~n27632;
  assign n27634 = ~i_hbusreq5 & ~n27633;
  assign n27635 = ~n26947 & ~n27634;
  assign n27636 = ~controllable_hgrant5 & ~n27635;
  assign n27637 = ~n12674 & ~n27636;
  assign n27638 = ~controllable_hmaster2 & ~n27637;
  assign n27639 = ~n14918 & ~n27638;
  assign n27640 = ~controllable_hmaster1 & ~n27639;
  assign n27641 = ~n14917 & ~n27640;
  assign n27642 = ~i_hbusreq6 & ~n27641;
  assign n27643 = ~n26946 & ~n27642;
  assign n27644 = ~controllable_hgrant6 & ~n27643;
  assign n27645 = ~n14849 & ~n27644;
  assign n27646 = controllable_hmaster0 & ~n27645;
  assign n27647 = ~n14957 & ~n27646;
  assign n27648 = i_hlock8 & ~n27647;
  assign n27649 = ~n14988 & ~n27646;
  assign n27650 = ~i_hlock8 & ~n27649;
  assign n27651 = ~n27648 & ~n27650;
  assign n27652 = ~i_hbusreq8 & ~n27651;
  assign n27653 = ~n27300 & ~n27652;
  assign n27654 = controllable_hmaster3 & ~n27653;
  assign n27655 = ~n15017 & ~n26783;
  assign n27656 = controllable_hmaster1 & ~n27655;
  assign n27657 = ~n15056 & ~n27656;
  assign n27658 = ~i_hbusreq6 & ~n27657;
  assign n27659 = ~n27332 & ~n27658;
  assign n27660 = ~controllable_hgrant6 & ~n27659;
  assign n27661 = ~n14995 & ~n27660;
  assign n27662 = controllable_hmaster0 & ~n27661;
  assign n27663 = ~n15145 & ~n27662;
  assign n27664 = ~i_hbusreq8 & ~n27663;
  assign n27665 = ~n27331 & ~n27664;
  assign n27666 = ~controllable_hmaster3 & ~n27665;
  assign n27667 = ~n27654 & ~n27666;
  assign n27668 = i_hlock7 & ~n27667;
  assign n27669 = ~n15017 & ~n26814;
  assign n27670 = controllable_hmaster1 & ~n27669;
  assign n27671 = ~n15056 & ~n27670;
  assign n27672 = ~i_hbusreq6 & ~n27671;
  assign n27673 = ~n27359 & ~n27672;
  assign n27674 = ~controllable_hgrant6 & ~n27673;
  assign n27675 = ~n15152 & ~n27674;
  assign n27676 = controllable_hmaster0 & ~n27675;
  assign n27677 = ~n15145 & ~n27676;
  assign n27678 = ~i_hbusreq8 & ~n27677;
  assign n27679 = ~n27358 & ~n27678;
  assign n27680 = ~controllable_hmaster3 & ~n27679;
  assign n27681 = ~n27654 & ~n27680;
  assign n27682 = ~i_hlock7 & ~n27681;
  assign n27683 = ~n27668 & ~n27682;
  assign n27684 = ~i_hbusreq7 & ~n27683;
  assign n27685 = ~n27299 & ~n27684;
  assign n27686 = n7924 & ~n27685;
  assign n27687 = ~n27624 & ~n27686;
  assign n27688 = n7920 & ~n27687;
  assign n27689 = ~n8640 & ~n27688;
  assign n27690 = ~n7728 & ~n27689;
  assign n27691 = ~n27592 & ~n27690;
  assign n27692 = ~n7723 & ~n27691;
  assign n27693 = ~n27590 & ~n27692;
  assign n27694 = ~n7714 & ~n27693;
  assign n27695 = ~n27589 & ~n27694;
  assign n27696 = ~n7705 & ~n27695;
  assign n27697 = ~n26887 & ~n27696;
  assign n27698 = n7808 & ~n27697;
  assign n27699 = ~n8650 & ~n27698;
  assign n27700 = n8195 & ~n27699;
  assign n27701 = ~n8196 & ~n27700;
  assign n27702 = ~n8193 & ~n27701;
  assign n27703 = ~n10055 & ~n26890;
  assign n27704 = ~controllable_hgrant6 & ~n27703;
  assign n27705 = ~n15193 & ~n27704;
  assign n27706 = controllable_hmaster0 & ~n27705;
  assign n27707 = ~n9099 & ~n27706;
  assign n27708 = ~controllable_hmaster3 & ~n27707;
  assign n27709 = ~n9093 & ~n27708;
  assign n27710 = i_hbusreq7 & ~n27709;
  assign n27711 = i_hbusreq8 & ~n27707;
  assign n27712 = i_hbusreq6 & ~n27703;
  assign n27713 = ~n10066 & ~n26903;
  assign n27714 = ~i_hbusreq6 & ~n27713;
  assign n27715 = ~n27712 & ~n27714;
  assign n27716 = ~controllable_hgrant6 & ~n27715;
  assign n27717 = ~n15206 & ~n27716;
  assign n27718 = controllable_hmaster0 & ~n27717;
  assign n27719 = ~n9127 & ~n27718;
  assign n27720 = ~i_hbusreq8 & ~n27719;
  assign n27721 = ~n27711 & ~n27720;
  assign n27722 = ~controllable_hmaster3 & ~n27721;
  assign n27723 = ~n9117 & ~n27722;
  assign n27724 = ~i_hbusreq7 & ~n27723;
  assign n27725 = ~n27710 & ~n27724;
  assign n27726 = ~n7924 & ~n27725;
  assign n27727 = ~n15196 & ~n26936;
  assign n27728 = ~controllable_hgrant6 & ~n27727;
  assign n27729 = ~n15193 & ~n27728;
  assign n27730 = controllable_hmaster0 & ~n27729;
  assign n27731 = ~n13682 & ~n27730;
  assign n27732 = ~controllable_hmaster3 & ~n27731;
  assign n27733 = ~n27088 & ~n27732;
  assign n27734 = i_hbusreq7 & ~n27733;
  assign n27735 = i_hbusreq8 & ~n27731;
  assign n27736 = i_hbusreq6 & ~n27727;
  assign n27737 = ~n15218 & ~n26980;
  assign n27738 = ~i_hbusreq6 & ~n27737;
  assign n27739 = ~n27736 & ~n27738;
  assign n27740 = ~controllable_hgrant6 & ~n27739;
  assign n27741 = ~n15206 & ~n27740;
  assign n27742 = controllable_hmaster0 & ~n27741;
  assign n27743 = ~n13728 & ~n27742;
  assign n27744 = ~i_hbusreq8 & ~n27743;
  assign n27745 = ~n27735 & ~n27744;
  assign n27746 = ~controllable_hmaster3 & ~n27745;
  assign n27747 = ~n27174 & ~n27746;
  assign n27748 = ~i_hbusreq7 & ~n27747;
  assign n27749 = ~n27734 & ~n27748;
  assign n27750 = n7924 & ~n27749;
  assign n27751 = ~n27726 & ~n27750;
  assign n27752 = ~n8214 & ~n27751;
  assign n27753 = ~n10082 & ~n26894;
  assign n27754 = ~controllable_hmaster3 & ~n27753;
  assign n27755 = ~n9093 & ~n27754;
  assign n27756 = i_hbusreq7 & ~n27755;
  assign n27757 = i_hbusreq8 & ~n27753;
  assign n27758 = ~n10094 & ~n26909;
  assign n27759 = ~i_hbusreq8 & ~n27758;
  assign n27760 = ~n27757 & ~n27759;
  assign n27761 = ~controllable_hmaster3 & ~n27760;
  assign n27762 = ~n9117 & ~n27761;
  assign n27763 = ~i_hbusreq7 & ~n27762;
  assign n27764 = ~n27756 & ~n27763;
  assign n27765 = ~n7924 & ~n27764;
  assign n27766 = ~n15247 & ~n26940;
  assign n27767 = ~controllable_hmaster3 & ~n27766;
  assign n27768 = ~n27088 & ~n27767;
  assign n27769 = i_hbusreq7 & ~n27768;
  assign n27770 = i_hbusreq8 & ~n27766;
  assign n27771 = ~n15274 & ~n26986;
  assign n27772 = ~i_hbusreq8 & ~n27771;
  assign n27773 = ~n27770 & ~n27772;
  assign n27774 = ~controllable_hmaster3 & ~n27773;
  assign n27775 = ~n27174 & ~n27774;
  assign n27776 = ~i_hbusreq7 & ~n27775;
  assign n27777 = ~n27769 & ~n27776;
  assign n27778 = n7924 & ~n27777;
  assign n27779 = ~n27765 & ~n27778;
  assign n27780 = n8214 & ~n27779;
  assign n27781 = ~n27752 & ~n27780;
  assign n27782 = ~n8202 & ~n27781;
  assign n27783 = ~n9193 & ~n26888;
  assign n27784 = controllable_hmaster1 & ~n27783;
  assign n27785 = ~n9096 & ~n27784;
  assign n27786 = ~controllable_hgrant6 & ~n27785;
  assign n27787 = ~n15293 & ~n27786;
  assign n27788 = controllable_hmaster0 & ~n27787;
  assign n27789 = ~n9099 & ~n27788;
  assign n27790 = ~controllable_hmaster3 & ~n27789;
  assign n27791 = ~n9093 & ~n27790;
  assign n27792 = i_hbusreq7 & ~n27791;
  assign n27793 = i_hbusreq8 & ~n27789;
  assign n27794 = i_hbusreq6 & ~n27785;
  assign n27795 = ~n9638 & ~n26901;
  assign n27796 = controllable_hmaster1 & ~n27795;
  assign n27797 = ~n9122 & ~n27796;
  assign n27798 = ~i_hbusreq6 & ~n27797;
  assign n27799 = ~n27794 & ~n27798;
  assign n27800 = ~controllable_hgrant6 & ~n27799;
  assign n27801 = ~n15306 & ~n27800;
  assign n27802 = controllable_hmaster0 & ~n27801;
  assign n27803 = ~n9127 & ~n27802;
  assign n27804 = ~i_hbusreq8 & ~n27803;
  assign n27805 = ~n27793 & ~n27804;
  assign n27806 = ~controllable_hmaster3 & ~n27805;
  assign n27807 = ~n9117 & ~n27806;
  assign n27808 = ~i_hbusreq7 & ~n27807;
  assign n27809 = ~n27792 & ~n27808;
  assign n27810 = ~n7924 & ~n27809;
  assign n27811 = ~n13862 & ~n26934;
  assign n27812 = controllable_hmaster1 & ~n27811;
  assign n27813 = ~n13677 & ~n27812;
  assign n27814 = ~controllable_hgrant6 & ~n27813;
  assign n27815 = ~n15293 & ~n27814;
  assign n27816 = controllable_hmaster0 & ~n27815;
  assign n27817 = ~n13682 & ~n27816;
  assign n27818 = ~controllable_hmaster3 & ~n27817;
  assign n27819 = ~n27088 & ~n27818;
  assign n27820 = i_hbusreq7 & ~n27819;
  assign n27821 = i_hbusreq8 & ~n27817;
  assign n27822 = i_hbusreq6 & ~n27813;
  assign n27823 = ~n15326 & ~n26978;
  assign n27824 = controllable_hmaster1 & ~n27823;
  assign n27825 = ~n13721 & ~n27824;
  assign n27826 = ~i_hbusreq6 & ~n27825;
  assign n27827 = ~n27822 & ~n27826;
  assign n27828 = ~controllable_hgrant6 & ~n27827;
  assign n27829 = ~n15306 & ~n27828;
  assign n27830 = controllable_hmaster0 & ~n27829;
  assign n27831 = ~n13728 & ~n27830;
  assign n27832 = ~i_hbusreq8 & ~n27831;
  assign n27833 = ~n27821 & ~n27832;
  assign n27834 = ~controllable_hmaster3 & ~n27833;
  assign n27835 = ~n27174 & ~n27834;
  assign n27836 = ~i_hbusreq7 & ~n27835;
  assign n27837 = ~n27820 & ~n27836;
  assign n27838 = n7924 & ~n27837;
  assign n27839 = ~n27810 & ~n27838;
  assign n27840 = ~n8214 & ~n27839;
  assign n27841 = ~n10134 & ~n26894;
  assign n27842 = ~controllable_hmaster3 & ~n27841;
  assign n27843 = ~n9093 & ~n27842;
  assign n27844 = i_hbusreq7 & ~n27843;
  assign n27845 = i_hbusreq8 & ~n27841;
  assign n27846 = ~n10146 & ~n26909;
  assign n27847 = ~i_hbusreq8 & ~n27846;
  assign n27848 = ~n27845 & ~n27847;
  assign n27849 = ~controllable_hmaster3 & ~n27848;
  assign n27850 = ~n9117 & ~n27849;
  assign n27851 = ~i_hbusreq7 & ~n27850;
  assign n27852 = ~n27844 & ~n27851;
  assign n27853 = ~n7924 & ~n27852;
  assign n27854 = ~n15357 & ~n26940;
  assign n27855 = ~controllable_hmaster3 & ~n27854;
  assign n27856 = ~n27088 & ~n27855;
  assign n27857 = i_hbusreq7 & ~n27856;
  assign n27858 = i_hbusreq8 & ~n27854;
  assign n27859 = ~n15392 & ~n26986;
  assign n27860 = ~i_hbusreq8 & ~n27859;
  assign n27861 = ~n27858 & ~n27860;
  assign n27862 = ~controllable_hmaster3 & ~n27861;
  assign n27863 = ~n27174 & ~n27862;
  assign n27864 = ~i_hbusreq7 & ~n27863;
  assign n27865 = ~n27857 & ~n27864;
  assign n27866 = n7924 & ~n27865;
  assign n27867 = ~n27853 & ~n27866;
  assign n27868 = n8214 & ~n27867;
  assign n27869 = ~n27840 & ~n27868;
  assign n27870 = n8202 & ~n27869;
  assign n27871 = ~n27782 & ~n27870;
  assign n27872 = n7920 & ~n27871;
  assign n27873 = ~n10014 & ~n27872;
  assign n27874 = n7728 & ~n27873;
  assign n27875 = ~n10162 & ~n27228;
  assign n27876 = ~i_hbusreq6 & ~n27875;
  assign n27877 = ~n27215 & ~n27876;
  assign n27878 = ~controllable_hgrant6 & ~n27877;
  assign n27879 = ~n15417 & ~n27878;
  assign n27880 = controllable_hmaster0 & ~n27879;
  assign n27881 = ~n9439 & ~n27880;
  assign n27882 = ~i_hbusreq8 & ~n27881;
  assign n27883 = ~n27214 & ~n27882;
  assign n27884 = ~controllable_hmaster3 & ~n27883;
  assign n27885 = ~n9517 & ~n27884;
  assign n27886 = i_hlock7 & ~n27885;
  assign n27887 = ~n10162 & ~n27255;
  assign n27888 = ~i_hbusreq6 & ~n27887;
  assign n27889 = ~n27242 & ~n27888;
  assign n27890 = ~controllable_hgrant6 & ~n27889;
  assign n27891 = ~n15440 & ~n27890;
  assign n27892 = controllable_hmaster0 & ~n27891;
  assign n27893 = ~n9439 & ~n27892;
  assign n27894 = ~i_hbusreq8 & ~n27893;
  assign n27895 = ~n27241 & ~n27894;
  assign n27896 = ~controllable_hmaster3 & ~n27895;
  assign n27897 = ~n9517 & ~n27896;
  assign n27898 = ~i_hlock7 & ~n27897;
  assign n27899 = ~n27886 & ~n27898;
  assign n27900 = ~i_hbusreq7 & ~n27899;
  assign n27901 = ~n27213 & ~n27900;
  assign n27902 = ~n7924 & ~n27901;
  assign n27903 = ~n15427 & ~n27345;
  assign n27904 = ~i_hbusreq6 & ~n27903;
  assign n27905 = ~n27332 & ~n27904;
  assign n27906 = ~controllable_hgrant6 & ~n27905;
  assign n27907 = ~n15417 & ~n27906;
  assign n27908 = controllable_hmaster0 & ~n27907;
  assign n27909 = ~n14685 & ~n27908;
  assign n27910 = ~i_hbusreq8 & ~n27909;
  assign n27911 = ~n27331 & ~n27910;
  assign n27912 = ~controllable_hmaster3 & ~n27911;
  assign n27913 = ~n27560 & ~n27912;
  assign n27914 = i_hlock7 & ~n27913;
  assign n27915 = ~n15427 & ~n27372;
  assign n27916 = ~i_hbusreq6 & ~n27915;
  assign n27917 = ~n27359 & ~n27916;
  assign n27918 = ~controllable_hgrant6 & ~n27917;
  assign n27919 = ~n15440 & ~n27918;
  assign n27920 = controllable_hmaster0 & ~n27919;
  assign n27921 = ~n14685 & ~n27920;
  assign n27922 = ~i_hbusreq8 & ~n27921;
  assign n27923 = ~n27358 & ~n27922;
  assign n27924 = ~controllable_hmaster3 & ~n27923;
  assign n27925 = ~n27560 & ~n27924;
  assign n27926 = ~i_hlock7 & ~n27925;
  assign n27927 = ~n27914 & ~n27926;
  assign n27928 = ~i_hbusreq7 & ~n27927;
  assign n27929 = ~n27299 & ~n27928;
  assign n27930 = n7924 & ~n27929;
  assign n27931 = ~n27902 & ~n27930;
  assign n27932 = ~n8214 & ~n27931;
  assign n27933 = ~n10196 & ~n27234;
  assign n27934 = ~i_hbusreq8 & ~n27933;
  assign n27935 = ~n27214 & ~n27934;
  assign n27936 = ~controllable_hmaster3 & ~n27935;
  assign n27937 = ~n9517 & ~n27936;
  assign n27938 = i_hlock7 & ~n27937;
  assign n27939 = ~n10196 & ~n27261;
  assign n27940 = ~i_hbusreq8 & ~n27939;
  assign n27941 = ~n27241 & ~n27940;
  assign n27942 = ~controllable_hmaster3 & ~n27941;
  assign n27943 = ~n9517 & ~n27942;
  assign n27944 = ~i_hlock7 & ~n27943;
  assign n27945 = ~n27938 & ~n27944;
  assign n27946 = ~i_hbusreq7 & ~n27945;
  assign n27947 = ~n27213 & ~n27946;
  assign n27948 = ~n7924 & ~n27947;
  assign n27949 = ~n15491 & ~n27351;
  assign n27950 = ~i_hbusreq8 & ~n27949;
  assign n27951 = ~n27331 & ~n27950;
  assign n27952 = ~controllable_hmaster3 & ~n27951;
  assign n27953 = ~n27560 & ~n27952;
  assign n27954 = i_hlock7 & ~n27953;
  assign n27955 = ~n15491 & ~n27378;
  assign n27956 = ~i_hbusreq8 & ~n27955;
  assign n27957 = ~n27358 & ~n27956;
  assign n27958 = ~controllable_hmaster3 & ~n27957;
  assign n27959 = ~n27560 & ~n27958;
  assign n27960 = ~i_hlock7 & ~n27959;
  assign n27961 = ~n27954 & ~n27960;
  assign n27962 = ~i_hbusreq7 & ~n27961;
  assign n27963 = ~n27299 & ~n27962;
  assign n27964 = n7924 & ~n27963;
  assign n27965 = ~n27948 & ~n27964;
  assign n27966 = n8214 & ~n27965;
  assign n27967 = ~n27932 & ~n27966;
  assign n27968 = ~n8202 & ~n27967;
  assign n27969 = ~n9638 & ~n27226;
  assign n27970 = controllable_hmaster1 & ~n27969;
  assign n27971 = ~n9360 & ~n27970;
  assign n27972 = ~i_hbusreq6 & ~n27971;
  assign n27973 = ~n27215 & ~n27972;
  assign n27974 = ~controllable_hgrant6 & ~n27973;
  assign n27975 = ~n15520 & ~n27974;
  assign n27976 = controllable_hmaster0 & ~n27975;
  assign n27977 = ~n9439 & ~n27976;
  assign n27978 = ~i_hbusreq8 & ~n27977;
  assign n27979 = ~n27214 & ~n27978;
  assign n27980 = ~controllable_hmaster3 & ~n27979;
  assign n27981 = ~n9517 & ~n27980;
  assign n27982 = i_hlock7 & ~n27981;
  assign n27983 = ~n9638 & ~n27253;
  assign n27984 = controllable_hmaster1 & ~n27983;
  assign n27985 = ~n9360 & ~n27984;
  assign n27986 = ~i_hbusreq6 & ~n27985;
  assign n27987 = ~n27242 & ~n27986;
  assign n27988 = ~controllable_hgrant6 & ~n27987;
  assign n27989 = ~n15553 & ~n27988;
  assign n27990 = controllable_hmaster0 & ~n27989;
  assign n27991 = ~n9439 & ~n27990;
  assign n27992 = ~i_hbusreq8 & ~n27991;
  assign n27993 = ~n27241 & ~n27992;
  assign n27994 = ~controllable_hmaster3 & ~n27993;
  assign n27995 = ~n9517 & ~n27994;
  assign n27996 = ~i_hlock7 & ~n27995;
  assign n27997 = ~n27982 & ~n27996;
  assign n27998 = ~i_hbusreq7 & ~n27997;
  assign n27999 = ~n27213 & ~n27998;
  assign n28000 = ~n7924 & ~n27999;
  assign n28001 = ~n15538 & ~n27343;
  assign n28002 = controllable_hmaster1 & ~n28001;
  assign n28003 = ~n14605 & ~n28002;
  assign n28004 = ~i_hbusreq6 & ~n28003;
  assign n28005 = ~n27332 & ~n28004;
  assign n28006 = ~controllable_hgrant6 & ~n28005;
  assign n28007 = ~n15520 & ~n28006;
  assign n28008 = controllable_hmaster0 & ~n28007;
  assign n28009 = ~n14685 & ~n28008;
  assign n28010 = ~i_hbusreq8 & ~n28009;
  assign n28011 = ~n27331 & ~n28010;
  assign n28012 = ~controllable_hmaster3 & ~n28011;
  assign n28013 = ~n27560 & ~n28012;
  assign n28014 = i_hlock7 & ~n28013;
  assign n28015 = ~n15538 & ~n27370;
  assign n28016 = controllable_hmaster1 & ~n28015;
  assign n28017 = ~n14605 & ~n28016;
  assign n28018 = ~i_hbusreq6 & ~n28017;
  assign n28019 = ~n27359 & ~n28018;
  assign n28020 = ~controllable_hgrant6 & ~n28019;
  assign n28021 = ~n15553 & ~n28020;
  assign n28022 = controllable_hmaster0 & ~n28021;
  assign n28023 = ~n14685 & ~n28022;
  assign n28024 = ~i_hbusreq8 & ~n28023;
  assign n28025 = ~n27358 & ~n28024;
  assign n28026 = ~controllable_hmaster3 & ~n28025;
  assign n28027 = ~n27560 & ~n28026;
  assign n28028 = ~i_hlock7 & ~n28027;
  assign n28029 = ~n28014 & ~n28028;
  assign n28030 = ~i_hbusreq7 & ~n28029;
  assign n28031 = ~n27299 & ~n28030;
  assign n28032 = n7924 & ~n28031;
  assign n28033 = ~n28000 & ~n28032;
  assign n28034 = ~n8214 & ~n28033;
  assign n28035 = ~n10254 & ~n27234;
  assign n28036 = ~i_hbusreq8 & ~n28035;
  assign n28037 = ~n27214 & ~n28036;
  assign n28038 = ~controllable_hmaster3 & ~n28037;
  assign n28039 = ~n9517 & ~n28038;
  assign n28040 = i_hlock7 & ~n28039;
  assign n28041 = ~n10254 & ~n27261;
  assign n28042 = ~i_hbusreq8 & ~n28041;
  assign n28043 = ~n27241 & ~n28042;
  assign n28044 = ~controllable_hmaster3 & ~n28043;
  assign n28045 = ~n9517 & ~n28044;
  assign n28046 = ~i_hlock7 & ~n28045;
  assign n28047 = ~n28040 & ~n28046;
  assign n28048 = ~i_hbusreq7 & ~n28047;
  assign n28049 = ~n27213 & ~n28048;
  assign n28050 = ~n7924 & ~n28049;
  assign n28051 = ~n15616 & ~n27351;
  assign n28052 = ~i_hbusreq8 & ~n28051;
  assign n28053 = ~n27331 & ~n28052;
  assign n28054 = ~controllable_hmaster3 & ~n28053;
  assign n28055 = ~n27560 & ~n28054;
  assign n28056 = i_hlock7 & ~n28055;
  assign n28057 = ~n15616 & ~n27378;
  assign n28058 = ~i_hbusreq8 & ~n28057;
  assign n28059 = ~n27358 & ~n28058;
  assign n28060 = ~controllable_hmaster3 & ~n28059;
  assign n28061 = ~n27560 & ~n28060;
  assign n28062 = ~i_hlock7 & ~n28061;
  assign n28063 = ~n28056 & ~n28062;
  assign n28064 = ~i_hbusreq7 & ~n28063;
  assign n28065 = ~n27299 & ~n28064;
  assign n28066 = n7924 & ~n28065;
  assign n28067 = ~n28050 & ~n28066;
  assign n28068 = n8214 & ~n28067;
  assign n28069 = ~n28034 & ~n28068;
  assign n28070 = n8202 & ~n28069;
  assign n28071 = ~n27968 & ~n28070;
  assign n28072 = n7920 & ~n28071;
  assign n28073 = ~n10014 & ~n28072;
  assign n28074 = ~n7728 & ~n28073;
  assign n28075 = ~n27874 & ~n28074;
  assign n28076 = n7723 & ~n28075;
  assign n28077 = ~n7723 & ~n28073;
  assign n28078 = ~n28076 & ~n28077;
  assign n28079 = n7714 & ~n28078;
  assign n28080 = n7723 & ~n28073;
  assign n28081 = ~n8640 & ~n28072;
  assign n28082 = n7728 & ~n28081;
  assign n28083 = ~n27690 & ~n28082;
  assign n28084 = ~n7723 & ~n28083;
  assign n28085 = ~n28080 & ~n28084;
  assign n28086 = ~n7714 & ~n28085;
  assign n28087 = ~n28079 & ~n28086;
  assign n28088 = ~n7705 & ~n28087;
  assign n28089 = ~n10052 & ~n28088;
  assign n28090 = n7808 & ~n28089;
  assign n28091 = ~n9908 & ~n28090;
  assign n28092 = ~n8195 & ~n28091;
  assign n28093 = n7924 & ~n27686;
  assign n28094 = ~n8214 & ~n28093;
  assign n28095 = controllable_hmaster3 & ~n8987;
  assign n28096 = ~n26896 & ~n28095;
  assign n28097 = i_hbusreq7 & ~n28096;
  assign n28098 = controllable_hmaster2 & ~n15696;
  assign n28099 = ~n10751 & ~n28098;
  assign n28100 = controllable_hmaster1 & ~n28099;
  assign n28101 = ~controllable_hmaster1 & ~n10750;
  assign n28102 = ~n28100 & ~n28101;
  assign n28103 = ~i_hbusreq6 & ~n28102;
  assign n28104 = ~n26900 & ~n28103;
  assign n28105 = ~controllable_hgrant6 & ~n28104;
  assign n28106 = ~n15812 & ~n28105;
  assign n28107 = controllable_hmaster0 & ~n28106;
  assign n28108 = ~n10782 & ~n28107;
  assign n28109 = ~i_hbusreq8 & ~n28108;
  assign n28110 = ~n26899 & ~n28109;
  assign n28111 = ~controllable_hmaster3 & ~n28110;
  assign n28112 = ~n10759 & ~n28111;
  assign n28113 = ~i_hbusreq7 & ~n28112;
  assign n28114 = ~n28097 & ~n28113;
  assign n28115 = ~n7924 & ~n28114;
  assign n28116 = controllable_hmaster3 & ~n13200;
  assign n28117 = ~n26942 & ~n28116;
  assign n28118 = i_hbusreq7 & ~n28117;
  assign n28119 = ~i_hbusreq8 & ~n15806;
  assign n28120 = ~n13297 & ~n28119;
  assign n28121 = controllable_hmaster3 & ~n28120;
  assign n28122 = controllable_hmaster2 & ~n15770;
  assign n28123 = ~n15799 & ~n28122;
  assign n28124 = controllable_hmaster1 & ~n28123;
  assign n28125 = ~controllable_hmaster1 & ~n15798;
  assign n28126 = ~n28124 & ~n28125;
  assign n28127 = ~i_hbusreq6 & ~n28126;
  assign n28128 = ~n26977 & ~n28127;
  assign n28129 = ~controllable_hgrant6 & ~n28128;
  assign n28130 = ~n15812 & ~n28129;
  assign n28131 = controllable_hmaster0 & ~n28130;
  assign n28132 = ~n15852 & ~n28131;
  assign n28133 = ~i_hbusreq8 & ~n28132;
  assign n28134 = ~n26976 & ~n28133;
  assign n28135 = ~controllable_hmaster3 & ~n28134;
  assign n28136 = ~n28121 & ~n28135;
  assign n28137 = ~i_hbusreq7 & ~n28136;
  assign n28138 = ~n28118 & ~n28137;
  assign n28139 = n7924 & ~n28138;
  assign n28140 = ~n28115 & ~n28139;
  assign n28141 = n8214 & ~n28140;
  assign n28142 = ~n28094 & ~n28141;
  assign n28143 = n8202 & ~n28142;
  assign n28144 = ~n10721 & ~n28143;
  assign n28145 = n7920 & ~n28144;
  assign n28146 = ~n10671 & ~n28145;
  assign n28147 = n7728 & ~n28146;
  assign n28148 = ~n10812 & ~n27686;
  assign n28149 = ~n8214 & ~n28148;
  assign n28150 = n8214 & ~n27687;
  assign n28151 = ~n28149 & ~n28150;
  assign n28152 = n8202 & ~n28151;
  assign n28153 = ~n10811 & ~n28152;
  assign n28154 = n7920 & ~n28153;
  assign n28155 = ~n10797 & ~n28154;
  assign n28156 = ~n7728 & ~n28155;
  assign n28157 = ~n28147 & ~n28156;
  assign n28158 = ~n7723 & ~n28157;
  assign n28159 = ~n7723 & ~n28158;
  assign n28160 = ~n7714 & ~n28159;
  assign n28161 = ~n7714 & ~n28160;
  assign n28162 = n7705 & ~n28161;
  assign n28163 = ~n10829 & ~n26890;
  assign n28164 = ~controllable_hgrant6 & ~n28163;
  assign n28165 = ~n15890 & ~n28164;
  assign n28166 = controllable_hmaster0 & ~n28165;
  assign n28167 = ~n9099 & ~n28166;
  assign n28168 = ~controllable_hmaster3 & ~n28167;
  assign n28169 = ~n9093 & ~n28168;
  assign n28170 = i_hbusreq7 & ~n28169;
  assign n28171 = i_hbusreq8 & ~n28167;
  assign n28172 = i_hbusreq6 & ~n28163;
  assign n28173 = ~n10839 & ~n26903;
  assign n28174 = ~i_hbusreq6 & ~n28173;
  assign n28175 = ~n28172 & ~n28174;
  assign n28176 = ~controllable_hgrant6 & ~n28175;
  assign n28177 = ~n15902 & ~n28176;
  assign n28178 = controllable_hmaster0 & ~n28177;
  assign n28179 = ~n9127 & ~n28178;
  assign n28180 = ~i_hbusreq8 & ~n28179;
  assign n28181 = ~n28171 & ~n28180;
  assign n28182 = ~controllable_hmaster3 & ~n28181;
  assign n28183 = ~n9117 & ~n28182;
  assign n28184 = ~i_hbusreq7 & ~n28183;
  assign n28185 = ~n28170 & ~n28184;
  assign n28186 = ~n7924 & ~n28185;
  assign n28187 = ~n15892 & ~n26936;
  assign n28188 = ~controllable_hgrant6 & ~n28187;
  assign n28189 = ~n15890 & ~n28188;
  assign n28190 = controllable_hmaster0 & ~n28189;
  assign n28191 = ~n13682 & ~n28190;
  assign n28192 = ~controllable_hmaster3 & ~n28191;
  assign n28193 = ~n27088 & ~n28192;
  assign n28194 = i_hbusreq7 & ~n28193;
  assign n28195 = i_hbusreq8 & ~n28191;
  assign n28196 = i_hbusreq6 & ~n28187;
  assign n28197 = ~n15927 & ~n26980;
  assign n28198 = ~i_hbusreq6 & ~n28197;
  assign n28199 = ~n28196 & ~n28198;
  assign n28200 = ~controllable_hgrant6 & ~n28199;
  assign n28201 = ~n15902 & ~n28200;
  assign n28202 = controllable_hmaster0 & ~n28201;
  assign n28203 = ~n13728 & ~n28202;
  assign n28204 = ~i_hbusreq8 & ~n28203;
  assign n28205 = ~n28195 & ~n28204;
  assign n28206 = ~controllable_hmaster3 & ~n28205;
  assign n28207 = ~n27174 & ~n28206;
  assign n28208 = ~i_hbusreq7 & ~n28207;
  assign n28209 = ~n28194 & ~n28208;
  assign n28210 = n7924 & ~n28209;
  assign n28211 = ~n28186 & ~n28210;
  assign n28212 = ~n8214 & ~n28211;
  assign n28213 = ~n10855 & ~n26894;
  assign n28214 = ~controllable_hmaster3 & ~n28213;
  assign n28215 = ~n9093 & ~n28214;
  assign n28216 = i_hbusreq7 & ~n28215;
  assign n28217 = i_hbusreq8 & ~n28213;
  assign n28218 = ~n10875 & ~n28107;
  assign n28219 = ~i_hbusreq8 & ~n28218;
  assign n28220 = ~n28217 & ~n28219;
  assign n28221 = ~controllable_hmaster3 & ~n28220;
  assign n28222 = ~n10867 & ~n28221;
  assign n28223 = ~i_hbusreq7 & ~n28222;
  assign n28224 = ~n28216 & ~n28223;
  assign n28225 = ~n7924 & ~n28224;
  assign n28226 = ~n15970 & ~n26940;
  assign n28227 = ~controllable_hmaster3 & ~n28226;
  assign n28228 = ~n27088 & ~n28227;
  assign n28229 = i_hbusreq7 & ~n28228;
  assign n28230 = ~i_hbusreq8 & ~n15989;
  assign n28231 = ~n27111 & ~n28230;
  assign n28232 = controllable_hmaster3 & ~n28231;
  assign n28233 = i_hbusreq8 & ~n28226;
  assign n28234 = ~n16005 & ~n28131;
  assign n28235 = ~i_hbusreq8 & ~n28234;
  assign n28236 = ~n28233 & ~n28235;
  assign n28237 = ~controllable_hmaster3 & ~n28236;
  assign n28238 = ~n28232 & ~n28237;
  assign n28239 = ~i_hbusreq7 & ~n28238;
  assign n28240 = ~n28229 & ~n28239;
  assign n28241 = n7924 & ~n28240;
  assign n28242 = ~n28225 & ~n28241;
  assign n28243 = n8214 & ~n28242;
  assign n28244 = ~n28212 & ~n28243;
  assign n28245 = ~n8202 & ~n28244;
  assign n28246 = n8202 & ~n27687;
  assign n28247 = ~n28245 & ~n28246;
  assign n28248 = n7920 & ~n28247;
  assign n28249 = ~n10797 & ~n28248;
  assign n28250 = n7728 & ~n28249;
  assign n28251 = ~n10892 & ~n27228;
  assign n28252 = ~i_hbusreq6 & ~n28251;
  assign n28253 = ~n27215 & ~n28252;
  assign n28254 = ~controllable_hgrant6 & ~n28253;
  assign n28255 = ~n16031 & ~n28254;
  assign n28256 = controllable_hmaster0 & ~n28255;
  assign n28257 = ~n9439 & ~n28256;
  assign n28258 = ~i_hbusreq8 & ~n28257;
  assign n28259 = ~n27214 & ~n28258;
  assign n28260 = ~controllable_hmaster3 & ~n28259;
  assign n28261 = ~n9517 & ~n28260;
  assign n28262 = i_hlock7 & ~n28261;
  assign n28263 = ~n10892 & ~n27255;
  assign n28264 = ~i_hbusreq6 & ~n28263;
  assign n28265 = ~n27242 & ~n28264;
  assign n28266 = ~controllable_hgrant6 & ~n28265;
  assign n28267 = ~n16068 & ~n28266;
  assign n28268 = controllable_hmaster0 & ~n28267;
  assign n28269 = ~n9439 & ~n28268;
  assign n28270 = ~i_hbusreq8 & ~n28269;
  assign n28271 = ~n27241 & ~n28270;
  assign n28272 = ~controllable_hmaster3 & ~n28271;
  assign n28273 = ~n9517 & ~n28272;
  assign n28274 = ~i_hlock7 & ~n28273;
  assign n28275 = ~n28262 & ~n28274;
  assign n28276 = ~i_hbusreq7 & ~n28275;
  assign n28277 = ~n27213 & ~n28276;
  assign n28278 = ~n7924 & ~n28277;
  assign n28279 = ~n16055 & ~n27345;
  assign n28280 = ~i_hbusreq6 & ~n28279;
  assign n28281 = ~n27332 & ~n28280;
  assign n28282 = ~controllable_hgrant6 & ~n28281;
  assign n28283 = ~n16031 & ~n28282;
  assign n28284 = controllable_hmaster0 & ~n28283;
  assign n28285 = ~n14685 & ~n28284;
  assign n28286 = ~i_hbusreq8 & ~n28285;
  assign n28287 = ~n27331 & ~n28286;
  assign n28288 = ~controllable_hmaster3 & ~n28287;
  assign n28289 = ~n27560 & ~n28288;
  assign n28290 = i_hlock7 & ~n28289;
  assign n28291 = ~n16055 & ~n27372;
  assign n28292 = ~i_hbusreq6 & ~n28291;
  assign n28293 = ~n27359 & ~n28292;
  assign n28294 = ~controllable_hgrant6 & ~n28293;
  assign n28295 = ~n16068 & ~n28294;
  assign n28296 = controllable_hmaster0 & ~n28295;
  assign n28297 = ~n14685 & ~n28296;
  assign n28298 = ~i_hbusreq8 & ~n28297;
  assign n28299 = ~n27358 & ~n28298;
  assign n28300 = ~controllable_hmaster3 & ~n28299;
  assign n28301 = ~n27560 & ~n28300;
  assign n28302 = ~i_hlock7 & ~n28301;
  assign n28303 = ~n28290 & ~n28302;
  assign n28304 = ~i_hbusreq7 & ~n28303;
  assign n28305 = ~n27299 & ~n28304;
  assign n28306 = n7924 & ~n28305;
  assign n28307 = ~n28278 & ~n28306;
  assign n28308 = ~n8214 & ~n28307;
  assign n28309 = ~n28150 & ~n28308;
  assign n28310 = ~n8202 & ~n28309;
  assign n28311 = ~n28246 & ~n28310;
  assign n28312 = n7920 & ~n28311;
  assign n28313 = ~n10797 & ~n28312;
  assign n28314 = ~n7728 & ~n28313;
  assign n28315 = ~n28250 & ~n28314;
  assign n28316 = n7723 & ~n28315;
  assign n28317 = ~n7723 & ~n28313;
  assign n28318 = ~n28316 & ~n28317;
  assign n28319 = n7714 & ~n28318;
  assign n28320 = n7723 & ~n28313;
  assign n28321 = ~n8640 & ~n28312;
  assign n28322 = n7728 & ~n28321;
  assign n28323 = ~n27690 & ~n28322;
  assign n28324 = ~n7723 & ~n28323;
  assign n28325 = ~n28320 & ~n28324;
  assign n28326 = ~n7714 & ~n28325;
  assign n28327 = ~n28319 & ~n28326;
  assign n28328 = ~n7705 & ~n28327;
  assign n28329 = ~n28162 & ~n28328;
  assign n28330 = n7808 & ~n28329;
  assign n28331 = ~n10670 & ~n28330;
  assign n28332 = n8195 & ~n28331;
  assign n28333 = ~n28092 & ~n28332;
  assign n28334 = n8193 & ~n28333;
  assign n28335 = ~n27702 & ~n28334;
  assign n28336 = n8191 & ~n28335;
  assign n28337 = ~n11068 & ~n26838;
  assign n28338 = n7728 & ~n28337;
  assign n28339 = ~n11071 & ~n26879;
  assign n28340 = ~n7728 & ~n28339;
  assign n28341 = ~n28338 & ~n28340;
  assign n28342 = ~n7723 & ~n28341;
  assign n28343 = ~n7723 & ~n28342;
  assign n28344 = ~n7714 & ~n28343;
  assign n28345 = ~n7714 & ~n28344;
  assign n28346 = n7705 & ~n28345;
  assign n28347 = ~n11071 & ~n27189;
  assign n28348 = n7728 & ~n28347;
  assign n28349 = ~n11071 & ~n27582;
  assign n28350 = ~n7728 & ~n28349;
  assign n28351 = ~n28348 & ~n28350;
  assign n28352 = n7723 & ~n28351;
  assign n28353 = ~n7723 & ~n28349;
  assign n28354 = ~n28352 & ~n28353;
  assign n28355 = n7714 & ~n28354;
  assign n28356 = n7723 & ~n28349;
  assign n28357 = ~n11057 & ~n27582;
  assign n28358 = n7728 & ~n28357;
  assign n28359 = ~n11057 & ~n27688;
  assign n28360 = ~n7728 & ~n28359;
  assign n28361 = ~n28358 & ~n28360;
  assign n28362 = ~n7723 & ~n28361;
  assign n28363 = ~n28356 & ~n28362;
  assign n28364 = ~n7714 & ~n28363;
  assign n28365 = ~n28355 & ~n28364;
  assign n28366 = ~n7705 & ~n28365;
  assign n28367 = ~n28346 & ~n28366;
  assign n28368 = n7808 & ~n28367;
  assign n28369 = ~n11067 & ~n28368;
  assign n28370 = n8195 & ~n28369;
  assign n28371 = ~n8196 & ~n28370;
  assign n28372 = ~n8193 & ~n28371;
  assign n28373 = ~n11057 & ~n28072;
  assign n28374 = n7728 & ~n28373;
  assign n28375 = ~n28360 & ~n28374;
  assign n28376 = ~n7723 & ~n28375;
  assign n28377 = ~n28080 & ~n28376;
  assign n28378 = ~n7714 & ~n28377;
  assign n28379 = ~n28079 & ~n28378;
  assign n28380 = ~n7705 & ~n28379;
  assign n28381 = ~n10052 & ~n28380;
  assign n28382 = n7808 & ~n28381;
  assign n28383 = ~n11113 & ~n28382;
  assign n28384 = ~n8195 & ~n28383;
  assign n28385 = ~n11196 & ~n28145;
  assign n28386 = n7728 & ~n28385;
  assign n28387 = ~n11199 & ~n28154;
  assign n28388 = ~n7728 & ~n28387;
  assign n28389 = ~n28386 & ~n28388;
  assign n28390 = ~n7723 & ~n28389;
  assign n28391 = ~n7723 & ~n28390;
  assign n28392 = ~n7714 & ~n28391;
  assign n28393 = ~n7714 & ~n28392;
  assign n28394 = n7705 & ~n28393;
  assign n28395 = ~n11199 & ~n28248;
  assign n28396 = n7728 & ~n28395;
  assign n28397 = ~n11199 & ~n28312;
  assign n28398 = ~n7728 & ~n28397;
  assign n28399 = ~n28396 & ~n28398;
  assign n28400 = n7723 & ~n28399;
  assign n28401 = ~n7723 & ~n28397;
  assign n28402 = ~n28400 & ~n28401;
  assign n28403 = n7714 & ~n28402;
  assign n28404 = n7723 & ~n28397;
  assign n28405 = ~n11057 & ~n28312;
  assign n28406 = n7728 & ~n28405;
  assign n28407 = ~n28360 & ~n28406;
  assign n28408 = ~n7723 & ~n28407;
  assign n28409 = ~n28404 & ~n28408;
  assign n28410 = ~n7714 & ~n28409;
  assign n28411 = ~n28403 & ~n28410;
  assign n28412 = ~n7705 & ~n28411;
  assign n28413 = ~n28394 & ~n28412;
  assign n28414 = n7808 & ~n28413;
  assign n28415 = ~n11195 & ~n28414;
  assign n28416 = n8195 & ~n28415;
  assign n28417 = ~n28384 & ~n28416;
  assign n28418 = n8193 & ~n28417;
  assign n28419 = ~n28372 & ~n28418;
  assign n28420 = ~n8191 & ~n28419;
  assign n28421 = ~n28336 & ~n28420;
  assign n28422 = n8188 & ~n28421;
  assign n28423 = ~n11402 & ~n26838;
  assign n28424 = n7728 & ~n28423;
  assign n28425 = ~n11405 & ~n26879;
  assign n28426 = ~n7728 & ~n28425;
  assign n28427 = ~n28424 & ~n28426;
  assign n28428 = ~n7723 & ~n28427;
  assign n28429 = ~n7723 & ~n28428;
  assign n28430 = ~n7714 & ~n28429;
  assign n28431 = ~n7714 & ~n28430;
  assign n28432 = n7705 & ~n28431;
  assign n28433 = ~n11405 & ~n27189;
  assign n28434 = n7728 & ~n28433;
  assign n28435 = ~n11405 & ~n27582;
  assign n28436 = ~n7728 & ~n28435;
  assign n28437 = ~n28434 & ~n28436;
  assign n28438 = n7723 & ~n28437;
  assign n28439 = ~n7723 & ~n28435;
  assign n28440 = ~n28438 & ~n28439;
  assign n28441 = n7714 & ~n28440;
  assign n28442 = n7723 & ~n28435;
  assign n28443 = ~n11391 & ~n27582;
  assign n28444 = n7728 & ~n28443;
  assign n28445 = ~n11391 & ~n27688;
  assign n28446 = ~n7728 & ~n28445;
  assign n28447 = ~n28444 & ~n28446;
  assign n28448 = ~n7723 & ~n28447;
  assign n28449 = ~n28442 & ~n28448;
  assign n28450 = ~n7714 & ~n28449;
  assign n28451 = ~n28441 & ~n28450;
  assign n28452 = ~n7705 & ~n28451;
  assign n28453 = ~n28432 & ~n28452;
  assign n28454 = n7808 & ~n28453;
  assign n28455 = ~n11401 & ~n28454;
  assign n28456 = n8195 & ~n28455;
  assign n28457 = ~n8196 & ~n28456;
  assign n28458 = ~n8193 & ~n28457;
  assign n28459 = ~n11391 & ~n28072;
  assign n28460 = n7728 & ~n28459;
  assign n28461 = ~n28446 & ~n28460;
  assign n28462 = ~n7723 & ~n28461;
  assign n28463 = ~n28080 & ~n28462;
  assign n28464 = ~n7714 & ~n28463;
  assign n28465 = ~n28079 & ~n28464;
  assign n28466 = ~n7705 & ~n28465;
  assign n28467 = ~n10052 & ~n28466;
  assign n28468 = n7808 & ~n28467;
  assign n28469 = ~n11447 & ~n28468;
  assign n28470 = ~n8195 & ~n28469;
  assign n28471 = ~n11536 & ~n28145;
  assign n28472 = n7728 & ~n28471;
  assign n28473 = ~n11539 & ~n28154;
  assign n28474 = ~n7728 & ~n28473;
  assign n28475 = ~n28472 & ~n28474;
  assign n28476 = ~n7723 & ~n28475;
  assign n28477 = ~n7723 & ~n28476;
  assign n28478 = ~n7714 & ~n28477;
  assign n28479 = ~n7714 & ~n28478;
  assign n28480 = n7705 & ~n28479;
  assign n28481 = ~n11539 & ~n28248;
  assign n28482 = n7728 & ~n28481;
  assign n28483 = ~n11539 & ~n28312;
  assign n28484 = ~n7728 & ~n28483;
  assign n28485 = ~n28482 & ~n28484;
  assign n28486 = n7723 & ~n28485;
  assign n28487 = ~n7723 & ~n28483;
  assign n28488 = ~n28486 & ~n28487;
  assign n28489 = n7714 & ~n28488;
  assign n28490 = n7723 & ~n28483;
  assign n28491 = ~n11391 & ~n28312;
  assign n28492 = n7728 & ~n28491;
  assign n28493 = ~n28446 & ~n28492;
  assign n28494 = ~n7723 & ~n28493;
  assign n28495 = ~n28490 & ~n28494;
  assign n28496 = ~n7714 & ~n28495;
  assign n28497 = ~n28489 & ~n28496;
  assign n28498 = ~n7705 & ~n28497;
  assign n28499 = ~n28480 & ~n28498;
  assign n28500 = n7808 & ~n28499;
  assign n28501 = ~n11535 & ~n28500;
  assign n28502 = n8195 & ~n28501;
  assign n28503 = ~n28470 & ~n28502;
  assign n28504 = n8193 & ~n28503;
  assign n28505 = ~n28458 & ~n28504;
  assign n28506 = n8191 & ~n28505;
  assign n28507 = ~n11622 & ~n26838;
  assign n28508 = n7728 & ~n28507;
  assign n28509 = ~n11625 & ~n26879;
  assign n28510 = ~n7728 & ~n28509;
  assign n28511 = ~n28508 & ~n28510;
  assign n28512 = ~n7723 & ~n28511;
  assign n28513 = ~n7723 & ~n28512;
  assign n28514 = ~n7714 & ~n28513;
  assign n28515 = ~n7714 & ~n28514;
  assign n28516 = n7705 & ~n28515;
  assign n28517 = ~n11625 & ~n27189;
  assign n28518 = n7728 & ~n28517;
  assign n28519 = ~n11625 & ~n27582;
  assign n28520 = ~n7728 & ~n28519;
  assign n28521 = ~n28518 & ~n28520;
  assign n28522 = n7723 & ~n28521;
  assign n28523 = ~n7723 & ~n28519;
  assign n28524 = ~n28522 & ~n28523;
  assign n28525 = n7714 & ~n28524;
  assign n28526 = n7723 & ~n28519;
  assign n28527 = ~n11611 & ~n27582;
  assign n28528 = n7728 & ~n28527;
  assign n28529 = ~n11611 & ~n27688;
  assign n28530 = ~n7728 & ~n28529;
  assign n28531 = ~n28528 & ~n28530;
  assign n28532 = ~n7723 & ~n28531;
  assign n28533 = ~n28526 & ~n28532;
  assign n28534 = ~n7714 & ~n28533;
  assign n28535 = ~n28525 & ~n28534;
  assign n28536 = ~n7705 & ~n28535;
  assign n28537 = ~n28516 & ~n28536;
  assign n28538 = n7808 & ~n28537;
  assign n28539 = ~n11621 & ~n28538;
  assign n28540 = n8195 & ~n28539;
  assign n28541 = ~n8196 & ~n28540;
  assign n28542 = ~n8193 & ~n28541;
  assign n28543 = ~n11611 & ~n28072;
  assign n28544 = n7728 & ~n28543;
  assign n28545 = ~n28530 & ~n28544;
  assign n28546 = ~n7723 & ~n28545;
  assign n28547 = ~n28080 & ~n28546;
  assign n28548 = ~n7714 & ~n28547;
  assign n28549 = ~n28079 & ~n28548;
  assign n28550 = ~n7705 & ~n28549;
  assign n28551 = ~n10052 & ~n28550;
  assign n28552 = n7808 & ~n28551;
  assign n28553 = ~n11667 & ~n28552;
  assign n28554 = ~n8195 & ~n28553;
  assign n28555 = ~n11728 & ~n28145;
  assign n28556 = n7728 & ~n28555;
  assign n28557 = ~n11731 & ~n28154;
  assign n28558 = ~n7728 & ~n28557;
  assign n28559 = ~n28556 & ~n28558;
  assign n28560 = ~n7723 & ~n28559;
  assign n28561 = ~n7723 & ~n28560;
  assign n28562 = ~n7714 & ~n28561;
  assign n28563 = ~n7714 & ~n28562;
  assign n28564 = n7705 & ~n28563;
  assign n28565 = ~n11731 & ~n28248;
  assign n28566 = n7728 & ~n28565;
  assign n28567 = ~n11731 & ~n28312;
  assign n28568 = ~n7728 & ~n28567;
  assign n28569 = ~n28566 & ~n28568;
  assign n28570 = n7723 & ~n28569;
  assign n28571 = ~n7723 & ~n28567;
  assign n28572 = ~n28570 & ~n28571;
  assign n28573 = n7714 & ~n28572;
  assign n28574 = n7723 & ~n28567;
  assign n28575 = ~n11611 & ~n28312;
  assign n28576 = n7728 & ~n28575;
  assign n28577 = ~n28530 & ~n28576;
  assign n28578 = ~n7723 & ~n28577;
  assign n28579 = ~n28574 & ~n28578;
  assign n28580 = ~n7714 & ~n28579;
  assign n28581 = ~n28573 & ~n28580;
  assign n28582 = ~n7705 & ~n28581;
  assign n28583 = ~n28564 & ~n28582;
  assign n28584 = n7808 & ~n28583;
  assign n28585 = ~n11727 & ~n28584;
  assign n28586 = n8195 & ~n28585;
  assign n28587 = ~n28554 & ~n28586;
  assign n28588 = n8193 & ~n28587;
  assign n28589 = ~n28542 & ~n28588;
  assign n28590 = ~n8191 & ~n28589;
  assign n28591 = ~n28506 & ~n28590;
  assign n28592 = ~n8188 & ~n28591;
  assign n28593 = ~n28422 & ~n28592;
  assign n28594 = n8185 & ~n28593;
  assign n28595 = controllable_hgrant6 & ~n8227;
  assign n28596 = controllable_hgrant5 & ~n8223;
  assign n28597 = controllable_hgrant4 & ~n8223;
  assign n28598 = ~controllable_hgrant4 & ~n16134;
  assign n28599 = ~n28597 & ~n28598;
  assign n28600 = ~controllable_hgrant5 & ~n28599;
  assign n28601 = ~n28596 & ~n28600;
  assign n28602 = controllable_hmaster2 & ~n28601;
  assign n28603 = controllable_hmaster2 & ~n28602;
  assign n28604 = controllable_hmaster1 & ~n28603;
  assign n28605 = controllable_hmaster1 & ~n28604;
  assign n28606 = ~controllable_hgrant6 & ~n28605;
  assign n28607 = ~n28595 & ~n28606;
  assign n28608 = controllable_hmaster0 & ~n28607;
  assign n28609 = controllable_hmaster0 & ~n28608;
  assign n28610 = ~controllable_hmaster3 & ~n28609;
  assign n28611 = ~controllable_hmaster3 & ~n28610;
  assign n28612 = i_hlock7 & ~n28611;
  assign n28613 = controllable_hgrant6 & ~n8241;
  assign n28614 = controllable_hgrant5 & ~n8237;
  assign n28615 = controllable_hgrant4 & ~n8237;
  assign n28616 = ~controllable_hgrant4 & ~n16152;
  assign n28617 = ~n28615 & ~n28616;
  assign n28618 = ~controllable_hgrant5 & ~n28617;
  assign n28619 = ~n28614 & ~n28618;
  assign n28620 = controllable_hmaster2 & ~n28619;
  assign n28621 = controllable_hmaster2 & ~n28620;
  assign n28622 = controllable_hmaster1 & ~n28621;
  assign n28623 = controllable_hmaster1 & ~n28622;
  assign n28624 = ~controllable_hgrant6 & ~n28623;
  assign n28625 = ~n28613 & ~n28624;
  assign n28626 = controllable_hmaster0 & ~n28625;
  assign n28627 = controllable_hmaster0 & ~n28626;
  assign n28628 = ~controllable_hmaster3 & ~n28627;
  assign n28629 = ~controllable_hmaster3 & ~n28628;
  assign n28630 = ~i_hlock7 & ~n28629;
  assign n28631 = ~n28612 & ~n28630;
  assign n28632 = i_hbusreq7 & ~n28631;
  assign n28633 = i_hbusreq8 & ~n28609;
  assign n28634 = controllable_hgrant6 & ~n11785;
  assign n28635 = i_hbusreq6 & ~n28605;
  assign n28636 = controllable_hgrant5 & ~n8277;
  assign n28637 = i_hbusreq5 & ~n28599;
  assign n28638 = controllable_hgrant4 & ~n8275;
  assign n28639 = i_hbusreq4 & ~n16134;
  assign n28640 = i_hbusreq9 & ~n16134;
  assign n28641 = ~i_hbusreq9 & ~n16201;
  assign n28642 = ~n28640 & ~n28641;
  assign n28643 = ~i_hbusreq4 & ~n28642;
  assign n28644 = ~n28639 & ~n28643;
  assign n28645 = ~controllable_hgrant4 & ~n28644;
  assign n28646 = ~n28638 & ~n28645;
  assign n28647 = ~i_hbusreq5 & ~n28646;
  assign n28648 = ~n28637 & ~n28647;
  assign n28649 = ~controllable_hgrant5 & ~n28648;
  assign n28650 = ~n28636 & ~n28649;
  assign n28651 = controllable_hmaster2 & ~n28650;
  assign n28652 = controllable_hmaster2 & ~n28651;
  assign n28653 = controllable_hmaster1 & ~n28652;
  assign n28654 = controllable_hmaster1 & ~n28653;
  assign n28655 = ~i_hbusreq6 & ~n28654;
  assign n28656 = ~n28635 & ~n28655;
  assign n28657 = ~controllable_hgrant6 & ~n28656;
  assign n28658 = ~n28634 & ~n28657;
  assign n28659 = controllable_hmaster0 & ~n28658;
  assign n28660 = controllable_hmaster0 & ~n28659;
  assign n28661 = ~i_hbusreq8 & ~n28660;
  assign n28662 = ~n28633 & ~n28661;
  assign n28663 = ~controllable_hmaster3 & ~n28662;
  assign n28664 = ~controllable_hmaster3 & ~n28663;
  assign n28665 = i_hlock7 & ~n28664;
  assign n28666 = i_hbusreq8 & ~n28627;
  assign n28667 = controllable_hgrant6 & ~n11796;
  assign n28668 = i_hbusreq6 & ~n28623;
  assign n28669 = controllable_hgrant5 & ~n8309;
  assign n28670 = i_hbusreq5 & ~n28617;
  assign n28671 = controllable_hgrant4 & ~n8307;
  assign n28672 = i_hbusreq4 & ~n16152;
  assign n28673 = i_hbusreq9 & ~n16152;
  assign n28674 = ~i_hbusreq9 & ~n16226;
  assign n28675 = ~n28673 & ~n28674;
  assign n28676 = ~i_hbusreq4 & ~n28675;
  assign n28677 = ~n28672 & ~n28676;
  assign n28678 = ~controllable_hgrant4 & ~n28677;
  assign n28679 = ~n28671 & ~n28678;
  assign n28680 = ~i_hbusreq5 & ~n28679;
  assign n28681 = ~n28670 & ~n28680;
  assign n28682 = ~controllable_hgrant5 & ~n28681;
  assign n28683 = ~n28669 & ~n28682;
  assign n28684 = controllable_hmaster2 & ~n28683;
  assign n28685 = controllable_hmaster2 & ~n28684;
  assign n28686 = controllable_hmaster1 & ~n28685;
  assign n28687 = controllable_hmaster1 & ~n28686;
  assign n28688 = ~i_hbusreq6 & ~n28687;
  assign n28689 = ~n28668 & ~n28688;
  assign n28690 = ~controllable_hgrant6 & ~n28689;
  assign n28691 = ~n28667 & ~n28690;
  assign n28692 = controllable_hmaster0 & ~n28691;
  assign n28693 = controllable_hmaster0 & ~n28692;
  assign n28694 = ~i_hbusreq8 & ~n28693;
  assign n28695 = ~n28666 & ~n28694;
  assign n28696 = ~controllable_hmaster3 & ~n28695;
  assign n28697 = ~controllable_hmaster3 & ~n28696;
  assign n28698 = ~i_hlock7 & ~n28697;
  assign n28699 = ~n28665 & ~n28698;
  assign n28700 = ~i_hbusreq7 & ~n28699;
  assign n28701 = ~n28632 & ~n28700;
  assign n28702 = n7924 & ~n28701;
  assign n28703 = n7924 & ~n28702;
  assign n28704 = ~n8214 & ~n28703;
  assign n28705 = ~n8330 & ~n28704;
  assign n28706 = n8202 & ~n28705;
  assign n28707 = n8202 & ~n28706;
  assign n28708 = n7728 & ~n28707;
  assign n28709 = ~n7743 & ~n28610;
  assign n28710 = i_hlock7 & ~n28709;
  assign n28711 = ~n7743 & ~n28628;
  assign n28712 = ~i_hlock7 & ~n28711;
  assign n28713 = ~n28710 & ~n28712;
  assign n28714 = i_hbusreq7 & ~n28713;
  assign n28715 = ~n7779 & ~n28663;
  assign n28716 = i_hlock7 & ~n28715;
  assign n28717 = ~n7779 & ~n28696;
  assign n28718 = ~i_hlock7 & ~n28717;
  assign n28719 = ~n28716 & ~n28718;
  assign n28720 = ~i_hbusreq7 & ~n28719;
  assign n28721 = ~n28714 & ~n28720;
  assign n28722 = n7924 & ~n28721;
  assign n28723 = ~n8337 & ~n28722;
  assign n28724 = ~n8214 & ~n28723;
  assign n28725 = ~n8345 & ~n28724;
  assign n28726 = n8202 & ~n28725;
  assign n28727 = ~n8335 & ~n28726;
  assign n28728 = ~n7728 & ~n28727;
  assign n28729 = ~n28708 & ~n28728;
  assign n28730 = ~n7723 & ~n28729;
  assign n28731 = ~n7723 & ~n28730;
  assign n28732 = ~n7714 & ~n28731;
  assign n28733 = ~n7714 & ~n28732;
  assign n28734 = n7705 & ~n28733;
  assign n28735 = n7723 & ~n28727;
  assign n28736 = controllable_hgrant6 & ~n11843;
  assign n28737 = ~n8373 & ~n28602;
  assign n28738 = controllable_hmaster1 & ~n28737;
  assign n28739 = ~n8399 & ~n28738;
  assign n28740 = ~controllable_hgrant6 & ~n28739;
  assign n28741 = ~n28736 & ~n28740;
  assign n28742 = controllable_hmaster0 & ~n28741;
  assign n28743 = ~n8461 & ~n28742;
  assign n28744 = ~controllable_hmaster3 & ~n28743;
  assign n28745 = ~n8362 & ~n28744;
  assign n28746 = i_hlock7 & ~n28745;
  assign n28747 = controllable_hgrant6 & ~n11851;
  assign n28748 = ~n8373 & ~n28620;
  assign n28749 = controllable_hmaster1 & ~n28748;
  assign n28750 = ~n8399 & ~n28749;
  assign n28751 = ~controllable_hgrant6 & ~n28750;
  assign n28752 = ~n28747 & ~n28751;
  assign n28753 = controllable_hmaster0 & ~n28752;
  assign n28754 = ~n8461 & ~n28753;
  assign n28755 = ~controllable_hmaster3 & ~n28754;
  assign n28756 = ~n8362 & ~n28755;
  assign n28757 = ~i_hlock7 & ~n28756;
  assign n28758 = ~n28746 & ~n28757;
  assign n28759 = i_hbusreq7 & ~n28758;
  assign n28760 = i_hbusreq8 & ~n28743;
  assign n28761 = controllable_hgrant6 & ~n11865;
  assign n28762 = i_hbusreq6 & ~n28739;
  assign n28763 = ~n8514 & ~n28651;
  assign n28764 = controllable_hmaster1 & ~n28763;
  assign n28765 = ~n8552 & ~n28764;
  assign n28766 = ~i_hbusreq6 & ~n28765;
  assign n28767 = ~n28762 & ~n28766;
  assign n28768 = ~controllable_hgrant6 & ~n28767;
  assign n28769 = ~n28761 & ~n28768;
  assign n28770 = controllable_hmaster0 & ~n28769;
  assign n28771 = ~n8630 & ~n28770;
  assign n28772 = ~i_hbusreq8 & ~n28771;
  assign n28773 = ~n28760 & ~n28772;
  assign n28774 = ~controllable_hmaster3 & ~n28773;
  assign n28775 = ~n8492 & ~n28774;
  assign n28776 = i_hlock7 & ~n28775;
  assign n28777 = i_hbusreq8 & ~n28754;
  assign n28778 = controllable_hgrant6 & ~n11879;
  assign n28779 = i_hbusreq6 & ~n28750;
  assign n28780 = ~n8514 & ~n28684;
  assign n28781 = controllable_hmaster1 & ~n28780;
  assign n28782 = ~n8552 & ~n28781;
  assign n28783 = ~i_hbusreq6 & ~n28782;
  assign n28784 = ~n28779 & ~n28783;
  assign n28785 = ~controllable_hgrant6 & ~n28784;
  assign n28786 = ~n28778 & ~n28785;
  assign n28787 = controllable_hmaster0 & ~n28786;
  assign n28788 = ~n8630 & ~n28787;
  assign n28789 = ~i_hbusreq8 & ~n28788;
  assign n28790 = ~n28777 & ~n28789;
  assign n28791 = ~controllable_hmaster3 & ~n28790;
  assign n28792 = ~n8492 & ~n28791;
  assign n28793 = ~i_hlock7 & ~n28792;
  assign n28794 = ~n28776 & ~n28793;
  assign n28795 = ~i_hbusreq7 & ~n28794;
  assign n28796 = ~n28759 & ~n28795;
  assign n28797 = n7924 & ~n28796;
  assign n28798 = ~n8337 & ~n28797;
  assign n28799 = ~n7920 & ~n28798;
  assign n28800 = n7920 & ~n28727;
  assign n28801 = ~n28799 & ~n28800;
  assign n28802 = ~n7723 & ~n28801;
  assign n28803 = ~n28735 & ~n28802;
  assign n28804 = n7714 & ~n28803;
  assign n28805 = ~n7714 & ~n28798;
  assign n28806 = ~n28804 & ~n28805;
  assign n28807 = ~n7705 & ~n28806;
  assign n28808 = ~n28734 & ~n28807;
  assign n28809 = ~n7808 & ~n28808;
  assign n28810 = ~n7920 & ~n28707;
  assign n28811 = i_hlock9 & ~n16740;
  assign n28812 = ~i_hlock9 & ~n16759;
  assign n28813 = ~n28811 & ~n28812;
  assign n28814 = ~controllable_hgrant4 & ~n28813;
  assign n28815 = ~n12609 & ~n28814;
  assign n28816 = ~controllable_hgrant5 & ~n28815;
  assign n28817 = ~n12608 & ~n28816;
  assign n28818 = ~controllable_hmaster2 & ~n28817;
  assign n28819 = ~controllable_hmaster2 & ~n28818;
  assign n28820 = ~controllable_hmaster1 & ~n28819;
  assign n28821 = ~controllable_hmaster1 & ~n28820;
  assign n28822 = ~controllable_hgrant6 & ~n28821;
  assign n28823 = ~n12607 & ~n28822;
  assign n28824 = controllable_hmaster0 & ~n28823;
  assign n28825 = controllable_hmaster0 & ~n28824;
  assign n28826 = controllable_hmaster3 & ~n28825;
  assign n28827 = controllable_hmaster3 & ~n28826;
  assign n28828 = i_hbusreq7 & ~n28827;
  assign n28829 = i_hbusreq8 & ~n28825;
  assign n28830 = i_hbusreq6 & ~n28821;
  assign n28831 = i_hbusreq5 & ~n28815;
  assign n28832 = i_hbusreq4 & ~n28813;
  assign n28833 = i_hbusreq9 & ~n28813;
  assign n28834 = i_hlock9 & ~n16826;
  assign n28835 = ~i_hlock9 & ~n16863;
  assign n28836 = ~n28834 & ~n28835;
  assign n28837 = ~i_hbusreq9 & ~n28836;
  assign n28838 = ~n28833 & ~n28837;
  assign n28839 = ~i_hbusreq4 & ~n28838;
  assign n28840 = ~n28832 & ~n28839;
  assign n28841 = ~controllable_hgrant4 & ~n28840;
  assign n28842 = ~n12676 & ~n28841;
  assign n28843 = ~i_hbusreq5 & ~n28842;
  assign n28844 = ~n28831 & ~n28843;
  assign n28845 = ~controllable_hgrant5 & ~n28844;
  assign n28846 = ~n12674 & ~n28845;
  assign n28847 = ~controllable_hmaster2 & ~n28846;
  assign n28848 = ~controllable_hmaster2 & ~n28847;
  assign n28849 = ~controllable_hmaster1 & ~n28848;
  assign n28850 = ~controllable_hmaster1 & ~n28849;
  assign n28851 = ~i_hbusreq6 & ~n28850;
  assign n28852 = ~n28830 & ~n28851;
  assign n28853 = ~controllable_hgrant6 & ~n28852;
  assign n28854 = ~n12672 & ~n28853;
  assign n28855 = controllable_hmaster0 & ~n28854;
  assign n28856 = controllable_hmaster0 & ~n28855;
  assign n28857 = ~i_hbusreq8 & ~n28856;
  assign n28858 = ~n28829 & ~n28857;
  assign n28859 = controllable_hmaster3 & ~n28858;
  assign n28860 = controllable_hmaster3 & ~n28859;
  assign n28861 = ~i_hbusreq7 & ~n28860;
  assign n28862 = ~n28828 & ~n28861;
  assign n28863 = ~n8214 & ~n28862;
  assign n28864 = ~n16892 & ~n28863;
  assign n28865 = ~n8202 & ~n28864;
  assign n28866 = ~controllable_hgrant4 & ~n16359;
  assign n28867 = ~n13408 & ~n28866;
  assign n28868 = ~controllable_hgrant5 & ~n28867;
  assign n28869 = ~n13407 & ~n28868;
  assign n28870 = controllable_hmaster2 & ~n28869;
  assign n28871 = controllable_hmaster2 & ~n28870;
  assign n28872 = controllable_hmaster1 & ~n28871;
  assign n28873 = controllable_hmaster1 & ~n28872;
  assign n28874 = ~controllable_hgrant6 & ~n28873;
  assign n28875 = ~n16895 & ~n28874;
  assign n28876 = controllable_hmaster0 & ~n28875;
  assign n28877 = controllable_hmaster0 & ~n28876;
  assign n28878 = ~controllable_hmaster3 & ~n28877;
  assign n28879 = ~controllable_hmaster3 & ~n28878;
  assign n28880 = i_hlock7 & ~n28879;
  assign n28881 = ~controllable_hgrant4 & ~n16365;
  assign n28882 = ~n13429 & ~n28881;
  assign n28883 = ~controllable_hgrant5 & ~n28882;
  assign n28884 = ~n13428 & ~n28883;
  assign n28885 = controllable_hmaster2 & ~n28884;
  assign n28886 = controllable_hmaster2 & ~n28885;
  assign n28887 = controllable_hmaster1 & ~n28886;
  assign n28888 = controllable_hmaster1 & ~n28887;
  assign n28889 = ~controllable_hgrant6 & ~n28888;
  assign n28890 = ~n16907 & ~n28889;
  assign n28891 = controllable_hmaster0 & ~n28890;
  assign n28892 = controllable_hmaster0 & ~n28891;
  assign n28893 = ~controllable_hmaster3 & ~n28892;
  assign n28894 = ~controllable_hmaster3 & ~n28893;
  assign n28895 = ~i_hlock7 & ~n28894;
  assign n28896 = ~n28880 & ~n28895;
  assign n28897 = i_hbusreq7 & ~n28896;
  assign n28898 = i_hbusreq8 & ~n28877;
  assign n28899 = i_hbusreq6 & ~n28873;
  assign n28900 = i_hbusreq5 & ~n28867;
  assign n28901 = i_hbusreq4 & ~n16359;
  assign n28902 = i_hbusreq9 & ~n16359;
  assign n28903 = ~i_hbusreq9 & ~n16427;
  assign n28904 = ~n28902 & ~n28903;
  assign n28905 = ~i_hbusreq4 & ~n28904;
  assign n28906 = ~n28901 & ~n28905;
  assign n28907 = ~controllable_hgrant4 & ~n28906;
  assign n28908 = ~n13524 & ~n28907;
  assign n28909 = ~i_hbusreq5 & ~n28908;
  assign n28910 = ~n28900 & ~n28909;
  assign n28911 = ~controllable_hgrant5 & ~n28910;
  assign n28912 = ~n13522 & ~n28911;
  assign n28913 = controllable_hmaster2 & ~n28912;
  assign n28914 = controllable_hmaster2 & ~n28913;
  assign n28915 = controllable_hmaster1 & ~n28914;
  assign n28916 = controllable_hmaster1 & ~n28915;
  assign n28917 = ~i_hbusreq6 & ~n28916;
  assign n28918 = ~n28899 & ~n28917;
  assign n28919 = ~controllable_hgrant6 & ~n28918;
  assign n28920 = ~n16922 & ~n28919;
  assign n28921 = controllable_hmaster0 & ~n28920;
  assign n28922 = controllable_hmaster0 & ~n28921;
  assign n28923 = ~i_hbusreq8 & ~n28922;
  assign n28924 = ~n28898 & ~n28923;
  assign n28925 = ~controllable_hmaster3 & ~n28924;
  assign n28926 = ~controllable_hmaster3 & ~n28925;
  assign n28927 = i_hlock7 & ~n28926;
  assign n28928 = i_hbusreq8 & ~n28892;
  assign n28929 = i_hbusreq6 & ~n28888;
  assign n28930 = i_hbusreq5 & ~n28882;
  assign n28931 = i_hbusreq4 & ~n16365;
  assign n28932 = i_hbusreq9 & ~n16365;
  assign n28933 = ~i_hbusreq9 & ~n16439;
  assign n28934 = ~n28932 & ~n28933;
  assign n28935 = ~i_hbusreq4 & ~n28934;
  assign n28936 = ~n28931 & ~n28935;
  assign n28937 = ~controllable_hgrant4 & ~n28936;
  assign n28938 = ~n13577 & ~n28937;
  assign n28939 = ~i_hbusreq5 & ~n28938;
  assign n28940 = ~n28930 & ~n28939;
  assign n28941 = ~controllable_hgrant5 & ~n28940;
  assign n28942 = ~n13575 & ~n28941;
  assign n28943 = controllable_hmaster2 & ~n28942;
  assign n28944 = controllable_hmaster2 & ~n28943;
  assign n28945 = controllable_hmaster1 & ~n28944;
  assign n28946 = controllable_hmaster1 & ~n28945;
  assign n28947 = ~i_hbusreq6 & ~n28946;
  assign n28948 = ~n28929 & ~n28947;
  assign n28949 = ~controllable_hgrant6 & ~n28948;
  assign n28950 = ~n16940 & ~n28949;
  assign n28951 = controllable_hmaster0 & ~n28950;
  assign n28952 = controllable_hmaster0 & ~n28951;
  assign n28953 = ~i_hbusreq8 & ~n28952;
  assign n28954 = ~n28928 & ~n28953;
  assign n28955 = ~controllable_hmaster3 & ~n28954;
  assign n28956 = ~controllable_hmaster3 & ~n28955;
  assign n28957 = ~i_hlock7 & ~n28956;
  assign n28958 = ~n28927 & ~n28957;
  assign n28959 = ~i_hbusreq7 & ~n28958;
  assign n28960 = ~n28897 & ~n28959;
  assign n28961 = ~n7924 & ~n28960;
  assign n28962 = ~controllable_hgrant4 & ~n16481;
  assign n28963 = ~controllable_hgrant4 & ~n28962;
  assign n28964 = ~controllable_hgrant5 & ~n28963;
  assign n28965 = ~controllable_hgrant5 & ~n28964;
  assign n28966 = ~controllable_hgrant6 & ~n28965;
  assign n28967 = ~controllable_hgrant6 & ~n28966;
  assign n28968 = controllable_hmaster3 & ~n28967;
  assign n28969 = ~controllable_hgrant4 & ~n16515;
  assign n28970 = ~n13408 & ~n28969;
  assign n28971 = ~controllable_hgrant5 & ~n28970;
  assign n28972 = ~n13407 & ~n28971;
  assign n28973 = controllable_hmaster2 & ~n28972;
  assign n28974 = ~controllable_hmaster2 & ~n28965;
  assign n28975 = ~n28973 & ~n28974;
  assign n28976 = controllable_hmaster1 & ~n28975;
  assign n28977 = ~controllable_hmaster1 & ~n28965;
  assign n28978 = ~n28976 & ~n28977;
  assign n28979 = ~controllable_hgrant6 & ~n28978;
  assign n28980 = ~n16895 & ~n28979;
  assign n28981 = controllable_hmaster0 & ~n28980;
  assign n28982 = ~controllable_hmaster0 & ~n28967;
  assign n28983 = ~n28981 & ~n28982;
  assign n28984 = ~controllable_hmaster3 & ~n28983;
  assign n28985 = ~n28968 & ~n28984;
  assign n28986 = i_hlock7 & ~n28985;
  assign n28987 = ~controllable_hgrant4 & ~n16495;
  assign n28988 = ~controllable_hgrant4 & ~n28987;
  assign n28989 = ~controllable_hgrant5 & ~n28988;
  assign n28990 = ~controllable_hgrant5 & ~n28989;
  assign n28991 = ~controllable_hgrant6 & ~n28990;
  assign n28992 = ~controllable_hgrant6 & ~n28991;
  assign n28993 = controllable_hmaster3 & ~n28992;
  assign n28994 = ~controllable_hgrant4 & ~n16529;
  assign n28995 = ~n13429 & ~n28994;
  assign n28996 = ~controllable_hgrant5 & ~n28995;
  assign n28997 = ~n13428 & ~n28996;
  assign n28998 = controllable_hmaster2 & ~n28997;
  assign n28999 = ~controllable_hmaster2 & ~n28990;
  assign n29000 = ~n28998 & ~n28999;
  assign n29001 = controllable_hmaster1 & ~n29000;
  assign n29002 = ~controllable_hmaster1 & ~n28990;
  assign n29003 = ~n29001 & ~n29002;
  assign n29004 = ~controllable_hgrant6 & ~n29003;
  assign n29005 = ~n16907 & ~n29004;
  assign n29006 = controllable_hmaster0 & ~n29005;
  assign n29007 = ~controllable_hmaster0 & ~n28992;
  assign n29008 = ~n29006 & ~n29007;
  assign n29009 = ~controllable_hmaster3 & ~n29008;
  assign n29010 = ~n28993 & ~n29009;
  assign n29011 = ~i_hlock7 & ~n29010;
  assign n29012 = ~n28986 & ~n29011;
  assign n29013 = i_hbusreq7 & ~n29012;
  assign n29014 = i_hbusreq8 & ~n28967;
  assign n29015 = i_hbusreq6 & ~n28965;
  assign n29016 = i_hbusreq5 & ~n28963;
  assign n29017 = i_hbusreq4 & ~n16481;
  assign n29018 = i_hbusreq9 & ~n16481;
  assign n29019 = ~i_hbusreq9 & ~n16589;
  assign n29020 = ~n29018 & ~n29019;
  assign n29021 = ~i_hbusreq4 & ~n29020;
  assign n29022 = ~n29017 & ~n29021;
  assign n29023 = ~controllable_hgrant4 & ~n29022;
  assign n29024 = ~controllable_hgrant4 & ~n29023;
  assign n29025 = ~i_hbusreq5 & ~n29024;
  assign n29026 = ~n29016 & ~n29025;
  assign n29027 = ~controllable_hgrant5 & ~n29026;
  assign n29028 = ~controllable_hgrant5 & ~n29027;
  assign n29029 = ~i_hbusreq6 & ~n29028;
  assign n29030 = ~n29015 & ~n29029;
  assign n29031 = ~controllable_hgrant6 & ~n29030;
  assign n29032 = ~controllable_hgrant6 & ~n29031;
  assign n29033 = ~i_hbusreq8 & ~n29032;
  assign n29034 = ~n29014 & ~n29033;
  assign n29035 = controllable_hmaster3 & ~n29034;
  assign n29036 = i_hbusreq8 & ~n28983;
  assign n29037 = i_hbusreq6 & ~n28978;
  assign n29038 = i_hbusreq5 & ~n28970;
  assign n29039 = i_hbusreq4 & ~n16515;
  assign n29040 = i_hbusreq9 & ~n16515;
  assign n29041 = ~i_hbusreq9 & ~n16658;
  assign n29042 = ~n29040 & ~n29041;
  assign n29043 = ~i_hbusreq4 & ~n29042;
  assign n29044 = ~n29039 & ~n29043;
  assign n29045 = ~controllable_hgrant4 & ~n29044;
  assign n29046 = ~n13524 & ~n29045;
  assign n29047 = ~i_hbusreq5 & ~n29046;
  assign n29048 = ~n29038 & ~n29047;
  assign n29049 = ~controllable_hgrant5 & ~n29048;
  assign n29050 = ~n13522 & ~n29049;
  assign n29051 = controllable_hmaster2 & ~n29050;
  assign n29052 = ~controllable_hmaster2 & ~n29028;
  assign n29053 = ~n29051 & ~n29052;
  assign n29054 = controllable_hmaster1 & ~n29053;
  assign n29055 = ~controllable_hmaster1 & ~n29028;
  assign n29056 = ~n29054 & ~n29055;
  assign n29057 = ~i_hbusreq6 & ~n29056;
  assign n29058 = ~n29037 & ~n29057;
  assign n29059 = ~controllable_hgrant6 & ~n29058;
  assign n29060 = ~n16922 & ~n29059;
  assign n29061 = controllable_hmaster0 & ~n29060;
  assign n29062 = ~controllable_hmaster0 & ~n29032;
  assign n29063 = ~n29061 & ~n29062;
  assign n29064 = ~i_hbusreq8 & ~n29063;
  assign n29065 = ~n29036 & ~n29064;
  assign n29066 = ~controllable_hmaster3 & ~n29065;
  assign n29067 = ~n29035 & ~n29066;
  assign n29068 = i_hlock7 & ~n29067;
  assign n29069 = i_hbusreq8 & ~n28992;
  assign n29070 = i_hbusreq6 & ~n28990;
  assign n29071 = i_hbusreq5 & ~n28988;
  assign n29072 = i_hbusreq4 & ~n16495;
  assign n29073 = i_hbusreq9 & ~n16495;
  assign n29074 = ~i_hbusreq9 & ~n16603;
  assign n29075 = ~n29073 & ~n29074;
  assign n29076 = ~i_hbusreq4 & ~n29075;
  assign n29077 = ~n29072 & ~n29076;
  assign n29078 = ~controllable_hgrant4 & ~n29077;
  assign n29079 = ~controllable_hgrant4 & ~n29078;
  assign n29080 = ~i_hbusreq5 & ~n29079;
  assign n29081 = ~n29071 & ~n29080;
  assign n29082 = ~controllable_hgrant5 & ~n29081;
  assign n29083 = ~controllable_hgrant5 & ~n29082;
  assign n29084 = ~i_hbusreq6 & ~n29083;
  assign n29085 = ~n29070 & ~n29084;
  assign n29086 = ~controllable_hgrant6 & ~n29085;
  assign n29087 = ~controllable_hgrant6 & ~n29086;
  assign n29088 = ~i_hbusreq8 & ~n29087;
  assign n29089 = ~n29069 & ~n29088;
  assign n29090 = controllable_hmaster3 & ~n29089;
  assign n29091 = i_hbusreq8 & ~n29008;
  assign n29092 = i_hbusreq6 & ~n29003;
  assign n29093 = i_hbusreq5 & ~n28995;
  assign n29094 = i_hbusreq4 & ~n16529;
  assign n29095 = i_hbusreq9 & ~n16529;
  assign n29096 = ~i_hbusreq9 & ~n16680;
  assign n29097 = ~n29095 & ~n29096;
  assign n29098 = ~i_hbusreq4 & ~n29097;
  assign n29099 = ~n29094 & ~n29098;
  assign n29100 = ~controllable_hgrant4 & ~n29099;
  assign n29101 = ~n13577 & ~n29100;
  assign n29102 = ~i_hbusreq5 & ~n29101;
  assign n29103 = ~n29093 & ~n29102;
  assign n29104 = ~controllable_hgrant5 & ~n29103;
  assign n29105 = ~n13575 & ~n29104;
  assign n29106 = controllable_hmaster2 & ~n29105;
  assign n29107 = ~controllable_hmaster2 & ~n29083;
  assign n29108 = ~n29106 & ~n29107;
  assign n29109 = controllable_hmaster1 & ~n29108;
  assign n29110 = ~controllable_hmaster1 & ~n29083;
  assign n29111 = ~n29109 & ~n29110;
  assign n29112 = ~i_hbusreq6 & ~n29111;
  assign n29113 = ~n29092 & ~n29112;
  assign n29114 = ~controllable_hgrant6 & ~n29113;
  assign n29115 = ~n16940 & ~n29114;
  assign n29116 = controllable_hmaster0 & ~n29115;
  assign n29117 = ~controllable_hmaster0 & ~n29087;
  assign n29118 = ~n29116 & ~n29117;
  assign n29119 = ~i_hbusreq8 & ~n29118;
  assign n29120 = ~n29091 & ~n29119;
  assign n29121 = ~controllable_hmaster3 & ~n29120;
  assign n29122 = ~n29090 & ~n29121;
  assign n29123 = ~i_hlock7 & ~n29122;
  assign n29124 = ~n29068 & ~n29123;
  assign n29125 = ~i_hbusreq7 & ~n29124;
  assign n29126 = ~n29013 & ~n29125;
  assign n29127 = n7924 & ~n29126;
  assign n29128 = ~n28961 & ~n29127;
  assign n29129 = ~n8214 & ~n29128;
  assign n29130 = ~n16990 & ~n29129;
  assign n29131 = n8202 & ~n29130;
  assign n29132 = ~n28865 & ~n29131;
  assign n29133 = n7920 & ~n29132;
  assign n29134 = ~n28810 & ~n29133;
  assign n29135 = n7728 & ~n29134;
  assign n29136 = ~n7920 & ~n28727;
  assign n29137 = ~n7739 & ~n28818;
  assign n29138 = ~controllable_hmaster1 & ~n29137;
  assign n29139 = ~n7738 & ~n29138;
  assign n29140 = ~controllable_hgrant6 & ~n29139;
  assign n29141 = ~n12977 & ~n29140;
  assign n29142 = controllable_hmaster0 & ~n29141;
  assign n29143 = ~n8882 & ~n29142;
  assign n29144 = controllable_hmaster3 & ~n29143;
  assign n29145 = controllable_hmaster3 & ~n29144;
  assign n29146 = i_hbusreq7 & ~n29145;
  assign n29147 = i_hbusreq8 & ~n29143;
  assign n29148 = i_hbusreq6 & ~n29139;
  assign n29149 = ~n7771 & ~n28847;
  assign n29150 = ~controllable_hmaster1 & ~n29149;
  assign n29151 = ~n7770 & ~n29150;
  assign n29152 = ~i_hbusreq6 & ~n29151;
  assign n29153 = ~n29148 & ~n29152;
  assign n29154 = ~controllable_hgrant6 & ~n29153;
  assign n29155 = ~n12989 & ~n29154;
  assign n29156 = controllable_hmaster0 & ~n29155;
  assign n29157 = ~n8895 & ~n29156;
  assign n29158 = ~i_hbusreq8 & ~n29157;
  assign n29159 = ~n29147 & ~n29158;
  assign n29160 = controllable_hmaster3 & ~n29159;
  assign n29161 = controllable_hmaster3 & ~n29160;
  assign n29162 = ~i_hbusreq7 & ~n29161;
  assign n29163 = ~n29146 & ~n29162;
  assign n29164 = ~n8214 & ~n29163;
  assign n29165 = ~n17279 & ~n29164;
  assign n29166 = ~n8202 & ~n29165;
  assign n29167 = ~n24262 & ~n28878;
  assign n29168 = i_hlock7 & ~n29167;
  assign n29169 = ~n24262 & ~n28893;
  assign n29170 = ~i_hlock7 & ~n29169;
  assign n29171 = ~n29168 & ~n29170;
  assign n29172 = i_hbusreq7 & ~n29171;
  assign n29173 = i_hbusreq8 & ~n17022;
  assign n29174 = ~i_hbusreq8 & ~n17078;
  assign n29175 = ~n29173 & ~n29174;
  assign n29176 = controllable_hmaster3 & ~n29175;
  assign n29177 = ~n28925 & ~n29176;
  assign n29178 = i_hlock7 & ~n29177;
  assign n29179 = ~n28955 & ~n29176;
  assign n29180 = ~i_hlock7 & ~n29179;
  assign n29181 = ~n29178 & ~n29180;
  assign n29182 = ~i_hbusreq7 & ~n29181;
  assign n29183 = ~n29172 & ~n29182;
  assign n29184 = ~n7924 & ~n29183;
  assign n29185 = ~controllable_hgrant4 & ~n17099;
  assign n29186 = ~n7811 & ~n29185;
  assign n29187 = ~controllable_hgrant5 & ~n29186;
  assign n29188 = ~n7810 & ~n29187;
  assign n29189 = controllable_hmaster1 & ~n29188;
  assign n29190 = controllable_hmaster2 & ~n29188;
  assign n29191 = ~n28974 & ~n29190;
  assign n29192 = ~controllable_hmaster1 & ~n29191;
  assign n29193 = ~n29189 & ~n29192;
  assign n29194 = ~controllable_hgrant6 & ~n29193;
  assign n29195 = ~n7809 & ~n29194;
  assign n29196 = controllable_hmaster3 & ~n29195;
  assign n29197 = ~n28984 & ~n29196;
  assign n29198 = i_hlock7 & ~n29197;
  assign n29199 = ~controllable_hgrant4 & ~n17107;
  assign n29200 = ~n7811 & ~n29199;
  assign n29201 = ~controllable_hgrant5 & ~n29200;
  assign n29202 = ~n7810 & ~n29201;
  assign n29203 = controllable_hmaster1 & ~n29202;
  assign n29204 = controllable_hmaster2 & ~n29202;
  assign n29205 = ~n28999 & ~n29204;
  assign n29206 = ~controllable_hmaster1 & ~n29205;
  assign n29207 = ~n29203 & ~n29206;
  assign n29208 = ~controllable_hgrant6 & ~n29207;
  assign n29209 = ~n7809 & ~n29208;
  assign n29210 = controllable_hmaster3 & ~n29209;
  assign n29211 = ~n29009 & ~n29210;
  assign n29212 = ~i_hlock7 & ~n29211;
  assign n29213 = ~n29198 & ~n29212;
  assign n29214 = i_hbusreq7 & ~n29213;
  assign n29215 = i_hbusreq8 & ~n29195;
  assign n29216 = i_hbusreq6 & ~n29193;
  assign n29217 = i_hbusreq5 & ~n29186;
  assign n29218 = i_hbusreq4 & ~n17099;
  assign n29219 = i_hbusreq9 & ~n17099;
  assign n29220 = ~i_hbusreq9 & ~n17168;
  assign n29221 = ~n29219 & ~n29220;
  assign n29222 = ~i_hbusreq4 & ~n29221;
  assign n29223 = ~n29218 & ~n29222;
  assign n29224 = ~controllable_hgrant4 & ~n29223;
  assign n29225 = ~n7848 & ~n29224;
  assign n29226 = ~i_hbusreq5 & ~n29225;
  assign n29227 = ~n29217 & ~n29226;
  assign n29228 = ~controllable_hgrant5 & ~n29227;
  assign n29229 = ~n7846 & ~n29228;
  assign n29230 = controllable_hmaster1 & ~n29229;
  assign n29231 = controllable_hmaster2 & ~n29229;
  assign n29232 = ~n29052 & ~n29231;
  assign n29233 = ~controllable_hmaster1 & ~n29232;
  assign n29234 = ~n29230 & ~n29233;
  assign n29235 = ~i_hbusreq6 & ~n29234;
  assign n29236 = ~n29216 & ~n29235;
  assign n29237 = ~controllable_hgrant6 & ~n29236;
  assign n29238 = ~n7844 & ~n29237;
  assign n29239 = ~i_hbusreq8 & ~n29238;
  assign n29240 = ~n29215 & ~n29239;
  assign n29241 = controllable_hmaster3 & ~n29240;
  assign n29242 = ~n29066 & ~n29241;
  assign n29243 = i_hlock7 & ~n29242;
  assign n29244 = i_hbusreq8 & ~n29209;
  assign n29245 = i_hbusreq6 & ~n29207;
  assign n29246 = i_hbusreq5 & ~n29200;
  assign n29247 = i_hbusreq4 & ~n17107;
  assign n29248 = i_hbusreq9 & ~n17107;
  assign n29249 = ~i_hbusreq9 & ~n17182;
  assign n29250 = ~n29248 & ~n29249;
  assign n29251 = ~i_hbusreq4 & ~n29250;
  assign n29252 = ~n29247 & ~n29251;
  assign n29253 = ~controllable_hgrant4 & ~n29252;
  assign n29254 = ~n7848 & ~n29253;
  assign n29255 = ~i_hbusreq5 & ~n29254;
  assign n29256 = ~n29246 & ~n29255;
  assign n29257 = ~controllable_hgrant5 & ~n29256;
  assign n29258 = ~n7846 & ~n29257;
  assign n29259 = controllable_hmaster1 & ~n29258;
  assign n29260 = controllable_hmaster2 & ~n29258;
  assign n29261 = ~n29107 & ~n29260;
  assign n29262 = ~controllable_hmaster1 & ~n29261;
  assign n29263 = ~n29259 & ~n29262;
  assign n29264 = ~i_hbusreq6 & ~n29263;
  assign n29265 = ~n29245 & ~n29264;
  assign n29266 = ~controllable_hgrant6 & ~n29265;
  assign n29267 = ~n7844 & ~n29266;
  assign n29268 = ~i_hbusreq8 & ~n29267;
  assign n29269 = ~n29244 & ~n29268;
  assign n29270 = controllable_hmaster3 & ~n29269;
  assign n29271 = ~n29121 & ~n29270;
  assign n29272 = ~i_hlock7 & ~n29271;
  assign n29273 = ~n29243 & ~n29272;
  assign n29274 = ~i_hbusreq7 & ~n29273;
  assign n29275 = ~n29214 & ~n29274;
  assign n29276 = n7924 & ~n29275;
  assign n29277 = ~n29184 & ~n29276;
  assign n29278 = ~n8214 & ~n29277;
  assign n29279 = ~n17301 & ~n29278;
  assign n29280 = n8202 & ~n29279;
  assign n29281 = ~n29166 & ~n29280;
  assign n29282 = n7920 & ~n29281;
  assign n29283 = ~n29136 & ~n29282;
  assign n29284 = ~n7728 & ~n29283;
  assign n29285 = ~n29135 & ~n29284;
  assign n29286 = ~n7723 & ~n29285;
  assign n29287 = ~n7723 & ~n29286;
  assign n29288 = ~n7714 & ~n29287;
  assign n29289 = ~n7714 & ~n29288;
  assign n29290 = n7705 & ~n29289;
  assign n29291 = ~n8358 & ~n28818;
  assign n29292 = ~controllable_hmaster1 & ~n29291;
  assign n29293 = ~n8357 & ~n29292;
  assign n29294 = ~controllable_hgrant6 & ~n29293;
  assign n29295 = ~n13122 & ~n29294;
  assign n29296 = controllable_hmaster0 & ~n29295;
  assign n29297 = ~n8992 & ~n29296;
  assign n29298 = controllable_hmaster3 & ~n29297;
  assign n29299 = ~n26896 & ~n29298;
  assign n29300 = i_hbusreq7 & ~n29299;
  assign n29301 = i_hbusreq8 & ~n29297;
  assign n29302 = i_hbusreq6 & ~n29293;
  assign n29303 = ~n8484 & ~n28847;
  assign n29304 = ~controllable_hmaster1 & ~n29303;
  assign n29305 = ~n8483 & ~n29304;
  assign n29306 = ~i_hbusreq6 & ~n29305;
  assign n29307 = ~n29302 & ~n29306;
  assign n29308 = ~controllable_hgrant6 & ~n29307;
  assign n29309 = ~n13134 & ~n29308;
  assign n29310 = controllable_hmaster0 & ~n29309;
  assign n29311 = ~n9030 & ~n29310;
  assign n29312 = ~i_hbusreq8 & ~n29311;
  assign n29313 = ~n29301 & ~n29312;
  assign n29314 = controllable_hmaster3 & ~n29313;
  assign n29315 = ~n26913 & ~n29314;
  assign n29316 = ~i_hbusreq7 & ~n29315;
  assign n29317 = ~n29300 & ~n29316;
  assign n29318 = ~n7924 & ~n29317;
  assign n29319 = i_hlock9 & ~n17771;
  assign n29320 = ~i_hlock9 & ~n17789;
  assign n29321 = ~n29319 & ~n29320;
  assign n29322 = ~controllable_hgrant4 & ~n29321;
  assign n29323 = ~n12609 & ~n29322;
  assign n29324 = ~controllable_hgrant5 & ~n29323;
  assign n29325 = ~n12608 & ~n29324;
  assign n29326 = ~controllable_hmaster2 & ~n29325;
  assign n29327 = ~n13168 & ~n29326;
  assign n29328 = ~controllable_hmaster1 & ~n29327;
  assign n29329 = ~n13167 & ~n29328;
  assign n29330 = ~controllable_hgrant6 & ~n29329;
  assign n29331 = ~n13122 & ~n29330;
  assign n29332 = controllable_hmaster0 & ~n29331;
  assign n29333 = ~n13195 & ~n29332;
  assign n29334 = controllable_hmaster3 & ~n29333;
  assign n29335 = ~n26942 & ~n29334;
  assign n29336 = i_hbusreq7 & ~n29335;
  assign n29337 = i_hbusreq8 & ~n29333;
  assign n29338 = i_hbusreq6 & ~n29329;
  assign n29339 = i_hbusreq5 & ~n29323;
  assign n29340 = i_hbusreq4 & ~n29321;
  assign n29341 = i_hbusreq9 & ~n29321;
  assign n29342 = i_hlock9 & ~n17840;
  assign n29343 = ~i_hlock9 & ~n17876;
  assign n29344 = ~n29342 & ~n29343;
  assign n29345 = ~i_hbusreq9 & ~n29344;
  assign n29346 = ~n29341 & ~n29345;
  assign n29347 = ~i_hbusreq4 & ~n29346;
  assign n29348 = ~n29340 & ~n29347;
  assign n29349 = ~controllable_hgrant4 & ~n29348;
  assign n29350 = ~n12676 & ~n29349;
  assign n29351 = ~i_hbusreq5 & ~n29350;
  assign n29352 = ~n29339 & ~n29351;
  assign n29353 = ~controllable_hgrant5 & ~n29352;
  assign n29354 = ~n12674 & ~n29353;
  assign n29355 = ~controllable_hmaster2 & ~n29354;
  assign n29356 = ~n13480 & ~n29355;
  assign n29357 = ~controllable_hmaster1 & ~n29356;
  assign n29358 = ~n13479 & ~n29357;
  assign n29359 = ~i_hbusreq6 & ~n29358;
  assign n29360 = ~n29338 & ~n29359;
  assign n29361 = ~controllable_hgrant6 & ~n29360;
  assign n29362 = ~n13134 & ~n29361;
  assign n29363 = controllable_hmaster0 & ~n29362;
  assign n29364 = ~n13710 & ~n29363;
  assign n29365 = ~i_hbusreq8 & ~n29364;
  assign n29366 = ~n29337 & ~n29365;
  assign n29367 = controllable_hmaster3 & ~n29366;
  assign n29368 = ~n26990 & ~n29367;
  assign n29369 = ~i_hbusreq7 & ~n29368;
  assign n29370 = ~n29336 & ~n29369;
  assign n29371 = n7924 & ~n29370;
  assign n29372 = ~n29318 & ~n29371;
  assign n29373 = ~n8214 & ~n29372;
  assign n29374 = ~n9046 & ~n17710;
  assign n29375 = i_hlock8 & ~n29374;
  assign n29376 = ~n9046 & ~n17718;
  assign n29377 = ~i_hlock8 & ~n29376;
  assign n29378 = ~n29375 & ~n29377;
  assign n29379 = controllable_hmaster3 & ~n29378;
  assign n29380 = ~n26896 & ~n29379;
  assign n29381 = i_hbusreq7 & ~n29380;
  assign n29382 = i_hbusreq8 & ~n29378;
  assign n29383 = ~n9064 & ~n17734;
  assign n29384 = i_hlock8 & ~n29383;
  assign n29385 = ~n9064 & ~n17745;
  assign n29386 = ~i_hlock8 & ~n29385;
  assign n29387 = ~n29384 & ~n29386;
  assign n29388 = ~i_hbusreq8 & ~n29387;
  assign n29389 = ~n29382 & ~n29388;
  assign n29390 = controllable_hmaster3 & ~n29389;
  assign n29391 = ~n26913 & ~n29390;
  assign n29392 = ~i_hbusreq7 & ~n29391;
  assign n29393 = ~n29381 & ~n29392;
  assign n29394 = ~n7924 & ~n29393;
  assign n29395 = ~n17782 & ~n27003;
  assign n29396 = i_hlock8 & ~n29395;
  assign n29397 = ~n17800 & ~n27003;
  assign n29398 = ~i_hlock8 & ~n29397;
  assign n29399 = ~n29396 & ~n29398;
  assign n29400 = controllable_hmaster3 & ~n29399;
  assign n29401 = ~n26942 & ~n29400;
  assign n29402 = i_hbusreq7 & ~n29401;
  assign n29403 = i_hbusreq8 & ~n29399;
  assign n29404 = ~n17859 & ~n27013;
  assign n29405 = i_hlock8 & ~n29404;
  assign n29406 = ~n17895 & ~n27013;
  assign n29407 = ~i_hlock8 & ~n29406;
  assign n29408 = ~n29405 & ~n29407;
  assign n29409 = ~i_hbusreq8 & ~n29408;
  assign n29410 = ~n29403 & ~n29409;
  assign n29411 = controllable_hmaster3 & ~n29410;
  assign n29412 = ~n26990 & ~n29411;
  assign n29413 = ~i_hbusreq7 & ~n29412;
  assign n29414 = ~n29402 & ~n29413;
  assign n29415 = n7924 & ~n29414;
  assign n29416 = ~n29394 & ~n29415;
  assign n29417 = n8214 & ~n29416;
  assign n29418 = ~n29373 & ~n29417;
  assign n29419 = ~n8202 & ~n29418;
  assign n29420 = controllable_hmaster3 & ~n17345;
  assign n29421 = ~n17340 & ~n28870;
  assign n29422 = controllable_hmaster1 & ~n29421;
  assign n29423 = ~controllable_hmaster1 & ~n17339;
  assign n29424 = ~n29422 & ~n29423;
  assign n29425 = ~controllable_hgrant6 & ~n29424;
  assign n29426 = ~n13673 & ~n29425;
  assign n29427 = controllable_hmaster0 & ~n29426;
  assign n29428 = ~controllable_hmaster0 & ~n17350;
  assign n29429 = ~n29427 & ~n29428;
  assign n29430 = ~controllable_hmaster3 & ~n29429;
  assign n29431 = ~n29420 & ~n29430;
  assign n29432 = i_hlock7 & ~n29431;
  assign n29433 = ~n17340 & ~n28885;
  assign n29434 = controllable_hmaster1 & ~n29433;
  assign n29435 = ~n29423 & ~n29434;
  assign n29436 = ~controllable_hgrant6 & ~n29435;
  assign n29437 = ~n13687 & ~n29436;
  assign n29438 = controllable_hmaster0 & ~n29437;
  assign n29439 = ~n29428 & ~n29438;
  assign n29440 = ~controllable_hmaster3 & ~n29439;
  assign n29441 = ~n29420 & ~n29440;
  assign n29442 = ~i_hlock7 & ~n29441;
  assign n29443 = ~n29432 & ~n29442;
  assign n29444 = i_hbusreq7 & ~n29443;
  assign n29445 = i_hbusreq8 & ~n17345;
  assign n29446 = ~i_hbusreq8 & ~n17442;
  assign n29447 = ~n29445 & ~n29446;
  assign n29448 = controllable_hmaster3 & ~n29447;
  assign n29449 = i_hbusreq8 & ~n29429;
  assign n29450 = i_hbusreq6 & ~n29424;
  assign n29451 = ~n17435 & ~n28913;
  assign n29452 = controllable_hmaster1 & ~n29451;
  assign n29453 = ~controllable_hmaster1 & ~n17434;
  assign n29454 = ~n29452 & ~n29453;
  assign n29455 = ~i_hbusreq6 & ~n29454;
  assign n29456 = ~n29450 & ~n29455;
  assign n29457 = ~controllable_hgrant6 & ~n29456;
  assign n29458 = ~n13716 & ~n29457;
  assign n29459 = controllable_hmaster0 & ~n29458;
  assign n29460 = ~controllable_hmaster0 & ~n17453;
  assign n29461 = ~n29459 & ~n29460;
  assign n29462 = ~i_hbusreq8 & ~n29461;
  assign n29463 = ~n29449 & ~n29462;
  assign n29464 = ~controllable_hmaster3 & ~n29463;
  assign n29465 = ~n29448 & ~n29464;
  assign n29466 = i_hlock7 & ~n29465;
  assign n29467 = i_hbusreq8 & ~n29439;
  assign n29468 = i_hbusreq6 & ~n29435;
  assign n29469 = ~n17435 & ~n28943;
  assign n29470 = controllable_hmaster1 & ~n29469;
  assign n29471 = ~n29453 & ~n29470;
  assign n29472 = ~i_hbusreq6 & ~n29471;
  assign n29473 = ~n29468 & ~n29472;
  assign n29474 = ~controllable_hgrant6 & ~n29473;
  assign n29475 = ~n13736 & ~n29474;
  assign n29476 = controllable_hmaster0 & ~n29475;
  assign n29477 = ~n29460 & ~n29476;
  assign n29478 = ~i_hbusreq8 & ~n29477;
  assign n29479 = ~n29467 & ~n29478;
  assign n29480 = ~controllable_hmaster3 & ~n29479;
  assign n29481 = ~n29448 & ~n29480;
  assign n29482 = ~i_hlock7 & ~n29481;
  assign n29483 = ~n29466 & ~n29482;
  assign n29484 = ~i_hbusreq7 & ~n29483;
  assign n29485 = ~n29444 & ~n29484;
  assign n29486 = ~n7924 & ~n29485;
  assign n29487 = ~controllable_hgrant4 & ~n17474;
  assign n29488 = ~n13153 & ~n29487;
  assign n29489 = ~controllable_hgrant5 & ~n29488;
  assign n29490 = ~n13152 & ~n29489;
  assign n29491 = controllable_hmaster1 & ~n29490;
  assign n29492 = controllable_hmaster2 & ~n29490;
  assign n29493 = ~controllable_hgrant4 & ~n17514;
  assign n29494 = ~n13177 & ~n29493;
  assign n29495 = ~controllable_hgrant5 & ~n29494;
  assign n29496 = ~n13176 & ~n29495;
  assign n29497 = ~controllable_hmaster2 & ~n29496;
  assign n29498 = ~n29492 & ~n29497;
  assign n29499 = ~controllable_hmaster1 & ~n29498;
  assign n29500 = ~n29491 & ~n29499;
  assign n29501 = ~controllable_hgrant6 & ~n29500;
  assign n29502 = ~n13175 & ~n29501;
  assign n29503 = controllable_hmaster3 & ~n29502;
  assign n29504 = ~n28973 & ~n29497;
  assign n29505 = controllable_hmaster1 & ~n29504;
  assign n29506 = ~controllable_hmaster1 & ~n29496;
  assign n29507 = ~n29505 & ~n29506;
  assign n29508 = ~controllable_hgrant6 & ~n29507;
  assign n29509 = ~n13673 & ~n29508;
  assign n29510 = controllable_hmaster0 & ~n29509;
  assign n29511 = ~controllable_hgrant6 & ~n29496;
  assign n29512 = ~n13198 & ~n29511;
  assign n29513 = ~controllable_hmaster0 & ~n29512;
  assign n29514 = ~n29510 & ~n29513;
  assign n29515 = ~controllable_hmaster3 & ~n29514;
  assign n29516 = ~n29503 & ~n29515;
  assign n29517 = i_hlock7 & ~n29516;
  assign n29518 = ~controllable_hgrant4 & ~n17490;
  assign n29519 = ~n13153 & ~n29518;
  assign n29520 = ~controllable_hgrant5 & ~n29519;
  assign n29521 = ~n13152 & ~n29520;
  assign n29522 = controllable_hmaster1 & ~n29521;
  assign n29523 = controllable_hmaster2 & ~n29521;
  assign n29524 = ~controllable_hgrant4 & ~n17522;
  assign n29525 = ~n13177 & ~n29524;
  assign n29526 = ~controllable_hgrant5 & ~n29525;
  assign n29527 = ~n13176 & ~n29526;
  assign n29528 = ~controllable_hmaster2 & ~n29527;
  assign n29529 = ~n29523 & ~n29528;
  assign n29530 = ~controllable_hmaster1 & ~n29529;
  assign n29531 = ~n29522 & ~n29530;
  assign n29532 = ~controllable_hgrant6 & ~n29531;
  assign n29533 = ~n13175 & ~n29532;
  assign n29534 = controllable_hmaster3 & ~n29533;
  assign n29535 = ~n28998 & ~n29528;
  assign n29536 = controllable_hmaster1 & ~n29535;
  assign n29537 = ~controllable_hmaster1 & ~n29527;
  assign n29538 = ~n29536 & ~n29537;
  assign n29539 = ~controllable_hgrant6 & ~n29538;
  assign n29540 = ~n13687 & ~n29539;
  assign n29541 = controllable_hmaster0 & ~n29540;
  assign n29542 = ~controllable_hgrant6 & ~n29527;
  assign n29543 = ~n13198 & ~n29542;
  assign n29544 = ~controllable_hmaster0 & ~n29543;
  assign n29545 = ~n29541 & ~n29544;
  assign n29546 = ~controllable_hmaster3 & ~n29545;
  assign n29547 = ~n29534 & ~n29546;
  assign n29548 = ~i_hlock7 & ~n29547;
  assign n29549 = ~n29517 & ~n29548;
  assign n29550 = i_hbusreq7 & ~n29549;
  assign n29551 = i_hbusreq8 & ~n29502;
  assign n29552 = i_hbusreq6 & ~n29500;
  assign n29553 = i_hbusreq5 & ~n29488;
  assign n29554 = i_hbusreq4 & ~n17474;
  assign n29555 = i_hbusreq9 & ~n17474;
  assign n29556 = ~i_hbusreq9 & ~n17575;
  assign n29557 = ~n29555 & ~n29556;
  assign n29558 = ~i_hbusreq4 & ~n29557;
  assign n29559 = ~n29554 & ~n29558;
  assign n29560 = ~controllable_hgrant4 & ~n29559;
  assign n29561 = ~n13208 & ~n29560;
  assign n29562 = ~i_hbusreq5 & ~n29561;
  assign n29563 = ~n29553 & ~n29562;
  assign n29564 = ~controllable_hgrant5 & ~n29563;
  assign n29565 = ~n13206 & ~n29564;
  assign n29566 = controllable_hmaster1 & ~n29565;
  assign n29567 = controllable_hmaster2 & ~n29565;
  assign n29568 = i_hbusreq5 & ~n29494;
  assign n29569 = i_hbusreq4 & ~n17514;
  assign n29570 = i_hbusreq9 & ~n17514;
  assign n29571 = ~i_hbusreq9 & ~n17650;
  assign n29572 = ~n29570 & ~n29571;
  assign n29573 = ~i_hbusreq4 & ~n29572;
  assign n29574 = ~n29569 & ~n29573;
  assign n29575 = ~controllable_hgrant4 & ~n29574;
  assign n29576 = ~n13258 & ~n29575;
  assign n29577 = ~i_hbusreq5 & ~n29576;
  assign n29578 = ~n29568 & ~n29577;
  assign n29579 = ~controllable_hgrant5 & ~n29578;
  assign n29580 = ~n13256 & ~n29579;
  assign n29581 = ~controllable_hmaster2 & ~n29580;
  assign n29582 = ~n29567 & ~n29581;
  assign n29583 = ~controllable_hmaster1 & ~n29582;
  assign n29584 = ~n29566 & ~n29583;
  assign n29585 = ~i_hbusreq6 & ~n29584;
  assign n29586 = ~n29552 & ~n29585;
  assign n29587 = ~controllable_hgrant6 & ~n29586;
  assign n29588 = ~n13254 & ~n29587;
  assign n29589 = ~i_hbusreq8 & ~n29588;
  assign n29590 = ~n29551 & ~n29589;
  assign n29591 = controllable_hmaster3 & ~n29590;
  assign n29592 = i_hbusreq8 & ~n29514;
  assign n29593 = i_hbusreq6 & ~n29507;
  assign n29594 = ~n29051 & ~n29581;
  assign n29595 = controllable_hmaster1 & ~n29594;
  assign n29596 = ~controllable_hmaster1 & ~n29580;
  assign n29597 = ~n29595 & ~n29596;
  assign n29598 = ~i_hbusreq6 & ~n29597;
  assign n29599 = ~n29593 & ~n29598;
  assign n29600 = ~controllable_hgrant6 & ~n29599;
  assign n29601 = ~n13716 & ~n29600;
  assign n29602 = controllable_hmaster0 & ~n29601;
  assign n29603 = i_hbusreq6 & ~n29496;
  assign n29604 = ~i_hbusreq6 & ~n29580;
  assign n29605 = ~n29603 & ~n29604;
  assign n29606 = ~controllable_hgrant6 & ~n29605;
  assign n29607 = ~n13298 & ~n29606;
  assign n29608 = ~controllable_hmaster0 & ~n29607;
  assign n29609 = ~n29602 & ~n29608;
  assign n29610 = ~i_hbusreq8 & ~n29609;
  assign n29611 = ~n29592 & ~n29610;
  assign n29612 = ~controllable_hmaster3 & ~n29611;
  assign n29613 = ~n29591 & ~n29612;
  assign n29614 = i_hlock7 & ~n29613;
  assign n29615 = i_hbusreq8 & ~n29533;
  assign n29616 = i_hbusreq6 & ~n29531;
  assign n29617 = i_hbusreq5 & ~n29519;
  assign n29618 = i_hbusreq4 & ~n17490;
  assign n29619 = i_hbusreq9 & ~n17490;
  assign n29620 = ~i_hbusreq9 & ~n17597;
  assign n29621 = ~n29619 & ~n29620;
  assign n29622 = ~i_hbusreq4 & ~n29621;
  assign n29623 = ~n29618 & ~n29622;
  assign n29624 = ~controllable_hgrant4 & ~n29623;
  assign n29625 = ~n13208 & ~n29624;
  assign n29626 = ~i_hbusreq5 & ~n29625;
  assign n29627 = ~n29617 & ~n29626;
  assign n29628 = ~controllable_hgrant5 & ~n29627;
  assign n29629 = ~n13206 & ~n29628;
  assign n29630 = controllable_hmaster1 & ~n29629;
  assign n29631 = controllable_hmaster2 & ~n29629;
  assign n29632 = i_hbusreq5 & ~n29525;
  assign n29633 = i_hbusreq4 & ~n17522;
  assign n29634 = i_hbusreq9 & ~n17522;
  assign n29635 = ~i_hbusreq9 & ~n17664;
  assign n29636 = ~n29634 & ~n29635;
  assign n29637 = ~i_hbusreq4 & ~n29636;
  assign n29638 = ~n29633 & ~n29637;
  assign n29639 = ~controllable_hgrant4 & ~n29638;
  assign n29640 = ~n13258 & ~n29639;
  assign n29641 = ~i_hbusreq5 & ~n29640;
  assign n29642 = ~n29632 & ~n29641;
  assign n29643 = ~controllable_hgrant5 & ~n29642;
  assign n29644 = ~n13256 & ~n29643;
  assign n29645 = ~controllable_hmaster2 & ~n29644;
  assign n29646 = ~n29631 & ~n29645;
  assign n29647 = ~controllable_hmaster1 & ~n29646;
  assign n29648 = ~n29630 & ~n29647;
  assign n29649 = ~i_hbusreq6 & ~n29648;
  assign n29650 = ~n29616 & ~n29649;
  assign n29651 = ~controllable_hgrant6 & ~n29650;
  assign n29652 = ~n13254 & ~n29651;
  assign n29653 = ~i_hbusreq8 & ~n29652;
  assign n29654 = ~n29615 & ~n29653;
  assign n29655 = controllable_hmaster3 & ~n29654;
  assign n29656 = i_hbusreq8 & ~n29545;
  assign n29657 = i_hbusreq6 & ~n29538;
  assign n29658 = ~n29106 & ~n29645;
  assign n29659 = controllable_hmaster1 & ~n29658;
  assign n29660 = ~controllable_hmaster1 & ~n29644;
  assign n29661 = ~n29659 & ~n29660;
  assign n29662 = ~i_hbusreq6 & ~n29661;
  assign n29663 = ~n29657 & ~n29662;
  assign n29664 = ~controllable_hgrant6 & ~n29663;
  assign n29665 = ~n13736 & ~n29664;
  assign n29666 = controllable_hmaster0 & ~n29665;
  assign n29667 = i_hbusreq6 & ~n29527;
  assign n29668 = ~i_hbusreq6 & ~n29644;
  assign n29669 = ~n29667 & ~n29668;
  assign n29670 = ~controllable_hgrant6 & ~n29669;
  assign n29671 = ~n13298 & ~n29670;
  assign n29672 = ~controllable_hmaster0 & ~n29671;
  assign n29673 = ~n29666 & ~n29672;
  assign n29674 = ~i_hbusreq8 & ~n29673;
  assign n29675 = ~n29656 & ~n29674;
  assign n29676 = ~controllable_hmaster3 & ~n29675;
  assign n29677 = ~n29655 & ~n29676;
  assign n29678 = ~i_hlock7 & ~n29677;
  assign n29679 = ~n29614 & ~n29678;
  assign n29680 = ~i_hbusreq7 & ~n29679;
  assign n29681 = ~n29550 & ~n29680;
  assign n29682 = n7924 & ~n29681;
  assign n29683 = ~n29486 & ~n29682;
  assign n29684 = ~n8214 & ~n29683;
  assign n29685 = ~n18037 & ~n26894;
  assign n29686 = ~controllable_hmaster3 & ~n29685;
  assign n29687 = ~n9093 & ~n29686;
  assign n29688 = i_hbusreq7 & ~n29687;
  assign n29689 = i_hbusreq8 & ~n29685;
  assign n29690 = ~n18051 & ~n26909;
  assign n29691 = ~i_hbusreq8 & ~n29690;
  assign n29692 = ~n29689 & ~n29691;
  assign n29693 = ~controllable_hmaster3 & ~n29692;
  assign n29694 = ~n9117 & ~n29693;
  assign n29695 = ~i_hbusreq7 & ~n29694;
  assign n29696 = ~n29688 & ~n29695;
  assign n29697 = ~n7924 & ~n29696;
  assign n29698 = ~n18065 & ~n26940;
  assign n29699 = ~controllable_hmaster3 & ~n29698;
  assign n29700 = ~n27088 & ~n29699;
  assign n29701 = i_hbusreq7 & ~n29700;
  assign n29702 = i_hbusreq8 & ~n29698;
  assign n29703 = ~n18079 & ~n26986;
  assign n29704 = ~i_hbusreq8 & ~n29703;
  assign n29705 = ~n29702 & ~n29704;
  assign n29706 = ~controllable_hmaster3 & ~n29705;
  assign n29707 = ~n27174 & ~n29706;
  assign n29708 = ~i_hbusreq7 & ~n29707;
  assign n29709 = ~n29701 & ~n29708;
  assign n29710 = n7924 & ~n29709;
  assign n29711 = ~n29697 & ~n29710;
  assign n29712 = n8214 & ~n29711;
  assign n29713 = ~n29684 & ~n29712;
  assign n29714 = n8202 & ~n29713;
  assign n29715 = ~n29419 & ~n29714;
  assign n29716 = n7920 & ~n29715;
  assign n29717 = ~n29136 & ~n29716;
  assign n29718 = n7728 & ~n29717;
  assign n29719 = ~n19182 & ~n28818;
  assign n29720 = ~controllable_hmaster1 & ~n29719;
  assign n29721 = ~n19181 & ~n29720;
  assign n29722 = ~controllable_hgrant6 & ~n29721;
  assign n29723 = ~n13122 & ~n29722;
  assign n29724 = controllable_hmaster0 & ~n29723;
  assign n29725 = ~n20274 & ~n29724;
  assign n29726 = i_hlock8 & ~n29725;
  assign n29727 = ~n20283 & ~n29724;
  assign n29728 = ~i_hlock8 & ~n29727;
  assign n29729 = ~n29726 & ~n29728;
  assign n29730 = controllable_hmaster3 & ~n29729;
  assign n29731 = ~controllable_hgrant4 & ~n19188;
  assign n29732 = ~n13408 & ~n29731;
  assign n29733 = ~controllable_hgrant5 & ~n29732;
  assign n29734 = ~n13407 & ~n29733;
  assign n29735 = controllable_hmaster2 & ~n29734;
  assign n29736 = ~n19249 & ~n29735;
  assign n29737 = controllable_hmaster1 & ~n29736;
  assign n29738 = ~n19275 & ~n29737;
  assign n29739 = ~controllable_hgrant6 & ~n29738;
  assign n29740 = ~n13849 & ~n29739;
  assign n29741 = controllable_hmaster0 & ~n29740;
  assign n29742 = ~n19324 & ~n29741;
  assign n29743 = ~controllable_hmaster3 & ~n29742;
  assign n29744 = ~n29730 & ~n29743;
  assign n29745 = i_hlock7 & ~n29744;
  assign n29746 = ~controllable_hgrant4 & ~n19194;
  assign n29747 = ~n13429 & ~n29746;
  assign n29748 = ~controllable_hgrant5 & ~n29747;
  assign n29749 = ~n13428 & ~n29748;
  assign n29750 = controllable_hmaster2 & ~n29749;
  assign n29751 = ~n19249 & ~n29750;
  assign n29752 = controllable_hmaster1 & ~n29751;
  assign n29753 = ~n19275 & ~n29752;
  assign n29754 = ~controllable_hgrant6 & ~n29753;
  assign n29755 = ~n13951 & ~n29754;
  assign n29756 = controllable_hmaster0 & ~n29755;
  assign n29757 = ~n19324 & ~n29756;
  assign n29758 = ~controllable_hmaster3 & ~n29757;
  assign n29759 = ~n29730 & ~n29758;
  assign n29760 = ~i_hlock7 & ~n29759;
  assign n29761 = ~n29745 & ~n29760;
  assign n29762 = i_hbusreq7 & ~n29761;
  assign n29763 = i_hbusreq8 & ~n29729;
  assign n29764 = i_hbusreq6 & ~n29721;
  assign n29765 = ~n19367 & ~n28847;
  assign n29766 = ~controllable_hmaster1 & ~n29765;
  assign n29767 = ~n19366 & ~n29766;
  assign n29768 = ~i_hbusreq6 & ~n29767;
  assign n29769 = ~n29764 & ~n29768;
  assign n29770 = ~controllable_hgrant6 & ~n29769;
  assign n29771 = ~n13818 & ~n29770;
  assign n29772 = controllable_hmaster0 & ~n29771;
  assign n29773 = ~n20320 & ~n29772;
  assign n29774 = i_hlock8 & ~n29773;
  assign n29775 = ~n20332 & ~n29772;
  assign n29776 = ~i_hlock8 & ~n29775;
  assign n29777 = ~n29774 & ~n29776;
  assign n29778 = ~i_hbusreq8 & ~n29777;
  assign n29779 = ~n29763 & ~n29778;
  assign n29780 = controllable_hmaster3 & ~n29779;
  assign n29781 = i_hbusreq8 & ~n29742;
  assign n29782 = i_hbusreq6 & ~n29738;
  assign n29783 = i_hbusreq5 & ~n29732;
  assign n29784 = i_hbusreq4 & ~n19188;
  assign n29785 = i_hbusreq9 & ~n19188;
  assign n29786 = ~i_hbusreq9 & ~n19382;
  assign n29787 = ~n29785 & ~n29786;
  assign n29788 = ~i_hbusreq4 & ~n29787;
  assign n29789 = ~n29784 & ~n29788;
  assign n29790 = ~controllable_hgrant4 & ~n29789;
  assign n29791 = ~n14021 & ~n29790;
  assign n29792 = ~i_hbusreq5 & ~n29791;
  assign n29793 = ~n29783 & ~n29792;
  assign n29794 = ~controllable_hgrant5 & ~n29793;
  assign n29795 = ~n14020 & ~n29794;
  assign n29796 = controllable_hmaster2 & ~n29795;
  assign n29797 = ~n19497 & ~n29796;
  assign n29798 = controllable_hmaster1 & ~n29797;
  assign n29799 = ~n19550 & ~n29798;
  assign n29800 = ~i_hbusreq6 & ~n29799;
  assign n29801 = ~n29782 & ~n29800;
  assign n29802 = ~controllable_hgrant6 & ~n29801;
  assign n29803 = ~n14094 & ~n29802;
  assign n29804 = controllable_hmaster0 & ~n29803;
  assign n29805 = ~n19644 & ~n29804;
  assign n29806 = ~i_hbusreq8 & ~n29805;
  assign n29807 = ~n29781 & ~n29806;
  assign n29808 = ~controllable_hmaster3 & ~n29807;
  assign n29809 = ~n29780 & ~n29808;
  assign n29810 = i_hlock7 & ~n29809;
  assign n29811 = i_hbusreq8 & ~n29757;
  assign n29812 = i_hbusreq6 & ~n29753;
  assign n29813 = i_hbusreq5 & ~n29747;
  assign n29814 = i_hbusreq4 & ~n19194;
  assign n29815 = i_hbusreq9 & ~n19194;
  assign n29816 = ~i_hbusreq9 & ~n19394;
  assign n29817 = ~n29815 & ~n29816;
  assign n29818 = ~i_hbusreq4 & ~n29817;
  assign n29819 = ~n29814 & ~n29818;
  assign n29820 = ~controllable_hgrant4 & ~n29819;
  assign n29821 = ~n14056 & ~n29820;
  assign n29822 = ~i_hbusreq5 & ~n29821;
  assign n29823 = ~n29813 & ~n29822;
  assign n29824 = ~controllable_hgrant5 & ~n29823;
  assign n29825 = ~n14055 & ~n29824;
  assign n29826 = controllable_hmaster2 & ~n29825;
  assign n29827 = ~n19497 & ~n29826;
  assign n29828 = controllable_hmaster1 & ~n29827;
  assign n29829 = ~n19550 & ~n29828;
  assign n29830 = ~i_hbusreq6 & ~n29829;
  assign n29831 = ~n29812 & ~n29830;
  assign n29832 = ~controllable_hgrant6 & ~n29831;
  assign n29833 = ~n14298 & ~n29832;
  assign n29834 = controllable_hmaster0 & ~n29833;
  assign n29835 = ~n19644 & ~n29834;
  assign n29836 = ~i_hbusreq8 & ~n29835;
  assign n29837 = ~n29811 & ~n29836;
  assign n29838 = ~controllable_hmaster3 & ~n29837;
  assign n29839 = ~n29780 & ~n29838;
  assign n29840 = ~i_hlock7 & ~n29839;
  assign n29841 = ~n29810 & ~n29840;
  assign n29842 = ~i_hbusreq7 & ~n29841;
  assign n29843 = ~n29762 & ~n29842;
  assign n29844 = ~n7924 & ~n29843;
  assign n29845 = i_hlock9 & ~n19718;
  assign n29846 = ~i_hlock9 & ~n19736;
  assign n29847 = ~n29845 & ~n29846;
  assign n29848 = ~controllable_hgrant4 & ~n29847;
  assign n29849 = ~n12609 & ~n29848;
  assign n29850 = ~controllable_hgrant5 & ~n29849;
  assign n29851 = ~n12608 & ~n29850;
  assign n29852 = ~controllable_hmaster2 & ~n29851;
  assign n29853 = ~n19683 & ~n29852;
  assign n29854 = ~controllable_hmaster1 & ~n29853;
  assign n29855 = ~n19682 & ~n29854;
  assign n29856 = ~controllable_hgrant6 & ~n29855;
  assign n29857 = ~n13122 & ~n29856;
  assign n29858 = controllable_hmaster0 & ~n29857;
  assign n29859 = ~n20381 & ~n29858;
  assign n29860 = i_hlock8 & ~n29859;
  assign n29861 = ~n20390 & ~n29858;
  assign n29862 = ~i_hlock8 & ~n29861;
  assign n29863 = ~n29860 & ~n29862;
  assign n29864 = controllable_hmaster3 & ~n29863;
  assign n29865 = ~controllable_hgrant4 & ~n19689;
  assign n29866 = ~n13408 & ~n29865;
  assign n29867 = ~controllable_hgrant5 & ~n29866;
  assign n29868 = ~n13407 & ~n29867;
  assign n29869 = controllable_hmaster2 & ~n29868;
  assign n29870 = ~n19774 & ~n29869;
  assign n29871 = controllable_hmaster1 & ~n29870;
  assign n29872 = ~n19800 & ~n29871;
  assign n29873 = ~controllable_hgrant6 & ~n29872;
  assign n29874 = ~n13849 & ~n29873;
  assign n29875 = controllable_hmaster0 & ~n29874;
  assign n29876 = ~n19849 & ~n29875;
  assign n29877 = ~controllable_hmaster3 & ~n29876;
  assign n29878 = ~n29864 & ~n29877;
  assign n29879 = i_hlock7 & ~n29878;
  assign n29880 = ~controllable_hgrant4 & ~n19695;
  assign n29881 = ~n13429 & ~n29880;
  assign n29882 = ~controllable_hgrant5 & ~n29881;
  assign n29883 = ~n13428 & ~n29882;
  assign n29884 = controllable_hmaster2 & ~n29883;
  assign n29885 = ~n19774 & ~n29884;
  assign n29886 = controllable_hmaster1 & ~n29885;
  assign n29887 = ~n19800 & ~n29886;
  assign n29888 = ~controllable_hgrant6 & ~n29887;
  assign n29889 = ~n13951 & ~n29888;
  assign n29890 = controllable_hmaster0 & ~n29889;
  assign n29891 = ~n19849 & ~n29890;
  assign n29892 = ~controllable_hmaster3 & ~n29891;
  assign n29893 = ~n29864 & ~n29892;
  assign n29894 = ~i_hlock7 & ~n29893;
  assign n29895 = ~n29879 & ~n29894;
  assign n29896 = i_hbusreq7 & ~n29895;
  assign n29897 = i_hbusreq8 & ~n29863;
  assign n29898 = i_hbusreq6 & ~n29855;
  assign n29899 = i_hbusreq5 & ~n29849;
  assign n29900 = i_hbusreq4 & ~n29847;
  assign n29901 = i_hbusreq9 & ~n29847;
  assign n29902 = i_hlock9 & ~n19974;
  assign n29903 = ~i_hlock9 & ~n20010;
  assign n29904 = ~n29902 & ~n29903;
  assign n29905 = ~i_hbusreq9 & ~n29904;
  assign n29906 = ~n29901 & ~n29905;
  assign n29907 = ~i_hbusreq4 & ~n29906;
  assign n29908 = ~n29900 & ~n29907;
  assign n29909 = ~controllable_hgrant4 & ~n29908;
  assign n29910 = ~n12676 & ~n29909;
  assign n29911 = ~i_hbusreq5 & ~n29910;
  assign n29912 = ~n29899 & ~n29911;
  assign n29913 = ~controllable_hgrant5 & ~n29912;
  assign n29914 = ~n12674 & ~n29913;
  assign n29915 = ~controllable_hmaster2 & ~n29914;
  assign n29916 = ~n19895 & ~n29915;
  assign n29917 = ~controllable_hmaster1 & ~n29916;
  assign n29918 = ~n19894 & ~n29917;
  assign n29919 = ~i_hbusreq6 & ~n29918;
  assign n29920 = ~n29898 & ~n29919;
  assign n29921 = ~controllable_hgrant6 & ~n29920;
  assign n29922 = ~n13818 & ~n29921;
  assign n29923 = controllable_hmaster0 & ~n29922;
  assign n29924 = ~n20429 & ~n29923;
  assign n29925 = i_hlock8 & ~n29924;
  assign n29926 = ~n20441 & ~n29923;
  assign n29927 = ~i_hlock8 & ~n29926;
  assign n29928 = ~n29925 & ~n29927;
  assign n29929 = ~i_hbusreq8 & ~n29928;
  assign n29930 = ~n29897 & ~n29929;
  assign n29931 = controllable_hmaster3 & ~n29930;
  assign n29932 = i_hbusreq8 & ~n29876;
  assign n29933 = i_hbusreq6 & ~n29872;
  assign n29934 = i_hbusreq5 & ~n29866;
  assign n29935 = i_hbusreq4 & ~n19689;
  assign n29936 = i_hbusreq9 & ~n19689;
  assign n29937 = ~i_hbusreq9 & ~n19910;
  assign n29938 = ~n29936 & ~n29937;
  assign n29939 = ~i_hbusreq4 & ~n29938;
  assign n29940 = ~n29935 & ~n29939;
  assign n29941 = ~controllable_hgrant4 & ~n29940;
  assign n29942 = ~n14021 & ~n29941;
  assign n29943 = ~i_hbusreq5 & ~n29942;
  assign n29944 = ~n29934 & ~n29943;
  assign n29945 = ~controllable_hgrant5 & ~n29944;
  assign n29946 = ~n14020 & ~n29945;
  assign n29947 = controllable_hmaster2 & ~n29946;
  assign n29948 = ~n20090 & ~n29947;
  assign n29949 = controllable_hmaster1 & ~n29948;
  assign n29950 = ~n20143 & ~n29949;
  assign n29951 = ~i_hbusreq6 & ~n29950;
  assign n29952 = ~n29933 & ~n29951;
  assign n29953 = ~controllable_hgrant6 & ~n29952;
  assign n29954 = ~n14094 & ~n29953;
  assign n29955 = controllable_hmaster0 & ~n29954;
  assign n29956 = ~n20237 & ~n29955;
  assign n29957 = ~i_hbusreq8 & ~n29956;
  assign n29958 = ~n29932 & ~n29957;
  assign n29959 = ~controllable_hmaster3 & ~n29958;
  assign n29960 = ~n29931 & ~n29959;
  assign n29961 = i_hlock7 & ~n29960;
  assign n29962 = i_hbusreq8 & ~n29891;
  assign n29963 = i_hbusreq6 & ~n29887;
  assign n29964 = i_hbusreq5 & ~n29881;
  assign n29965 = i_hbusreq4 & ~n19695;
  assign n29966 = i_hbusreq9 & ~n19695;
  assign n29967 = ~i_hbusreq9 & ~n19922;
  assign n29968 = ~n29966 & ~n29967;
  assign n29969 = ~i_hbusreq4 & ~n29968;
  assign n29970 = ~n29965 & ~n29969;
  assign n29971 = ~controllable_hgrant4 & ~n29970;
  assign n29972 = ~n14056 & ~n29971;
  assign n29973 = ~i_hbusreq5 & ~n29972;
  assign n29974 = ~n29964 & ~n29973;
  assign n29975 = ~controllable_hgrant5 & ~n29974;
  assign n29976 = ~n14055 & ~n29975;
  assign n29977 = controllable_hmaster2 & ~n29976;
  assign n29978 = ~n20090 & ~n29977;
  assign n29979 = controllable_hmaster1 & ~n29978;
  assign n29980 = ~n20143 & ~n29979;
  assign n29981 = ~i_hbusreq6 & ~n29980;
  assign n29982 = ~n29963 & ~n29981;
  assign n29983 = ~controllable_hgrant6 & ~n29982;
  assign n29984 = ~n14298 & ~n29983;
  assign n29985 = controllable_hmaster0 & ~n29984;
  assign n29986 = ~n20237 & ~n29985;
  assign n29987 = ~i_hbusreq8 & ~n29986;
  assign n29988 = ~n29962 & ~n29987;
  assign n29989 = ~controllable_hmaster3 & ~n29988;
  assign n29990 = ~n29931 & ~n29989;
  assign n29991 = ~i_hlock7 & ~n29990;
  assign n29992 = ~n29961 & ~n29991;
  assign n29993 = ~i_hbusreq7 & ~n29992;
  assign n29994 = ~n29896 & ~n29993;
  assign n29995 = n7924 & ~n29994;
  assign n29996 = ~n29844 & ~n29995;
  assign n29997 = ~n8214 & ~n29996;
  assign n29998 = i_hlock9 & ~n19231;
  assign n29999 = ~i_hlock9 & ~n19254;
  assign n30000 = ~n29998 & ~n29999;
  assign n30001 = ~controllable_hgrant4 & ~n30000;
  assign n30002 = ~n12609 & ~n30001;
  assign n30003 = ~controllable_hgrant5 & ~n30002;
  assign n30004 = ~n12608 & ~n30003;
  assign n30005 = ~controllable_hmaster2 & ~n30004;
  assign n30006 = ~n19182 & ~n30005;
  assign n30007 = ~controllable_hmaster1 & ~n30006;
  assign n30008 = ~n19181 & ~n30007;
  assign n30009 = ~controllable_hgrant6 & ~n30008;
  assign n30010 = ~n13122 & ~n30009;
  assign n30011 = controllable_hmaster0 & ~n30010;
  assign n30012 = ~n19213 & ~n30011;
  assign n30013 = i_hlock8 & ~n30012;
  assign n30014 = ~n19221 & ~n30011;
  assign n30015 = ~i_hlock8 & ~n30014;
  assign n30016 = ~n30013 & ~n30015;
  assign n30017 = controllable_hmaster3 & ~n30016;
  assign n30018 = ~n29743 & ~n30017;
  assign n30019 = i_hlock7 & ~n30018;
  assign n30020 = ~n29758 & ~n30017;
  assign n30021 = ~i_hlock7 & ~n30020;
  assign n30022 = ~n30019 & ~n30021;
  assign n30023 = i_hbusreq7 & ~n30022;
  assign n30024 = i_hbusreq8 & ~n30016;
  assign n30025 = i_hbusreq6 & ~n30008;
  assign n30026 = i_hbusreq5 & ~n30002;
  assign n30027 = i_hbusreq4 & ~n30000;
  assign n30028 = i_hbusreq9 & ~n30000;
  assign n30029 = i_hlock9 & ~n19458;
  assign n30030 = ~i_hlock9 & ~n19508;
  assign n30031 = ~n30029 & ~n30030;
  assign n30032 = ~i_hbusreq9 & ~n30031;
  assign n30033 = ~n30028 & ~n30032;
  assign n30034 = ~i_hbusreq4 & ~n30033;
  assign n30035 = ~n30027 & ~n30034;
  assign n30036 = ~controllable_hgrant4 & ~n30035;
  assign n30037 = ~n14322 & ~n30036;
  assign n30038 = ~i_hbusreq5 & ~n30037;
  assign n30039 = ~n30026 & ~n30038;
  assign n30040 = ~controllable_hgrant5 & ~n30039;
  assign n30041 = ~n14321 & ~n30040;
  assign n30042 = ~controllable_hmaster2 & ~n30041;
  assign n30043 = ~n19367 & ~n30042;
  assign n30044 = ~controllable_hmaster1 & ~n30043;
  assign n30045 = ~n19366 & ~n30044;
  assign n30046 = ~i_hbusreq6 & ~n30045;
  assign n30047 = ~n30025 & ~n30046;
  assign n30048 = ~controllable_hgrant6 & ~n30047;
  assign n30049 = ~n14320 & ~n30048;
  assign n30050 = controllable_hmaster0 & ~n30049;
  assign n30051 = ~n19424 & ~n30050;
  assign n30052 = i_hlock8 & ~n30051;
  assign n30053 = ~n19435 & ~n30050;
  assign n30054 = ~i_hlock8 & ~n30053;
  assign n30055 = ~n30052 & ~n30054;
  assign n30056 = ~i_hbusreq8 & ~n30055;
  assign n30057 = ~n30024 & ~n30056;
  assign n30058 = controllable_hmaster3 & ~n30057;
  assign n30059 = ~n29808 & ~n30058;
  assign n30060 = i_hlock7 & ~n30059;
  assign n30061 = ~n29838 & ~n30058;
  assign n30062 = ~i_hlock7 & ~n30061;
  assign n30063 = ~n30060 & ~n30062;
  assign n30064 = ~i_hbusreq7 & ~n30063;
  assign n30065 = ~n30023 & ~n30064;
  assign n30066 = ~n7924 & ~n30065;
  assign n30067 = i_hlock9 & ~n19756;
  assign n30068 = ~i_hlock9 & ~n19779;
  assign n30069 = ~n30067 & ~n30068;
  assign n30070 = ~controllable_hgrant4 & ~n30069;
  assign n30071 = ~n12609 & ~n30070;
  assign n30072 = ~controllable_hgrant5 & ~n30071;
  assign n30073 = ~n12608 & ~n30072;
  assign n30074 = ~controllable_hmaster2 & ~n30073;
  assign n30075 = ~n19683 & ~n30074;
  assign n30076 = ~controllable_hmaster1 & ~n30075;
  assign n30077 = ~n19682 & ~n30076;
  assign n30078 = ~controllable_hgrant6 & ~n30077;
  assign n30079 = ~n13122 & ~n30078;
  assign n30080 = controllable_hmaster0 & ~n30079;
  assign n30081 = ~n19729 & ~n30080;
  assign n30082 = i_hlock8 & ~n30081;
  assign n30083 = ~n19747 & ~n30080;
  assign n30084 = ~i_hlock8 & ~n30083;
  assign n30085 = ~n30082 & ~n30084;
  assign n30086 = controllable_hmaster3 & ~n30085;
  assign n30087 = ~n29877 & ~n30086;
  assign n30088 = i_hlock7 & ~n30087;
  assign n30089 = ~n29892 & ~n30086;
  assign n30090 = ~i_hlock7 & ~n30089;
  assign n30091 = ~n30088 & ~n30090;
  assign n30092 = i_hbusreq7 & ~n30091;
  assign n30093 = i_hbusreq8 & ~n30085;
  assign n30094 = i_hbusreq6 & ~n30077;
  assign n30095 = i_hbusreq5 & ~n30071;
  assign n30096 = i_hbusreq4 & ~n30069;
  assign n30097 = i_hbusreq9 & ~n30069;
  assign n30098 = i_hlock9 & ~n20051;
  assign n30099 = ~i_hlock9 & ~n20101;
  assign n30100 = ~n30098 & ~n30099;
  assign n30101 = ~i_hbusreq9 & ~n30100;
  assign n30102 = ~n30097 & ~n30101;
  assign n30103 = ~i_hbusreq4 & ~n30102;
  assign n30104 = ~n30096 & ~n30103;
  assign n30105 = ~controllable_hgrant4 & ~n30104;
  assign n30106 = ~n14322 & ~n30105;
  assign n30107 = ~i_hbusreq5 & ~n30106;
  assign n30108 = ~n30095 & ~n30107;
  assign n30109 = ~controllable_hgrant5 & ~n30108;
  assign n30110 = ~n14321 & ~n30109;
  assign n30111 = ~controllable_hmaster2 & ~n30110;
  assign n30112 = ~n19895 & ~n30111;
  assign n30113 = ~controllable_hmaster1 & ~n30112;
  assign n30114 = ~n19894 & ~n30113;
  assign n30115 = ~i_hbusreq6 & ~n30114;
  assign n30116 = ~n30094 & ~n30115;
  assign n30117 = ~controllable_hgrant6 & ~n30116;
  assign n30118 = ~n14320 & ~n30117;
  assign n30119 = controllable_hmaster0 & ~n30118;
  assign n30120 = ~n19993 & ~n30119;
  assign n30121 = i_hlock8 & ~n30120;
  assign n30122 = ~n20029 & ~n30119;
  assign n30123 = ~i_hlock8 & ~n30122;
  assign n30124 = ~n30121 & ~n30123;
  assign n30125 = ~i_hbusreq8 & ~n30124;
  assign n30126 = ~n30093 & ~n30125;
  assign n30127 = controllable_hmaster3 & ~n30126;
  assign n30128 = ~n29959 & ~n30127;
  assign n30129 = i_hlock7 & ~n30128;
  assign n30130 = ~n29989 & ~n30127;
  assign n30131 = ~i_hlock7 & ~n30130;
  assign n30132 = ~n30129 & ~n30131;
  assign n30133 = ~i_hbusreq7 & ~n30132;
  assign n30134 = ~n30092 & ~n30133;
  assign n30135 = n7924 & ~n30134;
  assign n30136 = ~n30066 & ~n30135;
  assign n30137 = n8214 & ~n30136;
  assign n30138 = ~n29997 & ~n30137;
  assign n30139 = ~n8202 & ~n30138;
  assign n30140 = ~n17324 & ~n28818;
  assign n30141 = ~controllable_hmaster1 & ~n30140;
  assign n30142 = ~n17323 & ~n30141;
  assign n30143 = ~controllable_hgrant6 & ~n30142;
  assign n30144 = ~n13122 & ~n30143;
  assign n30145 = controllable_hmaster0 & ~n30144;
  assign n30146 = ~n18101 & ~n30145;
  assign n30147 = i_hlock8 & ~n30146;
  assign n30148 = ~n18109 & ~n30145;
  assign n30149 = ~i_hlock8 & ~n30148;
  assign n30150 = ~n30147 & ~n30149;
  assign n30151 = controllable_hmaster3 & ~n30150;
  assign n30152 = ~n18123 & ~n28870;
  assign n30153 = controllable_hmaster1 & ~n30152;
  assign n30154 = ~n18145 & ~n30153;
  assign n30155 = ~controllable_hgrant6 & ~n30154;
  assign n30156 = ~n13849 & ~n30155;
  assign n30157 = controllable_hmaster0 & ~n30156;
  assign n30158 = ~n18191 & ~n30157;
  assign n30159 = ~controllable_hmaster3 & ~n30158;
  assign n30160 = ~n30151 & ~n30159;
  assign n30161 = i_hlock7 & ~n30160;
  assign n30162 = ~n18123 & ~n28885;
  assign n30163 = controllable_hmaster1 & ~n30162;
  assign n30164 = ~n18145 & ~n30163;
  assign n30165 = ~controllable_hgrant6 & ~n30164;
  assign n30166 = ~n13951 & ~n30165;
  assign n30167 = controllable_hmaster0 & ~n30166;
  assign n30168 = ~n18191 & ~n30167;
  assign n30169 = ~controllable_hmaster3 & ~n30168;
  assign n30170 = ~n30151 & ~n30169;
  assign n30171 = ~i_hlock7 & ~n30170;
  assign n30172 = ~n30161 & ~n30171;
  assign n30173 = i_hbusreq7 & ~n30172;
  assign n30174 = i_hbusreq8 & ~n30150;
  assign n30175 = i_hbusreq6 & ~n30142;
  assign n30176 = i_hlock9 & ~n18268;
  assign n30177 = ~i_hlock9 & ~n18299;
  assign n30178 = ~n30176 & ~n30177;
  assign n30179 = ~i_hbusreq9 & ~n30178;
  assign n30180 = ~n28833 & ~n30179;
  assign n30181 = ~i_hbusreq4 & ~n30180;
  assign n30182 = ~n28832 & ~n30181;
  assign n30183 = ~controllable_hgrant4 & ~n30182;
  assign n30184 = ~n14322 & ~n30183;
  assign n30185 = ~i_hbusreq5 & ~n30184;
  assign n30186 = ~n28831 & ~n30185;
  assign n30187 = ~controllable_hgrant5 & ~n30186;
  assign n30188 = ~n14321 & ~n30187;
  assign n30189 = ~controllable_hmaster2 & ~n30188;
  assign n30190 = ~n18248 & ~n30189;
  assign n30191 = ~controllable_hmaster1 & ~n30190;
  assign n30192 = ~n18247 & ~n30191;
  assign n30193 = ~i_hbusreq6 & ~n30192;
  assign n30194 = ~n30175 & ~n30193;
  assign n30195 = ~controllable_hgrant6 & ~n30194;
  assign n30196 = ~n14320 & ~n30195;
  assign n30197 = controllable_hmaster0 & ~n30196;
  assign n30198 = ~n18287 & ~n30197;
  assign n30199 = i_hlock8 & ~n30198;
  assign n30200 = ~n18318 & ~n30197;
  assign n30201 = ~i_hlock8 & ~n30200;
  assign n30202 = ~n30199 & ~n30201;
  assign n30203 = ~i_hbusreq8 & ~n30202;
  assign n30204 = ~n30174 & ~n30203;
  assign n30205 = controllable_hmaster3 & ~n30204;
  assign n30206 = i_hbusreq8 & ~n30158;
  assign n30207 = i_hbusreq6 & ~n30154;
  assign n30208 = ~n18349 & ~n28913;
  assign n30209 = controllable_hmaster1 & ~n30208;
  assign n30210 = ~n18389 & ~n30209;
  assign n30211 = ~i_hbusreq6 & ~n30210;
  assign n30212 = ~n30207 & ~n30211;
  assign n30213 = ~controllable_hgrant6 & ~n30212;
  assign n30214 = ~n14756 & ~n30213;
  assign n30215 = controllable_hmaster0 & ~n30214;
  assign n30216 = ~n18503 & ~n30215;
  assign n30217 = ~i_hbusreq8 & ~n30216;
  assign n30218 = ~n30206 & ~n30217;
  assign n30219 = ~controllable_hmaster3 & ~n30218;
  assign n30220 = ~n30205 & ~n30219;
  assign n30221 = i_hlock7 & ~n30220;
  assign n30222 = i_hbusreq8 & ~n30168;
  assign n30223 = i_hbusreq6 & ~n30164;
  assign n30224 = ~n18349 & ~n28943;
  assign n30225 = controllable_hmaster1 & ~n30224;
  assign n30226 = ~n18389 & ~n30225;
  assign n30227 = ~i_hbusreq6 & ~n30226;
  assign n30228 = ~n30223 & ~n30227;
  assign n30229 = ~controllable_hgrant6 & ~n30228;
  assign n30230 = ~n14772 & ~n30229;
  assign n30231 = controllable_hmaster0 & ~n30230;
  assign n30232 = ~n18503 & ~n30231;
  assign n30233 = ~i_hbusreq8 & ~n30232;
  assign n30234 = ~n30222 & ~n30233;
  assign n30235 = ~controllable_hmaster3 & ~n30234;
  assign n30236 = ~n30205 & ~n30235;
  assign n30237 = ~i_hlock7 & ~n30236;
  assign n30238 = ~n30221 & ~n30237;
  assign n30239 = ~i_hbusreq7 & ~n30238;
  assign n30240 = ~n30173 & ~n30239;
  assign n30241 = ~n7924 & ~n30240;
  assign n30242 = ~i_hlock9 & ~n18560;
  assign n30243 = ~n18535 & ~n30242;
  assign n30244 = ~controllable_hgrant4 & ~n30243;
  assign n30245 = ~n12609 & ~n30244;
  assign n30246 = ~controllable_hgrant5 & ~n30245;
  assign n30247 = ~n12608 & ~n30246;
  assign n30248 = ~controllable_hmaster2 & ~n30247;
  assign n30249 = ~n29492 & ~n30248;
  assign n30250 = ~controllable_hmaster1 & ~n30249;
  assign n30251 = ~n29491 & ~n30250;
  assign n30252 = ~controllable_hgrant6 & ~n30251;
  assign n30253 = ~n13122 & ~n30252;
  assign n30254 = controllable_hmaster0 & ~n30253;
  assign n30255 = ~controllable_hgrant4 & ~n18534;
  assign n30256 = ~n13408 & ~n30255;
  assign n30257 = ~controllable_hgrant5 & ~n30256;
  assign n30258 = ~n13407 & ~n30257;
  assign n30259 = ~controllable_hmaster2 & ~n30258;
  assign n30260 = ~n29492 & ~n30259;
  assign n30261 = ~controllable_hmaster1 & ~n30260;
  assign n30262 = ~n29491 & ~n30261;
  assign n30263 = ~controllable_hgrant6 & ~n30262;
  assign n30264 = ~n13406 & ~n30263;
  assign n30265 = ~controllable_hmaster0 & ~n30264;
  assign n30266 = ~n30254 & ~n30265;
  assign n30267 = i_hlock8 & ~n30266;
  assign n30268 = ~controllable_hgrant4 & ~n18560;
  assign n30269 = ~n13429 & ~n30268;
  assign n30270 = ~controllable_hgrant5 & ~n30269;
  assign n30271 = ~n13428 & ~n30270;
  assign n30272 = ~controllable_hmaster2 & ~n30271;
  assign n30273 = ~n29492 & ~n30272;
  assign n30274 = ~controllable_hmaster1 & ~n30273;
  assign n30275 = ~n29491 & ~n30274;
  assign n30276 = ~controllable_hgrant6 & ~n30275;
  assign n30277 = ~n13427 & ~n30276;
  assign n30278 = ~controllable_hmaster0 & ~n30277;
  assign n30279 = ~n30254 & ~n30278;
  assign n30280 = ~i_hlock8 & ~n30279;
  assign n30281 = ~n30267 & ~n30280;
  assign n30282 = controllable_hmaster3 & ~n30281;
  assign n30283 = ~controllable_hgrant4 & ~n18589;
  assign n30284 = ~n13851 & ~n30283;
  assign n30285 = ~controllable_hgrant5 & ~n30284;
  assign n30286 = ~n13850 & ~n30285;
  assign n30287 = ~controllable_hmaster2 & ~n30286;
  assign n30288 = ~n28973 & ~n30287;
  assign n30289 = controllable_hmaster1 & ~n30288;
  assign n30290 = i_hlock5 & ~n30256;
  assign n30291 = ~i_hlock5 & ~n30269;
  assign n30292 = ~n30290 & ~n30291;
  assign n30293 = ~controllable_hgrant5 & ~n30292;
  assign n30294 = ~n13865 & ~n30293;
  assign n30295 = controllable_hmaster2 & ~n30294;
  assign n30296 = ~controllable_hgrant4 & ~n18617;
  assign n30297 = ~n13873 & ~n30296;
  assign n30298 = ~controllable_hgrant5 & ~n30297;
  assign n30299 = ~n13872 & ~n30298;
  assign n30300 = ~controllable_hmaster2 & ~n30299;
  assign n30301 = ~n30295 & ~n30300;
  assign n30302 = ~controllable_hmaster1 & ~n30301;
  assign n30303 = ~n30289 & ~n30302;
  assign n30304 = ~controllable_hgrant6 & ~n30303;
  assign n30305 = ~n13849 & ~n30304;
  assign n30306 = controllable_hmaster0 & ~n30305;
  assign n30307 = controllable_hmaster2 & ~n30258;
  assign n30308 = ~controllable_hgrant4 & ~n18643;
  assign n30309 = ~n13896 & ~n30308;
  assign n30310 = ~controllable_hgrant5 & ~n30309;
  assign n30311 = ~n13895 & ~n30310;
  assign n30312 = ~controllable_hmaster2 & ~n30311;
  assign n30313 = ~n30307 & ~n30312;
  assign n30314 = controllable_hmaster1 & ~n30313;
  assign n30315 = i_hlock4 & ~n18534;
  assign n30316 = ~i_hlock4 & ~n18560;
  assign n30317 = ~n30315 & ~n30316;
  assign n30318 = ~controllable_hgrant4 & ~n30317;
  assign n30319 = ~n13912 & ~n30318;
  assign n30320 = ~controllable_hgrant5 & ~n30319;
  assign n30321 = ~n13911 & ~n30320;
  assign n30322 = controllable_hmaster2 & ~n30321;
  assign n30323 = ~controllable_hgrant4 & ~n18671;
  assign n30324 = ~n13922 & ~n30323;
  assign n30325 = ~controllable_hgrant5 & ~n30324;
  assign n30326 = ~n13921 & ~n30325;
  assign n30327 = ~controllable_hmaster2 & ~n30326;
  assign n30328 = ~n30322 & ~n30327;
  assign n30329 = ~controllable_hmaster1 & ~n30328;
  assign n30330 = ~n30314 & ~n30329;
  assign n30331 = i_hlock6 & ~n30330;
  assign n30332 = controllable_hmaster2 & ~n30271;
  assign n30333 = ~n30312 & ~n30332;
  assign n30334 = controllable_hmaster1 & ~n30333;
  assign n30335 = ~n30329 & ~n30334;
  assign n30336 = ~i_hlock6 & ~n30335;
  assign n30337 = ~n30331 & ~n30336;
  assign n30338 = ~controllable_hgrant6 & ~n30337;
  assign n30339 = ~n13894 & ~n30338;
  assign n30340 = ~controllable_hmaster0 & ~n30339;
  assign n30341 = ~n30306 & ~n30340;
  assign n30342 = ~controllable_hmaster3 & ~n30341;
  assign n30343 = ~n30282 & ~n30342;
  assign n30344 = i_hlock7 & ~n30343;
  assign n30345 = i_hlock9 & ~n18540;
  assign n30346 = ~n18567 & ~n30345;
  assign n30347 = ~controllable_hgrant4 & ~n30346;
  assign n30348 = ~n12609 & ~n30347;
  assign n30349 = ~controllable_hgrant5 & ~n30348;
  assign n30350 = ~n12608 & ~n30349;
  assign n30351 = ~controllable_hmaster2 & ~n30350;
  assign n30352 = ~n29523 & ~n30351;
  assign n30353 = ~controllable_hmaster1 & ~n30352;
  assign n30354 = ~n29522 & ~n30353;
  assign n30355 = ~controllable_hgrant6 & ~n30354;
  assign n30356 = ~n13122 & ~n30355;
  assign n30357 = controllable_hmaster0 & ~n30356;
  assign n30358 = ~controllable_hgrant4 & ~n18540;
  assign n30359 = ~n13408 & ~n30358;
  assign n30360 = ~controllable_hgrant5 & ~n30359;
  assign n30361 = ~n13407 & ~n30360;
  assign n30362 = ~controllable_hmaster2 & ~n30361;
  assign n30363 = ~n29523 & ~n30362;
  assign n30364 = ~controllable_hmaster1 & ~n30363;
  assign n30365 = ~n29522 & ~n30364;
  assign n30366 = ~controllable_hgrant6 & ~n30365;
  assign n30367 = ~n13406 & ~n30366;
  assign n30368 = ~controllable_hmaster0 & ~n30367;
  assign n30369 = ~n30357 & ~n30368;
  assign n30370 = i_hlock8 & ~n30369;
  assign n30371 = ~controllable_hgrant4 & ~n18566;
  assign n30372 = ~n13429 & ~n30371;
  assign n30373 = ~controllable_hgrant5 & ~n30372;
  assign n30374 = ~n13428 & ~n30373;
  assign n30375 = ~controllable_hmaster2 & ~n30374;
  assign n30376 = ~n29523 & ~n30375;
  assign n30377 = ~controllable_hmaster1 & ~n30376;
  assign n30378 = ~n29522 & ~n30377;
  assign n30379 = ~controllable_hgrant6 & ~n30378;
  assign n30380 = ~n13427 & ~n30379;
  assign n30381 = ~controllable_hmaster0 & ~n30380;
  assign n30382 = ~n30357 & ~n30381;
  assign n30383 = ~i_hlock8 & ~n30382;
  assign n30384 = ~n30370 & ~n30383;
  assign n30385 = controllable_hmaster3 & ~n30384;
  assign n30386 = ~controllable_hgrant4 & ~n18595;
  assign n30387 = ~n13851 & ~n30386;
  assign n30388 = ~controllable_hgrant5 & ~n30387;
  assign n30389 = ~n13850 & ~n30388;
  assign n30390 = ~controllable_hmaster2 & ~n30389;
  assign n30391 = ~n28998 & ~n30390;
  assign n30392 = controllable_hmaster1 & ~n30391;
  assign n30393 = i_hlock5 & ~n30359;
  assign n30394 = ~i_hlock5 & ~n30372;
  assign n30395 = ~n30393 & ~n30394;
  assign n30396 = ~controllable_hgrant5 & ~n30395;
  assign n30397 = ~n13865 & ~n30396;
  assign n30398 = controllable_hmaster2 & ~n30397;
  assign n30399 = ~controllable_hgrant4 & ~n18625;
  assign n30400 = ~n13873 & ~n30399;
  assign n30401 = ~controllable_hgrant5 & ~n30400;
  assign n30402 = ~n13872 & ~n30401;
  assign n30403 = ~controllable_hmaster2 & ~n30402;
  assign n30404 = ~n30398 & ~n30403;
  assign n30405 = ~controllable_hmaster1 & ~n30404;
  assign n30406 = ~n30392 & ~n30405;
  assign n30407 = ~controllable_hgrant6 & ~n30406;
  assign n30408 = ~n13951 & ~n30407;
  assign n30409 = controllable_hmaster0 & ~n30408;
  assign n30410 = controllable_hmaster2 & ~n30361;
  assign n30411 = ~controllable_hgrant4 & ~n18649;
  assign n30412 = ~n13896 & ~n30411;
  assign n30413 = ~controllable_hgrant5 & ~n30412;
  assign n30414 = ~n13895 & ~n30413;
  assign n30415 = ~controllable_hmaster2 & ~n30414;
  assign n30416 = ~n30410 & ~n30415;
  assign n30417 = controllable_hmaster1 & ~n30416;
  assign n30418 = i_hlock4 & ~n18540;
  assign n30419 = ~i_hlock4 & ~n18566;
  assign n30420 = ~n30418 & ~n30419;
  assign n30421 = ~controllable_hgrant4 & ~n30420;
  assign n30422 = ~n13912 & ~n30421;
  assign n30423 = ~controllable_hgrant5 & ~n30422;
  assign n30424 = ~n13911 & ~n30423;
  assign n30425 = controllable_hmaster2 & ~n30424;
  assign n30426 = ~controllable_hgrant4 & ~n18677;
  assign n30427 = ~n13922 & ~n30426;
  assign n30428 = ~controllable_hgrant5 & ~n30427;
  assign n30429 = ~n13921 & ~n30428;
  assign n30430 = ~controllable_hmaster2 & ~n30429;
  assign n30431 = ~n30425 & ~n30430;
  assign n30432 = ~controllable_hmaster1 & ~n30431;
  assign n30433 = ~n30417 & ~n30432;
  assign n30434 = i_hlock6 & ~n30433;
  assign n30435 = controllable_hmaster2 & ~n30374;
  assign n30436 = ~n30415 & ~n30435;
  assign n30437 = controllable_hmaster1 & ~n30436;
  assign n30438 = ~n30432 & ~n30437;
  assign n30439 = ~i_hlock6 & ~n30438;
  assign n30440 = ~n30434 & ~n30439;
  assign n30441 = ~controllable_hgrant6 & ~n30440;
  assign n30442 = ~n13894 & ~n30441;
  assign n30443 = ~controllable_hmaster0 & ~n30442;
  assign n30444 = ~n30409 & ~n30443;
  assign n30445 = ~controllable_hmaster3 & ~n30444;
  assign n30446 = ~n30385 & ~n30445;
  assign n30447 = ~i_hlock7 & ~n30446;
  assign n30448 = ~n30344 & ~n30447;
  assign n30449 = i_hbusreq7 & ~n30448;
  assign n30450 = i_hbusreq8 & ~n30281;
  assign n30451 = i_hbusreq6 & ~n30251;
  assign n30452 = ~i_hbusreq9 & ~n18745;
  assign n30453 = ~n29555 & ~n30452;
  assign n30454 = ~i_hbusreq4 & ~n30453;
  assign n30455 = ~n29554 & ~n30454;
  assign n30456 = ~controllable_hgrant4 & ~n30455;
  assign n30457 = ~n13966 & ~n30456;
  assign n30458 = ~i_hbusreq5 & ~n30457;
  assign n30459 = ~n29553 & ~n30458;
  assign n30460 = ~controllable_hgrant5 & ~n30459;
  assign n30461 = ~n13965 & ~n30460;
  assign n30462 = controllable_hmaster1 & ~n30461;
  assign n30463 = controllable_hmaster2 & ~n30461;
  assign n30464 = i_hbusreq5 & ~n30245;
  assign n30465 = i_hbusreq4 & ~n30243;
  assign n30466 = i_hbusreq9 & ~n30243;
  assign n30467 = ~i_hlock9 & ~n18863;
  assign n30468 = ~n18812 & ~n30467;
  assign n30469 = ~i_hbusreq9 & ~n30468;
  assign n30470 = ~n30466 & ~n30469;
  assign n30471 = ~i_hbusreq4 & ~n30470;
  assign n30472 = ~n30465 & ~n30471;
  assign n30473 = ~controllable_hgrant4 & ~n30472;
  assign n30474 = ~n14322 & ~n30473;
  assign n30475 = ~i_hbusreq5 & ~n30474;
  assign n30476 = ~n30464 & ~n30475;
  assign n30477 = ~controllable_hgrant5 & ~n30476;
  assign n30478 = ~n14321 & ~n30477;
  assign n30479 = ~controllable_hmaster2 & ~n30478;
  assign n30480 = ~n30463 & ~n30479;
  assign n30481 = ~controllable_hmaster1 & ~n30480;
  assign n30482 = ~n30462 & ~n30481;
  assign n30483 = ~i_hbusreq6 & ~n30482;
  assign n30484 = ~n30451 & ~n30483;
  assign n30485 = ~controllable_hgrant6 & ~n30484;
  assign n30486 = ~n14320 & ~n30485;
  assign n30487 = controllable_hmaster0 & ~n30486;
  assign n30488 = i_hbusreq6 & ~n30262;
  assign n30489 = i_hbusreq5 & ~n30256;
  assign n30490 = i_hbusreq4 & ~n18534;
  assign n30491 = i_hbusreq9 & ~n18534;
  assign n30492 = ~i_hbusreq9 & ~n18811;
  assign n30493 = ~n30491 & ~n30492;
  assign n30494 = ~i_hbusreq4 & ~n30493;
  assign n30495 = ~n30490 & ~n30494;
  assign n30496 = ~controllable_hgrant4 & ~n30495;
  assign n30497 = ~n14021 & ~n30496;
  assign n30498 = ~i_hbusreq5 & ~n30497;
  assign n30499 = ~n30489 & ~n30498;
  assign n30500 = ~controllable_hgrant5 & ~n30499;
  assign n30501 = ~n14020 & ~n30500;
  assign n30502 = ~controllable_hmaster2 & ~n30501;
  assign n30503 = ~n30463 & ~n30502;
  assign n30504 = ~controllable_hmaster1 & ~n30503;
  assign n30505 = ~n30462 & ~n30504;
  assign n30506 = ~i_hbusreq6 & ~n30505;
  assign n30507 = ~n30488 & ~n30506;
  assign n30508 = ~controllable_hgrant6 & ~n30507;
  assign n30509 = ~n14019 & ~n30508;
  assign n30510 = ~controllable_hmaster0 & ~n30509;
  assign n30511 = ~n30487 & ~n30510;
  assign n30512 = i_hlock8 & ~n30511;
  assign n30513 = i_hbusreq6 & ~n30275;
  assign n30514 = i_hbusreq5 & ~n30269;
  assign n30515 = i_hbusreq4 & ~n18560;
  assign n30516 = i_hbusreq9 & ~n18560;
  assign n30517 = ~i_hbusreq9 & ~n18863;
  assign n30518 = ~n30516 & ~n30517;
  assign n30519 = ~i_hbusreq4 & ~n30518;
  assign n30520 = ~n30515 & ~n30519;
  assign n30521 = ~controllable_hgrant4 & ~n30520;
  assign n30522 = ~n14056 & ~n30521;
  assign n30523 = ~i_hbusreq5 & ~n30522;
  assign n30524 = ~n30514 & ~n30523;
  assign n30525 = ~controllable_hgrant5 & ~n30524;
  assign n30526 = ~n14055 & ~n30525;
  assign n30527 = ~controllable_hmaster2 & ~n30526;
  assign n30528 = ~n30463 & ~n30527;
  assign n30529 = ~controllable_hmaster1 & ~n30528;
  assign n30530 = ~n30462 & ~n30529;
  assign n30531 = ~i_hbusreq6 & ~n30530;
  assign n30532 = ~n30513 & ~n30531;
  assign n30533 = ~controllable_hgrant6 & ~n30532;
  assign n30534 = ~n14054 & ~n30533;
  assign n30535 = ~controllable_hmaster0 & ~n30534;
  assign n30536 = ~n30487 & ~n30535;
  assign n30537 = ~i_hlock8 & ~n30536;
  assign n30538 = ~n30512 & ~n30537;
  assign n30539 = ~i_hbusreq8 & ~n30538;
  assign n30540 = ~n30450 & ~n30539;
  assign n30541 = controllable_hmaster3 & ~n30540;
  assign n30542 = i_hbusreq8 & ~n30341;
  assign n30543 = i_hbusreq6 & ~n30303;
  assign n30544 = i_hbusreq5 & ~n30284;
  assign n30545 = i_hbusreq4 & ~n18589;
  assign n30546 = i_hbusreq9 & ~n18589;
  assign n30547 = ~i_hbusreq9 & ~n18916;
  assign n30548 = ~n30546 & ~n30547;
  assign n30549 = ~i_hbusreq4 & ~n30548;
  assign n30550 = ~n30545 & ~n30549;
  assign n30551 = ~controllable_hgrant4 & ~n30550;
  assign n30552 = ~n14099 & ~n30551;
  assign n30553 = ~i_hbusreq5 & ~n30552;
  assign n30554 = ~n30544 & ~n30553;
  assign n30555 = ~controllable_hgrant5 & ~n30554;
  assign n30556 = ~n14097 & ~n30555;
  assign n30557 = ~controllable_hmaster2 & ~n30556;
  assign n30558 = ~n29051 & ~n30557;
  assign n30559 = controllable_hmaster1 & ~n30558;
  assign n30560 = i_hbusreq5 & ~n30292;
  assign n30561 = i_hlock5 & ~n30497;
  assign n30562 = ~i_hlock5 & ~n30522;
  assign n30563 = ~n30561 & ~n30562;
  assign n30564 = ~i_hbusreq5 & ~n30563;
  assign n30565 = ~n30560 & ~n30564;
  assign n30566 = ~controllable_hgrant5 & ~n30565;
  assign n30567 = ~n14124 & ~n30566;
  assign n30568 = controllable_hmaster2 & ~n30567;
  assign n30569 = i_hbusreq5 & ~n30297;
  assign n30570 = i_hbusreq4 & ~n18617;
  assign n30571 = i_hbusreq9 & ~n18617;
  assign n30572 = ~i_hbusreq9 & ~n18965;
  assign n30573 = ~n30571 & ~n30572;
  assign n30574 = ~i_hbusreq4 & ~n30573;
  assign n30575 = ~n30570 & ~n30574;
  assign n30576 = ~controllable_hgrant4 & ~n30575;
  assign n30577 = ~n14136 & ~n30576;
  assign n30578 = ~i_hbusreq5 & ~n30577;
  assign n30579 = ~n30569 & ~n30578;
  assign n30580 = ~controllable_hgrant5 & ~n30579;
  assign n30581 = ~n14134 & ~n30580;
  assign n30582 = ~controllable_hmaster2 & ~n30581;
  assign n30583 = ~n30568 & ~n30582;
  assign n30584 = ~controllable_hmaster1 & ~n30583;
  assign n30585 = ~n30559 & ~n30584;
  assign n30586 = ~i_hbusreq6 & ~n30585;
  assign n30587 = ~n30543 & ~n30586;
  assign n30588 = ~controllable_hgrant6 & ~n30587;
  assign n30589 = ~n14756 & ~n30588;
  assign n30590 = controllable_hmaster0 & ~n30589;
  assign n30591 = i_hbusreq6 & ~n30337;
  assign n30592 = controllable_hmaster2 & ~n30501;
  assign n30593 = i_hbusreq5 & ~n30309;
  assign n30594 = i_hbusreq4 & ~n18643;
  assign n30595 = i_hbusreq9 & ~n18643;
  assign n30596 = ~i_hbusreq9 & ~n19015;
  assign n30597 = ~n30595 & ~n30596;
  assign n30598 = ~i_hbusreq4 & ~n30597;
  assign n30599 = ~n30594 & ~n30598;
  assign n30600 = ~controllable_hgrant4 & ~n30599;
  assign n30601 = ~n14177 & ~n30600;
  assign n30602 = ~i_hbusreq5 & ~n30601;
  assign n30603 = ~n30593 & ~n30602;
  assign n30604 = ~controllable_hgrant5 & ~n30603;
  assign n30605 = ~n14175 & ~n30604;
  assign n30606 = ~controllable_hmaster2 & ~n30605;
  assign n30607 = ~n30592 & ~n30606;
  assign n30608 = controllable_hmaster1 & ~n30607;
  assign n30609 = i_hbusreq5 & ~n30319;
  assign n30610 = i_hbusreq4 & ~n30317;
  assign n30611 = i_hlock4 & ~n30493;
  assign n30612 = ~i_hlock4 & ~n30518;
  assign n30613 = ~n30611 & ~n30612;
  assign n30614 = ~i_hbusreq4 & ~n30613;
  assign n30615 = ~n30610 & ~n30614;
  assign n30616 = ~controllable_hgrant4 & ~n30615;
  assign n30617 = ~n14208 & ~n30616;
  assign n30618 = ~i_hbusreq5 & ~n30617;
  assign n30619 = ~n30609 & ~n30618;
  assign n30620 = ~controllable_hgrant5 & ~n30619;
  assign n30621 = ~n14206 & ~n30620;
  assign n30622 = controllable_hmaster2 & ~n30621;
  assign n30623 = i_hbusreq5 & ~n30324;
  assign n30624 = i_hbusreq4 & ~n18671;
  assign n30625 = i_hbusreq9 & ~n18671;
  assign n30626 = ~i_hbusreq9 & ~n19096;
  assign n30627 = ~n30625 & ~n30626;
  assign n30628 = ~i_hbusreq4 & ~n30627;
  assign n30629 = ~n30624 & ~n30628;
  assign n30630 = ~controllable_hgrant4 & ~n30629;
  assign n30631 = ~n14224 & ~n30630;
  assign n30632 = ~i_hbusreq5 & ~n30631;
  assign n30633 = ~n30623 & ~n30632;
  assign n30634 = ~controllable_hgrant5 & ~n30633;
  assign n30635 = ~n14222 & ~n30634;
  assign n30636 = ~controllable_hmaster2 & ~n30635;
  assign n30637 = ~n30622 & ~n30636;
  assign n30638 = ~controllable_hmaster1 & ~n30637;
  assign n30639 = ~n30608 & ~n30638;
  assign n30640 = i_hlock6 & ~n30639;
  assign n30641 = controllable_hmaster2 & ~n30526;
  assign n30642 = ~n30606 & ~n30641;
  assign n30643 = controllable_hmaster1 & ~n30642;
  assign n30644 = ~n30638 & ~n30643;
  assign n30645 = ~i_hlock6 & ~n30644;
  assign n30646 = ~n30640 & ~n30645;
  assign n30647 = ~i_hbusreq6 & ~n30646;
  assign n30648 = ~n30591 & ~n30647;
  assign n30649 = ~controllable_hgrant6 & ~n30648;
  assign n30650 = ~n14173 & ~n30649;
  assign n30651 = ~controllable_hmaster0 & ~n30650;
  assign n30652 = ~n30590 & ~n30651;
  assign n30653 = ~i_hbusreq8 & ~n30652;
  assign n30654 = ~n30542 & ~n30653;
  assign n30655 = ~controllable_hmaster3 & ~n30654;
  assign n30656 = ~n30541 & ~n30655;
  assign n30657 = i_hlock7 & ~n30656;
  assign n30658 = i_hbusreq8 & ~n30384;
  assign n30659 = i_hbusreq6 & ~n30354;
  assign n30660 = ~i_hbusreq9 & ~n18763;
  assign n30661 = ~n29619 & ~n30660;
  assign n30662 = ~i_hbusreq4 & ~n30661;
  assign n30663 = ~n29618 & ~n30662;
  assign n30664 = ~controllable_hgrant4 & ~n30663;
  assign n30665 = ~n13966 & ~n30664;
  assign n30666 = ~i_hbusreq5 & ~n30665;
  assign n30667 = ~n29617 & ~n30666;
  assign n30668 = ~controllable_hgrant5 & ~n30667;
  assign n30669 = ~n13965 & ~n30668;
  assign n30670 = controllable_hmaster1 & ~n30669;
  assign n30671 = controllable_hmaster2 & ~n30669;
  assign n30672 = i_hbusreq5 & ~n30348;
  assign n30673 = i_hbusreq4 & ~n30346;
  assign n30674 = i_hbusreq9 & ~n30346;
  assign n30675 = i_hlock9 & ~n18825;
  assign n30676 = ~n18876 & ~n30675;
  assign n30677 = ~i_hbusreq9 & ~n30676;
  assign n30678 = ~n30674 & ~n30677;
  assign n30679 = ~i_hbusreq4 & ~n30678;
  assign n30680 = ~n30673 & ~n30679;
  assign n30681 = ~controllable_hgrant4 & ~n30680;
  assign n30682 = ~n14322 & ~n30681;
  assign n30683 = ~i_hbusreq5 & ~n30682;
  assign n30684 = ~n30672 & ~n30683;
  assign n30685 = ~controllable_hgrant5 & ~n30684;
  assign n30686 = ~n14321 & ~n30685;
  assign n30687 = ~controllable_hmaster2 & ~n30686;
  assign n30688 = ~n30671 & ~n30687;
  assign n30689 = ~controllable_hmaster1 & ~n30688;
  assign n30690 = ~n30670 & ~n30689;
  assign n30691 = ~i_hbusreq6 & ~n30690;
  assign n30692 = ~n30659 & ~n30691;
  assign n30693 = ~controllable_hgrant6 & ~n30692;
  assign n30694 = ~n14320 & ~n30693;
  assign n30695 = controllable_hmaster0 & ~n30694;
  assign n30696 = i_hbusreq6 & ~n30365;
  assign n30697 = i_hbusreq5 & ~n30359;
  assign n30698 = i_hbusreq4 & ~n18540;
  assign n30699 = i_hbusreq9 & ~n18540;
  assign n30700 = ~i_hbusreq9 & ~n18825;
  assign n30701 = ~n30699 & ~n30700;
  assign n30702 = ~i_hbusreq4 & ~n30701;
  assign n30703 = ~n30698 & ~n30702;
  assign n30704 = ~controllable_hgrant4 & ~n30703;
  assign n30705 = ~n14021 & ~n30704;
  assign n30706 = ~i_hbusreq5 & ~n30705;
  assign n30707 = ~n30697 & ~n30706;
  assign n30708 = ~controllable_hgrant5 & ~n30707;
  assign n30709 = ~n14020 & ~n30708;
  assign n30710 = ~controllable_hmaster2 & ~n30709;
  assign n30711 = ~n30671 & ~n30710;
  assign n30712 = ~controllable_hmaster1 & ~n30711;
  assign n30713 = ~n30670 & ~n30712;
  assign n30714 = ~i_hbusreq6 & ~n30713;
  assign n30715 = ~n30696 & ~n30714;
  assign n30716 = ~controllable_hgrant6 & ~n30715;
  assign n30717 = ~n14019 & ~n30716;
  assign n30718 = ~controllable_hmaster0 & ~n30717;
  assign n30719 = ~n30695 & ~n30718;
  assign n30720 = i_hlock8 & ~n30719;
  assign n30721 = i_hbusreq6 & ~n30378;
  assign n30722 = i_hbusreq5 & ~n30372;
  assign n30723 = i_hbusreq4 & ~n18566;
  assign n30724 = i_hbusreq9 & ~n18566;
  assign n30725 = ~i_hbusreq9 & ~n18875;
  assign n30726 = ~n30724 & ~n30725;
  assign n30727 = ~i_hbusreq4 & ~n30726;
  assign n30728 = ~n30723 & ~n30727;
  assign n30729 = ~controllable_hgrant4 & ~n30728;
  assign n30730 = ~n14056 & ~n30729;
  assign n30731 = ~i_hbusreq5 & ~n30730;
  assign n30732 = ~n30722 & ~n30731;
  assign n30733 = ~controllable_hgrant5 & ~n30732;
  assign n30734 = ~n14055 & ~n30733;
  assign n30735 = ~controllable_hmaster2 & ~n30734;
  assign n30736 = ~n30671 & ~n30735;
  assign n30737 = ~controllable_hmaster1 & ~n30736;
  assign n30738 = ~n30670 & ~n30737;
  assign n30739 = ~i_hbusreq6 & ~n30738;
  assign n30740 = ~n30721 & ~n30739;
  assign n30741 = ~controllable_hgrant6 & ~n30740;
  assign n30742 = ~n14054 & ~n30741;
  assign n30743 = ~controllable_hmaster0 & ~n30742;
  assign n30744 = ~n30695 & ~n30743;
  assign n30745 = ~i_hlock8 & ~n30744;
  assign n30746 = ~n30720 & ~n30745;
  assign n30747 = ~i_hbusreq8 & ~n30746;
  assign n30748 = ~n30658 & ~n30747;
  assign n30749 = controllable_hmaster3 & ~n30748;
  assign n30750 = i_hbusreq8 & ~n30444;
  assign n30751 = i_hbusreq6 & ~n30406;
  assign n30752 = i_hbusreq5 & ~n30387;
  assign n30753 = i_hbusreq4 & ~n18595;
  assign n30754 = i_hbusreq9 & ~n18595;
  assign n30755 = ~i_hbusreq9 & ~n18925;
  assign n30756 = ~n30754 & ~n30755;
  assign n30757 = ~i_hbusreq4 & ~n30756;
  assign n30758 = ~n30753 & ~n30757;
  assign n30759 = ~controllable_hgrant4 & ~n30758;
  assign n30760 = ~n14099 & ~n30759;
  assign n30761 = ~i_hbusreq5 & ~n30760;
  assign n30762 = ~n30752 & ~n30761;
  assign n30763 = ~controllable_hgrant5 & ~n30762;
  assign n30764 = ~n14097 & ~n30763;
  assign n30765 = ~controllable_hmaster2 & ~n30764;
  assign n30766 = ~n29106 & ~n30765;
  assign n30767 = controllable_hmaster1 & ~n30766;
  assign n30768 = i_hbusreq5 & ~n30395;
  assign n30769 = i_hlock5 & ~n30705;
  assign n30770 = ~i_hlock5 & ~n30730;
  assign n30771 = ~n30769 & ~n30770;
  assign n30772 = ~i_hbusreq5 & ~n30771;
  assign n30773 = ~n30768 & ~n30772;
  assign n30774 = ~controllable_hgrant5 & ~n30773;
  assign n30775 = ~n14124 & ~n30774;
  assign n30776 = controllable_hmaster2 & ~n30775;
  assign n30777 = i_hbusreq5 & ~n30400;
  assign n30778 = i_hbusreq4 & ~n18625;
  assign n30779 = i_hbusreq9 & ~n18625;
  assign n30780 = ~i_hbusreq9 & ~n18979;
  assign n30781 = ~n30779 & ~n30780;
  assign n30782 = ~i_hbusreq4 & ~n30781;
  assign n30783 = ~n30778 & ~n30782;
  assign n30784 = ~controllable_hgrant4 & ~n30783;
  assign n30785 = ~n14136 & ~n30784;
  assign n30786 = ~i_hbusreq5 & ~n30785;
  assign n30787 = ~n30777 & ~n30786;
  assign n30788 = ~controllable_hgrant5 & ~n30787;
  assign n30789 = ~n14134 & ~n30788;
  assign n30790 = ~controllable_hmaster2 & ~n30789;
  assign n30791 = ~n30776 & ~n30790;
  assign n30792 = ~controllable_hmaster1 & ~n30791;
  assign n30793 = ~n30767 & ~n30792;
  assign n30794 = ~i_hbusreq6 & ~n30793;
  assign n30795 = ~n30751 & ~n30794;
  assign n30796 = ~controllable_hgrant6 & ~n30795;
  assign n30797 = ~n14772 & ~n30796;
  assign n30798 = controllable_hmaster0 & ~n30797;
  assign n30799 = i_hbusreq6 & ~n30440;
  assign n30800 = controllable_hmaster2 & ~n30709;
  assign n30801 = i_hbusreq5 & ~n30412;
  assign n30802 = i_hbusreq4 & ~n18649;
  assign n30803 = i_hbusreq9 & ~n18649;
  assign n30804 = ~i_hbusreq9 & ~n19027;
  assign n30805 = ~n30803 & ~n30804;
  assign n30806 = ~i_hbusreq4 & ~n30805;
  assign n30807 = ~n30802 & ~n30806;
  assign n30808 = ~controllable_hgrant4 & ~n30807;
  assign n30809 = ~n14177 & ~n30808;
  assign n30810 = ~i_hbusreq5 & ~n30809;
  assign n30811 = ~n30801 & ~n30810;
  assign n30812 = ~controllable_hgrant5 & ~n30811;
  assign n30813 = ~n14175 & ~n30812;
  assign n30814 = ~controllable_hmaster2 & ~n30813;
  assign n30815 = ~n30800 & ~n30814;
  assign n30816 = controllable_hmaster1 & ~n30815;
  assign n30817 = i_hbusreq5 & ~n30422;
  assign n30818 = i_hbusreq4 & ~n30420;
  assign n30819 = i_hlock4 & ~n30701;
  assign n30820 = ~i_hlock4 & ~n30726;
  assign n30821 = ~n30819 & ~n30820;
  assign n30822 = ~i_hbusreq4 & ~n30821;
  assign n30823 = ~n30818 & ~n30822;
  assign n30824 = ~controllable_hgrant4 & ~n30823;
  assign n30825 = ~n14208 & ~n30824;
  assign n30826 = ~i_hbusreq5 & ~n30825;
  assign n30827 = ~n30817 & ~n30826;
  assign n30828 = ~controllable_hgrant5 & ~n30827;
  assign n30829 = ~n14206 & ~n30828;
  assign n30830 = controllable_hmaster2 & ~n30829;
  assign n30831 = i_hbusreq5 & ~n30427;
  assign n30832 = i_hbusreq4 & ~n18677;
  assign n30833 = i_hbusreq9 & ~n18677;
  assign n30834 = ~i_hbusreq9 & ~n19116;
  assign n30835 = ~n30833 & ~n30834;
  assign n30836 = ~i_hbusreq4 & ~n30835;
  assign n30837 = ~n30832 & ~n30836;
  assign n30838 = ~controllable_hgrant4 & ~n30837;
  assign n30839 = ~n14224 & ~n30838;
  assign n30840 = ~i_hbusreq5 & ~n30839;
  assign n30841 = ~n30831 & ~n30840;
  assign n30842 = ~controllable_hgrant5 & ~n30841;
  assign n30843 = ~n14222 & ~n30842;
  assign n30844 = ~controllable_hmaster2 & ~n30843;
  assign n30845 = ~n30830 & ~n30844;
  assign n30846 = ~controllable_hmaster1 & ~n30845;
  assign n30847 = ~n30816 & ~n30846;
  assign n30848 = i_hlock6 & ~n30847;
  assign n30849 = controllable_hmaster2 & ~n30734;
  assign n30850 = ~n30814 & ~n30849;
  assign n30851 = controllable_hmaster1 & ~n30850;
  assign n30852 = ~n30846 & ~n30851;
  assign n30853 = ~i_hlock6 & ~n30852;
  assign n30854 = ~n30848 & ~n30853;
  assign n30855 = ~i_hbusreq6 & ~n30854;
  assign n30856 = ~n30799 & ~n30855;
  assign n30857 = ~controllable_hgrant6 & ~n30856;
  assign n30858 = ~n14173 & ~n30857;
  assign n30859 = ~controllable_hmaster0 & ~n30858;
  assign n30860 = ~n30798 & ~n30859;
  assign n30861 = ~i_hbusreq8 & ~n30860;
  assign n30862 = ~n30750 & ~n30861;
  assign n30863 = ~controllable_hmaster3 & ~n30862;
  assign n30864 = ~n30749 & ~n30863;
  assign n30865 = ~i_hlock7 & ~n30864;
  assign n30866 = ~n30657 & ~n30865;
  assign n30867 = ~i_hbusreq7 & ~n30866;
  assign n30868 = ~n30449 & ~n30867;
  assign n30869 = n7924 & ~n30868;
  assign n30870 = ~n30241 & ~n30869;
  assign n30871 = ~n8214 & ~n30870;
  assign n30872 = ~n20274 & ~n30011;
  assign n30873 = i_hlock8 & ~n30872;
  assign n30874 = ~n20283 & ~n30011;
  assign n30875 = ~i_hlock8 & ~n30874;
  assign n30876 = ~n30873 & ~n30875;
  assign n30877 = controllable_hmaster3 & ~n30876;
  assign n30878 = ~n20499 & ~n29741;
  assign n30879 = ~controllable_hmaster3 & ~n30878;
  assign n30880 = ~n30877 & ~n30879;
  assign n30881 = i_hlock7 & ~n30880;
  assign n30882 = ~n20499 & ~n29756;
  assign n30883 = ~controllable_hmaster3 & ~n30882;
  assign n30884 = ~n30877 & ~n30883;
  assign n30885 = ~i_hlock7 & ~n30884;
  assign n30886 = ~n30881 & ~n30885;
  assign n30887 = i_hbusreq7 & ~n30886;
  assign n30888 = i_hbusreq8 & ~n30876;
  assign n30889 = ~n20320 & ~n30050;
  assign n30890 = i_hlock8 & ~n30889;
  assign n30891 = ~n20332 & ~n30050;
  assign n30892 = ~i_hlock8 & ~n30891;
  assign n30893 = ~n30890 & ~n30892;
  assign n30894 = ~i_hbusreq8 & ~n30893;
  assign n30895 = ~n30888 & ~n30894;
  assign n30896 = controllable_hmaster3 & ~n30895;
  assign n30897 = i_hbusreq8 & ~n30878;
  assign n30898 = ~n20525 & ~n29804;
  assign n30899 = ~i_hbusreq8 & ~n30898;
  assign n30900 = ~n30897 & ~n30899;
  assign n30901 = ~controllable_hmaster3 & ~n30900;
  assign n30902 = ~n30896 & ~n30901;
  assign n30903 = i_hlock7 & ~n30902;
  assign n30904 = i_hbusreq8 & ~n30882;
  assign n30905 = ~n20525 & ~n29834;
  assign n30906 = ~i_hbusreq8 & ~n30905;
  assign n30907 = ~n30904 & ~n30906;
  assign n30908 = ~controllable_hmaster3 & ~n30907;
  assign n30909 = ~n30896 & ~n30908;
  assign n30910 = ~i_hlock7 & ~n30909;
  assign n30911 = ~n30903 & ~n30910;
  assign n30912 = ~i_hbusreq7 & ~n30911;
  assign n30913 = ~n30887 & ~n30912;
  assign n30914 = ~n7924 & ~n30913;
  assign n30915 = ~n20381 & ~n30080;
  assign n30916 = i_hlock8 & ~n30915;
  assign n30917 = ~n20390 & ~n30080;
  assign n30918 = ~i_hlock8 & ~n30917;
  assign n30919 = ~n30916 & ~n30918;
  assign n30920 = controllable_hmaster3 & ~n30919;
  assign n30921 = ~n20554 & ~n29875;
  assign n30922 = ~controllable_hmaster3 & ~n30921;
  assign n30923 = ~n30920 & ~n30922;
  assign n30924 = i_hlock7 & ~n30923;
  assign n30925 = ~n20554 & ~n29890;
  assign n30926 = ~controllable_hmaster3 & ~n30925;
  assign n30927 = ~n30920 & ~n30926;
  assign n30928 = ~i_hlock7 & ~n30927;
  assign n30929 = ~n30924 & ~n30928;
  assign n30930 = i_hbusreq7 & ~n30929;
  assign n30931 = i_hbusreq8 & ~n30919;
  assign n30932 = ~n20429 & ~n30119;
  assign n30933 = i_hlock8 & ~n30932;
  assign n30934 = ~n20441 & ~n30119;
  assign n30935 = ~i_hlock8 & ~n30934;
  assign n30936 = ~n30933 & ~n30935;
  assign n30937 = ~i_hbusreq8 & ~n30936;
  assign n30938 = ~n30931 & ~n30937;
  assign n30939 = controllable_hmaster3 & ~n30938;
  assign n30940 = i_hbusreq8 & ~n30921;
  assign n30941 = ~n20580 & ~n29955;
  assign n30942 = ~i_hbusreq8 & ~n30941;
  assign n30943 = ~n30940 & ~n30942;
  assign n30944 = ~controllable_hmaster3 & ~n30943;
  assign n30945 = ~n30939 & ~n30944;
  assign n30946 = i_hlock7 & ~n30945;
  assign n30947 = i_hbusreq8 & ~n30925;
  assign n30948 = ~n20580 & ~n29985;
  assign n30949 = ~i_hbusreq8 & ~n30948;
  assign n30950 = ~n30947 & ~n30949;
  assign n30951 = ~controllable_hmaster3 & ~n30950;
  assign n30952 = ~n30939 & ~n30951;
  assign n30953 = ~i_hlock7 & ~n30952;
  assign n30954 = ~n30946 & ~n30953;
  assign n30955 = ~i_hbusreq7 & ~n30954;
  assign n30956 = ~n30930 & ~n30955;
  assign n30957 = n7924 & ~n30956;
  assign n30958 = ~n30914 & ~n30957;
  assign n30959 = n8214 & ~n30958;
  assign n30960 = ~n30871 & ~n30959;
  assign n30961 = n8202 & ~n30960;
  assign n30962 = ~n30139 & ~n30961;
  assign n30963 = n7920 & ~n30962;
  assign n30964 = ~n29136 & ~n30963;
  assign n30965 = ~n7728 & ~n30964;
  assign n30966 = ~n29718 & ~n30965;
  assign n30967 = n7723 & ~n30966;
  assign n30968 = ~n7723 & ~n30964;
  assign n30969 = ~n30967 & ~n30968;
  assign n30970 = n7714 & ~n30969;
  assign n30971 = n7723 & ~n30964;
  assign n30972 = ~controllable_hgrant4 & ~n20622;
  assign n30973 = ~n13153 & ~n30972;
  assign n30974 = ~controllable_hgrant5 & ~n30973;
  assign n30975 = ~n13152 & ~n30974;
  assign n30976 = controllable_hmaster1 & ~n30975;
  assign n30977 = controllable_hmaster2 & ~n30975;
  assign n30978 = ~n30248 & ~n30977;
  assign n30979 = ~controllable_hmaster1 & ~n30978;
  assign n30980 = ~n30976 & ~n30979;
  assign n30981 = ~controllable_hgrant6 & ~n30980;
  assign n30982 = ~n13122 & ~n30981;
  assign n30983 = controllable_hmaster0 & ~n30982;
  assign n30984 = ~controllable_hgrant4 & ~n20705;
  assign n30985 = ~n13408 & ~n30984;
  assign n30986 = ~controllable_hgrant5 & ~n30985;
  assign n30987 = ~n13407 & ~n30986;
  assign n30988 = ~controllable_hmaster2 & ~n30987;
  assign n30989 = ~n30977 & ~n30988;
  assign n30990 = ~controllable_hmaster1 & ~n30989;
  assign n30991 = ~n30976 & ~n30990;
  assign n30992 = ~controllable_hgrant6 & ~n30991;
  assign n30993 = ~n13406 & ~n30992;
  assign n30994 = ~controllable_hmaster0 & ~n30993;
  assign n30995 = ~n30983 & ~n30994;
  assign n30996 = i_hlock8 & ~n30995;
  assign n30997 = ~controllable_hgrant4 & ~n20747;
  assign n30998 = ~n13429 & ~n30997;
  assign n30999 = ~controllable_hgrant5 & ~n30998;
  assign n31000 = ~n13428 & ~n30999;
  assign n31001 = ~controllable_hmaster2 & ~n31000;
  assign n31002 = ~n30977 & ~n31001;
  assign n31003 = ~controllable_hmaster1 & ~n31002;
  assign n31004 = ~n30976 & ~n31003;
  assign n31005 = ~controllable_hgrant6 & ~n31004;
  assign n31006 = ~n13427 & ~n31005;
  assign n31007 = ~controllable_hmaster0 & ~n31006;
  assign n31008 = ~n30983 & ~n31007;
  assign n31009 = ~i_hlock8 & ~n31008;
  assign n31010 = ~n30996 & ~n31009;
  assign n31011 = controllable_hmaster3 & ~n31010;
  assign n31012 = ~controllable_hgrant4 & ~n20654;
  assign n31013 = ~n13408 & ~n31012;
  assign n31014 = ~controllable_hgrant5 & ~n31013;
  assign n31015 = ~n13407 & ~n31014;
  assign n31016 = controllable_hmaster2 & ~n31015;
  assign n31017 = ~controllable_hgrant4 & ~n20726;
  assign n31018 = ~n13851 & ~n31017;
  assign n31019 = ~controllable_hgrant5 & ~n31018;
  assign n31020 = ~n13850 & ~n31019;
  assign n31021 = ~controllable_hmaster2 & ~n31020;
  assign n31022 = ~n31016 & ~n31021;
  assign n31023 = controllable_hmaster1 & ~n31022;
  assign n31024 = i_hlock5 & ~n30985;
  assign n31025 = ~i_hlock5 & ~n30998;
  assign n31026 = ~n31024 & ~n31025;
  assign n31027 = ~controllable_hgrant5 & ~n31026;
  assign n31028 = ~n13865 & ~n31027;
  assign n31029 = controllable_hmaster2 & ~n31028;
  assign n31030 = ~controllable_hgrant4 & ~n20766;
  assign n31031 = ~n13873 & ~n31030;
  assign n31032 = ~controllable_hgrant5 & ~n31031;
  assign n31033 = ~n13872 & ~n31032;
  assign n31034 = ~controllable_hmaster2 & ~n31033;
  assign n31035 = ~n31029 & ~n31034;
  assign n31036 = ~controllable_hmaster1 & ~n31035;
  assign n31037 = ~n31023 & ~n31036;
  assign n31038 = ~controllable_hgrant6 & ~n31037;
  assign n31039 = ~n13849 & ~n31038;
  assign n31040 = controllable_hmaster0 & ~n31039;
  assign n31041 = controllable_hmaster2 & ~n30987;
  assign n31042 = ~controllable_hgrant4 & ~n20792;
  assign n31043 = ~n13896 & ~n31042;
  assign n31044 = ~controllable_hgrant5 & ~n31043;
  assign n31045 = ~n13895 & ~n31044;
  assign n31046 = ~controllable_hmaster2 & ~n31045;
  assign n31047 = ~n31041 & ~n31046;
  assign n31048 = controllable_hmaster1 & ~n31047;
  assign n31049 = i_hlock4 & ~n20705;
  assign n31050 = ~i_hlock4 & ~n20747;
  assign n31051 = ~n31049 & ~n31050;
  assign n31052 = ~controllable_hgrant4 & ~n31051;
  assign n31053 = ~n13912 & ~n31052;
  assign n31054 = ~controllable_hgrant5 & ~n31053;
  assign n31055 = ~n13911 & ~n31054;
  assign n31056 = controllable_hmaster2 & ~n31055;
  assign n31057 = ~controllable_hgrant4 & ~n20820;
  assign n31058 = ~n13922 & ~n31057;
  assign n31059 = ~controllable_hgrant5 & ~n31058;
  assign n31060 = ~n13921 & ~n31059;
  assign n31061 = ~controllable_hmaster2 & ~n31060;
  assign n31062 = ~n31056 & ~n31061;
  assign n31063 = ~controllable_hmaster1 & ~n31062;
  assign n31064 = ~n31048 & ~n31063;
  assign n31065 = i_hlock6 & ~n31064;
  assign n31066 = controllable_hmaster2 & ~n31000;
  assign n31067 = ~n31046 & ~n31066;
  assign n31068 = controllable_hmaster1 & ~n31067;
  assign n31069 = ~n31063 & ~n31068;
  assign n31070 = ~i_hlock6 & ~n31069;
  assign n31071 = ~n31065 & ~n31070;
  assign n31072 = ~controllable_hgrant6 & ~n31071;
  assign n31073 = ~n13894 & ~n31072;
  assign n31074 = ~controllable_hmaster0 & ~n31073;
  assign n31075 = ~n31040 & ~n31074;
  assign n31076 = ~controllable_hmaster3 & ~n31075;
  assign n31077 = ~n31011 & ~n31076;
  assign n31078 = i_hlock7 & ~n31077;
  assign n31079 = ~controllable_hgrant4 & ~n20635;
  assign n31080 = ~n13153 & ~n31079;
  assign n31081 = ~controllable_hgrant5 & ~n31080;
  assign n31082 = ~n13152 & ~n31081;
  assign n31083 = controllable_hmaster1 & ~n31082;
  assign n31084 = controllable_hmaster2 & ~n31082;
  assign n31085 = ~n30351 & ~n31084;
  assign n31086 = ~controllable_hmaster1 & ~n31085;
  assign n31087 = ~n31083 & ~n31086;
  assign n31088 = ~controllable_hgrant6 & ~n31087;
  assign n31089 = ~n13122 & ~n31088;
  assign n31090 = controllable_hmaster0 & ~n31089;
  assign n31091 = ~controllable_hgrant4 & ~n20711;
  assign n31092 = ~n13408 & ~n31091;
  assign n31093 = ~controllable_hgrant5 & ~n31092;
  assign n31094 = ~n13407 & ~n31093;
  assign n31095 = ~controllable_hmaster2 & ~n31094;
  assign n31096 = ~n31084 & ~n31095;
  assign n31097 = ~controllable_hmaster1 & ~n31096;
  assign n31098 = ~n31083 & ~n31097;
  assign n31099 = ~controllable_hgrant6 & ~n31098;
  assign n31100 = ~n13406 & ~n31099;
  assign n31101 = ~controllable_hmaster0 & ~n31100;
  assign n31102 = ~n31090 & ~n31101;
  assign n31103 = i_hlock8 & ~n31102;
  assign n31104 = ~controllable_hgrant4 & ~n20750;
  assign n31105 = ~n13429 & ~n31104;
  assign n31106 = ~controllable_hgrant5 & ~n31105;
  assign n31107 = ~n13428 & ~n31106;
  assign n31108 = ~controllable_hmaster2 & ~n31107;
  assign n31109 = ~n31084 & ~n31108;
  assign n31110 = ~controllable_hmaster1 & ~n31109;
  assign n31111 = ~n31083 & ~n31110;
  assign n31112 = ~controllable_hgrant6 & ~n31111;
  assign n31113 = ~n13427 & ~n31112;
  assign n31114 = ~controllable_hmaster0 & ~n31113;
  assign n31115 = ~n31090 & ~n31114;
  assign n31116 = ~i_hlock8 & ~n31115;
  assign n31117 = ~n31103 & ~n31116;
  assign n31118 = controllable_hmaster3 & ~n31117;
  assign n31119 = ~controllable_hgrant4 & ~n20669;
  assign n31120 = ~n13429 & ~n31119;
  assign n31121 = ~controllable_hgrant5 & ~n31120;
  assign n31122 = ~n13428 & ~n31121;
  assign n31123 = controllable_hmaster2 & ~n31122;
  assign n31124 = ~controllable_hgrant4 & ~n20735;
  assign n31125 = ~n13851 & ~n31124;
  assign n31126 = ~controllable_hgrant5 & ~n31125;
  assign n31127 = ~n13850 & ~n31126;
  assign n31128 = ~controllable_hmaster2 & ~n31127;
  assign n31129 = ~n31123 & ~n31128;
  assign n31130 = controllable_hmaster1 & ~n31129;
  assign n31131 = i_hlock5 & ~n31092;
  assign n31132 = ~i_hlock5 & ~n31105;
  assign n31133 = ~n31131 & ~n31132;
  assign n31134 = ~controllable_hgrant5 & ~n31133;
  assign n31135 = ~n13865 & ~n31134;
  assign n31136 = controllable_hmaster2 & ~n31135;
  assign n31137 = ~controllable_hgrant4 & ~n20774;
  assign n31138 = ~n13873 & ~n31137;
  assign n31139 = ~controllable_hgrant5 & ~n31138;
  assign n31140 = ~n13872 & ~n31139;
  assign n31141 = ~controllable_hmaster2 & ~n31140;
  assign n31142 = ~n31136 & ~n31141;
  assign n31143 = ~controllable_hmaster1 & ~n31142;
  assign n31144 = ~n31130 & ~n31143;
  assign n31145 = ~controllable_hgrant6 & ~n31144;
  assign n31146 = ~n13951 & ~n31145;
  assign n31147 = controllable_hmaster0 & ~n31146;
  assign n31148 = controllable_hmaster2 & ~n31094;
  assign n31149 = ~controllable_hgrant4 & ~n20798;
  assign n31150 = ~n13896 & ~n31149;
  assign n31151 = ~controllable_hgrant5 & ~n31150;
  assign n31152 = ~n13895 & ~n31151;
  assign n31153 = ~controllable_hmaster2 & ~n31152;
  assign n31154 = ~n31148 & ~n31153;
  assign n31155 = controllable_hmaster1 & ~n31154;
  assign n31156 = i_hlock4 & ~n20711;
  assign n31157 = ~i_hlock4 & ~n20750;
  assign n31158 = ~n31156 & ~n31157;
  assign n31159 = ~controllable_hgrant4 & ~n31158;
  assign n31160 = ~n13912 & ~n31159;
  assign n31161 = ~controllable_hgrant5 & ~n31160;
  assign n31162 = ~n13911 & ~n31161;
  assign n31163 = controllable_hmaster2 & ~n31162;
  assign n31164 = ~controllable_hgrant4 & ~n20826;
  assign n31165 = ~n13922 & ~n31164;
  assign n31166 = ~controllable_hgrant5 & ~n31165;
  assign n31167 = ~n13921 & ~n31166;
  assign n31168 = ~controllable_hmaster2 & ~n31167;
  assign n31169 = ~n31163 & ~n31168;
  assign n31170 = ~controllable_hmaster1 & ~n31169;
  assign n31171 = ~n31155 & ~n31170;
  assign n31172 = i_hlock6 & ~n31171;
  assign n31173 = controllable_hmaster2 & ~n31107;
  assign n31174 = ~n31153 & ~n31173;
  assign n31175 = controllable_hmaster1 & ~n31174;
  assign n31176 = ~n31170 & ~n31175;
  assign n31177 = ~i_hlock6 & ~n31176;
  assign n31178 = ~n31172 & ~n31177;
  assign n31179 = ~controllable_hgrant6 & ~n31178;
  assign n31180 = ~n13894 & ~n31179;
  assign n31181 = ~controllable_hmaster0 & ~n31180;
  assign n31182 = ~n31147 & ~n31181;
  assign n31183 = ~controllable_hmaster3 & ~n31182;
  assign n31184 = ~n31118 & ~n31183;
  assign n31185 = ~i_hlock7 & ~n31184;
  assign n31186 = ~n31078 & ~n31185;
  assign n31187 = i_hbusreq7 & ~n31186;
  assign n31188 = i_hbusreq8 & ~n31010;
  assign n31189 = i_hbusreq6 & ~n30980;
  assign n31190 = i_hbusreq5 & ~n30973;
  assign n31191 = i_hbusreq4 & ~n20622;
  assign n31192 = i_hbusreq9 & ~n20622;
  assign n31193 = ~i_hbusreq9 & ~n20895;
  assign n31194 = ~n31192 & ~n31193;
  assign n31195 = ~i_hbusreq4 & ~n31194;
  assign n31196 = ~n31191 & ~n31195;
  assign n31197 = ~controllable_hgrant4 & ~n31196;
  assign n31198 = ~n13966 & ~n31197;
  assign n31199 = ~i_hbusreq5 & ~n31198;
  assign n31200 = ~n31190 & ~n31199;
  assign n31201 = ~controllable_hgrant5 & ~n31200;
  assign n31202 = ~n13965 & ~n31201;
  assign n31203 = controllable_hmaster1 & ~n31202;
  assign n31204 = controllable_hmaster2 & ~n31202;
  assign n31205 = ~i_hlock9 & ~n21081;
  assign n31206 = ~n21031 & ~n31205;
  assign n31207 = ~i_hbusreq9 & ~n31206;
  assign n31208 = ~n30466 & ~n31207;
  assign n31209 = ~i_hbusreq4 & ~n31208;
  assign n31210 = ~n30465 & ~n31209;
  assign n31211 = ~controllable_hgrant4 & ~n31210;
  assign n31212 = ~n12676 & ~n31211;
  assign n31213 = ~i_hbusreq5 & ~n31212;
  assign n31214 = ~n30464 & ~n31213;
  assign n31215 = ~controllable_hgrant5 & ~n31214;
  assign n31216 = ~n12674 & ~n31215;
  assign n31217 = ~controllable_hmaster2 & ~n31216;
  assign n31218 = ~n31204 & ~n31217;
  assign n31219 = ~controllable_hmaster1 & ~n31218;
  assign n31220 = ~n31203 & ~n31219;
  assign n31221 = ~i_hbusreq6 & ~n31220;
  assign n31222 = ~n31189 & ~n31221;
  assign n31223 = ~controllable_hgrant6 & ~n31222;
  assign n31224 = ~n13818 & ~n31223;
  assign n31225 = controllable_hmaster0 & ~n31224;
  assign n31226 = i_hbusreq6 & ~n30991;
  assign n31227 = i_hbusreq5 & ~n30985;
  assign n31228 = i_hbusreq4 & ~n20705;
  assign n31229 = i_hbusreq9 & ~n20705;
  assign n31230 = ~i_hbusreq9 & ~n21134;
  assign n31231 = ~n31229 & ~n31230;
  assign n31232 = ~i_hbusreq4 & ~n31231;
  assign n31233 = ~n31228 & ~n31232;
  assign n31234 = ~controllable_hgrant4 & ~n31233;
  assign n31235 = ~n14021 & ~n31234;
  assign n31236 = ~i_hbusreq5 & ~n31235;
  assign n31237 = ~n31227 & ~n31236;
  assign n31238 = ~controllable_hgrant5 & ~n31237;
  assign n31239 = ~n14020 & ~n31238;
  assign n31240 = ~controllable_hmaster2 & ~n31239;
  assign n31241 = ~n31204 & ~n31240;
  assign n31242 = ~controllable_hmaster1 & ~n31241;
  assign n31243 = ~n31203 & ~n31242;
  assign n31244 = ~i_hbusreq6 & ~n31243;
  assign n31245 = ~n31226 & ~n31244;
  assign n31246 = ~controllable_hgrant6 & ~n31245;
  assign n31247 = ~n14019 & ~n31246;
  assign n31248 = ~controllable_hmaster0 & ~n31247;
  assign n31249 = ~n31225 & ~n31248;
  assign n31250 = i_hlock8 & ~n31249;
  assign n31251 = i_hbusreq6 & ~n31004;
  assign n31252 = i_hbusreq5 & ~n30998;
  assign n31253 = i_hbusreq4 & ~n20747;
  assign n31254 = i_hbusreq9 & ~n20747;
  assign n31255 = ~i_hbusreq9 & ~n21215;
  assign n31256 = ~n31254 & ~n31255;
  assign n31257 = ~i_hbusreq4 & ~n31256;
  assign n31258 = ~n31253 & ~n31257;
  assign n31259 = ~controllable_hgrant4 & ~n31258;
  assign n31260 = ~n14056 & ~n31259;
  assign n31261 = ~i_hbusreq5 & ~n31260;
  assign n31262 = ~n31252 & ~n31261;
  assign n31263 = ~controllable_hgrant5 & ~n31262;
  assign n31264 = ~n14055 & ~n31263;
  assign n31265 = ~controllable_hmaster2 & ~n31264;
  assign n31266 = ~n31204 & ~n31265;
  assign n31267 = ~controllable_hmaster1 & ~n31266;
  assign n31268 = ~n31203 & ~n31267;
  assign n31269 = ~i_hbusreq6 & ~n31268;
  assign n31270 = ~n31251 & ~n31269;
  assign n31271 = ~controllable_hgrant6 & ~n31270;
  assign n31272 = ~n14054 & ~n31271;
  assign n31273 = ~controllable_hmaster0 & ~n31272;
  assign n31274 = ~n31225 & ~n31273;
  assign n31275 = ~i_hlock8 & ~n31274;
  assign n31276 = ~n31250 & ~n31275;
  assign n31277 = ~i_hbusreq8 & ~n31276;
  assign n31278 = ~n31188 & ~n31277;
  assign n31279 = controllable_hmaster3 & ~n31278;
  assign n31280 = i_hbusreq8 & ~n31075;
  assign n31281 = i_hbusreq6 & ~n31037;
  assign n31282 = i_hbusreq5 & ~n31013;
  assign n31283 = i_hbusreq4 & ~n20654;
  assign n31284 = i_hbusreq9 & ~n20654;
  assign n31285 = ~i_hbusreq9 & ~n20963;
  assign n31286 = ~n31284 & ~n31285;
  assign n31287 = ~i_hbusreq4 & ~n31286;
  assign n31288 = ~n31283 & ~n31287;
  assign n31289 = ~controllable_hgrant4 & ~n31288;
  assign n31290 = ~n14021 & ~n31289;
  assign n31291 = ~i_hbusreq5 & ~n31290;
  assign n31292 = ~n31282 & ~n31291;
  assign n31293 = ~controllable_hgrant5 & ~n31292;
  assign n31294 = ~n14020 & ~n31293;
  assign n31295 = controllable_hmaster2 & ~n31294;
  assign n31296 = i_hbusreq5 & ~n31018;
  assign n31297 = i_hbusreq4 & ~n20726;
  assign n31298 = i_hbusreq9 & ~n20726;
  assign n31299 = ~i_hbusreq9 & ~n21176;
  assign n31300 = ~n31298 & ~n31299;
  assign n31301 = ~i_hbusreq4 & ~n31300;
  assign n31302 = ~n31297 & ~n31301;
  assign n31303 = ~controllable_hgrant4 & ~n31302;
  assign n31304 = ~n14099 & ~n31303;
  assign n31305 = ~i_hbusreq5 & ~n31304;
  assign n31306 = ~n31296 & ~n31305;
  assign n31307 = ~controllable_hgrant5 & ~n31306;
  assign n31308 = ~n14097 & ~n31307;
  assign n31309 = ~controllable_hmaster2 & ~n31308;
  assign n31310 = ~n31295 & ~n31309;
  assign n31311 = controllable_hmaster1 & ~n31310;
  assign n31312 = i_hbusreq5 & ~n31026;
  assign n31313 = i_hlock5 & ~n31235;
  assign n31314 = ~i_hlock5 & ~n31260;
  assign n31315 = ~n31313 & ~n31314;
  assign n31316 = ~i_hbusreq5 & ~n31315;
  assign n31317 = ~n31312 & ~n31316;
  assign n31318 = ~controllable_hgrant5 & ~n31317;
  assign n31319 = ~n14124 & ~n31318;
  assign n31320 = controllable_hmaster2 & ~n31319;
  assign n31321 = i_hbusreq5 & ~n31031;
  assign n31322 = i_hbusreq4 & ~n20766;
  assign n31323 = i_hbusreq9 & ~n20766;
  assign n31324 = ~i_hbusreq9 & ~n21252;
  assign n31325 = ~n31323 & ~n31324;
  assign n31326 = ~i_hbusreq4 & ~n31325;
  assign n31327 = ~n31322 & ~n31326;
  assign n31328 = ~controllable_hgrant4 & ~n31327;
  assign n31329 = ~n14136 & ~n31328;
  assign n31330 = ~i_hbusreq5 & ~n31329;
  assign n31331 = ~n31321 & ~n31330;
  assign n31332 = ~controllable_hgrant5 & ~n31331;
  assign n31333 = ~n14134 & ~n31332;
  assign n31334 = ~controllable_hmaster2 & ~n31333;
  assign n31335 = ~n31320 & ~n31334;
  assign n31336 = ~controllable_hmaster1 & ~n31335;
  assign n31337 = ~n31311 & ~n31336;
  assign n31338 = ~i_hbusreq6 & ~n31337;
  assign n31339 = ~n31281 & ~n31338;
  assign n31340 = ~controllable_hgrant6 & ~n31339;
  assign n31341 = ~n14094 & ~n31340;
  assign n31342 = controllable_hmaster0 & ~n31341;
  assign n31343 = i_hbusreq6 & ~n31071;
  assign n31344 = controllable_hmaster2 & ~n31239;
  assign n31345 = i_hbusreq5 & ~n31043;
  assign n31346 = i_hbusreq4 & ~n20792;
  assign n31347 = i_hbusreq9 & ~n20792;
  assign n31348 = ~i_hbusreq9 & ~n21302;
  assign n31349 = ~n31347 & ~n31348;
  assign n31350 = ~i_hbusreq4 & ~n31349;
  assign n31351 = ~n31346 & ~n31350;
  assign n31352 = ~controllable_hgrant4 & ~n31351;
  assign n31353 = ~n14177 & ~n31352;
  assign n31354 = ~i_hbusreq5 & ~n31353;
  assign n31355 = ~n31345 & ~n31354;
  assign n31356 = ~controllable_hgrant5 & ~n31355;
  assign n31357 = ~n14175 & ~n31356;
  assign n31358 = ~controllable_hmaster2 & ~n31357;
  assign n31359 = ~n31344 & ~n31358;
  assign n31360 = controllable_hmaster1 & ~n31359;
  assign n31361 = i_hbusreq5 & ~n31053;
  assign n31362 = i_hbusreq4 & ~n31051;
  assign n31363 = i_hlock4 & ~n31231;
  assign n31364 = ~i_hlock4 & ~n31256;
  assign n31365 = ~n31363 & ~n31364;
  assign n31366 = ~i_hbusreq4 & ~n31365;
  assign n31367 = ~n31362 & ~n31366;
  assign n31368 = ~controllable_hgrant4 & ~n31367;
  assign n31369 = ~n14208 & ~n31368;
  assign n31370 = ~i_hbusreq5 & ~n31369;
  assign n31371 = ~n31361 & ~n31370;
  assign n31372 = ~controllable_hgrant5 & ~n31371;
  assign n31373 = ~n14206 & ~n31372;
  assign n31374 = controllable_hmaster2 & ~n31373;
  assign n31375 = i_hbusreq5 & ~n31058;
  assign n31376 = i_hbusreq4 & ~n20820;
  assign n31377 = i_hbusreq9 & ~n20820;
  assign n31378 = ~i_hbusreq9 & ~n21371;
  assign n31379 = ~n31377 & ~n31378;
  assign n31380 = ~i_hbusreq4 & ~n31379;
  assign n31381 = ~n31376 & ~n31380;
  assign n31382 = ~controllable_hgrant4 & ~n31381;
  assign n31383 = ~n14224 & ~n31382;
  assign n31384 = ~i_hbusreq5 & ~n31383;
  assign n31385 = ~n31375 & ~n31384;
  assign n31386 = ~controllable_hgrant5 & ~n31385;
  assign n31387 = ~n14222 & ~n31386;
  assign n31388 = ~controllable_hmaster2 & ~n31387;
  assign n31389 = ~n31374 & ~n31388;
  assign n31390 = ~controllable_hmaster1 & ~n31389;
  assign n31391 = ~n31360 & ~n31390;
  assign n31392 = i_hlock6 & ~n31391;
  assign n31393 = controllable_hmaster2 & ~n31264;
  assign n31394 = ~n31358 & ~n31393;
  assign n31395 = controllable_hmaster1 & ~n31394;
  assign n31396 = ~n31390 & ~n31395;
  assign n31397 = ~i_hlock6 & ~n31396;
  assign n31398 = ~n31392 & ~n31397;
  assign n31399 = ~i_hbusreq6 & ~n31398;
  assign n31400 = ~n31343 & ~n31399;
  assign n31401 = ~controllable_hgrant6 & ~n31400;
  assign n31402 = ~n14173 & ~n31401;
  assign n31403 = ~controllable_hmaster0 & ~n31402;
  assign n31404 = ~n31342 & ~n31403;
  assign n31405 = ~i_hbusreq8 & ~n31404;
  assign n31406 = ~n31280 & ~n31405;
  assign n31407 = ~controllable_hmaster3 & ~n31406;
  assign n31408 = ~n31279 & ~n31407;
  assign n31409 = i_hlock7 & ~n31408;
  assign n31410 = i_hbusreq8 & ~n31117;
  assign n31411 = i_hbusreq6 & ~n31087;
  assign n31412 = i_hbusreq5 & ~n31080;
  assign n31413 = i_hbusreq4 & ~n20635;
  assign n31414 = i_hbusreq9 & ~n20635;
  assign n31415 = ~i_hbusreq9 & ~n20917;
  assign n31416 = ~n31414 & ~n31415;
  assign n31417 = ~i_hbusreq4 & ~n31416;
  assign n31418 = ~n31413 & ~n31417;
  assign n31419 = ~controllable_hgrant4 & ~n31418;
  assign n31420 = ~n13966 & ~n31419;
  assign n31421 = ~i_hbusreq5 & ~n31420;
  assign n31422 = ~n31412 & ~n31421;
  assign n31423 = ~controllable_hgrant5 & ~n31422;
  assign n31424 = ~n13965 & ~n31423;
  assign n31425 = controllable_hmaster1 & ~n31424;
  assign n31426 = controllable_hmaster2 & ~n31424;
  assign n31427 = i_hlock9 & ~n21048;
  assign n31428 = ~n21092 & ~n31427;
  assign n31429 = ~i_hbusreq9 & ~n31428;
  assign n31430 = ~n30674 & ~n31429;
  assign n31431 = ~i_hbusreq4 & ~n31430;
  assign n31432 = ~n30673 & ~n31431;
  assign n31433 = ~controllable_hgrant4 & ~n31432;
  assign n31434 = ~n12676 & ~n31433;
  assign n31435 = ~i_hbusreq5 & ~n31434;
  assign n31436 = ~n30672 & ~n31435;
  assign n31437 = ~controllable_hgrant5 & ~n31436;
  assign n31438 = ~n12674 & ~n31437;
  assign n31439 = ~controllable_hmaster2 & ~n31438;
  assign n31440 = ~n31426 & ~n31439;
  assign n31441 = ~controllable_hmaster1 & ~n31440;
  assign n31442 = ~n31425 & ~n31441;
  assign n31443 = ~i_hbusreq6 & ~n31442;
  assign n31444 = ~n31411 & ~n31443;
  assign n31445 = ~controllable_hgrant6 & ~n31444;
  assign n31446 = ~n13818 & ~n31445;
  assign n31447 = controllable_hmaster0 & ~n31446;
  assign n31448 = i_hbusreq6 & ~n31098;
  assign n31449 = i_hbusreq5 & ~n31092;
  assign n31450 = i_hbusreq4 & ~n20711;
  assign n31451 = i_hbusreq9 & ~n20711;
  assign n31452 = ~i_hbusreq9 & ~n21146;
  assign n31453 = ~n31451 & ~n31452;
  assign n31454 = ~i_hbusreq4 & ~n31453;
  assign n31455 = ~n31450 & ~n31454;
  assign n31456 = ~controllable_hgrant4 & ~n31455;
  assign n31457 = ~n14021 & ~n31456;
  assign n31458 = ~i_hbusreq5 & ~n31457;
  assign n31459 = ~n31449 & ~n31458;
  assign n31460 = ~controllable_hgrant5 & ~n31459;
  assign n31461 = ~n14020 & ~n31460;
  assign n31462 = ~controllable_hmaster2 & ~n31461;
  assign n31463 = ~n31426 & ~n31462;
  assign n31464 = ~controllable_hmaster1 & ~n31463;
  assign n31465 = ~n31425 & ~n31464;
  assign n31466 = ~i_hbusreq6 & ~n31465;
  assign n31467 = ~n31448 & ~n31466;
  assign n31468 = ~controllable_hgrant6 & ~n31467;
  assign n31469 = ~n14019 & ~n31468;
  assign n31470 = ~controllable_hmaster0 & ~n31469;
  assign n31471 = ~n31447 & ~n31470;
  assign n31472 = i_hlock8 & ~n31471;
  assign n31473 = i_hbusreq6 & ~n31111;
  assign n31474 = i_hbusreq5 & ~n31105;
  assign n31475 = i_hbusreq4 & ~n20750;
  assign n31476 = i_hbusreq9 & ~n20750;
  assign n31477 = ~i_hbusreq9 & ~n21221;
  assign n31478 = ~n31476 & ~n31477;
  assign n31479 = ~i_hbusreq4 & ~n31478;
  assign n31480 = ~n31475 & ~n31479;
  assign n31481 = ~controllable_hgrant4 & ~n31480;
  assign n31482 = ~n14056 & ~n31481;
  assign n31483 = ~i_hbusreq5 & ~n31482;
  assign n31484 = ~n31474 & ~n31483;
  assign n31485 = ~controllable_hgrant5 & ~n31484;
  assign n31486 = ~n14055 & ~n31485;
  assign n31487 = ~controllable_hmaster2 & ~n31486;
  assign n31488 = ~n31426 & ~n31487;
  assign n31489 = ~controllable_hmaster1 & ~n31488;
  assign n31490 = ~n31425 & ~n31489;
  assign n31491 = ~i_hbusreq6 & ~n31490;
  assign n31492 = ~n31473 & ~n31491;
  assign n31493 = ~controllable_hgrant6 & ~n31492;
  assign n31494 = ~n14054 & ~n31493;
  assign n31495 = ~controllable_hmaster0 & ~n31494;
  assign n31496 = ~n31447 & ~n31495;
  assign n31497 = ~i_hlock8 & ~n31496;
  assign n31498 = ~n31472 & ~n31497;
  assign n31499 = ~i_hbusreq8 & ~n31498;
  assign n31500 = ~n31410 & ~n31499;
  assign n31501 = controllable_hmaster3 & ~n31500;
  assign n31502 = i_hbusreq8 & ~n31182;
  assign n31503 = i_hbusreq6 & ~n31144;
  assign n31504 = i_hbusreq5 & ~n31120;
  assign n31505 = i_hbusreq4 & ~n20669;
  assign n31506 = i_hbusreq9 & ~n20669;
  assign n31507 = ~i_hbusreq9 & ~n20985;
  assign n31508 = ~n31506 & ~n31507;
  assign n31509 = ~i_hbusreq4 & ~n31508;
  assign n31510 = ~n31505 & ~n31509;
  assign n31511 = ~controllable_hgrant4 & ~n31510;
  assign n31512 = ~n14056 & ~n31511;
  assign n31513 = ~i_hbusreq5 & ~n31512;
  assign n31514 = ~n31504 & ~n31513;
  assign n31515 = ~controllable_hgrant5 & ~n31514;
  assign n31516 = ~n14055 & ~n31515;
  assign n31517 = controllable_hmaster2 & ~n31516;
  assign n31518 = i_hbusreq5 & ~n31125;
  assign n31519 = i_hbusreq4 & ~n20735;
  assign n31520 = i_hbusreq9 & ~n20735;
  assign n31521 = ~i_hbusreq9 & ~n21191;
  assign n31522 = ~n31520 & ~n31521;
  assign n31523 = ~i_hbusreq4 & ~n31522;
  assign n31524 = ~n31519 & ~n31523;
  assign n31525 = ~controllable_hgrant4 & ~n31524;
  assign n31526 = ~n14099 & ~n31525;
  assign n31527 = ~i_hbusreq5 & ~n31526;
  assign n31528 = ~n31518 & ~n31527;
  assign n31529 = ~controllable_hgrant5 & ~n31528;
  assign n31530 = ~n14097 & ~n31529;
  assign n31531 = ~controllable_hmaster2 & ~n31530;
  assign n31532 = ~n31517 & ~n31531;
  assign n31533 = controllable_hmaster1 & ~n31532;
  assign n31534 = i_hbusreq5 & ~n31133;
  assign n31535 = i_hlock5 & ~n31457;
  assign n31536 = ~i_hlock5 & ~n31482;
  assign n31537 = ~n31535 & ~n31536;
  assign n31538 = ~i_hbusreq5 & ~n31537;
  assign n31539 = ~n31534 & ~n31538;
  assign n31540 = ~controllable_hgrant5 & ~n31539;
  assign n31541 = ~n14124 & ~n31540;
  assign n31542 = controllable_hmaster2 & ~n31541;
  assign n31543 = i_hbusreq5 & ~n31138;
  assign n31544 = i_hbusreq4 & ~n20774;
  assign n31545 = i_hbusreq9 & ~n20774;
  assign n31546 = ~i_hbusreq9 & ~n21266;
  assign n31547 = ~n31545 & ~n31546;
  assign n31548 = ~i_hbusreq4 & ~n31547;
  assign n31549 = ~n31544 & ~n31548;
  assign n31550 = ~controllable_hgrant4 & ~n31549;
  assign n31551 = ~n14136 & ~n31550;
  assign n31552 = ~i_hbusreq5 & ~n31551;
  assign n31553 = ~n31543 & ~n31552;
  assign n31554 = ~controllable_hgrant5 & ~n31553;
  assign n31555 = ~n14134 & ~n31554;
  assign n31556 = ~controllable_hmaster2 & ~n31555;
  assign n31557 = ~n31542 & ~n31556;
  assign n31558 = ~controllable_hmaster1 & ~n31557;
  assign n31559 = ~n31533 & ~n31558;
  assign n31560 = ~i_hbusreq6 & ~n31559;
  assign n31561 = ~n31503 & ~n31560;
  assign n31562 = ~controllable_hgrant6 & ~n31561;
  assign n31563 = ~n14298 & ~n31562;
  assign n31564 = controllable_hmaster0 & ~n31563;
  assign n31565 = i_hbusreq6 & ~n31178;
  assign n31566 = controllable_hmaster2 & ~n31461;
  assign n31567 = i_hbusreq5 & ~n31150;
  assign n31568 = i_hbusreq4 & ~n20798;
  assign n31569 = i_hbusreq9 & ~n20798;
  assign n31570 = ~i_hbusreq9 & ~n21314;
  assign n31571 = ~n31569 & ~n31570;
  assign n31572 = ~i_hbusreq4 & ~n31571;
  assign n31573 = ~n31568 & ~n31572;
  assign n31574 = ~controllable_hgrant4 & ~n31573;
  assign n31575 = ~n14177 & ~n31574;
  assign n31576 = ~i_hbusreq5 & ~n31575;
  assign n31577 = ~n31567 & ~n31576;
  assign n31578 = ~controllable_hgrant5 & ~n31577;
  assign n31579 = ~n14175 & ~n31578;
  assign n31580 = ~controllable_hmaster2 & ~n31579;
  assign n31581 = ~n31566 & ~n31580;
  assign n31582 = controllable_hmaster1 & ~n31581;
  assign n31583 = i_hbusreq5 & ~n31160;
  assign n31584 = i_hbusreq4 & ~n31158;
  assign n31585 = i_hlock4 & ~n31453;
  assign n31586 = ~i_hlock4 & ~n31478;
  assign n31587 = ~n31585 & ~n31586;
  assign n31588 = ~i_hbusreq4 & ~n31587;
  assign n31589 = ~n31584 & ~n31588;
  assign n31590 = ~controllable_hgrant4 & ~n31589;
  assign n31591 = ~n14208 & ~n31590;
  assign n31592 = ~i_hbusreq5 & ~n31591;
  assign n31593 = ~n31583 & ~n31592;
  assign n31594 = ~controllable_hgrant5 & ~n31593;
  assign n31595 = ~n14206 & ~n31594;
  assign n31596 = controllable_hmaster2 & ~n31595;
  assign n31597 = i_hbusreq5 & ~n31165;
  assign n31598 = i_hbusreq4 & ~n20826;
  assign n31599 = i_hbusreq9 & ~n20826;
  assign n31600 = ~i_hbusreq9 & ~n21391;
  assign n31601 = ~n31599 & ~n31600;
  assign n31602 = ~i_hbusreq4 & ~n31601;
  assign n31603 = ~n31598 & ~n31602;
  assign n31604 = ~controllable_hgrant4 & ~n31603;
  assign n31605 = ~n14224 & ~n31604;
  assign n31606 = ~i_hbusreq5 & ~n31605;
  assign n31607 = ~n31597 & ~n31606;
  assign n31608 = ~controllable_hgrant5 & ~n31607;
  assign n31609 = ~n14222 & ~n31608;
  assign n31610 = ~controllable_hmaster2 & ~n31609;
  assign n31611 = ~n31596 & ~n31610;
  assign n31612 = ~controllable_hmaster1 & ~n31611;
  assign n31613 = ~n31582 & ~n31612;
  assign n31614 = i_hlock6 & ~n31613;
  assign n31615 = controllable_hmaster2 & ~n31486;
  assign n31616 = ~n31580 & ~n31615;
  assign n31617 = controllable_hmaster1 & ~n31616;
  assign n31618 = ~n31612 & ~n31617;
  assign n31619 = ~i_hlock6 & ~n31618;
  assign n31620 = ~n31614 & ~n31619;
  assign n31621 = ~i_hbusreq6 & ~n31620;
  assign n31622 = ~n31565 & ~n31621;
  assign n31623 = ~controllable_hgrant6 & ~n31622;
  assign n31624 = ~n14173 & ~n31623;
  assign n31625 = ~controllable_hmaster0 & ~n31624;
  assign n31626 = ~n31564 & ~n31625;
  assign n31627 = ~i_hbusreq8 & ~n31626;
  assign n31628 = ~n31502 & ~n31627;
  assign n31629 = ~controllable_hmaster3 & ~n31628;
  assign n31630 = ~n31501 & ~n31629;
  assign n31631 = ~i_hlock7 & ~n31630;
  assign n31632 = ~n31409 & ~n31631;
  assign n31633 = ~i_hbusreq7 & ~n31632;
  assign n31634 = ~n31187 & ~n31633;
  assign n31635 = n7924 & ~n31634;
  assign n31636 = ~n29844 & ~n31635;
  assign n31637 = ~n8214 & ~n31636;
  assign n31638 = ~i_hlock9 & ~n20747;
  assign n31639 = ~n20706 & ~n31638;
  assign n31640 = ~controllable_hgrant4 & ~n31639;
  assign n31641 = ~n12609 & ~n31640;
  assign n31642 = ~controllable_hgrant5 & ~n31641;
  assign n31643 = ~n12608 & ~n31642;
  assign n31644 = ~controllable_hmaster2 & ~n31643;
  assign n31645 = ~n30977 & ~n31644;
  assign n31646 = ~controllable_hmaster1 & ~n31645;
  assign n31647 = ~n30976 & ~n31646;
  assign n31648 = ~controllable_hgrant6 & ~n31647;
  assign n31649 = ~n13122 & ~n31648;
  assign n31650 = controllable_hmaster0 & ~n31649;
  assign n31651 = ~n30259 & ~n30977;
  assign n31652 = ~controllable_hmaster1 & ~n31651;
  assign n31653 = ~n30976 & ~n31652;
  assign n31654 = ~controllable_hgrant6 & ~n31653;
  assign n31655 = ~n13406 & ~n31654;
  assign n31656 = ~controllable_hmaster0 & ~n31655;
  assign n31657 = ~n31650 & ~n31656;
  assign n31658 = i_hlock8 & ~n31657;
  assign n31659 = ~n30272 & ~n30977;
  assign n31660 = ~controllable_hmaster1 & ~n31659;
  assign n31661 = ~n30976 & ~n31660;
  assign n31662 = ~controllable_hgrant6 & ~n31661;
  assign n31663 = ~n13427 & ~n31662;
  assign n31664 = ~controllable_hmaster0 & ~n31663;
  assign n31665 = ~n31650 & ~n31664;
  assign n31666 = ~i_hlock8 & ~n31665;
  assign n31667 = ~n31658 & ~n31666;
  assign n31668 = controllable_hmaster3 & ~n31667;
  assign n31669 = ~n31076 & ~n31668;
  assign n31670 = i_hlock7 & ~n31669;
  assign n31671 = i_hlock9 & ~n20711;
  assign n31672 = ~n20751 & ~n31671;
  assign n31673 = ~controllable_hgrant4 & ~n31672;
  assign n31674 = ~n12609 & ~n31673;
  assign n31675 = ~controllable_hgrant5 & ~n31674;
  assign n31676 = ~n12608 & ~n31675;
  assign n31677 = ~controllable_hmaster2 & ~n31676;
  assign n31678 = ~n31084 & ~n31677;
  assign n31679 = ~controllable_hmaster1 & ~n31678;
  assign n31680 = ~n31083 & ~n31679;
  assign n31681 = ~controllable_hgrant6 & ~n31680;
  assign n31682 = ~n13122 & ~n31681;
  assign n31683 = controllable_hmaster0 & ~n31682;
  assign n31684 = ~n30362 & ~n31084;
  assign n31685 = ~controllable_hmaster1 & ~n31684;
  assign n31686 = ~n31083 & ~n31685;
  assign n31687 = ~controllable_hgrant6 & ~n31686;
  assign n31688 = ~n13406 & ~n31687;
  assign n31689 = ~controllable_hmaster0 & ~n31688;
  assign n31690 = ~n31683 & ~n31689;
  assign n31691 = i_hlock8 & ~n31690;
  assign n31692 = ~n30375 & ~n31084;
  assign n31693 = ~controllable_hmaster1 & ~n31692;
  assign n31694 = ~n31083 & ~n31693;
  assign n31695 = ~controllable_hgrant6 & ~n31694;
  assign n31696 = ~n13427 & ~n31695;
  assign n31697 = ~controllable_hmaster0 & ~n31696;
  assign n31698 = ~n31683 & ~n31697;
  assign n31699 = ~i_hlock8 & ~n31698;
  assign n31700 = ~n31691 & ~n31699;
  assign n31701 = controllable_hmaster3 & ~n31700;
  assign n31702 = ~n31183 & ~n31701;
  assign n31703 = ~i_hlock7 & ~n31702;
  assign n31704 = ~n31670 & ~n31703;
  assign n31705 = i_hbusreq7 & ~n31704;
  assign n31706 = i_hbusreq8 & ~n31667;
  assign n31707 = i_hbusreq6 & ~n31647;
  assign n31708 = i_hbusreq5 & ~n31641;
  assign n31709 = i_hbusreq4 & ~n31639;
  assign n31710 = i_hbusreq9 & ~n31639;
  assign n31711 = ~i_hlock9 & ~n21215;
  assign n31712 = ~n21135 & ~n31711;
  assign n31713 = ~i_hbusreq9 & ~n31712;
  assign n31714 = ~n31710 & ~n31713;
  assign n31715 = ~i_hbusreq4 & ~n31714;
  assign n31716 = ~n31709 & ~n31715;
  assign n31717 = ~controllable_hgrant4 & ~n31716;
  assign n31718 = ~n14322 & ~n31717;
  assign n31719 = ~i_hbusreq5 & ~n31718;
  assign n31720 = ~n31708 & ~n31719;
  assign n31721 = ~controllable_hgrant5 & ~n31720;
  assign n31722 = ~n14321 & ~n31721;
  assign n31723 = ~controllable_hmaster2 & ~n31722;
  assign n31724 = ~n31204 & ~n31723;
  assign n31725 = ~controllable_hmaster1 & ~n31724;
  assign n31726 = ~n31203 & ~n31725;
  assign n31727 = ~i_hbusreq6 & ~n31726;
  assign n31728 = ~n31707 & ~n31727;
  assign n31729 = ~controllable_hgrant6 & ~n31728;
  assign n31730 = ~n14320 & ~n31729;
  assign n31731 = controllable_hmaster0 & ~n31730;
  assign n31732 = i_hbusreq6 & ~n31653;
  assign n31733 = ~i_hbusreq9 & ~n21030;
  assign n31734 = ~n30491 & ~n31733;
  assign n31735 = ~i_hbusreq4 & ~n31734;
  assign n31736 = ~n30490 & ~n31735;
  assign n31737 = ~controllable_hgrant4 & ~n31736;
  assign n31738 = ~n13524 & ~n31737;
  assign n31739 = ~i_hbusreq5 & ~n31738;
  assign n31740 = ~n30489 & ~n31739;
  assign n31741 = ~controllable_hgrant5 & ~n31740;
  assign n31742 = ~n13522 & ~n31741;
  assign n31743 = ~controllable_hmaster2 & ~n31742;
  assign n31744 = ~n31204 & ~n31743;
  assign n31745 = ~controllable_hmaster1 & ~n31744;
  assign n31746 = ~n31203 & ~n31745;
  assign n31747 = ~i_hbusreq6 & ~n31746;
  assign n31748 = ~n31732 & ~n31747;
  assign n31749 = ~controllable_hgrant6 & ~n31748;
  assign n31750 = ~n14443 & ~n31749;
  assign n31751 = ~controllable_hmaster0 & ~n31750;
  assign n31752 = ~n31731 & ~n31751;
  assign n31753 = i_hlock8 & ~n31752;
  assign n31754 = i_hbusreq6 & ~n31661;
  assign n31755 = ~i_hbusreq9 & ~n21081;
  assign n31756 = ~n30516 & ~n31755;
  assign n31757 = ~i_hbusreq4 & ~n31756;
  assign n31758 = ~n30515 & ~n31757;
  assign n31759 = ~controllable_hgrant4 & ~n31758;
  assign n31760 = ~n13577 & ~n31759;
  assign n31761 = ~i_hbusreq5 & ~n31760;
  assign n31762 = ~n30514 & ~n31761;
  assign n31763 = ~controllable_hgrant5 & ~n31762;
  assign n31764 = ~n13575 & ~n31763;
  assign n31765 = ~controllable_hmaster2 & ~n31764;
  assign n31766 = ~n31204 & ~n31765;
  assign n31767 = ~controllable_hmaster1 & ~n31766;
  assign n31768 = ~n31203 & ~n31767;
  assign n31769 = ~i_hbusreq6 & ~n31768;
  assign n31770 = ~n31754 & ~n31769;
  assign n31771 = ~controllable_hgrant6 & ~n31770;
  assign n31772 = ~n14484 & ~n31771;
  assign n31773 = ~controllable_hmaster0 & ~n31772;
  assign n31774 = ~n31731 & ~n31773;
  assign n31775 = ~i_hlock8 & ~n31774;
  assign n31776 = ~n31753 & ~n31775;
  assign n31777 = ~i_hbusreq8 & ~n31776;
  assign n31778 = ~n31706 & ~n31777;
  assign n31779 = controllable_hmaster3 & ~n31778;
  assign n31780 = ~n31407 & ~n31779;
  assign n31781 = i_hlock7 & ~n31780;
  assign n31782 = i_hbusreq8 & ~n31700;
  assign n31783 = i_hbusreq6 & ~n31680;
  assign n31784 = i_hbusreq5 & ~n31674;
  assign n31785 = i_hbusreq4 & ~n31672;
  assign n31786 = i_hbusreq9 & ~n31672;
  assign n31787 = i_hlock9 & ~n21146;
  assign n31788 = ~n21222 & ~n31787;
  assign n31789 = ~i_hbusreq9 & ~n31788;
  assign n31790 = ~n31786 & ~n31789;
  assign n31791 = ~i_hbusreq4 & ~n31790;
  assign n31792 = ~n31785 & ~n31791;
  assign n31793 = ~controllable_hgrant4 & ~n31792;
  assign n31794 = ~n14322 & ~n31793;
  assign n31795 = ~i_hbusreq5 & ~n31794;
  assign n31796 = ~n31784 & ~n31795;
  assign n31797 = ~controllable_hgrant5 & ~n31796;
  assign n31798 = ~n14321 & ~n31797;
  assign n31799 = ~controllable_hmaster2 & ~n31798;
  assign n31800 = ~n31426 & ~n31799;
  assign n31801 = ~controllable_hmaster1 & ~n31800;
  assign n31802 = ~n31425 & ~n31801;
  assign n31803 = ~i_hbusreq6 & ~n31802;
  assign n31804 = ~n31783 & ~n31803;
  assign n31805 = ~controllable_hgrant6 & ~n31804;
  assign n31806 = ~n14320 & ~n31805;
  assign n31807 = controllable_hmaster0 & ~n31806;
  assign n31808 = i_hbusreq6 & ~n31686;
  assign n31809 = ~i_hbusreq9 & ~n21048;
  assign n31810 = ~n30699 & ~n31809;
  assign n31811 = ~i_hbusreq4 & ~n31810;
  assign n31812 = ~n30698 & ~n31811;
  assign n31813 = ~controllable_hgrant4 & ~n31812;
  assign n31814 = ~n13524 & ~n31813;
  assign n31815 = ~i_hbusreq5 & ~n31814;
  assign n31816 = ~n30697 & ~n31815;
  assign n31817 = ~controllable_hgrant5 & ~n31816;
  assign n31818 = ~n13522 & ~n31817;
  assign n31819 = ~controllable_hmaster2 & ~n31818;
  assign n31820 = ~n31426 & ~n31819;
  assign n31821 = ~controllable_hmaster1 & ~n31820;
  assign n31822 = ~n31425 & ~n31821;
  assign n31823 = ~i_hbusreq6 & ~n31822;
  assign n31824 = ~n31808 & ~n31823;
  assign n31825 = ~controllable_hgrant6 & ~n31824;
  assign n31826 = ~n14443 & ~n31825;
  assign n31827 = ~controllable_hmaster0 & ~n31826;
  assign n31828 = ~n31807 & ~n31827;
  assign n31829 = i_hlock8 & ~n31828;
  assign n31830 = i_hbusreq6 & ~n31694;
  assign n31831 = ~i_hbusreq9 & ~n21091;
  assign n31832 = ~n30724 & ~n31831;
  assign n31833 = ~i_hbusreq4 & ~n31832;
  assign n31834 = ~n30723 & ~n31833;
  assign n31835 = ~controllable_hgrant4 & ~n31834;
  assign n31836 = ~n13577 & ~n31835;
  assign n31837 = ~i_hbusreq5 & ~n31836;
  assign n31838 = ~n30722 & ~n31837;
  assign n31839 = ~controllable_hgrant5 & ~n31838;
  assign n31840 = ~n13575 & ~n31839;
  assign n31841 = ~controllable_hmaster2 & ~n31840;
  assign n31842 = ~n31426 & ~n31841;
  assign n31843 = ~controllable_hmaster1 & ~n31842;
  assign n31844 = ~n31425 & ~n31843;
  assign n31845 = ~i_hbusreq6 & ~n31844;
  assign n31846 = ~n31830 & ~n31845;
  assign n31847 = ~controllable_hgrant6 & ~n31846;
  assign n31848 = ~n14484 & ~n31847;
  assign n31849 = ~controllable_hmaster0 & ~n31848;
  assign n31850 = ~n31807 & ~n31849;
  assign n31851 = ~i_hlock8 & ~n31850;
  assign n31852 = ~n31829 & ~n31851;
  assign n31853 = ~i_hbusreq8 & ~n31852;
  assign n31854 = ~n31782 & ~n31853;
  assign n31855 = controllable_hmaster3 & ~n31854;
  assign n31856 = ~n31629 & ~n31855;
  assign n31857 = ~i_hlock7 & ~n31856;
  assign n31858 = ~n31781 & ~n31857;
  assign n31859 = ~i_hbusreq7 & ~n31858;
  assign n31860 = ~n31705 & ~n31859;
  assign n31861 = n7924 & ~n31860;
  assign n31862 = ~n30066 & ~n31861;
  assign n31863 = n8214 & ~n31862;
  assign n31864 = ~n31637 & ~n31863;
  assign n31865 = ~n8202 & ~n31864;
  assign n31866 = ~n30994 & ~n31650;
  assign n31867 = i_hlock8 & ~n31866;
  assign n31868 = ~n31007 & ~n31650;
  assign n31869 = ~i_hlock8 & ~n31868;
  assign n31870 = ~n31867 & ~n31869;
  assign n31871 = controllable_hmaster3 & ~n31870;
  assign n31872 = ~n30307 & ~n31046;
  assign n31873 = controllable_hmaster1 & ~n31872;
  assign n31874 = ~n31063 & ~n31873;
  assign n31875 = i_hlock6 & ~n31874;
  assign n31876 = ~n30332 & ~n31046;
  assign n31877 = controllable_hmaster1 & ~n31876;
  assign n31878 = ~n31063 & ~n31877;
  assign n31879 = ~i_hlock6 & ~n31878;
  assign n31880 = ~n31875 & ~n31879;
  assign n31881 = ~controllable_hgrant6 & ~n31880;
  assign n31882 = ~n13894 & ~n31881;
  assign n31883 = ~controllable_hmaster0 & ~n31882;
  assign n31884 = ~n31040 & ~n31883;
  assign n31885 = ~controllable_hmaster3 & ~n31884;
  assign n31886 = ~n31871 & ~n31885;
  assign n31887 = i_hlock7 & ~n31886;
  assign n31888 = ~n31101 & ~n31683;
  assign n31889 = i_hlock8 & ~n31888;
  assign n31890 = ~n31114 & ~n31683;
  assign n31891 = ~i_hlock8 & ~n31890;
  assign n31892 = ~n31889 & ~n31891;
  assign n31893 = controllable_hmaster3 & ~n31892;
  assign n31894 = ~n30410 & ~n31153;
  assign n31895 = controllable_hmaster1 & ~n31894;
  assign n31896 = ~n31170 & ~n31895;
  assign n31897 = i_hlock6 & ~n31896;
  assign n31898 = ~n30435 & ~n31153;
  assign n31899 = controllable_hmaster1 & ~n31898;
  assign n31900 = ~n31170 & ~n31899;
  assign n31901 = ~i_hlock6 & ~n31900;
  assign n31902 = ~n31897 & ~n31901;
  assign n31903 = ~controllable_hgrant6 & ~n31902;
  assign n31904 = ~n13894 & ~n31903;
  assign n31905 = ~controllable_hmaster0 & ~n31904;
  assign n31906 = ~n31147 & ~n31905;
  assign n31907 = ~controllable_hmaster3 & ~n31906;
  assign n31908 = ~n31893 & ~n31907;
  assign n31909 = ~i_hlock7 & ~n31908;
  assign n31910 = ~n31887 & ~n31909;
  assign n31911 = i_hbusreq7 & ~n31910;
  assign n31912 = i_hbusreq8 & ~n31870;
  assign n31913 = ~n31248 & ~n31731;
  assign n31914 = i_hlock8 & ~n31913;
  assign n31915 = ~n31273 & ~n31731;
  assign n31916 = ~i_hlock8 & ~n31915;
  assign n31917 = ~n31914 & ~n31916;
  assign n31918 = ~i_hbusreq8 & ~n31917;
  assign n31919 = ~n31912 & ~n31918;
  assign n31920 = controllable_hmaster3 & ~n31919;
  assign n31921 = i_hbusreq8 & ~n31884;
  assign n31922 = i_hbusreq6 & ~n31880;
  assign n31923 = controllable_hmaster2 & ~n31742;
  assign n31924 = ~n31358 & ~n31923;
  assign n31925 = controllable_hmaster1 & ~n31924;
  assign n31926 = ~n31390 & ~n31925;
  assign n31927 = i_hlock6 & ~n31926;
  assign n31928 = controllable_hmaster2 & ~n31764;
  assign n31929 = ~n31358 & ~n31928;
  assign n31930 = controllable_hmaster1 & ~n31929;
  assign n31931 = ~n31390 & ~n31930;
  assign n31932 = ~i_hlock6 & ~n31931;
  assign n31933 = ~n31927 & ~n31932;
  assign n31934 = ~i_hbusreq6 & ~n31933;
  assign n31935 = ~n31922 & ~n31934;
  assign n31936 = ~controllable_hgrant6 & ~n31935;
  assign n31937 = ~n14802 & ~n31936;
  assign n31938 = ~controllable_hmaster0 & ~n31937;
  assign n31939 = ~n31342 & ~n31938;
  assign n31940 = ~i_hbusreq8 & ~n31939;
  assign n31941 = ~n31921 & ~n31940;
  assign n31942 = ~controllable_hmaster3 & ~n31941;
  assign n31943 = ~n31920 & ~n31942;
  assign n31944 = i_hlock7 & ~n31943;
  assign n31945 = i_hbusreq8 & ~n31892;
  assign n31946 = ~n31470 & ~n31807;
  assign n31947 = i_hlock8 & ~n31946;
  assign n31948 = ~n31495 & ~n31807;
  assign n31949 = ~i_hlock8 & ~n31948;
  assign n31950 = ~n31947 & ~n31949;
  assign n31951 = ~i_hbusreq8 & ~n31950;
  assign n31952 = ~n31945 & ~n31951;
  assign n31953 = controllable_hmaster3 & ~n31952;
  assign n31954 = i_hbusreq8 & ~n31906;
  assign n31955 = i_hbusreq6 & ~n31902;
  assign n31956 = controllable_hmaster2 & ~n31818;
  assign n31957 = ~n31580 & ~n31956;
  assign n31958 = controllable_hmaster1 & ~n31957;
  assign n31959 = ~n31612 & ~n31958;
  assign n31960 = i_hlock6 & ~n31959;
  assign n31961 = controllable_hmaster2 & ~n31840;
  assign n31962 = ~n31580 & ~n31961;
  assign n31963 = controllable_hmaster1 & ~n31962;
  assign n31964 = ~n31612 & ~n31963;
  assign n31965 = ~i_hlock6 & ~n31964;
  assign n31966 = ~n31960 & ~n31965;
  assign n31967 = ~i_hbusreq6 & ~n31966;
  assign n31968 = ~n31955 & ~n31967;
  assign n31969 = ~controllable_hgrant6 & ~n31968;
  assign n31970 = ~n14802 & ~n31969;
  assign n31971 = ~controllable_hmaster0 & ~n31970;
  assign n31972 = ~n31564 & ~n31971;
  assign n31973 = ~i_hbusreq8 & ~n31972;
  assign n31974 = ~n31954 & ~n31973;
  assign n31975 = ~controllable_hmaster3 & ~n31974;
  assign n31976 = ~n31953 & ~n31975;
  assign n31977 = ~i_hlock7 & ~n31976;
  assign n31978 = ~n31944 & ~n31977;
  assign n31979 = ~i_hbusreq7 & ~n31978;
  assign n31980 = ~n31911 & ~n31979;
  assign n31981 = n7924 & ~n31980;
  assign n31982 = ~n30914 & ~n31981;
  assign n31983 = n8214 & ~n31982;
  assign n31984 = ~n30871 & ~n31983;
  assign n31985 = n8202 & ~n31984;
  assign n31986 = ~n31865 & ~n31985;
  assign n31987 = n7920 & ~n31986;
  assign n31988 = ~n28799 & ~n31987;
  assign n31989 = n7728 & ~n31988;
  assign n31990 = ~n21649 & ~n28847;
  assign n31991 = ~controllable_hmaster1 & ~n31990;
  assign n31992 = ~n21648 & ~n31991;
  assign n31993 = ~i_hbusreq6 & ~n31992;
  assign n31994 = ~n30175 & ~n31993;
  assign n31995 = ~controllable_hgrant6 & ~n31994;
  assign n31996 = ~n14849 & ~n31995;
  assign n31997 = controllable_hmaster0 & ~n31996;
  assign n31998 = ~n21665 & ~n31997;
  assign n31999 = i_hlock8 & ~n31998;
  assign n32000 = ~n21675 & ~n31997;
  assign n32001 = ~i_hlock8 & ~n32000;
  assign n32002 = ~n31999 & ~n32001;
  assign n32003 = ~i_hbusreq8 & ~n32002;
  assign n32004 = ~n30174 & ~n32003;
  assign n32005 = controllable_hmaster3 & ~n32004;
  assign n32006 = ~n21699 & ~n28913;
  assign n32007 = controllable_hmaster1 & ~n32006;
  assign n32008 = ~n21733 & ~n32007;
  assign n32009 = ~i_hbusreq6 & ~n32008;
  assign n32010 = ~n30207 & ~n32009;
  assign n32011 = ~controllable_hgrant6 & ~n32010;
  assign n32012 = ~n14995 & ~n32011;
  assign n32013 = controllable_hmaster0 & ~n32012;
  assign n32014 = ~n21809 & ~n32013;
  assign n32015 = ~i_hbusreq8 & ~n32014;
  assign n32016 = ~n30206 & ~n32015;
  assign n32017 = ~controllable_hmaster3 & ~n32016;
  assign n32018 = ~n32005 & ~n32017;
  assign n32019 = i_hlock7 & ~n32018;
  assign n32020 = ~n21699 & ~n28943;
  assign n32021 = controllable_hmaster1 & ~n32020;
  assign n32022 = ~n21733 & ~n32021;
  assign n32023 = ~i_hbusreq6 & ~n32022;
  assign n32024 = ~n30223 & ~n32023;
  assign n32025 = ~controllable_hgrant6 & ~n32024;
  assign n32026 = ~n15152 & ~n32025;
  assign n32027 = controllable_hmaster0 & ~n32026;
  assign n32028 = ~n21809 & ~n32027;
  assign n32029 = ~i_hbusreq8 & ~n32028;
  assign n32030 = ~n30222 & ~n32029;
  assign n32031 = ~controllable_hmaster3 & ~n32030;
  assign n32032 = ~n32005 & ~n32031;
  assign n32033 = ~i_hlock7 & ~n32032;
  assign n32034 = ~n32019 & ~n32033;
  assign n32035 = ~i_hbusreq7 & ~n32034;
  assign n32036 = ~n30173 & ~n32035;
  assign n32037 = ~n7924 & ~n32036;
  assign n32038 = ~i_hbusreq9 & ~n21866;
  assign n32039 = ~n29555 & ~n32038;
  assign n32040 = ~i_hbusreq4 & ~n32039;
  assign n32041 = ~n29554 & ~n32040;
  assign n32042 = ~controllable_hgrant4 & ~n32041;
  assign n32043 = ~n14875 & ~n32042;
  assign n32044 = ~i_hbusreq5 & ~n32043;
  assign n32045 = ~n29553 & ~n32044;
  assign n32046 = ~controllable_hgrant5 & ~n32045;
  assign n32047 = ~n14874 & ~n32046;
  assign n32048 = controllable_hmaster1 & ~n32047;
  assign n32049 = controllable_hmaster2 & ~n32047;
  assign n32050 = ~i_hlock9 & ~n21961;
  assign n32051 = ~n21918 & ~n32050;
  assign n32052 = ~i_hbusreq9 & ~n32051;
  assign n32053 = ~n30466 & ~n32052;
  assign n32054 = ~i_hbusreq4 & ~n32053;
  assign n32055 = ~n30465 & ~n32054;
  assign n32056 = ~controllable_hgrant4 & ~n32055;
  assign n32057 = ~n12676 & ~n32056;
  assign n32058 = ~i_hbusreq5 & ~n32057;
  assign n32059 = ~n30464 & ~n32058;
  assign n32060 = ~controllable_hgrant5 & ~n32059;
  assign n32061 = ~n12674 & ~n32060;
  assign n32062 = ~controllable_hmaster2 & ~n32061;
  assign n32063 = ~n32049 & ~n32062;
  assign n32064 = ~controllable_hmaster1 & ~n32063;
  assign n32065 = ~n32048 & ~n32064;
  assign n32066 = ~i_hbusreq6 & ~n32065;
  assign n32067 = ~n30451 & ~n32066;
  assign n32068 = ~controllable_hgrant6 & ~n32067;
  assign n32069 = ~n14849 & ~n32068;
  assign n32070 = controllable_hmaster0 & ~n32069;
  assign n32071 = ~i_hbusreq9 & ~n21917;
  assign n32072 = ~n30491 & ~n32071;
  assign n32073 = ~i_hbusreq4 & ~n32072;
  assign n32074 = ~n30490 & ~n32073;
  assign n32075 = ~controllable_hgrant4 & ~n32074;
  assign n32076 = ~n13524 & ~n32075;
  assign n32077 = ~i_hbusreq5 & ~n32076;
  assign n32078 = ~n30489 & ~n32077;
  assign n32079 = ~controllable_hgrant5 & ~n32078;
  assign n32080 = ~n13522 & ~n32079;
  assign n32081 = ~controllable_hmaster2 & ~n32080;
  assign n32082 = ~n32049 & ~n32081;
  assign n32083 = ~controllable_hmaster1 & ~n32082;
  assign n32084 = ~n32048 & ~n32083;
  assign n32085 = ~i_hbusreq6 & ~n32084;
  assign n32086 = ~n30488 & ~n32085;
  assign n32087 = ~controllable_hgrant6 & ~n32086;
  assign n32088 = ~n14927 & ~n32087;
  assign n32089 = ~controllable_hmaster0 & ~n32088;
  assign n32090 = ~n32070 & ~n32089;
  assign n32091 = i_hlock8 & ~n32090;
  assign n32092 = ~i_hbusreq9 & ~n21961;
  assign n32093 = ~n30516 & ~n32092;
  assign n32094 = ~i_hbusreq4 & ~n32093;
  assign n32095 = ~n30515 & ~n32094;
  assign n32096 = ~controllable_hgrant4 & ~n32095;
  assign n32097 = ~n13577 & ~n32096;
  assign n32098 = ~i_hbusreq5 & ~n32097;
  assign n32099 = ~n30514 & ~n32098;
  assign n32100 = ~controllable_hgrant5 & ~n32099;
  assign n32101 = ~n13575 & ~n32100;
  assign n32102 = ~controllable_hmaster2 & ~n32101;
  assign n32103 = ~n32049 & ~n32102;
  assign n32104 = ~controllable_hmaster1 & ~n32103;
  assign n32105 = ~n32048 & ~n32104;
  assign n32106 = ~i_hbusreq6 & ~n32105;
  assign n32107 = ~n30513 & ~n32106;
  assign n32108 = ~controllable_hgrant6 & ~n32107;
  assign n32109 = ~n14960 & ~n32108;
  assign n32110 = ~controllable_hmaster0 & ~n32109;
  assign n32111 = ~n32070 & ~n32110;
  assign n32112 = ~i_hlock8 & ~n32111;
  assign n32113 = ~n32091 & ~n32112;
  assign n32114 = ~i_hbusreq8 & ~n32113;
  assign n32115 = ~n30450 & ~n32114;
  assign n32116 = controllable_hmaster3 & ~n32115;
  assign n32117 = ~i_hbusreq9 & ~n22006;
  assign n32118 = ~n30546 & ~n32117;
  assign n32119 = ~i_hbusreq4 & ~n32118;
  assign n32120 = ~n30545 & ~n32119;
  assign n32121 = ~controllable_hgrant4 & ~n32120;
  assign n32122 = ~n14998 & ~n32121;
  assign n32123 = ~i_hbusreq5 & ~n32122;
  assign n32124 = ~n30544 & ~n32123;
  assign n32125 = ~controllable_hgrant5 & ~n32124;
  assign n32126 = ~n14997 & ~n32125;
  assign n32127 = ~controllable_hmaster2 & ~n32126;
  assign n32128 = ~n29051 & ~n32127;
  assign n32129 = controllable_hmaster1 & ~n32128;
  assign n32130 = i_hlock5 & ~n32076;
  assign n32131 = ~i_hlock5 & ~n32097;
  assign n32132 = ~n32130 & ~n32131;
  assign n32133 = ~i_hbusreq5 & ~n32132;
  assign n32134 = ~n30560 & ~n32133;
  assign n32135 = ~controllable_hgrant5 & ~n32134;
  assign n32136 = ~n15020 & ~n32135;
  assign n32137 = controllable_hmaster2 & ~n32136;
  assign n32138 = ~i_hbusreq9 & ~n22048;
  assign n32139 = ~n30571 & ~n32138;
  assign n32140 = ~i_hbusreq4 & ~n32139;
  assign n32141 = ~n30570 & ~n32140;
  assign n32142 = ~controllable_hgrant4 & ~n32141;
  assign n32143 = ~n15030 & ~n32142;
  assign n32144 = ~i_hbusreq5 & ~n32143;
  assign n32145 = ~n30569 & ~n32144;
  assign n32146 = ~controllable_hgrant5 & ~n32145;
  assign n32147 = ~n15029 & ~n32146;
  assign n32148 = ~controllable_hmaster2 & ~n32147;
  assign n32149 = ~n32137 & ~n32148;
  assign n32150 = ~controllable_hmaster1 & ~n32149;
  assign n32151 = ~n32129 & ~n32150;
  assign n32152 = ~i_hbusreq6 & ~n32151;
  assign n32153 = ~n30543 & ~n32152;
  assign n32154 = ~controllable_hgrant6 & ~n32153;
  assign n32155 = ~n14995 & ~n32154;
  assign n32156 = controllable_hmaster0 & ~n32155;
  assign n32157 = controllable_hmaster2 & ~n32080;
  assign n32158 = ~i_hbusreq9 & ~n22090;
  assign n32159 = ~n30595 & ~n32158;
  assign n32160 = ~i_hbusreq4 & ~n32159;
  assign n32161 = ~n30594 & ~n32160;
  assign n32162 = ~controllable_hgrant4 & ~n32161;
  assign n32163 = ~n15065 & ~n32162;
  assign n32164 = ~i_hbusreq5 & ~n32163;
  assign n32165 = ~n30593 & ~n32164;
  assign n32166 = ~controllable_hgrant5 & ~n32165;
  assign n32167 = ~n15064 & ~n32166;
  assign n32168 = ~controllable_hmaster2 & ~n32167;
  assign n32169 = ~n32157 & ~n32168;
  assign n32170 = controllable_hmaster1 & ~n32169;
  assign n32171 = i_hlock4 & ~n32072;
  assign n32172 = ~i_hlock4 & ~n32093;
  assign n32173 = ~n32171 & ~n32172;
  assign n32174 = ~i_hbusreq4 & ~n32173;
  assign n32175 = ~n30610 & ~n32174;
  assign n32176 = ~controllable_hgrant4 & ~n32175;
  assign n32177 = ~n15091 & ~n32176;
  assign n32178 = ~i_hbusreq5 & ~n32177;
  assign n32179 = ~n30609 & ~n32178;
  assign n32180 = ~controllable_hgrant5 & ~n32179;
  assign n32181 = ~n15090 & ~n32180;
  assign n32182 = controllable_hmaster2 & ~n32181;
  assign n32183 = ~i_hbusreq9 & ~n22145;
  assign n32184 = ~n30625 & ~n32183;
  assign n32185 = ~i_hbusreq4 & ~n32184;
  assign n32186 = ~n30624 & ~n32185;
  assign n32187 = ~controllable_hgrant4 & ~n32186;
  assign n32188 = ~n15105 & ~n32187;
  assign n32189 = ~i_hbusreq5 & ~n32188;
  assign n32190 = ~n30623 & ~n32189;
  assign n32191 = ~controllable_hgrant5 & ~n32190;
  assign n32192 = ~n15104 & ~n32191;
  assign n32193 = ~controllable_hmaster2 & ~n32192;
  assign n32194 = ~n32182 & ~n32193;
  assign n32195 = ~controllable_hmaster1 & ~n32194;
  assign n32196 = ~n32170 & ~n32195;
  assign n32197 = i_hlock6 & ~n32196;
  assign n32198 = controllable_hmaster2 & ~n32101;
  assign n32199 = ~n32168 & ~n32198;
  assign n32200 = controllable_hmaster1 & ~n32199;
  assign n32201 = ~n32195 & ~n32200;
  assign n32202 = ~i_hlock6 & ~n32201;
  assign n32203 = ~n32197 & ~n32202;
  assign n32204 = ~i_hbusreq6 & ~n32203;
  assign n32205 = ~n30591 & ~n32204;
  assign n32206 = ~controllable_hgrant6 & ~n32205;
  assign n32207 = ~n15063 & ~n32206;
  assign n32208 = ~controllable_hmaster0 & ~n32207;
  assign n32209 = ~n32156 & ~n32208;
  assign n32210 = ~i_hbusreq8 & ~n32209;
  assign n32211 = ~n30542 & ~n32210;
  assign n32212 = ~controllable_hmaster3 & ~n32211;
  assign n32213 = ~n32116 & ~n32212;
  assign n32214 = i_hlock7 & ~n32213;
  assign n32215 = ~i_hbusreq9 & ~n21884;
  assign n32216 = ~n29619 & ~n32215;
  assign n32217 = ~i_hbusreq4 & ~n32216;
  assign n32218 = ~n29618 & ~n32217;
  assign n32219 = ~controllable_hgrant4 & ~n32218;
  assign n32220 = ~n14875 & ~n32219;
  assign n32221 = ~i_hbusreq5 & ~n32220;
  assign n32222 = ~n29617 & ~n32221;
  assign n32223 = ~controllable_hgrant5 & ~n32222;
  assign n32224 = ~n14874 & ~n32223;
  assign n32225 = controllable_hmaster1 & ~n32224;
  assign n32226 = controllable_hmaster2 & ~n32224;
  assign n32227 = i_hlock9 & ~n21929;
  assign n32228 = ~n21972 & ~n32227;
  assign n32229 = ~i_hbusreq9 & ~n32228;
  assign n32230 = ~n30674 & ~n32229;
  assign n32231 = ~i_hbusreq4 & ~n32230;
  assign n32232 = ~n30673 & ~n32231;
  assign n32233 = ~controllable_hgrant4 & ~n32232;
  assign n32234 = ~n12676 & ~n32233;
  assign n32235 = ~i_hbusreq5 & ~n32234;
  assign n32236 = ~n30672 & ~n32235;
  assign n32237 = ~controllable_hgrant5 & ~n32236;
  assign n32238 = ~n12674 & ~n32237;
  assign n32239 = ~controllable_hmaster2 & ~n32238;
  assign n32240 = ~n32226 & ~n32239;
  assign n32241 = ~controllable_hmaster1 & ~n32240;
  assign n32242 = ~n32225 & ~n32241;
  assign n32243 = ~i_hbusreq6 & ~n32242;
  assign n32244 = ~n30659 & ~n32243;
  assign n32245 = ~controllable_hgrant6 & ~n32244;
  assign n32246 = ~n14849 & ~n32245;
  assign n32247 = controllable_hmaster0 & ~n32246;
  assign n32248 = ~i_hbusreq9 & ~n21929;
  assign n32249 = ~n30699 & ~n32248;
  assign n32250 = ~i_hbusreq4 & ~n32249;
  assign n32251 = ~n30698 & ~n32250;
  assign n32252 = ~controllable_hgrant4 & ~n32251;
  assign n32253 = ~n13524 & ~n32252;
  assign n32254 = ~i_hbusreq5 & ~n32253;
  assign n32255 = ~n30697 & ~n32254;
  assign n32256 = ~controllable_hgrant5 & ~n32255;
  assign n32257 = ~n13522 & ~n32256;
  assign n32258 = ~controllable_hmaster2 & ~n32257;
  assign n32259 = ~n32226 & ~n32258;
  assign n32260 = ~controllable_hmaster1 & ~n32259;
  assign n32261 = ~n32225 & ~n32260;
  assign n32262 = ~i_hbusreq6 & ~n32261;
  assign n32263 = ~n30696 & ~n32262;
  assign n32264 = ~controllable_hgrant6 & ~n32263;
  assign n32265 = ~n14927 & ~n32264;
  assign n32266 = ~controllable_hmaster0 & ~n32265;
  assign n32267 = ~n32247 & ~n32266;
  assign n32268 = i_hlock8 & ~n32267;
  assign n32269 = ~i_hbusreq9 & ~n21971;
  assign n32270 = ~n30724 & ~n32269;
  assign n32271 = ~i_hbusreq4 & ~n32270;
  assign n32272 = ~n30723 & ~n32271;
  assign n32273 = ~controllable_hgrant4 & ~n32272;
  assign n32274 = ~n13577 & ~n32273;
  assign n32275 = ~i_hbusreq5 & ~n32274;
  assign n32276 = ~n30722 & ~n32275;
  assign n32277 = ~controllable_hgrant5 & ~n32276;
  assign n32278 = ~n13575 & ~n32277;
  assign n32279 = ~controllable_hmaster2 & ~n32278;
  assign n32280 = ~n32226 & ~n32279;
  assign n32281 = ~controllable_hmaster1 & ~n32280;
  assign n32282 = ~n32225 & ~n32281;
  assign n32283 = ~i_hbusreq6 & ~n32282;
  assign n32284 = ~n30721 & ~n32283;
  assign n32285 = ~controllable_hgrant6 & ~n32284;
  assign n32286 = ~n14960 & ~n32285;
  assign n32287 = ~controllable_hmaster0 & ~n32286;
  assign n32288 = ~n32247 & ~n32287;
  assign n32289 = ~i_hlock8 & ~n32288;
  assign n32290 = ~n32268 & ~n32289;
  assign n32291 = ~i_hbusreq8 & ~n32290;
  assign n32292 = ~n30658 & ~n32291;
  assign n32293 = controllable_hmaster3 & ~n32292;
  assign n32294 = ~i_hbusreq9 & ~n22014;
  assign n32295 = ~n30754 & ~n32294;
  assign n32296 = ~i_hbusreq4 & ~n32295;
  assign n32297 = ~n30753 & ~n32296;
  assign n32298 = ~controllable_hgrant4 & ~n32297;
  assign n32299 = ~n14998 & ~n32298;
  assign n32300 = ~i_hbusreq5 & ~n32299;
  assign n32301 = ~n30752 & ~n32300;
  assign n32302 = ~controllable_hgrant5 & ~n32301;
  assign n32303 = ~n14997 & ~n32302;
  assign n32304 = ~controllable_hmaster2 & ~n32303;
  assign n32305 = ~n29106 & ~n32304;
  assign n32306 = controllable_hmaster1 & ~n32305;
  assign n32307 = i_hlock5 & ~n32253;
  assign n32308 = ~i_hlock5 & ~n32274;
  assign n32309 = ~n32307 & ~n32308;
  assign n32310 = ~i_hbusreq5 & ~n32309;
  assign n32311 = ~n30768 & ~n32310;
  assign n32312 = ~controllable_hgrant5 & ~n32311;
  assign n32313 = ~n15020 & ~n32312;
  assign n32314 = controllable_hmaster2 & ~n32313;
  assign n32315 = ~i_hbusreq9 & ~n22060;
  assign n32316 = ~n30779 & ~n32315;
  assign n32317 = ~i_hbusreq4 & ~n32316;
  assign n32318 = ~n30778 & ~n32317;
  assign n32319 = ~controllable_hgrant4 & ~n32318;
  assign n32320 = ~n15030 & ~n32319;
  assign n32321 = ~i_hbusreq5 & ~n32320;
  assign n32322 = ~n30777 & ~n32321;
  assign n32323 = ~controllable_hgrant5 & ~n32322;
  assign n32324 = ~n15029 & ~n32323;
  assign n32325 = ~controllable_hmaster2 & ~n32324;
  assign n32326 = ~n32314 & ~n32325;
  assign n32327 = ~controllable_hmaster1 & ~n32326;
  assign n32328 = ~n32306 & ~n32327;
  assign n32329 = ~i_hbusreq6 & ~n32328;
  assign n32330 = ~n30751 & ~n32329;
  assign n32331 = ~controllable_hgrant6 & ~n32330;
  assign n32332 = ~n15152 & ~n32331;
  assign n32333 = controllable_hmaster0 & ~n32332;
  assign n32334 = controllable_hmaster2 & ~n32257;
  assign n32335 = ~i_hbusreq9 & ~n22100;
  assign n32336 = ~n30803 & ~n32335;
  assign n32337 = ~i_hbusreq4 & ~n32336;
  assign n32338 = ~n30802 & ~n32337;
  assign n32339 = ~controllable_hgrant4 & ~n32338;
  assign n32340 = ~n15065 & ~n32339;
  assign n32341 = ~i_hbusreq5 & ~n32340;
  assign n32342 = ~n30801 & ~n32341;
  assign n32343 = ~controllable_hgrant5 & ~n32342;
  assign n32344 = ~n15064 & ~n32343;
  assign n32345 = ~controllable_hmaster2 & ~n32344;
  assign n32346 = ~n32334 & ~n32345;
  assign n32347 = controllable_hmaster1 & ~n32346;
  assign n32348 = i_hlock4 & ~n32249;
  assign n32349 = ~i_hlock4 & ~n32270;
  assign n32350 = ~n32348 & ~n32349;
  assign n32351 = ~i_hbusreq4 & ~n32350;
  assign n32352 = ~n30818 & ~n32351;
  assign n32353 = ~controllable_hgrant4 & ~n32352;
  assign n32354 = ~n15091 & ~n32353;
  assign n32355 = ~i_hbusreq5 & ~n32354;
  assign n32356 = ~n30817 & ~n32355;
  assign n32357 = ~controllable_hgrant5 & ~n32356;
  assign n32358 = ~n15090 & ~n32357;
  assign n32359 = controllable_hmaster2 & ~n32358;
  assign n32360 = ~i_hbusreq9 & ~n22157;
  assign n32361 = ~n30833 & ~n32360;
  assign n32362 = ~i_hbusreq4 & ~n32361;
  assign n32363 = ~n30832 & ~n32362;
  assign n32364 = ~controllable_hgrant4 & ~n32363;
  assign n32365 = ~n15105 & ~n32364;
  assign n32366 = ~i_hbusreq5 & ~n32365;
  assign n32367 = ~n30831 & ~n32366;
  assign n32368 = ~controllable_hgrant5 & ~n32367;
  assign n32369 = ~n15104 & ~n32368;
  assign n32370 = ~controllable_hmaster2 & ~n32369;
  assign n32371 = ~n32359 & ~n32370;
  assign n32372 = ~controllable_hmaster1 & ~n32371;
  assign n32373 = ~n32347 & ~n32372;
  assign n32374 = i_hlock6 & ~n32373;
  assign n32375 = controllable_hmaster2 & ~n32278;
  assign n32376 = ~n32345 & ~n32375;
  assign n32377 = controllable_hmaster1 & ~n32376;
  assign n32378 = ~n32372 & ~n32377;
  assign n32379 = ~i_hlock6 & ~n32378;
  assign n32380 = ~n32374 & ~n32379;
  assign n32381 = ~i_hbusreq6 & ~n32380;
  assign n32382 = ~n30799 & ~n32381;
  assign n32383 = ~controllable_hgrant6 & ~n32382;
  assign n32384 = ~n15063 & ~n32383;
  assign n32385 = ~controllable_hmaster0 & ~n32384;
  assign n32386 = ~n32333 & ~n32385;
  assign n32387 = ~i_hbusreq8 & ~n32386;
  assign n32388 = ~n30750 & ~n32387;
  assign n32389 = ~controllable_hmaster3 & ~n32388;
  assign n32390 = ~n32293 & ~n32389;
  assign n32391 = ~i_hlock7 & ~n32390;
  assign n32392 = ~n32214 & ~n32391;
  assign n32393 = ~i_hbusreq7 & ~n32392;
  assign n32394 = ~n30449 & ~n32393;
  assign n32395 = n7924 & ~n32394;
  assign n32396 = ~n32037 & ~n32395;
  assign n32397 = n7920 & ~n32396;
  assign n32398 = ~n28799 & ~n32397;
  assign n32399 = ~n7728 & ~n32398;
  assign n32400 = ~n31989 & ~n32399;
  assign n32401 = ~n7723 & ~n32400;
  assign n32402 = ~n30971 & ~n32401;
  assign n32403 = ~n7714 & ~n32402;
  assign n32404 = ~n30970 & ~n32403;
  assign n32405 = ~n7705 & ~n32404;
  assign n32406 = ~n29290 & ~n32405;
  assign n32407 = n7808 & ~n32406;
  assign n32408 = ~n28809 & ~n32407;
  assign n32409 = n8195 & ~n32408;
  assign n32410 = ~n8196 & ~n32409;
  assign n32411 = ~n8193 & ~n32410;
  assign n32412 = ~n9900 & ~n28799;
  assign n32413 = ~n7723 & ~n32412;
  assign n32414 = ~n9899 & ~n32413;
  assign n32415 = n7714 & ~n32414;
  assign n32416 = ~n28805 & ~n32415;
  assign n32417 = ~n7705 & ~n32416;
  assign n32418 = ~n9898 & ~n32417;
  assign n32419 = ~n7808 & ~n32418;
  assign n32420 = ~n22401 & ~n26890;
  assign n32421 = ~controllable_hgrant6 & ~n32420;
  assign n32422 = ~n15193 & ~n32421;
  assign n32423 = controllable_hmaster0 & ~n32422;
  assign n32424 = ~n9099 & ~n32423;
  assign n32425 = ~controllable_hmaster3 & ~n32424;
  assign n32426 = ~n9093 & ~n32425;
  assign n32427 = i_hbusreq7 & ~n32426;
  assign n32428 = i_hbusreq8 & ~n32424;
  assign n32429 = i_hbusreq6 & ~n32420;
  assign n32430 = ~n22413 & ~n26903;
  assign n32431 = ~i_hbusreq6 & ~n32430;
  assign n32432 = ~n32429 & ~n32431;
  assign n32433 = ~controllable_hgrant6 & ~n32432;
  assign n32434 = ~n15206 & ~n32433;
  assign n32435 = controllable_hmaster0 & ~n32434;
  assign n32436 = ~n9127 & ~n32435;
  assign n32437 = ~i_hbusreq8 & ~n32436;
  assign n32438 = ~n32428 & ~n32437;
  assign n32439 = ~controllable_hmaster3 & ~n32438;
  assign n32440 = ~n9117 & ~n32439;
  assign n32441 = ~i_hbusreq7 & ~n32440;
  assign n32442 = ~n32427 & ~n32441;
  assign n32443 = ~n7924 & ~n32442;
  assign n32444 = ~n22435 & ~n26936;
  assign n32445 = ~controllable_hgrant6 & ~n32444;
  assign n32446 = ~n15193 & ~n32445;
  assign n32447 = controllable_hmaster0 & ~n32446;
  assign n32448 = ~n13682 & ~n32447;
  assign n32449 = ~controllable_hmaster3 & ~n32448;
  assign n32450 = ~n27088 & ~n32449;
  assign n32451 = i_hbusreq7 & ~n32450;
  assign n32452 = i_hbusreq8 & ~n32448;
  assign n32453 = i_hbusreq6 & ~n32444;
  assign n32454 = ~n22456 & ~n26980;
  assign n32455 = ~i_hbusreq6 & ~n32454;
  assign n32456 = ~n32453 & ~n32455;
  assign n32457 = ~controllable_hgrant6 & ~n32456;
  assign n32458 = ~n15206 & ~n32457;
  assign n32459 = controllable_hmaster0 & ~n32458;
  assign n32460 = ~n13728 & ~n32459;
  assign n32461 = ~i_hbusreq8 & ~n32460;
  assign n32462 = ~n32452 & ~n32461;
  assign n32463 = ~controllable_hmaster3 & ~n32462;
  assign n32464 = ~n27174 & ~n32463;
  assign n32465 = ~i_hbusreq7 & ~n32464;
  assign n32466 = ~n32451 & ~n32465;
  assign n32467 = n7924 & ~n32466;
  assign n32468 = ~n32443 & ~n32467;
  assign n32469 = ~n8214 & ~n32468;
  assign n32470 = ~n22478 & ~n26894;
  assign n32471 = ~controllable_hmaster3 & ~n32470;
  assign n32472 = ~n9093 & ~n32471;
  assign n32473 = i_hbusreq7 & ~n32472;
  assign n32474 = i_hbusreq8 & ~n32470;
  assign n32475 = ~n22492 & ~n26909;
  assign n32476 = ~i_hbusreq8 & ~n32475;
  assign n32477 = ~n32474 & ~n32476;
  assign n32478 = ~controllable_hmaster3 & ~n32477;
  assign n32479 = ~n9117 & ~n32478;
  assign n32480 = ~i_hbusreq7 & ~n32479;
  assign n32481 = ~n32473 & ~n32480;
  assign n32482 = ~n7924 & ~n32481;
  assign n32483 = ~n22514 & ~n26940;
  assign n32484 = ~controllable_hmaster3 & ~n32483;
  assign n32485 = ~n27088 & ~n32484;
  assign n32486 = i_hbusreq7 & ~n32485;
  assign n32487 = i_hbusreq8 & ~n32483;
  assign n32488 = ~n22542 & ~n26986;
  assign n32489 = ~i_hbusreq8 & ~n32488;
  assign n32490 = ~n32487 & ~n32489;
  assign n32491 = ~controllable_hmaster3 & ~n32490;
  assign n32492 = ~n27174 & ~n32491;
  assign n32493 = ~i_hbusreq7 & ~n32492;
  assign n32494 = ~n32486 & ~n32493;
  assign n32495 = n7924 & ~n32494;
  assign n32496 = ~n32482 & ~n32495;
  assign n32497 = n8214 & ~n32496;
  assign n32498 = ~n32469 & ~n32497;
  assign n32499 = ~n8202 & ~n32498;
  assign n32500 = ~n18123 & ~n26888;
  assign n32501 = controllable_hmaster1 & ~n32500;
  assign n32502 = ~n9096 & ~n32501;
  assign n32503 = ~controllable_hgrant6 & ~n32502;
  assign n32504 = ~n15293 & ~n32503;
  assign n32505 = controllable_hmaster0 & ~n32504;
  assign n32506 = ~n9099 & ~n32505;
  assign n32507 = ~controllable_hmaster3 & ~n32506;
  assign n32508 = ~n9093 & ~n32507;
  assign n32509 = i_hbusreq7 & ~n32508;
  assign n32510 = i_hbusreq8 & ~n32506;
  assign n32511 = i_hbusreq6 & ~n32502;
  assign n32512 = ~n21699 & ~n26901;
  assign n32513 = controllable_hmaster1 & ~n32512;
  assign n32514 = ~n9122 & ~n32513;
  assign n32515 = ~i_hbusreq6 & ~n32514;
  assign n32516 = ~n32511 & ~n32515;
  assign n32517 = ~controllable_hgrant6 & ~n32516;
  assign n32518 = ~n15306 & ~n32517;
  assign n32519 = controllable_hmaster0 & ~n32518;
  assign n32520 = ~n9127 & ~n32519;
  assign n32521 = ~i_hbusreq8 & ~n32520;
  assign n32522 = ~n32510 & ~n32521;
  assign n32523 = ~controllable_hmaster3 & ~n32522;
  assign n32524 = ~n9117 & ~n32523;
  assign n32525 = ~i_hbusreq7 & ~n32524;
  assign n32526 = ~n32509 & ~n32525;
  assign n32527 = ~n7924 & ~n32526;
  assign n32528 = ~n22592 & ~n26934;
  assign n32529 = controllable_hmaster1 & ~n32528;
  assign n32530 = ~n13677 & ~n32529;
  assign n32531 = ~controllable_hgrant6 & ~n32530;
  assign n32532 = ~n15293 & ~n32531;
  assign n32533 = controllable_hmaster0 & ~n32532;
  assign n32534 = ~n13682 & ~n32533;
  assign n32535 = ~controllable_hmaster3 & ~n32534;
  assign n32536 = ~n27088 & ~n32535;
  assign n32537 = i_hbusreq7 & ~n32536;
  assign n32538 = i_hbusreq8 & ~n32534;
  assign n32539 = i_hbusreq6 & ~n32530;
  assign n32540 = ~n22626 & ~n26978;
  assign n32541 = controllable_hmaster1 & ~n32540;
  assign n32542 = ~n13721 & ~n32541;
  assign n32543 = ~i_hbusreq6 & ~n32542;
  assign n32544 = ~n32539 & ~n32543;
  assign n32545 = ~controllable_hgrant6 & ~n32544;
  assign n32546 = ~n15306 & ~n32545;
  assign n32547 = controllable_hmaster0 & ~n32546;
  assign n32548 = ~n13728 & ~n32547;
  assign n32549 = ~i_hbusreq8 & ~n32548;
  assign n32550 = ~n32538 & ~n32549;
  assign n32551 = ~controllable_hmaster3 & ~n32550;
  assign n32552 = ~n27174 & ~n32551;
  assign n32553 = ~i_hbusreq7 & ~n32552;
  assign n32554 = ~n32537 & ~n32553;
  assign n32555 = n7924 & ~n32554;
  assign n32556 = ~n32527 & ~n32555;
  assign n32557 = ~n8214 & ~n32556;
  assign n32558 = ~n22650 & ~n26894;
  assign n32559 = ~controllable_hmaster3 & ~n32558;
  assign n32560 = ~n9093 & ~n32559;
  assign n32561 = i_hbusreq7 & ~n32560;
  assign n32562 = i_hbusreq8 & ~n32558;
  assign n32563 = ~n22664 & ~n26909;
  assign n32564 = ~i_hbusreq8 & ~n32563;
  assign n32565 = ~n32562 & ~n32564;
  assign n32566 = ~controllable_hmaster3 & ~n32565;
  assign n32567 = ~n9117 & ~n32566;
  assign n32568 = ~i_hbusreq7 & ~n32567;
  assign n32569 = ~n32561 & ~n32568;
  assign n32570 = ~n7924 & ~n32569;
  assign n32571 = ~n22688 & ~n26940;
  assign n32572 = ~controllable_hmaster3 & ~n32571;
  assign n32573 = ~n27088 & ~n32572;
  assign n32574 = i_hbusreq7 & ~n32573;
  assign n32575 = i_hbusreq8 & ~n32571;
  assign n32576 = ~n22727 & ~n26986;
  assign n32577 = ~i_hbusreq8 & ~n32576;
  assign n32578 = ~n32575 & ~n32577;
  assign n32579 = ~controllable_hmaster3 & ~n32578;
  assign n32580 = ~n27174 & ~n32579;
  assign n32581 = ~i_hbusreq7 & ~n32580;
  assign n32582 = ~n32574 & ~n32581;
  assign n32583 = n7924 & ~n32582;
  assign n32584 = ~n32570 & ~n32583;
  assign n32585 = n8214 & ~n32584;
  assign n32586 = ~n32557 & ~n32585;
  assign n32587 = n8202 & ~n32586;
  assign n32588 = ~n32499 & ~n32587;
  assign n32589 = n7920 & ~n32588;
  assign n32590 = ~n10014 & ~n32589;
  assign n32591 = n7728 & ~n32590;
  assign n32592 = ~n22745 & ~n29737;
  assign n32593 = ~controllable_hgrant6 & ~n32592;
  assign n32594 = ~n13849 & ~n32593;
  assign n32595 = controllable_hmaster0 & ~n32594;
  assign n32596 = ~n19324 & ~n32595;
  assign n32597 = ~controllable_hmaster3 & ~n32596;
  assign n32598 = ~n30877 & ~n32597;
  assign n32599 = i_hlock7 & ~n32598;
  assign n32600 = ~n22745 & ~n29752;
  assign n32601 = ~controllable_hgrant6 & ~n32600;
  assign n32602 = ~n13951 & ~n32601;
  assign n32603 = controllable_hmaster0 & ~n32602;
  assign n32604 = ~n19324 & ~n32603;
  assign n32605 = ~controllable_hmaster3 & ~n32604;
  assign n32606 = ~n30877 & ~n32605;
  assign n32607 = ~i_hlock7 & ~n32606;
  assign n32608 = ~n32599 & ~n32607;
  assign n32609 = i_hbusreq7 & ~n32608;
  assign n32610 = i_hbusreq8 & ~n32596;
  assign n32611 = i_hbusreq6 & ~n32592;
  assign n32612 = ~n22767 & ~n29798;
  assign n32613 = ~i_hbusreq6 & ~n32612;
  assign n32614 = ~n32611 & ~n32613;
  assign n32615 = ~controllable_hgrant6 & ~n32614;
  assign n32616 = ~n15417 & ~n32615;
  assign n32617 = controllable_hmaster0 & ~n32616;
  assign n32618 = ~n19644 & ~n32617;
  assign n32619 = ~i_hbusreq8 & ~n32618;
  assign n32620 = ~n32610 & ~n32619;
  assign n32621 = ~controllable_hmaster3 & ~n32620;
  assign n32622 = ~n30896 & ~n32621;
  assign n32623 = i_hlock7 & ~n32622;
  assign n32624 = i_hbusreq8 & ~n32604;
  assign n32625 = i_hbusreq6 & ~n32600;
  assign n32626 = ~n22767 & ~n29828;
  assign n32627 = ~i_hbusreq6 & ~n32626;
  assign n32628 = ~n32625 & ~n32627;
  assign n32629 = ~controllable_hgrant6 & ~n32628;
  assign n32630 = ~n15440 & ~n32629;
  assign n32631 = controllable_hmaster0 & ~n32630;
  assign n32632 = ~n19644 & ~n32631;
  assign n32633 = ~i_hbusreq8 & ~n32632;
  assign n32634 = ~n32624 & ~n32633;
  assign n32635 = ~controllable_hmaster3 & ~n32634;
  assign n32636 = ~n30896 & ~n32635;
  assign n32637 = ~i_hlock7 & ~n32636;
  assign n32638 = ~n32623 & ~n32637;
  assign n32639 = ~i_hbusreq7 & ~n32638;
  assign n32640 = ~n32609 & ~n32639;
  assign n32641 = ~n7924 & ~n32640;
  assign n32642 = ~n22805 & ~n29871;
  assign n32643 = ~controllable_hgrant6 & ~n32642;
  assign n32644 = ~n13849 & ~n32643;
  assign n32645 = controllable_hmaster0 & ~n32644;
  assign n32646 = ~n19849 & ~n32645;
  assign n32647 = ~controllable_hmaster3 & ~n32646;
  assign n32648 = ~n30920 & ~n32647;
  assign n32649 = i_hlock7 & ~n32648;
  assign n32650 = ~n22805 & ~n29886;
  assign n32651 = ~controllable_hgrant6 & ~n32650;
  assign n32652 = ~n13951 & ~n32651;
  assign n32653 = controllable_hmaster0 & ~n32652;
  assign n32654 = ~n19849 & ~n32653;
  assign n32655 = ~controllable_hmaster3 & ~n32654;
  assign n32656 = ~n30920 & ~n32655;
  assign n32657 = ~i_hlock7 & ~n32656;
  assign n32658 = ~n32649 & ~n32657;
  assign n32659 = i_hbusreq7 & ~n32658;
  assign n32660 = i_hbusreq8 & ~n32646;
  assign n32661 = i_hbusreq6 & ~n32642;
  assign n32662 = ~n22836 & ~n29949;
  assign n32663 = ~i_hbusreq6 & ~n32662;
  assign n32664 = ~n32661 & ~n32663;
  assign n32665 = ~controllable_hgrant6 & ~n32664;
  assign n32666 = ~n15417 & ~n32665;
  assign n32667 = controllable_hmaster0 & ~n32666;
  assign n32668 = ~n20237 & ~n32667;
  assign n32669 = ~i_hbusreq8 & ~n32668;
  assign n32670 = ~n32660 & ~n32669;
  assign n32671 = ~controllable_hmaster3 & ~n32670;
  assign n32672 = ~n30939 & ~n32671;
  assign n32673 = i_hlock7 & ~n32672;
  assign n32674 = i_hbusreq8 & ~n32654;
  assign n32675 = i_hbusreq6 & ~n32650;
  assign n32676 = ~n22836 & ~n29979;
  assign n32677 = ~i_hbusreq6 & ~n32676;
  assign n32678 = ~n32675 & ~n32677;
  assign n32679 = ~controllable_hgrant6 & ~n32678;
  assign n32680 = ~n15440 & ~n32679;
  assign n32681 = controllable_hmaster0 & ~n32680;
  assign n32682 = ~n20237 & ~n32681;
  assign n32683 = ~i_hbusreq8 & ~n32682;
  assign n32684 = ~n32674 & ~n32683;
  assign n32685 = ~controllable_hmaster3 & ~n32684;
  assign n32686 = ~n30939 & ~n32685;
  assign n32687 = ~i_hlock7 & ~n32686;
  assign n32688 = ~n32673 & ~n32687;
  assign n32689 = ~i_hbusreq7 & ~n32688;
  assign n32690 = ~n32659 & ~n32689;
  assign n32691 = n7924 & ~n32690;
  assign n32692 = ~n32641 & ~n32691;
  assign n32693 = ~n8214 & ~n32692;
  assign n32694 = ~n22878 & ~n29741;
  assign n32695 = ~controllable_hmaster3 & ~n32694;
  assign n32696 = ~n30877 & ~n32695;
  assign n32697 = i_hlock7 & ~n32696;
  assign n32698 = ~n22878 & ~n29756;
  assign n32699 = ~controllable_hmaster3 & ~n32698;
  assign n32700 = ~n30877 & ~n32699;
  assign n32701 = ~i_hlock7 & ~n32700;
  assign n32702 = ~n32697 & ~n32701;
  assign n32703 = i_hbusreq7 & ~n32702;
  assign n32704 = i_hbusreq8 & ~n32694;
  assign n32705 = ~n22902 & ~n29804;
  assign n32706 = ~i_hbusreq8 & ~n32705;
  assign n32707 = ~n32704 & ~n32706;
  assign n32708 = ~controllable_hmaster3 & ~n32707;
  assign n32709 = ~n30896 & ~n32708;
  assign n32710 = i_hlock7 & ~n32709;
  assign n32711 = i_hbusreq8 & ~n32698;
  assign n32712 = ~n22902 & ~n29834;
  assign n32713 = ~i_hbusreq8 & ~n32712;
  assign n32714 = ~n32711 & ~n32713;
  assign n32715 = ~controllable_hmaster3 & ~n32714;
  assign n32716 = ~n30896 & ~n32715;
  assign n32717 = ~i_hlock7 & ~n32716;
  assign n32718 = ~n32710 & ~n32717;
  assign n32719 = ~i_hbusreq7 & ~n32718;
  assign n32720 = ~n32703 & ~n32719;
  assign n32721 = ~n7924 & ~n32720;
  assign n32722 = ~n22937 & ~n29875;
  assign n32723 = ~controllable_hmaster3 & ~n32722;
  assign n32724 = ~n30920 & ~n32723;
  assign n32725 = i_hlock7 & ~n32724;
  assign n32726 = ~n22937 & ~n29890;
  assign n32727 = ~controllable_hmaster3 & ~n32726;
  assign n32728 = ~n30920 & ~n32727;
  assign n32729 = ~i_hlock7 & ~n32728;
  assign n32730 = ~n32725 & ~n32729;
  assign n32731 = i_hbusreq7 & ~n32730;
  assign n32732 = i_hbusreq8 & ~n32722;
  assign n32733 = ~n22975 & ~n29955;
  assign n32734 = ~i_hbusreq8 & ~n32733;
  assign n32735 = ~n32732 & ~n32734;
  assign n32736 = ~controllable_hmaster3 & ~n32735;
  assign n32737 = ~n30939 & ~n32736;
  assign n32738 = i_hlock7 & ~n32737;
  assign n32739 = i_hbusreq8 & ~n32726;
  assign n32740 = ~n22975 & ~n29985;
  assign n32741 = ~i_hbusreq8 & ~n32740;
  assign n32742 = ~n32739 & ~n32741;
  assign n32743 = ~controllable_hmaster3 & ~n32742;
  assign n32744 = ~n30939 & ~n32743;
  assign n32745 = ~i_hlock7 & ~n32744;
  assign n32746 = ~n32738 & ~n32745;
  assign n32747 = ~i_hbusreq7 & ~n32746;
  assign n32748 = ~n32731 & ~n32747;
  assign n32749 = n7924 & ~n32748;
  assign n32750 = ~n32721 & ~n32749;
  assign n32751 = n8214 & ~n32750;
  assign n32752 = ~n32693 & ~n32751;
  assign n32753 = ~n8202 & ~n32752;
  assign n32754 = ~n18123 & ~n29735;
  assign n32755 = controllable_hmaster1 & ~n32754;
  assign n32756 = ~n19275 & ~n32755;
  assign n32757 = ~controllable_hgrant6 & ~n32756;
  assign n32758 = ~n13849 & ~n32757;
  assign n32759 = controllable_hmaster0 & ~n32758;
  assign n32760 = ~n19324 & ~n32759;
  assign n32761 = ~controllable_hmaster3 & ~n32760;
  assign n32762 = ~n30877 & ~n32761;
  assign n32763 = i_hlock7 & ~n32762;
  assign n32764 = ~n18123 & ~n29750;
  assign n32765 = controllable_hmaster1 & ~n32764;
  assign n32766 = ~n19275 & ~n32765;
  assign n32767 = ~controllable_hgrant6 & ~n32766;
  assign n32768 = ~n13951 & ~n32767;
  assign n32769 = controllable_hmaster0 & ~n32768;
  assign n32770 = ~n19324 & ~n32769;
  assign n32771 = ~controllable_hmaster3 & ~n32770;
  assign n32772 = ~n30877 & ~n32771;
  assign n32773 = ~i_hlock7 & ~n32772;
  assign n32774 = ~n32763 & ~n32773;
  assign n32775 = i_hbusreq7 & ~n32774;
  assign n32776 = i_hbusreq8 & ~n32760;
  assign n32777 = i_hbusreq6 & ~n32756;
  assign n32778 = ~n21699 & ~n29796;
  assign n32779 = controllable_hmaster1 & ~n32778;
  assign n32780 = ~n19550 & ~n32779;
  assign n32781 = ~i_hbusreq6 & ~n32780;
  assign n32782 = ~n32777 & ~n32781;
  assign n32783 = ~controllable_hgrant6 & ~n32782;
  assign n32784 = ~n15520 & ~n32783;
  assign n32785 = controllable_hmaster0 & ~n32784;
  assign n32786 = ~n19644 & ~n32785;
  assign n32787 = ~i_hbusreq8 & ~n32786;
  assign n32788 = ~n32776 & ~n32787;
  assign n32789 = ~controllable_hmaster3 & ~n32788;
  assign n32790 = ~n30896 & ~n32789;
  assign n32791 = i_hlock7 & ~n32790;
  assign n32792 = i_hbusreq8 & ~n32770;
  assign n32793 = i_hbusreq6 & ~n32766;
  assign n32794 = ~n21699 & ~n29826;
  assign n32795 = controllable_hmaster1 & ~n32794;
  assign n32796 = ~n19550 & ~n32795;
  assign n32797 = ~i_hbusreq6 & ~n32796;
  assign n32798 = ~n32793 & ~n32797;
  assign n32799 = ~controllable_hgrant6 & ~n32798;
  assign n32800 = ~n15553 & ~n32799;
  assign n32801 = controllable_hmaster0 & ~n32800;
  assign n32802 = ~n19644 & ~n32801;
  assign n32803 = ~i_hbusreq8 & ~n32802;
  assign n32804 = ~n32792 & ~n32803;
  assign n32805 = ~controllable_hmaster3 & ~n32804;
  assign n32806 = ~n30896 & ~n32805;
  assign n32807 = ~i_hlock7 & ~n32806;
  assign n32808 = ~n32791 & ~n32807;
  assign n32809 = ~i_hbusreq7 & ~n32808;
  assign n32810 = ~n32775 & ~n32809;
  assign n32811 = ~n7924 & ~n32810;
  assign n32812 = ~n23064 & ~n29869;
  assign n32813 = controllable_hmaster1 & ~n32812;
  assign n32814 = ~n19800 & ~n32813;
  assign n32815 = ~controllable_hgrant6 & ~n32814;
  assign n32816 = ~n13849 & ~n32815;
  assign n32817 = controllable_hmaster0 & ~n32816;
  assign n32818 = ~n19849 & ~n32817;
  assign n32819 = ~controllable_hmaster3 & ~n32818;
  assign n32820 = ~n30920 & ~n32819;
  assign n32821 = i_hlock7 & ~n32820;
  assign n32822 = ~n23064 & ~n29884;
  assign n32823 = controllable_hmaster1 & ~n32822;
  assign n32824 = ~n19800 & ~n32823;
  assign n32825 = ~controllable_hgrant6 & ~n32824;
  assign n32826 = ~n13951 & ~n32825;
  assign n32827 = controllable_hmaster0 & ~n32826;
  assign n32828 = ~n19849 & ~n32827;
  assign n32829 = ~controllable_hmaster3 & ~n32828;
  assign n32830 = ~n30920 & ~n32829;
  assign n32831 = ~i_hlock7 & ~n32830;
  assign n32832 = ~n32821 & ~n32831;
  assign n32833 = i_hbusreq7 & ~n32832;
  assign n32834 = i_hbusreq8 & ~n32818;
  assign n32835 = i_hbusreq6 & ~n32814;
  assign n32836 = ~n23110 & ~n29947;
  assign n32837 = controllable_hmaster1 & ~n32836;
  assign n32838 = ~n20143 & ~n32837;
  assign n32839 = ~i_hbusreq6 & ~n32838;
  assign n32840 = ~n32835 & ~n32839;
  assign n32841 = ~controllable_hgrant6 & ~n32840;
  assign n32842 = ~n15520 & ~n32841;
  assign n32843 = controllable_hmaster0 & ~n32842;
  assign n32844 = ~n20237 & ~n32843;
  assign n32845 = ~i_hbusreq8 & ~n32844;
  assign n32846 = ~n32834 & ~n32845;
  assign n32847 = ~controllable_hmaster3 & ~n32846;
  assign n32848 = ~n30939 & ~n32847;
  assign n32849 = i_hlock7 & ~n32848;
  assign n32850 = i_hbusreq8 & ~n32828;
  assign n32851 = i_hbusreq6 & ~n32824;
  assign n32852 = ~n23110 & ~n29977;
  assign n32853 = controllable_hmaster1 & ~n32852;
  assign n32854 = ~n20143 & ~n32853;
  assign n32855 = ~i_hbusreq6 & ~n32854;
  assign n32856 = ~n32851 & ~n32855;
  assign n32857 = ~controllable_hgrant6 & ~n32856;
  assign n32858 = ~n15553 & ~n32857;
  assign n32859 = controllable_hmaster0 & ~n32858;
  assign n32860 = ~n20237 & ~n32859;
  assign n32861 = ~i_hbusreq8 & ~n32860;
  assign n32862 = ~n32850 & ~n32861;
  assign n32863 = ~controllable_hmaster3 & ~n32862;
  assign n32864 = ~n30939 & ~n32863;
  assign n32865 = ~i_hlock7 & ~n32864;
  assign n32866 = ~n32849 & ~n32865;
  assign n32867 = ~i_hbusreq7 & ~n32866;
  assign n32868 = ~n32833 & ~n32867;
  assign n32869 = n7924 & ~n32868;
  assign n32870 = ~n32811 & ~n32869;
  assign n32871 = ~n8214 & ~n32870;
  assign n32872 = ~n23158 & ~n29741;
  assign n32873 = ~controllable_hmaster3 & ~n32872;
  assign n32874 = ~n30877 & ~n32873;
  assign n32875 = i_hlock7 & ~n32874;
  assign n32876 = ~n23158 & ~n29756;
  assign n32877 = ~controllable_hmaster3 & ~n32876;
  assign n32878 = ~n30877 & ~n32877;
  assign n32879 = ~i_hlock7 & ~n32878;
  assign n32880 = ~n32875 & ~n32879;
  assign n32881 = i_hbusreq7 & ~n32880;
  assign n32882 = i_hbusreq8 & ~n32872;
  assign n32883 = ~n23184 & ~n29804;
  assign n32884 = ~i_hbusreq8 & ~n32883;
  assign n32885 = ~n32882 & ~n32884;
  assign n32886 = ~controllable_hmaster3 & ~n32885;
  assign n32887 = ~n30896 & ~n32886;
  assign n32888 = i_hlock7 & ~n32887;
  assign n32889 = i_hbusreq8 & ~n32876;
  assign n32890 = ~n23184 & ~n29834;
  assign n32891 = ~i_hbusreq8 & ~n32890;
  assign n32892 = ~n32889 & ~n32891;
  assign n32893 = ~controllable_hmaster3 & ~n32892;
  assign n32894 = ~n30896 & ~n32893;
  assign n32895 = ~i_hlock7 & ~n32894;
  assign n32896 = ~n32888 & ~n32895;
  assign n32897 = ~i_hbusreq7 & ~n32896;
  assign n32898 = ~n32881 & ~n32897;
  assign n32899 = ~n7924 & ~n32898;
  assign n32900 = ~n23223 & ~n29875;
  assign n32901 = ~controllable_hmaster3 & ~n32900;
  assign n32902 = ~n30920 & ~n32901;
  assign n32903 = i_hlock7 & ~n32902;
  assign n32904 = ~n23223 & ~n29890;
  assign n32905 = ~controllable_hmaster3 & ~n32904;
  assign n32906 = ~n30920 & ~n32905;
  assign n32907 = ~i_hlock7 & ~n32906;
  assign n32908 = ~n32903 & ~n32907;
  assign n32909 = i_hbusreq7 & ~n32908;
  assign n32910 = i_hbusreq8 & ~n32900;
  assign n32911 = ~n23274 & ~n29955;
  assign n32912 = ~i_hbusreq8 & ~n32911;
  assign n32913 = ~n32910 & ~n32912;
  assign n32914 = ~controllable_hmaster3 & ~n32913;
  assign n32915 = ~n30939 & ~n32914;
  assign n32916 = i_hlock7 & ~n32915;
  assign n32917 = i_hbusreq8 & ~n32904;
  assign n32918 = ~n23274 & ~n29985;
  assign n32919 = ~i_hbusreq8 & ~n32918;
  assign n32920 = ~n32917 & ~n32919;
  assign n32921 = ~controllable_hmaster3 & ~n32920;
  assign n32922 = ~n30939 & ~n32921;
  assign n32923 = ~i_hlock7 & ~n32922;
  assign n32924 = ~n32916 & ~n32923;
  assign n32925 = ~i_hbusreq7 & ~n32924;
  assign n32926 = ~n32909 & ~n32925;
  assign n32927 = n7924 & ~n32926;
  assign n32928 = ~n32899 & ~n32927;
  assign n32929 = n8214 & ~n32928;
  assign n32930 = ~n32871 & ~n32929;
  assign n32931 = n8202 & ~n32930;
  assign n32932 = ~n32753 & ~n32931;
  assign n32933 = n7920 & ~n32932;
  assign n32934 = ~n10014 & ~n32933;
  assign n32935 = ~n7728 & ~n32934;
  assign n32936 = ~n32591 & ~n32935;
  assign n32937 = n7723 & ~n32936;
  assign n32938 = ~n7723 & ~n32934;
  assign n32939 = ~n32937 & ~n32938;
  assign n32940 = n7714 & ~n32939;
  assign n32941 = n7723 & ~n32934;
  assign n32942 = ~n30295 & ~n31034;
  assign n32943 = ~controllable_hmaster1 & ~n32942;
  assign n32944 = ~n31023 & ~n32943;
  assign n32945 = ~controllable_hgrant6 & ~n32944;
  assign n32946 = ~n13849 & ~n32945;
  assign n32947 = controllable_hmaster0 & ~n32946;
  assign n32948 = ~n31074 & ~n32947;
  assign n32949 = ~controllable_hmaster3 & ~n32948;
  assign n32950 = ~n31871 & ~n32949;
  assign n32951 = i_hlock7 & ~n32950;
  assign n32952 = ~n30398 & ~n31141;
  assign n32953 = ~controllable_hmaster1 & ~n32952;
  assign n32954 = ~n31130 & ~n32953;
  assign n32955 = ~controllable_hgrant6 & ~n32954;
  assign n32956 = ~n13951 & ~n32955;
  assign n32957 = controllable_hmaster0 & ~n32956;
  assign n32958 = ~n31181 & ~n32957;
  assign n32959 = ~controllable_hmaster3 & ~n32958;
  assign n32960 = ~n31893 & ~n32959;
  assign n32961 = ~i_hlock7 & ~n32960;
  assign n32962 = ~n32951 & ~n32961;
  assign n32963 = i_hbusreq7 & ~n32962;
  assign n32964 = i_hbusreq8 & ~n32948;
  assign n32965 = i_hbusreq6 & ~n32944;
  assign n32966 = i_hlock5 & ~n31738;
  assign n32967 = ~i_hlock5 & ~n31760;
  assign n32968 = ~n32966 & ~n32967;
  assign n32969 = ~i_hbusreq5 & ~n32968;
  assign n32970 = ~n30560 & ~n32969;
  assign n32971 = ~controllable_hgrant5 & ~n32970;
  assign n32972 = ~n15020 & ~n32971;
  assign n32973 = controllable_hmaster2 & ~n32972;
  assign n32974 = ~n31334 & ~n32973;
  assign n32975 = ~controllable_hmaster1 & ~n32974;
  assign n32976 = ~n31311 & ~n32975;
  assign n32977 = ~i_hbusreq6 & ~n32976;
  assign n32978 = ~n32965 & ~n32977;
  assign n32979 = ~controllable_hgrant6 & ~n32978;
  assign n32980 = ~n15417 & ~n32979;
  assign n32981 = controllable_hmaster0 & ~n32980;
  assign n32982 = ~n31403 & ~n32981;
  assign n32983 = ~i_hbusreq8 & ~n32982;
  assign n32984 = ~n32964 & ~n32983;
  assign n32985 = ~controllable_hmaster3 & ~n32984;
  assign n32986 = ~n31920 & ~n32985;
  assign n32987 = i_hlock7 & ~n32986;
  assign n32988 = i_hbusreq8 & ~n32958;
  assign n32989 = i_hbusreq6 & ~n32954;
  assign n32990 = i_hlock5 & ~n31814;
  assign n32991 = ~i_hlock5 & ~n31836;
  assign n32992 = ~n32990 & ~n32991;
  assign n32993 = ~i_hbusreq5 & ~n32992;
  assign n32994 = ~n30768 & ~n32993;
  assign n32995 = ~controllable_hgrant5 & ~n32994;
  assign n32996 = ~n15020 & ~n32995;
  assign n32997 = controllable_hmaster2 & ~n32996;
  assign n32998 = ~n31556 & ~n32997;
  assign n32999 = ~controllable_hmaster1 & ~n32998;
  assign n33000 = ~n31533 & ~n32999;
  assign n33001 = ~i_hbusreq6 & ~n33000;
  assign n33002 = ~n32989 & ~n33001;
  assign n33003 = ~controllable_hgrant6 & ~n33002;
  assign n33004 = ~n15440 & ~n33003;
  assign n33005 = controllable_hmaster0 & ~n33004;
  assign n33006 = ~n31625 & ~n33005;
  assign n33007 = ~i_hbusreq8 & ~n33006;
  assign n33008 = ~n32988 & ~n33007;
  assign n33009 = ~controllable_hmaster3 & ~n33008;
  assign n33010 = ~n31953 & ~n33009;
  assign n33011 = ~i_hlock7 & ~n33010;
  assign n33012 = ~n32987 & ~n33011;
  assign n33013 = ~i_hbusreq7 & ~n33012;
  assign n33014 = ~n32963 & ~n33013;
  assign n33015 = n7924 & ~n33014;
  assign n33016 = ~n32641 & ~n33015;
  assign n33017 = ~n8214 & ~n33016;
  assign n33018 = ~n30322 & ~n31061;
  assign n33019 = ~controllable_hmaster1 & ~n33018;
  assign n33020 = ~n31048 & ~n33019;
  assign n33021 = i_hlock6 & ~n33020;
  assign n33022 = ~n31068 & ~n33019;
  assign n33023 = ~i_hlock6 & ~n33022;
  assign n33024 = ~n33021 & ~n33023;
  assign n33025 = ~controllable_hgrant6 & ~n33024;
  assign n33026 = ~n13894 & ~n33025;
  assign n33027 = ~controllable_hmaster0 & ~n33026;
  assign n33028 = ~n31040 & ~n33027;
  assign n33029 = ~controllable_hmaster3 & ~n33028;
  assign n33030 = ~n31871 & ~n33029;
  assign n33031 = i_hlock7 & ~n33030;
  assign n33032 = ~n30425 & ~n31168;
  assign n33033 = ~controllable_hmaster1 & ~n33032;
  assign n33034 = ~n31155 & ~n33033;
  assign n33035 = i_hlock6 & ~n33034;
  assign n33036 = ~n31175 & ~n33033;
  assign n33037 = ~i_hlock6 & ~n33036;
  assign n33038 = ~n33035 & ~n33037;
  assign n33039 = ~controllable_hgrant6 & ~n33038;
  assign n33040 = ~n13894 & ~n33039;
  assign n33041 = ~controllable_hmaster0 & ~n33040;
  assign n33042 = ~n31147 & ~n33041;
  assign n33043 = ~controllable_hmaster3 & ~n33042;
  assign n33044 = ~n31893 & ~n33043;
  assign n33045 = ~i_hlock7 & ~n33044;
  assign n33046 = ~n33031 & ~n33045;
  assign n33047 = i_hbusreq7 & ~n33046;
  assign n33048 = i_hbusreq8 & ~n33028;
  assign n33049 = i_hbusreq6 & ~n33024;
  assign n33050 = i_hlock4 & ~n31734;
  assign n33051 = ~i_hlock4 & ~n31756;
  assign n33052 = ~n33050 & ~n33051;
  assign n33053 = ~i_hbusreq4 & ~n33052;
  assign n33054 = ~n30610 & ~n33053;
  assign n33055 = ~controllable_hgrant4 & ~n33054;
  assign n33056 = ~n15091 & ~n33055;
  assign n33057 = ~i_hbusreq5 & ~n33056;
  assign n33058 = ~n30609 & ~n33057;
  assign n33059 = ~controllable_hgrant5 & ~n33058;
  assign n33060 = ~n15090 & ~n33059;
  assign n33061 = controllable_hmaster2 & ~n33060;
  assign n33062 = ~n31388 & ~n33061;
  assign n33063 = ~controllable_hmaster1 & ~n33062;
  assign n33064 = ~n31360 & ~n33063;
  assign n33065 = i_hlock6 & ~n33064;
  assign n33066 = ~n31395 & ~n33063;
  assign n33067 = ~i_hlock6 & ~n33066;
  assign n33068 = ~n33065 & ~n33067;
  assign n33069 = ~i_hbusreq6 & ~n33068;
  assign n33070 = ~n33049 & ~n33069;
  assign n33071 = ~controllable_hgrant6 & ~n33070;
  assign n33072 = ~n15467 & ~n33071;
  assign n33073 = ~controllable_hmaster0 & ~n33072;
  assign n33074 = ~n31342 & ~n33073;
  assign n33075 = ~i_hbusreq8 & ~n33074;
  assign n33076 = ~n33048 & ~n33075;
  assign n33077 = ~controllable_hmaster3 & ~n33076;
  assign n33078 = ~n31920 & ~n33077;
  assign n33079 = i_hlock7 & ~n33078;
  assign n33080 = i_hbusreq8 & ~n33042;
  assign n33081 = i_hbusreq6 & ~n33038;
  assign n33082 = i_hlock4 & ~n31810;
  assign n33083 = ~i_hlock4 & ~n31832;
  assign n33084 = ~n33082 & ~n33083;
  assign n33085 = ~i_hbusreq4 & ~n33084;
  assign n33086 = ~n30818 & ~n33085;
  assign n33087 = ~controllable_hgrant4 & ~n33086;
  assign n33088 = ~n15091 & ~n33087;
  assign n33089 = ~i_hbusreq5 & ~n33088;
  assign n33090 = ~n30817 & ~n33089;
  assign n33091 = ~controllable_hgrant5 & ~n33090;
  assign n33092 = ~n15090 & ~n33091;
  assign n33093 = controllable_hmaster2 & ~n33092;
  assign n33094 = ~n31610 & ~n33093;
  assign n33095 = ~controllable_hmaster1 & ~n33094;
  assign n33096 = ~n31582 & ~n33095;
  assign n33097 = i_hlock6 & ~n33096;
  assign n33098 = ~n31617 & ~n33095;
  assign n33099 = ~i_hlock6 & ~n33098;
  assign n33100 = ~n33097 & ~n33099;
  assign n33101 = ~i_hbusreq6 & ~n33100;
  assign n33102 = ~n33081 & ~n33101;
  assign n33103 = ~controllable_hgrant6 & ~n33102;
  assign n33104 = ~n15467 & ~n33103;
  assign n33105 = ~controllable_hmaster0 & ~n33104;
  assign n33106 = ~n31564 & ~n33105;
  assign n33107 = ~i_hbusreq8 & ~n33106;
  assign n33108 = ~n33080 & ~n33107;
  assign n33109 = ~controllable_hmaster3 & ~n33108;
  assign n33110 = ~n31953 & ~n33109;
  assign n33111 = ~i_hlock7 & ~n33110;
  assign n33112 = ~n33079 & ~n33111;
  assign n33113 = ~i_hbusreq7 & ~n33112;
  assign n33114 = ~n33047 & ~n33113;
  assign n33115 = n7924 & ~n33114;
  assign n33116 = ~n32721 & ~n33115;
  assign n33117 = n8214 & ~n33116;
  assign n33118 = ~n33017 & ~n33117;
  assign n33119 = ~n8202 & ~n33118;
  assign n33120 = ~n30287 & ~n31016;
  assign n33121 = controllable_hmaster1 & ~n33120;
  assign n33122 = ~n31036 & ~n33121;
  assign n33123 = ~controllable_hgrant6 & ~n33122;
  assign n33124 = ~n13849 & ~n33123;
  assign n33125 = controllable_hmaster0 & ~n33124;
  assign n33126 = ~n31074 & ~n33125;
  assign n33127 = ~controllable_hmaster3 & ~n33126;
  assign n33128 = ~n31871 & ~n33127;
  assign n33129 = i_hlock7 & ~n33128;
  assign n33130 = ~n30390 & ~n31123;
  assign n33131 = controllable_hmaster1 & ~n33130;
  assign n33132 = ~n31143 & ~n33131;
  assign n33133 = ~controllable_hgrant6 & ~n33132;
  assign n33134 = ~n13951 & ~n33133;
  assign n33135 = controllable_hmaster0 & ~n33134;
  assign n33136 = ~n31181 & ~n33135;
  assign n33137 = ~controllable_hmaster3 & ~n33136;
  assign n33138 = ~n31893 & ~n33137;
  assign n33139 = ~i_hlock7 & ~n33138;
  assign n33140 = ~n33129 & ~n33139;
  assign n33141 = i_hbusreq7 & ~n33140;
  assign n33142 = i_hbusreq8 & ~n33126;
  assign n33143 = i_hbusreq6 & ~n33122;
  assign n33144 = ~i_hbusreq9 & ~n23467;
  assign n33145 = ~n30546 & ~n33144;
  assign n33146 = ~i_hbusreq4 & ~n33145;
  assign n33147 = ~n30545 & ~n33146;
  assign n33148 = ~controllable_hgrant4 & ~n33147;
  assign n33149 = ~n14998 & ~n33148;
  assign n33150 = ~i_hbusreq5 & ~n33149;
  assign n33151 = ~n30544 & ~n33150;
  assign n33152 = ~controllable_hgrant5 & ~n33151;
  assign n33153 = ~n14997 & ~n33152;
  assign n33154 = ~controllable_hmaster2 & ~n33153;
  assign n33155 = ~n31295 & ~n33154;
  assign n33156 = controllable_hmaster1 & ~n33155;
  assign n33157 = ~n31336 & ~n33156;
  assign n33158 = ~i_hbusreq6 & ~n33157;
  assign n33159 = ~n33143 & ~n33158;
  assign n33160 = ~controllable_hgrant6 & ~n33159;
  assign n33161 = ~n15520 & ~n33160;
  assign n33162 = controllable_hmaster0 & ~n33161;
  assign n33163 = ~n31403 & ~n33162;
  assign n33164 = ~i_hbusreq8 & ~n33163;
  assign n33165 = ~n33142 & ~n33164;
  assign n33166 = ~controllable_hmaster3 & ~n33165;
  assign n33167 = ~n31920 & ~n33166;
  assign n33168 = i_hlock7 & ~n33167;
  assign n33169 = i_hbusreq8 & ~n33136;
  assign n33170 = i_hbusreq6 & ~n33132;
  assign n33171 = ~i_hbusreq9 & ~n23475;
  assign n33172 = ~n30754 & ~n33171;
  assign n33173 = ~i_hbusreq4 & ~n33172;
  assign n33174 = ~n30753 & ~n33173;
  assign n33175 = ~controllable_hgrant4 & ~n33174;
  assign n33176 = ~n14998 & ~n33175;
  assign n33177 = ~i_hbusreq5 & ~n33176;
  assign n33178 = ~n30752 & ~n33177;
  assign n33179 = ~controllable_hgrant5 & ~n33178;
  assign n33180 = ~n14997 & ~n33179;
  assign n33181 = ~controllable_hmaster2 & ~n33180;
  assign n33182 = ~n31517 & ~n33181;
  assign n33183 = controllable_hmaster1 & ~n33182;
  assign n33184 = ~n31558 & ~n33183;
  assign n33185 = ~i_hbusreq6 & ~n33184;
  assign n33186 = ~n33170 & ~n33185;
  assign n33187 = ~controllable_hgrant6 & ~n33186;
  assign n33188 = ~n15553 & ~n33187;
  assign n33189 = controllable_hmaster0 & ~n33188;
  assign n33190 = ~n31625 & ~n33189;
  assign n33191 = ~i_hbusreq8 & ~n33190;
  assign n33192 = ~n33169 & ~n33191;
  assign n33193 = ~controllable_hmaster3 & ~n33192;
  assign n33194 = ~n31953 & ~n33193;
  assign n33195 = ~i_hlock7 & ~n33194;
  assign n33196 = ~n33168 & ~n33195;
  assign n33197 = ~i_hbusreq7 & ~n33196;
  assign n33198 = ~n33141 & ~n33197;
  assign n33199 = n7924 & ~n33198;
  assign n33200 = ~n32811 & ~n33199;
  assign n33201 = ~n8214 & ~n33200;
  assign n33202 = ~n30312 & ~n31041;
  assign n33203 = controllable_hmaster1 & ~n33202;
  assign n33204 = ~n31063 & ~n33203;
  assign n33205 = i_hlock6 & ~n33204;
  assign n33206 = ~n30312 & ~n31066;
  assign n33207 = controllable_hmaster1 & ~n33206;
  assign n33208 = ~n31063 & ~n33207;
  assign n33209 = ~i_hlock6 & ~n33208;
  assign n33210 = ~n33205 & ~n33209;
  assign n33211 = ~controllable_hgrant6 & ~n33210;
  assign n33212 = ~n13894 & ~n33211;
  assign n33213 = ~controllable_hmaster0 & ~n33212;
  assign n33214 = ~n31040 & ~n33213;
  assign n33215 = ~controllable_hmaster3 & ~n33214;
  assign n33216 = ~n31871 & ~n33215;
  assign n33217 = i_hlock7 & ~n33216;
  assign n33218 = ~n30415 & ~n31148;
  assign n33219 = controllable_hmaster1 & ~n33218;
  assign n33220 = ~n31170 & ~n33219;
  assign n33221 = i_hlock6 & ~n33220;
  assign n33222 = ~n30415 & ~n31173;
  assign n33223 = controllable_hmaster1 & ~n33222;
  assign n33224 = ~n31170 & ~n33223;
  assign n33225 = ~i_hlock6 & ~n33224;
  assign n33226 = ~n33221 & ~n33225;
  assign n33227 = ~controllable_hgrant6 & ~n33226;
  assign n33228 = ~n13894 & ~n33227;
  assign n33229 = ~controllable_hmaster0 & ~n33228;
  assign n33230 = ~n31147 & ~n33229;
  assign n33231 = ~controllable_hmaster3 & ~n33230;
  assign n33232 = ~n31893 & ~n33231;
  assign n33233 = ~i_hlock7 & ~n33232;
  assign n33234 = ~n33217 & ~n33233;
  assign n33235 = i_hbusreq7 & ~n33234;
  assign n33236 = i_hbusreq8 & ~n33214;
  assign n33237 = i_hbusreq6 & ~n33210;
  assign n33238 = ~i_hbusreq9 & ~n23557;
  assign n33239 = ~n30595 & ~n33238;
  assign n33240 = ~i_hbusreq4 & ~n33239;
  assign n33241 = ~n30594 & ~n33240;
  assign n33242 = ~controllable_hgrant4 & ~n33241;
  assign n33243 = ~n15065 & ~n33242;
  assign n33244 = ~i_hbusreq5 & ~n33243;
  assign n33245 = ~n30593 & ~n33244;
  assign n33246 = ~controllable_hgrant5 & ~n33245;
  assign n33247 = ~n15064 & ~n33246;
  assign n33248 = ~controllable_hmaster2 & ~n33247;
  assign n33249 = ~n31344 & ~n33248;
  assign n33250 = controllable_hmaster1 & ~n33249;
  assign n33251 = ~n31390 & ~n33250;
  assign n33252 = i_hlock6 & ~n33251;
  assign n33253 = ~n31393 & ~n33248;
  assign n33254 = controllable_hmaster1 & ~n33253;
  assign n33255 = ~n31390 & ~n33254;
  assign n33256 = ~i_hlock6 & ~n33255;
  assign n33257 = ~n33252 & ~n33256;
  assign n33258 = ~i_hbusreq6 & ~n33257;
  assign n33259 = ~n33237 & ~n33258;
  assign n33260 = ~controllable_hgrant6 & ~n33259;
  assign n33261 = ~n15582 & ~n33260;
  assign n33262 = ~controllable_hmaster0 & ~n33261;
  assign n33263 = ~n31342 & ~n33262;
  assign n33264 = ~i_hbusreq8 & ~n33263;
  assign n33265 = ~n33236 & ~n33264;
  assign n33266 = ~controllable_hmaster3 & ~n33265;
  assign n33267 = ~n31920 & ~n33266;
  assign n33268 = i_hlock7 & ~n33267;
  assign n33269 = i_hbusreq8 & ~n33230;
  assign n33270 = i_hbusreq6 & ~n33226;
  assign n33271 = ~i_hbusreq9 & ~n23567;
  assign n33272 = ~n30803 & ~n33271;
  assign n33273 = ~i_hbusreq4 & ~n33272;
  assign n33274 = ~n30802 & ~n33273;
  assign n33275 = ~controllable_hgrant4 & ~n33274;
  assign n33276 = ~n15065 & ~n33275;
  assign n33277 = ~i_hbusreq5 & ~n33276;
  assign n33278 = ~n30801 & ~n33277;
  assign n33279 = ~controllable_hgrant5 & ~n33278;
  assign n33280 = ~n15064 & ~n33279;
  assign n33281 = ~controllable_hmaster2 & ~n33280;
  assign n33282 = ~n31566 & ~n33281;
  assign n33283 = controllable_hmaster1 & ~n33282;
  assign n33284 = ~n31612 & ~n33283;
  assign n33285 = i_hlock6 & ~n33284;
  assign n33286 = ~n31615 & ~n33281;
  assign n33287 = controllable_hmaster1 & ~n33286;
  assign n33288 = ~n31612 & ~n33287;
  assign n33289 = ~i_hlock6 & ~n33288;
  assign n33290 = ~n33285 & ~n33289;
  assign n33291 = ~i_hbusreq6 & ~n33290;
  assign n33292 = ~n33270 & ~n33291;
  assign n33293 = ~controllable_hgrant6 & ~n33292;
  assign n33294 = ~n15582 & ~n33293;
  assign n33295 = ~controllable_hmaster0 & ~n33294;
  assign n33296 = ~n31564 & ~n33295;
  assign n33297 = ~i_hbusreq8 & ~n33296;
  assign n33298 = ~n33269 & ~n33297;
  assign n33299 = ~controllable_hmaster3 & ~n33298;
  assign n33300 = ~n31953 & ~n33299;
  assign n33301 = ~i_hlock7 & ~n33300;
  assign n33302 = ~n33268 & ~n33301;
  assign n33303 = ~i_hbusreq7 & ~n33302;
  assign n33304 = ~n33235 & ~n33303;
  assign n33305 = n7924 & ~n33304;
  assign n33306 = ~n32899 & ~n33305;
  assign n33307 = n8214 & ~n33306;
  assign n33308 = ~n33201 & ~n33307;
  assign n33309 = n8202 & ~n33308;
  assign n33310 = ~n33119 & ~n33309;
  assign n33311 = n7920 & ~n33310;
  assign n33312 = ~n28799 & ~n33311;
  assign n33313 = n7728 & ~n33312;
  assign n33314 = ~n32399 & ~n33313;
  assign n33315 = ~n7723 & ~n33314;
  assign n33316 = ~n32941 & ~n33315;
  assign n33317 = ~n7714 & ~n33316;
  assign n33318 = ~n32940 & ~n33317;
  assign n33319 = ~n7705 & ~n33318;
  assign n33320 = ~n22399 & ~n33319;
  assign n33321 = n7808 & ~n33320;
  assign n33322 = ~n32419 & ~n33321;
  assign n33323 = ~n8195 & ~n33322;
  assign n33324 = controllable_hgrant6 & ~n11963;
  assign n33325 = controllable_hgrant5 & ~n10380;
  assign n33326 = controllable_hgrant4 & ~n10380;
  assign n33327 = ~controllable_hgrant4 & ~n23639;
  assign n33328 = ~n33326 & ~n33327;
  assign n33329 = ~controllable_hgrant5 & ~n33328;
  assign n33330 = ~n33325 & ~n33329;
  assign n33331 = controllable_hmaster2 & ~n33330;
  assign n33332 = ~n10389 & ~n33331;
  assign n33333 = controllable_hmaster1 & ~n33332;
  assign n33334 = ~n10409 & ~n33333;
  assign n33335 = ~controllable_hgrant6 & ~n33334;
  assign n33336 = ~n33324 & ~n33335;
  assign n33337 = controllable_hmaster0 & ~n33336;
  assign n33338 = ~n10445 & ~n33337;
  assign n33339 = ~controllable_hmaster3 & ~n33338;
  assign n33340 = ~n10379 & ~n33339;
  assign n33341 = i_hlock7 & ~n33340;
  assign n33342 = controllable_hgrant6 & ~n11971;
  assign n33343 = controllable_hgrant5 & ~n10384;
  assign n33344 = controllable_hgrant4 & ~n10384;
  assign n33345 = ~controllable_hgrant4 & ~n23647;
  assign n33346 = ~n33344 & ~n33345;
  assign n33347 = ~controllable_hgrant5 & ~n33346;
  assign n33348 = ~n33343 & ~n33347;
  assign n33349 = controllable_hmaster2 & ~n33348;
  assign n33350 = ~n10389 & ~n33349;
  assign n33351 = controllable_hmaster1 & ~n33350;
  assign n33352 = ~n10409 & ~n33351;
  assign n33353 = ~controllable_hgrant6 & ~n33352;
  assign n33354 = ~n33342 & ~n33353;
  assign n33355 = controllable_hmaster0 & ~n33354;
  assign n33356 = ~n10445 & ~n33355;
  assign n33357 = ~controllable_hmaster3 & ~n33356;
  assign n33358 = ~n10379 & ~n33357;
  assign n33359 = ~i_hlock7 & ~n33358;
  assign n33360 = ~n33341 & ~n33359;
  assign n33361 = i_hbusreq7 & ~n33360;
  assign n33362 = i_hbusreq8 & ~n33338;
  assign n33363 = controllable_hgrant6 & ~n11985;
  assign n33364 = i_hbusreq6 & ~n33334;
  assign n33365 = controllable_hgrant5 & ~n10596;
  assign n33366 = i_hbusreq5 & ~n33328;
  assign n33367 = controllable_hgrant4 & ~n10501;
  assign n33368 = i_hbusreq4 & ~n23639;
  assign n33369 = i_hbusreq9 & ~n23639;
  assign n33370 = ~i_hbusreq9 & ~n23685;
  assign n33371 = ~n33369 & ~n33370;
  assign n33372 = ~i_hbusreq4 & ~n33371;
  assign n33373 = ~n33368 & ~n33372;
  assign n33374 = ~controllable_hgrant4 & ~n33373;
  assign n33375 = ~n33367 & ~n33374;
  assign n33376 = ~i_hbusreq5 & ~n33375;
  assign n33377 = ~n33366 & ~n33376;
  assign n33378 = ~controllable_hgrant5 & ~n33377;
  assign n33379 = ~n33365 & ~n33378;
  assign n33380 = controllable_hmaster2 & ~n33379;
  assign n33381 = ~n10489 & ~n33380;
  assign n33382 = controllable_hmaster1 & ~n33381;
  assign n33383 = ~n10545 & ~n33382;
  assign n33384 = ~i_hbusreq6 & ~n33383;
  assign n33385 = ~n33364 & ~n33384;
  assign n33386 = ~controllable_hgrant6 & ~n33385;
  assign n33387 = ~n33363 & ~n33386;
  assign n33388 = controllable_hmaster0 & ~n33387;
  assign n33389 = ~n10617 & ~n33388;
  assign n33390 = ~i_hbusreq8 & ~n33389;
  assign n33391 = ~n33362 & ~n33390;
  assign n33392 = ~controllable_hmaster3 & ~n33391;
  assign n33393 = ~n10459 & ~n33392;
  assign n33394 = i_hlock7 & ~n33393;
  assign n33395 = i_hbusreq8 & ~n33356;
  assign n33396 = controllable_hgrant6 & ~n11999;
  assign n33397 = i_hbusreq6 & ~n33352;
  assign n33398 = controllable_hgrant5 & ~n10606;
  assign n33399 = i_hbusreq5 & ~n33346;
  assign n33400 = controllable_hgrant4 & ~n10513;
  assign n33401 = i_hbusreq4 & ~n23647;
  assign n33402 = i_hbusreq9 & ~n23647;
  assign n33403 = ~i_hbusreq9 & ~n23699;
  assign n33404 = ~n33402 & ~n33403;
  assign n33405 = ~i_hbusreq4 & ~n33404;
  assign n33406 = ~n33401 & ~n33405;
  assign n33407 = ~controllable_hgrant4 & ~n33406;
  assign n33408 = ~n33400 & ~n33407;
  assign n33409 = ~i_hbusreq5 & ~n33408;
  assign n33410 = ~n33399 & ~n33409;
  assign n33411 = ~controllable_hgrant5 & ~n33410;
  assign n33412 = ~n33398 & ~n33411;
  assign n33413 = controllable_hmaster2 & ~n33412;
  assign n33414 = ~n10489 & ~n33413;
  assign n33415 = controllable_hmaster1 & ~n33414;
  assign n33416 = ~n10545 & ~n33415;
  assign n33417 = ~i_hbusreq6 & ~n33416;
  assign n33418 = ~n33397 & ~n33417;
  assign n33419 = ~controllable_hgrant6 & ~n33418;
  assign n33420 = ~n33396 & ~n33419;
  assign n33421 = controllable_hmaster0 & ~n33420;
  assign n33422 = ~n10617 & ~n33421;
  assign n33423 = ~i_hbusreq8 & ~n33422;
  assign n33424 = ~n33395 & ~n33423;
  assign n33425 = ~controllable_hmaster3 & ~n33424;
  assign n33426 = ~n10459 & ~n33425;
  assign n33427 = ~i_hlock7 & ~n33426;
  assign n33428 = ~n33394 & ~n33427;
  assign n33429 = ~i_hbusreq7 & ~n33428;
  assign n33430 = ~n33361 & ~n33429;
  assign n33431 = n7924 & ~n33430;
  assign n33432 = ~n10375 & ~n33431;
  assign n33433 = n8214 & ~n33432;
  assign n33434 = n8214 & ~n33433;
  assign n33435 = n8202 & ~n33434;
  assign n33436 = ~n10332 & ~n33435;
  assign n33437 = n7728 & ~n33436;
  assign n33438 = n8214 & ~n28798;
  assign n33439 = ~n8336 & ~n33438;
  assign n33440 = n8202 & ~n33439;
  assign n33441 = ~n10649 & ~n33440;
  assign n33442 = ~n7728 & ~n33441;
  assign n33443 = ~n33437 & ~n33442;
  assign n33444 = ~n7723 & ~n33443;
  assign n33445 = ~n7723 & ~n33444;
  assign n33446 = ~n7714 & ~n33445;
  assign n33447 = ~n7714 & ~n33446;
  assign n33448 = n7705 & ~n33447;
  assign n33449 = n7723 & ~n33441;
  assign n33450 = n7920 & ~n33441;
  assign n33451 = ~n28799 & ~n33450;
  assign n33452 = ~n7723 & ~n33451;
  assign n33453 = ~n33449 & ~n33452;
  assign n33454 = n7714 & ~n33453;
  assign n33455 = ~n28805 & ~n33454;
  assign n33456 = ~n7705 & ~n33455;
  assign n33457 = ~n33448 & ~n33456;
  assign n33458 = ~n7808 & ~n33457;
  assign n33459 = ~n7920 & ~n33436;
  assign n33460 = n7924 & ~n32395;
  assign n33461 = ~n8214 & ~n33460;
  assign n33462 = controllable_hmaster3 & ~n23853;
  assign n33463 = controllable_hmaster2 & ~n23841;
  assign n33464 = ~n17340 & ~n33463;
  assign n33465 = controllable_hmaster1 & ~n33464;
  assign n33466 = ~n29423 & ~n33465;
  assign n33467 = ~controllable_hgrant6 & ~n33466;
  assign n33468 = ~n13198 & ~n33467;
  assign n33469 = controllable_hmaster0 & ~n33468;
  assign n33470 = ~n29428 & ~n33469;
  assign n33471 = ~controllable_hmaster3 & ~n33470;
  assign n33472 = ~n33462 & ~n33471;
  assign n33473 = i_hbusreq7 & ~n33472;
  assign n33474 = i_hbusreq8 & ~n23853;
  assign n33475 = ~i_hbusreq8 & ~n23948;
  assign n33476 = ~n33474 & ~n33475;
  assign n33477 = controllable_hmaster3 & ~n33476;
  assign n33478 = i_hbusreq8 & ~n33470;
  assign n33479 = i_hbusreq6 & ~n33466;
  assign n33480 = controllable_hmaster2 & ~n23911;
  assign n33481 = ~n23941 & ~n33480;
  assign n33482 = controllable_hmaster1 & ~n33481;
  assign n33483 = ~controllable_hmaster1 & ~n23940;
  assign n33484 = ~n33482 & ~n33483;
  assign n33485 = ~i_hbusreq6 & ~n33484;
  assign n33486 = ~n33479 & ~n33485;
  assign n33487 = ~controllable_hgrant6 & ~n33486;
  assign n33488 = ~n15812 & ~n33487;
  assign n33489 = controllable_hmaster0 & ~n33488;
  assign n33490 = ~n23988 & ~n33489;
  assign n33491 = ~i_hbusreq8 & ~n33490;
  assign n33492 = ~n33478 & ~n33491;
  assign n33493 = ~controllable_hmaster3 & ~n33492;
  assign n33494 = ~n33477 & ~n33493;
  assign n33495 = ~i_hbusreq7 & ~n33494;
  assign n33496 = ~n33473 & ~n33495;
  assign n33497 = ~n7924 & ~n33496;
  assign n33498 = ~controllable_hgrant4 & ~n24001;
  assign n33499 = ~n13177 & ~n33498;
  assign n33500 = ~controllable_hgrant5 & ~n33499;
  assign n33501 = ~n13176 & ~n33500;
  assign n33502 = controllable_hmaster1 & ~n33501;
  assign n33503 = controllable_hmaster2 & ~n33501;
  assign n33504 = ~n29497 & ~n33503;
  assign n33505 = ~controllable_hmaster1 & ~n33504;
  assign n33506 = ~n33502 & ~n33505;
  assign n33507 = ~controllable_hgrant6 & ~n33506;
  assign n33508 = ~n13198 & ~n33507;
  assign n33509 = controllable_hmaster3 & ~n33508;
  assign n33510 = ~controllable_hgrant4 & ~n24020;
  assign n33511 = ~n13177 & ~n33510;
  assign n33512 = ~controllable_hgrant5 & ~n33511;
  assign n33513 = ~n13176 & ~n33512;
  assign n33514 = controllable_hmaster2 & ~n33513;
  assign n33515 = ~n29497 & ~n33514;
  assign n33516 = controllable_hmaster1 & ~n33515;
  assign n33517 = ~n29506 & ~n33516;
  assign n33518 = ~controllable_hgrant6 & ~n33517;
  assign n33519 = ~n13198 & ~n33518;
  assign n33520 = controllable_hmaster0 & ~n33519;
  assign n33521 = ~n29513 & ~n33520;
  assign n33522 = ~controllable_hmaster3 & ~n33521;
  assign n33523 = ~n33509 & ~n33522;
  assign n33524 = i_hlock7 & ~n33523;
  assign n33525 = ~controllable_hgrant4 & ~n24007;
  assign n33526 = ~n13177 & ~n33525;
  assign n33527 = ~controllable_hgrant5 & ~n33526;
  assign n33528 = ~n13176 & ~n33527;
  assign n33529 = controllable_hmaster1 & ~n33528;
  assign n33530 = controllable_hmaster2 & ~n33528;
  assign n33531 = ~n29528 & ~n33530;
  assign n33532 = ~controllable_hmaster1 & ~n33531;
  assign n33533 = ~n33529 & ~n33532;
  assign n33534 = ~controllable_hgrant6 & ~n33533;
  assign n33535 = ~n13198 & ~n33534;
  assign n33536 = controllable_hmaster3 & ~n33535;
  assign n33537 = ~controllable_hgrant4 & ~n24026;
  assign n33538 = ~n13177 & ~n33537;
  assign n33539 = ~controllable_hgrant5 & ~n33538;
  assign n33540 = ~n13176 & ~n33539;
  assign n33541 = controllable_hmaster2 & ~n33540;
  assign n33542 = ~n29528 & ~n33541;
  assign n33543 = controllable_hmaster1 & ~n33542;
  assign n33544 = ~n29537 & ~n33543;
  assign n33545 = ~controllable_hgrant6 & ~n33544;
  assign n33546 = ~n13198 & ~n33545;
  assign n33547 = controllable_hmaster0 & ~n33546;
  assign n33548 = ~n29544 & ~n33547;
  assign n33549 = ~controllable_hmaster3 & ~n33548;
  assign n33550 = ~n33536 & ~n33549;
  assign n33551 = ~i_hlock7 & ~n33550;
  assign n33552 = ~n33524 & ~n33551;
  assign n33553 = i_hbusreq7 & ~n33552;
  assign n33554 = i_hbusreq8 & ~n33508;
  assign n33555 = i_hbusreq6 & ~n33506;
  assign n33556 = i_hbusreq5 & ~n33499;
  assign n33557 = i_hbusreq4 & ~n24001;
  assign n33558 = i_hbusreq9 & ~n24001;
  assign n33559 = ~i_hbusreq9 & ~n24065;
  assign n33560 = ~n33558 & ~n33559;
  assign n33561 = ~i_hbusreq4 & ~n33560;
  assign n33562 = ~n33557 & ~n33561;
  assign n33563 = ~controllable_hgrant4 & ~n33562;
  assign n33564 = ~n15728 & ~n33563;
  assign n33565 = ~i_hbusreq5 & ~n33564;
  assign n33566 = ~n33556 & ~n33565;
  assign n33567 = ~controllable_hgrant5 & ~n33566;
  assign n33568 = ~n15727 & ~n33567;
  assign n33569 = controllable_hmaster1 & ~n33568;
  assign n33570 = controllable_hmaster2 & ~n33568;
  assign n33571 = ~i_hbusreq9 & ~n24148;
  assign n33572 = ~n29570 & ~n33571;
  assign n33573 = ~i_hbusreq4 & ~n33572;
  assign n33574 = ~n29569 & ~n33573;
  assign n33575 = ~controllable_hgrant4 & ~n33574;
  assign n33576 = ~n15675 & ~n33575;
  assign n33577 = ~i_hbusreq5 & ~n33576;
  assign n33578 = ~n29568 & ~n33577;
  assign n33579 = ~controllable_hgrant5 & ~n33578;
  assign n33580 = ~n15674 & ~n33579;
  assign n33581 = ~controllable_hmaster2 & ~n33580;
  assign n33582 = ~n33570 & ~n33581;
  assign n33583 = ~controllable_hmaster1 & ~n33582;
  assign n33584 = ~n33569 & ~n33583;
  assign n33585 = ~i_hbusreq6 & ~n33584;
  assign n33586 = ~n33555 & ~n33585;
  assign n33587 = ~controllable_hgrant6 & ~n33586;
  assign n33588 = ~n15672 & ~n33587;
  assign n33589 = ~i_hbusreq8 & ~n33588;
  assign n33590 = ~n33554 & ~n33589;
  assign n33591 = controllable_hmaster3 & ~n33590;
  assign n33592 = i_hbusreq8 & ~n33521;
  assign n33593 = i_hbusreq6 & ~n33517;
  assign n33594 = i_hbusreq5 & ~n33511;
  assign n33595 = i_hbusreq4 & ~n24020;
  assign n33596 = i_hbusreq9 & ~n24020;
  assign n33597 = ~i_hbusreq9 & ~n24105;
  assign n33598 = ~n33596 & ~n33597;
  assign n33599 = ~i_hbusreq4 & ~n33598;
  assign n33600 = ~n33595 & ~n33599;
  assign n33601 = ~controllable_hgrant4 & ~n33600;
  assign n33602 = ~n15675 & ~n33601;
  assign n33603 = ~i_hbusreq5 & ~n33602;
  assign n33604 = ~n33594 & ~n33603;
  assign n33605 = ~controllable_hgrant5 & ~n33604;
  assign n33606 = ~n15674 & ~n33605;
  assign n33607 = controllable_hmaster2 & ~n33606;
  assign n33608 = ~n33581 & ~n33607;
  assign n33609 = controllable_hmaster1 & ~n33608;
  assign n33610 = ~controllable_hmaster1 & ~n33580;
  assign n33611 = ~n33609 & ~n33610;
  assign n33612 = ~i_hbusreq6 & ~n33611;
  assign n33613 = ~n33593 & ~n33612;
  assign n33614 = ~controllable_hgrant6 & ~n33613;
  assign n33615 = ~n15812 & ~n33614;
  assign n33616 = controllable_hmaster0 & ~n33615;
  assign n33617 = controllable_hmaster1 & ~n33580;
  assign n33618 = controllable_hmaster2 & ~n33580;
  assign n33619 = ~i_hbusreq9 & ~n24199;
  assign n33620 = ~n29570 & ~n33619;
  assign n33621 = ~i_hbusreq4 & ~n33620;
  assign n33622 = ~n29569 & ~n33621;
  assign n33623 = ~controllable_hgrant4 & ~n33622;
  assign n33624 = ~n15822 & ~n33623;
  assign n33625 = ~i_hbusreq5 & ~n33624;
  assign n33626 = ~n29568 & ~n33625;
  assign n33627 = ~controllable_hgrant5 & ~n33626;
  assign n33628 = ~n15821 & ~n33627;
  assign n33629 = ~controllable_hmaster2 & ~n33628;
  assign n33630 = ~n33618 & ~n33629;
  assign n33631 = ~controllable_hmaster1 & ~n33630;
  assign n33632 = ~n33617 & ~n33631;
  assign n33633 = ~i_hbusreq6 & ~n33632;
  assign n33634 = ~n29603 & ~n33633;
  assign n33635 = ~controllable_hgrant6 & ~n33634;
  assign n33636 = ~n15818 & ~n33635;
  assign n33637 = ~controllable_hmaster0 & ~n33636;
  assign n33638 = ~n33616 & ~n33637;
  assign n33639 = ~i_hbusreq8 & ~n33638;
  assign n33640 = ~n33592 & ~n33639;
  assign n33641 = ~controllable_hmaster3 & ~n33640;
  assign n33642 = ~n33591 & ~n33641;
  assign n33643 = i_hlock7 & ~n33642;
  assign n33644 = i_hbusreq8 & ~n33535;
  assign n33645 = i_hbusreq6 & ~n33533;
  assign n33646 = i_hbusreq5 & ~n33526;
  assign n33647 = i_hbusreq4 & ~n24007;
  assign n33648 = i_hbusreq9 & ~n24007;
  assign n33649 = ~i_hbusreq9 & ~n24077;
  assign n33650 = ~n33648 & ~n33649;
  assign n33651 = ~i_hbusreq4 & ~n33650;
  assign n33652 = ~n33647 & ~n33651;
  assign n33653 = ~controllable_hgrant4 & ~n33652;
  assign n33654 = ~n15728 & ~n33653;
  assign n33655 = ~i_hbusreq5 & ~n33654;
  assign n33656 = ~n33646 & ~n33655;
  assign n33657 = ~controllable_hgrant5 & ~n33656;
  assign n33658 = ~n15727 & ~n33657;
  assign n33659 = controllable_hmaster1 & ~n33658;
  assign n33660 = controllable_hmaster2 & ~n33658;
  assign n33661 = ~i_hbusreq9 & ~n24158;
  assign n33662 = ~n29634 & ~n33661;
  assign n33663 = ~i_hbusreq4 & ~n33662;
  assign n33664 = ~n29633 & ~n33663;
  assign n33665 = ~controllable_hgrant4 & ~n33664;
  assign n33666 = ~n15675 & ~n33665;
  assign n33667 = ~i_hbusreq5 & ~n33666;
  assign n33668 = ~n29632 & ~n33667;
  assign n33669 = ~controllable_hgrant5 & ~n33668;
  assign n33670 = ~n15674 & ~n33669;
  assign n33671 = ~controllable_hmaster2 & ~n33670;
  assign n33672 = ~n33660 & ~n33671;
  assign n33673 = ~controllable_hmaster1 & ~n33672;
  assign n33674 = ~n33659 & ~n33673;
  assign n33675 = ~i_hbusreq6 & ~n33674;
  assign n33676 = ~n33645 & ~n33675;
  assign n33677 = ~controllable_hgrant6 & ~n33676;
  assign n33678 = ~n15672 & ~n33677;
  assign n33679 = ~i_hbusreq8 & ~n33678;
  assign n33680 = ~n33644 & ~n33679;
  assign n33681 = controllable_hmaster3 & ~n33680;
  assign n33682 = i_hbusreq8 & ~n33548;
  assign n33683 = i_hbusreq6 & ~n33544;
  assign n33684 = i_hbusreq5 & ~n33538;
  assign n33685 = i_hbusreq4 & ~n24026;
  assign n33686 = i_hbusreq9 & ~n24026;
  assign n33687 = ~i_hbusreq9 & ~n24117;
  assign n33688 = ~n33686 & ~n33687;
  assign n33689 = ~i_hbusreq4 & ~n33688;
  assign n33690 = ~n33685 & ~n33689;
  assign n33691 = ~controllable_hgrant4 & ~n33690;
  assign n33692 = ~n15675 & ~n33691;
  assign n33693 = ~i_hbusreq5 & ~n33692;
  assign n33694 = ~n33684 & ~n33693;
  assign n33695 = ~controllable_hgrant5 & ~n33694;
  assign n33696 = ~n15674 & ~n33695;
  assign n33697 = controllable_hmaster2 & ~n33696;
  assign n33698 = ~n33671 & ~n33697;
  assign n33699 = controllable_hmaster1 & ~n33698;
  assign n33700 = ~controllable_hmaster1 & ~n33670;
  assign n33701 = ~n33699 & ~n33700;
  assign n33702 = ~i_hbusreq6 & ~n33701;
  assign n33703 = ~n33683 & ~n33702;
  assign n33704 = ~controllable_hgrant6 & ~n33703;
  assign n33705 = ~n15812 & ~n33704;
  assign n33706 = controllable_hmaster0 & ~n33705;
  assign n33707 = controllable_hmaster1 & ~n33670;
  assign n33708 = controllable_hmaster2 & ~n33670;
  assign n33709 = ~i_hbusreq9 & ~n24209;
  assign n33710 = ~n29634 & ~n33709;
  assign n33711 = ~i_hbusreq4 & ~n33710;
  assign n33712 = ~n29633 & ~n33711;
  assign n33713 = ~controllable_hgrant4 & ~n33712;
  assign n33714 = ~n15822 & ~n33713;
  assign n33715 = ~i_hbusreq5 & ~n33714;
  assign n33716 = ~n29632 & ~n33715;
  assign n33717 = ~controllable_hgrant5 & ~n33716;
  assign n33718 = ~n15821 & ~n33717;
  assign n33719 = ~controllable_hmaster2 & ~n33718;
  assign n33720 = ~n33708 & ~n33719;
  assign n33721 = ~controllable_hmaster1 & ~n33720;
  assign n33722 = ~n33707 & ~n33721;
  assign n33723 = ~i_hbusreq6 & ~n33722;
  assign n33724 = ~n29667 & ~n33723;
  assign n33725 = ~controllable_hgrant6 & ~n33724;
  assign n33726 = ~n15818 & ~n33725;
  assign n33727 = ~controllable_hmaster0 & ~n33726;
  assign n33728 = ~n33706 & ~n33727;
  assign n33729 = ~i_hbusreq8 & ~n33728;
  assign n33730 = ~n33682 & ~n33729;
  assign n33731 = ~controllable_hmaster3 & ~n33730;
  assign n33732 = ~n33681 & ~n33731;
  assign n33733 = ~i_hlock7 & ~n33732;
  assign n33734 = ~n33643 & ~n33733;
  assign n33735 = ~i_hbusreq7 & ~n33734;
  assign n33736 = ~n33553 & ~n33735;
  assign n33737 = n7924 & ~n33736;
  assign n33738 = ~n33497 & ~n33737;
  assign n33739 = n8214 & ~n33738;
  assign n33740 = ~n33461 & ~n33739;
  assign n33741 = n8202 & ~n33740;
  assign n33742 = ~n23818 & ~n33741;
  assign n33743 = n7920 & ~n33742;
  assign n33744 = ~n33459 & ~n33743;
  assign n33745 = n7728 & ~n33744;
  assign n33746 = ~n7920 & ~n33441;
  assign n33747 = ~n24264 & ~n32395;
  assign n33748 = ~n8214 & ~n33747;
  assign n33749 = n8214 & ~n32396;
  assign n33750 = ~n33748 & ~n33749;
  assign n33751 = n8202 & ~n33750;
  assign n33752 = ~n24261 & ~n33751;
  assign n33753 = n7920 & ~n33752;
  assign n33754 = ~n33746 & ~n33753;
  assign n33755 = ~n7728 & ~n33754;
  assign n33756 = ~n33745 & ~n33755;
  assign n33757 = ~n7723 & ~n33756;
  assign n33758 = ~n7723 & ~n33757;
  assign n33759 = ~n7714 & ~n33758;
  assign n33760 = ~n7714 & ~n33759;
  assign n33761 = n7705 & ~n33760;
  assign n33762 = ~n24281 & ~n26890;
  assign n33763 = ~controllable_hgrant6 & ~n33762;
  assign n33764 = ~n15890 & ~n33763;
  assign n33765 = controllable_hmaster0 & ~n33764;
  assign n33766 = ~n9099 & ~n33765;
  assign n33767 = ~controllable_hmaster3 & ~n33766;
  assign n33768 = ~n9093 & ~n33767;
  assign n33769 = i_hbusreq7 & ~n33768;
  assign n33770 = i_hbusreq8 & ~n33766;
  assign n33771 = i_hbusreq6 & ~n33762;
  assign n33772 = ~n24293 & ~n26903;
  assign n33773 = ~i_hbusreq6 & ~n33772;
  assign n33774 = ~n33771 & ~n33773;
  assign n33775 = ~controllable_hgrant6 & ~n33774;
  assign n33776 = ~n15902 & ~n33775;
  assign n33777 = controllable_hmaster0 & ~n33776;
  assign n33778 = ~n9127 & ~n33777;
  assign n33779 = ~i_hbusreq8 & ~n33778;
  assign n33780 = ~n33770 & ~n33779;
  assign n33781 = ~controllable_hmaster3 & ~n33780;
  assign n33782 = ~n9117 & ~n33781;
  assign n33783 = ~i_hbusreq7 & ~n33782;
  assign n33784 = ~n33769 & ~n33783;
  assign n33785 = ~n7924 & ~n33784;
  assign n33786 = ~n24321 & ~n26936;
  assign n33787 = ~controllable_hgrant6 & ~n33786;
  assign n33788 = ~n15890 & ~n33787;
  assign n33789 = controllable_hmaster0 & ~n33788;
  assign n33790 = ~n13682 & ~n33789;
  assign n33791 = ~controllable_hmaster3 & ~n33790;
  assign n33792 = ~n27088 & ~n33791;
  assign n33793 = i_hbusreq7 & ~n33792;
  assign n33794 = i_hbusreq8 & ~n33790;
  assign n33795 = i_hbusreq6 & ~n33786;
  assign n33796 = ~n24360 & ~n26980;
  assign n33797 = ~i_hbusreq6 & ~n33796;
  assign n33798 = ~n33795 & ~n33797;
  assign n33799 = ~controllable_hgrant6 & ~n33798;
  assign n33800 = ~n15902 & ~n33799;
  assign n33801 = controllable_hmaster0 & ~n33800;
  assign n33802 = ~n13728 & ~n33801;
  assign n33803 = ~i_hbusreq8 & ~n33802;
  assign n33804 = ~n33794 & ~n33803;
  assign n33805 = ~controllable_hmaster3 & ~n33804;
  assign n33806 = ~n27174 & ~n33805;
  assign n33807 = ~i_hbusreq7 & ~n33806;
  assign n33808 = ~n33793 & ~n33807;
  assign n33809 = n7924 & ~n33808;
  assign n33810 = ~n33785 & ~n33809;
  assign n33811 = ~n8214 & ~n33810;
  assign n33812 = ~n24382 & ~n26894;
  assign n33813 = ~controllable_hmaster3 & ~n33812;
  assign n33814 = ~n9093 & ~n33813;
  assign n33815 = i_hbusreq7 & ~n33814;
  assign n33816 = i_hbusreq8 & ~n33812;
  assign n33817 = ~n24396 & ~n28107;
  assign n33818 = ~i_hbusreq8 & ~n33817;
  assign n33819 = ~n33816 & ~n33818;
  assign n33820 = ~controllable_hmaster3 & ~n33819;
  assign n33821 = ~n10867 & ~n33820;
  assign n33822 = ~i_hbusreq7 & ~n33821;
  assign n33823 = ~n33815 & ~n33822;
  assign n33824 = ~n7924 & ~n33823;
  assign n33825 = ~n24420 & ~n26940;
  assign n33826 = ~controllable_hmaster3 & ~n33825;
  assign n33827 = ~n27088 & ~n33826;
  assign n33828 = i_hbusreq7 & ~n33827;
  assign n33829 = i_hbusreq8 & ~n33825;
  assign n33830 = ~n24470 & ~n28131;
  assign n33831 = ~i_hbusreq8 & ~n33830;
  assign n33832 = ~n33829 & ~n33831;
  assign n33833 = ~controllable_hmaster3 & ~n33832;
  assign n33834 = ~n28232 & ~n33833;
  assign n33835 = ~i_hbusreq7 & ~n33834;
  assign n33836 = ~n33828 & ~n33835;
  assign n33837 = n7924 & ~n33836;
  assign n33838 = ~n33824 & ~n33837;
  assign n33839 = n8214 & ~n33838;
  assign n33840 = ~n33811 & ~n33839;
  assign n33841 = ~n8202 & ~n33840;
  assign n33842 = n8202 & ~n32396;
  assign n33843 = ~n33841 & ~n33842;
  assign n33844 = n7920 & ~n33843;
  assign n33845 = ~n33746 & ~n33844;
  assign n33846 = n7728 & ~n33845;
  assign n33847 = ~n24489 & ~n29737;
  assign n33848 = ~controllable_hgrant6 & ~n33847;
  assign n33849 = ~n13849 & ~n33848;
  assign n33850 = controllable_hmaster0 & ~n33849;
  assign n33851 = ~n19324 & ~n33850;
  assign n33852 = ~controllable_hmaster3 & ~n33851;
  assign n33853 = ~n30877 & ~n33852;
  assign n33854 = i_hlock7 & ~n33853;
  assign n33855 = ~n24489 & ~n29752;
  assign n33856 = ~controllable_hgrant6 & ~n33855;
  assign n33857 = ~n13951 & ~n33856;
  assign n33858 = controllable_hmaster0 & ~n33857;
  assign n33859 = ~n19324 & ~n33858;
  assign n33860 = ~controllable_hmaster3 & ~n33859;
  assign n33861 = ~n30877 & ~n33860;
  assign n33862 = ~i_hlock7 & ~n33861;
  assign n33863 = ~n33854 & ~n33862;
  assign n33864 = i_hbusreq7 & ~n33863;
  assign n33865 = i_hbusreq8 & ~n33851;
  assign n33866 = i_hbusreq6 & ~n33847;
  assign n33867 = ~n24511 & ~n29798;
  assign n33868 = ~i_hbusreq6 & ~n33867;
  assign n33869 = ~n33866 & ~n33868;
  assign n33870 = ~controllable_hgrant6 & ~n33869;
  assign n33871 = ~n16031 & ~n33870;
  assign n33872 = controllable_hmaster0 & ~n33871;
  assign n33873 = ~n19644 & ~n33872;
  assign n33874 = ~i_hbusreq8 & ~n33873;
  assign n33875 = ~n33865 & ~n33874;
  assign n33876 = ~controllable_hmaster3 & ~n33875;
  assign n33877 = ~n30896 & ~n33876;
  assign n33878 = i_hlock7 & ~n33877;
  assign n33879 = i_hbusreq8 & ~n33859;
  assign n33880 = i_hbusreq6 & ~n33855;
  assign n33881 = ~n24511 & ~n29828;
  assign n33882 = ~i_hbusreq6 & ~n33881;
  assign n33883 = ~n33880 & ~n33882;
  assign n33884 = ~controllable_hgrant6 & ~n33883;
  assign n33885 = ~n16068 & ~n33884;
  assign n33886 = controllable_hmaster0 & ~n33885;
  assign n33887 = ~n19644 & ~n33886;
  assign n33888 = ~i_hbusreq8 & ~n33887;
  assign n33889 = ~n33879 & ~n33888;
  assign n33890 = ~controllable_hmaster3 & ~n33889;
  assign n33891 = ~n30896 & ~n33890;
  assign n33892 = ~i_hlock7 & ~n33891;
  assign n33893 = ~n33878 & ~n33892;
  assign n33894 = ~i_hbusreq7 & ~n33893;
  assign n33895 = ~n33864 & ~n33894;
  assign n33896 = ~n7924 & ~n33895;
  assign n33897 = ~n24555 & ~n29871;
  assign n33898 = ~controllable_hgrant6 & ~n33897;
  assign n33899 = ~n13849 & ~n33898;
  assign n33900 = controllable_hmaster0 & ~n33899;
  assign n33901 = ~n19849 & ~n33900;
  assign n33902 = ~controllable_hmaster3 & ~n33901;
  assign n33903 = ~n30920 & ~n33902;
  assign n33904 = i_hlock7 & ~n33903;
  assign n33905 = ~n24555 & ~n29886;
  assign n33906 = ~controllable_hgrant6 & ~n33905;
  assign n33907 = ~n13951 & ~n33906;
  assign n33908 = controllable_hmaster0 & ~n33907;
  assign n33909 = ~n19849 & ~n33908;
  assign n33910 = ~controllable_hmaster3 & ~n33909;
  assign n33911 = ~n30920 & ~n33910;
  assign n33912 = ~i_hlock7 & ~n33911;
  assign n33913 = ~n33904 & ~n33912;
  assign n33914 = i_hbusreq7 & ~n33913;
  assign n33915 = i_hbusreq8 & ~n33901;
  assign n33916 = i_hbusreq6 & ~n33897;
  assign n33917 = ~n24604 & ~n29949;
  assign n33918 = ~i_hbusreq6 & ~n33917;
  assign n33919 = ~n33916 & ~n33918;
  assign n33920 = ~controllable_hgrant6 & ~n33919;
  assign n33921 = ~n16031 & ~n33920;
  assign n33922 = controllable_hmaster0 & ~n33921;
  assign n33923 = ~n20237 & ~n33922;
  assign n33924 = ~i_hbusreq8 & ~n33923;
  assign n33925 = ~n33915 & ~n33924;
  assign n33926 = ~controllable_hmaster3 & ~n33925;
  assign n33927 = ~n30939 & ~n33926;
  assign n33928 = i_hlock7 & ~n33927;
  assign n33929 = i_hbusreq8 & ~n33909;
  assign n33930 = i_hbusreq6 & ~n33905;
  assign n33931 = ~n24604 & ~n29979;
  assign n33932 = ~i_hbusreq6 & ~n33931;
  assign n33933 = ~n33930 & ~n33932;
  assign n33934 = ~controllable_hgrant6 & ~n33933;
  assign n33935 = ~n16068 & ~n33934;
  assign n33936 = controllable_hmaster0 & ~n33935;
  assign n33937 = ~n20237 & ~n33936;
  assign n33938 = ~i_hbusreq8 & ~n33937;
  assign n33939 = ~n33929 & ~n33938;
  assign n33940 = ~controllable_hmaster3 & ~n33939;
  assign n33941 = ~n30939 & ~n33940;
  assign n33942 = ~i_hlock7 & ~n33941;
  assign n33943 = ~n33928 & ~n33942;
  assign n33944 = ~i_hbusreq7 & ~n33943;
  assign n33945 = ~n33914 & ~n33944;
  assign n33946 = n7924 & ~n33945;
  assign n33947 = ~n33896 & ~n33946;
  assign n33948 = ~n8214 & ~n33947;
  assign n33949 = ~n24646 & ~n29741;
  assign n33950 = ~controllable_hmaster3 & ~n33949;
  assign n33951 = ~n30877 & ~n33950;
  assign n33952 = i_hlock7 & ~n33951;
  assign n33953 = ~n24646 & ~n29756;
  assign n33954 = ~controllable_hmaster3 & ~n33953;
  assign n33955 = ~n30877 & ~n33954;
  assign n33956 = ~i_hlock7 & ~n33955;
  assign n33957 = ~n33952 & ~n33956;
  assign n33958 = i_hbusreq7 & ~n33957;
  assign n33959 = i_hlock9 & ~n24750;
  assign n33960 = ~i_hlock9 & ~n24780;
  assign n33961 = ~n33959 & ~n33960;
  assign n33962 = ~i_hbusreq9 & ~n33961;
  assign n33963 = ~n30028 & ~n33962;
  assign n33964 = ~i_hbusreq4 & ~n33963;
  assign n33965 = ~n30027 & ~n33964;
  assign n33966 = ~controllable_hgrant4 & ~n33965;
  assign n33967 = ~n12676 & ~n33966;
  assign n33968 = ~i_hbusreq5 & ~n33967;
  assign n33969 = ~n30026 & ~n33968;
  assign n33970 = ~controllable_hgrant5 & ~n33969;
  assign n33971 = ~n12674 & ~n33970;
  assign n33972 = ~controllable_hmaster2 & ~n33971;
  assign n33973 = ~n24687 & ~n33972;
  assign n33974 = ~controllable_hmaster1 & ~n33973;
  assign n33975 = ~n24686 & ~n33974;
  assign n33976 = ~i_hbusreq6 & ~n33975;
  assign n33977 = ~n30025 & ~n33976;
  assign n33978 = ~controllable_hgrant6 & ~n33977;
  assign n33979 = ~n14849 & ~n33978;
  assign n33980 = controllable_hmaster0 & ~n33979;
  assign n33981 = ~n24769 & ~n33980;
  assign n33982 = i_hlock8 & ~n33981;
  assign n33983 = ~n24799 & ~n33980;
  assign n33984 = ~i_hlock8 & ~n33983;
  assign n33985 = ~n33982 & ~n33984;
  assign n33986 = ~i_hbusreq8 & ~n33985;
  assign n33987 = ~n30888 & ~n33986;
  assign n33988 = controllable_hmaster3 & ~n33987;
  assign n33989 = i_hbusreq8 & ~n33949;
  assign n33990 = ~i_hbusreq9 & ~n24708;
  assign n33991 = ~n29785 & ~n33990;
  assign n33992 = ~i_hbusreq4 & ~n33991;
  assign n33993 = ~n29784 & ~n33992;
  assign n33994 = ~controllable_hgrant4 & ~n33993;
  assign n33995 = ~n13524 & ~n33994;
  assign n33996 = ~i_hbusreq5 & ~n33995;
  assign n33997 = ~n29783 & ~n33996;
  assign n33998 = ~controllable_hgrant5 & ~n33997;
  assign n33999 = ~n13522 & ~n33998;
  assign n34000 = controllable_hmaster2 & ~n33999;
  assign n34001 = ~n24825 & ~n34000;
  assign n34002 = controllable_hmaster1 & ~n34001;
  assign n34003 = ~n24859 & ~n34002;
  assign n34004 = ~i_hbusreq6 & ~n34003;
  assign n34005 = ~n29782 & ~n34004;
  assign n34006 = ~controllable_hgrant6 & ~n34005;
  assign n34007 = ~n14995 & ~n34006;
  assign n34008 = controllable_hmaster0 & ~n34007;
  assign n34009 = ~n24915 & ~n34008;
  assign n34010 = ~i_hbusreq8 & ~n34009;
  assign n34011 = ~n33989 & ~n34010;
  assign n34012 = ~controllable_hmaster3 & ~n34011;
  assign n34013 = ~n33988 & ~n34012;
  assign n34014 = i_hlock7 & ~n34013;
  assign n34015 = i_hbusreq8 & ~n33953;
  assign n34016 = ~i_hbusreq9 & ~n24718;
  assign n34017 = ~n29815 & ~n34016;
  assign n34018 = ~i_hbusreq4 & ~n34017;
  assign n34019 = ~n29814 & ~n34018;
  assign n34020 = ~controllable_hgrant4 & ~n34019;
  assign n34021 = ~n13577 & ~n34020;
  assign n34022 = ~i_hbusreq5 & ~n34021;
  assign n34023 = ~n29813 & ~n34022;
  assign n34024 = ~controllable_hgrant5 & ~n34023;
  assign n34025 = ~n13575 & ~n34024;
  assign n34026 = controllable_hmaster2 & ~n34025;
  assign n34027 = ~n24825 & ~n34026;
  assign n34028 = controllable_hmaster1 & ~n34027;
  assign n34029 = ~n24859 & ~n34028;
  assign n34030 = ~i_hbusreq6 & ~n34029;
  assign n34031 = ~n29812 & ~n34030;
  assign n34032 = ~controllable_hgrant6 & ~n34031;
  assign n34033 = ~n15152 & ~n34032;
  assign n34034 = controllable_hmaster0 & ~n34033;
  assign n34035 = ~n24915 & ~n34034;
  assign n34036 = ~i_hbusreq8 & ~n34035;
  assign n34037 = ~n34015 & ~n34036;
  assign n34038 = ~controllable_hmaster3 & ~n34037;
  assign n34039 = ~n33988 & ~n34038;
  assign n34040 = ~i_hlock7 & ~n34039;
  assign n34041 = ~n34014 & ~n34040;
  assign n34042 = ~i_hbusreq7 & ~n34041;
  assign n34043 = ~n33958 & ~n34042;
  assign n34044 = ~n7924 & ~n34043;
  assign n34045 = ~n24960 & ~n29875;
  assign n34046 = ~controllable_hmaster3 & ~n34045;
  assign n34047 = ~n30920 & ~n34046;
  assign n34048 = i_hlock7 & ~n34047;
  assign n34049 = ~n24960 & ~n29890;
  assign n34050 = ~controllable_hmaster3 & ~n34049;
  assign n34051 = ~n30920 & ~n34050;
  assign n34052 = ~i_hlock7 & ~n34051;
  assign n34053 = ~n34048 & ~n34052;
  assign n34054 = i_hbusreq7 & ~n34053;
  assign n34055 = i_hlock9 & ~n25078;
  assign n34056 = ~i_hlock9 & ~n25108;
  assign n34057 = ~n34055 & ~n34056;
  assign n34058 = ~i_hbusreq9 & ~n34057;
  assign n34059 = ~n30097 & ~n34058;
  assign n34060 = ~i_hbusreq4 & ~n34059;
  assign n34061 = ~n30096 & ~n34060;
  assign n34062 = ~controllable_hgrant4 & ~n34061;
  assign n34063 = ~n12676 & ~n34062;
  assign n34064 = ~i_hbusreq5 & ~n34063;
  assign n34065 = ~n30095 & ~n34064;
  assign n34066 = ~controllable_hgrant5 & ~n34065;
  assign n34067 = ~n12674 & ~n34066;
  assign n34068 = ~controllable_hmaster2 & ~n34067;
  assign n34069 = ~n25015 & ~n34068;
  assign n34070 = ~controllable_hmaster1 & ~n34069;
  assign n34071 = ~n25014 & ~n34070;
  assign n34072 = ~i_hbusreq6 & ~n34071;
  assign n34073 = ~n30094 & ~n34072;
  assign n34074 = ~controllable_hgrant6 & ~n34073;
  assign n34075 = ~n14849 & ~n34074;
  assign n34076 = controllable_hmaster0 & ~n34075;
  assign n34077 = ~n25097 & ~n34076;
  assign n34078 = i_hlock8 & ~n34077;
  assign n34079 = ~n25127 & ~n34076;
  assign n34080 = ~i_hlock8 & ~n34079;
  assign n34081 = ~n34078 & ~n34080;
  assign n34082 = ~i_hbusreq8 & ~n34081;
  assign n34083 = ~n30931 & ~n34082;
  assign n34084 = controllable_hmaster3 & ~n34083;
  assign n34085 = i_hbusreq8 & ~n34045;
  assign n34086 = ~i_hbusreq9 & ~n25036;
  assign n34087 = ~n29936 & ~n34086;
  assign n34088 = ~i_hbusreq4 & ~n34087;
  assign n34089 = ~n29935 & ~n34088;
  assign n34090 = ~controllable_hgrant4 & ~n34089;
  assign n34091 = ~n13524 & ~n34090;
  assign n34092 = ~i_hbusreq5 & ~n34091;
  assign n34093 = ~n29934 & ~n34092;
  assign n34094 = ~controllable_hgrant5 & ~n34093;
  assign n34095 = ~n13522 & ~n34094;
  assign n34096 = controllable_hmaster2 & ~n34095;
  assign n34097 = ~n25153 & ~n34096;
  assign n34098 = controllable_hmaster1 & ~n34097;
  assign n34099 = ~n25187 & ~n34098;
  assign n34100 = ~i_hbusreq6 & ~n34099;
  assign n34101 = ~n29933 & ~n34100;
  assign n34102 = ~controllable_hgrant6 & ~n34101;
  assign n34103 = ~n14995 & ~n34102;
  assign n34104 = controllable_hmaster0 & ~n34103;
  assign n34105 = ~n25270 & ~n34104;
  assign n34106 = ~i_hbusreq8 & ~n34105;
  assign n34107 = ~n34085 & ~n34106;
  assign n34108 = ~controllable_hmaster3 & ~n34107;
  assign n34109 = ~n34084 & ~n34108;
  assign n34110 = i_hlock7 & ~n34109;
  assign n34111 = i_hbusreq8 & ~n34049;
  assign n34112 = ~i_hbusreq9 & ~n25046;
  assign n34113 = ~n29966 & ~n34112;
  assign n34114 = ~i_hbusreq4 & ~n34113;
  assign n34115 = ~n29965 & ~n34114;
  assign n34116 = ~controllable_hgrant4 & ~n34115;
  assign n34117 = ~n13577 & ~n34116;
  assign n34118 = ~i_hbusreq5 & ~n34117;
  assign n34119 = ~n29964 & ~n34118;
  assign n34120 = ~controllable_hgrant5 & ~n34119;
  assign n34121 = ~n13575 & ~n34120;
  assign n34122 = controllable_hmaster2 & ~n34121;
  assign n34123 = ~n25153 & ~n34122;
  assign n34124 = controllable_hmaster1 & ~n34123;
  assign n34125 = ~n25187 & ~n34124;
  assign n34126 = ~i_hbusreq6 & ~n34125;
  assign n34127 = ~n29963 & ~n34126;
  assign n34128 = ~controllable_hgrant6 & ~n34127;
  assign n34129 = ~n15152 & ~n34128;
  assign n34130 = controllable_hmaster0 & ~n34129;
  assign n34131 = ~n25270 & ~n34130;
  assign n34132 = ~i_hbusreq8 & ~n34131;
  assign n34133 = ~n34111 & ~n34132;
  assign n34134 = ~controllable_hmaster3 & ~n34133;
  assign n34135 = ~n34084 & ~n34134;
  assign n34136 = ~i_hlock7 & ~n34135;
  assign n34137 = ~n34110 & ~n34136;
  assign n34138 = ~i_hbusreq7 & ~n34137;
  assign n34139 = ~n34054 & ~n34138;
  assign n34140 = n7924 & ~n34139;
  assign n34141 = ~n34044 & ~n34140;
  assign n34142 = n8214 & ~n34141;
  assign n34143 = ~n33948 & ~n34142;
  assign n34144 = ~n8202 & ~n34143;
  assign n34145 = ~n33842 & ~n34144;
  assign n34146 = n7920 & ~n34145;
  assign n34147 = ~n33746 & ~n34146;
  assign n34148 = ~n7728 & ~n34147;
  assign n34149 = ~n33846 & ~n34148;
  assign n34150 = n7723 & ~n34149;
  assign n34151 = ~n7723 & ~n34147;
  assign n34152 = ~n34150 & ~n34151;
  assign n34153 = n7714 & ~n34152;
  assign n34154 = n7723 & ~n34147;
  assign n34155 = ~n30300 & ~n31029;
  assign n34156 = ~controllable_hmaster1 & ~n34155;
  assign n34157 = ~n31023 & ~n34156;
  assign n34158 = ~controllable_hgrant6 & ~n34157;
  assign n34159 = ~n13849 & ~n34158;
  assign n34160 = controllable_hmaster0 & ~n34159;
  assign n34161 = ~n31074 & ~n34160;
  assign n34162 = ~controllable_hmaster3 & ~n34161;
  assign n34163 = ~n31871 & ~n34162;
  assign n34164 = i_hlock7 & ~n34163;
  assign n34165 = ~n30403 & ~n31136;
  assign n34166 = ~controllable_hmaster1 & ~n34165;
  assign n34167 = ~n31130 & ~n34166;
  assign n34168 = ~controllable_hgrant6 & ~n34167;
  assign n34169 = ~n13951 & ~n34168;
  assign n34170 = controllable_hmaster0 & ~n34169;
  assign n34171 = ~n31181 & ~n34170;
  assign n34172 = ~controllable_hmaster3 & ~n34171;
  assign n34173 = ~n31893 & ~n34172;
  assign n34174 = ~i_hlock7 & ~n34173;
  assign n34175 = ~n34164 & ~n34174;
  assign n34176 = i_hbusreq7 & ~n34175;
  assign n34177 = i_hbusreq8 & ~n34161;
  assign n34178 = i_hbusreq6 & ~n34157;
  assign n34179 = ~i_hbusreq9 & ~n25342;
  assign n34180 = ~n30571 & ~n34179;
  assign n34181 = ~i_hbusreq4 & ~n34180;
  assign n34182 = ~n30570 & ~n34181;
  assign n34183 = ~controllable_hgrant4 & ~n34182;
  assign n34184 = ~n15030 & ~n34183;
  assign n34185 = ~i_hbusreq5 & ~n34184;
  assign n34186 = ~n30569 & ~n34185;
  assign n34187 = ~controllable_hgrant5 & ~n34186;
  assign n34188 = ~n15029 & ~n34187;
  assign n34189 = ~controllable_hmaster2 & ~n34188;
  assign n34190 = ~n31320 & ~n34189;
  assign n34191 = ~controllable_hmaster1 & ~n34190;
  assign n34192 = ~n31311 & ~n34191;
  assign n34193 = ~i_hbusreq6 & ~n34192;
  assign n34194 = ~n34178 & ~n34193;
  assign n34195 = ~controllable_hgrant6 & ~n34194;
  assign n34196 = ~n16031 & ~n34195;
  assign n34197 = controllable_hmaster0 & ~n34196;
  assign n34198 = ~n31403 & ~n34197;
  assign n34199 = ~i_hbusreq8 & ~n34198;
  assign n34200 = ~n34177 & ~n34199;
  assign n34201 = ~controllable_hmaster3 & ~n34200;
  assign n34202 = ~n31920 & ~n34201;
  assign n34203 = i_hlock7 & ~n34202;
  assign n34204 = i_hbusreq8 & ~n34171;
  assign n34205 = i_hbusreq6 & ~n34167;
  assign n34206 = ~i_hbusreq9 & ~n25354;
  assign n34207 = ~n30779 & ~n34206;
  assign n34208 = ~i_hbusreq4 & ~n34207;
  assign n34209 = ~n30778 & ~n34208;
  assign n34210 = ~controllable_hgrant4 & ~n34209;
  assign n34211 = ~n15030 & ~n34210;
  assign n34212 = ~i_hbusreq5 & ~n34211;
  assign n34213 = ~n30777 & ~n34212;
  assign n34214 = ~controllable_hgrant5 & ~n34213;
  assign n34215 = ~n15029 & ~n34214;
  assign n34216 = ~controllable_hmaster2 & ~n34215;
  assign n34217 = ~n31542 & ~n34216;
  assign n34218 = ~controllable_hmaster1 & ~n34217;
  assign n34219 = ~n31533 & ~n34218;
  assign n34220 = ~i_hbusreq6 & ~n34219;
  assign n34221 = ~n34205 & ~n34220;
  assign n34222 = ~controllable_hgrant6 & ~n34221;
  assign n34223 = ~n16068 & ~n34222;
  assign n34224 = controllable_hmaster0 & ~n34223;
  assign n34225 = ~n31625 & ~n34224;
  assign n34226 = ~i_hbusreq8 & ~n34225;
  assign n34227 = ~n34204 & ~n34226;
  assign n34228 = ~controllable_hmaster3 & ~n34227;
  assign n34229 = ~n31953 & ~n34228;
  assign n34230 = ~i_hlock7 & ~n34229;
  assign n34231 = ~n34203 & ~n34230;
  assign n34232 = ~i_hbusreq7 & ~n34231;
  assign n34233 = ~n34176 & ~n34232;
  assign n34234 = n7924 & ~n34233;
  assign n34235 = ~n33896 & ~n34234;
  assign n34236 = ~n8214 & ~n34235;
  assign n34237 = ~n30327 & ~n31056;
  assign n34238 = ~controllable_hmaster1 & ~n34237;
  assign n34239 = ~n31048 & ~n34238;
  assign n34240 = i_hlock6 & ~n34239;
  assign n34241 = ~n31068 & ~n34238;
  assign n34242 = ~i_hlock6 & ~n34241;
  assign n34243 = ~n34240 & ~n34242;
  assign n34244 = ~controllable_hgrant6 & ~n34243;
  assign n34245 = ~n13894 & ~n34244;
  assign n34246 = ~controllable_hmaster0 & ~n34245;
  assign n34247 = ~n31040 & ~n34246;
  assign n34248 = ~controllable_hmaster3 & ~n34247;
  assign n34249 = ~n31871 & ~n34248;
  assign n34250 = i_hlock7 & ~n34249;
  assign n34251 = ~n30430 & ~n31163;
  assign n34252 = ~controllable_hmaster1 & ~n34251;
  assign n34253 = ~n31155 & ~n34252;
  assign n34254 = i_hlock6 & ~n34253;
  assign n34255 = ~n31175 & ~n34252;
  assign n34256 = ~i_hlock6 & ~n34255;
  assign n34257 = ~n34254 & ~n34256;
  assign n34258 = ~controllable_hgrant6 & ~n34257;
  assign n34259 = ~n13894 & ~n34258;
  assign n34260 = ~controllable_hmaster0 & ~n34259;
  assign n34261 = ~n31147 & ~n34260;
  assign n34262 = ~controllable_hmaster3 & ~n34261;
  assign n34263 = ~n31893 & ~n34262;
  assign n34264 = ~i_hlock7 & ~n34263;
  assign n34265 = ~n34250 & ~n34264;
  assign n34266 = i_hbusreq7 & ~n34265;
  assign n34267 = ~i_hbusreq9 & ~n25444;
  assign n34268 = ~n31192 & ~n34267;
  assign n34269 = ~i_hbusreq4 & ~n34268;
  assign n34270 = ~n31191 & ~n34269;
  assign n34271 = ~controllable_hgrant4 & ~n34270;
  assign n34272 = ~n14875 & ~n34271;
  assign n34273 = ~i_hbusreq5 & ~n34272;
  assign n34274 = ~n31190 & ~n34273;
  assign n34275 = ~controllable_hgrant5 & ~n34274;
  assign n34276 = ~n14874 & ~n34275;
  assign n34277 = controllable_hmaster1 & ~n34276;
  assign n34278 = controllable_hmaster2 & ~n34276;
  assign n34279 = ~i_hlock9 & ~n25593;
  assign n34280 = ~n25550 & ~n34279;
  assign n34281 = ~i_hbusreq9 & ~n34280;
  assign n34282 = ~n31710 & ~n34281;
  assign n34283 = ~i_hbusreq4 & ~n34282;
  assign n34284 = ~n31709 & ~n34283;
  assign n34285 = ~controllable_hgrant4 & ~n34284;
  assign n34286 = ~n12676 & ~n34285;
  assign n34287 = ~i_hbusreq5 & ~n34286;
  assign n34288 = ~n31708 & ~n34287;
  assign n34289 = ~controllable_hgrant5 & ~n34288;
  assign n34290 = ~n12674 & ~n34289;
  assign n34291 = ~controllable_hmaster2 & ~n34290;
  assign n34292 = ~n34278 & ~n34291;
  assign n34293 = ~controllable_hmaster1 & ~n34292;
  assign n34294 = ~n34277 & ~n34293;
  assign n34295 = ~i_hbusreq6 & ~n34294;
  assign n34296 = ~n31707 & ~n34295;
  assign n34297 = ~controllable_hgrant6 & ~n34296;
  assign n34298 = ~n14849 & ~n34297;
  assign n34299 = controllable_hmaster0 & ~n34298;
  assign n34300 = ~i_hbusreq9 & ~n25549;
  assign n34301 = ~n31229 & ~n34300;
  assign n34302 = ~i_hbusreq4 & ~n34301;
  assign n34303 = ~n31228 & ~n34302;
  assign n34304 = ~controllable_hgrant4 & ~n34303;
  assign n34305 = ~n13524 & ~n34304;
  assign n34306 = ~i_hbusreq5 & ~n34305;
  assign n34307 = ~n31227 & ~n34306;
  assign n34308 = ~controllable_hgrant5 & ~n34307;
  assign n34309 = ~n13522 & ~n34308;
  assign n34310 = ~controllable_hmaster2 & ~n34309;
  assign n34311 = ~n34278 & ~n34310;
  assign n34312 = ~controllable_hmaster1 & ~n34311;
  assign n34313 = ~n34277 & ~n34312;
  assign n34314 = ~i_hbusreq6 & ~n34313;
  assign n34315 = ~n31226 & ~n34314;
  assign n34316 = ~controllable_hgrant6 & ~n34315;
  assign n34317 = ~n14927 & ~n34316;
  assign n34318 = ~controllable_hmaster0 & ~n34317;
  assign n34319 = ~n34299 & ~n34318;
  assign n34320 = i_hlock8 & ~n34319;
  assign n34321 = ~i_hbusreq9 & ~n25593;
  assign n34322 = ~n31254 & ~n34321;
  assign n34323 = ~i_hbusreq4 & ~n34322;
  assign n34324 = ~n31253 & ~n34323;
  assign n34325 = ~controllable_hgrant4 & ~n34324;
  assign n34326 = ~n13577 & ~n34325;
  assign n34327 = ~i_hbusreq5 & ~n34326;
  assign n34328 = ~n31252 & ~n34327;
  assign n34329 = ~controllable_hgrant5 & ~n34328;
  assign n34330 = ~n13575 & ~n34329;
  assign n34331 = ~controllable_hmaster2 & ~n34330;
  assign n34332 = ~n34278 & ~n34331;
  assign n34333 = ~controllable_hmaster1 & ~n34332;
  assign n34334 = ~n34277 & ~n34333;
  assign n34335 = ~i_hbusreq6 & ~n34334;
  assign n34336 = ~n31251 & ~n34335;
  assign n34337 = ~controllable_hgrant6 & ~n34336;
  assign n34338 = ~n14960 & ~n34337;
  assign n34339 = ~controllable_hmaster0 & ~n34338;
  assign n34340 = ~n34299 & ~n34339;
  assign n34341 = ~i_hlock8 & ~n34340;
  assign n34342 = ~n34320 & ~n34341;
  assign n34343 = ~i_hbusreq8 & ~n34342;
  assign n34344 = ~n31912 & ~n34343;
  assign n34345 = controllable_hmaster3 & ~n34344;
  assign n34346 = i_hbusreq8 & ~n34247;
  assign n34347 = ~i_hbusreq9 & ~n25499;
  assign n34348 = ~n31284 & ~n34347;
  assign n34349 = ~i_hbusreq4 & ~n34348;
  assign n34350 = ~n31283 & ~n34349;
  assign n34351 = ~controllable_hgrant4 & ~n34350;
  assign n34352 = ~n13524 & ~n34351;
  assign n34353 = ~i_hbusreq5 & ~n34352;
  assign n34354 = ~n31282 & ~n34353;
  assign n34355 = ~controllable_hgrant5 & ~n34354;
  assign n34356 = ~n13522 & ~n34355;
  assign n34357 = controllable_hmaster2 & ~n34356;
  assign n34358 = ~i_hbusreq9 & ~n25639;
  assign n34359 = ~n31298 & ~n34358;
  assign n34360 = ~i_hbusreq4 & ~n34359;
  assign n34361 = ~n31297 & ~n34360;
  assign n34362 = ~controllable_hgrant4 & ~n34361;
  assign n34363 = ~n14998 & ~n34362;
  assign n34364 = ~i_hbusreq5 & ~n34363;
  assign n34365 = ~n31296 & ~n34364;
  assign n34366 = ~controllable_hgrant5 & ~n34365;
  assign n34367 = ~n14997 & ~n34366;
  assign n34368 = ~controllable_hmaster2 & ~n34367;
  assign n34369 = ~n34357 & ~n34368;
  assign n34370 = controllable_hmaster1 & ~n34369;
  assign n34371 = i_hlock5 & ~n34305;
  assign n34372 = ~i_hlock5 & ~n34326;
  assign n34373 = ~n34371 & ~n34372;
  assign n34374 = ~i_hbusreq5 & ~n34373;
  assign n34375 = ~n31312 & ~n34374;
  assign n34376 = ~controllable_hgrant5 & ~n34375;
  assign n34377 = ~n15020 & ~n34376;
  assign n34378 = controllable_hmaster2 & ~n34377;
  assign n34379 = ~i_hbusreq9 & ~n25681;
  assign n34380 = ~n31323 & ~n34379;
  assign n34381 = ~i_hbusreq4 & ~n34380;
  assign n34382 = ~n31322 & ~n34381;
  assign n34383 = ~controllable_hgrant4 & ~n34382;
  assign n34384 = ~n15030 & ~n34383;
  assign n34385 = ~i_hbusreq5 & ~n34384;
  assign n34386 = ~n31321 & ~n34385;
  assign n34387 = ~controllable_hgrant5 & ~n34386;
  assign n34388 = ~n15029 & ~n34387;
  assign n34389 = ~controllable_hmaster2 & ~n34388;
  assign n34390 = ~n34378 & ~n34389;
  assign n34391 = ~controllable_hmaster1 & ~n34390;
  assign n34392 = ~n34370 & ~n34391;
  assign n34393 = ~i_hbusreq6 & ~n34392;
  assign n34394 = ~n31281 & ~n34393;
  assign n34395 = ~controllable_hgrant6 & ~n34394;
  assign n34396 = ~n14995 & ~n34395;
  assign n34397 = controllable_hmaster0 & ~n34396;
  assign n34398 = i_hbusreq6 & ~n34243;
  assign n34399 = controllable_hmaster2 & ~n34309;
  assign n34400 = ~i_hbusreq9 & ~n25724;
  assign n34401 = ~n31347 & ~n34400;
  assign n34402 = ~i_hbusreq4 & ~n34401;
  assign n34403 = ~n31346 & ~n34402;
  assign n34404 = ~controllable_hgrant4 & ~n34403;
  assign n34405 = ~n15065 & ~n34404;
  assign n34406 = ~i_hbusreq5 & ~n34405;
  assign n34407 = ~n31345 & ~n34406;
  assign n34408 = ~controllable_hgrant5 & ~n34407;
  assign n34409 = ~n15064 & ~n34408;
  assign n34410 = ~controllable_hmaster2 & ~n34409;
  assign n34411 = ~n34399 & ~n34410;
  assign n34412 = controllable_hmaster1 & ~n34411;
  assign n34413 = i_hlock4 & ~n34301;
  assign n34414 = ~i_hlock4 & ~n34322;
  assign n34415 = ~n34413 & ~n34414;
  assign n34416 = ~i_hbusreq4 & ~n34415;
  assign n34417 = ~n31362 & ~n34416;
  assign n34418 = ~controllable_hgrant4 & ~n34417;
  assign n34419 = ~n15091 & ~n34418;
  assign n34420 = ~i_hbusreq5 & ~n34419;
  assign n34421 = ~n31361 & ~n34420;
  assign n34422 = ~controllable_hgrant5 & ~n34421;
  assign n34423 = ~n15090 & ~n34422;
  assign n34424 = controllable_hmaster2 & ~n34423;
  assign n34425 = ~n32193 & ~n34424;
  assign n34426 = ~controllable_hmaster1 & ~n34425;
  assign n34427 = ~n34412 & ~n34426;
  assign n34428 = i_hlock6 & ~n34427;
  assign n34429 = controllable_hmaster2 & ~n34330;
  assign n34430 = ~n34410 & ~n34429;
  assign n34431 = controllable_hmaster1 & ~n34430;
  assign n34432 = ~n34426 & ~n34431;
  assign n34433 = ~i_hlock6 & ~n34432;
  assign n34434 = ~n34428 & ~n34433;
  assign n34435 = ~i_hbusreq6 & ~n34434;
  assign n34436 = ~n34398 & ~n34435;
  assign n34437 = ~controllable_hgrant6 & ~n34436;
  assign n34438 = ~n15063 & ~n34437;
  assign n34439 = ~controllable_hmaster0 & ~n34438;
  assign n34440 = ~n34397 & ~n34439;
  assign n34441 = ~i_hbusreq8 & ~n34440;
  assign n34442 = ~n34346 & ~n34441;
  assign n34443 = ~controllable_hmaster3 & ~n34442;
  assign n34444 = ~n34345 & ~n34443;
  assign n34445 = i_hlock7 & ~n34444;
  assign n34446 = ~i_hbusreq9 & ~n25462;
  assign n34447 = ~n31414 & ~n34446;
  assign n34448 = ~i_hbusreq4 & ~n34447;
  assign n34449 = ~n31413 & ~n34448;
  assign n34450 = ~controllable_hgrant4 & ~n34449;
  assign n34451 = ~n14875 & ~n34450;
  assign n34452 = ~i_hbusreq5 & ~n34451;
  assign n34453 = ~n31412 & ~n34452;
  assign n34454 = ~controllable_hgrant5 & ~n34453;
  assign n34455 = ~n14874 & ~n34454;
  assign n34456 = controllable_hmaster1 & ~n34455;
  assign n34457 = controllable_hmaster2 & ~n34455;
  assign n34458 = i_hlock9 & ~n25561;
  assign n34459 = ~n25604 & ~n34458;
  assign n34460 = ~i_hbusreq9 & ~n34459;
  assign n34461 = ~n31786 & ~n34460;
  assign n34462 = ~i_hbusreq4 & ~n34461;
  assign n34463 = ~n31785 & ~n34462;
  assign n34464 = ~controllable_hgrant4 & ~n34463;
  assign n34465 = ~n12676 & ~n34464;
  assign n34466 = ~i_hbusreq5 & ~n34465;
  assign n34467 = ~n31784 & ~n34466;
  assign n34468 = ~controllable_hgrant5 & ~n34467;
  assign n34469 = ~n12674 & ~n34468;
  assign n34470 = ~controllable_hmaster2 & ~n34469;
  assign n34471 = ~n34457 & ~n34470;
  assign n34472 = ~controllable_hmaster1 & ~n34471;
  assign n34473 = ~n34456 & ~n34472;
  assign n34474 = ~i_hbusreq6 & ~n34473;
  assign n34475 = ~n31783 & ~n34474;
  assign n34476 = ~controllable_hgrant6 & ~n34475;
  assign n34477 = ~n14849 & ~n34476;
  assign n34478 = controllable_hmaster0 & ~n34477;
  assign n34479 = ~i_hbusreq9 & ~n25561;
  assign n34480 = ~n31451 & ~n34479;
  assign n34481 = ~i_hbusreq4 & ~n34480;
  assign n34482 = ~n31450 & ~n34481;
  assign n34483 = ~controllable_hgrant4 & ~n34482;
  assign n34484 = ~n13524 & ~n34483;
  assign n34485 = ~i_hbusreq5 & ~n34484;
  assign n34486 = ~n31449 & ~n34485;
  assign n34487 = ~controllable_hgrant5 & ~n34486;
  assign n34488 = ~n13522 & ~n34487;
  assign n34489 = ~controllable_hmaster2 & ~n34488;
  assign n34490 = ~n34457 & ~n34489;
  assign n34491 = ~controllable_hmaster1 & ~n34490;
  assign n34492 = ~n34456 & ~n34491;
  assign n34493 = ~i_hbusreq6 & ~n34492;
  assign n34494 = ~n31448 & ~n34493;
  assign n34495 = ~controllable_hgrant6 & ~n34494;
  assign n34496 = ~n14927 & ~n34495;
  assign n34497 = ~controllable_hmaster0 & ~n34496;
  assign n34498 = ~n34478 & ~n34497;
  assign n34499 = i_hlock8 & ~n34498;
  assign n34500 = ~i_hbusreq9 & ~n25603;
  assign n34501 = ~n31476 & ~n34500;
  assign n34502 = ~i_hbusreq4 & ~n34501;
  assign n34503 = ~n31475 & ~n34502;
  assign n34504 = ~controllable_hgrant4 & ~n34503;
  assign n34505 = ~n13577 & ~n34504;
  assign n34506 = ~i_hbusreq5 & ~n34505;
  assign n34507 = ~n31474 & ~n34506;
  assign n34508 = ~controllable_hgrant5 & ~n34507;
  assign n34509 = ~n13575 & ~n34508;
  assign n34510 = ~controllable_hmaster2 & ~n34509;
  assign n34511 = ~n34457 & ~n34510;
  assign n34512 = ~controllable_hmaster1 & ~n34511;
  assign n34513 = ~n34456 & ~n34512;
  assign n34514 = ~i_hbusreq6 & ~n34513;
  assign n34515 = ~n31473 & ~n34514;
  assign n34516 = ~controllable_hgrant6 & ~n34515;
  assign n34517 = ~n14960 & ~n34516;
  assign n34518 = ~controllable_hmaster0 & ~n34517;
  assign n34519 = ~n34478 & ~n34518;
  assign n34520 = ~i_hlock8 & ~n34519;
  assign n34521 = ~n34499 & ~n34520;
  assign n34522 = ~i_hbusreq8 & ~n34521;
  assign n34523 = ~n31945 & ~n34522;
  assign n34524 = controllable_hmaster3 & ~n34523;
  assign n34525 = i_hbusreq8 & ~n34261;
  assign n34526 = ~i_hbusreq9 & ~n25517;
  assign n34527 = ~n31506 & ~n34526;
  assign n34528 = ~i_hbusreq4 & ~n34527;
  assign n34529 = ~n31505 & ~n34528;
  assign n34530 = ~controllable_hgrant4 & ~n34529;
  assign n34531 = ~n13577 & ~n34530;
  assign n34532 = ~i_hbusreq5 & ~n34531;
  assign n34533 = ~n31504 & ~n34532;
  assign n34534 = ~controllable_hgrant5 & ~n34533;
  assign n34535 = ~n13575 & ~n34534;
  assign n34536 = controllable_hmaster2 & ~n34535;
  assign n34537 = ~i_hbusreq9 & ~n25647;
  assign n34538 = ~n31520 & ~n34537;
  assign n34539 = ~i_hbusreq4 & ~n34538;
  assign n34540 = ~n31519 & ~n34539;
  assign n34541 = ~controllable_hgrant4 & ~n34540;
  assign n34542 = ~n14998 & ~n34541;
  assign n34543 = ~i_hbusreq5 & ~n34542;
  assign n34544 = ~n31518 & ~n34543;
  assign n34545 = ~controllable_hgrant5 & ~n34544;
  assign n34546 = ~n14997 & ~n34545;
  assign n34547 = ~controllable_hmaster2 & ~n34546;
  assign n34548 = ~n34536 & ~n34547;
  assign n34549 = controllable_hmaster1 & ~n34548;
  assign n34550 = i_hlock5 & ~n34484;
  assign n34551 = ~i_hlock5 & ~n34505;
  assign n34552 = ~n34550 & ~n34551;
  assign n34553 = ~i_hbusreq5 & ~n34552;
  assign n34554 = ~n31534 & ~n34553;
  assign n34555 = ~controllable_hgrant5 & ~n34554;
  assign n34556 = ~n15020 & ~n34555;
  assign n34557 = controllable_hmaster2 & ~n34556;
  assign n34558 = ~i_hbusreq9 & ~n25693;
  assign n34559 = ~n31545 & ~n34558;
  assign n34560 = ~i_hbusreq4 & ~n34559;
  assign n34561 = ~n31544 & ~n34560;
  assign n34562 = ~controllable_hgrant4 & ~n34561;
  assign n34563 = ~n15030 & ~n34562;
  assign n34564 = ~i_hbusreq5 & ~n34563;
  assign n34565 = ~n31543 & ~n34564;
  assign n34566 = ~controllable_hgrant5 & ~n34565;
  assign n34567 = ~n15029 & ~n34566;
  assign n34568 = ~controllable_hmaster2 & ~n34567;
  assign n34569 = ~n34557 & ~n34568;
  assign n34570 = ~controllable_hmaster1 & ~n34569;
  assign n34571 = ~n34549 & ~n34570;
  assign n34572 = ~i_hbusreq6 & ~n34571;
  assign n34573 = ~n31503 & ~n34572;
  assign n34574 = ~controllable_hgrant6 & ~n34573;
  assign n34575 = ~n15152 & ~n34574;
  assign n34576 = controllable_hmaster0 & ~n34575;
  assign n34577 = i_hbusreq6 & ~n34257;
  assign n34578 = controllable_hmaster2 & ~n34488;
  assign n34579 = ~i_hbusreq9 & ~n25734;
  assign n34580 = ~n31569 & ~n34579;
  assign n34581 = ~i_hbusreq4 & ~n34580;
  assign n34582 = ~n31568 & ~n34581;
  assign n34583 = ~controllable_hgrant4 & ~n34582;
  assign n34584 = ~n15065 & ~n34583;
  assign n34585 = ~i_hbusreq5 & ~n34584;
  assign n34586 = ~n31567 & ~n34585;
  assign n34587 = ~controllable_hgrant5 & ~n34586;
  assign n34588 = ~n15064 & ~n34587;
  assign n34589 = ~controllable_hmaster2 & ~n34588;
  assign n34590 = ~n34578 & ~n34589;
  assign n34591 = controllable_hmaster1 & ~n34590;
  assign n34592 = i_hlock4 & ~n34480;
  assign n34593 = ~i_hlock4 & ~n34501;
  assign n34594 = ~n34592 & ~n34593;
  assign n34595 = ~i_hbusreq4 & ~n34594;
  assign n34596 = ~n31584 & ~n34595;
  assign n34597 = ~controllable_hgrant4 & ~n34596;
  assign n34598 = ~n15091 & ~n34597;
  assign n34599 = ~i_hbusreq5 & ~n34598;
  assign n34600 = ~n31583 & ~n34599;
  assign n34601 = ~controllable_hgrant5 & ~n34600;
  assign n34602 = ~n15090 & ~n34601;
  assign n34603 = controllable_hmaster2 & ~n34602;
  assign n34604 = ~n32370 & ~n34603;
  assign n34605 = ~controllable_hmaster1 & ~n34604;
  assign n34606 = ~n34591 & ~n34605;
  assign n34607 = i_hlock6 & ~n34606;
  assign n34608 = controllable_hmaster2 & ~n34509;
  assign n34609 = ~n34589 & ~n34608;
  assign n34610 = controllable_hmaster1 & ~n34609;
  assign n34611 = ~n34605 & ~n34610;
  assign n34612 = ~i_hlock6 & ~n34611;
  assign n34613 = ~n34607 & ~n34612;
  assign n34614 = ~i_hbusreq6 & ~n34613;
  assign n34615 = ~n34577 & ~n34614;
  assign n34616 = ~controllable_hgrant6 & ~n34615;
  assign n34617 = ~n15063 & ~n34616;
  assign n34618 = ~controllable_hmaster0 & ~n34617;
  assign n34619 = ~n34576 & ~n34618;
  assign n34620 = ~i_hbusreq8 & ~n34619;
  assign n34621 = ~n34525 & ~n34620;
  assign n34622 = ~controllable_hmaster3 & ~n34621;
  assign n34623 = ~n34524 & ~n34622;
  assign n34624 = ~i_hlock7 & ~n34623;
  assign n34625 = ~n34445 & ~n34624;
  assign n34626 = ~i_hbusreq7 & ~n34625;
  assign n34627 = ~n34266 & ~n34626;
  assign n34628 = n7924 & ~n34627;
  assign n34629 = ~n34044 & ~n34628;
  assign n34630 = n8214 & ~n34629;
  assign n34631 = ~n34236 & ~n34630;
  assign n34632 = ~n8202 & ~n34631;
  assign n34633 = ~n33842 & ~n34632;
  assign n34634 = n7920 & ~n34633;
  assign n34635 = ~n28799 & ~n34634;
  assign n34636 = n7728 & ~n34635;
  assign n34637 = ~n32399 & ~n34636;
  assign n34638 = ~n7723 & ~n34637;
  assign n34639 = ~n34154 & ~n34638;
  assign n34640 = ~n7714 & ~n34639;
  assign n34641 = ~n34153 & ~n34640;
  assign n34642 = ~n7705 & ~n34641;
  assign n34643 = ~n33761 & ~n34642;
  assign n34644 = n7808 & ~n34643;
  assign n34645 = ~n33458 & ~n34644;
  assign n34646 = n8195 & ~n34645;
  assign n34647 = ~n33323 & ~n34646;
  assign n34648 = n8193 & ~n34647;
  assign n34649 = ~n32411 & ~n34648;
  assign n34650 = n8191 & ~n34649;
  assign n34651 = ~n10989 & ~n28706;
  assign n34652 = n7728 & ~n34651;
  assign n34653 = ~n11020 & ~n28726;
  assign n34654 = ~n7728 & ~n34653;
  assign n34655 = ~n34652 & ~n34654;
  assign n34656 = ~n7723 & ~n34655;
  assign n34657 = ~n7723 & ~n34656;
  assign n34658 = ~n7714 & ~n34657;
  assign n34659 = ~n7714 & ~n34658;
  assign n34660 = n7705 & ~n34659;
  assign n34661 = n7723 & ~n34653;
  assign n34662 = ~n11036 & ~n28744;
  assign n34663 = i_hlock7 & ~n34662;
  assign n34664 = ~n11036 & ~n28755;
  assign n34665 = ~i_hlock7 & ~n34664;
  assign n34666 = ~n34663 & ~n34665;
  assign n34667 = i_hbusreq7 & ~n34666;
  assign n34668 = ~n11051 & ~n28774;
  assign n34669 = i_hlock7 & ~n34668;
  assign n34670 = ~n11051 & ~n28791;
  assign n34671 = ~i_hlock7 & ~n34670;
  assign n34672 = ~n34669 & ~n34671;
  assign n34673 = ~i_hbusreq7 & ~n34672;
  assign n34674 = ~n34667 & ~n34673;
  assign n34675 = n7924 & ~n34674;
  assign n34676 = ~n8337 & ~n34675;
  assign n34677 = ~n7920 & ~n34676;
  assign n34678 = n7920 & ~n34653;
  assign n34679 = ~n34677 & ~n34678;
  assign n34680 = ~n7723 & ~n34679;
  assign n34681 = ~n34661 & ~n34680;
  assign n34682 = n7714 & ~n34681;
  assign n34683 = ~n7714 & ~n34676;
  assign n34684 = ~n34682 & ~n34683;
  assign n34685 = ~n7705 & ~n34684;
  assign n34686 = ~n34660 & ~n34685;
  assign n34687 = ~n7808 & ~n34686;
  assign n34688 = ~n7920 & ~n34651;
  assign n34689 = ~n29133 & ~n34688;
  assign n34690 = n7728 & ~n34689;
  assign n34691 = ~n7920 & ~n34653;
  assign n34692 = ~n29282 & ~n34691;
  assign n34693 = ~n7728 & ~n34692;
  assign n34694 = ~n34690 & ~n34693;
  assign n34695 = ~n7723 & ~n34694;
  assign n34696 = ~n7723 & ~n34695;
  assign n34697 = ~n7714 & ~n34696;
  assign n34698 = ~n7714 & ~n34697;
  assign n34699 = n7705 & ~n34698;
  assign n34700 = ~n29716 & ~n34691;
  assign n34701 = n7728 & ~n34700;
  assign n34702 = ~n30963 & ~n34691;
  assign n34703 = ~n7728 & ~n34702;
  assign n34704 = ~n34701 & ~n34703;
  assign n34705 = n7723 & ~n34704;
  assign n34706 = ~n7723 & ~n34702;
  assign n34707 = ~n34705 & ~n34706;
  assign n34708 = n7714 & ~n34707;
  assign n34709 = n7723 & ~n34702;
  assign n34710 = ~n31987 & ~n34677;
  assign n34711 = n7728 & ~n34710;
  assign n34712 = ~n32397 & ~n34677;
  assign n34713 = ~n7728 & ~n34712;
  assign n34714 = ~n34711 & ~n34713;
  assign n34715 = ~n7723 & ~n34714;
  assign n34716 = ~n34709 & ~n34715;
  assign n34717 = ~n7714 & ~n34716;
  assign n34718 = ~n34708 & ~n34717;
  assign n34719 = ~n7705 & ~n34718;
  assign n34720 = ~n34699 & ~n34719;
  assign n34721 = n7808 & ~n34720;
  assign n34722 = ~n34687 & ~n34721;
  assign n34723 = n8195 & ~n34722;
  assign n34724 = ~n8196 & ~n34723;
  assign n34725 = ~n8193 & ~n34724;
  assign n34726 = ~n9900 & ~n34677;
  assign n34727 = ~n7723 & ~n34726;
  assign n34728 = ~n9899 & ~n34727;
  assign n34729 = n7714 & ~n34728;
  assign n34730 = ~n34683 & ~n34729;
  assign n34731 = ~n7705 & ~n34730;
  assign n34732 = ~n9898 & ~n34731;
  assign n34733 = ~n7808 & ~n34732;
  assign n34734 = ~n33311 & ~n34677;
  assign n34735 = n7728 & ~n34734;
  assign n34736 = ~n34713 & ~n34735;
  assign n34737 = ~n7723 & ~n34736;
  assign n34738 = ~n32941 & ~n34737;
  assign n34739 = ~n7714 & ~n34738;
  assign n34740 = ~n32940 & ~n34739;
  assign n34741 = ~n7705 & ~n34740;
  assign n34742 = ~n22399 & ~n34741;
  assign n34743 = n7808 & ~n34742;
  assign n34744 = ~n34733 & ~n34743;
  assign n34745 = ~n8195 & ~n34744;
  assign n34746 = ~n11136 & ~n33339;
  assign n34747 = i_hlock7 & ~n34746;
  assign n34748 = ~n11136 & ~n33357;
  assign n34749 = ~i_hlock7 & ~n34748;
  assign n34750 = ~n34747 & ~n34749;
  assign n34751 = i_hbusreq7 & ~n34750;
  assign n34752 = ~n11164 & ~n33392;
  assign n34753 = i_hlock7 & ~n34752;
  assign n34754 = ~n11164 & ~n33425;
  assign n34755 = ~i_hlock7 & ~n34754;
  assign n34756 = ~n34753 & ~n34755;
  assign n34757 = ~i_hbusreq7 & ~n34756;
  assign n34758 = ~n34751 & ~n34757;
  assign n34759 = n7924 & ~n34758;
  assign n34760 = ~n10375 & ~n34759;
  assign n34761 = n8214 & ~n34760;
  assign n34762 = n8214 & ~n34761;
  assign n34763 = n8202 & ~n34762;
  assign n34764 = ~n10332 & ~n34763;
  assign n34765 = n7728 & ~n34764;
  assign n34766 = n8214 & ~n34676;
  assign n34767 = ~n8336 & ~n34766;
  assign n34768 = n8202 & ~n34767;
  assign n34769 = ~n10649 & ~n34768;
  assign n34770 = ~n7728 & ~n34769;
  assign n34771 = ~n34765 & ~n34770;
  assign n34772 = ~n7723 & ~n34771;
  assign n34773 = ~n7723 & ~n34772;
  assign n34774 = ~n7714 & ~n34773;
  assign n34775 = ~n7714 & ~n34774;
  assign n34776 = n7705 & ~n34775;
  assign n34777 = n7723 & ~n34769;
  assign n34778 = n7920 & ~n34769;
  assign n34779 = ~n34677 & ~n34778;
  assign n34780 = ~n7723 & ~n34779;
  assign n34781 = ~n34777 & ~n34780;
  assign n34782 = n7714 & ~n34781;
  assign n34783 = ~n34683 & ~n34782;
  assign n34784 = ~n7705 & ~n34783;
  assign n34785 = ~n34776 & ~n34784;
  assign n34786 = ~n7808 & ~n34785;
  assign n34787 = ~n7920 & ~n34764;
  assign n34788 = ~n33743 & ~n34787;
  assign n34789 = n7728 & ~n34788;
  assign n34790 = ~n7920 & ~n34769;
  assign n34791 = ~n33753 & ~n34790;
  assign n34792 = ~n7728 & ~n34791;
  assign n34793 = ~n34789 & ~n34792;
  assign n34794 = ~n7723 & ~n34793;
  assign n34795 = ~n7723 & ~n34794;
  assign n34796 = ~n7714 & ~n34795;
  assign n34797 = ~n7714 & ~n34796;
  assign n34798 = n7705 & ~n34797;
  assign n34799 = ~n33844 & ~n34790;
  assign n34800 = n7728 & ~n34799;
  assign n34801 = ~n34146 & ~n34790;
  assign n34802 = ~n7728 & ~n34801;
  assign n34803 = ~n34800 & ~n34802;
  assign n34804 = n7723 & ~n34803;
  assign n34805 = ~n7723 & ~n34801;
  assign n34806 = ~n34804 & ~n34805;
  assign n34807 = n7714 & ~n34806;
  assign n34808 = n7723 & ~n34801;
  assign n34809 = ~n34634 & ~n34677;
  assign n34810 = n7728 & ~n34809;
  assign n34811 = ~n34713 & ~n34810;
  assign n34812 = ~n7723 & ~n34811;
  assign n34813 = ~n34808 & ~n34812;
  assign n34814 = ~n7714 & ~n34813;
  assign n34815 = ~n34807 & ~n34814;
  assign n34816 = ~n7705 & ~n34815;
  assign n34817 = ~n34798 & ~n34816;
  assign n34818 = n7808 & ~n34817;
  assign n34819 = ~n34786 & ~n34818;
  assign n34820 = n8195 & ~n34819;
  assign n34821 = ~n34745 & ~n34820;
  assign n34822 = n8193 & ~n34821;
  assign n34823 = ~n34725 & ~n34822;
  assign n34824 = ~n8191 & ~n34823;
  assign n34825 = ~n34650 & ~n34824;
  assign n34826 = n8188 & ~n34825;
  assign n34827 = ~n11286 & ~n28706;
  assign n34828 = n7728 & ~n34827;
  assign n34829 = ~n11335 & ~n28726;
  assign n34830 = ~n7728 & ~n34829;
  assign n34831 = ~n34828 & ~n34830;
  assign n34832 = ~n7723 & ~n34831;
  assign n34833 = ~n7723 & ~n34832;
  assign n34834 = ~n7714 & ~n34833;
  assign n34835 = ~n7714 & ~n34834;
  assign n34836 = n7705 & ~n34835;
  assign n34837 = n7723 & ~n34829;
  assign n34838 = ~n11359 & ~n28744;
  assign n34839 = i_hlock7 & ~n34838;
  assign n34840 = ~n11359 & ~n28755;
  assign n34841 = ~i_hlock7 & ~n34840;
  assign n34842 = ~n34839 & ~n34841;
  assign n34843 = i_hbusreq7 & ~n34842;
  assign n34844 = ~n11385 & ~n28774;
  assign n34845 = i_hlock7 & ~n34844;
  assign n34846 = ~n11385 & ~n28791;
  assign n34847 = ~i_hlock7 & ~n34846;
  assign n34848 = ~n34845 & ~n34847;
  assign n34849 = ~i_hbusreq7 & ~n34848;
  assign n34850 = ~n34843 & ~n34849;
  assign n34851 = n7924 & ~n34850;
  assign n34852 = ~n8337 & ~n34851;
  assign n34853 = ~n7920 & ~n34852;
  assign n34854 = n7920 & ~n34829;
  assign n34855 = ~n34853 & ~n34854;
  assign n34856 = ~n7723 & ~n34855;
  assign n34857 = ~n34837 & ~n34856;
  assign n34858 = n7714 & ~n34857;
  assign n34859 = ~n7714 & ~n34852;
  assign n34860 = ~n34858 & ~n34859;
  assign n34861 = ~n7705 & ~n34860;
  assign n34862 = ~n34836 & ~n34861;
  assign n34863 = ~n7808 & ~n34862;
  assign n34864 = ~n7920 & ~n34827;
  assign n34865 = ~n29133 & ~n34864;
  assign n34866 = n7728 & ~n34865;
  assign n34867 = ~n7920 & ~n34829;
  assign n34868 = ~n29282 & ~n34867;
  assign n34869 = ~n7728 & ~n34868;
  assign n34870 = ~n34866 & ~n34869;
  assign n34871 = ~n7723 & ~n34870;
  assign n34872 = ~n7723 & ~n34871;
  assign n34873 = ~n7714 & ~n34872;
  assign n34874 = ~n7714 & ~n34873;
  assign n34875 = n7705 & ~n34874;
  assign n34876 = ~n29716 & ~n34867;
  assign n34877 = n7728 & ~n34876;
  assign n34878 = ~n30963 & ~n34867;
  assign n34879 = ~n7728 & ~n34878;
  assign n34880 = ~n34877 & ~n34879;
  assign n34881 = n7723 & ~n34880;
  assign n34882 = ~n7723 & ~n34878;
  assign n34883 = ~n34881 & ~n34882;
  assign n34884 = n7714 & ~n34883;
  assign n34885 = n7723 & ~n34878;
  assign n34886 = ~n31987 & ~n34853;
  assign n34887 = n7728 & ~n34886;
  assign n34888 = ~n32397 & ~n34853;
  assign n34889 = ~n7728 & ~n34888;
  assign n34890 = ~n34887 & ~n34889;
  assign n34891 = ~n7723 & ~n34890;
  assign n34892 = ~n34885 & ~n34891;
  assign n34893 = ~n7714 & ~n34892;
  assign n34894 = ~n34884 & ~n34893;
  assign n34895 = ~n7705 & ~n34894;
  assign n34896 = ~n34875 & ~n34895;
  assign n34897 = n7808 & ~n34896;
  assign n34898 = ~n34863 & ~n34897;
  assign n34899 = n8195 & ~n34898;
  assign n34900 = ~n8196 & ~n34899;
  assign n34901 = ~n8193 & ~n34900;
  assign n34902 = ~n9900 & ~n34853;
  assign n34903 = ~n7723 & ~n34902;
  assign n34904 = ~n9899 & ~n34903;
  assign n34905 = n7714 & ~n34904;
  assign n34906 = ~n34859 & ~n34905;
  assign n34907 = ~n7705 & ~n34906;
  assign n34908 = ~n9898 & ~n34907;
  assign n34909 = ~n7808 & ~n34908;
  assign n34910 = ~n33311 & ~n34853;
  assign n34911 = n7728 & ~n34910;
  assign n34912 = ~n34889 & ~n34911;
  assign n34913 = ~n7723 & ~n34912;
  assign n34914 = ~n32941 & ~n34913;
  assign n34915 = ~n7714 & ~n34914;
  assign n34916 = ~n32940 & ~n34915;
  assign n34917 = ~n7705 & ~n34916;
  assign n34918 = ~n22399 & ~n34917;
  assign n34919 = n7808 & ~n34918;
  assign n34920 = ~n34909 & ~n34919;
  assign n34921 = ~n8195 & ~n34920;
  assign n34922 = ~n11476 & ~n33339;
  assign n34923 = i_hlock7 & ~n34922;
  assign n34924 = ~n11476 & ~n33357;
  assign n34925 = ~i_hlock7 & ~n34924;
  assign n34926 = ~n34923 & ~n34925;
  assign n34927 = i_hbusreq7 & ~n34926;
  assign n34928 = ~n11504 & ~n33392;
  assign n34929 = i_hlock7 & ~n34928;
  assign n34930 = ~n11504 & ~n33425;
  assign n34931 = ~i_hlock7 & ~n34930;
  assign n34932 = ~n34929 & ~n34931;
  assign n34933 = ~i_hbusreq7 & ~n34932;
  assign n34934 = ~n34927 & ~n34933;
  assign n34935 = n7924 & ~n34934;
  assign n34936 = ~n10375 & ~n34935;
  assign n34937 = n8214 & ~n34936;
  assign n34938 = n8214 & ~n34937;
  assign n34939 = n8202 & ~n34938;
  assign n34940 = ~n10332 & ~n34939;
  assign n34941 = n7728 & ~n34940;
  assign n34942 = n8214 & ~n34852;
  assign n34943 = ~n8336 & ~n34942;
  assign n34944 = n8202 & ~n34943;
  assign n34945 = ~n10649 & ~n34944;
  assign n34946 = ~n7728 & ~n34945;
  assign n34947 = ~n34941 & ~n34946;
  assign n34948 = ~n7723 & ~n34947;
  assign n34949 = ~n7723 & ~n34948;
  assign n34950 = ~n7714 & ~n34949;
  assign n34951 = ~n7714 & ~n34950;
  assign n34952 = n7705 & ~n34951;
  assign n34953 = n7723 & ~n34945;
  assign n34954 = n7920 & ~n34945;
  assign n34955 = ~n34853 & ~n34954;
  assign n34956 = ~n7723 & ~n34955;
  assign n34957 = ~n34953 & ~n34956;
  assign n34958 = n7714 & ~n34957;
  assign n34959 = ~n34859 & ~n34958;
  assign n34960 = ~n7705 & ~n34959;
  assign n34961 = ~n34952 & ~n34960;
  assign n34962 = ~n7808 & ~n34961;
  assign n34963 = ~n7920 & ~n34940;
  assign n34964 = ~n33743 & ~n34963;
  assign n34965 = n7728 & ~n34964;
  assign n34966 = ~n7920 & ~n34945;
  assign n34967 = ~n33753 & ~n34966;
  assign n34968 = ~n7728 & ~n34967;
  assign n34969 = ~n34965 & ~n34968;
  assign n34970 = ~n7723 & ~n34969;
  assign n34971 = ~n7723 & ~n34970;
  assign n34972 = ~n7714 & ~n34971;
  assign n34973 = ~n7714 & ~n34972;
  assign n34974 = n7705 & ~n34973;
  assign n34975 = ~n33844 & ~n34966;
  assign n34976 = n7728 & ~n34975;
  assign n34977 = ~n34146 & ~n34966;
  assign n34978 = ~n7728 & ~n34977;
  assign n34979 = ~n34976 & ~n34978;
  assign n34980 = n7723 & ~n34979;
  assign n34981 = ~n7723 & ~n34977;
  assign n34982 = ~n34980 & ~n34981;
  assign n34983 = n7714 & ~n34982;
  assign n34984 = n7723 & ~n34977;
  assign n34985 = ~n34634 & ~n34853;
  assign n34986 = n7728 & ~n34985;
  assign n34987 = ~n34889 & ~n34986;
  assign n34988 = ~n7723 & ~n34987;
  assign n34989 = ~n34984 & ~n34988;
  assign n34990 = ~n7714 & ~n34989;
  assign n34991 = ~n34983 & ~n34990;
  assign n34992 = ~n7705 & ~n34991;
  assign n34993 = ~n34974 & ~n34992;
  assign n34994 = n7808 & ~n34993;
  assign n34995 = ~n34962 & ~n34994;
  assign n34996 = n8195 & ~n34995;
  assign n34997 = ~n34921 & ~n34996;
  assign n34998 = n8193 & ~n34997;
  assign n34999 = ~n34901 & ~n34998;
  assign n35000 = n8191 & ~n34999;
  assign n35001 = ~n11575 & ~n28706;
  assign n35002 = n7728 & ~n35001;
  assign n35003 = ~n11579 & ~n28726;
  assign n35004 = ~n7728 & ~n35003;
  assign n35005 = ~n35002 & ~n35004;
  assign n35006 = ~n7723 & ~n35005;
  assign n35007 = ~n7723 & ~n35006;
  assign n35008 = ~n7714 & ~n35007;
  assign n35009 = ~n7714 & ~n35008;
  assign n35010 = n7705 & ~n35009;
  assign n35011 = n7723 & ~n35003;
  assign n35012 = ~n11594 & ~n28744;
  assign n35013 = i_hlock7 & ~n35012;
  assign n35014 = ~n11594 & ~n28755;
  assign n35015 = ~i_hlock7 & ~n35014;
  assign n35016 = ~n35013 & ~n35015;
  assign n35017 = i_hbusreq7 & ~n35016;
  assign n35018 = ~n11605 & ~n28774;
  assign n35019 = i_hlock7 & ~n35018;
  assign n35020 = ~n11605 & ~n28791;
  assign n35021 = ~i_hlock7 & ~n35020;
  assign n35022 = ~n35019 & ~n35021;
  assign n35023 = ~i_hbusreq7 & ~n35022;
  assign n35024 = ~n35017 & ~n35023;
  assign n35025 = n7924 & ~n35024;
  assign n35026 = ~n8337 & ~n35025;
  assign n35027 = ~n7920 & ~n35026;
  assign n35028 = n7920 & ~n35003;
  assign n35029 = ~n35027 & ~n35028;
  assign n35030 = ~n7723 & ~n35029;
  assign n35031 = ~n35011 & ~n35030;
  assign n35032 = n7714 & ~n35031;
  assign n35033 = ~n7714 & ~n35026;
  assign n35034 = ~n35032 & ~n35033;
  assign n35035 = ~n7705 & ~n35034;
  assign n35036 = ~n35010 & ~n35035;
  assign n35037 = ~n7808 & ~n35036;
  assign n35038 = ~n7920 & ~n35001;
  assign n35039 = ~n29133 & ~n35038;
  assign n35040 = n7728 & ~n35039;
  assign n35041 = ~n7920 & ~n35003;
  assign n35042 = ~n29282 & ~n35041;
  assign n35043 = ~n7728 & ~n35042;
  assign n35044 = ~n35040 & ~n35043;
  assign n35045 = ~n7723 & ~n35044;
  assign n35046 = ~n7723 & ~n35045;
  assign n35047 = ~n7714 & ~n35046;
  assign n35048 = ~n7714 & ~n35047;
  assign n35049 = n7705 & ~n35048;
  assign n35050 = ~n29716 & ~n35041;
  assign n35051 = n7728 & ~n35050;
  assign n35052 = ~n30963 & ~n35041;
  assign n35053 = ~n7728 & ~n35052;
  assign n35054 = ~n35051 & ~n35053;
  assign n35055 = n7723 & ~n35054;
  assign n35056 = ~n7723 & ~n35052;
  assign n35057 = ~n35055 & ~n35056;
  assign n35058 = n7714 & ~n35057;
  assign n35059 = n7723 & ~n35052;
  assign n35060 = ~n31987 & ~n35027;
  assign n35061 = n7728 & ~n35060;
  assign n35062 = ~n32397 & ~n35027;
  assign n35063 = ~n7728 & ~n35062;
  assign n35064 = ~n35061 & ~n35063;
  assign n35065 = ~n7723 & ~n35064;
  assign n35066 = ~n35059 & ~n35065;
  assign n35067 = ~n7714 & ~n35066;
  assign n35068 = ~n35058 & ~n35067;
  assign n35069 = ~n7705 & ~n35068;
  assign n35070 = ~n35049 & ~n35069;
  assign n35071 = n7808 & ~n35070;
  assign n35072 = ~n35037 & ~n35071;
  assign n35073 = n8195 & ~n35072;
  assign n35074 = ~n8196 & ~n35073;
  assign n35075 = ~n8193 & ~n35074;
  assign n35076 = ~n9900 & ~n35027;
  assign n35077 = ~n7723 & ~n35076;
  assign n35078 = ~n9899 & ~n35077;
  assign n35079 = n7714 & ~n35078;
  assign n35080 = ~n35033 & ~n35079;
  assign n35081 = ~n7705 & ~n35080;
  assign n35082 = ~n9898 & ~n35081;
  assign n35083 = ~n7808 & ~n35082;
  assign n35084 = ~n33311 & ~n35027;
  assign n35085 = n7728 & ~n35084;
  assign n35086 = ~n35063 & ~n35085;
  assign n35087 = ~n7723 & ~n35086;
  assign n35088 = ~n32941 & ~n35087;
  assign n35089 = ~n7714 & ~n35088;
  assign n35090 = ~n32940 & ~n35089;
  assign n35091 = ~n7705 & ~n35090;
  assign n35092 = ~n22399 & ~n35091;
  assign n35093 = n7808 & ~n35092;
  assign n35094 = ~n35083 & ~n35093;
  assign n35095 = ~n8195 & ~n35094;
  assign n35096 = ~n11685 & ~n33339;
  assign n35097 = i_hlock7 & ~n35096;
  assign n35098 = ~n11685 & ~n33357;
  assign n35099 = ~i_hlock7 & ~n35098;
  assign n35100 = ~n35097 & ~n35099;
  assign n35101 = i_hbusreq7 & ~n35100;
  assign n35102 = ~n11696 & ~n33392;
  assign n35103 = i_hlock7 & ~n35102;
  assign n35104 = ~n11696 & ~n33425;
  assign n35105 = ~i_hlock7 & ~n35104;
  assign n35106 = ~n35103 & ~n35105;
  assign n35107 = ~i_hbusreq7 & ~n35106;
  assign n35108 = ~n35101 & ~n35107;
  assign n35109 = n7924 & ~n35108;
  assign n35110 = ~n10375 & ~n35109;
  assign n35111 = n8214 & ~n35110;
  assign n35112 = n8214 & ~n35111;
  assign n35113 = n8202 & ~n35112;
  assign n35114 = ~n10332 & ~n35113;
  assign n35115 = n7728 & ~n35114;
  assign n35116 = n8214 & ~n35026;
  assign n35117 = ~n8336 & ~n35116;
  assign n35118 = n8202 & ~n35117;
  assign n35119 = ~n10649 & ~n35118;
  assign n35120 = ~n7728 & ~n35119;
  assign n35121 = ~n35115 & ~n35120;
  assign n35122 = ~n7723 & ~n35121;
  assign n35123 = ~n7723 & ~n35122;
  assign n35124 = ~n7714 & ~n35123;
  assign n35125 = ~n7714 & ~n35124;
  assign n35126 = n7705 & ~n35125;
  assign n35127 = n7723 & ~n35119;
  assign n35128 = n7920 & ~n35119;
  assign n35129 = ~n35027 & ~n35128;
  assign n35130 = ~n7723 & ~n35129;
  assign n35131 = ~n35127 & ~n35130;
  assign n35132 = n7714 & ~n35131;
  assign n35133 = ~n35033 & ~n35132;
  assign n35134 = ~n7705 & ~n35133;
  assign n35135 = ~n35126 & ~n35134;
  assign n35136 = ~n7808 & ~n35135;
  assign n35137 = ~n7920 & ~n35114;
  assign n35138 = ~n33743 & ~n35137;
  assign n35139 = n7728 & ~n35138;
  assign n35140 = ~n7920 & ~n35119;
  assign n35141 = ~n33753 & ~n35140;
  assign n35142 = ~n7728 & ~n35141;
  assign n35143 = ~n35139 & ~n35142;
  assign n35144 = ~n7723 & ~n35143;
  assign n35145 = ~n7723 & ~n35144;
  assign n35146 = ~n7714 & ~n35145;
  assign n35147 = ~n7714 & ~n35146;
  assign n35148 = n7705 & ~n35147;
  assign n35149 = ~n33844 & ~n35140;
  assign n35150 = n7728 & ~n35149;
  assign n35151 = ~n34146 & ~n35140;
  assign n35152 = ~n7728 & ~n35151;
  assign n35153 = ~n35150 & ~n35152;
  assign n35154 = n7723 & ~n35153;
  assign n35155 = ~n7723 & ~n35151;
  assign n35156 = ~n35154 & ~n35155;
  assign n35157 = n7714 & ~n35156;
  assign n35158 = n7723 & ~n35151;
  assign n35159 = ~n34634 & ~n35027;
  assign n35160 = n7728 & ~n35159;
  assign n35161 = ~n35063 & ~n35160;
  assign n35162 = ~n7723 & ~n35161;
  assign n35163 = ~n35158 & ~n35162;
  assign n35164 = ~n7714 & ~n35163;
  assign n35165 = ~n35157 & ~n35164;
  assign n35166 = ~n7705 & ~n35165;
  assign n35167 = ~n35148 & ~n35166;
  assign n35168 = n7808 & ~n35167;
  assign n35169 = ~n35136 & ~n35168;
  assign n35170 = n8195 & ~n35169;
  assign n35171 = ~n35095 & ~n35170;
  assign n35172 = n8193 & ~n35171;
  assign n35173 = ~n35075 & ~n35172;
  assign n35174 = ~n8191 & ~n35173;
  assign n35175 = ~n35000 & ~n35174;
  assign n35176 = ~n8188 & ~n35175;
  assign n35177 = ~n34826 & ~n35176;
  assign n35178 = ~n8185 & ~n35177;
  assign n35179 = ~n28594 & ~n35178;
  assign n35180 = ~controllable_hgrant8 & ~n35179;
  assign n35181 = ~n12606 & ~n35180;
  assign n35182 = controllable_nhgrant0 & ~n35181;
  assign n35183 = ~n26632 & ~n35182;
  assign n35184 = controllable_hgrant7 & ~n35183;
  assign n35185 = ~controllable_hmaster2 & ~n26640;
  assign n35186 = ~controllable_hmaster2 & ~n35185;
  assign n35187 = ~controllable_hmaster1 & ~n35186;
  assign n35188 = ~controllable_hmaster1 & ~n35187;
  assign n35189 = ~controllable_hgrant6 & ~n35188;
  assign n35190 = ~n16722 & ~n35189;
  assign n35191 = ~controllable_hmaster0 & ~n35190;
  assign n35192 = ~controllable_hmaster0 & ~n35191;
  assign n35193 = i_hlock8 & ~n35192;
  assign n35194 = ~controllable_hmaster2 & ~n26655;
  assign n35195 = ~controllable_hmaster2 & ~n35194;
  assign n35196 = ~controllable_hmaster1 & ~n35195;
  assign n35197 = ~controllable_hmaster1 & ~n35196;
  assign n35198 = ~controllable_hgrant6 & ~n35197;
  assign n35199 = ~n16754 & ~n35198;
  assign n35200 = ~controllable_hmaster0 & ~n35199;
  assign n35201 = ~controllable_hmaster0 & ~n35200;
  assign n35202 = ~i_hlock8 & ~n35201;
  assign n35203 = ~n35193 & ~n35202;
  assign n35204 = controllable_hmaster3 & ~n35203;
  assign n35205 = controllable_hmaster3 & ~n35204;
  assign n35206 = i_hbusreq7 & ~n35205;
  assign n35207 = i_hbusreq8 & ~n35203;
  assign n35208 = i_hbusreq6 & ~n35188;
  assign n35209 = ~controllable_hmaster2 & ~n26683;
  assign n35210 = ~controllable_hmaster2 & ~n35209;
  assign n35211 = ~controllable_hmaster1 & ~n35210;
  assign n35212 = ~controllable_hmaster1 & ~n35211;
  assign n35213 = ~i_hbusreq6 & ~n35212;
  assign n35214 = ~n35208 & ~n35213;
  assign n35215 = ~controllable_hgrant6 & ~n35214;
  assign n35216 = ~n16778 & ~n35215;
  assign n35217 = ~controllable_hmaster0 & ~n35216;
  assign n35218 = ~controllable_hmaster0 & ~n35217;
  assign n35219 = i_hlock8 & ~n35218;
  assign n35220 = i_hbusreq6 & ~n35197;
  assign n35221 = ~controllable_hmaster2 & ~n26713;
  assign n35222 = ~controllable_hmaster2 & ~n35221;
  assign n35223 = ~controllable_hmaster1 & ~n35222;
  assign n35224 = ~controllable_hmaster1 & ~n35223;
  assign n35225 = ~i_hbusreq6 & ~n35224;
  assign n35226 = ~n35220 & ~n35225;
  assign n35227 = ~controllable_hgrant6 & ~n35226;
  assign n35228 = ~n16848 & ~n35227;
  assign n35229 = ~controllable_hmaster0 & ~n35228;
  assign n35230 = ~controllable_hmaster0 & ~n35229;
  assign n35231 = ~i_hlock8 & ~n35230;
  assign n35232 = ~n35219 & ~n35231;
  assign n35233 = ~i_hbusreq8 & ~n35232;
  assign n35234 = ~n35207 & ~n35233;
  assign n35235 = controllable_hmaster3 & ~n35234;
  assign n35236 = controllable_hmaster3 & ~n35235;
  assign n35237 = ~i_hbusreq7 & ~n35236;
  assign n35238 = ~n35206 & ~n35237;
  assign n35239 = ~n7924 & ~n35238;
  assign n35240 = controllable_hmaster0 & ~n12829;
  assign n35241 = ~controllable_hmaster2 & ~n26737;
  assign n35242 = ~n12798 & ~n35241;
  assign n35243 = ~controllable_hmaster1 & ~n35242;
  assign n35244 = ~n12797 & ~n35243;
  assign n35245 = ~controllable_hgrant6 & ~n35244;
  assign n35246 = ~n16722 & ~n35245;
  assign n35247 = ~controllable_hmaster0 & ~n35246;
  assign n35248 = ~n35240 & ~n35247;
  assign n35249 = i_hlock8 & ~n35248;
  assign n35250 = ~controllable_hmaster2 & ~n26753;
  assign n35251 = ~n12798 & ~n35250;
  assign n35252 = ~controllable_hmaster1 & ~n35251;
  assign n35253 = ~n12797 & ~n35252;
  assign n35254 = ~controllable_hgrant6 & ~n35253;
  assign n35255 = ~n16754 & ~n35254;
  assign n35256 = ~controllable_hmaster0 & ~n35255;
  assign n35257 = ~n35240 & ~n35256;
  assign n35258 = ~i_hlock8 & ~n35257;
  assign n35259 = ~n35249 & ~n35258;
  assign n35260 = controllable_hmaster3 & ~n35259;
  assign n35261 = ~n12833 & ~n35260;
  assign n35262 = i_hbusreq7 & ~n35261;
  assign n35263 = i_hbusreq8 & ~n35259;
  assign n35264 = controllable_hmaster0 & ~n12955;
  assign n35265 = i_hbusreq6 & ~n35244;
  assign n35266 = ~controllable_hmaster2 & ~n26782;
  assign n35267 = ~n12877 & ~n35266;
  assign n35268 = ~controllable_hmaster1 & ~n35267;
  assign n35269 = ~n12876 & ~n35268;
  assign n35270 = ~i_hbusreq6 & ~n35269;
  assign n35271 = ~n35265 & ~n35270;
  assign n35272 = ~controllable_hgrant6 & ~n35271;
  assign n35273 = ~n16778 & ~n35272;
  assign n35274 = ~controllable_hmaster0 & ~n35273;
  assign n35275 = ~n35264 & ~n35274;
  assign n35276 = i_hlock8 & ~n35275;
  assign n35277 = i_hbusreq6 & ~n35253;
  assign n35278 = ~controllable_hmaster2 & ~n26813;
  assign n35279 = ~n12877 & ~n35278;
  assign n35280 = ~controllable_hmaster1 & ~n35279;
  assign n35281 = ~n12876 & ~n35280;
  assign n35282 = ~i_hbusreq6 & ~n35281;
  assign n35283 = ~n35277 & ~n35282;
  assign n35284 = ~controllable_hgrant6 & ~n35283;
  assign n35285 = ~n16848 & ~n35284;
  assign n35286 = ~controllable_hmaster0 & ~n35285;
  assign n35287 = ~n35264 & ~n35286;
  assign n35288 = ~i_hlock8 & ~n35287;
  assign n35289 = ~n35276 & ~n35288;
  assign n35290 = ~i_hbusreq8 & ~n35289;
  assign n35291 = ~n35263 & ~n35290;
  assign n35292 = controllable_hmaster3 & ~n35291;
  assign n35293 = ~n12964 & ~n35292;
  assign n35294 = ~i_hbusreq7 & ~n35293;
  assign n35295 = ~n35262 & ~n35294;
  assign n35296 = n7924 & ~n35295;
  assign n35297 = ~n35239 & ~n35296;
  assign n35298 = n8214 & ~n35297;
  assign n35299 = ~n8725 & ~n35298;
  assign n35300 = ~n8202 & ~n35299;
  assign n35301 = ~n8872 & ~n35300;
  assign n35302 = n7920 & ~n35301;
  assign n35303 = ~n8651 & ~n35302;
  assign n35304 = n7728 & ~n35303;
  assign n35305 = ~n7739 & ~n35185;
  assign n35306 = ~controllable_hmaster1 & ~n35305;
  assign n35307 = ~n7738 & ~n35306;
  assign n35308 = ~controllable_hgrant6 & ~n35307;
  assign n35309 = ~n17225 & ~n35308;
  assign n35310 = ~controllable_hmaster0 & ~n35309;
  assign n35311 = ~n8904 & ~n35310;
  assign n35312 = i_hlock8 & ~n35311;
  assign n35313 = ~n7739 & ~n35194;
  assign n35314 = ~controllable_hmaster1 & ~n35313;
  assign n35315 = ~n7738 & ~n35314;
  assign n35316 = ~controllable_hgrant6 & ~n35315;
  assign n35317 = ~n17234 & ~n35316;
  assign n35318 = ~controllable_hmaster0 & ~n35317;
  assign n35319 = ~n8904 & ~n35318;
  assign n35320 = ~i_hlock8 & ~n35319;
  assign n35321 = ~n35312 & ~n35320;
  assign n35322 = controllable_hmaster3 & ~n35321;
  assign n35323 = controllable_hmaster3 & ~n35322;
  assign n35324 = i_hbusreq7 & ~n35323;
  assign n35325 = i_hbusreq8 & ~n35321;
  assign n35326 = i_hbusreq6 & ~n35307;
  assign n35327 = ~n7771 & ~n35209;
  assign n35328 = ~controllable_hmaster1 & ~n35327;
  assign n35329 = ~n7770 & ~n35328;
  assign n35330 = ~i_hbusreq6 & ~n35329;
  assign n35331 = ~n35326 & ~n35330;
  assign n35332 = ~controllable_hgrant6 & ~n35331;
  assign n35333 = ~n17248 & ~n35332;
  assign n35334 = ~controllable_hmaster0 & ~n35333;
  assign n35335 = ~n8922 & ~n35334;
  assign n35336 = i_hlock8 & ~n35335;
  assign n35337 = i_hbusreq6 & ~n35315;
  assign n35338 = ~n7771 & ~n35221;
  assign n35339 = ~controllable_hmaster1 & ~n35338;
  assign n35340 = ~n7770 & ~n35339;
  assign n35341 = ~i_hbusreq6 & ~n35340;
  assign n35342 = ~n35337 & ~n35341;
  assign n35343 = ~controllable_hgrant6 & ~n35342;
  assign n35344 = ~n17260 & ~n35343;
  assign n35345 = ~controllable_hmaster0 & ~n35344;
  assign n35346 = ~n8922 & ~n35345;
  assign n35347 = ~i_hlock8 & ~n35346;
  assign n35348 = ~n35336 & ~n35347;
  assign n35349 = ~i_hbusreq8 & ~n35348;
  assign n35350 = ~n35325 & ~n35349;
  assign n35351 = controllable_hmaster3 & ~n35350;
  assign n35352 = controllable_hmaster3 & ~n35351;
  assign n35353 = ~i_hbusreq7 & ~n35352;
  assign n35354 = ~n35324 & ~n35353;
  assign n35355 = ~n7924 & ~n35354;
  assign n35356 = controllable_hmaster0 & ~n13037;
  assign n35357 = ~n13025 & ~n35241;
  assign n35358 = ~controllable_hmaster1 & ~n35357;
  assign n35359 = ~n13024 & ~n35358;
  assign n35360 = ~controllable_hgrant6 & ~n35359;
  assign n35361 = ~n17225 & ~n35360;
  assign n35362 = ~controllable_hmaster0 & ~n35361;
  assign n35363 = ~n35356 & ~n35362;
  assign n35364 = i_hlock8 & ~n35363;
  assign n35365 = ~n13025 & ~n35250;
  assign n35366 = ~controllable_hmaster1 & ~n35365;
  assign n35367 = ~n13024 & ~n35366;
  assign n35368 = ~controllable_hgrant6 & ~n35367;
  assign n35369 = ~n17234 & ~n35368;
  assign n35370 = ~controllable_hmaster0 & ~n35369;
  assign n35371 = ~n35356 & ~n35370;
  assign n35372 = ~i_hlock8 & ~n35371;
  assign n35373 = ~n35364 & ~n35372;
  assign n35374 = controllable_hmaster3 & ~n35373;
  assign n35375 = ~n12833 & ~n35374;
  assign n35376 = i_hbusreq7 & ~n35375;
  assign n35377 = i_hbusreq8 & ~n35373;
  assign n35378 = controllable_hmaster0 & ~n13098;
  assign n35379 = i_hbusreq6 & ~n35359;
  assign n35380 = ~n13081 & ~n35266;
  assign n35381 = ~controllable_hmaster1 & ~n35380;
  assign n35382 = ~n13080 & ~n35381;
  assign n35383 = ~i_hbusreq6 & ~n35382;
  assign n35384 = ~n35379 & ~n35383;
  assign n35385 = ~controllable_hgrant6 & ~n35384;
  assign n35386 = ~n17248 & ~n35385;
  assign n35387 = ~controllable_hmaster0 & ~n35386;
  assign n35388 = ~n35378 & ~n35387;
  assign n35389 = i_hlock8 & ~n35388;
  assign n35390 = i_hbusreq6 & ~n35367;
  assign n35391 = ~n13081 & ~n35278;
  assign n35392 = ~controllable_hmaster1 & ~n35391;
  assign n35393 = ~n13080 & ~n35392;
  assign n35394 = ~i_hbusreq6 & ~n35393;
  assign n35395 = ~n35390 & ~n35394;
  assign n35396 = ~controllable_hgrant6 & ~n35395;
  assign n35397 = ~n17260 & ~n35396;
  assign n35398 = ~controllable_hmaster0 & ~n35397;
  assign n35399 = ~n35378 & ~n35398;
  assign n35400 = ~i_hlock8 & ~n35399;
  assign n35401 = ~n35389 & ~n35400;
  assign n35402 = ~i_hbusreq8 & ~n35401;
  assign n35403 = ~n35377 & ~n35402;
  assign n35404 = controllable_hmaster3 & ~n35403;
  assign n35405 = ~n12964 & ~n35404;
  assign n35406 = ~i_hbusreq7 & ~n35405;
  assign n35407 = ~n35376 & ~n35406;
  assign n35408 = n7924 & ~n35407;
  assign n35409 = ~n35355 & ~n35408;
  assign n35410 = n8214 & ~n35409;
  assign n35411 = ~n8903 & ~n35410;
  assign n35412 = ~n8202 & ~n35411;
  assign n35413 = ~n8972 & ~n35412;
  assign n35414 = n7920 & ~n35413;
  assign n35415 = ~n8877 & ~n35414;
  assign n35416 = ~n7728 & ~n35415;
  assign n35417 = ~n35304 & ~n35416;
  assign n35418 = ~n7723 & ~n35417;
  assign n35419 = ~n7723 & ~n35418;
  assign n35420 = ~n7714 & ~n35419;
  assign n35421 = ~n7714 & ~n35420;
  assign n35422 = n7705 & ~n35421;
  assign n35423 = ~controllable_hmaster0 & ~n13327;
  assign n35424 = ~n8986 & ~n35423;
  assign n35425 = controllable_hmaster3 & ~n35424;
  assign n35426 = ~n8995 & ~n35425;
  assign n35427 = i_hbusreq7 & ~n35426;
  assign n35428 = i_hbusreq8 & ~n35424;
  assign n35429 = ~controllable_hmaster0 & ~n13376;
  assign n35430 = ~n9005 & ~n35429;
  assign n35431 = ~i_hbusreq8 & ~n35430;
  assign n35432 = ~n35428 & ~n35431;
  assign n35433 = controllable_hmaster3 & ~n35432;
  assign n35434 = ~n9041 & ~n35433;
  assign n35435 = ~i_hbusreq7 & ~n35434;
  assign n35436 = ~n35427 & ~n35435;
  assign n35437 = ~n7924 & ~n35436;
  assign n35438 = ~controllable_hmaster0 & ~n13404;
  assign n35439 = ~n26931 & ~n35438;
  assign n35440 = controllable_hmaster3 & ~n35439;
  assign n35441 = ~n13201 & ~n35440;
  assign n35442 = i_hbusreq7 & ~n35441;
  assign n35443 = i_hbusreq8 & ~n35439;
  assign n35444 = ~controllable_hmaster0 & ~n13518;
  assign n35445 = ~n26971 & ~n35444;
  assign n35446 = ~i_hbusreq8 & ~n35445;
  assign n35447 = ~n35443 & ~n35446;
  assign n35448 = controllable_hmaster3 & ~n35447;
  assign n35449 = ~n13641 & ~n35448;
  assign n35450 = ~i_hbusreq7 & ~n35449;
  assign n35451 = ~n35442 & ~n35450;
  assign n35452 = n7924 & ~n35451;
  assign n35453 = ~n35437 & ~n35452;
  assign n35454 = ~n8214 & ~n35453;
  assign n35455 = ~n8358 & ~n35185;
  assign n35456 = ~controllable_hmaster1 & ~n35455;
  assign n35457 = ~n8357 & ~n35456;
  assign n35458 = ~controllable_hgrant6 & ~n35457;
  assign n35459 = ~n13406 & ~n35458;
  assign n35460 = ~controllable_hmaster0 & ~n35459;
  assign n35461 = ~n9046 & ~n35460;
  assign n35462 = i_hlock8 & ~n35461;
  assign n35463 = ~n8358 & ~n35194;
  assign n35464 = ~controllable_hmaster1 & ~n35463;
  assign n35465 = ~n8357 & ~n35464;
  assign n35466 = ~controllable_hgrant6 & ~n35465;
  assign n35467 = ~n13427 & ~n35466;
  assign n35468 = ~controllable_hmaster0 & ~n35467;
  assign n35469 = ~n9046 & ~n35468;
  assign n35470 = ~i_hlock8 & ~n35469;
  assign n35471 = ~n35462 & ~n35470;
  assign n35472 = controllable_hmaster3 & ~n35471;
  assign n35473 = ~n8995 & ~n35472;
  assign n35474 = i_hbusreq7 & ~n35473;
  assign n35475 = i_hbusreq8 & ~n35471;
  assign n35476 = i_hbusreq6 & ~n35457;
  assign n35477 = ~n8484 & ~n35209;
  assign n35478 = ~controllable_hmaster1 & ~n35477;
  assign n35479 = ~n8483 & ~n35478;
  assign n35480 = ~i_hbusreq6 & ~n35479;
  assign n35481 = ~n35476 & ~n35480;
  assign n35482 = ~controllable_hgrant6 & ~n35481;
  assign n35483 = ~n13520 & ~n35482;
  assign n35484 = ~controllable_hmaster0 & ~n35483;
  assign n35485 = ~n9064 & ~n35484;
  assign n35486 = i_hlock8 & ~n35485;
  assign n35487 = i_hbusreq6 & ~n35465;
  assign n35488 = ~n8484 & ~n35221;
  assign n35489 = ~controllable_hmaster1 & ~n35488;
  assign n35490 = ~n8483 & ~n35489;
  assign n35491 = ~i_hbusreq6 & ~n35490;
  assign n35492 = ~n35487 & ~n35491;
  assign n35493 = ~controllable_hgrant6 & ~n35492;
  assign n35494 = ~n13573 & ~n35493;
  assign n35495 = ~controllable_hmaster0 & ~n35494;
  assign n35496 = ~n9064 & ~n35495;
  assign n35497 = ~i_hlock8 & ~n35496;
  assign n35498 = ~n35486 & ~n35497;
  assign n35499 = ~i_hbusreq8 & ~n35498;
  assign n35500 = ~n35475 & ~n35499;
  assign n35501 = controllable_hmaster3 & ~n35500;
  assign n35502 = ~n9041 & ~n35501;
  assign n35503 = ~i_hbusreq7 & ~n35502;
  assign n35504 = ~n35474 & ~n35503;
  assign n35505 = ~n7924 & ~n35504;
  assign n35506 = ~n13168 & ~n35241;
  assign n35507 = ~controllable_hmaster1 & ~n35506;
  assign n35508 = ~n13167 & ~n35507;
  assign n35509 = ~controllable_hgrant6 & ~n35508;
  assign n35510 = ~n13406 & ~n35509;
  assign n35511 = ~controllable_hmaster0 & ~n35510;
  assign n35512 = ~n27003 & ~n35511;
  assign n35513 = i_hlock8 & ~n35512;
  assign n35514 = ~n13168 & ~n35250;
  assign n35515 = ~controllable_hmaster1 & ~n35514;
  assign n35516 = ~n13167 & ~n35515;
  assign n35517 = ~controllable_hgrant6 & ~n35516;
  assign n35518 = ~n13427 & ~n35517;
  assign n35519 = ~controllable_hmaster0 & ~n35518;
  assign n35520 = ~n27003 & ~n35519;
  assign n35521 = ~i_hlock8 & ~n35520;
  assign n35522 = ~n35513 & ~n35521;
  assign n35523 = controllable_hmaster3 & ~n35522;
  assign n35524 = ~n13201 & ~n35523;
  assign n35525 = i_hbusreq7 & ~n35524;
  assign n35526 = i_hbusreq8 & ~n35522;
  assign n35527 = controllable_hmaster0 & ~n13291;
  assign n35528 = i_hbusreq6 & ~n35508;
  assign n35529 = ~n13245 & ~n35266;
  assign n35530 = ~controllable_hmaster1 & ~n35529;
  assign n35531 = ~n13244 & ~n35530;
  assign n35532 = ~i_hbusreq6 & ~n35531;
  assign n35533 = ~n35528 & ~n35532;
  assign n35534 = ~controllable_hgrant6 & ~n35533;
  assign n35535 = ~n13520 & ~n35534;
  assign n35536 = ~controllable_hmaster0 & ~n35535;
  assign n35537 = ~n35527 & ~n35536;
  assign n35538 = i_hlock8 & ~n35537;
  assign n35539 = i_hbusreq6 & ~n35516;
  assign n35540 = ~n13245 & ~n35278;
  assign n35541 = ~controllable_hmaster1 & ~n35540;
  assign n35542 = ~n13244 & ~n35541;
  assign n35543 = ~i_hbusreq6 & ~n35542;
  assign n35544 = ~n35539 & ~n35543;
  assign n35545 = ~controllable_hgrant6 & ~n35544;
  assign n35546 = ~n13573 & ~n35545;
  assign n35547 = ~controllable_hmaster0 & ~n35546;
  assign n35548 = ~n35527 & ~n35547;
  assign n35549 = ~i_hlock8 & ~n35548;
  assign n35550 = ~n35538 & ~n35549;
  assign n35551 = ~i_hbusreq8 & ~n35550;
  assign n35552 = ~n35526 & ~n35551;
  assign n35553 = controllable_hmaster3 & ~n35552;
  assign n35554 = ~n13306 & ~n35553;
  assign n35555 = ~i_hbusreq7 & ~n35554;
  assign n35556 = ~n35525 & ~n35555;
  assign n35557 = n7924 & ~n35556;
  assign n35558 = ~n35505 & ~n35557;
  assign n35559 = n8214 & ~n35558;
  assign n35560 = ~n35454 & ~n35559;
  assign n35561 = ~n8202 & ~n35560;
  assign n35562 = ~n9046 & ~n35423;
  assign n35563 = controllable_hmaster3 & ~n35562;
  assign n35564 = ~n9101 & ~n35563;
  assign n35565 = i_hlock7 & ~n35564;
  assign n35566 = ~n9109 & ~n35563;
  assign n35567 = ~i_hlock7 & ~n35566;
  assign n35568 = ~n35565 & ~n35567;
  assign n35569 = i_hbusreq7 & ~n35568;
  assign n35570 = i_hbusreq8 & ~n35562;
  assign n35571 = ~n9064 & ~n35429;
  assign n35572 = ~i_hbusreq8 & ~n35571;
  assign n35573 = ~n35570 & ~n35572;
  assign n35574 = controllable_hmaster3 & ~n35573;
  assign n35575 = ~n9131 & ~n35574;
  assign n35576 = i_hlock7 & ~n35575;
  assign n35577 = ~n9145 & ~n35574;
  assign n35578 = ~i_hlock7 & ~n35577;
  assign n35579 = ~n35576 & ~n35578;
  assign n35580 = ~i_hbusreq7 & ~n35579;
  assign n35581 = ~n35569 & ~n35580;
  assign n35582 = ~n7924 & ~n35581;
  assign n35583 = ~n27003 & ~n35438;
  assign n35584 = controllable_hmaster3 & ~n35583;
  assign n35585 = ~n13684 & ~n35584;
  assign n35586 = i_hlock7 & ~n35585;
  assign n35587 = ~n13696 & ~n35584;
  assign n35588 = ~i_hlock7 & ~n35587;
  assign n35589 = ~n35586 & ~n35588;
  assign n35590 = i_hbusreq7 & ~n35589;
  assign n35591 = i_hbusreq8 & ~n35583;
  assign n35592 = ~n27013 & ~n35444;
  assign n35593 = ~i_hbusreq8 & ~n35592;
  assign n35594 = ~n35591 & ~n35593;
  assign n35595 = controllable_hmaster3 & ~n35594;
  assign n35596 = ~n13732 & ~n35595;
  assign n35597 = i_hlock7 & ~n35596;
  assign n35598 = ~n13750 & ~n35595;
  assign n35599 = ~i_hlock7 & ~n35598;
  assign n35600 = ~n35597 & ~n35599;
  assign n35601 = ~i_hbusreq7 & ~n35600;
  assign n35602 = ~n35590 & ~n35601;
  assign n35603 = n7924 & ~n35602;
  assign n35604 = ~n35582 & ~n35603;
  assign n35605 = ~n8214 & ~n35604;
  assign n35606 = ~n9158 & ~n35563;
  assign n35607 = i_hbusreq7 & ~n35606;
  assign n35608 = ~n9173 & ~n35574;
  assign n35609 = ~i_hbusreq7 & ~n35608;
  assign n35610 = ~n35607 & ~n35609;
  assign n35611 = ~n7924 & ~n35610;
  assign n35612 = ~n13774 & ~n35584;
  assign n35613 = i_hbusreq7 & ~n35612;
  assign n35614 = ~n13792 & ~n35595;
  assign n35615 = ~i_hbusreq7 & ~n35614;
  assign n35616 = ~n35613 & ~n35615;
  assign n35617 = n7924 & ~n35616;
  assign n35618 = ~n35611 & ~n35617;
  assign n35619 = n8214 & ~n35618;
  assign n35620 = ~n35605 & ~n35619;
  assign n35621 = n8202 & ~n35620;
  assign n35622 = ~n35561 & ~n35621;
  assign n35623 = n7920 & ~n35622;
  assign n35624 = ~n8877 & ~n35623;
  assign n35625 = n7728 & ~n35624;
  assign n35626 = ~n8986 & ~n35460;
  assign n35627 = i_hlock8 & ~n35626;
  assign n35628 = ~n8986 & ~n35468;
  assign n35629 = ~i_hlock8 & ~n35628;
  assign n35630 = ~n35627 & ~n35629;
  assign n35631 = controllable_hmaster3 & ~n35630;
  assign n35632 = ~n9235 & ~n35631;
  assign n35633 = i_hlock7 & ~n35632;
  assign n35634 = ~n9243 & ~n35631;
  assign n35635 = ~i_hlock7 & ~n35634;
  assign n35636 = ~n35633 & ~n35635;
  assign n35637 = i_hbusreq7 & ~n35636;
  assign n35638 = i_hbusreq8 & ~n35630;
  assign n35639 = ~controllable_hmaster2 & ~n27225;
  assign n35640 = ~n9260 & ~n35639;
  assign n35641 = ~controllable_hmaster1 & ~n35640;
  assign n35642 = ~n9259 & ~n35641;
  assign n35643 = ~i_hbusreq6 & ~n35642;
  assign n35644 = ~n35476 & ~n35643;
  assign n35645 = ~controllable_hgrant6 & ~n35644;
  assign n35646 = ~n14019 & ~n35645;
  assign n35647 = ~controllable_hmaster0 & ~n35646;
  assign n35648 = ~n9266 & ~n35647;
  assign n35649 = i_hlock8 & ~n35648;
  assign n35650 = ~controllable_hmaster2 & ~n27252;
  assign n35651 = ~n9260 & ~n35650;
  assign n35652 = ~controllable_hmaster1 & ~n35651;
  assign n35653 = ~n9259 & ~n35652;
  assign n35654 = ~i_hbusreq6 & ~n35653;
  assign n35655 = ~n35487 & ~n35654;
  assign n35656 = ~controllable_hgrant6 & ~n35655;
  assign n35657 = ~n14054 & ~n35656;
  assign n35658 = ~controllable_hmaster0 & ~n35657;
  assign n35659 = ~n9266 & ~n35658;
  assign n35660 = ~i_hlock8 & ~n35659;
  assign n35661 = ~n35649 & ~n35660;
  assign n35662 = ~i_hbusreq8 & ~n35661;
  assign n35663 = ~n35638 & ~n35662;
  assign n35664 = controllable_hmaster3 & ~n35663;
  assign n35665 = ~n9443 & ~n35664;
  assign n35666 = i_hlock7 & ~n35665;
  assign n35667 = ~n9457 & ~n35664;
  assign n35668 = ~i_hlock7 & ~n35667;
  assign n35669 = ~n35666 & ~n35668;
  assign n35670 = ~i_hbusreq7 & ~n35669;
  assign n35671 = ~n35637 & ~n35670;
  assign n35672 = ~n7924 & ~n35671;
  assign n35673 = ~n26931 & ~n35511;
  assign n35674 = i_hlock8 & ~n35673;
  assign n35675 = ~n26931 & ~n35519;
  assign n35676 = ~i_hlock8 & ~n35675;
  assign n35677 = ~n35674 & ~n35676;
  assign n35678 = controllable_hmaster3 & ~n35677;
  assign n35679 = ~n13948 & ~n35678;
  assign n35680 = i_hlock7 & ~n35679;
  assign n35681 = ~n13959 & ~n35678;
  assign n35682 = ~i_hlock7 & ~n35681;
  assign n35683 = ~n35680 & ~n35682;
  assign n35684 = i_hbusreq7 & ~n35683;
  assign n35685 = i_hbusreq8 & ~n35677;
  assign n35686 = ~controllable_hmaster2 & ~n27342;
  assign n35687 = ~n14401 & ~n35686;
  assign n35688 = ~controllable_hmaster1 & ~n35687;
  assign n35689 = ~n14400 & ~n35688;
  assign n35690 = ~i_hbusreq6 & ~n35689;
  assign n35691 = ~n35528 & ~n35690;
  assign n35692 = ~controllable_hgrant6 & ~n35691;
  assign n35693 = ~n14019 & ~n35692;
  assign n35694 = ~controllable_hmaster0 & ~n35693;
  assign n35695 = ~n27322 & ~n35694;
  assign n35696 = i_hlock8 & ~n35695;
  assign n35697 = ~controllable_hmaster2 & ~n27369;
  assign n35698 = ~n14401 & ~n35697;
  assign n35699 = ~controllable_hmaster1 & ~n35698;
  assign n35700 = ~n14400 & ~n35699;
  assign n35701 = ~i_hbusreq6 & ~n35700;
  assign n35702 = ~n35539 & ~n35701;
  assign n35703 = ~controllable_hgrant6 & ~n35702;
  assign n35704 = ~n14054 & ~n35703;
  assign n35705 = ~controllable_hmaster0 & ~n35704;
  assign n35706 = ~n27322 & ~n35705;
  assign n35707 = ~i_hlock8 & ~n35706;
  assign n35708 = ~n35696 & ~n35707;
  assign n35709 = ~i_hbusreq8 & ~n35708;
  assign n35710 = ~n35685 & ~n35709;
  assign n35711 = controllable_hmaster3 & ~n35710;
  assign n35712 = ~n14689 & ~n35711;
  assign n35713 = i_hlock7 & ~n35712;
  assign n35714 = ~n14703 & ~n35711;
  assign n35715 = ~i_hlock7 & ~n35714;
  assign n35716 = ~n35713 & ~n35715;
  assign n35717 = ~i_hbusreq7 & ~n35716;
  assign n35718 = ~n35684 & ~n35717;
  assign n35719 = n7924 & ~n35718;
  assign n35720 = ~n35672 & ~n35719;
  assign n35721 = ~n8214 & ~n35720;
  assign n35722 = ~n9260 & ~n35209;
  assign n35723 = ~controllable_hmaster1 & ~n35722;
  assign n35724 = ~n9259 & ~n35723;
  assign n35725 = ~i_hbusreq6 & ~n35724;
  assign n35726 = ~n35476 & ~n35725;
  assign n35727 = ~controllable_hgrant6 & ~n35726;
  assign n35728 = ~n14443 & ~n35727;
  assign n35729 = ~controllable_hmaster0 & ~n35728;
  assign n35730 = ~n9479 & ~n35729;
  assign n35731 = i_hlock8 & ~n35730;
  assign n35732 = ~n9260 & ~n35221;
  assign n35733 = ~controllable_hmaster1 & ~n35732;
  assign n35734 = ~n9259 & ~n35733;
  assign n35735 = ~i_hbusreq6 & ~n35734;
  assign n35736 = ~n35487 & ~n35735;
  assign n35737 = ~controllable_hgrant6 & ~n35736;
  assign n35738 = ~n14484 & ~n35737;
  assign n35739 = ~controllable_hmaster0 & ~n35738;
  assign n35740 = ~n9479 & ~n35739;
  assign n35741 = ~i_hlock8 & ~n35740;
  assign n35742 = ~n35731 & ~n35741;
  assign n35743 = ~i_hbusreq8 & ~n35742;
  assign n35744 = ~n35638 & ~n35743;
  assign n35745 = controllable_hmaster3 & ~n35744;
  assign n35746 = ~n9443 & ~n35745;
  assign n35747 = i_hlock7 & ~n35746;
  assign n35748 = ~n9457 & ~n35745;
  assign n35749 = ~i_hlock7 & ~n35748;
  assign n35750 = ~n35747 & ~n35749;
  assign n35751 = ~i_hbusreq7 & ~n35750;
  assign n35752 = ~n35637 & ~n35751;
  assign n35753 = ~n7924 & ~n35752;
  assign n35754 = ~n14010 & ~n35266;
  assign n35755 = ~controllable_hmaster1 & ~n35754;
  assign n35756 = ~n14009 & ~n35755;
  assign n35757 = ~i_hbusreq6 & ~n35756;
  assign n35758 = ~n35528 & ~n35757;
  assign n35759 = ~controllable_hgrant6 & ~n35758;
  assign n35760 = ~n14443 & ~n35759;
  assign n35761 = ~controllable_hmaster0 & ~n35760;
  assign n35762 = ~n27494 & ~n35761;
  assign n35763 = i_hlock8 & ~n35762;
  assign n35764 = ~n14010 & ~n35278;
  assign n35765 = ~controllable_hmaster1 & ~n35764;
  assign n35766 = ~n14009 & ~n35765;
  assign n35767 = ~i_hbusreq6 & ~n35766;
  assign n35768 = ~n35539 & ~n35767;
  assign n35769 = ~controllable_hgrant6 & ~n35768;
  assign n35770 = ~n14484 & ~n35769;
  assign n35771 = ~controllable_hmaster0 & ~n35770;
  assign n35772 = ~n27494 & ~n35771;
  assign n35773 = ~i_hlock8 & ~n35772;
  assign n35774 = ~n35763 & ~n35773;
  assign n35775 = ~i_hbusreq8 & ~n35774;
  assign n35776 = ~n35685 & ~n35775;
  assign n35777 = controllable_hmaster3 & ~n35776;
  assign n35778 = ~n14294 & ~n35777;
  assign n35779 = i_hlock7 & ~n35778;
  assign n35780 = ~n14311 & ~n35777;
  assign n35781 = ~i_hlock7 & ~n35780;
  assign n35782 = ~n35779 & ~n35781;
  assign n35783 = ~i_hbusreq7 & ~n35782;
  assign n35784 = ~n35684 & ~n35783;
  assign n35785 = n7924 & ~n35784;
  assign n35786 = ~n35753 & ~n35785;
  assign n35787 = n8214 & ~n35786;
  assign n35788 = ~n35721 & ~n35787;
  assign n35789 = ~n8202 & ~n35788;
  assign n35790 = ~n9479 & ~n35647;
  assign n35791 = i_hlock8 & ~n35790;
  assign n35792 = ~n9479 & ~n35658;
  assign n35793 = ~i_hlock8 & ~n35792;
  assign n35794 = ~n35791 & ~n35793;
  assign n35795 = ~i_hbusreq8 & ~n35794;
  assign n35796 = ~n35638 & ~n35795;
  assign n35797 = controllable_hmaster3 & ~n35796;
  assign n35798 = ~n9527 & ~n35797;
  assign n35799 = i_hlock7 & ~n35798;
  assign n35800 = ~n9539 & ~n35797;
  assign n35801 = ~i_hlock7 & ~n35800;
  assign n35802 = ~n35799 & ~n35801;
  assign n35803 = ~i_hbusreq7 & ~n35802;
  assign n35804 = ~n35637 & ~n35803;
  assign n35805 = ~n7924 & ~n35804;
  assign n35806 = ~n27420 & ~n35694;
  assign n35807 = i_hlock8 & ~n35806;
  assign n35808 = ~n27420 & ~n35705;
  assign n35809 = ~i_hlock8 & ~n35808;
  assign n35810 = ~n35807 & ~n35809;
  assign n35811 = ~i_hbusreq8 & ~n35810;
  assign n35812 = ~n35685 & ~n35811;
  assign n35813 = controllable_hmaster3 & ~n35812;
  assign n35814 = ~n14769 & ~n35813;
  assign n35815 = i_hlock7 & ~n35814;
  assign n35816 = ~n14785 & ~n35813;
  assign n35817 = ~i_hlock7 & ~n35816;
  assign n35818 = ~n35815 & ~n35817;
  assign n35819 = ~i_hbusreq7 & ~n35818;
  assign n35820 = ~n35684 & ~n35819;
  assign n35821 = n7924 & ~n35820;
  assign n35822 = ~n35805 & ~n35821;
  assign n35823 = ~n8214 & ~n35822;
  assign n35824 = ~n9561 & ~n35797;
  assign n35825 = i_hlock7 & ~n35824;
  assign n35826 = ~n9567 & ~n35797;
  assign n35827 = ~i_hlock7 & ~n35826;
  assign n35828 = ~n35825 & ~n35827;
  assign n35829 = ~i_hbusreq7 & ~n35828;
  assign n35830 = ~n35637 & ~n35829;
  assign n35831 = ~n7924 & ~n35830;
  assign n35832 = ~n14820 & ~n35813;
  assign n35833 = i_hlock7 & ~n35832;
  assign n35834 = ~n14826 & ~n35813;
  assign n35835 = ~i_hlock7 & ~n35834;
  assign n35836 = ~n35833 & ~n35835;
  assign n35837 = ~i_hbusreq7 & ~n35836;
  assign n35838 = ~n35684 & ~n35837;
  assign n35839 = n7924 & ~n35838;
  assign n35840 = ~n35831 & ~n35839;
  assign n35841 = n8214 & ~n35840;
  assign n35842 = ~n35823 & ~n35841;
  assign n35843 = n8202 & ~n35842;
  assign n35844 = ~n35789 & ~n35843;
  assign n35845 = n7920 & ~n35844;
  assign n35846 = ~n8877 & ~n35845;
  assign n35847 = ~n7728 & ~n35846;
  assign n35848 = ~n35625 & ~n35847;
  assign n35849 = n7723 & ~n35848;
  assign n35850 = ~n7723 & ~n35846;
  assign n35851 = ~n35849 & ~n35850;
  assign n35852 = n7714 & ~n35851;
  assign n35853 = n7723 & ~n35846;
  assign n35854 = ~n8640 & ~n35845;
  assign n35855 = n7728 & ~n35854;
  assign n35856 = ~n9600 & ~n35209;
  assign n35857 = ~controllable_hmaster1 & ~n35856;
  assign n35858 = ~n9599 & ~n35857;
  assign n35859 = ~i_hbusreq6 & ~n35858;
  assign n35860 = ~n35476 & ~n35859;
  assign n35861 = ~controllable_hgrant6 & ~n35860;
  assign n35862 = ~n14927 & ~n35861;
  assign n35863 = ~controllable_hmaster0 & ~n35862;
  assign n35864 = ~n9606 & ~n35863;
  assign n35865 = i_hlock8 & ~n35864;
  assign n35866 = ~n9600 & ~n35221;
  assign n35867 = ~controllable_hmaster1 & ~n35866;
  assign n35868 = ~n9599 & ~n35867;
  assign n35869 = ~i_hbusreq6 & ~n35868;
  assign n35870 = ~n35487 & ~n35869;
  assign n35871 = ~controllable_hgrant6 & ~n35870;
  assign n35872 = ~n14960 & ~n35871;
  assign n35873 = ~controllable_hmaster0 & ~n35872;
  assign n35874 = ~n9606 & ~n35873;
  assign n35875 = ~i_hlock8 & ~n35874;
  assign n35876 = ~n35865 & ~n35875;
  assign n35877 = ~i_hbusreq8 & ~n35876;
  assign n35878 = ~n35638 & ~n35877;
  assign n35879 = controllable_hmaster3 & ~n35878;
  assign n35880 = ~n9720 & ~n35879;
  assign n35881 = i_hlock7 & ~n35880;
  assign n35882 = ~n9732 & ~n35879;
  assign n35883 = ~i_hlock7 & ~n35882;
  assign n35884 = ~n35881 & ~n35883;
  assign n35885 = ~i_hbusreq7 & ~n35884;
  assign n35886 = ~n35637 & ~n35885;
  assign n35887 = ~n7924 & ~n35886;
  assign n35888 = ~n14918 & ~n35266;
  assign n35889 = ~controllable_hmaster1 & ~n35888;
  assign n35890 = ~n14917 & ~n35889;
  assign n35891 = ~i_hbusreq6 & ~n35890;
  assign n35892 = ~n35528 & ~n35891;
  assign n35893 = ~controllable_hgrant6 & ~n35892;
  assign n35894 = ~n14927 & ~n35893;
  assign n35895 = ~controllable_hmaster0 & ~n35894;
  assign n35896 = ~n27646 & ~n35895;
  assign n35897 = i_hlock8 & ~n35896;
  assign n35898 = ~n14918 & ~n35278;
  assign n35899 = ~controllable_hmaster1 & ~n35898;
  assign n35900 = ~n14917 & ~n35899;
  assign n35901 = ~i_hbusreq6 & ~n35900;
  assign n35902 = ~n35539 & ~n35901;
  assign n35903 = ~controllable_hgrant6 & ~n35902;
  assign n35904 = ~n14960 & ~n35903;
  assign n35905 = ~controllable_hmaster0 & ~n35904;
  assign n35906 = ~n27646 & ~n35905;
  assign n35907 = ~i_hlock8 & ~n35906;
  assign n35908 = ~n35897 & ~n35907;
  assign n35909 = ~i_hbusreq8 & ~n35908;
  assign n35910 = ~n35685 & ~n35909;
  assign n35911 = controllable_hmaster3 & ~n35910;
  assign n35912 = ~n15149 & ~n35911;
  assign n35913 = i_hlock7 & ~n35912;
  assign n35914 = ~n15164 & ~n35911;
  assign n35915 = ~i_hlock7 & ~n35914;
  assign n35916 = ~n35913 & ~n35915;
  assign n35917 = ~i_hbusreq7 & ~n35916;
  assign n35918 = ~n35684 & ~n35917;
  assign n35919 = n7924 & ~n35918;
  assign n35920 = ~n35887 & ~n35919;
  assign n35921 = n7920 & ~n35920;
  assign n35922 = ~n8640 & ~n35921;
  assign n35923 = ~n7728 & ~n35922;
  assign n35924 = ~n35855 & ~n35923;
  assign n35925 = ~n7723 & ~n35924;
  assign n35926 = ~n35853 & ~n35925;
  assign n35927 = ~n7714 & ~n35926;
  assign n35928 = ~n35852 & ~n35927;
  assign n35929 = ~n7705 & ~n35928;
  assign n35930 = ~n35422 & ~n35929;
  assign n35931 = n7808 & ~n35930;
  assign n35932 = ~n8650 & ~n35931;
  assign n35933 = n8195 & ~n35932;
  assign n35934 = ~n8196 & ~n35933;
  assign n35935 = ~n8193 & ~n35934;
  assign n35936 = ~n10059 & ~n35563;
  assign n35937 = i_hbusreq7 & ~n35936;
  assign n35938 = ~n10074 & ~n35574;
  assign n35939 = ~i_hbusreq7 & ~n35938;
  assign n35940 = ~n35937 & ~n35939;
  assign n35941 = ~n7924 & ~n35940;
  assign n35942 = ~n15202 & ~n35584;
  assign n35943 = i_hbusreq7 & ~n35942;
  assign n35944 = ~n15228 & ~n35595;
  assign n35945 = ~i_hbusreq7 & ~n35944;
  assign n35946 = ~n35943 & ~n35945;
  assign n35947 = n7924 & ~n35946;
  assign n35948 = ~n35941 & ~n35947;
  assign n35949 = ~n8214 & ~n35948;
  assign n35950 = ~n10084 & ~n35563;
  assign n35951 = i_hbusreq7 & ~n35950;
  assign n35952 = ~n10098 & ~n35574;
  assign n35953 = ~i_hbusreq7 & ~n35952;
  assign n35954 = ~n35951 & ~n35953;
  assign n35955 = ~n7924 & ~n35954;
  assign n35956 = ~n15249 & ~n35584;
  assign n35957 = i_hbusreq7 & ~n35956;
  assign n35958 = ~n15278 & ~n35595;
  assign n35959 = ~i_hbusreq7 & ~n35958;
  assign n35960 = ~n35957 & ~n35959;
  assign n35961 = n7924 & ~n35960;
  assign n35962 = ~n35955 & ~n35961;
  assign n35963 = n8214 & ~n35962;
  assign n35964 = ~n35949 & ~n35963;
  assign n35965 = ~n8202 & ~n35964;
  assign n35966 = ~n10111 & ~n35563;
  assign n35967 = i_hbusreq7 & ~n35966;
  assign n35968 = ~n10126 & ~n35574;
  assign n35969 = ~i_hbusreq7 & ~n35968;
  assign n35970 = ~n35967 & ~n35969;
  assign n35971 = ~n7924 & ~n35970;
  assign n35972 = ~n15302 & ~n35584;
  assign n35973 = i_hbusreq7 & ~n35972;
  assign n35974 = ~n15338 & ~n35595;
  assign n35975 = ~i_hbusreq7 & ~n35974;
  assign n35976 = ~n35973 & ~n35975;
  assign n35977 = n7924 & ~n35976;
  assign n35978 = ~n35971 & ~n35977;
  assign n35979 = ~n8214 & ~n35978;
  assign n35980 = ~n10136 & ~n35563;
  assign n35981 = i_hbusreq7 & ~n35980;
  assign n35982 = ~n10150 & ~n35574;
  assign n35983 = ~i_hbusreq7 & ~n35982;
  assign n35984 = ~n35981 & ~n35983;
  assign n35985 = ~n7924 & ~n35984;
  assign n35986 = ~n15359 & ~n35584;
  assign n35987 = i_hbusreq7 & ~n35986;
  assign n35988 = ~n15396 & ~n35595;
  assign n35989 = ~i_hbusreq7 & ~n35988;
  assign n35990 = ~n35987 & ~n35989;
  assign n35991 = n7924 & ~n35990;
  assign n35992 = ~n35985 & ~n35991;
  assign n35993 = n8214 & ~n35992;
  assign n35994 = ~n35979 & ~n35993;
  assign n35995 = n8202 & ~n35994;
  assign n35996 = ~n35965 & ~n35995;
  assign n35997 = n7920 & ~n35996;
  assign n35998 = ~n10014 & ~n35997;
  assign n35999 = n7728 & ~n35998;
  assign n36000 = ~n10170 & ~n35797;
  assign n36001 = i_hlock7 & ~n36000;
  assign n36002 = ~n10180 & ~n35797;
  assign n36003 = ~i_hlock7 & ~n36002;
  assign n36004 = ~n36001 & ~n36003;
  assign n36005 = ~i_hbusreq7 & ~n36004;
  assign n36006 = ~n35637 & ~n36005;
  assign n36007 = ~n7924 & ~n36006;
  assign n36008 = ~n15437 & ~n35813;
  assign n36009 = i_hlock7 & ~n36008;
  assign n36010 = ~n15450 & ~n35813;
  assign n36011 = ~i_hlock7 & ~n36010;
  assign n36012 = ~n36009 & ~n36011;
  assign n36013 = ~i_hbusreq7 & ~n36012;
  assign n36014 = ~n35684 & ~n36013;
  assign n36015 = n7924 & ~n36014;
  assign n36016 = ~n36007 & ~n36015;
  assign n36017 = ~n8214 & ~n36016;
  assign n36018 = ~n10200 & ~n35797;
  assign n36019 = i_hlock7 & ~n36018;
  assign n36020 = ~n10206 & ~n35797;
  assign n36021 = ~i_hlock7 & ~n36020;
  assign n36022 = ~n36019 & ~n36021;
  assign n36023 = ~i_hbusreq7 & ~n36022;
  assign n36024 = ~n35637 & ~n36023;
  assign n36025 = ~n7924 & ~n36024;
  assign n36026 = ~n15495 & ~n35813;
  assign n36027 = i_hlock7 & ~n36026;
  assign n36028 = ~n15501 & ~n35813;
  assign n36029 = ~i_hlock7 & ~n36028;
  assign n36030 = ~n36027 & ~n36029;
  assign n36031 = ~i_hbusreq7 & ~n36030;
  assign n36032 = ~n35684 & ~n36031;
  assign n36033 = n7924 & ~n36032;
  assign n36034 = ~n36025 & ~n36033;
  assign n36035 = n8214 & ~n36034;
  assign n36036 = ~n36017 & ~n36035;
  assign n36037 = ~n8202 & ~n36036;
  assign n36038 = ~n10224 & ~n35797;
  assign n36039 = i_hlock7 & ~n36038;
  assign n36040 = ~n10236 & ~n35797;
  assign n36041 = ~i_hlock7 & ~n36040;
  assign n36042 = ~n36039 & ~n36041;
  assign n36043 = ~i_hbusreq7 & ~n36042;
  assign n36044 = ~n35637 & ~n36043;
  assign n36045 = ~n7924 & ~n36044;
  assign n36046 = ~n15550 & ~n35813;
  assign n36047 = i_hlock7 & ~n36046;
  assign n36048 = ~n15565 & ~n35813;
  assign n36049 = ~i_hlock7 & ~n36048;
  assign n36050 = ~n36047 & ~n36049;
  assign n36051 = ~i_hbusreq7 & ~n36050;
  assign n36052 = ~n35684 & ~n36051;
  assign n36053 = n7924 & ~n36052;
  assign n36054 = ~n36045 & ~n36053;
  assign n36055 = ~n8214 & ~n36054;
  assign n36056 = ~n10258 & ~n35797;
  assign n36057 = i_hlock7 & ~n36056;
  assign n36058 = ~n10264 & ~n35797;
  assign n36059 = ~i_hlock7 & ~n36058;
  assign n36060 = ~n36057 & ~n36059;
  assign n36061 = ~i_hbusreq7 & ~n36060;
  assign n36062 = ~n35637 & ~n36061;
  assign n36063 = ~n7924 & ~n36062;
  assign n36064 = ~n15620 & ~n35813;
  assign n36065 = i_hlock7 & ~n36064;
  assign n36066 = ~n15626 & ~n35813;
  assign n36067 = ~i_hlock7 & ~n36066;
  assign n36068 = ~n36065 & ~n36067;
  assign n36069 = ~i_hbusreq7 & ~n36068;
  assign n36070 = ~n35684 & ~n36069;
  assign n36071 = n7924 & ~n36070;
  assign n36072 = ~n36063 & ~n36071;
  assign n36073 = n8214 & ~n36072;
  assign n36074 = ~n36055 & ~n36073;
  assign n36075 = n8202 & ~n36074;
  assign n36076 = ~n36037 & ~n36075;
  assign n36077 = n7920 & ~n36076;
  assign n36078 = ~n10014 & ~n36077;
  assign n36079 = ~n7728 & ~n36078;
  assign n36080 = ~n35999 & ~n36079;
  assign n36081 = n7723 & ~n36080;
  assign n36082 = ~n7723 & ~n36078;
  assign n36083 = ~n36081 & ~n36082;
  assign n36084 = n7714 & ~n36083;
  assign n36085 = n7723 & ~n36078;
  assign n36086 = ~n8640 & ~n36077;
  assign n36087 = n7728 & ~n36086;
  assign n36088 = ~n35923 & ~n36087;
  assign n36089 = ~n7723 & ~n36088;
  assign n36090 = ~n36085 & ~n36089;
  assign n36091 = ~n7714 & ~n36090;
  assign n36092 = ~n36084 & ~n36091;
  assign n36093 = ~n7705 & ~n36092;
  assign n36094 = ~n10052 & ~n36093;
  assign n36095 = n7808 & ~n36094;
  assign n36096 = ~n9908 & ~n36095;
  assign n36097 = ~n8195 & ~n36096;
  assign n36098 = n7924 & ~n35919;
  assign n36099 = ~n8214 & ~n36098;
  assign n36100 = ~controllable_hmaster0 & ~n15665;
  assign n36101 = ~n9152 & ~n36100;
  assign n36102 = controllable_hmaster3 & ~n36101;
  assign n36103 = ~n8995 & ~n36102;
  assign n36104 = i_hbusreq7 & ~n36103;
  assign n36105 = i_hbusreq8 & ~n36101;
  assign n36106 = controllable_hmaster0 & ~n10756;
  assign n36107 = ~controllable_hmaster0 & ~n15704;
  assign n36108 = ~n36106 & ~n36107;
  assign n36109 = ~i_hbusreq8 & ~n36108;
  assign n36110 = ~n36105 & ~n36109;
  assign n36111 = controllable_hmaster3 & ~n36110;
  assign n36112 = ~n10786 & ~n36111;
  assign n36113 = ~i_hbusreq7 & ~n36112;
  assign n36114 = ~n36104 & ~n36113;
  assign n36115 = ~n7924 & ~n36114;
  assign n36116 = ~controllable_hmaster0 & ~n15719;
  assign n36117 = ~n13765 & ~n36116;
  assign n36118 = controllable_hmaster3 & ~n36117;
  assign n36119 = ~n13201 & ~n36118;
  assign n36120 = i_hbusreq7 & ~n36119;
  assign n36121 = i_hbusreq8 & ~n36117;
  assign n36122 = controllable_hmaster0 & ~n15806;
  assign n36123 = ~controllable_hmaster0 & ~n15778;
  assign n36124 = ~n36122 & ~n36123;
  assign n36125 = ~i_hbusreq8 & ~n36124;
  assign n36126 = ~n36121 & ~n36125;
  assign n36127 = controllable_hmaster3 & ~n36126;
  assign n36128 = ~n15856 & ~n36127;
  assign n36129 = ~i_hbusreq7 & ~n36128;
  assign n36130 = ~n36120 & ~n36129;
  assign n36131 = n7924 & ~n36130;
  assign n36132 = ~n36115 & ~n36131;
  assign n36133 = n8214 & ~n36132;
  assign n36134 = ~n36099 & ~n36133;
  assign n36135 = n8202 & ~n36134;
  assign n36136 = ~n10721 & ~n36135;
  assign n36137 = n7920 & ~n36136;
  assign n36138 = ~n10671 & ~n36137;
  assign n36139 = n7728 & ~n36138;
  assign n36140 = ~n10812 & ~n35919;
  assign n36141 = ~n8214 & ~n36140;
  assign n36142 = n8214 & ~n35920;
  assign n36143 = ~n36141 & ~n36142;
  assign n36144 = n8202 & ~n36143;
  assign n36145 = ~n10811 & ~n36144;
  assign n36146 = n7920 & ~n36145;
  assign n36147 = ~n10797 & ~n36146;
  assign n36148 = ~n7728 & ~n36147;
  assign n36149 = ~n36139 & ~n36148;
  assign n36150 = ~n7723 & ~n36149;
  assign n36151 = ~n7723 & ~n36150;
  assign n36152 = ~n7714 & ~n36151;
  assign n36153 = ~n7714 & ~n36152;
  assign n36154 = n7705 & ~n36153;
  assign n36155 = ~n10833 & ~n35563;
  assign n36156 = i_hbusreq7 & ~n36155;
  assign n36157 = ~n10847 & ~n35574;
  assign n36158 = ~i_hbusreq7 & ~n36157;
  assign n36159 = ~n36156 & ~n36158;
  assign n36160 = ~n7924 & ~n36159;
  assign n36161 = ~n15898 & ~n35584;
  assign n36162 = i_hbusreq7 & ~n36161;
  assign n36163 = ~n15937 & ~n35595;
  assign n36164 = ~i_hbusreq7 & ~n36163;
  assign n36165 = ~n36162 & ~n36164;
  assign n36166 = n7924 & ~n36165;
  assign n36167 = ~n36160 & ~n36166;
  assign n36168 = ~n8214 & ~n36167;
  assign n36169 = ~n10857 & ~n35563;
  assign n36170 = i_hbusreq7 & ~n36169;
  assign n36171 = controllable_hmaster0 & ~n10864;
  assign n36172 = ~controllable_hmaster0 & ~n15953;
  assign n36173 = ~n36171 & ~n36172;
  assign n36174 = ~i_hbusreq8 & ~n36173;
  assign n36175 = ~n35570 & ~n36174;
  assign n36176 = controllable_hmaster3 & ~n36175;
  assign n36177 = ~n10879 & ~n36176;
  assign n36178 = ~i_hbusreq7 & ~n36177;
  assign n36179 = ~n36170 & ~n36178;
  assign n36180 = ~n7924 & ~n36179;
  assign n36181 = ~n15972 & ~n35584;
  assign n36182 = i_hbusreq7 & ~n36181;
  assign n36183 = controllable_hmaster0 & ~n15989;
  assign n36184 = ~controllable_hmaster0 & ~n15981;
  assign n36185 = ~n36183 & ~n36184;
  assign n36186 = ~i_hbusreq8 & ~n36185;
  assign n36187 = ~n35591 & ~n36186;
  assign n36188 = controllable_hmaster3 & ~n36187;
  assign n36189 = ~n16009 & ~n36188;
  assign n36190 = ~i_hbusreq7 & ~n36189;
  assign n36191 = ~n36182 & ~n36190;
  assign n36192 = n7924 & ~n36191;
  assign n36193 = ~n36180 & ~n36192;
  assign n36194 = n8214 & ~n36193;
  assign n36195 = ~n36168 & ~n36194;
  assign n36196 = ~n8202 & ~n36195;
  assign n36197 = n8202 & ~n35920;
  assign n36198 = ~n36196 & ~n36197;
  assign n36199 = n7920 & ~n36198;
  assign n36200 = ~n10797 & ~n36199;
  assign n36201 = n7728 & ~n36200;
  assign n36202 = ~n10900 & ~n35797;
  assign n36203 = i_hlock7 & ~n36202;
  assign n36204 = ~n10910 & ~n35797;
  assign n36205 = ~i_hlock7 & ~n36204;
  assign n36206 = ~n36203 & ~n36205;
  assign n36207 = ~i_hbusreq7 & ~n36206;
  assign n36208 = ~n35637 & ~n36207;
  assign n36209 = ~n7924 & ~n36208;
  assign n36210 = ~n16065 & ~n35813;
  assign n36211 = i_hlock7 & ~n36210;
  assign n36212 = ~n16078 & ~n35813;
  assign n36213 = ~i_hlock7 & ~n36212;
  assign n36214 = ~n36211 & ~n36213;
  assign n36215 = ~i_hbusreq7 & ~n36214;
  assign n36216 = ~n35684 & ~n36215;
  assign n36217 = n7924 & ~n36216;
  assign n36218 = ~n36209 & ~n36217;
  assign n36219 = ~n8214 & ~n36218;
  assign n36220 = ~n36142 & ~n36219;
  assign n36221 = ~n8202 & ~n36220;
  assign n36222 = ~n36197 & ~n36221;
  assign n36223 = n7920 & ~n36222;
  assign n36224 = ~n10797 & ~n36223;
  assign n36225 = ~n7728 & ~n36224;
  assign n36226 = ~n36201 & ~n36225;
  assign n36227 = n7723 & ~n36226;
  assign n36228 = ~n7723 & ~n36224;
  assign n36229 = ~n36227 & ~n36228;
  assign n36230 = n7714 & ~n36229;
  assign n36231 = n7723 & ~n36224;
  assign n36232 = ~n8640 & ~n36223;
  assign n36233 = n7728 & ~n36232;
  assign n36234 = ~n35923 & ~n36233;
  assign n36235 = ~n7723 & ~n36234;
  assign n36236 = ~n36231 & ~n36235;
  assign n36237 = ~n7714 & ~n36236;
  assign n36238 = ~n36230 & ~n36237;
  assign n36239 = ~n7705 & ~n36238;
  assign n36240 = ~n36154 & ~n36239;
  assign n36241 = n7808 & ~n36240;
  assign n36242 = ~n10670 & ~n36241;
  assign n36243 = n8195 & ~n36242;
  assign n36244 = ~n36097 & ~n36243;
  assign n36245 = n8193 & ~n36244;
  assign n36246 = ~n35935 & ~n36245;
  assign n36247 = n8191 & ~n36246;
  assign n36248 = ~n11068 & ~n35302;
  assign n36249 = n7728 & ~n36248;
  assign n36250 = ~n11071 & ~n35414;
  assign n36251 = ~n7728 & ~n36250;
  assign n36252 = ~n36249 & ~n36251;
  assign n36253 = ~n7723 & ~n36252;
  assign n36254 = ~n7723 & ~n36253;
  assign n36255 = ~n7714 & ~n36254;
  assign n36256 = ~n7714 & ~n36255;
  assign n36257 = n7705 & ~n36256;
  assign n36258 = ~n11071 & ~n35623;
  assign n36259 = n7728 & ~n36258;
  assign n36260 = ~n11071 & ~n35845;
  assign n36261 = ~n7728 & ~n36260;
  assign n36262 = ~n36259 & ~n36261;
  assign n36263 = n7723 & ~n36262;
  assign n36264 = ~n7723 & ~n36260;
  assign n36265 = ~n36263 & ~n36264;
  assign n36266 = n7714 & ~n36265;
  assign n36267 = n7723 & ~n36260;
  assign n36268 = ~n11057 & ~n35845;
  assign n36269 = n7728 & ~n36268;
  assign n36270 = ~n11057 & ~n35921;
  assign n36271 = ~n7728 & ~n36270;
  assign n36272 = ~n36269 & ~n36271;
  assign n36273 = ~n7723 & ~n36272;
  assign n36274 = ~n36267 & ~n36273;
  assign n36275 = ~n7714 & ~n36274;
  assign n36276 = ~n36266 & ~n36275;
  assign n36277 = ~n7705 & ~n36276;
  assign n36278 = ~n36257 & ~n36277;
  assign n36279 = n7808 & ~n36278;
  assign n36280 = ~n11067 & ~n36279;
  assign n36281 = n8195 & ~n36280;
  assign n36282 = ~n8196 & ~n36281;
  assign n36283 = ~n8193 & ~n36282;
  assign n36284 = ~n11057 & ~n36077;
  assign n36285 = n7728 & ~n36284;
  assign n36286 = ~n36271 & ~n36285;
  assign n36287 = ~n7723 & ~n36286;
  assign n36288 = ~n36085 & ~n36287;
  assign n36289 = ~n7714 & ~n36288;
  assign n36290 = ~n36084 & ~n36289;
  assign n36291 = ~n7705 & ~n36290;
  assign n36292 = ~n10052 & ~n36291;
  assign n36293 = n7808 & ~n36292;
  assign n36294 = ~n11113 & ~n36293;
  assign n36295 = ~n8195 & ~n36294;
  assign n36296 = ~n11196 & ~n36137;
  assign n36297 = n7728 & ~n36296;
  assign n36298 = ~n11199 & ~n36146;
  assign n36299 = ~n7728 & ~n36298;
  assign n36300 = ~n36297 & ~n36299;
  assign n36301 = ~n7723 & ~n36300;
  assign n36302 = ~n7723 & ~n36301;
  assign n36303 = ~n7714 & ~n36302;
  assign n36304 = ~n7714 & ~n36303;
  assign n36305 = n7705 & ~n36304;
  assign n36306 = ~n11199 & ~n36199;
  assign n36307 = n7728 & ~n36306;
  assign n36308 = ~n11199 & ~n36223;
  assign n36309 = ~n7728 & ~n36308;
  assign n36310 = ~n36307 & ~n36309;
  assign n36311 = n7723 & ~n36310;
  assign n36312 = ~n7723 & ~n36308;
  assign n36313 = ~n36311 & ~n36312;
  assign n36314 = n7714 & ~n36313;
  assign n36315 = n7723 & ~n36308;
  assign n36316 = ~n11057 & ~n36223;
  assign n36317 = n7728 & ~n36316;
  assign n36318 = ~n36271 & ~n36317;
  assign n36319 = ~n7723 & ~n36318;
  assign n36320 = ~n36315 & ~n36319;
  assign n36321 = ~n7714 & ~n36320;
  assign n36322 = ~n36314 & ~n36321;
  assign n36323 = ~n7705 & ~n36322;
  assign n36324 = ~n36305 & ~n36323;
  assign n36325 = n7808 & ~n36324;
  assign n36326 = ~n11195 & ~n36325;
  assign n36327 = n8195 & ~n36326;
  assign n36328 = ~n36295 & ~n36327;
  assign n36329 = n8193 & ~n36328;
  assign n36330 = ~n36283 & ~n36329;
  assign n36331 = ~n8191 & ~n36330;
  assign n36332 = ~n36247 & ~n36331;
  assign n36333 = n8188 & ~n36332;
  assign n36334 = controllable_hgrant6 & ~n11239;
  assign n36335 = ~controllable_hmaster2 & ~n28601;
  assign n36336 = ~controllable_hmaster2 & ~n36335;
  assign n36337 = ~controllable_hmaster1 & ~n36336;
  assign n36338 = ~controllable_hmaster1 & ~n36337;
  assign n36339 = ~controllable_hgrant6 & ~n36338;
  assign n36340 = ~n36334 & ~n36339;
  assign n36341 = ~controllable_hmaster0 & ~n36340;
  assign n36342 = ~controllable_hmaster0 & ~n36341;
  assign n36343 = i_hlock8 & ~n36342;
  assign n36344 = controllable_hgrant6 & ~n11246;
  assign n36345 = ~controllable_hmaster2 & ~n28619;
  assign n36346 = ~controllable_hmaster2 & ~n36345;
  assign n36347 = ~controllable_hmaster1 & ~n36346;
  assign n36348 = ~controllable_hmaster1 & ~n36347;
  assign n36349 = ~controllable_hgrant6 & ~n36348;
  assign n36350 = ~n36344 & ~n36349;
  assign n36351 = ~controllable_hmaster0 & ~n36350;
  assign n36352 = ~controllable_hmaster0 & ~n36351;
  assign n36353 = ~i_hlock8 & ~n36352;
  assign n36354 = ~n36343 & ~n36353;
  assign n36355 = controllable_hmaster3 & ~n36354;
  assign n36356 = controllable_hmaster3 & ~n36355;
  assign n36357 = i_hbusreq7 & ~n36356;
  assign n36358 = i_hbusreq8 & ~n36354;
  assign n36359 = controllable_hgrant6 & ~n11261;
  assign n36360 = i_hbusreq6 & ~n36338;
  assign n36361 = ~controllable_hmaster2 & ~n28650;
  assign n36362 = ~controllable_hmaster2 & ~n36361;
  assign n36363 = ~controllable_hmaster1 & ~n36362;
  assign n36364 = ~controllable_hmaster1 & ~n36363;
  assign n36365 = ~i_hbusreq6 & ~n36364;
  assign n36366 = ~n36360 & ~n36365;
  assign n36367 = ~controllable_hgrant6 & ~n36366;
  assign n36368 = ~n36359 & ~n36367;
  assign n36369 = ~controllable_hmaster0 & ~n36368;
  assign n36370 = ~controllable_hmaster0 & ~n36369;
  assign n36371 = i_hlock8 & ~n36370;
  assign n36372 = controllable_hgrant6 & ~n11271;
  assign n36373 = i_hbusreq6 & ~n36348;
  assign n36374 = ~controllable_hmaster2 & ~n28683;
  assign n36375 = ~controllable_hmaster2 & ~n36374;
  assign n36376 = ~controllable_hmaster1 & ~n36375;
  assign n36377 = ~controllable_hmaster1 & ~n36376;
  assign n36378 = ~i_hbusreq6 & ~n36377;
  assign n36379 = ~n36373 & ~n36378;
  assign n36380 = ~controllable_hgrant6 & ~n36379;
  assign n36381 = ~n36372 & ~n36380;
  assign n36382 = ~controllable_hmaster0 & ~n36381;
  assign n36383 = ~controllable_hmaster0 & ~n36382;
  assign n36384 = ~i_hlock8 & ~n36383;
  assign n36385 = ~n36371 & ~n36384;
  assign n36386 = ~i_hbusreq8 & ~n36385;
  assign n36387 = ~n36358 & ~n36386;
  assign n36388 = controllable_hmaster3 & ~n36387;
  assign n36389 = controllable_hmaster3 & ~n36388;
  assign n36390 = ~i_hbusreq7 & ~n36389;
  assign n36391 = ~n36357 & ~n36390;
  assign n36392 = n7924 & ~n36391;
  assign n36393 = n7924 & ~n36392;
  assign n36394 = n8214 & ~n36393;
  assign n36395 = n8214 & ~n36394;
  assign n36396 = ~n8202 & ~n36395;
  assign n36397 = ~n8332 & ~n36396;
  assign n36398 = n7728 & ~n36397;
  assign n36399 = controllable_hgrant6 & ~n11291;
  assign n36400 = ~n7739 & ~n36335;
  assign n36401 = ~controllable_hmaster1 & ~n36400;
  assign n36402 = ~n7738 & ~n36401;
  assign n36403 = ~controllable_hgrant6 & ~n36402;
  assign n36404 = ~n36399 & ~n36403;
  assign n36405 = ~controllable_hmaster0 & ~n36404;
  assign n36406 = ~n8904 & ~n36405;
  assign n36407 = i_hlock8 & ~n36406;
  assign n36408 = controllable_hgrant6 & ~n11297;
  assign n36409 = ~n7739 & ~n36345;
  assign n36410 = ~controllable_hmaster1 & ~n36409;
  assign n36411 = ~n7738 & ~n36410;
  assign n36412 = ~controllable_hgrant6 & ~n36411;
  assign n36413 = ~n36408 & ~n36412;
  assign n36414 = ~controllable_hmaster0 & ~n36413;
  assign n36415 = ~n8904 & ~n36414;
  assign n36416 = ~i_hlock8 & ~n36415;
  assign n36417 = ~n36407 & ~n36416;
  assign n36418 = controllable_hmaster3 & ~n36417;
  assign n36419 = controllable_hmaster3 & ~n36418;
  assign n36420 = i_hbusreq7 & ~n36419;
  assign n36421 = i_hbusreq8 & ~n36417;
  assign n36422 = controllable_hgrant6 & ~n11311;
  assign n36423 = i_hbusreq6 & ~n36402;
  assign n36424 = ~n7771 & ~n36361;
  assign n36425 = ~controllable_hmaster1 & ~n36424;
  assign n36426 = ~n7770 & ~n36425;
  assign n36427 = ~i_hbusreq6 & ~n36426;
  assign n36428 = ~n36423 & ~n36427;
  assign n36429 = ~controllable_hgrant6 & ~n36428;
  assign n36430 = ~n36422 & ~n36429;
  assign n36431 = ~controllable_hmaster0 & ~n36430;
  assign n36432 = ~n8922 & ~n36431;
  assign n36433 = i_hlock8 & ~n36432;
  assign n36434 = controllable_hgrant6 & ~n11320;
  assign n36435 = i_hbusreq6 & ~n36411;
  assign n36436 = ~n7771 & ~n36374;
  assign n36437 = ~controllable_hmaster1 & ~n36436;
  assign n36438 = ~n7770 & ~n36437;
  assign n36439 = ~i_hbusreq6 & ~n36438;
  assign n36440 = ~n36435 & ~n36439;
  assign n36441 = ~controllable_hgrant6 & ~n36440;
  assign n36442 = ~n36434 & ~n36441;
  assign n36443 = ~controllable_hmaster0 & ~n36442;
  assign n36444 = ~n8922 & ~n36443;
  assign n36445 = ~i_hlock8 & ~n36444;
  assign n36446 = ~n36433 & ~n36445;
  assign n36447 = ~i_hbusreq8 & ~n36446;
  assign n36448 = ~n36421 & ~n36447;
  assign n36449 = controllable_hmaster3 & ~n36448;
  assign n36450 = controllable_hmaster3 & ~n36449;
  assign n36451 = ~i_hbusreq7 & ~n36450;
  assign n36452 = ~n36420 & ~n36451;
  assign n36453 = n7924 & ~n36452;
  assign n36454 = ~n8337 & ~n36453;
  assign n36455 = n8214 & ~n36454;
  assign n36456 = ~n8336 & ~n36455;
  assign n36457 = ~n8202 & ~n36456;
  assign n36458 = ~n8347 & ~n36457;
  assign n36459 = ~n7728 & ~n36458;
  assign n36460 = ~n36398 & ~n36459;
  assign n36461 = ~n7723 & ~n36460;
  assign n36462 = ~n7723 & ~n36461;
  assign n36463 = ~n7714 & ~n36462;
  assign n36464 = ~n7714 & ~n36463;
  assign n36465 = n7705 & ~n36464;
  assign n36466 = n7723 & ~n36458;
  assign n36467 = controllable_hgrant6 & ~n11348;
  assign n36468 = ~n8358 & ~n36335;
  assign n36469 = ~controllable_hmaster1 & ~n36468;
  assign n36470 = ~n8357 & ~n36469;
  assign n36471 = ~controllable_hgrant6 & ~n36470;
  assign n36472 = ~n36467 & ~n36471;
  assign n36473 = ~controllable_hmaster0 & ~n36472;
  assign n36474 = ~n11345 & ~n36473;
  assign n36475 = i_hlock8 & ~n36474;
  assign n36476 = controllable_hgrant6 & ~n11354;
  assign n36477 = ~n8358 & ~n36345;
  assign n36478 = ~controllable_hmaster1 & ~n36477;
  assign n36479 = ~n8357 & ~n36478;
  assign n36480 = ~controllable_hgrant6 & ~n36479;
  assign n36481 = ~n36476 & ~n36480;
  assign n36482 = ~controllable_hmaster0 & ~n36481;
  assign n36483 = ~n11345 & ~n36482;
  assign n36484 = ~i_hlock8 & ~n36483;
  assign n36485 = ~n36475 & ~n36484;
  assign n36486 = controllable_hmaster3 & ~n36485;
  assign n36487 = ~n8463 & ~n36486;
  assign n36488 = i_hbusreq7 & ~n36487;
  assign n36489 = i_hbusreq8 & ~n36485;
  assign n36490 = controllable_hgrant6 & ~n11369;
  assign n36491 = i_hbusreq6 & ~n36470;
  assign n36492 = ~n8484 & ~n36361;
  assign n36493 = ~controllable_hmaster1 & ~n36492;
  assign n36494 = ~n8483 & ~n36493;
  assign n36495 = ~i_hbusreq6 & ~n36494;
  assign n36496 = ~n36491 & ~n36495;
  assign n36497 = ~controllable_hgrant6 & ~n36496;
  assign n36498 = ~n36490 & ~n36497;
  assign n36499 = ~controllable_hmaster0 & ~n36498;
  assign n36500 = ~n11363 & ~n36499;
  assign n36501 = i_hlock8 & ~n36500;
  assign n36502 = controllable_hgrant6 & ~n11378;
  assign n36503 = i_hbusreq6 & ~n36479;
  assign n36504 = ~n8484 & ~n36374;
  assign n36505 = ~controllable_hmaster1 & ~n36504;
  assign n36506 = ~n8483 & ~n36505;
  assign n36507 = ~i_hbusreq6 & ~n36506;
  assign n36508 = ~n36503 & ~n36507;
  assign n36509 = ~controllable_hgrant6 & ~n36508;
  assign n36510 = ~n36502 & ~n36509;
  assign n36511 = ~controllable_hmaster0 & ~n36510;
  assign n36512 = ~n11363 & ~n36511;
  assign n36513 = ~i_hlock8 & ~n36512;
  assign n36514 = ~n36501 & ~n36513;
  assign n36515 = ~i_hbusreq8 & ~n36514;
  assign n36516 = ~n36489 & ~n36515;
  assign n36517 = controllable_hmaster3 & ~n36516;
  assign n36518 = ~n8634 & ~n36517;
  assign n36519 = ~i_hbusreq7 & ~n36518;
  assign n36520 = ~n36488 & ~n36519;
  assign n36521 = n7924 & ~n36520;
  assign n36522 = ~n8337 & ~n36521;
  assign n36523 = ~n7920 & ~n36522;
  assign n36524 = n7920 & ~n36458;
  assign n36525 = ~n36523 & ~n36524;
  assign n36526 = ~n7723 & ~n36525;
  assign n36527 = ~n36466 & ~n36526;
  assign n36528 = n7714 & ~n36527;
  assign n36529 = ~n7714 & ~n36522;
  assign n36530 = ~n36528 & ~n36529;
  assign n36531 = ~n7705 & ~n36530;
  assign n36532 = ~n36465 & ~n36531;
  assign n36533 = ~n7808 & ~n36532;
  assign n36534 = ~n7920 & ~n36397;
  assign n36535 = ~controllable_hmaster2 & ~n28869;
  assign n36536 = ~controllable_hmaster2 & ~n36535;
  assign n36537 = ~controllable_hmaster1 & ~n36536;
  assign n36538 = ~controllable_hmaster1 & ~n36537;
  assign n36539 = ~controllable_hgrant6 & ~n36538;
  assign n36540 = ~n16722 & ~n36539;
  assign n36541 = ~controllable_hmaster0 & ~n36540;
  assign n36542 = ~controllable_hmaster0 & ~n36541;
  assign n36543 = i_hlock8 & ~n36542;
  assign n36544 = ~controllable_hmaster2 & ~n28884;
  assign n36545 = ~controllable_hmaster2 & ~n36544;
  assign n36546 = ~controllable_hmaster1 & ~n36545;
  assign n36547 = ~controllable_hmaster1 & ~n36546;
  assign n36548 = ~controllable_hgrant6 & ~n36547;
  assign n36549 = ~n16754 & ~n36548;
  assign n36550 = ~controllable_hmaster0 & ~n36549;
  assign n36551 = ~controllable_hmaster0 & ~n36550;
  assign n36552 = ~i_hlock8 & ~n36551;
  assign n36553 = ~n36543 & ~n36552;
  assign n36554 = controllable_hmaster3 & ~n36553;
  assign n36555 = controllable_hmaster3 & ~n36554;
  assign n36556 = i_hbusreq7 & ~n36555;
  assign n36557 = i_hbusreq8 & ~n36553;
  assign n36558 = i_hbusreq6 & ~n36538;
  assign n36559 = ~controllable_hmaster2 & ~n28912;
  assign n36560 = ~controllable_hmaster2 & ~n36559;
  assign n36561 = ~controllable_hmaster1 & ~n36560;
  assign n36562 = ~controllable_hmaster1 & ~n36561;
  assign n36563 = ~i_hbusreq6 & ~n36562;
  assign n36564 = ~n36558 & ~n36563;
  assign n36565 = ~controllable_hgrant6 & ~n36564;
  assign n36566 = ~n16778 & ~n36565;
  assign n36567 = ~controllable_hmaster0 & ~n36566;
  assign n36568 = ~controllable_hmaster0 & ~n36567;
  assign n36569 = i_hlock8 & ~n36568;
  assign n36570 = i_hbusreq6 & ~n36547;
  assign n36571 = ~controllable_hmaster2 & ~n28942;
  assign n36572 = ~controllable_hmaster2 & ~n36571;
  assign n36573 = ~controllable_hmaster1 & ~n36572;
  assign n36574 = ~controllable_hmaster1 & ~n36573;
  assign n36575 = ~i_hbusreq6 & ~n36574;
  assign n36576 = ~n36570 & ~n36575;
  assign n36577 = ~controllable_hgrant6 & ~n36576;
  assign n36578 = ~n16848 & ~n36577;
  assign n36579 = ~controllable_hmaster0 & ~n36578;
  assign n36580 = ~controllable_hmaster0 & ~n36579;
  assign n36581 = ~i_hlock8 & ~n36580;
  assign n36582 = ~n36569 & ~n36581;
  assign n36583 = ~i_hbusreq8 & ~n36582;
  assign n36584 = ~n36557 & ~n36583;
  assign n36585 = controllable_hmaster3 & ~n36584;
  assign n36586 = controllable_hmaster3 & ~n36585;
  assign n36587 = ~i_hbusreq7 & ~n36586;
  assign n36588 = ~n36556 & ~n36587;
  assign n36589 = ~n7924 & ~n36588;
  assign n36590 = controllable_hmaster0 & ~n28967;
  assign n36591 = controllable_hmaster1 & ~n28965;
  assign n36592 = controllable_hmaster2 & ~n28965;
  assign n36593 = ~controllable_hmaster2 & ~n28972;
  assign n36594 = ~n36592 & ~n36593;
  assign n36595 = ~controllable_hmaster1 & ~n36594;
  assign n36596 = ~n36591 & ~n36595;
  assign n36597 = ~controllable_hgrant6 & ~n36596;
  assign n36598 = ~n16722 & ~n36597;
  assign n36599 = ~controllable_hmaster0 & ~n36598;
  assign n36600 = ~n36590 & ~n36599;
  assign n36601 = i_hlock8 & ~n36600;
  assign n36602 = controllable_hmaster0 & ~n28992;
  assign n36603 = controllable_hmaster1 & ~n28990;
  assign n36604 = controllable_hmaster2 & ~n28990;
  assign n36605 = ~controllable_hmaster2 & ~n28997;
  assign n36606 = ~n36604 & ~n36605;
  assign n36607 = ~controllable_hmaster1 & ~n36606;
  assign n36608 = ~n36603 & ~n36607;
  assign n36609 = ~controllable_hgrant6 & ~n36608;
  assign n36610 = ~n16754 & ~n36609;
  assign n36611 = ~controllable_hmaster0 & ~n36610;
  assign n36612 = ~n36602 & ~n36611;
  assign n36613 = ~i_hlock8 & ~n36612;
  assign n36614 = ~n36601 & ~n36613;
  assign n36615 = controllable_hmaster3 & ~n36614;
  assign n36616 = i_hlock8 & ~n28967;
  assign n36617 = ~i_hlock8 & ~n28992;
  assign n36618 = ~n36616 & ~n36617;
  assign n36619 = ~controllable_hmaster3 & ~n36618;
  assign n36620 = ~n36615 & ~n36619;
  assign n36621 = i_hbusreq7 & ~n36620;
  assign n36622 = i_hbusreq8 & ~n36614;
  assign n36623 = controllable_hmaster0 & ~n29032;
  assign n36624 = i_hbusreq6 & ~n36596;
  assign n36625 = controllable_hmaster1 & ~n29028;
  assign n36626 = controllable_hmaster2 & ~n29028;
  assign n36627 = ~controllable_hmaster2 & ~n29050;
  assign n36628 = ~n36626 & ~n36627;
  assign n36629 = ~controllable_hmaster1 & ~n36628;
  assign n36630 = ~n36625 & ~n36629;
  assign n36631 = ~i_hbusreq6 & ~n36630;
  assign n36632 = ~n36624 & ~n36631;
  assign n36633 = ~controllable_hgrant6 & ~n36632;
  assign n36634 = ~n16778 & ~n36633;
  assign n36635 = ~controllable_hmaster0 & ~n36634;
  assign n36636 = ~n36623 & ~n36635;
  assign n36637 = i_hlock8 & ~n36636;
  assign n36638 = controllable_hmaster0 & ~n29087;
  assign n36639 = i_hbusreq6 & ~n36608;
  assign n36640 = controllable_hmaster1 & ~n29083;
  assign n36641 = controllable_hmaster2 & ~n29083;
  assign n36642 = ~controllable_hmaster2 & ~n29105;
  assign n36643 = ~n36641 & ~n36642;
  assign n36644 = ~controllable_hmaster1 & ~n36643;
  assign n36645 = ~n36640 & ~n36644;
  assign n36646 = ~i_hbusreq6 & ~n36645;
  assign n36647 = ~n36639 & ~n36646;
  assign n36648 = ~controllable_hgrant6 & ~n36647;
  assign n36649 = ~n16848 & ~n36648;
  assign n36650 = ~controllable_hmaster0 & ~n36649;
  assign n36651 = ~n36638 & ~n36650;
  assign n36652 = ~i_hlock8 & ~n36651;
  assign n36653 = ~n36637 & ~n36652;
  assign n36654 = ~i_hbusreq8 & ~n36653;
  assign n36655 = ~n36622 & ~n36654;
  assign n36656 = controllable_hmaster3 & ~n36655;
  assign n36657 = i_hbusreq8 & ~n36618;
  assign n36658 = i_hlock8 & ~n29032;
  assign n36659 = ~i_hlock8 & ~n29087;
  assign n36660 = ~n36658 & ~n36659;
  assign n36661 = ~i_hbusreq8 & ~n36660;
  assign n36662 = ~n36657 & ~n36661;
  assign n36663 = ~controllable_hmaster3 & ~n36662;
  assign n36664 = ~n36656 & ~n36663;
  assign n36665 = ~i_hbusreq7 & ~n36664;
  assign n36666 = ~n36621 & ~n36665;
  assign n36667 = n7924 & ~n36666;
  assign n36668 = ~n36589 & ~n36667;
  assign n36669 = n8214 & ~n36668;
  assign n36670 = ~n28863 & ~n36669;
  assign n36671 = ~n8202 & ~n36670;
  assign n36672 = ~n16992 & ~n36671;
  assign n36673 = n7920 & ~n36672;
  assign n36674 = ~n36534 & ~n36673;
  assign n36675 = n7728 & ~n36674;
  assign n36676 = ~n7920 & ~n36458;
  assign n36677 = controllable_hmaster0 & ~n17022;
  assign n36678 = ~n17011 & ~n36535;
  assign n36679 = ~controllable_hmaster1 & ~n36678;
  assign n36680 = ~n17010 & ~n36679;
  assign n36681 = ~controllable_hgrant6 & ~n36680;
  assign n36682 = ~n17225 & ~n36681;
  assign n36683 = ~controllable_hmaster0 & ~n36682;
  assign n36684 = ~n36677 & ~n36683;
  assign n36685 = i_hlock8 & ~n36684;
  assign n36686 = ~n17011 & ~n36544;
  assign n36687 = ~controllable_hmaster1 & ~n36686;
  assign n36688 = ~n17010 & ~n36687;
  assign n36689 = ~controllable_hgrant6 & ~n36688;
  assign n36690 = ~n17234 & ~n36689;
  assign n36691 = ~controllable_hmaster0 & ~n36690;
  assign n36692 = ~n36677 & ~n36691;
  assign n36693 = ~i_hlock8 & ~n36692;
  assign n36694 = ~n36685 & ~n36693;
  assign n36695 = controllable_hmaster3 & ~n36694;
  assign n36696 = controllable_hmaster3 & ~n36695;
  assign n36697 = i_hbusreq7 & ~n36696;
  assign n36698 = i_hbusreq8 & ~n36694;
  assign n36699 = controllable_hmaster0 & ~n17078;
  assign n36700 = i_hbusreq6 & ~n36680;
  assign n36701 = ~n17062 & ~n36559;
  assign n36702 = ~controllable_hmaster1 & ~n36701;
  assign n36703 = ~n17061 & ~n36702;
  assign n36704 = ~i_hbusreq6 & ~n36703;
  assign n36705 = ~n36700 & ~n36704;
  assign n36706 = ~controllable_hgrant6 & ~n36705;
  assign n36707 = ~n17248 & ~n36706;
  assign n36708 = ~controllable_hmaster0 & ~n36707;
  assign n36709 = ~n36699 & ~n36708;
  assign n36710 = i_hlock8 & ~n36709;
  assign n36711 = i_hbusreq6 & ~n36688;
  assign n36712 = ~n17062 & ~n36571;
  assign n36713 = ~controllable_hmaster1 & ~n36712;
  assign n36714 = ~n17061 & ~n36713;
  assign n36715 = ~i_hbusreq6 & ~n36714;
  assign n36716 = ~n36711 & ~n36715;
  assign n36717 = ~controllable_hgrant6 & ~n36716;
  assign n36718 = ~n17260 & ~n36717;
  assign n36719 = ~controllable_hmaster0 & ~n36718;
  assign n36720 = ~n36699 & ~n36719;
  assign n36721 = ~i_hlock8 & ~n36720;
  assign n36722 = ~n36710 & ~n36721;
  assign n36723 = ~i_hbusreq8 & ~n36722;
  assign n36724 = ~n36698 & ~n36723;
  assign n36725 = controllable_hmaster3 & ~n36724;
  assign n36726 = controllable_hmaster3 & ~n36725;
  assign n36727 = ~i_hbusreq7 & ~n36726;
  assign n36728 = ~n36697 & ~n36727;
  assign n36729 = ~n7924 & ~n36728;
  assign n36730 = controllable_hmaster0 & ~n29195;
  assign n36731 = ~n29190 & ~n36593;
  assign n36732 = ~controllable_hmaster1 & ~n36731;
  assign n36733 = ~n29189 & ~n36732;
  assign n36734 = ~controllable_hgrant6 & ~n36733;
  assign n36735 = ~n17225 & ~n36734;
  assign n36736 = ~controllable_hmaster0 & ~n36735;
  assign n36737 = ~n36730 & ~n36736;
  assign n36738 = i_hlock8 & ~n36737;
  assign n36739 = controllable_hmaster0 & ~n29209;
  assign n36740 = ~n29204 & ~n36605;
  assign n36741 = ~controllable_hmaster1 & ~n36740;
  assign n36742 = ~n29203 & ~n36741;
  assign n36743 = ~controllable_hgrant6 & ~n36742;
  assign n36744 = ~n17234 & ~n36743;
  assign n36745 = ~controllable_hmaster0 & ~n36744;
  assign n36746 = ~n36739 & ~n36745;
  assign n36747 = ~i_hlock8 & ~n36746;
  assign n36748 = ~n36738 & ~n36747;
  assign n36749 = controllable_hmaster3 & ~n36748;
  assign n36750 = ~n36619 & ~n36749;
  assign n36751 = i_hbusreq7 & ~n36750;
  assign n36752 = i_hbusreq8 & ~n36748;
  assign n36753 = controllable_hmaster0 & ~n29238;
  assign n36754 = i_hbusreq6 & ~n36733;
  assign n36755 = ~n29231 & ~n36627;
  assign n36756 = ~controllable_hmaster1 & ~n36755;
  assign n36757 = ~n29230 & ~n36756;
  assign n36758 = ~i_hbusreq6 & ~n36757;
  assign n36759 = ~n36754 & ~n36758;
  assign n36760 = ~controllable_hgrant6 & ~n36759;
  assign n36761 = ~n17248 & ~n36760;
  assign n36762 = ~controllable_hmaster0 & ~n36761;
  assign n36763 = ~n36753 & ~n36762;
  assign n36764 = i_hlock8 & ~n36763;
  assign n36765 = controllable_hmaster0 & ~n29267;
  assign n36766 = i_hbusreq6 & ~n36742;
  assign n36767 = ~n29260 & ~n36642;
  assign n36768 = ~controllable_hmaster1 & ~n36767;
  assign n36769 = ~n29259 & ~n36768;
  assign n36770 = ~i_hbusreq6 & ~n36769;
  assign n36771 = ~n36766 & ~n36770;
  assign n36772 = ~controllable_hgrant6 & ~n36771;
  assign n36773 = ~n17260 & ~n36772;
  assign n36774 = ~controllable_hmaster0 & ~n36773;
  assign n36775 = ~n36765 & ~n36774;
  assign n36776 = ~i_hlock8 & ~n36775;
  assign n36777 = ~n36764 & ~n36776;
  assign n36778 = ~i_hbusreq8 & ~n36777;
  assign n36779 = ~n36752 & ~n36778;
  assign n36780 = controllable_hmaster3 & ~n36779;
  assign n36781 = ~n36663 & ~n36780;
  assign n36782 = ~i_hbusreq7 & ~n36781;
  assign n36783 = ~n36751 & ~n36782;
  assign n36784 = n7924 & ~n36783;
  assign n36785 = ~n36729 & ~n36784;
  assign n36786 = n8214 & ~n36785;
  assign n36787 = ~n29164 & ~n36786;
  assign n36788 = ~n8202 & ~n36787;
  assign n36789 = ~n17303 & ~n36788;
  assign n36790 = n7920 & ~n36789;
  assign n36791 = ~n36676 & ~n36790;
  assign n36792 = ~n7728 & ~n36791;
  assign n36793 = ~n36675 & ~n36792;
  assign n36794 = ~n7723 & ~n36793;
  assign n36795 = ~n7723 & ~n36794;
  assign n36796 = ~n7714 & ~n36795;
  assign n36797 = ~n7714 & ~n36796;
  assign n36798 = n7705 & ~n36797;
  assign n36799 = ~n29296 & ~n35423;
  assign n36800 = controllable_hmaster3 & ~n36799;
  assign n36801 = ~n8995 & ~n36800;
  assign n36802 = i_hbusreq7 & ~n36801;
  assign n36803 = i_hbusreq8 & ~n36799;
  assign n36804 = ~n29310 & ~n35429;
  assign n36805 = ~i_hbusreq8 & ~n36804;
  assign n36806 = ~n36803 & ~n36805;
  assign n36807 = controllable_hmaster3 & ~n36806;
  assign n36808 = ~n9041 & ~n36807;
  assign n36809 = ~i_hbusreq7 & ~n36808;
  assign n36810 = ~n36802 & ~n36809;
  assign n36811 = ~n7924 & ~n36810;
  assign n36812 = ~n29332 & ~n35438;
  assign n36813 = controllable_hmaster3 & ~n36812;
  assign n36814 = ~n13201 & ~n36813;
  assign n36815 = i_hbusreq7 & ~n36814;
  assign n36816 = i_hbusreq8 & ~n36812;
  assign n36817 = ~n29363 & ~n35444;
  assign n36818 = ~i_hbusreq8 & ~n36817;
  assign n36819 = ~n36816 & ~n36818;
  assign n36820 = controllable_hmaster3 & ~n36819;
  assign n36821 = ~n13641 & ~n36820;
  assign n36822 = ~i_hbusreq7 & ~n36821;
  assign n36823 = ~n36815 & ~n36822;
  assign n36824 = n7924 & ~n36823;
  assign n36825 = ~n36811 & ~n36824;
  assign n36826 = ~n8214 & ~n36825;
  assign n36827 = controllable_hmaster0 & ~n17345;
  assign n36828 = ~n17324 & ~n36535;
  assign n36829 = ~controllable_hmaster1 & ~n36828;
  assign n36830 = ~n17323 & ~n36829;
  assign n36831 = ~controllable_hgrant6 & ~n36830;
  assign n36832 = ~n13406 & ~n36831;
  assign n36833 = ~controllable_hmaster0 & ~n36832;
  assign n36834 = ~n36827 & ~n36833;
  assign n36835 = i_hlock8 & ~n36834;
  assign n36836 = ~n17324 & ~n36544;
  assign n36837 = ~controllable_hmaster1 & ~n36836;
  assign n36838 = ~n17323 & ~n36837;
  assign n36839 = ~controllable_hgrant6 & ~n36838;
  assign n36840 = ~n13427 & ~n36839;
  assign n36841 = ~controllable_hmaster0 & ~n36840;
  assign n36842 = ~n36827 & ~n36841;
  assign n36843 = ~i_hlock8 & ~n36842;
  assign n36844 = ~n36835 & ~n36843;
  assign n36845 = controllable_hmaster3 & ~n36844;
  assign n36846 = ~n17351 & ~n36845;
  assign n36847 = i_hbusreq7 & ~n36846;
  assign n36848 = i_hbusreq8 & ~n36844;
  assign n36849 = controllable_hmaster0 & ~n17442;
  assign n36850 = i_hbusreq6 & ~n36830;
  assign n36851 = ~n17392 & ~n36559;
  assign n36852 = ~controllable_hmaster1 & ~n36851;
  assign n36853 = ~n17391 & ~n36852;
  assign n36854 = ~i_hbusreq6 & ~n36853;
  assign n36855 = ~n36850 & ~n36854;
  assign n36856 = ~controllable_hgrant6 & ~n36855;
  assign n36857 = ~n13520 & ~n36856;
  assign n36858 = ~controllable_hmaster0 & ~n36857;
  assign n36859 = ~n36849 & ~n36858;
  assign n36860 = i_hlock8 & ~n36859;
  assign n36861 = i_hbusreq6 & ~n36838;
  assign n36862 = ~n17392 & ~n36571;
  assign n36863 = ~controllable_hmaster1 & ~n36862;
  assign n36864 = ~n17391 & ~n36863;
  assign n36865 = ~i_hbusreq6 & ~n36864;
  assign n36866 = ~n36861 & ~n36865;
  assign n36867 = ~controllable_hgrant6 & ~n36866;
  assign n36868 = ~n13573 & ~n36867;
  assign n36869 = ~controllable_hmaster0 & ~n36868;
  assign n36870 = ~n36849 & ~n36869;
  assign n36871 = ~i_hlock8 & ~n36870;
  assign n36872 = ~n36860 & ~n36871;
  assign n36873 = ~i_hbusreq8 & ~n36872;
  assign n36874 = ~n36848 & ~n36873;
  assign n36875 = controllable_hmaster3 & ~n36874;
  assign n36876 = ~n17456 & ~n36875;
  assign n36877 = ~i_hbusreq7 & ~n36876;
  assign n36878 = ~n36847 & ~n36877;
  assign n36879 = ~n7924 & ~n36878;
  assign n36880 = controllable_hmaster0 & ~n29502;
  assign n36881 = ~n29492 & ~n36593;
  assign n36882 = ~controllable_hmaster1 & ~n36881;
  assign n36883 = ~n29491 & ~n36882;
  assign n36884 = ~controllable_hgrant6 & ~n36883;
  assign n36885 = ~n13406 & ~n36884;
  assign n36886 = ~controllable_hmaster0 & ~n36885;
  assign n36887 = ~n36880 & ~n36886;
  assign n36888 = i_hlock8 & ~n36887;
  assign n36889 = controllable_hmaster0 & ~n29533;
  assign n36890 = ~n29523 & ~n36605;
  assign n36891 = ~controllable_hmaster1 & ~n36890;
  assign n36892 = ~n29522 & ~n36891;
  assign n36893 = ~controllable_hgrant6 & ~n36892;
  assign n36894 = ~n13427 & ~n36893;
  assign n36895 = ~controllable_hmaster0 & ~n36894;
  assign n36896 = ~n36889 & ~n36895;
  assign n36897 = ~i_hlock8 & ~n36896;
  assign n36898 = ~n36888 & ~n36897;
  assign n36899 = controllable_hmaster3 & ~n36898;
  assign n36900 = i_hlock8 & ~n29512;
  assign n36901 = ~i_hlock8 & ~n29543;
  assign n36902 = ~n36900 & ~n36901;
  assign n36903 = ~controllable_hmaster3 & ~n36902;
  assign n36904 = ~n36899 & ~n36903;
  assign n36905 = i_hbusreq7 & ~n36904;
  assign n36906 = i_hbusreq8 & ~n36898;
  assign n36907 = controllable_hmaster0 & ~n29588;
  assign n36908 = i_hbusreq6 & ~n36883;
  assign n36909 = ~n29567 & ~n36627;
  assign n36910 = ~controllable_hmaster1 & ~n36909;
  assign n36911 = ~n29566 & ~n36910;
  assign n36912 = ~i_hbusreq6 & ~n36911;
  assign n36913 = ~n36908 & ~n36912;
  assign n36914 = ~controllable_hgrant6 & ~n36913;
  assign n36915 = ~n13520 & ~n36914;
  assign n36916 = ~controllable_hmaster0 & ~n36915;
  assign n36917 = ~n36907 & ~n36916;
  assign n36918 = i_hlock8 & ~n36917;
  assign n36919 = controllable_hmaster0 & ~n29652;
  assign n36920 = i_hbusreq6 & ~n36892;
  assign n36921 = ~n29631 & ~n36642;
  assign n36922 = ~controllable_hmaster1 & ~n36921;
  assign n36923 = ~n29630 & ~n36922;
  assign n36924 = ~i_hbusreq6 & ~n36923;
  assign n36925 = ~n36920 & ~n36924;
  assign n36926 = ~controllable_hgrant6 & ~n36925;
  assign n36927 = ~n13573 & ~n36926;
  assign n36928 = ~controllable_hmaster0 & ~n36927;
  assign n36929 = ~n36919 & ~n36928;
  assign n36930 = ~i_hlock8 & ~n36929;
  assign n36931 = ~n36918 & ~n36930;
  assign n36932 = ~i_hbusreq8 & ~n36931;
  assign n36933 = ~n36906 & ~n36932;
  assign n36934 = controllable_hmaster3 & ~n36933;
  assign n36935 = i_hbusreq8 & ~n36902;
  assign n36936 = i_hlock8 & ~n29607;
  assign n36937 = ~i_hlock8 & ~n29671;
  assign n36938 = ~n36936 & ~n36937;
  assign n36939 = ~i_hbusreq8 & ~n36938;
  assign n36940 = ~n36935 & ~n36939;
  assign n36941 = ~controllable_hmaster3 & ~n36940;
  assign n36942 = ~n36934 & ~n36941;
  assign n36943 = ~i_hbusreq7 & ~n36942;
  assign n36944 = ~n36905 & ~n36943;
  assign n36945 = n7924 & ~n36944;
  assign n36946 = ~n36879 & ~n36945;
  assign n36947 = n8214 & ~n36946;
  assign n36948 = ~n36826 & ~n36947;
  assign n36949 = ~n8202 & ~n36948;
  assign n36950 = ~n17917 & ~n35563;
  assign n36951 = i_hlock7 & ~n36950;
  assign n36952 = ~n17927 & ~n35563;
  assign n36953 = ~i_hlock7 & ~n36952;
  assign n36954 = ~n36951 & ~n36953;
  assign n36955 = i_hbusreq7 & ~n36954;
  assign n36956 = ~n17945 & ~n35574;
  assign n36957 = i_hlock7 & ~n36956;
  assign n36958 = ~n17961 & ~n35574;
  assign n36959 = ~i_hlock7 & ~n36958;
  assign n36960 = ~n36957 & ~n36959;
  assign n36961 = ~i_hbusreq7 & ~n36960;
  assign n36962 = ~n36955 & ~n36961;
  assign n36963 = ~n7924 & ~n36962;
  assign n36964 = ~n17976 & ~n35584;
  assign n36965 = i_hlock7 & ~n36964;
  assign n36966 = ~n17987 & ~n35584;
  assign n36967 = ~i_hlock7 & ~n36966;
  assign n36968 = ~n36965 & ~n36967;
  assign n36969 = i_hbusreq7 & ~n36968;
  assign n36970 = ~n18006 & ~n35595;
  assign n36971 = i_hlock7 & ~n36970;
  assign n36972 = ~n18023 & ~n35595;
  assign n36973 = ~i_hlock7 & ~n36972;
  assign n36974 = ~n36971 & ~n36973;
  assign n36975 = ~i_hbusreq7 & ~n36974;
  assign n36976 = ~n36969 & ~n36975;
  assign n36977 = n7924 & ~n36976;
  assign n36978 = ~n36963 & ~n36977;
  assign n36979 = ~n8214 & ~n36978;
  assign n36980 = ~n18039 & ~n35563;
  assign n36981 = i_hbusreq7 & ~n36980;
  assign n36982 = ~n18055 & ~n35574;
  assign n36983 = ~i_hbusreq7 & ~n36982;
  assign n36984 = ~n36981 & ~n36983;
  assign n36985 = ~n7924 & ~n36984;
  assign n36986 = ~n18067 & ~n35584;
  assign n36987 = i_hbusreq7 & ~n36986;
  assign n36988 = ~n18083 & ~n35595;
  assign n36989 = ~i_hbusreq7 & ~n36988;
  assign n36990 = ~n36987 & ~n36989;
  assign n36991 = n7924 & ~n36990;
  assign n36992 = ~n36985 & ~n36991;
  assign n36993 = n8214 & ~n36992;
  assign n36994 = ~n36979 & ~n36993;
  assign n36995 = n8202 & ~n36994;
  assign n36996 = ~n36949 & ~n36995;
  assign n36997 = n7920 & ~n36996;
  assign n36998 = ~n36676 & ~n36997;
  assign n36999 = n7728 & ~n36998;
  assign n37000 = ~controllable_hmaster2 & ~n29734;
  assign n37001 = ~n19182 & ~n37000;
  assign n37002 = ~controllable_hmaster1 & ~n37001;
  assign n37003 = ~n19181 & ~n37002;
  assign n37004 = ~controllable_hgrant6 & ~n37003;
  assign n37005 = ~n13406 & ~n37004;
  assign n37006 = ~controllable_hmaster0 & ~n37005;
  assign n37007 = ~n29724 & ~n37006;
  assign n37008 = i_hlock8 & ~n37007;
  assign n37009 = ~controllable_hmaster2 & ~n29749;
  assign n37010 = ~n19182 & ~n37009;
  assign n37011 = ~controllable_hmaster1 & ~n37010;
  assign n37012 = ~n19181 & ~n37011;
  assign n37013 = ~controllable_hgrant6 & ~n37012;
  assign n37014 = ~n13427 & ~n37013;
  assign n37015 = ~controllable_hmaster0 & ~n37014;
  assign n37016 = ~n29724 & ~n37015;
  assign n37017 = ~i_hlock8 & ~n37016;
  assign n37018 = ~n37008 & ~n37017;
  assign n37019 = controllable_hmaster3 & ~n37018;
  assign n37020 = ~n19326 & ~n37019;
  assign n37021 = i_hlock7 & ~n37020;
  assign n37022 = ~n19336 & ~n37019;
  assign n37023 = ~i_hlock7 & ~n37022;
  assign n37024 = ~n37021 & ~n37023;
  assign n37025 = i_hbusreq7 & ~n37024;
  assign n37026 = i_hbusreq8 & ~n37018;
  assign n37027 = i_hbusreq6 & ~n37003;
  assign n37028 = ~controllable_hmaster2 & ~n29795;
  assign n37029 = ~n19367 & ~n37028;
  assign n37030 = ~controllable_hmaster1 & ~n37029;
  assign n37031 = ~n19366 & ~n37030;
  assign n37032 = ~i_hbusreq6 & ~n37031;
  assign n37033 = ~n37027 & ~n37032;
  assign n37034 = ~controllable_hgrant6 & ~n37033;
  assign n37035 = ~n14019 & ~n37034;
  assign n37036 = ~controllable_hmaster0 & ~n37035;
  assign n37037 = ~n29772 & ~n37036;
  assign n37038 = i_hlock8 & ~n37037;
  assign n37039 = i_hbusreq6 & ~n37012;
  assign n37040 = ~controllable_hmaster2 & ~n29825;
  assign n37041 = ~n19367 & ~n37040;
  assign n37042 = ~controllable_hmaster1 & ~n37041;
  assign n37043 = ~n19366 & ~n37042;
  assign n37044 = ~i_hbusreq6 & ~n37043;
  assign n37045 = ~n37039 & ~n37044;
  assign n37046 = ~controllable_hgrant6 & ~n37045;
  assign n37047 = ~n14054 & ~n37046;
  assign n37048 = ~controllable_hmaster0 & ~n37047;
  assign n37049 = ~n29772 & ~n37048;
  assign n37050 = ~i_hlock8 & ~n37049;
  assign n37051 = ~n37038 & ~n37050;
  assign n37052 = ~i_hbusreq8 & ~n37051;
  assign n37053 = ~n37026 & ~n37052;
  assign n37054 = controllable_hmaster3 & ~n37053;
  assign n37055 = ~n19648 & ~n37054;
  assign n37056 = i_hlock7 & ~n37055;
  assign n37057 = ~n19664 & ~n37054;
  assign n37058 = ~i_hlock7 & ~n37057;
  assign n37059 = ~n37056 & ~n37058;
  assign n37060 = ~i_hbusreq7 & ~n37059;
  assign n37061 = ~n37025 & ~n37060;
  assign n37062 = ~n7924 & ~n37061;
  assign n37063 = ~controllable_hmaster2 & ~n29868;
  assign n37064 = ~n19683 & ~n37063;
  assign n37065 = ~controllable_hmaster1 & ~n37064;
  assign n37066 = ~n19682 & ~n37065;
  assign n37067 = ~controllable_hgrant6 & ~n37066;
  assign n37068 = ~n13406 & ~n37067;
  assign n37069 = ~controllable_hmaster0 & ~n37068;
  assign n37070 = ~n29858 & ~n37069;
  assign n37071 = i_hlock8 & ~n37070;
  assign n37072 = ~controllable_hmaster2 & ~n29883;
  assign n37073 = ~n19683 & ~n37072;
  assign n37074 = ~controllable_hmaster1 & ~n37073;
  assign n37075 = ~n19682 & ~n37074;
  assign n37076 = ~controllable_hgrant6 & ~n37075;
  assign n37077 = ~n13427 & ~n37076;
  assign n37078 = ~controllable_hmaster0 & ~n37077;
  assign n37079 = ~n29858 & ~n37078;
  assign n37080 = ~i_hlock8 & ~n37079;
  assign n37081 = ~n37071 & ~n37080;
  assign n37082 = controllable_hmaster3 & ~n37081;
  assign n37083 = ~n19851 & ~n37082;
  assign n37084 = i_hlock7 & ~n37083;
  assign n37085 = ~n19861 & ~n37082;
  assign n37086 = ~i_hlock7 & ~n37085;
  assign n37087 = ~n37084 & ~n37086;
  assign n37088 = i_hbusreq7 & ~n37087;
  assign n37089 = i_hbusreq8 & ~n37081;
  assign n37090 = i_hbusreq6 & ~n37066;
  assign n37091 = ~controllable_hmaster2 & ~n29946;
  assign n37092 = ~n19895 & ~n37091;
  assign n37093 = ~controllable_hmaster1 & ~n37092;
  assign n37094 = ~n19894 & ~n37093;
  assign n37095 = ~i_hbusreq6 & ~n37094;
  assign n37096 = ~n37090 & ~n37095;
  assign n37097 = ~controllable_hgrant6 & ~n37096;
  assign n37098 = ~n14019 & ~n37097;
  assign n37099 = ~controllable_hmaster0 & ~n37098;
  assign n37100 = ~n29923 & ~n37099;
  assign n37101 = i_hlock8 & ~n37100;
  assign n37102 = i_hbusreq6 & ~n37075;
  assign n37103 = ~controllable_hmaster2 & ~n29976;
  assign n37104 = ~n19895 & ~n37103;
  assign n37105 = ~controllable_hmaster1 & ~n37104;
  assign n37106 = ~n19894 & ~n37105;
  assign n37107 = ~i_hbusreq6 & ~n37106;
  assign n37108 = ~n37102 & ~n37107;
  assign n37109 = ~controllable_hgrant6 & ~n37108;
  assign n37110 = ~n14054 & ~n37109;
  assign n37111 = ~controllable_hmaster0 & ~n37110;
  assign n37112 = ~n29923 & ~n37111;
  assign n37113 = ~i_hlock8 & ~n37112;
  assign n37114 = ~n37101 & ~n37113;
  assign n37115 = ~i_hbusreq8 & ~n37114;
  assign n37116 = ~n37089 & ~n37115;
  assign n37117 = controllable_hmaster3 & ~n37116;
  assign n37118 = ~n20241 & ~n37117;
  assign n37119 = i_hlock7 & ~n37118;
  assign n37120 = ~n20257 & ~n37117;
  assign n37121 = ~i_hlock7 & ~n37120;
  assign n37122 = ~n37119 & ~n37121;
  assign n37123 = ~i_hbusreq7 & ~n37122;
  assign n37124 = ~n37088 & ~n37123;
  assign n37125 = n7924 & ~n37124;
  assign n37126 = ~n37062 & ~n37125;
  assign n37127 = ~n8214 & ~n37126;
  assign n37128 = ~n30145 & ~n36833;
  assign n37129 = i_hlock8 & ~n37128;
  assign n37130 = ~n30145 & ~n36841;
  assign n37131 = ~i_hlock8 & ~n37130;
  assign n37132 = ~n37129 & ~n37131;
  assign n37133 = controllable_hmaster3 & ~n37132;
  assign n37134 = ~n18193 & ~n37133;
  assign n37135 = i_hlock7 & ~n37134;
  assign n37136 = ~n18203 & ~n37133;
  assign n37137 = ~i_hlock7 & ~n37136;
  assign n37138 = ~n37135 & ~n37137;
  assign n37139 = i_hbusreq7 & ~n37138;
  assign n37140 = i_hbusreq8 & ~n37132;
  assign n37141 = ~n18248 & ~n36559;
  assign n37142 = ~controllable_hmaster1 & ~n37141;
  assign n37143 = ~n18247 & ~n37142;
  assign n37144 = ~i_hbusreq6 & ~n37143;
  assign n37145 = ~n36850 & ~n37144;
  assign n37146 = ~controllable_hgrant6 & ~n37145;
  assign n37147 = ~n14443 & ~n37146;
  assign n37148 = ~controllable_hmaster0 & ~n37147;
  assign n37149 = ~n30197 & ~n37148;
  assign n37150 = i_hlock8 & ~n37149;
  assign n37151 = ~n18248 & ~n36571;
  assign n37152 = ~controllable_hmaster1 & ~n37151;
  assign n37153 = ~n18247 & ~n37152;
  assign n37154 = ~i_hbusreq6 & ~n37153;
  assign n37155 = ~n36861 & ~n37154;
  assign n37156 = ~controllable_hgrant6 & ~n37155;
  assign n37157 = ~n14484 & ~n37156;
  assign n37158 = ~controllable_hmaster0 & ~n37157;
  assign n37159 = ~n30197 & ~n37158;
  assign n37160 = ~i_hlock8 & ~n37159;
  assign n37161 = ~n37150 & ~n37160;
  assign n37162 = ~i_hbusreq8 & ~n37161;
  assign n37163 = ~n37140 & ~n37162;
  assign n37164 = controllable_hmaster3 & ~n37163;
  assign n37165 = ~n18507 & ~n37164;
  assign n37166 = i_hlock7 & ~n37165;
  assign n37167 = ~n18523 & ~n37164;
  assign n37168 = ~i_hlock7 & ~n37167;
  assign n37169 = ~n37166 & ~n37168;
  assign n37170 = ~i_hbusreq7 & ~n37169;
  assign n37171 = ~n37139 & ~n37170;
  assign n37172 = ~n7924 & ~n37171;
  assign n37173 = ~n30254 & ~n36886;
  assign n37174 = i_hlock8 & ~n37173;
  assign n37175 = ~n30357 & ~n36895;
  assign n37176 = ~i_hlock8 & ~n37175;
  assign n37177 = ~n37174 & ~n37176;
  assign n37178 = controllable_hmaster3 & ~n37177;
  assign n37179 = ~n30287 & ~n30307;
  assign n37180 = controllable_hmaster1 & ~n37179;
  assign n37181 = ~n30302 & ~n37180;
  assign n37182 = ~controllable_hgrant6 & ~n37181;
  assign n37183 = ~n13849 & ~n37182;
  assign n37184 = controllable_hmaster0 & ~n37183;
  assign n37185 = ~n30340 & ~n37184;
  assign n37186 = i_hlock8 & ~n37185;
  assign n37187 = ~n30390 & ~n30410;
  assign n37188 = controllable_hmaster1 & ~n37187;
  assign n37189 = ~n30405 & ~n37188;
  assign n37190 = ~controllable_hgrant6 & ~n37189;
  assign n37191 = ~n13849 & ~n37190;
  assign n37192 = controllable_hmaster0 & ~n37191;
  assign n37193 = ~n30443 & ~n37192;
  assign n37194 = ~i_hlock8 & ~n37193;
  assign n37195 = ~n37186 & ~n37194;
  assign n37196 = ~controllable_hmaster3 & ~n37195;
  assign n37197 = ~n37178 & ~n37196;
  assign n37198 = i_hlock7 & ~n37197;
  assign n37199 = ~n30287 & ~n30332;
  assign n37200 = controllable_hmaster1 & ~n37199;
  assign n37201 = ~n30302 & ~n37200;
  assign n37202 = ~controllable_hgrant6 & ~n37201;
  assign n37203 = ~n13951 & ~n37202;
  assign n37204 = controllable_hmaster0 & ~n37203;
  assign n37205 = ~n30340 & ~n37204;
  assign n37206 = i_hlock8 & ~n37205;
  assign n37207 = ~n30390 & ~n30435;
  assign n37208 = controllable_hmaster1 & ~n37207;
  assign n37209 = ~n30405 & ~n37208;
  assign n37210 = ~controllable_hgrant6 & ~n37209;
  assign n37211 = ~n13951 & ~n37210;
  assign n37212 = controllable_hmaster0 & ~n37211;
  assign n37213 = ~n30443 & ~n37212;
  assign n37214 = ~i_hlock8 & ~n37213;
  assign n37215 = ~n37206 & ~n37214;
  assign n37216 = ~controllable_hmaster3 & ~n37215;
  assign n37217 = ~n37178 & ~n37216;
  assign n37218 = ~i_hlock7 & ~n37217;
  assign n37219 = ~n37198 & ~n37218;
  assign n37220 = i_hbusreq7 & ~n37219;
  assign n37221 = i_hbusreq8 & ~n37177;
  assign n37222 = ~n30463 & ~n36627;
  assign n37223 = ~controllable_hmaster1 & ~n37222;
  assign n37224 = ~n30462 & ~n37223;
  assign n37225 = ~i_hbusreq6 & ~n37224;
  assign n37226 = ~n36908 & ~n37225;
  assign n37227 = ~controllable_hgrant6 & ~n37226;
  assign n37228 = ~n14443 & ~n37227;
  assign n37229 = ~controllable_hmaster0 & ~n37228;
  assign n37230 = ~n30487 & ~n37229;
  assign n37231 = i_hlock8 & ~n37230;
  assign n37232 = ~n30671 & ~n36642;
  assign n37233 = ~controllable_hmaster1 & ~n37232;
  assign n37234 = ~n30670 & ~n37233;
  assign n37235 = ~i_hbusreq6 & ~n37234;
  assign n37236 = ~n36920 & ~n37235;
  assign n37237 = ~controllable_hgrant6 & ~n37236;
  assign n37238 = ~n14484 & ~n37237;
  assign n37239 = ~controllable_hmaster0 & ~n37238;
  assign n37240 = ~n30695 & ~n37239;
  assign n37241 = ~i_hlock8 & ~n37240;
  assign n37242 = ~n37231 & ~n37241;
  assign n37243 = ~i_hbusreq8 & ~n37242;
  assign n37244 = ~n37221 & ~n37243;
  assign n37245 = controllable_hmaster3 & ~n37244;
  assign n37246 = i_hbusreq8 & ~n37195;
  assign n37247 = i_hbusreq6 & ~n37181;
  assign n37248 = ~n30557 & ~n30592;
  assign n37249 = controllable_hmaster1 & ~n37248;
  assign n37250 = ~n30584 & ~n37249;
  assign n37251 = ~i_hbusreq6 & ~n37250;
  assign n37252 = ~n37247 & ~n37251;
  assign n37253 = ~controllable_hgrant6 & ~n37252;
  assign n37254 = ~n14094 & ~n37253;
  assign n37255 = controllable_hmaster0 & ~n37254;
  assign n37256 = ~n30651 & ~n37255;
  assign n37257 = i_hlock8 & ~n37256;
  assign n37258 = i_hbusreq6 & ~n37189;
  assign n37259 = ~n30765 & ~n30800;
  assign n37260 = controllable_hmaster1 & ~n37259;
  assign n37261 = ~n30792 & ~n37260;
  assign n37262 = ~i_hbusreq6 & ~n37261;
  assign n37263 = ~n37258 & ~n37262;
  assign n37264 = ~controllable_hgrant6 & ~n37263;
  assign n37265 = ~n14094 & ~n37264;
  assign n37266 = controllable_hmaster0 & ~n37265;
  assign n37267 = ~n30859 & ~n37266;
  assign n37268 = ~i_hlock8 & ~n37267;
  assign n37269 = ~n37257 & ~n37268;
  assign n37270 = ~i_hbusreq8 & ~n37269;
  assign n37271 = ~n37246 & ~n37270;
  assign n37272 = ~controllable_hmaster3 & ~n37271;
  assign n37273 = ~n37245 & ~n37272;
  assign n37274 = i_hlock7 & ~n37273;
  assign n37275 = i_hbusreq8 & ~n37215;
  assign n37276 = i_hbusreq6 & ~n37201;
  assign n37277 = ~n30557 & ~n30641;
  assign n37278 = controllable_hmaster1 & ~n37277;
  assign n37279 = ~n30584 & ~n37278;
  assign n37280 = ~i_hbusreq6 & ~n37279;
  assign n37281 = ~n37276 & ~n37280;
  assign n37282 = ~controllable_hgrant6 & ~n37281;
  assign n37283 = ~n14298 & ~n37282;
  assign n37284 = controllable_hmaster0 & ~n37283;
  assign n37285 = ~n30651 & ~n37284;
  assign n37286 = i_hlock8 & ~n37285;
  assign n37287 = i_hbusreq6 & ~n37209;
  assign n37288 = ~n30765 & ~n30849;
  assign n37289 = controllable_hmaster1 & ~n37288;
  assign n37290 = ~n30792 & ~n37289;
  assign n37291 = ~i_hbusreq6 & ~n37290;
  assign n37292 = ~n37287 & ~n37291;
  assign n37293 = ~controllable_hgrant6 & ~n37292;
  assign n37294 = ~n14298 & ~n37293;
  assign n37295 = controllable_hmaster0 & ~n37294;
  assign n37296 = ~n30859 & ~n37295;
  assign n37297 = ~i_hlock8 & ~n37296;
  assign n37298 = ~n37286 & ~n37297;
  assign n37299 = ~i_hbusreq8 & ~n37298;
  assign n37300 = ~n37275 & ~n37299;
  assign n37301 = ~controllable_hmaster3 & ~n37300;
  assign n37302 = ~n37245 & ~n37301;
  assign n37303 = ~i_hlock7 & ~n37302;
  assign n37304 = ~n37274 & ~n37303;
  assign n37305 = ~i_hbusreq7 & ~n37304;
  assign n37306 = ~n37220 & ~n37305;
  assign n37307 = n7924 & ~n37306;
  assign n37308 = ~n37172 & ~n37307;
  assign n37309 = n8214 & ~n37308;
  assign n37310 = ~n37127 & ~n37309;
  assign n37311 = ~n8202 & ~n37310;
  assign n37312 = ~n30011 & ~n37006;
  assign n37313 = i_hlock8 & ~n37312;
  assign n37314 = ~n30011 & ~n37015;
  assign n37315 = ~i_hlock8 & ~n37314;
  assign n37316 = ~n37313 & ~n37315;
  assign n37317 = controllable_hmaster3 & ~n37316;
  assign n37318 = ~n20295 & ~n37317;
  assign n37319 = i_hlock7 & ~n37318;
  assign n37320 = ~n20305 & ~n37317;
  assign n37321 = ~i_hlock7 & ~n37320;
  assign n37322 = ~n37319 & ~n37321;
  assign n37323 = i_hbusreq7 & ~n37322;
  assign n37324 = i_hbusreq8 & ~n37316;
  assign n37325 = ~n30050 & ~n37036;
  assign n37326 = i_hlock8 & ~n37325;
  assign n37327 = ~n30050 & ~n37048;
  assign n37328 = ~i_hlock8 & ~n37327;
  assign n37329 = ~n37326 & ~n37328;
  assign n37330 = ~i_hbusreq8 & ~n37329;
  assign n37331 = ~n37324 & ~n37330;
  assign n37332 = controllable_hmaster3 & ~n37331;
  assign n37333 = ~n20352 & ~n37332;
  assign n37334 = i_hlock7 & ~n37333;
  assign n37335 = ~n20368 & ~n37332;
  assign n37336 = ~i_hlock7 & ~n37335;
  assign n37337 = ~n37334 & ~n37336;
  assign n37338 = ~i_hbusreq7 & ~n37337;
  assign n37339 = ~n37323 & ~n37338;
  assign n37340 = ~n7924 & ~n37339;
  assign n37341 = ~n30080 & ~n37069;
  assign n37342 = i_hlock8 & ~n37341;
  assign n37343 = ~n30080 & ~n37078;
  assign n37344 = ~i_hlock8 & ~n37343;
  assign n37345 = ~n37342 & ~n37344;
  assign n37346 = controllable_hmaster3 & ~n37345;
  assign n37347 = ~n20403 & ~n37346;
  assign n37348 = i_hlock7 & ~n37347;
  assign n37349 = ~n20414 & ~n37346;
  assign n37350 = ~i_hlock7 & ~n37349;
  assign n37351 = ~n37348 & ~n37350;
  assign n37352 = i_hbusreq7 & ~n37351;
  assign n37353 = i_hbusreq8 & ~n37345;
  assign n37354 = ~n30119 & ~n37099;
  assign n37355 = i_hlock8 & ~n37354;
  assign n37356 = ~n30119 & ~n37111;
  assign n37357 = ~i_hlock8 & ~n37356;
  assign n37358 = ~n37355 & ~n37357;
  assign n37359 = ~i_hbusreq8 & ~n37358;
  assign n37360 = ~n37353 & ~n37359;
  assign n37361 = controllable_hmaster3 & ~n37360;
  assign n37362 = ~n20462 & ~n37361;
  assign n37363 = i_hlock7 & ~n37362;
  assign n37364 = ~n20479 & ~n37361;
  assign n37365 = ~i_hlock7 & ~n37364;
  assign n37366 = ~n37363 & ~n37365;
  assign n37367 = ~i_hbusreq7 & ~n37366;
  assign n37368 = ~n37352 & ~n37367;
  assign n37369 = n7924 & ~n37368;
  assign n37370 = ~n37340 & ~n37369;
  assign n37371 = ~n8214 & ~n37370;
  assign n37372 = ~n20501 & ~n37317;
  assign n37373 = i_hlock7 & ~n37372;
  assign n37374 = ~n20505 & ~n37317;
  assign n37375 = ~i_hlock7 & ~n37374;
  assign n37376 = ~n37373 & ~n37375;
  assign n37377 = i_hbusreq7 & ~n37376;
  assign n37378 = ~n20529 & ~n37332;
  assign n37379 = i_hlock7 & ~n37378;
  assign n37380 = ~n20536 & ~n37332;
  assign n37381 = ~i_hlock7 & ~n37380;
  assign n37382 = ~n37379 & ~n37381;
  assign n37383 = ~i_hbusreq7 & ~n37382;
  assign n37384 = ~n37377 & ~n37383;
  assign n37385 = ~n7924 & ~n37384;
  assign n37386 = ~n20556 & ~n37346;
  assign n37387 = i_hlock7 & ~n37386;
  assign n37388 = ~n20560 & ~n37346;
  assign n37389 = ~i_hlock7 & ~n37388;
  assign n37390 = ~n37387 & ~n37389;
  assign n37391 = i_hbusreq7 & ~n37390;
  assign n37392 = ~n20584 & ~n37361;
  assign n37393 = i_hlock7 & ~n37392;
  assign n37394 = ~n20591 & ~n37361;
  assign n37395 = ~i_hlock7 & ~n37394;
  assign n37396 = ~n37393 & ~n37395;
  assign n37397 = ~i_hbusreq7 & ~n37396;
  assign n37398 = ~n37391 & ~n37397;
  assign n37399 = n7924 & ~n37398;
  assign n37400 = ~n37385 & ~n37399;
  assign n37401 = n8214 & ~n37400;
  assign n37402 = ~n37371 & ~n37401;
  assign n37403 = n8202 & ~n37402;
  assign n37404 = ~n37311 & ~n37403;
  assign n37405 = n7920 & ~n37404;
  assign n37406 = ~n36676 & ~n37405;
  assign n37407 = ~n7728 & ~n37406;
  assign n37408 = ~n36999 & ~n37407;
  assign n37409 = n7723 & ~n37408;
  assign n37410 = ~n7723 & ~n37406;
  assign n37411 = ~n37409 & ~n37410;
  assign n37412 = n7714 & ~n37411;
  assign n37413 = n7723 & ~n37406;
  assign n37414 = ~controllable_hmaster2 & ~n31015;
  assign n37415 = ~n30977 & ~n37414;
  assign n37416 = ~controllable_hmaster1 & ~n37415;
  assign n37417 = ~n30976 & ~n37416;
  assign n37418 = ~controllable_hgrant6 & ~n37417;
  assign n37419 = ~n13406 & ~n37418;
  assign n37420 = ~controllable_hmaster0 & ~n37419;
  assign n37421 = ~n30983 & ~n37420;
  assign n37422 = i_hlock8 & ~n37421;
  assign n37423 = ~controllable_hmaster2 & ~n31122;
  assign n37424 = ~n31084 & ~n37423;
  assign n37425 = ~controllable_hmaster1 & ~n37424;
  assign n37426 = ~n31083 & ~n37425;
  assign n37427 = ~controllable_hgrant6 & ~n37426;
  assign n37428 = ~n13427 & ~n37427;
  assign n37429 = ~controllable_hmaster0 & ~n37428;
  assign n37430 = ~n31090 & ~n37429;
  assign n37431 = ~i_hlock8 & ~n37430;
  assign n37432 = ~n37422 & ~n37431;
  assign n37433 = controllable_hmaster3 & ~n37432;
  assign n37434 = ~n31021 & ~n31041;
  assign n37435 = controllable_hmaster1 & ~n37434;
  assign n37436 = ~n31036 & ~n37435;
  assign n37437 = ~controllable_hgrant6 & ~n37436;
  assign n37438 = ~n13849 & ~n37437;
  assign n37439 = controllable_hmaster0 & ~n37438;
  assign n37440 = ~n31074 & ~n37439;
  assign n37441 = i_hlock8 & ~n37440;
  assign n37442 = ~n31128 & ~n31148;
  assign n37443 = controllable_hmaster1 & ~n37442;
  assign n37444 = ~n31143 & ~n37443;
  assign n37445 = ~controllable_hgrant6 & ~n37444;
  assign n37446 = ~n13849 & ~n37445;
  assign n37447 = controllable_hmaster0 & ~n37446;
  assign n37448 = ~n31181 & ~n37447;
  assign n37449 = ~i_hlock8 & ~n37448;
  assign n37450 = ~n37441 & ~n37449;
  assign n37451 = ~controllable_hmaster3 & ~n37450;
  assign n37452 = ~n37433 & ~n37451;
  assign n37453 = i_hlock7 & ~n37452;
  assign n37454 = ~n31021 & ~n31066;
  assign n37455 = controllable_hmaster1 & ~n37454;
  assign n37456 = ~n31036 & ~n37455;
  assign n37457 = ~controllable_hgrant6 & ~n37456;
  assign n37458 = ~n13951 & ~n37457;
  assign n37459 = controllable_hmaster0 & ~n37458;
  assign n37460 = ~n31074 & ~n37459;
  assign n37461 = i_hlock8 & ~n37460;
  assign n37462 = ~n31128 & ~n31173;
  assign n37463 = controllable_hmaster1 & ~n37462;
  assign n37464 = ~n31143 & ~n37463;
  assign n37465 = ~controllable_hgrant6 & ~n37464;
  assign n37466 = ~n13951 & ~n37465;
  assign n37467 = controllable_hmaster0 & ~n37466;
  assign n37468 = ~n31181 & ~n37467;
  assign n37469 = ~i_hlock8 & ~n37468;
  assign n37470 = ~n37461 & ~n37469;
  assign n37471 = ~controllable_hmaster3 & ~n37470;
  assign n37472 = ~n37433 & ~n37471;
  assign n37473 = ~i_hlock7 & ~n37472;
  assign n37474 = ~n37453 & ~n37473;
  assign n37475 = i_hbusreq7 & ~n37474;
  assign n37476 = i_hbusreq8 & ~n37432;
  assign n37477 = i_hbusreq6 & ~n37417;
  assign n37478 = ~controllable_hmaster2 & ~n31294;
  assign n37479 = ~n31204 & ~n37478;
  assign n37480 = ~controllable_hmaster1 & ~n37479;
  assign n37481 = ~n31203 & ~n37480;
  assign n37482 = ~i_hbusreq6 & ~n37481;
  assign n37483 = ~n37477 & ~n37482;
  assign n37484 = ~controllable_hgrant6 & ~n37483;
  assign n37485 = ~n14019 & ~n37484;
  assign n37486 = ~controllable_hmaster0 & ~n37485;
  assign n37487 = ~n31225 & ~n37486;
  assign n37488 = i_hlock8 & ~n37487;
  assign n37489 = i_hbusreq6 & ~n37426;
  assign n37490 = ~controllable_hmaster2 & ~n31516;
  assign n37491 = ~n31426 & ~n37490;
  assign n37492 = ~controllable_hmaster1 & ~n37491;
  assign n37493 = ~n31425 & ~n37492;
  assign n37494 = ~i_hbusreq6 & ~n37493;
  assign n37495 = ~n37489 & ~n37494;
  assign n37496 = ~controllable_hgrant6 & ~n37495;
  assign n37497 = ~n14054 & ~n37496;
  assign n37498 = ~controllable_hmaster0 & ~n37497;
  assign n37499 = ~n31447 & ~n37498;
  assign n37500 = ~i_hlock8 & ~n37499;
  assign n37501 = ~n37488 & ~n37500;
  assign n37502 = ~i_hbusreq8 & ~n37501;
  assign n37503 = ~n37476 & ~n37502;
  assign n37504 = controllable_hmaster3 & ~n37503;
  assign n37505 = i_hbusreq8 & ~n37450;
  assign n37506 = i_hbusreq6 & ~n37436;
  assign n37507 = ~n31309 & ~n31344;
  assign n37508 = controllable_hmaster1 & ~n37507;
  assign n37509 = ~n31336 & ~n37508;
  assign n37510 = ~i_hbusreq6 & ~n37509;
  assign n37511 = ~n37506 & ~n37510;
  assign n37512 = ~controllable_hgrant6 & ~n37511;
  assign n37513 = ~n14094 & ~n37512;
  assign n37514 = controllable_hmaster0 & ~n37513;
  assign n37515 = ~n31403 & ~n37514;
  assign n37516 = i_hlock8 & ~n37515;
  assign n37517 = i_hbusreq6 & ~n37444;
  assign n37518 = ~n31531 & ~n31566;
  assign n37519 = controllable_hmaster1 & ~n37518;
  assign n37520 = ~n31558 & ~n37519;
  assign n37521 = ~i_hbusreq6 & ~n37520;
  assign n37522 = ~n37517 & ~n37521;
  assign n37523 = ~controllable_hgrant6 & ~n37522;
  assign n37524 = ~n14094 & ~n37523;
  assign n37525 = controllable_hmaster0 & ~n37524;
  assign n37526 = ~n31625 & ~n37525;
  assign n37527 = ~i_hlock8 & ~n37526;
  assign n37528 = ~n37516 & ~n37527;
  assign n37529 = ~i_hbusreq8 & ~n37528;
  assign n37530 = ~n37505 & ~n37529;
  assign n37531 = ~controllable_hmaster3 & ~n37530;
  assign n37532 = ~n37504 & ~n37531;
  assign n37533 = i_hlock7 & ~n37532;
  assign n37534 = i_hbusreq8 & ~n37470;
  assign n37535 = i_hbusreq6 & ~n37456;
  assign n37536 = ~n31309 & ~n31393;
  assign n37537 = controllable_hmaster1 & ~n37536;
  assign n37538 = ~n31336 & ~n37537;
  assign n37539 = ~i_hbusreq6 & ~n37538;
  assign n37540 = ~n37535 & ~n37539;
  assign n37541 = ~controllable_hgrant6 & ~n37540;
  assign n37542 = ~n14298 & ~n37541;
  assign n37543 = controllable_hmaster0 & ~n37542;
  assign n37544 = ~n31403 & ~n37543;
  assign n37545 = i_hlock8 & ~n37544;
  assign n37546 = i_hbusreq6 & ~n37464;
  assign n37547 = ~n31531 & ~n31615;
  assign n37548 = controllable_hmaster1 & ~n37547;
  assign n37549 = ~n31558 & ~n37548;
  assign n37550 = ~i_hbusreq6 & ~n37549;
  assign n37551 = ~n37546 & ~n37550;
  assign n37552 = ~controllable_hgrant6 & ~n37551;
  assign n37553 = ~n14298 & ~n37552;
  assign n37554 = controllable_hmaster0 & ~n37553;
  assign n37555 = ~n31625 & ~n37554;
  assign n37556 = ~i_hlock8 & ~n37555;
  assign n37557 = ~n37545 & ~n37556;
  assign n37558 = ~i_hbusreq8 & ~n37557;
  assign n37559 = ~n37534 & ~n37558;
  assign n37560 = ~controllable_hmaster3 & ~n37559;
  assign n37561 = ~n37504 & ~n37560;
  assign n37562 = ~i_hlock7 & ~n37561;
  assign n37563 = ~n37533 & ~n37562;
  assign n37564 = ~i_hbusreq7 & ~n37563;
  assign n37565 = ~n37475 & ~n37564;
  assign n37566 = n7924 & ~n37565;
  assign n37567 = ~n37062 & ~n37566;
  assign n37568 = ~n8214 & ~n37567;
  assign n37569 = ~n37309 & ~n37568;
  assign n37570 = ~n8202 & ~n37569;
  assign n37571 = ~n31650 & ~n37420;
  assign n37572 = i_hlock8 & ~n37571;
  assign n37573 = ~n31683 & ~n37429;
  assign n37574 = ~i_hlock8 & ~n37573;
  assign n37575 = ~n37572 & ~n37574;
  assign n37576 = controllable_hmaster3 & ~n37575;
  assign n37577 = ~n30307 & ~n31021;
  assign n37578 = controllable_hmaster1 & ~n37577;
  assign n37579 = ~n31036 & ~n37578;
  assign n37580 = ~controllable_hgrant6 & ~n37579;
  assign n37581 = ~n13849 & ~n37580;
  assign n37582 = controllable_hmaster0 & ~n37581;
  assign n37583 = ~n31074 & ~n37582;
  assign n37584 = i_hlock8 & ~n37583;
  assign n37585 = ~n30410 & ~n31128;
  assign n37586 = controllable_hmaster1 & ~n37585;
  assign n37587 = ~n31143 & ~n37586;
  assign n37588 = ~controllable_hgrant6 & ~n37587;
  assign n37589 = ~n13849 & ~n37588;
  assign n37590 = controllable_hmaster0 & ~n37589;
  assign n37591 = ~n31181 & ~n37590;
  assign n37592 = ~i_hlock8 & ~n37591;
  assign n37593 = ~n37584 & ~n37592;
  assign n37594 = ~controllable_hmaster3 & ~n37593;
  assign n37595 = ~n37576 & ~n37594;
  assign n37596 = i_hlock7 & ~n37595;
  assign n37597 = ~n30332 & ~n31021;
  assign n37598 = controllable_hmaster1 & ~n37597;
  assign n37599 = ~n31036 & ~n37598;
  assign n37600 = ~controllable_hgrant6 & ~n37599;
  assign n37601 = ~n13951 & ~n37600;
  assign n37602 = controllable_hmaster0 & ~n37601;
  assign n37603 = ~n31074 & ~n37602;
  assign n37604 = i_hlock8 & ~n37603;
  assign n37605 = ~n30435 & ~n31128;
  assign n37606 = controllable_hmaster1 & ~n37605;
  assign n37607 = ~n31143 & ~n37606;
  assign n37608 = ~controllable_hgrant6 & ~n37607;
  assign n37609 = ~n13951 & ~n37608;
  assign n37610 = controllable_hmaster0 & ~n37609;
  assign n37611 = ~n31181 & ~n37610;
  assign n37612 = ~i_hlock8 & ~n37611;
  assign n37613 = ~n37604 & ~n37612;
  assign n37614 = ~controllable_hmaster3 & ~n37613;
  assign n37615 = ~n37576 & ~n37614;
  assign n37616 = ~i_hlock7 & ~n37615;
  assign n37617 = ~n37596 & ~n37616;
  assign n37618 = i_hbusreq7 & ~n37617;
  assign n37619 = i_hbusreq8 & ~n37575;
  assign n37620 = ~n31731 & ~n37486;
  assign n37621 = i_hlock8 & ~n37620;
  assign n37622 = ~n31807 & ~n37498;
  assign n37623 = ~i_hlock8 & ~n37622;
  assign n37624 = ~n37621 & ~n37623;
  assign n37625 = ~i_hbusreq8 & ~n37624;
  assign n37626 = ~n37619 & ~n37625;
  assign n37627 = controllable_hmaster3 & ~n37626;
  assign n37628 = i_hbusreq8 & ~n37593;
  assign n37629 = i_hbusreq6 & ~n37579;
  assign n37630 = ~n31309 & ~n31923;
  assign n37631 = controllable_hmaster1 & ~n37630;
  assign n37632 = ~n31336 & ~n37631;
  assign n37633 = ~i_hbusreq6 & ~n37632;
  assign n37634 = ~n37629 & ~n37633;
  assign n37635 = ~controllable_hgrant6 & ~n37634;
  assign n37636 = ~n14756 & ~n37635;
  assign n37637 = controllable_hmaster0 & ~n37636;
  assign n37638 = ~n31403 & ~n37637;
  assign n37639 = i_hlock8 & ~n37638;
  assign n37640 = i_hbusreq6 & ~n37587;
  assign n37641 = ~n31531 & ~n31956;
  assign n37642 = controllable_hmaster1 & ~n37641;
  assign n37643 = ~n31558 & ~n37642;
  assign n37644 = ~i_hbusreq6 & ~n37643;
  assign n37645 = ~n37640 & ~n37644;
  assign n37646 = ~controllable_hgrant6 & ~n37645;
  assign n37647 = ~n14756 & ~n37646;
  assign n37648 = controllable_hmaster0 & ~n37647;
  assign n37649 = ~n31625 & ~n37648;
  assign n37650 = ~i_hlock8 & ~n37649;
  assign n37651 = ~n37639 & ~n37650;
  assign n37652 = ~i_hbusreq8 & ~n37651;
  assign n37653 = ~n37628 & ~n37652;
  assign n37654 = ~controllable_hmaster3 & ~n37653;
  assign n37655 = ~n37627 & ~n37654;
  assign n37656 = i_hlock7 & ~n37655;
  assign n37657 = i_hbusreq8 & ~n37613;
  assign n37658 = i_hbusreq6 & ~n37599;
  assign n37659 = ~n31309 & ~n31928;
  assign n37660 = controllable_hmaster1 & ~n37659;
  assign n37661 = ~n31336 & ~n37660;
  assign n37662 = ~i_hbusreq6 & ~n37661;
  assign n37663 = ~n37658 & ~n37662;
  assign n37664 = ~controllable_hgrant6 & ~n37663;
  assign n37665 = ~n14772 & ~n37664;
  assign n37666 = controllable_hmaster0 & ~n37665;
  assign n37667 = ~n31403 & ~n37666;
  assign n37668 = i_hlock8 & ~n37667;
  assign n37669 = i_hbusreq6 & ~n37607;
  assign n37670 = ~n31531 & ~n31961;
  assign n37671 = controllable_hmaster1 & ~n37670;
  assign n37672 = ~n31558 & ~n37671;
  assign n37673 = ~i_hbusreq6 & ~n37672;
  assign n37674 = ~n37669 & ~n37673;
  assign n37675 = ~controllable_hgrant6 & ~n37674;
  assign n37676 = ~n14772 & ~n37675;
  assign n37677 = controllable_hmaster0 & ~n37676;
  assign n37678 = ~n31625 & ~n37677;
  assign n37679 = ~i_hlock8 & ~n37678;
  assign n37680 = ~n37668 & ~n37679;
  assign n37681 = ~i_hbusreq8 & ~n37680;
  assign n37682 = ~n37657 & ~n37681;
  assign n37683 = ~controllable_hmaster3 & ~n37682;
  assign n37684 = ~n37627 & ~n37683;
  assign n37685 = ~i_hlock7 & ~n37684;
  assign n37686 = ~n37656 & ~n37685;
  assign n37687 = ~i_hbusreq7 & ~n37686;
  assign n37688 = ~n37618 & ~n37687;
  assign n37689 = n7924 & ~n37688;
  assign n37690 = ~n37340 & ~n37689;
  assign n37691 = ~n8214 & ~n37690;
  assign n37692 = ~n31883 & ~n37439;
  assign n37693 = i_hlock8 & ~n37692;
  assign n37694 = ~n31905 & ~n37447;
  assign n37695 = ~i_hlock8 & ~n37694;
  assign n37696 = ~n37693 & ~n37695;
  assign n37697 = ~controllable_hmaster3 & ~n37696;
  assign n37698 = ~n37576 & ~n37697;
  assign n37699 = i_hlock7 & ~n37698;
  assign n37700 = ~n31883 & ~n37459;
  assign n37701 = i_hlock8 & ~n37700;
  assign n37702 = ~n31905 & ~n37467;
  assign n37703 = ~i_hlock8 & ~n37702;
  assign n37704 = ~n37701 & ~n37703;
  assign n37705 = ~controllable_hmaster3 & ~n37704;
  assign n37706 = ~n37576 & ~n37705;
  assign n37707 = ~i_hlock7 & ~n37706;
  assign n37708 = ~n37699 & ~n37707;
  assign n37709 = i_hbusreq7 & ~n37708;
  assign n37710 = i_hbusreq8 & ~n37696;
  assign n37711 = ~n31938 & ~n37514;
  assign n37712 = i_hlock8 & ~n37711;
  assign n37713 = ~n31971 & ~n37525;
  assign n37714 = ~i_hlock8 & ~n37713;
  assign n37715 = ~n37712 & ~n37714;
  assign n37716 = ~i_hbusreq8 & ~n37715;
  assign n37717 = ~n37710 & ~n37716;
  assign n37718 = ~controllable_hmaster3 & ~n37717;
  assign n37719 = ~n37627 & ~n37718;
  assign n37720 = i_hlock7 & ~n37719;
  assign n37721 = i_hbusreq8 & ~n37704;
  assign n37722 = ~n31938 & ~n37543;
  assign n37723 = i_hlock8 & ~n37722;
  assign n37724 = ~n31971 & ~n37554;
  assign n37725 = ~i_hlock8 & ~n37724;
  assign n37726 = ~n37723 & ~n37725;
  assign n37727 = ~i_hbusreq8 & ~n37726;
  assign n37728 = ~n37721 & ~n37727;
  assign n37729 = ~controllable_hmaster3 & ~n37728;
  assign n37730 = ~n37627 & ~n37729;
  assign n37731 = ~i_hlock7 & ~n37730;
  assign n37732 = ~n37720 & ~n37731;
  assign n37733 = ~i_hbusreq7 & ~n37732;
  assign n37734 = ~n37709 & ~n37733;
  assign n37735 = n7924 & ~n37734;
  assign n37736 = ~n37385 & ~n37735;
  assign n37737 = n8214 & ~n37736;
  assign n37738 = ~n37691 & ~n37737;
  assign n37739 = n8202 & ~n37738;
  assign n37740 = ~n37570 & ~n37739;
  assign n37741 = n7920 & ~n37740;
  assign n37742 = ~n36523 & ~n37741;
  assign n37743 = n7728 & ~n37742;
  assign n37744 = ~n21649 & ~n36559;
  assign n37745 = ~controllable_hmaster1 & ~n37744;
  assign n37746 = ~n21648 & ~n37745;
  assign n37747 = ~i_hbusreq6 & ~n37746;
  assign n37748 = ~n36850 & ~n37747;
  assign n37749 = ~controllable_hgrant6 & ~n37748;
  assign n37750 = ~n14927 & ~n37749;
  assign n37751 = ~controllable_hmaster0 & ~n37750;
  assign n37752 = ~n31997 & ~n37751;
  assign n37753 = i_hlock8 & ~n37752;
  assign n37754 = ~n21649 & ~n36571;
  assign n37755 = ~controllable_hmaster1 & ~n37754;
  assign n37756 = ~n21648 & ~n37755;
  assign n37757 = ~i_hbusreq6 & ~n37756;
  assign n37758 = ~n36861 & ~n37757;
  assign n37759 = ~controllable_hgrant6 & ~n37758;
  assign n37760 = ~n14960 & ~n37759;
  assign n37761 = ~controllable_hmaster0 & ~n37760;
  assign n37762 = ~n31997 & ~n37761;
  assign n37763 = ~i_hlock8 & ~n37762;
  assign n37764 = ~n37753 & ~n37763;
  assign n37765 = ~i_hbusreq8 & ~n37764;
  assign n37766 = ~n37140 & ~n37765;
  assign n37767 = controllable_hmaster3 & ~n37766;
  assign n37768 = ~n21813 & ~n37767;
  assign n37769 = i_hlock7 & ~n37768;
  assign n37770 = ~n21827 & ~n37767;
  assign n37771 = ~i_hlock7 & ~n37770;
  assign n37772 = ~n37769 & ~n37771;
  assign n37773 = ~i_hbusreq7 & ~n37772;
  assign n37774 = ~n37139 & ~n37773;
  assign n37775 = ~n7924 & ~n37774;
  assign n37776 = ~n32049 & ~n36627;
  assign n37777 = ~controllable_hmaster1 & ~n37776;
  assign n37778 = ~n32048 & ~n37777;
  assign n37779 = ~i_hbusreq6 & ~n37778;
  assign n37780 = ~n36908 & ~n37779;
  assign n37781 = ~controllable_hgrant6 & ~n37780;
  assign n37782 = ~n14927 & ~n37781;
  assign n37783 = ~controllable_hmaster0 & ~n37782;
  assign n37784 = ~n32070 & ~n37783;
  assign n37785 = i_hlock8 & ~n37784;
  assign n37786 = ~n32226 & ~n36642;
  assign n37787 = ~controllable_hmaster1 & ~n37786;
  assign n37788 = ~n32225 & ~n37787;
  assign n37789 = ~i_hbusreq6 & ~n37788;
  assign n37790 = ~n36920 & ~n37789;
  assign n37791 = ~controllable_hgrant6 & ~n37790;
  assign n37792 = ~n14960 & ~n37791;
  assign n37793 = ~controllable_hmaster0 & ~n37792;
  assign n37794 = ~n32247 & ~n37793;
  assign n37795 = ~i_hlock8 & ~n37794;
  assign n37796 = ~n37785 & ~n37795;
  assign n37797 = ~i_hbusreq8 & ~n37796;
  assign n37798 = ~n37221 & ~n37797;
  assign n37799 = controllable_hmaster3 & ~n37798;
  assign n37800 = ~n32127 & ~n32157;
  assign n37801 = controllable_hmaster1 & ~n37800;
  assign n37802 = ~n32150 & ~n37801;
  assign n37803 = ~i_hbusreq6 & ~n37802;
  assign n37804 = ~n37247 & ~n37803;
  assign n37805 = ~controllable_hgrant6 & ~n37804;
  assign n37806 = ~n14995 & ~n37805;
  assign n37807 = controllable_hmaster0 & ~n37806;
  assign n37808 = ~n32208 & ~n37807;
  assign n37809 = i_hlock8 & ~n37808;
  assign n37810 = ~n32304 & ~n32334;
  assign n37811 = controllable_hmaster1 & ~n37810;
  assign n37812 = ~n32327 & ~n37811;
  assign n37813 = ~i_hbusreq6 & ~n37812;
  assign n37814 = ~n37258 & ~n37813;
  assign n37815 = ~controllable_hgrant6 & ~n37814;
  assign n37816 = ~n14995 & ~n37815;
  assign n37817 = controllable_hmaster0 & ~n37816;
  assign n37818 = ~n32385 & ~n37817;
  assign n37819 = ~i_hlock8 & ~n37818;
  assign n37820 = ~n37809 & ~n37819;
  assign n37821 = ~i_hbusreq8 & ~n37820;
  assign n37822 = ~n37246 & ~n37821;
  assign n37823 = ~controllable_hmaster3 & ~n37822;
  assign n37824 = ~n37799 & ~n37823;
  assign n37825 = i_hlock7 & ~n37824;
  assign n37826 = ~n32127 & ~n32198;
  assign n37827 = controllable_hmaster1 & ~n37826;
  assign n37828 = ~n32150 & ~n37827;
  assign n37829 = ~i_hbusreq6 & ~n37828;
  assign n37830 = ~n37276 & ~n37829;
  assign n37831 = ~controllable_hgrant6 & ~n37830;
  assign n37832 = ~n15152 & ~n37831;
  assign n37833 = controllable_hmaster0 & ~n37832;
  assign n37834 = ~n32208 & ~n37833;
  assign n37835 = i_hlock8 & ~n37834;
  assign n37836 = ~n32304 & ~n32375;
  assign n37837 = controllable_hmaster1 & ~n37836;
  assign n37838 = ~n32327 & ~n37837;
  assign n37839 = ~i_hbusreq6 & ~n37838;
  assign n37840 = ~n37287 & ~n37839;
  assign n37841 = ~controllable_hgrant6 & ~n37840;
  assign n37842 = ~n15152 & ~n37841;
  assign n37843 = controllable_hmaster0 & ~n37842;
  assign n37844 = ~n32385 & ~n37843;
  assign n37845 = ~i_hlock8 & ~n37844;
  assign n37846 = ~n37835 & ~n37845;
  assign n37847 = ~i_hbusreq8 & ~n37846;
  assign n37848 = ~n37275 & ~n37847;
  assign n37849 = ~controllable_hmaster3 & ~n37848;
  assign n37850 = ~n37799 & ~n37849;
  assign n37851 = ~i_hlock7 & ~n37850;
  assign n37852 = ~n37825 & ~n37851;
  assign n37853 = ~i_hbusreq7 & ~n37852;
  assign n37854 = ~n37220 & ~n37853;
  assign n37855 = n7924 & ~n37854;
  assign n37856 = ~n37775 & ~n37855;
  assign n37857 = n7920 & ~n37856;
  assign n37858 = ~n36523 & ~n37857;
  assign n37859 = ~n7728 & ~n37858;
  assign n37860 = ~n37743 & ~n37859;
  assign n37861 = ~n7723 & ~n37860;
  assign n37862 = ~n37413 & ~n37861;
  assign n37863 = ~n7714 & ~n37862;
  assign n37864 = ~n37412 & ~n37863;
  assign n37865 = ~n7705 & ~n37864;
  assign n37866 = ~n36798 & ~n37865;
  assign n37867 = n7808 & ~n37866;
  assign n37868 = ~n36533 & ~n37867;
  assign n37869 = n8195 & ~n37868;
  assign n37870 = ~n8196 & ~n37869;
  assign n37871 = ~n8193 & ~n37870;
  assign n37872 = ~n9900 & ~n36523;
  assign n37873 = ~n7723 & ~n37872;
  assign n37874 = ~n9899 & ~n37873;
  assign n37875 = n7714 & ~n37874;
  assign n37876 = ~n36529 & ~n37875;
  assign n37877 = ~n7705 & ~n37876;
  assign n37878 = ~n9898 & ~n37877;
  assign n37879 = ~n7808 & ~n37878;
  assign n37880 = ~n22407 & ~n35563;
  assign n37881 = i_hbusreq7 & ~n37880;
  assign n37882 = ~n22423 & ~n35574;
  assign n37883 = ~i_hbusreq7 & ~n37882;
  assign n37884 = ~n37881 & ~n37883;
  assign n37885 = ~n7924 & ~n37884;
  assign n37886 = ~n22441 & ~n35584;
  assign n37887 = i_hbusreq7 & ~n37886;
  assign n37888 = ~n22466 & ~n35595;
  assign n37889 = ~i_hbusreq7 & ~n37888;
  assign n37890 = ~n37887 & ~n37889;
  assign n37891 = n7924 & ~n37890;
  assign n37892 = ~n37885 & ~n37891;
  assign n37893 = ~n8214 & ~n37892;
  assign n37894 = ~n22480 & ~n35563;
  assign n37895 = i_hbusreq7 & ~n37894;
  assign n37896 = ~n22496 & ~n35574;
  assign n37897 = ~i_hbusreq7 & ~n37896;
  assign n37898 = ~n37895 & ~n37897;
  assign n37899 = ~n7924 & ~n37898;
  assign n37900 = ~n22516 & ~n35584;
  assign n37901 = i_hbusreq7 & ~n37900;
  assign n37902 = ~n22546 & ~n35595;
  assign n37903 = ~i_hbusreq7 & ~n37902;
  assign n37904 = ~n37901 & ~n37903;
  assign n37905 = n7924 & ~n37904;
  assign n37906 = ~n37899 & ~n37905;
  assign n37907 = n8214 & ~n37906;
  assign n37908 = ~n37893 & ~n37907;
  assign n37909 = ~n8202 & ~n37908;
  assign n37910 = ~n22562 & ~n35563;
  assign n37911 = i_hbusreq7 & ~n37910;
  assign n37912 = ~n22578 & ~n35574;
  assign n37913 = ~i_hbusreq7 & ~n37912;
  assign n37914 = ~n37911 & ~n37913;
  assign n37915 = ~n7924 & ~n37914;
  assign n37916 = ~n22600 & ~n35584;
  assign n37917 = i_hbusreq7 & ~n37916;
  assign n37918 = ~n22638 & ~n35595;
  assign n37919 = ~i_hbusreq7 & ~n37918;
  assign n37920 = ~n37917 & ~n37919;
  assign n37921 = n7924 & ~n37920;
  assign n37922 = ~n37915 & ~n37921;
  assign n37923 = ~n8214 & ~n37922;
  assign n37924 = ~n22652 & ~n35563;
  assign n37925 = i_hbusreq7 & ~n37924;
  assign n37926 = ~n22668 & ~n35574;
  assign n37927 = ~i_hbusreq7 & ~n37926;
  assign n37928 = ~n37925 & ~n37927;
  assign n37929 = ~n7924 & ~n37928;
  assign n37930 = ~n22690 & ~n35584;
  assign n37931 = i_hbusreq7 & ~n37930;
  assign n37932 = ~n22731 & ~n35595;
  assign n37933 = ~i_hbusreq7 & ~n37932;
  assign n37934 = ~n37931 & ~n37933;
  assign n37935 = n7924 & ~n37934;
  assign n37936 = ~n37929 & ~n37935;
  assign n37937 = n8214 & ~n37936;
  assign n37938 = ~n37923 & ~n37937;
  assign n37939 = n8202 & ~n37938;
  assign n37940 = ~n37909 & ~n37939;
  assign n37941 = n7920 & ~n37940;
  assign n37942 = ~n10014 & ~n37941;
  assign n37943 = n7728 & ~n37942;
  assign n37944 = ~n22751 & ~n37317;
  assign n37945 = i_hlock7 & ~n37944;
  assign n37946 = ~n22759 & ~n37317;
  assign n37947 = ~i_hlock7 & ~n37946;
  assign n37948 = ~n37945 & ~n37947;
  assign n37949 = i_hbusreq7 & ~n37948;
  assign n37950 = ~n22777 & ~n37332;
  assign n37951 = i_hlock7 & ~n37950;
  assign n37952 = ~n22791 & ~n37332;
  assign n37953 = ~i_hlock7 & ~n37952;
  assign n37954 = ~n37951 & ~n37953;
  assign n37955 = ~i_hbusreq7 & ~n37954;
  assign n37956 = ~n37949 & ~n37955;
  assign n37957 = ~n7924 & ~n37956;
  assign n37958 = ~n22811 & ~n37346;
  assign n37959 = i_hlock7 & ~n37958;
  assign n37960 = ~n22819 & ~n37346;
  assign n37961 = ~i_hlock7 & ~n37960;
  assign n37962 = ~n37959 & ~n37961;
  assign n37963 = i_hbusreq7 & ~n37962;
  assign n37964 = ~n22846 & ~n37361;
  assign n37965 = i_hlock7 & ~n37964;
  assign n37966 = ~n22860 & ~n37361;
  assign n37967 = ~i_hlock7 & ~n37966;
  assign n37968 = ~n37965 & ~n37967;
  assign n37969 = ~i_hbusreq7 & ~n37968;
  assign n37970 = ~n37963 & ~n37969;
  assign n37971 = n7924 & ~n37970;
  assign n37972 = ~n37957 & ~n37971;
  assign n37973 = ~n8214 & ~n37972;
  assign n37974 = ~n22880 & ~n37317;
  assign n37975 = i_hlock7 & ~n37974;
  assign n37976 = ~n22884 & ~n37317;
  assign n37977 = ~i_hlock7 & ~n37976;
  assign n37978 = ~n37975 & ~n37977;
  assign n37979 = i_hbusreq7 & ~n37978;
  assign n37980 = ~n22906 & ~n37332;
  assign n37981 = i_hlock7 & ~n37980;
  assign n37982 = ~n22913 & ~n37332;
  assign n37983 = ~i_hlock7 & ~n37982;
  assign n37984 = ~n37981 & ~n37983;
  assign n37985 = ~i_hbusreq7 & ~n37984;
  assign n37986 = ~n37979 & ~n37985;
  assign n37987 = ~n7924 & ~n37986;
  assign n37988 = ~n22939 & ~n37346;
  assign n37989 = i_hlock7 & ~n37988;
  assign n37990 = ~n22943 & ~n37346;
  assign n37991 = ~i_hlock7 & ~n37990;
  assign n37992 = ~n37989 & ~n37991;
  assign n37993 = i_hbusreq7 & ~n37992;
  assign n37994 = ~n22979 & ~n37361;
  assign n37995 = i_hlock7 & ~n37994;
  assign n37996 = ~n22986 & ~n37361;
  assign n37997 = ~i_hlock7 & ~n37996;
  assign n37998 = ~n37995 & ~n37997;
  assign n37999 = ~i_hbusreq7 & ~n37998;
  assign n38000 = ~n37993 & ~n37999;
  assign n38001 = n7924 & ~n38000;
  assign n38002 = ~n37987 & ~n38001;
  assign n38003 = n8214 & ~n38002;
  assign n38004 = ~n37973 & ~n38003;
  assign n38005 = ~n8202 & ~n38004;
  assign n38006 = ~n23004 & ~n37317;
  assign n38007 = i_hlock7 & ~n38006;
  assign n38008 = ~n23014 & ~n37317;
  assign n38009 = ~i_hlock7 & ~n38008;
  assign n38010 = ~n38007 & ~n38009;
  assign n38011 = i_hbusreq7 & ~n38010;
  assign n38012 = ~n23032 & ~n37332;
  assign n38013 = i_hlock7 & ~n38012;
  assign n38014 = ~n23048 & ~n37332;
  assign n38015 = ~i_hlock7 & ~n38014;
  assign n38016 = ~n38013 & ~n38015;
  assign n38017 = ~i_hbusreq7 & ~n38016;
  assign n38018 = ~n38011 & ~n38017;
  assign n38019 = ~n7924 & ~n38018;
  assign n38020 = ~n23072 & ~n37346;
  assign n38021 = i_hlock7 & ~n38020;
  assign n38022 = ~n23082 & ~n37346;
  assign n38023 = ~i_hlock7 & ~n38022;
  assign n38024 = ~n38021 & ~n38023;
  assign n38025 = i_hbusreq7 & ~n38024;
  assign n38026 = ~n23122 & ~n37361;
  assign n38027 = i_hlock7 & ~n38026;
  assign n38028 = ~n23138 & ~n37361;
  assign n38029 = ~i_hlock7 & ~n38028;
  assign n38030 = ~n38027 & ~n38029;
  assign n38031 = ~i_hbusreq7 & ~n38030;
  assign n38032 = ~n38025 & ~n38031;
  assign n38033 = n7924 & ~n38032;
  assign n38034 = ~n38019 & ~n38033;
  assign n38035 = ~n8214 & ~n38034;
  assign n38036 = ~n23160 & ~n37317;
  assign n38037 = i_hlock7 & ~n38036;
  assign n38038 = ~n23164 & ~n37317;
  assign n38039 = ~i_hlock7 & ~n38038;
  assign n38040 = ~n38037 & ~n38039;
  assign n38041 = i_hbusreq7 & ~n38040;
  assign n38042 = ~n23188 & ~n37332;
  assign n38043 = i_hlock7 & ~n38042;
  assign n38044 = ~n23195 & ~n37332;
  assign n38045 = ~i_hlock7 & ~n38044;
  assign n38046 = ~n38043 & ~n38045;
  assign n38047 = ~i_hbusreq7 & ~n38046;
  assign n38048 = ~n38041 & ~n38047;
  assign n38049 = ~n7924 & ~n38048;
  assign n38050 = ~n23225 & ~n37346;
  assign n38051 = i_hlock7 & ~n38050;
  assign n38052 = ~n23229 & ~n37346;
  assign n38053 = ~i_hlock7 & ~n38052;
  assign n38054 = ~n38051 & ~n38053;
  assign n38055 = i_hbusreq7 & ~n38054;
  assign n38056 = ~n23278 & ~n37361;
  assign n38057 = i_hlock7 & ~n38056;
  assign n38058 = ~n23285 & ~n37361;
  assign n38059 = ~i_hlock7 & ~n38058;
  assign n38060 = ~n38057 & ~n38059;
  assign n38061 = ~i_hbusreq7 & ~n38060;
  assign n38062 = ~n38055 & ~n38061;
  assign n38063 = n7924 & ~n38062;
  assign n38064 = ~n38049 & ~n38063;
  assign n38065 = n8214 & ~n38064;
  assign n38066 = ~n38035 & ~n38065;
  assign n38067 = n8202 & ~n38066;
  assign n38068 = ~n38005 & ~n38067;
  assign n38069 = n7920 & ~n38068;
  assign n38070 = ~n10014 & ~n38069;
  assign n38071 = ~n7728 & ~n38070;
  assign n38072 = ~n37943 & ~n38071;
  assign n38073 = n7723 & ~n38072;
  assign n38074 = ~n7723 & ~n38070;
  assign n38075 = ~n38073 & ~n38074;
  assign n38076 = n7714 & ~n38075;
  assign n38077 = n7723 & ~n38070;
  assign n38078 = ~n32943 & ~n37435;
  assign n38079 = ~controllable_hgrant6 & ~n38078;
  assign n38080 = ~n13849 & ~n38079;
  assign n38081 = controllable_hmaster0 & ~n38080;
  assign n38082 = ~n31074 & ~n38081;
  assign n38083 = i_hlock8 & ~n38082;
  assign n38084 = ~n32953 & ~n37443;
  assign n38085 = ~controllable_hgrant6 & ~n38084;
  assign n38086 = ~n13849 & ~n38085;
  assign n38087 = controllable_hmaster0 & ~n38086;
  assign n38088 = ~n31181 & ~n38087;
  assign n38089 = ~i_hlock8 & ~n38088;
  assign n38090 = ~n38083 & ~n38089;
  assign n38091 = ~controllable_hmaster3 & ~n38090;
  assign n38092 = ~n37576 & ~n38091;
  assign n38093 = i_hlock7 & ~n38092;
  assign n38094 = ~n32943 & ~n37455;
  assign n38095 = ~controllable_hgrant6 & ~n38094;
  assign n38096 = ~n13951 & ~n38095;
  assign n38097 = controllable_hmaster0 & ~n38096;
  assign n38098 = ~n31074 & ~n38097;
  assign n38099 = i_hlock8 & ~n38098;
  assign n38100 = ~n32953 & ~n37463;
  assign n38101 = ~controllable_hgrant6 & ~n38100;
  assign n38102 = ~n13951 & ~n38101;
  assign n38103 = controllable_hmaster0 & ~n38102;
  assign n38104 = ~n31181 & ~n38103;
  assign n38105 = ~i_hlock8 & ~n38104;
  assign n38106 = ~n38099 & ~n38105;
  assign n38107 = ~controllable_hmaster3 & ~n38106;
  assign n38108 = ~n37576 & ~n38107;
  assign n38109 = ~i_hlock7 & ~n38108;
  assign n38110 = ~n38093 & ~n38109;
  assign n38111 = i_hbusreq7 & ~n38110;
  assign n38112 = i_hbusreq8 & ~n38090;
  assign n38113 = i_hbusreq6 & ~n38078;
  assign n38114 = ~n32975 & ~n37508;
  assign n38115 = ~i_hbusreq6 & ~n38114;
  assign n38116 = ~n38113 & ~n38115;
  assign n38117 = ~controllable_hgrant6 & ~n38116;
  assign n38118 = ~n15417 & ~n38117;
  assign n38119 = controllable_hmaster0 & ~n38118;
  assign n38120 = ~n31403 & ~n38119;
  assign n38121 = i_hlock8 & ~n38120;
  assign n38122 = i_hbusreq6 & ~n38084;
  assign n38123 = ~n32999 & ~n37519;
  assign n38124 = ~i_hbusreq6 & ~n38123;
  assign n38125 = ~n38122 & ~n38124;
  assign n38126 = ~controllable_hgrant6 & ~n38125;
  assign n38127 = ~n15417 & ~n38126;
  assign n38128 = controllable_hmaster0 & ~n38127;
  assign n38129 = ~n31625 & ~n38128;
  assign n38130 = ~i_hlock8 & ~n38129;
  assign n38131 = ~n38121 & ~n38130;
  assign n38132 = ~i_hbusreq8 & ~n38131;
  assign n38133 = ~n38112 & ~n38132;
  assign n38134 = ~controllable_hmaster3 & ~n38133;
  assign n38135 = ~n37627 & ~n38134;
  assign n38136 = i_hlock7 & ~n38135;
  assign n38137 = i_hbusreq8 & ~n38106;
  assign n38138 = i_hbusreq6 & ~n38094;
  assign n38139 = ~n32975 & ~n37537;
  assign n38140 = ~i_hbusreq6 & ~n38139;
  assign n38141 = ~n38138 & ~n38140;
  assign n38142 = ~controllable_hgrant6 & ~n38141;
  assign n38143 = ~n15440 & ~n38142;
  assign n38144 = controllable_hmaster0 & ~n38143;
  assign n38145 = ~n31403 & ~n38144;
  assign n38146 = i_hlock8 & ~n38145;
  assign n38147 = i_hbusreq6 & ~n38100;
  assign n38148 = ~n32999 & ~n37548;
  assign n38149 = ~i_hbusreq6 & ~n38148;
  assign n38150 = ~n38147 & ~n38149;
  assign n38151 = ~controllable_hgrant6 & ~n38150;
  assign n38152 = ~n15440 & ~n38151;
  assign n38153 = controllable_hmaster0 & ~n38152;
  assign n38154 = ~n31625 & ~n38153;
  assign n38155 = ~i_hlock8 & ~n38154;
  assign n38156 = ~n38146 & ~n38155;
  assign n38157 = ~i_hbusreq8 & ~n38156;
  assign n38158 = ~n38137 & ~n38157;
  assign n38159 = ~controllable_hmaster3 & ~n38158;
  assign n38160 = ~n37627 & ~n38159;
  assign n38161 = ~i_hlock7 & ~n38160;
  assign n38162 = ~n38136 & ~n38161;
  assign n38163 = ~i_hbusreq7 & ~n38162;
  assign n38164 = ~n38111 & ~n38163;
  assign n38165 = n7924 & ~n38164;
  assign n38166 = ~n37957 & ~n38165;
  assign n38167 = ~n8214 & ~n38166;
  assign n38168 = ~n33027 & ~n37439;
  assign n38169 = i_hlock8 & ~n38168;
  assign n38170 = ~n33041 & ~n37447;
  assign n38171 = ~i_hlock8 & ~n38170;
  assign n38172 = ~n38169 & ~n38171;
  assign n38173 = ~controllable_hmaster3 & ~n38172;
  assign n38174 = ~n37576 & ~n38173;
  assign n38175 = i_hlock7 & ~n38174;
  assign n38176 = ~n33027 & ~n37459;
  assign n38177 = i_hlock8 & ~n38176;
  assign n38178 = ~n33041 & ~n37467;
  assign n38179 = ~i_hlock8 & ~n38178;
  assign n38180 = ~n38177 & ~n38179;
  assign n38181 = ~controllable_hmaster3 & ~n38180;
  assign n38182 = ~n37576 & ~n38181;
  assign n38183 = ~i_hlock7 & ~n38182;
  assign n38184 = ~n38175 & ~n38183;
  assign n38185 = i_hbusreq7 & ~n38184;
  assign n38186 = i_hbusreq8 & ~n38172;
  assign n38187 = ~n33073 & ~n37514;
  assign n38188 = i_hlock8 & ~n38187;
  assign n38189 = ~n33105 & ~n37525;
  assign n38190 = ~i_hlock8 & ~n38189;
  assign n38191 = ~n38188 & ~n38190;
  assign n38192 = ~i_hbusreq8 & ~n38191;
  assign n38193 = ~n38186 & ~n38192;
  assign n38194 = ~controllable_hmaster3 & ~n38193;
  assign n38195 = ~n37627 & ~n38194;
  assign n38196 = i_hlock7 & ~n38195;
  assign n38197 = i_hbusreq8 & ~n38180;
  assign n38198 = ~n33073 & ~n37543;
  assign n38199 = i_hlock8 & ~n38198;
  assign n38200 = ~n33105 & ~n37554;
  assign n38201 = ~i_hlock8 & ~n38200;
  assign n38202 = ~n38199 & ~n38201;
  assign n38203 = ~i_hbusreq8 & ~n38202;
  assign n38204 = ~n38197 & ~n38203;
  assign n38205 = ~controllable_hmaster3 & ~n38204;
  assign n38206 = ~n37627 & ~n38205;
  assign n38207 = ~i_hlock7 & ~n38206;
  assign n38208 = ~n38196 & ~n38207;
  assign n38209 = ~i_hbusreq7 & ~n38208;
  assign n38210 = ~n38185 & ~n38209;
  assign n38211 = n7924 & ~n38210;
  assign n38212 = ~n37987 & ~n38211;
  assign n38213 = n8214 & ~n38212;
  assign n38214 = ~n38167 & ~n38213;
  assign n38215 = ~n8202 & ~n38214;
  assign n38216 = ~n30287 & ~n31041;
  assign n38217 = controllable_hmaster1 & ~n38216;
  assign n38218 = ~n31036 & ~n38217;
  assign n38219 = ~controllable_hgrant6 & ~n38218;
  assign n38220 = ~n13849 & ~n38219;
  assign n38221 = controllable_hmaster0 & ~n38220;
  assign n38222 = ~n31074 & ~n38221;
  assign n38223 = i_hlock8 & ~n38222;
  assign n38224 = ~n30390 & ~n31148;
  assign n38225 = controllable_hmaster1 & ~n38224;
  assign n38226 = ~n31143 & ~n38225;
  assign n38227 = ~controllable_hgrant6 & ~n38226;
  assign n38228 = ~n13849 & ~n38227;
  assign n38229 = controllable_hmaster0 & ~n38228;
  assign n38230 = ~n31181 & ~n38229;
  assign n38231 = ~i_hlock8 & ~n38230;
  assign n38232 = ~n38223 & ~n38231;
  assign n38233 = ~controllable_hmaster3 & ~n38232;
  assign n38234 = ~n37576 & ~n38233;
  assign n38235 = i_hlock7 & ~n38234;
  assign n38236 = ~n30287 & ~n31066;
  assign n38237 = controllable_hmaster1 & ~n38236;
  assign n38238 = ~n31036 & ~n38237;
  assign n38239 = ~controllable_hgrant6 & ~n38238;
  assign n38240 = ~n13951 & ~n38239;
  assign n38241 = controllable_hmaster0 & ~n38240;
  assign n38242 = ~n31074 & ~n38241;
  assign n38243 = i_hlock8 & ~n38242;
  assign n38244 = ~n30390 & ~n31173;
  assign n38245 = controllable_hmaster1 & ~n38244;
  assign n38246 = ~n31143 & ~n38245;
  assign n38247 = ~controllable_hgrant6 & ~n38246;
  assign n38248 = ~n13951 & ~n38247;
  assign n38249 = controllable_hmaster0 & ~n38248;
  assign n38250 = ~n31181 & ~n38249;
  assign n38251 = ~i_hlock8 & ~n38250;
  assign n38252 = ~n38243 & ~n38251;
  assign n38253 = ~controllable_hmaster3 & ~n38252;
  assign n38254 = ~n37576 & ~n38253;
  assign n38255 = ~i_hlock7 & ~n38254;
  assign n38256 = ~n38235 & ~n38255;
  assign n38257 = i_hbusreq7 & ~n38256;
  assign n38258 = i_hbusreq8 & ~n38232;
  assign n38259 = i_hbusreq6 & ~n38218;
  assign n38260 = ~n31344 & ~n33154;
  assign n38261 = controllable_hmaster1 & ~n38260;
  assign n38262 = ~n31336 & ~n38261;
  assign n38263 = ~i_hbusreq6 & ~n38262;
  assign n38264 = ~n38259 & ~n38263;
  assign n38265 = ~controllable_hgrant6 & ~n38264;
  assign n38266 = ~n15520 & ~n38265;
  assign n38267 = controllable_hmaster0 & ~n38266;
  assign n38268 = ~n31403 & ~n38267;
  assign n38269 = i_hlock8 & ~n38268;
  assign n38270 = i_hbusreq6 & ~n38226;
  assign n38271 = ~n31566 & ~n33181;
  assign n38272 = controllable_hmaster1 & ~n38271;
  assign n38273 = ~n31558 & ~n38272;
  assign n38274 = ~i_hbusreq6 & ~n38273;
  assign n38275 = ~n38270 & ~n38274;
  assign n38276 = ~controllable_hgrant6 & ~n38275;
  assign n38277 = ~n15520 & ~n38276;
  assign n38278 = controllable_hmaster0 & ~n38277;
  assign n38279 = ~n31625 & ~n38278;
  assign n38280 = ~i_hlock8 & ~n38279;
  assign n38281 = ~n38269 & ~n38280;
  assign n38282 = ~i_hbusreq8 & ~n38281;
  assign n38283 = ~n38258 & ~n38282;
  assign n38284 = ~controllable_hmaster3 & ~n38283;
  assign n38285 = ~n37627 & ~n38284;
  assign n38286 = i_hlock7 & ~n38285;
  assign n38287 = i_hbusreq8 & ~n38252;
  assign n38288 = i_hbusreq6 & ~n38238;
  assign n38289 = ~n31393 & ~n33154;
  assign n38290 = controllable_hmaster1 & ~n38289;
  assign n38291 = ~n31336 & ~n38290;
  assign n38292 = ~i_hbusreq6 & ~n38291;
  assign n38293 = ~n38288 & ~n38292;
  assign n38294 = ~controllable_hgrant6 & ~n38293;
  assign n38295 = ~n15553 & ~n38294;
  assign n38296 = controllable_hmaster0 & ~n38295;
  assign n38297 = ~n31403 & ~n38296;
  assign n38298 = i_hlock8 & ~n38297;
  assign n38299 = i_hbusreq6 & ~n38246;
  assign n38300 = ~n31615 & ~n33181;
  assign n38301 = controllable_hmaster1 & ~n38300;
  assign n38302 = ~n31558 & ~n38301;
  assign n38303 = ~i_hbusreq6 & ~n38302;
  assign n38304 = ~n38299 & ~n38303;
  assign n38305 = ~controllable_hgrant6 & ~n38304;
  assign n38306 = ~n15553 & ~n38305;
  assign n38307 = controllable_hmaster0 & ~n38306;
  assign n38308 = ~n31625 & ~n38307;
  assign n38309 = ~i_hlock8 & ~n38308;
  assign n38310 = ~n38298 & ~n38309;
  assign n38311 = ~i_hbusreq8 & ~n38310;
  assign n38312 = ~n38287 & ~n38311;
  assign n38313 = ~controllable_hmaster3 & ~n38312;
  assign n38314 = ~n37627 & ~n38313;
  assign n38315 = ~i_hlock7 & ~n38314;
  assign n38316 = ~n38286 & ~n38315;
  assign n38317 = ~i_hbusreq7 & ~n38316;
  assign n38318 = ~n38257 & ~n38317;
  assign n38319 = n7924 & ~n38318;
  assign n38320 = ~n38019 & ~n38319;
  assign n38321 = ~n8214 & ~n38320;
  assign n38322 = ~n33213 & ~n37439;
  assign n38323 = i_hlock8 & ~n38322;
  assign n38324 = ~n33229 & ~n37447;
  assign n38325 = ~i_hlock8 & ~n38324;
  assign n38326 = ~n38323 & ~n38325;
  assign n38327 = ~controllable_hmaster3 & ~n38326;
  assign n38328 = ~n37576 & ~n38327;
  assign n38329 = i_hlock7 & ~n38328;
  assign n38330 = ~n33213 & ~n37459;
  assign n38331 = i_hlock8 & ~n38330;
  assign n38332 = ~n33229 & ~n37467;
  assign n38333 = ~i_hlock8 & ~n38332;
  assign n38334 = ~n38331 & ~n38333;
  assign n38335 = ~controllable_hmaster3 & ~n38334;
  assign n38336 = ~n37576 & ~n38335;
  assign n38337 = ~i_hlock7 & ~n38336;
  assign n38338 = ~n38329 & ~n38337;
  assign n38339 = i_hbusreq7 & ~n38338;
  assign n38340 = i_hbusreq8 & ~n38326;
  assign n38341 = ~n33262 & ~n37514;
  assign n38342 = i_hlock8 & ~n38341;
  assign n38343 = ~n33295 & ~n37525;
  assign n38344 = ~i_hlock8 & ~n38343;
  assign n38345 = ~n38342 & ~n38344;
  assign n38346 = ~i_hbusreq8 & ~n38345;
  assign n38347 = ~n38340 & ~n38346;
  assign n38348 = ~controllable_hmaster3 & ~n38347;
  assign n38349 = ~n37627 & ~n38348;
  assign n38350 = i_hlock7 & ~n38349;
  assign n38351 = i_hbusreq8 & ~n38334;
  assign n38352 = ~n33262 & ~n37543;
  assign n38353 = i_hlock8 & ~n38352;
  assign n38354 = ~n33295 & ~n37554;
  assign n38355 = ~i_hlock8 & ~n38354;
  assign n38356 = ~n38353 & ~n38355;
  assign n38357 = ~i_hbusreq8 & ~n38356;
  assign n38358 = ~n38351 & ~n38357;
  assign n38359 = ~controllable_hmaster3 & ~n38358;
  assign n38360 = ~n37627 & ~n38359;
  assign n38361 = ~i_hlock7 & ~n38360;
  assign n38362 = ~n38350 & ~n38361;
  assign n38363 = ~i_hbusreq7 & ~n38362;
  assign n38364 = ~n38339 & ~n38363;
  assign n38365 = n7924 & ~n38364;
  assign n38366 = ~n38049 & ~n38365;
  assign n38367 = n8214 & ~n38366;
  assign n38368 = ~n38321 & ~n38367;
  assign n38369 = n8202 & ~n38368;
  assign n38370 = ~n38215 & ~n38369;
  assign n38371 = n7920 & ~n38370;
  assign n38372 = ~n36523 & ~n38371;
  assign n38373 = n7728 & ~n38372;
  assign n38374 = ~n37859 & ~n38373;
  assign n38375 = ~n7723 & ~n38374;
  assign n38376 = ~n38077 & ~n38375;
  assign n38377 = ~n7714 & ~n38376;
  assign n38378 = ~n38076 & ~n38377;
  assign n38379 = ~n7705 & ~n38378;
  assign n38380 = ~n22399 & ~n38379;
  assign n38381 = n7808 & ~n38380;
  assign n38382 = ~n37879 & ~n38381;
  assign n38383 = ~n8195 & ~n38382;
  assign n38384 = controllable_hgrant6 & ~n11464;
  assign n38385 = ~controllable_hmaster2 & ~n33330;
  assign n38386 = ~n10105 & ~n38385;
  assign n38387 = ~controllable_hmaster1 & ~n38386;
  assign n38388 = ~n10053 & ~n38387;
  assign n38389 = ~controllable_hgrant6 & ~n38388;
  assign n38390 = ~n38384 & ~n38389;
  assign n38391 = ~controllable_hmaster0 & ~n38390;
  assign n38392 = ~n11460 & ~n38391;
  assign n38393 = i_hlock8 & ~n38392;
  assign n38394 = controllable_hgrant6 & ~n11471;
  assign n38395 = ~controllable_hmaster2 & ~n33348;
  assign n38396 = ~n10105 & ~n38395;
  assign n38397 = ~controllable_hmaster1 & ~n38396;
  assign n38398 = ~n10053 & ~n38397;
  assign n38399 = ~controllable_hgrant6 & ~n38398;
  assign n38400 = ~n38394 & ~n38399;
  assign n38401 = ~controllable_hmaster0 & ~n38400;
  assign n38402 = ~n11460 & ~n38401;
  assign n38403 = ~i_hlock8 & ~n38402;
  assign n38404 = ~n38393 & ~n38403;
  assign n38405 = controllable_hmaster3 & ~n38404;
  assign n38406 = ~n10447 & ~n38405;
  assign n38407 = i_hbusreq7 & ~n38406;
  assign n38408 = i_hbusreq8 & ~n38404;
  assign n38409 = controllable_hgrant6 & ~n11487;
  assign n38410 = i_hbusreq6 & ~n38388;
  assign n38411 = ~controllable_hmaster2 & ~n33379;
  assign n38412 = ~n10116 & ~n38411;
  assign n38413 = ~controllable_hmaster1 & ~n38412;
  assign n38414 = ~n10064 & ~n38413;
  assign n38415 = ~i_hbusreq6 & ~n38414;
  assign n38416 = ~n38410 & ~n38415;
  assign n38417 = ~controllable_hgrant6 & ~n38416;
  assign n38418 = ~n38409 & ~n38417;
  assign n38419 = ~controllable_hmaster0 & ~n38418;
  assign n38420 = ~n11480 & ~n38419;
  assign n38421 = i_hlock8 & ~n38420;
  assign n38422 = controllable_hgrant6 & ~n11497;
  assign n38423 = i_hbusreq6 & ~n38398;
  assign n38424 = ~controllable_hmaster2 & ~n33412;
  assign n38425 = ~n10116 & ~n38424;
  assign n38426 = ~controllable_hmaster1 & ~n38425;
  assign n38427 = ~n10064 & ~n38426;
  assign n38428 = ~i_hbusreq6 & ~n38427;
  assign n38429 = ~n38423 & ~n38428;
  assign n38430 = ~controllable_hgrant6 & ~n38429;
  assign n38431 = ~n38422 & ~n38430;
  assign n38432 = ~controllable_hmaster0 & ~n38431;
  assign n38433 = ~n11480 & ~n38432;
  assign n38434 = ~i_hlock8 & ~n38433;
  assign n38435 = ~n38421 & ~n38434;
  assign n38436 = ~i_hbusreq8 & ~n38435;
  assign n38437 = ~n38408 & ~n38436;
  assign n38438 = controllable_hmaster3 & ~n38437;
  assign n38439 = ~n10621 & ~n38438;
  assign n38440 = ~i_hbusreq7 & ~n38439;
  assign n38441 = ~n38407 & ~n38440;
  assign n38442 = n7924 & ~n38441;
  assign n38443 = ~n10375 & ~n38442;
  assign n38444 = n8214 & ~n38443;
  assign n38445 = n8214 & ~n38444;
  assign n38446 = n8202 & ~n38445;
  assign n38447 = ~n10332 & ~n38446;
  assign n38448 = n7728 & ~n38447;
  assign n38449 = n8214 & ~n36522;
  assign n38450 = ~n8336 & ~n38449;
  assign n38451 = n8202 & ~n38450;
  assign n38452 = ~n10649 & ~n38451;
  assign n38453 = ~n7728 & ~n38452;
  assign n38454 = ~n38448 & ~n38453;
  assign n38455 = ~n7723 & ~n38454;
  assign n38456 = ~n7723 & ~n38455;
  assign n38457 = ~n7714 & ~n38456;
  assign n38458 = ~n7714 & ~n38457;
  assign n38459 = n7705 & ~n38458;
  assign n38460 = n7723 & ~n38452;
  assign n38461 = n7920 & ~n38452;
  assign n38462 = ~n36523 & ~n38461;
  assign n38463 = ~n7723 & ~n38462;
  assign n38464 = ~n38460 & ~n38463;
  assign n38465 = n7714 & ~n38464;
  assign n38466 = ~n36529 & ~n38465;
  assign n38467 = ~n7705 & ~n38466;
  assign n38468 = ~n38459 & ~n38467;
  assign n38469 = ~n7808 & ~n38468;
  assign n38470 = ~n7920 & ~n38447;
  assign n38471 = n7924 & ~n37855;
  assign n38472 = ~n8214 & ~n38471;
  assign n38473 = controllable_hmaster0 & ~n23853;
  assign n38474 = ~controllable_hmaster0 & ~n23847;
  assign n38475 = ~n38473 & ~n38474;
  assign n38476 = controllable_hmaster3 & ~n38475;
  assign n38477 = ~n17351 & ~n38476;
  assign n38478 = i_hbusreq7 & ~n38477;
  assign n38479 = i_hbusreq8 & ~n38475;
  assign n38480 = controllable_hmaster0 & ~n23948;
  assign n38481 = ~controllable_hmaster0 & ~n23919;
  assign n38482 = ~n38480 & ~n38481;
  assign n38483 = ~i_hbusreq8 & ~n38482;
  assign n38484 = ~n38479 & ~n38483;
  assign n38485 = controllable_hmaster3 & ~n38484;
  assign n38486 = ~n23992 & ~n38485;
  assign n38487 = ~i_hbusreq7 & ~n38486;
  assign n38488 = ~n38478 & ~n38487;
  assign n38489 = ~n7924 & ~n38488;
  assign n38490 = controllable_hmaster0 & ~n33508;
  assign n38491 = ~controllable_hmaster2 & ~n33513;
  assign n38492 = ~n33503 & ~n38491;
  assign n38493 = ~controllable_hmaster1 & ~n38492;
  assign n38494 = ~n33502 & ~n38493;
  assign n38495 = ~controllable_hgrant6 & ~n38494;
  assign n38496 = ~n13198 & ~n38495;
  assign n38497 = ~controllable_hmaster0 & ~n38496;
  assign n38498 = ~n38490 & ~n38497;
  assign n38499 = i_hlock8 & ~n38498;
  assign n38500 = controllable_hmaster0 & ~n33535;
  assign n38501 = ~controllable_hmaster2 & ~n33540;
  assign n38502 = ~n33530 & ~n38501;
  assign n38503 = ~controllable_hmaster1 & ~n38502;
  assign n38504 = ~n33529 & ~n38503;
  assign n38505 = ~controllable_hgrant6 & ~n38504;
  assign n38506 = ~n13198 & ~n38505;
  assign n38507 = ~controllable_hmaster0 & ~n38506;
  assign n38508 = ~n38500 & ~n38507;
  assign n38509 = ~i_hlock8 & ~n38508;
  assign n38510 = ~n38499 & ~n38509;
  assign n38511 = controllable_hmaster3 & ~n38510;
  assign n38512 = ~n36903 & ~n38511;
  assign n38513 = i_hbusreq7 & ~n38512;
  assign n38514 = i_hbusreq8 & ~n38510;
  assign n38515 = controllable_hmaster0 & ~n33588;
  assign n38516 = i_hbusreq6 & ~n38494;
  assign n38517 = ~controllable_hmaster2 & ~n33606;
  assign n38518 = ~n33570 & ~n38517;
  assign n38519 = ~controllable_hmaster1 & ~n38518;
  assign n38520 = ~n33569 & ~n38519;
  assign n38521 = ~i_hbusreq6 & ~n38520;
  assign n38522 = ~n38516 & ~n38521;
  assign n38523 = ~controllable_hgrant6 & ~n38522;
  assign n38524 = ~n15672 & ~n38523;
  assign n38525 = ~controllable_hmaster0 & ~n38524;
  assign n38526 = ~n38515 & ~n38525;
  assign n38527 = i_hlock8 & ~n38526;
  assign n38528 = controllable_hmaster0 & ~n33678;
  assign n38529 = i_hbusreq6 & ~n38504;
  assign n38530 = ~controllable_hmaster2 & ~n33696;
  assign n38531 = ~n33660 & ~n38530;
  assign n38532 = ~controllable_hmaster1 & ~n38531;
  assign n38533 = ~n33659 & ~n38532;
  assign n38534 = ~i_hbusreq6 & ~n38533;
  assign n38535 = ~n38529 & ~n38534;
  assign n38536 = ~controllable_hgrant6 & ~n38535;
  assign n38537 = ~n15672 & ~n38536;
  assign n38538 = ~controllable_hmaster0 & ~n38537;
  assign n38539 = ~n38528 & ~n38538;
  assign n38540 = ~i_hlock8 & ~n38539;
  assign n38541 = ~n38527 & ~n38540;
  assign n38542 = ~i_hbusreq8 & ~n38541;
  assign n38543 = ~n38514 & ~n38542;
  assign n38544 = controllable_hmaster3 & ~n38543;
  assign n38545 = ~i_hbusreq6 & ~n33580;
  assign n38546 = ~n29603 & ~n38545;
  assign n38547 = ~controllable_hgrant6 & ~n38546;
  assign n38548 = ~n15812 & ~n38547;
  assign n38549 = controllable_hmaster0 & ~n38548;
  assign n38550 = ~n33637 & ~n38549;
  assign n38551 = i_hlock8 & ~n38550;
  assign n38552 = ~i_hbusreq6 & ~n33670;
  assign n38553 = ~n29667 & ~n38552;
  assign n38554 = ~controllable_hgrant6 & ~n38553;
  assign n38555 = ~n15812 & ~n38554;
  assign n38556 = controllable_hmaster0 & ~n38555;
  assign n38557 = ~n33727 & ~n38556;
  assign n38558 = ~i_hlock8 & ~n38557;
  assign n38559 = ~n38551 & ~n38558;
  assign n38560 = ~i_hbusreq8 & ~n38559;
  assign n38561 = ~n36935 & ~n38560;
  assign n38562 = ~controllable_hmaster3 & ~n38561;
  assign n38563 = ~n38544 & ~n38562;
  assign n38564 = ~i_hbusreq7 & ~n38563;
  assign n38565 = ~n38513 & ~n38564;
  assign n38566 = n7924 & ~n38565;
  assign n38567 = ~n38489 & ~n38566;
  assign n38568 = n8214 & ~n38567;
  assign n38569 = ~n38472 & ~n38568;
  assign n38570 = n8202 & ~n38569;
  assign n38571 = ~n23818 & ~n38570;
  assign n38572 = n7920 & ~n38571;
  assign n38573 = ~n38470 & ~n38572;
  assign n38574 = n7728 & ~n38573;
  assign n38575 = ~n7920 & ~n38452;
  assign n38576 = ~n24264 & ~n37855;
  assign n38577 = ~n8214 & ~n38576;
  assign n38578 = n8214 & ~n37856;
  assign n38579 = ~n38577 & ~n38578;
  assign n38580 = n8202 & ~n38579;
  assign n38581 = ~n24261 & ~n38580;
  assign n38582 = n7920 & ~n38581;
  assign n38583 = ~n38575 & ~n38582;
  assign n38584 = ~n7728 & ~n38583;
  assign n38585 = ~n38574 & ~n38584;
  assign n38586 = ~n7723 & ~n38585;
  assign n38587 = ~n7723 & ~n38586;
  assign n38588 = ~n7714 & ~n38587;
  assign n38589 = ~n7714 & ~n38588;
  assign n38590 = n7705 & ~n38589;
  assign n38591 = ~n24287 & ~n35563;
  assign n38592 = i_hbusreq7 & ~n38591;
  assign n38593 = ~n24303 & ~n35574;
  assign n38594 = ~i_hbusreq7 & ~n38593;
  assign n38595 = ~n38592 & ~n38594;
  assign n38596 = ~n7924 & ~n38595;
  assign n38597 = ~n24327 & ~n35584;
  assign n38598 = i_hbusreq7 & ~n38597;
  assign n38599 = ~n24370 & ~n35595;
  assign n38600 = ~i_hbusreq7 & ~n38599;
  assign n38601 = ~n38598 & ~n38600;
  assign n38602 = n7924 & ~n38601;
  assign n38603 = ~n38596 & ~n38602;
  assign n38604 = ~n8214 & ~n38603;
  assign n38605 = ~n24384 & ~n35563;
  assign n38606 = i_hbusreq7 & ~n38605;
  assign n38607 = ~n24400 & ~n36176;
  assign n38608 = ~i_hbusreq7 & ~n38607;
  assign n38609 = ~n38606 & ~n38608;
  assign n38610 = ~n7924 & ~n38609;
  assign n38611 = ~n24422 & ~n35584;
  assign n38612 = i_hbusreq7 & ~n38611;
  assign n38613 = ~n24474 & ~n36188;
  assign n38614 = ~i_hbusreq7 & ~n38613;
  assign n38615 = ~n38612 & ~n38614;
  assign n38616 = n7924 & ~n38615;
  assign n38617 = ~n38610 & ~n38616;
  assign n38618 = n8214 & ~n38617;
  assign n38619 = ~n38604 & ~n38618;
  assign n38620 = ~n8202 & ~n38619;
  assign n38621 = n8202 & ~n37856;
  assign n38622 = ~n38620 & ~n38621;
  assign n38623 = n7920 & ~n38622;
  assign n38624 = ~n38575 & ~n38623;
  assign n38625 = n7728 & ~n38624;
  assign n38626 = ~n24495 & ~n37317;
  assign n38627 = i_hlock7 & ~n38626;
  assign n38628 = ~n24503 & ~n37317;
  assign n38629 = ~i_hlock7 & ~n38628;
  assign n38630 = ~n38627 & ~n38629;
  assign n38631 = i_hbusreq7 & ~n38630;
  assign n38632 = ~n24521 & ~n37332;
  assign n38633 = i_hlock7 & ~n38632;
  assign n38634 = ~n24535 & ~n37332;
  assign n38635 = ~i_hlock7 & ~n38634;
  assign n38636 = ~n38633 & ~n38635;
  assign n38637 = ~i_hbusreq7 & ~n38636;
  assign n38638 = ~n38631 & ~n38637;
  assign n38639 = ~n7924 & ~n38638;
  assign n38640 = ~n24561 & ~n37346;
  assign n38641 = i_hlock7 & ~n38640;
  assign n38642 = ~n24569 & ~n37346;
  assign n38643 = ~i_hlock7 & ~n38642;
  assign n38644 = ~n38641 & ~n38643;
  assign n38645 = i_hbusreq7 & ~n38644;
  assign n38646 = ~n24614 & ~n37361;
  assign n38647 = i_hlock7 & ~n38646;
  assign n38648 = ~n24628 & ~n37361;
  assign n38649 = ~i_hlock7 & ~n38648;
  assign n38650 = ~n38647 & ~n38649;
  assign n38651 = ~i_hbusreq7 & ~n38650;
  assign n38652 = ~n38645 & ~n38651;
  assign n38653 = n7924 & ~n38652;
  assign n38654 = ~n38639 & ~n38653;
  assign n38655 = ~n8214 & ~n38654;
  assign n38656 = ~n24648 & ~n37317;
  assign n38657 = i_hlock7 & ~n38656;
  assign n38658 = ~n24652 & ~n37317;
  assign n38659 = ~i_hlock7 & ~n38658;
  assign n38660 = ~n38657 & ~n38659;
  assign n38661 = i_hbusreq7 & ~n38660;
  assign n38662 = ~controllable_hmaster2 & ~n33999;
  assign n38663 = ~n24687 & ~n38662;
  assign n38664 = ~controllable_hmaster1 & ~n38663;
  assign n38665 = ~n24686 & ~n38664;
  assign n38666 = ~i_hbusreq6 & ~n38665;
  assign n38667 = ~n37027 & ~n38666;
  assign n38668 = ~controllable_hgrant6 & ~n38667;
  assign n38669 = ~n14927 & ~n38668;
  assign n38670 = ~controllable_hmaster0 & ~n38669;
  assign n38671 = ~n33980 & ~n38670;
  assign n38672 = i_hlock8 & ~n38671;
  assign n38673 = ~controllable_hmaster2 & ~n34025;
  assign n38674 = ~n24687 & ~n38673;
  assign n38675 = ~controllable_hmaster1 & ~n38674;
  assign n38676 = ~n24686 & ~n38675;
  assign n38677 = ~i_hbusreq6 & ~n38676;
  assign n38678 = ~n37039 & ~n38677;
  assign n38679 = ~controllable_hgrant6 & ~n38678;
  assign n38680 = ~n14960 & ~n38679;
  assign n38681 = ~controllable_hmaster0 & ~n38680;
  assign n38682 = ~n33980 & ~n38681;
  assign n38683 = ~i_hlock8 & ~n38682;
  assign n38684 = ~n38672 & ~n38683;
  assign n38685 = ~i_hbusreq8 & ~n38684;
  assign n38686 = ~n37324 & ~n38685;
  assign n38687 = controllable_hmaster3 & ~n38686;
  assign n38688 = ~n24919 & ~n38687;
  assign n38689 = i_hlock7 & ~n38688;
  assign n38690 = ~n24934 & ~n38687;
  assign n38691 = ~i_hlock7 & ~n38690;
  assign n38692 = ~n38689 & ~n38691;
  assign n38693 = ~i_hbusreq7 & ~n38692;
  assign n38694 = ~n38661 & ~n38693;
  assign n38695 = ~n7924 & ~n38694;
  assign n38696 = ~n24962 & ~n37346;
  assign n38697 = i_hlock7 & ~n38696;
  assign n38698 = ~n24966 & ~n37346;
  assign n38699 = ~i_hlock7 & ~n38698;
  assign n38700 = ~n38697 & ~n38699;
  assign n38701 = i_hbusreq7 & ~n38700;
  assign n38702 = ~controllable_hmaster2 & ~n34095;
  assign n38703 = ~n25015 & ~n38702;
  assign n38704 = ~controllable_hmaster1 & ~n38703;
  assign n38705 = ~n25014 & ~n38704;
  assign n38706 = ~i_hbusreq6 & ~n38705;
  assign n38707 = ~n37090 & ~n38706;
  assign n38708 = ~controllable_hgrant6 & ~n38707;
  assign n38709 = ~n14927 & ~n38708;
  assign n38710 = ~controllable_hmaster0 & ~n38709;
  assign n38711 = ~n34076 & ~n38710;
  assign n38712 = i_hlock8 & ~n38711;
  assign n38713 = ~controllable_hmaster2 & ~n34121;
  assign n38714 = ~n25015 & ~n38713;
  assign n38715 = ~controllable_hmaster1 & ~n38714;
  assign n38716 = ~n25014 & ~n38715;
  assign n38717 = ~i_hbusreq6 & ~n38716;
  assign n38718 = ~n37102 & ~n38717;
  assign n38719 = ~controllable_hgrant6 & ~n38718;
  assign n38720 = ~n14960 & ~n38719;
  assign n38721 = ~controllable_hmaster0 & ~n38720;
  assign n38722 = ~n34076 & ~n38721;
  assign n38723 = ~i_hlock8 & ~n38722;
  assign n38724 = ~n38712 & ~n38723;
  assign n38725 = ~i_hbusreq8 & ~n38724;
  assign n38726 = ~n37353 & ~n38725;
  assign n38727 = controllable_hmaster3 & ~n38726;
  assign n38728 = ~n25274 & ~n38727;
  assign n38729 = i_hlock7 & ~n38728;
  assign n38730 = ~n25289 & ~n38727;
  assign n38731 = ~i_hlock7 & ~n38730;
  assign n38732 = ~n38729 & ~n38731;
  assign n38733 = ~i_hbusreq7 & ~n38732;
  assign n38734 = ~n38701 & ~n38733;
  assign n38735 = n7924 & ~n38734;
  assign n38736 = ~n38695 & ~n38735;
  assign n38737 = n8214 & ~n38736;
  assign n38738 = ~n38655 & ~n38737;
  assign n38739 = ~n8202 & ~n38738;
  assign n38740 = ~n38621 & ~n38739;
  assign n38741 = n7920 & ~n38740;
  assign n38742 = ~n38575 & ~n38741;
  assign n38743 = ~n7728 & ~n38742;
  assign n38744 = ~n38625 & ~n38743;
  assign n38745 = n7723 & ~n38744;
  assign n38746 = ~n7723 & ~n38742;
  assign n38747 = ~n38745 & ~n38746;
  assign n38748 = n7714 & ~n38747;
  assign n38749 = n7723 & ~n38742;
  assign n38750 = ~n34156 & ~n37435;
  assign n38751 = ~controllable_hgrant6 & ~n38750;
  assign n38752 = ~n13849 & ~n38751;
  assign n38753 = controllable_hmaster0 & ~n38752;
  assign n38754 = ~n31074 & ~n38753;
  assign n38755 = i_hlock8 & ~n38754;
  assign n38756 = ~n34166 & ~n37443;
  assign n38757 = ~controllable_hgrant6 & ~n38756;
  assign n38758 = ~n13849 & ~n38757;
  assign n38759 = controllable_hmaster0 & ~n38758;
  assign n38760 = ~n31181 & ~n38759;
  assign n38761 = ~i_hlock8 & ~n38760;
  assign n38762 = ~n38755 & ~n38761;
  assign n38763 = ~controllable_hmaster3 & ~n38762;
  assign n38764 = ~n37576 & ~n38763;
  assign n38765 = i_hlock7 & ~n38764;
  assign n38766 = ~n34156 & ~n37455;
  assign n38767 = ~controllable_hgrant6 & ~n38766;
  assign n38768 = ~n13951 & ~n38767;
  assign n38769 = controllable_hmaster0 & ~n38768;
  assign n38770 = ~n31074 & ~n38769;
  assign n38771 = i_hlock8 & ~n38770;
  assign n38772 = ~n34166 & ~n37463;
  assign n38773 = ~controllable_hgrant6 & ~n38772;
  assign n38774 = ~n13951 & ~n38773;
  assign n38775 = controllable_hmaster0 & ~n38774;
  assign n38776 = ~n31181 & ~n38775;
  assign n38777 = ~i_hlock8 & ~n38776;
  assign n38778 = ~n38771 & ~n38777;
  assign n38779 = ~controllable_hmaster3 & ~n38778;
  assign n38780 = ~n37576 & ~n38779;
  assign n38781 = ~i_hlock7 & ~n38780;
  assign n38782 = ~n38765 & ~n38781;
  assign n38783 = i_hbusreq7 & ~n38782;
  assign n38784 = i_hbusreq8 & ~n38762;
  assign n38785 = i_hbusreq6 & ~n38750;
  assign n38786 = ~n34191 & ~n37508;
  assign n38787 = ~i_hbusreq6 & ~n38786;
  assign n38788 = ~n38785 & ~n38787;
  assign n38789 = ~controllable_hgrant6 & ~n38788;
  assign n38790 = ~n16031 & ~n38789;
  assign n38791 = controllable_hmaster0 & ~n38790;
  assign n38792 = ~n31403 & ~n38791;
  assign n38793 = i_hlock8 & ~n38792;
  assign n38794 = i_hbusreq6 & ~n38756;
  assign n38795 = ~n34218 & ~n37519;
  assign n38796 = ~i_hbusreq6 & ~n38795;
  assign n38797 = ~n38794 & ~n38796;
  assign n38798 = ~controllable_hgrant6 & ~n38797;
  assign n38799 = ~n16031 & ~n38798;
  assign n38800 = controllable_hmaster0 & ~n38799;
  assign n38801 = ~n31625 & ~n38800;
  assign n38802 = ~i_hlock8 & ~n38801;
  assign n38803 = ~n38793 & ~n38802;
  assign n38804 = ~i_hbusreq8 & ~n38803;
  assign n38805 = ~n38784 & ~n38804;
  assign n38806 = ~controllable_hmaster3 & ~n38805;
  assign n38807 = ~n37627 & ~n38806;
  assign n38808 = i_hlock7 & ~n38807;
  assign n38809 = i_hbusreq8 & ~n38778;
  assign n38810 = i_hbusreq6 & ~n38766;
  assign n38811 = ~n34191 & ~n37537;
  assign n38812 = ~i_hbusreq6 & ~n38811;
  assign n38813 = ~n38810 & ~n38812;
  assign n38814 = ~controllable_hgrant6 & ~n38813;
  assign n38815 = ~n16068 & ~n38814;
  assign n38816 = controllable_hmaster0 & ~n38815;
  assign n38817 = ~n31403 & ~n38816;
  assign n38818 = i_hlock8 & ~n38817;
  assign n38819 = i_hbusreq6 & ~n38772;
  assign n38820 = ~n34218 & ~n37548;
  assign n38821 = ~i_hbusreq6 & ~n38820;
  assign n38822 = ~n38819 & ~n38821;
  assign n38823 = ~controllable_hgrant6 & ~n38822;
  assign n38824 = ~n16068 & ~n38823;
  assign n38825 = controllable_hmaster0 & ~n38824;
  assign n38826 = ~n31625 & ~n38825;
  assign n38827 = ~i_hlock8 & ~n38826;
  assign n38828 = ~n38818 & ~n38827;
  assign n38829 = ~i_hbusreq8 & ~n38828;
  assign n38830 = ~n38809 & ~n38829;
  assign n38831 = ~controllable_hmaster3 & ~n38830;
  assign n38832 = ~n37627 & ~n38831;
  assign n38833 = ~i_hlock7 & ~n38832;
  assign n38834 = ~n38808 & ~n38833;
  assign n38835 = ~i_hbusreq7 & ~n38834;
  assign n38836 = ~n38783 & ~n38835;
  assign n38837 = n7924 & ~n38836;
  assign n38838 = ~n38639 & ~n38837;
  assign n38839 = ~n8214 & ~n38838;
  assign n38840 = ~n34246 & ~n37439;
  assign n38841 = i_hlock8 & ~n38840;
  assign n38842 = ~n34260 & ~n37447;
  assign n38843 = ~i_hlock8 & ~n38842;
  assign n38844 = ~n38841 & ~n38843;
  assign n38845 = ~controllable_hmaster3 & ~n38844;
  assign n38846 = ~n37576 & ~n38845;
  assign n38847 = i_hlock7 & ~n38846;
  assign n38848 = ~n34246 & ~n37459;
  assign n38849 = i_hlock8 & ~n38848;
  assign n38850 = ~n34260 & ~n37467;
  assign n38851 = ~i_hlock8 & ~n38850;
  assign n38852 = ~n38849 & ~n38851;
  assign n38853 = ~controllable_hmaster3 & ~n38852;
  assign n38854 = ~n37576 & ~n38853;
  assign n38855 = ~i_hlock7 & ~n38854;
  assign n38856 = ~n38847 & ~n38855;
  assign n38857 = i_hbusreq7 & ~n38856;
  assign n38858 = ~controllable_hmaster2 & ~n34356;
  assign n38859 = ~n34278 & ~n38858;
  assign n38860 = ~controllable_hmaster1 & ~n38859;
  assign n38861 = ~n34277 & ~n38860;
  assign n38862 = ~i_hbusreq6 & ~n38861;
  assign n38863 = ~n37477 & ~n38862;
  assign n38864 = ~controllable_hgrant6 & ~n38863;
  assign n38865 = ~n14927 & ~n38864;
  assign n38866 = ~controllable_hmaster0 & ~n38865;
  assign n38867 = ~n34299 & ~n38866;
  assign n38868 = i_hlock8 & ~n38867;
  assign n38869 = ~controllable_hmaster2 & ~n34535;
  assign n38870 = ~n34457 & ~n38869;
  assign n38871 = ~controllable_hmaster1 & ~n38870;
  assign n38872 = ~n34456 & ~n38871;
  assign n38873 = ~i_hbusreq6 & ~n38872;
  assign n38874 = ~n37489 & ~n38873;
  assign n38875 = ~controllable_hgrant6 & ~n38874;
  assign n38876 = ~n14960 & ~n38875;
  assign n38877 = ~controllable_hmaster0 & ~n38876;
  assign n38878 = ~n34478 & ~n38877;
  assign n38879 = ~i_hlock8 & ~n38878;
  assign n38880 = ~n38868 & ~n38879;
  assign n38881 = ~i_hbusreq8 & ~n38880;
  assign n38882 = ~n37619 & ~n38881;
  assign n38883 = controllable_hmaster3 & ~n38882;
  assign n38884 = i_hbusreq8 & ~n38844;
  assign n38885 = ~n34368 & ~n34399;
  assign n38886 = controllable_hmaster1 & ~n38885;
  assign n38887 = ~n34391 & ~n38886;
  assign n38888 = ~i_hbusreq6 & ~n38887;
  assign n38889 = ~n37506 & ~n38888;
  assign n38890 = ~controllable_hgrant6 & ~n38889;
  assign n38891 = ~n14995 & ~n38890;
  assign n38892 = controllable_hmaster0 & ~n38891;
  assign n38893 = ~n34439 & ~n38892;
  assign n38894 = i_hlock8 & ~n38893;
  assign n38895 = ~n34547 & ~n34578;
  assign n38896 = controllable_hmaster1 & ~n38895;
  assign n38897 = ~n34570 & ~n38896;
  assign n38898 = ~i_hbusreq6 & ~n38897;
  assign n38899 = ~n37517 & ~n38898;
  assign n38900 = ~controllable_hgrant6 & ~n38899;
  assign n38901 = ~n14995 & ~n38900;
  assign n38902 = controllable_hmaster0 & ~n38901;
  assign n38903 = ~n34618 & ~n38902;
  assign n38904 = ~i_hlock8 & ~n38903;
  assign n38905 = ~n38894 & ~n38904;
  assign n38906 = ~i_hbusreq8 & ~n38905;
  assign n38907 = ~n38884 & ~n38906;
  assign n38908 = ~controllable_hmaster3 & ~n38907;
  assign n38909 = ~n38883 & ~n38908;
  assign n38910 = i_hlock7 & ~n38909;
  assign n38911 = i_hbusreq8 & ~n38852;
  assign n38912 = ~n34368 & ~n34429;
  assign n38913 = controllable_hmaster1 & ~n38912;
  assign n38914 = ~n34391 & ~n38913;
  assign n38915 = ~i_hbusreq6 & ~n38914;
  assign n38916 = ~n37535 & ~n38915;
  assign n38917 = ~controllable_hgrant6 & ~n38916;
  assign n38918 = ~n15152 & ~n38917;
  assign n38919 = controllable_hmaster0 & ~n38918;
  assign n38920 = ~n34439 & ~n38919;
  assign n38921 = i_hlock8 & ~n38920;
  assign n38922 = ~n34547 & ~n34608;
  assign n38923 = controllable_hmaster1 & ~n38922;
  assign n38924 = ~n34570 & ~n38923;
  assign n38925 = ~i_hbusreq6 & ~n38924;
  assign n38926 = ~n37546 & ~n38925;
  assign n38927 = ~controllable_hgrant6 & ~n38926;
  assign n38928 = ~n15152 & ~n38927;
  assign n38929 = controllable_hmaster0 & ~n38928;
  assign n38930 = ~n34618 & ~n38929;
  assign n38931 = ~i_hlock8 & ~n38930;
  assign n38932 = ~n38921 & ~n38931;
  assign n38933 = ~i_hbusreq8 & ~n38932;
  assign n38934 = ~n38911 & ~n38933;
  assign n38935 = ~controllable_hmaster3 & ~n38934;
  assign n38936 = ~n38883 & ~n38935;
  assign n38937 = ~i_hlock7 & ~n38936;
  assign n38938 = ~n38910 & ~n38937;
  assign n38939 = ~i_hbusreq7 & ~n38938;
  assign n38940 = ~n38857 & ~n38939;
  assign n38941 = n7924 & ~n38940;
  assign n38942 = ~n38695 & ~n38941;
  assign n38943 = n8214 & ~n38942;
  assign n38944 = ~n38839 & ~n38943;
  assign n38945 = ~n8202 & ~n38944;
  assign n38946 = ~n38621 & ~n38945;
  assign n38947 = n7920 & ~n38946;
  assign n38948 = ~n36523 & ~n38947;
  assign n38949 = n7728 & ~n38948;
  assign n38950 = ~n37859 & ~n38949;
  assign n38951 = ~n7723 & ~n38950;
  assign n38952 = ~n38749 & ~n38951;
  assign n38953 = ~n7714 & ~n38952;
  assign n38954 = ~n38748 & ~n38953;
  assign n38955 = ~n7705 & ~n38954;
  assign n38956 = ~n38590 & ~n38955;
  assign n38957 = n7808 & ~n38956;
  assign n38958 = ~n38469 & ~n38957;
  assign n38959 = n8195 & ~n38958;
  assign n38960 = ~n38383 & ~n38959;
  assign n38961 = n8193 & ~n38960;
  assign n38962 = ~n37871 & ~n38961;
  assign n38963 = n8191 & ~n38962;
  assign n38964 = ~n10987 & ~n36394;
  assign n38965 = ~n8202 & ~n38964;
  assign n38966 = ~n8332 & ~n38965;
  assign n38967 = n7728 & ~n38966;
  assign n38968 = ~n11017 & ~n36455;
  assign n38969 = ~n8202 & ~n38968;
  assign n38970 = ~n8347 & ~n38969;
  assign n38971 = ~n7728 & ~n38970;
  assign n38972 = ~n38967 & ~n38971;
  assign n38973 = ~n7723 & ~n38972;
  assign n38974 = ~n7723 & ~n38973;
  assign n38975 = ~n7714 & ~n38974;
  assign n38976 = ~n7714 & ~n38975;
  assign n38977 = n7705 & ~n38976;
  assign n38978 = n7723 & ~n38970;
  assign n38979 = ~n11033 & ~n36473;
  assign n38980 = i_hlock8 & ~n38979;
  assign n38981 = ~n11033 & ~n36482;
  assign n38982 = ~i_hlock8 & ~n38981;
  assign n38983 = ~n38980 & ~n38982;
  assign n38984 = controllable_hmaster3 & ~n38983;
  assign n38985 = ~n8463 & ~n38984;
  assign n38986 = i_hbusreq7 & ~n38985;
  assign n38987 = i_hbusreq8 & ~n38983;
  assign n38988 = ~n11046 & ~n36499;
  assign n38989 = i_hlock8 & ~n38988;
  assign n38990 = ~n11046 & ~n36511;
  assign n38991 = ~i_hlock8 & ~n38990;
  assign n38992 = ~n38989 & ~n38991;
  assign n38993 = ~i_hbusreq8 & ~n38992;
  assign n38994 = ~n38987 & ~n38993;
  assign n38995 = controllable_hmaster3 & ~n38994;
  assign n38996 = ~n8634 & ~n38995;
  assign n38997 = ~i_hbusreq7 & ~n38996;
  assign n38998 = ~n38986 & ~n38997;
  assign n38999 = n7924 & ~n38998;
  assign n39000 = ~n8337 & ~n38999;
  assign n39001 = ~n7920 & ~n39000;
  assign n39002 = n7920 & ~n38970;
  assign n39003 = ~n39001 & ~n39002;
  assign n39004 = ~n7723 & ~n39003;
  assign n39005 = ~n38978 & ~n39004;
  assign n39006 = n7714 & ~n39005;
  assign n39007 = ~n7714 & ~n39000;
  assign n39008 = ~n39006 & ~n39007;
  assign n39009 = ~n7705 & ~n39008;
  assign n39010 = ~n38977 & ~n39009;
  assign n39011 = ~n7808 & ~n39010;
  assign n39012 = ~n7920 & ~n38966;
  assign n39013 = ~n36673 & ~n39012;
  assign n39014 = n7728 & ~n39013;
  assign n39015 = ~n7920 & ~n38970;
  assign n39016 = ~n36790 & ~n39015;
  assign n39017 = ~n7728 & ~n39016;
  assign n39018 = ~n39014 & ~n39017;
  assign n39019 = ~n7723 & ~n39018;
  assign n39020 = ~n7723 & ~n39019;
  assign n39021 = ~n7714 & ~n39020;
  assign n39022 = ~n7714 & ~n39021;
  assign n39023 = n7705 & ~n39022;
  assign n39024 = ~n36997 & ~n39015;
  assign n39025 = n7728 & ~n39024;
  assign n39026 = ~n37405 & ~n39015;
  assign n39027 = ~n7728 & ~n39026;
  assign n39028 = ~n39025 & ~n39027;
  assign n39029 = n7723 & ~n39028;
  assign n39030 = ~n7723 & ~n39026;
  assign n39031 = ~n39029 & ~n39030;
  assign n39032 = n7714 & ~n39031;
  assign n39033 = n7723 & ~n39026;
  assign n39034 = ~n37741 & ~n39001;
  assign n39035 = n7728 & ~n39034;
  assign n39036 = ~n37857 & ~n39001;
  assign n39037 = ~n7728 & ~n39036;
  assign n39038 = ~n39035 & ~n39037;
  assign n39039 = ~n7723 & ~n39038;
  assign n39040 = ~n39033 & ~n39039;
  assign n39041 = ~n7714 & ~n39040;
  assign n39042 = ~n39032 & ~n39041;
  assign n39043 = ~n7705 & ~n39042;
  assign n39044 = ~n39023 & ~n39043;
  assign n39045 = n7808 & ~n39044;
  assign n39046 = ~n39011 & ~n39045;
  assign n39047 = n8195 & ~n39046;
  assign n39048 = ~n8196 & ~n39047;
  assign n39049 = ~n8193 & ~n39048;
  assign n39050 = ~n9900 & ~n39001;
  assign n39051 = ~n7723 & ~n39050;
  assign n39052 = ~n9899 & ~n39051;
  assign n39053 = n7714 & ~n39052;
  assign n39054 = ~n39007 & ~n39053;
  assign n39055 = ~n7705 & ~n39054;
  assign n39056 = ~n9898 & ~n39055;
  assign n39057 = ~n7808 & ~n39056;
  assign n39058 = ~n38371 & ~n39001;
  assign n39059 = n7728 & ~n39058;
  assign n39060 = ~n39037 & ~n39059;
  assign n39061 = ~n7723 & ~n39060;
  assign n39062 = ~n38077 & ~n39061;
  assign n39063 = ~n7714 & ~n39062;
  assign n39064 = ~n38076 & ~n39063;
  assign n39065 = ~n7705 & ~n39064;
  assign n39066 = ~n22399 & ~n39065;
  assign n39067 = n7808 & ~n39066;
  assign n39068 = ~n39057 & ~n39067;
  assign n39069 = ~n8195 & ~n39068;
  assign n39070 = ~n11133 & ~n38391;
  assign n39071 = i_hlock8 & ~n39070;
  assign n39072 = ~n11133 & ~n38401;
  assign n39073 = ~i_hlock8 & ~n39072;
  assign n39074 = ~n39071 & ~n39073;
  assign n39075 = controllable_hmaster3 & ~n39074;
  assign n39076 = ~n10447 & ~n39075;
  assign n39077 = i_hbusreq7 & ~n39076;
  assign n39078 = i_hbusreq8 & ~n39074;
  assign n39079 = ~n11159 & ~n38419;
  assign n39080 = i_hlock8 & ~n39079;
  assign n39081 = ~n11159 & ~n38432;
  assign n39082 = ~i_hlock8 & ~n39081;
  assign n39083 = ~n39080 & ~n39082;
  assign n39084 = ~i_hbusreq8 & ~n39083;
  assign n39085 = ~n39078 & ~n39084;
  assign n39086 = controllable_hmaster3 & ~n39085;
  assign n39087 = ~n10621 & ~n39086;
  assign n39088 = ~i_hbusreq7 & ~n39087;
  assign n39089 = ~n39077 & ~n39088;
  assign n39090 = n7924 & ~n39089;
  assign n39091 = ~n10375 & ~n39090;
  assign n39092 = n8214 & ~n39091;
  assign n39093 = n8214 & ~n39092;
  assign n39094 = n8202 & ~n39093;
  assign n39095 = ~n10332 & ~n39094;
  assign n39096 = n7728 & ~n39095;
  assign n39097 = n8214 & ~n39000;
  assign n39098 = ~n8336 & ~n39097;
  assign n39099 = n8202 & ~n39098;
  assign n39100 = ~n10649 & ~n39099;
  assign n39101 = ~n7728 & ~n39100;
  assign n39102 = ~n39096 & ~n39101;
  assign n39103 = ~n7723 & ~n39102;
  assign n39104 = ~n7723 & ~n39103;
  assign n39105 = ~n7714 & ~n39104;
  assign n39106 = ~n7714 & ~n39105;
  assign n39107 = n7705 & ~n39106;
  assign n39108 = n7723 & ~n39100;
  assign n39109 = n7920 & ~n39100;
  assign n39110 = ~n39001 & ~n39109;
  assign n39111 = ~n7723 & ~n39110;
  assign n39112 = ~n39108 & ~n39111;
  assign n39113 = n7714 & ~n39112;
  assign n39114 = ~n39007 & ~n39113;
  assign n39115 = ~n7705 & ~n39114;
  assign n39116 = ~n39107 & ~n39115;
  assign n39117 = ~n7808 & ~n39116;
  assign n39118 = ~n7920 & ~n39095;
  assign n39119 = ~n38572 & ~n39118;
  assign n39120 = n7728 & ~n39119;
  assign n39121 = ~n7920 & ~n39100;
  assign n39122 = ~n38582 & ~n39121;
  assign n39123 = ~n7728 & ~n39122;
  assign n39124 = ~n39120 & ~n39123;
  assign n39125 = ~n7723 & ~n39124;
  assign n39126 = ~n7723 & ~n39125;
  assign n39127 = ~n7714 & ~n39126;
  assign n39128 = ~n7714 & ~n39127;
  assign n39129 = n7705 & ~n39128;
  assign n39130 = ~n38623 & ~n39121;
  assign n39131 = n7728 & ~n39130;
  assign n39132 = ~n38741 & ~n39121;
  assign n39133 = ~n7728 & ~n39132;
  assign n39134 = ~n39131 & ~n39133;
  assign n39135 = n7723 & ~n39134;
  assign n39136 = ~n7723 & ~n39132;
  assign n39137 = ~n39135 & ~n39136;
  assign n39138 = n7714 & ~n39137;
  assign n39139 = n7723 & ~n39132;
  assign n39140 = ~n38947 & ~n39001;
  assign n39141 = n7728 & ~n39140;
  assign n39142 = ~n39037 & ~n39141;
  assign n39143 = ~n7723 & ~n39142;
  assign n39144 = ~n39139 & ~n39143;
  assign n39145 = ~n7714 & ~n39144;
  assign n39146 = ~n39138 & ~n39145;
  assign n39147 = ~n7705 & ~n39146;
  assign n39148 = ~n39129 & ~n39147;
  assign n39149 = n7808 & ~n39148;
  assign n39150 = ~n39117 & ~n39149;
  assign n39151 = n8195 & ~n39150;
  assign n39152 = ~n39069 & ~n39151;
  assign n39153 = n8193 & ~n39152;
  assign n39154 = ~n39049 & ~n39153;
  assign n39155 = ~n8191 & ~n39154;
  assign n39156 = ~n38963 & ~n39155;
  assign n39157 = ~n8188 & ~n39156;
  assign n39158 = ~n36333 & ~n39157;
  assign n39159 = n8185 & ~n39158;
  assign n39160 = ~n11903 & ~n35302;
  assign n39161 = n7728 & ~n39160;
  assign n39162 = ~n11906 & ~n35414;
  assign n39163 = ~n7728 & ~n39162;
  assign n39164 = ~n39161 & ~n39163;
  assign n39165 = ~n7723 & ~n39164;
  assign n39166 = ~n7723 & ~n39165;
  assign n39167 = ~n7714 & ~n39166;
  assign n39168 = ~n7714 & ~n39167;
  assign n39169 = n7705 & ~n39168;
  assign n39170 = ~n11906 & ~n35623;
  assign n39171 = n7728 & ~n39170;
  assign n39172 = ~n11906 & ~n35845;
  assign n39173 = ~n7728 & ~n39172;
  assign n39174 = ~n39171 & ~n39173;
  assign n39175 = n7723 & ~n39174;
  assign n39176 = ~n7723 & ~n39172;
  assign n39177 = ~n39175 & ~n39176;
  assign n39178 = n7714 & ~n39177;
  assign n39179 = n7723 & ~n39172;
  assign n39180 = ~n11892 & ~n35845;
  assign n39181 = n7728 & ~n39180;
  assign n39182 = ~n11892 & ~n35921;
  assign n39183 = ~n7728 & ~n39182;
  assign n39184 = ~n39181 & ~n39183;
  assign n39185 = ~n7723 & ~n39184;
  assign n39186 = ~n39179 & ~n39185;
  assign n39187 = ~n7714 & ~n39186;
  assign n39188 = ~n39178 & ~n39187;
  assign n39189 = ~n7705 & ~n39188;
  assign n39190 = ~n39169 & ~n39189;
  assign n39191 = n7808 & ~n39190;
  assign n39192 = ~n11902 & ~n39191;
  assign n39193 = n8195 & ~n39192;
  assign n39194 = ~n8196 & ~n39193;
  assign n39195 = ~n8193 & ~n39194;
  assign n39196 = ~n11892 & ~n36077;
  assign n39197 = n7728 & ~n39196;
  assign n39198 = ~n39183 & ~n39197;
  assign n39199 = ~n7723 & ~n39198;
  assign n39200 = ~n36085 & ~n39199;
  assign n39201 = ~n7714 & ~n39200;
  assign n39202 = ~n36084 & ~n39201;
  assign n39203 = ~n7705 & ~n39202;
  assign n39204 = ~n10052 & ~n39203;
  assign n39205 = n7808 & ~n39204;
  assign n39206 = ~n11948 & ~n39205;
  assign n39207 = ~n8195 & ~n39206;
  assign n39208 = ~n12038 & ~n36137;
  assign n39209 = n7728 & ~n39208;
  assign n39210 = ~n12041 & ~n36146;
  assign n39211 = ~n7728 & ~n39210;
  assign n39212 = ~n39209 & ~n39211;
  assign n39213 = ~n7723 & ~n39212;
  assign n39214 = ~n7723 & ~n39213;
  assign n39215 = ~n7714 & ~n39214;
  assign n39216 = ~n7714 & ~n39215;
  assign n39217 = n7705 & ~n39216;
  assign n39218 = ~n12041 & ~n36199;
  assign n39219 = n7728 & ~n39218;
  assign n39220 = ~n12041 & ~n36223;
  assign n39221 = ~n7728 & ~n39220;
  assign n39222 = ~n39219 & ~n39221;
  assign n39223 = n7723 & ~n39222;
  assign n39224 = ~n7723 & ~n39220;
  assign n39225 = ~n39223 & ~n39224;
  assign n39226 = n7714 & ~n39225;
  assign n39227 = n7723 & ~n39220;
  assign n39228 = ~n11892 & ~n36223;
  assign n39229 = n7728 & ~n39228;
  assign n39230 = ~n39183 & ~n39229;
  assign n39231 = ~n7723 & ~n39230;
  assign n39232 = ~n39227 & ~n39231;
  assign n39233 = ~n7714 & ~n39232;
  assign n39234 = ~n39226 & ~n39233;
  assign n39235 = ~n7705 & ~n39234;
  assign n39236 = ~n39217 & ~n39235;
  assign n39237 = n7808 & ~n39236;
  assign n39238 = ~n12037 & ~n39237;
  assign n39239 = n8195 & ~n39238;
  assign n39240 = ~n39207 & ~n39239;
  assign n39241 = n8193 & ~n39240;
  assign n39242 = ~n39195 & ~n39241;
  assign n39243 = n8191 & ~n39242;
  assign n39244 = ~n12113 & ~n35302;
  assign n39245 = n7728 & ~n39244;
  assign n39246 = ~n12116 & ~n35414;
  assign n39247 = ~n7728 & ~n39246;
  assign n39248 = ~n39245 & ~n39247;
  assign n39249 = ~n7723 & ~n39248;
  assign n39250 = ~n7723 & ~n39249;
  assign n39251 = ~n7714 & ~n39250;
  assign n39252 = ~n7714 & ~n39251;
  assign n39253 = n7705 & ~n39252;
  assign n39254 = ~n12116 & ~n35623;
  assign n39255 = n7728 & ~n39254;
  assign n39256 = ~n12116 & ~n35845;
  assign n39257 = ~n7728 & ~n39256;
  assign n39258 = ~n39255 & ~n39257;
  assign n39259 = n7723 & ~n39258;
  assign n39260 = ~n7723 & ~n39256;
  assign n39261 = ~n39259 & ~n39260;
  assign n39262 = n7714 & ~n39261;
  assign n39263 = n7723 & ~n39256;
  assign n39264 = ~n12102 & ~n35845;
  assign n39265 = n7728 & ~n39264;
  assign n39266 = ~n12102 & ~n35921;
  assign n39267 = ~n7728 & ~n39266;
  assign n39268 = ~n39265 & ~n39267;
  assign n39269 = ~n7723 & ~n39268;
  assign n39270 = ~n39263 & ~n39269;
  assign n39271 = ~n7714 & ~n39270;
  assign n39272 = ~n39262 & ~n39271;
  assign n39273 = ~n7705 & ~n39272;
  assign n39274 = ~n39253 & ~n39273;
  assign n39275 = n7808 & ~n39274;
  assign n39276 = ~n12112 & ~n39275;
  assign n39277 = n8195 & ~n39276;
  assign n39278 = ~n8196 & ~n39277;
  assign n39279 = ~n8193 & ~n39278;
  assign n39280 = ~n12102 & ~n36077;
  assign n39281 = n7728 & ~n39280;
  assign n39282 = ~n39267 & ~n39281;
  assign n39283 = ~n7723 & ~n39282;
  assign n39284 = ~n36085 & ~n39283;
  assign n39285 = ~n7714 & ~n39284;
  assign n39286 = ~n36084 & ~n39285;
  assign n39287 = ~n7705 & ~n39286;
  assign n39288 = ~n10052 & ~n39287;
  assign n39289 = n7808 & ~n39288;
  assign n39290 = ~n12158 & ~n39289;
  assign n39291 = ~n8195 & ~n39290;
  assign n39292 = ~n12212 & ~n36137;
  assign n39293 = n7728 & ~n39292;
  assign n39294 = ~n12215 & ~n36146;
  assign n39295 = ~n7728 & ~n39294;
  assign n39296 = ~n39293 & ~n39295;
  assign n39297 = ~n7723 & ~n39296;
  assign n39298 = ~n7723 & ~n39297;
  assign n39299 = ~n7714 & ~n39298;
  assign n39300 = ~n7714 & ~n39299;
  assign n39301 = n7705 & ~n39300;
  assign n39302 = ~n12215 & ~n36199;
  assign n39303 = n7728 & ~n39302;
  assign n39304 = ~n12215 & ~n36223;
  assign n39305 = ~n7728 & ~n39304;
  assign n39306 = ~n39303 & ~n39305;
  assign n39307 = n7723 & ~n39306;
  assign n39308 = ~n7723 & ~n39304;
  assign n39309 = ~n39307 & ~n39308;
  assign n39310 = n7714 & ~n39309;
  assign n39311 = n7723 & ~n39304;
  assign n39312 = ~n12102 & ~n36223;
  assign n39313 = n7728 & ~n39312;
  assign n39314 = ~n39267 & ~n39313;
  assign n39315 = ~n7723 & ~n39314;
  assign n39316 = ~n39311 & ~n39315;
  assign n39317 = ~n7714 & ~n39316;
  assign n39318 = ~n39310 & ~n39317;
  assign n39319 = ~n7705 & ~n39318;
  assign n39320 = ~n39301 & ~n39319;
  assign n39321 = n7808 & ~n39320;
  assign n39322 = ~n12211 & ~n39321;
  assign n39323 = n8195 & ~n39322;
  assign n39324 = ~n39291 & ~n39323;
  assign n39325 = n8193 & ~n39324;
  assign n39326 = ~n39279 & ~n39325;
  assign n39327 = ~n8191 & ~n39326;
  assign n39328 = ~n39243 & ~n39327;
  assign n39329 = n8188 & ~n39328;
  assign n39330 = ~n11811 & ~n36396;
  assign n39331 = n7728 & ~n39330;
  assign n39332 = ~n11831 & ~n36457;
  assign n39333 = ~n7728 & ~n39332;
  assign n39334 = ~n39331 & ~n39333;
  assign n39335 = ~n7723 & ~n39334;
  assign n39336 = ~n7723 & ~n39335;
  assign n39337 = ~n7714 & ~n39336;
  assign n39338 = ~n7714 & ~n39337;
  assign n39339 = n7705 & ~n39338;
  assign n39340 = n7723 & ~n39332;
  assign n39341 = ~n11846 & ~n36486;
  assign n39342 = i_hlock7 & ~n39341;
  assign n39343 = ~n11854 & ~n36486;
  assign n39344 = ~i_hlock7 & ~n39343;
  assign n39345 = ~n39342 & ~n39344;
  assign n39346 = i_hbusreq7 & ~n39345;
  assign n39347 = ~n11870 & ~n36517;
  assign n39348 = i_hlock7 & ~n39347;
  assign n39349 = ~n11884 & ~n36517;
  assign n39350 = ~i_hlock7 & ~n39349;
  assign n39351 = ~n39348 & ~n39350;
  assign n39352 = ~i_hbusreq7 & ~n39351;
  assign n39353 = ~n39346 & ~n39352;
  assign n39354 = n7924 & ~n39353;
  assign n39355 = ~n8337 & ~n39354;
  assign n39356 = ~n7920 & ~n39355;
  assign n39357 = n7920 & ~n39332;
  assign n39358 = ~n39356 & ~n39357;
  assign n39359 = ~n7723 & ~n39358;
  assign n39360 = ~n39340 & ~n39359;
  assign n39361 = n7714 & ~n39360;
  assign n39362 = ~n7714 & ~n39355;
  assign n39363 = ~n39361 & ~n39362;
  assign n39364 = ~n7705 & ~n39363;
  assign n39365 = ~n39339 & ~n39364;
  assign n39366 = ~n7808 & ~n39365;
  assign n39367 = ~n7920 & ~n39330;
  assign n39368 = ~n36673 & ~n39367;
  assign n39369 = n7728 & ~n39368;
  assign n39370 = ~n7920 & ~n39332;
  assign n39371 = ~n36790 & ~n39370;
  assign n39372 = ~n7728 & ~n39371;
  assign n39373 = ~n39369 & ~n39372;
  assign n39374 = ~n7723 & ~n39373;
  assign n39375 = ~n7723 & ~n39374;
  assign n39376 = ~n7714 & ~n39375;
  assign n39377 = ~n7714 & ~n39376;
  assign n39378 = n7705 & ~n39377;
  assign n39379 = ~n36997 & ~n39370;
  assign n39380 = n7728 & ~n39379;
  assign n39381 = ~n37405 & ~n39370;
  assign n39382 = ~n7728 & ~n39381;
  assign n39383 = ~n39380 & ~n39382;
  assign n39384 = n7723 & ~n39383;
  assign n39385 = ~n7723 & ~n39381;
  assign n39386 = ~n39384 & ~n39385;
  assign n39387 = n7714 & ~n39386;
  assign n39388 = n7723 & ~n39381;
  assign n39389 = ~n37741 & ~n39356;
  assign n39390 = n7728 & ~n39389;
  assign n39391 = ~n37857 & ~n39356;
  assign n39392 = ~n7728 & ~n39391;
  assign n39393 = ~n39390 & ~n39392;
  assign n39394 = ~n7723 & ~n39393;
  assign n39395 = ~n39388 & ~n39394;
  assign n39396 = ~n7714 & ~n39395;
  assign n39397 = ~n39387 & ~n39396;
  assign n39398 = ~n7705 & ~n39397;
  assign n39399 = ~n39378 & ~n39398;
  assign n39400 = n7808 & ~n39399;
  assign n39401 = ~n39366 & ~n39400;
  assign n39402 = n8195 & ~n39401;
  assign n39403 = ~n8196 & ~n39402;
  assign n39404 = ~n8193 & ~n39403;
  assign n39405 = ~n9900 & ~n39356;
  assign n39406 = ~n7723 & ~n39405;
  assign n39407 = ~n9899 & ~n39406;
  assign n39408 = n7714 & ~n39407;
  assign n39409 = ~n39362 & ~n39408;
  assign n39410 = ~n7705 & ~n39409;
  assign n39411 = ~n9898 & ~n39410;
  assign n39412 = ~n7808 & ~n39411;
  assign n39413 = ~n38371 & ~n39356;
  assign n39414 = n7728 & ~n39413;
  assign n39415 = ~n39392 & ~n39414;
  assign n39416 = ~n7723 & ~n39415;
  assign n39417 = ~n38077 & ~n39416;
  assign n39418 = ~n7714 & ~n39417;
  assign n39419 = ~n38076 & ~n39418;
  assign n39420 = ~n7705 & ~n39419;
  assign n39421 = ~n22399 & ~n39420;
  assign n39422 = n7808 & ~n39421;
  assign n39423 = ~n39412 & ~n39422;
  assign n39424 = ~n8195 & ~n39423;
  assign n39425 = ~n11966 & ~n38405;
  assign n39426 = i_hlock7 & ~n39425;
  assign n39427 = ~n11974 & ~n38405;
  assign n39428 = ~i_hlock7 & ~n39427;
  assign n39429 = ~n39426 & ~n39428;
  assign n39430 = i_hbusreq7 & ~n39429;
  assign n39431 = ~n11990 & ~n38438;
  assign n39432 = i_hlock7 & ~n39431;
  assign n39433 = ~n12004 & ~n38438;
  assign n39434 = ~i_hlock7 & ~n39433;
  assign n39435 = ~n39432 & ~n39434;
  assign n39436 = ~i_hbusreq7 & ~n39435;
  assign n39437 = ~n39430 & ~n39436;
  assign n39438 = n7924 & ~n39437;
  assign n39439 = ~n10375 & ~n39438;
  assign n39440 = n8214 & ~n39439;
  assign n39441 = n8214 & ~n39440;
  assign n39442 = n8202 & ~n39441;
  assign n39443 = ~n10332 & ~n39442;
  assign n39444 = n7728 & ~n39443;
  assign n39445 = n8214 & ~n39355;
  assign n39446 = ~n8336 & ~n39445;
  assign n39447 = n8202 & ~n39446;
  assign n39448 = ~n10649 & ~n39447;
  assign n39449 = ~n7728 & ~n39448;
  assign n39450 = ~n39444 & ~n39449;
  assign n39451 = ~n7723 & ~n39450;
  assign n39452 = ~n7723 & ~n39451;
  assign n39453 = ~n7714 & ~n39452;
  assign n39454 = ~n7714 & ~n39453;
  assign n39455 = n7705 & ~n39454;
  assign n39456 = n7723 & ~n39448;
  assign n39457 = n7920 & ~n39448;
  assign n39458 = ~n39356 & ~n39457;
  assign n39459 = ~n7723 & ~n39458;
  assign n39460 = ~n39456 & ~n39459;
  assign n39461 = n7714 & ~n39460;
  assign n39462 = ~n39362 & ~n39461;
  assign n39463 = ~n7705 & ~n39462;
  assign n39464 = ~n39455 & ~n39463;
  assign n39465 = ~n7808 & ~n39464;
  assign n39466 = ~n7920 & ~n39443;
  assign n39467 = ~n38572 & ~n39466;
  assign n39468 = n7728 & ~n39467;
  assign n39469 = ~n7920 & ~n39448;
  assign n39470 = ~n38582 & ~n39469;
  assign n39471 = ~n7728 & ~n39470;
  assign n39472 = ~n39468 & ~n39471;
  assign n39473 = ~n7723 & ~n39472;
  assign n39474 = ~n7723 & ~n39473;
  assign n39475 = ~n7714 & ~n39474;
  assign n39476 = ~n7714 & ~n39475;
  assign n39477 = n7705 & ~n39476;
  assign n39478 = ~n38623 & ~n39469;
  assign n39479 = n7728 & ~n39478;
  assign n39480 = ~n38741 & ~n39469;
  assign n39481 = ~n7728 & ~n39480;
  assign n39482 = ~n39479 & ~n39481;
  assign n39483 = n7723 & ~n39482;
  assign n39484 = ~n7723 & ~n39480;
  assign n39485 = ~n39483 & ~n39484;
  assign n39486 = n7714 & ~n39485;
  assign n39487 = n7723 & ~n39480;
  assign n39488 = ~n38947 & ~n39356;
  assign n39489 = n7728 & ~n39488;
  assign n39490 = ~n39392 & ~n39489;
  assign n39491 = ~n7723 & ~n39490;
  assign n39492 = ~n39487 & ~n39491;
  assign n39493 = ~n7714 & ~n39492;
  assign n39494 = ~n39486 & ~n39493;
  assign n39495 = ~n7705 & ~n39494;
  assign n39496 = ~n39477 & ~n39495;
  assign n39497 = n7808 & ~n39496;
  assign n39498 = ~n39465 & ~n39497;
  assign n39499 = n8195 & ~n39498;
  assign n39500 = ~n39424 & ~n39499;
  assign n39501 = n8193 & ~n39500;
  assign n39502 = ~n39404 & ~n39501;
  assign n39503 = n8191 & ~n39502;
  assign n39504 = ~n11811 & ~n38965;
  assign n39505 = n7728 & ~n39504;
  assign n39506 = ~n11831 & ~n38969;
  assign n39507 = ~n7728 & ~n39506;
  assign n39508 = ~n39505 & ~n39507;
  assign n39509 = ~n7723 & ~n39508;
  assign n39510 = ~n7723 & ~n39509;
  assign n39511 = ~n7714 & ~n39510;
  assign n39512 = ~n7714 & ~n39511;
  assign n39513 = n7705 & ~n39512;
  assign n39514 = n7723 & ~n39506;
  assign n39515 = ~n11846 & ~n38984;
  assign n39516 = i_hlock7 & ~n39515;
  assign n39517 = ~n11854 & ~n38984;
  assign n39518 = ~i_hlock7 & ~n39517;
  assign n39519 = ~n39516 & ~n39518;
  assign n39520 = i_hbusreq7 & ~n39519;
  assign n39521 = ~n11870 & ~n38995;
  assign n39522 = i_hlock7 & ~n39521;
  assign n39523 = ~n11884 & ~n38995;
  assign n39524 = ~i_hlock7 & ~n39523;
  assign n39525 = ~n39522 & ~n39524;
  assign n39526 = ~i_hbusreq7 & ~n39525;
  assign n39527 = ~n39520 & ~n39526;
  assign n39528 = n7924 & ~n39527;
  assign n39529 = ~n8337 & ~n39528;
  assign n39530 = ~n7920 & ~n39529;
  assign n39531 = n7920 & ~n39506;
  assign n39532 = ~n39530 & ~n39531;
  assign n39533 = ~n7723 & ~n39532;
  assign n39534 = ~n39514 & ~n39533;
  assign n39535 = n7714 & ~n39534;
  assign n39536 = ~n7714 & ~n39529;
  assign n39537 = ~n39535 & ~n39536;
  assign n39538 = ~n7705 & ~n39537;
  assign n39539 = ~n39513 & ~n39538;
  assign n39540 = ~n7808 & ~n39539;
  assign n39541 = ~n7920 & ~n39504;
  assign n39542 = ~n36673 & ~n39541;
  assign n39543 = n7728 & ~n39542;
  assign n39544 = ~n7920 & ~n39506;
  assign n39545 = ~n36790 & ~n39544;
  assign n39546 = ~n7728 & ~n39545;
  assign n39547 = ~n39543 & ~n39546;
  assign n39548 = ~n7723 & ~n39547;
  assign n39549 = ~n7723 & ~n39548;
  assign n39550 = ~n7714 & ~n39549;
  assign n39551 = ~n7714 & ~n39550;
  assign n39552 = n7705 & ~n39551;
  assign n39553 = ~n36997 & ~n39544;
  assign n39554 = n7728 & ~n39553;
  assign n39555 = ~n37405 & ~n39544;
  assign n39556 = ~n7728 & ~n39555;
  assign n39557 = ~n39554 & ~n39556;
  assign n39558 = n7723 & ~n39557;
  assign n39559 = ~n7723 & ~n39555;
  assign n39560 = ~n39558 & ~n39559;
  assign n39561 = n7714 & ~n39560;
  assign n39562 = n7723 & ~n39555;
  assign n39563 = ~n37741 & ~n39530;
  assign n39564 = n7728 & ~n39563;
  assign n39565 = ~n37857 & ~n39530;
  assign n39566 = ~n7728 & ~n39565;
  assign n39567 = ~n39564 & ~n39566;
  assign n39568 = ~n7723 & ~n39567;
  assign n39569 = ~n39562 & ~n39568;
  assign n39570 = ~n7714 & ~n39569;
  assign n39571 = ~n39561 & ~n39570;
  assign n39572 = ~n7705 & ~n39571;
  assign n39573 = ~n39552 & ~n39572;
  assign n39574 = n7808 & ~n39573;
  assign n39575 = ~n39540 & ~n39574;
  assign n39576 = n8195 & ~n39575;
  assign n39577 = ~n8196 & ~n39576;
  assign n39578 = ~n8193 & ~n39577;
  assign n39579 = ~n9900 & ~n39530;
  assign n39580 = ~n7723 & ~n39579;
  assign n39581 = ~n9899 & ~n39580;
  assign n39582 = n7714 & ~n39581;
  assign n39583 = ~n39536 & ~n39582;
  assign n39584 = ~n7705 & ~n39583;
  assign n39585 = ~n9898 & ~n39584;
  assign n39586 = ~n7808 & ~n39585;
  assign n39587 = ~n38371 & ~n39530;
  assign n39588 = n7728 & ~n39587;
  assign n39589 = ~n39566 & ~n39588;
  assign n39590 = ~n7723 & ~n39589;
  assign n39591 = ~n38077 & ~n39590;
  assign n39592 = ~n7714 & ~n39591;
  assign n39593 = ~n38076 & ~n39592;
  assign n39594 = ~n7705 & ~n39593;
  assign n39595 = ~n22399 & ~n39594;
  assign n39596 = n7808 & ~n39595;
  assign n39597 = ~n39586 & ~n39596;
  assign n39598 = ~n8195 & ~n39597;
  assign n39599 = ~n11966 & ~n39075;
  assign n39600 = i_hlock7 & ~n39599;
  assign n39601 = ~n11974 & ~n39075;
  assign n39602 = ~i_hlock7 & ~n39601;
  assign n39603 = ~n39600 & ~n39602;
  assign n39604 = i_hbusreq7 & ~n39603;
  assign n39605 = ~n11990 & ~n39086;
  assign n39606 = i_hlock7 & ~n39605;
  assign n39607 = ~n12004 & ~n39086;
  assign n39608 = ~i_hlock7 & ~n39607;
  assign n39609 = ~n39606 & ~n39608;
  assign n39610 = ~i_hbusreq7 & ~n39609;
  assign n39611 = ~n39604 & ~n39610;
  assign n39612 = n7924 & ~n39611;
  assign n39613 = ~n10375 & ~n39612;
  assign n39614 = n8214 & ~n39613;
  assign n39615 = n8214 & ~n39614;
  assign n39616 = n8202 & ~n39615;
  assign n39617 = ~n10332 & ~n39616;
  assign n39618 = n7728 & ~n39617;
  assign n39619 = n8214 & ~n39529;
  assign n39620 = ~n8336 & ~n39619;
  assign n39621 = n8202 & ~n39620;
  assign n39622 = ~n10649 & ~n39621;
  assign n39623 = ~n7728 & ~n39622;
  assign n39624 = ~n39618 & ~n39623;
  assign n39625 = ~n7723 & ~n39624;
  assign n39626 = ~n7723 & ~n39625;
  assign n39627 = ~n7714 & ~n39626;
  assign n39628 = ~n7714 & ~n39627;
  assign n39629 = n7705 & ~n39628;
  assign n39630 = n7723 & ~n39622;
  assign n39631 = n7920 & ~n39622;
  assign n39632 = ~n39530 & ~n39631;
  assign n39633 = ~n7723 & ~n39632;
  assign n39634 = ~n39630 & ~n39633;
  assign n39635 = n7714 & ~n39634;
  assign n39636 = ~n39536 & ~n39635;
  assign n39637 = ~n7705 & ~n39636;
  assign n39638 = ~n39629 & ~n39637;
  assign n39639 = ~n7808 & ~n39638;
  assign n39640 = ~n7920 & ~n39617;
  assign n39641 = ~n38572 & ~n39640;
  assign n39642 = n7728 & ~n39641;
  assign n39643 = ~n7920 & ~n39622;
  assign n39644 = ~n38582 & ~n39643;
  assign n39645 = ~n7728 & ~n39644;
  assign n39646 = ~n39642 & ~n39645;
  assign n39647 = ~n7723 & ~n39646;
  assign n39648 = ~n7723 & ~n39647;
  assign n39649 = ~n7714 & ~n39648;
  assign n39650 = ~n7714 & ~n39649;
  assign n39651 = n7705 & ~n39650;
  assign n39652 = ~n38623 & ~n39643;
  assign n39653 = n7728 & ~n39652;
  assign n39654 = ~n38741 & ~n39643;
  assign n39655 = ~n7728 & ~n39654;
  assign n39656 = ~n39653 & ~n39655;
  assign n39657 = n7723 & ~n39656;
  assign n39658 = ~n7723 & ~n39654;
  assign n39659 = ~n39657 & ~n39658;
  assign n39660 = n7714 & ~n39659;
  assign n39661 = n7723 & ~n39654;
  assign n39662 = ~n38947 & ~n39530;
  assign n39663 = n7728 & ~n39662;
  assign n39664 = ~n39566 & ~n39663;
  assign n39665 = ~n7723 & ~n39664;
  assign n39666 = ~n39661 & ~n39665;
  assign n39667 = ~n7714 & ~n39666;
  assign n39668 = ~n39660 & ~n39667;
  assign n39669 = ~n7705 & ~n39668;
  assign n39670 = ~n39651 & ~n39669;
  assign n39671 = n7808 & ~n39670;
  assign n39672 = ~n39639 & ~n39671;
  assign n39673 = n8195 & ~n39672;
  assign n39674 = ~n39598 & ~n39673;
  assign n39675 = n8193 & ~n39674;
  assign n39676 = ~n39578 & ~n39675;
  assign n39677 = ~n8191 & ~n39676;
  assign n39678 = ~n39503 & ~n39677;
  assign n39679 = ~n8188 & ~n39678;
  assign n39680 = ~n39329 & ~n39679;
  assign n39681 = ~n8185 & ~n39680;
  assign n39682 = ~n39159 & ~n39681;
  assign n39683 = controllable_hgrant8 & ~n39682;
  assign n39684 = ~n8172 & ~n8195;
  assign n39685 = ~n8217 & ~n28605;
  assign n39686 = ~n8217 & ~n39685;
  assign n39687 = i_hlock6 & ~n39686;
  assign n39688 = ~n8217 & ~n28623;
  assign n39689 = ~n8217 & ~n39688;
  assign n39690 = ~i_hlock6 & ~n39689;
  assign n39691 = ~n39687 & ~n39690;
  assign n39692 = controllable_hgrant6 & ~n39691;
  assign n39693 = ~controllable_hgrant6 & ~n8245;
  assign n39694 = ~n39692 & ~n39693;
  assign n39695 = ~controllable_hmaster0 & ~n39694;
  assign n39696 = ~controllable_hmaster0 & ~n39695;
  assign n39697 = ~controllable_hmaster3 & ~n39696;
  assign n39698 = ~controllable_hmaster3 & ~n39697;
  assign n39699 = i_hbusreq7 & ~n39698;
  assign n39700 = i_hbusreq8 & ~n39696;
  assign n39701 = i_hbusreq6 & ~n39691;
  assign n39702 = ~n8217 & ~n28654;
  assign n39703 = ~n8217 & ~n39702;
  assign n39704 = i_hlock6 & ~n39703;
  assign n39705 = ~n8217 & ~n28687;
  assign n39706 = ~n8217 & ~n39705;
  assign n39707 = ~i_hlock6 & ~n39706;
  assign n39708 = ~n39704 & ~n39707;
  assign n39709 = ~i_hbusreq6 & ~n39708;
  assign n39710 = ~n39701 & ~n39709;
  assign n39711 = controllable_hgrant6 & ~n39710;
  assign n39712 = ~controllable_hgrant6 & ~n8319;
  assign n39713 = ~n39711 & ~n39712;
  assign n39714 = ~controllable_hmaster0 & ~n39713;
  assign n39715 = ~controllable_hmaster0 & ~n39714;
  assign n39716 = ~i_hbusreq8 & ~n39715;
  assign n39717 = ~n39700 & ~n39716;
  assign n39718 = ~controllable_hmaster3 & ~n39717;
  assign n39719 = ~controllable_hmaster3 & ~n39718;
  assign n39720 = ~i_hbusreq7 & ~n39719;
  assign n39721 = ~n39699 & ~n39720;
  assign n39722 = n7924 & ~n39721;
  assign n39723 = n7924 & ~n39722;
  assign n39724 = n8214 & ~n39723;
  assign n39725 = n8214 & ~n39724;
  assign n39726 = n8202 & ~n39725;
  assign n39727 = n8202 & ~n39726;
  assign n39728 = n7728 & ~n39727;
  assign n39729 = ~n7904 & ~n8202;
  assign n39730 = ~n7904 & ~n8214;
  assign n39731 = ~n7904 & ~n7924;
  assign n39732 = ~n7840 & ~n39697;
  assign n39733 = i_hbusreq7 & ~n39732;
  assign n39734 = ~n7901 & ~n39718;
  assign n39735 = ~i_hbusreq7 & ~n39734;
  assign n39736 = ~n39733 & ~n39735;
  assign n39737 = n7924 & ~n39736;
  assign n39738 = ~n39731 & ~n39737;
  assign n39739 = n8214 & ~n39738;
  assign n39740 = ~n39730 & ~n39739;
  assign n39741 = n8202 & ~n39740;
  assign n39742 = ~n39729 & ~n39741;
  assign n39743 = ~n7728 & ~n39742;
  assign n39744 = ~n39728 & ~n39743;
  assign n39745 = ~n7723 & ~n39744;
  assign n39746 = ~n7723 & ~n39745;
  assign n39747 = ~n7714 & ~n39746;
  assign n39748 = ~n7714 & ~n39747;
  assign n39749 = n7705 & ~n39748;
  assign n39750 = n7723 & ~n39742;
  assign n39751 = controllable_hgrant6 & ~n8361;
  assign n39752 = ~controllable_hgrant1 & ~n7822;
  assign n39753 = ~n13155 & ~n39752;
  assign n39754 = ~controllable_hgrant3 & ~n39753;
  assign n39755 = ~n13154 & ~n39754;
  assign n39756 = ~controllable_hgrant4 & ~n39755;
  assign n39757 = ~n13153 & ~n39756;
  assign n39758 = ~controllable_hgrant5 & ~n39757;
  assign n39759 = ~n13152 & ~n39758;
  assign n39760 = controllable_hmaster1 & ~n39759;
  assign n39761 = controllable_hmaster2 & ~n39759;
  assign n39762 = controllable_hmaster2 & ~n39761;
  assign n39763 = ~controllable_hmaster1 & ~n39762;
  assign n39764 = ~n39760 & ~n39763;
  assign n39765 = ~controllable_hgrant6 & ~n39764;
  assign n39766 = ~n39751 & ~n39765;
  assign n39767 = controllable_hmaster3 & ~n39766;
  assign n39768 = controllable_hgrant6 & ~n8400;
  assign n39769 = controllable_hgrant5 & ~n8372;
  assign n39770 = controllable_hgrant4 & ~n8372;
  assign n39771 = ~n8365 & ~n16132;
  assign n39772 = ~n8365 & ~n39771;
  assign n39773 = i_hlock3 & ~n39772;
  assign n39774 = ~n8365 & ~n16150;
  assign n39775 = ~n8365 & ~n39774;
  assign n39776 = ~i_hlock3 & ~n39775;
  assign n39777 = ~n39773 & ~n39776;
  assign n39778 = controllable_hgrant3 & ~n39777;
  assign n39779 = ~controllable_hgrant3 & ~n8372;
  assign n39780 = ~n39778 & ~n39779;
  assign n39781 = ~controllable_hgrant4 & ~n39780;
  assign n39782 = ~n39770 & ~n39781;
  assign n39783 = ~controllable_hgrant5 & ~n39782;
  assign n39784 = ~n39769 & ~n39783;
  assign n39785 = ~controllable_hmaster2 & ~n39784;
  assign n39786 = ~controllable_hmaster2 & ~n39785;
  assign n39787 = controllable_hmaster1 & ~n39786;
  assign n39788 = ~n8378 & ~n28599;
  assign n39789 = ~n8378 & ~n39788;
  assign n39790 = i_hlock5 & ~n39789;
  assign n39791 = ~n8378 & ~n28617;
  assign n39792 = ~n8378 & ~n39791;
  assign n39793 = ~i_hlock5 & ~n39792;
  assign n39794 = ~n39790 & ~n39793;
  assign n39795 = controllable_hgrant5 & ~n39794;
  assign n39796 = ~controllable_hgrant5 & ~n8385;
  assign n39797 = ~n39795 & ~n39796;
  assign n39798 = controllable_hmaster2 & ~n39797;
  assign n39799 = controllable_hgrant5 & ~n8396;
  assign n39800 = controllable_hgrant4 & ~n8396;
  assign n39801 = controllable_hgrant3 & ~n8396;
  assign n39802 = ~n8389 & ~n16130;
  assign n39803 = ~n8389 & ~n39802;
  assign n39804 = i_hlock1 & ~n39803;
  assign n39805 = ~n8389 & ~n16148;
  assign n39806 = ~n8389 & ~n39805;
  assign n39807 = ~i_hlock1 & ~n39806;
  assign n39808 = ~n39804 & ~n39807;
  assign n39809 = controllable_hgrant1 & ~n39808;
  assign n39810 = ~controllable_hgrant1 & ~n8396;
  assign n39811 = ~n39809 & ~n39810;
  assign n39812 = ~controllable_hgrant3 & ~n39811;
  assign n39813 = ~n39801 & ~n39812;
  assign n39814 = ~controllable_hgrant4 & ~n39813;
  assign n39815 = ~n39800 & ~n39814;
  assign n39816 = ~controllable_hgrant5 & ~n39815;
  assign n39817 = ~n39799 & ~n39816;
  assign n39818 = ~controllable_hmaster2 & ~n39817;
  assign n39819 = ~n39798 & ~n39818;
  assign n39820 = ~controllable_hmaster1 & ~n39819;
  assign n39821 = ~n39787 & ~n39820;
  assign n39822 = ~controllable_hgrant6 & ~n39821;
  assign n39823 = ~n39768 & ~n39822;
  assign n39824 = controllable_hmaster0 & ~n39823;
  assign n39825 = ~n8421 & ~n28602;
  assign n39826 = controllable_hmaster1 & ~n39825;
  assign n39827 = ~n8445 & ~n39826;
  assign n39828 = ~n8217 & ~n39827;
  assign n39829 = ~n8447 & ~n39828;
  assign n39830 = i_hlock6 & ~n39829;
  assign n39831 = ~n8421 & ~n28620;
  assign n39832 = controllable_hmaster1 & ~n39831;
  assign n39833 = ~n8445 & ~n39832;
  assign n39834 = ~n8217 & ~n39833;
  assign n39835 = ~n8447 & ~n39834;
  assign n39836 = ~i_hlock6 & ~n39835;
  assign n39837 = ~n39830 & ~n39836;
  assign n39838 = controllable_hgrant6 & ~n39837;
  assign n39839 = controllable_hgrant5 & ~n8420;
  assign n39840 = controllable_hgrant4 & ~n8420;
  assign n39841 = controllable_hgrant3 & ~n8420;
  assign n39842 = controllable_hgrant1 & ~n8420;
  assign n39843 = controllable_hmastlock & n8404;
  assign n39844 = controllable_hmastlock & ~n39843;
  assign n39845 = controllable_locked & ~n39844;
  assign n39846 = controllable_ndecide & n8404;
  assign n39847 = controllable_ndecide & ~n39846;
  assign n39848 = ~controllable_hmastlock & ~n39847;
  assign n39849 = ~n8409 & ~n39848;
  assign n39850 = ~controllable_locked & ~n39849;
  assign n39851 = ~n39845 & ~n39850;
  assign n39852 = i_hlock2 & ~n39851;
  assign n39853 = controllable_hmastlock & ~n39847;
  assign n39854 = ~n8412 & ~n39853;
  assign n39855 = controllable_locked & ~n39854;
  assign n39856 = ~controllable_hmastlock & n8404;
  assign n39857 = ~controllable_hmastlock & ~n39856;
  assign n39858 = ~controllable_locked & ~n39857;
  assign n39859 = ~n39855 & ~n39858;
  assign n39860 = ~i_hlock2 & ~n39859;
  assign n39861 = ~n39852 & ~n39860;
  assign n39862 = controllable_hgrant2 & ~n39861;
  assign n39863 = ~controllable_hgrant2 & ~n8415;
  assign n39864 = ~n39862 & ~n39863;
  assign n39865 = ~n7733 & ~n39864;
  assign n39866 = ~n7733 & ~n39865;
  assign n39867 = ~n7928 & ~n39866;
  assign n39868 = n7928 & ~n39864;
  assign n39869 = ~n39867 & ~n39868;
  assign n39870 = ~controllable_hgrant1 & ~n39869;
  assign n39871 = ~n39842 & ~n39870;
  assign n39872 = ~controllable_hgrant3 & ~n39871;
  assign n39873 = ~n39841 & ~n39872;
  assign n39874 = ~controllable_hgrant4 & ~n39873;
  assign n39875 = ~n39840 & ~n39874;
  assign n39876 = ~controllable_hgrant5 & ~n39875;
  assign n39877 = ~n39839 & ~n39876;
  assign n39878 = ~controllable_hmaster2 & ~n39877;
  assign n39879 = ~controllable_hmaster2 & ~n39878;
  assign n39880 = controllable_hmaster1 & ~n39879;
  assign n39881 = controllable_hgrant5 & ~n8433;
  assign n39882 = ~n8426 & ~n16134;
  assign n39883 = ~n8426 & ~n39882;
  assign n39884 = i_hlock4 & ~n39883;
  assign n39885 = ~n8426 & ~n16152;
  assign n39886 = ~n8426 & ~n39885;
  assign n39887 = ~i_hlock4 & ~n39886;
  assign n39888 = ~n39884 & ~n39887;
  assign n39889 = controllable_hgrant4 & ~n39888;
  assign n39890 = ~controllable_hgrant4 & ~n8433;
  assign n39891 = ~n39889 & ~n39890;
  assign n39892 = ~controllable_hgrant5 & ~n39891;
  assign n39893 = ~n39881 & ~n39892;
  assign n39894 = controllable_hmaster2 & ~n39893;
  assign n39895 = ~n8443 & ~n39894;
  assign n39896 = ~controllable_hmaster1 & ~n39895;
  assign n39897 = ~n39880 & ~n39896;
  assign n39898 = n8217 & ~n39897;
  assign n39899 = ~n8224 & ~n39878;
  assign n39900 = controllable_hmaster1 & ~n39899;
  assign n39901 = ~n39896 & ~n39900;
  assign n39902 = ~n8217 & ~n39901;
  assign n39903 = ~n39898 & ~n39902;
  assign n39904 = i_hlock6 & ~n39903;
  assign n39905 = ~n8238 & ~n39878;
  assign n39906 = controllable_hmaster1 & ~n39905;
  assign n39907 = ~n39896 & ~n39906;
  assign n39908 = ~n8217 & ~n39907;
  assign n39909 = ~n39898 & ~n39908;
  assign n39910 = ~i_hlock6 & ~n39909;
  assign n39911 = ~n39904 & ~n39910;
  assign n39912 = ~controllable_hgrant6 & ~n39911;
  assign n39913 = ~n39838 & ~n39912;
  assign n39914 = ~controllable_hmaster0 & ~n39913;
  assign n39915 = ~n39824 & ~n39914;
  assign n39916 = ~controllable_hmaster3 & ~n39915;
  assign n39917 = ~n39767 & ~n39916;
  assign n39918 = i_hbusreq7 & ~n39917;
  assign n39919 = i_hbusreq8 & ~n39766;
  assign n39920 = controllable_hgrant6 & ~n8489;
  assign n39921 = i_hbusreq6 & ~n39764;
  assign n39922 = i_hbusreq5 & ~n39757;
  assign n39923 = i_hbusreq4 & ~n39755;
  assign n39924 = i_hbusreq9 & ~n39755;
  assign n39925 = i_hbusreq3 & ~n39753;
  assign n39926 = i_hbusreq1 & ~n7822;
  assign n39927 = ~i_hbusreq1 & ~n7869;
  assign n39928 = ~n39926 & ~n39927;
  assign n39929 = ~controllable_hgrant1 & ~n39928;
  assign n39930 = ~n13213 & ~n39929;
  assign n39931 = ~i_hbusreq3 & ~n39930;
  assign n39932 = ~n39925 & ~n39931;
  assign n39933 = ~controllable_hgrant3 & ~n39932;
  assign n39934 = ~n13211 & ~n39933;
  assign n39935 = ~i_hbusreq9 & ~n39934;
  assign n39936 = ~n39924 & ~n39935;
  assign n39937 = ~i_hbusreq4 & ~n39936;
  assign n39938 = ~n39923 & ~n39937;
  assign n39939 = ~controllable_hgrant4 & ~n39938;
  assign n39940 = ~n13208 & ~n39939;
  assign n39941 = ~i_hbusreq5 & ~n39940;
  assign n39942 = ~n39922 & ~n39941;
  assign n39943 = ~controllable_hgrant5 & ~n39942;
  assign n39944 = ~n13206 & ~n39943;
  assign n39945 = controllable_hmaster1 & ~n39944;
  assign n39946 = controllable_hmaster2 & ~n39944;
  assign n39947 = controllable_hmaster2 & ~n39946;
  assign n39948 = ~controllable_hmaster1 & ~n39947;
  assign n39949 = ~n39945 & ~n39948;
  assign n39950 = ~i_hbusreq6 & ~n39949;
  assign n39951 = ~n39921 & ~n39950;
  assign n39952 = ~controllable_hgrant6 & ~n39951;
  assign n39953 = ~n39920 & ~n39952;
  assign n39954 = ~i_hbusreq8 & ~n39953;
  assign n39955 = ~n39919 & ~n39954;
  assign n39956 = controllable_hmaster3 & ~n39955;
  assign n39957 = i_hbusreq8 & ~n39915;
  assign n39958 = controllable_hgrant6 & ~n8555;
  assign n39959 = i_hbusreq6 & ~n39821;
  assign n39960 = controllable_hgrant5 & ~n8513;
  assign n39961 = i_hbusreq5 & ~n39782;
  assign n39962 = controllable_hgrant4 & ~n8511;
  assign n39963 = i_hbusreq4 & ~n39780;
  assign n39964 = i_hbusreq9 & ~n39780;
  assign n39965 = i_hbusreq3 & ~n39777;
  assign n39966 = ~n8365 & ~n16197;
  assign n39967 = ~n8365 & ~n39966;
  assign n39968 = i_hlock3 & ~n39967;
  assign n39969 = ~n8365 & ~n16222;
  assign n39970 = ~n8365 & ~n39969;
  assign n39971 = ~i_hlock3 & ~n39970;
  assign n39972 = ~n39968 & ~n39971;
  assign n39973 = ~i_hbusreq3 & ~n39972;
  assign n39974 = ~n39965 & ~n39973;
  assign n39975 = controllable_hgrant3 & ~n39974;
  assign n39976 = ~controllable_hgrant3 & ~n8507;
  assign n39977 = ~n39975 & ~n39976;
  assign n39978 = ~i_hbusreq9 & ~n39977;
  assign n39979 = ~n39964 & ~n39978;
  assign n39980 = ~i_hbusreq4 & ~n39979;
  assign n39981 = ~n39963 & ~n39980;
  assign n39982 = ~controllable_hgrant4 & ~n39981;
  assign n39983 = ~n39962 & ~n39982;
  assign n39984 = ~i_hbusreq5 & ~n39983;
  assign n39985 = ~n39961 & ~n39984;
  assign n39986 = ~controllable_hgrant5 & ~n39985;
  assign n39987 = ~n39960 & ~n39986;
  assign n39988 = ~controllable_hmaster2 & ~n39987;
  assign n39989 = ~controllable_hmaster2 & ~n39988;
  assign n39990 = controllable_hmaster1 & ~n39989;
  assign n39991 = i_hbusreq5 & ~n39794;
  assign n39992 = ~n8378 & ~n28646;
  assign n39993 = ~n8378 & ~n39992;
  assign n39994 = i_hlock5 & ~n39993;
  assign n39995 = ~n8378 & ~n28679;
  assign n39996 = ~n8378 & ~n39995;
  assign n39997 = ~i_hlock5 & ~n39996;
  assign n39998 = ~n39994 & ~n39997;
  assign n39999 = ~i_hbusreq5 & ~n39998;
  assign n40000 = ~n39991 & ~n39999;
  assign n40001 = controllable_hgrant5 & ~n40000;
  assign n40002 = ~controllable_hgrant5 & ~n8526;
  assign n40003 = ~n40001 & ~n40002;
  assign n40004 = controllable_hmaster2 & ~n40003;
  assign n40005 = controllable_hgrant5 & ~n8549;
  assign n40006 = i_hbusreq5 & ~n39815;
  assign n40007 = controllable_hgrant4 & ~n8547;
  assign n40008 = i_hbusreq4 & ~n39813;
  assign n40009 = i_hbusreq9 & ~n39813;
  assign n40010 = controllable_hgrant3 & ~n8543;
  assign n40011 = i_hbusreq3 & ~n39811;
  assign n40012 = i_hbusreq1 & ~n39808;
  assign n40013 = ~n8389 & ~n16193;
  assign n40014 = ~n8389 & ~n40013;
  assign n40015 = i_hlock1 & ~n40014;
  assign n40016 = ~n8389 & ~n16218;
  assign n40017 = ~n8389 & ~n40016;
  assign n40018 = ~i_hlock1 & ~n40017;
  assign n40019 = ~n40015 & ~n40018;
  assign n40020 = ~i_hbusreq1 & ~n40019;
  assign n40021 = ~n40012 & ~n40020;
  assign n40022 = controllable_hgrant1 & ~n40021;
  assign n40023 = ~controllable_hgrant1 & ~n8541;
  assign n40024 = ~n40022 & ~n40023;
  assign n40025 = ~i_hbusreq3 & ~n40024;
  assign n40026 = ~n40011 & ~n40025;
  assign n40027 = ~controllable_hgrant3 & ~n40026;
  assign n40028 = ~n40010 & ~n40027;
  assign n40029 = ~i_hbusreq9 & ~n40028;
  assign n40030 = ~n40009 & ~n40029;
  assign n40031 = ~i_hbusreq4 & ~n40030;
  assign n40032 = ~n40008 & ~n40031;
  assign n40033 = ~controllable_hgrant4 & ~n40032;
  assign n40034 = ~n40007 & ~n40033;
  assign n40035 = ~i_hbusreq5 & ~n40034;
  assign n40036 = ~n40006 & ~n40035;
  assign n40037 = ~controllable_hgrant5 & ~n40036;
  assign n40038 = ~n40005 & ~n40037;
  assign n40039 = ~controllable_hmaster2 & ~n40038;
  assign n40040 = ~n40004 & ~n40039;
  assign n40041 = ~controllable_hmaster1 & ~n40040;
  assign n40042 = ~n39990 & ~n40041;
  assign n40043 = ~i_hbusreq6 & ~n40042;
  assign n40044 = ~n39959 & ~n40043;
  assign n40045 = ~controllable_hgrant6 & ~n40044;
  assign n40046 = ~n39958 & ~n40045;
  assign n40047 = controllable_hmaster0 & ~n40046;
  assign n40048 = i_hbusreq6 & ~n39837;
  assign n40049 = ~n8588 & ~n28651;
  assign n40050 = controllable_hmaster1 & ~n40049;
  assign n40051 = ~n8612 & ~n40050;
  assign n40052 = ~n8217 & ~n40051;
  assign n40053 = ~n8614 & ~n40052;
  assign n40054 = i_hlock6 & ~n40053;
  assign n40055 = ~n8588 & ~n28684;
  assign n40056 = controllable_hmaster1 & ~n40055;
  assign n40057 = ~n8612 & ~n40056;
  assign n40058 = ~n8217 & ~n40057;
  assign n40059 = ~n8614 & ~n40058;
  assign n40060 = ~i_hlock6 & ~n40059;
  assign n40061 = ~n40054 & ~n40060;
  assign n40062 = ~i_hbusreq6 & ~n40061;
  assign n40063 = ~n40048 & ~n40062;
  assign n40064 = controllable_hgrant6 & ~n40063;
  assign n40065 = i_hbusreq6 & ~n39911;
  assign n40066 = controllable_hgrant5 & ~n8587;
  assign n40067 = i_hbusreq5 & ~n39875;
  assign n40068 = controllable_hgrant4 & ~n8585;
  assign n40069 = i_hbusreq4 & ~n39873;
  assign n40070 = i_hbusreq9 & ~n39873;
  assign n40071 = controllable_hgrant3 & ~n8581;
  assign n40072 = i_hbusreq3 & ~n39871;
  assign n40073 = controllable_hgrant1 & ~n8579;
  assign n40074 = i_hbusreq1 & ~n39869;
  assign n40075 = i_hbusreq2 & ~n39861;
  assign n40076 = i_hbusreq0 & ~n39851;
  assign n40077 = controllable_hmastlock & ~n39853;
  assign n40078 = controllable_locked & ~n40077;
  assign n40079 = ~controllable_hmastlock & ~n39848;
  assign n40080 = ~controllable_locked & ~n40079;
  assign n40081 = ~n40078 & ~n40080;
  assign n40082 = ~i_hbusreq0 & ~n40081;
  assign n40083 = ~n40076 & ~n40082;
  assign n40084 = i_hlock2 & ~n40083;
  assign n40085 = i_hbusreq0 & ~n39859;
  assign n40086 = ~n40082 & ~n40085;
  assign n40087 = ~i_hlock2 & ~n40086;
  assign n40088 = ~n40084 & ~n40087;
  assign n40089 = ~i_hbusreq2 & ~n40088;
  assign n40090 = ~n40075 & ~n40089;
  assign n40091 = controllable_hgrant2 & ~n40090;
  assign n40092 = ~controllable_hgrant2 & ~n8572;
  assign n40093 = ~n40091 & ~n40092;
  assign n40094 = ~n7733 & ~n40093;
  assign n40095 = ~n7733 & ~n40094;
  assign n40096 = ~n7928 & ~n40095;
  assign n40097 = n7928 & ~n40093;
  assign n40098 = ~n40096 & ~n40097;
  assign n40099 = ~i_hbusreq1 & ~n40098;
  assign n40100 = ~n40074 & ~n40099;
  assign n40101 = ~controllable_hgrant1 & ~n40100;
  assign n40102 = ~n40073 & ~n40101;
  assign n40103 = ~i_hbusreq3 & ~n40102;
  assign n40104 = ~n40072 & ~n40103;
  assign n40105 = ~controllable_hgrant3 & ~n40104;
  assign n40106 = ~n40071 & ~n40105;
  assign n40107 = ~i_hbusreq9 & ~n40106;
  assign n40108 = ~n40070 & ~n40107;
  assign n40109 = ~i_hbusreq4 & ~n40108;
  assign n40110 = ~n40069 & ~n40109;
  assign n40111 = ~controllable_hgrant4 & ~n40110;
  assign n40112 = ~n40068 & ~n40111;
  assign n40113 = ~i_hbusreq5 & ~n40112;
  assign n40114 = ~n40067 & ~n40113;
  assign n40115 = ~controllable_hgrant5 & ~n40114;
  assign n40116 = ~n40066 & ~n40115;
  assign n40117 = ~controllable_hmaster2 & ~n40116;
  assign n40118 = ~controllable_hmaster2 & ~n40117;
  assign n40119 = controllable_hmaster1 & ~n40118;
  assign n40120 = controllable_hgrant5 & ~n8609;
  assign n40121 = i_hbusreq5 & ~n39891;
  assign n40122 = i_hbusreq4 & ~n39888;
  assign n40123 = i_hbusreq9 & ~n39883;
  assign n40124 = ~n8426 & ~n16201;
  assign n40125 = ~n8426 & ~n40124;
  assign n40126 = ~i_hbusreq9 & ~n40125;
  assign n40127 = ~n40123 & ~n40126;
  assign n40128 = i_hlock4 & ~n40127;
  assign n40129 = i_hbusreq9 & ~n39886;
  assign n40130 = ~n8426 & ~n16226;
  assign n40131 = ~n8426 & ~n40130;
  assign n40132 = ~i_hbusreq9 & ~n40131;
  assign n40133 = ~n40129 & ~n40132;
  assign n40134 = ~i_hlock4 & ~n40133;
  assign n40135 = ~n40128 & ~n40134;
  assign n40136 = ~i_hbusreq4 & ~n40135;
  assign n40137 = ~n40122 & ~n40136;
  assign n40138 = controllable_hgrant4 & ~n40137;
  assign n40139 = ~controllable_hgrant4 & ~n8607;
  assign n40140 = ~n40138 & ~n40139;
  assign n40141 = ~i_hbusreq5 & ~n40140;
  assign n40142 = ~n40121 & ~n40141;
  assign n40143 = ~controllable_hgrant5 & ~n40142;
  assign n40144 = ~n40120 & ~n40143;
  assign n40145 = controllable_hmaster2 & ~n40144;
  assign n40146 = ~n8443 & ~n40145;
  assign n40147 = ~controllable_hmaster1 & ~n40146;
  assign n40148 = ~n40119 & ~n40147;
  assign n40149 = n8217 & ~n40148;
  assign n40150 = ~n8278 & ~n40117;
  assign n40151 = controllable_hmaster1 & ~n40150;
  assign n40152 = ~n40147 & ~n40151;
  assign n40153 = ~n8217 & ~n40152;
  assign n40154 = ~n40149 & ~n40153;
  assign n40155 = i_hlock6 & ~n40154;
  assign n40156 = ~n8310 & ~n40117;
  assign n40157 = controllable_hmaster1 & ~n40156;
  assign n40158 = ~n40147 & ~n40157;
  assign n40159 = ~n8217 & ~n40158;
  assign n40160 = ~n40149 & ~n40159;
  assign n40161 = ~i_hlock6 & ~n40160;
  assign n40162 = ~n40155 & ~n40161;
  assign n40163 = ~i_hbusreq6 & ~n40162;
  assign n40164 = ~n40065 & ~n40163;
  assign n40165 = ~controllable_hgrant6 & ~n40164;
  assign n40166 = ~n40064 & ~n40165;
  assign n40167 = ~controllable_hmaster0 & ~n40166;
  assign n40168 = ~n40047 & ~n40167;
  assign n40169 = ~i_hbusreq8 & ~n40168;
  assign n40170 = ~n39957 & ~n40169;
  assign n40171 = ~controllable_hmaster3 & ~n40170;
  assign n40172 = ~n39956 & ~n40171;
  assign n40173 = ~i_hbusreq7 & ~n40172;
  assign n40174 = ~n39918 & ~n40173;
  assign n40175 = n7924 & ~n40174;
  assign n40176 = ~n39731 & ~n40175;
  assign n40177 = ~n7920 & ~n40176;
  assign n40178 = n7920 & ~n39742;
  assign n40179 = ~n40177 & ~n40178;
  assign n40180 = ~n7723 & ~n40179;
  assign n40181 = ~n39750 & ~n40180;
  assign n40182 = n7714 & ~n40181;
  assign n40183 = ~n7714 & ~n40176;
  assign n40184 = ~n40182 & ~n40183;
  assign n40185 = ~n7705 & ~n40184;
  assign n40186 = ~n39749 & ~n40185;
  assign n40187 = ~n7808 & ~n40186;
  assign n40188 = ~n7920 & ~n39727;
  assign n40189 = n8217 & ~n8661;
  assign n40190 = ~n8217 & ~n28821;
  assign n40191 = ~n40189 & ~n40190;
  assign n40192 = controllable_hgrant6 & ~n40191;
  assign n40193 = n8378 & ~n8657;
  assign n40194 = ~n8378 & ~n28815;
  assign n40195 = ~n40193 & ~n40194;
  assign n40196 = controllable_hgrant5 & ~n40195;
  assign n40197 = n8426 & ~n8653;
  assign n40198 = ~n8426 & ~n16740;
  assign n40199 = ~n40197 & ~n40198;
  assign n40200 = i_hlock9 & ~n40199;
  assign n40201 = n8426 & ~n8655;
  assign n40202 = ~n8426 & ~n16759;
  assign n40203 = ~n40201 & ~n40202;
  assign n40204 = ~i_hlock9 & ~n40203;
  assign n40205 = ~n40200 & ~n40204;
  assign n40206 = controllable_hgrant4 & ~n40205;
  assign n40207 = n8365 & ~n8653;
  assign n40208 = ~n8365 & ~n16738;
  assign n40209 = ~n40207 & ~n40208;
  assign n40210 = controllable_hgrant3 & ~n40209;
  assign n40211 = n8389 & ~n8653;
  assign n40212 = ~n8389 & ~n16736;
  assign n40213 = ~n40211 & ~n40212;
  assign n40214 = controllable_hgrant1 & ~n40213;
  assign n40215 = controllable_ndecide & ~n8406;
  assign n40216 = ~n7734 & ~n40215;
  assign n40217 = ~controllable_locked & ~n40216;
  assign n40218 = ~n13008 & ~n40217;
  assign n40219 = controllable_hgrant2 & ~n40218;
  assign n40220 = ~n16998 & ~n40219;
  assign n40221 = ~n7733 & ~n40220;
  assign n40222 = ~controllable_hmastlock & ~n40216;
  assign n40223 = ~n7818 & ~n40222;
  assign n40224 = controllable_locked & ~n40223;
  assign n40225 = ~n40217 & ~n40224;
  assign n40226 = controllable_hgrant2 & ~n40225;
  assign n40227 = ~n16998 & ~n40226;
  assign n40228 = n7733 & ~n40227;
  assign n40229 = ~n40221 & ~n40228;
  assign n40230 = n7928 & ~n40229;
  assign n40231 = ~n8221 & ~n40230;
  assign n40232 = ~controllable_hgrant1 & ~n40231;
  assign n40233 = ~n40214 & ~n40232;
  assign n40234 = ~controllable_hgrant3 & ~n40233;
  assign n40235 = ~n40210 & ~n40234;
  assign n40236 = i_hlock9 & ~n40235;
  assign n40237 = n8365 & ~n8655;
  assign n40238 = ~n8365 & ~n16757;
  assign n40239 = ~n40237 & ~n40238;
  assign n40240 = controllable_hgrant3 & ~n40239;
  assign n40241 = n8389 & ~n8655;
  assign n40242 = ~n8389 & ~n16755;
  assign n40243 = ~n40241 & ~n40242;
  assign n40244 = controllable_hgrant1 & ~n40243;
  assign n40245 = ~n8235 & ~n40230;
  assign n40246 = ~controllable_hgrant1 & ~n40245;
  assign n40247 = ~n40244 & ~n40246;
  assign n40248 = ~controllable_hgrant3 & ~n40247;
  assign n40249 = ~n40240 & ~n40248;
  assign n40250 = ~i_hlock9 & ~n40249;
  assign n40251 = ~n40236 & ~n40250;
  assign n40252 = ~controllable_hgrant4 & ~n40251;
  assign n40253 = ~n40206 & ~n40252;
  assign n40254 = ~controllable_hgrant5 & ~n40253;
  assign n40255 = ~n40196 & ~n40254;
  assign n40256 = ~controllable_hmaster2 & ~n40255;
  assign n40257 = ~controllable_hmaster2 & ~n40256;
  assign n40258 = ~controllable_hmaster1 & ~n40257;
  assign n40259 = ~controllable_hmaster1 & ~n40258;
  assign n40260 = ~controllable_hgrant6 & ~n40259;
  assign n40261 = ~n40192 & ~n40260;
  assign n40262 = controllable_hmaster0 & ~n40261;
  assign n40263 = controllable_hmaster0 & ~n40262;
  assign n40264 = controllable_hmaster3 & ~n40263;
  assign n40265 = controllable_hmaster3 & ~n40264;
  assign n40266 = i_hbusreq7 & ~n40265;
  assign n40267 = i_hbusreq8 & ~n40263;
  assign n40268 = i_hbusreq6 & ~n40191;
  assign n40269 = n8217 & ~n8714;
  assign n40270 = ~n8217 & ~n28850;
  assign n40271 = ~n40269 & ~n40270;
  assign n40272 = ~i_hbusreq6 & ~n40271;
  assign n40273 = ~n40268 & ~n40272;
  assign n40274 = controllable_hgrant6 & ~n40273;
  assign n40275 = i_hbusreq6 & ~n40259;
  assign n40276 = i_hbusreq5 & ~n40195;
  assign n40277 = n8378 & ~n8708;
  assign n40278 = ~n8378 & ~n28842;
  assign n40279 = ~n40277 & ~n40278;
  assign n40280 = ~i_hbusreq5 & ~n40279;
  assign n40281 = ~n40276 & ~n40280;
  assign n40282 = controllable_hgrant5 & ~n40281;
  assign n40283 = i_hbusreq5 & ~n40253;
  assign n40284 = i_hbusreq4 & ~n40205;
  assign n40285 = i_hbusreq9 & ~n40205;
  assign n40286 = n8426 & ~n8694;
  assign n40287 = ~n8426 & ~n16826;
  assign n40288 = ~n40286 & ~n40287;
  assign n40289 = i_hlock9 & ~n40288;
  assign n40290 = n8426 & ~n8702;
  assign n40291 = ~n8426 & ~n16863;
  assign n40292 = ~n40290 & ~n40291;
  assign n40293 = ~i_hlock9 & ~n40292;
  assign n40294 = ~n40289 & ~n40293;
  assign n40295 = ~i_hbusreq9 & ~n40294;
  assign n40296 = ~n40285 & ~n40295;
  assign n40297 = ~i_hbusreq4 & ~n40296;
  assign n40298 = ~n40284 & ~n40297;
  assign n40299 = controllable_hgrant4 & ~n40298;
  assign n40300 = i_hbusreq4 & ~n40251;
  assign n40301 = i_hbusreq9 & ~n40251;
  assign n40302 = i_hbusreq3 & ~n40209;
  assign n40303 = n8365 & ~n8692;
  assign n40304 = ~n8365 & ~n16822;
  assign n40305 = ~n40303 & ~n40304;
  assign n40306 = ~i_hbusreq3 & ~n40305;
  assign n40307 = ~n40302 & ~n40306;
  assign n40308 = controllable_hgrant3 & ~n40307;
  assign n40309 = i_hbusreq3 & ~n40233;
  assign n40310 = i_hbusreq1 & ~n40213;
  assign n40311 = n8389 & ~n8690;
  assign n40312 = ~n8389 & ~n16818;
  assign n40313 = ~n40311 & ~n40312;
  assign n40314 = ~i_hbusreq1 & ~n40313;
  assign n40315 = ~n40310 & ~n40314;
  assign n40316 = controllable_hgrant1 & ~n40315;
  assign n40317 = i_hbusreq1 & ~n40231;
  assign n40318 = i_hbusreq2 & ~n40218;
  assign n40319 = i_hbusreq0 & ~n40218;
  assign n40320 = controllable_ndecide & ~n40215;
  assign n40321 = ~controllable_locked & ~n40320;
  assign n40322 = ~controllable_locked & ~n40321;
  assign n40323 = i_hlock0 & ~n40322;
  assign n40324 = ~i_hlock0 & ~n40218;
  assign n40325 = ~n40323 & ~n40324;
  assign n40326 = ~i_hbusreq0 & ~n40325;
  assign n40327 = ~n40319 & ~n40326;
  assign n40328 = ~i_hbusreq2 & ~n40327;
  assign n40329 = ~n40318 & ~n40328;
  assign n40330 = controllable_hgrant2 & ~n40329;
  assign n40331 = ~n18216 & ~n40330;
  assign n40332 = ~n7733 & ~n40331;
  assign n40333 = i_hbusreq2 & ~n40225;
  assign n40334 = i_hbusreq0 & ~n40225;
  assign n40335 = ~controllable_hmastlock & ~n40222;
  assign n40336 = controllable_locked & ~n40335;
  assign n40337 = controllable_hmastlock & ~n40320;
  assign n40338 = ~n40222 & ~n40337;
  assign n40339 = ~controllable_locked & ~n40338;
  assign n40340 = ~n40336 & ~n40339;
  assign n40341 = i_hlock0 & ~n40340;
  assign n40342 = ~i_hlock0 & ~n40225;
  assign n40343 = ~n40341 & ~n40342;
  assign n40344 = ~i_hbusreq0 & ~n40343;
  assign n40345 = ~n40334 & ~n40344;
  assign n40346 = ~i_hbusreq2 & ~n40345;
  assign n40347 = ~n40333 & ~n40346;
  assign n40348 = controllable_hgrant2 & ~n40347;
  assign n40349 = i_hlock0 & ~n16803;
  assign n40350 = ~n18210 & ~n40349;
  assign n40351 = ~i_hbusreq0 & ~n40350;
  assign n40352 = ~n8106 & ~n40351;
  assign n40353 = ~i_hbusreq2 & ~n40352;
  assign n40354 = ~n8105 & ~n40353;
  assign n40355 = ~controllable_hgrant2 & ~n40354;
  assign n40356 = ~n40348 & ~n40355;
  assign n40357 = n7733 & ~n40356;
  assign n40358 = ~n40332 & ~n40357;
  assign n40359 = n7928 & ~n40358;
  assign n40360 = ~n8265 & ~n40359;
  assign n40361 = ~i_hbusreq1 & ~n40360;
  assign n40362 = ~n40317 & ~n40361;
  assign n40363 = ~controllable_hgrant1 & ~n40362;
  assign n40364 = ~n40316 & ~n40363;
  assign n40365 = ~i_hbusreq3 & ~n40364;
  assign n40366 = ~n40309 & ~n40365;
  assign n40367 = ~controllable_hgrant3 & ~n40366;
  assign n40368 = ~n40308 & ~n40367;
  assign n40369 = i_hlock9 & ~n40368;
  assign n40370 = i_hbusreq3 & ~n40239;
  assign n40371 = n8365 & ~n8700;
  assign n40372 = ~n8365 & ~n16859;
  assign n40373 = ~n40371 & ~n40372;
  assign n40374 = ~i_hbusreq3 & ~n40373;
  assign n40375 = ~n40370 & ~n40374;
  assign n40376 = controllable_hgrant3 & ~n40375;
  assign n40377 = i_hbusreq3 & ~n40247;
  assign n40378 = i_hbusreq1 & ~n40243;
  assign n40379 = n8389 & ~n8698;
  assign n40380 = ~n8389 & ~n16855;
  assign n40381 = ~n40379 & ~n40380;
  assign n40382 = ~i_hbusreq1 & ~n40381;
  assign n40383 = ~n40378 & ~n40382;
  assign n40384 = controllable_hgrant1 & ~n40383;
  assign n40385 = i_hbusreq1 & ~n40245;
  assign n40386 = ~n8297 & ~n40359;
  assign n40387 = ~i_hbusreq1 & ~n40386;
  assign n40388 = ~n40385 & ~n40387;
  assign n40389 = ~controllable_hgrant1 & ~n40388;
  assign n40390 = ~n40384 & ~n40389;
  assign n40391 = ~i_hbusreq3 & ~n40390;
  assign n40392 = ~n40377 & ~n40391;
  assign n40393 = ~controllable_hgrant3 & ~n40392;
  assign n40394 = ~n40376 & ~n40393;
  assign n40395 = ~i_hlock9 & ~n40394;
  assign n40396 = ~n40369 & ~n40395;
  assign n40397 = ~i_hbusreq9 & ~n40396;
  assign n40398 = ~n40301 & ~n40397;
  assign n40399 = ~i_hbusreq4 & ~n40398;
  assign n40400 = ~n40300 & ~n40399;
  assign n40401 = ~controllable_hgrant4 & ~n40400;
  assign n40402 = ~n40299 & ~n40401;
  assign n40403 = ~i_hbusreq5 & ~n40402;
  assign n40404 = ~n40283 & ~n40403;
  assign n40405 = ~controllable_hgrant5 & ~n40404;
  assign n40406 = ~n40282 & ~n40405;
  assign n40407 = ~controllable_hmaster2 & ~n40406;
  assign n40408 = ~controllable_hmaster2 & ~n40407;
  assign n40409 = ~controllable_hmaster1 & ~n40408;
  assign n40410 = ~controllable_hmaster1 & ~n40409;
  assign n40411 = ~i_hbusreq6 & ~n40410;
  assign n40412 = ~n40275 & ~n40411;
  assign n40413 = ~controllable_hgrant6 & ~n40412;
  assign n40414 = ~n40274 & ~n40413;
  assign n40415 = controllable_hmaster0 & ~n40414;
  assign n40416 = controllable_hmaster0 & ~n40415;
  assign n40417 = ~i_hbusreq8 & ~n40416;
  assign n40418 = ~n40267 & ~n40417;
  assign n40419 = controllable_hmaster3 & ~n40418;
  assign n40420 = controllable_hmaster3 & ~n40419;
  assign n40421 = ~i_hbusreq7 & ~n40420;
  assign n40422 = ~n40266 & ~n40421;
  assign n40423 = ~n8214 & ~n40422;
  assign n40424 = n8217 & ~n8729;
  assign n40425 = ~n8217 & ~n16748;
  assign n40426 = ~n40424 & ~n40425;
  assign n40427 = controllable_hgrant6 & ~n40426;
  assign n40428 = n8378 & ~n8653;
  assign n40429 = ~n8378 & ~n16742;
  assign n40430 = ~n40428 & ~n40429;
  assign n40431 = controllable_hgrant5 & ~n40430;
  assign n40432 = controllable_hgrant4 & ~n40199;
  assign n40433 = ~controllable_hgrant4 & ~n40235;
  assign n40434 = ~n40432 & ~n40433;
  assign n40435 = ~controllable_hgrant5 & ~n40434;
  assign n40436 = ~n40431 & ~n40435;
  assign n40437 = ~controllable_hmaster2 & ~n40436;
  assign n40438 = ~controllable_hmaster2 & ~n40437;
  assign n40439 = ~controllable_hmaster1 & ~n40438;
  assign n40440 = ~controllable_hmaster1 & ~n40439;
  assign n40441 = ~controllable_hgrant6 & ~n40440;
  assign n40442 = ~n40427 & ~n40441;
  assign n40443 = ~controllable_hmaster0 & ~n40442;
  assign n40444 = ~controllable_hmaster0 & ~n40443;
  assign n40445 = i_hlock8 & ~n40444;
  assign n40446 = n8217 & ~n8736;
  assign n40447 = ~n8217 & ~n16767;
  assign n40448 = ~n40446 & ~n40447;
  assign n40449 = controllable_hgrant6 & ~n40448;
  assign n40450 = n8378 & ~n8655;
  assign n40451 = ~n8378 & ~n16761;
  assign n40452 = ~n40450 & ~n40451;
  assign n40453 = controllable_hgrant5 & ~n40452;
  assign n40454 = controllable_hgrant4 & ~n40203;
  assign n40455 = ~controllable_hgrant4 & ~n40249;
  assign n40456 = ~n40454 & ~n40455;
  assign n40457 = ~controllable_hgrant5 & ~n40456;
  assign n40458 = ~n40453 & ~n40457;
  assign n40459 = ~controllable_hmaster2 & ~n40458;
  assign n40460 = ~controllable_hmaster2 & ~n40459;
  assign n40461 = ~controllable_hmaster1 & ~n40460;
  assign n40462 = ~controllable_hmaster1 & ~n40461;
  assign n40463 = ~controllable_hgrant6 & ~n40462;
  assign n40464 = ~n40449 & ~n40463;
  assign n40465 = ~controllable_hmaster0 & ~n40464;
  assign n40466 = ~controllable_hmaster0 & ~n40465;
  assign n40467 = ~i_hlock8 & ~n40466;
  assign n40468 = ~n40445 & ~n40467;
  assign n40469 = controllable_hmaster3 & ~n40468;
  assign n40470 = controllable_hmaster3 & ~n40469;
  assign n40471 = i_hbusreq7 & ~n40470;
  assign n40472 = i_hbusreq8 & ~n40468;
  assign n40473 = i_hbusreq6 & ~n40426;
  assign n40474 = n8217 & ~n8758;
  assign n40475 = ~n8217 & ~n16840;
  assign n40476 = ~n40474 & ~n40475;
  assign n40477 = ~i_hbusreq6 & ~n40476;
  assign n40478 = ~n40473 & ~n40477;
  assign n40479 = controllable_hgrant6 & ~n40478;
  assign n40480 = i_hbusreq6 & ~n40440;
  assign n40481 = i_hbusreq5 & ~n40430;
  assign n40482 = n8378 & ~n8752;
  assign n40483 = ~n8378 & ~n16832;
  assign n40484 = ~n40482 & ~n40483;
  assign n40485 = ~i_hbusreq5 & ~n40484;
  assign n40486 = ~n40481 & ~n40485;
  assign n40487 = controllable_hgrant5 & ~n40486;
  assign n40488 = i_hbusreq5 & ~n40434;
  assign n40489 = i_hbusreq4 & ~n40199;
  assign n40490 = i_hbusreq9 & ~n40199;
  assign n40491 = ~i_hbusreq9 & ~n40288;
  assign n40492 = ~n40490 & ~n40491;
  assign n40493 = ~i_hbusreq4 & ~n40492;
  assign n40494 = ~n40489 & ~n40493;
  assign n40495 = controllable_hgrant4 & ~n40494;
  assign n40496 = i_hbusreq4 & ~n40235;
  assign n40497 = i_hbusreq9 & ~n40235;
  assign n40498 = ~i_hbusreq9 & ~n40368;
  assign n40499 = ~n40497 & ~n40498;
  assign n40500 = ~i_hbusreq4 & ~n40499;
  assign n40501 = ~n40496 & ~n40500;
  assign n40502 = ~controllable_hgrant4 & ~n40501;
  assign n40503 = ~n40495 & ~n40502;
  assign n40504 = ~i_hbusreq5 & ~n40503;
  assign n40505 = ~n40488 & ~n40504;
  assign n40506 = ~controllable_hgrant5 & ~n40505;
  assign n40507 = ~n40487 & ~n40506;
  assign n40508 = ~controllable_hmaster2 & ~n40507;
  assign n40509 = ~controllable_hmaster2 & ~n40508;
  assign n40510 = ~controllable_hmaster1 & ~n40509;
  assign n40511 = ~controllable_hmaster1 & ~n40510;
  assign n40512 = ~i_hbusreq6 & ~n40511;
  assign n40513 = ~n40480 & ~n40512;
  assign n40514 = ~controllable_hgrant6 & ~n40513;
  assign n40515 = ~n40479 & ~n40514;
  assign n40516 = ~controllable_hmaster0 & ~n40515;
  assign n40517 = ~controllable_hmaster0 & ~n40516;
  assign n40518 = i_hlock8 & ~n40517;
  assign n40519 = i_hbusreq6 & ~n40448;
  assign n40520 = n8217 & ~n8777;
  assign n40521 = ~n8217 & ~n16877;
  assign n40522 = ~n40520 & ~n40521;
  assign n40523 = ~i_hbusreq6 & ~n40522;
  assign n40524 = ~n40519 & ~n40523;
  assign n40525 = controllable_hgrant6 & ~n40524;
  assign n40526 = i_hbusreq6 & ~n40462;
  assign n40527 = i_hbusreq5 & ~n40452;
  assign n40528 = n8378 & ~n8771;
  assign n40529 = ~n8378 & ~n16869;
  assign n40530 = ~n40528 & ~n40529;
  assign n40531 = ~i_hbusreq5 & ~n40530;
  assign n40532 = ~n40527 & ~n40531;
  assign n40533 = controllable_hgrant5 & ~n40532;
  assign n40534 = i_hbusreq5 & ~n40456;
  assign n40535 = i_hbusreq4 & ~n40203;
  assign n40536 = i_hbusreq9 & ~n40203;
  assign n40537 = ~i_hbusreq9 & ~n40292;
  assign n40538 = ~n40536 & ~n40537;
  assign n40539 = ~i_hbusreq4 & ~n40538;
  assign n40540 = ~n40535 & ~n40539;
  assign n40541 = controllable_hgrant4 & ~n40540;
  assign n40542 = i_hbusreq4 & ~n40249;
  assign n40543 = i_hbusreq9 & ~n40249;
  assign n40544 = ~i_hbusreq9 & ~n40394;
  assign n40545 = ~n40543 & ~n40544;
  assign n40546 = ~i_hbusreq4 & ~n40545;
  assign n40547 = ~n40542 & ~n40546;
  assign n40548 = ~controllable_hgrant4 & ~n40547;
  assign n40549 = ~n40541 & ~n40548;
  assign n40550 = ~i_hbusreq5 & ~n40549;
  assign n40551 = ~n40534 & ~n40550;
  assign n40552 = ~controllable_hgrant5 & ~n40551;
  assign n40553 = ~n40533 & ~n40552;
  assign n40554 = ~controllable_hmaster2 & ~n40553;
  assign n40555 = ~controllable_hmaster2 & ~n40554;
  assign n40556 = ~controllable_hmaster1 & ~n40555;
  assign n40557 = ~controllable_hmaster1 & ~n40556;
  assign n40558 = ~i_hbusreq6 & ~n40557;
  assign n40559 = ~n40526 & ~n40558;
  assign n40560 = ~controllable_hgrant6 & ~n40559;
  assign n40561 = ~n40525 & ~n40560;
  assign n40562 = ~controllable_hmaster0 & ~n40561;
  assign n40563 = ~controllable_hmaster0 & ~n40562;
  assign n40564 = ~i_hlock8 & ~n40563;
  assign n40565 = ~n40518 & ~n40564;
  assign n40566 = ~i_hbusreq8 & ~n40565;
  assign n40567 = ~n40472 & ~n40566;
  assign n40568 = controllable_hmaster3 & ~n40567;
  assign n40569 = controllable_hmaster3 & ~n40568;
  assign n40570 = ~i_hbusreq7 & ~n40569;
  assign n40571 = ~n40471 & ~n40570;
  assign n40572 = n8214 & ~n40571;
  assign n40573 = ~n40423 & ~n40572;
  assign n40574 = ~n8202 & ~n40573;
  assign n40575 = n8217 & ~n8796;
  assign n40576 = ~n8217 & ~n16899;
  assign n40577 = ~n40575 & ~n40576;
  assign n40578 = controllable_hgrant6 & ~n40577;
  assign n40579 = controllable_hmaster2 & ~n40436;
  assign n40580 = controllable_hmaster2 & ~n40579;
  assign n40581 = controllable_hmaster1 & ~n40580;
  assign n40582 = controllable_hmaster1 & ~n40581;
  assign n40583 = ~controllable_hgrant6 & ~n40582;
  assign n40584 = ~n40578 & ~n40583;
  assign n40585 = controllable_hmaster0 & ~n40584;
  assign n40586 = controllable_hmaster0 & ~n40585;
  assign n40587 = ~controllable_hmaster3 & ~n40586;
  assign n40588 = ~controllable_hmaster3 & ~n40587;
  assign n40589 = i_hlock7 & ~n40588;
  assign n40590 = n8217 & ~n8805;
  assign n40591 = ~n8217 & ~n16911;
  assign n40592 = ~n40590 & ~n40591;
  assign n40593 = controllable_hgrant6 & ~n40592;
  assign n40594 = controllable_hmaster2 & ~n40458;
  assign n40595 = controllable_hmaster2 & ~n40594;
  assign n40596 = controllable_hmaster1 & ~n40595;
  assign n40597 = controllable_hmaster1 & ~n40596;
  assign n40598 = ~controllable_hgrant6 & ~n40597;
  assign n40599 = ~n40593 & ~n40598;
  assign n40600 = controllable_hmaster0 & ~n40599;
  assign n40601 = controllable_hmaster0 & ~n40600;
  assign n40602 = ~controllable_hmaster3 & ~n40601;
  assign n40603 = ~controllable_hmaster3 & ~n40602;
  assign n40604 = ~i_hlock7 & ~n40603;
  assign n40605 = ~n40589 & ~n40604;
  assign n40606 = i_hbusreq7 & ~n40605;
  assign n40607 = i_hbusreq8 & ~n40586;
  assign n40608 = i_hbusreq6 & ~n40577;
  assign n40609 = n8217 & ~n8818;
  assign n40610 = ~n8217 & ~n16927;
  assign n40611 = ~n40609 & ~n40610;
  assign n40612 = ~i_hbusreq6 & ~n40611;
  assign n40613 = ~n40608 & ~n40612;
  assign n40614 = controllable_hgrant6 & ~n40613;
  assign n40615 = i_hbusreq6 & ~n40582;
  assign n40616 = controllable_hmaster2 & ~n40507;
  assign n40617 = controllable_hmaster2 & ~n40616;
  assign n40618 = controllable_hmaster1 & ~n40617;
  assign n40619 = controllable_hmaster1 & ~n40618;
  assign n40620 = ~i_hbusreq6 & ~n40619;
  assign n40621 = ~n40615 & ~n40620;
  assign n40622 = ~controllable_hgrant6 & ~n40621;
  assign n40623 = ~n40614 & ~n40622;
  assign n40624 = controllable_hmaster0 & ~n40623;
  assign n40625 = controllable_hmaster0 & ~n40624;
  assign n40626 = ~i_hbusreq8 & ~n40625;
  assign n40627 = ~n40607 & ~n40626;
  assign n40628 = ~controllable_hmaster3 & ~n40627;
  assign n40629 = ~controllable_hmaster3 & ~n40628;
  assign n40630 = i_hlock7 & ~n40629;
  assign n40631 = i_hbusreq8 & ~n40601;
  assign n40632 = i_hbusreq6 & ~n40592;
  assign n40633 = n8217 & ~n8833;
  assign n40634 = ~n8217 & ~n16945;
  assign n40635 = ~n40633 & ~n40634;
  assign n40636 = ~i_hbusreq6 & ~n40635;
  assign n40637 = ~n40632 & ~n40636;
  assign n40638 = controllable_hgrant6 & ~n40637;
  assign n40639 = i_hbusreq6 & ~n40597;
  assign n40640 = controllable_hmaster2 & ~n40553;
  assign n40641 = controllable_hmaster2 & ~n40640;
  assign n40642 = controllable_hmaster1 & ~n40641;
  assign n40643 = controllable_hmaster1 & ~n40642;
  assign n40644 = ~i_hbusreq6 & ~n40643;
  assign n40645 = ~n40639 & ~n40644;
  assign n40646 = ~controllable_hgrant6 & ~n40645;
  assign n40647 = ~n40638 & ~n40646;
  assign n40648 = controllable_hmaster0 & ~n40647;
  assign n40649 = controllable_hmaster0 & ~n40648;
  assign n40650 = ~i_hbusreq8 & ~n40649;
  assign n40651 = ~n40631 & ~n40650;
  assign n40652 = ~controllable_hmaster3 & ~n40651;
  assign n40653 = ~controllable_hmaster3 & ~n40652;
  assign n40654 = ~i_hlock7 & ~n40653;
  assign n40655 = ~n40630 & ~n40654;
  assign n40656 = ~i_hbusreq7 & ~n40655;
  assign n40657 = ~n40606 & ~n40656;
  assign n40658 = ~n8214 & ~n40657;
  assign n40659 = n8217 & ~n26644;
  assign n40660 = ~n8217 & ~n28873;
  assign n40661 = ~n40659 & ~n40660;
  assign n40662 = i_hlock6 & ~n40661;
  assign n40663 = n8217 & ~n26659;
  assign n40664 = ~n8217 & ~n28888;
  assign n40665 = ~n40663 & ~n40664;
  assign n40666 = ~i_hlock6 & ~n40665;
  assign n40667 = ~n40662 & ~n40666;
  assign n40668 = controllable_hgrant6 & ~n40667;
  assign n40669 = i_hlock6 & ~n40582;
  assign n40670 = ~i_hlock6 & ~n40597;
  assign n40671 = ~n40669 & ~n40670;
  assign n40672 = ~controllable_hgrant6 & ~n40671;
  assign n40673 = ~n40668 & ~n40672;
  assign n40674 = ~controllable_hmaster0 & ~n40673;
  assign n40675 = ~controllable_hmaster0 & ~n40674;
  assign n40676 = ~controllable_hmaster3 & ~n40675;
  assign n40677 = ~controllable_hmaster3 & ~n40676;
  assign n40678 = i_hbusreq7 & ~n40677;
  assign n40679 = i_hbusreq8 & ~n40675;
  assign n40680 = i_hbusreq6 & ~n40667;
  assign n40681 = n8217 & ~n26687;
  assign n40682 = ~n8217 & ~n28916;
  assign n40683 = ~n40681 & ~n40682;
  assign n40684 = i_hlock6 & ~n40683;
  assign n40685 = n8217 & ~n26717;
  assign n40686 = ~n8217 & ~n28946;
  assign n40687 = ~n40685 & ~n40686;
  assign n40688 = ~i_hlock6 & ~n40687;
  assign n40689 = ~n40684 & ~n40688;
  assign n40690 = ~i_hbusreq6 & ~n40689;
  assign n40691 = ~n40680 & ~n40690;
  assign n40692 = controllable_hgrant6 & ~n40691;
  assign n40693 = i_hbusreq6 & ~n40671;
  assign n40694 = i_hlock6 & ~n40619;
  assign n40695 = ~i_hlock6 & ~n40643;
  assign n40696 = ~n40694 & ~n40695;
  assign n40697 = ~i_hbusreq6 & ~n40696;
  assign n40698 = ~n40693 & ~n40697;
  assign n40699 = ~controllable_hgrant6 & ~n40698;
  assign n40700 = ~n40692 & ~n40699;
  assign n40701 = ~controllable_hmaster0 & ~n40700;
  assign n40702 = ~controllable_hmaster0 & ~n40701;
  assign n40703 = ~i_hbusreq8 & ~n40702;
  assign n40704 = ~n40679 & ~n40703;
  assign n40705 = ~controllable_hmaster3 & ~n40704;
  assign n40706 = ~controllable_hmaster3 & ~n40705;
  assign n40707 = ~i_hbusreq7 & ~n40706;
  assign n40708 = ~n40678 & ~n40707;
  assign n40709 = ~n7924 & ~n40708;
  assign n40710 = n8217 & ~n12796;
  assign n40711 = ~n8217 & ~n28965;
  assign n40712 = ~n40710 & ~n40711;
  assign n40713 = i_hlock6 & ~n40712;
  assign n40714 = ~n8217 & ~n28990;
  assign n40715 = ~n40710 & ~n40714;
  assign n40716 = ~i_hlock6 & ~n40715;
  assign n40717 = ~n40713 & ~n40716;
  assign n40718 = controllable_hgrant6 & ~n40717;
  assign n40719 = controllable_hgrant6 & ~n40718;
  assign n40720 = controllable_hmaster3 & ~n40719;
  assign n40721 = controllable_hmaster0 & ~n40719;
  assign n40722 = n8217 & ~n26742;
  assign n40723 = ~n8217 & ~n28978;
  assign n40724 = ~n40722 & ~n40723;
  assign n40725 = i_hlock6 & ~n40724;
  assign n40726 = n8217 & ~n26757;
  assign n40727 = ~n8217 & ~n29003;
  assign n40728 = ~n40726 & ~n40727;
  assign n40729 = ~i_hlock6 & ~n40728;
  assign n40730 = ~n40725 & ~n40729;
  assign n40731 = controllable_hgrant6 & ~n40730;
  assign n40732 = ~n40672 & ~n40731;
  assign n40733 = ~controllable_hmaster0 & ~n40732;
  assign n40734 = ~n40721 & ~n40733;
  assign n40735 = ~controllable_hmaster3 & ~n40734;
  assign n40736 = ~n40720 & ~n40735;
  assign n40737 = i_hbusreq7 & ~n40736;
  assign n40738 = i_hbusreq8 & ~n40719;
  assign n40739 = i_hbusreq6 & ~n40717;
  assign n40740 = n8217 & ~n12875;
  assign n40741 = ~n8217 & ~n29028;
  assign n40742 = ~n40740 & ~n40741;
  assign n40743 = i_hlock6 & ~n40742;
  assign n40744 = ~n8217 & ~n29083;
  assign n40745 = ~n40740 & ~n40744;
  assign n40746 = ~i_hlock6 & ~n40745;
  assign n40747 = ~n40743 & ~n40746;
  assign n40748 = ~i_hbusreq6 & ~n40747;
  assign n40749 = ~n40739 & ~n40748;
  assign n40750 = controllable_hgrant6 & ~n40749;
  assign n40751 = controllable_hgrant6 & ~n40750;
  assign n40752 = ~i_hbusreq8 & ~n40751;
  assign n40753 = ~n40738 & ~n40752;
  assign n40754 = controllable_hmaster3 & ~n40753;
  assign n40755 = i_hbusreq8 & ~n40734;
  assign n40756 = controllable_hmaster0 & ~n40751;
  assign n40757 = i_hbusreq6 & ~n40730;
  assign n40758 = n8217 & ~n26787;
  assign n40759 = ~n8217 & ~n29056;
  assign n40760 = ~n40758 & ~n40759;
  assign n40761 = i_hlock6 & ~n40760;
  assign n40762 = n8217 & ~n26817;
  assign n40763 = ~n8217 & ~n29111;
  assign n40764 = ~n40762 & ~n40763;
  assign n40765 = ~i_hlock6 & ~n40764;
  assign n40766 = ~n40761 & ~n40765;
  assign n40767 = ~i_hbusreq6 & ~n40766;
  assign n40768 = ~n40757 & ~n40767;
  assign n40769 = controllable_hgrant6 & ~n40768;
  assign n40770 = ~n40699 & ~n40769;
  assign n40771 = ~controllable_hmaster0 & ~n40770;
  assign n40772 = ~n40756 & ~n40771;
  assign n40773 = ~i_hbusreq8 & ~n40772;
  assign n40774 = ~n40755 & ~n40773;
  assign n40775 = ~controllable_hmaster3 & ~n40774;
  assign n40776 = ~n40754 & ~n40775;
  assign n40777 = ~i_hbusreq7 & ~n40776;
  assign n40778 = ~n40737 & ~n40777;
  assign n40779 = n7924 & ~n40778;
  assign n40780 = ~n40709 & ~n40779;
  assign n40781 = n8214 & ~n40780;
  assign n40782 = ~n40658 & ~n40781;
  assign n40783 = n8202 & ~n40782;
  assign n40784 = ~n40574 & ~n40783;
  assign n40785 = n7920 & ~n40784;
  assign n40786 = ~n40188 & ~n40785;
  assign n40787 = n7728 & ~n40786;
  assign n40788 = ~n7920 & ~n39742;
  assign n40789 = n8217 & ~n8880;
  assign n40790 = ~n8217 & ~n29139;
  assign n40791 = ~n40789 & ~n40790;
  assign n40792 = controllable_hgrant6 & ~n40791;
  assign n40793 = ~n7951 & ~n40256;
  assign n40794 = ~controllable_hmaster1 & ~n40793;
  assign n40795 = ~n7950 & ~n40794;
  assign n40796 = ~controllable_hgrant6 & ~n40795;
  assign n40797 = ~n40792 & ~n40796;
  assign n40798 = controllable_hmaster0 & ~n40797;
  assign n40799 = ~controllable_hmaster0 & ~n7956;
  assign n40800 = ~n40798 & ~n40799;
  assign n40801 = controllable_hmaster3 & ~n40800;
  assign n40802 = controllable_hmaster3 & ~n40801;
  assign n40803 = i_hbusreq7 & ~n40802;
  assign n40804 = i_hbusreq8 & ~n40800;
  assign n40805 = i_hbusreq6 & ~n40791;
  assign n40806 = n8217 & ~n8891;
  assign n40807 = ~n8217 & ~n29151;
  assign n40808 = ~n40806 & ~n40807;
  assign n40809 = ~i_hbusreq6 & ~n40808;
  assign n40810 = ~n40805 & ~n40809;
  assign n40811 = controllable_hgrant6 & ~n40810;
  assign n40812 = i_hbusreq6 & ~n40795;
  assign n40813 = ~n8008 & ~n40407;
  assign n40814 = ~controllable_hmaster1 & ~n40813;
  assign n40815 = ~n8007 & ~n40814;
  assign n40816 = ~i_hbusreq6 & ~n40815;
  assign n40817 = ~n40812 & ~n40816;
  assign n40818 = ~controllable_hgrant6 & ~n40817;
  assign n40819 = ~n40811 & ~n40818;
  assign n40820 = controllable_hmaster0 & ~n40819;
  assign n40821 = ~controllable_hmaster0 & ~n8015;
  assign n40822 = ~n40820 & ~n40821;
  assign n40823 = ~i_hbusreq8 & ~n40822;
  assign n40824 = ~n40804 & ~n40823;
  assign n40825 = controllable_hmaster3 & ~n40824;
  assign n40826 = controllable_hmaster3 & ~n40825;
  assign n40827 = ~i_hbusreq7 & ~n40826;
  assign n40828 = ~n40803 & ~n40827;
  assign n40829 = ~n7924 & ~n40828;
  assign n40830 = ~n7733 & n40219;
  assign n40831 = ~n40228 & ~n40830;
  assign n40832 = n7928 & ~n40831;
  assign n40833 = ~n8221 & ~n40832;
  assign n40834 = ~controllable_hgrant1 & ~n40833;
  assign n40835 = ~n40214 & ~n40834;
  assign n40836 = ~controllable_hgrant3 & ~n40835;
  assign n40837 = ~n40210 & ~n40836;
  assign n40838 = i_hlock9 & ~n40837;
  assign n40839 = ~n8235 & ~n40832;
  assign n40840 = ~controllable_hgrant1 & ~n40839;
  assign n40841 = ~n40244 & ~n40840;
  assign n40842 = ~controllable_hgrant3 & ~n40841;
  assign n40843 = ~n40240 & ~n40842;
  assign n40844 = ~i_hlock9 & ~n40843;
  assign n40845 = ~n40838 & ~n40844;
  assign n40846 = ~controllable_hgrant4 & ~n40845;
  assign n40847 = ~n40206 & ~n40846;
  assign n40848 = ~controllable_hgrant5 & ~n40847;
  assign n40849 = ~n40196 & ~n40848;
  assign n40850 = ~controllable_hmaster2 & ~n40849;
  assign n40851 = ~n8036 & ~n40850;
  assign n40852 = ~controllable_hmaster1 & ~n40851;
  assign n40853 = ~n8035 & ~n40852;
  assign n40854 = ~controllable_hgrant6 & ~n40853;
  assign n40855 = ~n40792 & ~n40854;
  assign n40856 = controllable_hmaster0 & ~n40855;
  assign n40857 = ~controllable_hmaster0 & ~n8056;
  assign n40858 = ~n40856 & ~n40857;
  assign n40859 = controllable_hmaster3 & ~n40858;
  assign n40860 = ~n8060 & ~n40859;
  assign n40861 = i_hbusreq7 & ~n40860;
  assign n40862 = i_hbusreq8 & ~n40858;
  assign n40863 = i_hbusreq6 & ~n40853;
  assign n40864 = i_hbusreq5 & ~n40847;
  assign n40865 = i_hbusreq4 & ~n40845;
  assign n40866 = i_hbusreq9 & ~n40845;
  assign n40867 = i_hbusreq3 & ~n40835;
  assign n40868 = i_hbusreq1 & ~n40833;
  assign n40869 = i_hlock0 & controllable_ndecide;
  assign n40870 = ~i_hlock0 & ~n12782;
  assign n40871 = ~n40869 & ~n40870;
  assign n40872 = ~i_hbusreq0 & ~n40871;
  assign n40873 = ~i_hbusreq0 & ~n40872;
  assign n40874 = ~i_hbusreq2 & ~n40873;
  assign n40875 = ~i_hbusreq2 & ~n40874;
  assign n40876 = ~controllable_hgrant2 & n40875;
  assign n40877 = ~n40330 & ~n40876;
  assign n40878 = ~n7733 & ~n40877;
  assign n40879 = ~n40357 & ~n40878;
  assign n40880 = n7928 & ~n40879;
  assign n40881 = ~n8265 & ~n40880;
  assign n40882 = ~i_hbusreq1 & ~n40881;
  assign n40883 = ~n40868 & ~n40882;
  assign n40884 = ~controllable_hgrant1 & ~n40883;
  assign n40885 = ~n40316 & ~n40884;
  assign n40886 = ~i_hbusreq3 & ~n40885;
  assign n40887 = ~n40867 & ~n40886;
  assign n40888 = ~controllable_hgrant3 & ~n40887;
  assign n40889 = ~n40308 & ~n40888;
  assign n40890 = i_hlock9 & ~n40889;
  assign n40891 = i_hbusreq3 & ~n40841;
  assign n40892 = i_hbusreq1 & ~n40839;
  assign n40893 = ~n8297 & ~n40880;
  assign n40894 = ~i_hbusreq1 & ~n40893;
  assign n40895 = ~n40892 & ~n40894;
  assign n40896 = ~controllable_hgrant1 & ~n40895;
  assign n40897 = ~n40384 & ~n40896;
  assign n40898 = ~i_hbusreq3 & ~n40897;
  assign n40899 = ~n40891 & ~n40898;
  assign n40900 = ~controllable_hgrant3 & ~n40899;
  assign n40901 = ~n40376 & ~n40900;
  assign n40902 = ~i_hlock9 & ~n40901;
  assign n40903 = ~n40890 & ~n40902;
  assign n40904 = ~i_hbusreq9 & ~n40903;
  assign n40905 = ~n40866 & ~n40904;
  assign n40906 = ~i_hbusreq4 & ~n40905;
  assign n40907 = ~n40865 & ~n40906;
  assign n40908 = ~controllable_hgrant4 & ~n40907;
  assign n40909 = ~n40299 & ~n40908;
  assign n40910 = ~i_hbusreq5 & ~n40909;
  assign n40911 = ~n40864 & ~n40910;
  assign n40912 = ~controllable_hgrant5 & ~n40911;
  assign n40913 = ~n40282 & ~n40912;
  assign n40914 = ~controllable_hmaster2 & ~n40913;
  assign n40915 = ~n8099 & ~n40914;
  assign n40916 = ~controllable_hmaster1 & ~n40915;
  assign n40917 = ~n8098 & ~n40916;
  assign n40918 = ~i_hbusreq6 & ~n40917;
  assign n40919 = ~n40863 & ~n40918;
  assign n40920 = ~controllable_hgrant6 & ~n40919;
  assign n40921 = ~n40811 & ~n40920;
  assign n40922 = controllable_hmaster0 & ~n40921;
  assign n40923 = ~controllable_hmaster0 & ~n8142;
  assign n40924 = ~n40922 & ~n40923;
  assign n40925 = ~i_hbusreq8 & ~n40924;
  assign n40926 = ~n40862 & ~n40925;
  assign n40927 = controllable_hmaster3 & ~n40926;
  assign n40928 = ~n8154 & ~n40927;
  assign n40929 = ~i_hbusreq7 & ~n40928;
  assign n40930 = ~n40861 & ~n40929;
  assign n40931 = n7924 & ~n40930;
  assign n40932 = ~n40829 & ~n40931;
  assign n40933 = ~n8214 & ~n40932;
  assign n40934 = controllable_hmaster0 & ~n7956;
  assign n40935 = n8217 & ~n8907;
  assign n40936 = ~n8217 & ~n17228;
  assign n40937 = ~n40935 & ~n40936;
  assign n40938 = controllable_hgrant6 & ~n40937;
  assign n40939 = ~n7951 & ~n40437;
  assign n40940 = ~controllable_hmaster1 & ~n40939;
  assign n40941 = ~n7950 & ~n40940;
  assign n40942 = ~controllable_hgrant6 & ~n40941;
  assign n40943 = ~n40938 & ~n40942;
  assign n40944 = ~controllable_hmaster0 & ~n40943;
  assign n40945 = ~n40934 & ~n40944;
  assign n40946 = i_hlock8 & ~n40945;
  assign n40947 = n8217 & ~n8913;
  assign n40948 = ~n8217 & ~n17237;
  assign n40949 = ~n40947 & ~n40948;
  assign n40950 = controllable_hgrant6 & ~n40949;
  assign n40951 = ~n7951 & ~n40459;
  assign n40952 = ~controllable_hmaster1 & ~n40951;
  assign n40953 = ~n7950 & ~n40952;
  assign n40954 = ~controllable_hgrant6 & ~n40953;
  assign n40955 = ~n40950 & ~n40954;
  assign n40956 = ~controllable_hmaster0 & ~n40955;
  assign n40957 = ~n40934 & ~n40956;
  assign n40958 = ~i_hlock8 & ~n40957;
  assign n40959 = ~n40946 & ~n40958;
  assign n40960 = controllable_hmaster3 & ~n40959;
  assign n40961 = controllable_hmaster3 & ~n40960;
  assign n40962 = i_hbusreq7 & ~n40961;
  assign n40963 = i_hbusreq8 & ~n40959;
  assign n40964 = controllable_hmaster0 & ~n8015;
  assign n40965 = i_hbusreq6 & ~n40937;
  assign n40966 = n8217 & ~n8926;
  assign n40967 = ~n8217 & ~n17252;
  assign n40968 = ~n40966 & ~n40967;
  assign n40969 = ~i_hbusreq6 & ~n40968;
  assign n40970 = ~n40965 & ~n40969;
  assign n40971 = controllable_hgrant6 & ~n40970;
  assign n40972 = i_hbusreq6 & ~n40941;
  assign n40973 = ~n8008 & ~n40508;
  assign n40974 = ~controllable_hmaster1 & ~n40973;
  assign n40975 = ~n8007 & ~n40974;
  assign n40976 = ~i_hbusreq6 & ~n40975;
  assign n40977 = ~n40972 & ~n40976;
  assign n40978 = ~controllable_hgrant6 & ~n40977;
  assign n40979 = ~n40971 & ~n40978;
  assign n40980 = ~controllable_hmaster0 & ~n40979;
  assign n40981 = ~n40964 & ~n40980;
  assign n40982 = i_hlock8 & ~n40981;
  assign n40983 = i_hbusreq6 & ~n40949;
  assign n40984 = n8217 & ~n8935;
  assign n40985 = ~n8217 & ~n17264;
  assign n40986 = ~n40984 & ~n40985;
  assign n40987 = ~i_hbusreq6 & ~n40986;
  assign n40988 = ~n40983 & ~n40987;
  assign n40989 = controllable_hgrant6 & ~n40988;
  assign n40990 = i_hbusreq6 & ~n40953;
  assign n40991 = ~n8008 & ~n40554;
  assign n40992 = ~controllable_hmaster1 & ~n40991;
  assign n40993 = ~n8007 & ~n40992;
  assign n40994 = ~i_hbusreq6 & ~n40993;
  assign n40995 = ~n40990 & ~n40994;
  assign n40996 = ~controllable_hgrant6 & ~n40995;
  assign n40997 = ~n40989 & ~n40996;
  assign n40998 = ~controllable_hmaster0 & ~n40997;
  assign n40999 = ~n40964 & ~n40998;
  assign n41000 = ~i_hlock8 & ~n40999;
  assign n41001 = ~n40982 & ~n41000;
  assign n41002 = ~i_hbusreq8 & ~n41001;
  assign n41003 = ~n40963 & ~n41002;
  assign n41004 = controllable_hmaster3 & ~n41003;
  assign n41005 = controllable_hmaster3 & ~n41004;
  assign n41006 = ~i_hbusreq7 & ~n41005;
  assign n41007 = ~n40962 & ~n41006;
  assign n41008 = ~n7924 & ~n41007;
  assign n41009 = controllable_hmaster0 & ~n8056;
  assign n41010 = ~controllable_hgrant4 & ~n40837;
  assign n41011 = ~n40432 & ~n41010;
  assign n41012 = ~controllable_hgrant5 & ~n41011;
  assign n41013 = ~n40431 & ~n41012;
  assign n41014 = ~controllable_hmaster2 & ~n41013;
  assign n41015 = ~n8036 & ~n41014;
  assign n41016 = ~controllable_hmaster1 & ~n41015;
  assign n41017 = ~n8035 & ~n41016;
  assign n41018 = ~controllable_hgrant6 & ~n41017;
  assign n41019 = ~n40938 & ~n41018;
  assign n41020 = ~controllable_hmaster0 & ~n41019;
  assign n41021 = ~n41009 & ~n41020;
  assign n41022 = i_hlock8 & ~n41021;
  assign n41023 = ~controllable_hgrant4 & ~n40843;
  assign n41024 = ~n40454 & ~n41023;
  assign n41025 = ~controllable_hgrant5 & ~n41024;
  assign n41026 = ~n40453 & ~n41025;
  assign n41027 = ~controllable_hmaster2 & ~n41026;
  assign n41028 = ~n8036 & ~n41027;
  assign n41029 = ~controllable_hmaster1 & ~n41028;
  assign n41030 = ~n8035 & ~n41029;
  assign n41031 = ~controllable_hgrant6 & ~n41030;
  assign n41032 = ~n40950 & ~n41031;
  assign n41033 = ~controllable_hmaster0 & ~n41032;
  assign n41034 = ~n41009 & ~n41033;
  assign n41035 = ~i_hlock8 & ~n41034;
  assign n41036 = ~n41022 & ~n41035;
  assign n41037 = controllable_hmaster3 & ~n41036;
  assign n41038 = ~n8060 & ~n41037;
  assign n41039 = i_hbusreq7 & ~n41038;
  assign n41040 = i_hbusreq8 & ~n41036;
  assign n41041 = controllable_hmaster0 & ~n8142;
  assign n41042 = i_hbusreq6 & ~n41017;
  assign n41043 = i_hbusreq5 & ~n41011;
  assign n41044 = i_hbusreq4 & ~n40837;
  assign n41045 = i_hbusreq9 & ~n40837;
  assign n41046 = ~i_hbusreq9 & ~n40889;
  assign n41047 = ~n41045 & ~n41046;
  assign n41048 = ~i_hbusreq4 & ~n41047;
  assign n41049 = ~n41044 & ~n41048;
  assign n41050 = ~controllable_hgrant4 & ~n41049;
  assign n41051 = ~n40495 & ~n41050;
  assign n41052 = ~i_hbusreq5 & ~n41051;
  assign n41053 = ~n41043 & ~n41052;
  assign n41054 = ~controllable_hgrant5 & ~n41053;
  assign n41055 = ~n40487 & ~n41054;
  assign n41056 = ~controllable_hmaster2 & ~n41055;
  assign n41057 = ~n8099 & ~n41056;
  assign n41058 = ~controllable_hmaster1 & ~n41057;
  assign n41059 = ~n8098 & ~n41058;
  assign n41060 = ~i_hbusreq6 & ~n41059;
  assign n41061 = ~n41042 & ~n41060;
  assign n41062 = ~controllable_hgrant6 & ~n41061;
  assign n41063 = ~n40971 & ~n41062;
  assign n41064 = ~controllable_hmaster0 & ~n41063;
  assign n41065 = ~n41041 & ~n41064;
  assign n41066 = i_hlock8 & ~n41065;
  assign n41067 = i_hbusreq6 & ~n41030;
  assign n41068 = i_hbusreq5 & ~n41024;
  assign n41069 = i_hbusreq4 & ~n40843;
  assign n41070 = i_hbusreq9 & ~n40843;
  assign n41071 = ~i_hbusreq9 & ~n40901;
  assign n41072 = ~n41070 & ~n41071;
  assign n41073 = ~i_hbusreq4 & ~n41072;
  assign n41074 = ~n41069 & ~n41073;
  assign n41075 = ~controllable_hgrant4 & ~n41074;
  assign n41076 = ~n40541 & ~n41075;
  assign n41077 = ~i_hbusreq5 & ~n41076;
  assign n41078 = ~n41068 & ~n41077;
  assign n41079 = ~controllable_hgrant5 & ~n41078;
  assign n41080 = ~n40533 & ~n41079;
  assign n41081 = ~controllable_hmaster2 & ~n41080;
  assign n41082 = ~n8099 & ~n41081;
  assign n41083 = ~controllable_hmaster1 & ~n41082;
  assign n41084 = ~n8098 & ~n41083;
  assign n41085 = ~i_hbusreq6 & ~n41084;
  assign n41086 = ~n41067 & ~n41085;
  assign n41087 = ~controllable_hgrant6 & ~n41086;
  assign n41088 = ~n40989 & ~n41087;
  assign n41089 = ~controllable_hmaster0 & ~n41088;
  assign n41090 = ~n41041 & ~n41089;
  assign n41091 = ~i_hlock8 & ~n41090;
  assign n41092 = ~n41066 & ~n41091;
  assign n41093 = ~i_hbusreq8 & ~n41092;
  assign n41094 = ~n41040 & ~n41093;
  assign n41095 = controllable_hmaster3 & ~n41094;
  assign n41096 = ~n8154 & ~n41095;
  assign n41097 = ~i_hbusreq7 & ~n41096;
  assign n41098 = ~n41039 & ~n41097;
  assign n41099 = n7924 & ~n41098;
  assign n41100 = ~n41008 & ~n41099;
  assign n41101 = n8214 & ~n41100;
  assign n41102 = ~n40933 & ~n41101;
  assign n41103 = ~n8202 & ~n41102;
  assign n41104 = ~n7957 & ~n40587;
  assign n41105 = i_hlock7 & ~n41104;
  assign n41106 = ~n7957 & ~n40602;
  assign n41107 = ~i_hlock7 & ~n41106;
  assign n41108 = ~n41105 & ~n41107;
  assign n41109 = i_hbusreq7 & ~n41108;
  assign n41110 = ~n8018 & ~n40628;
  assign n41111 = i_hlock7 & ~n41110;
  assign n41112 = ~n8018 & ~n40652;
  assign n41113 = ~i_hlock7 & ~n41112;
  assign n41114 = ~n41111 & ~n41113;
  assign n41115 = ~i_hbusreq7 & ~n41114;
  assign n41116 = ~n41109 & ~n41115;
  assign n41117 = ~n7924 & ~n41116;
  assign n41118 = controllable_hmaster2 & ~n41013;
  assign n41119 = ~n8051 & ~n41118;
  assign n41120 = controllable_hmaster1 & ~n41119;
  assign n41121 = ~controllable_hmaster1 & ~n8050;
  assign n41122 = ~n41120 & ~n41121;
  assign n41123 = ~controllable_hgrant6 & ~n41122;
  assign n41124 = ~n40578 & ~n41123;
  assign n41125 = controllable_hmaster0 & ~n41124;
  assign n41126 = ~controllable_hmaster0 & ~n8059;
  assign n41127 = ~n41125 & ~n41126;
  assign n41128 = ~controllable_hmaster3 & ~n41127;
  assign n41129 = ~n8057 & ~n41128;
  assign n41130 = i_hlock7 & ~n41129;
  assign n41131 = controllable_hmaster2 & ~n41026;
  assign n41132 = ~n8051 & ~n41131;
  assign n41133 = controllable_hmaster1 & ~n41132;
  assign n41134 = ~n41121 & ~n41133;
  assign n41135 = ~controllable_hgrant6 & ~n41134;
  assign n41136 = ~n40593 & ~n41135;
  assign n41137 = controllable_hmaster0 & ~n41136;
  assign n41138 = ~n41126 & ~n41137;
  assign n41139 = ~controllable_hmaster3 & ~n41138;
  assign n41140 = ~n8057 & ~n41139;
  assign n41141 = ~i_hlock7 & ~n41140;
  assign n41142 = ~n41130 & ~n41141;
  assign n41143 = i_hbusreq7 & ~n41142;
  assign n41144 = i_hbusreq8 & ~n41127;
  assign n41145 = i_hbusreq6 & ~n41122;
  assign n41146 = controllable_hmaster2 & ~n41055;
  assign n41147 = ~n8135 & ~n41146;
  assign n41148 = controllable_hmaster1 & ~n41147;
  assign n41149 = ~controllable_hmaster1 & ~n8134;
  assign n41150 = ~n41148 & ~n41149;
  assign n41151 = ~i_hbusreq6 & ~n41150;
  assign n41152 = ~n41145 & ~n41151;
  assign n41153 = ~controllable_hgrant6 & ~n41152;
  assign n41154 = ~n40614 & ~n41153;
  assign n41155 = controllable_hmaster0 & ~n41154;
  assign n41156 = ~controllable_hmaster0 & ~n8151;
  assign n41157 = ~n41155 & ~n41156;
  assign n41158 = ~i_hbusreq8 & ~n41157;
  assign n41159 = ~n41144 & ~n41158;
  assign n41160 = ~controllable_hmaster3 & ~n41159;
  assign n41161 = ~n8145 & ~n41160;
  assign n41162 = i_hlock7 & ~n41161;
  assign n41163 = i_hbusreq8 & ~n41138;
  assign n41164 = i_hbusreq6 & ~n41134;
  assign n41165 = controllable_hmaster2 & ~n41080;
  assign n41166 = ~n8135 & ~n41165;
  assign n41167 = controllable_hmaster1 & ~n41166;
  assign n41168 = ~n41149 & ~n41167;
  assign n41169 = ~i_hbusreq6 & ~n41168;
  assign n41170 = ~n41164 & ~n41169;
  assign n41171 = ~controllable_hgrant6 & ~n41170;
  assign n41172 = ~n40638 & ~n41171;
  assign n41173 = controllable_hmaster0 & ~n41172;
  assign n41174 = ~n41156 & ~n41173;
  assign n41175 = ~i_hbusreq8 & ~n41174;
  assign n41176 = ~n41163 & ~n41175;
  assign n41177 = ~controllable_hmaster3 & ~n41176;
  assign n41178 = ~n8145 & ~n41177;
  assign n41179 = ~i_hlock7 & ~n41178;
  assign n41180 = ~n41162 & ~n41179;
  assign n41181 = ~i_hbusreq7 & ~n41180;
  assign n41182 = ~n41143 & ~n41181;
  assign n41183 = n7924 & ~n41182;
  assign n41184 = ~n41117 & ~n41183;
  assign n41185 = ~n8214 & ~n41184;
  assign n41186 = ~n7742 & n8217;
  assign n41187 = ~n8217 & ~n17020;
  assign n41188 = ~n41186 & ~n41187;
  assign n41189 = controllable_hgrant6 & ~n41188;
  assign n41190 = ~n7955 & ~n41189;
  assign n41191 = controllable_hmaster3 & ~n41190;
  assign n41192 = ~n40676 & ~n41191;
  assign n41193 = i_hbusreq7 & ~n41192;
  assign n41194 = i_hbusreq8 & ~n41190;
  assign n41195 = i_hbusreq6 & ~n41188;
  assign n41196 = ~n7774 & n8217;
  assign n41197 = ~n8217 & ~n17074;
  assign n41198 = ~n41196 & ~n41197;
  assign n41199 = ~i_hbusreq6 & ~n41198;
  assign n41200 = ~n41195 & ~n41199;
  assign n41201 = controllable_hgrant6 & ~n41200;
  assign n41202 = ~n8014 & ~n41201;
  assign n41203 = ~i_hbusreq8 & ~n41202;
  assign n41204 = ~n41194 & ~n41203;
  assign n41205 = controllable_hmaster3 & ~n41204;
  assign n41206 = ~n40705 & ~n41205;
  assign n41207 = ~i_hbusreq7 & ~n41206;
  assign n41208 = ~n41193 & ~n41207;
  assign n41209 = ~n7924 & ~n41208;
  assign n41210 = n8217 & ~n13035;
  assign n41211 = ~n8217 & ~n29193;
  assign n41212 = ~n41210 & ~n41211;
  assign n41213 = i_hlock6 & ~n41212;
  assign n41214 = ~n8217 & ~n29207;
  assign n41215 = ~n41210 & ~n41214;
  assign n41216 = ~i_hlock6 & ~n41215;
  assign n41217 = ~n41213 & ~n41216;
  assign n41218 = controllable_hgrant6 & ~n41217;
  assign n41219 = ~n8055 & ~n41218;
  assign n41220 = controllable_hmaster3 & ~n41219;
  assign n41221 = ~n8058 & ~n40718;
  assign n41222 = controllable_hmaster0 & ~n41221;
  assign n41223 = i_hlock6 & ~n41122;
  assign n41224 = ~i_hlock6 & ~n41134;
  assign n41225 = ~n41223 & ~n41224;
  assign n41226 = ~controllable_hgrant6 & ~n41225;
  assign n41227 = ~n40731 & ~n41226;
  assign n41228 = ~controllable_hmaster0 & ~n41227;
  assign n41229 = ~n41222 & ~n41228;
  assign n41230 = ~controllable_hmaster3 & ~n41229;
  assign n41231 = ~n41220 & ~n41230;
  assign n41232 = i_hbusreq7 & ~n41231;
  assign n41233 = i_hbusreq8 & ~n41219;
  assign n41234 = i_hbusreq6 & ~n41217;
  assign n41235 = n8217 & ~n13094;
  assign n41236 = ~n8217 & ~n29234;
  assign n41237 = ~n41235 & ~n41236;
  assign n41238 = i_hlock6 & ~n41237;
  assign n41239 = ~n8217 & ~n29263;
  assign n41240 = ~n41235 & ~n41239;
  assign n41241 = ~i_hlock6 & ~n41240;
  assign n41242 = ~n41238 & ~n41241;
  assign n41243 = ~i_hbusreq6 & ~n41242;
  assign n41244 = ~n41234 & ~n41243;
  assign n41245 = controllable_hgrant6 & ~n41244;
  assign n41246 = ~n8141 & ~n41245;
  assign n41247 = ~i_hbusreq8 & ~n41246;
  assign n41248 = ~n41233 & ~n41247;
  assign n41249 = controllable_hmaster3 & ~n41248;
  assign n41250 = i_hbusreq8 & ~n41229;
  assign n41251 = ~n8150 & ~n40750;
  assign n41252 = controllable_hmaster0 & ~n41251;
  assign n41253 = i_hbusreq6 & ~n41225;
  assign n41254 = i_hlock6 & ~n41150;
  assign n41255 = ~i_hlock6 & ~n41168;
  assign n41256 = ~n41254 & ~n41255;
  assign n41257 = ~i_hbusreq6 & ~n41256;
  assign n41258 = ~n41253 & ~n41257;
  assign n41259 = ~controllable_hgrant6 & ~n41258;
  assign n41260 = ~n40769 & ~n41259;
  assign n41261 = ~controllable_hmaster0 & ~n41260;
  assign n41262 = ~n41252 & ~n41261;
  assign n41263 = ~i_hbusreq8 & ~n41262;
  assign n41264 = ~n41250 & ~n41263;
  assign n41265 = ~controllable_hmaster3 & ~n41264;
  assign n41266 = ~n41249 & ~n41265;
  assign n41267 = ~i_hbusreq7 & ~n41266;
  assign n41268 = ~n41232 & ~n41267;
  assign n41269 = n7924 & ~n41268;
  assign n41270 = ~n41209 & ~n41269;
  assign n41271 = n8214 & ~n41270;
  assign n41272 = ~n41185 & ~n41271;
  assign n41273 = n8202 & ~n41272;
  assign n41274 = ~n41103 & ~n41273;
  assign n41275 = n7920 & ~n41274;
  assign n41276 = ~n40788 & ~n41275;
  assign n41277 = ~n7728 & ~n41276;
  assign n41278 = ~n40787 & ~n41277;
  assign n41279 = ~n7723 & ~n41278;
  assign n41280 = ~n7723 & ~n41279;
  assign n41281 = ~n7714 & ~n41280;
  assign n41282 = ~n7714 & ~n41281;
  assign n41283 = n7705 & ~n41282;
  assign n41284 = n8217 & ~n8985;
  assign n41285 = ~n8217 & ~n29293;
  assign n41286 = ~n41284 & ~n41285;
  assign n41287 = controllable_hgrant6 & ~n41286;
  assign n41288 = n7733 & ~n12629;
  assign n41289 = ~n7823 & ~n41288;
  assign n41290 = ~n7928 & ~n41289;
  assign n41291 = ~n7938 & ~n41288;
  assign n41292 = n7928 & ~n41291;
  assign n41293 = ~n41290 & ~n41292;
  assign n41294 = ~controllable_hgrant1 & ~n41293;
  assign n41295 = ~n13155 & ~n41294;
  assign n41296 = ~controllable_hgrant3 & ~n41295;
  assign n41297 = ~n13154 & ~n41296;
  assign n41298 = ~controllable_hgrant4 & ~n41297;
  assign n41299 = ~n13153 & ~n41298;
  assign n41300 = ~controllable_hgrant5 & ~n41299;
  assign n41301 = ~n13152 & ~n41300;
  assign n41302 = controllable_hmaster1 & ~n41301;
  assign n41303 = controllable_hmaster2 & ~n41301;
  assign n41304 = ~n40256 & ~n41303;
  assign n41305 = ~controllable_hmaster1 & ~n41304;
  assign n41306 = ~n41302 & ~n41305;
  assign n41307 = ~controllable_hgrant6 & ~n41306;
  assign n41308 = ~n41287 & ~n41307;
  assign n41309 = controllable_hmaster0 & ~n41308;
  assign n41310 = ~n8988 & ~n41303;
  assign n41311 = ~controllable_hmaster1 & ~n41310;
  assign n41312 = ~n41302 & ~n41311;
  assign n41313 = ~controllable_hgrant6 & ~n41312;
  assign n41314 = ~n13175 & ~n41313;
  assign n41315 = ~controllable_hmaster0 & ~n41314;
  assign n41316 = ~n41309 & ~n41315;
  assign n41317 = controllable_hmaster3 & ~n41316;
  assign n41318 = controllable_hgrant3 & ~n13315;
  assign n41319 = ~controllable_hgrant3 & ~n8987;
  assign n41320 = ~n41318 & ~n41319;
  assign n41321 = ~controllable_hgrant4 & ~n41320;
  assign n41322 = ~n13177 & ~n41321;
  assign n41323 = ~controllable_hgrant5 & ~n41322;
  assign n41324 = ~n13176 & ~n41323;
  assign n41325 = ~controllable_hmaster2 & ~n41324;
  assign n41326 = ~n10105 & ~n41325;
  assign n41327 = controllable_hmaster1 & ~n41326;
  assign n41328 = controllable_hgrant5 & ~n13319;
  assign n41329 = ~controllable_hgrant5 & ~n8987;
  assign n41330 = ~n41328 & ~n41329;
  assign n41331 = controllable_hmaster2 & ~n41330;
  assign n41332 = controllable_hgrant1 & ~n13313;
  assign n41333 = ~controllable_hgrant1 & ~n8987;
  assign n41334 = ~n41332 & ~n41333;
  assign n41335 = ~controllable_hgrant3 & ~n41334;
  assign n41336 = ~n13178 & ~n41335;
  assign n41337 = ~controllable_hgrant4 & ~n41336;
  assign n41338 = ~n13177 & ~n41337;
  assign n41339 = ~controllable_hgrant5 & ~n41338;
  assign n41340 = ~n13176 & ~n41339;
  assign n41341 = ~controllable_hmaster2 & ~n41340;
  assign n41342 = ~n41331 & ~n41341;
  assign n41343 = ~controllable_hmaster1 & ~n41342;
  assign n41344 = ~n41327 & ~n41343;
  assign n41345 = ~controllable_hgrant6 & ~n41344;
  assign n41346 = ~n13198 & ~n41345;
  assign n41347 = controllable_hmaster0 & ~n41346;
  assign n41348 = controllable_hgrant6 & ~n26891;
  assign n41349 = controllable_hgrant2 & ~n12627;
  assign n41350 = ~controllable_hgrant2 & ~n7735;
  assign n41351 = ~n41349 & ~n41350;
  assign n41352 = n7928 & ~n41351;
  assign n41353 = n7928 & ~n41352;
  assign n41354 = ~controllable_hgrant1 & ~n41353;
  assign n41355 = ~n13179 & ~n41354;
  assign n41356 = ~controllable_hgrant3 & ~n41355;
  assign n41357 = ~n13178 & ~n41356;
  assign n41358 = ~controllable_hgrant4 & ~n41357;
  assign n41359 = ~n13177 & ~n41358;
  assign n41360 = ~controllable_hgrant5 & ~n41359;
  assign n41361 = ~n13176 & ~n41360;
  assign n41362 = ~controllable_hmaster2 & ~n41361;
  assign n41363 = ~n10105 & ~n41362;
  assign n41364 = controllable_hmaster1 & ~n41363;
  assign n41365 = controllable_hgrant4 & ~n13317;
  assign n41366 = ~controllable_hgrant4 & ~n8987;
  assign n41367 = ~n41365 & ~n41366;
  assign n41368 = ~controllable_hgrant5 & ~n41367;
  assign n41369 = ~n13176 & ~n41368;
  assign n41370 = controllable_hmaster2 & ~n41369;
  assign n41371 = ~n8988 & ~n41370;
  assign n41372 = ~controllable_hmaster1 & ~n41371;
  assign n41373 = ~n41364 & ~n41372;
  assign n41374 = ~controllable_hgrant6 & ~n41373;
  assign n41375 = ~n41348 & ~n41374;
  assign n41376 = ~controllable_hmaster0 & ~n41375;
  assign n41377 = ~n41347 & ~n41376;
  assign n41378 = ~controllable_hmaster3 & ~n41377;
  assign n41379 = ~n41317 & ~n41378;
  assign n41380 = i_hbusreq7 & ~n41379;
  assign n41381 = i_hbusreq8 & ~n41316;
  assign n41382 = i_hbusreq6 & ~n41286;
  assign n41383 = n8217 & ~n9002;
  assign n41384 = ~n8217 & ~n29305;
  assign n41385 = ~n41383 & ~n41384;
  assign n41386 = ~i_hbusreq6 & ~n41385;
  assign n41387 = ~n41382 & ~n41386;
  assign n41388 = controllable_hgrant6 & ~n41387;
  assign n41389 = i_hbusreq6 & ~n41306;
  assign n41390 = i_hbusreq5 & ~n41299;
  assign n41391 = i_hbusreq4 & ~n41297;
  assign n41392 = i_hbusreq9 & ~n41297;
  assign n41393 = i_hbusreq3 & ~n41295;
  assign n41394 = i_hbusreq1 & ~n41293;
  assign n41395 = n7733 & ~n13348;
  assign n41396 = ~n7870 & ~n41395;
  assign n41397 = ~n7928 & ~n41396;
  assign n41398 = ~n7985 & ~n41395;
  assign n41399 = n7928 & ~n41398;
  assign n41400 = ~n41397 & ~n41399;
  assign n41401 = ~i_hbusreq1 & ~n41400;
  assign n41402 = ~n41394 & ~n41401;
  assign n41403 = ~controllable_hgrant1 & ~n41402;
  assign n41404 = ~n13213 & ~n41403;
  assign n41405 = ~i_hbusreq3 & ~n41404;
  assign n41406 = ~n41393 & ~n41405;
  assign n41407 = ~controllable_hgrant3 & ~n41406;
  assign n41408 = ~n13211 & ~n41407;
  assign n41409 = ~i_hbusreq9 & ~n41408;
  assign n41410 = ~n41392 & ~n41409;
  assign n41411 = ~i_hbusreq4 & ~n41410;
  assign n41412 = ~n41391 & ~n41411;
  assign n41413 = ~controllable_hgrant4 & ~n41412;
  assign n41414 = ~n13208 & ~n41413;
  assign n41415 = ~i_hbusreq5 & ~n41414;
  assign n41416 = ~n41390 & ~n41415;
  assign n41417 = ~controllable_hgrant5 & ~n41416;
  assign n41418 = ~n13206 & ~n41417;
  assign n41419 = controllable_hmaster1 & ~n41418;
  assign n41420 = controllable_hmaster2 & ~n41418;
  assign n41421 = ~n40407 & ~n41420;
  assign n41422 = ~controllable_hmaster1 & ~n41421;
  assign n41423 = ~n41419 & ~n41422;
  assign n41424 = ~i_hbusreq6 & ~n41423;
  assign n41425 = ~n41389 & ~n41424;
  assign n41426 = ~controllable_hgrant6 & ~n41425;
  assign n41427 = ~n41388 & ~n41426;
  assign n41428 = controllable_hmaster0 & ~n41427;
  assign n41429 = i_hbusreq6 & ~n41312;
  assign n41430 = ~n9024 & ~n41420;
  assign n41431 = ~controllable_hmaster1 & ~n41430;
  assign n41432 = ~n41419 & ~n41431;
  assign n41433 = ~i_hbusreq6 & ~n41432;
  assign n41434 = ~n41429 & ~n41433;
  assign n41435 = ~controllable_hgrant6 & ~n41434;
  assign n41436 = ~n13254 & ~n41435;
  assign n41437 = ~controllable_hmaster0 & ~n41436;
  assign n41438 = ~n41428 & ~n41437;
  assign n41439 = ~i_hbusreq8 & ~n41438;
  assign n41440 = ~n41381 & ~n41439;
  assign n41441 = controllable_hmaster3 & ~n41440;
  assign n41442 = i_hbusreq8 & ~n41377;
  assign n41443 = i_hbusreq6 & ~n41344;
  assign n41444 = i_hbusreq5 & ~n41322;
  assign n41445 = i_hbusreq4 & ~n41320;
  assign n41446 = i_hbusreq9 & ~n41320;
  assign n41447 = controllable_hgrant3 & ~n13356;
  assign n41448 = ~controllable_hgrant3 & ~n9017;
  assign n41449 = ~n41447 & ~n41448;
  assign n41450 = ~i_hbusreq9 & ~n41449;
  assign n41451 = ~n41446 & ~n41450;
  assign n41452 = ~i_hbusreq4 & ~n41451;
  assign n41453 = ~n41445 & ~n41452;
  assign n41454 = ~controllable_hgrant4 & ~n41453;
  assign n41455 = ~n13258 & ~n41454;
  assign n41456 = ~i_hbusreq5 & ~n41455;
  assign n41457 = ~n41444 & ~n41456;
  assign n41458 = ~controllable_hgrant5 & ~n41457;
  assign n41459 = ~n13256 & ~n41458;
  assign n41460 = ~controllable_hmaster2 & ~n41459;
  assign n41461 = ~n10116 & ~n41460;
  assign n41462 = controllable_hmaster1 & ~n41461;
  assign n41463 = controllable_hgrant5 & ~n13366;
  assign n41464 = ~controllable_hgrant5 & ~n9023;
  assign n41465 = ~n41463 & ~n41464;
  assign n41466 = controllable_hmaster2 & ~n41465;
  assign n41467 = i_hbusreq5 & ~n41338;
  assign n41468 = i_hbusreq4 & ~n41336;
  assign n41469 = i_hbusreq9 & ~n41336;
  assign n41470 = i_hbusreq3 & ~n41334;
  assign n41471 = controllable_hgrant1 & ~n13352;
  assign n41472 = ~controllable_hgrant1 & ~n9015;
  assign n41473 = ~n41471 & ~n41472;
  assign n41474 = ~i_hbusreq3 & ~n41473;
  assign n41475 = ~n41470 & ~n41474;
  assign n41476 = ~controllable_hgrant3 & ~n41475;
  assign n41477 = ~n13261 & ~n41476;
  assign n41478 = ~i_hbusreq9 & ~n41477;
  assign n41479 = ~n41469 & ~n41478;
  assign n41480 = ~i_hbusreq4 & ~n41479;
  assign n41481 = ~n41468 & ~n41480;
  assign n41482 = ~controllable_hgrant4 & ~n41481;
  assign n41483 = ~n13258 & ~n41482;
  assign n41484 = ~i_hbusreq5 & ~n41483;
  assign n41485 = ~n41467 & ~n41484;
  assign n41486 = ~controllable_hgrant5 & ~n41485;
  assign n41487 = ~n13256 & ~n41486;
  assign n41488 = ~controllable_hmaster2 & ~n41487;
  assign n41489 = ~n41466 & ~n41488;
  assign n41490 = ~controllable_hmaster1 & ~n41489;
  assign n41491 = ~n41462 & ~n41490;
  assign n41492 = ~i_hbusreq6 & ~n41491;
  assign n41493 = ~n41443 & ~n41492;
  assign n41494 = ~controllable_hgrant6 & ~n41493;
  assign n41495 = ~n13298 & ~n41494;
  assign n41496 = controllable_hmaster0 & ~n41495;
  assign n41497 = controllable_hgrant6 & ~n26906;
  assign n41498 = i_hbusreq6 & ~n41373;
  assign n41499 = i_hbusreq5 & ~n41359;
  assign n41500 = i_hbusreq4 & ~n41357;
  assign n41501 = i_hbusreq9 & ~n41357;
  assign n41502 = i_hbusreq3 & ~n41355;
  assign n41503 = i_hbusreq1 & ~n41353;
  assign n41504 = controllable_hgrant2 & ~n13346;
  assign n41505 = ~controllable_hgrant2 & ~n7757;
  assign n41506 = ~n41504 & ~n41505;
  assign n41507 = n7928 & ~n41506;
  assign n41508 = n7928 & ~n41507;
  assign n41509 = ~i_hbusreq1 & ~n41508;
  assign n41510 = ~n41503 & ~n41509;
  assign n41511 = ~controllable_hgrant1 & ~n41510;
  assign n41512 = ~n13263 & ~n41511;
  assign n41513 = ~i_hbusreq3 & ~n41512;
  assign n41514 = ~n41502 & ~n41513;
  assign n41515 = ~controllable_hgrant3 & ~n41514;
  assign n41516 = ~n13261 & ~n41515;
  assign n41517 = ~i_hbusreq9 & ~n41516;
  assign n41518 = ~n41501 & ~n41517;
  assign n41519 = ~i_hbusreq4 & ~n41518;
  assign n41520 = ~n41500 & ~n41519;
  assign n41521 = ~controllable_hgrant4 & ~n41520;
  assign n41522 = ~n13258 & ~n41521;
  assign n41523 = ~i_hbusreq5 & ~n41522;
  assign n41524 = ~n41499 & ~n41523;
  assign n41525 = ~controllable_hgrant5 & ~n41524;
  assign n41526 = ~n13256 & ~n41525;
  assign n41527 = ~controllable_hmaster2 & ~n41526;
  assign n41528 = ~n10116 & ~n41527;
  assign n41529 = controllable_hmaster1 & ~n41528;
  assign n41530 = i_hbusreq5 & ~n41367;
  assign n41531 = controllable_hgrant4 & ~n13362;
  assign n41532 = ~controllable_hgrant4 & ~n9021;
  assign n41533 = ~n41531 & ~n41532;
  assign n41534 = ~i_hbusreq5 & ~n41533;
  assign n41535 = ~n41530 & ~n41534;
  assign n41536 = ~controllable_hgrant5 & ~n41535;
  assign n41537 = ~n13256 & ~n41536;
  assign n41538 = controllable_hmaster2 & ~n41537;
  assign n41539 = ~n9024 & ~n41538;
  assign n41540 = ~controllable_hmaster1 & ~n41539;
  assign n41541 = ~n41529 & ~n41540;
  assign n41542 = ~i_hbusreq6 & ~n41541;
  assign n41543 = ~n41498 & ~n41542;
  assign n41544 = ~controllable_hgrant6 & ~n41543;
  assign n41545 = ~n41497 & ~n41544;
  assign n41546 = ~controllable_hmaster0 & ~n41545;
  assign n41547 = ~n41496 & ~n41546;
  assign n41548 = ~i_hbusreq8 & ~n41547;
  assign n41549 = ~n41442 & ~n41548;
  assign n41550 = ~controllable_hmaster3 & ~n41549;
  assign n41551 = ~n41441 & ~n41550;
  assign n41552 = ~i_hbusreq7 & ~n41551;
  assign n41553 = ~n41380 & ~n41552;
  assign n41554 = ~n7924 & ~n41553;
  assign n41555 = n8217 & ~n26928;
  assign n41556 = ~n8217 & ~n29329;
  assign n41557 = ~n41555 & ~n41556;
  assign n41558 = controllable_hgrant6 & ~n41557;
  assign n41559 = controllable_hgrant5 & ~n13164;
  assign n41560 = controllable_hgrant4 & ~n13162;
  assign n41561 = controllable_hgrant3 & ~n13160;
  assign n41562 = controllable_hgrant1 & ~n13158;
  assign n41563 = controllable_hgrant2 & ~n13009;
  assign n41564 = ~n7733 & n41563;
  assign n41565 = ~n12801 & ~n41563;
  assign n41566 = n7733 & ~n41565;
  assign n41567 = ~n41564 & ~n41566;
  assign n41568 = n7928 & ~n41567;
  assign n41569 = ~n41290 & ~n41568;
  assign n41570 = ~controllable_hgrant1 & ~n41569;
  assign n41571 = ~n41562 & ~n41570;
  assign n41572 = ~controllable_hgrant3 & ~n41571;
  assign n41573 = ~n41561 & ~n41572;
  assign n41574 = ~controllable_hgrant4 & ~n41573;
  assign n41575 = ~n41560 & ~n41574;
  assign n41576 = ~controllable_hgrant5 & ~n41575;
  assign n41577 = ~n41559 & ~n41576;
  assign n41578 = controllable_hmaster1 & ~n41577;
  assign n41579 = controllable_hmaster2 & ~n41577;
  assign n41580 = n8378 & ~n26922;
  assign n41581 = ~n8378 & ~n29323;
  assign n41582 = ~n41580 & ~n41581;
  assign n41583 = controllable_hgrant5 & ~n41582;
  assign n41584 = n8426 & ~n13413;
  assign n41585 = ~n8426 & ~n17771;
  assign n41586 = ~n41584 & ~n41585;
  assign n41587 = i_hlock9 & ~n41586;
  assign n41588 = n8426 & ~n13434;
  assign n41589 = ~n8426 & ~n17789;
  assign n41590 = ~n41588 & ~n41589;
  assign n41591 = ~i_hlock9 & ~n41590;
  assign n41592 = ~n41587 & ~n41591;
  assign n41593 = controllable_hgrant4 & ~n41592;
  assign n41594 = n8365 & ~n13411;
  assign n41595 = ~n8365 & ~n17769;
  assign n41596 = ~n41594 & ~n41595;
  assign n41597 = controllable_hgrant3 & ~n41596;
  assign n41598 = n8389 & ~n13409;
  assign n41599 = ~n8389 & ~n17767;
  assign n41600 = ~n41598 & ~n41599;
  assign n41601 = controllable_hgrant1 & ~n41600;
  assign n41602 = ~controllable_locked & n40215;
  assign n41603 = ~n13008 & ~n41602;
  assign n41604 = controllable_hgrant2 & ~n41603;
  assign n41605 = ~n7733 & n41604;
  assign n41606 = ~n40224 & ~n41602;
  assign n41607 = controllable_hgrant2 & ~n41606;
  assign n41608 = ~n17089 & ~n17756;
  assign n41609 = ~controllable_hgrant2 & ~n41608;
  assign n41610 = ~n41607 & ~n41609;
  assign n41611 = n7733 & ~n41610;
  assign n41612 = ~n41605 & ~n41611;
  assign n41613 = n7928 & ~n41612;
  assign n41614 = ~n8221 & ~n41613;
  assign n41615 = ~controllable_hgrant1 & ~n41614;
  assign n41616 = ~n41601 & ~n41615;
  assign n41617 = ~controllable_hgrant3 & ~n41616;
  assign n41618 = ~n41597 & ~n41617;
  assign n41619 = i_hlock9 & ~n41618;
  assign n41620 = n8365 & ~n13432;
  assign n41621 = ~n8365 & ~n17787;
  assign n41622 = ~n41620 & ~n41621;
  assign n41623 = controllable_hgrant3 & ~n41622;
  assign n41624 = n8389 & ~n13430;
  assign n41625 = ~n8389 & ~n17785;
  assign n41626 = ~n41624 & ~n41625;
  assign n41627 = controllable_hgrant1 & ~n41626;
  assign n41628 = ~n8235 & ~n41613;
  assign n41629 = ~controllable_hgrant1 & ~n41628;
  assign n41630 = ~n41627 & ~n41629;
  assign n41631 = ~controllable_hgrant3 & ~n41630;
  assign n41632 = ~n41623 & ~n41631;
  assign n41633 = ~i_hlock9 & ~n41632;
  assign n41634 = ~n41619 & ~n41633;
  assign n41635 = ~controllable_hgrant4 & ~n41634;
  assign n41636 = ~n41593 & ~n41635;
  assign n41637 = ~controllable_hgrant5 & ~n41636;
  assign n41638 = ~n41583 & ~n41637;
  assign n41639 = ~controllable_hmaster2 & ~n41638;
  assign n41640 = ~n41579 & ~n41639;
  assign n41641 = ~controllable_hmaster1 & ~n41640;
  assign n41642 = ~n41578 & ~n41641;
  assign n41643 = ~controllable_hgrant6 & ~n41642;
  assign n41644 = ~n41558 & ~n41643;
  assign n41645 = controllable_hmaster0 & ~n41644;
  assign n41646 = controllable_hgrant6 & ~n13192;
  assign n41647 = controllable_hgrant5 & ~n13186;
  assign n41648 = controllable_hgrant4 & ~n13184;
  assign n41649 = controllable_hgrant3 & ~n13182;
  assign n41650 = controllable_hgrant1 & ~n13180;
  assign n41651 = ~controllable_hgrant2 & n7971;
  assign n41652 = ~n41563 & ~n41651;
  assign n41653 = ~n7733 & ~n41652;
  assign n41654 = n7733 & ~n13009;
  assign n41655 = ~n41653 & ~n41654;
  assign n41656 = n7928 & ~n41655;
  assign n41657 = n7928 & ~n41656;
  assign n41658 = ~controllable_hgrant1 & ~n41657;
  assign n41659 = ~n41650 & ~n41658;
  assign n41660 = ~controllable_hgrant3 & ~n41659;
  assign n41661 = ~n41649 & ~n41660;
  assign n41662 = ~controllable_hgrant4 & ~n41661;
  assign n41663 = ~n41648 & ~n41662;
  assign n41664 = ~controllable_hgrant5 & ~n41663;
  assign n41665 = ~n41647 & ~n41664;
  assign n41666 = ~controllable_hmaster2 & ~n41665;
  assign n41667 = ~n41579 & ~n41666;
  assign n41668 = ~controllable_hmaster1 & ~n41667;
  assign n41669 = ~n41578 & ~n41668;
  assign n41670 = ~controllable_hgrant6 & ~n41669;
  assign n41671 = ~n41646 & ~n41670;
  assign n41672 = ~controllable_hmaster0 & ~n41671;
  assign n41673 = ~n41645 & ~n41672;
  assign n41674 = controllable_hmaster3 & ~n41673;
  assign n41675 = controllable_hgrant6 & ~n13188;
  assign n41676 = controllable_hmaster2 & ~n41665;
  assign n41677 = controllable_hgrant3 & ~n13392;
  assign n41678 = ~n41660 & ~n41677;
  assign n41679 = ~controllable_hgrant4 & ~n41678;
  assign n41680 = ~n41648 & ~n41679;
  assign n41681 = ~controllable_hgrant5 & ~n41680;
  assign n41682 = ~n41647 & ~n41681;
  assign n41683 = ~controllable_hmaster2 & ~n41682;
  assign n41684 = ~n41676 & ~n41683;
  assign n41685 = controllable_hmaster1 & ~n41684;
  assign n41686 = controllable_hgrant5 & ~n13396;
  assign n41687 = ~n41664 & ~n41686;
  assign n41688 = controllable_hmaster2 & ~n41687;
  assign n41689 = controllable_hgrant1 & ~n13390;
  assign n41690 = ~n41658 & ~n41689;
  assign n41691 = ~controllable_hgrant3 & ~n41690;
  assign n41692 = ~n41649 & ~n41691;
  assign n41693 = ~controllable_hgrant4 & ~n41692;
  assign n41694 = ~n41648 & ~n41693;
  assign n41695 = ~controllable_hgrant5 & ~n41694;
  assign n41696 = ~n41647 & ~n41695;
  assign n41697 = ~controllable_hmaster2 & ~n41696;
  assign n41698 = ~n41688 & ~n41697;
  assign n41699 = ~controllable_hmaster1 & ~n41698;
  assign n41700 = ~n41685 & ~n41699;
  assign n41701 = ~controllable_hgrant6 & ~n41700;
  assign n41702 = ~n41675 & ~n41701;
  assign n41703 = controllable_hmaster0 & ~n41702;
  assign n41704 = controllable_hgrant6 & ~n26937;
  assign n41705 = controllable_hgrant2 & ~n12800;
  assign n41706 = ~n41651 & ~n41705;
  assign n41707 = ~n7733 & ~n41706;
  assign n41708 = ~n13010 & ~n41705;
  assign n41709 = n7733 & ~n41708;
  assign n41710 = ~n41707 & ~n41709;
  assign n41711 = n7928 & ~n41710;
  assign n41712 = n7928 & ~n41711;
  assign n41713 = ~controllable_hgrant1 & ~n41712;
  assign n41714 = ~n41650 & ~n41713;
  assign n41715 = ~controllable_hgrant3 & ~n41714;
  assign n41716 = ~n41649 & ~n41715;
  assign n41717 = ~controllable_hgrant4 & ~n41716;
  assign n41718 = ~n41648 & ~n41717;
  assign n41719 = ~controllable_hgrant5 & ~n41718;
  assign n41720 = ~n41647 & ~n41719;
  assign n41721 = ~controllable_hmaster2 & ~n41720;
  assign n41722 = ~n41676 & ~n41721;
  assign n41723 = controllable_hmaster1 & ~n41722;
  assign n41724 = controllable_hgrant4 & ~n13394;
  assign n41725 = ~n41662 & ~n41724;
  assign n41726 = ~controllable_hgrant5 & ~n41725;
  assign n41727 = ~n41647 & ~n41726;
  assign n41728 = controllable_hmaster2 & ~n41727;
  assign n41729 = ~n41666 & ~n41728;
  assign n41730 = ~controllable_hmaster1 & ~n41729;
  assign n41731 = ~n41723 & ~n41730;
  assign n41732 = ~controllable_hgrant6 & ~n41731;
  assign n41733 = ~n41704 & ~n41732;
  assign n41734 = ~controllable_hmaster0 & ~n41733;
  assign n41735 = ~n41703 & ~n41734;
  assign n41736 = ~controllable_hmaster3 & ~n41735;
  assign n41737 = ~n41674 & ~n41736;
  assign n41738 = i_hbusreq7 & ~n41737;
  assign n41739 = i_hbusreq8 & ~n41673;
  assign n41740 = i_hbusreq6 & ~n41557;
  assign n41741 = n8217 & ~n26966;
  assign n41742 = ~n8217 & ~n29358;
  assign n41743 = ~n41741 & ~n41742;
  assign n41744 = ~i_hbusreq6 & ~n41743;
  assign n41745 = ~n41740 & ~n41744;
  assign n41746 = controllable_hgrant6 & ~n41745;
  assign n41747 = i_hbusreq6 & ~n41642;
  assign n41748 = controllable_hgrant5 & ~n13476;
  assign n41749 = i_hbusreq5 & ~n41575;
  assign n41750 = controllable_hgrant4 & ~n13472;
  assign n41751 = i_hbusreq4 & ~n41573;
  assign n41752 = i_hbusreq9 & ~n41573;
  assign n41753 = controllable_hgrant3 & ~n13466;
  assign n41754 = i_hbusreq3 & ~n41571;
  assign n41755 = controllable_hgrant1 & ~n13462;
  assign n41756 = i_hbusreq1 & ~n41569;
  assign n41757 = controllable_hgrant2 & ~n13456;
  assign n41758 = ~n8074 & ~n41757;
  assign n41759 = ~n7733 & ~n41758;
  assign n41760 = ~n13489 & ~n41757;
  assign n41761 = n7733 & ~n41760;
  assign n41762 = ~n41759 & ~n41761;
  assign n41763 = n7928 & ~n41762;
  assign n41764 = ~n41397 & ~n41763;
  assign n41765 = ~i_hbusreq1 & ~n41764;
  assign n41766 = ~n41756 & ~n41765;
  assign n41767 = ~controllable_hgrant1 & ~n41766;
  assign n41768 = ~n41755 & ~n41767;
  assign n41769 = ~i_hbusreq3 & ~n41768;
  assign n41770 = ~n41754 & ~n41769;
  assign n41771 = ~controllable_hgrant3 & ~n41770;
  assign n41772 = ~n41753 & ~n41771;
  assign n41773 = ~i_hbusreq9 & ~n41772;
  assign n41774 = ~n41752 & ~n41773;
  assign n41775 = ~i_hbusreq4 & ~n41774;
  assign n41776 = ~n41751 & ~n41775;
  assign n41777 = ~controllable_hgrant4 & ~n41776;
  assign n41778 = ~n41750 & ~n41777;
  assign n41779 = ~i_hbusreq5 & ~n41778;
  assign n41780 = ~n41749 & ~n41779;
  assign n41781 = ~controllable_hgrant5 & ~n41780;
  assign n41782 = ~n41748 & ~n41781;
  assign n41783 = controllable_hmaster1 & ~n41782;
  assign n41784 = controllable_hmaster2 & ~n41782;
  assign n41785 = i_hbusreq5 & ~n41582;
  assign n41786 = n8378 & ~n26958;
  assign n41787 = ~n8378 & ~n29350;
  assign n41788 = ~n41786 & ~n41787;
  assign n41789 = ~i_hbusreq5 & ~n41788;
  assign n41790 = ~n41785 & ~n41789;
  assign n41791 = controllable_hgrant5 & ~n41790;
  assign n41792 = i_hbusreq5 & ~n41636;
  assign n41793 = i_hbusreq4 & ~n41592;
  assign n41794 = i_hbusreq9 & ~n41592;
  assign n41795 = n8426 & ~n13551;
  assign n41796 = ~n8426 & ~n17840;
  assign n41797 = ~n41795 & ~n41796;
  assign n41798 = i_hlock9 & ~n41797;
  assign n41799 = n8426 & ~n13590;
  assign n41800 = ~n8426 & ~n17876;
  assign n41801 = ~n41799 & ~n41800;
  assign n41802 = ~i_hlock9 & ~n41801;
  assign n41803 = ~n41798 & ~n41802;
  assign n41804 = ~i_hbusreq9 & ~n41803;
  assign n41805 = ~n41794 & ~n41804;
  assign n41806 = ~i_hbusreq4 & ~n41805;
  assign n41807 = ~n41793 & ~n41806;
  assign n41808 = controllable_hgrant4 & ~n41807;
  assign n41809 = i_hbusreq4 & ~n41634;
  assign n41810 = i_hbusreq9 & ~n41634;
  assign n41811 = i_hbusreq3 & ~n41596;
  assign n41812 = n8365 & ~n13547;
  assign n41813 = ~n8365 & ~n17836;
  assign n41814 = ~n41812 & ~n41813;
  assign n41815 = ~i_hbusreq3 & ~n41814;
  assign n41816 = ~n41811 & ~n41815;
  assign n41817 = controllable_hgrant3 & ~n41816;
  assign n41818 = i_hbusreq3 & ~n41616;
  assign n41819 = i_hbusreq1 & ~n41600;
  assign n41820 = n8389 & ~n13543;
  assign n41821 = ~n8389 & ~n17832;
  assign n41822 = ~n41820 & ~n41821;
  assign n41823 = ~i_hbusreq1 & ~n41822;
  assign n41824 = ~n41819 & ~n41823;
  assign n41825 = controllable_hgrant1 & ~n41824;
  assign n41826 = i_hbusreq1 & ~n41614;
  assign n41827 = i_hbusreq2 & ~n41603;
  assign n41828 = i_hbusreq0 & ~n41603;
  assign n41829 = ~n40326 & ~n41828;
  assign n41830 = ~i_hbusreq2 & ~n41829;
  assign n41831 = ~n41827 & ~n41830;
  assign n41832 = controllable_hgrant2 & ~n41831;
  assign n41833 = ~n40876 & ~n41832;
  assign n41834 = ~n7733 & ~n41833;
  assign n41835 = i_hbusreq2 & ~n41606;
  assign n41836 = i_hbusreq0 & ~n41606;
  assign n41837 = ~n40344 & ~n41836;
  assign n41838 = ~i_hbusreq2 & ~n41837;
  assign n41839 = ~n41835 & ~n41838;
  assign n41840 = controllable_hgrant2 & ~n41839;
  assign n41841 = i_hbusreq2 & ~n41608;
  assign n41842 = i_hbusreq0 & ~n41608;
  assign n41843 = ~n40351 & ~n41842;
  assign n41844 = ~i_hbusreq2 & ~n41843;
  assign n41845 = ~n41841 & ~n41844;
  assign n41846 = ~controllable_hgrant2 & ~n41845;
  assign n41847 = ~n41840 & ~n41846;
  assign n41848 = n7733 & ~n41847;
  assign n41849 = ~n41834 & ~n41848;
  assign n41850 = n7928 & ~n41849;
  assign n41851 = ~n8265 & ~n41850;
  assign n41852 = ~i_hbusreq1 & ~n41851;
  assign n41853 = ~n41826 & ~n41852;
  assign n41854 = ~controllable_hgrant1 & ~n41853;
  assign n41855 = ~n41825 & ~n41854;
  assign n41856 = ~i_hbusreq3 & ~n41855;
  assign n41857 = ~n41818 & ~n41856;
  assign n41858 = ~controllable_hgrant3 & ~n41857;
  assign n41859 = ~n41817 & ~n41858;
  assign n41860 = i_hlock9 & ~n41859;
  assign n41861 = i_hbusreq3 & ~n41622;
  assign n41862 = n8365 & ~n13586;
  assign n41863 = ~n8365 & ~n17872;
  assign n41864 = ~n41862 & ~n41863;
  assign n41865 = ~i_hbusreq3 & ~n41864;
  assign n41866 = ~n41861 & ~n41865;
  assign n41867 = controllable_hgrant3 & ~n41866;
  assign n41868 = i_hbusreq3 & ~n41630;
  assign n41869 = i_hbusreq1 & ~n41626;
  assign n41870 = n8389 & ~n13582;
  assign n41871 = ~n8389 & ~n17868;
  assign n41872 = ~n41870 & ~n41871;
  assign n41873 = ~i_hbusreq1 & ~n41872;
  assign n41874 = ~n41869 & ~n41873;
  assign n41875 = controllable_hgrant1 & ~n41874;
  assign n41876 = i_hbusreq1 & ~n41628;
  assign n41877 = ~n8297 & ~n41850;
  assign n41878 = ~i_hbusreq1 & ~n41877;
  assign n41879 = ~n41876 & ~n41878;
  assign n41880 = ~controllable_hgrant1 & ~n41879;
  assign n41881 = ~n41875 & ~n41880;
  assign n41882 = ~i_hbusreq3 & ~n41881;
  assign n41883 = ~n41868 & ~n41882;
  assign n41884 = ~controllable_hgrant3 & ~n41883;
  assign n41885 = ~n41867 & ~n41884;
  assign n41886 = ~i_hlock9 & ~n41885;
  assign n41887 = ~n41860 & ~n41886;
  assign n41888 = ~i_hbusreq9 & ~n41887;
  assign n41889 = ~n41810 & ~n41888;
  assign n41890 = ~i_hbusreq4 & ~n41889;
  assign n41891 = ~n41809 & ~n41890;
  assign n41892 = ~controllable_hgrant4 & ~n41891;
  assign n41893 = ~n41808 & ~n41892;
  assign n41894 = ~i_hbusreq5 & ~n41893;
  assign n41895 = ~n41792 & ~n41894;
  assign n41896 = ~controllable_hgrant5 & ~n41895;
  assign n41897 = ~n41791 & ~n41896;
  assign n41898 = ~controllable_hmaster2 & ~n41897;
  assign n41899 = ~n41784 & ~n41898;
  assign n41900 = ~controllable_hmaster1 & ~n41899;
  assign n41901 = ~n41783 & ~n41900;
  assign n41902 = ~i_hbusreq6 & ~n41901;
  assign n41903 = ~n41747 & ~n41902;
  assign n41904 = ~controllable_hgrant6 & ~n41903;
  assign n41905 = ~n41746 & ~n41904;
  assign n41906 = controllable_hmaster0 & ~n41905;
  assign n41907 = controllable_hgrant6 & ~n13707;
  assign n41908 = i_hbusreq6 & ~n41669;
  assign n41909 = controllable_hgrant5 & ~n13632;
  assign n41910 = i_hbusreq5 & ~n41663;
  assign n41911 = controllable_hgrant4 & ~n13628;
  assign n41912 = i_hbusreq4 & ~n41661;
  assign n41913 = i_hbusreq9 & ~n41661;
  assign n41914 = controllable_hgrant3 & ~n13622;
  assign n41915 = i_hbusreq3 & ~n41659;
  assign n41916 = controllable_hgrant1 & ~n13618;
  assign n41917 = i_hbusreq1 & ~n41657;
  assign n41918 = i_hbusreq2 & ~n7971;
  assign n41919 = i_hbusreq0 & ~n7971;
  assign n41920 = ~n8107 & ~n41919;
  assign n41921 = ~i_hbusreq2 & ~n41920;
  assign n41922 = ~n41918 & ~n41921;
  assign n41923 = ~controllable_hgrant2 & n41922;
  assign n41924 = ~n41757 & ~n41923;
  assign n41925 = ~n7733 & ~n41924;
  assign n41926 = n7733 & ~n13456;
  assign n41927 = ~n41925 & ~n41926;
  assign n41928 = n7928 & ~n41927;
  assign n41929 = n7928 & ~n41928;
  assign n41930 = ~i_hbusreq1 & ~n41929;
  assign n41931 = ~n41917 & ~n41930;
  assign n41932 = ~controllable_hgrant1 & ~n41931;
  assign n41933 = ~n41916 & ~n41932;
  assign n41934 = ~i_hbusreq3 & ~n41933;
  assign n41935 = ~n41915 & ~n41934;
  assign n41936 = ~controllable_hgrant3 & ~n41935;
  assign n41937 = ~n41914 & ~n41936;
  assign n41938 = ~i_hbusreq9 & ~n41937;
  assign n41939 = ~n41913 & ~n41938;
  assign n41940 = ~i_hbusreq4 & ~n41939;
  assign n41941 = ~n41912 & ~n41940;
  assign n41942 = ~controllable_hgrant4 & ~n41941;
  assign n41943 = ~n41911 & ~n41942;
  assign n41944 = ~i_hbusreq5 & ~n41943;
  assign n41945 = ~n41910 & ~n41944;
  assign n41946 = ~controllable_hgrant5 & ~n41945;
  assign n41947 = ~n41909 & ~n41946;
  assign n41948 = ~controllable_hmaster2 & ~n41947;
  assign n41949 = ~n41784 & ~n41948;
  assign n41950 = ~controllable_hmaster1 & ~n41949;
  assign n41951 = ~n41783 & ~n41950;
  assign n41952 = ~i_hbusreq6 & ~n41951;
  assign n41953 = ~n41908 & ~n41952;
  assign n41954 = ~controllable_hgrant6 & ~n41953;
  assign n41955 = ~n41907 & ~n41954;
  assign n41956 = ~controllable_hmaster0 & ~n41955;
  assign n41957 = ~n41906 & ~n41956;
  assign n41958 = ~i_hbusreq8 & ~n41957;
  assign n41959 = ~n41739 & ~n41958;
  assign n41960 = controllable_hmaster3 & ~n41959;
  assign n41961 = i_hbusreq8 & ~n41735;
  assign n41962 = controllable_hgrant6 & ~n13636;
  assign n41963 = i_hbusreq6 & ~n41700;
  assign n41964 = controllable_hmaster2 & ~n41947;
  assign n41965 = i_hbusreq5 & ~n41680;
  assign n41966 = i_hbusreq4 & ~n41678;
  assign n41967 = i_hbusreq9 & ~n41678;
  assign n41968 = controllable_hgrant3 & ~n13498;
  assign n41969 = ~n41936 & ~n41968;
  assign n41970 = ~i_hbusreq9 & ~n41969;
  assign n41971 = ~n41967 & ~n41970;
  assign n41972 = ~i_hbusreq4 & ~n41971;
  assign n41973 = ~n41966 & ~n41972;
  assign n41974 = ~controllable_hgrant4 & ~n41973;
  assign n41975 = ~n41911 & ~n41974;
  assign n41976 = ~i_hbusreq5 & ~n41975;
  assign n41977 = ~n41965 & ~n41976;
  assign n41978 = ~controllable_hgrant5 & ~n41977;
  assign n41979 = ~n41909 & ~n41978;
  assign n41980 = ~controllable_hmaster2 & ~n41979;
  assign n41981 = ~n41964 & ~n41980;
  assign n41982 = controllable_hmaster1 & ~n41981;
  assign n41983 = controllable_hgrant5 & ~n13508;
  assign n41984 = ~n41946 & ~n41983;
  assign n41985 = controllable_hmaster2 & ~n41984;
  assign n41986 = i_hbusreq5 & ~n41694;
  assign n41987 = i_hbusreq4 & ~n41692;
  assign n41988 = i_hbusreq9 & ~n41692;
  assign n41989 = i_hbusreq3 & ~n41690;
  assign n41990 = controllable_hgrant1 & ~n13494;
  assign n41991 = ~n41932 & ~n41990;
  assign n41992 = ~i_hbusreq3 & ~n41991;
  assign n41993 = ~n41989 & ~n41992;
  assign n41994 = ~controllable_hgrant3 & ~n41993;
  assign n41995 = ~n41914 & ~n41994;
  assign n41996 = ~i_hbusreq9 & ~n41995;
  assign n41997 = ~n41988 & ~n41996;
  assign n41998 = ~i_hbusreq4 & ~n41997;
  assign n41999 = ~n41987 & ~n41998;
  assign n42000 = ~controllable_hgrant4 & ~n41999;
  assign n42001 = ~n41911 & ~n42000;
  assign n42002 = ~i_hbusreq5 & ~n42001;
  assign n42003 = ~n41986 & ~n42002;
  assign n42004 = ~controllable_hgrant5 & ~n42003;
  assign n42005 = ~n41909 & ~n42004;
  assign n42006 = ~controllable_hmaster2 & ~n42005;
  assign n42007 = ~n41985 & ~n42006;
  assign n42008 = ~controllable_hmaster1 & ~n42007;
  assign n42009 = ~n41982 & ~n42008;
  assign n42010 = ~i_hbusreq6 & ~n42009;
  assign n42011 = ~n41963 & ~n42010;
  assign n42012 = ~controllable_hgrant6 & ~n42011;
  assign n42013 = ~n41962 & ~n42012;
  assign n42014 = controllable_hmaster0 & ~n42013;
  assign n42015 = controllable_hgrant6 & ~n26983;
  assign n42016 = i_hbusreq6 & ~n41731;
  assign n42017 = i_hbusreq5 & ~n41718;
  assign n42018 = i_hbusreq4 & ~n41716;
  assign n42019 = i_hbusreq9 & ~n41716;
  assign n42020 = i_hbusreq3 & ~n41714;
  assign n42021 = i_hbusreq1 & ~n41712;
  assign n42022 = controllable_hgrant2 & ~n13488;
  assign n42023 = ~n41923 & ~n42022;
  assign n42024 = ~n7733 & ~n42023;
  assign n42025 = ~n13457 & ~n42022;
  assign n42026 = n7733 & ~n42025;
  assign n42027 = ~n42024 & ~n42026;
  assign n42028 = n7928 & ~n42027;
  assign n42029 = n7928 & ~n42028;
  assign n42030 = ~i_hbusreq1 & ~n42029;
  assign n42031 = ~n42021 & ~n42030;
  assign n42032 = ~controllable_hgrant1 & ~n42031;
  assign n42033 = ~n41916 & ~n42032;
  assign n42034 = ~i_hbusreq3 & ~n42033;
  assign n42035 = ~n42020 & ~n42034;
  assign n42036 = ~controllable_hgrant3 & ~n42035;
  assign n42037 = ~n41914 & ~n42036;
  assign n42038 = ~i_hbusreq9 & ~n42037;
  assign n42039 = ~n42019 & ~n42038;
  assign n42040 = ~i_hbusreq4 & ~n42039;
  assign n42041 = ~n42018 & ~n42040;
  assign n42042 = ~controllable_hgrant4 & ~n42041;
  assign n42043 = ~n41911 & ~n42042;
  assign n42044 = ~i_hbusreq5 & ~n42043;
  assign n42045 = ~n42017 & ~n42044;
  assign n42046 = ~controllable_hgrant5 & ~n42045;
  assign n42047 = ~n41909 & ~n42046;
  assign n42048 = ~controllable_hmaster2 & ~n42047;
  assign n42049 = ~n41964 & ~n42048;
  assign n42050 = controllable_hmaster1 & ~n42049;
  assign n42051 = i_hbusreq5 & ~n41725;
  assign n42052 = controllable_hgrant4 & ~n13504;
  assign n42053 = ~n41942 & ~n42052;
  assign n42054 = ~i_hbusreq5 & ~n42053;
  assign n42055 = ~n42051 & ~n42054;
  assign n42056 = ~controllable_hgrant5 & ~n42055;
  assign n42057 = ~n41909 & ~n42056;
  assign n42058 = controllable_hmaster2 & ~n42057;
  assign n42059 = ~n41948 & ~n42058;
  assign n42060 = ~controllable_hmaster1 & ~n42059;
  assign n42061 = ~n42050 & ~n42060;
  assign n42062 = ~i_hbusreq6 & ~n42061;
  assign n42063 = ~n42016 & ~n42062;
  assign n42064 = ~controllable_hgrant6 & ~n42063;
  assign n42065 = ~n42015 & ~n42064;
  assign n42066 = ~controllable_hmaster0 & ~n42065;
  assign n42067 = ~n42014 & ~n42066;
  assign n42068 = ~i_hbusreq8 & ~n42067;
  assign n42069 = ~n41961 & ~n42068;
  assign n42070 = ~controllable_hmaster3 & ~n42069;
  assign n42071 = ~n41960 & ~n42070;
  assign n42072 = ~i_hbusreq7 & ~n42071;
  assign n42073 = ~n41738 & ~n42072;
  assign n42074 = n7924 & ~n42073;
  assign n42075 = ~n41554 & ~n42074;
  assign n42076 = ~n8214 & ~n42075;
  assign n42077 = controllable_hmaster0 & ~n41314;
  assign n42078 = n8217 & ~n9049;
  assign n42079 = ~n8217 & ~n17707;
  assign n42080 = ~n42078 & ~n42079;
  assign n42081 = controllable_hgrant6 & ~n42080;
  assign n42082 = ~n40437 & ~n41303;
  assign n42083 = ~controllable_hmaster1 & ~n42082;
  assign n42084 = ~n41302 & ~n42083;
  assign n42085 = ~controllable_hgrant6 & ~n42084;
  assign n42086 = ~n42081 & ~n42085;
  assign n42087 = ~controllable_hmaster0 & ~n42086;
  assign n42088 = ~n42077 & ~n42087;
  assign n42089 = i_hlock8 & ~n42088;
  assign n42090 = n8217 & ~n9055;
  assign n42091 = ~n8217 & ~n17715;
  assign n42092 = ~n42090 & ~n42091;
  assign n42093 = controllable_hgrant6 & ~n42092;
  assign n42094 = ~n40459 & ~n41303;
  assign n42095 = ~controllable_hmaster1 & ~n42094;
  assign n42096 = ~n41302 & ~n42095;
  assign n42097 = ~controllable_hgrant6 & ~n42096;
  assign n42098 = ~n42093 & ~n42097;
  assign n42099 = ~controllable_hmaster0 & ~n42098;
  assign n42100 = ~n42077 & ~n42099;
  assign n42101 = ~i_hlock8 & ~n42100;
  assign n42102 = ~n42089 & ~n42101;
  assign n42103 = controllable_hmaster3 & ~n42102;
  assign n42104 = ~n41378 & ~n42103;
  assign n42105 = i_hbusreq7 & ~n42104;
  assign n42106 = i_hbusreq8 & ~n42102;
  assign n42107 = controllable_hmaster0 & ~n41436;
  assign n42108 = i_hbusreq6 & ~n42080;
  assign n42109 = n8217 & ~n9068;
  assign n42110 = ~n8217 & ~n17729;
  assign n42111 = ~n42109 & ~n42110;
  assign n42112 = ~i_hbusreq6 & ~n42111;
  assign n42113 = ~n42108 & ~n42112;
  assign n42114 = controllable_hgrant6 & ~n42113;
  assign n42115 = i_hbusreq6 & ~n42084;
  assign n42116 = ~n40508 & ~n41420;
  assign n42117 = ~controllable_hmaster1 & ~n42116;
  assign n42118 = ~n41419 & ~n42117;
  assign n42119 = ~i_hbusreq6 & ~n42118;
  assign n42120 = ~n42115 & ~n42119;
  assign n42121 = ~controllable_hgrant6 & ~n42120;
  assign n42122 = ~n42114 & ~n42121;
  assign n42123 = ~controllable_hmaster0 & ~n42122;
  assign n42124 = ~n42107 & ~n42123;
  assign n42125 = i_hlock8 & ~n42124;
  assign n42126 = i_hbusreq6 & ~n42092;
  assign n42127 = n8217 & ~n9077;
  assign n42128 = ~n8217 & ~n17740;
  assign n42129 = ~n42127 & ~n42128;
  assign n42130 = ~i_hbusreq6 & ~n42129;
  assign n42131 = ~n42126 & ~n42130;
  assign n42132 = controllable_hgrant6 & ~n42131;
  assign n42133 = i_hbusreq6 & ~n42096;
  assign n42134 = ~n40554 & ~n41420;
  assign n42135 = ~controllable_hmaster1 & ~n42134;
  assign n42136 = ~n41419 & ~n42135;
  assign n42137 = ~i_hbusreq6 & ~n42136;
  assign n42138 = ~n42133 & ~n42137;
  assign n42139 = ~controllable_hgrant6 & ~n42138;
  assign n42140 = ~n42132 & ~n42139;
  assign n42141 = ~controllable_hmaster0 & ~n42140;
  assign n42142 = ~n42107 & ~n42141;
  assign n42143 = ~i_hlock8 & ~n42142;
  assign n42144 = ~n42125 & ~n42143;
  assign n42145 = ~i_hbusreq8 & ~n42144;
  assign n42146 = ~n42106 & ~n42145;
  assign n42147 = controllable_hmaster3 & ~n42146;
  assign n42148 = ~n41550 & ~n42147;
  assign n42149 = ~i_hbusreq7 & ~n42148;
  assign n42150 = ~n42105 & ~n42149;
  assign n42151 = ~n7924 & ~n42150;
  assign n42152 = controllable_hmaster0 & ~n41671;
  assign n42153 = n8217 & ~n13421;
  assign n42154 = ~n8217 & ~n17779;
  assign n42155 = ~n42153 & ~n42154;
  assign n42156 = controllable_hgrant6 & ~n42155;
  assign n42157 = n8378 & ~n13415;
  assign n42158 = ~n8378 & ~n17773;
  assign n42159 = ~n42157 & ~n42158;
  assign n42160 = controllable_hgrant5 & ~n42159;
  assign n42161 = controllable_hgrant4 & ~n41586;
  assign n42162 = ~controllable_hgrant4 & ~n41618;
  assign n42163 = ~n42161 & ~n42162;
  assign n42164 = ~controllable_hgrant5 & ~n42163;
  assign n42165 = ~n42160 & ~n42164;
  assign n42166 = ~controllable_hmaster2 & ~n42165;
  assign n42167 = ~n41579 & ~n42166;
  assign n42168 = ~controllable_hmaster1 & ~n42167;
  assign n42169 = ~n41578 & ~n42168;
  assign n42170 = ~controllable_hgrant6 & ~n42169;
  assign n42171 = ~n42156 & ~n42170;
  assign n42172 = ~controllable_hmaster0 & ~n42171;
  assign n42173 = ~n42152 & ~n42172;
  assign n42174 = i_hlock8 & ~n42173;
  assign n42175 = n8217 & ~n13442;
  assign n42176 = ~n8217 & ~n17797;
  assign n42177 = ~n42175 & ~n42176;
  assign n42178 = controllable_hgrant6 & ~n42177;
  assign n42179 = n8378 & ~n13436;
  assign n42180 = ~n8378 & ~n17791;
  assign n42181 = ~n42179 & ~n42180;
  assign n42182 = controllable_hgrant5 & ~n42181;
  assign n42183 = controllable_hgrant4 & ~n41590;
  assign n42184 = ~controllable_hgrant4 & ~n41632;
  assign n42185 = ~n42183 & ~n42184;
  assign n42186 = ~controllable_hgrant5 & ~n42185;
  assign n42187 = ~n42182 & ~n42186;
  assign n42188 = ~controllable_hmaster2 & ~n42187;
  assign n42189 = ~n41579 & ~n42188;
  assign n42190 = ~controllable_hmaster1 & ~n42189;
  assign n42191 = ~n41578 & ~n42190;
  assign n42192 = ~controllable_hgrant6 & ~n42191;
  assign n42193 = ~n42178 & ~n42192;
  assign n42194 = ~controllable_hmaster0 & ~n42193;
  assign n42195 = ~n42152 & ~n42194;
  assign n42196 = ~i_hlock8 & ~n42195;
  assign n42197 = ~n42174 & ~n42196;
  assign n42198 = controllable_hmaster3 & ~n42197;
  assign n42199 = ~n41736 & ~n42198;
  assign n42200 = i_hbusreq7 & ~n42199;
  assign n42201 = i_hbusreq8 & ~n42197;
  assign n42202 = controllable_hmaster0 & ~n41955;
  assign n42203 = i_hbusreq6 & ~n42155;
  assign n42204 = n8217 & ~n13565;
  assign n42205 = ~n8217 & ~n17854;
  assign n42206 = ~n42204 & ~n42205;
  assign n42207 = ~i_hbusreq6 & ~n42206;
  assign n42208 = ~n42203 & ~n42207;
  assign n42209 = controllable_hgrant6 & ~n42208;
  assign n42210 = i_hbusreq6 & ~n42169;
  assign n42211 = i_hbusreq5 & ~n42159;
  assign n42212 = n8378 & ~n13557;
  assign n42213 = ~n8378 & ~n17846;
  assign n42214 = ~n42212 & ~n42213;
  assign n42215 = ~i_hbusreq5 & ~n42214;
  assign n42216 = ~n42211 & ~n42215;
  assign n42217 = controllable_hgrant5 & ~n42216;
  assign n42218 = i_hbusreq5 & ~n42163;
  assign n42219 = i_hbusreq4 & ~n41586;
  assign n42220 = i_hbusreq9 & ~n41586;
  assign n42221 = ~i_hbusreq9 & ~n41797;
  assign n42222 = ~n42220 & ~n42221;
  assign n42223 = ~i_hbusreq4 & ~n42222;
  assign n42224 = ~n42219 & ~n42223;
  assign n42225 = controllable_hgrant4 & ~n42224;
  assign n42226 = i_hbusreq4 & ~n41618;
  assign n42227 = i_hbusreq9 & ~n41618;
  assign n42228 = ~i_hbusreq9 & ~n41859;
  assign n42229 = ~n42227 & ~n42228;
  assign n42230 = ~i_hbusreq4 & ~n42229;
  assign n42231 = ~n42226 & ~n42230;
  assign n42232 = ~controllable_hgrant4 & ~n42231;
  assign n42233 = ~n42225 & ~n42232;
  assign n42234 = ~i_hbusreq5 & ~n42233;
  assign n42235 = ~n42218 & ~n42234;
  assign n42236 = ~controllable_hgrant5 & ~n42235;
  assign n42237 = ~n42217 & ~n42236;
  assign n42238 = ~controllable_hmaster2 & ~n42237;
  assign n42239 = ~n41784 & ~n42238;
  assign n42240 = ~controllable_hmaster1 & ~n42239;
  assign n42241 = ~n41783 & ~n42240;
  assign n42242 = ~i_hbusreq6 & ~n42241;
  assign n42243 = ~n42210 & ~n42242;
  assign n42244 = ~controllable_hgrant6 & ~n42243;
  assign n42245 = ~n42209 & ~n42244;
  assign n42246 = ~controllable_hmaster0 & ~n42245;
  assign n42247 = ~n42202 & ~n42246;
  assign n42248 = i_hlock8 & ~n42247;
  assign n42249 = i_hbusreq6 & ~n42177;
  assign n42250 = n8217 & ~n13604;
  assign n42251 = ~n8217 & ~n17890;
  assign n42252 = ~n42250 & ~n42251;
  assign n42253 = ~i_hbusreq6 & ~n42252;
  assign n42254 = ~n42249 & ~n42253;
  assign n42255 = controllable_hgrant6 & ~n42254;
  assign n42256 = i_hbusreq6 & ~n42191;
  assign n42257 = i_hbusreq5 & ~n42181;
  assign n42258 = n8378 & ~n13596;
  assign n42259 = ~n8378 & ~n17882;
  assign n42260 = ~n42258 & ~n42259;
  assign n42261 = ~i_hbusreq5 & ~n42260;
  assign n42262 = ~n42257 & ~n42261;
  assign n42263 = controllable_hgrant5 & ~n42262;
  assign n42264 = i_hbusreq5 & ~n42185;
  assign n42265 = i_hbusreq4 & ~n41590;
  assign n42266 = i_hbusreq9 & ~n41590;
  assign n42267 = ~i_hbusreq9 & ~n41801;
  assign n42268 = ~n42266 & ~n42267;
  assign n42269 = ~i_hbusreq4 & ~n42268;
  assign n42270 = ~n42265 & ~n42269;
  assign n42271 = controllable_hgrant4 & ~n42270;
  assign n42272 = i_hbusreq4 & ~n41632;
  assign n42273 = i_hbusreq9 & ~n41632;
  assign n42274 = ~i_hbusreq9 & ~n41885;
  assign n42275 = ~n42273 & ~n42274;
  assign n42276 = ~i_hbusreq4 & ~n42275;
  assign n42277 = ~n42272 & ~n42276;
  assign n42278 = ~controllable_hgrant4 & ~n42277;
  assign n42279 = ~n42271 & ~n42278;
  assign n42280 = ~i_hbusreq5 & ~n42279;
  assign n42281 = ~n42264 & ~n42280;
  assign n42282 = ~controllable_hgrant5 & ~n42281;
  assign n42283 = ~n42263 & ~n42282;
  assign n42284 = ~controllable_hmaster2 & ~n42283;
  assign n42285 = ~n41784 & ~n42284;
  assign n42286 = ~controllable_hmaster1 & ~n42285;
  assign n42287 = ~n41783 & ~n42286;
  assign n42288 = ~i_hbusreq6 & ~n42287;
  assign n42289 = ~n42256 & ~n42288;
  assign n42290 = ~controllable_hgrant6 & ~n42289;
  assign n42291 = ~n42255 & ~n42290;
  assign n42292 = ~controllable_hmaster0 & ~n42291;
  assign n42293 = ~n42202 & ~n42292;
  assign n42294 = ~i_hlock8 & ~n42293;
  assign n42295 = ~n42248 & ~n42294;
  assign n42296 = ~i_hbusreq8 & ~n42295;
  assign n42297 = ~n42201 & ~n42296;
  assign n42298 = controllable_hmaster3 & ~n42297;
  assign n42299 = ~n42070 & ~n42298;
  assign n42300 = ~i_hbusreq7 & ~n42299;
  assign n42301 = ~n42200 & ~n42300;
  assign n42302 = n7924 & ~n42301;
  assign n42303 = ~n42151 & ~n42302;
  assign n42304 = n8214 & ~n42303;
  assign n42305 = ~n42076 & ~n42304;
  assign n42306 = ~n8202 & ~n42305;
  assign n42307 = controllable_hmaster3 & ~n41314;
  assign n42308 = n8217 & ~n9097;
  assign n42309 = ~n8217 & ~n17912;
  assign n42310 = ~n42308 & ~n42309;
  assign n42311 = controllable_hgrant6 & ~n42310;
  assign n42312 = ~n40579 & ~n41325;
  assign n42313 = controllable_hmaster1 & ~n42312;
  assign n42314 = ~n41343 & ~n42313;
  assign n42315 = ~controllable_hgrant6 & ~n42314;
  assign n42316 = ~n42311 & ~n42315;
  assign n42317 = controllable_hmaster0 & ~n42316;
  assign n42318 = ~n41376 & ~n42317;
  assign n42319 = ~controllable_hmaster3 & ~n42318;
  assign n42320 = ~n42307 & ~n42319;
  assign n42321 = i_hlock7 & ~n42320;
  assign n42322 = n8217 & ~n9106;
  assign n42323 = ~n8217 & ~n17922;
  assign n42324 = ~n42322 & ~n42323;
  assign n42325 = controllable_hgrant6 & ~n42324;
  assign n42326 = ~n40594 & ~n41325;
  assign n42327 = controllable_hmaster1 & ~n42326;
  assign n42328 = ~n41343 & ~n42327;
  assign n42329 = ~controllable_hgrant6 & ~n42328;
  assign n42330 = ~n42325 & ~n42329;
  assign n42331 = controllable_hmaster0 & ~n42330;
  assign n42332 = ~n41376 & ~n42331;
  assign n42333 = ~controllable_hmaster3 & ~n42332;
  assign n42334 = ~n42307 & ~n42333;
  assign n42335 = ~i_hlock7 & ~n42334;
  assign n42336 = ~n42321 & ~n42335;
  assign n42337 = i_hbusreq7 & ~n42336;
  assign n42338 = i_hbusreq8 & ~n41314;
  assign n42339 = ~i_hbusreq8 & ~n41436;
  assign n42340 = ~n42338 & ~n42339;
  assign n42341 = controllable_hmaster3 & ~n42340;
  assign n42342 = i_hbusreq8 & ~n42318;
  assign n42343 = i_hbusreq6 & ~n42310;
  assign n42344 = n8217 & ~n9123;
  assign n42345 = ~n8217 & ~n17936;
  assign n42346 = ~n42344 & ~n42345;
  assign n42347 = ~i_hbusreq6 & ~n42346;
  assign n42348 = ~n42343 & ~n42347;
  assign n42349 = controllable_hgrant6 & ~n42348;
  assign n42350 = i_hbusreq6 & ~n42314;
  assign n42351 = ~n40616 & ~n41460;
  assign n42352 = controllable_hmaster1 & ~n42351;
  assign n42353 = ~n41490 & ~n42352;
  assign n42354 = ~i_hbusreq6 & ~n42353;
  assign n42355 = ~n42350 & ~n42354;
  assign n42356 = ~controllable_hgrant6 & ~n42355;
  assign n42357 = ~n42349 & ~n42356;
  assign n42358 = controllable_hmaster0 & ~n42357;
  assign n42359 = ~n41546 & ~n42358;
  assign n42360 = ~i_hbusreq8 & ~n42359;
  assign n42361 = ~n42342 & ~n42360;
  assign n42362 = ~controllable_hmaster3 & ~n42361;
  assign n42363 = ~n42341 & ~n42362;
  assign n42364 = i_hlock7 & ~n42363;
  assign n42365 = i_hbusreq8 & ~n42332;
  assign n42366 = i_hbusreq6 & ~n42324;
  assign n42367 = n8217 & ~n9138;
  assign n42368 = ~n8217 & ~n17952;
  assign n42369 = ~n42367 & ~n42368;
  assign n42370 = ~i_hbusreq6 & ~n42369;
  assign n42371 = ~n42366 & ~n42370;
  assign n42372 = controllable_hgrant6 & ~n42371;
  assign n42373 = i_hbusreq6 & ~n42328;
  assign n42374 = ~n40640 & ~n41460;
  assign n42375 = controllable_hmaster1 & ~n42374;
  assign n42376 = ~n41490 & ~n42375;
  assign n42377 = ~i_hbusreq6 & ~n42376;
  assign n42378 = ~n42373 & ~n42377;
  assign n42379 = ~controllable_hgrant6 & ~n42378;
  assign n42380 = ~n42372 & ~n42379;
  assign n42381 = controllable_hmaster0 & ~n42380;
  assign n42382 = ~n41546 & ~n42381;
  assign n42383 = ~i_hbusreq8 & ~n42382;
  assign n42384 = ~n42365 & ~n42383;
  assign n42385 = ~controllable_hmaster3 & ~n42384;
  assign n42386 = ~n42341 & ~n42385;
  assign n42387 = ~i_hlock7 & ~n42386;
  assign n42388 = ~n42364 & ~n42387;
  assign n42389 = ~i_hbusreq7 & ~n42388;
  assign n42390 = ~n42337 & ~n42389;
  assign n42391 = ~n7924 & ~n42390;
  assign n42392 = controllable_hmaster3 & ~n41671;
  assign n42393 = n8217 & ~n13678;
  assign n42394 = ~n8217 & ~n17971;
  assign n42395 = ~n42393 & ~n42394;
  assign n42396 = controllable_hgrant6 & ~n42395;
  assign n42397 = controllable_hmaster2 & ~n42165;
  assign n42398 = ~n41683 & ~n42397;
  assign n42399 = controllable_hmaster1 & ~n42398;
  assign n42400 = ~n41699 & ~n42399;
  assign n42401 = ~controllable_hgrant6 & ~n42400;
  assign n42402 = ~n42396 & ~n42401;
  assign n42403 = controllable_hmaster0 & ~n42402;
  assign n42404 = ~n41734 & ~n42403;
  assign n42405 = ~controllable_hmaster3 & ~n42404;
  assign n42406 = ~n42392 & ~n42405;
  assign n42407 = i_hlock7 & ~n42406;
  assign n42408 = n8217 & ~n13691;
  assign n42409 = ~n8217 & ~n17982;
  assign n42410 = ~n42408 & ~n42409;
  assign n42411 = controllable_hgrant6 & ~n42410;
  assign n42412 = controllable_hmaster2 & ~n42187;
  assign n42413 = ~n41683 & ~n42412;
  assign n42414 = controllable_hmaster1 & ~n42413;
  assign n42415 = ~n41699 & ~n42414;
  assign n42416 = ~controllable_hgrant6 & ~n42415;
  assign n42417 = ~n42411 & ~n42416;
  assign n42418 = controllable_hmaster0 & ~n42417;
  assign n42419 = ~n41734 & ~n42418;
  assign n42420 = ~controllable_hmaster3 & ~n42419;
  assign n42421 = ~n42392 & ~n42420;
  assign n42422 = ~i_hlock7 & ~n42421;
  assign n42423 = ~n42407 & ~n42422;
  assign n42424 = i_hbusreq7 & ~n42423;
  assign n42425 = i_hbusreq8 & ~n41671;
  assign n42426 = ~i_hbusreq8 & ~n41955;
  assign n42427 = ~n42425 & ~n42426;
  assign n42428 = controllable_hmaster3 & ~n42427;
  assign n42429 = i_hbusreq8 & ~n42404;
  assign n42430 = i_hbusreq6 & ~n42395;
  assign n42431 = n8217 & ~n13722;
  assign n42432 = ~n8217 & ~n17997;
  assign n42433 = ~n42431 & ~n42432;
  assign n42434 = ~i_hbusreq6 & ~n42433;
  assign n42435 = ~n42430 & ~n42434;
  assign n42436 = controllable_hgrant6 & ~n42435;
  assign n42437 = i_hbusreq6 & ~n42400;
  assign n42438 = controllable_hmaster2 & ~n42237;
  assign n42439 = ~n41980 & ~n42438;
  assign n42440 = controllable_hmaster1 & ~n42439;
  assign n42441 = ~n42008 & ~n42440;
  assign n42442 = ~i_hbusreq6 & ~n42441;
  assign n42443 = ~n42437 & ~n42442;
  assign n42444 = ~controllable_hgrant6 & ~n42443;
  assign n42445 = ~n42436 & ~n42444;
  assign n42446 = controllable_hmaster0 & ~n42445;
  assign n42447 = ~n42066 & ~n42446;
  assign n42448 = ~i_hbusreq8 & ~n42447;
  assign n42449 = ~n42429 & ~n42448;
  assign n42450 = ~controllable_hmaster3 & ~n42449;
  assign n42451 = ~n42428 & ~n42450;
  assign n42452 = i_hlock7 & ~n42451;
  assign n42453 = i_hbusreq8 & ~n42419;
  assign n42454 = i_hbusreq6 & ~n42410;
  assign n42455 = n8217 & ~n13741;
  assign n42456 = ~n8217 & ~n18014;
  assign n42457 = ~n42455 & ~n42456;
  assign n42458 = ~i_hbusreq6 & ~n42457;
  assign n42459 = ~n42454 & ~n42458;
  assign n42460 = controllable_hgrant6 & ~n42459;
  assign n42461 = i_hbusreq6 & ~n42415;
  assign n42462 = controllable_hmaster2 & ~n42283;
  assign n42463 = ~n41980 & ~n42462;
  assign n42464 = controllable_hmaster1 & ~n42463;
  assign n42465 = ~n42008 & ~n42464;
  assign n42466 = ~i_hbusreq6 & ~n42465;
  assign n42467 = ~n42461 & ~n42466;
  assign n42468 = ~controllable_hgrant6 & ~n42467;
  assign n42469 = ~n42460 & ~n42468;
  assign n42470 = controllable_hmaster0 & ~n42469;
  assign n42471 = ~n42066 & ~n42470;
  assign n42472 = ~i_hbusreq8 & ~n42471;
  assign n42473 = ~n42453 & ~n42472;
  assign n42474 = ~controllable_hmaster3 & ~n42473;
  assign n42475 = ~n42428 & ~n42474;
  assign n42476 = ~i_hlock7 & ~n42475;
  assign n42477 = ~n42452 & ~n42476;
  assign n42478 = ~i_hbusreq7 & ~n42477;
  assign n42479 = ~n42424 & ~n42478;
  assign n42480 = n7924 & ~n42479;
  assign n42481 = ~n42391 & ~n42480;
  assign n42482 = ~n8214 & ~n42481;
  assign n42483 = n8217 & ~n8991;
  assign n42484 = ~n8217 & ~n17343;
  assign n42485 = ~n42483 & ~n42484;
  assign n42486 = controllable_hgrant6 & ~n42485;
  assign n42487 = ~n41313 & ~n42486;
  assign n42488 = controllable_hmaster3 & ~n42487;
  assign n42489 = n8217 & ~n8987;
  assign n42490 = ~n8217 & ~n17339;
  assign n42491 = ~n42489 & ~n42490;
  assign n42492 = controllable_hgrant6 & ~n42491;
  assign n42493 = ~n41345 & ~n42492;
  assign n42494 = controllable_hmaster0 & ~n42493;
  assign n42495 = n8217 & ~n27032;
  assign n42496 = ~n8217 & ~n29424;
  assign n42497 = ~n42495 & ~n42496;
  assign n42498 = i_hlock6 & ~n42497;
  assign n42499 = n8217 & ~n27042;
  assign n42500 = ~n8217 & ~n29435;
  assign n42501 = ~n42499 & ~n42500;
  assign n42502 = ~i_hlock6 & ~n42501;
  assign n42503 = ~n42498 & ~n42502;
  assign n42504 = controllable_hgrant6 & ~n42503;
  assign n42505 = ~n40579 & ~n41362;
  assign n42506 = controllable_hmaster1 & ~n42505;
  assign n42507 = ~n41372 & ~n42506;
  assign n42508 = i_hlock6 & ~n42507;
  assign n42509 = ~n40594 & ~n41362;
  assign n42510 = controllable_hmaster1 & ~n42509;
  assign n42511 = ~n41372 & ~n42510;
  assign n42512 = ~i_hlock6 & ~n42511;
  assign n42513 = ~n42508 & ~n42512;
  assign n42514 = ~controllable_hgrant6 & ~n42513;
  assign n42515 = ~n42504 & ~n42514;
  assign n42516 = ~controllable_hmaster0 & ~n42515;
  assign n42517 = ~n42494 & ~n42516;
  assign n42518 = ~controllable_hmaster3 & ~n42517;
  assign n42519 = ~n42488 & ~n42518;
  assign n42520 = i_hbusreq7 & ~n42519;
  assign n42521 = i_hbusreq8 & ~n42487;
  assign n42522 = i_hbusreq6 & ~n42485;
  assign n42523 = n8217 & ~n9027;
  assign n42524 = ~n8217 & ~n17438;
  assign n42525 = ~n42523 & ~n42524;
  assign n42526 = ~i_hbusreq6 & ~n42525;
  assign n42527 = ~n42522 & ~n42526;
  assign n42528 = controllable_hgrant6 & ~n42527;
  assign n42529 = ~n41435 & ~n42528;
  assign n42530 = ~i_hbusreq8 & ~n42529;
  assign n42531 = ~n42521 & ~n42530;
  assign n42532 = controllable_hmaster3 & ~n42531;
  assign n42533 = i_hbusreq8 & ~n42517;
  assign n42534 = i_hbusreq6 & ~n42491;
  assign n42535 = n8217 & ~n9023;
  assign n42536 = ~n8217 & ~n17434;
  assign n42537 = ~n42535 & ~n42536;
  assign n42538 = ~i_hbusreq6 & ~n42537;
  assign n42539 = ~n42534 & ~n42538;
  assign n42540 = controllable_hgrant6 & ~n42539;
  assign n42541 = ~n41494 & ~n42540;
  assign n42542 = controllable_hmaster0 & ~n42541;
  assign n42543 = i_hbusreq6 & ~n42503;
  assign n42544 = n8217 & ~n27056;
  assign n42545 = ~n8217 & ~n29454;
  assign n42546 = ~n42544 & ~n42545;
  assign n42547 = i_hlock6 & ~n42546;
  assign n42548 = n8217 & ~n27072;
  assign n42549 = ~n8217 & ~n29471;
  assign n42550 = ~n42548 & ~n42549;
  assign n42551 = ~i_hlock6 & ~n42550;
  assign n42552 = ~n42547 & ~n42551;
  assign n42553 = ~i_hbusreq6 & ~n42552;
  assign n42554 = ~n42543 & ~n42553;
  assign n42555 = controllable_hgrant6 & ~n42554;
  assign n42556 = i_hbusreq6 & ~n42513;
  assign n42557 = ~n40616 & ~n41527;
  assign n42558 = controllable_hmaster1 & ~n42557;
  assign n42559 = ~n41540 & ~n42558;
  assign n42560 = i_hlock6 & ~n42559;
  assign n42561 = ~n40640 & ~n41527;
  assign n42562 = controllable_hmaster1 & ~n42561;
  assign n42563 = ~n41540 & ~n42562;
  assign n42564 = ~i_hlock6 & ~n42563;
  assign n42565 = ~n42560 & ~n42564;
  assign n42566 = ~i_hbusreq6 & ~n42565;
  assign n42567 = ~n42556 & ~n42566;
  assign n42568 = ~controllable_hgrant6 & ~n42567;
  assign n42569 = ~n42555 & ~n42568;
  assign n42570 = ~controllable_hmaster0 & ~n42569;
  assign n42571 = ~n42542 & ~n42570;
  assign n42572 = ~i_hbusreq8 & ~n42571;
  assign n42573 = ~n42533 & ~n42572;
  assign n42574 = ~controllable_hmaster3 & ~n42573;
  assign n42575 = ~n42532 & ~n42574;
  assign n42576 = ~i_hbusreq7 & ~n42575;
  assign n42577 = ~n42520 & ~n42576;
  assign n42578 = ~n7924 & ~n42577;
  assign n42579 = n8217 & ~n13192;
  assign n42580 = ~n8217 & ~n29500;
  assign n42581 = ~n42579 & ~n42580;
  assign n42582 = i_hlock6 & ~n42581;
  assign n42583 = ~n8217 & ~n29531;
  assign n42584 = ~n42579 & ~n42583;
  assign n42585 = ~i_hlock6 & ~n42584;
  assign n42586 = ~n42582 & ~n42585;
  assign n42587 = controllable_hgrant6 & ~n42586;
  assign n42588 = ~n41670 & ~n42587;
  assign n42589 = controllable_hmaster3 & ~n42588;
  assign n42590 = n8217 & ~n13188;
  assign n42591 = ~n8217 & ~n29496;
  assign n42592 = ~n42590 & ~n42591;
  assign n42593 = i_hlock6 & ~n42592;
  assign n42594 = ~n8217 & ~n29527;
  assign n42595 = ~n42590 & ~n42594;
  assign n42596 = ~i_hlock6 & ~n42595;
  assign n42597 = ~n42593 & ~n42596;
  assign n42598 = controllable_hgrant6 & ~n42597;
  assign n42599 = ~n41701 & ~n42598;
  assign n42600 = controllable_hmaster0 & ~n42599;
  assign n42601 = n8217 & ~n27091;
  assign n42602 = ~n8217 & ~n29507;
  assign n42603 = ~n42601 & ~n42602;
  assign n42604 = i_hlock6 & ~n42603;
  assign n42605 = n8217 & ~n27101;
  assign n42606 = ~n8217 & ~n29538;
  assign n42607 = ~n42605 & ~n42606;
  assign n42608 = ~i_hlock6 & ~n42607;
  assign n42609 = ~n42604 & ~n42608;
  assign n42610 = controllable_hgrant6 & ~n42609;
  assign n42611 = ~n41721 & ~n42397;
  assign n42612 = controllable_hmaster1 & ~n42611;
  assign n42613 = ~n41730 & ~n42612;
  assign n42614 = i_hlock6 & ~n42613;
  assign n42615 = ~n41721 & ~n42412;
  assign n42616 = controllable_hmaster1 & ~n42615;
  assign n42617 = ~n41730 & ~n42616;
  assign n42618 = ~i_hlock6 & ~n42617;
  assign n42619 = ~n42614 & ~n42618;
  assign n42620 = ~controllable_hgrant6 & ~n42619;
  assign n42621 = ~n42610 & ~n42620;
  assign n42622 = ~controllable_hmaster0 & ~n42621;
  assign n42623 = ~n42600 & ~n42622;
  assign n42624 = ~controllable_hmaster3 & ~n42623;
  assign n42625 = ~n42589 & ~n42624;
  assign n42626 = i_hbusreq7 & ~n42625;
  assign n42627 = i_hbusreq8 & ~n42588;
  assign n42628 = i_hbusreq6 & ~n42586;
  assign n42629 = n8217 & ~n13287;
  assign n42630 = ~n8217 & ~n29584;
  assign n42631 = ~n42629 & ~n42630;
  assign n42632 = i_hlock6 & ~n42631;
  assign n42633 = ~n8217 & ~n29648;
  assign n42634 = ~n42629 & ~n42633;
  assign n42635 = ~i_hlock6 & ~n42634;
  assign n42636 = ~n42632 & ~n42635;
  assign n42637 = ~i_hbusreq6 & ~n42636;
  assign n42638 = ~n42628 & ~n42637;
  assign n42639 = controllable_hgrant6 & ~n42638;
  assign n42640 = ~n41954 & ~n42639;
  assign n42641 = ~i_hbusreq8 & ~n42640;
  assign n42642 = ~n42627 & ~n42641;
  assign n42643 = controllable_hmaster3 & ~n42642;
  assign n42644 = i_hbusreq8 & ~n42623;
  assign n42645 = i_hbusreq6 & ~n42597;
  assign n42646 = n8217 & ~n13283;
  assign n42647 = ~n8217 & ~n29580;
  assign n42648 = ~n42646 & ~n42647;
  assign n42649 = i_hlock6 & ~n42648;
  assign n42650 = ~n8217 & ~n29644;
  assign n42651 = ~n42646 & ~n42650;
  assign n42652 = ~i_hlock6 & ~n42651;
  assign n42653 = ~n42649 & ~n42652;
  assign n42654 = ~i_hbusreq6 & ~n42653;
  assign n42655 = ~n42645 & ~n42654;
  assign n42656 = controllable_hgrant6 & ~n42655;
  assign n42657 = ~n42012 & ~n42656;
  assign n42658 = controllable_hmaster0 & ~n42657;
  assign n42659 = i_hbusreq6 & ~n42609;
  assign n42660 = n8217 & ~n27120;
  assign n42661 = ~n8217 & ~n29597;
  assign n42662 = ~n42660 & ~n42661;
  assign n42663 = i_hlock6 & ~n42662;
  assign n42664 = n8217 & ~n27137;
  assign n42665 = ~n8217 & ~n29661;
  assign n42666 = ~n42664 & ~n42665;
  assign n42667 = ~i_hlock6 & ~n42666;
  assign n42668 = ~n42663 & ~n42667;
  assign n42669 = ~i_hbusreq6 & ~n42668;
  assign n42670 = ~n42659 & ~n42669;
  assign n42671 = controllable_hgrant6 & ~n42670;
  assign n42672 = i_hbusreq6 & ~n42619;
  assign n42673 = ~n42048 & ~n42438;
  assign n42674 = controllable_hmaster1 & ~n42673;
  assign n42675 = ~n42060 & ~n42674;
  assign n42676 = i_hlock6 & ~n42675;
  assign n42677 = ~n42048 & ~n42462;
  assign n42678 = controllable_hmaster1 & ~n42677;
  assign n42679 = ~n42060 & ~n42678;
  assign n42680 = ~i_hlock6 & ~n42679;
  assign n42681 = ~n42676 & ~n42680;
  assign n42682 = ~i_hbusreq6 & ~n42681;
  assign n42683 = ~n42672 & ~n42682;
  assign n42684 = ~controllable_hgrant6 & ~n42683;
  assign n42685 = ~n42671 & ~n42684;
  assign n42686 = ~controllable_hmaster0 & ~n42685;
  assign n42687 = ~n42658 & ~n42686;
  assign n42688 = ~i_hbusreq8 & ~n42687;
  assign n42689 = ~n42644 & ~n42688;
  assign n42690 = ~controllable_hmaster3 & ~n42689;
  assign n42691 = ~n42643 & ~n42690;
  assign n42692 = ~i_hbusreq7 & ~n42691;
  assign n42693 = ~n42626 & ~n42692;
  assign n42694 = n7924 & ~n42693;
  assign n42695 = ~n42578 & ~n42694;
  assign n42696 = n8214 & ~n42695;
  assign n42697 = ~n42482 & ~n42696;
  assign n42698 = n8202 & ~n42697;
  assign n42699 = ~n42306 & ~n42698;
  assign n42700 = n7920 & ~n42699;
  assign n42701 = ~n40788 & ~n42700;
  assign n42702 = n7728 & ~n42701;
  assign n42703 = ~n8217 & ~n29721;
  assign n42704 = ~n41284 & ~n42703;
  assign n42705 = controllable_hgrant6 & ~n42704;
  assign n42706 = ~n7735 & n8378;
  assign n42707 = ~n8378 & ~n19178;
  assign n42708 = ~n42706 & ~n42707;
  assign n42709 = controllable_hgrant5 & ~n42708;
  assign n42710 = ~n7735 & n8426;
  assign n42711 = ~n8426 & ~n19176;
  assign n42712 = ~n42710 & ~n42711;
  assign n42713 = controllable_hgrant4 & ~n42712;
  assign n42714 = ~n7735 & n8365;
  assign n42715 = ~n8365 & ~n19174;
  assign n42716 = ~n42714 & ~n42715;
  assign n42717 = controllable_hgrant3 & ~n42716;
  assign n42718 = ~n7735 & n8389;
  assign n42719 = ~n8389 & ~n16725;
  assign n42720 = ~n42718 & ~n42719;
  assign n42721 = controllable_hgrant1 & ~n42720;
  assign n42722 = ~n16349 & ~n40219;
  assign n42723 = ~n7928 & ~n42722;
  assign n42724 = ~n7936 & ~n40219;
  assign n42725 = ~n7733 & ~n42724;
  assign n42726 = n7733 & ~n42722;
  assign n42727 = ~n42725 & ~n42726;
  assign n42728 = n7928 & ~n42727;
  assign n42729 = ~n42723 & ~n42728;
  assign n42730 = ~controllable_hgrant1 & ~n42729;
  assign n42731 = ~n42721 & ~n42730;
  assign n42732 = ~controllable_hgrant3 & ~n42731;
  assign n42733 = ~n42717 & ~n42732;
  assign n42734 = ~controllable_hgrant4 & ~n42733;
  assign n42735 = ~n42713 & ~n42734;
  assign n42736 = ~controllable_hgrant5 & ~n42735;
  assign n42737 = ~n42709 & ~n42736;
  assign n42738 = controllable_hmaster1 & ~n42737;
  assign n42739 = controllable_hmaster2 & ~n42737;
  assign n42740 = ~n40256 & ~n42739;
  assign n42741 = ~controllable_hmaster1 & ~n42740;
  assign n42742 = ~n42738 & ~n42741;
  assign n42743 = ~controllable_hgrant6 & ~n42742;
  assign n42744 = ~n42705 & ~n42743;
  assign n42745 = controllable_hmaster0 & ~n42744;
  assign n42746 = ~n8217 & ~n20271;
  assign n42747 = ~n42078 & ~n42746;
  assign n42748 = controllable_hgrant6 & ~n42747;
  assign n42749 = ~n8378 & ~n19233;
  assign n42750 = ~n40428 & ~n42749;
  assign n42751 = controllable_hgrant5 & ~n42750;
  assign n42752 = ~n8426 & ~n19231;
  assign n42753 = ~n40197 & ~n42752;
  assign n42754 = controllable_hgrant4 & ~n42753;
  assign n42755 = ~n8365 & ~n19229;
  assign n42756 = ~n40207 & ~n42755;
  assign n42757 = controllable_hgrant3 & ~n42756;
  assign n42758 = ~n8389 & ~n19227;
  assign n42759 = ~n40211 & ~n42758;
  assign n42760 = controllable_hgrant1 & ~n42759;
  assign n42761 = ~n16724 & ~n40219;
  assign n42762 = n7928 & ~n42761;
  assign n42763 = ~n8221 & ~n42762;
  assign n42764 = ~controllable_hgrant1 & ~n42763;
  assign n42765 = ~n42760 & ~n42764;
  assign n42766 = ~controllable_hgrant3 & ~n42765;
  assign n42767 = ~n42757 & ~n42766;
  assign n42768 = ~controllable_hgrant4 & ~n42767;
  assign n42769 = ~n42754 & ~n42768;
  assign n42770 = ~controllable_hgrant5 & ~n42769;
  assign n42771 = ~n42751 & ~n42770;
  assign n42772 = ~controllable_hmaster2 & ~n42771;
  assign n42773 = ~n42739 & ~n42772;
  assign n42774 = ~controllable_hmaster1 & ~n42773;
  assign n42775 = ~n42738 & ~n42774;
  assign n42776 = ~controllable_hgrant6 & ~n42775;
  assign n42777 = ~n42748 & ~n42776;
  assign n42778 = ~controllable_hmaster0 & ~n42777;
  assign n42779 = ~n42745 & ~n42778;
  assign n42780 = i_hlock8 & ~n42779;
  assign n42781 = ~n8217 & ~n20280;
  assign n42782 = ~n42090 & ~n42781;
  assign n42783 = controllable_hgrant6 & ~n42782;
  assign n42784 = ~n8378 & ~n19256;
  assign n42785 = ~n40450 & ~n42784;
  assign n42786 = controllable_hgrant5 & ~n42785;
  assign n42787 = ~n8426 & ~n19254;
  assign n42788 = ~n40201 & ~n42787;
  assign n42789 = controllable_hgrant4 & ~n42788;
  assign n42790 = ~n8365 & ~n19240;
  assign n42791 = ~n40237 & ~n42790;
  assign n42792 = controllable_hgrant3 & ~n42791;
  assign n42793 = ~n8389 & ~n19238;
  assign n42794 = ~n40241 & ~n42793;
  assign n42795 = controllable_hgrant1 & ~n42794;
  assign n42796 = ~n8235 & ~n42762;
  assign n42797 = ~controllable_hgrant1 & ~n42796;
  assign n42798 = ~n42795 & ~n42797;
  assign n42799 = ~controllable_hgrant3 & ~n42798;
  assign n42800 = ~n42792 & ~n42799;
  assign n42801 = ~controllable_hgrant4 & ~n42800;
  assign n42802 = ~n42789 & ~n42801;
  assign n42803 = ~controllable_hgrant5 & ~n42802;
  assign n42804 = ~n42786 & ~n42803;
  assign n42805 = ~controllable_hmaster2 & ~n42804;
  assign n42806 = ~n42739 & ~n42805;
  assign n42807 = ~controllable_hmaster1 & ~n42806;
  assign n42808 = ~n42738 & ~n42807;
  assign n42809 = ~controllable_hgrant6 & ~n42808;
  assign n42810 = ~n42783 & ~n42809;
  assign n42811 = ~controllable_hmaster0 & ~n42810;
  assign n42812 = ~n42745 & ~n42811;
  assign n42813 = ~i_hlock8 & ~n42812;
  assign n42814 = ~n42780 & ~n42813;
  assign n42815 = controllable_hmaster3 & ~n42814;
  assign n42816 = n8217 & ~n9206;
  assign n42817 = ~n8217 & ~n19276;
  assign n42818 = ~n42816 & ~n42817;
  assign n42819 = controllable_hgrant6 & ~n42818;
  assign n42820 = controllable_hmaster2 & ~n42771;
  assign n42821 = n8378 & ~n9192;
  assign n42822 = ~n8378 & ~n19246;
  assign n42823 = ~n42821 & ~n42822;
  assign n42824 = controllable_hgrant5 & ~n42823;
  assign n42825 = n8426 & ~n9192;
  assign n42826 = ~n8426 & ~n19244;
  assign n42827 = ~n42825 & ~n42826;
  assign n42828 = controllable_hgrant4 & ~n42827;
  assign n42829 = n8365 & ~n12633;
  assign n42830 = ~n8365 & ~n19186;
  assign n42831 = ~n42829 & ~n42830;
  assign n42832 = i_hlock3 & ~n42831;
  assign n42833 = n8365 & ~n12651;
  assign n42834 = ~n8365 & ~n19192;
  assign n42835 = ~n42833 & ~n42834;
  assign n42836 = ~i_hlock3 & ~n42835;
  assign n42837 = ~n42832 & ~n42836;
  assign n42838 = controllable_hgrant3 & ~n42837;
  assign n42839 = i_hlock3 & ~n42765;
  assign n42840 = ~i_hlock3 & ~n42798;
  assign n42841 = ~n42839 & ~n42840;
  assign n42842 = ~controllable_hgrant3 & ~n42841;
  assign n42843 = ~n42838 & ~n42842;
  assign n42844 = ~controllable_hgrant4 & ~n42843;
  assign n42845 = ~n42828 & ~n42844;
  assign n42846 = ~controllable_hgrant5 & ~n42845;
  assign n42847 = ~n42824 & ~n42846;
  assign n42848 = ~controllable_hmaster2 & ~n42847;
  assign n42849 = ~n42820 & ~n42848;
  assign n42850 = controllable_hmaster1 & ~n42849;
  assign n42851 = n8378 & ~n26638;
  assign n42852 = ~n8378 & ~n29732;
  assign n42853 = ~n42851 & ~n42852;
  assign n42854 = i_hlock5 & ~n42853;
  assign n42855 = n8378 & ~n26653;
  assign n42856 = ~n8378 & ~n29747;
  assign n42857 = ~n42855 & ~n42856;
  assign n42858 = ~i_hlock5 & ~n42857;
  assign n42859 = ~n42854 & ~n42858;
  assign n42860 = controllable_hgrant5 & ~n42859;
  assign n42861 = i_hlock5 & ~n42769;
  assign n42862 = ~i_hlock5 & ~n42802;
  assign n42863 = ~n42861 & ~n42862;
  assign n42864 = ~controllable_hgrant5 & ~n42863;
  assign n42865 = ~n42860 & ~n42864;
  assign n42866 = controllable_hmaster2 & ~n42865;
  assign n42867 = n8378 & ~n9202;
  assign n42868 = ~n8378 & ~n19270;
  assign n42869 = ~n42867 & ~n42868;
  assign n42870 = controllable_hgrant5 & ~n42869;
  assign n42871 = n8426 & ~n9202;
  assign n42872 = ~n8426 & ~n19268;
  assign n42873 = ~n42871 & ~n42872;
  assign n42874 = controllable_hgrant4 & ~n42873;
  assign n42875 = n8365 & ~n9202;
  assign n42876 = ~n8365 & ~n19266;
  assign n42877 = ~n42875 & ~n42876;
  assign n42878 = controllable_hgrant3 & ~n42877;
  assign n42879 = n8389 & ~n12631;
  assign n42880 = ~n8389 & ~n19184;
  assign n42881 = ~n42879 & ~n42880;
  assign n42882 = i_hlock1 & ~n42881;
  assign n42883 = n8389 & ~n12649;
  assign n42884 = ~n8389 & ~n19190;
  assign n42885 = ~n42883 & ~n42884;
  assign n42886 = ~i_hlock1 & ~n42885;
  assign n42887 = ~n42882 & ~n42886;
  assign n42888 = controllable_hgrant1 & ~n42887;
  assign n42889 = i_hlock1 & ~n42763;
  assign n42890 = ~i_hlock1 & ~n42796;
  assign n42891 = ~n42889 & ~n42890;
  assign n42892 = ~controllable_hgrant1 & ~n42891;
  assign n42893 = ~n42888 & ~n42892;
  assign n42894 = ~controllable_hgrant3 & ~n42893;
  assign n42895 = ~n42878 & ~n42894;
  assign n42896 = ~controllable_hgrant4 & ~n42895;
  assign n42897 = ~n42874 & ~n42896;
  assign n42898 = ~controllable_hgrant5 & ~n42897;
  assign n42899 = ~n42870 & ~n42898;
  assign n42900 = ~controllable_hmaster2 & ~n42899;
  assign n42901 = ~n42866 & ~n42900;
  assign n42902 = ~controllable_hmaster1 & ~n42901;
  assign n42903 = ~n42850 & ~n42902;
  assign n42904 = ~controllable_hgrant6 & ~n42903;
  assign n42905 = ~n42819 & ~n42904;
  assign n42906 = controllable_hmaster0 & ~n42905;
  assign n42907 = ~n9215 & ~n26641;
  assign n42908 = controllable_hmaster1 & ~n42907;
  assign n42909 = ~n9225 & ~n42908;
  assign n42910 = n8217 & ~n42909;
  assign n42911 = ~n19289 & ~n29735;
  assign n42912 = controllable_hmaster1 & ~n42911;
  assign n42913 = ~n19311 & ~n42912;
  assign n42914 = ~n8217 & ~n42913;
  assign n42915 = ~n42910 & ~n42914;
  assign n42916 = i_hlock6 & ~n42915;
  assign n42917 = ~n9215 & ~n26656;
  assign n42918 = controllable_hmaster1 & ~n42917;
  assign n42919 = ~n9225 & ~n42918;
  assign n42920 = n8217 & ~n42919;
  assign n42921 = ~n19289 & ~n29750;
  assign n42922 = controllable_hmaster1 & ~n42921;
  assign n42923 = ~n19311 & ~n42922;
  assign n42924 = ~n8217 & ~n42923;
  assign n42925 = ~n42920 & ~n42924;
  assign n42926 = ~i_hlock6 & ~n42925;
  assign n42927 = ~n42916 & ~n42926;
  assign n42928 = controllable_hgrant6 & ~n42927;
  assign n42929 = n8378 & ~n9214;
  assign n42930 = ~n8378 & ~n19286;
  assign n42931 = ~n42929 & ~n42930;
  assign n42932 = controllable_hgrant5 & ~n42931;
  assign n42933 = n8426 & ~n9214;
  assign n42934 = ~n8426 & ~n19284;
  assign n42935 = ~n42933 & ~n42934;
  assign n42936 = controllable_hgrant4 & ~n42935;
  assign n42937 = n8365 & ~n9214;
  assign n42938 = ~n8365 & ~n19282;
  assign n42939 = ~n42937 & ~n42938;
  assign n42940 = controllable_hgrant3 & ~n42939;
  assign n42941 = n8389 & ~n9214;
  assign n42942 = ~n8389 & ~n19280;
  assign n42943 = ~n42941 & ~n42942;
  assign n42944 = controllable_hgrant1 & ~n42943;
  assign n42945 = controllable_hmastlock & n39846;
  assign n42946 = controllable_hmastlock & ~n42945;
  assign n42947 = controllable_locked & ~n42946;
  assign n42948 = ~n7818 & ~n39848;
  assign n42949 = ~controllable_locked & ~n42948;
  assign n42950 = ~n42947 & ~n42949;
  assign n42951 = i_hlock2 & ~n42950;
  assign n42952 = ~n8231 & ~n39853;
  assign n42953 = controllable_locked & ~n42952;
  assign n42954 = ~controllable_hmastlock & n39846;
  assign n42955 = ~controllable_hmastlock & ~n42954;
  assign n42956 = ~controllable_locked & ~n42955;
  assign n42957 = ~n42953 & ~n42956;
  assign n42958 = ~i_hlock2 & ~n42957;
  assign n42959 = ~n42951 & ~n42958;
  assign n42960 = controllable_hgrant2 & ~n42959;
  assign n42961 = ~controllable_hgrant2 & ~n9210;
  assign n42962 = ~n42960 & ~n42961;
  assign n42963 = ~n7733 & ~n42962;
  assign n42964 = ~n7733 & ~n42963;
  assign n42965 = ~n7928 & ~n42964;
  assign n42966 = ~n8231 & ~n42945;
  assign n42967 = controllable_locked & ~n42966;
  assign n42968 = controllable_hmastlock & ~n40216;
  assign n42969 = ~n42954 & ~n42968;
  assign n42970 = ~controllable_locked & ~n42969;
  assign n42971 = ~n42967 & ~n42970;
  assign n42972 = controllable_hgrant2 & ~n42971;
  assign n42973 = ~n16724 & ~n42972;
  assign n42974 = n7928 & ~n42973;
  assign n42975 = ~n42965 & ~n42974;
  assign n42976 = ~controllable_hgrant1 & ~n42975;
  assign n42977 = ~n42944 & ~n42976;
  assign n42978 = ~controllable_hgrant3 & ~n42977;
  assign n42979 = ~n42940 & ~n42978;
  assign n42980 = ~controllable_hgrant4 & ~n42979;
  assign n42981 = ~n42936 & ~n42980;
  assign n42982 = ~controllable_hgrant5 & ~n42981;
  assign n42983 = ~n42932 & ~n42982;
  assign n42984 = ~controllable_hmaster2 & ~n42983;
  assign n42985 = ~n42820 & ~n42984;
  assign n42986 = controllable_hmaster1 & ~n42985;
  assign n42987 = n8378 & ~n9220;
  assign n42988 = ~n8378 & ~n19296;
  assign n42989 = ~n42987 & ~n42988;
  assign n42990 = controllable_hgrant5 & ~n42989;
  assign n42991 = n8426 & ~n12635;
  assign n42992 = ~n8426 & ~n19188;
  assign n42993 = ~n42991 & ~n42992;
  assign n42994 = i_hlock4 & ~n42993;
  assign n42995 = n8426 & ~n12653;
  assign n42996 = ~n8426 & ~n19194;
  assign n42997 = ~n42995 & ~n42996;
  assign n42998 = ~i_hlock4 & ~n42997;
  assign n42999 = ~n42994 & ~n42998;
  assign n43000 = controllable_hgrant4 & ~n42999;
  assign n43001 = i_hlock4 & ~n42767;
  assign n43002 = ~i_hlock4 & ~n42800;
  assign n43003 = ~n43001 & ~n43002;
  assign n43004 = ~controllable_hgrant4 & ~n43003;
  assign n43005 = ~n43000 & ~n43004;
  assign n43006 = ~controllable_hgrant5 & ~n43005;
  assign n43007 = ~n42990 & ~n43006;
  assign n43008 = controllable_hmaster2 & ~n43007;
  assign n43009 = n8378 & ~n9222;
  assign n43010 = ~n8378 & ~n19306;
  assign n43011 = ~n43009 & ~n43010;
  assign n43012 = controllable_hgrant5 & ~n43011;
  assign n43013 = n8426 & ~n9222;
  assign n43014 = ~n8426 & ~n19304;
  assign n43015 = ~n43013 & ~n43014;
  assign n43016 = controllable_hgrant4 & ~n43015;
  assign n43017 = n8365 & ~n9222;
  assign n43018 = ~n8365 & ~n19302;
  assign n43019 = ~n43017 & ~n43018;
  assign n43020 = controllable_hgrant3 & ~n43019;
  assign n43021 = n8389 & ~n9222;
  assign n43022 = ~n8389 & ~n19300;
  assign n43023 = ~n43021 & ~n43022;
  assign n43024 = controllable_hgrant1 & ~n43023;
  assign n43025 = ~n8440 & ~n42762;
  assign n43026 = ~controllable_hgrant1 & ~n43025;
  assign n43027 = ~n43024 & ~n43026;
  assign n43028 = ~controllable_hgrant3 & ~n43027;
  assign n43029 = ~n43020 & ~n43028;
  assign n43030 = ~controllable_hgrant4 & ~n43029;
  assign n43031 = ~n43016 & ~n43030;
  assign n43032 = ~controllable_hgrant5 & ~n43031;
  assign n43033 = ~n43012 & ~n43032;
  assign n43034 = ~controllable_hmaster2 & ~n43033;
  assign n43035 = ~n43008 & ~n43034;
  assign n43036 = ~controllable_hmaster1 & ~n43035;
  assign n43037 = ~n42986 & ~n43036;
  assign n43038 = i_hlock6 & ~n43037;
  assign n43039 = controllable_hmaster2 & ~n42804;
  assign n43040 = ~n42984 & ~n43039;
  assign n43041 = controllable_hmaster1 & ~n43040;
  assign n43042 = ~n43036 & ~n43041;
  assign n43043 = ~i_hlock6 & ~n43042;
  assign n43044 = ~n43038 & ~n43043;
  assign n43045 = ~controllable_hgrant6 & ~n43044;
  assign n43046 = ~n42928 & ~n43045;
  assign n43047 = ~controllable_hmaster0 & ~n43046;
  assign n43048 = ~n42906 & ~n43047;
  assign n43049 = ~controllable_hmaster3 & ~n43048;
  assign n43050 = ~n42815 & ~n43049;
  assign n43051 = i_hlock7 & ~n43050;
  assign n43052 = n8217 & ~n9240;
  assign n43053 = ~n8217 & ~n19331;
  assign n43054 = ~n43052 & ~n43053;
  assign n43055 = controllable_hgrant6 & ~n43054;
  assign n43056 = ~n42848 & ~n43039;
  assign n43057 = controllable_hmaster1 & ~n43056;
  assign n43058 = ~n42902 & ~n43057;
  assign n43059 = ~controllable_hgrant6 & ~n43058;
  assign n43060 = ~n43055 & ~n43059;
  assign n43061 = controllable_hmaster0 & ~n43060;
  assign n43062 = ~n43047 & ~n43061;
  assign n43063 = ~controllable_hmaster3 & ~n43062;
  assign n43064 = ~n42815 & ~n43063;
  assign n43065 = ~i_hlock7 & ~n43064;
  assign n43066 = ~n43051 & ~n43065;
  assign n43067 = i_hbusreq7 & ~n43066;
  assign n43068 = i_hbusreq8 & ~n42814;
  assign n43069 = i_hbusreq6 & ~n42704;
  assign n43070 = n8217 & ~n9263;
  assign n43071 = ~n8217 & ~n29767;
  assign n43072 = ~n43070 & ~n43071;
  assign n43073 = ~i_hbusreq6 & ~n43072;
  assign n43074 = ~n43069 & ~n43073;
  assign n43075 = controllable_hgrant6 & ~n43074;
  assign n43076 = i_hbusreq6 & ~n42742;
  assign n43077 = i_hbusreq5 & ~n42708;
  assign n43078 = n8378 & ~n9256;
  assign n43079 = ~n8378 & ~n19361;
  assign n43080 = ~n43078 & ~n43079;
  assign n43081 = ~i_hbusreq5 & ~n43080;
  assign n43082 = ~n43077 & ~n43081;
  assign n43083 = controllable_hgrant5 & ~n43082;
  assign n43084 = i_hbusreq5 & ~n42735;
  assign n43085 = i_hbusreq4 & ~n42712;
  assign n43086 = i_hbusreq9 & ~n42712;
  assign n43087 = n8426 & ~n9252;
  assign n43088 = ~n8426 & ~n19355;
  assign n43089 = ~n43087 & ~n43088;
  assign n43090 = ~i_hbusreq9 & ~n43089;
  assign n43091 = ~n43086 & ~n43090;
  assign n43092 = ~i_hbusreq4 & ~n43091;
  assign n43093 = ~n43085 & ~n43092;
  assign n43094 = controllable_hgrant4 & ~n43093;
  assign n43095 = i_hbusreq4 & ~n42733;
  assign n43096 = i_hbusreq9 & ~n42733;
  assign n43097 = i_hbusreq3 & ~n42716;
  assign n43098 = n8365 & ~n9250;
  assign n43099 = ~n8365 & ~n19351;
  assign n43100 = ~n43098 & ~n43099;
  assign n43101 = ~i_hbusreq3 & ~n43100;
  assign n43102 = ~n43097 & ~n43101;
  assign n43103 = controllable_hgrant3 & ~n43102;
  assign n43104 = i_hbusreq3 & ~n42731;
  assign n43105 = i_hbusreq1 & ~n42720;
  assign n43106 = n8389 & ~n8679;
  assign n43107 = ~n8389 & ~n16797;
  assign n43108 = ~n43106 & ~n43107;
  assign n43109 = ~i_hbusreq1 & ~n43108;
  assign n43110 = ~n43105 & ~n43109;
  assign n43111 = controllable_hgrant1 & ~n43110;
  assign n43112 = i_hbusreq1 & ~n42729;
  assign n43113 = ~n16400 & ~n40330;
  assign n43114 = ~n7928 & ~n43113;
  assign n43115 = i_hlock0 & ~n7978;
  assign n43116 = ~n16408 & ~n43115;
  assign n43117 = ~i_hbusreq0 & ~n43116;
  assign n43118 = ~n7969 & ~n43117;
  assign n43119 = ~i_hbusreq2 & ~n43118;
  assign n43120 = ~n7968 & ~n43119;
  assign n43121 = ~controllable_hgrant2 & n43120;
  assign n43122 = ~n40330 & ~n43121;
  assign n43123 = ~n7733 & ~n43122;
  assign n43124 = n7733 & ~n43113;
  assign n43125 = ~n43123 & ~n43124;
  assign n43126 = n7928 & ~n43125;
  assign n43127 = ~n43114 & ~n43126;
  assign n43128 = ~i_hbusreq1 & ~n43127;
  assign n43129 = ~n43112 & ~n43128;
  assign n43130 = ~controllable_hgrant1 & ~n43129;
  assign n43131 = ~n43111 & ~n43130;
  assign n43132 = ~i_hbusreq3 & ~n43131;
  assign n43133 = ~n43104 & ~n43132;
  assign n43134 = ~controllable_hgrant3 & ~n43133;
  assign n43135 = ~n43103 & ~n43134;
  assign n43136 = ~i_hbusreq9 & ~n43135;
  assign n43137 = ~n43096 & ~n43136;
  assign n43138 = ~i_hbusreq4 & ~n43137;
  assign n43139 = ~n43095 & ~n43138;
  assign n43140 = ~controllable_hgrant4 & ~n43139;
  assign n43141 = ~n43094 & ~n43140;
  assign n43142 = ~i_hbusreq5 & ~n43141;
  assign n43143 = ~n43084 & ~n43142;
  assign n43144 = ~controllable_hgrant5 & ~n43143;
  assign n43145 = ~n43083 & ~n43144;
  assign n43146 = controllable_hmaster1 & ~n43145;
  assign n43147 = controllable_hmaster2 & ~n43145;
  assign n43148 = ~n40407 & ~n43147;
  assign n43149 = ~controllable_hmaster1 & ~n43148;
  assign n43150 = ~n43146 & ~n43149;
  assign n43151 = ~i_hbusreq6 & ~n43150;
  assign n43152 = ~n43076 & ~n43151;
  assign n43153 = ~controllable_hgrant6 & ~n43152;
  assign n43154 = ~n43075 & ~n43153;
  assign n43155 = controllable_hmaster0 & ~n43154;
  assign n43156 = i_hbusreq6 & ~n42747;
  assign n43157 = n8217 & ~n9282;
  assign n43158 = ~n8217 & ~n20315;
  assign n43159 = ~n43157 & ~n43158;
  assign n43160 = ~i_hbusreq6 & ~n43159;
  assign n43161 = ~n43156 & ~n43160;
  assign n43162 = controllable_hgrant6 & ~n43161;
  assign n43163 = i_hbusreq6 & ~n42775;
  assign n43164 = i_hbusreq5 & ~n42750;
  assign n43165 = n8378 & ~n9276;
  assign n43166 = ~n8378 & ~n19464;
  assign n43167 = ~n43165 & ~n43166;
  assign n43168 = ~i_hbusreq5 & ~n43167;
  assign n43169 = ~n43164 & ~n43168;
  assign n43170 = controllable_hgrant5 & ~n43169;
  assign n43171 = i_hbusreq5 & ~n42769;
  assign n43172 = i_hbusreq4 & ~n42753;
  assign n43173 = i_hbusreq9 & ~n42753;
  assign n43174 = n8426 & ~n9272;
  assign n43175 = ~n8426 & ~n19458;
  assign n43176 = ~n43174 & ~n43175;
  assign n43177 = ~i_hbusreq9 & ~n43176;
  assign n43178 = ~n43173 & ~n43177;
  assign n43179 = ~i_hbusreq4 & ~n43178;
  assign n43180 = ~n43172 & ~n43179;
  assign n43181 = controllable_hgrant4 & ~n43180;
  assign n43182 = i_hbusreq4 & ~n42767;
  assign n43183 = i_hbusreq9 & ~n42767;
  assign n43184 = i_hbusreq3 & ~n42756;
  assign n43185 = n8365 & ~n9270;
  assign n43186 = ~n8365 & ~n19454;
  assign n43187 = ~n43185 & ~n43186;
  assign n43188 = ~i_hbusreq3 & ~n43187;
  assign n43189 = ~n43184 & ~n43188;
  assign n43190 = controllable_hgrant3 & ~n43189;
  assign n43191 = i_hbusreq3 & ~n42765;
  assign n43192 = i_hbusreq1 & ~n42759;
  assign n43193 = n8389 & ~n9268;
  assign n43194 = ~n8389 & ~n19450;
  assign n43195 = ~n43193 & ~n43194;
  assign n43196 = ~i_hbusreq1 & ~n43195;
  assign n43197 = ~n43192 & ~n43196;
  assign n43198 = controllable_hgrant1 & ~n43197;
  assign n43199 = i_hbusreq1 & ~n42763;
  assign n43200 = ~n16796 & ~n40330;
  assign n43201 = n7928 & ~n43200;
  assign n43202 = ~n8265 & ~n43201;
  assign n43203 = ~i_hbusreq1 & ~n43202;
  assign n43204 = ~n43199 & ~n43203;
  assign n43205 = ~controllable_hgrant1 & ~n43204;
  assign n43206 = ~n43198 & ~n43205;
  assign n43207 = ~i_hbusreq3 & ~n43206;
  assign n43208 = ~n43191 & ~n43207;
  assign n43209 = ~controllable_hgrant3 & ~n43208;
  assign n43210 = ~n43190 & ~n43209;
  assign n43211 = ~i_hbusreq9 & ~n43210;
  assign n43212 = ~n43183 & ~n43211;
  assign n43213 = ~i_hbusreq4 & ~n43212;
  assign n43214 = ~n43182 & ~n43213;
  assign n43215 = ~controllable_hgrant4 & ~n43214;
  assign n43216 = ~n43181 & ~n43215;
  assign n43217 = ~i_hbusreq5 & ~n43216;
  assign n43218 = ~n43171 & ~n43217;
  assign n43219 = ~controllable_hgrant5 & ~n43218;
  assign n43220 = ~n43170 & ~n43219;
  assign n43221 = ~controllable_hmaster2 & ~n43220;
  assign n43222 = ~n43147 & ~n43221;
  assign n43223 = ~controllable_hmaster1 & ~n43222;
  assign n43224 = ~n43146 & ~n43223;
  assign n43225 = ~i_hbusreq6 & ~n43224;
  assign n43226 = ~n43163 & ~n43225;
  assign n43227 = ~controllable_hgrant6 & ~n43226;
  assign n43228 = ~n43162 & ~n43227;
  assign n43229 = ~controllable_hmaster0 & ~n43228;
  assign n43230 = ~n43155 & ~n43229;
  assign n43231 = i_hlock8 & ~n43230;
  assign n43232 = i_hbusreq6 & ~n42782;
  assign n43233 = n8217 & ~n9302;
  assign n43234 = ~n8217 & ~n20327;
  assign n43235 = ~n43233 & ~n43234;
  assign n43236 = ~i_hbusreq6 & ~n43235;
  assign n43237 = ~n43232 & ~n43236;
  assign n43238 = controllable_hgrant6 & ~n43237;
  assign n43239 = i_hbusreq6 & ~n42808;
  assign n43240 = i_hbusreq5 & ~n42785;
  assign n43241 = n8378 & ~n9296;
  assign n43242 = ~n8378 & ~n19514;
  assign n43243 = ~n43241 & ~n43242;
  assign n43244 = ~i_hbusreq5 & ~n43243;
  assign n43245 = ~n43240 & ~n43244;
  assign n43246 = controllable_hgrant5 & ~n43245;
  assign n43247 = i_hbusreq5 & ~n42802;
  assign n43248 = i_hbusreq4 & ~n42788;
  assign n43249 = i_hbusreq9 & ~n42788;
  assign n43250 = n8426 & ~n9292;
  assign n43251 = ~n8426 & ~n19508;
  assign n43252 = ~n43250 & ~n43251;
  assign n43253 = ~i_hbusreq9 & ~n43252;
  assign n43254 = ~n43249 & ~n43253;
  assign n43255 = ~i_hbusreq4 & ~n43254;
  assign n43256 = ~n43248 & ~n43255;
  assign n43257 = controllable_hgrant4 & ~n43256;
  assign n43258 = i_hbusreq4 & ~n42800;
  assign n43259 = i_hbusreq9 & ~n42800;
  assign n43260 = i_hbusreq3 & ~n42791;
  assign n43261 = n8365 & ~n9290;
  assign n43262 = ~n8365 & ~n19480;
  assign n43263 = ~n43261 & ~n43262;
  assign n43264 = ~i_hbusreq3 & ~n43263;
  assign n43265 = ~n43260 & ~n43264;
  assign n43266 = controllable_hgrant3 & ~n43265;
  assign n43267 = i_hbusreq3 & ~n42798;
  assign n43268 = i_hbusreq1 & ~n42794;
  assign n43269 = n8389 & ~n9288;
  assign n43270 = ~n8389 & ~n19476;
  assign n43271 = ~n43269 & ~n43270;
  assign n43272 = ~i_hbusreq1 & ~n43271;
  assign n43273 = ~n43268 & ~n43272;
  assign n43274 = controllable_hgrant1 & ~n43273;
  assign n43275 = i_hbusreq1 & ~n42796;
  assign n43276 = ~n8297 & ~n43201;
  assign n43277 = ~i_hbusreq1 & ~n43276;
  assign n43278 = ~n43275 & ~n43277;
  assign n43279 = ~controllable_hgrant1 & ~n43278;
  assign n43280 = ~n43274 & ~n43279;
  assign n43281 = ~i_hbusreq3 & ~n43280;
  assign n43282 = ~n43267 & ~n43281;
  assign n43283 = ~controllable_hgrant3 & ~n43282;
  assign n43284 = ~n43266 & ~n43283;
  assign n43285 = ~i_hbusreq9 & ~n43284;
  assign n43286 = ~n43259 & ~n43285;
  assign n43287 = ~i_hbusreq4 & ~n43286;
  assign n43288 = ~n43258 & ~n43287;
  assign n43289 = ~controllable_hgrant4 & ~n43288;
  assign n43290 = ~n43257 & ~n43289;
  assign n43291 = ~i_hbusreq5 & ~n43290;
  assign n43292 = ~n43247 & ~n43291;
  assign n43293 = ~controllable_hgrant5 & ~n43292;
  assign n43294 = ~n43246 & ~n43293;
  assign n43295 = ~controllable_hmaster2 & ~n43294;
  assign n43296 = ~n43147 & ~n43295;
  assign n43297 = ~controllable_hmaster1 & ~n43296;
  assign n43298 = ~n43146 & ~n43297;
  assign n43299 = ~i_hbusreq6 & ~n43298;
  assign n43300 = ~n43239 & ~n43299;
  assign n43301 = ~controllable_hgrant6 & ~n43300;
  assign n43302 = ~n43238 & ~n43301;
  assign n43303 = ~controllable_hmaster0 & ~n43302;
  assign n43304 = ~n43155 & ~n43303;
  assign n43305 = ~i_hlock8 & ~n43304;
  assign n43306 = ~n43231 & ~n43305;
  assign n43307 = ~i_hbusreq8 & ~n43306;
  assign n43308 = ~n43068 & ~n43307;
  assign n43309 = controllable_hmaster3 & ~n43308;
  assign n43310 = i_hbusreq8 & ~n43048;
  assign n43311 = i_hbusreq6 & ~n42818;
  assign n43312 = n8217 & ~n9361;
  assign n43313 = ~n8217 & ~n19551;
  assign n43314 = ~n43312 & ~n43313;
  assign n43315 = ~i_hbusreq6 & ~n43314;
  assign n43316 = ~n43311 & ~n43315;
  assign n43317 = controllable_hgrant6 & ~n43316;
  assign n43318 = i_hbusreq6 & ~n42903;
  assign n43319 = controllable_hmaster2 & ~n43220;
  assign n43320 = i_hbusreq5 & ~n42823;
  assign n43321 = n8378 & ~n9327;
  assign n43322 = ~n8378 & ~n19492;
  assign n43323 = ~n43321 & ~n43322;
  assign n43324 = ~i_hbusreq5 & ~n43323;
  assign n43325 = ~n43320 & ~n43324;
  assign n43326 = controllable_hgrant5 & ~n43325;
  assign n43327 = i_hbusreq5 & ~n42845;
  assign n43328 = i_hbusreq4 & ~n42827;
  assign n43329 = i_hbusreq9 & ~n42827;
  assign n43330 = n8426 & ~n9323;
  assign n43331 = ~n8426 & ~n19486;
  assign n43332 = ~n43330 & ~n43331;
  assign n43333 = ~i_hbusreq9 & ~n43332;
  assign n43334 = ~n43329 & ~n43333;
  assign n43335 = ~i_hbusreq4 & ~n43334;
  assign n43336 = ~n43328 & ~n43335;
  assign n43337 = controllable_hgrant4 & ~n43336;
  assign n43338 = i_hbusreq4 & ~n42843;
  assign n43339 = i_hbusreq9 & ~n42843;
  assign n43340 = i_hbusreq3 & ~n42837;
  assign n43341 = n8365 & ~n14328;
  assign n43342 = ~n8365 & ~n19378;
  assign n43343 = ~n43341 & ~n43342;
  assign n43344 = i_hlock3 & ~n43343;
  assign n43345 = n8365 & ~n14338;
  assign n43346 = ~n8365 & ~n19390;
  assign n43347 = ~n43345 & ~n43346;
  assign n43348 = ~i_hlock3 & ~n43347;
  assign n43349 = ~n43344 & ~n43348;
  assign n43350 = ~i_hbusreq3 & ~n43349;
  assign n43351 = ~n43340 & ~n43350;
  assign n43352 = controllable_hgrant3 & ~n43351;
  assign n43353 = i_hbusreq3 & ~n42841;
  assign n43354 = i_hlock3 & ~n43206;
  assign n43355 = ~i_hlock3 & ~n43280;
  assign n43356 = ~n43354 & ~n43355;
  assign n43357 = ~i_hbusreq3 & ~n43356;
  assign n43358 = ~n43353 & ~n43357;
  assign n43359 = ~controllable_hgrant3 & ~n43358;
  assign n43360 = ~n43352 & ~n43359;
  assign n43361 = ~i_hbusreq9 & ~n43360;
  assign n43362 = ~n43339 & ~n43361;
  assign n43363 = ~i_hbusreq4 & ~n43362;
  assign n43364 = ~n43338 & ~n43363;
  assign n43365 = ~controllable_hgrant4 & ~n43364;
  assign n43366 = ~n43337 & ~n43365;
  assign n43367 = ~i_hbusreq5 & ~n43366;
  assign n43368 = ~n43327 & ~n43367;
  assign n43369 = ~controllable_hgrant5 & ~n43368;
  assign n43370 = ~n43326 & ~n43369;
  assign n43371 = ~controllable_hmaster2 & ~n43370;
  assign n43372 = ~n43319 & ~n43371;
  assign n43373 = controllable_hmaster1 & ~n43372;
  assign n43374 = i_hbusreq5 & ~n42859;
  assign n43375 = n8378 & ~n27221;
  assign n43376 = ~n8378 & ~n29791;
  assign n43377 = ~n43375 & ~n43376;
  assign n43378 = i_hlock5 & ~n43377;
  assign n43379 = n8378 & ~n27248;
  assign n43380 = ~n8378 & ~n29821;
  assign n43381 = ~n43379 & ~n43380;
  assign n43382 = ~i_hlock5 & ~n43381;
  assign n43383 = ~n43378 & ~n43382;
  assign n43384 = ~i_hbusreq5 & ~n43383;
  assign n43385 = ~n43374 & ~n43384;
  assign n43386 = controllable_hgrant5 & ~n43385;
  assign n43387 = i_hbusreq5 & ~n42863;
  assign n43388 = i_hlock5 & ~n43216;
  assign n43389 = ~i_hlock5 & ~n43290;
  assign n43390 = ~n43388 & ~n43389;
  assign n43391 = ~i_hbusreq5 & ~n43390;
  assign n43392 = ~n43387 & ~n43391;
  assign n43393 = ~controllable_hgrant5 & ~n43392;
  assign n43394 = ~n43386 & ~n43393;
  assign n43395 = controllable_hmaster2 & ~n43394;
  assign n43396 = i_hbusreq5 & ~n42869;
  assign n43397 = n8378 & ~n9355;
  assign n43398 = ~n8378 & ~n19543;
  assign n43399 = ~n43397 & ~n43398;
  assign n43400 = ~i_hbusreq5 & ~n43399;
  assign n43401 = ~n43396 & ~n43400;
  assign n43402 = controllable_hgrant5 & ~n43401;
  assign n43403 = i_hbusreq5 & ~n42897;
  assign n43404 = i_hbusreq4 & ~n42873;
  assign n43405 = i_hbusreq9 & ~n42873;
  assign n43406 = n8426 & ~n9351;
  assign n43407 = ~n8426 & ~n19537;
  assign n43408 = ~n43406 & ~n43407;
  assign n43409 = ~i_hbusreq9 & ~n43408;
  assign n43410 = ~n43405 & ~n43409;
  assign n43411 = ~i_hbusreq4 & ~n43410;
  assign n43412 = ~n43404 & ~n43411;
  assign n43413 = controllable_hgrant4 & ~n43412;
  assign n43414 = i_hbusreq4 & ~n42895;
  assign n43415 = i_hbusreq9 & ~n42895;
  assign n43416 = i_hbusreq3 & ~n42877;
  assign n43417 = n8365 & ~n9349;
  assign n43418 = ~n8365 & ~n19533;
  assign n43419 = ~n43417 & ~n43418;
  assign n43420 = ~i_hbusreq3 & ~n43419;
  assign n43421 = ~n43416 & ~n43420;
  assign n43422 = controllable_hgrant3 & ~n43421;
  assign n43423 = i_hbusreq3 & ~n42893;
  assign n43424 = i_hbusreq1 & ~n42887;
  assign n43425 = n8389 & ~n14324;
  assign n43426 = ~n8389 & ~n19374;
  assign n43427 = ~n43425 & ~n43426;
  assign n43428 = i_hlock1 & ~n43427;
  assign n43429 = n8389 & ~n14334;
  assign n43430 = ~n8389 & ~n19386;
  assign n43431 = ~n43429 & ~n43430;
  assign n43432 = ~i_hlock1 & ~n43431;
  assign n43433 = ~n43428 & ~n43432;
  assign n43434 = ~i_hbusreq1 & ~n43433;
  assign n43435 = ~n43424 & ~n43434;
  assign n43436 = controllable_hgrant1 & ~n43435;
  assign n43437 = i_hbusreq1 & ~n42891;
  assign n43438 = i_hlock1 & ~n43202;
  assign n43439 = ~i_hlock1 & ~n43276;
  assign n43440 = ~n43438 & ~n43439;
  assign n43441 = ~i_hbusreq1 & ~n43440;
  assign n43442 = ~n43437 & ~n43441;
  assign n43443 = ~controllable_hgrant1 & ~n43442;
  assign n43444 = ~n43436 & ~n43443;
  assign n43445 = ~i_hbusreq3 & ~n43444;
  assign n43446 = ~n43423 & ~n43445;
  assign n43447 = ~controllable_hgrant3 & ~n43446;
  assign n43448 = ~n43422 & ~n43447;
  assign n43449 = ~i_hbusreq9 & ~n43448;
  assign n43450 = ~n43415 & ~n43449;
  assign n43451 = ~i_hbusreq4 & ~n43450;
  assign n43452 = ~n43414 & ~n43451;
  assign n43453 = ~controllable_hgrant4 & ~n43452;
  assign n43454 = ~n43413 & ~n43453;
  assign n43455 = ~i_hbusreq5 & ~n43454;
  assign n43456 = ~n43403 & ~n43455;
  assign n43457 = ~controllable_hgrant5 & ~n43456;
  assign n43458 = ~n43402 & ~n43457;
  assign n43459 = ~controllable_hmaster2 & ~n43458;
  assign n43460 = ~n43395 & ~n43459;
  assign n43461 = ~controllable_hmaster1 & ~n43460;
  assign n43462 = ~n43373 & ~n43461;
  assign n43463 = ~i_hbusreq6 & ~n43462;
  assign n43464 = ~n43318 & ~n43463;
  assign n43465 = ~controllable_hgrant6 & ~n43464;
  assign n43466 = ~n43317 & ~n43465;
  assign n43467 = controllable_hmaster0 & ~n43466;
  assign n43468 = i_hbusreq6 & ~n42927;
  assign n43469 = ~n9391 & ~n27226;
  assign n43470 = controllable_hmaster1 & ~n43469;
  assign n43471 = ~n9428 & ~n43470;
  assign n43472 = n8217 & ~n43471;
  assign n43473 = ~n19582 & ~n29796;
  assign n43474 = controllable_hmaster1 & ~n43473;
  assign n43475 = ~n19626 & ~n43474;
  assign n43476 = ~n8217 & ~n43475;
  assign n43477 = ~n43472 & ~n43476;
  assign n43478 = i_hlock6 & ~n43477;
  assign n43479 = ~n9391 & ~n27253;
  assign n43480 = controllable_hmaster1 & ~n43479;
  assign n43481 = ~n9428 & ~n43480;
  assign n43482 = n8217 & ~n43481;
  assign n43483 = ~n19582 & ~n29826;
  assign n43484 = controllable_hmaster1 & ~n43483;
  assign n43485 = ~n19626 & ~n43484;
  assign n43486 = ~n8217 & ~n43485;
  assign n43487 = ~n43482 & ~n43486;
  assign n43488 = ~i_hlock6 & ~n43487;
  assign n43489 = ~n43478 & ~n43488;
  assign n43490 = ~i_hbusreq6 & ~n43489;
  assign n43491 = ~n43468 & ~n43490;
  assign n43492 = controllable_hgrant6 & ~n43491;
  assign n43493 = i_hbusreq6 & ~n43044;
  assign n43494 = i_hbusreq5 & ~n42931;
  assign n43495 = n8378 & ~n9388;
  assign n43496 = ~n8378 & ~n19577;
  assign n43497 = ~n43495 & ~n43496;
  assign n43498 = ~i_hbusreq5 & ~n43497;
  assign n43499 = ~n43494 & ~n43498;
  assign n43500 = controllable_hgrant5 & ~n43499;
  assign n43501 = i_hbusreq5 & ~n42981;
  assign n43502 = i_hbusreq4 & ~n42935;
  assign n43503 = i_hbusreq9 & ~n42935;
  assign n43504 = n8426 & ~n9384;
  assign n43505 = ~n8426 & ~n19571;
  assign n43506 = ~n43504 & ~n43505;
  assign n43507 = ~i_hbusreq9 & ~n43506;
  assign n43508 = ~n43503 & ~n43507;
  assign n43509 = ~i_hbusreq4 & ~n43508;
  assign n43510 = ~n43502 & ~n43509;
  assign n43511 = controllable_hgrant4 & ~n43510;
  assign n43512 = i_hbusreq4 & ~n42979;
  assign n43513 = i_hbusreq9 & ~n42979;
  assign n43514 = i_hbusreq3 & ~n42939;
  assign n43515 = n8365 & ~n9382;
  assign n43516 = ~n8365 & ~n19567;
  assign n43517 = ~n43515 & ~n43516;
  assign n43518 = ~i_hbusreq3 & ~n43517;
  assign n43519 = ~n43514 & ~n43518;
  assign n43520 = controllable_hgrant3 & ~n43519;
  assign n43521 = i_hbusreq3 & ~n42977;
  assign n43522 = i_hbusreq1 & ~n42943;
  assign n43523 = n8389 & ~n9380;
  assign n43524 = ~n8389 & ~n19563;
  assign n43525 = ~n43523 & ~n43524;
  assign n43526 = ~i_hbusreq1 & ~n43525;
  assign n43527 = ~n43522 & ~n43526;
  assign n43528 = controllable_hgrant1 & ~n43527;
  assign n43529 = i_hbusreq1 & ~n42975;
  assign n43530 = i_hbusreq2 & ~n42959;
  assign n43531 = i_hbusreq0 & ~n42950;
  assign n43532 = ~n40082 & ~n43531;
  assign n43533 = i_hlock2 & ~n43532;
  assign n43534 = i_hbusreq0 & ~n42957;
  assign n43535 = ~n40082 & ~n43534;
  assign n43536 = ~i_hlock2 & ~n43535;
  assign n43537 = ~n43533 & ~n43536;
  assign n43538 = ~i_hbusreq2 & ~n43537;
  assign n43539 = ~n43530 & ~n43538;
  assign n43540 = controllable_hgrant2 & ~n43539;
  assign n43541 = ~controllable_hgrant2 & ~n9376;
  assign n43542 = ~n43540 & ~n43541;
  assign n43543 = ~n7733 & ~n43542;
  assign n43544 = ~n7733 & ~n43543;
  assign n43545 = ~n7928 & ~n43544;
  assign n43546 = i_hbusreq2 & ~n42971;
  assign n43547 = i_hbusreq0 & ~n42971;
  assign n43548 = ~n39848 & ~n40337;
  assign n43549 = ~controllable_locked & ~n43548;
  assign n43550 = ~n40078 & ~n43549;
  assign n43551 = i_hlock0 & ~n43550;
  assign n43552 = ~i_hlock0 & ~n42971;
  assign n43553 = ~n43551 & ~n43552;
  assign n43554 = ~i_hbusreq0 & ~n43553;
  assign n43555 = ~n43547 & ~n43554;
  assign n43556 = ~i_hbusreq2 & ~n43555;
  assign n43557 = ~n43546 & ~n43556;
  assign n43558 = controllable_hgrant2 & ~n43557;
  assign n43559 = ~n16796 & ~n43558;
  assign n43560 = n7928 & ~n43559;
  assign n43561 = ~n43545 & ~n43560;
  assign n43562 = ~i_hbusreq1 & ~n43561;
  assign n43563 = ~n43529 & ~n43562;
  assign n43564 = ~controllable_hgrant1 & ~n43563;
  assign n43565 = ~n43528 & ~n43564;
  assign n43566 = ~i_hbusreq3 & ~n43565;
  assign n43567 = ~n43521 & ~n43566;
  assign n43568 = ~controllable_hgrant3 & ~n43567;
  assign n43569 = ~n43520 & ~n43568;
  assign n43570 = ~i_hbusreq9 & ~n43569;
  assign n43571 = ~n43513 & ~n43570;
  assign n43572 = ~i_hbusreq4 & ~n43571;
  assign n43573 = ~n43512 & ~n43572;
  assign n43574 = ~controllable_hgrant4 & ~n43573;
  assign n43575 = ~n43511 & ~n43574;
  assign n43576 = ~i_hbusreq5 & ~n43575;
  assign n43577 = ~n43501 & ~n43576;
  assign n43578 = ~controllable_hgrant5 & ~n43577;
  assign n43579 = ~n43500 & ~n43578;
  assign n43580 = ~controllable_hmaster2 & ~n43579;
  assign n43581 = ~n43319 & ~n43580;
  assign n43582 = controllable_hmaster1 & ~n43581;
  assign n43583 = i_hbusreq5 & ~n42989;
  assign n43584 = n8378 & ~n9400;
  assign n43585 = ~n8378 & ~n19593;
  assign n43586 = ~n43584 & ~n43585;
  assign n43587 = ~i_hbusreq5 & ~n43586;
  assign n43588 = ~n43583 & ~n43587;
  assign n43589 = controllable_hgrant5 & ~n43588;
  assign n43590 = i_hbusreq5 & ~n43005;
  assign n43591 = i_hbusreq4 & ~n42999;
  assign n43592 = i_hbusreq9 & ~n42993;
  assign n43593 = n8426 & ~n14332;
  assign n43594 = ~n8426 & ~n19382;
  assign n43595 = ~n43593 & ~n43594;
  assign n43596 = ~i_hbusreq9 & ~n43595;
  assign n43597 = ~n43592 & ~n43596;
  assign n43598 = i_hlock4 & ~n43597;
  assign n43599 = i_hbusreq9 & ~n42997;
  assign n43600 = n8426 & ~n14342;
  assign n43601 = ~n8426 & ~n19394;
  assign n43602 = ~n43600 & ~n43601;
  assign n43603 = ~i_hbusreq9 & ~n43602;
  assign n43604 = ~n43599 & ~n43603;
  assign n43605 = ~i_hlock4 & ~n43604;
  assign n43606 = ~n43598 & ~n43605;
  assign n43607 = ~i_hbusreq4 & ~n43606;
  assign n43608 = ~n43591 & ~n43607;
  assign n43609 = controllable_hgrant4 & ~n43608;
  assign n43610 = i_hbusreq4 & ~n43003;
  assign n43611 = i_hlock4 & ~n43212;
  assign n43612 = ~i_hlock4 & ~n43286;
  assign n43613 = ~n43611 & ~n43612;
  assign n43614 = ~i_hbusreq4 & ~n43613;
  assign n43615 = ~n43610 & ~n43614;
  assign n43616 = ~controllable_hgrant4 & ~n43615;
  assign n43617 = ~n43609 & ~n43616;
  assign n43618 = ~i_hbusreq5 & ~n43617;
  assign n43619 = ~n43590 & ~n43618;
  assign n43620 = ~controllable_hgrant5 & ~n43619;
  assign n43621 = ~n43589 & ~n43620;
  assign n43622 = controllable_hmaster2 & ~n43621;
  assign n43623 = i_hbusreq5 & ~n43011;
  assign n43624 = n8378 & ~n9423;
  assign n43625 = ~n8378 & ~n19619;
  assign n43626 = ~n43624 & ~n43625;
  assign n43627 = ~i_hbusreq5 & ~n43626;
  assign n43628 = ~n43623 & ~n43627;
  assign n43629 = controllable_hgrant5 & ~n43628;
  assign n43630 = i_hbusreq5 & ~n43031;
  assign n43631 = i_hbusreq4 & ~n43015;
  assign n43632 = i_hbusreq9 & ~n43015;
  assign n43633 = n8426 & ~n9419;
  assign n43634 = ~n8426 & ~n19613;
  assign n43635 = ~n43633 & ~n43634;
  assign n43636 = ~i_hbusreq9 & ~n43635;
  assign n43637 = ~n43632 & ~n43636;
  assign n43638 = ~i_hbusreq4 & ~n43637;
  assign n43639 = ~n43631 & ~n43638;
  assign n43640 = controllable_hgrant4 & ~n43639;
  assign n43641 = i_hbusreq4 & ~n43029;
  assign n43642 = i_hbusreq9 & ~n43029;
  assign n43643 = i_hbusreq3 & ~n43019;
  assign n43644 = n8365 & ~n9417;
  assign n43645 = ~n8365 & ~n19609;
  assign n43646 = ~n43644 & ~n43645;
  assign n43647 = ~i_hbusreq3 & ~n43646;
  assign n43648 = ~n43643 & ~n43647;
  assign n43649 = controllable_hgrant3 & ~n43648;
  assign n43650 = i_hbusreq3 & ~n43027;
  assign n43651 = i_hbusreq1 & ~n43023;
  assign n43652 = n8389 & ~n9415;
  assign n43653 = ~n8389 & ~n19605;
  assign n43654 = ~n43652 & ~n43653;
  assign n43655 = ~i_hbusreq1 & ~n43654;
  assign n43656 = ~n43651 & ~n43655;
  assign n43657 = controllable_hgrant1 & ~n43656;
  assign n43658 = i_hbusreq1 & ~n43025;
  assign n43659 = ~controllable_hmastlock & ~n40320;
  assign n43660 = ~n42968 & ~n43659;
  assign n43661 = ~controllable_locked & ~n43660;
  assign n43662 = ~n14240 & ~n43661;
  assign n43663 = i_hlock0 & ~n43662;
  assign n43664 = ~n40324 & ~n43663;
  assign n43665 = ~i_hbusreq0 & ~n43664;
  assign n43666 = ~n40319 & ~n43665;
  assign n43667 = ~i_hbusreq2 & ~n43666;
  assign n43668 = ~n40318 & ~n43667;
  assign n43669 = controllable_hgrant2 & ~n43668;
  assign n43670 = ~n18452 & ~n43669;
  assign n43671 = n7928 & ~n43670;
  assign n43672 = ~n8440 & ~n43671;
  assign n43673 = ~i_hbusreq1 & ~n43672;
  assign n43674 = ~n43658 & ~n43673;
  assign n43675 = ~controllable_hgrant1 & ~n43674;
  assign n43676 = ~n43657 & ~n43675;
  assign n43677 = ~i_hbusreq3 & ~n43676;
  assign n43678 = ~n43650 & ~n43677;
  assign n43679 = ~controllable_hgrant3 & ~n43678;
  assign n43680 = ~n43649 & ~n43679;
  assign n43681 = ~i_hbusreq9 & ~n43680;
  assign n43682 = ~n43642 & ~n43681;
  assign n43683 = ~i_hbusreq4 & ~n43682;
  assign n43684 = ~n43641 & ~n43683;
  assign n43685 = ~controllable_hgrant4 & ~n43684;
  assign n43686 = ~n43640 & ~n43685;
  assign n43687 = ~i_hbusreq5 & ~n43686;
  assign n43688 = ~n43630 & ~n43687;
  assign n43689 = ~controllable_hgrant5 & ~n43688;
  assign n43690 = ~n43629 & ~n43689;
  assign n43691 = ~controllable_hmaster2 & ~n43690;
  assign n43692 = ~n43622 & ~n43691;
  assign n43693 = ~controllable_hmaster1 & ~n43692;
  assign n43694 = ~n43582 & ~n43693;
  assign n43695 = i_hlock6 & ~n43694;
  assign n43696 = controllable_hmaster2 & ~n43294;
  assign n43697 = ~n43580 & ~n43696;
  assign n43698 = controllable_hmaster1 & ~n43697;
  assign n43699 = ~n43693 & ~n43698;
  assign n43700 = ~i_hlock6 & ~n43699;
  assign n43701 = ~n43695 & ~n43700;
  assign n43702 = ~i_hbusreq6 & ~n43701;
  assign n43703 = ~n43493 & ~n43702;
  assign n43704 = ~controllable_hgrant6 & ~n43703;
  assign n43705 = ~n43492 & ~n43704;
  assign n43706 = ~controllable_hmaster0 & ~n43705;
  assign n43707 = ~n43467 & ~n43706;
  assign n43708 = ~i_hbusreq8 & ~n43707;
  assign n43709 = ~n43310 & ~n43708;
  assign n43710 = ~controllable_hmaster3 & ~n43709;
  assign n43711 = ~n43309 & ~n43710;
  assign n43712 = i_hlock7 & ~n43711;
  assign n43713 = i_hbusreq8 & ~n43062;
  assign n43714 = i_hbusreq6 & ~n43054;
  assign n43715 = n8217 & ~n9450;
  assign n43716 = ~n8217 & ~n19655;
  assign n43717 = ~n43715 & ~n43716;
  assign n43718 = ~i_hbusreq6 & ~n43717;
  assign n43719 = ~n43714 & ~n43718;
  assign n43720 = controllable_hgrant6 & ~n43719;
  assign n43721 = i_hbusreq6 & ~n43058;
  assign n43722 = ~n43371 & ~n43696;
  assign n43723 = controllable_hmaster1 & ~n43722;
  assign n43724 = ~n43461 & ~n43723;
  assign n43725 = ~i_hbusreq6 & ~n43724;
  assign n43726 = ~n43721 & ~n43725;
  assign n43727 = ~controllable_hgrant6 & ~n43726;
  assign n43728 = ~n43720 & ~n43727;
  assign n43729 = controllable_hmaster0 & ~n43728;
  assign n43730 = ~n43706 & ~n43729;
  assign n43731 = ~i_hbusreq8 & ~n43730;
  assign n43732 = ~n43713 & ~n43731;
  assign n43733 = ~controllable_hmaster3 & ~n43732;
  assign n43734 = ~n43309 & ~n43733;
  assign n43735 = ~i_hlock7 & ~n43734;
  assign n43736 = ~n43712 & ~n43735;
  assign n43737 = ~i_hbusreq7 & ~n43736;
  assign n43738 = ~n43067 & ~n43737;
  assign n43739 = ~n7924 & ~n43738;
  assign n43740 = ~n8217 & ~n29855;
  assign n43741 = ~n41555 & ~n43740;
  assign n43742 = controllable_hgrant6 & ~n43741;
  assign n43743 = n8378 & ~n13164;
  assign n43744 = ~n8378 & ~n19679;
  assign n43745 = ~n43743 & ~n43744;
  assign n43746 = controllable_hgrant5 & ~n43745;
  assign n43747 = n8426 & ~n13162;
  assign n43748 = ~n8426 & ~n19677;
  assign n43749 = ~n43747 & ~n43748;
  assign n43750 = controllable_hgrant4 & ~n43749;
  assign n43751 = n8365 & ~n13160;
  assign n43752 = ~n8365 & ~n19675;
  assign n43753 = ~n43751 & ~n43752;
  assign n43754 = controllable_hgrant3 & ~n43753;
  assign n43755 = n8389 & ~n13158;
  assign n43756 = ~n8389 & ~n19673;
  assign n43757 = ~n43755 & ~n43756;
  assign n43758 = controllable_hgrant1 & ~n43757;
  assign n43759 = ~controllable_locked & n39846;
  assign n43760 = ~n13008 & ~n43759;
  assign n43761 = controllable_hgrant2 & ~n43760;
  assign n43762 = ~n7733 & n43761;
  assign n43763 = ~n16505 & ~n43761;
  assign n43764 = n7733 & ~n43763;
  assign n43765 = ~n43762 & ~n43764;
  assign n43766 = n7928 & ~n43765;
  assign n43767 = ~n42723 & ~n43766;
  assign n43768 = ~controllable_hgrant1 & ~n43767;
  assign n43769 = ~n43758 & ~n43768;
  assign n43770 = ~controllable_hgrant3 & ~n43769;
  assign n43771 = ~n43754 & ~n43770;
  assign n43772 = ~controllable_hgrant4 & ~n43771;
  assign n43773 = ~n43750 & ~n43772;
  assign n43774 = ~controllable_hgrant5 & ~n43773;
  assign n43775 = ~n43746 & ~n43774;
  assign n43776 = controllable_hmaster1 & ~n43775;
  assign n43777 = controllable_hmaster2 & ~n43775;
  assign n43778 = ~n8378 & ~n29849;
  assign n43779 = ~n41580 & ~n43778;
  assign n43780 = controllable_hgrant5 & ~n43779;
  assign n43781 = ~n8426 & ~n19718;
  assign n43782 = ~n41584 & ~n43781;
  assign n43783 = i_hlock9 & ~n43782;
  assign n43784 = ~n8426 & ~n19736;
  assign n43785 = ~n41588 & ~n43784;
  assign n43786 = ~i_hlock9 & ~n43785;
  assign n43787 = ~n43783 & ~n43786;
  assign n43788 = controllable_hgrant4 & ~n43787;
  assign n43789 = ~n8365 & ~n19716;
  assign n43790 = ~n41594 & ~n43789;
  assign n43791 = controllable_hgrant3 & ~n43790;
  assign n43792 = ~n8389 & ~n19714;
  assign n43793 = ~n41598 & ~n43792;
  assign n43794 = controllable_hgrant1 & ~n43793;
  assign n43795 = ~n40224 & ~n43759;
  assign n43796 = controllable_hgrant2 & ~n43795;
  assign n43797 = ~n17090 & ~n43796;
  assign n43798 = n7733 & ~n43797;
  assign n43799 = ~n43762 & ~n43798;
  assign n43800 = n7928 & ~n43799;
  assign n43801 = ~n8221 & ~n43800;
  assign n43802 = ~controllable_hgrant1 & ~n43801;
  assign n43803 = ~n43794 & ~n43802;
  assign n43804 = ~controllable_hgrant3 & ~n43803;
  assign n43805 = ~n43791 & ~n43804;
  assign n43806 = i_hlock9 & ~n43805;
  assign n43807 = ~n8365 & ~n19734;
  assign n43808 = ~n41620 & ~n43807;
  assign n43809 = controllable_hgrant3 & ~n43808;
  assign n43810 = ~n8389 & ~n19732;
  assign n43811 = ~n41624 & ~n43810;
  assign n43812 = controllable_hgrant1 & ~n43811;
  assign n43813 = ~n8235 & ~n43800;
  assign n43814 = ~controllable_hgrant1 & ~n43813;
  assign n43815 = ~n43812 & ~n43814;
  assign n43816 = ~controllable_hgrant3 & ~n43815;
  assign n43817 = ~n43809 & ~n43816;
  assign n43818 = ~i_hlock9 & ~n43817;
  assign n43819 = ~n43806 & ~n43818;
  assign n43820 = ~controllable_hgrant4 & ~n43819;
  assign n43821 = ~n43788 & ~n43820;
  assign n43822 = ~controllable_hgrant5 & ~n43821;
  assign n43823 = ~n43780 & ~n43822;
  assign n43824 = ~controllable_hmaster2 & ~n43823;
  assign n43825 = ~n43777 & ~n43824;
  assign n43826 = ~controllable_hmaster1 & ~n43825;
  assign n43827 = ~n43776 & ~n43826;
  assign n43828 = ~controllable_hgrant6 & ~n43827;
  assign n43829 = ~n43742 & ~n43828;
  assign n43830 = controllable_hmaster0 & ~n43829;
  assign n43831 = ~n8217 & ~n20378;
  assign n43832 = ~n42153 & ~n43831;
  assign n43833 = controllable_hgrant6 & ~n43832;
  assign n43834 = ~n8378 & ~n19758;
  assign n43835 = ~n42157 & ~n43834;
  assign n43836 = controllable_hgrant5 & ~n43835;
  assign n43837 = ~n8426 & ~n19756;
  assign n43838 = ~n41584 & ~n43837;
  assign n43839 = controllable_hgrant4 & ~n43838;
  assign n43840 = ~n8365 & ~n19754;
  assign n43841 = ~n41594 & ~n43840;
  assign n43842 = controllable_hgrant3 & ~n43841;
  assign n43843 = ~n8389 & ~n19752;
  assign n43844 = ~n41598 & ~n43843;
  assign n43845 = controllable_hgrant1 & ~n43844;
  assign n43846 = ~n20613 & ~n43761;
  assign n43847 = ~n7733 & ~n43846;
  assign n43848 = ~n17505 & ~n43761;
  assign n43849 = n7733 & ~n43848;
  assign n43850 = ~n43847 & ~n43849;
  assign n43851 = n7928 & ~n43850;
  assign n43852 = ~n8221 & ~n43851;
  assign n43853 = ~controllable_hgrant1 & ~n43852;
  assign n43854 = ~n43845 & ~n43853;
  assign n43855 = ~controllable_hgrant3 & ~n43854;
  assign n43856 = ~n43842 & ~n43855;
  assign n43857 = ~controllable_hgrant4 & ~n43856;
  assign n43858 = ~n43839 & ~n43857;
  assign n43859 = ~controllable_hgrant5 & ~n43858;
  assign n43860 = ~n43836 & ~n43859;
  assign n43861 = ~controllable_hmaster2 & ~n43860;
  assign n43862 = ~n43777 & ~n43861;
  assign n43863 = ~controllable_hmaster1 & ~n43862;
  assign n43864 = ~n43776 & ~n43863;
  assign n43865 = ~controllable_hgrant6 & ~n43864;
  assign n43866 = ~n43833 & ~n43865;
  assign n43867 = ~controllable_hmaster0 & ~n43866;
  assign n43868 = ~n43830 & ~n43867;
  assign n43869 = i_hlock8 & ~n43868;
  assign n43870 = ~n8217 & ~n20387;
  assign n43871 = ~n42175 & ~n43870;
  assign n43872 = controllable_hgrant6 & ~n43871;
  assign n43873 = ~n8378 & ~n19781;
  assign n43874 = ~n42179 & ~n43873;
  assign n43875 = controllable_hgrant5 & ~n43874;
  assign n43876 = ~n8426 & ~n19779;
  assign n43877 = ~n41588 & ~n43876;
  assign n43878 = controllable_hgrant4 & ~n43877;
  assign n43879 = ~n8365 & ~n19765;
  assign n43880 = ~n41620 & ~n43879;
  assign n43881 = controllable_hgrant3 & ~n43880;
  assign n43882 = ~n8389 & ~n19763;
  assign n43883 = ~n41624 & ~n43882;
  assign n43884 = controllable_hgrant1 & ~n43883;
  assign n43885 = ~n8235 & ~n43851;
  assign n43886 = ~controllable_hgrant1 & ~n43885;
  assign n43887 = ~n43884 & ~n43886;
  assign n43888 = ~controllable_hgrant3 & ~n43887;
  assign n43889 = ~n43881 & ~n43888;
  assign n43890 = ~controllable_hgrant4 & ~n43889;
  assign n43891 = ~n43878 & ~n43890;
  assign n43892 = ~controllable_hgrant5 & ~n43891;
  assign n43893 = ~n43875 & ~n43892;
  assign n43894 = ~controllable_hmaster2 & ~n43893;
  assign n43895 = ~n43777 & ~n43894;
  assign n43896 = ~controllable_hmaster1 & ~n43895;
  assign n43897 = ~n43776 & ~n43896;
  assign n43898 = ~controllable_hgrant6 & ~n43897;
  assign n43899 = ~n43872 & ~n43898;
  assign n43900 = ~controllable_hmaster0 & ~n43899;
  assign n43901 = ~n43830 & ~n43900;
  assign n43902 = ~i_hlock8 & ~n43901;
  assign n43903 = ~n43869 & ~n43902;
  assign n43904 = controllable_hmaster3 & ~n43903;
  assign n43905 = n8217 & ~n13890;
  assign n43906 = ~n8217 & ~n19801;
  assign n43907 = ~n43905 & ~n43906;
  assign n43908 = controllable_hgrant6 & ~n43907;
  assign n43909 = controllable_hmaster2 & ~n43860;
  assign n43910 = n8378 & ~n13859;
  assign n43911 = ~n8378 & ~n19771;
  assign n43912 = ~n43910 & ~n43911;
  assign n43913 = controllable_hgrant5 & ~n43912;
  assign n43914 = n8426 & ~n13857;
  assign n43915 = ~n8426 & ~n19769;
  assign n43916 = ~n43914 & ~n43915;
  assign n43917 = controllable_hgrant4 & ~n43916;
  assign n43918 = n8365 & ~n12806;
  assign n43919 = ~n8365 & ~n19687;
  assign n43920 = ~n43918 & ~n43919;
  assign n43921 = i_hlock3 & ~n43920;
  assign n43922 = n8365 & ~n12812;
  assign n43923 = ~n8365 & ~n19693;
  assign n43924 = ~n43922 & ~n43923;
  assign n43925 = ~i_hlock3 & ~n43924;
  assign n43926 = ~n43921 & ~n43925;
  assign n43927 = controllable_hgrant3 & ~n43926;
  assign n43928 = i_hlock3 & ~n43854;
  assign n43929 = ~i_hlock3 & ~n43887;
  assign n43930 = ~n43928 & ~n43929;
  assign n43931 = ~controllable_hgrant3 & ~n43930;
  assign n43932 = ~n43927 & ~n43931;
  assign n43933 = ~controllable_hgrant4 & ~n43932;
  assign n43934 = ~n43917 & ~n43933;
  assign n43935 = ~controllable_hgrant5 & ~n43934;
  assign n43936 = ~n43913 & ~n43935;
  assign n43937 = ~controllable_hmaster2 & ~n43936;
  assign n43938 = ~n43909 & ~n43937;
  assign n43939 = controllable_hmaster1 & ~n43938;
  assign n43940 = n8378 & ~n26735;
  assign n43941 = ~n8378 & ~n29866;
  assign n43942 = ~n43940 & ~n43941;
  assign n43943 = i_hlock5 & ~n43942;
  assign n43944 = n8378 & ~n26751;
  assign n43945 = ~n8378 & ~n29881;
  assign n43946 = ~n43944 & ~n43945;
  assign n43947 = ~i_hlock5 & ~n43946;
  assign n43948 = ~n43943 & ~n43947;
  assign n43949 = controllable_hgrant5 & ~n43948;
  assign n43950 = i_hlock5 & ~n43858;
  assign n43951 = ~i_hlock5 & ~n43891;
  assign n43952 = ~n43950 & ~n43951;
  assign n43953 = ~controllable_hgrant5 & ~n43952;
  assign n43954 = ~n43949 & ~n43953;
  assign n43955 = controllable_hmaster2 & ~n43954;
  assign n43956 = n8378 & ~n13884;
  assign n43957 = ~n8378 & ~n19795;
  assign n43958 = ~n43956 & ~n43957;
  assign n43959 = controllable_hgrant5 & ~n43958;
  assign n43960 = n8426 & ~n13882;
  assign n43961 = ~n8426 & ~n19793;
  assign n43962 = ~n43960 & ~n43961;
  assign n43963 = controllable_hgrant4 & ~n43962;
  assign n43964 = n8365 & ~n13880;
  assign n43965 = ~n8365 & ~n19791;
  assign n43966 = ~n43964 & ~n43965;
  assign n43967 = controllable_hgrant3 & ~n43966;
  assign n43968 = n8389 & ~n12804;
  assign n43969 = ~n8389 & ~n19685;
  assign n43970 = ~n43968 & ~n43969;
  assign n43971 = i_hlock1 & ~n43970;
  assign n43972 = n8389 & ~n12810;
  assign n43973 = ~n8389 & ~n19691;
  assign n43974 = ~n43972 & ~n43973;
  assign n43975 = ~i_hlock1 & ~n43974;
  assign n43976 = ~n43971 & ~n43975;
  assign n43977 = controllable_hgrant1 & ~n43976;
  assign n43978 = i_hlock1 & ~n43852;
  assign n43979 = ~i_hlock1 & ~n43885;
  assign n43980 = ~n43978 & ~n43979;
  assign n43981 = ~controllable_hgrant1 & ~n43980;
  assign n43982 = ~n43977 & ~n43981;
  assign n43983 = ~controllable_hgrant3 & ~n43982;
  assign n43984 = ~n43967 & ~n43983;
  assign n43985 = ~controllable_hgrant4 & ~n43984;
  assign n43986 = ~n43963 & ~n43985;
  assign n43987 = ~controllable_hgrant5 & ~n43986;
  assign n43988 = ~n43959 & ~n43987;
  assign n43989 = ~controllable_hmaster2 & ~n43988;
  assign n43990 = ~n43955 & ~n43989;
  assign n43991 = ~controllable_hmaster1 & ~n43990;
  assign n43992 = ~n43939 & ~n43991;
  assign n43993 = ~controllable_hgrant6 & ~n43992;
  assign n43994 = ~n43908 & ~n43993;
  assign n43995 = controllable_hmaster0 & ~n43994;
  assign n43996 = ~n13908 & ~n26738;
  assign n43997 = controllable_hmaster1 & ~n43996;
  assign n43998 = ~n13936 & ~n43997;
  assign n43999 = n8217 & ~n43998;
  assign n44000 = ~n19814 & ~n29869;
  assign n44001 = controllable_hmaster1 & ~n44000;
  assign n44002 = ~n19836 & ~n44001;
  assign n44003 = ~n8217 & ~n44002;
  assign n44004 = ~n43999 & ~n44003;
  assign n44005 = i_hlock6 & ~n44004;
  assign n44006 = ~n13908 & ~n26754;
  assign n44007 = controllable_hmaster1 & ~n44006;
  assign n44008 = ~n13936 & ~n44007;
  assign n44009 = n8217 & ~n44008;
  assign n44010 = ~n19814 & ~n29884;
  assign n44011 = controllable_hmaster1 & ~n44010;
  assign n44012 = ~n19836 & ~n44011;
  assign n44013 = ~n8217 & ~n44012;
  assign n44014 = ~n44009 & ~n44013;
  assign n44015 = ~i_hlock6 & ~n44014;
  assign n44016 = ~n44005 & ~n44015;
  assign n44017 = controllable_hgrant6 & ~n44016;
  assign n44018 = n8378 & ~n13905;
  assign n44019 = ~n8378 & ~n19811;
  assign n44020 = ~n44018 & ~n44019;
  assign n44021 = controllable_hgrant5 & ~n44020;
  assign n44022 = n8426 & ~n13903;
  assign n44023 = ~n8426 & ~n19809;
  assign n44024 = ~n44022 & ~n44023;
  assign n44025 = controllable_hgrant4 & ~n44024;
  assign n44026 = n8365 & ~n13901;
  assign n44027 = ~n8365 & ~n19807;
  assign n44028 = ~n44026 & ~n44027;
  assign n44029 = controllable_hgrant3 & ~n44028;
  assign n44030 = n8389 & ~n13899;
  assign n44031 = ~n8389 & ~n19805;
  assign n44032 = ~n44030 & ~n44031;
  assign n44033 = controllable_hgrant1 & ~n44032;
  assign n44034 = ~n42967 & ~n43759;
  assign n44035 = controllable_hgrant2 & ~n44034;
  assign n44036 = ~n20613 & ~n44035;
  assign n44037 = ~n7733 & ~n44036;
  assign n44038 = ~n17505 & ~n44035;
  assign n44039 = n7733 & ~n44038;
  assign n44040 = ~n44037 & ~n44039;
  assign n44041 = n7928 & ~n44040;
  assign n44042 = ~n42965 & ~n44041;
  assign n44043 = ~controllable_hgrant1 & ~n44042;
  assign n44044 = ~n44033 & ~n44043;
  assign n44045 = ~controllable_hgrant3 & ~n44044;
  assign n44046 = ~n44029 & ~n44045;
  assign n44047 = ~controllable_hgrant4 & ~n44046;
  assign n44048 = ~n44025 & ~n44047;
  assign n44049 = ~controllable_hgrant5 & ~n44048;
  assign n44050 = ~n44021 & ~n44049;
  assign n44051 = ~controllable_hmaster2 & ~n44050;
  assign n44052 = ~n43909 & ~n44051;
  assign n44053 = controllable_hmaster1 & ~n44052;
  assign n44054 = n8378 & ~n13917;
  assign n44055 = ~n8378 & ~n19821;
  assign n44056 = ~n44054 & ~n44055;
  assign n44057 = controllable_hgrant5 & ~n44056;
  assign n44058 = n8426 & ~n12808;
  assign n44059 = ~n8426 & ~n19689;
  assign n44060 = ~n44058 & ~n44059;
  assign n44061 = i_hlock4 & ~n44060;
  assign n44062 = n8426 & ~n12814;
  assign n44063 = ~n8426 & ~n19695;
  assign n44064 = ~n44062 & ~n44063;
  assign n44065 = ~i_hlock4 & ~n44064;
  assign n44066 = ~n44061 & ~n44065;
  assign n44067 = controllable_hgrant4 & ~n44066;
  assign n44068 = i_hlock4 & ~n43856;
  assign n44069 = ~i_hlock4 & ~n43889;
  assign n44070 = ~n44068 & ~n44069;
  assign n44071 = ~controllable_hgrant4 & ~n44070;
  assign n44072 = ~n44067 & ~n44071;
  assign n44073 = ~controllable_hgrant5 & ~n44072;
  assign n44074 = ~n44057 & ~n44073;
  assign n44075 = controllable_hmaster2 & ~n44074;
  assign n44076 = n8378 & ~n13931;
  assign n44077 = ~n8378 & ~n19831;
  assign n44078 = ~n44076 & ~n44077;
  assign n44079 = controllable_hgrant5 & ~n44078;
  assign n44080 = n8426 & ~n13929;
  assign n44081 = ~n8426 & ~n19829;
  assign n44082 = ~n44080 & ~n44081;
  assign n44083 = controllable_hgrant4 & ~n44082;
  assign n44084 = n8365 & ~n13927;
  assign n44085 = ~n8365 & ~n19827;
  assign n44086 = ~n44084 & ~n44085;
  assign n44087 = controllable_hgrant3 & ~n44086;
  assign n44088 = n8389 & ~n13925;
  assign n44089 = ~n8389 & ~n19825;
  assign n44090 = ~n44088 & ~n44089;
  assign n44091 = controllable_hgrant1 & ~n44090;
  assign n44092 = ~n8440 & ~n43851;
  assign n44093 = ~controllable_hgrant1 & ~n44092;
  assign n44094 = ~n44091 & ~n44093;
  assign n44095 = ~controllable_hgrant3 & ~n44094;
  assign n44096 = ~n44087 & ~n44095;
  assign n44097 = ~controllable_hgrant4 & ~n44096;
  assign n44098 = ~n44083 & ~n44097;
  assign n44099 = ~controllable_hgrant5 & ~n44098;
  assign n44100 = ~n44079 & ~n44099;
  assign n44101 = ~controllable_hmaster2 & ~n44100;
  assign n44102 = ~n44075 & ~n44101;
  assign n44103 = ~controllable_hmaster1 & ~n44102;
  assign n44104 = ~n44053 & ~n44103;
  assign n44105 = i_hlock6 & ~n44104;
  assign n44106 = controllable_hmaster2 & ~n43893;
  assign n44107 = ~n44051 & ~n44106;
  assign n44108 = controllable_hmaster1 & ~n44107;
  assign n44109 = ~n44103 & ~n44108;
  assign n44110 = ~i_hlock6 & ~n44109;
  assign n44111 = ~n44105 & ~n44110;
  assign n44112 = ~controllable_hgrant6 & ~n44111;
  assign n44113 = ~n44017 & ~n44112;
  assign n44114 = ~controllable_hmaster0 & ~n44113;
  assign n44115 = ~n43995 & ~n44114;
  assign n44116 = ~controllable_hmaster3 & ~n44115;
  assign n44117 = ~n43904 & ~n44116;
  assign n44118 = i_hlock7 & ~n44117;
  assign n44119 = n8217 & ~n13954;
  assign n44120 = ~n8217 & ~n19856;
  assign n44121 = ~n44119 & ~n44120;
  assign n44122 = controllable_hgrant6 & ~n44121;
  assign n44123 = ~n43937 & ~n44106;
  assign n44124 = controllable_hmaster1 & ~n44123;
  assign n44125 = ~n43991 & ~n44124;
  assign n44126 = ~controllable_hgrant6 & ~n44125;
  assign n44127 = ~n44122 & ~n44126;
  assign n44128 = controllable_hmaster0 & ~n44127;
  assign n44129 = ~n44114 & ~n44128;
  assign n44130 = ~controllable_hmaster3 & ~n44129;
  assign n44131 = ~n43904 & ~n44130;
  assign n44132 = ~i_hlock7 & ~n44131;
  assign n44133 = ~n44118 & ~n44132;
  assign n44134 = i_hbusreq7 & ~n44133;
  assign n44135 = i_hbusreq8 & ~n43903;
  assign n44136 = i_hbusreq6 & ~n43741;
  assign n44137 = n8217 & ~n27317;
  assign n44138 = ~n8217 & ~n29918;
  assign n44139 = ~n44137 & ~n44138;
  assign n44140 = ~i_hbusreq6 & ~n44139;
  assign n44141 = ~n44136 & ~n44140;
  assign n44142 = controllable_hgrant6 & ~n44141;
  assign n44143 = i_hbusreq6 & ~n43827;
  assign n44144 = i_hbusreq5 & ~n43745;
  assign n44145 = n8378 & ~n14395;
  assign n44146 = ~n8378 & ~n19889;
  assign n44147 = ~n44145 & ~n44146;
  assign n44148 = ~i_hbusreq5 & ~n44147;
  assign n44149 = ~n44144 & ~n44148;
  assign n44150 = controllable_hgrant5 & ~n44149;
  assign n44151 = i_hbusreq5 & ~n43773;
  assign n44152 = i_hbusreq4 & ~n43749;
  assign n44153 = i_hbusreq9 & ~n43749;
  assign n44154 = n8426 & ~n14389;
  assign n44155 = ~n8426 & ~n19883;
  assign n44156 = ~n44154 & ~n44155;
  assign n44157 = ~i_hbusreq9 & ~n44156;
  assign n44158 = ~n44153 & ~n44157;
  assign n44159 = ~i_hbusreq4 & ~n44158;
  assign n44160 = ~n44152 & ~n44159;
  assign n44161 = controllable_hgrant4 & ~n44160;
  assign n44162 = i_hbusreq4 & ~n43771;
  assign n44163 = i_hbusreq9 & ~n43771;
  assign n44164 = i_hbusreq3 & ~n43753;
  assign n44165 = n8365 & ~n14385;
  assign n44166 = ~n8365 & ~n19879;
  assign n44167 = ~n44165 & ~n44166;
  assign n44168 = ~i_hbusreq3 & ~n44167;
  assign n44169 = ~n44164 & ~n44168;
  assign n44170 = controllable_hgrant3 & ~n44169;
  assign n44171 = i_hbusreq3 & ~n43769;
  assign n44172 = i_hbusreq1 & ~n43757;
  assign n44173 = n8389 & ~n14381;
  assign n44174 = ~n8389 & ~n19875;
  assign n44175 = ~n44173 & ~n44174;
  assign n44176 = ~i_hbusreq1 & ~n44175;
  assign n44177 = ~n44172 & ~n44176;
  assign n44178 = controllable_hgrant1 & ~n44177;
  assign n44179 = i_hbusreq1 & ~n43767;
  assign n44180 = i_hbusreq2 & ~n43760;
  assign n44181 = i_hbusreq0 & ~n43760;
  assign n44182 = ~controllable_locked & ~n39847;
  assign n44183 = ~controllable_locked & ~n44182;
  assign n44184 = i_hlock0 & ~n44183;
  assign n44185 = ~i_hlock0 & ~n43760;
  assign n44186 = ~n44184 & ~n44185;
  assign n44187 = ~i_hbusreq0 & ~n44186;
  assign n44188 = ~n44181 & ~n44187;
  assign n44189 = ~i_hbusreq2 & ~n44188;
  assign n44190 = ~n44180 & ~n44189;
  assign n44191 = controllable_hgrant2 & ~n44190;
  assign n44192 = ~n16639 & ~n40869;
  assign n44193 = ~i_hbusreq0 & ~n44192;
  assign n44194 = ~i_hbusreq0 & ~n44193;
  assign n44195 = ~i_hbusreq2 & ~n44194;
  assign n44196 = ~i_hbusreq2 & ~n44195;
  assign n44197 = ~controllable_hgrant2 & n44196;
  assign n44198 = ~n44191 & ~n44197;
  assign n44199 = ~n7733 & ~n44198;
  assign n44200 = ~n16633 & ~n44191;
  assign n44201 = n7733 & ~n44200;
  assign n44202 = ~n44199 & ~n44201;
  assign n44203 = n7928 & ~n44202;
  assign n44204 = ~n43114 & ~n44203;
  assign n44205 = ~i_hbusreq1 & ~n44204;
  assign n44206 = ~n44179 & ~n44205;
  assign n44207 = ~controllable_hgrant1 & ~n44206;
  assign n44208 = ~n44178 & ~n44207;
  assign n44209 = ~i_hbusreq3 & ~n44208;
  assign n44210 = ~n44171 & ~n44209;
  assign n44211 = ~controllable_hgrant3 & ~n44210;
  assign n44212 = ~n44170 & ~n44211;
  assign n44213 = ~i_hbusreq9 & ~n44212;
  assign n44214 = ~n44163 & ~n44213;
  assign n44215 = ~i_hbusreq4 & ~n44214;
  assign n44216 = ~n44162 & ~n44215;
  assign n44217 = ~controllable_hgrant4 & ~n44216;
  assign n44218 = ~n44161 & ~n44217;
  assign n44219 = ~i_hbusreq5 & ~n44218;
  assign n44220 = ~n44151 & ~n44219;
  assign n44221 = ~controllable_hgrant5 & ~n44220;
  assign n44222 = ~n44150 & ~n44221;
  assign n44223 = controllable_hmaster1 & ~n44222;
  assign n44224 = controllable_hmaster2 & ~n44222;
  assign n44225 = i_hbusreq5 & ~n43779;
  assign n44226 = n8378 & ~n27309;
  assign n44227 = ~n8378 & ~n29910;
  assign n44228 = ~n44226 & ~n44227;
  assign n44229 = ~i_hbusreq5 & ~n44228;
  assign n44230 = ~n44225 & ~n44229;
  assign n44231 = controllable_hgrant5 & ~n44230;
  assign n44232 = i_hbusreq5 & ~n43821;
  assign n44233 = i_hbusreq4 & ~n43787;
  assign n44234 = i_hbusreq9 & ~n43787;
  assign n44235 = n8426 & ~n14462;
  assign n44236 = ~n8426 & ~n19974;
  assign n44237 = ~n44235 & ~n44236;
  assign n44238 = i_hlock9 & ~n44237;
  assign n44239 = n8426 & ~n14493;
  assign n44240 = ~n8426 & ~n20010;
  assign n44241 = ~n44239 & ~n44240;
  assign n44242 = ~i_hlock9 & ~n44241;
  assign n44243 = ~n44238 & ~n44242;
  assign n44244 = ~i_hbusreq9 & ~n44243;
  assign n44245 = ~n44234 & ~n44244;
  assign n44246 = ~i_hbusreq4 & ~n44245;
  assign n44247 = ~n44233 & ~n44246;
  assign n44248 = controllable_hgrant4 & ~n44247;
  assign n44249 = i_hbusreq4 & ~n43819;
  assign n44250 = i_hbusreq9 & ~n43819;
  assign n44251 = i_hbusreq3 & ~n43790;
  assign n44252 = n8365 & ~n14458;
  assign n44253 = ~n8365 & ~n19970;
  assign n44254 = ~n44252 & ~n44253;
  assign n44255 = ~i_hbusreq3 & ~n44254;
  assign n44256 = ~n44251 & ~n44255;
  assign n44257 = controllable_hgrant3 & ~n44256;
  assign n44258 = i_hbusreq3 & ~n43803;
  assign n44259 = i_hbusreq1 & ~n43793;
  assign n44260 = n8389 & ~n14454;
  assign n44261 = ~n8389 & ~n19966;
  assign n44262 = ~n44260 & ~n44261;
  assign n44263 = ~i_hbusreq1 & ~n44262;
  assign n44264 = ~n44259 & ~n44263;
  assign n44265 = controllable_hgrant1 & ~n44264;
  assign n44266 = i_hbusreq1 & ~n43801;
  assign n44267 = controllable_locked & ~n12782;
  assign n44268 = controllable_locked & ~n44267;
  assign n44269 = ~i_hlock0 & ~n44268;
  assign n44270 = ~n40869 & ~n44269;
  assign n44271 = ~i_hbusreq0 & ~n44270;
  assign n44272 = ~i_hbusreq0 & ~n44271;
  assign n44273 = ~i_hbusreq2 & ~n44272;
  assign n44274 = ~i_hbusreq2 & ~n44273;
  assign n44275 = ~controllable_hgrant2 & n44274;
  assign n44276 = ~n44191 & ~n44275;
  assign n44277 = ~n7733 & ~n44276;
  assign n44278 = i_hbusreq2 & ~n43795;
  assign n44279 = i_hbusreq0 & ~n43795;
  assign n44280 = ~n7734 & ~n39846;
  assign n44281 = ~controllable_hmastlock & ~n44280;
  assign n44282 = ~n39853 & ~n44281;
  assign n44283 = ~controllable_locked & ~n44282;
  assign n44284 = ~n40336 & ~n44283;
  assign n44285 = i_hlock0 & ~n44284;
  assign n44286 = ~i_hlock0 & ~n43795;
  assign n44287 = ~n44285 & ~n44286;
  assign n44288 = ~i_hbusreq0 & ~n44287;
  assign n44289 = ~n44279 & ~n44288;
  assign n44290 = ~i_hbusreq2 & ~n44289;
  assign n44291 = ~n44278 & ~n44290;
  assign n44292 = controllable_hgrant2 & ~n44291;
  assign n44293 = controllable_locked & ~n16803;
  assign n44294 = ~n19952 & ~n44293;
  assign n44295 = i_hlock0 & ~n44294;
  assign n44296 = ~n18716 & ~n44295;
  assign n44297 = ~i_hbusreq0 & ~n44296;
  assign n44298 = ~n17142 & ~n44297;
  assign n44299 = ~i_hbusreq2 & ~n44298;
  assign n44300 = ~n17141 & ~n44299;
  assign n44301 = ~controllable_hgrant2 & ~n44300;
  assign n44302 = ~n44292 & ~n44301;
  assign n44303 = n7733 & ~n44302;
  assign n44304 = ~n44277 & ~n44303;
  assign n44305 = n7928 & ~n44304;
  assign n44306 = ~n8265 & ~n44305;
  assign n44307 = ~i_hbusreq1 & ~n44306;
  assign n44308 = ~n44266 & ~n44307;
  assign n44309 = ~controllable_hgrant1 & ~n44308;
  assign n44310 = ~n44265 & ~n44309;
  assign n44311 = ~i_hbusreq3 & ~n44310;
  assign n44312 = ~n44258 & ~n44311;
  assign n44313 = ~controllable_hgrant3 & ~n44312;
  assign n44314 = ~n44257 & ~n44313;
  assign n44315 = i_hlock9 & ~n44314;
  assign n44316 = i_hbusreq3 & ~n43808;
  assign n44317 = n8365 & ~n14489;
  assign n44318 = ~n8365 & ~n20006;
  assign n44319 = ~n44317 & ~n44318;
  assign n44320 = ~i_hbusreq3 & ~n44319;
  assign n44321 = ~n44316 & ~n44320;
  assign n44322 = controllable_hgrant3 & ~n44321;
  assign n44323 = i_hbusreq3 & ~n43815;
  assign n44324 = i_hbusreq1 & ~n43811;
  assign n44325 = n8389 & ~n14485;
  assign n44326 = ~n8389 & ~n20002;
  assign n44327 = ~n44325 & ~n44326;
  assign n44328 = ~i_hbusreq1 & ~n44327;
  assign n44329 = ~n44324 & ~n44328;
  assign n44330 = controllable_hgrant1 & ~n44329;
  assign n44331 = i_hbusreq1 & ~n43813;
  assign n44332 = ~n8297 & ~n44305;
  assign n44333 = ~i_hbusreq1 & ~n44332;
  assign n44334 = ~n44331 & ~n44333;
  assign n44335 = ~controllable_hgrant1 & ~n44334;
  assign n44336 = ~n44330 & ~n44335;
  assign n44337 = ~i_hbusreq3 & ~n44336;
  assign n44338 = ~n44323 & ~n44337;
  assign n44339 = ~controllable_hgrant3 & ~n44338;
  assign n44340 = ~n44322 & ~n44339;
  assign n44341 = ~i_hlock9 & ~n44340;
  assign n44342 = ~n44315 & ~n44341;
  assign n44343 = ~i_hbusreq9 & ~n44342;
  assign n44344 = ~n44250 & ~n44343;
  assign n44345 = ~i_hbusreq4 & ~n44344;
  assign n44346 = ~n44249 & ~n44345;
  assign n44347 = ~controllable_hgrant4 & ~n44346;
  assign n44348 = ~n44248 & ~n44347;
  assign n44349 = ~i_hbusreq5 & ~n44348;
  assign n44350 = ~n44232 & ~n44349;
  assign n44351 = ~controllable_hgrant5 & ~n44350;
  assign n44352 = ~n44231 & ~n44351;
  assign n44353 = ~controllable_hmaster2 & ~n44352;
  assign n44354 = ~n44224 & ~n44353;
  assign n44355 = ~controllable_hmaster1 & ~n44354;
  assign n44356 = ~n44223 & ~n44355;
  assign n44357 = ~i_hbusreq6 & ~n44356;
  assign n44358 = ~n44143 & ~n44357;
  assign n44359 = ~controllable_hgrant6 & ~n44358;
  assign n44360 = ~n44142 & ~n44359;
  assign n44361 = controllable_hmaster0 & ~n44360;
  assign n44362 = i_hbusreq6 & ~n43832;
  assign n44363 = n8217 & ~n14733;
  assign n44364 = ~n8217 & ~n20424;
  assign n44365 = ~n44363 & ~n44364;
  assign n44366 = ~i_hbusreq6 & ~n44365;
  assign n44367 = ~n44362 & ~n44366;
  assign n44368 = controllable_hgrant6 & ~n44367;
  assign n44369 = i_hbusreq6 & ~n43864;
  assign n44370 = i_hbusreq5 & ~n43835;
  assign n44371 = n8378 & ~n14533;
  assign n44372 = ~n8378 & ~n20057;
  assign n44373 = ~n44371 & ~n44372;
  assign n44374 = ~i_hbusreq5 & ~n44373;
  assign n44375 = ~n44370 & ~n44374;
  assign n44376 = controllable_hgrant5 & ~n44375;
  assign n44377 = i_hbusreq5 & ~n43858;
  assign n44378 = i_hbusreq4 & ~n43838;
  assign n44379 = i_hbusreq9 & ~n43838;
  assign n44380 = n8426 & ~n14527;
  assign n44381 = ~n8426 & ~n20051;
  assign n44382 = ~n44380 & ~n44381;
  assign n44383 = ~i_hbusreq9 & ~n44382;
  assign n44384 = ~n44379 & ~n44383;
  assign n44385 = ~i_hbusreq4 & ~n44384;
  assign n44386 = ~n44378 & ~n44385;
  assign n44387 = controllable_hgrant4 & ~n44386;
  assign n44388 = i_hbusreq4 & ~n43856;
  assign n44389 = i_hbusreq9 & ~n43856;
  assign n44390 = i_hbusreq3 & ~n43841;
  assign n44391 = n8365 & ~n14523;
  assign n44392 = ~n8365 & ~n20047;
  assign n44393 = ~n44391 & ~n44392;
  assign n44394 = ~i_hbusreq3 & ~n44393;
  assign n44395 = ~n44390 & ~n44394;
  assign n44396 = controllable_hgrant3 & ~n44395;
  assign n44397 = i_hbusreq3 & ~n43854;
  assign n44398 = i_hbusreq1 & ~n43844;
  assign n44399 = n8389 & ~n14519;
  assign n44400 = ~n8389 & ~n20043;
  assign n44401 = ~n44399 & ~n44400;
  assign n44402 = ~i_hbusreq1 & ~n44401;
  assign n44403 = ~n44398 & ~n44402;
  assign n44404 = controllable_hgrant1 & ~n44403;
  assign n44405 = i_hbusreq1 & ~n43852;
  assign n44406 = ~n20882 & ~n44191;
  assign n44407 = ~n7733 & ~n44406;
  assign n44408 = ~n18798 & ~n44191;
  assign n44409 = n7733 & ~n44408;
  assign n44410 = ~n44407 & ~n44409;
  assign n44411 = n7928 & ~n44410;
  assign n44412 = ~n8265 & ~n44411;
  assign n44413 = ~i_hbusreq1 & ~n44412;
  assign n44414 = ~n44405 & ~n44413;
  assign n44415 = ~controllable_hgrant1 & ~n44414;
  assign n44416 = ~n44404 & ~n44415;
  assign n44417 = ~i_hbusreq3 & ~n44416;
  assign n44418 = ~n44397 & ~n44417;
  assign n44419 = ~controllable_hgrant3 & ~n44418;
  assign n44420 = ~n44396 & ~n44419;
  assign n44421 = ~i_hbusreq9 & ~n44420;
  assign n44422 = ~n44389 & ~n44421;
  assign n44423 = ~i_hbusreq4 & ~n44422;
  assign n44424 = ~n44388 & ~n44423;
  assign n44425 = ~controllable_hgrant4 & ~n44424;
  assign n44426 = ~n44387 & ~n44425;
  assign n44427 = ~i_hbusreq5 & ~n44426;
  assign n44428 = ~n44377 & ~n44427;
  assign n44429 = ~controllable_hgrant5 & ~n44428;
  assign n44430 = ~n44376 & ~n44429;
  assign n44431 = ~controllable_hmaster2 & ~n44430;
  assign n44432 = ~n44224 & ~n44431;
  assign n44433 = ~controllable_hmaster1 & ~n44432;
  assign n44434 = ~n44223 & ~n44433;
  assign n44435 = ~i_hbusreq6 & ~n44434;
  assign n44436 = ~n44369 & ~n44435;
  assign n44437 = ~controllable_hgrant6 & ~n44436;
  assign n44438 = ~n44368 & ~n44437;
  assign n44439 = ~controllable_hmaster0 & ~n44438;
  assign n44440 = ~n44361 & ~n44439;
  assign n44441 = i_hlock8 & ~n44440;
  assign n44442 = i_hbusreq6 & ~n43871;
  assign n44443 = n8217 & ~n14744;
  assign n44444 = ~n8217 & ~n20436;
  assign n44445 = ~n44443 & ~n44444;
  assign n44446 = ~i_hbusreq6 & ~n44445;
  assign n44447 = ~n44442 & ~n44446;
  assign n44448 = controllable_hgrant6 & ~n44447;
  assign n44449 = i_hbusreq6 & ~n43897;
  assign n44450 = i_hbusreq5 & ~n43874;
  assign n44451 = n8378 & ~n14574;
  assign n44452 = ~n8378 & ~n20107;
  assign n44453 = ~n44451 & ~n44452;
  assign n44454 = ~i_hbusreq5 & ~n44453;
  assign n44455 = ~n44450 & ~n44454;
  assign n44456 = controllable_hgrant5 & ~n44455;
  assign n44457 = i_hbusreq5 & ~n43891;
  assign n44458 = i_hbusreq4 & ~n43877;
  assign n44459 = i_hbusreq9 & ~n43877;
  assign n44460 = n8426 & ~n14568;
  assign n44461 = ~n8426 & ~n20101;
  assign n44462 = ~n44460 & ~n44461;
  assign n44463 = ~i_hbusreq9 & ~n44462;
  assign n44464 = ~n44459 & ~n44463;
  assign n44465 = ~i_hbusreq4 & ~n44464;
  assign n44466 = ~n44458 & ~n44465;
  assign n44467 = controllable_hgrant4 & ~n44466;
  assign n44468 = i_hbusreq4 & ~n43889;
  assign n44469 = i_hbusreq9 & ~n43889;
  assign n44470 = i_hbusreq3 & ~n43880;
  assign n44471 = n8365 & ~n14544;
  assign n44472 = ~n8365 & ~n20073;
  assign n44473 = ~n44471 & ~n44472;
  assign n44474 = ~i_hbusreq3 & ~n44473;
  assign n44475 = ~n44470 & ~n44474;
  assign n44476 = controllable_hgrant3 & ~n44475;
  assign n44477 = i_hbusreq3 & ~n43887;
  assign n44478 = i_hbusreq1 & ~n43883;
  assign n44479 = n8389 & ~n14540;
  assign n44480 = ~n8389 & ~n20069;
  assign n44481 = ~n44479 & ~n44480;
  assign n44482 = ~i_hbusreq1 & ~n44481;
  assign n44483 = ~n44478 & ~n44482;
  assign n44484 = controllable_hgrant1 & ~n44483;
  assign n44485 = i_hbusreq1 & ~n43885;
  assign n44486 = ~n8297 & ~n44411;
  assign n44487 = ~i_hbusreq1 & ~n44486;
  assign n44488 = ~n44485 & ~n44487;
  assign n44489 = ~controllable_hgrant1 & ~n44488;
  assign n44490 = ~n44484 & ~n44489;
  assign n44491 = ~i_hbusreq3 & ~n44490;
  assign n44492 = ~n44477 & ~n44491;
  assign n44493 = ~controllable_hgrant3 & ~n44492;
  assign n44494 = ~n44476 & ~n44493;
  assign n44495 = ~i_hbusreq9 & ~n44494;
  assign n44496 = ~n44469 & ~n44495;
  assign n44497 = ~i_hbusreq4 & ~n44496;
  assign n44498 = ~n44468 & ~n44497;
  assign n44499 = ~controllable_hgrant4 & ~n44498;
  assign n44500 = ~n44467 & ~n44499;
  assign n44501 = ~i_hbusreq5 & ~n44500;
  assign n44502 = ~n44457 & ~n44501;
  assign n44503 = ~controllable_hgrant5 & ~n44502;
  assign n44504 = ~n44456 & ~n44503;
  assign n44505 = ~controllable_hmaster2 & ~n44504;
  assign n44506 = ~n44224 & ~n44505;
  assign n44507 = ~controllable_hmaster1 & ~n44506;
  assign n44508 = ~n44223 & ~n44507;
  assign n44509 = ~i_hbusreq6 & ~n44508;
  assign n44510 = ~n44449 & ~n44509;
  assign n44511 = ~controllable_hgrant6 & ~n44510;
  assign n44512 = ~n44448 & ~n44511;
  assign n44513 = ~controllable_hmaster0 & ~n44512;
  assign n44514 = ~n44361 & ~n44513;
  assign n44515 = ~i_hlock8 & ~n44514;
  assign n44516 = ~n44441 & ~n44515;
  assign n44517 = ~i_hbusreq8 & ~n44516;
  assign n44518 = ~n44135 & ~n44517;
  assign n44519 = controllable_hmaster3 & ~n44518;
  assign n44520 = i_hbusreq8 & ~n44115;
  assign n44521 = i_hbusreq6 & ~n43907;
  assign n44522 = n8217 & ~n14606;
  assign n44523 = ~n8217 & ~n20144;
  assign n44524 = ~n44522 & ~n44523;
  assign n44525 = ~i_hbusreq6 & ~n44524;
  assign n44526 = ~n44521 & ~n44525;
  assign n44527 = controllable_hgrant6 & ~n44526;
  assign n44528 = i_hbusreq6 & ~n43992;
  assign n44529 = controllable_hmaster2 & ~n44430;
  assign n44530 = i_hbusreq5 & ~n43912;
  assign n44531 = n8378 & ~n14556;
  assign n44532 = ~n8378 & ~n20085;
  assign n44533 = ~n44531 & ~n44532;
  assign n44534 = ~i_hbusreq5 & ~n44533;
  assign n44535 = ~n44530 & ~n44534;
  assign n44536 = controllable_hgrant5 & ~n44535;
  assign n44537 = i_hbusreq5 & ~n43934;
  assign n44538 = i_hbusreq4 & ~n43916;
  assign n44539 = i_hbusreq9 & ~n43916;
  assign n44540 = n8426 & ~n14550;
  assign n44541 = ~n8426 & ~n20079;
  assign n44542 = ~n44540 & ~n44541;
  assign n44543 = ~i_hbusreq9 & ~n44542;
  assign n44544 = ~n44539 & ~n44543;
  assign n44545 = ~i_hbusreq4 & ~n44544;
  assign n44546 = ~n44538 & ~n44545;
  assign n44547 = controllable_hgrant4 & ~n44546;
  assign n44548 = i_hbusreq4 & ~n43932;
  assign n44549 = i_hbusreq9 & ~n43932;
  assign n44550 = i_hbusreq3 & ~n43926;
  assign n44551 = n8365 & ~n14407;
  assign n44552 = ~n8365 & ~n19906;
  assign n44553 = ~n44551 & ~n44552;
  assign n44554 = i_hlock3 & ~n44553;
  assign n44555 = n8365 & ~n14417;
  assign n44556 = ~n8365 & ~n19918;
  assign n44557 = ~n44555 & ~n44556;
  assign n44558 = ~i_hlock3 & ~n44557;
  assign n44559 = ~n44554 & ~n44558;
  assign n44560 = ~i_hbusreq3 & ~n44559;
  assign n44561 = ~n44550 & ~n44560;
  assign n44562 = controllable_hgrant3 & ~n44561;
  assign n44563 = i_hbusreq3 & ~n43930;
  assign n44564 = i_hlock3 & ~n44416;
  assign n44565 = ~i_hlock3 & ~n44490;
  assign n44566 = ~n44564 & ~n44565;
  assign n44567 = ~i_hbusreq3 & ~n44566;
  assign n44568 = ~n44563 & ~n44567;
  assign n44569 = ~controllable_hgrant3 & ~n44568;
  assign n44570 = ~n44562 & ~n44569;
  assign n44571 = ~i_hbusreq9 & ~n44570;
  assign n44572 = ~n44549 & ~n44571;
  assign n44573 = ~i_hbusreq4 & ~n44572;
  assign n44574 = ~n44548 & ~n44573;
  assign n44575 = ~controllable_hgrant4 & ~n44574;
  assign n44576 = ~n44547 & ~n44575;
  assign n44577 = ~i_hbusreq5 & ~n44576;
  assign n44578 = ~n44537 & ~n44577;
  assign n44579 = ~controllable_hgrant5 & ~n44578;
  assign n44580 = ~n44536 & ~n44579;
  assign n44581 = ~controllable_hmaster2 & ~n44580;
  assign n44582 = ~n44529 & ~n44581;
  assign n44583 = controllable_hmaster1 & ~n44582;
  assign n44584 = i_hbusreq5 & ~n43948;
  assign n44585 = n8378 & ~n27338;
  assign n44586 = ~n8378 & ~n29942;
  assign n44587 = ~n44585 & ~n44586;
  assign n44588 = i_hlock5 & ~n44587;
  assign n44589 = n8378 & ~n27365;
  assign n44590 = ~n8378 & ~n29972;
  assign n44591 = ~n44589 & ~n44590;
  assign n44592 = ~i_hlock5 & ~n44591;
  assign n44593 = ~n44588 & ~n44592;
  assign n44594 = ~i_hbusreq5 & ~n44593;
  assign n44595 = ~n44584 & ~n44594;
  assign n44596 = controllable_hgrant5 & ~n44595;
  assign n44597 = i_hbusreq5 & ~n43952;
  assign n44598 = i_hlock5 & ~n44426;
  assign n44599 = ~i_hlock5 & ~n44500;
  assign n44600 = ~n44598 & ~n44599;
  assign n44601 = ~i_hbusreq5 & ~n44600;
  assign n44602 = ~n44597 & ~n44601;
  assign n44603 = ~controllable_hgrant5 & ~n44602;
  assign n44604 = ~n44596 & ~n44603;
  assign n44605 = controllable_hmaster2 & ~n44604;
  assign n44606 = i_hbusreq5 & ~n43958;
  assign n44607 = n8378 & ~n14598;
  assign n44608 = ~n8378 & ~n20136;
  assign n44609 = ~n44607 & ~n44608;
  assign n44610 = ~i_hbusreq5 & ~n44609;
  assign n44611 = ~n44606 & ~n44610;
  assign n44612 = controllable_hgrant5 & ~n44611;
  assign n44613 = i_hbusreq5 & ~n43986;
  assign n44614 = i_hbusreq4 & ~n43962;
  assign n44615 = i_hbusreq9 & ~n43962;
  assign n44616 = n8426 & ~n14592;
  assign n44617 = ~n8426 & ~n20130;
  assign n44618 = ~n44616 & ~n44617;
  assign n44619 = ~i_hbusreq9 & ~n44618;
  assign n44620 = ~n44615 & ~n44619;
  assign n44621 = ~i_hbusreq4 & ~n44620;
  assign n44622 = ~n44614 & ~n44621;
  assign n44623 = controllable_hgrant4 & ~n44622;
  assign n44624 = i_hbusreq4 & ~n43984;
  assign n44625 = i_hbusreq9 & ~n43984;
  assign n44626 = i_hbusreq3 & ~n43966;
  assign n44627 = n8365 & ~n14588;
  assign n44628 = ~n8365 & ~n20126;
  assign n44629 = ~n44627 & ~n44628;
  assign n44630 = ~i_hbusreq3 & ~n44629;
  assign n44631 = ~n44626 & ~n44630;
  assign n44632 = controllable_hgrant3 & ~n44631;
  assign n44633 = i_hbusreq3 & ~n43982;
  assign n44634 = i_hbusreq1 & ~n43976;
  assign n44635 = n8389 & ~n14403;
  assign n44636 = ~n8389 & ~n19902;
  assign n44637 = ~n44635 & ~n44636;
  assign n44638 = i_hlock1 & ~n44637;
  assign n44639 = n8389 & ~n14413;
  assign n44640 = ~n8389 & ~n19914;
  assign n44641 = ~n44639 & ~n44640;
  assign n44642 = ~i_hlock1 & ~n44641;
  assign n44643 = ~n44638 & ~n44642;
  assign n44644 = ~i_hbusreq1 & ~n44643;
  assign n44645 = ~n44634 & ~n44644;
  assign n44646 = controllable_hgrant1 & ~n44645;
  assign n44647 = i_hbusreq1 & ~n43980;
  assign n44648 = i_hlock1 & ~n44412;
  assign n44649 = ~i_hlock1 & ~n44486;
  assign n44650 = ~n44648 & ~n44649;
  assign n44651 = ~i_hbusreq1 & ~n44650;
  assign n44652 = ~n44647 & ~n44651;
  assign n44653 = ~controllable_hgrant1 & ~n44652;
  assign n44654 = ~n44646 & ~n44653;
  assign n44655 = ~i_hbusreq3 & ~n44654;
  assign n44656 = ~n44633 & ~n44655;
  assign n44657 = ~controllable_hgrant3 & ~n44656;
  assign n44658 = ~n44632 & ~n44657;
  assign n44659 = ~i_hbusreq9 & ~n44658;
  assign n44660 = ~n44625 & ~n44659;
  assign n44661 = ~i_hbusreq4 & ~n44660;
  assign n44662 = ~n44624 & ~n44661;
  assign n44663 = ~controllable_hgrant4 & ~n44662;
  assign n44664 = ~n44623 & ~n44663;
  assign n44665 = ~i_hbusreq5 & ~n44664;
  assign n44666 = ~n44613 & ~n44665;
  assign n44667 = ~controllable_hgrant5 & ~n44666;
  assign n44668 = ~n44612 & ~n44667;
  assign n44669 = ~controllable_hmaster2 & ~n44668;
  assign n44670 = ~n44605 & ~n44669;
  assign n44671 = ~controllable_hmaster1 & ~n44670;
  assign n44672 = ~n44583 & ~n44671;
  assign n44673 = ~i_hbusreq6 & ~n44672;
  assign n44674 = ~n44528 & ~n44673;
  assign n44675 = ~controllable_hgrant6 & ~n44674;
  assign n44676 = ~n44527 & ~n44675;
  assign n44677 = controllable_hmaster0 & ~n44676;
  assign n44678 = i_hbusreq6 & ~n44016;
  assign n44679 = ~n14631 & ~n27343;
  assign n44680 = controllable_hmaster1 & ~n44679;
  assign n44681 = ~n14668 & ~n44680;
  assign n44682 = n8217 & ~n44681;
  assign n44683 = ~n20175 & ~n29947;
  assign n44684 = controllable_hmaster1 & ~n44683;
  assign n44685 = ~n20219 & ~n44684;
  assign n44686 = ~n8217 & ~n44685;
  assign n44687 = ~n44682 & ~n44686;
  assign n44688 = i_hlock6 & ~n44687;
  assign n44689 = ~n14631 & ~n27370;
  assign n44690 = controllable_hmaster1 & ~n44689;
  assign n44691 = ~n14668 & ~n44690;
  assign n44692 = n8217 & ~n44691;
  assign n44693 = ~n20175 & ~n29977;
  assign n44694 = controllable_hmaster1 & ~n44693;
  assign n44695 = ~n20219 & ~n44694;
  assign n44696 = ~n8217 & ~n44695;
  assign n44697 = ~n44692 & ~n44696;
  assign n44698 = ~i_hlock6 & ~n44697;
  assign n44699 = ~n44688 & ~n44698;
  assign n44700 = ~i_hbusreq6 & ~n44699;
  assign n44701 = ~n44678 & ~n44700;
  assign n44702 = controllable_hgrant6 & ~n44701;
  assign n44703 = i_hbusreq6 & ~n44111;
  assign n44704 = i_hbusreq5 & ~n44020;
  assign n44705 = n8378 & ~n14626;
  assign n44706 = ~n8378 & ~n20170;
  assign n44707 = ~n44705 & ~n44706;
  assign n44708 = ~i_hbusreq5 & ~n44707;
  assign n44709 = ~n44704 & ~n44708;
  assign n44710 = controllable_hgrant5 & ~n44709;
  assign n44711 = i_hbusreq5 & ~n44048;
  assign n44712 = i_hbusreq4 & ~n44024;
  assign n44713 = i_hbusreq9 & ~n44024;
  assign n44714 = n8426 & ~n14620;
  assign n44715 = ~n8426 & ~n20164;
  assign n44716 = ~n44714 & ~n44715;
  assign n44717 = ~i_hbusreq9 & ~n44716;
  assign n44718 = ~n44713 & ~n44717;
  assign n44719 = ~i_hbusreq4 & ~n44718;
  assign n44720 = ~n44712 & ~n44719;
  assign n44721 = controllable_hgrant4 & ~n44720;
  assign n44722 = i_hbusreq4 & ~n44046;
  assign n44723 = i_hbusreq9 & ~n44046;
  assign n44724 = i_hbusreq3 & ~n44028;
  assign n44725 = n8365 & ~n14616;
  assign n44726 = ~n8365 & ~n20160;
  assign n44727 = ~n44725 & ~n44726;
  assign n44728 = ~i_hbusreq3 & ~n44727;
  assign n44729 = ~n44724 & ~n44728;
  assign n44730 = controllable_hgrant3 & ~n44729;
  assign n44731 = i_hbusreq3 & ~n44044;
  assign n44732 = i_hbusreq1 & ~n44032;
  assign n44733 = n8389 & ~n14612;
  assign n44734 = ~n8389 & ~n20156;
  assign n44735 = ~n44733 & ~n44734;
  assign n44736 = ~i_hbusreq1 & ~n44735;
  assign n44737 = ~n44732 & ~n44736;
  assign n44738 = controllable_hgrant1 & ~n44737;
  assign n44739 = i_hbusreq1 & ~n44042;
  assign n44740 = i_hbusreq2 & ~n44034;
  assign n44741 = i_hbusreq0 & ~n44034;
  assign n44742 = ~n40078 & ~n44182;
  assign n44743 = i_hlock0 & ~n44742;
  assign n44744 = ~i_hlock0 & ~n44034;
  assign n44745 = ~n44743 & ~n44744;
  assign n44746 = ~i_hbusreq0 & ~n44745;
  assign n44747 = ~n44741 & ~n44746;
  assign n44748 = ~i_hbusreq2 & ~n44747;
  assign n44749 = ~n44740 & ~n44748;
  assign n44750 = controllable_hgrant2 & ~n44749;
  assign n44751 = ~n20882 & ~n44750;
  assign n44752 = ~n7733 & ~n44751;
  assign n44753 = ~n18798 & ~n44750;
  assign n44754 = n7733 & ~n44753;
  assign n44755 = ~n44752 & ~n44754;
  assign n44756 = n7928 & ~n44755;
  assign n44757 = ~n43545 & ~n44756;
  assign n44758 = ~i_hbusreq1 & ~n44757;
  assign n44759 = ~n44739 & ~n44758;
  assign n44760 = ~controllable_hgrant1 & ~n44759;
  assign n44761 = ~n44738 & ~n44760;
  assign n44762 = ~i_hbusreq3 & ~n44761;
  assign n44763 = ~n44731 & ~n44762;
  assign n44764 = ~controllable_hgrant3 & ~n44763;
  assign n44765 = ~n44730 & ~n44764;
  assign n44766 = ~i_hbusreq9 & ~n44765;
  assign n44767 = ~n44723 & ~n44766;
  assign n44768 = ~i_hbusreq4 & ~n44767;
  assign n44769 = ~n44722 & ~n44768;
  assign n44770 = ~controllable_hgrant4 & ~n44769;
  assign n44771 = ~n44721 & ~n44770;
  assign n44772 = ~i_hbusreq5 & ~n44771;
  assign n44773 = ~n44711 & ~n44772;
  assign n44774 = ~controllable_hgrant5 & ~n44773;
  assign n44775 = ~n44710 & ~n44774;
  assign n44776 = ~controllable_hmaster2 & ~n44775;
  assign n44777 = ~n44529 & ~n44776;
  assign n44778 = controllable_hmaster1 & ~n44777;
  assign n44779 = i_hbusreq5 & ~n44056;
  assign n44780 = n8378 & ~n14640;
  assign n44781 = ~n8378 & ~n20186;
  assign n44782 = ~n44780 & ~n44781;
  assign n44783 = ~i_hbusreq5 & ~n44782;
  assign n44784 = ~n44779 & ~n44783;
  assign n44785 = controllable_hgrant5 & ~n44784;
  assign n44786 = i_hbusreq5 & ~n44072;
  assign n44787 = i_hbusreq4 & ~n44066;
  assign n44788 = i_hbusreq9 & ~n44060;
  assign n44789 = n8426 & ~n14411;
  assign n44790 = ~n8426 & ~n19910;
  assign n44791 = ~n44789 & ~n44790;
  assign n44792 = ~i_hbusreq9 & ~n44791;
  assign n44793 = ~n44788 & ~n44792;
  assign n44794 = i_hlock4 & ~n44793;
  assign n44795 = i_hbusreq9 & ~n44064;
  assign n44796 = n8426 & ~n14421;
  assign n44797 = ~n8426 & ~n19922;
  assign n44798 = ~n44796 & ~n44797;
  assign n44799 = ~i_hbusreq9 & ~n44798;
  assign n44800 = ~n44795 & ~n44799;
  assign n44801 = ~i_hlock4 & ~n44800;
  assign n44802 = ~n44794 & ~n44801;
  assign n44803 = ~i_hbusreq4 & ~n44802;
  assign n44804 = ~n44787 & ~n44803;
  assign n44805 = controllable_hgrant4 & ~n44804;
  assign n44806 = i_hbusreq4 & ~n44070;
  assign n44807 = i_hlock4 & ~n44422;
  assign n44808 = ~i_hlock4 & ~n44496;
  assign n44809 = ~n44807 & ~n44808;
  assign n44810 = ~i_hbusreq4 & ~n44809;
  assign n44811 = ~n44806 & ~n44810;
  assign n44812 = ~controllable_hgrant4 & ~n44811;
  assign n44813 = ~n44805 & ~n44812;
  assign n44814 = ~i_hbusreq5 & ~n44813;
  assign n44815 = ~n44786 & ~n44814;
  assign n44816 = ~controllable_hgrant5 & ~n44815;
  assign n44817 = ~n44785 & ~n44816;
  assign n44818 = controllable_hmaster2 & ~n44817;
  assign n44819 = i_hbusreq5 & ~n44078;
  assign n44820 = n8378 & ~n14661;
  assign n44821 = ~n8378 & ~n20212;
  assign n44822 = ~n44820 & ~n44821;
  assign n44823 = ~i_hbusreq5 & ~n44822;
  assign n44824 = ~n44819 & ~n44823;
  assign n44825 = controllable_hgrant5 & ~n44824;
  assign n44826 = i_hbusreq5 & ~n44098;
  assign n44827 = i_hbusreq4 & ~n44082;
  assign n44828 = i_hbusreq9 & ~n44082;
  assign n44829 = n8426 & ~n14655;
  assign n44830 = ~n8426 & ~n20206;
  assign n44831 = ~n44829 & ~n44830;
  assign n44832 = ~i_hbusreq9 & ~n44831;
  assign n44833 = ~n44828 & ~n44832;
  assign n44834 = ~i_hbusreq4 & ~n44833;
  assign n44835 = ~n44827 & ~n44834;
  assign n44836 = controllable_hgrant4 & ~n44835;
  assign n44837 = i_hbusreq4 & ~n44096;
  assign n44838 = i_hbusreq9 & ~n44096;
  assign n44839 = i_hbusreq3 & ~n44086;
  assign n44840 = n8365 & ~n14651;
  assign n44841 = ~n8365 & ~n20202;
  assign n44842 = ~n44840 & ~n44841;
  assign n44843 = ~i_hbusreq3 & ~n44842;
  assign n44844 = ~n44839 & ~n44843;
  assign n44845 = controllable_hgrant3 & ~n44844;
  assign n44846 = i_hbusreq3 & ~n44094;
  assign n44847 = i_hbusreq1 & ~n44090;
  assign n44848 = n8389 & ~n14647;
  assign n44849 = ~n8389 & ~n20198;
  assign n44850 = ~n44848 & ~n44849;
  assign n44851 = ~i_hbusreq1 & ~n44850;
  assign n44852 = ~n44847 & ~n44851;
  assign n44853 = controllable_hgrant1 & ~n44852;
  assign n44854 = i_hbusreq1 & ~n44092;
  assign n44855 = controllable_hmastlock & ~n44280;
  assign n44856 = ~n39848 & ~n44855;
  assign n44857 = ~controllable_locked & ~n44856;
  assign n44858 = ~n14240 & ~n44857;
  assign n44859 = i_hlock0 & ~n44858;
  assign n44860 = ~n44185 & ~n44859;
  assign n44861 = ~i_hbusreq0 & ~n44860;
  assign n44862 = ~n44181 & ~n44861;
  assign n44863 = ~i_hbusreq2 & ~n44862;
  assign n44864 = ~n44180 & ~n44863;
  assign n44865 = controllable_hgrant2 & ~n44864;
  assign n44866 = ~n21358 & ~n44865;
  assign n44867 = ~n7733 & ~n44866;
  assign n44868 = ~n19070 & ~n44865;
  assign n44869 = n7733 & ~n44868;
  assign n44870 = ~n44867 & ~n44869;
  assign n44871 = n7928 & ~n44870;
  assign n44872 = ~n8440 & ~n44871;
  assign n44873 = ~i_hbusreq1 & ~n44872;
  assign n44874 = ~n44854 & ~n44873;
  assign n44875 = ~controllable_hgrant1 & ~n44874;
  assign n44876 = ~n44853 & ~n44875;
  assign n44877 = ~i_hbusreq3 & ~n44876;
  assign n44878 = ~n44846 & ~n44877;
  assign n44879 = ~controllable_hgrant3 & ~n44878;
  assign n44880 = ~n44845 & ~n44879;
  assign n44881 = ~i_hbusreq9 & ~n44880;
  assign n44882 = ~n44838 & ~n44881;
  assign n44883 = ~i_hbusreq4 & ~n44882;
  assign n44884 = ~n44837 & ~n44883;
  assign n44885 = ~controllable_hgrant4 & ~n44884;
  assign n44886 = ~n44836 & ~n44885;
  assign n44887 = ~i_hbusreq5 & ~n44886;
  assign n44888 = ~n44826 & ~n44887;
  assign n44889 = ~controllable_hgrant5 & ~n44888;
  assign n44890 = ~n44825 & ~n44889;
  assign n44891 = ~controllable_hmaster2 & ~n44890;
  assign n44892 = ~n44818 & ~n44891;
  assign n44893 = ~controllable_hmaster1 & ~n44892;
  assign n44894 = ~n44778 & ~n44893;
  assign n44895 = i_hlock6 & ~n44894;
  assign n44896 = controllable_hmaster2 & ~n44504;
  assign n44897 = ~n44776 & ~n44896;
  assign n44898 = controllable_hmaster1 & ~n44897;
  assign n44899 = ~n44893 & ~n44898;
  assign n44900 = ~i_hlock6 & ~n44899;
  assign n44901 = ~n44895 & ~n44900;
  assign n44902 = ~i_hbusreq6 & ~n44901;
  assign n44903 = ~n44703 & ~n44902;
  assign n44904 = ~controllable_hgrant6 & ~n44903;
  assign n44905 = ~n44702 & ~n44904;
  assign n44906 = ~controllable_hmaster0 & ~n44905;
  assign n44907 = ~n44677 & ~n44906;
  assign n44908 = ~i_hbusreq8 & ~n44907;
  assign n44909 = ~n44520 & ~n44908;
  assign n44910 = ~controllable_hmaster3 & ~n44909;
  assign n44911 = ~n44519 & ~n44910;
  assign n44912 = i_hlock7 & ~n44911;
  assign n44913 = i_hbusreq8 & ~n44129;
  assign n44914 = i_hbusreq6 & ~n44121;
  assign n44915 = n8217 & ~n14694;
  assign n44916 = ~n8217 & ~n20248;
  assign n44917 = ~n44915 & ~n44916;
  assign n44918 = ~i_hbusreq6 & ~n44917;
  assign n44919 = ~n44914 & ~n44918;
  assign n44920 = controllable_hgrant6 & ~n44919;
  assign n44921 = i_hbusreq6 & ~n44125;
  assign n44922 = ~n44581 & ~n44896;
  assign n44923 = controllable_hmaster1 & ~n44922;
  assign n44924 = ~n44671 & ~n44923;
  assign n44925 = ~i_hbusreq6 & ~n44924;
  assign n44926 = ~n44921 & ~n44925;
  assign n44927 = ~controllable_hgrant6 & ~n44926;
  assign n44928 = ~n44920 & ~n44927;
  assign n44929 = controllable_hmaster0 & ~n44928;
  assign n44930 = ~n44906 & ~n44929;
  assign n44931 = ~i_hbusreq8 & ~n44930;
  assign n44932 = ~n44913 & ~n44931;
  assign n44933 = ~controllable_hmaster3 & ~n44932;
  assign n44934 = ~n44519 & ~n44933;
  assign n44935 = ~i_hlock7 & ~n44934;
  assign n44936 = ~n44912 & ~n44935;
  assign n44937 = ~i_hbusreq7 & ~n44936;
  assign n44938 = ~n44134 & ~n44937;
  assign n44939 = n7924 & ~n44938;
  assign n44940 = ~n43739 & ~n44939;
  assign n44941 = ~n8214 & ~n44940;
  assign n44942 = ~n8217 & ~n30008;
  assign n44943 = ~n41284 & ~n44942;
  assign n44944 = controllable_hgrant6 & ~n44943;
  assign n44945 = ~n8378 & ~n30002;
  assign n44946 = ~n40193 & ~n44945;
  assign n44947 = controllable_hgrant5 & ~n44946;
  assign n44948 = i_hlock9 & ~n42753;
  assign n44949 = ~i_hlock9 & ~n42788;
  assign n44950 = ~n44948 & ~n44949;
  assign n44951 = controllable_hgrant4 & ~n44950;
  assign n44952 = i_hlock9 & ~n42767;
  assign n44953 = ~i_hlock9 & ~n42800;
  assign n44954 = ~n44952 & ~n44953;
  assign n44955 = ~controllable_hgrant4 & ~n44954;
  assign n44956 = ~n44951 & ~n44955;
  assign n44957 = ~controllable_hgrant5 & ~n44956;
  assign n44958 = ~n44947 & ~n44957;
  assign n44959 = ~controllable_hmaster2 & ~n44958;
  assign n44960 = ~n42739 & ~n44959;
  assign n44961 = ~controllable_hmaster1 & ~n44960;
  assign n44962 = ~n42738 & ~n44961;
  assign n44963 = ~controllable_hgrant6 & ~n44962;
  assign n44964 = ~n44944 & ~n44963;
  assign n44965 = controllable_hmaster0 & ~n44964;
  assign n44966 = ~n8217 & ~n19210;
  assign n44967 = ~n42078 & ~n44966;
  assign n44968 = controllable_hgrant6 & ~n44967;
  assign n44969 = ~n40437 & ~n42739;
  assign n44970 = ~controllable_hmaster1 & ~n44969;
  assign n44971 = ~n42738 & ~n44970;
  assign n44972 = ~controllable_hgrant6 & ~n44971;
  assign n44973 = ~n44968 & ~n44972;
  assign n44974 = ~controllable_hmaster0 & ~n44973;
  assign n44975 = ~n44965 & ~n44974;
  assign n44976 = i_hlock8 & ~n44975;
  assign n44977 = ~n8217 & ~n19218;
  assign n44978 = ~n42090 & ~n44977;
  assign n44979 = controllable_hgrant6 & ~n44978;
  assign n44980 = ~n40459 & ~n42739;
  assign n44981 = ~controllable_hmaster1 & ~n44980;
  assign n44982 = ~n42738 & ~n44981;
  assign n44983 = ~controllable_hgrant6 & ~n44982;
  assign n44984 = ~n44979 & ~n44983;
  assign n44985 = ~controllable_hmaster0 & ~n44984;
  assign n44986 = ~n44965 & ~n44985;
  assign n44987 = ~i_hlock8 & ~n44986;
  assign n44988 = ~n44976 & ~n44987;
  assign n44989 = controllable_hmaster3 & ~n44988;
  assign n44990 = ~n43049 & ~n44989;
  assign n44991 = i_hlock7 & ~n44990;
  assign n44992 = ~n43063 & ~n44989;
  assign n44993 = ~i_hlock7 & ~n44992;
  assign n44994 = ~n44991 & ~n44993;
  assign n44995 = i_hbusreq7 & ~n44994;
  assign n44996 = i_hbusreq8 & ~n44988;
  assign n44997 = i_hbusreq6 & ~n44943;
  assign n44998 = n8217 & ~n9476;
  assign n44999 = ~n8217 & ~n30045;
  assign n45000 = ~n44998 & ~n44999;
  assign n45001 = ~i_hbusreq6 & ~n45000;
  assign n45002 = ~n44997 & ~n45001;
  assign n45003 = controllable_hgrant6 & ~n45002;
  assign n45004 = i_hbusreq6 & ~n44962;
  assign n45005 = i_hbusreq5 & ~n44946;
  assign n45006 = n8378 & ~n9470;
  assign n45007 = ~n8378 & ~n30037;
  assign n45008 = ~n45006 & ~n45007;
  assign n45009 = ~i_hbusreq5 & ~n45008;
  assign n45010 = ~n45005 & ~n45009;
  assign n45011 = controllable_hgrant5 & ~n45010;
  assign n45012 = i_hbusreq5 & ~n44956;
  assign n45013 = i_hbusreq4 & ~n44950;
  assign n45014 = i_hbusreq9 & ~n44950;
  assign n45015 = i_hlock9 & ~n43176;
  assign n45016 = ~i_hlock9 & ~n43252;
  assign n45017 = ~n45015 & ~n45016;
  assign n45018 = ~i_hbusreq9 & ~n45017;
  assign n45019 = ~n45014 & ~n45018;
  assign n45020 = ~i_hbusreq4 & ~n45019;
  assign n45021 = ~n45013 & ~n45020;
  assign n45022 = controllable_hgrant4 & ~n45021;
  assign n45023 = i_hbusreq4 & ~n44954;
  assign n45024 = i_hbusreq9 & ~n44954;
  assign n45025 = i_hlock9 & ~n43210;
  assign n45026 = ~i_hlock9 & ~n43284;
  assign n45027 = ~n45025 & ~n45026;
  assign n45028 = ~i_hbusreq9 & ~n45027;
  assign n45029 = ~n45024 & ~n45028;
  assign n45030 = ~i_hbusreq4 & ~n45029;
  assign n45031 = ~n45023 & ~n45030;
  assign n45032 = ~controllable_hgrant4 & ~n45031;
  assign n45033 = ~n45022 & ~n45032;
  assign n45034 = ~i_hbusreq5 & ~n45033;
  assign n45035 = ~n45012 & ~n45034;
  assign n45036 = ~controllable_hgrant5 & ~n45035;
  assign n45037 = ~n45011 & ~n45036;
  assign n45038 = ~controllable_hmaster2 & ~n45037;
  assign n45039 = ~n43147 & ~n45038;
  assign n45040 = ~controllable_hmaster1 & ~n45039;
  assign n45041 = ~n43146 & ~n45040;
  assign n45042 = ~i_hbusreq6 & ~n45041;
  assign n45043 = ~n45004 & ~n45042;
  assign n45044 = ~controllable_hgrant6 & ~n45043;
  assign n45045 = ~n45003 & ~n45044;
  assign n45046 = controllable_hmaster0 & ~n45045;
  assign n45047 = i_hbusreq6 & ~n44967;
  assign n45048 = n8217 & ~n9482;
  assign n45049 = ~n8217 & ~n19419;
  assign n45050 = ~n45048 & ~n45049;
  assign n45051 = ~i_hbusreq6 & ~n45050;
  assign n45052 = ~n45047 & ~n45051;
  assign n45053 = controllable_hgrant6 & ~n45052;
  assign n45054 = i_hbusreq6 & ~n44971;
  assign n45055 = ~n40508 & ~n43147;
  assign n45056 = ~controllable_hmaster1 & ~n45055;
  assign n45057 = ~n43146 & ~n45056;
  assign n45058 = ~i_hbusreq6 & ~n45057;
  assign n45059 = ~n45054 & ~n45058;
  assign n45060 = ~controllable_hgrant6 & ~n45059;
  assign n45061 = ~n45053 & ~n45060;
  assign n45062 = ~controllable_hmaster0 & ~n45061;
  assign n45063 = ~n45046 & ~n45062;
  assign n45064 = i_hlock8 & ~n45063;
  assign n45065 = i_hbusreq6 & ~n44978;
  assign n45066 = n8217 & ~n9490;
  assign n45067 = ~n8217 & ~n19430;
  assign n45068 = ~n45066 & ~n45067;
  assign n45069 = ~i_hbusreq6 & ~n45068;
  assign n45070 = ~n45065 & ~n45069;
  assign n45071 = controllable_hgrant6 & ~n45070;
  assign n45072 = i_hbusreq6 & ~n44982;
  assign n45073 = ~n40554 & ~n43147;
  assign n45074 = ~controllable_hmaster1 & ~n45073;
  assign n45075 = ~n43146 & ~n45074;
  assign n45076 = ~i_hbusreq6 & ~n45075;
  assign n45077 = ~n45072 & ~n45076;
  assign n45078 = ~controllable_hgrant6 & ~n45077;
  assign n45079 = ~n45071 & ~n45078;
  assign n45080 = ~controllable_hmaster0 & ~n45079;
  assign n45081 = ~n45046 & ~n45080;
  assign n45082 = ~i_hlock8 & ~n45081;
  assign n45083 = ~n45064 & ~n45082;
  assign n45084 = ~i_hbusreq8 & ~n45083;
  assign n45085 = ~n44996 & ~n45084;
  assign n45086 = controllable_hmaster3 & ~n45085;
  assign n45087 = ~n43710 & ~n45086;
  assign n45088 = i_hlock7 & ~n45087;
  assign n45089 = ~n43733 & ~n45086;
  assign n45090 = ~i_hlock7 & ~n45089;
  assign n45091 = ~n45088 & ~n45090;
  assign n45092 = ~i_hbusreq7 & ~n45091;
  assign n45093 = ~n44995 & ~n45092;
  assign n45094 = ~n7924 & ~n45093;
  assign n45095 = ~n8217 & ~n30077;
  assign n45096 = ~n41555 & ~n45095;
  assign n45097 = controllable_hgrant6 & ~n45096;
  assign n45098 = ~n8378 & ~n30071;
  assign n45099 = ~n41580 & ~n45098;
  assign n45100 = controllable_hgrant5 & ~n45099;
  assign n45101 = i_hlock9 & ~n43838;
  assign n45102 = ~i_hlock9 & ~n43877;
  assign n45103 = ~n45101 & ~n45102;
  assign n45104 = controllable_hgrant4 & ~n45103;
  assign n45105 = i_hlock9 & ~n43856;
  assign n45106 = ~i_hlock9 & ~n43889;
  assign n45107 = ~n45105 & ~n45106;
  assign n45108 = ~controllable_hgrant4 & ~n45107;
  assign n45109 = ~n45104 & ~n45108;
  assign n45110 = ~controllable_hgrant5 & ~n45109;
  assign n45111 = ~n45100 & ~n45110;
  assign n45112 = ~controllable_hmaster2 & ~n45111;
  assign n45113 = ~n43777 & ~n45112;
  assign n45114 = ~controllable_hmaster1 & ~n45113;
  assign n45115 = ~n43776 & ~n45114;
  assign n45116 = ~controllable_hgrant6 & ~n45115;
  assign n45117 = ~n45097 & ~n45116;
  assign n45118 = controllable_hmaster0 & ~n45117;
  assign n45119 = ~n8217 & ~n19726;
  assign n45120 = ~n42153 & ~n45119;
  assign n45121 = controllable_hgrant6 & ~n45120;
  assign n45122 = ~n8378 & ~n19720;
  assign n45123 = ~n42157 & ~n45122;
  assign n45124 = controllable_hgrant5 & ~n45123;
  assign n45125 = controllable_hgrant4 & ~n43782;
  assign n45126 = ~controllable_hgrant4 & ~n43805;
  assign n45127 = ~n45125 & ~n45126;
  assign n45128 = ~controllable_hgrant5 & ~n45127;
  assign n45129 = ~n45124 & ~n45128;
  assign n45130 = ~controllable_hmaster2 & ~n45129;
  assign n45131 = ~n43777 & ~n45130;
  assign n45132 = ~controllable_hmaster1 & ~n45131;
  assign n45133 = ~n43776 & ~n45132;
  assign n45134 = ~controllable_hgrant6 & ~n45133;
  assign n45135 = ~n45121 & ~n45134;
  assign n45136 = ~controllable_hmaster0 & ~n45135;
  assign n45137 = ~n45118 & ~n45136;
  assign n45138 = i_hlock8 & ~n45137;
  assign n45139 = ~n8217 & ~n19744;
  assign n45140 = ~n42175 & ~n45139;
  assign n45141 = controllable_hgrant6 & ~n45140;
  assign n45142 = ~n8378 & ~n19738;
  assign n45143 = ~n42179 & ~n45142;
  assign n45144 = controllable_hgrant5 & ~n45143;
  assign n45145 = controllable_hgrant4 & ~n43785;
  assign n45146 = ~controllable_hgrant4 & ~n43817;
  assign n45147 = ~n45145 & ~n45146;
  assign n45148 = ~controllable_hgrant5 & ~n45147;
  assign n45149 = ~n45144 & ~n45148;
  assign n45150 = ~controllable_hmaster2 & ~n45149;
  assign n45151 = ~n43777 & ~n45150;
  assign n45152 = ~controllable_hmaster1 & ~n45151;
  assign n45153 = ~n43776 & ~n45152;
  assign n45154 = ~controllable_hgrant6 & ~n45153;
  assign n45155 = ~n45141 & ~n45154;
  assign n45156 = ~controllable_hmaster0 & ~n45155;
  assign n45157 = ~n45118 & ~n45156;
  assign n45158 = ~i_hlock8 & ~n45157;
  assign n45159 = ~n45138 & ~n45158;
  assign n45160 = controllable_hmaster3 & ~n45159;
  assign n45161 = ~n44116 & ~n45160;
  assign n45162 = i_hlock7 & ~n45161;
  assign n45163 = ~n44130 & ~n45160;
  assign n45164 = ~i_hlock7 & ~n45163;
  assign n45165 = ~n45162 & ~n45164;
  assign n45166 = i_hbusreq7 & ~n45165;
  assign n45167 = i_hbusreq8 & ~n45159;
  assign n45168 = i_hbusreq6 & ~n45096;
  assign n45169 = n8217 & ~n27415;
  assign n45170 = ~n8217 & ~n30114;
  assign n45171 = ~n45169 & ~n45170;
  assign n45172 = ~i_hbusreq6 & ~n45171;
  assign n45173 = ~n45168 & ~n45172;
  assign n45174 = controllable_hgrant6 & ~n45173;
  assign n45175 = i_hbusreq6 & ~n45115;
  assign n45176 = i_hbusreq5 & ~n45099;
  assign n45177 = n8378 & ~n27407;
  assign n45178 = ~n8378 & ~n30106;
  assign n45179 = ~n45177 & ~n45178;
  assign n45180 = ~i_hbusreq5 & ~n45179;
  assign n45181 = ~n45176 & ~n45180;
  assign n45182 = controllable_hgrant5 & ~n45181;
  assign n45183 = i_hbusreq5 & ~n45109;
  assign n45184 = i_hbusreq4 & ~n45103;
  assign n45185 = i_hbusreq9 & ~n45103;
  assign n45186 = i_hlock9 & ~n44382;
  assign n45187 = ~i_hlock9 & ~n44462;
  assign n45188 = ~n45186 & ~n45187;
  assign n45189 = ~i_hbusreq9 & ~n45188;
  assign n45190 = ~n45185 & ~n45189;
  assign n45191 = ~i_hbusreq4 & ~n45190;
  assign n45192 = ~n45184 & ~n45191;
  assign n45193 = controllable_hgrant4 & ~n45192;
  assign n45194 = i_hbusreq4 & ~n45107;
  assign n45195 = i_hbusreq9 & ~n45107;
  assign n45196 = i_hlock9 & ~n44420;
  assign n45197 = ~i_hlock9 & ~n44494;
  assign n45198 = ~n45196 & ~n45197;
  assign n45199 = ~i_hbusreq9 & ~n45198;
  assign n45200 = ~n45195 & ~n45199;
  assign n45201 = ~i_hbusreq4 & ~n45200;
  assign n45202 = ~n45194 & ~n45201;
  assign n45203 = ~controllable_hgrant4 & ~n45202;
  assign n45204 = ~n45193 & ~n45203;
  assign n45205 = ~i_hbusreq5 & ~n45204;
  assign n45206 = ~n45183 & ~n45205;
  assign n45207 = ~controllable_hgrant5 & ~n45206;
  assign n45208 = ~n45182 & ~n45207;
  assign n45209 = ~controllable_hmaster2 & ~n45208;
  assign n45210 = ~n44224 & ~n45209;
  assign n45211 = ~controllable_hmaster1 & ~n45210;
  assign n45212 = ~n44223 & ~n45211;
  assign n45213 = ~i_hbusreq6 & ~n45212;
  assign n45214 = ~n45175 & ~n45213;
  assign n45215 = ~controllable_hgrant6 & ~n45214;
  assign n45216 = ~n45174 & ~n45215;
  assign n45217 = controllable_hmaster0 & ~n45216;
  assign n45218 = i_hbusreq6 & ~n45120;
  assign n45219 = n8217 & ~n14476;
  assign n45220 = ~n8217 & ~n19988;
  assign n45221 = ~n45219 & ~n45220;
  assign n45222 = ~i_hbusreq6 & ~n45221;
  assign n45223 = ~n45218 & ~n45222;
  assign n45224 = controllable_hgrant6 & ~n45223;
  assign n45225 = i_hbusreq6 & ~n45133;
  assign n45226 = i_hbusreq5 & ~n45123;
  assign n45227 = n8378 & ~n14468;
  assign n45228 = ~n8378 & ~n19980;
  assign n45229 = ~n45227 & ~n45228;
  assign n45230 = ~i_hbusreq5 & ~n45229;
  assign n45231 = ~n45226 & ~n45230;
  assign n45232 = controllable_hgrant5 & ~n45231;
  assign n45233 = i_hbusreq5 & ~n45127;
  assign n45234 = i_hbusreq4 & ~n43782;
  assign n45235 = i_hbusreq9 & ~n43782;
  assign n45236 = ~i_hbusreq9 & ~n44237;
  assign n45237 = ~n45235 & ~n45236;
  assign n45238 = ~i_hbusreq4 & ~n45237;
  assign n45239 = ~n45234 & ~n45238;
  assign n45240 = controllable_hgrant4 & ~n45239;
  assign n45241 = i_hbusreq4 & ~n43805;
  assign n45242 = i_hbusreq9 & ~n43805;
  assign n45243 = ~i_hbusreq9 & ~n44314;
  assign n45244 = ~n45242 & ~n45243;
  assign n45245 = ~i_hbusreq4 & ~n45244;
  assign n45246 = ~n45241 & ~n45245;
  assign n45247 = ~controllable_hgrant4 & ~n45246;
  assign n45248 = ~n45240 & ~n45247;
  assign n45249 = ~i_hbusreq5 & ~n45248;
  assign n45250 = ~n45233 & ~n45249;
  assign n45251 = ~controllable_hgrant5 & ~n45250;
  assign n45252 = ~n45232 & ~n45251;
  assign n45253 = ~controllable_hmaster2 & ~n45252;
  assign n45254 = ~n44224 & ~n45253;
  assign n45255 = ~controllable_hmaster1 & ~n45254;
  assign n45256 = ~n44223 & ~n45255;
  assign n45257 = ~i_hbusreq6 & ~n45256;
  assign n45258 = ~n45225 & ~n45257;
  assign n45259 = ~controllable_hgrant6 & ~n45258;
  assign n45260 = ~n45224 & ~n45259;
  assign n45261 = ~controllable_hmaster0 & ~n45260;
  assign n45262 = ~n45217 & ~n45261;
  assign n45263 = i_hlock8 & ~n45262;
  assign n45264 = i_hbusreq6 & ~n45140;
  assign n45265 = n8217 & ~n14507;
  assign n45266 = ~n8217 & ~n20024;
  assign n45267 = ~n45265 & ~n45266;
  assign n45268 = ~i_hbusreq6 & ~n45267;
  assign n45269 = ~n45264 & ~n45268;
  assign n45270 = controllable_hgrant6 & ~n45269;
  assign n45271 = i_hbusreq6 & ~n45153;
  assign n45272 = i_hbusreq5 & ~n45143;
  assign n45273 = n8378 & ~n14499;
  assign n45274 = ~n8378 & ~n20016;
  assign n45275 = ~n45273 & ~n45274;
  assign n45276 = ~i_hbusreq5 & ~n45275;
  assign n45277 = ~n45272 & ~n45276;
  assign n45278 = controllable_hgrant5 & ~n45277;
  assign n45279 = i_hbusreq5 & ~n45147;
  assign n45280 = i_hbusreq4 & ~n43785;
  assign n45281 = i_hbusreq9 & ~n43785;
  assign n45282 = ~i_hbusreq9 & ~n44241;
  assign n45283 = ~n45281 & ~n45282;
  assign n45284 = ~i_hbusreq4 & ~n45283;
  assign n45285 = ~n45280 & ~n45284;
  assign n45286 = controllable_hgrant4 & ~n45285;
  assign n45287 = i_hbusreq4 & ~n43817;
  assign n45288 = i_hbusreq9 & ~n43817;
  assign n45289 = ~i_hbusreq9 & ~n44340;
  assign n45290 = ~n45288 & ~n45289;
  assign n45291 = ~i_hbusreq4 & ~n45290;
  assign n45292 = ~n45287 & ~n45291;
  assign n45293 = ~controllable_hgrant4 & ~n45292;
  assign n45294 = ~n45286 & ~n45293;
  assign n45295 = ~i_hbusreq5 & ~n45294;
  assign n45296 = ~n45279 & ~n45295;
  assign n45297 = ~controllable_hgrant5 & ~n45296;
  assign n45298 = ~n45278 & ~n45297;
  assign n45299 = ~controllable_hmaster2 & ~n45298;
  assign n45300 = ~n44224 & ~n45299;
  assign n45301 = ~controllable_hmaster1 & ~n45300;
  assign n45302 = ~n44223 & ~n45301;
  assign n45303 = ~i_hbusreq6 & ~n45302;
  assign n45304 = ~n45271 & ~n45303;
  assign n45305 = ~controllable_hgrant6 & ~n45304;
  assign n45306 = ~n45270 & ~n45305;
  assign n45307 = ~controllable_hmaster0 & ~n45306;
  assign n45308 = ~n45217 & ~n45307;
  assign n45309 = ~i_hlock8 & ~n45308;
  assign n45310 = ~n45263 & ~n45309;
  assign n45311 = ~i_hbusreq8 & ~n45310;
  assign n45312 = ~n45167 & ~n45311;
  assign n45313 = controllable_hmaster3 & ~n45312;
  assign n45314 = ~n44910 & ~n45313;
  assign n45315 = i_hlock7 & ~n45314;
  assign n45316 = ~n44933 & ~n45313;
  assign n45317 = ~i_hlock7 & ~n45316;
  assign n45318 = ~n45315 & ~n45317;
  assign n45319 = ~i_hbusreq7 & ~n45318;
  assign n45320 = ~n45166 & ~n45319;
  assign n45321 = n7924 & ~n45320;
  assign n45322 = ~n45094 & ~n45321;
  assign n45323 = n8214 & ~n45322;
  assign n45324 = ~n44941 & ~n45323;
  assign n45325 = ~n8202 & ~n45324;
  assign n45326 = ~n42778 & ~n44965;
  assign n45327 = i_hlock8 & ~n45326;
  assign n45328 = ~n42811 & ~n44965;
  assign n45329 = ~i_hlock8 & ~n45328;
  assign n45330 = ~n45327 & ~n45329;
  assign n45331 = controllable_hmaster3 & ~n45330;
  assign n45332 = ~n8217 & ~n20290;
  assign n45333 = ~n42816 & ~n45332;
  assign n45334 = controllable_hgrant6 & ~n45333;
  assign n45335 = ~n40579 & ~n42848;
  assign n45336 = controllable_hmaster1 & ~n45335;
  assign n45337 = ~n42902 & ~n45336;
  assign n45338 = ~controllable_hgrant6 & ~n45337;
  assign n45339 = ~n45334 & ~n45338;
  assign n45340 = controllable_hmaster0 & ~n45339;
  assign n45341 = ~n43047 & ~n45340;
  assign n45342 = ~controllable_hmaster3 & ~n45341;
  assign n45343 = ~n45331 & ~n45342;
  assign n45344 = i_hlock7 & ~n45343;
  assign n45345 = ~n8217 & ~n20300;
  assign n45346 = ~n43052 & ~n45345;
  assign n45347 = controllable_hgrant6 & ~n45346;
  assign n45348 = ~n40594 & ~n42848;
  assign n45349 = controllable_hmaster1 & ~n45348;
  assign n45350 = ~n42902 & ~n45349;
  assign n45351 = ~controllable_hgrant6 & ~n45350;
  assign n45352 = ~n45347 & ~n45351;
  assign n45353 = controllable_hmaster0 & ~n45352;
  assign n45354 = ~n43047 & ~n45353;
  assign n45355 = ~controllable_hmaster3 & ~n45354;
  assign n45356 = ~n45331 & ~n45355;
  assign n45357 = ~i_hlock7 & ~n45356;
  assign n45358 = ~n45344 & ~n45357;
  assign n45359 = i_hbusreq7 & ~n45358;
  assign n45360 = i_hbusreq8 & ~n45330;
  assign n45361 = ~n43229 & ~n45046;
  assign n45362 = i_hlock8 & ~n45361;
  assign n45363 = ~n43303 & ~n45046;
  assign n45364 = ~i_hlock8 & ~n45363;
  assign n45365 = ~n45362 & ~n45364;
  assign n45366 = ~i_hbusreq8 & ~n45365;
  assign n45367 = ~n45360 & ~n45366;
  assign n45368 = controllable_hmaster3 & ~n45367;
  assign n45369 = i_hbusreq8 & ~n45341;
  assign n45370 = i_hbusreq6 & ~n45333;
  assign n45371 = n8217 & ~n9520;
  assign n45372 = ~n8217 & ~n20343;
  assign n45373 = ~n45371 & ~n45372;
  assign n45374 = ~i_hbusreq6 & ~n45373;
  assign n45375 = ~n45370 & ~n45374;
  assign n45376 = controllable_hgrant6 & ~n45375;
  assign n45377 = i_hbusreq6 & ~n45337;
  assign n45378 = ~n40616 & ~n43371;
  assign n45379 = controllable_hmaster1 & ~n45378;
  assign n45380 = ~n43461 & ~n45379;
  assign n45381 = ~i_hbusreq6 & ~n45380;
  assign n45382 = ~n45377 & ~n45381;
  assign n45383 = ~controllable_hgrant6 & ~n45382;
  assign n45384 = ~n45376 & ~n45383;
  assign n45385 = controllable_hmaster0 & ~n45384;
  assign n45386 = ~n43706 & ~n45385;
  assign n45387 = ~i_hbusreq8 & ~n45386;
  assign n45388 = ~n45369 & ~n45387;
  assign n45389 = ~controllable_hmaster3 & ~n45388;
  assign n45390 = ~n45368 & ~n45389;
  assign n45391 = i_hlock7 & ~n45390;
  assign n45392 = i_hbusreq8 & ~n45354;
  assign n45393 = i_hbusreq6 & ~n45346;
  assign n45394 = n8217 & ~n9532;
  assign n45395 = ~n8217 & ~n20359;
  assign n45396 = ~n45394 & ~n45395;
  assign n45397 = ~i_hbusreq6 & ~n45396;
  assign n45398 = ~n45393 & ~n45397;
  assign n45399 = controllable_hgrant6 & ~n45398;
  assign n45400 = i_hbusreq6 & ~n45350;
  assign n45401 = ~n40640 & ~n43371;
  assign n45402 = controllable_hmaster1 & ~n45401;
  assign n45403 = ~n43461 & ~n45402;
  assign n45404 = ~i_hbusreq6 & ~n45403;
  assign n45405 = ~n45400 & ~n45404;
  assign n45406 = ~controllable_hgrant6 & ~n45405;
  assign n45407 = ~n45399 & ~n45406;
  assign n45408 = controllable_hmaster0 & ~n45407;
  assign n45409 = ~n43706 & ~n45408;
  assign n45410 = ~i_hbusreq8 & ~n45409;
  assign n45411 = ~n45392 & ~n45410;
  assign n45412 = ~controllable_hmaster3 & ~n45411;
  assign n45413 = ~n45368 & ~n45412;
  assign n45414 = ~i_hlock7 & ~n45413;
  assign n45415 = ~n45391 & ~n45414;
  assign n45416 = ~i_hbusreq7 & ~n45415;
  assign n45417 = ~n45359 & ~n45416;
  assign n45418 = ~n7924 & ~n45417;
  assign n45419 = ~n43867 & ~n45118;
  assign n45420 = i_hlock8 & ~n45419;
  assign n45421 = ~n43900 & ~n45118;
  assign n45422 = ~i_hlock8 & ~n45421;
  assign n45423 = ~n45420 & ~n45422;
  assign n45424 = controllable_hmaster3 & ~n45423;
  assign n45425 = ~n8217 & ~n20398;
  assign n45426 = ~n43905 & ~n45425;
  assign n45427 = controllable_hgrant6 & ~n45426;
  assign n45428 = controllable_hmaster2 & ~n45129;
  assign n45429 = ~n43937 & ~n45428;
  assign n45430 = controllable_hmaster1 & ~n45429;
  assign n45431 = ~n43991 & ~n45430;
  assign n45432 = ~controllable_hgrant6 & ~n45431;
  assign n45433 = ~n45427 & ~n45432;
  assign n45434 = controllable_hmaster0 & ~n45433;
  assign n45435 = ~n44114 & ~n45434;
  assign n45436 = ~controllable_hmaster3 & ~n45435;
  assign n45437 = ~n45424 & ~n45436;
  assign n45438 = i_hlock7 & ~n45437;
  assign n45439 = ~n8217 & ~n20409;
  assign n45440 = ~n44119 & ~n45439;
  assign n45441 = controllable_hgrant6 & ~n45440;
  assign n45442 = controllable_hmaster2 & ~n45149;
  assign n45443 = ~n43937 & ~n45442;
  assign n45444 = controllable_hmaster1 & ~n45443;
  assign n45445 = ~n43991 & ~n45444;
  assign n45446 = ~controllable_hgrant6 & ~n45445;
  assign n45447 = ~n45441 & ~n45446;
  assign n45448 = controllable_hmaster0 & ~n45447;
  assign n45449 = ~n44114 & ~n45448;
  assign n45450 = ~controllable_hmaster3 & ~n45449;
  assign n45451 = ~n45424 & ~n45450;
  assign n45452 = ~i_hlock7 & ~n45451;
  assign n45453 = ~n45438 & ~n45452;
  assign n45454 = i_hbusreq7 & ~n45453;
  assign n45455 = i_hbusreq8 & ~n45423;
  assign n45456 = ~n44439 & ~n45217;
  assign n45457 = i_hlock8 & ~n45456;
  assign n45458 = ~n44513 & ~n45217;
  assign n45459 = ~i_hlock8 & ~n45458;
  assign n45460 = ~n45457 & ~n45459;
  assign n45461 = ~i_hbusreq8 & ~n45460;
  assign n45462 = ~n45455 & ~n45461;
  assign n45463 = controllable_hmaster3 & ~n45462;
  assign n45464 = i_hbusreq8 & ~n45435;
  assign n45465 = i_hbusreq6 & ~n45426;
  assign n45466 = n8217 & ~n14760;
  assign n45467 = ~n8217 & ~n20453;
  assign n45468 = ~n45466 & ~n45467;
  assign n45469 = ~i_hbusreq6 & ~n45468;
  assign n45470 = ~n45465 & ~n45469;
  assign n45471 = controllable_hgrant6 & ~n45470;
  assign n45472 = i_hbusreq6 & ~n45431;
  assign n45473 = controllable_hmaster2 & ~n45252;
  assign n45474 = ~n44581 & ~n45473;
  assign n45475 = controllable_hmaster1 & ~n45474;
  assign n45476 = ~n44671 & ~n45475;
  assign n45477 = ~i_hbusreq6 & ~n45476;
  assign n45478 = ~n45472 & ~n45477;
  assign n45479 = ~controllable_hgrant6 & ~n45478;
  assign n45480 = ~n45471 & ~n45479;
  assign n45481 = controllable_hmaster0 & ~n45480;
  assign n45482 = ~n44906 & ~n45481;
  assign n45483 = ~i_hbusreq8 & ~n45482;
  assign n45484 = ~n45464 & ~n45483;
  assign n45485 = ~controllable_hmaster3 & ~n45484;
  assign n45486 = ~n45463 & ~n45485;
  assign n45487 = i_hlock7 & ~n45486;
  assign n45488 = i_hbusreq8 & ~n45449;
  assign n45489 = i_hbusreq6 & ~n45440;
  assign n45490 = n8217 & ~n14776;
  assign n45491 = ~n8217 & ~n20470;
  assign n45492 = ~n45490 & ~n45491;
  assign n45493 = ~i_hbusreq6 & ~n45492;
  assign n45494 = ~n45489 & ~n45493;
  assign n45495 = controllable_hgrant6 & ~n45494;
  assign n45496 = i_hbusreq6 & ~n45445;
  assign n45497 = controllable_hmaster2 & ~n45298;
  assign n45498 = ~n44581 & ~n45497;
  assign n45499 = controllable_hmaster1 & ~n45498;
  assign n45500 = ~n44671 & ~n45499;
  assign n45501 = ~i_hbusreq6 & ~n45500;
  assign n45502 = ~n45496 & ~n45501;
  assign n45503 = ~controllable_hgrant6 & ~n45502;
  assign n45504 = ~n45495 & ~n45503;
  assign n45505 = controllable_hmaster0 & ~n45504;
  assign n45506 = ~n44906 & ~n45505;
  assign n45507 = ~i_hbusreq8 & ~n45506;
  assign n45508 = ~n45488 & ~n45507;
  assign n45509 = ~controllable_hmaster3 & ~n45508;
  assign n45510 = ~n45463 & ~n45509;
  assign n45511 = ~i_hlock7 & ~n45510;
  assign n45512 = ~n45487 & ~n45511;
  assign n45513 = ~i_hbusreq7 & ~n45512;
  assign n45514 = ~n45454 & ~n45513;
  assign n45515 = n7924 & ~n45514;
  assign n45516 = ~n45418 & ~n45515;
  assign n45517 = ~n8214 & ~n45516;
  assign n45518 = ~n8217 & ~n30142;
  assign n45519 = ~n41284 & ~n45518;
  assign n45520 = controllable_hgrant6 & ~n45519;
  assign n45521 = ~n44963 & ~n45520;
  assign n45522 = controllable_hmaster0 & ~n45521;
  assign n45523 = ~n8217 & ~n18098;
  assign n45524 = ~n42078 & ~n45523;
  assign n45525 = controllable_hgrant6 & ~n45524;
  assign n45526 = ~n42776 & ~n45525;
  assign n45527 = ~controllable_hmaster0 & ~n45526;
  assign n45528 = ~n45522 & ~n45527;
  assign n45529 = i_hlock8 & ~n45528;
  assign n45530 = ~n8217 & ~n18106;
  assign n45531 = ~n42090 & ~n45530;
  assign n45532 = controllable_hgrant6 & ~n45531;
  assign n45533 = ~n42809 & ~n45532;
  assign n45534 = ~controllable_hmaster0 & ~n45533;
  assign n45535 = ~n45522 & ~n45534;
  assign n45536 = ~i_hlock8 & ~n45535;
  assign n45537 = ~n45529 & ~n45536;
  assign n45538 = controllable_hmaster3 & ~n45537;
  assign n45539 = ~n8217 & ~n18146;
  assign n45540 = ~n42816 & ~n45539;
  assign n45541 = controllable_hgrant6 & ~n45540;
  assign n45542 = ~n42904 & ~n45541;
  assign n45543 = controllable_hmaster0 & ~n45542;
  assign n45544 = ~n18159 & ~n28870;
  assign n45545 = controllable_hmaster1 & ~n45544;
  assign n45546 = ~n18181 & ~n45545;
  assign n45547 = ~n8217 & ~n45546;
  assign n45548 = ~n42910 & ~n45547;
  assign n45549 = i_hlock6 & ~n45548;
  assign n45550 = ~n18159 & ~n28885;
  assign n45551 = controllable_hmaster1 & ~n45550;
  assign n45552 = ~n18181 & ~n45551;
  assign n45553 = ~n8217 & ~n45552;
  assign n45554 = ~n42920 & ~n45553;
  assign n45555 = ~i_hlock6 & ~n45554;
  assign n45556 = ~n45549 & ~n45555;
  assign n45557 = controllable_hgrant6 & ~n45556;
  assign n45558 = ~n40579 & ~n42984;
  assign n45559 = controllable_hmaster1 & ~n45558;
  assign n45560 = ~n43036 & ~n45559;
  assign n45561 = i_hlock6 & ~n45560;
  assign n45562 = ~n40594 & ~n42984;
  assign n45563 = controllable_hmaster1 & ~n45562;
  assign n45564 = ~n43036 & ~n45563;
  assign n45565 = ~i_hlock6 & ~n45564;
  assign n45566 = ~n45561 & ~n45565;
  assign n45567 = ~controllable_hgrant6 & ~n45566;
  assign n45568 = ~n45557 & ~n45567;
  assign n45569 = ~controllable_hmaster0 & ~n45568;
  assign n45570 = ~n45543 & ~n45569;
  assign n45571 = ~controllable_hmaster3 & ~n45570;
  assign n45572 = ~n45538 & ~n45571;
  assign n45573 = i_hlock7 & ~n45572;
  assign n45574 = ~n8217 & ~n18198;
  assign n45575 = ~n43052 & ~n45574;
  assign n45576 = controllable_hgrant6 & ~n45575;
  assign n45577 = ~n43059 & ~n45576;
  assign n45578 = controllable_hmaster0 & ~n45577;
  assign n45579 = ~n45569 & ~n45578;
  assign n45580 = ~controllable_hmaster3 & ~n45579;
  assign n45581 = ~n45538 & ~n45580;
  assign n45582 = ~i_hlock7 & ~n45581;
  assign n45583 = ~n45573 & ~n45582;
  assign n45584 = i_hbusreq7 & ~n45583;
  assign n45585 = i_hbusreq8 & ~n45537;
  assign n45586 = i_hbusreq6 & ~n45519;
  assign n45587 = ~n8217 & ~n30192;
  assign n45588 = ~n44998 & ~n45587;
  assign n45589 = ~i_hbusreq6 & ~n45588;
  assign n45590 = ~n45586 & ~n45589;
  assign n45591 = controllable_hgrant6 & ~n45590;
  assign n45592 = ~n45044 & ~n45591;
  assign n45593 = controllable_hmaster0 & ~n45592;
  assign n45594 = i_hbusreq6 & ~n45524;
  assign n45595 = ~n8217 & ~n18282;
  assign n45596 = ~n43157 & ~n45595;
  assign n45597 = ~i_hbusreq6 & ~n45596;
  assign n45598 = ~n45594 & ~n45597;
  assign n45599 = controllable_hgrant6 & ~n45598;
  assign n45600 = ~n43227 & ~n45599;
  assign n45601 = ~controllable_hmaster0 & ~n45600;
  assign n45602 = ~n45593 & ~n45601;
  assign n45603 = i_hlock8 & ~n45602;
  assign n45604 = i_hbusreq6 & ~n45531;
  assign n45605 = ~n8217 & ~n18313;
  assign n45606 = ~n43233 & ~n45605;
  assign n45607 = ~i_hbusreq6 & ~n45606;
  assign n45608 = ~n45604 & ~n45607;
  assign n45609 = controllable_hgrant6 & ~n45608;
  assign n45610 = ~n43301 & ~n45609;
  assign n45611 = ~controllable_hmaster0 & ~n45610;
  assign n45612 = ~n45593 & ~n45611;
  assign n45613 = ~i_hlock8 & ~n45612;
  assign n45614 = ~n45603 & ~n45613;
  assign n45615 = ~i_hbusreq8 & ~n45614;
  assign n45616 = ~n45585 & ~n45615;
  assign n45617 = controllable_hmaster3 & ~n45616;
  assign n45618 = i_hbusreq8 & ~n45570;
  assign n45619 = i_hbusreq6 & ~n45540;
  assign n45620 = ~n8217 & ~n18390;
  assign n45621 = ~n43312 & ~n45620;
  assign n45622 = ~i_hbusreq6 & ~n45621;
  assign n45623 = ~n45619 & ~n45622;
  assign n45624 = controllable_hgrant6 & ~n45623;
  assign n45625 = ~n43465 & ~n45624;
  assign n45626 = controllable_hmaster0 & ~n45625;
  assign n45627 = i_hbusreq6 & ~n45556;
  assign n45628 = ~n9391 & ~n26684;
  assign n45629 = controllable_hmaster1 & ~n45628;
  assign n45630 = ~n9428 & ~n45629;
  assign n45631 = n8217 & ~n45630;
  assign n45632 = ~n18421 & ~n28913;
  assign n45633 = controllable_hmaster1 & ~n45632;
  assign n45634 = ~n18490 & ~n45633;
  assign n45635 = ~n8217 & ~n45634;
  assign n45636 = ~n45631 & ~n45635;
  assign n45637 = i_hlock6 & ~n45636;
  assign n45638 = ~n9391 & ~n26714;
  assign n45639 = controllable_hmaster1 & ~n45638;
  assign n45640 = ~n9428 & ~n45639;
  assign n45641 = n8217 & ~n45640;
  assign n45642 = ~n18421 & ~n28943;
  assign n45643 = controllable_hmaster1 & ~n45642;
  assign n45644 = ~n18490 & ~n45643;
  assign n45645 = ~n8217 & ~n45644;
  assign n45646 = ~n45641 & ~n45645;
  assign n45647 = ~i_hlock6 & ~n45646;
  assign n45648 = ~n45637 & ~n45647;
  assign n45649 = ~i_hbusreq6 & ~n45648;
  assign n45650 = ~n45627 & ~n45649;
  assign n45651 = controllable_hgrant6 & ~n45650;
  assign n45652 = i_hbusreq6 & ~n45566;
  assign n45653 = ~n40616 & ~n43580;
  assign n45654 = controllable_hmaster1 & ~n45653;
  assign n45655 = ~n43693 & ~n45654;
  assign n45656 = i_hlock6 & ~n45655;
  assign n45657 = ~n40640 & ~n43580;
  assign n45658 = controllable_hmaster1 & ~n45657;
  assign n45659 = ~n43693 & ~n45658;
  assign n45660 = ~i_hlock6 & ~n45659;
  assign n45661 = ~n45656 & ~n45660;
  assign n45662 = ~i_hbusreq6 & ~n45661;
  assign n45663 = ~n45652 & ~n45662;
  assign n45664 = ~controllable_hgrant6 & ~n45663;
  assign n45665 = ~n45651 & ~n45664;
  assign n45666 = ~controllable_hmaster0 & ~n45665;
  assign n45667 = ~n45626 & ~n45666;
  assign n45668 = ~i_hbusreq8 & ~n45667;
  assign n45669 = ~n45618 & ~n45668;
  assign n45670 = ~controllable_hmaster3 & ~n45669;
  assign n45671 = ~n45617 & ~n45670;
  assign n45672 = i_hlock7 & ~n45671;
  assign n45673 = i_hbusreq8 & ~n45579;
  assign n45674 = i_hbusreq6 & ~n45575;
  assign n45675 = ~n8217 & ~n18514;
  assign n45676 = ~n43715 & ~n45675;
  assign n45677 = ~i_hbusreq6 & ~n45676;
  assign n45678 = ~n45674 & ~n45677;
  assign n45679 = controllable_hgrant6 & ~n45678;
  assign n45680 = ~n43727 & ~n45679;
  assign n45681 = controllable_hmaster0 & ~n45680;
  assign n45682 = ~n45666 & ~n45681;
  assign n45683 = ~i_hbusreq8 & ~n45682;
  assign n45684 = ~n45673 & ~n45683;
  assign n45685 = ~controllable_hmaster3 & ~n45684;
  assign n45686 = ~n45617 & ~n45685;
  assign n45687 = ~i_hlock7 & ~n45686;
  assign n45688 = ~n45672 & ~n45687;
  assign n45689 = ~i_hbusreq7 & ~n45688;
  assign n45690 = ~n45584 & ~n45689;
  assign n45691 = ~n7924 & ~n45690;
  assign n45692 = ~n8217 & ~n30251;
  assign n45693 = ~n41555 & ~n45692;
  assign n45694 = i_hlock6 & ~n45693;
  assign n45695 = ~n8217 & ~n30354;
  assign n45696 = ~n41555 & ~n45695;
  assign n45697 = ~i_hlock6 & ~n45696;
  assign n45698 = ~n45694 & ~n45697;
  assign n45699 = controllable_hgrant6 & ~n45698;
  assign n45700 = ~n45116 & ~n45699;
  assign n45701 = controllable_hmaster0 & ~n45700;
  assign n45702 = ~n8217 & ~n30262;
  assign n45703 = ~n42153 & ~n45702;
  assign n45704 = i_hlock6 & ~n45703;
  assign n45705 = ~n8217 & ~n30365;
  assign n45706 = ~n42153 & ~n45705;
  assign n45707 = ~i_hlock6 & ~n45706;
  assign n45708 = ~n45704 & ~n45707;
  assign n45709 = controllable_hgrant6 & ~n45708;
  assign n45710 = ~n43865 & ~n45709;
  assign n45711 = ~controllable_hmaster0 & ~n45710;
  assign n45712 = ~n45701 & ~n45711;
  assign n45713 = i_hlock8 & ~n45712;
  assign n45714 = ~n8217 & ~n30275;
  assign n45715 = ~n42175 & ~n45714;
  assign n45716 = i_hlock6 & ~n45715;
  assign n45717 = ~n8217 & ~n30378;
  assign n45718 = ~n42175 & ~n45717;
  assign n45719 = ~i_hlock6 & ~n45718;
  assign n45720 = ~n45716 & ~n45719;
  assign n45721 = controllable_hgrant6 & ~n45720;
  assign n45722 = ~n43898 & ~n45721;
  assign n45723 = ~controllable_hmaster0 & ~n45722;
  assign n45724 = ~n45701 & ~n45723;
  assign n45725 = ~i_hlock8 & ~n45724;
  assign n45726 = ~n45713 & ~n45725;
  assign n45727 = controllable_hmaster3 & ~n45726;
  assign n45728 = ~n8217 & ~n37181;
  assign n45729 = ~n43905 & ~n45728;
  assign n45730 = i_hlock6 & ~n45729;
  assign n45731 = ~n8217 & ~n37189;
  assign n45732 = ~n43905 & ~n45731;
  assign n45733 = ~i_hlock6 & ~n45732;
  assign n45734 = ~n45730 & ~n45733;
  assign n45735 = controllable_hgrant6 & ~n45734;
  assign n45736 = ~n43993 & ~n45735;
  assign n45737 = controllable_hmaster0 & ~n45736;
  assign n45738 = ~n28973 & ~n30312;
  assign n45739 = controllable_hmaster1 & ~n45738;
  assign n45740 = ~n30329 & ~n45739;
  assign n45741 = ~n8217 & ~n45740;
  assign n45742 = ~n43999 & ~n45741;
  assign n45743 = i_hlock6 & ~n45742;
  assign n45744 = ~n28998 & ~n30415;
  assign n45745 = controllable_hmaster1 & ~n45744;
  assign n45746 = ~n30432 & ~n45745;
  assign n45747 = ~n8217 & ~n45746;
  assign n45748 = ~n44009 & ~n45747;
  assign n45749 = ~i_hlock6 & ~n45748;
  assign n45750 = ~n45743 & ~n45749;
  assign n45751 = controllable_hgrant6 & ~n45750;
  assign n45752 = ~n44051 & ~n45428;
  assign n45753 = controllable_hmaster1 & ~n45752;
  assign n45754 = ~n44103 & ~n45753;
  assign n45755 = i_hlock6 & ~n45754;
  assign n45756 = ~n44051 & ~n45442;
  assign n45757 = controllable_hmaster1 & ~n45756;
  assign n45758 = ~n44103 & ~n45757;
  assign n45759 = ~i_hlock6 & ~n45758;
  assign n45760 = ~n45755 & ~n45759;
  assign n45761 = ~controllable_hgrant6 & ~n45760;
  assign n45762 = ~n45751 & ~n45761;
  assign n45763 = ~controllable_hmaster0 & ~n45762;
  assign n45764 = ~n45737 & ~n45763;
  assign n45765 = ~controllable_hmaster3 & ~n45764;
  assign n45766 = ~n45727 & ~n45765;
  assign n45767 = i_hlock7 & ~n45766;
  assign n45768 = ~n8217 & ~n37201;
  assign n45769 = ~n44119 & ~n45768;
  assign n45770 = i_hlock6 & ~n45769;
  assign n45771 = ~n8217 & ~n37209;
  assign n45772 = ~n44119 & ~n45771;
  assign n45773 = ~i_hlock6 & ~n45772;
  assign n45774 = ~n45770 & ~n45773;
  assign n45775 = controllable_hgrant6 & ~n45774;
  assign n45776 = ~n44126 & ~n45775;
  assign n45777 = controllable_hmaster0 & ~n45776;
  assign n45778 = ~n45763 & ~n45777;
  assign n45779 = ~controllable_hmaster3 & ~n45778;
  assign n45780 = ~n45727 & ~n45779;
  assign n45781 = ~i_hlock7 & ~n45780;
  assign n45782 = ~n45767 & ~n45781;
  assign n45783 = i_hbusreq7 & ~n45782;
  assign n45784 = i_hbusreq8 & ~n45726;
  assign n45785 = i_hbusreq6 & ~n45698;
  assign n45786 = n8217 & ~n27489;
  assign n45787 = ~n8217 & ~n30482;
  assign n45788 = ~n45786 & ~n45787;
  assign n45789 = i_hlock6 & ~n45788;
  assign n45790 = ~n8217 & ~n30690;
  assign n45791 = ~n45786 & ~n45790;
  assign n45792 = ~i_hlock6 & ~n45791;
  assign n45793 = ~n45789 & ~n45792;
  assign n45794 = ~i_hbusreq6 & ~n45793;
  assign n45795 = ~n45785 & ~n45794;
  assign n45796 = controllable_hgrant6 & ~n45795;
  assign n45797 = ~n45215 & ~n45796;
  assign n45798 = controllable_hmaster0 & ~n45797;
  assign n45799 = i_hbusreq6 & ~n45708;
  assign n45800 = n8217 & ~n14046;
  assign n45801 = ~n8217 & ~n30505;
  assign n45802 = ~n45800 & ~n45801;
  assign n45803 = i_hlock6 & ~n45802;
  assign n45804 = ~n8217 & ~n30713;
  assign n45805 = ~n45800 & ~n45804;
  assign n45806 = ~i_hlock6 & ~n45805;
  assign n45807 = ~n45803 & ~n45806;
  assign n45808 = ~i_hbusreq6 & ~n45807;
  assign n45809 = ~n45799 & ~n45808;
  assign n45810 = controllable_hgrant6 & ~n45809;
  assign n45811 = ~n44437 & ~n45810;
  assign n45812 = ~controllable_hmaster0 & ~n45811;
  assign n45813 = ~n45798 & ~n45812;
  assign n45814 = i_hlock8 & ~n45813;
  assign n45815 = i_hbusreq6 & ~n45720;
  assign n45816 = n8217 & ~n14081;
  assign n45817 = ~n8217 & ~n30530;
  assign n45818 = ~n45816 & ~n45817;
  assign n45819 = i_hlock6 & ~n45818;
  assign n45820 = ~n8217 & ~n30738;
  assign n45821 = ~n45816 & ~n45820;
  assign n45822 = ~i_hlock6 & ~n45821;
  assign n45823 = ~n45819 & ~n45822;
  assign n45824 = ~i_hbusreq6 & ~n45823;
  assign n45825 = ~n45815 & ~n45824;
  assign n45826 = controllable_hgrant6 & ~n45825;
  assign n45827 = ~n44511 & ~n45826;
  assign n45828 = ~controllable_hmaster0 & ~n45827;
  assign n45829 = ~n45798 & ~n45828;
  assign n45830 = ~i_hlock8 & ~n45829;
  assign n45831 = ~n45814 & ~n45830;
  assign n45832 = ~i_hbusreq8 & ~n45831;
  assign n45833 = ~n45784 & ~n45832;
  assign n45834 = controllable_hmaster3 & ~n45833;
  assign n45835 = i_hbusreq8 & ~n45764;
  assign n45836 = i_hbusreq6 & ~n45734;
  assign n45837 = n8217 & ~n14167;
  assign n45838 = ~n8217 & ~n37250;
  assign n45839 = ~n45837 & ~n45838;
  assign n45840 = i_hlock6 & ~n45839;
  assign n45841 = ~n8217 & ~n37261;
  assign n45842 = ~n45837 & ~n45841;
  assign n45843 = ~i_hlock6 & ~n45842;
  assign n45844 = ~n45840 & ~n45843;
  assign n45845 = ~i_hbusreq6 & ~n45844;
  assign n45846 = ~n45836 & ~n45845;
  assign n45847 = controllable_hgrant6 & ~n45846;
  assign n45848 = ~n44675 & ~n45847;
  assign n45849 = controllable_hmaster0 & ~n45848;
  assign n45850 = i_hbusreq6 & ~n45750;
  assign n45851 = ~n14203 & ~n26783;
  assign n45852 = controllable_hmaster1 & ~n45851;
  assign n45853 = ~n14277 & ~n45852;
  assign n45854 = n8217 & ~n45853;
  assign n45855 = ~n29051 & ~n30606;
  assign n45856 = controllable_hmaster1 & ~n45855;
  assign n45857 = ~n30638 & ~n45856;
  assign n45858 = ~n8217 & ~n45857;
  assign n45859 = ~n45854 & ~n45858;
  assign n45860 = i_hlock6 & ~n45859;
  assign n45861 = ~n14203 & ~n26814;
  assign n45862 = controllable_hmaster1 & ~n45861;
  assign n45863 = ~n14277 & ~n45862;
  assign n45864 = n8217 & ~n45863;
  assign n45865 = ~n29106 & ~n30814;
  assign n45866 = controllable_hmaster1 & ~n45865;
  assign n45867 = ~n30846 & ~n45866;
  assign n45868 = ~n8217 & ~n45867;
  assign n45869 = ~n45864 & ~n45868;
  assign n45870 = ~i_hlock6 & ~n45869;
  assign n45871 = ~n45860 & ~n45870;
  assign n45872 = ~i_hbusreq6 & ~n45871;
  assign n45873 = ~n45850 & ~n45872;
  assign n45874 = controllable_hgrant6 & ~n45873;
  assign n45875 = i_hbusreq6 & ~n45760;
  assign n45876 = ~n44776 & ~n45473;
  assign n45877 = controllable_hmaster1 & ~n45876;
  assign n45878 = ~n44893 & ~n45877;
  assign n45879 = i_hlock6 & ~n45878;
  assign n45880 = ~n44776 & ~n45497;
  assign n45881 = controllable_hmaster1 & ~n45880;
  assign n45882 = ~n44893 & ~n45881;
  assign n45883 = ~i_hlock6 & ~n45882;
  assign n45884 = ~n45879 & ~n45883;
  assign n45885 = ~i_hbusreq6 & ~n45884;
  assign n45886 = ~n45875 & ~n45885;
  assign n45887 = ~controllable_hgrant6 & ~n45886;
  assign n45888 = ~n45874 & ~n45887;
  assign n45889 = ~controllable_hmaster0 & ~n45888;
  assign n45890 = ~n45849 & ~n45889;
  assign n45891 = ~i_hbusreq8 & ~n45890;
  assign n45892 = ~n45835 & ~n45891;
  assign n45893 = ~controllable_hmaster3 & ~n45892;
  assign n45894 = ~n45834 & ~n45893;
  assign n45895 = i_hlock7 & ~n45894;
  assign n45896 = i_hbusreq8 & ~n45778;
  assign n45897 = i_hbusreq6 & ~n45774;
  assign n45898 = n8217 & ~n14302;
  assign n45899 = ~n8217 & ~n37279;
  assign n45900 = ~n45898 & ~n45899;
  assign n45901 = i_hlock6 & ~n45900;
  assign n45902 = ~n8217 & ~n37290;
  assign n45903 = ~n45898 & ~n45902;
  assign n45904 = ~i_hlock6 & ~n45903;
  assign n45905 = ~n45901 & ~n45904;
  assign n45906 = ~i_hbusreq6 & ~n45905;
  assign n45907 = ~n45897 & ~n45906;
  assign n45908 = controllable_hgrant6 & ~n45907;
  assign n45909 = ~n44927 & ~n45908;
  assign n45910 = controllable_hmaster0 & ~n45909;
  assign n45911 = ~n45889 & ~n45910;
  assign n45912 = ~i_hbusreq8 & ~n45911;
  assign n45913 = ~n45896 & ~n45912;
  assign n45914 = ~controllable_hmaster3 & ~n45913;
  assign n45915 = ~n45834 & ~n45914;
  assign n45916 = ~i_hlock7 & ~n45915;
  assign n45917 = ~n45895 & ~n45916;
  assign n45918 = ~i_hbusreq7 & ~n45917;
  assign n45919 = ~n45783 & ~n45918;
  assign n45920 = n7924 & ~n45919;
  assign n45921 = ~n45691 & ~n45920;
  assign n45922 = n8214 & ~n45921;
  assign n45923 = ~n45517 & ~n45922;
  assign n45924 = n8202 & ~n45923;
  assign n45925 = ~n45325 & ~n45924;
  assign n45926 = n7920 & ~n45925;
  assign n45927 = ~n40788 & ~n45926;
  assign n45928 = ~n7728 & ~n45927;
  assign n45929 = ~n42702 & ~n45928;
  assign n45930 = n7723 & ~n45929;
  assign n45931 = ~n7723 & ~n45927;
  assign n45932 = ~n45930 & ~n45931;
  assign n45933 = n7714 & ~n45932;
  assign n45934 = n7723 & ~n45927;
  assign n45935 = ~n8217 & ~n30980;
  assign n45936 = ~n41555 & ~n45935;
  assign n45937 = i_hlock6 & ~n45936;
  assign n45938 = ~n8217 & ~n31087;
  assign n45939 = ~n41555 & ~n45938;
  assign n45940 = ~i_hlock6 & ~n45939;
  assign n45941 = ~n45937 & ~n45940;
  assign n45942 = controllable_hgrant6 & ~n45941;
  assign n45943 = ~n8378 & ~n30973;
  assign n45944 = ~n43743 & ~n45943;
  assign n45945 = i_hlock5 & ~n45944;
  assign n45946 = ~n8378 & ~n31080;
  assign n45947 = ~n43743 & ~n45946;
  assign n45948 = ~i_hlock5 & ~n45947;
  assign n45949 = ~n45945 & ~n45948;
  assign n45950 = controllable_hgrant5 & ~n45949;
  assign n45951 = ~n8426 & ~n20622;
  assign n45952 = ~n43747 & ~n45951;
  assign n45953 = i_hlock4 & ~n45952;
  assign n45954 = ~n8426 & ~n20635;
  assign n45955 = ~n43747 & ~n45954;
  assign n45956 = ~i_hlock4 & ~n45955;
  assign n45957 = ~n45953 & ~n45956;
  assign n45958 = controllable_hgrant4 & ~n45957;
  assign n45959 = ~n8365 & ~n20620;
  assign n45960 = ~n43751 & ~n45959;
  assign n45961 = i_hlock3 & ~n45960;
  assign n45962 = ~n8365 & ~n20633;
  assign n45963 = ~n43751 & ~n45962;
  assign n45964 = ~i_hlock3 & ~n45963;
  assign n45965 = ~n45961 & ~n45964;
  assign n45966 = controllable_hgrant3 & ~n45965;
  assign n45967 = ~n8389 & ~n20618;
  assign n45968 = ~n43755 & ~n45967;
  assign n45969 = i_hlock1 & ~n45968;
  assign n45970 = ~n8389 & ~n20631;
  assign n45971 = ~n43755 & ~n45970;
  assign n45972 = ~i_hlock1 & ~n45971;
  assign n45973 = ~n45969 & ~n45972;
  assign n45974 = controllable_hgrant1 & ~n45973;
  assign n45975 = ~i_hready & ~n8404;
  assign n45976 = ~n8404 & ~n45975;
  assign n45977 = controllable_ndecide & ~n45976;
  assign n45978 = i_hready & n8404;
  assign n45979 = ~controllable_ndecide & n45978;
  assign n45980 = ~n45977 & ~n45979;
  assign n45981 = controllable_locked & ~n45980;
  assign n45982 = ~n43759 & ~n45981;
  assign n45983 = i_hlock2 & ~n45982;
  assign n45984 = ~n7734 & ~n45977;
  assign n45985 = controllable_locked & ~n45984;
  assign n45986 = ~n43759 & ~n45985;
  assign n45987 = ~i_hlock2 & ~n45986;
  assign n45988 = ~n45983 & ~n45987;
  assign n45989 = controllable_hgrant2 & ~n45988;
  assign n45990 = ~n20645 & ~n45989;
  assign n45991 = n7733 & ~n45990;
  assign n45992 = ~n43762 & ~n45991;
  assign n45993 = n7928 & ~n45992;
  assign n45994 = ~n42723 & ~n45993;
  assign n45995 = ~controllable_hgrant1 & ~n45994;
  assign n45996 = ~n45974 & ~n45995;
  assign n45997 = ~controllable_hgrant3 & ~n45996;
  assign n45998 = ~n45966 & ~n45997;
  assign n45999 = ~controllable_hgrant4 & ~n45998;
  assign n46000 = ~n45958 & ~n45999;
  assign n46001 = ~controllable_hgrant5 & ~n46000;
  assign n46002 = ~n45950 & ~n46001;
  assign n46003 = controllable_hmaster1 & ~n46002;
  assign n46004 = controllable_hmaster2 & ~n46002;
  assign n46005 = ~n8378 & ~n30245;
  assign n46006 = ~n41580 & ~n46005;
  assign n46007 = i_hlock5 & ~n46006;
  assign n46008 = ~n8378 & ~n30348;
  assign n46009 = ~n41580 & ~n46008;
  assign n46010 = ~i_hlock5 & ~n46009;
  assign n46011 = ~n46007 & ~n46010;
  assign n46012 = controllable_hgrant5 & ~n46011;
  assign n46013 = ~n8426 & ~n18534;
  assign n46014 = ~n41584 & ~n46013;
  assign n46015 = i_hlock9 & ~n46014;
  assign n46016 = ~n8426 & ~n18560;
  assign n46017 = ~n41588 & ~n46016;
  assign n46018 = ~i_hlock9 & ~n46017;
  assign n46019 = ~n46015 & ~n46018;
  assign n46020 = i_hlock4 & ~n46019;
  assign n46021 = ~n8426 & ~n18540;
  assign n46022 = ~n41584 & ~n46021;
  assign n46023 = i_hlock9 & ~n46022;
  assign n46024 = ~n8426 & ~n18566;
  assign n46025 = ~n41588 & ~n46024;
  assign n46026 = ~i_hlock9 & ~n46025;
  assign n46027 = ~n46023 & ~n46026;
  assign n46028 = ~i_hlock4 & ~n46027;
  assign n46029 = ~n46020 & ~n46028;
  assign n46030 = controllable_hgrant4 & ~n46029;
  assign n46031 = ~n8365 & ~n18532;
  assign n46032 = ~n41594 & ~n46031;
  assign n46033 = i_hlock3 & ~n46032;
  assign n46034 = ~n8365 & ~n18538;
  assign n46035 = ~n41594 & ~n46034;
  assign n46036 = ~i_hlock3 & ~n46035;
  assign n46037 = ~n46033 & ~n46036;
  assign n46038 = controllable_hgrant3 & ~n46037;
  assign n46039 = ~n8389 & ~n18530;
  assign n46040 = ~n41598 & ~n46039;
  assign n46041 = i_hlock1 & ~n46040;
  assign n46042 = ~n8389 & ~n18536;
  assign n46043 = ~n41598 & ~n46042;
  assign n46044 = ~i_hlock1 & ~n46043;
  assign n46045 = ~n46041 & ~n46044;
  assign n46046 = controllable_hgrant1 & ~n46045;
  assign n46047 = controllable_hmastlock & ~n45980;
  assign n46048 = ~n39846 & ~n45979;
  assign n46049 = ~controllable_hmastlock & ~n46048;
  assign n46050 = ~n46047 & ~n46049;
  assign n46051 = controllable_locked & ~n46050;
  assign n46052 = ~n43759 & ~n46051;
  assign n46053 = i_hlock2 & ~n46052;
  assign n46054 = controllable_hmastlock & ~n45984;
  assign n46055 = ~n44281 & ~n46054;
  assign n46056 = controllable_locked & ~n46055;
  assign n46057 = ~n43759 & ~n46056;
  assign n46058 = ~i_hlock2 & ~n46057;
  assign n46059 = ~n46053 & ~n46058;
  assign n46060 = controllable_hgrant2 & ~n46059;
  assign n46061 = n7733 & n46060;
  assign n46062 = ~n43762 & ~n46061;
  assign n46063 = n7928 & ~n46062;
  assign n46064 = ~n8221 & ~n46063;
  assign n46065 = ~controllable_hgrant1 & ~n46064;
  assign n46066 = ~n46046 & ~n46065;
  assign n46067 = ~controllable_hgrant3 & ~n46066;
  assign n46068 = ~n46038 & ~n46067;
  assign n46069 = i_hlock9 & ~n46068;
  assign n46070 = ~n8365 & ~n18558;
  assign n46071 = ~n41620 & ~n46070;
  assign n46072 = i_hlock3 & ~n46071;
  assign n46073 = ~n8365 & ~n18564;
  assign n46074 = ~n41620 & ~n46073;
  assign n46075 = ~i_hlock3 & ~n46074;
  assign n46076 = ~n46072 & ~n46075;
  assign n46077 = controllable_hgrant3 & ~n46076;
  assign n46078 = ~n8389 & ~n18556;
  assign n46079 = ~n41624 & ~n46078;
  assign n46080 = i_hlock1 & ~n46079;
  assign n46081 = ~n8389 & ~n18562;
  assign n46082 = ~n41624 & ~n46081;
  assign n46083 = ~i_hlock1 & ~n46082;
  assign n46084 = ~n46080 & ~n46083;
  assign n46085 = controllable_hgrant1 & ~n46084;
  assign n46086 = ~n8235 & ~n46063;
  assign n46087 = ~controllable_hgrant1 & ~n46086;
  assign n46088 = ~n46085 & ~n46087;
  assign n46089 = ~controllable_hgrant3 & ~n46088;
  assign n46090 = ~n46077 & ~n46089;
  assign n46091 = ~i_hlock9 & ~n46090;
  assign n46092 = ~n46069 & ~n46091;
  assign n46093 = ~controllable_hgrant4 & ~n46092;
  assign n46094 = ~n46030 & ~n46093;
  assign n46095 = ~controllable_hgrant5 & ~n46094;
  assign n46096 = ~n46012 & ~n46095;
  assign n46097 = ~controllable_hmaster2 & ~n46096;
  assign n46098 = ~n46004 & ~n46097;
  assign n46099 = ~controllable_hmaster1 & ~n46098;
  assign n46100 = ~n46003 & ~n46099;
  assign n46101 = ~controllable_hgrant6 & ~n46100;
  assign n46102 = ~n45942 & ~n46101;
  assign n46103 = controllable_hmaster0 & ~n46102;
  assign n46104 = ~n8217 & ~n30991;
  assign n46105 = ~n42153 & ~n46104;
  assign n46106 = i_hlock6 & ~n46105;
  assign n46107 = ~n8217 & ~n31098;
  assign n46108 = ~n42153 & ~n46107;
  assign n46109 = ~i_hlock6 & ~n46108;
  assign n46110 = ~n46106 & ~n46109;
  assign n46111 = controllable_hgrant6 & ~n46110;
  assign n46112 = ~n8378 & ~n30985;
  assign n46113 = ~n42157 & ~n46112;
  assign n46114 = i_hlock5 & ~n46113;
  assign n46115 = ~n8378 & ~n31092;
  assign n46116 = ~n42157 & ~n46115;
  assign n46117 = ~i_hlock5 & ~n46116;
  assign n46118 = ~n46114 & ~n46117;
  assign n46119 = controllable_hgrant5 & ~n46118;
  assign n46120 = ~n8426 & ~n20705;
  assign n46121 = ~n41584 & ~n46120;
  assign n46122 = i_hlock4 & ~n46121;
  assign n46123 = ~n8426 & ~n20711;
  assign n46124 = ~n41584 & ~n46123;
  assign n46125 = ~i_hlock4 & ~n46124;
  assign n46126 = ~n46122 & ~n46125;
  assign n46127 = controllable_hgrant4 & ~n46126;
  assign n46128 = ~n8365 & ~n20703;
  assign n46129 = ~n41594 & ~n46128;
  assign n46130 = i_hlock3 & ~n46129;
  assign n46131 = ~n8365 & ~n20709;
  assign n46132 = ~n41594 & ~n46131;
  assign n46133 = ~i_hlock3 & ~n46132;
  assign n46134 = ~n46130 & ~n46133;
  assign n46135 = controllable_hgrant3 & ~n46134;
  assign n46136 = ~n8389 & ~n20701;
  assign n46137 = ~n41598 & ~n46136;
  assign n46138 = i_hlock1 & ~n46137;
  assign n46139 = ~n8389 & ~n20707;
  assign n46140 = ~n41598 & ~n46139;
  assign n46141 = ~i_hlock1 & ~n46140;
  assign n46142 = ~n46138 & ~n46141;
  assign n46143 = controllable_hgrant1 & ~n46142;
  assign n46144 = ~n20613 & ~n45989;
  assign n46145 = n7733 & ~n46144;
  assign n46146 = ~n43847 & ~n46145;
  assign n46147 = n7928 & ~n46146;
  assign n46148 = ~n8221 & ~n46147;
  assign n46149 = ~controllable_hgrant1 & ~n46148;
  assign n46150 = ~n46143 & ~n46149;
  assign n46151 = ~controllable_hgrant3 & ~n46150;
  assign n46152 = ~n46135 & ~n46151;
  assign n46153 = ~controllable_hgrant4 & ~n46152;
  assign n46154 = ~n46127 & ~n46153;
  assign n46155 = ~controllable_hgrant5 & ~n46154;
  assign n46156 = ~n46119 & ~n46155;
  assign n46157 = ~controllable_hmaster2 & ~n46156;
  assign n46158 = ~n46004 & ~n46157;
  assign n46159 = ~controllable_hmaster1 & ~n46158;
  assign n46160 = ~n46003 & ~n46159;
  assign n46161 = ~controllable_hgrant6 & ~n46160;
  assign n46162 = ~n46111 & ~n46161;
  assign n46163 = ~controllable_hmaster0 & ~n46162;
  assign n46164 = ~n46103 & ~n46163;
  assign n46165 = i_hlock8 & ~n46164;
  assign n46166 = ~n8217 & ~n31004;
  assign n46167 = ~n42175 & ~n46166;
  assign n46168 = i_hlock6 & ~n46167;
  assign n46169 = ~n8217 & ~n31111;
  assign n46170 = ~n42175 & ~n46169;
  assign n46171 = ~i_hlock6 & ~n46170;
  assign n46172 = ~n46168 & ~n46171;
  assign n46173 = controllable_hgrant6 & ~n46172;
  assign n46174 = ~n8378 & ~n30998;
  assign n46175 = ~n42179 & ~n46174;
  assign n46176 = i_hlock5 & ~n46175;
  assign n46177 = ~n8378 & ~n31105;
  assign n46178 = ~n42179 & ~n46177;
  assign n46179 = ~i_hlock5 & ~n46178;
  assign n46180 = ~n46176 & ~n46179;
  assign n46181 = controllable_hgrant5 & ~n46180;
  assign n46182 = ~n8426 & ~n20747;
  assign n46183 = ~n41588 & ~n46182;
  assign n46184 = i_hlock4 & ~n46183;
  assign n46185 = ~n8426 & ~n20750;
  assign n46186 = ~n41588 & ~n46185;
  assign n46187 = ~i_hlock4 & ~n46186;
  assign n46188 = ~n46184 & ~n46187;
  assign n46189 = controllable_hgrant4 & ~n46188;
  assign n46190 = ~n8365 & ~n20722;
  assign n46191 = ~n41620 & ~n46190;
  assign n46192 = i_hlock3 & ~n46191;
  assign n46193 = ~n8365 & ~n20731;
  assign n46194 = ~n41620 & ~n46193;
  assign n46195 = ~i_hlock3 & ~n46194;
  assign n46196 = ~n46192 & ~n46195;
  assign n46197 = controllable_hgrant3 & ~n46196;
  assign n46198 = ~n8389 & ~n20720;
  assign n46199 = ~n41624 & ~n46198;
  assign n46200 = i_hlock1 & ~n46199;
  assign n46201 = ~n8389 & ~n20729;
  assign n46202 = ~n41624 & ~n46201;
  assign n46203 = ~i_hlock1 & ~n46202;
  assign n46204 = ~n46200 & ~n46203;
  assign n46205 = controllable_hgrant1 & ~n46204;
  assign n46206 = ~n8235 & ~n46147;
  assign n46207 = ~controllable_hgrant1 & ~n46206;
  assign n46208 = ~n46205 & ~n46207;
  assign n46209 = ~controllable_hgrant3 & ~n46208;
  assign n46210 = ~n46197 & ~n46209;
  assign n46211 = ~controllable_hgrant4 & ~n46210;
  assign n46212 = ~n46189 & ~n46211;
  assign n46213 = ~controllable_hgrant5 & ~n46212;
  assign n46214 = ~n46181 & ~n46213;
  assign n46215 = ~controllable_hmaster2 & ~n46214;
  assign n46216 = ~n46004 & ~n46215;
  assign n46217 = ~controllable_hmaster1 & ~n46216;
  assign n46218 = ~n46003 & ~n46217;
  assign n46219 = ~controllable_hgrant6 & ~n46218;
  assign n46220 = ~n46173 & ~n46219;
  assign n46221 = ~controllable_hmaster0 & ~n46220;
  assign n46222 = ~n46103 & ~n46221;
  assign n46223 = ~i_hlock8 & ~n46222;
  assign n46224 = ~n46165 & ~n46223;
  assign n46225 = controllable_hmaster3 & ~n46224;
  assign n46226 = ~n8217 & ~n37436;
  assign n46227 = ~n43905 & ~n46226;
  assign n46228 = i_hlock6 & ~n46227;
  assign n46229 = ~n8217 & ~n37444;
  assign n46230 = ~n43905 & ~n46229;
  assign n46231 = ~i_hlock6 & ~n46230;
  assign n46232 = ~n46228 & ~n46231;
  assign n46233 = controllable_hgrant6 & ~n46232;
  assign n46234 = controllable_hmaster2 & ~n46156;
  assign n46235 = ~n8378 & ~n31018;
  assign n46236 = ~n43910 & ~n46235;
  assign n46237 = i_hlock5 & ~n46236;
  assign n46238 = ~n8378 & ~n31125;
  assign n46239 = ~n43910 & ~n46238;
  assign n46240 = ~i_hlock5 & ~n46239;
  assign n46241 = ~n46237 & ~n46240;
  assign n46242 = controllable_hgrant5 & ~n46241;
  assign n46243 = ~n8426 & ~n20726;
  assign n46244 = ~n43914 & ~n46243;
  assign n46245 = i_hlock4 & ~n46244;
  assign n46246 = ~n8426 & ~n20735;
  assign n46247 = ~n43914 & ~n46246;
  assign n46248 = ~i_hlock4 & ~n46247;
  assign n46249 = ~n46245 & ~n46248;
  assign n46250 = controllable_hgrant4 & ~n46249;
  assign n46251 = ~n8365 & ~n20652;
  assign n46252 = ~n43918 & ~n46251;
  assign n46253 = i_hlock3 & ~n46252;
  assign n46254 = ~n8365 & ~n20667;
  assign n46255 = ~n43922 & ~n46254;
  assign n46256 = ~i_hlock3 & ~n46255;
  assign n46257 = ~n46253 & ~n46256;
  assign n46258 = controllable_hgrant3 & ~n46257;
  assign n46259 = i_hlock3 & ~n46150;
  assign n46260 = ~i_hlock3 & ~n46208;
  assign n46261 = ~n46259 & ~n46260;
  assign n46262 = ~controllable_hgrant3 & ~n46261;
  assign n46263 = ~n46258 & ~n46262;
  assign n46264 = ~controllable_hgrant4 & ~n46263;
  assign n46265 = ~n46250 & ~n46264;
  assign n46266 = ~controllable_hgrant5 & ~n46265;
  assign n46267 = ~n46242 & ~n46266;
  assign n46268 = ~controllable_hmaster2 & ~n46267;
  assign n46269 = ~n46234 & ~n46268;
  assign n46270 = controllable_hmaster1 & ~n46269;
  assign n46271 = ~n8378 & ~n31013;
  assign n46272 = ~n43940 & ~n46271;
  assign n46273 = i_hlock5 & ~n46272;
  assign n46274 = ~n8378 & ~n31120;
  assign n46275 = ~n43944 & ~n46274;
  assign n46276 = ~i_hlock5 & ~n46275;
  assign n46277 = ~n46273 & ~n46276;
  assign n46278 = controllable_hgrant5 & ~n46277;
  assign n46279 = i_hlock5 & ~n46154;
  assign n46280 = ~i_hlock5 & ~n46212;
  assign n46281 = ~n46279 & ~n46280;
  assign n46282 = ~controllable_hgrant5 & ~n46281;
  assign n46283 = ~n46278 & ~n46282;
  assign n46284 = controllable_hmaster2 & ~n46283;
  assign n46285 = ~n8378 & ~n31031;
  assign n46286 = ~n43956 & ~n46285;
  assign n46287 = i_hlock5 & ~n46286;
  assign n46288 = ~n8378 & ~n31138;
  assign n46289 = ~n43956 & ~n46288;
  assign n46290 = ~i_hlock5 & ~n46289;
  assign n46291 = ~n46287 & ~n46290;
  assign n46292 = controllable_hgrant5 & ~n46291;
  assign n46293 = ~n8426 & ~n20766;
  assign n46294 = ~n43960 & ~n46293;
  assign n46295 = i_hlock4 & ~n46294;
  assign n46296 = ~n8426 & ~n20774;
  assign n46297 = ~n43960 & ~n46296;
  assign n46298 = ~i_hlock4 & ~n46297;
  assign n46299 = ~n46295 & ~n46298;
  assign n46300 = controllable_hgrant4 & ~n46299;
  assign n46301 = ~n8365 & ~n20764;
  assign n46302 = ~n43964 & ~n46301;
  assign n46303 = i_hlock3 & ~n46302;
  assign n46304 = ~n8365 & ~n20772;
  assign n46305 = ~n43964 & ~n46304;
  assign n46306 = ~i_hlock3 & ~n46305;
  assign n46307 = ~n46303 & ~n46306;
  assign n46308 = controllable_hgrant3 & ~n46307;
  assign n46309 = ~n8389 & ~n20650;
  assign n46310 = ~n43968 & ~n46309;
  assign n46311 = i_hlock1 & ~n46310;
  assign n46312 = ~n8389 & ~n20665;
  assign n46313 = ~n43972 & ~n46312;
  assign n46314 = ~i_hlock1 & ~n46313;
  assign n46315 = ~n46311 & ~n46314;
  assign n46316 = controllable_hgrant1 & ~n46315;
  assign n46317 = i_hlock1 & ~n46148;
  assign n46318 = ~i_hlock1 & ~n46206;
  assign n46319 = ~n46317 & ~n46318;
  assign n46320 = ~controllable_hgrant1 & ~n46319;
  assign n46321 = ~n46316 & ~n46320;
  assign n46322 = ~controllable_hgrant3 & ~n46321;
  assign n46323 = ~n46308 & ~n46322;
  assign n46324 = ~controllable_hgrant4 & ~n46323;
  assign n46325 = ~n46300 & ~n46324;
  assign n46326 = ~controllable_hgrant5 & ~n46325;
  assign n46327 = ~n46292 & ~n46326;
  assign n46328 = ~controllable_hmaster2 & ~n46327;
  assign n46329 = ~n46284 & ~n46328;
  assign n46330 = ~controllable_hmaster1 & ~n46329;
  assign n46331 = ~n46270 & ~n46330;
  assign n46332 = ~controllable_hgrant6 & ~n46331;
  assign n46333 = ~n46233 & ~n46332;
  assign n46334 = controllable_hmaster0 & ~n46333;
  assign n46335 = ~n31016 & ~n31046;
  assign n46336 = controllable_hmaster1 & ~n46335;
  assign n46337 = ~n31063 & ~n46336;
  assign n46338 = ~n8217 & ~n46337;
  assign n46339 = ~n43999 & ~n46338;
  assign n46340 = i_hlock6 & ~n46339;
  assign n46341 = ~n31123 & ~n31153;
  assign n46342 = controllable_hmaster1 & ~n46341;
  assign n46343 = ~n31170 & ~n46342;
  assign n46344 = ~n8217 & ~n46343;
  assign n46345 = ~n44009 & ~n46344;
  assign n46346 = ~i_hlock6 & ~n46345;
  assign n46347 = ~n46340 & ~n46346;
  assign n46348 = controllable_hgrant6 & ~n46347;
  assign n46349 = ~n8378 & ~n31043;
  assign n46350 = ~n44018 & ~n46349;
  assign n46351 = i_hlock5 & ~n46350;
  assign n46352 = ~n8378 & ~n31150;
  assign n46353 = ~n44018 & ~n46352;
  assign n46354 = ~i_hlock5 & ~n46353;
  assign n46355 = ~n46351 & ~n46354;
  assign n46356 = controllable_hgrant5 & ~n46355;
  assign n46357 = ~n8426 & ~n20792;
  assign n46358 = ~n44022 & ~n46357;
  assign n46359 = i_hlock4 & ~n46358;
  assign n46360 = ~n8426 & ~n20798;
  assign n46361 = ~n44022 & ~n46360;
  assign n46362 = ~i_hlock4 & ~n46361;
  assign n46363 = ~n46359 & ~n46362;
  assign n46364 = controllable_hgrant4 & ~n46363;
  assign n46365 = ~n8365 & ~n20790;
  assign n46366 = ~n44026 & ~n46365;
  assign n46367 = i_hlock3 & ~n46366;
  assign n46368 = ~n8365 & ~n20796;
  assign n46369 = ~n44026 & ~n46368;
  assign n46370 = ~i_hlock3 & ~n46369;
  assign n46371 = ~n46367 & ~n46370;
  assign n46372 = controllable_hgrant3 & ~n46371;
  assign n46373 = ~n8389 & ~n20788;
  assign n46374 = ~n44030 & ~n46373;
  assign n46375 = i_hlock1 & ~n46374;
  assign n46376 = ~n8389 & ~n20794;
  assign n46377 = ~n44030 & ~n46376;
  assign n46378 = ~i_hlock1 & ~n46377;
  assign n46379 = ~n46375 & ~n46378;
  assign n46380 = controllable_hgrant1 & ~n46379;
  assign n46381 = ~controllable_hmastlock & ~n45980;
  assign n46382 = ~n42945 & ~n46381;
  assign n46383 = controllable_locked & ~n46382;
  assign n46384 = ~n43759 & ~n46383;
  assign n46385 = i_hlock2 & ~n46384;
  assign n46386 = ~controllable_hmastlock & ~n45984;
  assign n46387 = ~n42945 & ~n46386;
  assign n46388 = controllable_locked & ~n46387;
  assign n46389 = ~n43759 & ~n46388;
  assign n46390 = ~i_hlock2 & ~n46389;
  assign n46391 = ~n46385 & ~n46390;
  assign n46392 = controllable_hgrant2 & ~n46391;
  assign n46393 = ~n20613 & ~n46392;
  assign n46394 = n7733 & ~n46393;
  assign n46395 = ~n44037 & ~n46394;
  assign n46396 = n7928 & ~n46395;
  assign n46397 = ~n42965 & ~n46396;
  assign n46398 = ~controllable_hgrant1 & ~n46397;
  assign n46399 = ~n46380 & ~n46398;
  assign n46400 = ~controllable_hgrant3 & ~n46399;
  assign n46401 = ~n46372 & ~n46400;
  assign n46402 = ~controllable_hgrant4 & ~n46401;
  assign n46403 = ~n46364 & ~n46402;
  assign n46404 = ~controllable_hgrant5 & ~n46403;
  assign n46405 = ~n46356 & ~n46404;
  assign n46406 = ~controllable_hmaster2 & ~n46405;
  assign n46407 = ~n46234 & ~n46406;
  assign n46408 = controllable_hmaster1 & ~n46407;
  assign n46409 = ~n8378 & ~n31053;
  assign n46410 = ~n44054 & ~n46409;
  assign n46411 = i_hlock5 & ~n46410;
  assign n46412 = ~n8378 & ~n31160;
  assign n46413 = ~n44054 & ~n46412;
  assign n46414 = ~i_hlock5 & ~n46413;
  assign n46415 = ~n46411 & ~n46414;
  assign n46416 = controllable_hgrant5 & ~n46415;
  assign n46417 = ~n8426 & ~n20654;
  assign n46418 = ~n44058 & ~n46417;
  assign n46419 = i_hlock4 & ~n46418;
  assign n46420 = ~n8426 & ~n20669;
  assign n46421 = ~n44062 & ~n46420;
  assign n46422 = ~i_hlock4 & ~n46421;
  assign n46423 = ~n46419 & ~n46422;
  assign n46424 = controllable_hgrant4 & ~n46423;
  assign n46425 = i_hlock4 & ~n46152;
  assign n46426 = ~i_hlock4 & ~n46210;
  assign n46427 = ~n46425 & ~n46426;
  assign n46428 = ~controllable_hgrant4 & ~n46427;
  assign n46429 = ~n46424 & ~n46428;
  assign n46430 = ~controllable_hgrant5 & ~n46429;
  assign n46431 = ~n46416 & ~n46430;
  assign n46432 = controllable_hmaster2 & ~n46431;
  assign n46433 = ~n8378 & ~n31058;
  assign n46434 = ~n44076 & ~n46433;
  assign n46435 = i_hlock5 & ~n46434;
  assign n46436 = ~n8378 & ~n31165;
  assign n46437 = ~n44076 & ~n46436;
  assign n46438 = ~i_hlock5 & ~n46437;
  assign n46439 = ~n46435 & ~n46438;
  assign n46440 = controllable_hgrant5 & ~n46439;
  assign n46441 = ~n8426 & ~n20820;
  assign n46442 = ~n44080 & ~n46441;
  assign n46443 = i_hlock4 & ~n46442;
  assign n46444 = ~n8426 & ~n20826;
  assign n46445 = ~n44080 & ~n46444;
  assign n46446 = ~i_hlock4 & ~n46445;
  assign n46447 = ~n46443 & ~n46446;
  assign n46448 = controllable_hgrant4 & ~n46447;
  assign n46449 = ~n8365 & ~n20818;
  assign n46450 = ~n44084 & ~n46449;
  assign n46451 = i_hlock3 & ~n46450;
  assign n46452 = ~n8365 & ~n20824;
  assign n46453 = ~n44084 & ~n46452;
  assign n46454 = ~i_hlock3 & ~n46453;
  assign n46455 = ~n46451 & ~n46454;
  assign n46456 = controllable_hgrant3 & ~n46455;
  assign n46457 = ~n8389 & ~n20816;
  assign n46458 = ~n44088 & ~n46457;
  assign n46459 = i_hlock1 & ~n46458;
  assign n46460 = ~n8389 & ~n20822;
  assign n46461 = ~n44088 & ~n46460;
  assign n46462 = ~i_hlock1 & ~n46461;
  assign n46463 = ~n46459 & ~n46462;
  assign n46464 = controllable_hgrant1 & ~n46463;
  assign n46465 = ~n8440 & ~n46147;
  assign n46466 = ~controllable_hgrant1 & ~n46465;
  assign n46467 = ~n46464 & ~n46466;
  assign n46468 = ~controllable_hgrant3 & ~n46467;
  assign n46469 = ~n46456 & ~n46468;
  assign n46470 = ~controllable_hgrant4 & ~n46469;
  assign n46471 = ~n46448 & ~n46470;
  assign n46472 = ~controllable_hgrant5 & ~n46471;
  assign n46473 = ~n46440 & ~n46472;
  assign n46474 = ~controllable_hmaster2 & ~n46473;
  assign n46475 = ~n46432 & ~n46474;
  assign n46476 = ~controllable_hmaster1 & ~n46475;
  assign n46477 = ~n46408 & ~n46476;
  assign n46478 = i_hlock6 & ~n46477;
  assign n46479 = controllable_hmaster2 & ~n46214;
  assign n46480 = ~n46406 & ~n46479;
  assign n46481 = controllable_hmaster1 & ~n46480;
  assign n46482 = ~n46476 & ~n46481;
  assign n46483 = ~i_hlock6 & ~n46482;
  assign n46484 = ~n46478 & ~n46483;
  assign n46485 = ~controllable_hgrant6 & ~n46484;
  assign n46486 = ~n46348 & ~n46485;
  assign n46487 = ~controllable_hmaster0 & ~n46486;
  assign n46488 = ~n46334 & ~n46487;
  assign n46489 = ~controllable_hmaster3 & ~n46488;
  assign n46490 = ~n46225 & ~n46489;
  assign n46491 = i_hlock7 & ~n46490;
  assign n46492 = ~n8217 & ~n37456;
  assign n46493 = ~n44119 & ~n46492;
  assign n46494 = i_hlock6 & ~n46493;
  assign n46495 = ~n8217 & ~n37464;
  assign n46496 = ~n44119 & ~n46495;
  assign n46497 = ~i_hlock6 & ~n46496;
  assign n46498 = ~n46494 & ~n46497;
  assign n46499 = controllable_hgrant6 & ~n46498;
  assign n46500 = ~n46268 & ~n46479;
  assign n46501 = controllable_hmaster1 & ~n46500;
  assign n46502 = ~n46330 & ~n46501;
  assign n46503 = ~controllable_hgrant6 & ~n46502;
  assign n46504 = ~n46499 & ~n46503;
  assign n46505 = controllable_hmaster0 & ~n46504;
  assign n46506 = ~n46487 & ~n46505;
  assign n46507 = ~controllable_hmaster3 & ~n46506;
  assign n46508 = ~n46225 & ~n46507;
  assign n46509 = ~i_hlock7 & ~n46508;
  assign n46510 = ~n46491 & ~n46509;
  assign n46511 = i_hbusreq7 & ~n46510;
  assign n46512 = i_hbusreq8 & ~n46224;
  assign n46513 = i_hbusreq6 & ~n45941;
  assign n46514 = ~n8217 & ~n31220;
  assign n46515 = ~n44137 & ~n46514;
  assign n46516 = i_hlock6 & ~n46515;
  assign n46517 = ~n8217 & ~n31442;
  assign n46518 = ~n44137 & ~n46517;
  assign n46519 = ~i_hlock6 & ~n46518;
  assign n46520 = ~n46516 & ~n46519;
  assign n46521 = ~i_hbusreq6 & ~n46520;
  assign n46522 = ~n46513 & ~n46521;
  assign n46523 = controllable_hgrant6 & ~n46522;
  assign n46524 = i_hbusreq6 & ~n46100;
  assign n46525 = i_hbusreq5 & ~n45949;
  assign n46526 = ~n8378 & ~n31198;
  assign n46527 = ~n44145 & ~n46526;
  assign n46528 = i_hlock5 & ~n46527;
  assign n46529 = ~n8378 & ~n31420;
  assign n46530 = ~n44145 & ~n46529;
  assign n46531 = ~i_hlock5 & ~n46530;
  assign n46532 = ~n46528 & ~n46531;
  assign n46533 = ~i_hbusreq5 & ~n46532;
  assign n46534 = ~n46525 & ~n46533;
  assign n46535 = controllable_hgrant5 & ~n46534;
  assign n46536 = i_hbusreq5 & ~n46000;
  assign n46537 = i_hbusreq4 & ~n45957;
  assign n46538 = i_hbusreq9 & ~n45952;
  assign n46539 = ~n8426 & ~n20895;
  assign n46540 = ~n44154 & ~n46539;
  assign n46541 = ~i_hbusreq9 & ~n46540;
  assign n46542 = ~n46538 & ~n46541;
  assign n46543 = i_hlock4 & ~n46542;
  assign n46544 = i_hbusreq9 & ~n45955;
  assign n46545 = ~n8426 & ~n20917;
  assign n46546 = ~n44154 & ~n46545;
  assign n46547 = ~i_hbusreq9 & ~n46546;
  assign n46548 = ~n46544 & ~n46547;
  assign n46549 = ~i_hlock4 & ~n46548;
  assign n46550 = ~n46543 & ~n46549;
  assign n46551 = ~i_hbusreq4 & ~n46550;
  assign n46552 = ~n46537 & ~n46551;
  assign n46553 = controllable_hgrant4 & ~n46552;
  assign n46554 = i_hbusreq4 & ~n45998;
  assign n46555 = i_hbusreq9 & ~n45998;
  assign n46556 = i_hbusreq3 & ~n45965;
  assign n46557 = ~n8365 & ~n20891;
  assign n46558 = ~n44165 & ~n46557;
  assign n46559 = i_hlock3 & ~n46558;
  assign n46560 = ~n8365 & ~n20913;
  assign n46561 = ~n44165 & ~n46560;
  assign n46562 = ~i_hlock3 & ~n46561;
  assign n46563 = ~n46559 & ~n46562;
  assign n46564 = ~i_hbusreq3 & ~n46563;
  assign n46565 = ~n46556 & ~n46564;
  assign n46566 = controllable_hgrant3 & ~n46565;
  assign n46567 = i_hbusreq3 & ~n45996;
  assign n46568 = i_hbusreq1 & ~n45973;
  assign n46569 = ~n8389 & ~n20887;
  assign n46570 = ~n44173 & ~n46569;
  assign n46571 = i_hlock1 & ~n46570;
  assign n46572 = ~n8389 & ~n20909;
  assign n46573 = ~n44173 & ~n46572;
  assign n46574 = ~i_hlock1 & ~n46573;
  assign n46575 = ~n46571 & ~n46574;
  assign n46576 = ~i_hbusreq1 & ~n46575;
  assign n46577 = ~n46568 & ~n46576;
  assign n46578 = controllable_hgrant1 & ~n46577;
  assign n46579 = i_hbusreq1 & ~n45994;
  assign n46580 = i_hbusreq2 & ~n45988;
  assign n46581 = i_hbusreq0 & ~n45982;
  assign n46582 = controllable_ndecide & ~n45977;
  assign n46583 = controllable_locked & ~n46582;
  assign n46584 = ~n44182 & ~n46583;
  assign n46585 = i_hlock0 & ~n46584;
  assign n46586 = ~i_hlock0 & ~n45986;
  assign n46587 = ~n46585 & ~n46586;
  assign n46588 = ~i_hbusreq0 & ~n46587;
  assign n46589 = ~n46581 & ~n46588;
  assign n46590 = i_hlock2 & ~n46589;
  assign n46591 = i_hbusreq0 & ~n45986;
  assign n46592 = ~n46588 & ~n46591;
  assign n46593 = ~i_hlock2 & ~n46592;
  assign n46594 = ~n46590 & ~n46593;
  assign n46595 = ~i_hbusreq2 & ~n46594;
  assign n46596 = ~n46580 & ~n46595;
  assign n46597 = controllable_hgrant2 & ~n46596;
  assign n46598 = ~n20950 & ~n46597;
  assign n46599 = n7733 & ~n46598;
  assign n46600 = ~n44199 & ~n46599;
  assign n46601 = n7928 & ~n46600;
  assign n46602 = ~n43114 & ~n46601;
  assign n46603 = ~i_hbusreq1 & ~n46602;
  assign n46604 = ~n46579 & ~n46603;
  assign n46605 = ~controllable_hgrant1 & ~n46604;
  assign n46606 = ~n46578 & ~n46605;
  assign n46607 = ~i_hbusreq3 & ~n46606;
  assign n46608 = ~n46567 & ~n46607;
  assign n46609 = ~controllable_hgrant3 & ~n46608;
  assign n46610 = ~n46566 & ~n46609;
  assign n46611 = ~i_hbusreq9 & ~n46610;
  assign n46612 = ~n46555 & ~n46611;
  assign n46613 = ~i_hbusreq4 & ~n46612;
  assign n46614 = ~n46554 & ~n46613;
  assign n46615 = ~controllable_hgrant4 & ~n46614;
  assign n46616 = ~n46553 & ~n46615;
  assign n46617 = ~i_hbusreq5 & ~n46616;
  assign n46618 = ~n46536 & ~n46617;
  assign n46619 = ~controllable_hgrant5 & ~n46618;
  assign n46620 = ~n46535 & ~n46619;
  assign n46621 = controllable_hmaster1 & ~n46620;
  assign n46622 = controllable_hmaster2 & ~n46620;
  assign n46623 = i_hbusreq5 & ~n46011;
  assign n46624 = ~n8378 & ~n31212;
  assign n46625 = ~n44226 & ~n46624;
  assign n46626 = i_hlock5 & ~n46625;
  assign n46627 = ~n8378 & ~n31434;
  assign n46628 = ~n44226 & ~n46627;
  assign n46629 = ~i_hlock5 & ~n46628;
  assign n46630 = ~n46626 & ~n46629;
  assign n46631 = ~i_hbusreq5 & ~n46630;
  assign n46632 = ~n46623 & ~n46631;
  assign n46633 = controllable_hgrant5 & ~n46632;
  assign n46634 = i_hbusreq5 & ~n46094;
  assign n46635 = i_hbusreq4 & ~n46029;
  assign n46636 = i_hbusreq9 & ~n46019;
  assign n46637 = ~n8426 & ~n21030;
  assign n46638 = ~n44235 & ~n46637;
  assign n46639 = i_hlock9 & ~n46638;
  assign n46640 = ~n8426 & ~n21081;
  assign n46641 = ~n44239 & ~n46640;
  assign n46642 = ~i_hlock9 & ~n46641;
  assign n46643 = ~n46639 & ~n46642;
  assign n46644 = ~i_hbusreq9 & ~n46643;
  assign n46645 = ~n46636 & ~n46644;
  assign n46646 = i_hlock4 & ~n46645;
  assign n46647 = i_hbusreq9 & ~n46027;
  assign n46648 = ~n8426 & ~n21048;
  assign n46649 = ~n44235 & ~n46648;
  assign n46650 = i_hlock9 & ~n46649;
  assign n46651 = ~n8426 & ~n21091;
  assign n46652 = ~n44239 & ~n46651;
  assign n46653 = ~i_hlock9 & ~n46652;
  assign n46654 = ~n46650 & ~n46653;
  assign n46655 = ~i_hbusreq9 & ~n46654;
  assign n46656 = ~n46647 & ~n46655;
  assign n46657 = ~i_hlock4 & ~n46656;
  assign n46658 = ~n46646 & ~n46657;
  assign n46659 = ~i_hbusreq4 & ~n46658;
  assign n46660 = ~n46635 & ~n46659;
  assign n46661 = controllable_hgrant4 & ~n46660;
  assign n46662 = i_hbusreq4 & ~n46092;
  assign n46663 = i_hbusreq9 & ~n46092;
  assign n46664 = i_hbusreq3 & ~n46037;
  assign n46665 = ~n8365 & ~n21026;
  assign n46666 = ~n44252 & ~n46665;
  assign n46667 = i_hlock3 & ~n46666;
  assign n46668 = ~n8365 & ~n21044;
  assign n46669 = ~n44252 & ~n46668;
  assign n46670 = ~i_hlock3 & ~n46669;
  assign n46671 = ~n46667 & ~n46670;
  assign n46672 = ~i_hbusreq3 & ~n46671;
  assign n46673 = ~n46664 & ~n46672;
  assign n46674 = controllable_hgrant3 & ~n46673;
  assign n46675 = i_hbusreq3 & ~n46066;
  assign n46676 = i_hbusreq1 & ~n46045;
  assign n46677 = ~n8389 & ~n21022;
  assign n46678 = ~n44260 & ~n46677;
  assign n46679 = i_hlock1 & ~n46678;
  assign n46680 = ~n8389 & ~n21040;
  assign n46681 = ~n44260 & ~n46680;
  assign n46682 = ~i_hlock1 & ~n46681;
  assign n46683 = ~n46679 & ~n46682;
  assign n46684 = ~i_hbusreq1 & ~n46683;
  assign n46685 = ~n46676 & ~n46684;
  assign n46686 = controllable_hgrant1 & ~n46685;
  assign n46687 = i_hbusreq1 & ~n46064;
  assign n46688 = i_hbusreq2 & ~n46059;
  assign n46689 = i_hbusreq0 & ~n46052;
  assign n46690 = controllable_hmastlock & ~n46582;
  assign n46691 = ~n44281 & ~n46690;
  assign n46692 = controllable_locked & ~n46691;
  assign n46693 = ~n44283 & ~n46692;
  assign n46694 = i_hlock0 & ~n46693;
  assign n46695 = ~i_hlock0 & ~n46057;
  assign n46696 = ~n46694 & ~n46695;
  assign n46697 = ~i_hbusreq0 & ~n46696;
  assign n46698 = ~n46689 & ~n46697;
  assign n46699 = i_hlock2 & ~n46698;
  assign n46700 = i_hbusreq0 & ~n46057;
  assign n46701 = ~n46697 & ~n46700;
  assign n46702 = ~i_hlock2 & ~n46701;
  assign n46703 = ~n46699 & ~n46702;
  assign n46704 = ~i_hbusreq2 & ~n46703;
  assign n46705 = ~n46688 & ~n46704;
  assign n46706 = controllable_hgrant2 & ~n46705;
  assign n46707 = i_hlock0 & ~n14242;
  assign n46708 = ~n44269 & ~n46707;
  assign n46709 = ~i_hbusreq0 & ~n46708;
  assign n46710 = ~i_hbusreq0 & ~n46709;
  assign n46711 = ~i_hbusreq2 & ~n46710;
  assign n46712 = ~i_hbusreq2 & ~n46711;
  assign n46713 = ~controllable_hgrant2 & n46712;
  assign n46714 = ~n46706 & ~n46713;
  assign n46715 = n7733 & ~n46714;
  assign n46716 = ~n44277 & ~n46715;
  assign n46717 = n7928 & ~n46716;
  assign n46718 = ~n8265 & ~n46717;
  assign n46719 = ~i_hbusreq1 & ~n46718;
  assign n46720 = ~n46687 & ~n46719;
  assign n46721 = ~controllable_hgrant1 & ~n46720;
  assign n46722 = ~n46686 & ~n46721;
  assign n46723 = ~i_hbusreq3 & ~n46722;
  assign n46724 = ~n46675 & ~n46723;
  assign n46725 = ~controllable_hgrant3 & ~n46724;
  assign n46726 = ~n46674 & ~n46725;
  assign n46727 = i_hlock9 & ~n46726;
  assign n46728 = i_hbusreq3 & ~n46076;
  assign n46729 = ~n8365 & ~n21077;
  assign n46730 = ~n44317 & ~n46729;
  assign n46731 = i_hlock3 & ~n46730;
  assign n46732 = ~n8365 & ~n21087;
  assign n46733 = ~n44317 & ~n46732;
  assign n46734 = ~i_hlock3 & ~n46733;
  assign n46735 = ~n46731 & ~n46734;
  assign n46736 = ~i_hbusreq3 & ~n46735;
  assign n46737 = ~n46728 & ~n46736;
  assign n46738 = controllable_hgrant3 & ~n46737;
  assign n46739 = i_hbusreq3 & ~n46088;
  assign n46740 = i_hbusreq1 & ~n46084;
  assign n46741 = ~n8389 & ~n21073;
  assign n46742 = ~n44325 & ~n46741;
  assign n46743 = i_hlock1 & ~n46742;
  assign n46744 = ~n8389 & ~n21083;
  assign n46745 = ~n44325 & ~n46744;
  assign n46746 = ~i_hlock1 & ~n46745;
  assign n46747 = ~n46743 & ~n46746;
  assign n46748 = ~i_hbusreq1 & ~n46747;
  assign n46749 = ~n46740 & ~n46748;
  assign n46750 = controllable_hgrant1 & ~n46749;
  assign n46751 = i_hbusreq1 & ~n46086;
  assign n46752 = ~n8297 & ~n46717;
  assign n46753 = ~i_hbusreq1 & ~n46752;
  assign n46754 = ~n46751 & ~n46753;
  assign n46755 = ~controllable_hgrant1 & ~n46754;
  assign n46756 = ~n46750 & ~n46755;
  assign n46757 = ~i_hbusreq3 & ~n46756;
  assign n46758 = ~n46739 & ~n46757;
  assign n46759 = ~controllable_hgrant3 & ~n46758;
  assign n46760 = ~n46738 & ~n46759;
  assign n46761 = ~i_hlock9 & ~n46760;
  assign n46762 = ~n46727 & ~n46761;
  assign n46763 = ~i_hbusreq9 & ~n46762;
  assign n46764 = ~n46663 & ~n46763;
  assign n46765 = ~i_hbusreq4 & ~n46764;
  assign n46766 = ~n46662 & ~n46765;
  assign n46767 = ~controllable_hgrant4 & ~n46766;
  assign n46768 = ~n46661 & ~n46767;
  assign n46769 = ~i_hbusreq5 & ~n46768;
  assign n46770 = ~n46634 & ~n46769;
  assign n46771 = ~controllable_hgrant5 & ~n46770;
  assign n46772 = ~n46633 & ~n46771;
  assign n46773 = ~controllable_hmaster2 & ~n46772;
  assign n46774 = ~n46622 & ~n46773;
  assign n46775 = ~controllable_hmaster1 & ~n46774;
  assign n46776 = ~n46621 & ~n46775;
  assign n46777 = ~i_hbusreq6 & ~n46776;
  assign n46778 = ~n46524 & ~n46777;
  assign n46779 = ~controllable_hgrant6 & ~n46778;
  assign n46780 = ~n46523 & ~n46779;
  assign n46781 = controllable_hmaster0 & ~n46780;
  assign n46782 = i_hbusreq6 & ~n46110;
  assign n46783 = ~n8217 & ~n31243;
  assign n46784 = ~n44363 & ~n46783;
  assign n46785 = i_hlock6 & ~n46784;
  assign n46786 = ~n8217 & ~n31465;
  assign n46787 = ~n44363 & ~n46786;
  assign n46788 = ~i_hlock6 & ~n46787;
  assign n46789 = ~n46785 & ~n46788;
  assign n46790 = ~i_hbusreq6 & ~n46789;
  assign n46791 = ~n46782 & ~n46790;
  assign n46792 = controllable_hgrant6 & ~n46791;
  assign n46793 = i_hbusreq6 & ~n46160;
  assign n46794 = i_hbusreq5 & ~n46118;
  assign n46795 = ~n8378 & ~n31235;
  assign n46796 = ~n44371 & ~n46795;
  assign n46797 = i_hlock5 & ~n46796;
  assign n46798 = ~n8378 & ~n31457;
  assign n46799 = ~n44371 & ~n46798;
  assign n46800 = ~i_hlock5 & ~n46799;
  assign n46801 = ~n46797 & ~n46800;
  assign n46802 = ~i_hbusreq5 & ~n46801;
  assign n46803 = ~n46794 & ~n46802;
  assign n46804 = controllable_hgrant5 & ~n46803;
  assign n46805 = i_hbusreq5 & ~n46154;
  assign n46806 = i_hbusreq4 & ~n46126;
  assign n46807 = i_hbusreq9 & ~n46121;
  assign n46808 = ~n8426 & ~n21134;
  assign n46809 = ~n44380 & ~n46808;
  assign n46810 = ~i_hbusreq9 & ~n46809;
  assign n46811 = ~n46807 & ~n46810;
  assign n46812 = i_hlock4 & ~n46811;
  assign n46813 = i_hbusreq9 & ~n46124;
  assign n46814 = ~n8426 & ~n21146;
  assign n46815 = ~n44380 & ~n46814;
  assign n46816 = ~i_hbusreq9 & ~n46815;
  assign n46817 = ~n46813 & ~n46816;
  assign n46818 = ~i_hlock4 & ~n46817;
  assign n46819 = ~n46812 & ~n46818;
  assign n46820 = ~i_hbusreq4 & ~n46819;
  assign n46821 = ~n46806 & ~n46820;
  assign n46822 = controllable_hgrant4 & ~n46821;
  assign n46823 = i_hbusreq4 & ~n46152;
  assign n46824 = i_hbusreq9 & ~n46152;
  assign n46825 = i_hbusreq3 & ~n46134;
  assign n46826 = ~n8365 & ~n21130;
  assign n46827 = ~n44391 & ~n46826;
  assign n46828 = i_hlock3 & ~n46827;
  assign n46829 = ~n8365 & ~n21142;
  assign n46830 = ~n44391 & ~n46829;
  assign n46831 = ~i_hlock3 & ~n46830;
  assign n46832 = ~n46828 & ~n46831;
  assign n46833 = ~i_hbusreq3 & ~n46832;
  assign n46834 = ~n46825 & ~n46833;
  assign n46835 = controllable_hgrant3 & ~n46834;
  assign n46836 = i_hbusreq3 & ~n46150;
  assign n46837 = i_hbusreq1 & ~n46142;
  assign n46838 = ~n8389 & ~n21126;
  assign n46839 = ~n44399 & ~n46838;
  assign n46840 = i_hlock1 & ~n46839;
  assign n46841 = ~n8389 & ~n21138;
  assign n46842 = ~n44399 & ~n46841;
  assign n46843 = ~i_hlock1 & ~n46842;
  assign n46844 = ~n46840 & ~n46843;
  assign n46845 = ~i_hbusreq1 & ~n46844;
  assign n46846 = ~n46837 & ~n46845;
  assign n46847 = controllable_hgrant1 & ~n46846;
  assign n46848 = i_hbusreq1 & ~n46148;
  assign n46849 = ~n20882 & ~n46597;
  assign n46850 = n7733 & ~n46849;
  assign n46851 = ~n44407 & ~n46850;
  assign n46852 = n7928 & ~n46851;
  assign n46853 = ~n8265 & ~n46852;
  assign n46854 = ~i_hbusreq1 & ~n46853;
  assign n46855 = ~n46848 & ~n46854;
  assign n46856 = ~controllable_hgrant1 & ~n46855;
  assign n46857 = ~n46847 & ~n46856;
  assign n46858 = ~i_hbusreq3 & ~n46857;
  assign n46859 = ~n46836 & ~n46858;
  assign n46860 = ~controllable_hgrant3 & ~n46859;
  assign n46861 = ~n46835 & ~n46860;
  assign n46862 = ~i_hbusreq9 & ~n46861;
  assign n46863 = ~n46824 & ~n46862;
  assign n46864 = ~i_hbusreq4 & ~n46863;
  assign n46865 = ~n46823 & ~n46864;
  assign n46866 = ~controllable_hgrant4 & ~n46865;
  assign n46867 = ~n46822 & ~n46866;
  assign n46868 = ~i_hbusreq5 & ~n46867;
  assign n46869 = ~n46805 & ~n46868;
  assign n46870 = ~controllable_hgrant5 & ~n46869;
  assign n46871 = ~n46804 & ~n46870;
  assign n46872 = ~controllable_hmaster2 & ~n46871;
  assign n46873 = ~n46622 & ~n46872;
  assign n46874 = ~controllable_hmaster1 & ~n46873;
  assign n46875 = ~n46621 & ~n46874;
  assign n46876 = ~i_hbusreq6 & ~n46875;
  assign n46877 = ~n46793 & ~n46876;
  assign n46878 = ~controllable_hgrant6 & ~n46877;
  assign n46879 = ~n46792 & ~n46878;
  assign n46880 = ~controllable_hmaster0 & ~n46879;
  assign n46881 = ~n46781 & ~n46880;
  assign n46882 = i_hlock8 & ~n46881;
  assign n46883 = i_hbusreq6 & ~n46172;
  assign n46884 = ~n8217 & ~n31268;
  assign n46885 = ~n44443 & ~n46884;
  assign n46886 = i_hlock6 & ~n46885;
  assign n46887 = ~n8217 & ~n31490;
  assign n46888 = ~n44443 & ~n46887;
  assign n46889 = ~i_hlock6 & ~n46888;
  assign n46890 = ~n46886 & ~n46889;
  assign n46891 = ~i_hbusreq6 & ~n46890;
  assign n46892 = ~n46883 & ~n46891;
  assign n46893 = controllable_hgrant6 & ~n46892;
  assign n46894 = i_hbusreq6 & ~n46218;
  assign n46895 = i_hbusreq5 & ~n46180;
  assign n46896 = ~n8378 & ~n31260;
  assign n46897 = ~n44451 & ~n46896;
  assign n46898 = i_hlock5 & ~n46897;
  assign n46899 = ~n8378 & ~n31482;
  assign n46900 = ~n44451 & ~n46899;
  assign n46901 = ~i_hlock5 & ~n46900;
  assign n46902 = ~n46898 & ~n46901;
  assign n46903 = ~i_hbusreq5 & ~n46902;
  assign n46904 = ~n46895 & ~n46903;
  assign n46905 = controllable_hgrant5 & ~n46904;
  assign n46906 = i_hbusreq5 & ~n46212;
  assign n46907 = i_hbusreq4 & ~n46188;
  assign n46908 = i_hbusreq9 & ~n46183;
  assign n46909 = ~n8426 & ~n21215;
  assign n46910 = ~n44460 & ~n46909;
  assign n46911 = ~i_hbusreq9 & ~n46910;
  assign n46912 = ~n46908 & ~n46911;
  assign n46913 = i_hlock4 & ~n46912;
  assign n46914 = i_hbusreq9 & ~n46186;
  assign n46915 = ~n8426 & ~n21221;
  assign n46916 = ~n44460 & ~n46915;
  assign n46917 = ~i_hbusreq9 & ~n46916;
  assign n46918 = ~n46914 & ~n46917;
  assign n46919 = ~i_hlock4 & ~n46918;
  assign n46920 = ~n46913 & ~n46919;
  assign n46921 = ~i_hbusreq4 & ~n46920;
  assign n46922 = ~n46907 & ~n46921;
  assign n46923 = controllable_hgrant4 & ~n46922;
  assign n46924 = i_hbusreq4 & ~n46210;
  assign n46925 = i_hbusreq9 & ~n46210;
  assign n46926 = i_hbusreq3 & ~n46196;
  assign n46927 = ~n8365 & ~n21170;
  assign n46928 = ~n44471 & ~n46927;
  assign n46929 = i_hlock3 & ~n46928;
  assign n46930 = ~n8365 & ~n21185;
  assign n46931 = ~n44471 & ~n46930;
  assign n46932 = ~i_hlock3 & ~n46931;
  assign n46933 = ~n46929 & ~n46932;
  assign n46934 = ~i_hbusreq3 & ~n46933;
  assign n46935 = ~n46926 & ~n46934;
  assign n46936 = controllable_hgrant3 & ~n46935;
  assign n46937 = i_hbusreq3 & ~n46208;
  assign n46938 = i_hbusreq1 & ~n46204;
  assign n46939 = ~n8389 & ~n21166;
  assign n46940 = ~n44479 & ~n46939;
  assign n46941 = i_hlock1 & ~n46940;
  assign n46942 = ~n8389 & ~n21181;
  assign n46943 = ~n44479 & ~n46942;
  assign n46944 = ~i_hlock1 & ~n46943;
  assign n46945 = ~n46941 & ~n46944;
  assign n46946 = ~i_hbusreq1 & ~n46945;
  assign n46947 = ~n46938 & ~n46946;
  assign n46948 = controllable_hgrant1 & ~n46947;
  assign n46949 = i_hbusreq1 & ~n46206;
  assign n46950 = ~n8297 & ~n46852;
  assign n46951 = ~i_hbusreq1 & ~n46950;
  assign n46952 = ~n46949 & ~n46951;
  assign n46953 = ~controllable_hgrant1 & ~n46952;
  assign n46954 = ~n46948 & ~n46953;
  assign n46955 = ~i_hbusreq3 & ~n46954;
  assign n46956 = ~n46937 & ~n46955;
  assign n46957 = ~controllable_hgrant3 & ~n46956;
  assign n46958 = ~n46936 & ~n46957;
  assign n46959 = ~i_hbusreq9 & ~n46958;
  assign n46960 = ~n46925 & ~n46959;
  assign n46961 = ~i_hbusreq4 & ~n46960;
  assign n46962 = ~n46924 & ~n46961;
  assign n46963 = ~controllable_hgrant4 & ~n46962;
  assign n46964 = ~n46923 & ~n46963;
  assign n46965 = ~i_hbusreq5 & ~n46964;
  assign n46966 = ~n46906 & ~n46965;
  assign n46967 = ~controllable_hgrant5 & ~n46966;
  assign n46968 = ~n46905 & ~n46967;
  assign n46969 = ~controllable_hmaster2 & ~n46968;
  assign n46970 = ~n46622 & ~n46969;
  assign n46971 = ~controllable_hmaster1 & ~n46970;
  assign n46972 = ~n46621 & ~n46971;
  assign n46973 = ~i_hbusreq6 & ~n46972;
  assign n46974 = ~n46894 & ~n46973;
  assign n46975 = ~controllable_hgrant6 & ~n46974;
  assign n46976 = ~n46893 & ~n46975;
  assign n46977 = ~controllable_hmaster0 & ~n46976;
  assign n46978 = ~n46781 & ~n46977;
  assign n46979 = ~i_hlock8 & ~n46978;
  assign n46980 = ~n46882 & ~n46979;
  assign n46981 = ~i_hbusreq8 & ~n46980;
  assign n46982 = ~n46512 & ~n46981;
  assign n46983 = controllable_hmaster3 & ~n46982;
  assign n46984 = i_hbusreq8 & ~n46488;
  assign n46985 = i_hbusreq6 & ~n46232;
  assign n46986 = ~n8217 & ~n37509;
  assign n46987 = ~n44522 & ~n46986;
  assign n46988 = i_hlock6 & ~n46987;
  assign n46989 = ~n8217 & ~n37520;
  assign n46990 = ~n44522 & ~n46989;
  assign n46991 = ~i_hlock6 & ~n46990;
  assign n46992 = ~n46988 & ~n46991;
  assign n46993 = ~i_hbusreq6 & ~n46992;
  assign n46994 = ~n46985 & ~n46993;
  assign n46995 = controllable_hgrant6 & ~n46994;
  assign n46996 = i_hbusreq6 & ~n46331;
  assign n46997 = controllable_hmaster2 & ~n46871;
  assign n46998 = i_hbusreq5 & ~n46241;
  assign n46999 = ~n8378 & ~n31304;
  assign n47000 = ~n44531 & ~n46999;
  assign n47001 = i_hlock5 & ~n47000;
  assign n47002 = ~n8378 & ~n31526;
  assign n47003 = ~n44531 & ~n47002;
  assign n47004 = ~i_hlock5 & ~n47003;
  assign n47005 = ~n47001 & ~n47004;
  assign n47006 = ~i_hbusreq5 & ~n47005;
  assign n47007 = ~n46998 & ~n47006;
  assign n47008 = controllable_hgrant5 & ~n47007;
  assign n47009 = i_hbusreq5 & ~n46265;
  assign n47010 = i_hbusreq4 & ~n46249;
  assign n47011 = i_hbusreq9 & ~n46244;
  assign n47012 = ~n8426 & ~n21176;
  assign n47013 = ~n44540 & ~n47012;
  assign n47014 = ~i_hbusreq9 & ~n47013;
  assign n47015 = ~n47011 & ~n47014;
  assign n47016 = i_hlock4 & ~n47015;
  assign n47017 = i_hbusreq9 & ~n46247;
  assign n47018 = ~n8426 & ~n21191;
  assign n47019 = ~n44540 & ~n47018;
  assign n47020 = ~i_hbusreq9 & ~n47019;
  assign n47021 = ~n47017 & ~n47020;
  assign n47022 = ~i_hlock4 & ~n47021;
  assign n47023 = ~n47016 & ~n47022;
  assign n47024 = ~i_hbusreq4 & ~n47023;
  assign n47025 = ~n47010 & ~n47024;
  assign n47026 = controllable_hgrant4 & ~n47025;
  assign n47027 = i_hbusreq4 & ~n46263;
  assign n47028 = i_hbusreq9 & ~n46263;
  assign n47029 = i_hbusreq3 & ~n46257;
  assign n47030 = ~n8365 & ~n20959;
  assign n47031 = ~n44551 & ~n47030;
  assign n47032 = i_hlock3 & ~n47031;
  assign n47033 = ~n8365 & ~n20981;
  assign n47034 = ~n44555 & ~n47033;
  assign n47035 = ~i_hlock3 & ~n47034;
  assign n47036 = ~n47032 & ~n47035;
  assign n47037 = ~i_hbusreq3 & ~n47036;
  assign n47038 = ~n47029 & ~n47037;
  assign n47039 = controllable_hgrant3 & ~n47038;
  assign n47040 = i_hbusreq3 & ~n46261;
  assign n47041 = i_hlock3 & ~n46857;
  assign n47042 = ~i_hlock3 & ~n46954;
  assign n47043 = ~n47041 & ~n47042;
  assign n47044 = ~i_hbusreq3 & ~n47043;
  assign n47045 = ~n47040 & ~n47044;
  assign n47046 = ~controllable_hgrant3 & ~n47045;
  assign n47047 = ~n47039 & ~n47046;
  assign n47048 = ~i_hbusreq9 & ~n47047;
  assign n47049 = ~n47028 & ~n47048;
  assign n47050 = ~i_hbusreq4 & ~n47049;
  assign n47051 = ~n47027 & ~n47050;
  assign n47052 = ~controllable_hgrant4 & ~n47051;
  assign n47053 = ~n47026 & ~n47052;
  assign n47054 = ~i_hbusreq5 & ~n47053;
  assign n47055 = ~n47009 & ~n47054;
  assign n47056 = ~controllable_hgrant5 & ~n47055;
  assign n47057 = ~n47008 & ~n47056;
  assign n47058 = ~controllable_hmaster2 & ~n47057;
  assign n47059 = ~n46997 & ~n47058;
  assign n47060 = controllable_hmaster1 & ~n47059;
  assign n47061 = i_hbusreq5 & ~n46277;
  assign n47062 = ~n8378 & ~n31290;
  assign n47063 = ~n44585 & ~n47062;
  assign n47064 = i_hlock5 & ~n47063;
  assign n47065 = ~n8378 & ~n31512;
  assign n47066 = ~n44589 & ~n47065;
  assign n47067 = ~i_hlock5 & ~n47066;
  assign n47068 = ~n47064 & ~n47067;
  assign n47069 = ~i_hbusreq5 & ~n47068;
  assign n47070 = ~n47061 & ~n47069;
  assign n47071 = controllable_hgrant5 & ~n47070;
  assign n47072 = i_hbusreq5 & ~n46281;
  assign n47073 = i_hlock5 & ~n46867;
  assign n47074 = ~i_hlock5 & ~n46964;
  assign n47075 = ~n47073 & ~n47074;
  assign n47076 = ~i_hbusreq5 & ~n47075;
  assign n47077 = ~n47072 & ~n47076;
  assign n47078 = ~controllable_hgrant5 & ~n47077;
  assign n47079 = ~n47071 & ~n47078;
  assign n47080 = controllable_hmaster2 & ~n47079;
  assign n47081 = i_hbusreq5 & ~n46291;
  assign n47082 = ~n8378 & ~n31329;
  assign n47083 = ~n44607 & ~n47082;
  assign n47084 = i_hlock5 & ~n47083;
  assign n47085 = ~n8378 & ~n31551;
  assign n47086 = ~n44607 & ~n47085;
  assign n47087 = ~i_hlock5 & ~n47086;
  assign n47088 = ~n47084 & ~n47087;
  assign n47089 = ~i_hbusreq5 & ~n47088;
  assign n47090 = ~n47081 & ~n47089;
  assign n47091 = controllable_hgrant5 & ~n47090;
  assign n47092 = i_hbusreq5 & ~n46325;
  assign n47093 = i_hbusreq4 & ~n46299;
  assign n47094 = i_hbusreq9 & ~n46294;
  assign n47095 = ~n8426 & ~n21252;
  assign n47096 = ~n44616 & ~n47095;
  assign n47097 = ~i_hbusreq9 & ~n47096;
  assign n47098 = ~n47094 & ~n47097;
  assign n47099 = i_hlock4 & ~n47098;
  assign n47100 = i_hbusreq9 & ~n46297;
  assign n47101 = ~n8426 & ~n21266;
  assign n47102 = ~n44616 & ~n47101;
  assign n47103 = ~i_hbusreq9 & ~n47102;
  assign n47104 = ~n47100 & ~n47103;
  assign n47105 = ~i_hlock4 & ~n47104;
  assign n47106 = ~n47099 & ~n47105;
  assign n47107 = ~i_hbusreq4 & ~n47106;
  assign n47108 = ~n47093 & ~n47107;
  assign n47109 = controllable_hgrant4 & ~n47108;
  assign n47110 = i_hbusreq4 & ~n46323;
  assign n47111 = i_hbusreq9 & ~n46323;
  assign n47112 = i_hbusreq3 & ~n46307;
  assign n47113 = ~n8365 & ~n21248;
  assign n47114 = ~n44627 & ~n47113;
  assign n47115 = i_hlock3 & ~n47114;
  assign n47116 = ~n8365 & ~n21262;
  assign n47117 = ~n44627 & ~n47116;
  assign n47118 = ~i_hlock3 & ~n47117;
  assign n47119 = ~n47115 & ~n47118;
  assign n47120 = ~i_hbusreq3 & ~n47119;
  assign n47121 = ~n47112 & ~n47120;
  assign n47122 = controllable_hgrant3 & ~n47121;
  assign n47123 = i_hbusreq3 & ~n46321;
  assign n47124 = i_hbusreq1 & ~n46315;
  assign n47125 = ~n8389 & ~n20955;
  assign n47126 = ~n44635 & ~n47125;
  assign n47127 = i_hlock1 & ~n47126;
  assign n47128 = ~n8389 & ~n20977;
  assign n47129 = ~n44639 & ~n47128;
  assign n47130 = ~i_hlock1 & ~n47129;
  assign n47131 = ~n47127 & ~n47130;
  assign n47132 = ~i_hbusreq1 & ~n47131;
  assign n47133 = ~n47124 & ~n47132;
  assign n47134 = controllable_hgrant1 & ~n47133;
  assign n47135 = i_hbusreq1 & ~n46319;
  assign n47136 = i_hlock1 & ~n46853;
  assign n47137 = ~i_hlock1 & ~n46950;
  assign n47138 = ~n47136 & ~n47137;
  assign n47139 = ~i_hbusreq1 & ~n47138;
  assign n47140 = ~n47135 & ~n47139;
  assign n47141 = ~controllable_hgrant1 & ~n47140;
  assign n47142 = ~n47134 & ~n47141;
  assign n47143 = ~i_hbusreq3 & ~n47142;
  assign n47144 = ~n47123 & ~n47143;
  assign n47145 = ~controllable_hgrant3 & ~n47144;
  assign n47146 = ~n47122 & ~n47145;
  assign n47147 = ~i_hbusreq9 & ~n47146;
  assign n47148 = ~n47111 & ~n47147;
  assign n47149 = ~i_hbusreq4 & ~n47148;
  assign n47150 = ~n47110 & ~n47149;
  assign n47151 = ~controllable_hgrant4 & ~n47150;
  assign n47152 = ~n47109 & ~n47151;
  assign n47153 = ~i_hbusreq5 & ~n47152;
  assign n47154 = ~n47092 & ~n47153;
  assign n47155 = ~controllable_hgrant5 & ~n47154;
  assign n47156 = ~n47091 & ~n47155;
  assign n47157 = ~controllable_hmaster2 & ~n47156;
  assign n47158 = ~n47080 & ~n47157;
  assign n47159 = ~controllable_hmaster1 & ~n47158;
  assign n47160 = ~n47060 & ~n47159;
  assign n47161 = ~i_hbusreq6 & ~n47160;
  assign n47162 = ~n46996 & ~n47161;
  assign n47163 = ~controllable_hgrant6 & ~n47162;
  assign n47164 = ~n46995 & ~n47163;
  assign n47165 = controllable_hmaster0 & ~n47164;
  assign n47166 = i_hbusreq6 & ~n46347;
  assign n47167 = ~n31295 & ~n31358;
  assign n47168 = controllable_hmaster1 & ~n47167;
  assign n47169 = ~n31390 & ~n47168;
  assign n47170 = ~n8217 & ~n47169;
  assign n47171 = ~n44682 & ~n47170;
  assign n47172 = i_hlock6 & ~n47171;
  assign n47173 = ~n31517 & ~n31580;
  assign n47174 = controllable_hmaster1 & ~n47173;
  assign n47175 = ~n31612 & ~n47174;
  assign n47176 = ~n8217 & ~n47175;
  assign n47177 = ~n44692 & ~n47176;
  assign n47178 = ~i_hlock6 & ~n47177;
  assign n47179 = ~n47172 & ~n47178;
  assign n47180 = ~i_hbusreq6 & ~n47179;
  assign n47181 = ~n47166 & ~n47180;
  assign n47182 = controllable_hgrant6 & ~n47181;
  assign n47183 = i_hbusreq6 & ~n46484;
  assign n47184 = i_hbusreq5 & ~n46355;
  assign n47185 = ~n8378 & ~n31353;
  assign n47186 = ~n44705 & ~n47185;
  assign n47187 = i_hlock5 & ~n47186;
  assign n47188 = ~n8378 & ~n31575;
  assign n47189 = ~n44705 & ~n47188;
  assign n47190 = ~i_hlock5 & ~n47189;
  assign n47191 = ~n47187 & ~n47190;
  assign n47192 = ~i_hbusreq5 & ~n47191;
  assign n47193 = ~n47184 & ~n47192;
  assign n47194 = controllable_hgrant5 & ~n47193;
  assign n47195 = i_hbusreq5 & ~n46403;
  assign n47196 = i_hbusreq4 & ~n46363;
  assign n47197 = i_hbusreq9 & ~n46358;
  assign n47198 = ~n8426 & ~n21302;
  assign n47199 = ~n44714 & ~n47198;
  assign n47200 = ~i_hbusreq9 & ~n47199;
  assign n47201 = ~n47197 & ~n47200;
  assign n47202 = i_hlock4 & ~n47201;
  assign n47203 = i_hbusreq9 & ~n46361;
  assign n47204 = ~n8426 & ~n21314;
  assign n47205 = ~n44714 & ~n47204;
  assign n47206 = ~i_hbusreq9 & ~n47205;
  assign n47207 = ~n47203 & ~n47206;
  assign n47208 = ~i_hlock4 & ~n47207;
  assign n47209 = ~n47202 & ~n47208;
  assign n47210 = ~i_hbusreq4 & ~n47209;
  assign n47211 = ~n47196 & ~n47210;
  assign n47212 = controllable_hgrant4 & ~n47211;
  assign n47213 = i_hbusreq4 & ~n46401;
  assign n47214 = i_hbusreq9 & ~n46401;
  assign n47215 = i_hbusreq3 & ~n46371;
  assign n47216 = ~n8365 & ~n21298;
  assign n47217 = ~n44725 & ~n47216;
  assign n47218 = i_hlock3 & ~n47217;
  assign n47219 = ~n8365 & ~n21310;
  assign n47220 = ~n44725 & ~n47219;
  assign n47221 = ~i_hlock3 & ~n47220;
  assign n47222 = ~n47218 & ~n47221;
  assign n47223 = ~i_hbusreq3 & ~n47222;
  assign n47224 = ~n47215 & ~n47223;
  assign n47225 = controllable_hgrant3 & ~n47224;
  assign n47226 = i_hbusreq3 & ~n46399;
  assign n47227 = i_hbusreq1 & ~n46379;
  assign n47228 = ~n8389 & ~n21294;
  assign n47229 = ~n44733 & ~n47228;
  assign n47230 = i_hlock1 & ~n47229;
  assign n47231 = ~n8389 & ~n21306;
  assign n47232 = ~n44733 & ~n47231;
  assign n47233 = ~i_hlock1 & ~n47232;
  assign n47234 = ~n47230 & ~n47233;
  assign n47235 = ~i_hbusreq1 & ~n47234;
  assign n47236 = ~n47227 & ~n47235;
  assign n47237 = controllable_hgrant1 & ~n47236;
  assign n47238 = i_hbusreq1 & ~n46397;
  assign n47239 = i_hbusreq2 & ~n46391;
  assign n47240 = i_hbusreq0 & ~n46384;
  assign n47241 = ~controllable_hmastlock & ~n46582;
  assign n47242 = ~n39853 & ~n47241;
  assign n47243 = controllable_locked & ~n47242;
  assign n47244 = ~n44182 & ~n47243;
  assign n47245 = i_hlock0 & ~n47244;
  assign n47246 = ~i_hlock0 & ~n46389;
  assign n47247 = ~n47245 & ~n47246;
  assign n47248 = ~i_hbusreq0 & ~n47247;
  assign n47249 = ~n47240 & ~n47248;
  assign n47250 = i_hlock2 & ~n47249;
  assign n47251 = i_hbusreq0 & ~n46389;
  assign n47252 = ~n47248 & ~n47251;
  assign n47253 = ~i_hlock2 & ~n47252;
  assign n47254 = ~n47250 & ~n47253;
  assign n47255 = ~i_hbusreq2 & ~n47254;
  assign n47256 = ~n47239 & ~n47255;
  assign n47257 = controllable_hgrant2 & ~n47256;
  assign n47258 = ~n20882 & ~n47257;
  assign n47259 = n7733 & ~n47258;
  assign n47260 = ~n44752 & ~n47259;
  assign n47261 = n7928 & ~n47260;
  assign n47262 = ~n43545 & ~n47261;
  assign n47263 = ~i_hbusreq1 & ~n47262;
  assign n47264 = ~n47238 & ~n47263;
  assign n47265 = ~controllable_hgrant1 & ~n47264;
  assign n47266 = ~n47237 & ~n47265;
  assign n47267 = ~i_hbusreq3 & ~n47266;
  assign n47268 = ~n47226 & ~n47267;
  assign n47269 = ~controllable_hgrant3 & ~n47268;
  assign n47270 = ~n47225 & ~n47269;
  assign n47271 = ~i_hbusreq9 & ~n47270;
  assign n47272 = ~n47214 & ~n47271;
  assign n47273 = ~i_hbusreq4 & ~n47272;
  assign n47274 = ~n47213 & ~n47273;
  assign n47275 = ~controllable_hgrant4 & ~n47274;
  assign n47276 = ~n47212 & ~n47275;
  assign n47277 = ~i_hbusreq5 & ~n47276;
  assign n47278 = ~n47195 & ~n47277;
  assign n47279 = ~controllable_hgrant5 & ~n47278;
  assign n47280 = ~n47194 & ~n47279;
  assign n47281 = ~controllable_hmaster2 & ~n47280;
  assign n47282 = ~n46997 & ~n47281;
  assign n47283 = controllable_hmaster1 & ~n47282;
  assign n47284 = i_hbusreq5 & ~n46415;
  assign n47285 = ~n8378 & ~n31369;
  assign n47286 = ~n44780 & ~n47285;
  assign n47287 = i_hlock5 & ~n47286;
  assign n47288 = ~n8378 & ~n31591;
  assign n47289 = ~n44780 & ~n47288;
  assign n47290 = ~i_hlock5 & ~n47289;
  assign n47291 = ~n47287 & ~n47290;
  assign n47292 = ~i_hbusreq5 & ~n47291;
  assign n47293 = ~n47284 & ~n47292;
  assign n47294 = controllable_hgrant5 & ~n47293;
  assign n47295 = i_hbusreq5 & ~n46429;
  assign n47296 = i_hbusreq4 & ~n46423;
  assign n47297 = i_hbusreq9 & ~n46418;
  assign n47298 = ~n8426 & ~n20963;
  assign n47299 = ~n44789 & ~n47298;
  assign n47300 = ~i_hbusreq9 & ~n47299;
  assign n47301 = ~n47297 & ~n47300;
  assign n47302 = i_hlock4 & ~n47301;
  assign n47303 = i_hbusreq9 & ~n46421;
  assign n47304 = ~n8426 & ~n20985;
  assign n47305 = ~n44796 & ~n47304;
  assign n47306 = ~i_hbusreq9 & ~n47305;
  assign n47307 = ~n47303 & ~n47306;
  assign n47308 = ~i_hlock4 & ~n47307;
  assign n47309 = ~n47302 & ~n47308;
  assign n47310 = ~i_hbusreq4 & ~n47309;
  assign n47311 = ~n47296 & ~n47310;
  assign n47312 = controllable_hgrant4 & ~n47311;
  assign n47313 = i_hbusreq4 & ~n46427;
  assign n47314 = i_hlock4 & ~n46863;
  assign n47315 = ~i_hlock4 & ~n46960;
  assign n47316 = ~n47314 & ~n47315;
  assign n47317 = ~i_hbusreq4 & ~n47316;
  assign n47318 = ~n47313 & ~n47317;
  assign n47319 = ~controllable_hgrant4 & ~n47318;
  assign n47320 = ~n47312 & ~n47319;
  assign n47321 = ~i_hbusreq5 & ~n47320;
  assign n47322 = ~n47295 & ~n47321;
  assign n47323 = ~controllable_hgrant5 & ~n47322;
  assign n47324 = ~n47294 & ~n47323;
  assign n47325 = controllable_hmaster2 & ~n47324;
  assign n47326 = i_hbusreq5 & ~n46439;
  assign n47327 = ~n8378 & ~n31383;
  assign n47328 = ~n44820 & ~n47327;
  assign n47329 = i_hlock5 & ~n47328;
  assign n47330 = ~n8378 & ~n31605;
  assign n47331 = ~n44820 & ~n47330;
  assign n47332 = ~i_hlock5 & ~n47331;
  assign n47333 = ~n47329 & ~n47332;
  assign n47334 = ~i_hbusreq5 & ~n47333;
  assign n47335 = ~n47326 & ~n47334;
  assign n47336 = controllable_hgrant5 & ~n47335;
  assign n47337 = i_hbusreq5 & ~n46471;
  assign n47338 = i_hbusreq4 & ~n46447;
  assign n47339 = i_hbusreq9 & ~n46442;
  assign n47340 = ~n8426 & ~n21371;
  assign n47341 = ~n44829 & ~n47340;
  assign n47342 = ~i_hbusreq9 & ~n47341;
  assign n47343 = ~n47339 & ~n47342;
  assign n47344 = i_hlock4 & ~n47343;
  assign n47345 = i_hbusreq9 & ~n46445;
  assign n47346 = ~n8426 & ~n21391;
  assign n47347 = ~n44829 & ~n47346;
  assign n47348 = ~i_hbusreq9 & ~n47347;
  assign n47349 = ~n47345 & ~n47348;
  assign n47350 = ~i_hlock4 & ~n47349;
  assign n47351 = ~n47344 & ~n47350;
  assign n47352 = ~i_hbusreq4 & ~n47351;
  assign n47353 = ~n47338 & ~n47352;
  assign n47354 = controllable_hgrant4 & ~n47353;
  assign n47355 = i_hbusreq4 & ~n46469;
  assign n47356 = i_hbusreq9 & ~n46469;
  assign n47357 = i_hbusreq3 & ~n46455;
  assign n47358 = ~n8365 & ~n21367;
  assign n47359 = ~n44840 & ~n47358;
  assign n47360 = i_hlock3 & ~n47359;
  assign n47361 = ~n8365 & ~n21387;
  assign n47362 = ~n44840 & ~n47361;
  assign n47363 = ~i_hlock3 & ~n47362;
  assign n47364 = ~n47360 & ~n47363;
  assign n47365 = ~i_hbusreq3 & ~n47364;
  assign n47366 = ~n47357 & ~n47365;
  assign n47367 = controllable_hgrant3 & ~n47366;
  assign n47368 = i_hbusreq3 & ~n46467;
  assign n47369 = i_hbusreq1 & ~n46463;
  assign n47370 = ~n8389 & ~n21363;
  assign n47371 = ~n44848 & ~n47370;
  assign n47372 = i_hlock1 & ~n47371;
  assign n47373 = ~n8389 & ~n21383;
  assign n47374 = ~n44848 & ~n47373;
  assign n47375 = ~i_hlock1 & ~n47374;
  assign n47376 = ~n47372 & ~n47375;
  assign n47377 = ~i_hbusreq1 & ~n47376;
  assign n47378 = ~n47369 & ~n47377;
  assign n47379 = controllable_hgrant1 & ~n47378;
  assign n47380 = i_hbusreq1 & ~n46465;
  assign n47381 = ~n46054 & ~n47241;
  assign n47382 = controllable_locked & ~n47381;
  assign n47383 = ~n44857 & ~n47382;
  assign n47384 = i_hlock0 & ~n47383;
  assign n47385 = ~n46586 & ~n47384;
  assign n47386 = ~i_hbusreq0 & ~n47385;
  assign n47387 = ~n46581 & ~n47386;
  assign n47388 = i_hlock2 & ~n47387;
  assign n47389 = ~n46591 & ~n47386;
  assign n47390 = ~i_hlock2 & ~n47389;
  assign n47391 = ~n47388 & ~n47390;
  assign n47392 = ~i_hbusreq2 & ~n47391;
  assign n47393 = ~n46580 & ~n47392;
  assign n47394 = controllable_hgrant2 & ~n47393;
  assign n47395 = ~n21358 & ~n47394;
  assign n47396 = n7733 & ~n47395;
  assign n47397 = ~n44867 & ~n47396;
  assign n47398 = n7928 & ~n47397;
  assign n47399 = ~n8440 & ~n47398;
  assign n47400 = ~i_hbusreq1 & ~n47399;
  assign n47401 = ~n47380 & ~n47400;
  assign n47402 = ~controllable_hgrant1 & ~n47401;
  assign n47403 = ~n47379 & ~n47402;
  assign n47404 = ~i_hbusreq3 & ~n47403;
  assign n47405 = ~n47368 & ~n47404;
  assign n47406 = ~controllable_hgrant3 & ~n47405;
  assign n47407 = ~n47367 & ~n47406;
  assign n47408 = ~i_hbusreq9 & ~n47407;
  assign n47409 = ~n47356 & ~n47408;
  assign n47410 = ~i_hbusreq4 & ~n47409;
  assign n47411 = ~n47355 & ~n47410;
  assign n47412 = ~controllable_hgrant4 & ~n47411;
  assign n47413 = ~n47354 & ~n47412;
  assign n47414 = ~i_hbusreq5 & ~n47413;
  assign n47415 = ~n47337 & ~n47414;
  assign n47416 = ~controllable_hgrant5 & ~n47415;
  assign n47417 = ~n47336 & ~n47416;
  assign n47418 = ~controllable_hmaster2 & ~n47417;
  assign n47419 = ~n47325 & ~n47418;
  assign n47420 = ~controllable_hmaster1 & ~n47419;
  assign n47421 = ~n47283 & ~n47420;
  assign n47422 = i_hlock6 & ~n47421;
  assign n47423 = controllable_hmaster2 & ~n46968;
  assign n47424 = ~n47281 & ~n47423;
  assign n47425 = controllable_hmaster1 & ~n47424;
  assign n47426 = ~n47420 & ~n47425;
  assign n47427 = ~i_hlock6 & ~n47426;
  assign n47428 = ~n47422 & ~n47427;
  assign n47429 = ~i_hbusreq6 & ~n47428;
  assign n47430 = ~n47183 & ~n47429;
  assign n47431 = ~controllable_hgrant6 & ~n47430;
  assign n47432 = ~n47182 & ~n47431;
  assign n47433 = ~controllable_hmaster0 & ~n47432;
  assign n47434 = ~n47165 & ~n47433;
  assign n47435 = ~i_hbusreq8 & ~n47434;
  assign n47436 = ~n46984 & ~n47435;
  assign n47437 = ~controllable_hmaster3 & ~n47436;
  assign n47438 = ~n46983 & ~n47437;
  assign n47439 = i_hlock7 & ~n47438;
  assign n47440 = i_hbusreq8 & ~n46506;
  assign n47441 = i_hbusreq6 & ~n46498;
  assign n47442 = ~n8217 & ~n37538;
  assign n47443 = ~n44915 & ~n47442;
  assign n47444 = i_hlock6 & ~n47443;
  assign n47445 = ~n8217 & ~n37549;
  assign n47446 = ~n44915 & ~n47445;
  assign n47447 = ~i_hlock6 & ~n47446;
  assign n47448 = ~n47444 & ~n47447;
  assign n47449 = ~i_hbusreq6 & ~n47448;
  assign n47450 = ~n47441 & ~n47449;
  assign n47451 = controllable_hgrant6 & ~n47450;
  assign n47452 = i_hbusreq6 & ~n46502;
  assign n47453 = ~n47058 & ~n47423;
  assign n47454 = controllable_hmaster1 & ~n47453;
  assign n47455 = ~n47159 & ~n47454;
  assign n47456 = ~i_hbusreq6 & ~n47455;
  assign n47457 = ~n47452 & ~n47456;
  assign n47458 = ~controllable_hgrant6 & ~n47457;
  assign n47459 = ~n47451 & ~n47458;
  assign n47460 = controllable_hmaster0 & ~n47459;
  assign n47461 = ~n47433 & ~n47460;
  assign n47462 = ~i_hbusreq8 & ~n47461;
  assign n47463 = ~n47440 & ~n47462;
  assign n47464 = ~controllable_hmaster3 & ~n47463;
  assign n47465 = ~n46983 & ~n47464;
  assign n47466 = ~i_hlock7 & ~n47465;
  assign n47467 = ~n47439 & ~n47466;
  assign n47468 = ~i_hbusreq7 & ~n47467;
  assign n47469 = ~n46511 & ~n47468;
  assign n47470 = n7924 & ~n47469;
  assign n47471 = ~n43739 & ~n47470;
  assign n47472 = ~n8214 & ~n47471;
  assign n47473 = ~n8217 & ~n31647;
  assign n47474 = ~n41555 & ~n47473;
  assign n47475 = i_hlock6 & ~n47474;
  assign n47476 = ~n8217 & ~n31680;
  assign n47477 = ~n41555 & ~n47476;
  assign n47478 = ~i_hlock6 & ~n47477;
  assign n47479 = ~n47475 & ~n47478;
  assign n47480 = controllable_hgrant6 & ~n47479;
  assign n47481 = ~n8378 & ~n31641;
  assign n47482 = ~n41580 & ~n47481;
  assign n47483 = i_hlock5 & ~n47482;
  assign n47484 = ~n8378 & ~n31674;
  assign n47485 = ~n41580 & ~n47484;
  assign n47486 = ~i_hlock5 & ~n47485;
  assign n47487 = ~n47483 & ~n47486;
  assign n47488 = controllable_hgrant5 & ~n47487;
  assign n47489 = i_hlock9 & ~n46121;
  assign n47490 = ~i_hlock9 & ~n46183;
  assign n47491 = ~n47489 & ~n47490;
  assign n47492 = i_hlock4 & ~n47491;
  assign n47493 = i_hlock9 & ~n46124;
  assign n47494 = ~i_hlock9 & ~n46186;
  assign n47495 = ~n47493 & ~n47494;
  assign n47496 = ~i_hlock4 & ~n47495;
  assign n47497 = ~n47492 & ~n47496;
  assign n47498 = controllable_hgrant4 & ~n47497;
  assign n47499 = i_hlock9 & ~n46152;
  assign n47500 = ~i_hlock9 & ~n46210;
  assign n47501 = ~n47499 & ~n47500;
  assign n47502 = ~controllable_hgrant4 & ~n47501;
  assign n47503 = ~n47498 & ~n47502;
  assign n47504 = ~controllable_hgrant5 & ~n47503;
  assign n47505 = ~n47488 & ~n47504;
  assign n47506 = ~controllable_hmaster2 & ~n47505;
  assign n47507 = ~n46004 & ~n47506;
  assign n47508 = ~controllable_hmaster1 & ~n47507;
  assign n47509 = ~n46003 & ~n47508;
  assign n47510 = ~controllable_hgrant6 & ~n47509;
  assign n47511 = ~n47480 & ~n47510;
  assign n47512 = controllable_hmaster0 & ~n47511;
  assign n47513 = ~n8217 & ~n31653;
  assign n47514 = ~n42153 & ~n47513;
  assign n47515 = i_hlock6 & ~n47514;
  assign n47516 = ~n8217 & ~n31686;
  assign n47517 = ~n42153 & ~n47516;
  assign n47518 = ~i_hlock6 & ~n47517;
  assign n47519 = ~n47515 & ~n47518;
  assign n47520 = controllable_hgrant6 & ~n47519;
  assign n47521 = ~n8378 & ~n30256;
  assign n47522 = ~n42157 & ~n47521;
  assign n47523 = i_hlock5 & ~n47522;
  assign n47524 = ~n8378 & ~n30359;
  assign n47525 = ~n42157 & ~n47524;
  assign n47526 = ~i_hlock5 & ~n47525;
  assign n47527 = ~n47523 & ~n47526;
  assign n47528 = controllable_hgrant5 & ~n47527;
  assign n47529 = i_hlock4 & ~n46014;
  assign n47530 = ~i_hlock4 & ~n46022;
  assign n47531 = ~n47529 & ~n47530;
  assign n47532 = controllable_hgrant4 & ~n47531;
  assign n47533 = ~controllable_hgrant4 & ~n46068;
  assign n47534 = ~n47532 & ~n47533;
  assign n47535 = ~controllable_hgrant5 & ~n47534;
  assign n47536 = ~n47528 & ~n47535;
  assign n47537 = ~controllable_hmaster2 & ~n47536;
  assign n47538 = ~n46004 & ~n47537;
  assign n47539 = ~controllable_hmaster1 & ~n47538;
  assign n47540 = ~n46003 & ~n47539;
  assign n47541 = ~controllable_hgrant6 & ~n47540;
  assign n47542 = ~n47520 & ~n47541;
  assign n47543 = ~controllable_hmaster0 & ~n47542;
  assign n47544 = ~n47512 & ~n47543;
  assign n47545 = i_hlock8 & ~n47544;
  assign n47546 = ~n8217 & ~n31661;
  assign n47547 = ~n42175 & ~n47546;
  assign n47548 = i_hlock6 & ~n47547;
  assign n47549 = ~n8217 & ~n31694;
  assign n47550 = ~n42175 & ~n47549;
  assign n47551 = ~i_hlock6 & ~n47550;
  assign n47552 = ~n47548 & ~n47551;
  assign n47553 = controllable_hgrant6 & ~n47552;
  assign n47554 = ~n8378 & ~n30269;
  assign n47555 = ~n42179 & ~n47554;
  assign n47556 = i_hlock5 & ~n47555;
  assign n47557 = ~n8378 & ~n30372;
  assign n47558 = ~n42179 & ~n47557;
  assign n47559 = ~i_hlock5 & ~n47558;
  assign n47560 = ~n47556 & ~n47559;
  assign n47561 = controllable_hgrant5 & ~n47560;
  assign n47562 = i_hlock4 & ~n46017;
  assign n47563 = ~i_hlock4 & ~n46025;
  assign n47564 = ~n47562 & ~n47563;
  assign n47565 = controllable_hgrant4 & ~n47564;
  assign n47566 = ~controllable_hgrant4 & ~n46090;
  assign n47567 = ~n47565 & ~n47566;
  assign n47568 = ~controllable_hgrant5 & ~n47567;
  assign n47569 = ~n47561 & ~n47568;
  assign n47570 = ~controllable_hmaster2 & ~n47569;
  assign n47571 = ~n46004 & ~n47570;
  assign n47572 = ~controllable_hmaster1 & ~n47571;
  assign n47573 = ~n46003 & ~n47572;
  assign n47574 = ~controllable_hgrant6 & ~n47573;
  assign n47575 = ~n47553 & ~n47574;
  assign n47576 = ~controllable_hmaster0 & ~n47575;
  assign n47577 = ~n47512 & ~n47576;
  assign n47578 = ~i_hlock8 & ~n47577;
  assign n47579 = ~n47545 & ~n47578;
  assign n47580 = controllable_hmaster3 & ~n47579;
  assign n47581 = ~n46489 & ~n47580;
  assign n47582 = i_hlock7 & ~n47581;
  assign n47583 = ~n46507 & ~n47580;
  assign n47584 = ~i_hlock7 & ~n47583;
  assign n47585 = ~n47582 & ~n47584;
  assign n47586 = i_hbusreq7 & ~n47585;
  assign n47587 = i_hbusreq8 & ~n47579;
  assign n47588 = i_hbusreq6 & ~n47479;
  assign n47589 = ~n8217 & ~n31726;
  assign n47590 = ~n45169 & ~n47589;
  assign n47591 = i_hlock6 & ~n47590;
  assign n47592 = ~n8217 & ~n31802;
  assign n47593 = ~n45169 & ~n47592;
  assign n47594 = ~i_hlock6 & ~n47593;
  assign n47595 = ~n47591 & ~n47594;
  assign n47596 = ~i_hbusreq6 & ~n47595;
  assign n47597 = ~n47588 & ~n47596;
  assign n47598 = controllable_hgrant6 & ~n47597;
  assign n47599 = i_hbusreq6 & ~n47509;
  assign n47600 = i_hbusreq5 & ~n47487;
  assign n47601 = ~n8378 & ~n31718;
  assign n47602 = ~n45177 & ~n47601;
  assign n47603 = i_hlock5 & ~n47602;
  assign n47604 = ~n8378 & ~n31794;
  assign n47605 = ~n45177 & ~n47604;
  assign n47606 = ~i_hlock5 & ~n47605;
  assign n47607 = ~n47603 & ~n47606;
  assign n47608 = ~i_hbusreq5 & ~n47607;
  assign n47609 = ~n47600 & ~n47608;
  assign n47610 = controllable_hgrant5 & ~n47609;
  assign n47611 = i_hbusreq5 & ~n47503;
  assign n47612 = i_hbusreq4 & ~n47497;
  assign n47613 = i_hbusreq9 & ~n47491;
  assign n47614 = i_hlock9 & ~n46809;
  assign n47615 = ~i_hlock9 & ~n46910;
  assign n47616 = ~n47614 & ~n47615;
  assign n47617 = ~i_hbusreq9 & ~n47616;
  assign n47618 = ~n47613 & ~n47617;
  assign n47619 = i_hlock4 & ~n47618;
  assign n47620 = i_hbusreq9 & ~n47495;
  assign n47621 = i_hlock9 & ~n46815;
  assign n47622 = ~i_hlock9 & ~n46916;
  assign n47623 = ~n47621 & ~n47622;
  assign n47624 = ~i_hbusreq9 & ~n47623;
  assign n47625 = ~n47620 & ~n47624;
  assign n47626 = ~i_hlock4 & ~n47625;
  assign n47627 = ~n47619 & ~n47626;
  assign n47628 = ~i_hbusreq4 & ~n47627;
  assign n47629 = ~n47612 & ~n47628;
  assign n47630 = controllable_hgrant4 & ~n47629;
  assign n47631 = i_hbusreq4 & ~n47501;
  assign n47632 = i_hbusreq9 & ~n47501;
  assign n47633 = i_hlock9 & ~n46861;
  assign n47634 = ~i_hlock9 & ~n46958;
  assign n47635 = ~n47633 & ~n47634;
  assign n47636 = ~i_hbusreq9 & ~n47635;
  assign n47637 = ~n47632 & ~n47636;
  assign n47638 = ~i_hbusreq4 & ~n47637;
  assign n47639 = ~n47631 & ~n47638;
  assign n47640 = ~controllable_hgrant4 & ~n47639;
  assign n47641 = ~n47630 & ~n47640;
  assign n47642 = ~i_hbusreq5 & ~n47641;
  assign n47643 = ~n47611 & ~n47642;
  assign n47644 = ~controllable_hgrant5 & ~n47643;
  assign n47645 = ~n47610 & ~n47644;
  assign n47646 = ~controllable_hmaster2 & ~n47645;
  assign n47647 = ~n46622 & ~n47646;
  assign n47648 = ~controllable_hmaster1 & ~n47647;
  assign n47649 = ~n46621 & ~n47648;
  assign n47650 = ~i_hbusreq6 & ~n47649;
  assign n47651 = ~n47599 & ~n47650;
  assign n47652 = ~controllable_hgrant6 & ~n47651;
  assign n47653 = ~n47598 & ~n47652;
  assign n47654 = controllable_hmaster0 & ~n47653;
  assign n47655 = i_hbusreq6 & ~n47519;
  assign n47656 = ~n8217 & ~n31746;
  assign n47657 = ~n45219 & ~n47656;
  assign n47658 = i_hlock6 & ~n47657;
  assign n47659 = ~n8217 & ~n31822;
  assign n47660 = ~n45219 & ~n47659;
  assign n47661 = ~i_hlock6 & ~n47660;
  assign n47662 = ~n47658 & ~n47661;
  assign n47663 = ~i_hbusreq6 & ~n47662;
  assign n47664 = ~n47655 & ~n47663;
  assign n47665 = controllable_hgrant6 & ~n47664;
  assign n47666 = i_hbusreq6 & ~n47540;
  assign n47667 = i_hbusreq5 & ~n47527;
  assign n47668 = ~n8378 & ~n31738;
  assign n47669 = ~n45227 & ~n47668;
  assign n47670 = i_hlock5 & ~n47669;
  assign n47671 = ~n8378 & ~n31814;
  assign n47672 = ~n45227 & ~n47671;
  assign n47673 = ~i_hlock5 & ~n47672;
  assign n47674 = ~n47670 & ~n47673;
  assign n47675 = ~i_hbusreq5 & ~n47674;
  assign n47676 = ~n47667 & ~n47675;
  assign n47677 = controllable_hgrant5 & ~n47676;
  assign n47678 = i_hbusreq5 & ~n47534;
  assign n47679 = i_hbusreq4 & ~n47531;
  assign n47680 = i_hbusreq9 & ~n46014;
  assign n47681 = ~i_hbusreq9 & ~n46638;
  assign n47682 = ~n47680 & ~n47681;
  assign n47683 = i_hlock4 & ~n47682;
  assign n47684 = i_hbusreq9 & ~n46022;
  assign n47685 = ~i_hbusreq9 & ~n46649;
  assign n47686 = ~n47684 & ~n47685;
  assign n47687 = ~i_hlock4 & ~n47686;
  assign n47688 = ~n47683 & ~n47687;
  assign n47689 = ~i_hbusreq4 & ~n47688;
  assign n47690 = ~n47679 & ~n47689;
  assign n47691 = controllable_hgrant4 & ~n47690;
  assign n47692 = i_hbusreq4 & ~n46068;
  assign n47693 = i_hbusreq9 & ~n46068;
  assign n47694 = ~i_hbusreq9 & ~n46726;
  assign n47695 = ~n47693 & ~n47694;
  assign n47696 = ~i_hbusreq4 & ~n47695;
  assign n47697 = ~n47692 & ~n47696;
  assign n47698 = ~controllable_hgrant4 & ~n47697;
  assign n47699 = ~n47691 & ~n47698;
  assign n47700 = ~i_hbusreq5 & ~n47699;
  assign n47701 = ~n47678 & ~n47700;
  assign n47702 = ~controllable_hgrant5 & ~n47701;
  assign n47703 = ~n47677 & ~n47702;
  assign n47704 = ~controllable_hmaster2 & ~n47703;
  assign n47705 = ~n46622 & ~n47704;
  assign n47706 = ~controllable_hmaster1 & ~n47705;
  assign n47707 = ~n46621 & ~n47706;
  assign n47708 = ~i_hbusreq6 & ~n47707;
  assign n47709 = ~n47666 & ~n47708;
  assign n47710 = ~controllable_hgrant6 & ~n47709;
  assign n47711 = ~n47665 & ~n47710;
  assign n47712 = ~controllable_hmaster0 & ~n47711;
  assign n47713 = ~n47654 & ~n47712;
  assign n47714 = i_hlock8 & ~n47713;
  assign n47715 = i_hbusreq6 & ~n47552;
  assign n47716 = ~n8217 & ~n31768;
  assign n47717 = ~n45265 & ~n47716;
  assign n47718 = i_hlock6 & ~n47717;
  assign n47719 = ~n8217 & ~n31844;
  assign n47720 = ~n45265 & ~n47719;
  assign n47721 = ~i_hlock6 & ~n47720;
  assign n47722 = ~n47718 & ~n47721;
  assign n47723 = ~i_hbusreq6 & ~n47722;
  assign n47724 = ~n47715 & ~n47723;
  assign n47725 = controllable_hgrant6 & ~n47724;
  assign n47726 = i_hbusreq6 & ~n47573;
  assign n47727 = i_hbusreq5 & ~n47560;
  assign n47728 = ~n8378 & ~n31760;
  assign n47729 = ~n45273 & ~n47728;
  assign n47730 = i_hlock5 & ~n47729;
  assign n47731 = ~n8378 & ~n31836;
  assign n47732 = ~n45273 & ~n47731;
  assign n47733 = ~i_hlock5 & ~n47732;
  assign n47734 = ~n47730 & ~n47733;
  assign n47735 = ~i_hbusreq5 & ~n47734;
  assign n47736 = ~n47727 & ~n47735;
  assign n47737 = controllable_hgrant5 & ~n47736;
  assign n47738 = i_hbusreq5 & ~n47567;
  assign n47739 = i_hbusreq4 & ~n47564;
  assign n47740 = i_hbusreq9 & ~n46017;
  assign n47741 = ~i_hbusreq9 & ~n46641;
  assign n47742 = ~n47740 & ~n47741;
  assign n47743 = i_hlock4 & ~n47742;
  assign n47744 = i_hbusreq9 & ~n46025;
  assign n47745 = ~i_hbusreq9 & ~n46652;
  assign n47746 = ~n47744 & ~n47745;
  assign n47747 = ~i_hlock4 & ~n47746;
  assign n47748 = ~n47743 & ~n47747;
  assign n47749 = ~i_hbusreq4 & ~n47748;
  assign n47750 = ~n47739 & ~n47749;
  assign n47751 = controllable_hgrant4 & ~n47750;
  assign n47752 = i_hbusreq4 & ~n46090;
  assign n47753 = i_hbusreq9 & ~n46090;
  assign n47754 = ~i_hbusreq9 & ~n46760;
  assign n47755 = ~n47753 & ~n47754;
  assign n47756 = ~i_hbusreq4 & ~n47755;
  assign n47757 = ~n47752 & ~n47756;
  assign n47758 = ~controllable_hgrant4 & ~n47757;
  assign n47759 = ~n47751 & ~n47758;
  assign n47760 = ~i_hbusreq5 & ~n47759;
  assign n47761 = ~n47738 & ~n47760;
  assign n47762 = ~controllable_hgrant5 & ~n47761;
  assign n47763 = ~n47737 & ~n47762;
  assign n47764 = ~controllable_hmaster2 & ~n47763;
  assign n47765 = ~n46622 & ~n47764;
  assign n47766 = ~controllable_hmaster1 & ~n47765;
  assign n47767 = ~n46621 & ~n47766;
  assign n47768 = ~i_hbusreq6 & ~n47767;
  assign n47769 = ~n47726 & ~n47768;
  assign n47770 = ~controllable_hgrant6 & ~n47769;
  assign n47771 = ~n47725 & ~n47770;
  assign n47772 = ~controllable_hmaster0 & ~n47771;
  assign n47773 = ~n47654 & ~n47772;
  assign n47774 = ~i_hlock8 & ~n47773;
  assign n47775 = ~n47714 & ~n47774;
  assign n47776 = ~i_hbusreq8 & ~n47775;
  assign n47777 = ~n47587 & ~n47776;
  assign n47778 = controllable_hmaster3 & ~n47777;
  assign n47779 = ~n47437 & ~n47778;
  assign n47780 = i_hlock7 & ~n47779;
  assign n47781 = ~n47464 & ~n47778;
  assign n47782 = ~i_hlock7 & ~n47781;
  assign n47783 = ~n47780 & ~n47782;
  assign n47784 = ~i_hbusreq7 & ~n47783;
  assign n47785 = ~n47586 & ~n47784;
  assign n47786 = n7924 & ~n47785;
  assign n47787 = ~n45094 & ~n47786;
  assign n47788 = n8214 & ~n47787;
  assign n47789 = ~n47472 & ~n47788;
  assign n47790 = ~n8202 & ~n47789;
  assign n47791 = ~n46163 & ~n47512;
  assign n47792 = i_hlock8 & ~n47791;
  assign n47793 = ~n46221 & ~n47512;
  assign n47794 = ~i_hlock8 & ~n47793;
  assign n47795 = ~n47792 & ~n47794;
  assign n47796 = controllable_hmaster3 & ~n47795;
  assign n47797 = ~n8217 & ~n37579;
  assign n47798 = ~n43905 & ~n47797;
  assign n47799 = i_hlock6 & ~n47798;
  assign n47800 = ~n8217 & ~n37587;
  assign n47801 = ~n43905 & ~n47800;
  assign n47802 = ~i_hlock6 & ~n47801;
  assign n47803 = ~n47799 & ~n47802;
  assign n47804 = controllable_hgrant6 & ~n47803;
  assign n47805 = controllable_hmaster2 & ~n47536;
  assign n47806 = ~n46268 & ~n47805;
  assign n47807 = controllable_hmaster1 & ~n47806;
  assign n47808 = ~n46330 & ~n47807;
  assign n47809 = ~controllable_hgrant6 & ~n47808;
  assign n47810 = ~n47804 & ~n47809;
  assign n47811 = controllable_hmaster0 & ~n47810;
  assign n47812 = ~n46487 & ~n47811;
  assign n47813 = ~controllable_hmaster3 & ~n47812;
  assign n47814 = ~n47796 & ~n47813;
  assign n47815 = i_hlock7 & ~n47814;
  assign n47816 = ~n8217 & ~n37599;
  assign n47817 = ~n44119 & ~n47816;
  assign n47818 = i_hlock6 & ~n47817;
  assign n47819 = ~n8217 & ~n37607;
  assign n47820 = ~n44119 & ~n47819;
  assign n47821 = ~i_hlock6 & ~n47820;
  assign n47822 = ~n47818 & ~n47821;
  assign n47823 = controllable_hgrant6 & ~n47822;
  assign n47824 = controllable_hmaster2 & ~n47569;
  assign n47825 = ~n46268 & ~n47824;
  assign n47826 = controllable_hmaster1 & ~n47825;
  assign n47827 = ~n46330 & ~n47826;
  assign n47828 = ~controllable_hgrant6 & ~n47827;
  assign n47829 = ~n47823 & ~n47828;
  assign n47830 = controllable_hmaster0 & ~n47829;
  assign n47831 = ~n46487 & ~n47830;
  assign n47832 = ~controllable_hmaster3 & ~n47831;
  assign n47833 = ~n47796 & ~n47832;
  assign n47834 = ~i_hlock7 & ~n47833;
  assign n47835 = ~n47815 & ~n47834;
  assign n47836 = i_hbusreq7 & ~n47835;
  assign n47837 = i_hbusreq8 & ~n47795;
  assign n47838 = ~n46880 & ~n47654;
  assign n47839 = i_hlock8 & ~n47838;
  assign n47840 = ~n46977 & ~n47654;
  assign n47841 = ~i_hlock8 & ~n47840;
  assign n47842 = ~n47839 & ~n47841;
  assign n47843 = ~i_hbusreq8 & ~n47842;
  assign n47844 = ~n47837 & ~n47843;
  assign n47845 = controllable_hmaster3 & ~n47844;
  assign n47846 = i_hbusreq8 & ~n47812;
  assign n47847 = i_hbusreq6 & ~n47803;
  assign n47848 = ~n8217 & ~n37632;
  assign n47849 = ~n45466 & ~n47848;
  assign n47850 = i_hlock6 & ~n47849;
  assign n47851 = ~n8217 & ~n37643;
  assign n47852 = ~n45466 & ~n47851;
  assign n47853 = ~i_hlock6 & ~n47852;
  assign n47854 = ~n47850 & ~n47853;
  assign n47855 = ~i_hbusreq6 & ~n47854;
  assign n47856 = ~n47847 & ~n47855;
  assign n47857 = controllable_hgrant6 & ~n47856;
  assign n47858 = i_hbusreq6 & ~n47808;
  assign n47859 = controllable_hmaster2 & ~n47703;
  assign n47860 = ~n47058 & ~n47859;
  assign n47861 = controllable_hmaster1 & ~n47860;
  assign n47862 = ~n47159 & ~n47861;
  assign n47863 = ~i_hbusreq6 & ~n47862;
  assign n47864 = ~n47858 & ~n47863;
  assign n47865 = ~controllable_hgrant6 & ~n47864;
  assign n47866 = ~n47857 & ~n47865;
  assign n47867 = controllable_hmaster0 & ~n47866;
  assign n47868 = ~n47433 & ~n47867;
  assign n47869 = ~i_hbusreq8 & ~n47868;
  assign n47870 = ~n47846 & ~n47869;
  assign n47871 = ~controllable_hmaster3 & ~n47870;
  assign n47872 = ~n47845 & ~n47871;
  assign n47873 = i_hlock7 & ~n47872;
  assign n47874 = i_hbusreq8 & ~n47831;
  assign n47875 = i_hbusreq6 & ~n47822;
  assign n47876 = ~n8217 & ~n37661;
  assign n47877 = ~n45490 & ~n47876;
  assign n47878 = i_hlock6 & ~n47877;
  assign n47879 = ~n8217 & ~n37672;
  assign n47880 = ~n45490 & ~n47879;
  assign n47881 = ~i_hlock6 & ~n47880;
  assign n47882 = ~n47878 & ~n47881;
  assign n47883 = ~i_hbusreq6 & ~n47882;
  assign n47884 = ~n47875 & ~n47883;
  assign n47885 = controllable_hgrant6 & ~n47884;
  assign n47886 = i_hbusreq6 & ~n47827;
  assign n47887 = controllable_hmaster2 & ~n47763;
  assign n47888 = ~n47058 & ~n47887;
  assign n47889 = controllable_hmaster1 & ~n47888;
  assign n47890 = ~n47159 & ~n47889;
  assign n47891 = ~i_hbusreq6 & ~n47890;
  assign n47892 = ~n47886 & ~n47891;
  assign n47893 = ~controllable_hgrant6 & ~n47892;
  assign n47894 = ~n47885 & ~n47893;
  assign n47895 = controllable_hmaster0 & ~n47894;
  assign n47896 = ~n47433 & ~n47895;
  assign n47897 = ~i_hbusreq8 & ~n47896;
  assign n47898 = ~n47874 & ~n47897;
  assign n47899 = ~controllable_hmaster3 & ~n47898;
  assign n47900 = ~n47845 & ~n47899;
  assign n47901 = ~i_hlock7 & ~n47900;
  assign n47902 = ~n47873 & ~n47901;
  assign n47903 = ~i_hbusreq7 & ~n47902;
  assign n47904 = ~n47836 & ~n47903;
  assign n47905 = n7924 & ~n47904;
  assign n47906 = ~n45418 & ~n47905;
  assign n47907 = ~n8214 & ~n47906;
  assign n47908 = ~n45699 & ~n47510;
  assign n47909 = controllable_hmaster0 & ~n47908;
  assign n47910 = ~n45709 & ~n46161;
  assign n47911 = ~controllable_hmaster0 & ~n47910;
  assign n47912 = ~n47909 & ~n47911;
  assign n47913 = i_hlock8 & ~n47912;
  assign n47914 = ~n45721 & ~n46219;
  assign n47915 = ~controllable_hmaster0 & ~n47914;
  assign n47916 = ~n47909 & ~n47915;
  assign n47917 = ~i_hlock8 & ~n47916;
  assign n47918 = ~n47913 & ~n47917;
  assign n47919 = controllable_hmaster3 & ~n47918;
  assign n47920 = ~n45735 & ~n46332;
  assign n47921 = controllable_hmaster0 & ~n47920;
  assign n47922 = ~n46406 & ~n47805;
  assign n47923 = controllable_hmaster1 & ~n47922;
  assign n47924 = ~n46476 & ~n47923;
  assign n47925 = i_hlock6 & ~n47924;
  assign n47926 = ~n46406 & ~n47824;
  assign n47927 = controllable_hmaster1 & ~n47926;
  assign n47928 = ~n46476 & ~n47927;
  assign n47929 = ~i_hlock6 & ~n47928;
  assign n47930 = ~n47925 & ~n47929;
  assign n47931 = ~controllable_hgrant6 & ~n47930;
  assign n47932 = ~n45751 & ~n47931;
  assign n47933 = ~controllable_hmaster0 & ~n47932;
  assign n47934 = ~n47921 & ~n47933;
  assign n47935 = ~controllable_hmaster3 & ~n47934;
  assign n47936 = ~n47919 & ~n47935;
  assign n47937 = i_hlock7 & ~n47936;
  assign n47938 = ~n45775 & ~n46503;
  assign n47939 = controllable_hmaster0 & ~n47938;
  assign n47940 = ~n47933 & ~n47939;
  assign n47941 = ~controllable_hmaster3 & ~n47940;
  assign n47942 = ~n47919 & ~n47941;
  assign n47943 = ~i_hlock7 & ~n47942;
  assign n47944 = ~n47937 & ~n47943;
  assign n47945 = i_hbusreq7 & ~n47944;
  assign n47946 = i_hbusreq8 & ~n47918;
  assign n47947 = ~n45796 & ~n47652;
  assign n47948 = controllable_hmaster0 & ~n47947;
  assign n47949 = ~n45810 & ~n46878;
  assign n47950 = ~controllable_hmaster0 & ~n47949;
  assign n47951 = ~n47948 & ~n47950;
  assign n47952 = i_hlock8 & ~n47951;
  assign n47953 = ~n45826 & ~n46975;
  assign n47954 = ~controllable_hmaster0 & ~n47953;
  assign n47955 = ~n47948 & ~n47954;
  assign n47956 = ~i_hlock8 & ~n47955;
  assign n47957 = ~n47952 & ~n47956;
  assign n47958 = ~i_hbusreq8 & ~n47957;
  assign n47959 = ~n47946 & ~n47958;
  assign n47960 = controllable_hmaster3 & ~n47959;
  assign n47961 = i_hbusreq8 & ~n47934;
  assign n47962 = ~n45847 & ~n47163;
  assign n47963 = controllable_hmaster0 & ~n47962;
  assign n47964 = i_hbusreq6 & ~n47930;
  assign n47965 = ~n47281 & ~n47859;
  assign n47966 = controllable_hmaster1 & ~n47965;
  assign n47967 = ~n47420 & ~n47966;
  assign n47968 = i_hlock6 & ~n47967;
  assign n47969 = ~n47281 & ~n47887;
  assign n47970 = controllable_hmaster1 & ~n47969;
  assign n47971 = ~n47420 & ~n47970;
  assign n47972 = ~i_hlock6 & ~n47971;
  assign n47973 = ~n47968 & ~n47972;
  assign n47974 = ~i_hbusreq6 & ~n47973;
  assign n47975 = ~n47964 & ~n47974;
  assign n47976 = ~controllable_hgrant6 & ~n47975;
  assign n47977 = ~n45874 & ~n47976;
  assign n47978 = ~controllable_hmaster0 & ~n47977;
  assign n47979 = ~n47963 & ~n47978;
  assign n47980 = ~i_hbusreq8 & ~n47979;
  assign n47981 = ~n47961 & ~n47980;
  assign n47982 = ~controllable_hmaster3 & ~n47981;
  assign n47983 = ~n47960 & ~n47982;
  assign n47984 = i_hlock7 & ~n47983;
  assign n47985 = i_hbusreq8 & ~n47940;
  assign n47986 = ~n45908 & ~n47458;
  assign n47987 = controllable_hmaster0 & ~n47986;
  assign n47988 = ~n47978 & ~n47987;
  assign n47989 = ~i_hbusreq8 & ~n47988;
  assign n47990 = ~n47985 & ~n47989;
  assign n47991 = ~controllable_hmaster3 & ~n47990;
  assign n47992 = ~n47960 & ~n47991;
  assign n47993 = ~i_hlock7 & ~n47992;
  assign n47994 = ~n47984 & ~n47993;
  assign n47995 = ~i_hbusreq7 & ~n47994;
  assign n47996 = ~n47945 & ~n47995;
  assign n47997 = n7924 & ~n47996;
  assign n47998 = ~n45691 & ~n47997;
  assign n47999 = n8214 & ~n47998;
  assign n48000 = ~n47907 & ~n47999;
  assign n48001 = n8202 & ~n48000;
  assign n48002 = ~n47790 & ~n48001;
  assign n48003 = n7920 & ~n48002;
  assign n48004 = ~n40177 & ~n48003;
  assign n48005 = n7728 & ~n48004;
  assign n48006 = ~n8378 & ~n17320;
  assign n48007 = ~n42706 & ~n48006;
  assign n48008 = controllable_hgrant5 & ~n48007;
  assign n48009 = ~n8426 & ~n17318;
  assign n48010 = ~n42710 & ~n48009;
  assign n48011 = controllable_hgrant4 & ~n48010;
  assign n48012 = ~n8365 & ~n17316;
  assign n48013 = ~n42714 & ~n48012;
  assign n48014 = controllable_hgrant3 & ~n48013;
  assign n48015 = ~n8389 & ~n17314;
  assign n48016 = ~n42718 & ~n48015;
  assign n48017 = controllable_hgrant1 & ~n48016;
  assign n48018 = controllable_hgrant2 & ~n40216;
  assign n48019 = ~n7936 & ~n48018;
  assign n48020 = ~n7733 & ~n48019;
  assign n48021 = ~n7936 & ~n40226;
  assign n48022 = n7733 & ~n48021;
  assign n48023 = ~n48020 & ~n48022;
  assign n48024 = ~controllable_hgrant1 & ~n48023;
  assign n48025 = ~n48017 & ~n48024;
  assign n48026 = ~controllable_hgrant3 & ~n48025;
  assign n48027 = ~n48014 & ~n48026;
  assign n48028 = ~controllable_hgrant4 & ~n48027;
  assign n48029 = ~n48011 & ~n48028;
  assign n48030 = ~controllable_hgrant5 & ~n48029;
  assign n48031 = ~n48008 & ~n48030;
  assign n48032 = controllable_hmaster1 & ~n48031;
  assign n48033 = controllable_hmaster2 & ~n48031;
  assign n48034 = ~n40256 & ~n48033;
  assign n48035 = ~controllable_hmaster1 & ~n48034;
  assign n48036 = ~n48032 & ~n48035;
  assign n48037 = ~controllable_hgrant6 & ~n48036;
  assign n48038 = ~n45520 & ~n48037;
  assign n48039 = controllable_hmaster0 & ~n48038;
  assign n48040 = ~n40437 & ~n48033;
  assign n48041 = ~controllable_hmaster1 & ~n48040;
  assign n48042 = ~n48032 & ~n48041;
  assign n48043 = ~controllable_hgrant6 & ~n48042;
  assign n48044 = ~n45525 & ~n48043;
  assign n48045 = ~controllable_hmaster0 & ~n48044;
  assign n48046 = ~n48039 & ~n48045;
  assign n48047 = i_hlock8 & ~n48046;
  assign n48048 = ~n40459 & ~n48033;
  assign n48049 = ~controllable_hmaster1 & ~n48048;
  assign n48050 = ~n48032 & ~n48049;
  assign n48051 = ~controllable_hgrant6 & ~n48050;
  assign n48052 = ~n45532 & ~n48051;
  assign n48053 = ~controllable_hmaster0 & ~n48052;
  assign n48054 = ~n48039 & ~n48053;
  assign n48055 = ~i_hlock8 & ~n48054;
  assign n48056 = ~n48047 & ~n48055;
  assign n48057 = controllable_hmaster3 & ~n48056;
  assign n48058 = ~n8378 & ~n18120;
  assign n48059 = ~n42821 & ~n48058;
  assign n48060 = controllable_hgrant5 & ~n48059;
  assign n48061 = ~n8426 & ~n18118;
  assign n48062 = ~n42825 & ~n48061;
  assign n48063 = controllable_hgrant4 & ~n48062;
  assign n48064 = ~n8365 & ~n16357;
  assign n48065 = ~n42829 & ~n48064;
  assign n48066 = i_hlock3 & ~n48065;
  assign n48067 = ~n8365 & ~n16363;
  assign n48068 = ~n42833 & ~n48067;
  assign n48069 = ~i_hlock3 & ~n48068;
  assign n48070 = ~n48066 & ~n48069;
  assign n48071 = controllable_hgrant3 & ~n48070;
  assign n48072 = i_hlock3 & ~n40233;
  assign n48073 = ~i_hlock3 & ~n40247;
  assign n48074 = ~n48072 & ~n48073;
  assign n48075 = ~controllable_hgrant3 & ~n48074;
  assign n48076 = ~n48071 & ~n48075;
  assign n48077 = ~controllable_hgrant4 & ~n48076;
  assign n48078 = ~n48063 & ~n48077;
  assign n48079 = ~controllable_hgrant5 & ~n48078;
  assign n48080 = ~n48060 & ~n48079;
  assign n48081 = ~controllable_hmaster2 & ~n48080;
  assign n48082 = ~n40579 & ~n48081;
  assign n48083 = controllable_hmaster1 & ~n48082;
  assign n48084 = ~n8378 & ~n28867;
  assign n48085 = ~n42851 & ~n48084;
  assign n48086 = i_hlock5 & ~n48085;
  assign n48087 = ~n8378 & ~n28882;
  assign n48088 = ~n42855 & ~n48087;
  assign n48089 = ~i_hlock5 & ~n48088;
  assign n48090 = ~n48086 & ~n48089;
  assign n48091 = controllable_hgrant5 & ~n48090;
  assign n48092 = i_hlock5 & ~n40434;
  assign n48093 = ~i_hlock5 & ~n40456;
  assign n48094 = ~n48092 & ~n48093;
  assign n48095 = ~controllable_hgrant5 & ~n48094;
  assign n48096 = ~n48091 & ~n48095;
  assign n48097 = controllable_hmaster2 & ~n48096;
  assign n48098 = ~n8378 & ~n18140;
  assign n48099 = ~n42867 & ~n48098;
  assign n48100 = controllable_hgrant5 & ~n48099;
  assign n48101 = ~n8426 & ~n18138;
  assign n48102 = ~n42871 & ~n48101;
  assign n48103 = controllable_hgrant4 & ~n48102;
  assign n48104 = ~n8365 & ~n18136;
  assign n48105 = ~n42875 & ~n48104;
  assign n48106 = controllable_hgrant3 & ~n48105;
  assign n48107 = ~n8389 & ~n16355;
  assign n48108 = ~n42879 & ~n48107;
  assign n48109 = i_hlock1 & ~n48108;
  assign n48110 = ~n8389 & ~n16361;
  assign n48111 = ~n42883 & ~n48110;
  assign n48112 = ~i_hlock1 & ~n48111;
  assign n48113 = ~n48109 & ~n48112;
  assign n48114 = controllable_hgrant1 & ~n48113;
  assign n48115 = i_hlock1 & ~n40231;
  assign n48116 = ~i_hlock1 & ~n40245;
  assign n48117 = ~n48115 & ~n48116;
  assign n48118 = ~controllable_hgrant1 & ~n48117;
  assign n48119 = ~n48114 & ~n48118;
  assign n48120 = ~controllable_hgrant3 & ~n48119;
  assign n48121 = ~n48106 & ~n48120;
  assign n48122 = ~controllable_hgrant4 & ~n48121;
  assign n48123 = ~n48103 & ~n48122;
  assign n48124 = ~controllable_hgrant5 & ~n48123;
  assign n48125 = ~n48100 & ~n48124;
  assign n48126 = ~controllable_hmaster2 & ~n48125;
  assign n48127 = ~n48097 & ~n48126;
  assign n48128 = ~controllable_hmaster1 & ~n48127;
  assign n48129 = ~n48083 & ~n48128;
  assign n48130 = ~controllable_hgrant6 & ~n48129;
  assign n48131 = ~n45541 & ~n48130;
  assign n48132 = controllable_hmaster0 & ~n48131;
  assign n48133 = ~n8378 & ~n18156;
  assign n48134 = ~n42929 & ~n48133;
  assign n48135 = controllable_hgrant5 & ~n48134;
  assign n48136 = ~n8426 & ~n18154;
  assign n48137 = ~n42933 & ~n48136;
  assign n48138 = controllable_hgrant4 & ~n48137;
  assign n48139 = ~n8365 & ~n18152;
  assign n48140 = ~n42937 & ~n48139;
  assign n48141 = controllable_hgrant3 & ~n48140;
  assign n48142 = ~n8389 & ~n18150;
  assign n48143 = ~n42941 & ~n48142;
  assign n48144 = controllable_hgrant1 & ~n48143;
  assign n48145 = ~n16998 & ~n42972;
  assign n48146 = ~n7733 & ~n48145;
  assign n48147 = ~n40222 & ~n42945;
  assign n48148 = controllable_locked & ~n48147;
  assign n48149 = ~n42970 & ~n48148;
  assign n48150 = controllable_hgrant2 & ~n48149;
  assign n48151 = ~n16998 & ~n48150;
  assign n48152 = n7733 & ~n48151;
  assign n48153 = ~n48146 & ~n48152;
  assign n48154 = n7928 & ~n48153;
  assign n48155 = ~n42965 & ~n48154;
  assign n48156 = ~controllable_hgrant1 & ~n48155;
  assign n48157 = ~n48144 & ~n48156;
  assign n48158 = ~controllable_hgrant3 & ~n48157;
  assign n48159 = ~n48141 & ~n48158;
  assign n48160 = ~controllable_hgrant4 & ~n48159;
  assign n48161 = ~n48138 & ~n48160;
  assign n48162 = ~controllable_hgrant5 & ~n48161;
  assign n48163 = ~n48135 & ~n48162;
  assign n48164 = ~controllable_hmaster2 & ~n48163;
  assign n48165 = ~n40579 & ~n48164;
  assign n48166 = controllable_hmaster1 & ~n48165;
  assign n48167 = ~n8378 & ~n18166;
  assign n48168 = ~n42987 & ~n48167;
  assign n48169 = controllable_hgrant5 & ~n48168;
  assign n48170 = ~n8426 & ~n16359;
  assign n48171 = ~n42991 & ~n48170;
  assign n48172 = i_hlock4 & ~n48171;
  assign n48173 = ~n8426 & ~n16365;
  assign n48174 = ~n42995 & ~n48173;
  assign n48175 = ~i_hlock4 & ~n48174;
  assign n48176 = ~n48172 & ~n48175;
  assign n48177 = controllable_hgrant4 & ~n48176;
  assign n48178 = i_hlock4 & ~n40235;
  assign n48179 = ~i_hlock4 & ~n40249;
  assign n48180 = ~n48178 & ~n48179;
  assign n48181 = ~controllable_hgrant4 & ~n48180;
  assign n48182 = ~n48177 & ~n48181;
  assign n48183 = ~controllable_hgrant5 & ~n48182;
  assign n48184 = ~n48169 & ~n48183;
  assign n48185 = controllable_hmaster2 & ~n48184;
  assign n48186 = ~n8378 & ~n18176;
  assign n48187 = ~n43009 & ~n48186;
  assign n48188 = controllable_hgrant5 & ~n48187;
  assign n48189 = ~n8426 & ~n18174;
  assign n48190 = ~n43013 & ~n48189;
  assign n48191 = controllable_hgrant4 & ~n48190;
  assign n48192 = ~n8365 & ~n18172;
  assign n48193 = ~n43017 & ~n48192;
  assign n48194 = controllable_hgrant3 & ~n48193;
  assign n48195 = ~n8389 & ~n18170;
  assign n48196 = ~n43021 & ~n48195;
  assign n48197 = controllable_hgrant1 & ~n48196;
  assign n48198 = ~n8440 & ~n40230;
  assign n48199 = ~controllable_hgrant1 & ~n48198;
  assign n48200 = ~n48197 & ~n48199;
  assign n48201 = ~controllable_hgrant3 & ~n48200;
  assign n48202 = ~n48194 & ~n48201;
  assign n48203 = ~controllable_hgrant4 & ~n48202;
  assign n48204 = ~n48191 & ~n48203;
  assign n48205 = ~controllable_hgrant5 & ~n48204;
  assign n48206 = ~n48188 & ~n48205;
  assign n48207 = ~controllable_hmaster2 & ~n48206;
  assign n48208 = ~n48185 & ~n48207;
  assign n48209 = ~controllable_hmaster1 & ~n48208;
  assign n48210 = ~n48166 & ~n48209;
  assign n48211 = i_hlock6 & ~n48210;
  assign n48212 = ~n40594 & ~n48164;
  assign n48213 = controllable_hmaster1 & ~n48212;
  assign n48214 = ~n48209 & ~n48213;
  assign n48215 = ~i_hlock6 & ~n48214;
  assign n48216 = ~n48211 & ~n48215;
  assign n48217 = ~controllable_hgrant6 & ~n48216;
  assign n48218 = ~n45557 & ~n48217;
  assign n48219 = ~controllable_hmaster0 & ~n48218;
  assign n48220 = ~n48132 & ~n48219;
  assign n48221 = ~controllable_hmaster3 & ~n48220;
  assign n48222 = ~n48057 & ~n48221;
  assign n48223 = i_hlock7 & ~n48222;
  assign n48224 = ~n40594 & ~n48081;
  assign n48225 = controllable_hmaster1 & ~n48224;
  assign n48226 = ~n48128 & ~n48225;
  assign n48227 = ~controllable_hgrant6 & ~n48226;
  assign n48228 = ~n45576 & ~n48227;
  assign n48229 = controllable_hmaster0 & ~n48228;
  assign n48230 = ~n48219 & ~n48229;
  assign n48231 = ~controllable_hmaster3 & ~n48230;
  assign n48232 = ~n48057 & ~n48231;
  assign n48233 = ~i_hlock7 & ~n48232;
  assign n48234 = ~n48223 & ~n48233;
  assign n48235 = i_hbusreq7 & ~n48234;
  assign n48236 = i_hbusreq8 & ~n48056;
  assign n48237 = n8217 & ~n9603;
  assign n48238 = ~n8217 & ~n31992;
  assign n48239 = ~n48237 & ~n48238;
  assign n48240 = ~i_hbusreq6 & ~n48239;
  assign n48241 = ~n45586 & ~n48240;
  assign n48242 = controllable_hgrant6 & ~n48241;
  assign n48243 = i_hbusreq6 & ~n48036;
  assign n48244 = i_hbusreq5 & ~n48007;
  assign n48245 = n8378 & ~n9596;
  assign n48246 = ~n8378 & ~n21643;
  assign n48247 = ~n48245 & ~n48246;
  assign n48248 = ~i_hbusreq5 & ~n48247;
  assign n48249 = ~n48244 & ~n48248;
  assign n48250 = controllable_hgrant5 & ~n48249;
  assign n48251 = i_hbusreq5 & ~n48029;
  assign n48252 = i_hbusreq4 & ~n48010;
  assign n48253 = i_hbusreq9 & ~n48010;
  assign n48254 = n8426 & ~n9592;
  assign n48255 = ~n8426 & ~n21637;
  assign n48256 = ~n48254 & ~n48255;
  assign n48257 = ~i_hbusreq9 & ~n48256;
  assign n48258 = ~n48253 & ~n48257;
  assign n48259 = ~i_hbusreq4 & ~n48258;
  assign n48260 = ~n48252 & ~n48259;
  assign n48261 = controllable_hgrant4 & ~n48260;
  assign n48262 = i_hbusreq4 & ~n48027;
  assign n48263 = i_hbusreq9 & ~n48027;
  assign n48264 = i_hbusreq3 & ~n48013;
  assign n48265 = n8365 & ~n9590;
  assign n48266 = ~n8365 & ~n21633;
  assign n48267 = ~n48265 & ~n48266;
  assign n48268 = ~i_hbusreq3 & ~n48267;
  assign n48269 = ~n48264 & ~n48268;
  assign n48270 = controllable_hgrant3 & ~n48269;
  assign n48271 = i_hbusreq3 & ~n48025;
  assign n48272 = i_hbusreq1 & ~n48016;
  assign n48273 = n8389 & ~n9588;
  assign n48274 = ~n8389 & ~n21629;
  assign n48275 = ~n48273 & ~n48274;
  assign n48276 = ~i_hbusreq1 & ~n48275;
  assign n48277 = ~n48272 & ~n48276;
  assign n48278 = controllable_hgrant1 & ~n48277;
  assign n48279 = i_hbusreq1 & ~n48023;
  assign n48280 = ~n16414 & ~n40348;
  assign n48281 = n7733 & ~n48280;
  assign n48282 = ~n48020 & ~n48281;
  assign n48283 = ~i_hbusreq1 & ~n48282;
  assign n48284 = ~n48279 & ~n48283;
  assign n48285 = ~controllable_hgrant1 & ~n48284;
  assign n48286 = ~n48278 & ~n48285;
  assign n48287 = ~i_hbusreq3 & ~n48286;
  assign n48288 = ~n48271 & ~n48287;
  assign n48289 = ~controllable_hgrant3 & ~n48288;
  assign n48290 = ~n48270 & ~n48289;
  assign n48291 = ~i_hbusreq9 & ~n48290;
  assign n48292 = ~n48263 & ~n48291;
  assign n48293 = ~i_hbusreq4 & ~n48292;
  assign n48294 = ~n48262 & ~n48293;
  assign n48295 = ~controllable_hgrant4 & ~n48294;
  assign n48296 = ~n48261 & ~n48295;
  assign n48297 = ~i_hbusreq5 & ~n48296;
  assign n48298 = ~n48251 & ~n48297;
  assign n48299 = ~controllable_hgrant5 & ~n48298;
  assign n48300 = ~n48250 & ~n48299;
  assign n48301 = controllable_hmaster1 & ~n48300;
  assign n48302 = controllable_hmaster2 & ~n48300;
  assign n48303 = ~n40407 & ~n48302;
  assign n48304 = ~controllable_hmaster1 & ~n48303;
  assign n48305 = ~n48301 & ~n48304;
  assign n48306 = ~i_hbusreq6 & ~n48305;
  assign n48307 = ~n48243 & ~n48306;
  assign n48308 = ~controllable_hgrant6 & ~n48307;
  assign n48309 = ~n48242 & ~n48308;
  assign n48310 = controllable_hmaster0 & ~n48309;
  assign n48311 = n8217 & ~n9609;
  assign n48312 = ~n8217 & ~n21660;
  assign n48313 = ~n48311 & ~n48312;
  assign n48314 = ~i_hbusreq6 & ~n48313;
  assign n48315 = ~n45594 & ~n48314;
  assign n48316 = controllable_hgrant6 & ~n48315;
  assign n48317 = i_hbusreq6 & ~n48042;
  assign n48318 = ~n40508 & ~n48302;
  assign n48319 = ~controllable_hmaster1 & ~n48318;
  assign n48320 = ~n48301 & ~n48319;
  assign n48321 = ~i_hbusreq6 & ~n48320;
  assign n48322 = ~n48317 & ~n48321;
  assign n48323 = ~controllable_hgrant6 & ~n48322;
  assign n48324 = ~n48316 & ~n48323;
  assign n48325 = ~controllable_hmaster0 & ~n48324;
  assign n48326 = ~n48310 & ~n48325;
  assign n48327 = i_hlock8 & ~n48326;
  assign n48328 = n8217 & ~n9617;
  assign n48329 = ~n8217 & ~n21670;
  assign n48330 = ~n48328 & ~n48329;
  assign n48331 = ~i_hbusreq6 & ~n48330;
  assign n48332 = ~n45604 & ~n48331;
  assign n48333 = controllable_hgrant6 & ~n48332;
  assign n48334 = i_hbusreq6 & ~n48050;
  assign n48335 = ~n40554 & ~n48302;
  assign n48336 = ~controllable_hmaster1 & ~n48335;
  assign n48337 = ~n48301 & ~n48336;
  assign n48338 = ~i_hbusreq6 & ~n48337;
  assign n48339 = ~n48334 & ~n48338;
  assign n48340 = ~controllable_hgrant6 & ~n48339;
  assign n48341 = ~n48333 & ~n48340;
  assign n48342 = ~controllable_hmaster0 & ~n48341;
  assign n48343 = ~n48310 & ~n48342;
  assign n48344 = ~i_hlock8 & ~n48343;
  assign n48345 = ~n48327 & ~n48344;
  assign n48346 = ~i_hbusreq8 & ~n48345;
  assign n48347 = ~n48236 & ~n48346;
  assign n48348 = controllable_hmaster3 & ~n48347;
  assign n48349 = i_hbusreq8 & ~n48220;
  assign n48350 = n8217 & ~n9663;
  assign n48351 = ~n8217 & ~n21734;
  assign n48352 = ~n48350 & ~n48351;
  assign n48353 = ~i_hbusreq6 & ~n48352;
  assign n48354 = ~n45619 & ~n48353;
  assign n48355 = controllable_hgrant6 & ~n48354;
  assign n48356 = i_hbusreq6 & ~n48129;
  assign n48357 = i_hbusreq5 & ~n48059;
  assign n48358 = n8378 & ~n9635;
  assign n48359 = ~n8378 & ~n21694;
  assign n48360 = ~n48358 & ~n48359;
  assign n48361 = ~i_hbusreq5 & ~n48360;
  assign n48362 = ~n48357 & ~n48361;
  assign n48363 = controllable_hgrant5 & ~n48362;
  assign n48364 = i_hbusreq5 & ~n48078;
  assign n48365 = i_hbusreq4 & ~n48062;
  assign n48366 = i_hbusreq9 & ~n48062;
  assign n48367 = n8426 & ~n9631;
  assign n48368 = ~n8426 & ~n21688;
  assign n48369 = ~n48367 & ~n48368;
  assign n48370 = ~i_hbusreq9 & ~n48369;
  assign n48371 = ~n48366 & ~n48370;
  assign n48372 = ~i_hbusreq4 & ~n48371;
  assign n48373 = ~n48365 & ~n48372;
  assign n48374 = controllable_hgrant4 & ~n48373;
  assign n48375 = i_hbusreq4 & ~n48076;
  assign n48376 = i_hbusreq9 & ~n48076;
  assign n48377 = i_hbusreq3 & ~n48070;
  assign n48378 = n8365 & ~n12722;
  assign n48379 = ~n8365 & ~n16423;
  assign n48380 = ~n48378 & ~n48379;
  assign n48381 = i_hlock3 & ~n48380;
  assign n48382 = n8365 & ~n12747;
  assign n48383 = ~n8365 & ~n16435;
  assign n48384 = ~n48382 & ~n48383;
  assign n48385 = ~i_hlock3 & ~n48384;
  assign n48386 = ~n48381 & ~n48385;
  assign n48387 = ~i_hbusreq3 & ~n48386;
  assign n48388 = ~n48377 & ~n48387;
  assign n48389 = controllable_hgrant3 & ~n48388;
  assign n48390 = i_hbusreq3 & ~n48074;
  assign n48391 = i_hlock3 & ~n40364;
  assign n48392 = ~i_hlock3 & ~n40390;
  assign n48393 = ~n48391 & ~n48392;
  assign n48394 = ~i_hbusreq3 & ~n48393;
  assign n48395 = ~n48390 & ~n48394;
  assign n48396 = ~controllable_hgrant3 & ~n48395;
  assign n48397 = ~n48389 & ~n48396;
  assign n48398 = ~i_hbusreq9 & ~n48397;
  assign n48399 = ~n48376 & ~n48398;
  assign n48400 = ~i_hbusreq4 & ~n48399;
  assign n48401 = ~n48375 & ~n48400;
  assign n48402 = ~controllable_hgrant4 & ~n48401;
  assign n48403 = ~n48374 & ~n48402;
  assign n48404 = ~i_hbusreq5 & ~n48403;
  assign n48405 = ~n48364 & ~n48404;
  assign n48406 = ~controllable_hgrant5 & ~n48405;
  assign n48407 = ~n48363 & ~n48406;
  assign n48408 = ~controllable_hmaster2 & ~n48407;
  assign n48409 = ~n40616 & ~n48408;
  assign n48410 = controllable_hmaster1 & ~n48409;
  assign n48411 = i_hbusreq5 & ~n48090;
  assign n48412 = n8378 & ~n26679;
  assign n48413 = ~n8378 & ~n28908;
  assign n48414 = ~n48412 & ~n48413;
  assign n48415 = i_hlock5 & ~n48414;
  assign n48416 = n8378 & ~n26709;
  assign n48417 = ~n8378 & ~n28938;
  assign n48418 = ~n48416 & ~n48417;
  assign n48419 = ~i_hlock5 & ~n48418;
  assign n48420 = ~n48415 & ~n48419;
  assign n48421 = ~i_hbusreq5 & ~n48420;
  assign n48422 = ~n48411 & ~n48421;
  assign n48423 = controllable_hgrant5 & ~n48422;
  assign n48424 = i_hbusreq5 & ~n48094;
  assign n48425 = i_hlock5 & ~n40503;
  assign n48426 = ~i_hlock5 & ~n40549;
  assign n48427 = ~n48425 & ~n48426;
  assign n48428 = ~i_hbusreq5 & ~n48427;
  assign n48429 = ~n48424 & ~n48428;
  assign n48430 = ~controllable_hgrant5 & ~n48429;
  assign n48431 = ~n48423 & ~n48430;
  assign n48432 = controllable_hmaster2 & ~n48431;
  assign n48433 = i_hbusreq5 & ~n48099;
  assign n48434 = n8378 & ~n9657;
  assign n48435 = ~n8378 & ~n21726;
  assign n48436 = ~n48434 & ~n48435;
  assign n48437 = ~i_hbusreq5 & ~n48436;
  assign n48438 = ~n48433 & ~n48437;
  assign n48439 = controllable_hgrant5 & ~n48438;
  assign n48440 = i_hbusreq5 & ~n48123;
  assign n48441 = i_hbusreq4 & ~n48102;
  assign n48442 = i_hbusreq9 & ~n48102;
  assign n48443 = n8426 & ~n9653;
  assign n48444 = ~n8426 & ~n21720;
  assign n48445 = ~n48443 & ~n48444;
  assign n48446 = ~i_hbusreq9 & ~n48445;
  assign n48447 = ~n48442 & ~n48446;
  assign n48448 = ~i_hbusreq4 & ~n48447;
  assign n48449 = ~n48441 & ~n48448;
  assign n48450 = controllable_hgrant4 & ~n48449;
  assign n48451 = i_hbusreq4 & ~n48121;
  assign n48452 = i_hbusreq9 & ~n48121;
  assign n48453 = i_hbusreq3 & ~n48105;
  assign n48454 = n8365 & ~n9651;
  assign n48455 = ~n8365 & ~n21716;
  assign n48456 = ~n48454 & ~n48455;
  assign n48457 = ~i_hbusreq3 & ~n48456;
  assign n48458 = ~n48453 & ~n48457;
  assign n48459 = controllable_hgrant3 & ~n48458;
  assign n48460 = i_hbusreq3 & ~n48119;
  assign n48461 = i_hbusreq1 & ~n48113;
  assign n48462 = n8389 & ~n12718;
  assign n48463 = ~n8389 & ~n16419;
  assign n48464 = ~n48462 & ~n48463;
  assign n48465 = i_hlock1 & ~n48464;
  assign n48466 = n8389 & ~n12743;
  assign n48467 = ~n8389 & ~n16431;
  assign n48468 = ~n48466 & ~n48467;
  assign n48469 = ~i_hlock1 & ~n48468;
  assign n48470 = ~n48465 & ~n48469;
  assign n48471 = ~i_hbusreq1 & ~n48470;
  assign n48472 = ~n48461 & ~n48471;
  assign n48473 = controllable_hgrant1 & ~n48472;
  assign n48474 = i_hbusreq1 & ~n48117;
  assign n48475 = i_hlock1 & ~n40360;
  assign n48476 = ~i_hlock1 & ~n40386;
  assign n48477 = ~n48475 & ~n48476;
  assign n48478 = ~i_hbusreq1 & ~n48477;
  assign n48479 = ~n48474 & ~n48478;
  assign n48480 = ~controllable_hgrant1 & ~n48479;
  assign n48481 = ~n48473 & ~n48480;
  assign n48482 = ~i_hbusreq3 & ~n48481;
  assign n48483 = ~n48460 & ~n48482;
  assign n48484 = ~controllable_hgrant3 & ~n48483;
  assign n48485 = ~n48459 & ~n48484;
  assign n48486 = ~i_hbusreq9 & ~n48485;
  assign n48487 = ~n48452 & ~n48486;
  assign n48488 = ~i_hbusreq4 & ~n48487;
  assign n48489 = ~n48451 & ~n48488;
  assign n48490 = ~controllable_hgrant4 & ~n48489;
  assign n48491 = ~n48450 & ~n48490;
  assign n48492 = ~i_hbusreq5 & ~n48491;
  assign n48493 = ~n48440 & ~n48492;
  assign n48494 = ~controllable_hgrant5 & ~n48493;
  assign n48495 = ~n48439 & ~n48494;
  assign n48496 = ~controllable_hmaster2 & ~n48495;
  assign n48497 = ~n48432 & ~n48496;
  assign n48498 = ~controllable_hmaster1 & ~n48497;
  assign n48499 = ~n48410 & ~n48498;
  assign n48500 = ~i_hbusreq6 & ~n48499;
  assign n48501 = ~n48356 & ~n48500;
  assign n48502 = ~controllable_hgrant6 & ~n48501;
  assign n48503 = ~n48355 & ~n48502;
  assign n48504 = controllable_hmaster0 & ~n48503;
  assign n48505 = ~n9678 & ~n26684;
  assign n48506 = controllable_hmaster1 & ~n48505;
  assign n48507 = ~n9706 & ~n48506;
  assign n48508 = n8217 & ~n48507;
  assign n48509 = ~n21759 & ~n28913;
  assign n48510 = controllable_hmaster1 & ~n48509;
  assign n48511 = ~n21797 & ~n48510;
  assign n48512 = ~n8217 & ~n48511;
  assign n48513 = ~n48508 & ~n48512;
  assign n48514 = i_hlock6 & ~n48513;
  assign n48515 = ~n9678 & ~n26714;
  assign n48516 = controllable_hmaster1 & ~n48515;
  assign n48517 = ~n9706 & ~n48516;
  assign n48518 = n8217 & ~n48517;
  assign n48519 = ~n21759 & ~n28943;
  assign n48520 = controllable_hmaster1 & ~n48519;
  assign n48521 = ~n21797 & ~n48520;
  assign n48522 = ~n8217 & ~n48521;
  assign n48523 = ~n48518 & ~n48522;
  assign n48524 = ~i_hlock6 & ~n48523;
  assign n48525 = ~n48514 & ~n48524;
  assign n48526 = ~i_hbusreq6 & ~n48525;
  assign n48527 = ~n45627 & ~n48526;
  assign n48528 = controllable_hgrant6 & ~n48527;
  assign n48529 = i_hbusreq6 & ~n48216;
  assign n48530 = i_hbusreq5 & ~n48134;
  assign n48531 = n8378 & ~n9675;
  assign n48532 = ~n8378 & ~n21754;
  assign n48533 = ~n48531 & ~n48532;
  assign n48534 = ~i_hbusreq5 & ~n48533;
  assign n48535 = ~n48530 & ~n48534;
  assign n48536 = controllable_hgrant5 & ~n48535;
  assign n48537 = i_hbusreq5 & ~n48161;
  assign n48538 = i_hbusreq4 & ~n48137;
  assign n48539 = i_hbusreq9 & ~n48137;
  assign n48540 = n8426 & ~n9671;
  assign n48541 = ~n8426 & ~n21748;
  assign n48542 = ~n48540 & ~n48541;
  assign n48543 = ~i_hbusreq9 & ~n48542;
  assign n48544 = ~n48539 & ~n48543;
  assign n48545 = ~i_hbusreq4 & ~n48544;
  assign n48546 = ~n48538 & ~n48545;
  assign n48547 = controllable_hgrant4 & ~n48546;
  assign n48548 = i_hbusreq4 & ~n48159;
  assign n48549 = i_hbusreq9 & ~n48159;
  assign n48550 = i_hbusreq3 & ~n48140;
  assign n48551 = n8365 & ~n9669;
  assign n48552 = ~n8365 & ~n21744;
  assign n48553 = ~n48551 & ~n48552;
  assign n48554 = ~i_hbusreq3 & ~n48553;
  assign n48555 = ~n48550 & ~n48554;
  assign n48556 = controllable_hgrant3 & ~n48555;
  assign n48557 = i_hbusreq3 & ~n48157;
  assign n48558 = i_hbusreq1 & ~n48143;
  assign n48559 = n8389 & ~n9667;
  assign n48560 = ~n8389 & ~n21740;
  assign n48561 = ~n48559 & ~n48560;
  assign n48562 = ~i_hbusreq1 & ~n48561;
  assign n48563 = ~n48558 & ~n48562;
  assign n48564 = controllable_hgrant1 & ~n48563;
  assign n48565 = i_hbusreq1 & ~n48155;
  assign n48566 = ~n18216 & ~n43558;
  assign n48567 = ~n7733 & ~n48566;
  assign n48568 = i_hbusreq2 & ~n48149;
  assign n48569 = i_hbusreq0 & ~n48149;
  assign n48570 = ~n39853 & ~n40222;
  assign n48571 = controllable_locked & ~n48570;
  assign n48572 = ~n40337 & ~n42954;
  assign n48573 = ~controllable_locked & ~n48572;
  assign n48574 = ~n48571 & ~n48573;
  assign n48575 = i_hlock0 & ~n48574;
  assign n48576 = ~i_hlock0 & ~n48149;
  assign n48577 = ~n48575 & ~n48576;
  assign n48578 = ~i_hbusreq0 & ~n48577;
  assign n48579 = ~n48569 & ~n48578;
  assign n48580 = ~i_hbusreq2 & ~n48579;
  assign n48581 = ~n48568 & ~n48580;
  assign n48582 = controllable_hgrant2 & ~n48581;
  assign n48583 = ~n40355 & ~n48582;
  assign n48584 = n7733 & ~n48583;
  assign n48585 = ~n48567 & ~n48584;
  assign n48586 = n7928 & ~n48585;
  assign n48587 = ~n43545 & ~n48586;
  assign n48588 = ~i_hbusreq1 & ~n48587;
  assign n48589 = ~n48565 & ~n48588;
  assign n48590 = ~controllable_hgrant1 & ~n48589;
  assign n48591 = ~n48564 & ~n48590;
  assign n48592 = ~i_hbusreq3 & ~n48591;
  assign n48593 = ~n48557 & ~n48592;
  assign n48594 = ~controllable_hgrant3 & ~n48593;
  assign n48595 = ~n48556 & ~n48594;
  assign n48596 = ~i_hbusreq9 & ~n48595;
  assign n48597 = ~n48549 & ~n48596;
  assign n48598 = ~i_hbusreq4 & ~n48597;
  assign n48599 = ~n48548 & ~n48598;
  assign n48600 = ~controllable_hgrant4 & ~n48599;
  assign n48601 = ~n48547 & ~n48600;
  assign n48602 = ~i_hbusreq5 & ~n48601;
  assign n48603 = ~n48537 & ~n48602;
  assign n48604 = ~controllable_hgrant5 & ~n48603;
  assign n48605 = ~n48536 & ~n48604;
  assign n48606 = ~controllable_hmaster2 & ~n48605;
  assign n48607 = ~n40616 & ~n48606;
  assign n48608 = controllable_hmaster1 & ~n48607;
  assign n48609 = i_hbusreq5 & ~n48168;
  assign n48610 = n8378 & ~n9685;
  assign n48611 = ~n8378 & ~n21768;
  assign n48612 = ~n48610 & ~n48611;
  assign n48613 = ~i_hbusreq5 & ~n48612;
  assign n48614 = ~n48609 & ~n48613;
  assign n48615 = controllable_hgrant5 & ~n48614;
  assign n48616 = i_hbusreq5 & ~n48182;
  assign n48617 = i_hbusreq4 & ~n48176;
  assign n48618 = i_hbusreq9 & ~n48171;
  assign n48619 = n8426 & ~n12726;
  assign n48620 = ~n8426 & ~n16427;
  assign n48621 = ~n48619 & ~n48620;
  assign n48622 = ~i_hbusreq9 & ~n48621;
  assign n48623 = ~n48618 & ~n48622;
  assign n48624 = i_hlock4 & ~n48623;
  assign n48625 = i_hbusreq9 & ~n48174;
  assign n48626 = n8426 & ~n12751;
  assign n48627 = ~n8426 & ~n16439;
  assign n48628 = ~n48626 & ~n48627;
  assign n48629 = ~i_hbusreq9 & ~n48628;
  assign n48630 = ~n48625 & ~n48629;
  assign n48631 = ~i_hlock4 & ~n48630;
  assign n48632 = ~n48624 & ~n48631;
  assign n48633 = ~i_hbusreq4 & ~n48632;
  assign n48634 = ~n48617 & ~n48633;
  assign n48635 = controllable_hgrant4 & ~n48634;
  assign n48636 = i_hbusreq4 & ~n48180;
  assign n48637 = i_hlock4 & ~n40499;
  assign n48638 = ~i_hlock4 & ~n40545;
  assign n48639 = ~n48637 & ~n48638;
  assign n48640 = ~i_hbusreq4 & ~n48639;
  assign n48641 = ~n48636 & ~n48640;
  assign n48642 = ~controllable_hgrant4 & ~n48641;
  assign n48643 = ~n48635 & ~n48642;
  assign n48644 = ~i_hbusreq5 & ~n48643;
  assign n48645 = ~n48616 & ~n48644;
  assign n48646 = ~controllable_hgrant5 & ~n48645;
  assign n48647 = ~n48615 & ~n48646;
  assign n48648 = controllable_hmaster2 & ~n48647;
  assign n48649 = i_hbusreq5 & ~n48187;
  assign n48650 = n8378 & ~n9701;
  assign n48651 = ~n8378 & ~n21790;
  assign n48652 = ~n48650 & ~n48651;
  assign n48653 = ~i_hbusreq5 & ~n48652;
  assign n48654 = ~n48649 & ~n48653;
  assign n48655 = controllable_hgrant5 & ~n48654;
  assign n48656 = i_hbusreq5 & ~n48204;
  assign n48657 = i_hbusreq4 & ~n48190;
  assign n48658 = i_hbusreq9 & ~n48190;
  assign n48659 = n8426 & ~n9697;
  assign n48660 = ~n8426 & ~n21784;
  assign n48661 = ~n48659 & ~n48660;
  assign n48662 = ~i_hbusreq9 & ~n48661;
  assign n48663 = ~n48658 & ~n48662;
  assign n48664 = ~i_hbusreq4 & ~n48663;
  assign n48665 = ~n48657 & ~n48664;
  assign n48666 = controllable_hgrant4 & ~n48665;
  assign n48667 = i_hbusreq4 & ~n48202;
  assign n48668 = i_hbusreq9 & ~n48202;
  assign n48669 = i_hbusreq3 & ~n48193;
  assign n48670 = n8365 & ~n9695;
  assign n48671 = ~n8365 & ~n21780;
  assign n48672 = ~n48670 & ~n48671;
  assign n48673 = ~i_hbusreq3 & ~n48672;
  assign n48674 = ~n48669 & ~n48673;
  assign n48675 = controllable_hgrant3 & ~n48674;
  assign n48676 = i_hbusreq3 & ~n48200;
  assign n48677 = i_hbusreq1 & ~n48196;
  assign n48678 = n8389 & ~n9693;
  assign n48679 = ~n8389 & ~n21776;
  assign n48680 = ~n48678 & ~n48679;
  assign n48681 = ~i_hbusreq1 & ~n48680;
  assign n48682 = ~n48677 & ~n48681;
  assign n48683 = controllable_hgrant1 & ~n48682;
  assign n48684 = i_hbusreq1 & ~n48198;
  assign n48685 = i_hlock0 & ~n18443;
  assign n48686 = ~n18210 & ~n48685;
  assign n48687 = ~i_hbusreq0 & ~n48686;
  assign n48688 = ~n8106 & ~n48687;
  assign n48689 = ~i_hbusreq2 & ~n48688;
  assign n48690 = ~n8105 & ~n48689;
  assign n48691 = ~controllable_hgrant2 & ~n48690;
  assign n48692 = ~n43669 & ~n48691;
  assign n48693 = ~n7733 & ~n48692;
  assign n48694 = ~n40228 & ~n48693;
  assign n48695 = n7928 & ~n48694;
  assign n48696 = ~n8440 & ~n48695;
  assign n48697 = ~i_hbusreq1 & ~n48696;
  assign n48698 = ~n48684 & ~n48697;
  assign n48699 = ~controllable_hgrant1 & ~n48698;
  assign n48700 = ~n48683 & ~n48699;
  assign n48701 = ~i_hbusreq3 & ~n48700;
  assign n48702 = ~n48676 & ~n48701;
  assign n48703 = ~controllable_hgrant3 & ~n48702;
  assign n48704 = ~n48675 & ~n48703;
  assign n48705 = ~i_hbusreq9 & ~n48704;
  assign n48706 = ~n48668 & ~n48705;
  assign n48707 = ~i_hbusreq4 & ~n48706;
  assign n48708 = ~n48667 & ~n48707;
  assign n48709 = ~controllable_hgrant4 & ~n48708;
  assign n48710 = ~n48666 & ~n48709;
  assign n48711 = ~i_hbusreq5 & ~n48710;
  assign n48712 = ~n48656 & ~n48711;
  assign n48713 = ~controllable_hgrant5 & ~n48712;
  assign n48714 = ~n48655 & ~n48713;
  assign n48715 = ~controllable_hmaster2 & ~n48714;
  assign n48716 = ~n48648 & ~n48715;
  assign n48717 = ~controllable_hmaster1 & ~n48716;
  assign n48718 = ~n48608 & ~n48717;
  assign n48719 = i_hlock6 & ~n48718;
  assign n48720 = ~n40640 & ~n48606;
  assign n48721 = controllable_hmaster1 & ~n48720;
  assign n48722 = ~n48717 & ~n48721;
  assign n48723 = ~i_hlock6 & ~n48722;
  assign n48724 = ~n48719 & ~n48723;
  assign n48725 = ~i_hbusreq6 & ~n48724;
  assign n48726 = ~n48529 & ~n48725;
  assign n48727 = ~controllable_hgrant6 & ~n48726;
  assign n48728 = ~n48528 & ~n48727;
  assign n48729 = ~controllable_hmaster0 & ~n48728;
  assign n48730 = ~n48504 & ~n48729;
  assign n48731 = ~i_hbusreq8 & ~n48730;
  assign n48732 = ~n48349 & ~n48731;
  assign n48733 = ~controllable_hmaster3 & ~n48732;
  assign n48734 = ~n48348 & ~n48733;
  assign n48735 = i_hlock7 & ~n48734;
  assign n48736 = i_hbusreq8 & ~n48230;
  assign n48737 = n8217 & ~n9725;
  assign n48738 = ~n8217 & ~n21818;
  assign n48739 = ~n48737 & ~n48738;
  assign n48740 = ~i_hbusreq6 & ~n48739;
  assign n48741 = ~n45674 & ~n48740;
  assign n48742 = controllable_hgrant6 & ~n48741;
  assign n48743 = i_hbusreq6 & ~n48226;
  assign n48744 = ~n40640 & ~n48408;
  assign n48745 = controllable_hmaster1 & ~n48744;
  assign n48746 = ~n48498 & ~n48745;
  assign n48747 = ~i_hbusreq6 & ~n48746;
  assign n48748 = ~n48743 & ~n48747;
  assign n48749 = ~controllable_hgrant6 & ~n48748;
  assign n48750 = ~n48742 & ~n48749;
  assign n48751 = controllable_hmaster0 & ~n48750;
  assign n48752 = ~n48729 & ~n48751;
  assign n48753 = ~i_hbusreq8 & ~n48752;
  assign n48754 = ~n48736 & ~n48753;
  assign n48755 = ~controllable_hmaster3 & ~n48754;
  assign n48756 = ~n48348 & ~n48755;
  assign n48757 = ~i_hlock7 & ~n48756;
  assign n48758 = ~n48735 & ~n48757;
  assign n48759 = ~i_hbusreq7 & ~n48758;
  assign n48760 = ~n48235 & ~n48759;
  assign n48761 = ~n7924 & ~n48760;
  assign n48762 = ~n8378 & ~n29488;
  assign n48763 = ~n43743 & ~n48762;
  assign n48764 = i_hlock5 & ~n48763;
  assign n48765 = ~n8378 & ~n29519;
  assign n48766 = ~n43743 & ~n48765;
  assign n48767 = ~i_hlock5 & ~n48766;
  assign n48768 = ~n48764 & ~n48767;
  assign n48769 = controllable_hgrant5 & ~n48768;
  assign n48770 = ~n8426 & ~n17474;
  assign n48771 = ~n43747 & ~n48770;
  assign n48772 = i_hlock4 & ~n48771;
  assign n48773 = ~n8426 & ~n17490;
  assign n48774 = ~n43747 & ~n48773;
  assign n48775 = ~i_hlock4 & ~n48774;
  assign n48776 = ~n48772 & ~n48775;
  assign n48777 = controllable_hgrant4 & ~n48776;
  assign n48778 = ~n8365 & ~n17472;
  assign n48779 = ~n43751 & ~n48778;
  assign n48780 = i_hlock3 & ~n48779;
  assign n48781 = ~n8365 & ~n17488;
  assign n48782 = ~n43751 & ~n48781;
  assign n48783 = ~i_hlock3 & ~n48782;
  assign n48784 = ~n48780 & ~n48783;
  assign n48785 = controllable_hgrant3 & ~n48784;
  assign n48786 = ~n8389 & ~n17470;
  assign n48787 = ~n43755 & ~n48786;
  assign n48788 = i_hlock1 & ~n48787;
  assign n48789 = ~n8389 & ~n17486;
  assign n48790 = ~n43755 & ~n48789;
  assign n48791 = ~i_hlock1 & ~n48790;
  assign n48792 = ~n48788 & ~n48791;
  assign n48793 = controllable_hgrant1 & ~n48792;
  assign n48794 = ~n7928 & ~n48023;
  assign n48795 = controllable_locked & ~n40216;
  assign n48796 = ~n43759 & ~n48795;
  assign n48797 = controllable_hgrant2 & ~n48796;
  assign n48798 = ~n7733 & n48797;
  assign n48799 = ~n46061 & ~n48798;
  assign n48800 = n7928 & ~n48799;
  assign n48801 = ~n48794 & ~n48800;
  assign n48802 = ~controllable_hgrant1 & ~n48801;
  assign n48803 = ~n48793 & ~n48802;
  assign n48804 = ~controllable_hgrant3 & ~n48803;
  assign n48805 = ~n48785 & ~n48804;
  assign n48806 = ~controllable_hgrant4 & ~n48805;
  assign n48807 = ~n48777 & ~n48806;
  assign n48808 = ~controllable_hgrant5 & ~n48807;
  assign n48809 = ~n48769 & ~n48808;
  assign n48810 = controllable_hmaster1 & ~n48809;
  assign n48811 = controllable_hmaster2 & ~n48809;
  assign n48812 = ~n46097 & ~n48811;
  assign n48813 = ~controllable_hmaster1 & ~n48812;
  assign n48814 = ~n48810 & ~n48813;
  assign n48815 = ~controllable_hgrant6 & ~n48814;
  assign n48816 = ~n45699 & ~n48815;
  assign n48817 = controllable_hmaster0 & ~n48816;
  assign n48818 = ~n47537 & ~n48811;
  assign n48819 = ~controllable_hmaster1 & ~n48818;
  assign n48820 = ~n48810 & ~n48819;
  assign n48821 = ~controllable_hgrant6 & ~n48820;
  assign n48822 = ~n45709 & ~n48821;
  assign n48823 = ~controllable_hmaster0 & ~n48822;
  assign n48824 = ~n48817 & ~n48823;
  assign n48825 = i_hlock8 & ~n48824;
  assign n48826 = ~n47570 & ~n48811;
  assign n48827 = ~controllable_hmaster1 & ~n48826;
  assign n48828 = ~n48810 & ~n48827;
  assign n48829 = ~controllable_hgrant6 & ~n48828;
  assign n48830 = ~n45721 & ~n48829;
  assign n48831 = ~controllable_hmaster0 & ~n48830;
  assign n48832 = ~n48817 & ~n48831;
  assign n48833 = ~i_hlock8 & ~n48832;
  assign n48834 = ~n48825 & ~n48833;
  assign n48835 = controllable_hmaster3 & ~n48834;
  assign n48836 = ~n8378 & ~n30284;
  assign n48837 = ~n43910 & ~n48836;
  assign n48838 = i_hlock5 & ~n48837;
  assign n48839 = ~n8378 & ~n30387;
  assign n48840 = ~n43910 & ~n48839;
  assign n48841 = ~i_hlock5 & ~n48840;
  assign n48842 = ~n48838 & ~n48841;
  assign n48843 = controllable_hgrant5 & ~n48842;
  assign n48844 = ~n8426 & ~n18589;
  assign n48845 = ~n43914 & ~n48844;
  assign n48846 = i_hlock4 & ~n48845;
  assign n48847 = ~n8426 & ~n18595;
  assign n48848 = ~n43914 & ~n48847;
  assign n48849 = ~i_hlock4 & ~n48848;
  assign n48850 = ~n48846 & ~n48849;
  assign n48851 = controllable_hgrant4 & ~n48850;
  assign n48852 = ~n8365 & ~n16513;
  assign n48853 = ~n43918 & ~n48852;
  assign n48854 = i_hlock3 & ~n48853;
  assign n48855 = ~n8365 & ~n16527;
  assign n48856 = ~n43922 & ~n48855;
  assign n48857 = ~i_hlock3 & ~n48856;
  assign n48858 = ~n48854 & ~n48857;
  assign n48859 = controllable_hgrant3 & ~n48858;
  assign n48860 = i_hlock3 & ~n46066;
  assign n48861 = ~i_hlock3 & ~n46088;
  assign n48862 = ~n48860 & ~n48861;
  assign n48863 = ~controllable_hgrant3 & ~n48862;
  assign n48864 = ~n48859 & ~n48863;
  assign n48865 = ~controllable_hgrant4 & ~n48864;
  assign n48866 = ~n48851 & ~n48865;
  assign n48867 = ~controllable_hgrant5 & ~n48866;
  assign n48868 = ~n48843 & ~n48867;
  assign n48869 = ~controllable_hmaster2 & ~n48868;
  assign n48870 = ~n47805 & ~n48869;
  assign n48871 = controllable_hmaster1 & ~n48870;
  assign n48872 = ~n8378 & ~n28970;
  assign n48873 = ~n43940 & ~n48872;
  assign n48874 = i_hlock5 & ~n48873;
  assign n48875 = ~n8378 & ~n28995;
  assign n48876 = ~n43944 & ~n48875;
  assign n48877 = ~i_hlock5 & ~n48876;
  assign n48878 = ~n48874 & ~n48877;
  assign n48879 = controllable_hgrant5 & ~n48878;
  assign n48880 = i_hlock5 & ~n47534;
  assign n48881 = ~i_hlock5 & ~n47567;
  assign n48882 = ~n48880 & ~n48881;
  assign n48883 = ~controllable_hgrant5 & ~n48882;
  assign n48884 = ~n48879 & ~n48883;
  assign n48885 = controllable_hmaster2 & ~n48884;
  assign n48886 = ~n8378 & ~n30297;
  assign n48887 = ~n43956 & ~n48886;
  assign n48888 = i_hlock5 & ~n48887;
  assign n48889 = ~n8378 & ~n30400;
  assign n48890 = ~n43956 & ~n48889;
  assign n48891 = ~i_hlock5 & ~n48890;
  assign n48892 = ~n48888 & ~n48891;
  assign n48893 = controllable_hgrant5 & ~n48892;
  assign n48894 = ~n8426 & ~n18617;
  assign n48895 = ~n43960 & ~n48894;
  assign n48896 = i_hlock4 & ~n48895;
  assign n48897 = ~n8426 & ~n18625;
  assign n48898 = ~n43960 & ~n48897;
  assign n48899 = ~i_hlock4 & ~n48898;
  assign n48900 = ~n48896 & ~n48899;
  assign n48901 = controllable_hgrant4 & ~n48900;
  assign n48902 = ~n8365 & ~n18615;
  assign n48903 = ~n43964 & ~n48902;
  assign n48904 = i_hlock3 & ~n48903;
  assign n48905 = ~n8365 & ~n18623;
  assign n48906 = ~n43964 & ~n48905;
  assign n48907 = ~i_hlock3 & ~n48906;
  assign n48908 = ~n48904 & ~n48907;
  assign n48909 = controllable_hgrant3 & ~n48908;
  assign n48910 = ~n8389 & ~n16511;
  assign n48911 = ~n43968 & ~n48910;
  assign n48912 = i_hlock1 & ~n48911;
  assign n48913 = ~n8389 & ~n16525;
  assign n48914 = ~n43972 & ~n48913;
  assign n48915 = ~i_hlock1 & ~n48914;
  assign n48916 = ~n48912 & ~n48915;
  assign n48917 = controllable_hgrant1 & ~n48916;
  assign n48918 = i_hlock1 & ~n46064;
  assign n48919 = ~i_hlock1 & ~n46086;
  assign n48920 = ~n48918 & ~n48919;
  assign n48921 = ~controllable_hgrant1 & ~n48920;
  assign n48922 = ~n48917 & ~n48921;
  assign n48923 = ~controllable_hgrant3 & ~n48922;
  assign n48924 = ~n48909 & ~n48923;
  assign n48925 = ~controllable_hgrant4 & ~n48924;
  assign n48926 = ~n48901 & ~n48925;
  assign n48927 = ~controllable_hgrant5 & ~n48926;
  assign n48928 = ~n48893 & ~n48927;
  assign n48929 = ~controllable_hmaster2 & ~n48928;
  assign n48930 = ~n48885 & ~n48929;
  assign n48931 = ~controllable_hmaster1 & ~n48930;
  assign n48932 = ~n48871 & ~n48931;
  assign n48933 = ~controllable_hgrant6 & ~n48932;
  assign n48934 = ~n45735 & ~n48933;
  assign n48935 = controllable_hmaster0 & ~n48934;
  assign n48936 = ~n8378 & ~n30309;
  assign n48937 = ~n44018 & ~n48936;
  assign n48938 = i_hlock5 & ~n48937;
  assign n48939 = ~n8378 & ~n30412;
  assign n48940 = ~n44018 & ~n48939;
  assign n48941 = ~i_hlock5 & ~n48940;
  assign n48942 = ~n48938 & ~n48941;
  assign n48943 = controllable_hgrant5 & ~n48942;
  assign n48944 = ~n8426 & ~n18643;
  assign n48945 = ~n44022 & ~n48944;
  assign n48946 = i_hlock4 & ~n48945;
  assign n48947 = ~n8426 & ~n18649;
  assign n48948 = ~n44022 & ~n48947;
  assign n48949 = ~i_hlock4 & ~n48948;
  assign n48950 = ~n48946 & ~n48949;
  assign n48951 = controllable_hgrant4 & ~n48950;
  assign n48952 = ~n8365 & ~n18641;
  assign n48953 = ~n44026 & ~n48952;
  assign n48954 = i_hlock3 & ~n48953;
  assign n48955 = ~n8365 & ~n18647;
  assign n48956 = ~n44026 & ~n48955;
  assign n48957 = ~i_hlock3 & ~n48956;
  assign n48958 = ~n48954 & ~n48957;
  assign n48959 = controllable_hgrant3 & ~n48958;
  assign n48960 = ~n8389 & ~n18639;
  assign n48961 = ~n44030 & ~n48960;
  assign n48962 = i_hlock1 & ~n48961;
  assign n48963 = ~n8389 & ~n18645;
  assign n48964 = ~n44030 & ~n48963;
  assign n48965 = ~i_hlock1 & ~n48964;
  assign n48966 = ~n48962 & ~n48965;
  assign n48967 = controllable_hgrant1 & ~n48966;
  assign n48968 = ~n7733 & n44035;
  assign n48969 = ~n42945 & ~n46049;
  assign n48970 = controllable_locked & ~n48969;
  assign n48971 = ~n43759 & ~n48970;
  assign n48972 = i_hlock2 & ~n48971;
  assign n48973 = ~n42945 & ~n44281;
  assign n48974 = controllable_locked & ~n48973;
  assign n48975 = ~n43759 & ~n48974;
  assign n48976 = ~i_hlock2 & ~n48975;
  assign n48977 = ~n48972 & ~n48976;
  assign n48978 = controllable_hgrant2 & ~n48977;
  assign n48979 = n7733 & n48978;
  assign n48980 = ~n48968 & ~n48979;
  assign n48981 = n7928 & ~n48980;
  assign n48982 = ~n42965 & ~n48981;
  assign n48983 = ~controllable_hgrant1 & ~n48982;
  assign n48984 = ~n48967 & ~n48983;
  assign n48985 = ~controllable_hgrant3 & ~n48984;
  assign n48986 = ~n48959 & ~n48985;
  assign n48987 = ~controllable_hgrant4 & ~n48986;
  assign n48988 = ~n48951 & ~n48987;
  assign n48989 = ~controllable_hgrant5 & ~n48988;
  assign n48990 = ~n48943 & ~n48989;
  assign n48991 = ~controllable_hmaster2 & ~n48990;
  assign n48992 = ~n47805 & ~n48991;
  assign n48993 = controllable_hmaster1 & ~n48992;
  assign n48994 = ~n8378 & ~n30319;
  assign n48995 = ~n44054 & ~n48994;
  assign n48996 = i_hlock5 & ~n48995;
  assign n48997 = ~n8378 & ~n30422;
  assign n48998 = ~n44054 & ~n48997;
  assign n48999 = ~i_hlock5 & ~n48998;
  assign n49000 = ~n48996 & ~n48999;
  assign n49001 = controllable_hgrant5 & ~n49000;
  assign n49002 = ~n8426 & ~n16515;
  assign n49003 = ~n44058 & ~n49002;
  assign n49004 = i_hlock4 & ~n49003;
  assign n49005 = ~n8426 & ~n16529;
  assign n49006 = ~n44062 & ~n49005;
  assign n49007 = ~i_hlock4 & ~n49006;
  assign n49008 = ~n49004 & ~n49007;
  assign n49009 = controllable_hgrant4 & ~n49008;
  assign n49010 = i_hlock4 & ~n46068;
  assign n49011 = ~i_hlock4 & ~n46090;
  assign n49012 = ~n49010 & ~n49011;
  assign n49013 = ~controllable_hgrant4 & ~n49012;
  assign n49014 = ~n49009 & ~n49013;
  assign n49015 = ~controllable_hgrant5 & ~n49014;
  assign n49016 = ~n49001 & ~n49015;
  assign n49017 = controllable_hmaster2 & ~n49016;
  assign n49018 = ~n8378 & ~n30324;
  assign n49019 = ~n44076 & ~n49018;
  assign n49020 = i_hlock5 & ~n49019;
  assign n49021 = ~n8378 & ~n30427;
  assign n49022 = ~n44076 & ~n49021;
  assign n49023 = ~i_hlock5 & ~n49022;
  assign n49024 = ~n49020 & ~n49023;
  assign n49025 = controllable_hgrant5 & ~n49024;
  assign n49026 = ~n8426 & ~n18671;
  assign n49027 = ~n44080 & ~n49026;
  assign n49028 = i_hlock4 & ~n49027;
  assign n49029 = ~n8426 & ~n18677;
  assign n49030 = ~n44080 & ~n49029;
  assign n49031 = ~i_hlock4 & ~n49030;
  assign n49032 = ~n49028 & ~n49031;
  assign n49033 = controllable_hgrant4 & ~n49032;
  assign n49034 = ~n8365 & ~n18669;
  assign n49035 = ~n44084 & ~n49034;
  assign n49036 = i_hlock3 & ~n49035;
  assign n49037 = ~n8365 & ~n18675;
  assign n49038 = ~n44084 & ~n49037;
  assign n49039 = ~i_hlock3 & ~n49038;
  assign n49040 = ~n49036 & ~n49039;
  assign n49041 = controllable_hgrant3 & ~n49040;
  assign n49042 = ~n8389 & ~n18667;
  assign n49043 = ~n44088 & ~n49042;
  assign n49044 = i_hlock1 & ~n49043;
  assign n49045 = ~n8389 & ~n18673;
  assign n49046 = ~n44088 & ~n49045;
  assign n49047 = ~i_hlock1 & ~n49046;
  assign n49048 = ~n49044 & ~n49047;
  assign n49049 = controllable_hgrant1 & ~n49048;
  assign n49050 = ~n8440 & ~n46063;
  assign n49051 = ~controllable_hgrant1 & ~n49050;
  assign n49052 = ~n49049 & ~n49051;
  assign n49053 = ~controllable_hgrant3 & ~n49052;
  assign n49054 = ~n49041 & ~n49053;
  assign n49055 = ~controllable_hgrant4 & ~n49054;
  assign n49056 = ~n49033 & ~n49055;
  assign n49057 = ~controllable_hgrant5 & ~n49056;
  assign n49058 = ~n49025 & ~n49057;
  assign n49059 = ~controllable_hmaster2 & ~n49058;
  assign n49060 = ~n49017 & ~n49059;
  assign n49061 = ~controllable_hmaster1 & ~n49060;
  assign n49062 = ~n48993 & ~n49061;
  assign n49063 = i_hlock6 & ~n49062;
  assign n49064 = ~n47824 & ~n48991;
  assign n49065 = controllable_hmaster1 & ~n49064;
  assign n49066 = ~n49061 & ~n49065;
  assign n49067 = ~i_hlock6 & ~n49066;
  assign n49068 = ~n49063 & ~n49067;
  assign n49069 = ~controllable_hgrant6 & ~n49068;
  assign n49070 = ~n45751 & ~n49069;
  assign n49071 = ~controllable_hmaster0 & ~n49070;
  assign n49072 = ~n48935 & ~n49071;
  assign n49073 = ~controllable_hmaster3 & ~n49072;
  assign n49074 = ~n48835 & ~n49073;
  assign n49075 = i_hlock7 & ~n49074;
  assign n49076 = ~n47824 & ~n48869;
  assign n49077 = controllable_hmaster1 & ~n49076;
  assign n49078 = ~n48931 & ~n49077;
  assign n49079 = ~controllable_hgrant6 & ~n49078;
  assign n49080 = ~n45775 & ~n49079;
  assign n49081 = controllable_hmaster0 & ~n49080;
  assign n49082 = ~n49071 & ~n49081;
  assign n49083 = ~controllable_hmaster3 & ~n49082;
  assign n49084 = ~n48835 & ~n49083;
  assign n49085 = ~i_hlock7 & ~n49084;
  assign n49086 = ~n49075 & ~n49085;
  assign n49087 = i_hbusreq7 & ~n49086;
  assign n49088 = i_hbusreq8 & ~n48834;
  assign n49089 = n8217 & ~n27641;
  assign n49090 = ~n8217 & ~n32065;
  assign n49091 = ~n49089 & ~n49090;
  assign n49092 = i_hlock6 & ~n49091;
  assign n49093 = ~n8217 & ~n32242;
  assign n49094 = ~n49089 & ~n49093;
  assign n49095 = ~i_hlock6 & ~n49094;
  assign n49096 = ~n49092 & ~n49095;
  assign n49097 = ~i_hbusreq6 & ~n49096;
  assign n49098 = ~n45785 & ~n49097;
  assign n49099 = controllable_hgrant6 & ~n49098;
  assign n49100 = i_hbusreq6 & ~n48814;
  assign n49101 = i_hbusreq5 & ~n48768;
  assign n49102 = n8378 & ~n14912;
  assign n49103 = ~n8378 & ~n32043;
  assign n49104 = ~n49102 & ~n49103;
  assign n49105 = i_hlock5 & ~n49104;
  assign n49106 = ~n8378 & ~n32220;
  assign n49107 = ~n49102 & ~n49106;
  assign n49108 = ~i_hlock5 & ~n49107;
  assign n49109 = ~n49105 & ~n49108;
  assign n49110 = ~i_hbusreq5 & ~n49109;
  assign n49111 = ~n49101 & ~n49110;
  assign n49112 = controllable_hgrant5 & ~n49111;
  assign n49113 = i_hbusreq5 & ~n48807;
  assign n49114 = i_hbusreq4 & ~n48776;
  assign n49115 = i_hbusreq9 & ~n48771;
  assign n49116 = n8426 & ~n14906;
  assign n49117 = ~n8426 & ~n21866;
  assign n49118 = ~n49116 & ~n49117;
  assign n49119 = ~i_hbusreq9 & ~n49118;
  assign n49120 = ~n49115 & ~n49119;
  assign n49121 = i_hlock4 & ~n49120;
  assign n49122 = i_hbusreq9 & ~n48774;
  assign n49123 = ~n8426 & ~n21884;
  assign n49124 = ~n49116 & ~n49123;
  assign n49125 = ~i_hbusreq9 & ~n49124;
  assign n49126 = ~n49122 & ~n49125;
  assign n49127 = ~i_hlock4 & ~n49126;
  assign n49128 = ~n49121 & ~n49127;
  assign n49129 = ~i_hbusreq4 & ~n49128;
  assign n49130 = ~n49114 & ~n49129;
  assign n49131 = controllable_hgrant4 & ~n49130;
  assign n49132 = i_hbusreq4 & ~n48805;
  assign n49133 = i_hbusreq9 & ~n48805;
  assign n49134 = i_hbusreq3 & ~n48784;
  assign n49135 = n8365 & ~n14902;
  assign n49136 = ~n8365 & ~n21862;
  assign n49137 = ~n49135 & ~n49136;
  assign n49138 = i_hlock3 & ~n49137;
  assign n49139 = ~n8365 & ~n21880;
  assign n49140 = ~n49135 & ~n49139;
  assign n49141 = ~i_hlock3 & ~n49140;
  assign n49142 = ~n49138 & ~n49141;
  assign n49143 = ~i_hbusreq3 & ~n49142;
  assign n49144 = ~n49134 & ~n49143;
  assign n49145 = controllable_hgrant3 & ~n49144;
  assign n49146 = i_hbusreq3 & ~n48803;
  assign n49147 = i_hbusreq1 & ~n48792;
  assign n49148 = n8389 & ~n14898;
  assign n49149 = ~n8389 & ~n21858;
  assign n49150 = ~n49148 & ~n49149;
  assign n49151 = i_hlock1 & ~n49150;
  assign n49152 = ~n8389 & ~n21876;
  assign n49153 = ~n49148 & ~n49152;
  assign n49154 = ~i_hlock1 & ~n49153;
  assign n49155 = ~n49151 & ~n49154;
  assign n49156 = ~i_hbusreq1 & ~n49155;
  assign n49157 = ~n49147 & ~n49156;
  assign n49158 = controllable_hgrant1 & ~n49157;
  assign n49159 = i_hbusreq1 & ~n48801;
  assign n49160 = ~n7928 & ~n48282;
  assign n49161 = i_hbusreq2 & ~n48796;
  assign n49162 = i_hbusreq0 & ~n48796;
  assign n49163 = ~controllable_locked & ~n44280;
  assign n49164 = ~n48795 & ~n49163;
  assign n49165 = i_hlock0 & ~n49164;
  assign n49166 = ~i_hlock0 & ~n48796;
  assign n49167 = ~n49165 & ~n49166;
  assign n49168 = ~i_hbusreq0 & ~n49167;
  assign n49169 = ~n49162 & ~n49168;
  assign n49170 = ~i_hbusreq2 & ~n49169;
  assign n49171 = ~n49161 & ~n49170;
  assign n49172 = controllable_hgrant2 & ~n49171;
  assign n49173 = ~i_hbusreq0 & ~n16519;
  assign n49174 = ~i_hbusreq0 & ~n49173;
  assign n49175 = ~i_hbusreq2 & ~n49174;
  assign n49176 = ~i_hbusreq2 & ~n49175;
  assign n49177 = ~controllable_hgrant2 & n49176;
  assign n49178 = ~n49172 & ~n49177;
  assign n49179 = ~n7733 & ~n49178;
  assign n49180 = ~n12781 & ~n39846;
  assign n49181 = controllable_hmastlock & ~n49180;
  assign n49182 = ~n42954 & ~n49181;
  assign n49183 = ~controllable_locked & ~n49182;
  assign n49184 = ~n46692 & ~n49183;
  assign n49185 = i_hlock0 & ~n49184;
  assign n49186 = ~n46695 & ~n49185;
  assign n49187 = ~i_hbusreq0 & ~n49186;
  assign n49188 = ~n46689 & ~n49187;
  assign n49189 = i_hlock2 & ~n49188;
  assign n49190 = ~n46700 & ~n49187;
  assign n49191 = ~i_hlock2 & ~n49190;
  assign n49192 = ~n49189 & ~n49191;
  assign n49193 = ~i_hbusreq2 & ~n49192;
  assign n49194 = ~n46688 & ~n49193;
  assign n49195 = controllable_hgrant2 & ~n49194;
  assign n49196 = ~n16645 & ~n49195;
  assign n49197 = n7733 & ~n49196;
  assign n49198 = ~n49179 & ~n49197;
  assign n49199 = n7928 & ~n49198;
  assign n49200 = ~n49160 & ~n49199;
  assign n49201 = ~i_hbusreq1 & ~n49200;
  assign n49202 = ~n49159 & ~n49201;
  assign n49203 = ~controllable_hgrant1 & ~n49202;
  assign n49204 = ~n49158 & ~n49203;
  assign n49205 = ~i_hbusreq3 & ~n49204;
  assign n49206 = ~n49146 & ~n49205;
  assign n49207 = ~controllable_hgrant3 & ~n49206;
  assign n49208 = ~n49145 & ~n49207;
  assign n49209 = ~i_hbusreq9 & ~n49208;
  assign n49210 = ~n49133 & ~n49209;
  assign n49211 = ~i_hbusreq4 & ~n49210;
  assign n49212 = ~n49132 & ~n49211;
  assign n49213 = ~controllable_hgrant4 & ~n49212;
  assign n49214 = ~n49131 & ~n49213;
  assign n49215 = ~i_hbusreq5 & ~n49214;
  assign n49216 = ~n49113 & ~n49215;
  assign n49217 = ~controllable_hgrant5 & ~n49216;
  assign n49218 = ~n49112 & ~n49217;
  assign n49219 = controllable_hmaster1 & ~n49218;
  assign n49220 = controllable_hmaster2 & ~n49218;
  assign n49221 = n8378 & ~n27633;
  assign n49222 = ~n8378 & ~n32057;
  assign n49223 = ~n49221 & ~n49222;
  assign n49224 = i_hlock5 & ~n49223;
  assign n49225 = ~n8378 & ~n32234;
  assign n49226 = ~n49221 & ~n49225;
  assign n49227 = ~i_hlock5 & ~n49226;
  assign n49228 = ~n49224 & ~n49227;
  assign n49229 = ~i_hbusreq5 & ~n49228;
  assign n49230 = ~n46623 & ~n49229;
  assign n49231 = controllable_hgrant5 & ~n49230;
  assign n49232 = n8426 & ~n14938;
  assign n49233 = ~n8426 & ~n21917;
  assign n49234 = ~n49232 & ~n49233;
  assign n49235 = i_hlock9 & ~n49234;
  assign n49236 = n8426 & ~n14969;
  assign n49237 = ~n8426 & ~n21961;
  assign n49238 = ~n49236 & ~n49237;
  assign n49239 = ~i_hlock9 & ~n49238;
  assign n49240 = ~n49235 & ~n49239;
  assign n49241 = ~i_hbusreq9 & ~n49240;
  assign n49242 = ~n46636 & ~n49241;
  assign n49243 = i_hlock4 & ~n49242;
  assign n49244 = ~n8426 & ~n21929;
  assign n49245 = ~n49232 & ~n49244;
  assign n49246 = i_hlock9 & ~n49245;
  assign n49247 = ~n8426 & ~n21971;
  assign n49248 = ~n49236 & ~n49247;
  assign n49249 = ~i_hlock9 & ~n49248;
  assign n49250 = ~n49246 & ~n49249;
  assign n49251 = ~i_hbusreq9 & ~n49250;
  assign n49252 = ~n46647 & ~n49251;
  assign n49253 = ~i_hlock4 & ~n49252;
  assign n49254 = ~n49243 & ~n49253;
  assign n49255 = ~i_hbusreq4 & ~n49254;
  assign n49256 = ~n46635 & ~n49255;
  assign n49257 = controllable_hgrant4 & ~n49256;
  assign n49258 = n8365 & ~n14934;
  assign n49259 = ~n8365 & ~n21913;
  assign n49260 = ~n49258 & ~n49259;
  assign n49261 = i_hlock3 & ~n49260;
  assign n49262 = ~n8365 & ~n21925;
  assign n49263 = ~n49258 & ~n49262;
  assign n49264 = ~i_hlock3 & ~n49263;
  assign n49265 = ~n49261 & ~n49264;
  assign n49266 = ~i_hbusreq3 & ~n49265;
  assign n49267 = ~n46664 & ~n49266;
  assign n49268 = controllable_hgrant3 & ~n49267;
  assign n49269 = n8389 & ~n14930;
  assign n49270 = ~n8389 & ~n21909;
  assign n49271 = ~n49269 & ~n49270;
  assign n49272 = i_hlock1 & ~n49271;
  assign n49273 = ~n8389 & ~n21921;
  assign n49274 = ~n49269 & ~n49273;
  assign n49275 = ~i_hlock1 & ~n49274;
  assign n49276 = ~n49272 & ~n49275;
  assign n49277 = ~i_hbusreq1 & ~n49276;
  assign n49278 = ~n46676 & ~n49277;
  assign n49279 = controllable_hgrant1 & ~n49278;
  assign n49280 = controllable_locked & controllable_ndecide;
  assign n49281 = ~n17556 & ~n49280;
  assign n49282 = i_hlock0 & ~n49281;
  assign n49283 = ~n44269 & ~n49282;
  assign n49284 = ~i_hbusreq0 & ~n49283;
  assign n49285 = ~i_hbusreq0 & ~n49284;
  assign n49286 = ~i_hbusreq2 & ~n49285;
  assign n49287 = ~i_hbusreq2 & ~n49286;
  assign n49288 = ~controllable_hgrant2 & n49287;
  assign n49289 = ~n44191 & ~n49288;
  assign n49290 = ~n7733 & ~n49289;
  assign n49291 = ~n16638 & ~n44269;
  assign n49292 = ~i_hbusreq0 & ~n49291;
  assign n49293 = ~i_hbusreq0 & ~n49292;
  assign n49294 = ~i_hbusreq2 & ~n49293;
  assign n49295 = ~i_hbusreq2 & ~n49294;
  assign n49296 = ~controllable_hgrant2 & n49295;
  assign n49297 = ~n49195 & ~n49296;
  assign n49298 = n7733 & ~n49297;
  assign n49299 = ~n49290 & ~n49298;
  assign n49300 = n7928 & ~n49299;
  assign n49301 = ~n8265 & ~n49300;
  assign n49302 = ~i_hbusreq1 & ~n49301;
  assign n49303 = ~n46687 & ~n49302;
  assign n49304 = ~controllable_hgrant1 & ~n49303;
  assign n49305 = ~n49279 & ~n49304;
  assign n49306 = ~i_hbusreq3 & ~n49305;
  assign n49307 = ~n46675 & ~n49306;
  assign n49308 = ~controllable_hgrant3 & ~n49307;
  assign n49309 = ~n49268 & ~n49308;
  assign n49310 = i_hlock9 & ~n49309;
  assign n49311 = n8365 & ~n14965;
  assign n49312 = ~n8365 & ~n21957;
  assign n49313 = ~n49311 & ~n49312;
  assign n49314 = i_hlock3 & ~n49313;
  assign n49315 = ~n8365 & ~n21967;
  assign n49316 = ~n49311 & ~n49315;
  assign n49317 = ~i_hlock3 & ~n49316;
  assign n49318 = ~n49314 & ~n49317;
  assign n49319 = ~i_hbusreq3 & ~n49318;
  assign n49320 = ~n46728 & ~n49319;
  assign n49321 = controllable_hgrant3 & ~n49320;
  assign n49322 = n8389 & ~n14961;
  assign n49323 = ~n8389 & ~n21953;
  assign n49324 = ~n49322 & ~n49323;
  assign n49325 = i_hlock1 & ~n49324;
  assign n49326 = ~n8389 & ~n21963;
  assign n49327 = ~n49322 & ~n49326;
  assign n49328 = ~i_hlock1 & ~n49327;
  assign n49329 = ~n49325 & ~n49328;
  assign n49330 = ~i_hbusreq1 & ~n49329;
  assign n49331 = ~n46740 & ~n49330;
  assign n49332 = controllable_hgrant1 & ~n49331;
  assign n49333 = ~n8297 & ~n49300;
  assign n49334 = ~i_hbusreq1 & ~n49333;
  assign n49335 = ~n46751 & ~n49334;
  assign n49336 = ~controllable_hgrant1 & ~n49335;
  assign n49337 = ~n49332 & ~n49336;
  assign n49338 = ~i_hbusreq3 & ~n49337;
  assign n49339 = ~n46739 & ~n49338;
  assign n49340 = ~controllable_hgrant3 & ~n49339;
  assign n49341 = ~n49321 & ~n49340;
  assign n49342 = ~i_hlock9 & ~n49341;
  assign n49343 = ~n49310 & ~n49342;
  assign n49344 = ~i_hbusreq9 & ~n49343;
  assign n49345 = ~n46663 & ~n49344;
  assign n49346 = ~i_hbusreq4 & ~n49345;
  assign n49347 = ~n46662 & ~n49346;
  assign n49348 = ~controllable_hgrant4 & ~n49347;
  assign n49349 = ~n49257 & ~n49348;
  assign n49350 = ~i_hbusreq5 & ~n49349;
  assign n49351 = ~n46634 & ~n49350;
  assign n49352 = ~controllable_hgrant5 & ~n49351;
  assign n49353 = ~n49231 & ~n49352;
  assign n49354 = ~controllable_hmaster2 & ~n49353;
  assign n49355 = ~n49220 & ~n49354;
  assign n49356 = ~controllable_hmaster1 & ~n49355;
  assign n49357 = ~n49219 & ~n49356;
  assign n49358 = ~i_hbusreq6 & ~n49357;
  assign n49359 = ~n49100 & ~n49358;
  assign n49360 = ~controllable_hgrant6 & ~n49359;
  assign n49361 = ~n49099 & ~n49360;
  assign n49362 = controllable_hmaster0 & ~n49361;
  assign n49363 = n8217 & ~n14952;
  assign n49364 = ~n8217 & ~n32084;
  assign n49365 = ~n49363 & ~n49364;
  assign n49366 = i_hlock6 & ~n49365;
  assign n49367 = ~n8217 & ~n32261;
  assign n49368 = ~n49363 & ~n49367;
  assign n49369 = ~i_hlock6 & ~n49368;
  assign n49370 = ~n49366 & ~n49369;
  assign n49371 = ~i_hbusreq6 & ~n49370;
  assign n49372 = ~n45799 & ~n49371;
  assign n49373 = controllable_hgrant6 & ~n49372;
  assign n49374 = i_hbusreq6 & ~n48820;
  assign n49375 = n8378 & ~n14944;
  assign n49376 = ~n8378 & ~n32076;
  assign n49377 = ~n49375 & ~n49376;
  assign n49378 = i_hlock5 & ~n49377;
  assign n49379 = ~n8378 & ~n32253;
  assign n49380 = ~n49375 & ~n49379;
  assign n49381 = ~i_hlock5 & ~n49380;
  assign n49382 = ~n49378 & ~n49381;
  assign n49383 = ~i_hbusreq5 & ~n49382;
  assign n49384 = ~n47667 & ~n49383;
  assign n49385 = controllable_hgrant5 & ~n49384;
  assign n49386 = ~i_hbusreq9 & ~n49234;
  assign n49387 = ~n47680 & ~n49386;
  assign n49388 = i_hlock4 & ~n49387;
  assign n49389 = ~i_hbusreq9 & ~n49245;
  assign n49390 = ~n47684 & ~n49389;
  assign n49391 = ~i_hlock4 & ~n49390;
  assign n49392 = ~n49388 & ~n49391;
  assign n49393 = ~i_hbusreq4 & ~n49392;
  assign n49394 = ~n47679 & ~n49393;
  assign n49395 = controllable_hgrant4 & ~n49394;
  assign n49396 = ~i_hbusreq9 & ~n49309;
  assign n49397 = ~n47693 & ~n49396;
  assign n49398 = ~i_hbusreq4 & ~n49397;
  assign n49399 = ~n47692 & ~n49398;
  assign n49400 = ~controllable_hgrant4 & ~n49399;
  assign n49401 = ~n49395 & ~n49400;
  assign n49402 = ~i_hbusreq5 & ~n49401;
  assign n49403 = ~n47678 & ~n49402;
  assign n49404 = ~controllable_hgrant5 & ~n49403;
  assign n49405 = ~n49385 & ~n49404;
  assign n49406 = ~controllable_hmaster2 & ~n49405;
  assign n49407 = ~n49220 & ~n49406;
  assign n49408 = ~controllable_hmaster1 & ~n49407;
  assign n49409 = ~n49219 & ~n49408;
  assign n49410 = ~i_hbusreq6 & ~n49409;
  assign n49411 = ~n49374 & ~n49410;
  assign n49412 = ~controllable_hgrant6 & ~n49411;
  assign n49413 = ~n49373 & ~n49412;
  assign n49414 = ~controllable_hmaster0 & ~n49413;
  assign n49415 = ~n49362 & ~n49414;
  assign n49416 = i_hlock8 & ~n49415;
  assign n49417 = n8217 & ~n14983;
  assign n49418 = ~n8217 & ~n32105;
  assign n49419 = ~n49417 & ~n49418;
  assign n49420 = i_hlock6 & ~n49419;
  assign n49421 = ~n8217 & ~n32282;
  assign n49422 = ~n49417 & ~n49421;
  assign n49423 = ~i_hlock6 & ~n49422;
  assign n49424 = ~n49420 & ~n49423;
  assign n49425 = ~i_hbusreq6 & ~n49424;
  assign n49426 = ~n45815 & ~n49425;
  assign n49427 = controllable_hgrant6 & ~n49426;
  assign n49428 = i_hbusreq6 & ~n48828;
  assign n49429 = n8378 & ~n14975;
  assign n49430 = ~n8378 & ~n32097;
  assign n49431 = ~n49429 & ~n49430;
  assign n49432 = i_hlock5 & ~n49431;
  assign n49433 = ~n8378 & ~n32274;
  assign n49434 = ~n49429 & ~n49433;
  assign n49435 = ~i_hlock5 & ~n49434;
  assign n49436 = ~n49432 & ~n49435;
  assign n49437 = ~i_hbusreq5 & ~n49436;
  assign n49438 = ~n47727 & ~n49437;
  assign n49439 = controllable_hgrant5 & ~n49438;
  assign n49440 = ~i_hbusreq9 & ~n49238;
  assign n49441 = ~n47740 & ~n49440;
  assign n49442 = i_hlock4 & ~n49441;
  assign n49443 = ~i_hbusreq9 & ~n49248;
  assign n49444 = ~n47744 & ~n49443;
  assign n49445 = ~i_hlock4 & ~n49444;
  assign n49446 = ~n49442 & ~n49445;
  assign n49447 = ~i_hbusreq4 & ~n49446;
  assign n49448 = ~n47739 & ~n49447;
  assign n49449 = controllable_hgrant4 & ~n49448;
  assign n49450 = ~i_hbusreq9 & ~n49341;
  assign n49451 = ~n47753 & ~n49450;
  assign n49452 = ~i_hbusreq4 & ~n49451;
  assign n49453 = ~n47752 & ~n49452;
  assign n49454 = ~controllable_hgrant4 & ~n49453;
  assign n49455 = ~n49449 & ~n49454;
  assign n49456 = ~i_hbusreq5 & ~n49455;
  assign n49457 = ~n47738 & ~n49456;
  assign n49458 = ~controllable_hgrant5 & ~n49457;
  assign n49459 = ~n49439 & ~n49458;
  assign n49460 = ~controllable_hmaster2 & ~n49459;
  assign n49461 = ~n49220 & ~n49460;
  assign n49462 = ~controllable_hmaster1 & ~n49461;
  assign n49463 = ~n49219 & ~n49462;
  assign n49464 = ~i_hbusreq6 & ~n49463;
  assign n49465 = ~n49428 & ~n49464;
  assign n49466 = ~controllable_hgrant6 & ~n49465;
  assign n49467 = ~n49427 & ~n49466;
  assign n49468 = ~controllable_hmaster0 & ~n49467;
  assign n49469 = ~n49362 & ~n49468;
  assign n49470 = ~i_hlock8 & ~n49469;
  assign n49471 = ~n49416 & ~n49470;
  assign n49472 = ~i_hbusreq8 & ~n49471;
  assign n49473 = ~n49088 & ~n49472;
  assign n49474 = controllable_hmaster3 & ~n49473;
  assign n49475 = i_hbusreq8 & ~n49072;
  assign n49476 = n8217 & ~n15057;
  assign n49477 = ~n8217 & ~n37802;
  assign n49478 = ~n49476 & ~n49477;
  assign n49479 = i_hlock6 & ~n49478;
  assign n49480 = ~n8217 & ~n37812;
  assign n49481 = ~n49476 & ~n49480;
  assign n49482 = ~i_hlock6 & ~n49481;
  assign n49483 = ~n49479 & ~n49482;
  assign n49484 = ~i_hbusreq6 & ~n49483;
  assign n49485 = ~n45836 & ~n49484;
  assign n49486 = controllable_hgrant6 & ~n49485;
  assign n49487 = i_hbusreq6 & ~n48932;
  assign n49488 = controllable_hmaster2 & ~n49405;
  assign n49489 = i_hbusreq5 & ~n48842;
  assign n49490 = n8378 & ~n15012;
  assign n49491 = ~n8378 & ~n32122;
  assign n49492 = ~n49490 & ~n49491;
  assign n49493 = i_hlock5 & ~n49492;
  assign n49494 = ~n8378 & ~n32299;
  assign n49495 = ~n49490 & ~n49494;
  assign n49496 = ~i_hlock5 & ~n49495;
  assign n49497 = ~n49493 & ~n49496;
  assign n49498 = ~i_hbusreq5 & ~n49497;
  assign n49499 = ~n49489 & ~n49498;
  assign n49500 = controllable_hgrant5 & ~n49499;
  assign n49501 = i_hbusreq5 & ~n48866;
  assign n49502 = i_hbusreq4 & ~n48850;
  assign n49503 = i_hbusreq9 & ~n48845;
  assign n49504 = n8426 & ~n15006;
  assign n49505 = ~n8426 & ~n22006;
  assign n49506 = ~n49504 & ~n49505;
  assign n49507 = ~i_hbusreq9 & ~n49506;
  assign n49508 = ~n49503 & ~n49507;
  assign n49509 = i_hlock4 & ~n49508;
  assign n49510 = i_hbusreq9 & ~n48848;
  assign n49511 = ~n8426 & ~n22014;
  assign n49512 = ~n49504 & ~n49511;
  assign n49513 = ~i_hbusreq9 & ~n49512;
  assign n49514 = ~n49510 & ~n49513;
  assign n49515 = ~i_hlock4 & ~n49514;
  assign n49516 = ~n49509 & ~n49515;
  assign n49517 = ~i_hbusreq4 & ~n49516;
  assign n49518 = ~n49502 & ~n49517;
  assign n49519 = controllable_hgrant4 & ~n49518;
  assign n49520 = i_hbusreq4 & ~n48864;
  assign n49521 = i_hbusreq9 & ~n48864;
  assign n49522 = i_hbusreq3 & ~n48858;
  assign n49523 = n8365 & ~n12913;
  assign n49524 = ~n8365 & ~n16654;
  assign n49525 = ~n49523 & ~n49524;
  assign n49526 = i_hlock3 & ~n49525;
  assign n49527 = n8365 & ~n12925;
  assign n49528 = ~n8365 & ~n16676;
  assign n49529 = ~n49527 & ~n49528;
  assign n49530 = ~i_hlock3 & ~n49529;
  assign n49531 = ~n49526 & ~n49530;
  assign n49532 = ~i_hbusreq3 & ~n49531;
  assign n49533 = ~n49522 & ~n49532;
  assign n49534 = controllable_hgrant3 & ~n49533;
  assign n49535 = i_hbusreq3 & ~n48862;
  assign n49536 = i_hlock3 & ~n49305;
  assign n49537 = ~i_hlock3 & ~n49337;
  assign n49538 = ~n49536 & ~n49537;
  assign n49539 = ~i_hbusreq3 & ~n49538;
  assign n49540 = ~n49535 & ~n49539;
  assign n49541 = ~controllable_hgrant3 & ~n49540;
  assign n49542 = ~n49534 & ~n49541;
  assign n49543 = ~i_hbusreq9 & ~n49542;
  assign n49544 = ~n49521 & ~n49543;
  assign n49545 = ~i_hbusreq4 & ~n49544;
  assign n49546 = ~n49520 & ~n49545;
  assign n49547 = ~controllable_hgrant4 & ~n49546;
  assign n49548 = ~n49519 & ~n49547;
  assign n49549 = ~i_hbusreq5 & ~n49548;
  assign n49550 = ~n49501 & ~n49549;
  assign n49551 = ~controllable_hgrant5 & ~n49550;
  assign n49552 = ~n49500 & ~n49551;
  assign n49553 = ~controllable_hmaster2 & ~n49552;
  assign n49554 = ~n49488 & ~n49553;
  assign n49555 = controllable_hmaster1 & ~n49554;
  assign n49556 = i_hbusreq5 & ~n48878;
  assign n49557 = n8378 & ~n26778;
  assign n49558 = ~n8378 & ~n29046;
  assign n49559 = ~n49557 & ~n49558;
  assign n49560 = i_hlock5 & ~n49559;
  assign n49561 = n8378 & ~n26809;
  assign n49562 = ~n8378 & ~n29101;
  assign n49563 = ~n49561 & ~n49562;
  assign n49564 = ~i_hlock5 & ~n49563;
  assign n49565 = ~n49560 & ~n49564;
  assign n49566 = ~i_hbusreq5 & ~n49565;
  assign n49567 = ~n49556 & ~n49566;
  assign n49568 = controllable_hgrant5 & ~n49567;
  assign n49569 = i_hbusreq5 & ~n48882;
  assign n49570 = i_hlock5 & ~n49401;
  assign n49571 = ~i_hlock5 & ~n49455;
  assign n49572 = ~n49570 & ~n49571;
  assign n49573 = ~i_hbusreq5 & ~n49572;
  assign n49574 = ~n49569 & ~n49573;
  assign n49575 = ~controllable_hgrant5 & ~n49574;
  assign n49576 = ~n49568 & ~n49575;
  assign n49577 = controllable_hmaster2 & ~n49576;
  assign n49578 = i_hbusreq5 & ~n48892;
  assign n49579 = n8378 & ~n15049;
  assign n49580 = ~n8378 & ~n32143;
  assign n49581 = ~n49579 & ~n49580;
  assign n49582 = i_hlock5 & ~n49581;
  assign n49583 = ~n8378 & ~n32320;
  assign n49584 = ~n49579 & ~n49583;
  assign n49585 = ~i_hlock5 & ~n49584;
  assign n49586 = ~n49582 & ~n49585;
  assign n49587 = ~i_hbusreq5 & ~n49586;
  assign n49588 = ~n49578 & ~n49587;
  assign n49589 = controllable_hgrant5 & ~n49588;
  assign n49590 = i_hbusreq5 & ~n48926;
  assign n49591 = i_hbusreq4 & ~n48900;
  assign n49592 = i_hbusreq9 & ~n48895;
  assign n49593 = n8426 & ~n15043;
  assign n49594 = ~n8426 & ~n22048;
  assign n49595 = ~n49593 & ~n49594;
  assign n49596 = ~i_hbusreq9 & ~n49595;
  assign n49597 = ~n49592 & ~n49596;
  assign n49598 = i_hlock4 & ~n49597;
  assign n49599 = i_hbusreq9 & ~n48898;
  assign n49600 = ~n8426 & ~n22060;
  assign n49601 = ~n49593 & ~n49600;
  assign n49602 = ~i_hbusreq9 & ~n49601;
  assign n49603 = ~n49599 & ~n49602;
  assign n49604 = ~i_hlock4 & ~n49603;
  assign n49605 = ~n49598 & ~n49604;
  assign n49606 = ~i_hbusreq4 & ~n49605;
  assign n49607 = ~n49591 & ~n49606;
  assign n49608 = controllable_hgrant4 & ~n49607;
  assign n49609 = i_hbusreq4 & ~n48924;
  assign n49610 = i_hbusreq9 & ~n48924;
  assign n49611 = i_hbusreq3 & ~n48908;
  assign n49612 = n8365 & ~n15039;
  assign n49613 = ~n8365 & ~n22044;
  assign n49614 = ~n49612 & ~n49613;
  assign n49615 = i_hlock3 & ~n49614;
  assign n49616 = ~n8365 & ~n22056;
  assign n49617 = ~n49612 & ~n49616;
  assign n49618 = ~i_hlock3 & ~n49617;
  assign n49619 = ~n49615 & ~n49618;
  assign n49620 = ~i_hbusreq3 & ~n49619;
  assign n49621 = ~n49611 & ~n49620;
  assign n49622 = controllable_hgrant3 & ~n49621;
  assign n49623 = i_hbusreq3 & ~n48922;
  assign n49624 = i_hbusreq1 & ~n48916;
  assign n49625 = n8389 & ~n12909;
  assign n49626 = ~n8389 & ~n16650;
  assign n49627 = ~n49625 & ~n49626;
  assign n49628 = i_hlock1 & ~n49627;
  assign n49629 = n8389 & ~n12921;
  assign n49630 = ~n8389 & ~n16672;
  assign n49631 = ~n49629 & ~n49630;
  assign n49632 = ~i_hlock1 & ~n49631;
  assign n49633 = ~n49628 & ~n49632;
  assign n49634 = ~i_hbusreq1 & ~n49633;
  assign n49635 = ~n49624 & ~n49634;
  assign n49636 = controllable_hgrant1 & ~n49635;
  assign n49637 = i_hbusreq1 & ~n48920;
  assign n49638 = i_hlock1 & ~n49301;
  assign n49639 = ~i_hlock1 & ~n49333;
  assign n49640 = ~n49638 & ~n49639;
  assign n49641 = ~i_hbusreq1 & ~n49640;
  assign n49642 = ~n49637 & ~n49641;
  assign n49643 = ~controllable_hgrant1 & ~n49642;
  assign n49644 = ~n49636 & ~n49643;
  assign n49645 = ~i_hbusreq3 & ~n49644;
  assign n49646 = ~n49623 & ~n49645;
  assign n49647 = ~controllable_hgrant3 & ~n49646;
  assign n49648 = ~n49622 & ~n49647;
  assign n49649 = ~i_hbusreq9 & ~n49648;
  assign n49650 = ~n49610 & ~n49649;
  assign n49651 = ~i_hbusreq4 & ~n49650;
  assign n49652 = ~n49609 & ~n49651;
  assign n49653 = ~controllable_hgrant4 & ~n49652;
  assign n49654 = ~n49608 & ~n49653;
  assign n49655 = ~i_hbusreq5 & ~n49654;
  assign n49656 = ~n49590 & ~n49655;
  assign n49657 = ~controllable_hgrant5 & ~n49656;
  assign n49658 = ~n49589 & ~n49657;
  assign n49659 = ~controllable_hmaster2 & ~n49658;
  assign n49660 = ~n49577 & ~n49659;
  assign n49661 = ~controllable_hmaster1 & ~n49660;
  assign n49662 = ~n49555 & ~n49661;
  assign n49663 = ~i_hbusreq6 & ~n49662;
  assign n49664 = ~n49487 & ~n49663;
  assign n49665 = ~controllable_hgrant6 & ~n49664;
  assign n49666 = ~n49486 & ~n49665;
  assign n49667 = controllable_hmaster0 & ~n49666;
  assign n49668 = ~n15087 & ~n26783;
  assign n49669 = controllable_hmaster1 & ~n49668;
  assign n49670 = ~n15132 & ~n49669;
  assign n49671 = n8217 & ~n49670;
  assign n49672 = ~n29051 & ~n32168;
  assign n49673 = controllable_hmaster1 & ~n49672;
  assign n49674 = ~n32195 & ~n49673;
  assign n49675 = ~n8217 & ~n49674;
  assign n49676 = ~n49671 & ~n49675;
  assign n49677 = i_hlock6 & ~n49676;
  assign n49678 = ~n15087 & ~n26814;
  assign n49679 = controllable_hmaster1 & ~n49678;
  assign n49680 = ~n15132 & ~n49679;
  assign n49681 = n8217 & ~n49680;
  assign n49682 = ~n29106 & ~n32345;
  assign n49683 = controllable_hmaster1 & ~n49682;
  assign n49684 = ~n32372 & ~n49683;
  assign n49685 = ~n8217 & ~n49684;
  assign n49686 = ~n49681 & ~n49685;
  assign n49687 = ~i_hlock6 & ~n49686;
  assign n49688 = ~n49677 & ~n49687;
  assign n49689 = ~i_hbusreq6 & ~n49688;
  assign n49690 = ~n45850 & ~n49689;
  assign n49691 = controllable_hgrant6 & ~n49690;
  assign n49692 = i_hbusreq6 & ~n49068;
  assign n49693 = i_hbusreq5 & ~n48942;
  assign n49694 = n8378 & ~n15082;
  assign n49695 = ~n8378 & ~n32163;
  assign n49696 = ~n49694 & ~n49695;
  assign n49697 = i_hlock5 & ~n49696;
  assign n49698 = ~n8378 & ~n32340;
  assign n49699 = ~n49694 & ~n49698;
  assign n49700 = ~i_hlock5 & ~n49699;
  assign n49701 = ~n49697 & ~n49700;
  assign n49702 = ~i_hbusreq5 & ~n49701;
  assign n49703 = ~n49693 & ~n49702;
  assign n49704 = controllable_hgrant5 & ~n49703;
  assign n49705 = i_hbusreq5 & ~n48988;
  assign n49706 = i_hbusreq4 & ~n48950;
  assign n49707 = i_hbusreq9 & ~n48945;
  assign n49708 = n8426 & ~n15076;
  assign n49709 = ~n8426 & ~n22090;
  assign n49710 = ~n49708 & ~n49709;
  assign n49711 = ~i_hbusreq9 & ~n49710;
  assign n49712 = ~n49707 & ~n49711;
  assign n49713 = i_hlock4 & ~n49712;
  assign n49714 = i_hbusreq9 & ~n48948;
  assign n49715 = ~n8426 & ~n22100;
  assign n49716 = ~n49708 & ~n49715;
  assign n49717 = ~i_hbusreq9 & ~n49716;
  assign n49718 = ~n49714 & ~n49717;
  assign n49719 = ~i_hlock4 & ~n49718;
  assign n49720 = ~n49713 & ~n49719;
  assign n49721 = ~i_hbusreq4 & ~n49720;
  assign n49722 = ~n49706 & ~n49721;
  assign n49723 = controllable_hgrant4 & ~n49722;
  assign n49724 = i_hbusreq4 & ~n48986;
  assign n49725 = i_hbusreq9 & ~n48986;
  assign n49726 = i_hbusreq3 & ~n48958;
  assign n49727 = n8365 & ~n15072;
  assign n49728 = ~n8365 & ~n22086;
  assign n49729 = ~n49727 & ~n49728;
  assign n49730 = i_hlock3 & ~n49729;
  assign n49731 = ~n8365 & ~n22096;
  assign n49732 = ~n49727 & ~n49731;
  assign n49733 = ~i_hlock3 & ~n49732;
  assign n49734 = ~n49730 & ~n49733;
  assign n49735 = ~i_hbusreq3 & ~n49734;
  assign n49736 = ~n49726 & ~n49735;
  assign n49737 = controllable_hgrant3 & ~n49736;
  assign n49738 = i_hbusreq3 & ~n48984;
  assign n49739 = i_hbusreq1 & ~n48966;
  assign n49740 = n8389 & ~n15068;
  assign n49741 = ~n8389 & ~n22082;
  assign n49742 = ~n49740 & ~n49741;
  assign n49743 = i_hlock1 & ~n49742;
  assign n49744 = ~n8389 & ~n22092;
  assign n49745 = ~n49740 & ~n49744;
  assign n49746 = ~i_hlock1 & ~n49745;
  assign n49747 = ~n49743 & ~n49746;
  assign n49748 = ~i_hbusreq1 & ~n49747;
  assign n49749 = ~n49739 & ~n49748;
  assign n49750 = controllable_hgrant1 & ~n49749;
  assign n49751 = i_hbusreq1 & ~n48982;
  assign n49752 = ~n44750 & ~n49288;
  assign n49753 = ~n7733 & ~n49752;
  assign n49754 = i_hbusreq2 & ~n48977;
  assign n49755 = i_hbusreq0 & ~n48971;
  assign n49756 = controllable_locked & ~n44282;
  assign n49757 = ~n49183 & ~n49756;
  assign n49758 = i_hlock0 & ~n49757;
  assign n49759 = ~i_hlock0 & ~n48975;
  assign n49760 = ~n49758 & ~n49759;
  assign n49761 = ~i_hbusreq0 & ~n49760;
  assign n49762 = ~n49755 & ~n49761;
  assign n49763 = i_hlock2 & ~n49762;
  assign n49764 = i_hbusreq0 & ~n48975;
  assign n49765 = ~n49761 & ~n49764;
  assign n49766 = ~i_hlock2 & ~n49765;
  assign n49767 = ~n49763 & ~n49766;
  assign n49768 = ~i_hbusreq2 & ~n49767;
  assign n49769 = ~n49754 & ~n49768;
  assign n49770 = controllable_hgrant2 & ~n49769;
  assign n49771 = ~n49296 & ~n49770;
  assign n49772 = n7733 & ~n49771;
  assign n49773 = ~n49753 & ~n49772;
  assign n49774 = n7928 & ~n49773;
  assign n49775 = ~n43545 & ~n49774;
  assign n49776 = ~i_hbusreq1 & ~n49775;
  assign n49777 = ~n49751 & ~n49776;
  assign n49778 = ~controllable_hgrant1 & ~n49777;
  assign n49779 = ~n49750 & ~n49778;
  assign n49780 = ~i_hbusreq3 & ~n49779;
  assign n49781 = ~n49738 & ~n49780;
  assign n49782 = ~controllable_hgrant3 & ~n49781;
  assign n49783 = ~n49737 & ~n49782;
  assign n49784 = ~i_hbusreq9 & ~n49783;
  assign n49785 = ~n49725 & ~n49784;
  assign n49786 = ~i_hbusreq4 & ~n49785;
  assign n49787 = ~n49724 & ~n49786;
  assign n49788 = ~controllable_hgrant4 & ~n49787;
  assign n49789 = ~n49723 & ~n49788;
  assign n49790 = ~i_hbusreq5 & ~n49789;
  assign n49791 = ~n49705 & ~n49790;
  assign n49792 = ~controllable_hgrant5 & ~n49791;
  assign n49793 = ~n49704 & ~n49792;
  assign n49794 = ~controllable_hmaster2 & ~n49793;
  assign n49795 = ~n49488 & ~n49794;
  assign n49796 = controllable_hmaster1 & ~n49795;
  assign n49797 = i_hbusreq5 & ~n49000;
  assign n49798 = n8378 & ~n15098;
  assign n49799 = ~n8378 & ~n32177;
  assign n49800 = ~n49798 & ~n49799;
  assign n49801 = i_hlock5 & ~n49800;
  assign n49802 = ~n8378 & ~n32354;
  assign n49803 = ~n49798 & ~n49802;
  assign n49804 = ~i_hlock5 & ~n49803;
  assign n49805 = ~n49801 & ~n49804;
  assign n49806 = ~i_hbusreq5 & ~n49805;
  assign n49807 = ~n49797 & ~n49806;
  assign n49808 = controllable_hgrant5 & ~n49807;
  assign n49809 = i_hbusreq5 & ~n49014;
  assign n49810 = i_hbusreq4 & ~n49008;
  assign n49811 = i_hbusreq9 & ~n49003;
  assign n49812 = n8426 & ~n12917;
  assign n49813 = ~n8426 & ~n16658;
  assign n49814 = ~n49812 & ~n49813;
  assign n49815 = ~i_hbusreq9 & ~n49814;
  assign n49816 = ~n49811 & ~n49815;
  assign n49817 = i_hlock4 & ~n49816;
  assign n49818 = i_hbusreq9 & ~n49006;
  assign n49819 = n8426 & ~n12929;
  assign n49820 = ~n8426 & ~n16680;
  assign n49821 = ~n49819 & ~n49820;
  assign n49822 = ~i_hbusreq9 & ~n49821;
  assign n49823 = ~n49818 & ~n49822;
  assign n49824 = ~i_hlock4 & ~n49823;
  assign n49825 = ~n49817 & ~n49824;
  assign n49826 = ~i_hbusreq4 & ~n49825;
  assign n49827 = ~n49810 & ~n49826;
  assign n49828 = controllable_hgrant4 & ~n49827;
  assign n49829 = i_hbusreq4 & ~n49012;
  assign n49830 = i_hlock4 & ~n49397;
  assign n49831 = ~i_hlock4 & ~n49451;
  assign n49832 = ~n49830 & ~n49831;
  assign n49833 = ~i_hbusreq4 & ~n49832;
  assign n49834 = ~n49829 & ~n49833;
  assign n49835 = ~controllable_hgrant4 & ~n49834;
  assign n49836 = ~n49828 & ~n49835;
  assign n49837 = ~i_hbusreq5 & ~n49836;
  assign n49838 = ~n49809 & ~n49837;
  assign n49839 = ~controllable_hgrant5 & ~n49838;
  assign n49840 = ~n49808 & ~n49839;
  assign n49841 = controllable_hmaster2 & ~n49840;
  assign n49842 = i_hbusreq5 & ~n49024;
  assign n49843 = n8378 & ~n15125;
  assign n49844 = ~n8378 & ~n32188;
  assign n49845 = ~n49843 & ~n49844;
  assign n49846 = i_hlock5 & ~n49845;
  assign n49847 = ~n8378 & ~n32365;
  assign n49848 = ~n49843 & ~n49847;
  assign n49849 = ~i_hlock5 & ~n49848;
  assign n49850 = ~n49846 & ~n49849;
  assign n49851 = ~i_hbusreq5 & ~n49850;
  assign n49852 = ~n49842 & ~n49851;
  assign n49853 = controllable_hgrant5 & ~n49852;
  assign n49854 = i_hbusreq5 & ~n49056;
  assign n49855 = i_hbusreq4 & ~n49032;
  assign n49856 = i_hbusreq9 & ~n49027;
  assign n49857 = n8426 & ~n15119;
  assign n49858 = ~n8426 & ~n22145;
  assign n49859 = ~n49857 & ~n49858;
  assign n49860 = ~i_hbusreq9 & ~n49859;
  assign n49861 = ~n49856 & ~n49860;
  assign n49862 = i_hlock4 & ~n49861;
  assign n49863 = i_hbusreq9 & ~n49030;
  assign n49864 = ~n8426 & ~n22157;
  assign n49865 = ~n49857 & ~n49864;
  assign n49866 = ~i_hbusreq9 & ~n49865;
  assign n49867 = ~n49863 & ~n49866;
  assign n49868 = ~i_hlock4 & ~n49867;
  assign n49869 = ~n49862 & ~n49868;
  assign n49870 = ~i_hbusreq4 & ~n49869;
  assign n49871 = ~n49855 & ~n49870;
  assign n49872 = controllable_hgrant4 & ~n49871;
  assign n49873 = i_hbusreq4 & ~n49054;
  assign n49874 = i_hbusreq9 & ~n49054;
  assign n49875 = i_hbusreq3 & ~n49040;
  assign n49876 = n8365 & ~n15115;
  assign n49877 = ~n8365 & ~n22141;
  assign n49878 = ~n49876 & ~n49877;
  assign n49879 = i_hlock3 & ~n49878;
  assign n49880 = ~n8365 & ~n22153;
  assign n49881 = ~n49876 & ~n49880;
  assign n49882 = ~i_hlock3 & ~n49881;
  assign n49883 = ~n49879 & ~n49882;
  assign n49884 = ~i_hbusreq3 & ~n49883;
  assign n49885 = ~n49875 & ~n49884;
  assign n49886 = controllable_hgrant3 & ~n49885;
  assign n49887 = i_hbusreq3 & ~n49052;
  assign n49888 = i_hbusreq1 & ~n49048;
  assign n49889 = n8389 & ~n15111;
  assign n49890 = ~n8389 & ~n22137;
  assign n49891 = ~n49889 & ~n49890;
  assign n49892 = i_hlock1 & ~n49891;
  assign n49893 = ~n8389 & ~n22149;
  assign n49894 = ~n49889 & ~n49893;
  assign n49895 = ~i_hlock1 & ~n49894;
  assign n49896 = ~n49892 & ~n49895;
  assign n49897 = ~i_hbusreq1 & ~n49896;
  assign n49898 = ~n49888 & ~n49897;
  assign n49899 = controllable_hgrant1 & ~n49898;
  assign n49900 = i_hbusreq1 & ~n49050;
  assign n49901 = controllable_locked & ~n12895;
  assign n49902 = ~n19075 & ~n49901;
  assign n49903 = i_hlock0 & ~n49902;
  assign n49904 = ~n44269 & ~n49903;
  assign n49905 = ~i_hbusreq0 & ~n49904;
  assign n49906 = ~i_hbusreq0 & ~n49905;
  assign n49907 = ~i_hbusreq2 & ~n49906;
  assign n49908 = ~i_hbusreq2 & ~n49907;
  assign n49909 = ~controllable_hgrant2 & n49908;
  assign n49910 = ~n44865 & ~n49909;
  assign n49911 = ~n7733 & ~n49910;
  assign n49912 = ~i_hbusreq0 & ~n46057;
  assign n49913 = ~n46689 & ~n49912;
  assign n49914 = i_hlock2 & ~n49913;
  assign n49915 = ~n46058 & ~n49914;
  assign n49916 = ~i_hbusreq2 & ~n49915;
  assign n49917 = ~n46688 & ~n49916;
  assign n49918 = controllable_hgrant2 & ~n49917;
  assign n49919 = ~i_hbusreq0 & ~n44268;
  assign n49920 = ~i_hbusreq0 & ~n49919;
  assign n49921 = ~i_hbusreq2 & ~n49920;
  assign n49922 = ~i_hbusreq2 & ~n49921;
  assign n49923 = ~controllable_hgrant2 & n49922;
  assign n49924 = ~n49918 & ~n49923;
  assign n49925 = n7733 & ~n49924;
  assign n49926 = ~n49911 & ~n49925;
  assign n49927 = n7928 & ~n49926;
  assign n49928 = ~n8440 & ~n49927;
  assign n49929 = ~i_hbusreq1 & ~n49928;
  assign n49930 = ~n49900 & ~n49929;
  assign n49931 = ~controllable_hgrant1 & ~n49930;
  assign n49932 = ~n49899 & ~n49931;
  assign n49933 = ~i_hbusreq3 & ~n49932;
  assign n49934 = ~n49887 & ~n49933;
  assign n49935 = ~controllable_hgrant3 & ~n49934;
  assign n49936 = ~n49886 & ~n49935;
  assign n49937 = ~i_hbusreq9 & ~n49936;
  assign n49938 = ~n49874 & ~n49937;
  assign n49939 = ~i_hbusreq4 & ~n49938;
  assign n49940 = ~n49873 & ~n49939;
  assign n49941 = ~controllable_hgrant4 & ~n49940;
  assign n49942 = ~n49872 & ~n49941;
  assign n49943 = ~i_hbusreq5 & ~n49942;
  assign n49944 = ~n49854 & ~n49943;
  assign n49945 = ~controllable_hgrant5 & ~n49944;
  assign n49946 = ~n49853 & ~n49945;
  assign n49947 = ~controllable_hmaster2 & ~n49946;
  assign n49948 = ~n49841 & ~n49947;
  assign n49949 = ~controllable_hmaster1 & ~n49948;
  assign n49950 = ~n49796 & ~n49949;
  assign n49951 = i_hlock6 & ~n49950;
  assign n49952 = controllable_hmaster2 & ~n49459;
  assign n49953 = ~n49794 & ~n49952;
  assign n49954 = controllable_hmaster1 & ~n49953;
  assign n49955 = ~n49949 & ~n49954;
  assign n49956 = ~i_hlock6 & ~n49955;
  assign n49957 = ~n49951 & ~n49956;
  assign n49958 = ~i_hbusreq6 & ~n49957;
  assign n49959 = ~n49692 & ~n49958;
  assign n49960 = ~controllable_hgrant6 & ~n49959;
  assign n49961 = ~n49691 & ~n49960;
  assign n49962 = ~controllable_hmaster0 & ~n49961;
  assign n49963 = ~n49667 & ~n49962;
  assign n49964 = ~i_hbusreq8 & ~n49963;
  assign n49965 = ~n49475 & ~n49964;
  assign n49966 = ~controllable_hmaster3 & ~n49965;
  assign n49967 = ~n49474 & ~n49966;
  assign n49968 = i_hlock7 & ~n49967;
  assign n49969 = i_hbusreq8 & ~n49082;
  assign n49970 = n8217 & ~n15155;
  assign n49971 = ~n8217 & ~n37828;
  assign n49972 = ~n49970 & ~n49971;
  assign n49973 = i_hlock6 & ~n49972;
  assign n49974 = ~n8217 & ~n37838;
  assign n49975 = ~n49970 & ~n49974;
  assign n49976 = ~i_hlock6 & ~n49975;
  assign n49977 = ~n49973 & ~n49976;
  assign n49978 = ~i_hbusreq6 & ~n49977;
  assign n49979 = ~n45897 & ~n49978;
  assign n49980 = controllable_hgrant6 & ~n49979;
  assign n49981 = i_hbusreq6 & ~n49078;
  assign n49982 = ~n49553 & ~n49952;
  assign n49983 = controllable_hmaster1 & ~n49982;
  assign n49984 = ~n49661 & ~n49983;
  assign n49985 = ~i_hbusreq6 & ~n49984;
  assign n49986 = ~n49981 & ~n49985;
  assign n49987 = ~controllable_hgrant6 & ~n49986;
  assign n49988 = ~n49980 & ~n49987;
  assign n49989 = controllable_hmaster0 & ~n49988;
  assign n49990 = ~n49962 & ~n49989;
  assign n49991 = ~i_hbusreq8 & ~n49990;
  assign n49992 = ~n49969 & ~n49991;
  assign n49993 = ~controllable_hmaster3 & ~n49992;
  assign n49994 = ~n49474 & ~n49993;
  assign n49995 = ~i_hlock7 & ~n49994;
  assign n49996 = ~n49968 & ~n49995;
  assign n49997 = ~i_hbusreq7 & ~n49996;
  assign n49998 = ~n49087 & ~n49997;
  assign n49999 = n7924 & ~n49998;
  assign n50000 = ~n48761 & ~n49999;
  assign n50001 = n7920 & ~n50000;
  assign n50002 = ~n40177 & ~n50001;
  assign n50003 = ~n7728 & ~n50002;
  assign n50004 = ~n48005 & ~n50003;
  assign n50005 = ~n7723 & ~n50004;
  assign n50006 = ~n45934 & ~n50005;
  assign n50007 = ~n7714 & ~n50006;
  assign n50008 = ~n45933 & ~n50007;
  assign n50009 = ~n7705 & ~n50008;
  assign n50010 = ~n41283 & ~n50009;
  assign n50011 = n7808 & ~n50010;
  assign n50012 = ~n40187 & ~n50011;
  assign n50013 = n8195 & ~n50012;
  assign n50014 = ~n39684 & ~n50013;
  assign n50015 = ~n8193 & ~n50014;
  assign n50016 = controllable_hgrant6 & ~n9755;
  assign n50017 = controllable_hmaster2 & ~n39798;
  assign n50018 = ~controllable_hmaster1 & ~n50017;
  assign n50019 = ~controllable_hmaster1 & ~n50018;
  assign n50020 = ~controllable_hgrant6 & ~n50019;
  assign n50021 = ~n50016 & ~n50020;
  assign n50022 = controllable_hmaster0 & ~n50021;
  assign n50023 = controllable_hmaster0 & ~n50022;
  assign n50024 = ~controllable_hmaster3 & ~n50023;
  assign n50025 = ~controllable_hmaster3 & ~n50024;
  assign n50026 = i_hbusreq7 & ~n50025;
  assign n50027 = i_hbusreq8 & ~n50023;
  assign n50028 = controllable_hgrant6 & ~n9767;
  assign n50029 = i_hbusreq6 & ~n50019;
  assign n50030 = controllable_hmaster2 & ~n40004;
  assign n50031 = ~controllable_hmaster1 & ~n50030;
  assign n50032 = ~controllable_hmaster1 & ~n50031;
  assign n50033 = ~i_hbusreq6 & ~n50032;
  assign n50034 = ~n50029 & ~n50033;
  assign n50035 = ~controllable_hgrant6 & ~n50034;
  assign n50036 = ~n50028 & ~n50035;
  assign n50037 = controllable_hmaster0 & ~n50036;
  assign n50038 = controllable_hmaster0 & ~n50037;
  assign n50039 = ~i_hbusreq8 & ~n50038;
  assign n50040 = ~n50027 & ~n50039;
  assign n50041 = ~controllable_hmaster3 & ~n50040;
  assign n50042 = ~controllable_hmaster3 & ~n50041;
  assign n50043 = ~i_hbusreq7 & ~n50042;
  assign n50044 = ~n50026 & ~n50043;
  assign n50045 = n7924 & ~n50044;
  assign n50046 = n7924 & ~n50045;
  assign n50047 = ~n8214 & ~n50046;
  assign n50048 = controllable_hgrant6 & ~n9781;
  assign n50049 = controllable_hmaster2 & ~n39894;
  assign n50050 = ~controllable_hmaster1 & ~n50049;
  assign n50051 = ~controllable_hmaster1 & ~n50050;
  assign n50052 = ~controllable_hgrant6 & ~n50051;
  assign n50053 = ~n50048 & ~n50052;
  assign n50054 = ~controllable_hmaster0 & ~n50053;
  assign n50055 = ~controllable_hmaster0 & ~n50054;
  assign n50056 = ~controllable_hmaster3 & ~n50055;
  assign n50057 = ~controllable_hmaster3 & ~n50056;
  assign n50058 = i_hbusreq7 & ~n50057;
  assign n50059 = i_hbusreq8 & ~n50055;
  assign n50060 = controllable_hgrant6 & ~n9793;
  assign n50061 = i_hbusreq6 & ~n50051;
  assign n50062 = controllable_hmaster2 & ~n40145;
  assign n50063 = ~controllable_hmaster1 & ~n50062;
  assign n50064 = ~controllable_hmaster1 & ~n50063;
  assign n50065 = ~i_hbusreq6 & ~n50064;
  assign n50066 = ~n50061 & ~n50065;
  assign n50067 = ~controllable_hgrant6 & ~n50066;
  assign n50068 = ~n50060 & ~n50067;
  assign n50069 = ~controllable_hmaster0 & ~n50068;
  assign n50070 = ~controllable_hmaster0 & ~n50069;
  assign n50071 = ~i_hbusreq8 & ~n50070;
  assign n50072 = ~n50059 & ~n50071;
  assign n50073 = ~controllable_hmaster3 & ~n50072;
  assign n50074 = ~controllable_hmaster3 & ~n50073;
  assign n50075 = ~i_hbusreq7 & ~n50074;
  assign n50076 = ~n50058 & ~n50075;
  assign n50077 = n7924 & ~n50076;
  assign n50078 = n7924 & ~n50077;
  assign n50079 = n8214 & ~n50078;
  assign n50080 = ~n50047 & ~n50079;
  assign n50081 = ~n8202 & ~n50080;
  assign n50082 = controllable_hgrant6 & ~n9807;
  assign n50083 = controllable_hmaster1 & ~n39787;
  assign n50084 = ~controllable_hgrant6 & ~n50083;
  assign n50085 = ~n50082 & ~n50084;
  assign n50086 = controllable_hmaster0 & ~n50085;
  assign n50087 = controllable_hmaster0 & ~n50086;
  assign n50088 = ~controllable_hmaster3 & ~n50087;
  assign n50089 = ~controllable_hmaster3 & ~n50088;
  assign n50090 = i_hbusreq7 & ~n50089;
  assign n50091 = i_hbusreq8 & ~n50087;
  assign n50092 = controllable_hgrant6 & ~n9817;
  assign n50093 = i_hbusreq6 & ~n50083;
  assign n50094 = controllable_hmaster1 & ~n39990;
  assign n50095 = ~i_hbusreq6 & ~n50094;
  assign n50096 = ~n50093 & ~n50095;
  assign n50097 = ~controllable_hgrant6 & ~n50096;
  assign n50098 = ~n50092 & ~n50097;
  assign n50099 = controllable_hmaster0 & ~n50098;
  assign n50100 = controllable_hmaster0 & ~n50099;
  assign n50101 = ~i_hbusreq8 & ~n50100;
  assign n50102 = ~n50091 & ~n50101;
  assign n50103 = ~controllable_hmaster3 & ~n50102;
  assign n50104 = ~controllable_hmaster3 & ~n50103;
  assign n50105 = ~i_hbusreq7 & ~n50104;
  assign n50106 = ~n50090 & ~n50105;
  assign n50107 = n7924 & ~n50106;
  assign n50108 = n7924 & ~n50107;
  assign n50109 = ~n8214 & ~n50108;
  assign n50110 = controllable_hgrant6 & ~n9829;
  assign n50111 = controllable_hmaster1 & ~n39880;
  assign n50112 = ~controllable_hgrant6 & ~n50111;
  assign n50113 = ~n50110 & ~n50112;
  assign n50114 = ~controllable_hmaster0 & ~n50113;
  assign n50115 = ~controllable_hmaster0 & ~n50114;
  assign n50116 = ~controllable_hmaster3 & ~n50115;
  assign n50117 = ~controllable_hmaster3 & ~n50116;
  assign n50118 = i_hbusreq7 & ~n50117;
  assign n50119 = i_hbusreq8 & ~n50115;
  assign n50120 = controllable_hgrant6 & ~n9839;
  assign n50121 = i_hbusreq6 & ~n50111;
  assign n50122 = controllable_hmaster1 & ~n40119;
  assign n50123 = ~i_hbusreq6 & ~n50122;
  assign n50124 = ~n50121 & ~n50123;
  assign n50125 = ~controllable_hgrant6 & ~n50124;
  assign n50126 = ~n50120 & ~n50125;
  assign n50127 = ~controllable_hmaster0 & ~n50126;
  assign n50128 = ~controllable_hmaster0 & ~n50127;
  assign n50129 = ~i_hbusreq8 & ~n50128;
  assign n50130 = ~n50119 & ~n50129;
  assign n50131 = ~controllable_hmaster3 & ~n50130;
  assign n50132 = ~controllable_hmaster3 & ~n50131;
  assign n50133 = ~i_hbusreq7 & ~n50132;
  assign n50134 = ~n50118 & ~n50133;
  assign n50135 = n7924 & ~n50134;
  assign n50136 = n7924 & ~n50135;
  assign n50137 = n8214 & ~n50136;
  assign n50138 = ~n50109 & ~n50137;
  assign n50139 = n8202 & ~n50138;
  assign n50140 = ~n50081 & ~n50139;
  assign n50141 = n7728 & ~n50140;
  assign n50142 = ~n7840 & ~n50024;
  assign n50143 = i_hbusreq7 & ~n50142;
  assign n50144 = ~n7901 & ~n50041;
  assign n50145 = ~i_hbusreq7 & ~n50144;
  assign n50146 = ~n50143 & ~n50145;
  assign n50147 = n7924 & ~n50146;
  assign n50148 = ~n39731 & ~n50147;
  assign n50149 = ~n8214 & ~n50148;
  assign n50150 = ~n7840 & ~n50056;
  assign n50151 = i_hbusreq7 & ~n50150;
  assign n50152 = ~n7901 & ~n50073;
  assign n50153 = ~i_hbusreq7 & ~n50152;
  assign n50154 = ~n50151 & ~n50153;
  assign n50155 = n7924 & ~n50154;
  assign n50156 = ~n39731 & ~n50155;
  assign n50157 = n8214 & ~n50156;
  assign n50158 = ~n50149 & ~n50157;
  assign n50159 = ~n8202 & ~n50158;
  assign n50160 = ~n7840 & ~n50088;
  assign n50161 = i_hbusreq7 & ~n50160;
  assign n50162 = ~n7901 & ~n50103;
  assign n50163 = ~i_hbusreq7 & ~n50162;
  assign n50164 = ~n50161 & ~n50163;
  assign n50165 = n7924 & ~n50164;
  assign n50166 = ~n39731 & ~n50165;
  assign n50167 = ~n8214 & ~n50166;
  assign n50168 = ~n7840 & ~n50116;
  assign n50169 = i_hbusreq7 & ~n50168;
  assign n50170 = ~n7901 & ~n50131;
  assign n50171 = ~i_hbusreq7 & ~n50170;
  assign n50172 = ~n50169 & ~n50171;
  assign n50173 = n7924 & ~n50172;
  assign n50174 = ~n39731 & ~n50173;
  assign n50175 = n8214 & ~n50174;
  assign n50176 = ~n50167 & ~n50175;
  assign n50177 = n8202 & ~n50176;
  assign n50178 = ~n50159 & ~n50177;
  assign n50179 = ~n7728 & ~n50178;
  assign n50180 = ~n50141 & ~n50179;
  assign n50181 = ~n7723 & ~n50180;
  assign n50182 = ~n7723 & ~n50181;
  assign n50183 = ~n7714 & ~n50182;
  assign n50184 = ~n7714 & ~n50183;
  assign n50185 = n7705 & ~n50184;
  assign n50186 = n7723 & ~n50178;
  assign n50187 = n7920 & ~n50178;
  assign n50188 = ~n40177 & ~n50187;
  assign n50189 = ~n7723 & ~n50188;
  assign n50190 = ~n50186 & ~n50189;
  assign n50191 = n7714 & ~n50190;
  assign n50192 = ~n40183 & ~n50191;
  assign n50193 = ~n7705 & ~n50192;
  assign n50194 = ~n50185 & ~n50193;
  assign n50195 = ~n7808 & ~n50194;
  assign n50196 = ~n7920 & ~n50140;
  assign n50197 = n8217 & ~n9912;
  assign n50198 = ~n8217 & ~n22237;
  assign n50199 = ~n50197 & ~n50198;
  assign n50200 = controllable_hgrant6 & ~n50199;
  assign n50201 = controllable_hmaster2 & ~n48097;
  assign n50202 = ~controllable_hmaster1 & ~n50201;
  assign n50203 = ~controllable_hmaster1 & ~n50202;
  assign n50204 = ~controllable_hgrant6 & ~n50203;
  assign n50205 = ~n50200 & ~n50204;
  assign n50206 = controllable_hmaster0 & ~n50205;
  assign n50207 = controllable_hmaster0 & ~n50206;
  assign n50208 = ~controllable_hmaster3 & ~n50207;
  assign n50209 = ~controllable_hmaster3 & ~n50208;
  assign n50210 = i_hbusreq7 & ~n50209;
  assign n50211 = i_hbusreq8 & ~n50207;
  assign n50212 = i_hbusreq6 & ~n50199;
  assign n50213 = n8217 & ~n9922;
  assign n50214 = ~n8217 & ~n22250;
  assign n50215 = ~n50213 & ~n50214;
  assign n50216 = ~i_hbusreq6 & ~n50215;
  assign n50217 = ~n50212 & ~n50216;
  assign n50218 = controllable_hgrant6 & ~n50217;
  assign n50219 = i_hbusreq6 & ~n50203;
  assign n50220 = controllable_hmaster2 & ~n48432;
  assign n50221 = ~controllable_hmaster1 & ~n50220;
  assign n50222 = ~controllable_hmaster1 & ~n50221;
  assign n50223 = ~i_hbusreq6 & ~n50222;
  assign n50224 = ~n50219 & ~n50223;
  assign n50225 = ~controllable_hgrant6 & ~n50224;
  assign n50226 = ~n50218 & ~n50225;
  assign n50227 = controllable_hmaster0 & ~n50226;
  assign n50228 = controllable_hmaster0 & ~n50227;
  assign n50229 = ~i_hbusreq8 & ~n50228;
  assign n50230 = ~n50211 & ~n50229;
  assign n50231 = ~controllable_hmaster3 & ~n50230;
  assign n50232 = ~controllable_hmaster3 & ~n50231;
  assign n50233 = ~i_hbusreq7 & ~n50232;
  assign n50234 = ~n50210 & ~n50233;
  assign n50235 = ~n7924 & ~n50234;
  assign n50236 = n8378 & ~n12794;
  assign n50237 = ~n8378 & ~n28963;
  assign n50238 = ~n50236 & ~n50237;
  assign n50239 = i_hlock5 & ~n50238;
  assign n50240 = ~n8378 & ~n28988;
  assign n50241 = ~n50236 & ~n50240;
  assign n50242 = ~i_hlock5 & ~n50241;
  assign n50243 = ~n50239 & ~n50242;
  assign n50244 = controllable_hgrant5 & ~n50243;
  assign n50245 = controllable_hgrant5 & ~n50244;
  assign n50246 = ~controllable_hgrant6 & ~n50245;
  assign n50247 = ~controllable_hgrant6 & ~n50246;
  assign n50248 = controllable_hmaster3 & ~n50247;
  assign n50249 = controllable_hmaster1 & ~n50245;
  assign n50250 = ~n48095 & ~n48879;
  assign n50251 = controllable_hmaster2 & ~n50250;
  assign n50252 = ~controllable_hmaster2 & ~n50245;
  assign n50253 = ~n50251 & ~n50252;
  assign n50254 = ~controllable_hmaster1 & ~n50253;
  assign n50255 = ~n50249 & ~n50254;
  assign n50256 = ~controllable_hgrant6 & ~n50255;
  assign n50257 = ~n50200 & ~n50256;
  assign n50258 = controllable_hmaster0 & ~n50257;
  assign n50259 = ~controllable_hmaster0 & ~n50247;
  assign n50260 = ~n50258 & ~n50259;
  assign n50261 = ~controllable_hmaster3 & ~n50260;
  assign n50262 = ~n50248 & ~n50261;
  assign n50263 = i_hbusreq7 & ~n50262;
  assign n50264 = i_hbusreq8 & ~n50247;
  assign n50265 = i_hbusreq6 & ~n50245;
  assign n50266 = i_hbusreq5 & ~n50243;
  assign n50267 = n8378 & ~n12871;
  assign n50268 = ~n8378 & ~n29024;
  assign n50269 = ~n50267 & ~n50268;
  assign n50270 = i_hlock5 & ~n50269;
  assign n50271 = ~n8378 & ~n29079;
  assign n50272 = ~n50267 & ~n50271;
  assign n50273 = ~i_hlock5 & ~n50272;
  assign n50274 = ~n50270 & ~n50273;
  assign n50275 = ~i_hbusreq5 & ~n50274;
  assign n50276 = ~n50266 & ~n50275;
  assign n50277 = controllable_hgrant5 & ~n50276;
  assign n50278 = controllable_hgrant5 & ~n50277;
  assign n50279 = ~i_hbusreq6 & ~n50278;
  assign n50280 = ~n50265 & ~n50279;
  assign n50281 = ~controllable_hgrant6 & ~n50280;
  assign n50282 = ~controllable_hgrant6 & ~n50281;
  assign n50283 = ~i_hbusreq8 & ~n50282;
  assign n50284 = ~n50264 & ~n50283;
  assign n50285 = controllable_hmaster3 & ~n50284;
  assign n50286 = i_hbusreq8 & ~n50260;
  assign n50287 = i_hbusreq6 & ~n50255;
  assign n50288 = controllable_hmaster1 & ~n50278;
  assign n50289 = ~n48430 & ~n49568;
  assign n50290 = controllable_hmaster2 & ~n50289;
  assign n50291 = ~controllable_hmaster2 & ~n50278;
  assign n50292 = ~n50290 & ~n50291;
  assign n50293 = ~controllable_hmaster1 & ~n50292;
  assign n50294 = ~n50288 & ~n50293;
  assign n50295 = ~i_hbusreq6 & ~n50294;
  assign n50296 = ~n50287 & ~n50295;
  assign n50297 = ~controllable_hgrant6 & ~n50296;
  assign n50298 = ~n50218 & ~n50297;
  assign n50299 = controllable_hmaster0 & ~n50298;
  assign n50300 = ~controllable_hmaster0 & ~n50282;
  assign n50301 = ~n50299 & ~n50300;
  assign n50302 = ~i_hbusreq8 & ~n50301;
  assign n50303 = ~n50286 & ~n50302;
  assign n50304 = ~controllable_hmaster3 & ~n50303;
  assign n50305 = ~n50285 & ~n50304;
  assign n50306 = ~i_hbusreq7 & ~n50305;
  assign n50307 = ~n50263 & ~n50306;
  assign n50308 = n7924 & ~n50307;
  assign n50309 = ~n50235 & ~n50308;
  assign n50310 = ~n8214 & ~n50309;
  assign n50311 = n8217 & ~n9936;
  assign n50312 = ~n8217 & ~n22267;
  assign n50313 = ~n50311 & ~n50312;
  assign n50314 = controllable_hgrant6 & ~n50313;
  assign n50315 = controllable_hmaster2 & ~n48185;
  assign n50316 = ~controllable_hmaster1 & ~n50315;
  assign n50317 = ~controllable_hmaster1 & ~n50316;
  assign n50318 = ~controllable_hgrant6 & ~n50317;
  assign n50319 = ~n50314 & ~n50318;
  assign n50320 = ~controllable_hmaster0 & ~n50319;
  assign n50321 = ~controllable_hmaster0 & ~n50320;
  assign n50322 = ~controllable_hmaster3 & ~n50321;
  assign n50323 = ~controllable_hmaster3 & ~n50322;
  assign n50324 = i_hbusreq7 & ~n50323;
  assign n50325 = i_hbusreq8 & ~n50321;
  assign n50326 = i_hbusreq6 & ~n50313;
  assign n50327 = n8217 & ~n9946;
  assign n50328 = ~n8217 & ~n22280;
  assign n50329 = ~n50327 & ~n50328;
  assign n50330 = ~i_hbusreq6 & ~n50329;
  assign n50331 = ~n50326 & ~n50330;
  assign n50332 = controllable_hgrant6 & ~n50331;
  assign n50333 = i_hbusreq6 & ~n50317;
  assign n50334 = controllable_hmaster2 & ~n48648;
  assign n50335 = ~controllable_hmaster1 & ~n50334;
  assign n50336 = ~controllable_hmaster1 & ~n50335;
  assign n50337 = ~i_hbusreq6 & ~n50336;
  assign n50338 = ~n50333 & ~n50337;
  assign n50339 = ~controllable_hgrant6 & ~n50338;
  assign n50340 = ~n50332 & ~n50339;
  assign n50341 = ~controllable_hmaster0 & ~n50340;
  assign n50342 = ~controllable_hmaster0 & ~n50341;
  assign n50343 = ~i_hbusreq8 & ~n50342;
  assign n50344 = ~n50325 & ~n50343;
  assign n50345 = ~controllable_hmaster3 & ~n50344;
  assign n50346 = ~controllable_hmaster3 & ~n50345;
  assign n50347 = ~i_hbusreq7 & ~n50346;
  assign n50348 = ~n50324 & ~n50347;
  assign n50349 = ~n7924 & ~n50348;
  assign n50350 = n8426 & ~n12792;
  assign n50351 = ~n8426 & ~n16481;
  assign n50352 = ~n50350 & ~n50351;
  assign n50353 = i_hlock4 & ~n50352;
  assign n50354 = ~n8426 & ~n16495;
  assign n50355 = ~n50350 & ~n50354;
  assign n50356 = ~i_hlock4 & ~n50355;
  assign n50357 = ~n50353 & ~n50356;
  assign n50358 = controllable_hgrant4 & ~n50357;
  assign n50359 = controllable_hgrant4 & ~n50358;
  assign n50360 = ~controllable_hgrant5 & ~n50359;
  assign n50361 = ~controllable_hgrant5 & ~n50360;
  assign n50362 = ~controllable_hgrant6 & ~n50361;
  assign n50363 = ~controllable_hgrant6 & ~n50362;
  assign n50364 = controllable_hmaster3 & ~n50363;
  assign n50365 = controllable_hmaster0 & ~n50363;
  assign n50366 = controllable_hmaster1 & ~n50361;
  assign n50367 = ~n48181 & ~n49009;
  assign n50368 = ~controllable_hgrant5 & ~n50367;
  assign n50369 = ~n48169 & ~n50368;
  assign n50370 = controllable_hmaster2 & ~n50369;
  assign n50371 = ~controllable_hmaster2 & ~n50361;
  assign n50372 = ~n50370 & ~n50371;
  assign n50373 = ~controllable_hmaster1 & ~n50372;
  assign n50374 = ~n50366 & ~n50373;
  assign n50375 = ~controllable_hgrant6 & ~n50374;
  assign n50376 = ~n50314 & ~n50375;
  assign n50377 = ~controllable_hmaster0 & ~n50376;
  assign n50378 = ~n50365 & ~n50377;
  assign n50379 = ~controllable_hmaster3 & ~n50378;
  assign n50380 = ~n50364 & ~n50379;
  assign n50381 = i_hbusreq7 & ~n50380;
  assign n50382 = i_hbusreq8 & ~n50363;
  assign n50383 = i_hbusreq6 & ~n50361;
  assign n50384 = i_hbusreq5 & ~n50359;
  assign n50385 = i_hbusreq4 & ~n50357;
  assign n50386 = i_hbusreq9 & ~n50352;
  assign n50387 = n8426 & ~n12865;
  assign n50388 = ~n8426 & ~n16589;
  assign n50389 = ~n50387 & ~n50388;
  assign n50390 = ~i_hbusreq9 & ~n50389;
  assign n50391 = ~n50386 & ~n50390;
  assign n50392 = i_hlock4 & ~n50391;
  assign n50393 = i_hbusreq9 & ~n50355;
  assign n50394 = ~n8426 & ~n16603;
  assign n50395 = ~n50387 & ~n50394;
  assign n50396 = ~i_hbusreq9 & ~n50395;
  assign n50397 = ~n50393 & ~n50396;
  assign n50398 = ~i_hlock4 & ~n50397;
  assign n50399 = ~n50392 & ~n50398;
  assign n50400 = ~i_hbusreq4 & ~n50399;
  assign n50401 = ~n50385 & ~n50400;
  assign n50402 = controllable_hgrant4 & ~n50401;
  assign n50403 = controllable_hgrant4 & ~n50402;
  assign n50404 = ~i_hbusreq5 & ~n50403;
  assign n50405 = ~n50384 & ~n50404;
  assign n50406 = ~controllable_hgrant5 & ~n50405;
  assign n50407 = ~controllable_hgrant5 & ~n50406;
  assign n50408 = ~i_hbusreq6 & ~n50407;
  assign n50409 = ~n50383 & ~n50408;
  assign n50410 = ~controllable_hgrant6 & ~n50409;
  assign n50411 = ~controllable_hgrant6 & ~n50410;
  assign n50412 = ~i_hbusreq8 & ~n50411;
  assign n50413 = ~n50382 & ~n50412;
  assign n50414 = controllable_hmaster3 & ~n50413;
  assign n50415 = i_hbusreq8 & ~n50378;
  assign n50416 = controllable_hmaster0 & ~n50411;
  assign n50417 = i_hbusreq6 & ~n50374;
  assign n50418 = controllable_hmaster1 & ~n50407;
  assign n50419 = i_hbusreq5 & ~n50367;
  assign n50420 = ~n48642 & ~n49828;
  assign n50421 = ~i_hbusreq5 & ~n50420;
  assign n50422 = ~n50419 & ~n50421;
  assign n50423 = ~controllable_hgrant5 & ~n50422;
  assign n50424 = ~n48615 & ~n50423;
  assign n50425 = controllable_hmaster2 & ~n50424;
  assign n50426 = ~controllable_hmaster2 & ~n50407;
  assign n50427 = ~n50425 & ~n50426;
  assign n50428 = ~controllable_hmaster1 & ~n50427;
  assign n50429 = ~n50418 & ~n50428;
  assign n50430 = ~i_hbusreq6 & ~n50429;
  assign n50431 = ~n50417 & ~n50430;
  assign n50432 = ~controllable_hgrant6 & ~n50431;
  assign n50433 = ~n50332 & ~n50432;
  assign n50434 = ~controllable_hmaster0 & ~n50433;
  assign n50435 = ~n50416 & ~n50434;
  assign n50436 = ~i_hbusreq8 & ~n50435;
  assign n50437 = ~n50415 & ~n50436;
  assign n50438 = ~controllable_hmaster3 & ~n50437;
  assign n50439 = ~n50414 & ~n50438;
  assign n50440 = ~i_hbusreq7 & ~n50439;
  assign n50441 = ~n50381 & ~n50440;
  assign n50442 = n7924 & ~n50441;
  assign n50443 = ~n50349 & ~n50442;
  assign n50444 = n8214 & ~n50443;
  assign n50445 = ~n50310 & ~n50444;
  assign n50446 = ~n8202 & ~n50445;
  assign n50447 = n8217 & ~n9962;
  assign n50448 = ~n8217 & ~n22299;
  assign n50449 = ~n50447 & ~n50448;
  assign n50450 = controllable_hgrant6 & ~n50449;
  assign n50451 = ~controllable_hmaster2 & ~n48081;
  assign n50452 = controllable_hmaster1 & ~n50451;
  assign n50453 = controllable_hmaster1 & ~n50452;
  assign n50454 = ~controllable_hgrant6 & ~n50453;
  assign n50455 = ~n50450 & ~n50454;
  assign n50456 = controllable_hmaster0 & ~n50455;
  assign n50457 = controllable_hmaster0 & ~n50456;
  assign n50458 = ~controllable_hmaster3 & ~n50457;
  assign n50459 = ~controllable_hmaster3 & ~n50458;
  assign n50460 = i_hbusreq7 & ~n50459;
  assign n50461 = i_hbusreq8 & ~n50457;
  assign n50462 = i_hbusreq6 & ~n50449;
  assign n50463 = n8217 & ~n9972;
  assign n50464 = ~n8217 & ~n22312;
  assign n50465 = ~n50463 & ~n50464;
  assign n50466 = ~i_hbusreq6 & ~n50465;
  assign n50467 = ~n50462 & ~n50466;
  assign n50468 = controllable_hgrant6 & ~n50467;
  assign n50469 = i_hbusreq6 & ~n50453;
  assign n50470 = ~controllable_hmaster2 & ~n48408;
  assign n50471 = controllable_hmaster1 & ~n50470;
  assign n50472 = controllable_hmaster1 & ~n50471;
  assign n50473 = ~i_hbusreq6 & ~n50472;
  assign n50474 = ~n50469 & ~n50473;
  assign n50475 = ~controllable_hgrant6 & ~n50474;
  assign n50476 = ~n50468 & ~n50475;
  assign n50477 = controllable_hmaster0 & ~n50476;
  assign n50478 = controllable_hmaster0 & ~n50477;
  assign n50479 = ~i_hbusreq8 & ~n50478;
  assign n50480 = ~n50461 & ~n50479;
  assign n50481 = ~controllable_hmaster3 & ~n50480;
  assign n50482 = ~controllable_hmaster3 & ~n50481;
  assign n50483 = ~i_hbusreq7 & ~n50482;
  assign n50484 = ~n50460 & ~n50483;
  assign n50485 = ~n7924 & ~n50484;
  assign n50486 = n8365 & ~n12790;
  assign n50487 = ~n8365 & ~n16479;
  assign n50488 = ~n50486 & ~n50487;
  assign n50489 = i_hlock3 & ~n50488;
  assign n50490 = ~n8365 & ~n16493;
  assign n50491 = ~n50486 & ~n50490;
  assign n50492 = ~i_hlock3 & ~n50491;
  assign n50493 = ~n50489 & ~n50492;
  assign n50494 = controllable_hgrant3 & ~n50493;
  assign n50495 = controllable_hgrant3 & ~n50494;
  assign n50496 = ~controllable_hgrant4 & ~n50495;
  assign n50497 = ~controllable_hgrant4 & ~n50496;
  assign n50498 = ~controllable_hgrant5 & ~n50497;
  assign n50499 = ~controllable_hgrant5 & ~n50498;
  assign n50500 = ~controllable_hgrant6 & ~n50499;
  assign n50501 = ~controllable_hgrant6 & ~n50500;
  assign n50502 = controllable_hmaster3 & ~n50501;
  assign n50503 = controllable_hmaster2 & ~n50499;
  assign n50504 = ~n48075 & ~n48859;
  assign n50505 = ~controllable_hgrant4 & ~n50504;
  assign n50506 = ~n48063 & ~n50505;
  assign n50507 = ~controllable_hgrant5 & ~n50506;
  assign n50508 = ~n48060 & ~n50507;
  assign n50509 = ~controllable_hmaster2 & ~n50508;
  assign n50510 = ~n50503 & ~n50509;
  assign n50511 = controllable_hmaster1 & ~n50510;
  assign n50512 = ~controllable_hmaster1 & ~n50499;
  assign n50513 = ~n50511 & ~n50512;
  assign n50514 = ~controllable_hgrant6 & ~n50513;
  assign n50515 = ~n50450 & ~n50514;
  assign n50516 = controllable_hmaster0 & ~n50515;
  assign n50517 = ~controllable_hmaster0 & ~n50501;
  assign n50518 = ~n50516 & ~n50517;
  assign n50519 = ~controllable_hmaster3 & ~n50518;
  assign n50520 = ~n50502 & ~n50519;
  assign n50521 = i_hbusreq7 & ~n50520;
  assign n50522 = i_hbusreq8 & ~n50501;
  assign n50523 = i_hbusreq6 & ~n50499;
  assign n50524 = i_hbusreq5 & ~n50497;
  assign n50525 = i_hbusreq4 & ~n50495;
  assign n50526 = i_hbusreq9 & ~n50495;
  assign n50527 = i_hbusreq3 & ~n50493;
  assign n50528 = n8365 & ~n12861;
  assign n50529 = ~n8365 & ~n16585;
  assign n50530 = ~n50528 & ~n50529;
  assign n50531 = i_hlock3 & ~n50530;
  assign n50532 = ~n8365 & ~n16599;
  assign n50533 = ~n50528 & ~n50532;
  assign n50534 = ~i_hlock3 & ~n50533;
  assign n50535 = ~n50531 & ~n50534;
  assign n50536 = ~i_hbusreq3 & ~n50535;
  assign n50537 = ~n50527 & ~n50536;
  assign n50538 = controllable_hgrant3 & ~n50537;
  assign n50539 = controllable_hgrant3 & ~n50538;
  assign n50540 = ~i_hbusreq9 & ~n50539;
  assign n50541 = ~n50526 & ~n50540;
  assign n50542 = ~i_hbusreq4 & ~n50541;
  assign n50543 = ~n50525 & ~n50542;
  assign n50544 = ~controllable_hgrant4 & ~n50543;
  assign n50545 = ~controllable_hgrant4 & ~n50544;
  assign n50546 = ~i_hbusreq5 & ~n50545;
  assign n50547 = ~n50524 & ~n50546;
  assign n50548 = ~controllable_hgrant5 & ~n50547;
  assign n50549 = ~controllable_hgrant5 & ~n50548;
  assign n50550 = ~i_hbusreq6 & ~n50549;
  assign n50551 = ~n50523 & ~n50550;
  assign n50552 = ~controllable_hgrant6 & ~n50551;
  assign n50553 = ~controllable_hgrant6 & ~n50552;
  assign n50554 = ~i_hbusreq8 & ~n50553;
  assign n50555 = ~n50522 & ~n50554;
  assign n50556 = controllable_hmaster3 & ~n50555;
  assign n50557 = i_hbusreq8 & ~n50518;
  assign n50558 = i_hbusreq6 & ~n50513;
  assign n50559 = controllable_hmaster2 & ~n50549;
  assign n50560 = i_hbusreq5 & ~n50506;
  assign n50561 = i_hbusreq4 & ~n50504;
  assign n50562 = i_hbusreq9 & ~n50504;
  assign n50563 = ~n48396 & ~n49534;
  assign n50564 = ~i_hbusreq9 & ~n50563;
  assign n50565 = ~n50562 & ~n50564;
  assign n50566 = ~i_hbusreq4 & ~n50565;
  assign n50567 = ~n50561 & ~n50566;
  assign n50568 = ~controllable_hgrant4 & ~n50567;
  assign n50569 = ~n48374 & ~n50568;
  assign n50570 = ~i_hbusreq5 & ~n50569;
  assign n50571 = ~n50560 & ~n50570;
  assign n50572 = ~controllable_hgrant5 & ~n50571;
  assign n50573 = ~n48363 & ~n50572;
  assign n50574 = ~controllable_hmaster2 & ~n50573;
  assign n50575 = ~n50559 & ~n50574;
  assign n50576 = controllable_hmaster1 & ~n50575;
  assign n50577 = ~controllable_hmaster1 & ~n50549;
  assign n50578 = ~n50576 & ~n50577;
  assign n50579 = ~i_hbusreq6 & ~n50578;
  assign n50580 = ~n50558 & ~n50579;
  assign n50581 = ~controllable_hgrant6 & ~n50580;
  assign n50582 = ~n50468 & ~n50581;
  assign n50583 = controllable_hmaster0 & ~n50582;
  assign n50584 = ~controllable_hmaster0 & ~n50553;
  assign n50585 = ~n50583 & ~n50584;
  assign n50586 = ~i_hbusreq8 & ~n50585;
  assign n50587 = ~n50557 & ~n50586;
  assign n50588 = ~controllable_hmaster3 & ~n50587;
  assign n50589 = ~n50556 & ~n50588;
  assign n50590 = ~i_hbusreq7 & ~n50589;
  assign n50591 = ~n50521 & ~n50590;
  assign n50592 = n7924 & ~n50591;
  assign n50593 = ~n50485 & ~n50592;
  assign n50594 = ~n8214 & ~n50593;
  assign n50595 = n8217 & ~n9986;
  assign n50596 = ~n8217 & ~n22329;
  assign n50597 = ~n50595 & ~n50596;
  assign n50598 = controllable_hgrant6 & ~n50597;
  assign n50599 = ~controllable_hmaster2 & ~n48164;
  assign n50600 = controllable_hmaster1 & ~n50599;
  assign n50601 = controllable_hmaster1 & ~n50600;
  assign n50602 = ~controllable_hgrant6 & ~n50601;
  assign n50603 = ~n50598 & ~n50602;
  assign n50604 = ~controllable_hmaster0 & ~n50603;
  assign n50605 = ~controllable_hmaster0 & ~n50604;
  assign n50606 = ~controllable_hmaster3 & ~n50605;
  assign n50607 = ~controllable_hmaster3 & ~n50606;
  assign n50608 = i_hbusreq7 & ~n50607;
  assign n50609 = i_hbusreq8 & ~n50605;
  assign n50610 = i_hbusreq6 & ~n50597;
  assign n50611 = n8217 & ~n9996;
  assign n50612 = ~n8217 & ~n22342;
  assign n50613 = ~n50611 & ~n50612;
  assign n50614 = ~i_hbusreq6 & ~n50613;
  assign n50615 = ~n50610 & ~n50614;
  assign n50616 = controllable_hgrant6 & ~n50615;
  assign n50617 = i_hbusreq6 & ~n50601;
  assign n50618 = ~controllable_hmaster2 & ~n48606;
  assign n50619 = controllable_hmaster1 & ~n50618;
  assign n50620 = controllable_hmaster1 & ~n50619;
  assign n50621 = ~i_hbusreq6 & ~n50620;
  assign n50622 = ~n50617 & ~n50621;
  assign n50623 = ~controllable_hgrant6 & ~n50622;
  assign n50624 = ~n50616 & ~n50623;
  assign n50625 = ~controllable_hmaster0 & ~n50624;
  assign n50626 = ~controllable_hmaster0 & ~n50625;
  assign n50627 = ~i_hbusreq8 & ~n50626;
  assign n50628 = ~n50609 & ~n50627;
  assign n50629 = ~controllable_hmaster3 & ~n50628;
  assign n50630 = ~controllable_hmaster3 & ~n50629;
  assign n50631 = ~i_hbusreq7 & ~n50630;
  assign n50632 = ~n50608 & ~n50631;
  assign n50633 = ~n7924 & ~n50632;
  assign n50634 = ~n12781 & ~n45977;
  assign n50635 = ~controllable_locked & ~n50634;
  assign n50636 = ~controllable_locked & ~n50635;
  assign n50637 = controllable_hgrant2 & ~n50636;
  assign n50638 = controllable_hgrant2 & ~n50637;
  assign n50639 = ~n7733 & ~n50638;
  assign n50640 = controllable_locked & ~n45976;
  assign n50641 = ~n50635 & ~n50640;
  assign n50642 = i_hlock2 & ~n50641;
  assign n50643 = ~n46583 & ~n50635;
  assign n50644 = ~i_hlock2 & ~n50643;
  assign n50645 = ~n50642 & ~n50644;
  assign n50646 = controllable_hgrant2 & ~n50645;
  assign n50647 = controllable_hgrant2 & ~n50646;
  assign n50648 = n7733 & ~n50647;
  assign n50649 = ~n50639 & ~n50648;
  assign n50650 = n7928 & ~n50649;
  assign n50651 = n7928 & ~n50650;
  assign n50652 = ~controllable_hgrant1 & ~n50651;
  assign n50653 = ~controllable_hgrant1 & ~n50652;
  assign n50654 = ~controllable_hgrant3 & ~n50653;
  assign n50655 = ~controllable_hgrant3 & ~n50654;
  assign n50656 = ~controllable_hgrant4 & ~n50655;
  assign n50657 = ~controllable_hgrant4 & ~n50656;
  assign n50658 = ~controllable_hgrant5 & ~n50657;
  assign n50659 = ~controllable_hgrant5 & ~n50658;
  assign n50660 = ~controllable_hgrant6 & ~n50659;
  assign n50661 = ~controllable_hgrant6 & ~n50660;
  assign n50662 = controllable_hmaster3 & ~n50661;
  assign n50663 = controllable_hmaster0 & ~n50661;
  assign n50664 = controllable_hmaster2 & ~n50659;
  assign n50665 = ~n16998 & ~n44035;
  assign n50666 = ~n7733 & ~n50665;
  assign n50667 = ~n16998 & ~n48978;
  assign n50668 = n7733 & ~n50667;
  assign n50669 = ~n50666 & ~n50668;
  assign n50670 = n7928 & ~n50669;
  assign n50671 = ~n42965 & ~n50670;
  assign n50672 = ~controllable_hgrant1 & ~n50671;
  assign n50673 = ~n48144 & ~n50672;
  assign n50674 = ~controllable_hgrant3 & ~n50673;
  assign n50675 = ~n48141 & ~n50674;
  assign n50676 = ~controllable_hgrant4 & ~n50675;
  assign n50677 = ~n48138 & ~n50676;
  assign n50678 = ~controllable_hgrant5 & ~n50677;
  assign n50679 = ~n48135 & ~n50678;
  assign n50680 = ~controllable_hmaster2 & ~n50679;
  assign n50681 = ~n50664 & ~n50680;
  assign n50682 = controllable_hmaster1 & ~n50681;
  assign n50683 = ~controllable_hmaster1 & ~n50659;
  assign n50684 = ~n50682 & ~n50683;
  assign n50685 = ~controllable_hgrant6 & ~n50684;
  assign n50686 = ~n50598 & ~n50685;
  assign n50687 = ~controllable_hmaster0 & ~n50686;
  assign n50688 = ~n50663 & ~n50687;
  assign n50689 = ~controllable_hmaster3 & ~n50688;
  assign n50690 = ~n50662 & ~n50689;
  assign n50691 = i_hbusreq7 & ~n50690;
  assign n50692 = i_hbusreq8 & ~n50661;
  assign n50693 = i_hbusreq6 & ~n50659;
  assign n50694 = i_hbusreq5 & ~n50657;
  assign n50695 = i_hbusreq4 & ~n50655;
  assign n50696 = i_hbusreq9 & ~n50655;
  assign n50697 = i_hbusreq3 & ~n50653;
  assign n50698 = i_hbusreq1 & ~n50651;
  assign n50699 = i_hbusreq2 & ~n50636;
  assign n50700 = i_hbusreq0 & ~n50636;
  assign n50701 = ~controllable_locked & ~n46582;
  assign n50702 = ~controllable_locked & ~n50701;
  assign n50703 = i_hlock0 & ~n50702;
  assign n50704 = ~i_hlock0 & ~n50636;
  assign n50705 = ~n50703 & ~n50704;
  assign n50706 = ~i_hbusreq0 & ~n50705;
  assign n50707 = ~n50700 & ~n50706;
  assign n50708 = ~i_hbusreq2 & ~n50707;
  assign n50709 = ~n50699 & ~n50708;
  assign n50710 = controllable_hgrant2 & ~n50709;
  assign n50711 = controllable_hgrant2 & ~n50710;
  assign n50712 = ~n7733 & ~n50711;
  assign n50713 = i_hbusreq2 & ~n50645;
  assign n50714 = i_hbusreq0 & ~n50641;
  assign n50715 = ~i_hbusreq0 & ~n50643;
  assign n50716 = ~n50714 & ~n50715;
  assign n50717 = i_hlock2 & ~n50716;
  assign n50718 = ~n50644 & ~n50717;
  assign n50719 = ~i_hbusreq2 & ~n50718;
  assign n50720 = ~n50713 & ~n50719;
  assign n50721 = controllable_hgrant2 & ~n50720;
  assign n50722 = controllable_hgrant2 & ~n50721;
  assign n50723 = n7733 & ~n50722;
  assign n50724 = ~n50712 & ~n50723;
  assign n50725 = n7928 & ~n50724;
  assign n50726 = n7928 & ~n50725;
  assign n50727 = ~i_hbusreq1 & ~n50726;
  assign n50728 = ~n50698 & ~n50727;
  assign n50729 = ~controllable_hgrant1 & ~n50728;
  assign n50730 = ~controllable_hgrant1 & ~n50729;
  assign n50731 = ~i_hbusreq3 & ~n50730;
  assign n50732 = ~n50697 & ~n50731;
  assign n50733 = ~controllable_hgrant3 & ~n50732;
  assign n50734 = ~controllable_hgrant3 & ~n50733;
  assign n50735 = ~i_hbusreq9 & ~n50734;
  assign n50736 = ~n50696 & ~n50735;
  assign n50737 = ~i_hbusreq4 & ~n50736;
  assign n50738 = ~n50695 & ~n50737;
  assign n50739 = ~controllable_hgrant4 & ~n50738;
  assign n50740 = ~controllable_hgrant4 & ~n50739;
  assign n50741 = ~i_hbusreq5 & ~n50740;
  assign n50742 = ~n50694 & ~n50741;
  assign n50743 = ~controllable_hgrant5 & ~n50742;
  assign n50744 = ~controllable_hgrant5 & ~n50743;
  assign n50745 = ~i_hbusreq6 & ~n50744;
  assign n50746 = ~n50693 & ~n50745;
  assign n50747 = ~controllable_hgrant6 & ~n50746;
  assign n50748 = ~controllable_hgrant6 & ~n50747;
  assign n50749 = ~i_hbusreq8 & ~n50748;
  assign n50750 = ~n50692 & ~n50749;
  assign n50751 = controllable_hmaster3 & ~n50750;
  assign n50752 = i_hbusreq8 & ~n50688;
  assign n50753 = controllable_hmaster0 & ~n50748;
  assign n50754 = i_hbusreq6 & ~n50684;
  assign n50755 = controllable_hmaster2 & ~n50744;
  assign n50756 = i_hbusreq5 & ~n50677;
  assign n50757 = i_hbusreq4 & ~n50675;
  assign n50758 = i_hbusreq9 & ~n50675;
  assign n50759 = i_hbusreq3 & ~n50673;
  assign n50760 = i_hbusreq1 & ~n50671;
  assign n50761 = ~n18216 & ~n44750;
  assign n50762 = ~n7733 & ~n50761;
  assign n50763 = ~n40355 & ~n49770;
  assign n50764 = n7733 & ~n50763;
  assign n50765 = ~n50762 & ~n50764;
  assign n50766 = n7928 & ~n50765;
  assign n50767 = ~n43545 & ~n50766;
  assign n50768 = ~i_hbusreq1 & ~n50767;
  assign n50769 = ~n50760 & ~n50768;
  assign n50770 = ~controllable_hgrant1 & ~n50769;
  assign n50771 = ~n48564 & ~n50770;
  assign n50772 = ~i_hbusreq3 & ~n50771;
  assign n50773 = ~n50759 & ~n50772;
  assign n50774 = ~controllable_hgrant3 & ~n50773;
  assign n50775 = ~n48556 & ~n50774;
  assign n50776 = ~i_hbusreq9 & ~n50775;
  assign n50777 = ~n50758 & ~n50776;
  assign n50778 = ~i_hbusreq4 & ~n50777;
  assign n50779 = ~n50757 & ~n50778;
  assign n50780 = ~controllable_hgrant4 & ~n50779;
  assign n50781 = ~n48547 & ~n50780;
  assign n50782 = ~i_hbusreq5 & ~n50781;
  assign n50783 = ~n50756 & ~n50782;
  assign n50784 = ~controllable_hgrant5 & ~n50783;
  assign n50785 = ~n48536 & ~n50784;
  assign n50786 = ~controllable_hmaster2 & ~n50785;
  assign n50787 = ~n50755 & ~n50786;
  assign n50788 = controllable_hmaster1 & ~n50787;
  assign n50789 = ~controllable_hmaster1 & ~n50744;
  assign n50790 = ~n50788 & ~n50789;
  assign n50791 = ~i_hbusreq6 & ~n50790;
  assign n50792 = ~n50754 & ~n50791;
  assign n50793 = ~controllable_hgrant6 & ~n50792;
  assign n50794 = ~n50616 & ~n50793;
  assign n50795 = ~controllable_hmaster0 & ~n50794;
  assign n50796 = ~n50753 & ~n50795;
  assign n50797 = ~i_hbusreq8 & ~n50796;
  assign n50798 = ~n50752 & ~n50797;
  assign n50799 = ~controllable_hmaster3 & ~n50798;
  assign n50800 = ~n50751 & ~n50799;
  assign n50801 = ~i_hbusreq7 & ~n50800;
  assign n50802 = ~n50691 & ~n50801;
  assign n50803 = n7924 & ~n50802;
  assign n50804 = ~n50633 & ~n50803;
  assign n50805 = n8214 & ~n50804;
  assign n50806 = ~n50594 & ~n50805;
  assign n50807 = n8202 & ~n50806;
  assign n50808 = ~n50446 & ~n50807;
  assign n50809 = n7920 & ~n50808;
  assign n50810 = ~n50196 & ~n50809;
  assign n50811 = n7728 & ~n50810;
  assign n50812 = ~n7920 & ~n50178;
  assign n50813 = ~n7737 & n8378;
  assign n50814 = ~n8378 & ~n17007;
  assign n50815 = ~n50813 & ~n50814;
  assign n50816 = controllable_hgrant5 & ~n50815;
  assign n50817 = ~n7948 & ~n50816;
  assign n50818 = controllable_hmaster1 & ~n50817;
  assign n50819 = controllable_hmaster2 & ~n50817;
  assign n50820 = controllable_hmaster2 & ~n50819;
  assign n50821 = ~controllable_hmaster1 & ~n50820;
  assign n50822 = ~n50818 & ~n50821;
  assign n50823 = ~controllable_hgrant6 & ~n50822;
  assign n50824 = ~n7809 & ~n50823;
  assign n50825 = controllable_hmaster3 & ~n50824;
  assign n50826 = ~n50208 & ~n50825;
  assign n50827 = i_hbusreq7 & ~n50826;
  assign n50828 = i_hbusreq8 & ~n50824;
  assign n50829 = i_hbusreq6 & ~n50822;
  assign n50830 = i_hbusreq5 & ~n50815;
  assign n50831 = ~n7767 & n8378;
  assign n50832 = ~n8378 & ~n17056;
  assign n50833 = ~n50831 & ~n50832;
  assign n50834 = ~i_hbusreq5 & ~n50833;
  assign n50835 = ~n50830 & ~n50834;
  assign n50836 = controllable_hgrant5 & ~n50835;
  assign n50837 = ~n8005 & ~n50836;
  assign n50838 = controllable_hmaster1 & ~n50837;
  assign n50839 = controllable_hmaster2 & ~n50837;
  assign n50840 = controllable_hmaster2 & ~n50839;
  assign n50841 = ~controllable_hmaster1 & ~n50840;
  assign n50842 = ~n50838 & ~n50841;
  assign n50843 = ~i_hbusreq6 & ~n50842;
  assign n50844 = ~n50829 & ~n50843;
  assign n50845 = ~controllable_hgrant6 & ~n50844;
  assign n50846 = ~n7844 & ~n50845;
  assign n50847 = ~i_hbusreq8 & ~n50846;
  assign n50848 = ~n50828 & ~n50847;
  assign n50849 = controllable_hmaster3 & ~n50848;
  assign n50850 = ~n50231 & ~n50849;
  assign n50851 = ~i_hbusreq7 & ~n50850;
  assign n50852 = ~n50827 & ~n50851;
  assign n50853 = ~n7924 & ~n50852;
  assign n50854 = n8378 & ~n13021;
  assign n50855 = ~n8378 & ~n29186;
  assign n50856 = ~n50854 & ~n50855;
  assign n50857 = i_hlock5 & ~n50856;
  assign n50858 = ~n8378 & ~n29200;
  assign n50859 = ~n50854 & ~n50858;
  assign n50860 = ~i_hlock5 & ~n50859;
  assign n50861 = ~n50857 & ~n50860;
  assign n50862 = controllable_hgrant5 & ~n50861;
  assign n50863 = ~n8033 & ~n50862;
  assign n50864 = controllable_hmaster1 & ~n50863;
  assign n50865 = controllable_hmaster2 & ~n50863;
  assign n50866 = ~n8049 & ~n50244;
  assign n50867 = ~controllable_hmaster2 & ~n50866;
  assign n50868 = ~n50865 & ~n50867;
  assign n50869 = ~controllable_hmaster1 & ~n50868;
  assign n50870 = ~n50864 & ~n50869;
  assign n50871 = ~controllable_hgrant6 & ~n50870;
  assign n50872 = ~n7809 & ~n50871;
  assign n50873 = controllable_hmaster3 & ~n50872;
  assign n50874 = controllable_hmaster1 & ~n50866;
  assign n50875 = i_hlock5 & ~n41011;
  assign n50876 = ~i_hlock5 & ~n41024;
  assign n50877 = ~n50875 & ~n50876;
  assign n50878 = ~controllable_hgrant5 & ~n50877;
  assign n50879 = ~n48879 & ~n50878;
  assign n50880 = controllable_hmaster2 & ~n50879;
  assign n50881 = ~n50867 & ~n50880;
  assign n50882 = ~controllable_hmaster1 & ~n50881;
  assign n50883 = ~n50874 & ~n50882;
  assign n50884 = ~controllable_hgrant6 & ~n50883;
  assign n50885 = ~n50200 & ~n50884;
  assign n50886 = controllable_hmaster0 & ~n50885;
  assign n50887 = ~controllable_hgrant6 & ~n50866;
  assign n50888 = ~controllable_hgrant6 & ~n50887;
  assign n50889 = ~controllable_hmaster0 & ~n50888;
  assign n50890 = ~n50886 & ~n50889;
  assign n50891 = ~controllable_hmaster3 & ~n50890;
  assign n50892 = ~n50873 & ~n50891;
  assign n50893 = i_hbusreq7 & ~n50892;
  assign n50894 = i_hbusreq8 & ~n50872;
  assign n50895 = i_hbusreq6 & ~n50870;
  assign n50896 = i_hbusreq5 & ~n50861;
  assign n50897 = n8378 & ~n13075;
  assign n50898 = ~n8378 & ~n29225;
  assign n50899 = ~n50897 & ~n50898;
  assign n50900 = i_hlock5 & ~n50899;
  assign n50901 = ~n8378 & ~n29254;
  assign n50902 = ~n50897 & ~n50901;
  assign n50903 = ~i_hlock5 & ~n50902;
  assign n50904 = ~n50900 & ~n50903;
  assign n50905 = ~i_hbusreq5 & ~n50904;
  assign n50906 = ~n50896 & ~n50905;
  assign n50907 = controllable_hgrant5 & ~n50906;
  assign n50908 = ~n8096 & ~n50907;
  assign n50909 = controllable_hmaster1 & ~n50908;
  assign n50910 = controllable_hmaster2 & ~n50908;
  assign n50911 = ~n8133 & ~n50277;
  assign n50912 = ~controllable_hmaster2 & ~n50911;
  assign n50913 = ~n50910 & ~n50912;
  assign n50914 = ~controllable_hmaster1 & ~n50913;
  assign n50915 = ~n50909 & ~n50914;
  assign n50916 = ~i_hbusreq6 & ~n50915;
  assign n50917 = ~n50895 & ~n50916;
  assign n50918 = ~controllable_hgrant6 & ~n50917;
  assign n50919 = ~n7844 & ~n50918;
  assign n50920 = ~i_hbusreq8 & ~n50919;
  assign n50921 = ~n50894 & ~n50920;
  assign n50922 = controllable_hmaster3 & ~n50921;
  assign n50923 = i_hbusreq8 & ~n50890;
  assign n50924 = i_hbusreq6 & ~n50883;
  assign n50925 = controllable_hmaster1 & ~n50911;
  assign n50926 = i_hbusreq5 & ~n50877;
  assign n50927 = i_hlock5 & ~n41051;
  assign n50928 = ~i_hlock5 & ~n41076;
  assign n50929 = ~n50927 & ~n50928;
  assign n50930 = ~i_hbusreq5 & ~n50929;
  assign n50931 = ~n50926 & ~n50930;
  assign n50932 = ~controllable_hgrant5 & ~n50931;
  assign n50933 = ~n49568 & ~n50932;
  assign n50934 = controllable_hmaster2 & ~n50933;
  assign n50935 = ~n50912 & ~n50934;
  assign n50936 = ~controllable_hmaster1 & ~n50935;
  assign n50937 = ~n50925 & ~n50936;
  assign n50938 = ~i_hbusreq6 & ~n50937;
  assign n50939 = ~n50924 & ~n50938;
  assign n50940 = ~controllable_hgrant6 & ~n50939;
  assign n50941 = ~n50218 & ~n50940;
  assign n50942 = controllable_hmaster0 & ~n50941;
  assign n50943 = i_hbusreq6 & ~n50866;
  assign n50944 = ~i_hbusreq6 & ~n50911;
  assign n50945 = ~n50943 & ~n50944;
  assign n50946 = ~controllable_hgrant6 & ~n50945;
  assign n50947 = ~controllable_hgrant6 & ~n50946;
  assign n50948 = ~controllable_hmaster0 & ~n50947;
  assign n50949 = ~n50942 & ~n50948;
  assign n50950 = ~i_hbusreq8 & ~n50949;
  assign n50951 = ~n50923 & ~n50950;
  assign n50952 = ~controllable_hmaster3 & ~n50951;
  assign n50953 = ~n50922 & ~n50952;
  assign n50954 = ~i_hbusreq7 & ~n50953;
  assign n50955 = ~n50893 & ~n50954;
  assign n50956 = n7924 & ~n50955;
  assign n50957 = ~n50853 & ~n50956;
  assign n50958 = ~n8214 & ~n50957;
  assign n50959 = ~n7737 & n8426;
  assign n50960 = ~n8426 & ~n17005;
  assign n50961 = ~n50959 & ~n50960;
  assign n50962 = controllable_hgrant4 & ~n50961;
  assign n50963 = ~n7946 & ~n50962;
  assign n50964 = ~controllable_hgrant5 & ~n50963;
  assign n50965 = ~n7810 & ~n50964;
  assign n50966 = controllable_hmaster1 & ~n50965;
  assign n50967 = controllable_hmaster2 & ~n50965;
  assign n50968 = controllable_hmaster2 & ~n50967;
  assign n50969 = ~controllable_hmaster1 & ~n50968;
  assign n50970 = ~n50966 & ~n50969;
  assign n50971 = ~controllable_hgrant6 & ~n50970;
  assign n50972 = ~n7809 & ~n50971;
  assign n50973 = controllable_hmaster3 & ~n50972;
  assign n50974 = ~n50322 & ~n50973;
  assign n50975 = i_hbusreq7 & ~n50974;
  assign n50976 = i_hbusreq8 & ~n50972;
  assign n50977 = i_hbusreq6 & ~n50970;
  assign n50978 = i_hbusreq5 & ~n50963;
  assign n50979 = i_hbusreq4 & ~n50961;
  assign n50980 = i_hbusreq9 & ~n50961;
  assign n50981 = ~n7763 & n8426;
  assign n50982 = ~n8426 & ~n17050;
  assign n50983 = ~n50981 & ~n50982;
  assign n50984 = ~i_hbusreq9 & ~n50983;
  assign n50985 = ~n50980 & ~n50984;
  assign n50986 = ~i_hbusreq4 & ~n50985;
  assign n50987 = ~n50979 & ~n50986;
  assign n50988 = controllable_hgrant4 & ~n50987;
  assign n50989 = ~n8001 & ~n50988;
  assign n50990 = ~i_hbusreq5 & ~n50989;
  assign n50991 = ~n50978 & ~n50990;
  assign n50992 = ~controllable_hgrant5 & ~n50991;
  assign n50993 = ~n7846 & ~n50992;
  assign n50994 = controllable_hmaster1 & ~n50993;
  assign n50995 = controllable_hmaster2 & ~n50993;
  assign n50996 = controllable_hmaster2 & ~n50995;
  assign n50997 = ~controllable_hmaster1 & ~n50996;
  assign n50998 = ~n50994 & ~n50997;
  assign n50999 = ~i_hbusreq6 & ~n50998;
  assign n51000 = ~n50977 & ~n50999;
  assign n51001 = ~controllable_hgrant6 & ~n51000;
  assign n51002 = ~n7844 & ~n51001;
  assign n51003 = ~i_hbusreq8 & ~n51002;
  assign n51004 = ~n50976 & ~n51003;
  assign n51005 = controllable_hmaster3 & ~n51004;
  assign n51006 = ~n50345 & ~n51005;
  assign n51007 = ~i_hbusreq7 & ~n51006;
  assign n51008 = ~n50975 & ~n51007;
  assign n51009 = ~n7924 & ~n51008;
  assign n51010 = n8426 & ~n13019;
  assign n51011 = ~n8426 & ~n17099;
  assign n51012 = ~n51010 & ~n51011;
  assign n51013 = i_hlock4 & ~n51012;
  assign n51014 = ~n8426 & ~n17107;
  assign n51015 = ~n51010 & ~n51014;
  assign n51016 = ~i_hlock4 & ~n51015;
  assign n51017 = ~n51013 & ~n51016;
  assign n51018 = controllable_hgrant4 & ~n51017;
  assign n51019 = ~n8031 & ~n51018;
  assign n51020 = ~controllable_hgrant5 & ~n51019;
  assign n51021 = ~n7810 & ~n51020;
  assign n51022 = controllable_hmaster1 & ~n51021;
  assign n51023 = controllable_hmaster2 & ~n51021;
  assign n51024 = ~n8047 & ~n50358;
  assign n51025 = ~controllable_hgrant5 & ~n51024;
  assign n51026 = ~controllable_hgrant5 & ~n51025;
  assign n51027 = ~controllable_hmaster2 & ~n51026;
  assign n51028 = ~n51023 & ~n51027;
  assign n51029 = ~controllable_hmaster1 & ~n51028;
  assign n51030 = ~n51022 & ~n51029;
  assign n51031 = ~controllable_hgrant6 & ~n51030;
  assign n51032 = ~n7809 & ~n51031;
  assign n51033 = controllable_hmaster3 & ~n51032;
  assign n51034 = ~controllable_hgrant6 & ~n51026;
  assign n51035 = ~controllable_hgrant6 & ~n51034;
  assign n51036 = controllable_hmaster0 & ~n51035;
  assign n51037 = controllable_hmaster1 & ~n51026;
  assign n51038 = i_hlock4 & ~n40837;
  assign n51039 = ~i_hlock4 & ~n40843;
  assign n51040 = ~n51038 & ~n51039;
  assign n51041 = ~controllable_hgrant4 & ~n51040;
  assign n51042 = ~n49009 & ~n51041;
  assign n51043 = ~controllable_hgrant5 & ~n51042;
  assign n51044 = ~n48169 & ~n51043;
  assign n51045 = controllable_hmaster2 & ~n51044;
  assign n51046 = ~n51027 & ~n51045;
  assign n51047 = ~controllable_hmaster1 & ~n51046;
  assign n51048 = ~n51037 & ~n51047;
  assign n51049 = ~controllable_hgrant6 & ~n51048;
  assign n51050 = ~n50314 & ~n51049;
  assign n51051 = ~controllable_hmaster0 & ~n51050;
  assign n51052 = ~n51036 & ~n51051;
  assign n51053 = ~controllable_hmaster3 & ~n51052;
  assign n51054 = ~n51033 & ~n51053;
  assign n51055 = i_hbusreq7 & ~n51054;
  assign n51056 = i_hbusreq8 & ~n51032;
  assign n51057 = i_hbusreq6 & ~n51030;
  assign n51058 = i_hbusreq5 & ~n51019;
  assign n51059 = i_hbusreq4 & ~n51017;
  assign n51060 = i_hbusreq9 & ~n51012;
  assign n51061 = n8426 & ~n13069;
  assign n51062 = ~n8426 & ~n17168;
  assign n51063 = ~n51061 & ~n51062;
  assign n51064 = ~i_hbusreq9 & ~n51063;
  assign n51065 = ~n51060 & ~n51064;
  assign n51066 = i_hlock4 & ~n51065;
  assign n51067 = i_hbusreq9 & ~n51015;
  assign n51068 = ~n8426 & ~n17182;
  assign n51069 = ~n51061 & ~n51068;
  assign n51070 = ~i_hbusreq9 & ~n51069;
  assign n51071 = ~n51067 & ~n51070;
  assign n51072 = ~i_hlock4 & ~n51071;
  assign n51073 = ~n51066 & ~n51072;
  assign n51074 = ~i_hbusreq4 & ~n51073;
  assign n51075 = ~n51059 & ~n51074;
  assign n51076 = controllable_hgrant4 & ~n51075;
  assign n51077 = ~n8092 & ~n51076;
  assign n51078 = ~i_hbusreq5 & ~n51077;
  assign n51079 = ~n51058 & ~n51078;
  assign n51080 = ~controllable_hgrant5 & ~n51079;
  assign n51081 = ~n7846 & ~n51080;
  assign n51082 = controllable_hmaster1 & ~n51081;
  assign n51083 = controllable_hmaster2 & ~n51081;
  assign n51084 = i_hbusreq5 & ~n51024;
  assign n51085 = ~n8129 & ~n50402;
  assign n51086 = ~i_hbusreq5 & ~n51085;
  assign n51087 = ~n51084 & ~n51086;
  assign n51088 = ~controllable_hgrant5 & ~n51087;
  assign n51089 = ~controllable_hgrant5 & ~n51088;
  assign n51090 = ~controllable_hmaster2 & ~n51089;
  assign n51091 = ~n51083 & ~n51090;
  assign n51092 = ~controllable_hmaster1 & ~n51091;
  assign n51093 = ~n51082 & ~n51092;
  assign n51094 = ~i_hbusreq6 & ~n51093;
  assign n51095 = ~n51057 & ~n51094;
  assign n51096 = ~controllable_hgrant6 & ~n51095;
  assign n51097 = ~n7844 & ~n51096;
  assign n51098 = ~i_hbusreq8 & ~n51097;
  assign n51099 = ~n51056 & ~n51098;
  assign n51100 = controllable_hmaster3 & ~n51099;
  assign n51101 = i_hbusreq8 & ~n51052;
  assign n51102 = i_hbusreq6 & ~n51026;
  assign n51103 = ~i_hbusreq6 & ~n51089;
  assign n51104 = ~n51102 & ~n51103;
  assign n51105 = ~controllable_hgrant6 & ~n51104;
  assign n51106 = ~controllable_hgrant6 & ~n51105;
  assign n51107 = controllable_hmaster0 & ~n51106;
  assign n51108 = i_hbusreq6 & ~n51048;
  assign n51109 = controllable_hmaster1 & ~n51089;
  assign n51110 = i_hbusreq5 & ~n51042;
  assign n51111 = i_hbusreq4 & ~n51040;
  assign n51112 = i_hlock4 & ~n41047;
  assign n51113 = ~i_hlock4 & ~n41072;
  assign n51114 = ~n51112 & ~n51113;
  assign n51115 = ~i_hbusreq4 & ~n51114;
  assign n51116 = ~n51111 & ~n51115;
  assign n51117 = ~controllable_hgrant4 & ~n51116;
  assign n51118 = ~n49828 & ~n51117;
  assign n51119 = ~i_hbusreq5 & ~n51118;
  assign n51120 = ~n51110 & ~n51119;
  assign n51121 = ~controllable_hgrant5 & ~n51120;
  assign n51122 = ~n48615 & ~n51121;
  assign n51123 = controllable_hmaster2 & ~n51122;
  assign n51124 = ~n51090 & ~n51123;
  assign n51125 = ~controllable_hmaster1 & ~n51124;
  assign n51126 = ~n51109 & ~n51125;
  assign n51127 = ~i_hbusreq6 & ~n51126;
  assign n51128 = ~n51108 & ~n51127;
  assign n51129 = ~controllable_hgrant6 & ~n51128;
  assign n51130 = ~n50332 & ~n51129;
  assign n51131 = ~controllable_hmaster0 & ~n51130;
  assign n51132 = ~n51107 & ~n51131;
  assign n51133 = ~i_hbusreq8 & ~n51132;
  assign n51134 = ~n51101 & ~n51133;
  assign n51135 = ~controllable_hmaster3 & ~n51134;
  assign n51136 = ~n51100 & ~n51135;
  assign n51137 = ~i_hbusreq7 & ~n51136;
  assign n51138 = ~n51055 & ~n51137;
  assign n51139 = n7924 & ~n51138;
  assign n51140 = ~n51009 & ~n51139;
  assign n51141 = n8214 & ~n51140;
  assign n51142 = ~n50958 & ~n51141;
  assign n51143 = ~n8202 & ~n51142;
  assign n51144 = ~n7737 & n8365;
  assign n51145 = ~n8365 & ~n17003;
  assign n51146 = ~n51144 & ~n51145;
  assign n51147 = controllable_hgrant3 & ~n51146;
  assign n51148 = ~n7944 & ~n51147;
  assign n51149 = ~controllable_hgrant4 & ~n51148;
  assign n51150 = ~n7811 & ~n51149;
  assign n51151 = ~controllable_hgrant5 & ~n51150;
  assign n51152 = ~n7810 & ~n51151;
  assign n51153 = controllable_hmaster1 & ~n51152;
  assign n51154 = controllable_hmaster2 & ~n51152;
  assign n51155 = controllable_hmaster2 & ~n51154;
  assign n51156 = ~controllable_hmaster1 & ~n51155;
  assign n51157 = ~n51153 & ~n51156;
  assign n51158 = ~controllable_hgrant6 & ~n51157;
  assign n51159 = ~n7809 & ~n51158;
  assign n51160 = controllable_hmaster3 & ~n51159;
  assign n51161 = ~n50458 & ~n51160;
  assign n51162 = i_hbusreq7 & ~n51161;
  assign n51163 = i_hbusreq8 & ~n51159;
  assign n51164 = i_hbusreq6 & ~n51157;
  assign n51165 = i_hbusreq5 & ~n51150;
  assign n51166 = i_hbusreq4 & ~n51148;
  assign n51167 = i_hbusreq9 & ~n51148;
  assign n51168 = i_hbusreq3 & ~n51146;
  assign n51169 = ~n7761 & n8365;
  assign n51170 = ~n8365 & ~n17046;
  assign n51171 = ~n51169 & ~n51170;
  assign n51172 = ~i_hbusreq3 & ~n51171;
  assign n51173 = ~n51168 & ~n51172;
  assign n51174 = controllable_hgrant3 & ~n51173;
  assign n51175 = ~n7995 & ~n51174;
  assign n51176 = ~i_hbusreq9 & ~n51175;
  assign n51177 = ~n51167 & ~n51176;
  assign n51178 = ~i_hbusreq4 & ~n51177;
  assign n51179 = ~n51166 & ~n51178;
  assign n51180 = ~controllable_hgrant4 & ~n51179;
  assign n51181 = ~n7848 & ~n51180;
  assign n51182 = ~i_hbusreq5 & ~n51181;
  assign n51183 = ~n51165 & ~n51182;
  assign n51184 = ~controllable_hgrant5 & ~n51183;
  assign n51185 = ~n7846 & ~n51184;
  assign n51186 = controllable_hmaster1 & ~n51185;
  assign n51187 = controllable_hmaster2 & ~n51185;
  assign n51188 = controllable_hmaster2 & ~n51187;
  assign n51189 = ~controllable_hmaster1 & ~n51188;
  assign n51190 = ~n51186 & ~n51189;
  assign n51191 = ~i_hbusreq6 & ~n51190;
  assign n51192 = ~n51164 & ~n51191;
  assign n51193 = ~controllable_hgrant6 & ~n51192;
  assign n51194 = ~n7844 & ~n51193;
  assign n51195 = ~i_hbusreq8 & ~n51194;
  assign n51196 = ~n51163 & ~n51195;
  assign n51197 = controllable_hmaster3 & ~n51196;
  assign n51198 = ~n50481 & ~n51197;
  assign n51199 = ~i_hbusreq7 & ~n51198;
  assign n51200 = ~n51162 & ~n51199;
  assign n51201 = ~n7924 & ~n51200;
  assign n51202 = n8365 & ~n13017;
  assign n51203 = ~n8365 & ~n17097;
  assign n51204 = ~n51202 & ~n51203;
  assign n51205 = i_hlock3 & ~n51204;
  assign n51206 = ~n8365 & ~n17105;
  assign n51207 = ~n51202 & ~n51206;
  assign n51208 = ~i_hlock3 & ~n51207;
  assign n51209 = ~n51205 & ~n51208;
  assign n51210 = controllable_hgrant3 & ~n51209;
  assign n51211 = ~n8029 & ~n51210;
  assign n51212 = ~controllable_hgrant4 & ~n51211;
  assign n51213 = ~n7811 & ~n51212;
  assign n51214 = ~controllable_hgrant5 & ~n51213;
  assign n51215 = ~n7810 & ~n51214;
  assign n51216 = controllable_hmaster1 & ~n51215;
  assign n51217 = controllable_hmaster2 & ~n51215;
  assign n51218 = ~n8045 & ~n50494;
  assign n51219 = ~controllable_hgrant4 & ~n51218;
  assign n51220 = ~controllable_hgrant4 & ~n51219;
  assign n51221 = ~controllable_hgrant5 & ~n51220;
  assign n51222 = ~controllable_hgrant5 & ~n51221;
  assign n51223 = ~controllable_hmaster2 & ~n51222;
  assign n51224 = ~n51217 & ~n51223;
  assign n51225 = ~controllable_hmaster1 & ~n51224;
  assign n51226 = ~n51216 & ~n51225;
  assign n51227 = ~controllable_hgrant6 & ~n51226;
  assign n51228 = ~n7809 & ~n51227;
  assign n51229 = controllable_hmaster3 & ~n51228;
  assign n51230 = controllable_hmaster2 & ~n51222;
  assign n51231 = i_hlock3 & ~n40835;
  assign n51232 = ~i_hlock3 & ~n40841;
  assign n51233 = ~n51231 & ~n51232;
  assign n51234 = ~controllable_hgrant3 & ~n51233;
  assign n51235 = ~n48859 & ~n51234;
  assign n51236 = ~controllable_hgrant4 & ~n51235;
  assign n51237 = ~n48063 & ~n51236;
  assign n51238 = ~controllable_hgrant5 & ~n51237;
  assign n51239 = ~n48060 & ~n51238;
  assign n51240 = ~controllable_hmaster2 & ~n51239;
  assign n51241 = ~n51230 & ~n51240;
  assign n51242 = controllable_hmaster1 & ~n51241;
  assign n51243 = ~controllable_hmaster1 & ~n51222;
  assign n51244 = ~n51242 & ~n51243;
  assign n51245 = ~controllable_hgrant6 & ~n51244;
  assign n51246 = ~n50450 & ~n51245;
  assign n51247 = controllable_hmaster0 & ~n51246;
  assign n51248 = ~controllable_hgrant6 & ~n51222;
  assign n51249 = ~controllable_hgrant6 & ~n51248;
  assign n51250 = ~controllable_hmaster0 & ~n51249;
  assign n51251 = ~n51247 & ~n51250;
  assign n51252 = ~controllable_hmaster3 & ~n51251;
  assign n51253 = ~n51229 & ~n51252;
  assign n51254 = i_hbusreq7 & ~n51253;
  assign n51255 = i_hbusreq8 & ~n51228;
  assign n51256 = i_hbusreq6 & ~n51226;
  assign n51257 = i_hbusreq5 & ~n51213;
  assign n51258 = i_hbusreq4 & ~n51211;
  assign n51259 = i_hbusreq9 & ~n51211;
  assign n51260 = i_hbusreq3 & ~n51209;
  assign n51261 = n8365 & ~n13065;
  assign n51262 = ~n8365 & ~n17164;
  assign n51263 = ~n51261 & ~n51262;
  assign n51264 = i_hlock3 & ~n51263;
  assign n51265 = ~n8365 & ~n17178;
  assign n51266 = ~n51261 & ~n51265;
  assign n51267 = ~i_hlock3 & ~n51266;
  assign n51268 = ~n51264 & ~n51267;
  assign n51269 = ~i_hbusreq3 & ~n51268;
  assign n51270 = ~n51260 & ~n51269;
  assign n51271 = controllable_hgrant3 & ~n51270;
  assign n51272 = ~n8086 & ~n51271;
  assign n51273 = ~i_hbusreq9 & ~n51272;
  assign n51274 = ~n51259 & ~n51273;
  assign n51275 = ~i_hbusreq4 & ~n51274;
  assign n51276 = ~n51258 & ~n51275;
  assign n51277 = ~controllable_hgrant4 & ~n51276;
  assign n51278 = ~n7848 & ~n51277;
  assign n51279 = ~i_hbusreq5 & ~n51278;
  assign n51280 = ~n51257 & ~n51279;
  assign n51281 = ~controllable_hgrant5 & ~n51280;
  assign n51282 = ~n7846 & ~n51281;
  assign n51283 = controllable_hmaster1 & ~n51282;
  assign n51284 = controllable_hmaster2 & ~n51282;
  assign n51285 = i_hbusreq5 & ~n51220;
  assign n51286 = i_hbusreq4 & ~n51218;
  assign n51287 = i_hbusreq9 & ~n51218;
  assign n51288 = ~n8123 & ~n50538;
  assign n51289 = ~i_hbusreq9 & ~n51288;
  assign n51290 = ~n51287 & ~n51289;
  assign n51291 = ~i_hbusreq4 & ~n51290;
  assign n51292 = ~n51286 & ~n51291;
  assign n51293 = ~controllable_hgrant4 & ~n51292;
  assign n51294 = ~controllable_hgrant4 & ~n51293;
  assign n51295 = ~i_hbusreq5 & ~n51294;
  assign n51296 = ~n51285 & ~n51295;
  assign n51297 = ~controllable_hgrant5 & ~n51296;
  assign n51298 = ~controllable_hgrant5 & ~n51297;
  assign n51299 = ~controllable_hmaster2 & ~n51298;
  assign n51300 = ~n51284 & ~n51299;
  assign n51301 = ~controllable_hmaster1 & ~n51300;
  assign n51302 = ~n51283 & ~n51301;
  assign n51303 = ~i_hbusreq6 & ~n51302;
  assign n51304 = ~n51256 & ~n51303;
  assign n51305 = ~controllable_hgrant6 & ~n51304;
  assign n51306 = ~n7844 & ~n51305;
  assign n51307 = ~i_hbusreq8 & ~n51306;
  assign n51308 = ~n51255 & ~n51307;
  assign n51309 = controllable_hmaster3 & ~n51308;
  assign n51310 = i_hbusreq8 & ~n51251;
  assign n51311 = i_hbusreq6 & ~n51244;
  assign n51312 = controllable_hmaster2 & ~n51298;
  assign n51313 = i_hbusreq5 & ~n51237;
  assign n51314 = i_hbusreq4 & ~n51235;
  assign n51315 = i_hbusreq9 & ~n51235;
  assign n51316 = i_hbusreq3 & ~n51233;
  assign n51317 = i_hlock3 & ~n40885;
  assign n51318 = ~i_hlock3 & ~n40897;
  assign n51319 = ~n51317 & ~n51318;
  assign n51320 = ~i_hbusreq3 & ~n51319;
  assign n51321 = ~n51316 & ~n51320;
  assign n51322 = ~controllable_hgrant3 & ~n51321;
  assign n51323 = ~n49534 & ~n51322;
  assign n51324 = ~i_hbusreq9 & ~n51323;
  assign n51325 = ~n51315 & ~n51324;
  assign n51326 = ~i_hbusreq4 & ~n51325;
  assign n51327 = ~n51314 & ~n51326;
  assign n51328 = ~controllable_hgrant4 & ~n51327;
  assign n51329 = ~n48374 & ~n51328;
  assign n51330 = ~i_hbusreq5 & ~n51329;
  assign n51331 = ~n51313 & ~n51330;
  assign n51332 = ~controllable_hgrant5 & ~n51331;
  assign n51333 = ~n48363 & ~n51332;
  assign n51334 = ~controllable_hmaster2 & ~n51333;
  assign n51335 = ~n51312 & ~n51334;
  assign n51336 = controllable_hmaster1 & ~n51335;
  assign n51337 = ~controllable_hmaster1 & ~n51298;
  assign n51338 = ~n51336 & ~n51337;
  assign n51339 = ~i_hbusreq6 & ~n51338;
  assign n51340 = ~n51311 & ~n51339;
  assign n51341 = ~controllable_hgrant6 & ~n51340;
  assign n51342 = ~n50468 & ~n51341;
  assign n51343 = controllable_hmaster0 & ~n51342;
  assign n51344 = i_hbusreq6 & ~n51222;
  assign n51345 = ~i_hbusreq6 & ~n51298;
  assign n51346 = ~n51344 & ~n51345;
  assign n51347 = ~controllable_hgrant6 & ~n51346;
  assign n51348 = ~controllable_hgrant6 & ~n51347;
  assign n51349 = ~controllable_hmaster0 & ~n51348;
  assign n51350 = ~n51343 & ~n51349;
  assign n51351 = ~i_hbusreq8 & ~n51350;
  assign n51352 = ~n51310 & ~n51351;
  assign n51353 = ~controllable_hmaster3 & ~n51352;
  assign n51354 = ~n51309 & ~n51353;
  assign n51355 = ~i_hbusreq7 & ~n51354;
  assign n51356 = ~n51254 & ~n51355;
  assign n51357 = n7924 & ~n51356;
  assign n51358 = ~n51201 & ~n51357;
  assign n51359 = ~n8214 & ~n51358;
  assign n51360 = ~n7821 & ~n48018;
  assign n51361 = ~n7733 & ~n51360;
  assign n51362 = ~n7733 & ~n51361;
  assign n51363 = ~n7928 & ~n51362;
  assign n51364 = ~n7733 & ~n48020;
  assign n51365 = n7928 & ~n51364;
  assign n51366 = ~n51363 & ~n51365;
  assign n51367 = ~controllable_hgrant1 & ~n51366;
  assign n51368 = ~n7813 & ~n51367;
  assign n51369 = ~controllable_hgrant3 & ~n51368;
  assign n51370 = ~n7812 & ~n51369;
  assign n51371 = ~controllable_hgrant4 & ~n51370;
  assign n51372 = ~n7811 & ~n51371;
  assign n51373 = ~controllable_hgrant5 & ~n51372;
  assign n51374 = ~n7810 & ~n51373;
  assign n51375 = controllable_hmaster1 & ~n51374;
  assign n51376 = controllable_hmaster2 & ~n51374;
  assign n51377 = controllable_hmaster2 & ~n51376;
  assign n51378 = ~controllable_hmaster1 & ~n51377;
  assign n51379 = ~n51375 & ~n51378;
  assign n51380 = ~controllable_hgrant6 & ~n51379;
  assign n51381 = ~n7809 & ~n51380;
  assign n51382 = controllable_hmaster3 & ~n51381;
  assign n51383 = ~n50606 & ~n51382;
  assign n51384 = i_hbusreq7 & ~n51383;
  assign n51385 = i_hbusreq8 & ~n51381;
  assign n51386 = i_hbusreq6 & ~n51379;
  assign n51387 = i_hbusreq5 & ~n51372;
  assign n51388 = i_hbusreq4 & ~n51370;
  assign n51389 = i_hbusreq9 & ~n51370;
  assign n51390 = i_hbusreq3 & ~n51368;
  assign n51391 = i_hbusreq1 & ~n51366;
  assign n51392 = i_hbusreq2 & ~n40216;
  assign n51393 = i_hbusreq0 & ~n40216;
  assign n51394 = ~i_hbusreq0 & ~n40320;
  assign n51395 = ~n51393 & ~n51394;
  assign n51396 = ~i_hbusreq2 & ~n51395;
  assign n51397 = ~n51392 & ~n51396;
  assign n51398 = controllable_hgrant2 & ~n51397;
  assign n51399 = ~n7868 & ~n51398;
  assign n51400 = ~n7733 & ~n51399;
  assign n51401 = ~n7733 & ~n51400;
  assign n51402 = ~n7928 & ~n51401;
  assign n51403 = ~n7983 & ~n51398;
  assign n51404 = ~n7733 & ~n51403;
  assign n51405 = ~n7733 & ~n51404;
  assign n51406 = n7928 & ~n51405;
  assign n51407 = ~n51402 & ~n51406;
  assign n51408 = ~i_hbusreq1 & ~n51407;
  assign n51409 = ~n51391 & ~n51408;
  assign n51410 = ~controllable_hgrant1 & ~n51409;
  assign n51411 = ~n7853 & ~n51410;
  assign n51412 = ~i_hbusreq3 & ~n51411;
  assign n51413 = ~n51390 & ~n51412;
  assign n51414 = ~controllable_hgrant3 & ~n51413;
  assign n51415 = ~n7851 & ~n51414;
  assign n51416 = ~i_hbusreq9 & ~n51415;
  assign n51417 = ~n51389 & ~n51416;
  assign n51418 = ~i_hbusreq4 & ~n51417;
  assign n51419 = ~n51388 & ~n51418;
  assign n51420 = ~controllable_hgrant4 & ~n51419;
  assign n51421 = ~n7848 & ~n51420;
  assign n51422 = ~i_hbusreq5 & ~n51421;
  assign n51423 = ~n51387 & ~n51422;
  assign n51424 = ~controllable_hgrant5 & ~n51423;
  assign n51425 = ~n7846 & ~n51424;
  assign n51426 = controllable_hmaster1 & ~n51425;
  assign n51427 = controllable_hmaster2 & ~n51425;
  assign n51428 = controllable_hmaster2 & ~n51427;
  assign n51429 = ~controllable_hmaster1 & ~n51428;
  assign n51430 = ~n51426 & ~n51429;
  assign n51431 = ~i_hbusreq6 & ~n51430;
  assign n51432 = ~n51386 & ~n51431;
  assign n51433 = ~controllable_hgrant6 & ~n51432;
  assign n51434 = ~n7844 & ~n51433;
  assign n51435 = ~i_hbusreq8 & ~n51434;
  assign n51436 = ~n51385 & ~n51435;
  assign n51437 = controllable_hmaster3 & ~n51436;
  assign n51438 = ~n50629 & ~n51437;
  assign n51439 = ~i_hbusreq7 & ~n51438;
  assign n51440 = ~n51384 & ~n51439;
  assign n51441 = ~n7924 & ~n51440;
  assign n51442 = ~n48798 & ~n50648;
  assign n51443 = n7928 & ~n51442;
  assign n51444 = ~n51363 & ~n51443;
  assign n51445 = ~controllable_hgrant1 & ~n51444;
  assign n51446 = ~n7813 & ~n51445;
  assign n51447 = ~controllable_hgrant3 & ~n51446;
  assign n51448 = ~n7812 & ~n51447;
  assign n51449 = ~controllable_hgrant4 & ~n51448;
  assign n51450 = ~n7811 & ~n51449;
  assign n51451 = ~controllable_hgrant5 & ~n51450;
  assign n51452 = ~n7810 & ~n51451;
  assign n51453 = controllable_hmaster1 & ~n51452;
  assign n51454 = controllable_hmaster2 & ~n51452;
  assign n51455 = ~n8037 & ~n50637;
  assign n51456 = ~n7733 & ~n51455;
  assign n51457 = ~n50648 & ~n51456;
  assign n51458 = n7928 & ~n51457;
  assign n51459 = n7928 & ~n51458;
  assign n51460 = ~controllable_hgrant1 & ~n51459;
  assign n51461 = ~controllable_hgrant1 & ~n51460;
  assign n51462 = ~controllable_hgrant3 & ~n51461;
  assign n51463 = ~controllable_hgrant3 & ~n51462;
  assign n51464 = ~controllable_hgrant4 & ~n51463;
  assign n51465 = ~controllable_hgrant4 & ~n51464;
  assign n51466 = ~controllable_hgrant5 & ~n51465;
  assign n51467 = ~controllable_hgrant5 & ~n51466;
  assign n51468 = ~controllable_hmaster2 & ~n51467;
  assign n51469 = ~n51454 & ~n51468;
  assign n51470 = ~controllable_hmaster1 & ~n51469;
  assign n51471 = ~n51453 & ~n51470;
  assign n51472 = ~controllable_hgrant6 & ~n51471;
  assign n51473 = ~n7809 & ~n51472;
  assign n51474 = controllable_hmaster3 & ~n51473;
  assign n51475 = ~controllable_hgrant6 & ~n51467;
  assign n51476 = ~controllable_hgrant6 & ~n51475;
  assign n51477 = controllable_hmaster0 & ~n51476;
  assign n51478 = controllable_hmaster2 & ~n51467;
  assign n51479 = ~n48968 & ~n50668;
  assign n51480 = n7928 & ~n51479;
  assign n51481 = ~n42965 & ~n51480;
  assign n51482 = ~controllable_hgrant1 & ~n51481;
  assign n51483 = ~n48144 & ~n51482;
  assign n51484 = ~controllable_hgrant3 & ~n51483;
  assign n51485 = ~n48141 & ~n51484;
  assign n51486 = ~controllable_hgrant4 & ~n51485;
  assign n51487 = ~n48138 & ~n51486;
  assign n51488 = ~controllable_hgrant5 & ~n51487;
  assign n51489 = ~n48135 & ~n51488;
  assign n51490 = ~controllable_hmaster2 & ~n51489;
  assign n51491 = ~n51478 & ~n51490;
  assign n51492 = controllable_hmaster1 & ~n51491;
  assign n51493 = ~controllable_hmaster1 & ~n51467;
  assign n51494 = ~n51492 & ~n51493;
  assign n51495 = ~controllable_hgrant6 & ~n51494;
  assign n51496 = ~n50598 & ~n51495;
  assign n51497 = ~controllable_hmaster0 & ~n51496;
  assign n51498 = ~n51477 & ~n51497;
  assign n51499 = ~controllable_hmaster3 & ~n51498;
  assign n51500 = ~n51474 & ~n51499;
  assign n51501 = i_hbusreq7 & ~n51500;
  assign n51502 = i_hbusreq8 & ~n51473;
  assign n51503 = i_hbusreq6 & ~n51471;
  assign n51504 = i_hbusreq5 & ~n51450;
  assign n51505 = i_hbusreq4 & ~n51448;
  assign n51506 = i_hbusreq9 & ~n51448;
  assign n51507 = i_hbusreq3 & ~n51446;
  assign n51508 = i_hbusreq1 & ~n51444;
  assign n51509 = controllable_locked & ~n40320;
  assign n51510 = ~n44182 & ~n51509;
  assign n51511 = i_hlock0 & ~n51510;
  assign n51512 = ~controllable_locked & ~n49180;
  assign n51513 = ~n51509 & ~n51512;
  assign n51514 = ~i_hlock0 & ~n51513;
  assign n51515 = ~n51511 & ~n51514;
  assign n51516 = ~i_hbusreq0 & ~n51515;
  assign n51517 = ~n49162 & ~n51516;
  assign n51518 = ~i_hbusreq2 & ~n51517;
  assign n51519 = ~n49161 & ~n51518;
  assign n51520 = controllable_hgrant2 & ~n51519;
  assign n51521 = ~n8074 & ~n51520;
  assign n51522 = ~n7733 & ~n51521;
  assign n51523 = ~n50723 & ~n51522;
  assign n51524 = n7928 & ~n51523;
  assign n51525 = ~n51402 & ~n51524;
  assign n51526 = ~i_hbusreq1 & ~n51525;
  assign n51527 = ~n51508 & ~n51526;
  assign n51528 = ~controllable_hgrant1 & ~n51527;
  assign n51529 = ~n7853 & ~n51528;
  assign n51530 = ~i_hbusreq3 & ~n51529;
  assign n51531 = ~n51507 & ~n51530;
  assign n51532 = ~controllable_hgrant3 & ~n51531;
  assign n51533 = ~n7851 & ~n51532;
  assign n51534 = ~i_hbusreq9 & ~n51533;
  assign n51535 = ~n51506 & ~n51534;
  assign n51536 = ~i_hbusreq4 & ~n51535;
  assign n51537 = ~n51505 & ~n51536;
  assign n51538 = ~controllable_hgrant4 & ~n51537;
  assign n51539 = ~n7848 & ~n51538;
  assign n51540 = ~i_hbusreq5 & ~n51539;
  assign n51541 = ~n51504 & ~n51540;
  assign n51542 = ~controllable_hgrant5 & ~n51541;
  assign n51543 = ~n7846 & ~n51542;
  assign n51544 = controllable_hmaster1 & ~n51543;
  assign n51545 = controllable_hmaster2 & ~n51543;
  assign n51546 = i_hbusreq5 & ~n51465;
  assign n51547 = i_hbusreq4 & ~n51463;
  assign n51548 = i_hbusreq9 & ~n51463;
  assign n51549 = i_hbusreq3 & ~n51461;
  assign n51550 = i_hbusreq1 & ~n51459;
  assign n51551 = ~n8111 & ~n50710;
  assign n51552 = ~n7733 & ~n51551;
  assign n51553 = ~n50723 & ~n51552;
  assign n51554 = n7928 & ~n51553;
  assign n51555 = n7928 & ~n51554;
  assign n51556 = ~i_hbusreq1 & ~n51555;
  assign n51557 = ~n51550 & ~n51556;
  assign n51558 = ~controllable_hgrant1 & ~n51557;
  assign n51559 = ~controllable_hgrant1 & ~n51558;
  assign n51560 = ~i_hbusreq3 & ~n51559;
  assign n51561 = ~n51549 & ~n51560;
  assign n51562 = ~controllable_hgrant3 & ~n51561;
  assign n51563 = ~controllable_hgrant3 & ~n51562;
  assign n51564 = ~i_hbusreq9 & ~n51563;
  assign n51565 = ~n51548 & ~n51564;
  assign n51566 = ~i_hbusreq4 & ~n51565;
  assign n51567 = ~n51547 & ~n51566;
  assign n51568 = ~controllable_hgrant4 & ~n51567;
  assign n51569 = ~controllable_hgrant4 & ~n51568;
  assign n51570 = ~i_hbusreq5 & ~n51569;
  assign n51571 = ~n51546 & ~n51570;
  assign n51572 = ~controllable_hgrant5 & ~n51571;
  assign n51573 = ~controllable_hgrant5 & ~n51572;
  assign n51574 = ~controllable_hmaster2 & ~n51573;
  assign n51575 = ~n51545 & ~n51574;
  assign n51576 = ~controllable_hmaster1 & ~n51575;
  assign n51577 = ~n51544 & ~n51576;
  assign n51578 = ~i_hbusreq6 & ~n51577;
  assign n51579 = ~n51503 & ~n51578;
  assign n51580 = ~controllable_hgrant6 & ~n51579;
  assign n51581 = ~n7844 & ~n51580;
  assign n51582 = ~i_hbusreq8 & ~n51581;
  assign n51583 = ~n51502 & ~n51582;
  assign n51584 = controllable_hmaster3 & ~n51583;
  assign n51585 = i_hbusreq8 & ~n51498;
  assign n51586 = i_hbusreq6 & ~n51467;
  assign n51587 = ~i_hbusreq6 & ~n51573;
  assign n51588 = ~n51586 & ~n51587;
  assign n51589 = ~controllable_hgrant6 & ~n51588;
  assign n51590 = ~controllable_hgrant6 & ~n51589;
  assign n51591 = controllable_hmaster0 & ~n51590;
  assign n51592 = i_hbusreq6 & ~n51494;
  assign n51593 = controllable_hmaster2 & ~n51573;
  assign n51594 = i_hbusreq5 & ~n51487;
  assign n51595 = i_hbusreq4 & ~n51485;
  assign n51596 = i_hbusreq9 & ~n51485;
  assign n51597 = i_hbusreq3 & ~n51483;
  assign n51598 = i_hbusreq1 & ~n51481;
  assign n51599 = ~n40876 & ~n44750;
  assign n51600 = ~n7733 & ~n51599;
  assign n51601 = ~n50764 & ~n51600;
  assign n51602 = n7928 & ~n51601;
  assign n51603 = ~n43545 & ~n51602;
  assign n51604 = ~i_hbusreq1 & ~n51603;
  assign n51605 = ~n51598 & ~n51604;
  assign n51606 = ~controllable_hgrant1 & ~n51605;
  assign n51607 = ~n48564 & ~n51606;
  assign n51608 = ~i_hbusreq3 & ~n51607;
  assign n51609 = ~n51597 & ~n51608;
  assign n51610 = ~controllable_hgrant3 & ~n51609;
  assign n51611 = ~n48556 & ~n51610;
  assign n51612 = ~i_hbusreq9 & ~n51611;
  assign n51613 = ~n51596 & ~n51612;
  assign n51614 = ~i_hbusreq4 & ~n51613;
  assign n51615 = ~n51595 & ~n51614;
  assign n51616 = ~controllable_hgrant4 & ~n51615;
  assign n51617 = ~n48547 & ~n51616;
  assign n51618 = ~i_hbusreq5 & ~n51617;
  assign n51619 = ~n51594 & ~n51618;
  assign n51620 = ~controllable_hgrant5 & ~n51619;
  assign n51621 = ~n48536 & ~n51620;
  assign n51622 = ~controllable_hmaster2 & ~n51621;
  assign n51623 = ~n51593 & ~n51622;
  assign n51624 = controllable_hmaster1 & ~n51623;
  assign n51625 = ~controllable_hmaster1 & ~n51573;
  assign n51626 = ~n51624 & ~n51625;
  assign n51627 = ~i_hbusreq6 & ~n51626;
  assign n51628 = ~n51592 & ~n51627;
  assign n51629 = ~controllable_hgrant6 & ~n51628;
  assign n51630 = ~n50616 & ~n51629;
  assign n51631 = ~controllable_hmaster0 & ~n51630;
  assign n51632 = ~n51591 & ~n51631;
  assign n51633 = ~i_hbusreq8 & ~n51632;
  assign n51634 = ~n51585 & ~n51633;
  assign n51635 = ~controllable_hmaster3 & ~n51634;
  assign n51636 = ~n51584 & ~n51635;
  assign n51637 = ~i_hbusreq7 & ~n51636;
  assign n51638 = ~n51501 & ~n51637;
  assign n51639 = n7924 & ~n51638;
  assign n51640 = ~n51441 & ~n51639;
  assign n51641 = n8214 & ~n51640;
  assign n51642 = ~n51359 & ~n51641;
  assign n51643 = n8202 & ~n51642;
  assign n51644 = ~n51143 & ~n51643;
  assign n51645 = n7920 & ~n51644;
  assign n51646 = ~n50812 & ~n51645;
  assign n51647 = ~n7728 & ~n51646;
  assign n51648 = ~n50811 & ~n51647;
  assign n51649 = ~n7723 & ~n51648;
  assign n51650 = ~n7723 & ~n51649;
  assign n51651 = ~n7714 & ~n51650;
  assign n51652 = ~n7714 & ~n51651;
  assign n51653 = n7705 & ~n51652;
  assign n51654 = ~n41300 & ~n48008;
  assign n51655 = controllable_hmaster1 & ~n51654;
  assign n51656 = controllable_hmaster2 & ~n51654;
  assign n51657 = n8378 & ~n8987;
  assign n51658 = ~n8378 & ~n17337;
  assign n51659 = ~n51657 & ~n51658;
  assign n51660 = controllable_hgrant5 & ~n51659;
  assign n51661 = ~n41329 & ~n51660;
  assign n51662 = ~controllable_hmaster2 & ~n51661;
  assign n51663 = ~n51656 & ~n51662;
  assign n51664 = ~controllable_hmaster1 & ~n51663;
  assign n51665 = ~n51655 & ~n51664;
  assign n51666 = ~controllable_hgrant6 & ~n51665;
  assign n51667 = ~n13175 & ~n51666;
  assign n51668 = controllable_hmaster3 & ~n51667;
  assign n51669 = n8217 & ~n10056;
  assign n51670 = ~n8217 & ~n22402;
  assign n51671 = ~n51669 & ~n51670;
  assign n51672 = controllable_hgrant6 & ~n51671;
  assign n51673 = controllable_hmaster2 & ~n51661;
  assign n51674 = ~n41323 & ~n51660;
  assign n51675 = ~controllable_hmaster2 & ~n51674;
  assign n51676 = ~n51673 & ~n51675;
  assign n51677 = controllable_hmaster1 & ~n51676;
  assign n51678 = ~n41339 & ~n51660;
  assign n51679 = ~controllable_hmaster2 & ~n51678;
  assign n51680 = ~n48097 & ~n51679;
  assign n51681 = ~controllable_hmaster1 & ~n51680;
  assign n51682 = ~n51677 & ~n51681;
  assign n51683 = ~controllable_hgrant6 & ~n51682;
  assign n51684 = ~n51672 & ~n51683;
  assign n51685 = controllable_hmaster0 & ~n51684;
  assign n51686 = ~n41360 & ~n51660;
  assign n51687 = ~controllable_hmaster2 & ~n51686;
  assign n51688 = ~n51673 & ~n51687;
  assign n51689 = controllable_hmaster1 & ~n51688;
  assign n51690 = ~n41368 & ~n51660;
  assign n51691 = controllable_hmaster2 & ~n51690;
  assign n51692 = ~n51662 & ~n51691;
  assign n51693 = ~controllable_hmaster1 & ~n51692;
  assign n51694 = ~n51689 & ~n51693;
  assign n51695 = ~controllable_hgrant6 & ~n51694;
  assign n51696 = ~n41348 & ~n51695;
  assign n51697 = ~controllable_hmaster0 & ~n51696;
  assign n51698 = ~n51685 & ~n51697;
  assign n51699 = ~controllable_hmaster3 & ~n51698;
  assign n51700 = ~n51668 & ~n51699;
  assign n51701 = i_hbusreq7 & ~n51700;
  assign n51702 = i_hbusreq8 & ~n51667;
  assign n51703 = i_hbusreq6 & ~n51665;
  assign n51704 = n8378 & ~n8480;
  assign n51705 = ~n8378 & ~n17386;
  assign n51706 = ~n51704 & ~n51705;
  assign n51707 = ~i_hbusreq5 & ~n51706;
  assign n51708 = ~n48244 & ~n51707;
  assign n51709 = controllable_hgrant5 & ~n51708;
  assign n51710 = ~n41417 & ~n51709;
  assign n51711 = controllable_hmaster1 & ~n51710;
  assign n51712 = controllable_hmaster2 & ~n51710;
  assign n51713 = i_hbusreq5 & ~n51659;
  assign n51714 = n8378 & ~n9021;
  assign n51715 = ~n8378 & ~n17430;
  assign n51716 = ~n51714 & ~n51715;
  assign n51717 = ~i_hbusreq5 & ~n51716;
  assign n51718 = ~n51713 & ~n51717;
  assign n51719 = controllable_hgrant5 & ~n51718;
  assign n51720 = ~n41464 & ~n51719;
  assign n51721 = ~controllable_hmaster2 & ~n51720;
  assign n51722 = ~n51712 & ~n51721;
  assign n51723 = ~controllable_hmaster1 & ~n51722;
  assign n51724 = ~n51711 & ~n51723;
  assign n51725 = ~i_hbusreq6 & ~n51724;
  assign n51726 = ~n51703 & ~n51725;
  assign n51727 = ~controllable_hgrant6 & ~n51726;
  assign n51728 = ~n13254 & ~n51727;
  assign n51729 = ~i_hbusreq8 & ~n51728;
  assign n51730 = ~n51702 & ~n51729;
  assign n51731 = controllable_hmaster3 & ~n51730;
  assign n51732 = i_hbusreq8 & ~n51698;
  assign n51733 = i_hbusreq6 & ~n51671;
  assign n51734 = n8217 & ~n10067;
  assign n51735 = ~n8217 & ~n22414;
  assign n51736 = ~n51734 & ~n51735;
  assign n51737 = ~i_hbusreq6 & ~n51736;
  assign n51738 = ~n51733 & ~n51737;
  assign n51739 = controllable_hgrant6 & ~n51738;
  assign n51740 = i_hbusreq6 & ~n51682;
  assign n51741 = controllable_hmaster2 & ~n51720;
  assign n51742 = ~n41458 & ~n51719;
  assign n51743 = ~controllable_hmaster2 & ~n51742;
  assign n51744 = ~n51741 & ~n51743;
  assign n51745 = controllable_hmaster1 & ~n51744;
  assign n51746 = ~n41486 & ~n51719;
  assign n51747 = ~controllable_hmaster2 & ~n51746;
  assign n51748 = ~n48432 & ~n51747;
  assign n51749 = ~controllable_hmaster1 & ~n51748;
  assign n51750 = ~n51745 & ~n51749;
  assign n51751 = ~i_hbusreq6 & ~n51750;
  assign n51752 = ~n51740 & ~n51751;
  assign n51753 = ~controllable_hgrant6 & ~n51752;
  assign n51754 = ~n51739 & ~n51753;
  assign n51755 = controllable_hmaster0 & ~n51754;
  assign n51756 = i_hbusreq6 & ~n51694;
  assign n51757 = ~n41525 & ~n51719;
  assign n51758 = ~controllable_hmaster2 & ~n51757;
  assign n51759 = ~n51741 & ~n51758;
  assign n51760 = controllable_hmaster1 & ~n51759;
  assign n51761 = ~n41536 & ~n51719;
  assign n51762 = controllable_hmaster2 & ~n51761;
  assign n51763 = ~n51721 & ~n51762;
  assign n51764 = ~controllable_hmaster1 & ~n51763;
  assign n51765 = ~n51760 & ~n51764;
  assign n51766 = ~i_hbusreq6 & ~n51765;
  assign n51767 = ~n51756 & ~n51766;
  assign n51768 = ~controllable_hgrant6 & ~n51767;
  assign n51769 = ~n41497 & ~n51768;
  assign n51770 = ~controllable_hmaster0 & ~n51769;
  assign n51771 = ~n51755 & ~n51770;
  assign n51772 = ~i_hbusreq8 & ~n51771;
  assign n51773 = ~n51732 & ~n51772;
  assign n51774 = ~controllable_hmaster3 & ~n51773;
  assign n51775 = ~n51731 & ~n51774;
  assign n51776 = ~i_hbusreq7 & ~n51775;
  assign n51777 = ~n51701 & ~n51776;
  assign n51778 = ~n7924 & ~n51777;
  assign n51779 = ~n41576 & ~n48769;
  assign n51780 = controllable_hmaster1 & ~n51779;
  assign n51781 = controllable_hmaster2 & ~n51779;
  assign n51782 = n8378 & ~n13186;
  assign n51783 = ~n8378 & ~n29494;
  assign n51784 = ~n51782 & ~n51783;
  assign n51785 = i_hlock5 & ~n51784;
  assign n51786 = ~n8378 & ~n29525;
  assign n51787 = ~n51782 & ~n51786;
  assign n51788 = ~i_hlock5 & ~n51787;
  assign n51789 = ~n51785 & ~n51788;
  assign n51790 = controllable_hgrant5 & ~n51789;
  assign n51791 = ~n41664 & ~n51790;
  assign n51792 = ~controllable_hmaster2 & ~n51791;
  assign n51793 = ~n51781 & ~n51792;
  assign n51794 = ~controllable_hmaster1 & ~n51793;
  assign n51795 = ~n51780 & ~n51794;
  assign n51796 = ~controllable_hgrant6 & ~n51795;
  assign n51797 = ~n41646 & ~n51796;
  assign n51798 = controllable_hmaster3 & ~n51797;
  assign n51799 = n8217 & ~n15197;
  assign n51800 = ~n8217 & ~n22436;
  assign n51801 = ~n51799 & ~n51800;
  assign n51802 = controllable_hgrant6 & ~n51801;
  assign n51803 = controllable_hmaster2 & ~n51791;
  assign n51804 = ~n41681 & ~n51790;
  assign n51805 = ~controllable_hmaster2 & ~n51804;
  assign n51806 = ~n51803 & ~n51805;
  assign n51807 = controllable_hmaster1 & ~n51806;
  assign n51808 = i_hlock5 & ~n42163;
  assign n51809 = ~i_hlock5 & ~n42185;
  assign n51810 = ~n51808 & ~n51809;
  assign n51811 = ~controllable_hgrant5 & ~n51810;
  assign n51812 = ~n48879 & ~n51811;
  assign n51813 = controllable_hmaster2 & ~n51812;
  assign n51814 = ~n41695 & ~n51790;
  assign n51815 = ~controllable_hmaster2 & ~n51814;
  assign n51816 = ~n51813 & ~n51815;
  assign n51817 = ~controllable_hmaster1 & ~n51816;
  assign n51818 = ~n51807 & ~n51817;
  assign n51819 = ~controllable_hgrant6 & ~n51818;
  assign n51820 = ~n51802 & ~n51819;
  assign n51821 = controllable_hmaster0 & ~n51820;
  assign n51822 = ~n41719 & ~n51790;
  assign n51823 = ~controllable_hmaster2 & ~n51822;
  assign n51824 = ~n51803 & ~n51823;
  assign n51825 = controllable_hmaster1 & ~n51824;
  assign n51826 = ~n41726 & ~n51790;
  assign n51827 = controllable_hmaster2 & ~n51826;
  assign n51828 = ~n51792 & ~n51827;
  assign n51829 = ~controllable_hmaster1 & ~n51828;
  assign n51830 = ~n51825 & ~n51829;
  assign n51831 = ~controllable_hgrant6 & ~n51830;
  assign n51832 = ~n41704 & ~n51831;
  assign n51833 = ~controllable_hmaster0 & ~n51832;
  assign n51834 = ~n51821 & ~n51833;
  assign n51835 = ~controllable_hmaster3 & ~n51834;
  assign n51836 = ~n51798 & ~n51835;
  assign n51837 = i_hbusreq7 & ~n51836;
  assign n51838 = i_hbusreq8 & ~n51797;
  assign n51839 = i_hbusreq6 & ~n51795;
  assign n51840 = n8378 & ~n13239;
  assign n51841 = ~n8378 & ~n29561;
  assign n51842 = ~n51840 & ~n51841;
  assign n51843 = i_hlock5 & ~n51842;
  assign n51844 = ~n8378 & ~n29625;
  assign n51845 = ~n51840 & ~n51844;
  assign n51846 = ~i_hlock5 & ~n51845;
  assign n51847 = ~n51843 & ~n51846;
  assign n51848 = ~i_hbusreq5 & ~n51847;
  assign n51849 = ~n49101 & ~n51848;
  assign n51850 = controllable_hgrant5 & ~n51849;
  assign n51851 = ~n41781 & ~n51850;
  assign n51852 = controllable_hmaster1 & ~n51851;
  assign n51853 = controllable_hmaster2 & ~n51851;
  assign n51854 = i_hbusreq5 & ~n51789;
  assign n51855 = n8378 & ~n13279;
  assign n51856 = ~n8378 & ~n29576;
  assign n51857 = ~n51855 & ~n51856;
  assign n51858 = i_hlock5 & ~n51857;
  assign n51859 = ~n8378 & ~n29640;
  assign n51860 = ~n51855 & ~n51859;
  assign n51861 = ~i_hlock5 & ~n51860;
  assign n51862 = ~n51858 & ~n51861;
  assign n51863 = ~i_hbusreq5 & ~n51862;
  assign n51864 = ~n51854 & ~n51863;
  assign n51865 = controllable_hgrant5 & ~n51864;
  assign n51866 = ~n41946 & ~n51865;
  assign n51867 = ~controllable_hmaster2 & ~n51866;
  assign n51868 = ~n51853 & ~n51867;
  assign n51869 = ~controllable_hmaster1 & ~n51868;
  assign n51870 = ~n51852 & ~n51869;
  assign n51871 = ~i_hbusreq6 & ~n51870;
  assign n51872 = ~n51839 & ~n51871;
  assign n51873 = ~controllable_hgrant6 & ~n51872;
  assign n51874 = ~n41907 & ~n51873;
  assign n51875 = ~i_hbusreq8 & ~n51874;
  assign n51876 = ~n51838 & ~n51875;
  assign n51877 = controllable_hmaster3 & ~n51876;
  assign n51878 = i_hbusreq8 & ~n51834;
  assign n51879 = i_hbusreq6 & ~n51801;
  assign n51880 = n8217 & ~n15219;
  assign n51881 = ~n8217 & ~n22457;
  assign n51882 = ~n51880 & ~n51881;
  assign n51883 = ~i_hbusreq6 & ~n51882;
  assign n51884 = ~n51879 & ~n51883;
  assign n51885 = controllable_hgrant6 & ~n51884;
  assign n51886 = i_hbusreq6 & ~n51818;
  assign n51887 = controllable_hmaster2 & ~n51866;
  assign n51888 = ~n41978 & ~n51865;
  assign n51889 = ~controllable_hmaster2 & ~n51888;
  assign n51890 = ~n51887 & ~n51889;
  assign n51891 = controllable_hmaster1 & ~n51890;
  assign n51892 = i_hbusreq5 & ~n51810;
  assign n51893 = i_hlock5 & ~n42233;
  assign n51894 = ~i_hlock5 & ~n42279;
  assign n51895 = ~n51893 & ~n51894;
  assign n51896 = ~i_hbusreq5 & ~n51895;
  assign n51897 = ~n51892 & ~n51896;
  assign n51898 = ~controllable_hgrant5 & ~n51897;
  assign n51899 = ~n49568 & ~n51898;
  assign n51900 = controllable_hmaster2 & ~n51899;
  assign n51901 = ~n42004 & ~n51865;
  assign n51902 = ~controllable_hmaster2 & ~n51901;
  assign n51903 = ~n51900 & ~n51902;
  assign n51904 = ~controllable_hmaster1 & ~n51903;
  assign n51905 = ~n51891 & ~n51904;
  assign n51906 = ~i_hbusreq6 & ~n51905;
  assign n51907 = ~n51886 & ~n51906;
  assign n51908 = ~controllable_hgrant6 & ~n51907;
  assign n51909 = ~n51885 & ~n51908;
  assign n51910 = controllable_hmaster0 & ~n51909;
  assign n51911 = i_hbusreq6 & ~n51830;
  assign n51912 = ~n42046 & ~n51865;
  assign n51913 = ~controllable_hmaster2 & ~n51912;
  assign n51914 = ~n51887 & ~n51913;
  assign n51915 = controllable_hmaster1 & ~n51914;
  assign n51916 = ~n42056 & ~n51865;
  assign n51917 = controllable_hmaster2 & ~n51916;
  assign n51918 = ~n51867 & ~n51917;
  assign n51919 = ~controllable_hmaster1 & ~n51918;
  assign n51920 = ~n51915 & ~n51919;
  assign n51921 = ~i_hbusreq6 & ~n51920;
  assign n51922 = ~n51911 & ~n51921;
  assign n51923 = ~controllable_hgrant6 & ~n51922;
  assign n51924 = ~n42015 & ~n51923;
  assign n51925 = ~controllable_hmaster0 & ~n51924;
  assign n51926 = ~n51910 & ~n51925;
  assign n51927 = ~i_hbusreq8 & ~n51926;
  assign n51928 = ~n51878 & ~n51927;
  assign n51929 = ~controllable_hmaster3 & ~n51928;
  assign n51930 = ~n51877 & ~n51929;
  assign n51931 = ~i_hbusreq7 & ~n51930;
  assign n51932 = ~n51837 & ~n51931;
  assign n51933 = n7924 & ~n51932;
  assign n51934 = ~n51778 & ~n51933;
  assign n51935 = ~n8214 & ~n51934;
  assign n51936 = ~n41298 & ~n48011;
  assign n51937 = ~controllable_hgrant5 & ~n51936;
  assign n51938 = ~n13152 & ~n51937;
  assign n51939 = controllable_hmaster1 & ~n51938;
  assign n51940 = controllable_hmaster2 & ~n51938;
  assign n51941 = n8426 & ~n8987;
  assign n51942 = ~n8426 & ~n17335;
  assign n51943 = ~n51941 & ~n51942;
  assign n51944 = controllable_hgrant4 & ~n51943;
  assign n51945 = ~n41366 & ~n51944;
  assign n51946 = ~controllable_hgrant5 & ~n51945;
  assign n51947 = ~n13176 & ~n51946;
  assign n51948 = ~controllable_hmaster2 & ~n51947;
  assign n51949 = ~n51940 & ~n51948;
  assign n51950 = ~controllable_hmaster1 & ~n51949;
  assign n51951 = ~n51939 & ~n51950;
  assign n51952 = ~controllable_hgrant6 & ~n51951;
  assign n51953 = ~n13175 & ~n51952;
  assign n51954 = controllable_hmaster3 & ~n51953;
  assign n51955 = controllable_hmaster2 & ~n51947;
  assign n51956 = ~n41321 & ~n51944;
  assign n51957 = ~controllable_hgrant5 & ~n51956;
  assign n51958 = ~n13176 & ~n51957;
  assign n51959 = ~controllable_hmaster2 & ~n51958;
  assign n51960 = ~n51955 & ~n51959;
  assign n51961 = controllable_hmaster1 & ~n51960;
  assign n51962 = ~n41328 & ~n51946;
  assign n51963 = controllable_hmaster2 & ~n51962;
  assign n51964 = ~n41337 & ~n51944;
  assign n51965 = ~controllable_hgrant5 & ~n51964;
  assign n51966 = ~n13176 & ~n51965;
  assign n51967 = ~controllable_hmaster2 & ~n51966;
  assign n51968 = ~n51963 & ~n51967;
  assign n51969 = ~controllable_hmaster1 & ~n51968;
  assign n51970 = ~n51961 & ~n51969;
  assign n51971 = ~controllable_hgrant6 & ~n51970;
  assign n51972 = ~n13198 & ~n51971;
  assign n51973 = controllable_hmaster0 & ~n51972;
  assign n51974 = ~n10080 & ~n26890;
  assign n51975 = n8217 & ~n51974;
  assign n51976 = ~n22474 & ~n26890;
  assign n51977 = ~n8217 & ~n51976;
  assign n51978 = ~n51975 & ~n51977;
  assign n51979 = controllable_hgrant6 & ~n51978;
  assign n51980 = ~n41358 & ~n51944;
  assign n51981 = ~controllable_hgrant5 & ~n51980;
  assign n51982 = ~n13176 & ~n51981;
  assign n51983 = ~controllable_hmaster2 & ~n51982;
  assign n51984 = ~n51955 & ~n51983;
  assign n51985 = controllable_hmaster1 & ~n51984;
  assign n51986 = ~n48185 & ~n51948;
  assign n51987 = ~controllable_hmaster1 & ~n51986;
  assign n51988 = ~n51985 & ~n51987;
  assign n51989 = ~controllable_hgrant6 & ~n51988;
  assign n51990 = ~n51979 & ~n51989;
  assign n51991 = ~controllable_hmaster0 & ~n51990;
  assign n51992 = ~n51973 & ~n51991;
  assign n51993 = ~controllable_hmaster3 & ~n51992;
  assign n51994 = ~n51954 & ~n51993;
  assign n51995 = i_hbusreq7 & ~n51994;
  assign n51996 = i_hbusreq8 & ~n51953;
  assign n51997 = i_hbusreq6 & ~n51951;
  assign n51998 = i_hbusreq5 & ~n51936;
  assign n51999 = n8426 & ~n8476;
  assign n52000 = ~n8426 & ~n17380;
  assign n52001 = ~n51999 & ~n52000;
  assign n52002 = ~i_hbusreq9 & ~n52001;
  assign n52003 = ~n48253 & ~n52002;
  assign n52004 = ~i_hbusreq4 & ~n52003;
  assign n52005 = ~n48252 & ~n52004;
  assign n52006 = controllable_hgrant4 & ~n52005;
  assign n52007 = ~n41413 & ~n52006;
  assign n52008 = ~i_hbusreq5 & ~n52007;
  assign n52009 = ~n51998 & ~n52008;
  assign n52010 = ~controllable_hgrant5 & ~n52009;
  assign n52011 = ~n13206 & ~n52010;
  assign n52012 = controllable_hmaster1 & ~n52011;
  assign n52013 = controllable_hmaster2 & ~n52011;
  assign n52014 = i_hbusreq5 & ~n51945;
  assign n52015 = i_hbusreq4 & ~n51943;
  assign n52016 = i_hbusreq9 & ~n51943;
  assign n52017 = n8426 & ~n9017;
  assign n52018 = ~n8426 & ~n17424;
  assign n52019 = ~n52017 & ~n52018;
  assign n52020 = ~i_hbusreq9 & ~n52019;
  assign n52021 = ~n52016 & ~n52020;
  assign n52022 = ~i_hbusreq4 & ~n52021;
  assign n52023 = ~n52015 & ~n52022;
  assign n52024 = controllable_hgrant4 & ~n52023;
  assign n52025 = ~n41532 & ~n52024;
  assign n52026 = ~i_hbusreq5 & ~n52025;
  assign n52027 = ~n52014 & ~n52026;
  assign n52028 = ~controllable_hgrant5 & ~n52027;
  assign n52029 = ~n13256 & ~n52028;
  assign n52030 = ~controllable_hmaster2 & ~n52029;
  assign n52031 = ~n52013 & ~n52030;
  assign n52032 = ~controllable_hmaster1 & ~n52031;
  assign n52033 = ~n52012 & ~n52032;
  assign n52034 = ~i_hbusreq6 & ~n52033;
  assign n52035 = ~n51997 & ~n52034;
  assign n52036 = ~controllable_hgrant6 & ~n52035;
  assign n52037 = ~n13254 & ~n52036;
  assign n52038 = ~i_hbusreq8 & ~n52037;
  assign n52039 = ~n51996 & ~n52038;
  assign n52040 = controllable_hmaster3 & ~n52039;
  assign n52041 = i_hbusreq8 & ~n51992;
  assign n52042 = i_hbusreq6 & ~n51970;
  assign n52043 = controllable_hmaster2 & ~n52029;
  assign n52044 = i_hbusreq5 & ~n51956;
  assign n52045 = ~n41454 & ~n52024;
  assign n52046 = ~i_hbusreq5 & ~n52045;
  assign n52047 = ~n52044 & ~n52046;
  assign n52048 = ~controllable_hgrant5 & ~n52047;
  assign n52049 = ~n13256 & ~n52048;
  assign n52050 = ~controllable_hmaster2 & ~n52049;
  assign n52051 = ~n52043 & ~n52050;
  assign n52052 = controllable_hmaster1 & ~n52051;
  assign n52053 = ~n41463 & ~n52028;
  assign n52054 = controllable_hmaster2 & ~n52053;
  assign n52055 = i_hbusreq5 & ~n51964;
  assign n52056 = ~n41482 & ~n52024;
  assign n52057 = ~i_hbusreq5 & ~n52056;
  assign n52058 = ~n52055 & ~n52057;
  assign n52059 = ~controllable_hgrant5 & ~n52058;
  assign n52060 = ~n13256 & ~n52059;
  assign n52061 = ~controllable_hmaster2 & ~n52060;
  assign n52062 = ~n52054 & ~n52061;
  assign n52063 = ~controllable_hmaster1 & ~n52062;
  assign n52064 = ~n52052 & ~n52063;
  assign n52065 = ~i_hbusreq6 & ~n52064;
  assign n52066 = ~n52042 & ~n52065;
  assign n52067 = ~controllable_hgrant6 & ~n52066;
  assign n52068 = ~n13298 & ~n52067;
  assign n52069 = controllable_hmaster0 & ~n52068;
  assign n52070 = i_hbusreq6 & ~n51978;
  assign n52071 = ~n10090 & ~n26903;
  assign n52072 = n8217 & ~n52071;
  assign n52073 = ~n22486 & ~n26903;
  assign n52074 = ~n8217 & ~n52073;
  assign n52075 = ~n52072 & ~n52074;
  assign n52076 = ~i_hbusreq6 & ~n52075;
  assign n52077 = ~n52070 & ~n52076;
  assign n52078 = controllable_hgrant6 & ~n52077;
  assign n52079 = i_hbusreq6 & ~n51988;
  assign n52080 = i_hbusreq5 & ~n51980;
  assign n52081 = ~n41521 & ~n52024;
  assign n52082 = ~i_hbusreq5 & ~n52081;
  assign n52083 = ~n52080 & ~n52082;
  assign n52084 = ~controllable_hgrant5 & ~n52083;
  assign n52085 = ~n13256 & ~n52084;
  assign n52086 = ~controllable_hmaster2 & ~n52085;
  assign n52087 = ~n52043 & ~n52086;
  assign n52088 = controllable_hmaster1 & ~n52087;
  assign n52089 = ~n48648 & ~n52030;
  assign n52090 = ~controllable_hmaster1 & ~n52089;
  assign n52091 = ~n52088 & ~n52090;
  assign n52092 = ~i_hbusreq6 & ~n52091;
  assign n52093 = ~n52079 & ~n52092;
  assign n52094 = ~controllable_hgrant6 & ~n52093;
  assign n52095 = ~n52078 & ~n52094;
  assign n52096 = ~controllable_hmaster0 & ~n52095;
  assign n52097 = ~n52069 & ~n52096;
  assign n52098 = ~i_hbusreq8 & ~n52097;
  assign n52099 = ~n52041 & ~n52098;
  assign n52100 = ~controllable_hmaster3 & ~n52099;
  assign n52101 = ~n52040 & ~n52100;
  assign n52102 = ~i_hbusreq7 & ~n52101;
  assign n52103 = ~n51995 & ~n52102;
  assign n52104 = ~n7924 & ~n52103;
  assign n52105 = ~n41574 & ~n48777;
  assign n52106 = ~controllable_hgrant5 & ~n52105;
  assign n52107 = ~n41559 & ~n52106;
  assign n52108 = controllable_hmaster1 & ~n52107;
  assign n52109 = controllable_hmaster2 & ~n52107;
  assign n52110 = n8426 & ~n13184;
  assign n52111 = ~n8426 & ~n17514;
  assign n52112 = ~n52110 & ~n52111;
  assign n52113 = i_hlock4 & ~n52112;
  assign n52114 = ~n8426 & ~n17522;
  assign n52115 = ~n52110 & ~n52114;
  assign n52116 = ~i_hlock4 & ~n52115;
  assign n52117 = ~n52113 & ~n52116;
  assign n52118 = controllable_hgrant4 & ~n52117;
  assign n52119 = ~n41662 & ~n52118;
  assign n52120 = ~controllable_hgrant5 & ~n52119;
  assign n52121 = ~n41647 & ~n52120;
  assign n52122 = ~controllable_hmaster2 & ~n52121;
  assign n52123 = ~n52109 & ~n52122;
  assign n52124 = ~controllable_hmaster1 & ~n52123;
  assign n52125 = ~n52108 & ~n52124;
  assign n52126 = ~controllable_hgrant6 & ~n52125;
  assign n52127 = ~n41646 & ~n52126;
  assign n52128 = controllable_hmaster3 & ~n52127;
  assign n52129 = controllable_hmaster2 & ~n52121;
  assign n52130 = ~n41679 & ~n52118;
  assign n52131 = ~controllable_hgrant5 & ~n52130;
  assign n52132 = ~n41647 & ~n52131;
  assign n52133 = ~controllable_hmaster2 & ~n52132;
  assign n52134 = ~n52129 & ~n52133;
  assign n52135 = controllable_hmaster1 & ~n52134;
  assign n52136 = ~n41686 & ~n52120;
  assign n52137 = controllable_hmaster2 & ~n52136;
  assign n52138 = ~n41693 & ~n52118;
  assign n52139 = ~controllable_hgrant5 & ~n52138;
  assign n52140 = ~n41647 & ~n52139;
  assign n52141 = ~controllable_hmaster2 & ~n52140;
  assign n52142 = ~n52137 & ~n52141;
  assign n52143 = ~controllable_hmaster1 & ~n52142;
  assign n52144 = ~n52135 & ~n52143;
  assign n52145 = ~controllable_hgrant6 & ~n52144;
  assign n52146 = ~n41675 & ~n52145;
  assign n52147 = controllable_hmaster0 & ~n52146;
  assign n52148 = ~n15243 & ~n26936;
  assign n52149 = n8217 & ~n52148;
  assign n52150 = ~n22510 & ~n26936;
  assign n52151 = ~n8217 & ~n52150;
  assign n52152 = ~n52149 & ~n52151;
  assign n52153 = controllable_hgrant6 & ~n52152;
  assign n52154 = ~n41717 & ~n52118;
  assign n52155 = ~controllable_hgrant5 & ~n52154;
  assign n52156 = ~n41647 & ~n52155;
  assign n52157 = ~controllable_hmaster2 & ~n52156;
  assign n52158 = ~n52129 & ~n52157;
  assign n52159 = controllable_hmaster1 & ~n52158;
  assign n52160 = ~n8378 & ~n22505;
  assign n52161 = ~n44054 & ~n52160;
  assign n52162 = controllable_hgrant5 & ~n52161;
  assign n52163 = i_hlock4 & ~n41618;
  assign n52164 = ~i_hlock4 & ~n41632;
  assign n52165 = ~n52163 & ~n52164;
  assign n52166 = ~controllable_hgrant4 & ~n52165;
  assign n52167 = ~n49009 & ~n52166;
  assign n52168 = ~controllable_hgrant5 & ~n52167;
  assign n52169 = ~n52162 & ~n52168;
  assign n52170 = controllable_hmaster2 & ~n52169;
  assign n52171 = ~n52122 & ~n52170;
  assign n52172 = ~controllable_hmaster1 & ~n52171;
  assign n52173 = ~n52159 & ~n52172;
  assign n52174 = ~controllable_hgrant6 & ~n52173;
  assign n52175 = ~n52153 & ~n52174;
  assign n52176 = ~controllable_hmaster0 & ~n52175;
  assign n52177 = ~n52147 & ~n52176;
  assign n52178 = ~controllable_hmaster3 & ~n52177;
  assign n52179 = ~n52128 & ~n52178;
  assign n52180 = i_hbusreq7 & ~n52179;
  assign n52181 = i_hbusreq8 & ~n52127;
  assign n52182 = i_hbusreq6 & ~n52125;
  assign n52183 = i_hbusreq5 & ~n52105;
  assign n52184 = n8426 & ~n13233;
  assign n52185 = ~n8426 & ~n17575;
  assign n52186 = ~n52184 & ~n52185;
  assign n52187 = ~i_hbusreq9 & ~n52186;
  assign n52188 = ~n49115 & ~n52187;
  assign n52189 = i_hlock4 & ~n52188;
  assign n52190 = ~n8426 & ~n17597;
  assign n52191 = ~n52184 & ~n52190;
  assign n52192 = ~i_hbusreq9 & ~n52191;
  assign n52193 = ~n49122 & ~n52192;
  assign n52194 = ~i_hlock4 & ~n52193;
  assign n52195 = ~n52189 & ~n52194;
  assign n52196 = ~i_hbusreq4 & ~n52195;
  assign n52197 = ~n49114 & ~n52196;
  assign n52198 = controllable_hgrant4 & ~n52197;
  assign n52199 = ~n41777 & ~n52198;
  assign n52200 = ~i_hbusreq5 & ~n52199;
  assign n52201 = ~n52183 & ~n52200;
  assign n52202 = ~controllable_hgrant5 & ~n52201;
  assign n52203 = ~n41748 & ~n52202;
  assign n52204 = controllable_hmaster1 & ~n52203;
  assign n52205 = controllable_hmaster2 & ~n52203;
  assign n52206 = i_hbusreq5 & ~n52119;
  assign n52207 = i_hbusreq4 & ~n52117;
  assign n52208 = i_hbusreq9 & ~n52112;
  assign n52209 = n8426 & ~n13273;
  assign n52210 = ~n8426 & ~n17650;
  assign n52211 = ~n52209 & ~n52210;
  assign n52212 = ~i_hbusreq9 & ~n52211;
  assign n52213 = ~n52208 & ~n52212;
  assign n52214 = i_hlock4 & ~n52213;
  assign n52215 = i_hbusreq9 & ~n52115;
  assign n52216 = ~n8426 & ~n17664;
  assign n52217 = ~n52209 & ~n52216;
  assign n52218 = ~i_hbusreq9 & ~n52217;
  assign n52219 = ~n52215 & ~n52218;
  assign n52220 = ~i_hlock4 & ~n52219;
  assign n52221 = ~n52214 & ~n52220;
  assign n52222 = ~i_hbusreq4 & ~n52221;
  assign n52223 = ~n52207 & ~n52222;
  assign n52224 = controllable_hgrant4 & ~n52223;
  assign n52225 = ~n41942 & ~n52224;
  assign n52226 = ~i_hbusreq5 & ~n52225;
  assign n52227 = ~n52206 & ~n52226;
  assign n52228 = ~controllable_hgrant5 & ~n52227;
  assign n52229 = ~n41909 & ~n52228;
  assign n52230 = ~controllable_hmaster2 & ~n52229;
  assign n52231 = ~n52205 & ~n52230;
  assign n52232 = ~controllable_hmaster1 & ~n52231;
  assign n52233 = ~n52204 & ~n52232;
  assign n52234 = ~i_hbusreq6 & ~n52233;
  assign n52235 = ~n52182 & ~n52234;
  assign n52236 = ~controllable_hgrant6 & ~n52235;
  assign n52237 = ~n41907 & ~n52236;
  assign n52238 = ~i_hbusreq8 & ~n52237;
  assign n52239 = ~n52181 & ~n52238;
  assign n52240 = controllable_hmaster3 & ~n52239;
  assign n52241 = i_hbusreq8 & ~n52177;
  assign n52242 = i_hbusreq6 & ~n52144;
  assign n52243 = controllable_hmaster2 & ~n52229;
  assign n52244 = i_hbusreq5 & ~n52130;
  assign n52245 = ~n41974 & ~n52224;
  assign n52246 = ~i_hbusreq5 & ~n52245;
  assign n52247 = ~n52244 & ~n52246;
  assign n52248 = ~controllable_hgrant5 & ~n52247;
  assign n52249 = ~n41909 & ~n52248;
  assign n52250 = ~controllable_hmaster2 & ~n52249;
  assign n52251 = ~n52243 & ~n52250;
  assign n52252 = controllable_hmaster1 & ~n52251;
  assign n52253 = ~n41983 & ~n52228;
  assign n52254 = controllable_hmaster2 & ~n52253;
  assign n52255 = i_hbusreq5 & ~n52138;
  assign n52256 = ~n42000 & ~n52224;
  assign n52257 = ~i_hbusreq5 & ~n52256;
  assign n52258 = ~n52255 & ~n52257;
  assign n52259 = ~controllable_hgrant5 & ~n52258;
  assign n52260 = ~n41909 & ~n52259;
  assign n52261 = ~controllable_hmaster2 & ~n52260;
  assign n52262 = ~n52254 & ~n52261;
  assign n52263 = ~controllable_hmaster1 & ~n52262;
  assign n52264 = ~n52252 & ~n52263;
  assign n52265 = ~i_hbusreq6 & ~n52264;
  assign n52266 = ~n52242 & ~n52265;
  assign n52267 = ~controllable_hgrant6 & ~n52266;
  assign n52268 = ~n41962 & ~n52267;
  assign n52269 = controllable_hmaster0 & ~n52268;
  assign n52270 = i_hbusreq6 & ~n52152;
  assign n52271 = ~n15268 & ~n26980;
  assign n52272 = n8217 & ~n52271;
  assign n52273 = ~n22536 & ~n26980;
  assign n52274 = ~n8217 & ~n52273;
  assign n52275 = ~n52272 & ~n52274;
  assign n52276 = ~i_hbusreq6 & ~n52275;
  assign n52277 = ~n52270 & ~n52276;
  assign n52278 = controllable_hgrant6 & ~n52277;
  assign n52279 = i_hbusreq6 & ~n52173;
  assign n52280 = i_hbusreq5 & ~n52154;
  assign n52281 = ~n42042 & ~n52224;
  assign n52282 = ~i_hbusreq5 & ~n52281;
  assign n52283 = ~n52280 & ~n52282;
  assign n52284 = ~controllable_hgrant5 & ~n52283;
  assign n52285 = ~n41909 & ~n52284;
  assign n52286 = ~controllable_hmaster2 & ~n52285;
  assign n52287 = ~n52243 & ~n52286;
  assign n52288 = controllable_hmaster1 & ~n52287;
  assign n52289 = i_hbusreq5 & ~n52161;
  assign n52290 = n8378 & ~n15261;
  assign n52291 = ~n8378 & ~n22529;
  assign n52292 = ~n52290 & ~n52291;
  assign n52293 = ~i_hbusreq5 & ~n52292;
  assign n52294 = ~n52289 & ~n52293;
  assign n52295 = controllable_hgrant5 & ~n52294;
  assign n52296 = i_hbusreq5 & ~n52167;
  assign n52297 = i_hbusreq4 & ~n52165;
  assign n52298 = i_hlock4 & ~n42229;
  assign n52299 = ~i_hlock4 & ~n42275;
  assign n52300 = ~n52298 & ~n52299;
  assign n52301 = ~i_hbusreq4 & ~n52300;
  assign n52302 = ~n52297 & ~n52301;
  assign n52303 = ~controllable_hgrant4 & ~n52302;
  assign n52304 = ~n49828 & ~n52303;
  assign n52305 = ~i_hbusreq5 & ~n52304;
  assign n52306 = ~n52296 & ~n52305;
  assign n52307 = ~controllable_hgrant5 & ~n52306;
  assign n52308 = ~n52295 & ~n52307;
  assign n52309 = controllable_hmaster2 & ~n52308;
  assign n52310 = ~n52230 & ~n52309;
  assign n52311 = ~controllable_hmaster1 & ~n52310;
  assign n52312 = ~n52288 & ~n52311;
  assign n52313 = ~i_hbusreq6 & ~n52312;
  assign n52314 = ~n52279 & ~n52313;
  assign n52315 = ~controllable_hgrant6 & ~n52314;
  assign n52316 = ~n52278 & ~n52315;
  assign n52317 = ~controllable_hmaster0 & ~n52316;
  assign n52318 = ~n52269 & ~n52317;
  assign n52319 = ~i_hbusreq8 & ~n52318;
  assign n52320 = ~n52241 & ~n52319;
  assign n52321 = ~controllable_hmaster3 & ~n52320;
  assign n52322 = ~n52240 & ~n52321;
  assign n52323 = ~i_hbusreq7 & ~n52322;
  assign n52324 = ~n52180 & ~n52323;
  assign n52325 = n7924 & ~n52324;
  assign n52326 = ~n52104 & ~n52325;
  assign n52327 = n8214 & ~n52326;
  assign n52328 = ~n51935 & ~n52327;
  assign n52329 = ~n8202 & ~n52328;
  assign n52330 = ~n41296 & ~n48014;
  assign n52331 = ~controllable_hgrant4 & ~n52330;
  assign n52332 = ~n13153 & ~n52331;
  assign n52333 = ~controllable_hgrant5 & ~n52332;
  assign n52334 = ~n13152 & ~n52333;
  assign n52335 = controllable_hmaster1 & ~n52334;
  assign n52336 = controllable_hmaster2 & ~n52334;
  assign n52337 = n8365 & ~n8987;
  assign n52338 = ~n8365 & ~n17333;
  assign n52339 = ~n52337 & ~n52338;
  assign n52340 = controllable_hgrant3 & ~n52339;
  assign n52341 = ~n41319 & ~n52340;
  assign n52342 = ~controllable_hgrant4 & ~n52341;
  assign n52343 = ~n13177 & ~n52342;
  assign n52344 = ~controllable_hgrant5 & ~n52343;
  assign n52345 = ~n13176 & ~n52344;
  assign n52346 = ~controllable_hmaster2 & ~n52345;
  assign n52347 = ~n52336 & ~n52346;
  assign n52348 = ~controllable_hmaster1 & ~n52347;
  assign n52349 = ~n52335 & ~n52348;
  assign n52350 = ~controllable_hgrant6 & ~n52349;
  assign n52351 = ~n13175 & ~n52350;
  assign n52352 = controllable_hmaster3 & ~n52351;
  assign n52353 = n8217 & ~n10108;
  assign n52354 = ~n8217 & ~n22557;
  assign n52355 = ~n52353 & ~n52354;
  assign n52356 = controllable_hgrant6 & ~n52355;
  assign n52357 = controllable_hmaster2 & ~n52345;
  assign n52358 = ~n48081 & ~n52357;
  assign n52359 = controllable_hmaster1 & ~n52358;
  assign n52360 = ~n41328 & ~n52344;
  assign n52361 = controllable_hmaster2 & ~n52360;
  assign n52362 = ~n41335 & ~n52340;
  assign n52363 = ~controllable_hgrant4 & ~n52362;
  assign n52364 = ~n13177 & ~n52363;
  assign n52365 = ~controllable_hgrant5 & ~n52364;
  assign n52366 = ~n13176 & ~n52365;
  assign n52367 = ~controllable_hmaster2 & ~n52366;
  assign n52368 = ~n52361 & ~n52367;
  assign n52369 = ~controllable_hmaster1 & ~n52368;
  assign n52370 = ~n52359 & ~n52369;
  assign n52371 = ~controllable_hgrant6 & ~n52370;
  assign n52372 = ~n52356 & ~n52371;
  assign n52373 = controllable_hmaster0 & ~n52372;
  assign n52374 = ~n41356 & ~n52340;
  assign n52375 = ~controllable_hgrant4 & ~n52374;
  assign n52376 = ~n13177 & ~n52375;
  assign n52377 = ~controllable_hgrant5 & ~n52376;
  assign n52378 = ~n13176 & ~n52377;
  assign n52379 = ~controllable_hmaster2 & ~n52378;
  assign n52380 = ~n52357 & ~n52379;
  assign n52381 = controllable_hmaster1 & ~n52380;
  assign n52382 = ~n41365 & ~n52342;
  assign n52383 = ~controllable_hgrant5 & ~n52382;
  assign n52384 = ~n13176 & ~n52383;
  assign n52385 = controllable_hmaster2 & ~n52384;
  assign n52386 = ~n52346 & ~n52385;
  assign n52387 = ~controllable_hmaster1 & ~n52386;
  assign n52388 = ~n52381 & ~n52387;
  assign n52389 = ~controllable_hgrant6 & ~n52388;
  assign n52390 = ~n41348 & ~n52389;
  assign n52391 = ~controllable_hmaster0 & ~n52390;
  assign n52392 = ~n52373 & ~n52391;
  assign n52393 = ~controllable_hmaster3 & ~n52392;
  assign n52394 = ~n52352 & ~n52393;
  assign n52395 = i_hbusreq7 & ~n52394;
  assign n52396 = i_hbusreq8 & ~n52351;
  assign n52397 = i_hbusreq6 & ~n52349;
  assign n52398 = i_hbusreq5 & ~n52332;
  assign n52399 = i_hbusreq4 & ~n52330;
  assign n52400 = i_hbusreq9 & ~n52330;
  assign n52401 = n8365 & ~n8474;
  assign n52402 = ~n8365 & ~n17376;
  assign n52403 = ~n52401 & ~n52402;
  assign n52404 = ~i_hbusreq3 & ~n52403;
  assign n52405 = ~n48264 & ~n52404;
  assign n52406 = controllable_hgrant3 & ~n52405;
  assign n52407 = ~n41407 & ~n52406;
  assign n52408 = ~i_hbusreq9 & ~n52407;
  assign n52409 = ~n52400 & ~n52408;
  assign n52410 = ~i_hbusreq4 & ~n52409;
  assign n52411 = ~n52399 & ~n52410;
  assign n52412 = ~controllable_hgrant4 & ~n52411;
  assign n52413 = ~n13208 & ~n52412;
  assign n52414 = ~i_hbusreq5 & ~n52413;
  assign n52415 = ~n52398 & ~n52414;
  assign n52416 = ~controllable_hgrant5 & ~n52415;
  assign n52417 = ~n13206 & ~n52416;
  assign n52418 = controllable_hmaster1 & ~n52417;
  assign n52419 = controllable_hmaster2 & ~n52417;
  assign n52420 = i_hbusreq5 & ~n52343;
  assign n52421 = i_hbusreq4 & ~n52341;
  assign n52422 = i_hbusreq9 & ~n52341;
  assign n52423 = i_hbusreq3 & ~n52339;
  assign n52424 = n8365 & ~n9015;
  assign n52425 = ~n8365 & ~n17420;
  assign n52426 = ~n52424 & ~n52425;
  assign n52427 = ~i_hbusreq3 & ~n52426;
  assign n52428 = ~n52423 & ~n52427;
  assign n52429 = controllable_hgrant3 & ~n52428;
  assign n52430 = ~n41448 & ~n52429;
  assign n52431 = ~i_hbusreq9 & ~n52430;
  assign n52432 = ~n52422 & ~n52431;
  assign n52433 = ~i_hbusreq4 & ~n52432;
  assign n52434 = ~n52421 & ~n52433;
  assign n52435 = ~controllable_hgrant4 & ~n52434;
  assign n52436 = ~n13258 & ~n52435;
  assign n52437 = ~i_hbusreq5 & ~n52436;
  assign n52438 = ~n52420 & ~n52437;
  assign n52439 = ~controllable_hgrant5 & ~n52438;
  assign n52440 = ~n13256 & ~n52439;
  assign n52441 = ~controllable_hmaster2 & ~n52440;
  assign n52442 = ~n52419 & ~n52441;
  assign n52443 = ~controllable_hmaster1 & ~n52442;
  assign n52444 = ~n52418 & ~n52443;
  assign n52445 = ~i_hbusreq6 & ~n52444;
  assign n52446 = ~n52397 & ~n52445;
  assign n52447 = ~controllable_hgrant6 & ~n52446;
  assign n52448 = ~n13254 & ~n52447;
  assign n52449 = ~i_hbusreq8 & ~n52448;
  assign n52450 = ~n52396 & ~n52449;
  assign n52451 = controllable_hmaster3 & ~n52450;
  assign n52452 = i_hbusreq8 & ~n52392;
  assign n52453 = i_hbusreq6 & ~n52355;
  assign n52454 = n8217 & ~n10119;
  assign n52455 = ~n8217 & ~n22569;
  assign n52456 = ~n52454 & ~n52455;
  assign n52457 = ~i_hbusreq6 & ~n52456;
  assign n52458 = ~n52453 & ~n52457;
  assign n52459 = controllable_hgrant6 & ~n52458;
  assign n52460 = i_hbusreq6 & ~n52370;
  assign n52461 = controllable_hmaster2 & ~n52440;
  assign n52462 = ~n48408 & ~n52461;
  assign n52463 = controllable_hmaster1 & ~n52462;
  assign n52464 = ~n41463 & ~n52439;
  assign n52465 = controllable_hmaster2 & ~n52464;
  assign n52466 = i_hbusreq5 & ~n52364;
  assign n52467 = i_hbusreq4 & ~n52362;
  assign n52468 = i_hbusreq9 & ~n52362;
  assign n52469 = ~n41476 & ~n52429;
  assign n52470 = ~i_hbusreq9 & ~n52469;
  assign n52471 = ~n52468 & ~n52470;
  assign n52472 = ~i_hbusreq4 & ~n52471;
  assign n52473 = ~n52467 & ~n52472;
  assign n52474 = ~controllable_hgrant4 & ~n52473;
  assign n52475 = ~n13258 & ~n52474;
  assign n52476 = ~i_hbusreq5 & ~n52475;
  assign n52477 = ~n52466 & ~n52476;
  assign n52478 = ~controllable_hgrant5 & ~n52477;
  assign n52479 = ~n13256 & ~n52478;
  assign n52480 = ~controllable_hmaster2 & ~n52479;
  assign n52481 = ~n52465 & ~n52480;
  assign n52482 = ~controllable_hmaster1 & ~n52481;
  assign n52483 = ~n52463 & ~n52482;
  assign n52484 = ~i_hbusreq6 & ~n52483;
  assign n52485 = ~n52460 & ~n52484;
  assign n52486 = ~controllable_hgrant6 & ~n52485;
  assign n52487 = ~n52459 & ~n52486;
  assign n52488 = controllable_hmaster0 & ~n52487;
  assign n52489 = i_hbusreq6 & ~n52388;
  assign n52490 = i_hbusreq5 & ~n52376;
  assign n52491 = i_hbusreq4 & ~n52374;
  assign n52492 = i_hbusreq9 & ~n52374;
  assign n52493 = ~n41515 & ~n52429;
  assign n52494 = ~i_hbusreq9 & ~n52493;
  assign n52495 = ~n52492 & ~n52494;
  assign n52496 = ~i_hbusreq4 & ~n52495;
  assign n52497 = ~n52491 & ~n52496;
  assign n52498 = ~controllable_hgrant4 & ~n52497;
  assign n52499 = ~n13258 & ~n52498;
  assign n52500 = ~i_hbusreq5 & ~n52499;
  assign n52501 = ~n52490 & ~n52500;
  assign n52502 = ~controllable_hgrant5 & ~n52501;
  assign n52503 = ~n13256 & ~n52502;
  assign n52504 = ~controllable_hmaster2 & ~n52503;
  assign n52505 = ~n52461 & ~n52504;
  assign n52506 = controllable_hmaster1 & ~n52505;
  assign n52507 = i_hbusreq5 & ~n52382;
  assign n52508 = ~n41531 & ~n52435;
  assign n52509 = ~i_hbusreq5 & ~n52508;
  assign n52510 = ~n52507 & ~n52509;
  assign n52511 = ~controllable_hgrant5 & ~n52510;
  assign n52512 = ~n13256 & ~n52511;
  assign n52513 = controllable_hmaster2 & ~n52512;
  assign n52514 = ~n52441 & ~n52513;
  assign n52515 = ~controllable_hmaster1 & ~n52514;
  assign n52516 = ~n52506 & ~n52515;
  assign n52517 = ~i_hbusreq6 & ~n52516;
  assign n52518 = ~n52489 & ~n52517;
  assign n52519 = ~controllable_hgrant6 & ~n52518;
  assign n52520 = ~n41497 & ~n52519;
  assign n52521 = ~controllable_hmaster0 & ~n52520;
  assign n52522 = ~n52488 & ~n52521;
  assign n52523 = ~i_hbusreq8 & ~n52522;
  assign n52524 = ~n52452 & ~n52523;
  assign n52525 = ~controllable_hmaster3 & ~n52524;
  assign n52526 = ~n52451 & ~n52525;
  assign n52527 = ~i_hbusreq7 & ~n52526;
  assign n52528 = ~n52395 & ~n52527;
  assign n52529 = ~n7924 & ~n52528;
  assign n52530 = ~n41572 & ~n48785;
  assign n52531 = ~controllable_hgrant4 & ~n52530;
  assign n52532 = ~n41560 & ~n52531;
  assign n52533 = ~controllable_hgrant5 & ~n52532;
  assign n52534 = ~n41559 & ~n52533;
  assign n52535 = controllable_hmaster1 & ~n52534;
  assign n52536 = controllable_hmaster2 & ~n52534;
  assign n52537 = n8365 & ~n13182;
  assign n52538 = ~n8365 & ~n17512;
  assign n52539 = ~n52537 & ~n52538;
  assign n52540 = i_hlock3 & ~n52539;
  assign n52541 = ~n8365 & ~n17520;
  assign n52542 = ~n52537 & ~n52541;
  assign n52543 = ~i_hlock3 & ~n52542;
  assign n52544 = ~n52540 & ~n52543;
  assign n52545 = controllable_hgrant3 & ~n52544;
  assign n52546 = ~n41660 & ~n52545;
  assign n52547 = ~controllable_hgrant4 & ~n52546;
  assign n52548 = ~n41648 & ~n52547;
  assign n52549 = ~controllable_hgrant5 & ~n52548;
  assign n52550 = ~n41647 & ~n52549;
  assign n52551 = ~controllable_hmaster2 & ~n52550;
  assign n52552 = ~n52536 & ~n52551;
  assign n52553 = ~controllable_hmaster1 & ~n52552;
  assign n52554 = ~n52535 & ~n52553;
  assign n52555 = ~controllable_hgrant6 & ~n52554;
  assign n52556 = ~n41646 & ~n52555;
  assign n52557 = controllable_hmaster3 & ~n52556;
  assign n52558 = n8217 & ~n15297;
  assign n52559 = ~n8217 & ~n22595;
  assign n52560 = ~n52558 & ~n52559;
  assign n52561 = controllable_hgrant6 & ~n52560;
  assign n52562 = controllable_hmaster2 & ~n52550;
  assign n52563 = ~n8378 & ~n22589;
  assign n52564 = ~n43910 & ~n52563;
  assign n52565 = controllable_hgrant5 & ~n52564;
  assign n52566 = ~n8426 & ~n22587;
  assign n52567 = ~n43914 & ~n52566;
  assign n52568 = controllable_hgrant4 & ~n52567;
  assign n52569 = i_hlock3 & ~n41616;
  assign n52570 = ~i_hlock3 & ~n41630;
  assign n52571 = ~n52569 & ~n52570;
  assign n52572 = ~controllable_hgrant3 & ~n52571;
  assign n52573 = ~n48859 & ~n52572;
  assign n52574 = ~controllable_hgrant4 & ~n52573;
  assign n52575 = ~n52568 & ~n52574;
  assign n52576 = ~controllable_hgrant5 & ~n52575;
  assign n52577 = ~n52565 & ~n52576;
  assign n52578 = ~controllable_hmaster2 & ~n52577;
  assign n52579 = ~n52562 & ~n52578;
  assign n52580 = controllable_hmaster1 & ~n52579;
  assign n52581 = ~n41686 & ~n52549;
  assign n52582 = controllable_hmaster2 & ~n52581;
  assign n52583 = ~n41691 & ~n52545;
  assign n52584 = ~controllable_hgrant4 & ~n52583;
  assign n52585 = ~n41648 & ~n52584;
  assign n52586 = ~controllable_hgrant5 & ~n52585;
  assign n52587 = ~n41647 & ~n52586;
  assign n52588 = ~controllable_hmaster2 & ~n52587;
  assign n52589 = ~n52582 & ~n52588;
  assign n52590 = ~controllable_hmaster1 & ~n52589;
  assign n52591 = ~n52580 & ~n52590;
  assign n52592 = ~controllable_hgrant6 & ~n52591;
  assign n52593 = ~n52561 & ~n52592;
  assign n52594 = controllable_hmaster0 & ~n52593;
  assign n52595 = ~n41715 & ~n52545;
  assign n52596 = ~controllable_hgrant4 & ~n52595;
  assign n52597 = ~n41648 & ~n52596;
  assign n52598 = ~controllable_hgrant5 & ~n52597;
  assign n52599 = ~n41647 & ~n52598;
  assign n52600 = ~controllable_hmaster2 & ~n52599;
  assign n52601 = ~n52562 & ~n52600;
  assign n52602 = controllable_hmaster1 & ~n52601;
  assign n52603 = ~n41724 & ~n52547;
  assign n52604 = ~controllable_hgrant5 & ~n52603;
  assign n52605 = ~n41647 & ~n52604;
  assign n52606 = controllable_hmaster2 & ~n52605;
  assign n52607 = ~n52551 & ~n52606;
  assign n52608 = ~controllable_hmaster1 & ~n52607;
  assign n52609 = ~n52602 & ~n52608;
  assign n52610 = ~controllable_hgrant6 & ~n52609;
  assign n52611 = ~n41704 & ~n52610;
  assign n52612 = ~controllable_hmaster0 & ~n52611;
  assign n52613 = ~n52594 & ~n52612;
  assign n52614 = ~controllable_hmaster3 & ~n52613;
  assign n52615 = ~n52557 & ~n52614;
  assign n52616 = i_hbusreq7 & ~n52615;
  assign n52617 = i_hbusreq8 & ~n52556;
  assign n52618 = i_hbusreq6 & ~n52554;
  assign n52619 = i_hbusreq5 & ~n52532;
  assign n52620 = i_hbusreq4 & ~n52530;
  assign n52621 = i_hbusreq9 & ~n52530;
  assign n52622 = n8365 & ~n13229;
  assign n52623 = ~n8365 & ~n17571;
  assign n52624 = ~n52622 & ~n52623;
  assign n52625 = i_hlock3 & ~n52624;
  assign n52626 = ~n8365 & ~n17593;
  assign n52627 = ~n52622 & ~n52626;
  assign n52628 = ~i_hlock3 & ~n52627;
  assign n52629 = ~n52625 & ~n52628;
  assign n52630 = ~i_hbusreq3 & ~n52629;
  assign n52631 = ~n49134 & ~n52630;
  assign n52632 = controllable_hgrant3 & ~n52631;
  assign n52633 = ~n41771 & ~n52632;
  assign n52634 = ~i_hbusreq9 & ~n52633;
  assign n52635 = ~n52621 & ~n52634;
  assign n52636 = ~i_hbusreq4 & ~n52635;
  assign n52637 = ~n52620 & ~n52636;
  assign n52638 = ~controllable_hgrant4 & ~n52637;
  assign n52639 = ~n41750 & ~n52638;
  assign n52640 = ~i_hbusreq5 & ~n52639;
  assign n52641 = ~n52619 & ~n52640;
  assign n52642 = ~controllable_hgrant5 & ~n52641;
  assign n52643 = ~n41748 & ~n52642;
  assign n52644 = controllable_hmaster1 & ~n52643;
  assign n52645 = controllable_hmaster2 & ~n52643;
  assign n52646 = i_hbusreq5 & ~n52548;
  assign n52647 = i_hbusreq4 & ~n52546;
  assign n52648 = i_hbusreq9 & ~n52546;
  assign n52649 = i_hbusreq3 & ~n52544;
  assign n52650 = n8365 & ~n13269;
  assign n52651 = ~n8365 & ~n17646;
  assign n52652 = ~n52650 & ~n52651;
  assign n52653 = i_hlock3 & ~n52652;
  assign n52654 = ~n8365 & ~n17660;
  assign n52655 = ~n52650 & ~n52654;
  assign n52656 = ~i_hlock3 & ~n52655;
  assign n52657 = ~n52653 & ~n52656;
  assign n52658 = ~i_hbusreq3 & ~n52657;
  assign n52659 = ~n52649 & ~n52658;
  assign n52660 = controllable_hgrant3 & ~n52659;
  assign n52661 = ~n41936 & ~n52660;
  assign n52662 = ~i_hbusreq9 & ~n52661;
  assign n52663 = ~n52648 & ~n52662;
  assign n52664 = ~i_hbusreq4 & ~n52663;
  assign n52665 = ~n52647 & ~n52664;
  assign n52666 = ~controllable_hgrant4 & ~n52665;
  assign n52667 = ~n41911 & ~n52666;
  assign n52668 = ~i_hbusreq5 & ~n52667;
  assign n52669 = ~n52646 & ~n52668;
  assign n52670 = ~controllable_hgrant5 & ~n52669;
  assign n52671 = ~n41909 & ~n52670;
  assign n52672 = ~controllable_hmaster2 & ~n52671;
  assign n52673 = ~n52645 & ~n52672;
  assign n52674 = ~controllable_hmaster1 & ~n52673;
  assign n52675 = ~n52644 & ~n52674;
  assign n52676 = ~i_hbusreq6 & ~n52675;
  assign n52677 = ~n52618 & ~n52676;
  assign n52678 = ~controllable_hgrant6 & ~n52677;
  assign n52679 = ~n41907 & ~n52678;
  assign n52680 = ~i_hbusreq8 & ~n52679;
  assign n52681 = ~n52617 & ~n52680;
  assign n52682 = controllable_hmaster3 & ~n52681;
  assign n52683 = i_hbusreq8 & ~n52613;
  assign n52684 = i_hbusreq6 & ~n52560;
  assign n52685 = n8217 & ~n15329;
  assign n52686 = ~n8217 & ~n22629;
  assign n52687 = ~n52685 & ~n52686;
  assign n52688 = ~i_hbusreq6 & ~n52687;
  assign n52689 = ~n52684 & ~n52688;
  assign n52690 = controllable_hgrant6 & ~n52689;
  assign n52691 = i_hbusreq6 & ~n52591;
  assign n52692 = controllable_hmaster2 & ~n52671;
  assign n52693 = i_hbusreq5 & ~n52564;
  assign n52694 = n8378 & ~n15321;
  assign n52695 = ~n8378 & ~n22621;
  assign n52696 = ~n52694 & ~n52695;
  assign n52697 = ~i_hbusreq5 & ~n52696;
  assign n52698 = ~n52693 & ~n52697;
  assign n52699 = controllable_hgrant5 & ~n52698;
  assign n52700 = i_hbusreq5 & ~n52575;
  assign n52701 = i_hbusreq4 & ~n52567;
  assign n52702 = i_hbusreq9 & ~n52567;
  assign n52703 = n8426 & ~n15315;
  assign n52704 = ~n8426 & ~n22615;
  assign n52705 = ~n52703 & ~n52704;
  assign n52706 = ~i_hbusreq9 & ~n52705;
  assign n52707 = ~n52702 & ~n52706;
  assign n52708 = ~i_hbusreq4 & ~n52707;
  assign n52709 = ~n52701 & ~n52708;
  assign n52710 = controllable_hgrant4 & ~n52709;
  assign n52711 = i_hbusreq4 & ~n52573;
  assign n52712 = i_hbusreq9 & ~n52573;
  assign n52713 = i_hbusreq3 & ~n52571;
  assign n52714 = i_hlock3 & ~n41855;
  assign n52715 = ~i_hlock3 & ~n41881;
  assign n52716 = ~n52714 & ~n52715;
  assign n52717 = ~i_hbusreq3 & ~n52716;
  assign n52718 = ~n52713 & ~n52717;
  assign n52719 = ~controllable_hgrant3 & ~n52718;
  assign n52720 = ~n49534 & ~n52719;
  assign n52721 = ~i_hbusreq9 & ~n52720;
  assign n52722 = ~n52712 & ~n52721;
  assign n52723 = ~i_hbusreq4 & ~n52722;
  assign n52724 = ~n52711 & ~n52723;
  assign n52725 = ~controllable_hgrant4 & ~n52724;
  assign n52726 = ~n52710 & ~n52725;
  assign n52727 = ~i_hbusreq5 & ~n52726;
  assign n52728 = ~n52700 & ~n52727;
  assign n52729 = ~controllable_hgrant5 & ~n52728;
  assign n52730 = ~n52699 & ~n52729;
  assign n52731 = ~controllable_hmaster2 & ~n52730;
  assign n52732 = ~n52692 & ~n52731;
  assign n52733 = controllable_hmaster1 & ~n52732;
  assign n52734 = ~n41983 & ~n52670;
  assign n52735 = controllable_hmaster2 & ~n52734;
  assign n52736 = i_hbusreq5 & ~n52585;
  assign n52737 = i_hbusreq4 & ~n52583;
  assign n52738 = i_hbusreq9 & ~n52583;
  assign n52739 = ~n41994 & ~n52660;
  assign n52740 = ~i_hbusreq9 & ~n52739;
  assign n52741 = ~n52738 & ~n52740;
  assign n52742 = ~i_hbusreq4 & ~n52741;
  assign n52743 = ~n52737 & ~n52742;
  assign n52744 = ~controllable_hgrant4 & ~n52743;
  assign n52745 = ~n41911 & ~n52744;
  assign n52746 = ~i_hbusreq5 & ~n52745;
  assign n52747 = ~n52736 & ~n52746;
  assign n52748 = ~controllable_hgrant5 & ~n52747;
  assign n52749 = ~n41909 & ~n52748;
  assign n52750 = ~controllable_hmaster2 & ~n52749;
  assign n52751 = ~n52735 & ~n52750;
  assign n52752 = ~controllable_hmaster1 & ~n52751;
  assign n52753 = ~n52733 & ~n52752;
  assign n52754 = ~i_hbusreq6 & ~n52753;
  assign n52755 = ~n52691 & ~n52754;
  assign n52756 = ~controllable_hgrant6 & ~n52755;
  assign n52757 = ~n52690 & ~n52756;
  assign n52758 = controllable_hmaster0 & ~n52757;
  assign n52759 = i_hbusreq6 & ~n52609;
  assign n52760 = i_hbusreq5 & ~n52597;
  assign n52761 = i_hbusreq4 & ~n52595;
  assign n52762 = i_hbusreq9 & ~n52595;
  assign n52763 = ~n42036 & ~n52660;
  assign n52764 = ~i_hbusreq9 & ~n52763;
  assign n52765 = ~n52762 & ~n52764;
  assign n52766 = ~i_hbusreq4 & ~n52765;
  assign n52767 = ~n52761 & ~n52766;
  assign n52768 = ~controllable_hgrant4 & ~n52767;
  assign n52769 = ~n41911 & ~n52768;
  assign n52770 = ~i_hbusreq5 & ~n52769;
  assign n52771 = ~n52760 & ~n52770;
  assign n52772 = ~controllable_hgrant5 & ~n52771;
  assign n52773 = ~n41909 & ~n52772;
  assign n52774 = ~controllable_hmaster2 & ~n52773;
  assign n52775 = ~n52692 & ~n52774;
  assign n52776 = controllable_hmaster1 & ~n52775;
  assign n52777 = i_hbusreq5 & ~n52603;
  assign n52778 = ~n42052 & ~n52666;
  assign n52779 = ~i_hbusreq5 & ~n52778;
  assign n52780 = ~n52777 & ~n52779;
  assign n52781 = ~controllable_hgrant5 & ~n52780;
  assign n52782 = ~n41909 & ~n52781;
  assign n52783 = controllable_hmaster2 & ~n52782;
  assign n52784 = ~n52672 & ~n52783;
  assign n52785 = ~controllable_hmaster1 & ~n52784;
  assign n52786 = ~n52776 & ~n52785;
  assign n52787 = ~i_hbusreq6 & ~n52786;
  assign n52788 = ~n52759 & ~n52787;
  assign n52789 = ~controllable_hgrant6 & ~n52788;
  assign n52790 = ~n42015 & ~n52789;
  assign n52791 = ~controllable_hmaster0 & ~n52790;
  assign n52792 = ~n52758 & ~n52791;
  assign n52793 = ~i_hbusreq8 & ~n52792;
  assign n52794 = ~n52683 & ~n52793;
  assign n52795 = ~controllable_hmaster3 & ~n52794;
  assign n52796 = ~n52682 & ~n52795;
  assign n52797 = ~i_hbusreq7 & ~n52796;
  assign n52798 = ~n52616 & ~n52797;
  assign n52799 = n7924 & ~n52798;
  assign n52800 = ~n52529 & ~n52799;
  assign n52801 = ~n8214 & ~n52800;
  assign n52802 = ~n12628 & ~n40226;
  assign n52803 = n7733 & ~n52802;
  assign n52804 = ~n51361 & ~n52803;
  assign n52805 = ~n7928 & ~n52804;
  assign n52806 = ~n48020 & ~n52803;
  assign n52807 = n7928 & ~n52806;
  assign n52808 = ~n52805 & ~n52807;
  assign n52809 = ~controllable_hgrant1 & ~n52808;
  assign n52810 = ~n13155 & ~n52809;
  assign n52811 = ~controllable_hgrant3 & ~n52810;
  assign n52812 = ~n13154 & ~n52811;
  assign n52813 = ~controllable_hgrant4 & ~n52812;
  assign n52814 = ~n13153 & ~n52813;
  assign n52815 = ~controllable_hgrant5 & ~n52814;
  assign n52816 = ~n13152 & ~n52815;
  assign n52817 = controllable_hmaster1 & ~n52816;
  assign n52818 = controllable_hmaster2 & ~n52816;
  assign n52819 = ~n40219 & ~n41350;
  assign n52820 = ~n7733 & ~n52819;
  assign n52821 = ~n40226 & ~n41350;
  assign n52822 = n7733 & ~n52821;
  assign n52823 = ~n52820 & ~n52822;
  assign n52824 = n7928 & ~n52823;
  assign n52825 = n7928 & ~n52824;
  assign n52826 = ~controllable_hgrant1 & ~n52825;
  assign n52827 = ~n13179 & ~n52826;
  assign n52828 = ~controllable_hgrant3 & ~n52827;
  assign n52829 = ~n13178 & ~n52828;
  assign n52830 = ~controllable_hgrant4 & ~n52829;
  assign n52831 = ~n13177 & ~n52830;
  assign n52832 = ~controllable_hgrant5 & ~n52831;
  assign n52833 = ~n13176 & ~n52832;
  assign n52834 = ~controllable_hmaster2 & ~n52833;
  assign n52835 = ~n52818 & ~n52834;
  assign n52836 = ~controllable_hmaster1 & ~n52835;
  assign n52837 = ~n52817 & ~n52836;
  assign n52838 = ~controllable_hgrant6 & ~n52837;
  assign n52839 = ~n13175 & ~n52838;
  assign n52840 = controllable_hmaster3 & ~n52839;
  assign n52841 = controllable_hmaster2 & ~n52833;
  assign n52842 = ~n41318 & ~n52828;
  assign n52843 = ~controllable_hgrant4 & ~n52842;
  assign n52844 = ~n13177 & ~n52843;
  assign n52845 = ~controllable_hgrant5 & ~n52844;
  assign n52846 = ~n13176 & ~n52845;
  assign n52847 = ~controllable_hmaster2 & ~n52846;
  assign n52848 = ~n52841 & ~n52847;
  assign n52849 = controllable_hmaster1 & ~n52848;
  assign n52850 = ~n41328 & ~n52832;
  assign n52851 = controllable_hmaster2 & ~n52850;
  assign n52852 = ~n41332 & ~n52826;
  assign n52853 = ~controllable_hgrant3 & ~n52852;
  assign n52854 = ~n13178 & ~n52853;
  assign n52855 = ~controllable_hgrant4 & ~n52854;
  assign n52856 = ~n13177 & ~n52855;
  assign n52857 = ~controllable_hgrant5 & ~n52856;
  assign n52858 = ~n13176 & ~n52857;
  assign n52859 = ~controllable_hmaster2 & ~n52858;
  assign n52860 = ~n52851 & ~n52859;
  assign n52861 = ~controllable_hmaster1 & ~n52860;
  assign n52862 = ~n52849 & ~n52861;
  assign n52863 = ~controllable_hgrant6 & ~n52862;
  assign n52864 = ~n13198 & ~n52863;
  assign n52865 = controllable_hmaster0 & ~n52864;
  assign n52866 = ~n9215 & ~n26888;
  assign n52867 = controllable_hmaster1 & ~n52866;
  assign n52868 = ~n9096 & ~n52867;
  assign n52869 = n8217 & ~n52868;
  assign n52870 = ~n18159 & ~n26888;
  assign n52871 = controllable_hmaster1 & ~n52870;
  assign n52872 = ~n9096 & ~n52871;
  assign n52873 = ~n8217 & ~n52872;
  assign n52874 = ~n52869 & ~n52873;
  assign n52875 = controllable_hgrant6 & ~n52874;
  assign n52876 = ~n48164 & ~n52841;
  assign n52877 = controllable_hmaster1 & ~n52876;
  assign n52878 = ~n41365 & ~n52830;
  assign n52879 = ~controllable_hgrant5 & ~n52878;
  assign n52880 = ~n13176 & ~n52879;
  assign n52881 = controllable_hmaster2 & ~n52880;
  assign n52882 = ~n52834 & ~n52881;
  assign n52883 = ~controllable_hmaster1 & ~n52882;
  assign n52884 = ~n52877 & ~n52883;
  assign n52885 = ~controllable_hgrant6 & ~n52884;
  assign n52886 = ~n52875 & ~n52885;
  assign n52887 = ~controllable_hmaster0 & ~n52886;
  assign n52888 = ~n52865 & ~n52887;
  assign n52889 = ~controllable_hmaster3 & ~n52888;
  assign n52890 = ~n52840 & ~n52889;
  assign n52891 = i_hbusreq7 & ~n52890;
  assign n52892 = i_hbusreq8 & ~n52839;
  assign n52893 = i_hbusreq6 & ~n52837;
  assign n52894 = i_hbusreq5 & ~n52814;
  assign n52895 = i_hbusreq4 & ~n52812;
  assign n52896 = i_hbusreq9 & ~n52812;
  assign n52897 = i_hbusreq3 & ~n52810;
  assign n52898 = i_hbusreq1 & ~n52808;
  assign n52899 = ~controllable_hmastlock & ~n43659;
  assign n52900 = controllable_locked & ~n52899;
  assign n52901 = ~n40321 & ~n52900;
  assign n52902 = ~i_hbusreq0 & ~n52901;
  assign n52903 = ~n40334 & ~n52902;
  assign n52904 = ~i_hbusreq2 & ~n52903;
  assign n52905 = ~n40333 & ~n52904;
  assign n52906 = controllable_hgrant2 & ~n52905;
  assign n52907 = ~n13347 & ~n52906;
  assign n52908 = n7733 & ~n52907;
  assign n52909 = ~n51400 & ~n52908;
  assign n52910 = ~n7928 & ~n52909;
  assign n52911 = ~n51404 & ~n52908;
  assign n52912 = n7928 & ~n52911;
  assign n52913 = ~n52910 & ~n52912;
  assign n52914 = ~i_hbusreq1 & ~n52913;
  assign n52915 = ~n52898 & ~n52914;
  assign n52916 = ~controllable_hgrant1 & ~n52915;
  assign n52917 = ~n13213 & ~n52916;
  assign n52918 = ~i_hbusreq3 & ~n52917;
  assign n52919 = ~n52897 & ~n52918;
  assign n52920 = ~controllable_hgrant3 & ~n52919;
  assign n52921 = ~n13211 & ~n52920;
  assign n52922 = ~i_hbusreq9 & ~n52921;
  assign n52923 = ~n52896 & ~n52922;
  assign n52924 = ~i_hbusreq4 & ~n52923;
  assign n52925 = ~n52895 & ~n52924;
  assign n52926 = ~controllable_hgrant4 & ~n52925;
  assign n52927 = ~n13208 & ~n52926;
  assign n52928 = ~i_hbusreq5 & ~n52927;
  assign n52929 = ~n52894 & ~n52928;
  assign n52930 = ~controllable_hgrant5 & ~n52929;
  assign n52931 = ~n13206 & ~n52930;
  assign n52932 = controllable_hmaster1 & ~n52931;
  assign n52933 = controllable_hmaster2 & ~n52931;
  assign n52934 = i_hbusreq5 & ~n52831;
  assign n52935 = i_hbusreq4 & ~n52829;
  assign n52936 = i_hbusreq9 & ~n52829;
  assign n52937 = i_hbusreq3 & ~n52827;
  assign n52938 = i_hbusreq1 & ~n52825;
  assign n52939 = ~i_hbusreq0 & ~n40322;
  assign n52940 = ~n40319 & ~n52939;
  assign n52941 = ~i_hbusreq2 & ~n52940;
  assign n52942 = ~n40318 & ~n52941;
  assign n52943 = controllable_hgrant2 & ~n52942;
  assign n52944 = ~n41505 & ~n52943;
  assign n52945 = ~n7733 & ~n52944;
  assign n52946 = ~n41505 & ~n52906;
  assign n52947 = n7733 & ~n52946;
  assign n52948 = ~n52945 & ~n52947;
  assign n52949 = n7928 & ~n52948;
  assign n52950 = n7928 & ~n52949;
  assign n52951 = ~i_hbusreq1 & ~n52950;
  assign n52952 = ~n52938 & ~n52951;
  assign n52953 = ~controllable_hgrant1 & ~n52952;
  assign n52954 = ~n13263 & ~n52953;
  assign n52955 = ~i_hbusreq3 & ~n52954;
  assign n52956 = ~n52937 & ~n52955;
  assign n52957 = ~controllable_hgrant3 & ~n52956;
  assign n52958 = ~n13261 & ~n52957;
  assign n52959 = ~i_hbusreq9 & ~n52958;
  assign n52960 = ~n52936 & ~n52959;
  assign n52961 = ~i_hbusreq4 & ~n52960;
  assign n52962 = ~n52935 & ~n52961;
  assign n52963 = ~controllable_hgrant4 & ~n52962;
  assign n52964 = ~n13258 & ~n52963;
  assign n52965 = ~i_hbusreq5 & ~n52964;
  assign n52966 = ~n52934 & ~n52965;
  assign n52967 = ~controllable_hgrant5 & ~n52966;
  assign n52968 = ~n13256 & ~n52967;
  assign n52969 = ~controllable_hmaster2 & ~n52968;
  assign n52970 = ~n52933 & ~n52969;
  assign n52971 = ~controllable_hmaster1 & ~n52970;
  assign n52972 = ~n52932 & ~n52971;
  assign n52973 = ~i_hbusreq6 & ~n52972;
  assign n52974 = ~n52893 & ~n52973;
  assign n52975 = ~controllable_hgrant6 & ~n52974;
  assign n52976 = ~n13254 & ~n52975;
  assign n52977 = ~i_hbusreq8 & ~n52976;
  assign n52978 = ~n52892 & ~n52977;
  assign n52979 = controllable_hmaster3 & ~n52978;
  assign n52980 = i_hbusreq8 & ~n52888;
  assign n52981 = i_hbusreq6 & ~n52862;
  assign n52982 = controllable_hmaster2 & ~n52968;
  assign n52983 = i_hbusreq5 & ~n52844;
  assign n52984 = i_hbusreq4 & ~n52842;
  assign n52985 = i_hbusreq9 & ~n52842;
  assign n52986 = ~n41447 & ~n52957;
  assign n52987 = ~i_hbusreq9 & ~n52986;
  assign n52988 = ~n52985 & ~n52987;
  assign n52989 = ~i_hbusreq4 & ~n52988;
  assign n52990 = ~n52984 & ~n52989;
  assign n52991 = ~controllable_hgrant4 & ~n52990;
  assign n52992 = ~n13258 & ~n52991;
  assign n52993 = ~i_hbusreq5 & ~n52992;
  assign n52994 = ~n52983 & ~n52993;
  assign n52995 = ~controllable_hgrant5 & ~n52994;
  assign n52996 = ~n13256 & ~n52995;
  assign n52997 = ~controllable_hmaster2 & ~n52996;
  assign n52998 = ~n52982 & ~n52997;
  assign n52999 = controllable_hmaster1 & ~n52998;
  assign n53000 = ~n41463 & ~n52967;
  assign n53001 = controllable_hmaster2 & ~n53000;
  assign n53002 = i_hbusreq5 & ~n52856;
  assign n53003 = i_hbusreq4 & ~n52854;
  assign n53004 = i_hbusreq9 & ~n52854;
  assign n53005 = i_hbusreq3 & ~n52852;
  assign n53006 = ~n41471 & ~n52953;
  assign n53007 = ~i_hbusreq3 & ~n53006;
  assign n53008 = ~n53005 & ~n53007;
  assign n53009 = ~controllable_hgrant3 & ~n53008;
  assign n53010 = ~n13261 & ~n53009;
  assign n53011 = ~i_hbusreq9 & ~n53010;
  assign n53012 = ~n53004 & ~n53011;
  assign n53013 = ~i_hbusreq4 & ~n53012;
  assign n53014 = ~n53003 & ~n53013;
  assign n53015 = ~controllable_hgrant4 & ~n53014;
  assign n53016 = ~n13258 & ~n53015;
  assign n53017 = ~i_hbusreq5 & ~n53016;
  assign n53018 = ~n53002 & ~n53017;
  assign n53019 = ~controllable_hgrant5 & ~n53018;
  assign n53020 = ~n13256 & ~n53019;
  assign n53021 = ~controllable_hmaster2 & ~n53020;
  assign n53022 = ~n53001 & ~n53021;
  assign n53023 = ~controllable_hmaster1 & ~n53022;
  assign n53024 = ~n52999 & ~n53023;
  assign n53025 = ~i_hbusreq6 & ~n53024;
  assign n53026 = ~n52981 & ~n53025;
  assign n53027 = ~controllable_hgrant6 & ~n53026;
  assign n53028 = ~n13298 & ~n53027;
  assign n53029 = controllable_hmaster0 & ~n53028;
  assign n53030 = i_hbusreq6 & ~n52874;
  assign n53031 = ~n9678 & ~n26901;
  assign n53032 = controllable_hmaster1 & ~n53031;
  assign n53033 = ~n9122 & ~n53032;
  assign n53034 = n8217 & ~n53033;
  assign n53035 = ~n21759 & ~n26901;
  assign n53036 = controllable_hmaster1 & ~n53035;
  assign n53037 = ~n9122 & ~n53036;
  assign n53038 = ~n8217 & ~n53037;
  assign n53039 = ~n53034 & ~n53038;
  assign n53040 = ~i_hbusreq6 & ~n53039;
  assign n53041 = ~n53030 & ~n53040;
  assign n53042 = controllable_hgrant6 & ~n53041;
  assign n53043 = i_hbusreq6 & ~n52884;
  assign n53044 = ~n48606 & ~n52982;
  assign n53045 = controllable_hmaster1 & ~n53044;
  assign n53046 = i_hbusreq5 & ~n52878;
  assign n53047 = ~n41531 & ~n52963;
  assign n53048 = ~i_hbusreq5 & ~n53047;
  assign n53049 = ~n53046 & ~n53048;
  assign n53050 = ~controllable_hgrant5 & ~n53049;
  assign n53051 = ~n13256 & ~n53050;
  assign n53052 = controllable_hmaster2 & ~n53051;
  assign n53053 = ~n52969 & ~n53052;
  assign n53054 = ~controllable_hmaster1 & ~n53053;
  assign n53055 = ~n53045 & ~n53054;
  assign n53056 = ~i_hbusreq6 & ~n53055;
  assign n53057 = ~n53043 & ~n53056;
  assign n53058 = ~controllable_hgrant6 & ~n53057;
  assign n53059 = ~n53042 & ~n53058;
  assign n53060 = ~controllable_hmaster0 & ~n53059;
  assign n53061 = ~n53029 & ~n53060;
  assign n53062 = ~i_hbusreq8 & ~n53061;
  assign n53063 = ~n52980 & ~n53062;
  assign n53064 = ~controllable_hmaster3 & ~n53063;
  assign n53065 = ~n52979 & ~n53064;
  assign n53066 = ~i_hbusreq7 & ~n53065;
  assign n53067 = ~n52891 & ~n53066;
  assign n53068 = ~n7924 & ~n53067;
  assign n53069 = ~n12801 & ~n46060;
  assign n53070 = n7733 & ~n53069;
  assign n53071 = ~n48798 & ~n53070;
  assign n53072 = n7928 & ~n53071;
  assign n53073 = ~n52805 & ~n53072;
  assign n53074 = ~controllable_hgrant1 & ~n53073;
  assign n53075 = ~n41562 & ~n53074;
  assign n53076 = ~controllable_hgrant3 & ~n53075;
  assign n53077 = ~n41561 & ~n53076;
  assign n53078 = ~controllable_hgrant4 & ~n53077;
  assign n53079 = ~n41560 & ~n53078;
  assign n53080 = ~controllable_hgrant5 & ~n53079;
  assign n53081 = ~n41559 & ~n53080;
  assign n53082 = controllable_hmaster1 & ~n53081;
  assign n53083 = controllable_hmaster2 & ~n53081;
  assign n53084 = ~n41651 & ~n43761;
  assign n53085 = ~n7733 & ~n53084;
  assign n53086 = ~n13010 & ~n46060;
  assign n53087 = n7733 & ~n53086;
  assign n53088 = ~n53085 & ~n53087;
  assign n53089 = n7928 & ~n53088;
  assign n53090 = n7928 & ~n53089;
  assign n53091 = ~controllable_hgrant1 & ~n53090;
  assign n53092 = ~n41650 & ~n53091;
  assign n53093 = ~controllable_hgrant3 & ~n53092;
  assign n53094 = ~n41649 & ~n53093;
  assign n53095 = ~controllable_hgrant4 & ~n53094;
  assign n53096 = ~n41648 & ~n53095;
  assign n53097 = ~controllable_hgrant5 & ~n53096;
  assign n53098 = ~n41647 & ~n53097;
  assign n53099 = ~controllable_hmaster2 & ~n53098;
  assign n53100 = ~n53083 & ~n53099;
  assign n53101 = ~controllable_hmaster1 & ~n53100;
  assign n53102 = ~n53082 & ~n53101;
  assign n53103 = ~controllable_hgrant6 & ~n53102;
  assign n53104 = ~n41646 & ~n53103;
  assign n53105 = controllable_hmaster3 & ~n53104;
  assign n53106 = controllable_hmaster2 & ~n53098;
  assign n53107 = ~n41677 & ~n53093;
  assign n53108 = ~controllable_hgrant4 & ~n53107;
  assign n53109 = ~n41648 & ~n53108;
  assign n53110 = ~controllable_hgrant5 & ~n53109;
  assign n53111 = ~n41647 & ~n53110;
  assign n53112 = ~controllable_hmaster2 & ~n53111;
  assign n53113 = ~n53106 & ~n53112;
  assign n53114 = controllable_hmaster1 & ~n53113;
  assign n53115 = ~n41686 & ~n53097;
  assign n53116 = controllable_hmaster2 & ~n53115;
  assign n53117 = ~n41689 & ~n53091;
  assign n53118 = ~controllable_hgrant3 & ~n53117;
  assign n53119 = ~n41649 & ~n53118;
  assign n53120 = ~controllable_hgrant4 & ~n53119;
  assign n53121 = ~n41648 & ~n53120;
  assign n53122 = ~controllable_hgrant5 & ~n53121;
  assign n53123 = ~n41647 & ~n53122;
  assign n53124 = ~controllable_hmaster2 & ~n53123;
  assign n53125 = ~n53116 & ~n53124;
  assign n53126 = ~controllable_hmaster1 & ~n53125;
  assign n53127 = ~n53114 & ~n53126;
  assign n53128 = ~controllable_hgrant6 & ~n53127;
  assign n53129 = ~n41675 & ~n53128;
  assign n53130 = controllable_hmaster0 & ~n53129;
  assign n53131 = ~n13908 & ~n26934;
  assign n53132 = controllable_hmaster1 & ~n53131;
  assign n53133 = ~n13677 & ~n53132;
  assign n53134 = n8217 & ~n53133;
  assign n53135 = ~n22682 & ~n26934;
  assign n53136 = controllable_hmaster1 & ~n53135;
  assign n53137 = ~n13677 & ~n53136;
  assign n53138 = ~n8217 & ~n53137;
  assign n53139 = ~n53134 & ~n53138;
  assign n53140 = controllable_hgrant6 & ~n53139;
  assign n53141 = ~n8378 & ~n22679;
  assign n53142 = ~n44018 & ~n53141;
  assign n53143 = controllable_hgrant5 & ~n53142;
  assign n53144 = ~n8426 & ~n22677;
  assign n53145 = ~n44022 & ~n53144;
  assign n53146 = controllable_hgrant4 & ~n53145;
  assign n53147 = ~n8365 & ~n22675;
  assign n53148 = ~n44026 & ~n53147;
  assign n53149 = controllable_hgrant3 & ~n53148;
  assign n53150 = ~n8389 & ~n22673;
  assign n53151 = ~n44030 & ~n53150;
  assign n53152 = controllable_hgrant1 & ~n53151;
  assign n53153 = ~n41609 & ~n48978;
  assign n53154 = n7733 & ~n53153;
  assign n53155 = ~n48968 & ~n53154;
  assign n53156 = n7928 & ~n53155;
  assign n53157 = ~n42965 & ~n53156;
  assign n53158 = ~controllable_hgrant1 & ~n53157;
  assign n53159 = ~n53152 & ~n53158;
  assign n53160 = ~controllable_hgrant3 & ~n53159;
  assign n53161 = ~n53149 & ~n53160;
  assign n53162 = ~controllable_hgrant4 & ~n53161;
  assign n53163 = ~n53146 & ~n53162;
  assign n53164 = ~controllable_hgrant5 & ~n53163;
  assign n53165 = ~n53143 & ~n53164;
  assign n53166 = ~controllable_hmaster2 & ~n53165;
  assign n53167 = ~n53106 & ~n53166;
  assign n53168 = controllable_hmaster1 & ~n53167;
  assign n53169 = ~n41724 & ~n53095;
  assign n53170 = ~controllable_hgrant5 & ~n53169;
  assign n53171 = ~n41647 & ~n53170;
  assign n53172 = controllable_hmaster2 & ~n53171;
  assign n53173 = ~n53099 & ~n53172;
  assign n53174 = ~controllable_hmaster1 & ~n53173;
  assign n53175 = ~n53168 & ~n53174;
  assign n53176 = ~controllable_hgrant6 & ~n53175;
  assign n53177 = ~n53140 & ~n53176;
  assign n53178 = ~controllable_hmaster0 & ~n53177;
  assign n53179 = ~n53130 & ~n53178;
  assign n53180 = ~controllable_hmaster3 & ~n53179;
  assign n53181 = ~n53105 & ~n53180;
  assign n53182 = i_hbusreq7 & ~n53181;
  assign n53183 = i_hbusreq8 & ~n53104;
  assign n53184 = i_hbusreq6 & ~n53102;
  assign n53185 = i_hbusreq5 & ~n53079;
  assign n53186 = i_hbusreq4 & ~n53077;
  assign n53187 = i_hbusreq9 & ~n53077;
  assign n53188 = i_hbusreq3 & ~n53075;
  assign n53189 = i_hbusreq1 & ~n53073;
  assign n53190 = ~n39848 & ~n46690;
  assign n53191 = controllable_locked & ~n53190;
  assign n53192 = ~n51512 & ~n53191;
  assign n53193 = ~i_hbusreq0 & ~n53192;
  assign n53194 = ~n46689 & ~n53193;
  assign n53195 = i_hlock2 & ~n53194;
  assign n53196 = ~n46700 & ~n53193;
  assign n53197 = ~i_hlock2 & ~n53196;
  assign n53198 = ~n53195 & ~n53197;
  assign n53199 = ~i_hbusreq2 & ~n53198;
  assign n53200 = ~n46688 & ~n53199;
  assign n53201 = controllable_hgrant2 & ~n53200;
  assign n53202 = ~n13489 & ~n53201;
  assign n53203 = n7733 & ~n53202;
  assign n53204 = ~n51522 & ~n53203;
  assign n53205 = n7928 & ~n53204;
  assign n53206 = ~n52910 & ~n53205;
  assign n53207 = ~i_hbusreq1 & ~n53206;
  assign n53208 = ~n53189 & ~n53207;
  assign n53209 = ~controllable_hgrant1 & ~n53208;
  assign n53210 = ~n41755 & ~n53209;
  assign n53211 = ~i_hbusreq3 & ~n53210;
  assign n53212 = ~n53188 & ~n53211;
  assign n53213 = ~controllable_hgrant3 & ~n53212;
  assign n53214 = ~n41753 & ~n53213;
  assign n53215 = ~i_hbusreq9 & ~n53214;
  assign n53216 = ~n53187 & ~n53215;
  assign n53217 = ~i_hbusreq4 & ~n53216;
  assign n53218 = ~n53186 & ~n53217;
  assign n53219 = ~controllable_hgrant4 & ~n53218;
  assign n53220 = ~n41750 & ~n53219;
  assign n53221 = ~i_hbusreq5 & ~n53220;
  assign n53222 = ~n53185 & ~n53221;
  assign n53223 = ~controllable_hgrant5 & ~n53222;
  assign n53224 = ~n41748 & ~n53223;
  assign n53225 = controllable_hmaster1 & ~n53224;
  assign n53226 = controllable_hmaster2 & ~n53224;
  assign n53227 = i_hbusreq5 & ~n53096;
  assign n53228 = i_hbusreq4 & ~n53094;
  assign n53229 = i_hbusreq9 & ~n53094;
  assign n53230 = i_hbusreq3 & ~n53092;
  assign n53231 = i_hbusreq1 & ~n53090;
  assign n53232 = ~controllable_locked & ~n51512;
  assign n53233 = ~i_hlock0 & ~n53232;
  assign n53234 = ~n44184 & ~n53233;
  assign n53235 = ~i_hbusreq0 & ~n53234;
  assign n53236 = ~n44181 & ~n53235;
  assign n53237 = ~i_hbusreq2 & ~n53236;
  assign n53238 = ~n44180 & ~n53237;
  assign n53239 = controllable_hgrant2 & ~n53238;
  assign n53240 = ~n41923 & ~n53239;
  assign n53241 = ~n7733 & ~n53240;
  assign n53242 = ~n13457 & ~n53201;
  assign n53243 = n7733 & ~n53242;
  assign n53244 = ~n53241 & ~n53243;
  assign n53245 = n7928 & ~n53244;
  assign n53246 = n7928 & ~n53245;
  assign n53247 = ~i_hbusreq1 & ~n53246;
  assign n53248 = ~n53231 & ~n53247;
  assign n53249 = ~controllable_hgrant1 & ~n53248;
  assign n53250 = ~n41916 & ~n53249;
  assign n53251 = ~i_hbusreq3 & ~n53250;
  assign n53252 = ~n53230 & ~n53251;
  assign n53253 = ~controllable_hgrant3 & ~n53252;
  assign n53254 = ~n41914 & ~n53253;
  assign n53255 = ~i_hbusreq9 & ~n53254;
  assign n53256 = ~n53229 & ~n53255;
  assign n53257 = ~i_hbusreq4 & ~n53256;
  assign n53258 = ~n53228 & ~n53257;
  assign n53259 = ~controllable_hgrant4 & ~n53258;
  assign n53260 = ~n41911 & ~n53259;
  assign n53261 = ~i_hbusreq5 & ~n53260;
  assign n53262 = ~n53227 & ~n53261;
  assign n53263 = ~controllable_hgrant5 & ~n53262;
  assign n53264 = ~n41909 & ~n53263;
  assign n53265 = ~controllable_hmaster2 & ~n53264;
  assign n53266 = ~n53226 & ~n53265;
  assign n53267 = ~controllable_hmaster1 & ~n53266;
  assign n53268 = ~n53225 & ~n53267;
  assign n53269 = ~i_hbusreq6 & ~n53268;
  assign n53270 = ~n53184 & ~n53269;
  assign n53271 = ~controllable_hgrant6 & ~n53270;
  assign n53272 = ~n41907 & ~n53271;
  assign n53273 = ~i_hbusreq8 & ~n53272;
  assign n53274 = ~n53183 & ~n53273;
  assign n53275 = controllable_hmaster3 & ~n53274;
  assign n53276 = i_hbusreq8 & ~n53179;
  assign n53277 = i_hbusreq6 & ~n53127;
  assign n53278 = controllable_hmaster2 & ~n53264;
  assign n53279 = i_hbusreq5 & ~n53109;
  assign n53280 = i_hbusreq4 & ~n53107;
  assign n53281 = i_hbusreq9 & ~n53107;
  assign n53282 = ~n41968 & ~n53253;
  assign n53283 = ~i_hbusreq9 & ~n53282;
  assign n53284 = ~n53281 & ~n53283;
  assign n53285 = ~i_hbusreq4 & ~n53284;
  assign n53286 = ~n53280 & ~n53285;
  assign n53287 = ~controllable_hgrant4 & ~n53286;
  assign n53288 = ~n41911 & ~n53287;
  assign n53289 = ~i_hbusreq5 & ~n53288;
  assign n53290 = ~n53279 & ~n53289;
  assign n53291 = ~controllable_hgrant5 & ~n53290;
  assign n53292 = ~n41909 & ~n53291;
  assign n53293 = ~controllable_hmaster2 & ~n53292;
  assign n53294 = ~n53278 & ~n53293;
  assign n53295 = controllable_hmaster1 & ~n53294;
  assign n53296 = ~n41983 & ~n53263;
  assign n53297 = controllable_hmaster2 & ~n53296;
  assign n53298 = i_hbusreq5 & ~n53121;
  assign n53299 = i_hbusreq4 & ~n53119;
  assign n53300 = i_hbusreq9 & ~n53119;
  assign n53301 = i_hbusreq3 & ~n53117;
  assign n53302 = ~n41990 & ~n53249;
  assign n53303 = ~i_hbusreq3 & ~n53302;
  assign n53304 = ~n53301 & ~n53303;
  assign n53305 = ~controllable_hgrant3 & ~n53304;
  assign n53306 = ~n41914 & ~n53305;
  assign n53307 = ~i_hbusreq9 & ~n53306;
  assign n53308 = ~n53300 & ~n53307;
  assign n53309 = ~i_hbusreq4 & ~n53308;
  assign n53310 = ~n53299 & ~n53309;
  assign n53311 = ~controllable_hgrant4 & ~n53310;
  assign n53312 = ~n41911 & ~n53311;
  assign n53313 = ~i_hbusreq5 & ~n53312;
  assign n53314 = ~n53298 & ~n53313;
  assign n53315 = ~controllable_hgrant5 & ~n53314;
  assign n53316 = ~n41909 & ~n53315;
  assign n53317 = ~controllable_hmaster2 & ~n53316;
  assign n53318 = ~n53297 & ~n53317;
  assign n53319 = ~controllable_hmaster1 & ~n53318;
  assign n53320 = ~n53295 & ~n53319;
  assign n53321 = ~i_hbusreq6 & ~n53320;
  assign n53322 = ~n53277 & ~n53321;
  assign n53323 = ~controllable_hgrant6 & ~n53322;
  assign n53324 = ~n41962 & ~n53323;
  assign n53325 = controllable_hmaster0 & ~n53324;
  assign n53326 = i_hbusreq6 & ~n53139;
  assign n53327 = ~n15384 & ~n26978;
  assign n53328 = controllable_hmaster1 & ~n53327;
  assign n53329 = ~n13721 & ~n53328;
  assign n53330 = n8217 & ~n53329;
  assign n53331 = ~n22719 & ~n26978;
  assign n53332 = controllable_hmaster1 & ~n53331;
  assign n53333 = ~n13721 & ~n53332;
  assign n53334 = ~n8217 & ~n53333;
  assign n53335 = ~n53330 & ~n53334;
  assign n53336 = ~i_hbusreq6 & ~n53335;
  assign n53337 = ~n53326 & ~n53336;
  assign n53338 = controllable_hgrant6 & ~n53337;
  assign n53339 = i_hbusreq6 & ~n53175;
  assign n53340 = i_hbusreq5 & ~n53142;
  assign n53341 = n8378 & ~n15379;
  assign n53342 = ~n8378 & ~n22714;
  assign n53343 = ~n53341 & ~n53342;
  assign n53344 = ~i_hbusreq5 & ~n53343;
  assign n53345 = ~n53340 & ~n53344;
  assign n53346 = controllable_hgrant5 & ~n53345;
  assign n53347 = i_hbusreq5 & ~n53163;
  assign n53348 = i_hbusreq4 & ~n53145;
  assign n53349 = i_hbusreq9 & ~n53145;
  assign n53350 = n8426 & ~n15373;
  assign n53351 = ~n8426 & ~n22708;
  assign n53352 = ~n53350 & ~n53351;
  assign n53353 = ~i_hbusreq9 & ~n53352;
  assign n53354 = ~n53349 & ~n53353;
  assign n53355 = ~i_hbusreq4 & ~n53354;
  assign n53356 = ~n53348 & ~n53355;
  assign n53357 = controllable_hgrant4 & ~n53356;
  assign n53358 = i_hbusreq4 & ~n53161;
  assign n53359 = i_hbusreq9 & ~n53161;
  assign n53360 = i_hbusreq3 & ~n53148;
  assign n53361 = n8365 & ~n15369;
  assign n53362 = ~n8365 & ~n22704;
  assign n53363 = ~n53361 & ~n53362;
  assign n53364 = ~i_hbusreq3 & ~n53363;
  assign n53365 = ~n53360 & ~n53364;
  assign n53366 = controllable_hgrant3 & ~n53365;
  assign n53367 = i_hbusreq3 & ~n53159;
  assign n53368 = i_hbusreq1 & ~n53151;
  assign n53369 = n8389 & ~n15365;
  assign n53370 = ~n8389 & ~n22700;
  assign n53371 = ~n53369 & ~n53370;
  assign n53372 = ~i_hbusreq1 & ~n53371;
  assign n53373 = ~n53368 & ~n53372;
  assign n53374 = controllable_hgrant1 & ~n53373;
  assign n53375 = i_hbusreq1 & ~n53157;
  assign n53376 = ~n41846 & ~n49770;
  assign n53377 = n7733 & ~n53376;
  assign n53378 = ~n51600 & ~n53377;
  assign n53379 = n7928 & ~n53378;
  assign n53380 = ~n43545 & ~n53379;
  assign n53381 = ~i_hbusreq1 & ~n53380;
  assign n53382 = ~n53375 & ~n53381;
  assign n53383 = ~controllable_hgrant1 & ~n53382;
  assign n53384 = ~n53374 & ~n53383;
  assign n53385 = ~i_hbusreq3 & ~n53384;
  assign n53386 = ~n53367 & ~n53385;
  assign n53387 = ~controllable_hgrant3 & ~n53386;
  assign n53388 = ~n53366 & ~n53387;
  assign n53389 = ~i_hbusreq9 & ~n53388;
  assign n53390 = ~n53359 & ~n53389;
  assign n53391 = ~i_hbusreq4 & ~n53390;
  assign n53392 = ~n53358 & ~n53391;
  assign n53393 = ~controllable_hgrant4 & ~n53392;
  assign n53394 = ~n53357 & ~n53393;
  assign n53395 = ~i_hbusreq5 & ~n53394;
  assign n53396 = ~n53347 & ~n53395;
  assign n53397 = ~controllable_hgrant5 & ~n53396;
  assign n53398 = ~n53346 & ~n53397;
  assign n53399 = ~controllable_hmaster2 & ~n53398;
  assign n53400 = ~n53278 & ~n53399;
  assign n53401 = controllable_hmaster1 & ~n53400;
  assign n53402 = i_hbusreq5 & ~n53169;
  assign n53403 = ~n42052 & ~n53259;
  assign n53404 = ~i_hbusreq5 & ~n53403;
  assign n53405 = ~n53402 & ~n53404;
  assign n53406 = ~controllable_hgrant5 & ~n53405;
  assign n53407 = ~n41909 & ~n53406;
  assign n53408 = controllable_hmaster2 & ~n53407;
  assign n53409 = ~n53265 & ~n53408;
  assign n53410 = ~controllable_hmaster1 & ~n53409;
  assign n53411 = ~n53401 & ~n53410;
  assign n53412 = ~i_hbusreq6 & ~n53411;
  assign n53413 = ~n53339 & ~n53412;
  assign n53414 = ~controllable_hgrant6 & ~n53413;
  assign n53415 = ~n53338 & ~n53414;
  assign n53416 = ~controllable_hmaster0 & ~n53415;
  assign n53417 = ~n53325 & ~n53416;
  assign n53418 = ~i_hbusreq8 & ~n53417;
  assign n53419 = ~n53276 & ~n53418;
  assign n53420 = ~controllable_hmaster3 & ~n53419;
  assign n53421 = ~n53275 & ~n53420;
  assign n53422 = ~i_hbusreq7 & ~n53421;
  assign n53423 = ~n53182 & ~n53422;
  assign n53424 = n7924 & ~n53423;
  assign n53425 = ~n53068 & ~n53424;
  assign n53426 = n8214 & ~n53425;
  assign n53427 = ~n52801 & ~n53426;
  assign n53428 = n8202 & ~n53427;
  assign n53429 = ~n52329 & ~n53428;
  assign n53430 = n7920 & ~n53429;
  assign n53431 = ~n50812 & ~n53430;
  assign n53432 = n7728 & ~n53431;
  assign n53433 = ~n42736 & ~n48008;
  assign n53434 = controllable_hmaster1 & ~n53433;
  assign n53435 = controllable_hmaster2 & ~n53433;
  assign n53436 = ~n40196 & ~n44957;
  assign n53437 = ~controllable_hmaster2 & ~n53436;
  assign n53438 = ~n53435 & ~n53437;
  assign n53439 = ~controllable_hmaster1 & ~n53438;
  assign n53440 = ~n53434 & ~n53439;
  assign n53441 = ~controllable_hgrant6 & ~n53440;
  assign n53442 = ~n44944 & ~n53441;
  assign n53443 = controllable_hmaster0 & ~n53442;
  assign n53444 = ~n40431 & ~n42770;
  assign n53445 = ~controllable_hmaster2 & ~n53444;
  assign n53446 = ~n53435 & ~n53445;
  assign n53447 = ~controllable_hmaster1 & ~n53446;
  assign n53448 = ~n53434 & ~n53447;
  assign n53449 = ~controllable_hgrant6 & ~n53448;
  assign n53450 = ~n42748 & ~n53449;
  assign n53451 = ~controllable_hmaster0 & ~n53450;
  assign n53452 = ~n53443 & ~n53451;
  assign n53453 = i_hlock8 & ~n53452;
  assign n53454 = ~n40453 & ~n42803;
  assign n53455 = ~controllable_hmaster2 & ~n53454;
  assign n53456 = ~n53435 & ~n53455;
  assign n53457 = ~controllable_hmaster1 & ~n53456;
  assign n53458 = ~n53434 & ~n53457;
  assign n53459 = ~controllable_hgrant6 & ~n53458;
  assign n53460 = ~n42783 & ~n53459;
  assign n53461 = ~controllable_hmaster0 & ~n53460;
  assign n53462 = ~n53443 & ~n53461;
  assign n53463 = ~i_hlock8 & ~n53462;
  assign n53464 = ~n53453 & ~n53463;
  assign n53465 = controllable_hmaster3 & ~n53464;
  assign n53466 = ~n8217 & ~n22746;
  assign n53467 = ~n42816 & ~n53466;
  assign n53468 = controllable_hgrant6 & ~n53467;
  assign n53469 = controllable_hmaster2 & ~n53444;
  assign n53470 = ~n42846 & ~n48060;
  assign n53471 = ~controllable_hmaster2 & ~n53470;
  assign n53472 = ~n53469 & ~n53471;
  assign n53473 = controllable_hmaster1 & ~n53472;
  assign n53474 = ~n42898 & ~n48100;
  assign n53475 = ~controllable_hmaster2 & ~n53474;
  assign n53476 = ~n48097 & ~n53475;
  assign n53477 = ~controllable_hmaster1 & ~n53476;
  assign n53478 = ~n53473 & ~n53477;
  assign n53479 = ~controllable_hgrant6 & ~n53478;
  assign n53480 = ~n53468 & ~n53479;
  assign n53481 = controllable_hmaster0 & ~n53480;
  assign n53482 = ~n42982 & ~n48135;
  assign n53483 = ~controllable_hmaster2 & ~n53482;
  assign n53484 = ~n53469 & ~n53483;
  assign n53485 = controllable_hmaster1 & ~n53484;
  assign n53486 = ~n43006 & ~n48169;
  assign n53487 = controllable_hmaster2 & ~n53486;
  assign n53488 = ~n43032 & ~n48188;
  assign n53489 = ~controllable_hmaster2 & ~n53488;
  assign n53490 = ~n53487 & ~n53489;
  assign n53491 = ~controllable_hmaster1 & ~n53490;
  assign n53492 = ~n53485 & ~n53491;
  assign n53493 = i_hlock6 & ~n53492;
  assign n53494 = controllable_hmaster2 & ~n53454;
  assign n53495 = ~n53483 & ~n53494;
  assign n53496 = controllable_hmaster1 & ~n53495;
  assign n53497 = ~n53491 & ~n53496;
  assign n53498 = ~i_hlock6 & ~n53497;
  assign n53499 = ~n53493 & ~n53498;
  assign n53500 = ~controllable_hgrant6 & ~n53499;
  assign n53501 = ~n42928 & ~n53500;
  assign n53502 = ~controllable_hmaster0 & ~n53501;
  assign n53503 = ~n53481 & ~n53502;
  assign n53504 = ~controllable_hmaster3 & ~n53503;
  assign n53505 = ~n53465 & ~n53504;
  assign n53506 = i_hlock7 & ~n53505;
  assign n53507 = ~n8217 & ~n22754;
  assign n53508 = ~n43052 & ~n53507;
  assign n53509 = controllable_hgrant6 & ~n53508;
  assign n53510 = ~n53471 & ~n53494;
  assign n53511 = controllable_hmaster1 & ~n53510;
  assign n53512 = ~n53477 & ~n53511;
  assign n53513 = ~controllable_hgrant6 & ~n53512;
  assign n53514 = ~n53509 & ~n53513;
  assign n53515 = controllable_hmaster0 & ~n53514;
  assign n53516 = ~n53502 & ~n53515;
  assign n53517 = ~controllable_hmaster3 & ~n53516;
  assign n53518 = ~n53465 & ~n53517;
  assign n53519 = ~i_hlock7 & ~n53518;
  assign n53520 = ~n53506 & ~n53519;
  assign n53521 = i_hbusreq7 & ~n53520;
  assign n53522 = i_hbusreq8 & ~n53464;
  assign n53523 = i_hbusreq6 & ~n53440;
  assign n53524 = ~n8378 & ~n18242;
  assign n53525 = ~n43078 & ~n53524;
  assign n53526 = ~i_hbusreq5 & ~n53525;
  assign n53527 = ~n48244 & ~n53526;
  assign n53528 = controllable_hgrant5 & ~n53527;
  assign n53529 = ~n43144 & ~n53528;
  assign n53530 = controllable_hmaster1 & ~n53529;
  assign n53531 = controllable_hmaster2 & ~n53529;
  assign n53532 = ~n8378 & ~n30184;
  assign n53533 = ~n45006 & ~n53532;
  assign n53534 = ~i_hbusreq5 & ~n53533;
  assign n53535 = ~n40276 & ~n53534;
  assign n53536 = controllable_hgrant5 & ~n53535;
  assign n53537 = ~n45036 & ~n53536;
  assign n53538 = ~controllable_hmaster2 & ~n53537;
  assign n53539 = ~n53531 & ~n53538;
  assign n53540 = ~controllable_hmaster1 & ~n53539;
  assign n53541 = ~n53530 & ~n53540;
  assign n53542 = ~i_hbusreq6 & ~n53541;
  assign n53543 = ~n53523 & ~n53542;
  assign n53544 = ~controllable_hgrant6 & ~n53543;
  assign n53545 = ~n45003 & ~n53544;
  assign n53546 = controllable_hmaster0 & ~n53545;
  assign n53547 = i_hbusreq6 & ~n53448;
  assign n53548 = ~n8378 & ~n18274;
  assign n53549 = ~n43165 & ~n53548;
  assign n53550 = ~i_hbusreq5 & ~n53549;
  assign n53551 = ~n40481 & ~n53550;
  assign n53552 = controllable_hgrant5 & ~n53551;
  assign n53553 = ~n43219 & ~n53552;
  assign n53554 = ~controllable_hmaster2 & ~n53553;
  assign n53555 = ~n53531 & ~n53554;
  assign n53556 = ~controllable_hmaster1 & ~n53555;
  assign n53557 = ~n53530 & ~n53556;
  assign n53558 = ~i_hbusreq6 & ~n53557;
  assign n53559 = ~n53547 & ~n53558;
  assign n53560 = ~controllable_hgrant6 & ~n53559;
  assign n53561 = ~n43162 & ~n53560;
  assign n53562 = ~controllable_hmaster0 & ~n53561;
  assign n53563 = ~n53546 & ~n53562;
  assign n53564 = i_hlock8 & ~n53563;
  assign n53565 = i_hbusreq6 & ~n53458;
  assign n53566 = ~n8378 & ~n18305;
  assign n53567 = ~n43241 & ~n53566;
  assign n53568 = ~i_hbusreq5 & ~n53567;
  assign n53569 = ~n40527 & ~n53568;
  assign n53570 = controllable_hgrant5 & ~n53569;
  assign n53571 = ~n43293 & ~n53570;
  assign n53572 = ~controllable_hmaster2 & ~n53571;
  assign n53573 = ~n53531 & ~n53572;
  assign n53574 = ~controllable_hmaster1 & ~n53573;
  assign n53575 = ~n53530 & ~n53574;
  assign n53576 = ~i_hbusreq6 & ~n53575;
  assign n53577 = ~n53565 & ~n53576;
  assign n53578 = ~controllable_hgrant6 & ~n53577;
  assign n53579 = ~n43238 & ~n53578;
  assign n53580 = ~controllable_hmaster0 & ~n53579;
  assign n53581 = ~n53546 & ~n53580;
  assign n53582 = ~i_hlock8 & ~n53581;
  assign n53583 = ~n53564 & ~n53582;
  assign n53584 = ~i_hbusreq8 & ~n53583;
  assign n53585 = ~n53522 & ~n53584;
  assign n53586 = controllable_hmaster3 & ~n53585;
  assign n53587 = i_hbusreq8 & ~n53503;
  assign n53588 = i_hbusreq6 & ~n53467;
  assign n53589 = n8217 & ~n10163;
  assign n53590 = ~n8217 & ~n22768;
  assign n53591 = ~n53589 & ~n53590;
  assign n53592 = ~i_hbusreq6 & ~n53591;
  assign n53593 = ~n53588 & ~n53592;
  assign n53594 = controllable_hgrant6 & ~n53593;
  assign n53595 = i_hbusreq6 & ~n53478;
  assign n53596 = controllable_hmaster2 & ~n53553;
  assign n53597 = ~n8378 & ~n18344;
  assign n53598 = ~n43321 & ~n53597;
  assign n53599 = ~i_hbusreq5 & ~n53598;
  assign n53600 = ~n48357 & ~n53599;
  assign n53601 = controllable_hgrant5 & ~n53600;
  assign n53602 = ~n43369 & ~n53601;
  assign n53603 = ~controllable_hmaster2 & ~n53602;
  assign n53604 = ~n53596 & ~n53603;
  assign n53605 = controllable_hmaster1 & ~n53604;
  assign n53606 = ~n8378 & ~n18382;
  assign n53607 = ~n43397 & ~n53606;
  assign n53608 = ~i_hbusreq5 & ~n53607;
  assign n53609 = ~n48433 & ~n53608;
  assign n53610 = controllable_hgrant5 & ~n53609;
  assign n53611 = ~n43457 & ~n53610;
  assign n53612 = ~controllable_hmaster2 & ~n53611;
  assign n53613 = ~n48432 & ~n53612;
  assign n53614 = ~controllable_hmaster1 & ~n53613;
  assign n53615 = ~n53605 & ~n53614;
  assign n53616 = ~i_hbusreq6 & ~n53615;
  assign n53617 = ~n53595 & ~n53616;
  assign n53618 = ~controllable_hgrant6 & ~n53617;
  assign n53619 = ~n53594 & ~n53618;
  assign n53620 = controllable_hmaster0 & ~n53619;
  assign n53621 = i_hbusreq6 & ~n53499;
  assign n53622 = ~n8378 & ~n18416;
  assign n53623 = ~n43495 & ~n53622;
  assign n53624 = ~i_hbusreq5 & ~n53623;
  assign n53625 = ~n48530 & ~n53624;
  assign n53626 = controllable_hgrant5 & ~n53625;
  assign n53627 = ~n43578 & ~n53626;
  assign n53628 = ~controllable_hmaster2 & ~n53627;
  assign n53629 = ~n53596 & ~n53628;
  assign n53630 = controllable_hmaster1 & ~n53629;
  assign n53631 = ~n8378 & ~n18432;
  assign n53632 = ~n43584 & ~n53631;
  assign n53633 = ~i_hbusreq5 & ~n53632;
  assign n53634 = ~n48609 & ~n53633;
  assign n53635 = controllable_hgrant5 & ~n53634;
  assign n53636 = ~n43620 & ~n53635;
  assign n53637 = controllable_hmaster2 & ~n53636;
  assign n53638 = ~n8378 & ~n18483;
  assign n53639 = ~n43624 & ~n53638;
  assign n53640 = ~i_hbusreq5 & ~n53639;
  assign n53641 = ~n48649 & ~n53640;
  assign n53642 = controllable_hgrant5 & ~n53641;
  assign n53643 = ~n43689 & ~n53642;
  assign n53644 = ~controllable_hmaster2 & ~n53643;
  assign n53645 = ~n53637 & ~n53644;
  assign n53646 = ~controllable_hmaster1 & ~n53645;
  assign n53647 = ~n53630 & ~n53646;
  assign n53648 = i_hlock6 & ~n53647;
  assign n53649 = controllable_hmaster2 & ~n53571;
  assign n53650 = ~n53628 & ~n53649;
  assign n53651 = controllable_hmaster1 & ~n53650;
  assign n53652 = ~n53646 & ~n53651;
  assign n53653 = ~i_hlock6 & ~n53652;
  assign n53654 = ~n53648 & ~n53653;
  assign n53655 = ~i_hbusreq6 & ~n53654;
  assign n53656 = ~n53621 & ~n53655;
  assign n53657 = ~controllable_hgrant6 & ~n53656;
  assign n53658 = ~n43492 & ~n53657;
  assign n53659 = ~controllable_hmaster0 & ~n53658;
  assign n53660 = ~n53620 & ~n53659;
  assign n53661 = ~i_hbusreq8 & ~n53660;
  assign n53662 = ~n53587 & ~n53661;
  assign n53663 = ~controllable_hmaster3 & ~n53662;
  assign n53664 = ~n53586 & ~n53663;
  assign n53665 = i_hlock7 & ~n53664;
  assign n53666 = i_hbusreq8 & ~n53516;
  assign n53667 = i_hbusreq6 & ~n53508;
  assign n53668 = n8217 & ~n10173;
  assign n53669 = ~n8217 & ~n22782;
  assign n53670 = ~n53668 & ~n53669;
  assign n53671 = ~i_hbusreq6 & ~n53670;
  assign n53672 = ~n53667 & ~n53671;
  assign n53673 = controllable_hgrant6 & ~n53672;
  assign n53674 = i_hbusreq6 & ~n53512;
  assign n53675 = ~n53603 & ~n53649;
  assign n53676 = controllable_hmaster1 & ~n53675;
  assign n53677 = ~n53614 & ~n53676;
  assign n53678 = ~i_hbusreq6 & ~n53677;
  assign n53679 = ~n53674 & ~n53678;
  assign n53680 = ~controllable_hgrant6 & ~n53679;
  assign n53681 = ~n53673 & ~n53680;
  assign n53682 = controllable_hmaster0 & ~n53681;
  assign n53683 = ~n53659 & ~n53682;
  assign n53684 = ~i_hbusreq8 & ~n53683;
  assign n53685 = ~n53666 & ~n53684;
  assign n53686 = ~controllable_hmaster3 & ~n53685;
  assign n53687 = ~n53586 & ~n53686;
  assign n53688 = ~i_hlock7 & ~n53687;
  assign n53689 = ~n53665 & ~n53688;
  assign n53690 = ~i_hbusreq7 & ~n53689;
  assign n53691 = ~n53521 & ~n53690;
  assign n53692 = ~n7924 & ~n53691;
  assign n53693 = ~n43774 & ~n48769;
  assign n53694 = controllable_hmaster1 & ~n53693;
  assign n53695 = controllable_hmaster2 & ~n53693;
  assign n53696 = ~n45110 & ~n46012;
  assign n53697 = ~controllable_hmaster2 & ~n53696;
  assign n53698 = ~n53695 & ~n53697;
  assign n53699 = ~controllable_hmaster1 & ~n53698;
  assign n53700 = ~n53694 & ~n53699;
  assign n53701 = ~controllable_hgrant6 & ~n53700;
  assign n53702 = ~n45097 & ~n53701;
  assign n53703 = controllable_hmaster0 & ~n53702;
  assign n53704 = ~n43859 & ~n47528;
  assign n53705 = ~controllable_hmaster2 & ~n53704;
  assign n53706 = ~n53695 & ~n53705;
  assign n53707 = ~controllable_hmaster1 & ~n53706;
  assign n53708 = ~n53694 & ~n53707;
  assign n53709 = ~controllable_hgrant6 & ~n53708;
  assign n53710 = ~n43833 & ~n53709;
  assign n53711 = ~controllable_hmaster0 & ~n53710;
  assign n53712 = ~n53703 & ~n53711;
  assign n53713 = i_hlock8 & ~n53712;
  assign n53714 = ~n43892 & ~n47561;
  assign n53715 = ~controllable_hmaster2 & ~n53714;
  assign n53716 = ~n53695 & ~n53715;
  assign n53717 = ~controllable_hmaster1 & ~n53716;
  assign n53718 = ~n53694 & ~n53717;
  assign n53719 = ~controllable_hgrant6 & ~n53718;
  assign n53720 = ~n43872 & ~n53719;
  assign n53721 = ~controllable_hmaster0 & ~n53720;
  assign n53722 = ~n53703 & ~n53721;
  assign n53723 = ~i_hlock8 & ~n53722;
  assign n53724 = ~n53713 & ~n53723;
  assign n53725 = controllable_hmaster3 & ~n53724;
  assign n53726 = ~n8217 & ~n22806;
  assign n53727 = ~n43905 & ~n53726;
  assign n53728 = controllable_hgrant6 & ~n53727;
  assign n53729 = controllable_hmaster2 & ~n53704;
  assign n53730 = ~n43935 & ~n48843;
  assign n53731 = ~controllable_hmaster2 & ~n53730;
  assign n53732 = ~n53729 & ~n53731;
  assign n53733 = controllable_hmaster1 & ~n53732;
  assign n53734 = i_hlock5 & ~n45127;
  assign n53735 = ~i_hlock5 & ~n45147;
  assign n53736 = ~n53734 & ~n53735;
  assign n53737 = ~controllable_hgrant5 & ~n53736;
  assign n53738 = ~n48879 & ~n53737;
  assign n53739 = controllable_hmaster2 & ~n53738;
  assign n53740 = ~n43987 & ~n48893;
  assign n53741 = ~controllable_hmaster2 & ~n53740;
  assign n53742 = ~n53739 & ~n53741;
  assign n53743 = ~controllable_hmaster1 & ~n53742;
  assign n53744 = ~n53733 & ~n53743;
  assign n53745 = ~controllable_hgrant6 & ~n53744;
  assign n53746 = ~n53728 & ~n53745;
  assign n53747 = controllable_hmaster0 & ~n53746;
  assign n53748 = ~n44049 & ~n48943;
  assign n53749 = ~controllable_hmaster2 & ~n53748;
  assign n53750 = ~n53729 & ~n53749;
  assign n53751 = controllable_hmaster1 & ~n53750;
  assign n53752 = ~n44073 & ~n49001;
  assign n53753 = controllable_hmaster2 & ~n53752;
  assign n53754 = ~n44099 & ~n49025;
  assign n53755 = ~controllable_hmaster2 & ~n53754;
  assign n53756 = ~n53753 & ~n53755;
  assign n53757 = ~controllable_hmaster1 & ~n53756;
  assign n53758 = ~n53751 & ~n53757;
  assign n53759 = i_hlock6 & ~n53758;
  assign n53760 = controllable_hmaster2 & ~n53714;
  assign n53761 = ~n53749 & ~n53760;
  assign n53762 = controllable_hmaster1 & ~n53761;
  assign n53763 = ~n53757 & ~n53762;
  assign n53764 = ~i_hlock6 & ~n53763;
  assign n53765 = ~n53759 & ~n53764;
  assign n53766 = ~controllable_hgrant6 & ~n53765;
  assign n53767 = ~n44017 & ~n53766;
  assign n53768 = ~controllable_hmaster0 & ~n53767;
  assign n53769 = ~n53747 & ~n53768;
  assign n53770 = ~controllable_hmaster3 & ~n53769;
  assign n53771 = ~n53725 & ~n53770;
  assign n53772 = i_hlock7 & ~n53771;
  assign n53773 = ~n8217 & ~n22814;
  assign n53774 = ~n44119 & ~n53773;
  assign n53775 = controllable_hgrant6 & ~n53774;
  assign n53776 = ~n53731 & ~n53760;
  assign n53777 = controllable_hmaster1 & ~n53776;
  assign n53778 = ~n53743 & ~n53777;
  assign n53779 = ~controllable_hgrant6 & ~n53778;
  assign n53780 = ~n53775 & ~n53779;
  assign n53781 = controllable_hmaster0 & ~n53780;
  assign n53782 = ~n53768 & ~n53781;
  assign n53783 = ~controllable_hmaster3 & ~n53782;
  assign n53784 = ~n53725 & ~n53783;
  assign n53785 = ~i_hlock7 & ~n53784;
  assign n53786 = ~n53772 & ~n53785;
  assign n53787 = i_hbusreq7 & ~n53786;
  assign n53788 = i_hbusreq8 & ~n53724;
  assign n53789 = i_hbusreq6 & ~n53700;
  assign n53790 = n8378 & ~n14004;
  assign n53791 = ~n8378 & ~n30457;
  assign n53792 = ~n53790 & ~n53791;
  assign n53793 = i_hlock5 & ~n53792;
  assign n53794 = ~n8378 & ~n30665;
  assign n53795 = ~n53790 & ~n53794;
  assign n53796 = ~i_hlock5 & ~n53795;
  assign n53797 = ~n53793 & ~n53796;
  assign n53798 = ~i_hbusreq5 & ~n53797;
  assign n53799 = ~n49101 & ~n53798;
  assign n53800 = controllable_hgrant5 & ~n53799;
  assign n53801 = ~n44221 & ~n53800;
  assign n53802 = controllable_hmaster1 & ~n53801;
  assign n53803 = controllable_hmaster2 & ~n53801;
  assign n53804 = n8378 & ~n27481;
  assign n53805 = ~n8378 & ~n30474;
  assign n53806 = ~n53804 & ~n53805;
  assign n53807 = i_hlock5 & ~n53806;
  assign n53808 = ~n8378 & ~n30682;
  assign n53809 = ~n53804 & ~n53808;
  assign n53810 = ~i_hlock5 & ~n53809;
  assign n53811 = ~n53807 & ~n53810;
  assign n53812 = ~i_hbusreq5 & ~n53811;
  assign n53813 = ~n46623 & ~n53812;
  assign n53814 = controllable_hgrant5 & ~n53813;
  assign n53815 = ~n45207 & ~n53814;
  assign n53816 = ~controllable_hmaster2 & ~n53815;
  assign n53817 = ~n53803 & ~n53816;
  assign n53818 = ~controllable_hmaster1 & ~n53817;
  assign n53819 = ~n53802 & ~n53818;
  assign n53820 = ~i_hbusreq6 & ~n53819;
  assign n53821 = ~n53789 & ~n53820;
  assign n53822 = ~controllable_hgrant6 & ~n53821;
  assign n53823 = ~n45174 & ~n53822;
  assign n53824 = controllable_hmaster0 & ~n53823;
  assign n53825 = i_hbusreq6 & ~n53708;
  assign n53826 = n8378 & ~n14038;
  assign n53827 = ~n8378 & ~n30497;
  assign n53828 = ~n53826 & ~n53827;
  assign n53829 = i_hlock5 & ~n53828;
  assign n53830 = ~n8378 & ~n30705;
  assign n53831 = ~n53826 & ~n53830;
  assign n53832 = ~i_hlock5 & ~n53831;
  assign n53833 = ~n53829 & ~n53832;
  assign n53834 = ~i_hbusreq5 & ~n53833;
  assign n53835 = ~n47667 & ~n53834;
  assign n53836 = controllable_hgrant5 & ~n53835;
  assign n53837 = ~n44429 & ~n53836;
  assign n53838 = ~controllable_hmaster2 & ~n53837;
  assign n53839 = ~n53803 & ~n53838;
  assign n53840 = ~controllable_hmaster1 & ~n53839;
  assign n53841 = ~n53802 & ~n53840;
  assign n53842 = ~i_hbusreq6 & ~n53841;
  assign n53843 = ~n53825 & ~n53842;
  assign n53844 = ~controllable_hgrant6 & ~n53843;
  assign n53845 = ~n44368 & ~n53844;
  assign n53846 = ~controllable_hmaster0 & ~n53845;
  assign n53847 = ~n53824 & ~n53846;
  assign n53848 = i_hlock8 & ~n53847;
  assign n53849 = i_hbusreq6 & ~n53718;
  assign n53850 = n8378 & ~n14073;
  assign n53851 = ~n8378 & ~n30522;
  assign n53852 = ~n53850 & ~n53851;
  assign n53853 = i_hlock5 & ~n53852;
  assign n53854 = ~n8378 & ~n30730;
  assign n53855 = ~n53850 & ~n53854;
  assign n53856 = ~i_hlock5 & ~n53855;
  assign n53857 = ~n53853 & ~n53856;
  assign n53858 = ~i_hbusreq5 & ~n53857;
  assign n53859 = ~n47727 & ~n53858;
  assign n53860 = controllable_hgrant5 & ~n53859;
  assign n53861 = ~n44503 & ~n53860;
  assign n53862 = ~controllable_hmaster2 & ~n53861;
  assign n53863 = ~n53803 & ~n53862;
  assign n53864 = ~controllable_hmaster1 & ~n53863;
  assign n53865 = ~n53802 & ~n53864;
  assign n53866 = ~i_hbusreq6 & ~n53865;
  assign n53867 = ~n53849 & ~n53866;
  assign n53868 = ~controllable_hgrant6 & ~n53867;
  assign n53869 = ~n44448 & ~n53868;
  assign n53870 = ~controllable_hmaster0 & ~n53869;
  assign n53871 = ~n53824 & ~n53870;
  assign n53872 = ~i_hlock8 & ~n53871;
  assign n53873 = ~n53848 & ~n53872;
  assign n53874 = ~i_hbusreq8 & ~n53873;
  assign n53875 = ~n53788 & ~n53874;
  assign n53876 = controllable_hmaster3 & ~n53875;
  assign n53877 = i_hbusreq8 & ~n53769;
  assign n53878 = i_hbusreq6 & ~n53727;
  assign n53879 = n8217 & ~n15428;
  assign n53880 = ~n8217 & ~n22837;
  assign n53881 = ~n53879 & ~n53880;
  assign n53882 = ~i_hbusreq6 & ~n53881;
  assign n53883 = ~n53878 & ~n53882;
  assign n53884 = controllable_hgrant6 & ~n53883;
  assign n53885 = i_hbusreq6 & ~n53744;
  assign n53886 = controllable_hmaster2 & ~n53837;
  assign n53887 = n8378 & ~n14116;
  assign n53888 = ~n8378 & ~n30552;
  assign n53889 = ~n53887 & ~n53888;
  assign n53890 = i_hlock5 & ~n53889;
  assign n53891 = ~n8378 & ~n30760;
  assign n53892 = ~n53887 & ~n53891;
  assign n53893 = ~i_hlock5 & ~n53892;
  assign n53894 = ~n53890 & ~n53893;
  assign n53895 = ~i_hbusreq5 & ~n53894;
  assign n53896 = ~n49489 & ~n53895;
  assign n53897 = controllable_hgrant5 & ~n53896;
  assign n53898 = ~n44579 & ~n53897;
  assign n53899 = ~controllable_hmaster2 & ~n53898;
  assign n53900 = ~n53886 & ~n53899;
  assign n53901 = controllable_hmaster1 & ~n53900;
  assign n53902 = i_hbusreq5 & ~n53736;
  assign n53903 = i_hlock5 & ~n45248;
  assign n53904 = ~i_hlock5 & ~n45294;
  assign n53905 = ~n53903 & ~n53904;
  assign n53906 = ~i_hbusreq5 & ~n53905;
  assign n53907 = ~n53902 & ~n53906;
  assign n53908 = ~controllable_hgrant5 & ~n53907;
  assign n53909 = ~n49568 & ~n53908;
  assign n53910 = controllable_hmaster2 & ~n53909;
  assign n53911 = n8378 & ~n14159;
  assign n53912 = ~n8378 & ~n30577;
  assign n53913 = ~n53911 & ~n53912;
  assign n53914 = i_hlock5 & ~n53913;
  assign n53915 = ~n8378 & ~n30785;
  assign n53916 = ~n53911 & ~n53915;
  assign n53917 = ~i_hlock5 & ~n53916;
  assign n53918 = ~n53914 & ~n53917;
  assign n53919 = ~i_hbusreq5 & ~n53918;
  assign n53920 = ~n49578 & ~n53919;
  assign n53921 = controllable_hgrant5 & ~n53920;
  assign n53922 = ~n44667 & ~n53921;
  assign n53923 = ~controllable_hmaster2 & ~n53922;
  assign n53924 = ~n53910 & ~n53923;
  assign n53925 = ~controllable_hmaster1 & ~n53924;
  assign n53926 = ~n53901 & ~n53925;
  assign n53927 = ~i_hbusreq6 & ~n53926;
  assign n53928 = ~n53885 & ~n53927;
  assign n53929 = ~controllable_hgrant6 & ~n53928;
  assign n53930 = ~n53884 & ~n53929;
  assign n53931 = controllable_hmaster0 & ~n53930;
  assign n53932 = i_hbusreq6 & ~n53765;
  assign n53933 = n8378 & ~n14198;
  assign n53934 = ~n8378 & ~n30601;
  assign n53935 = ~n53933 & ~n53934;
  assign n53936 = i_hlock5 & ~n53935;
  assign n53937 = ~n8378 & ~n30809;
  assign n53938 = ~n53933 & ~n53937;
  assign n53939 = ~i_hlock5 & ~n53938;
  assign n53940 = ~n53936 & ~n53939;
  assign n53941 = ~i_hbusreq5 & ~n53940;
  assign n53942 = ~n49693 & ~n53941;
  assign n53943 = controllable_hgrant5 & ~n53942;
  assign n53944 = ~n44774 & ~n53943;
  assign n53945 = ~controllable_hmaster2 & ~n53944;
  assign n53946 = ~n53886 & ~n53945;
  assign n53947 = controllable_hmaster1 & ~n53946;
  assign n53948 = n8378 & ~n14216;
  assign n53949 = ~n8378 & ~n30617;
  assign n53950 = ~n53948 & ~n53949;
  assign n53951 = i_hlock5 & ~n53950;
  assign n53952 = ~n8378 & ~n30825;
  assign n53953 = ~n53948 & ~n53952;
  assign n53954 = ~i_hlock5 & ~n53953;
  assign n53955 = ~n53951 & ~n53954;
  assign n53956 = ~i_hbusreq5 & ~n53955;
  assign n53957 = ~n49797 & ~n53956;
  assign n53958 = controllable_hgrant5 & ~n53957;
  assign n53959 = ~n44816 & ~n53958;
  assign n53960 = controllable_hmaster2 & ~n53959;
  assign n53961 = n8378 & ~n14270;
  assign n53962 = ~n8378 & ~n30631;
  assign n53963 = ~n53961 & ~n53962;
  assign n53964 = i_hlock5 & ~n53963;
  assign n53965 = ~n8378 & ~n30839;
  assign n53966 = ~n53961 & ~n53965;
  assign n53967 = ~i_hlock5 & ~n53966;
  assign n53968 = ~n53964 & ~n53967;
  assign n53969 = ~i_hbusreq5 & ~n53968;
  assign n53970 = ~n49842 & ~n53969;
  assign n53971 = controllable_hgrant5 & ~n53970;
  assign n53972 = ~n44889 & ~n53971;
  assign n53973 = ~controllable_hmaster2 & ~n53972;
  assign n53974 = ~n53960 & ~n53973;
  assign n53975 = ~controllable_hmaster1 & ~n53974;
  assign n53976 = ~n53947 & ~n53975;
  assign n53977 = i_hlock6 & ~n53976;
  assign n53978 = controllable_hmaster2 & ~n53861;
  assign n53979 = ~n53945 & ~n53978;
  assign n53980 = controllable_hmaster1 & ~n53979;
  assign n53981 = ~n53975 & ~n53980;
  assign n53982 = ~i_hlock6 & ~n53981;
  assign n53983 = ~n53977 & ~n53982;
  assign n53984 = ~i_hbusreq6 & ~n53983;
  assign n53985 = ~n53932 & ~n53984;
  assign n53986 = ~controllable_hgrant6 & ~n53985;
  assign n53987 = ~n44702 & ~n53986;
  assign n53988 = ~controllable_hmaster0 & ~n53987;
  assign n53989 = ~n53931 & ~n53988;
  assign n53990 = ~i_hbusreq8 & ~n53989;
  assign n53991 = ~n53877 & ~n53990;
  assign n53992 = ~controllable_hmaster3 & ~n53991;
  assign n53993 = ~n53876 & ~n53992;
  assign n53994 = i_hlock7 & ~n53993;
  assign n53995 = i_hbusreq8 & ~n53782;
  assign n53996 = i_hbusreq6 & ~n53774;
  assign n53997 = n8217 & ~n15441;
  assign n53998 = ~n8217 & ~n22851;
  assign n53999 = ~n53997 & ~n53998;
  assign n54000 = ~i_hbusreq6 & ~n53999;
  assign n54001 = ~n53996 & ~n54000;
  assign n54002 = controllable_hgrant6 & ~n54001;
  assign n54003 = i_hbusreq6 & ~n53778;
  assign n54004 = ~n53899 & ~n53978;
  assign n54005 = controllable_hmaster1 & ~n54004;
  assign n54006 = ~n53925 & ~n54005;
  assign n54007 = ~i_hbusreq6 & ~n54006;
  assign n54008 = ~n54003 & ~n54007;
  assign n54009 = ~controllable_hgrant6 & ~n54008;
  assign n54010 = ~n54002 & ~n54009;
  assign n54011 = controllable_hmaster0 & ~n54010;
  assign n54012 = ~n53988 & ~n54011;
  assign n54013 = ~i_hbusreq8 & ~n54012;
  assign n54014 = ~n53995 & ~n54013;
  assign n54015 = ~controllable_hmaster3 & ~n54014;
  assign n54016 = ~n53876 & ~n54015;
  assign n54017 = ~i_hlock7 & ~n54016;
  assign n54018 = ~n53994 & ~n54017;
  assign n54019 = ~i_hbusreq7 & ~n54018;
  assign n54020 = ~n53787 & ~n54019;
  assign n54021 = n7924 & ~n54020;
  assign n54022 = ~n53692 & ~n54021;
  assign n54023 = ~n8214 & ~n54022;
  assign n54024 = ~n42734 & ~n48011;
  assign n54025 = ~controllable_hgrant5 & ~n54024;
  assign n54026 = ~n42709 & ~n54025;
  assign n54027 = controllable_hmaster1 & ~n54026;
  assign n54028 = controllable_hmaster2 & ~n54026;
  assign n54029 = ~n40206 & ~n44955;
  assign n54030 = ~controllable_hgrant5 & ~n54029;
  assign n54031 = ~n44947 & ~n54030;
  assign n54032 = ~controllable_hmaster2 & ~n54031;
  assign n54033 = ~n54028 & ~n54032;
  assign n54034 = ~controllable_hmaster1 & ~n54033;
  assign n54035 = ~n54027 & ~n54034;
  assign n54036 = ~controllable_hgrant6 & ~n54035;
  assign n54037 = ~n44944 & ~n54036;
  assign n54038 = controllable_hmaster0 & ~n54037;
  assign n54039 = ~n40432 & ~n42768;
  assign n54040 = ~controllable_hgrant5 & ~n54039;
  assign n54041 = ~n42751 & ~n54040;
  assign n54042 = ~controllable_hmaster2 & ~n54041;
  assign n54043 = ~n54028 & ~n54042;
  assign n54044 = ~controllable_hmaster1 & ~n54043;
  assign n54045 = ~n54027 & ~n54044;
  assign n54046 = ~controllable_hgrant6 & ~n54045;
  assign n54047 = ~n42748 & ~n54046;
  assign n54048 = ~controllable_hmaster0 & ~n54047;
  assign n54049 = ~n54038 & ~n54048;
  assign n54050 = i_hlock8 & ~n54049;
  assign n54051 = ~n40454 & ~n42801;
  assign n54052 = ~controllable_hgrant5 & ~n54051;
  assign n54053 = ~n42786 & ~n54052;
  assign n54054 = ~controllable_hmaster2 & ~n54053;
  assign n54055 = ~n54028 & ~n54054;
  assign n54056 = ~controllable_hmaster1 & ~n54055;
  assign n54057 = ~n54027 & ~n54056;
  assign n54058 = ~controllable_hgrant6 & ~n54057;
  assign n54059 = ~n42783 & ~n54058;
  assign n54060 = ~controllable_hmaster0 & ~n54059;
  assign n54061 = ~n54038 & ~n54060;
  assign n54062 = ~i_hlock8 & ~n54061;
  assign n54063 = ~n54050 & ~n54062;
  assign n54064 = controllable_hmaster3 & ~n54063;
  assign n54065 = controllable_hmaster2 & ~n54041;
  assign n54066 = ~n42844 & ~n48063;
  assign n54067 = ~controllable_hgrant5 & ~n54066;
  assign n54068 = ~n42824 & ~n54067;
  assign n54069 = ~controllable_hmaster2 & ~n54068;
  assign n54070 = ~n54065 & ~n54069;
  assign n54071 = controllable_hmaster1 & ~n54070;
  assign n54072 = i_hlock5 & ~n54039;
  assign n54073 = ~i_hlock5 & ~n54051;
  assign n54074 = ~n54072 & ~n54073;
  assign n54075 = ~controllable_hgrant5 & ~n54074;
  assign n54076 = ~n42860 & ~n54075;
  assign n54077 = controllable_hmaster2 & ~n54076;
  assign n54078 = ~n42896 & ~n48103;
  assign n54079 = ~controllable_hgrant5 & ~n54078;
  assign n54080 = ~n42870 & ~n54079;
  assign n54081 = ~controllable_hmaster2 & ~n54080;
  assign n54082 = ~n54077 & ~n54081;
  assign n54083 = ~controllable_hmaster1 & ~n54082;
  assign n54084 = ~n54071 & ~n54083;
  assign n54085 = ~controllable_hgrant6 & ~n54084;
  assign n54086 = ~n42819 & ~n54085;
  assign n54087 = controllable_hmaster0 & ~n54086;
  assign n54088 = ~n22870 & ~n42912;
  assign n54089 = ~n8217 & ~n54088;
  assign n54090 = ~n42910 & ~n54089;
  assign n54091 = i_hlock6 & ~n54090;
  assign n54092 = ~n22870 & ~n42922;
  assign n54093 = ~n8217 & ~n54092;
  assign n54094 = ~n42920 & ~n54093;
  assign n54095 = ~i_hlock6 & ~n54094;
  assign n54096 = ~n54091 & ~n54095;
  assign n54097 = controllable_hgrant6 & ~n54096;
  assign n54098 = ~n42980 & ~n48138;
  assign n54099 = ~controllable_hgrant5 & ~n54098;
  assign n54100 = ~n42932 & ~n54099;
  assign n54101 = ~controllable_hmaster2 & ~n54100;
  assign n54102 = ~n54065 & ~n54101;
  assign n54103 = controllable_hmaster1 & ~n54102;
  assign n54104 = ~n43030 & ~n48191;
  assign n54105 = ~controllable_hgrant5 & ~n54104;
  assign n54106 = ~n43012 & ~n54105;
  assign n54107 = ~controllable_hmaster2 & ~n54106;
  assign n54108 = ~n48185 & ~n54107;
  assign n54109 = ~controllable_hmaster1 & ~n54108;
  assign n54110 = ~n54103 & ~n54109;
  assign n54111 = i_hlock6 & ~n54110;
  assign n54112 = controllable_hmaster2 & ~n54053;
  assign n54113 = ~n54101 & ~n54112;
  assign n54114 = controllable_hmaster1 & ~n54113;
  assign n54115 = ~n54109 & ~n54114;
  assign n54116 = ~i_hlock6 & ~n54115;
  assign n54117 = ~n54111 & ~n54116;
  assign n54118 = ~controllable_hgrant6 & ~n54117;
  assign n54119 = ~n54097 & ~n54118;
  assign n54120 = ~controllable_hmaster0 & ~n54119;
  assign n54121 = ~n54087 & ~n54120;
  assign n54122 = ~controllable_hmaster3 & ~n54121;
  assign n54123 = ~n54064 & ~n54122;
  assign n54124 = i_hlock7 & ~n54123;
  assign n54125 = ~n54069 & ~n54112;
  assign n54126 = controllable_hmaster1 & ~n54125;
  assign n54127 = ~n54083 & ~n54126;
  assign n54128 = ~controllable_hgrant6 & ~n54127;
  assign n54129 = ~n43055 & ~n54128;
  assign n54130 = controllable_hmaster0 & ~n54129;
  assign n54131 = ~n54120 & ~n54130;
  assign n54132 = ~controllable_hmaster3 & ~n54131;
  assign n54133 = ~n54064 & ~n54132;
  assign n54134 = ~i_hlock7 & ~n54133;
  assign n54135 = ~n54124 & ~n54134;
  assign n54136 = i_hbusreq7 & ~n54135;
  assign n54137 = i_hbusreq8 & ~n54063;
  assign n54138 = i_hbusreq6 & ~n54035;
  assign n54139 = i_hbusreq5 & ~n54024;
  assign n54140 = ~n8426 & ~n18236;
  assign n54141 = ~n43087 & ~n54140;
  assign n54142 = ~i_hbusreq9 & ~n54141;
  assign n54143 = ~n48253 & ~n54142;
  assign n54144 = ~i_hbusreq4 & ~n54143;
  assign n54145 = ~n48252 & ~n54144;
  assign n54146 = controllable_hgrant4 & ~n54145;
  assign n54147 = ~n43140 & ~n54146;
  assign n54148 = ~i_hbusreq5 & ~n54147;
  assign n54149 = ~n54139 & ~n54148;
  assign n54150 = ~controllable_hgrant5 & ~n54149;
  assign n54151 = ~n43083 & ~n54150;
  assign n54152 = controllable_hmaster1 & ~n54151;
  assign n54153 = controllable_hmaster2 & ~n54151;
  assign n54154 = i_hbusreq5 & ~n54029;
  assign n54155 = ~n8426 & ~n18268;
  assign n54156 = ~n43174 & ~n54155;
  assign n54157 = i_hlock9 & ~n54156;
  assign n54158 = ~n8426 & ~n18299;
  assign n54159 = ~n43250 & ~n54158;
  assign n54160 = ~i_hlock9 & ~n54159;
  assign n54161 = ~n54157 & ~n54160;
  assign n54162 = ~i_hbusreq9 & ~n54161;
  assign n54163 = ~n40285 & ~n54162;
  assign n54164 = ~i_hbusreq4 & ~n54163;
  assign n54165 = ~n40284 & ~n54164;
  assign n54166 = controllable_hgrant4 & ~n54165;
  assign n54167 = ~n45032 & ~n54166;
  assign n54168 = ~i_hbusreq5 & ~n54167;
  assign n54169 = ~n54154 & ~n54168;
  assign n54170 = ~controllable_hgrant5 & ~n54169;
  assign n54171 = ~n45011 & ~n54170;
  assign n54172 = ~controllable_hmaster2 & ~n54171;
  assign n54173 = ~n54153 & ~n54172;
  assign n54174 = ~controllable_hmaster1 & ~n54173;
  assign n54175 = ~n54152 & ~n54174;
  assign n54176 = ~i_hbusreq6 & ~n54175;
  assign n54177 = ~n54138 & ~n54176;
  assign n54178 = ~controllable_hgrant6 & ~n54177;
  assign n54179 = ~n45003 & ~n54178;
  assign n54180 = controllable_hmaster0 & ~n54179;
  assign n54181 = i_hbusreq6 & ~n54045;
  assign n54182 = i_hbusreq5 & ~n54039;
  assign n54183 = ~i_hbusreq9 & ~n54156;
  assign n54184 = ~n40490 & ~n54183;
  assign n54185 = ~i_hbusreq4 & ~n54184;
  assign n54186 = ~n40489 & ~n54185;
  assign n54187 = controllable_hgrant4 & ~n54186;
  assign n54188 = ~n43215 & ~n54187;
  assign n54189 = ~i_hbusreq5 & ~n54188;
  assign n54190 = ~n54182 & ~n54189;
  assign n54191 = ~controllable_hgrant5 & ~n54190;
  assign n54192 = ~n43170 & ~n54191;
  assign n54193 = ~controllable_hmaster2 & ~n54192;
  assign n54194 = ~n54153 & ~n54193;
  assign n54195 = ~controllable_hmaster1 & ~n54194;
  assign n54196 = ~n54152 & ~n54195;
  assign n54197 = ~i_hbusreq6 & ~n54196;
  assign n54198 = ~n54181 & ~n54197;
  assign n54199 = ~controllable_hgrant6 & ~n54198;
  assign n54200 = ~n43162 & ~n54199;
  assign n54201 = ~controllable_hmaster0 & ~n54200;
  assign n54202 = ~n54180 & ~n54201;
  assign n54203 = i_hlock8 & ~n54202;
  assign n54204 = i_hbusreq6 & ~n54057;
  assign n54205 = i_hbusreq5 & ~n54051;
  assign n54206 = ~i_hbusreq9 & ~n54159;
  assign n54207 = ~n40536 & ~n54206;
  assign n54208 = ~i_hbusreq4 & ~n54207;
  assign n54209 = ~n40535 & ~n54208;
  assign n54210 = controllable_hgrant4 & ~n54209;
  assign n54211 = ~n43289 & ~n54210;
  assign n54212 = ~i_hbusreq5 & ~n54211;
  assign n54213 = ~n54205 & ~n54212;
  assign n54214 = ~controllable_hgrant5 & ~n54213;
  assign n54215 = ~n43246 & ~n54214;
  assign n54216 = ~controllable_hmaster2 & ~n54215;
  assign n54217 = ~n54153 & ~n54216;
  assign n54218 = ~controllable_hmaster1 & ~n54217;
  assign n54219 = ~n54152 & ~n54218;
  assign n54220 = ~i_hbusreq6 & ~n54219;
  assign n54221 = ~n54204 & ~n54220;
  assign n54222 = ~controllable_hgrant6 & ~n54221;
  assign n54223 = ~n43238 & ~n54222;
  assign n54224 = ~controllable_hmaster0 & ~n54223;
  assign n54225 = ~n54180 & ~n54224;
  assign n54226 = ~i_hlock8 & ~n54225;
  assign n54227 = ~n54203 & ~n54226;
  assign n54228 = ~i_hbusreq8 & ~n54227;
  assign n54229 = ~n54137 & ~n54228;
  assign n54230 = controllable_hmaster3 & ~n54229;
  assign n54231 = i_hbusreq8 & ~n54121;
  assign n54232 = i_hbusreq6 & ~n54084;
  assign n54233 = controllable_hmaster2 & ~n54192;
  assign n54234 = i_hbusreq5 & ~n54066;
  assign n54235 = ~n8426 & ~n18338;
  assign n54236 = ~n43330 & ~n54235;
  assign n54237 = ~i_hbusreq9 & ~n54236;
  assign n54238 = ~n48366 & ~n54237;
  assign n54239 = ~i_hbusreq4 & ~n54238;
  assign n54240 = ~n48365 & ~n54239;
  assign n54241 = controllable_hgrant4 & ~n54240;
  assign n54242 = ~n43365 & ~n54241;
  assign n54243 = ~i_hbusreq5 & ~n54242;
  assign n54244 = ~n54234 & ~n54243;
  assign n54245 = ~controllable_hgrant5 & ~n54244;
  assign n54246 = ~n43326 & ~n54245;
  assign n54247 = ~controllable_hmaster2 & ~n54246;
  assign n54248 = ~n54233 & ~n54247;
  assign n54249 = controllable_hmaster1 & ~n54248;
  assign n54250 = i_hbusreq5 & ~n54074;
  assign n54251 = i_hlock5 & ~n54188;
  assign n54252 = ~i_hlock5 & ~n54211;
  assign n54253 = ~n54251 & ~n54252;
  assign n54254 = ~i_hbusreq5 & ~n54253;
  assign n54255 = ~n54250 & ~n54254;
  assign n54256 = ~controllable_hgrant5 & ~n54255;
  assign n54257 = ~n43386 & ~n54256;
  assign n54258 = controllable_hmaster2 & ~n54257;
  assign n54259 = i_hbusreq5 & ~n54078;
  assign n54260 = ~n8426 & ~n18376;
  assign n54261 = ~n43406 & ~n54260;
  assign n54262 = ~i_hbusreq9 & ~n54261;
  assign n54263 = ~n48442 & ~n54262;
  assign n54264 = ~i_hbusreq4 & ~n54263;
  assign n54265 = ~n48441 & ~n54264;
  assign n54266 = controllable_hgrant4 & ~n54265;
  assign n54267 = ~n43453 & ~n54266;
  assign n54268 = ~i_hbusreq5 & ~n54267;
  assign n54269 = ~n54259 & ~n54268;
  assign n54270 = ~controllable_hgrant5 & ~n54269;
  assign n54271 = ~n43402 & ~n54270;
  assign n54272 = ~controllable_hmaster2 & ~n54271;
  assign n54273 = ~n54258 & ~n54272;
  assign n54274 = ~controllable_hmaster1 & ~n54273;
  assign n54275 = ~n54249 & ~n54274;
  assign n54276 = ~i_hbusreq6 & ~n54275;
  assign n54277 = ~n54232 & ~n54276;
  assign n54278 = ~controllable_hgrant6 & ~n54277;
  assign n54279 = ~n43317 & ~n54278;
  assign n54280 = controllable_hmaster0 & ~n54279;
  assign n54281 = i_hbusreq6 & ~n54096;
  assign n54282 = ~n10188 & ~n43470;
  assign n54283 = n8217 & ~n54282;
  assign n54284 = ~n22892 & ~n43474;
  assign n54285 = ~n8217 & ~n54284;
  assign n54286 = ~n54283 & ~n54285;
  assign n54287 = i_hlock6 & ~n54286;
  assign n54288 = ~n10188 & ~n43480;
  assign n54289 = n8217 & ~n54288;
  assign n54290 = ~n22892 & ~n43484;
  assign n54291 = ~n8217 & ~n54290;
  assign n54292 = ~n54289 & ~n54291;
  assign n54293 = ~i_hlock6 & ~n54292;
  assign n54294 = ~n54287 & ~n54293;
  assign n54295 = ~i_hbusreq6 & ~n54294;
  assign n54296 = ~n54281 & ~n54295;
  assign n54297 = controllable_hgrant6 & ~n54296;
  assign n54298 = i_hbusreq6 & ~n54117;
  assign n54299 = i_hbusreq5 & ~n54098;
  assign n54300 = ~n8426 & ~n18410;
  assign n54301 = ~n43504 & ~n54300;
  assign n54302 = ~i_hbusreq9 & ~n54301;
  assign n54303 = ~n48539 & ~n54302;
  assign n54304 = ~i_hbusreq4 & ~n54303;
  assign n54305 = ~n48538 & ~n54304;
  assign n54306 = controllable_hgrant4 & ~n54305;
  assign n54307 = ~n43574 & ~n54306;
  assign n54308 = ~i_hbusreq5 & ~n54307;
  assign n54309 = ~n54299 & ~n54308;
  assign n54310 = ~controllable_hgrant5 & ~n54309;
  assign n54311 = ~n43500 & ~n54310;
  assign n54312 = ~controllable_hmaster2 & ~n54311;
  assign n54313 = ~n54233 & ~n54312;
  assign n54314 = controllable_hmaster1 & ~n54313;
  assign n54315 = i_hbusreq5 & ~n54104;
  assign n54316 = ~n8426 & ~n18477;
  assign n54317 = ~n43633 & ~n54316;
  assign n54318 = ~i_hbusreq9 & ~n54317;
  assign n54319 = ~n48658 & ~n54318;
  assign n54320 = ~i_hbusreq4 & ~n54319;
  assign n54321 = ~n48657 & ~n54320;
  assign n54322 = controllable_hgrant4 & ~n54321;
  assign n54323 = ~n43685 & ~n54322;
  assign n54324 = ~i_hbusreq5 & ~n54323;
  assign n54325 = ~n54315 & ~n54324;
  assign n54326 = ~controllable_hgrant5 & ~n54325;
  assign n54327 = ~n43629 & ~n54326;
  assign n54328 = ~controllable_hmaster2 & ~n54327;
  assign n54329 = ~n48648 & ~n54328;
  assign n54330 = ~controllable_hmaster1 & ~n54329;
  assign n54331 = ~n54314 & ~n54330;
  assign n54332 = i_hlock6 & ~n54331;
  assign n54333 = controllable_hmaster2 & ~n54215;
  assign n54334 = ~n54312 & ~n54333;
  assign n54335 = controllable_hmaster1 & ~n54334;
  assign n54336 = ~n54330 & ~n54335;
  assign n54337 = ~i_hlock6 & ~n54336;
  assign n54338 = ~n54332 & ~n54337;
  assign n54339 = ~i_hbusreq6 & ~n54338;
  assign n54340 = ~n54298 & ~n54339;
  assign n54341 = ~controllable_hgrant6 & ~n54340;
  assign n54342 = ~n54297 & ~n54341;
  assign n54343 = ~controllable_hmaster0 & ~n54342;
  assign n54344 = ~n54280 & ~n54343;
  assign n54345 = ~i_hbusreq8 & ~n54344;
  assign n54346 = ~n54231 & ~n54345;
  assign n54347 = ~controllable_hmaster3 & ~n54346;
  assign n54348 = ~n54230 & ~n54347;
  assign n54349 = i_hlock7 & ~n54348;
  assign n54350 = i_hbusreq8 & ~n54131;
  assign n54351 = i_hbusreq6 & ~n54127;
  assign n54352 = ~n54247 & ~n54333;
  assign n54353 = controllable_hmaster1 & ~n54352;
  assign n54354 = ~n54274 & ~n54353;
  assign n54355 = ~i_hbusreq6 & ~n54354;
  assign n54356 = ~n54351 & ~n54355;
  assign n54357 = ~controllable_hgrant6 & ~n54356;
  assign n54358 = ~n43720 & ~n54357;
  assign n54359 = controllable_hmaster0 & ~n54358;
  assign n54360 = ~n54343 & ~n54359;
  assign n54361 = ~i_hbusreq8 & ~n54360;
  assign n54362 = ~n54350 & ~n54361;
  assign n54363 = ~controllable_hmaster3 & ~n54362;
  assign n54364 = ~n54230 & ~n54363;
  assign n54365 = ~i_hlock7 & ~n54364;
  assign n54366 = ~n54349 & ~n54365;
  assign n54367 = ~i_hbusreq7 & ~n54366;
  assign n54368 = ~n54136 & ~n54367;
  assign n54369 = ~n7924 & ~n54368;
  assign n54370 = ~n43772 & ~n48777;
  assign n54371 = ~controllable_hgrant5 & ~n54370;
  assign n54372 = ~n43746 & ~n54371;
  assign n54373 = controllable_hmaster1 & ~n54372;
  assign n54374 = controllable_hmaster2 & ~n54372;
  assign n54375 = ~n45108 & ~n46030;
  assign n54376 = ~controllable_hgrant5 & ~n54375;
  assign n54377 = ~n45100 & ~n54376;
  assign n54378 = ~controllable_hmaster2 & ~n54377;
  assign n54379 = ~n54374 & ~n54378;
  assign n54380 = ~controllable_hmaster1 & ~n54379;
  assign n54381 = ~n54373 & ~n54380;
  assign n54382 = ~controllable_hgrant6 & ~n54381;
  assign n54383 = ~n45097 & ~n54382;
  assign n54384 = controllable_hmaster0 & ~n54383;
  assign n54385 = ~n43857 & ~n47532;
  assign n54386 = ~controllable_hgrant5 & ~n54385;
  assign n54387 = ~n43836 & ~n54386;
  assign n54388 = ~controllable_hmaster2 & ~n54387;
  assign n54389 = ~n54374 & ~n54388;
  assign n54390 = ~controllable_hmaster1 & ~n54389;
  assign n54391 = ~n54373 & ~n54390;
  assign n54392 = ~controllable_hgrant6 & ~n54391;
  assign n54393 = ~n43833 & ~n54392;
  assign n54394 = ~controllable_hmaster0 & ~n54393;
  assign n54395 = ~n54384 & ~n54394;
  assign n54396 = i_hlock8 & ~n54395;
  assign n54397 = ~n43890 & ~n47565;
  assign n54398 = ~controllable_hgrant5 & ~n54397;
  assign n54399 = ~n43875 & ~n54398;
  assign n54400 = ~controllable_hmaster2 & ~n54399;
  assign n54401 = ~n54374 & ~n54400;
  assign n54402 = ~controllable_hmaster1 & ~n54401;
  assign n54403 = ~n54373 & ~n54402;
  assign n54404 = ~controllable_hgrant6 & ~n54403;
  assign n54405 = ~n43872 & ~n54404;
  assign n54406 = ~controllable_hmaster0 & ~n54405;
  assign n54407 = ~n54384 & ~n54406;
  assign n54408 = ~i_hlock8 & ~n54407;
  assign n54409 = ~n54396 & ~n54408;
  assign n54410 = controllable_hmaster3 & ~n54409;
  assign n54411 = controllable_hmaster2 & ~n54387;
  assign n54412 = ~n43933 & ~n48851;
  assign n54413 = ~controllable_hgrant5 & ~n54412;
  assign n54414 = ~n43913 & ~n54413;
  assign n54415 = ~controllable_hmaster2 & ~n54414;
  assign n54416 = ~n54411 & ~n54415;
  assign n54417 = controllable_hmaster1 & ~n54416;
  assign n54418 = i_hlock5 & ~n54385;
  assign n54419 = ~i_hlock5 & ~n54397;
  assign n54420 = ~n54418 & ~n54419;
  assign n54421 = ~controllable_hgrant5 & ~n54420;
  assign n54422 = ~n43949 & ~n54421;
  assign n54423 = controllable_hmaster2 & ~n54422;
  assign n54424 = ~n43985 & ~n48901;
  assign n54425 = ~controllable_hgrant5 & ~n54424;
  assign n54426 = ~n43959 & ~n54425;
  assign n54427 = ~controllable_hmaster2 & ~n54426;
  assign n54428 = ~n54423 & ~n54427;
  assign n54429 = ~controllable_hmaster1 & ~n54428;
  assign n54430 = ~n54417 & ~n54429;
  assign n54431 = ~controllable_hgrant6 & ~n54430;
  assign n54432 = ~n43908 & ~n54431;
  assign n54433 = controllable_hmaster0 & ~n54432;
  assign n54434 = ~n22929 & ~n44001;
  assign n54435 = ~n8217 & ~n54434;
  assign n54436 = ~n43999 & ~n54435;
  assign n54437 = i_hlock6 & ~n54436;
  assign n54438 = ~n22929 & ~n44011;
  assign n54439 = ~n8217 & ~n54438;
  assign n54440 = ~n44009 & ~n54439;
  assign n54441 = ~i_hlock6 & ~n54440;
  assign n54442 = ~n54437 & ~n54441;
  assign n54443 = controllable_hgrant6 & ~n54442;
  assign n54444 = ~n44047 & ~n48951;
  assign n54445 = ~controllable_hgrant5 & ~n54444;
  assign n54446 = ~n44021 & ~n54445;
  assign n54447 = ~controllable_hmaster2 & ~n54446;
  assign n54448 = ~n54411 & ~n54447;
  assign n54449 = controllable_hmaster1 & ~n54448;
  assign n54450 = ~n8378 & ~n22924;
  assign n54451 = ~n44054 & ~n54450;
  assign n54452 = controllable_hgrant5 & ~n54451;
  assign n54453 = i_hlock4 & ~n43805;
  assign n54454 = ~i_hlock4 & ~n43817;
  assign n54455 = ~n54453 & ~n54454;
  assign n54456 = ~controllable_hgrant4 & ~n54455;
  assign n54457 = ~n49009 & ~n54456;
  assign n54458 = ~controllable_hgrant5 & ~n54457;
  assign n54459 = ~n54452 & ~n54458;
  assign n54460 = controllable_hmaster2 & ~n54459;
  assign n54461 = ~n44097 & ~n49033;
  assign n54462 = ~controllable_hgrant5 & ~n54461;
  assign n54463 = ~n44079 & ~n54462;
  assign n54464 = ~controllable_hmaster2 & ~n54463;
  assign n54465 = ~n54460 & ~n54464;
  assign n54466 = ~controllable_hmaster1 & ~n54465;
  assign n54467 = ~n54449 & ~n54466;
  assign n54468 = i_hlock6 & ~n54467;
  assign n54469 = controllable_hmaster2 & ~n54399;
  assign n54470 = ~n54447 & ~n54469;
  assign n54471 = controllable_hmaster1 & ~n54470;
  assign n54472 = ~n54466 & ~n54471;
  assign n54473 = ~i_hlock6 & ~n54472;
  assign n54474 = ~n54468 & ~n54473;
  assign n54475 = ~controllable_hgrant6 & ~n54474;
  assign n54476 = ~n54443 & ~n54475;
  assign n54477 = ~controllable_hmaster0 & ~n54476;
  assign n54478 = ~n54433 & ~n54477;
  assign n54479 = ~controllable_hmaster3 & ~n54478;
  assign n54480 = ~n54410 & ~n54479;
  assign n54481 = i_hlock7 & ~n54480;
  assign n54482 = ~n54415 & ~n54469;
  assign n54483 = controllable_hmaster1 & ~n54482;
  assign n54484 = ~n54429 & ~n54483;
  assign n54485 = ~controllable_hgrant6 & ~n54484;
  assign n54486 = ~n44122 & ~n54485;
  assign n54487 = controllable_hmaster0 & ~n54486;
  assign n54488 = ~n54477 & ~n54487;
  assign n54489 = ~controllable_hmaster3 & ~n54488;
  assign n54490 = ~n54410 & ~n54489;
  assign n54491 = ~i_hlock7 & ~n54490;
  assign n54492 = ~n54481 & ~n54491;
  assign n54493 = i_hbusreq7 & ~n54492;
  assign n54494 = i_hbusreq8 & ~n54409;
  assign n54495 = i_hbusreq6 & ~n54381;
  assign n54496 = i_hbusreq5 & ~n54370;
  assign n54497 = n8426 & ~n13998;
  assign n54498 = ~n8426 & ~n18745;
  assign n54499 = ~n54497 & ~n54498;
  assign n54500 = ~i_hbusreq9 & ~n54499;
  assign n54501 = ~n49115 & ~n54500;
  assign n54502 = i_hlock4 & ~n54501;
  assign n54503 = ~n8426 & ~n18763;
  assign n54504 = ~n54497 & ~n54503;
  assign n54505 = ~i_hbusreq9 & ~n54504;
  assign n54506 = ~n49122 & ~n54505;
  assign n54507 = ~i_hlock4 & ~n54506;
  assign n54508 = ~n54502 & ~n54507;
  assign n54509 = ~i_hbusreq4 & ~n54508;
  assign n54510 = ~n49114 & ~n54509;
  assign n54511 = controllable_hgrant4 & ~n54510;
  assign n54512 = ~n44217 & ~n54511;
  assign n54513 = ~i_hbusreq5 & ~n54512;
  assign n54514 = ~n54496 & ~n54513;
  assign n54515 = ~controllable_hgrant5 & ~n54514;
  assign n54516 = ~n44150 & ~n54515;
  assign n54517 = controllable_hmaster1 & ~n54516;
  assign n54518 = controllable_hmaster2 & ~n54516;
  assign n54519 = i_hbusreq5 & ~n54375;
  assign n54520 = n8426 & ~n14032;
  assign n54521 = ~n8426 & ~n18811;
  assign n54522 = ~n54520 & ~n54521;
  assign n54523 = i_hlock9 & ~n54522;
  assign n54524 = n8426 & ~n14067;
  assign n54525 = ~n8426 & ~n18863;
  assign n54526 = ~n54524 & ~n54525;
  assign n54527 = ~i_hlock9 & ~n54526;
  assign n54528 = ~n54523 & ~n54527;
  assign n54529 = ~i_hbusreq9 & ~n54528;
  assign n54530 = ~n46636 & ~n54529;
  assign n54531 = i_hlock4 & ~n54530;
  assign n54532 = ~n8426 & ~n18825;
  assign n54533 = ~n54520 & ~n54532;
  assign n54534 = i_hlock9 & ~n54533;
  assign n54535 = ~n8426 & ~n18875;
  assign n54536 = ~n54524 & ~n54535;
  assign n54537 = ~i_hlock9 & ~n54536;
  assign n54538 = ~n54534 & ~n54537;
  assign n54539 = ~i_hbusreq9 & ~n54538;
  assign n54540 = ~n46647 & ~n54539;
  assign n54541 = ~i_hlock4 & ~n54540;
  assign n54542 = ~n54531 & ~n54541;
  assign n54543 = ~i_hbusreq4 & ~n54542;
  assign n54544 = ~n46635 & ~n54543;
  assign n54545 = controllable_hgrant4 & ~n54544;
  assign n54546 = ~n45203 & ~n54545;
  assign n54547 = ~i_hbusreq5 & ~n54546;
  assign n54548 = ~n54519 & ~n54547;
  assign n54549 = ~controllable_hgrant5 & ~n54548;
  assign n54550 = ~n45182 & ~n54549;
  assign n54551 = ~controllable_hmaster2 & ~n54550;
  assign n54552 = ~n54518 & ~n54551;
  assign n54553 = ~controllable_hmaster1 & ~n54552;
  assign n54554 = ~n54517 & ~n54553;
  assign n54555 = ~i_hbusreq6 & ~n54554;
  assign n54556 = ~n54495 & ~n54555;
  assign n54557 = ~controllable_hgrant6 & ~n54556;
  assign n54558 = ~n45174 & ~n54557;
  assign n54559 = controllable_hmaster0 & ~n54558;
  assign n54560 = i_hbusreq6 & ~n54391;
  assign n54561 = i_hbusreq5 & ~n54385;
  assign n54562 = ~i_hbusreq9 & ~n54522;
  assign n54563 = ~n47680 & ~n54562;
  assign n54564 = i_hlock4 & ~n54563;
  assign n54565 = ~i_hbusreq9 & ~n54533;
  assign n54566 = ~n47684 & ~n54565;
  assign n54567 = ~i_hlock4 & ~n54566;
  assign n54568 = ~n54564 & ~n54567;
  assign n54569 = ~i_hbusreq4 & ~n54568;
  assign n54570 = ~n47679 & ~n54569;
  assign n54571 = controllable_hgrant4 & ~n54570;
  assign n54572 = ~n44425 & ~n54571;
  assign n54573 = ~i_hbusreq5 & ~n54572;
  assign n54574 = ~n54561 & ~n54573;
  assign n54575 = ~controllable_hgrant5 & ~n54574;
  assign n54576 = ~n44376 & ~n54575;
  assign n54577 = ~controllable_hmaster2 & ~n54576;
  assign n54578 = ~n54518 & ~n54577;
  assign n54579 = ~controllable_hmaster1 & ~n54578;
  assign n54580 = ~n54517 & ~n54579;
  assign n54581 = ~i_hbusreq6 & ~n54580;
  assign n54582 = ~n54560 & ~n54581;
  assign n54583 = ~controllable_hgrant6 & ~n54582;
  assign n54584 = ~n44368 & ~n54583;
  assign n54585 = ~controllable_hmaster0 & ~n54584;
  assign n54586 = ~n54559 & ~n54585;
  assign n54587 = i_hlock8 & ~n54586;
  assign n54588 = i_hbusreq6 & ~n54403;
  assign n54589 = i_hbusreq5 & ~n54397;
  assign n54590 = ~i_hbusreq9 & ~n54526;
  assign n54591 = ~n47740 & ~n54590;
  assign n54592 = i_hlock4 & ~n54591;
  assign n54593 = ~i_hbusreq9 & ~n54536;
  assign n54594 = ~n47744 & ~n54593;
  assign n54595 = ~i_hlock4 & ~n54594;
  assign n54596 = ~n54592 & ~n54595;
  assign n54597 = ~i_hbusreq4 & ~n54596;
  assign n54598 = ~n47739 & ~n54597;
  assign n54599 = controllable_hgrant4 & ~n54598;
  assign n54600 = ~n44499 & ~n54599;
  assign n54601 = ~i_hbusreq5 & ~n54600;
  assign n54602 = ~n54589 & ~n54601;
  assign n54603 = ~controllable_hgrant5 & ~n54602;
  assign n54604 = ~n44456 & ~n54603;
  assign n54605 = ~controllable_hmaster2 & ~n54604;
  assign n54606 = ~n54518 & ~n54605;
  assign n54607 = ~controllable_hmaster1 & ~n54606;
  assign n54608 = ~n54517 & ~n54607;
  assign n54609 = ~i_hbusreq6 & ~n54608;
  assign n54610 = ~n54588 & ~n54609;
  assign n54611 = ~controllable_hgrant6 & ~n54610;
  assign n54612 = ~n44448 & ~n54611;
  assign n54613 = ~controllable_hmaster0 & ~n54612;
  assign n54614 = ~n54559 & ~n54613;
  assign n54615 = ~i_hlock8 & ~n54614;
  assign n54616 = ~n54587 & ~n54615;
  assign n54617 = ~i_hbusreq8 & ~n54616;
  assign n54618 = ~n54494 & ~n54617;
  assign n54619 = controllable_hmaster3 & ~n54618;
  assign n54620 = i_hbusreq8 & ~n54478;
  assign n54621 = i_hbusreq6 & ~n54430;
  assign n54622 = controllable_hmaster2 & ~n54576;
  assign n54623 = i_hbusreq5 & ~n54412;
  assign n54624 = n8426 & ~n14110;
  assign n54625 = ~n8426 & ~n18916;
  assign n54626 = ~n54624 & ~n54625;
  assign n54627 = ~i_hbusreq9 & ~n54626;
  assign n54628 = ~n49503 & ~n54627;
  assign n54629 = i_hlock4 & ~n54628;
  assign n54630 = ~n8426 & ~n18925;
  assign n54631 = ~n54624 & ~n54630;
  assign n54632 = ~i_hbusreq9 & ~n54631;
  assign n54633 = ~n49510 & ~n54632;
  assign n54634 = ~i_hlock4 & ~n54633;
  assign n54635 = ~n54629 & ~n54634;
  assign n54636 = ~i_hbusreq4 & ~n54635;
  assign n54637 = ~n49502 & ~n54636;
  assign n54638 = controllable_hgrant4 & ~n54637;
  assign n54639 = ~n44575 & ~n54638;
  assign n54640 = ~i_hbusreq5 & ~n54639;
  assign n54641 = ~n54623 & ~n54640;
  assign n54642 = ~controllable_hgrant5 & ~n54641;
  assign n54643 = ~n44536 & ~n54642;
  assign n54644 = ~controllable_hmaster2 & ~n54643;
  assign n54645 = ~n54622 & ~n54644;
  assign n54646 = controllable_hmaster1 & ~n54645;
  assign n54647 = i_hbusreq5 & ~n54420;
  assign n54648 = i_hlock5 & ~n54572;
  assign n54649 = ~i_hlock5 & ~n54600;
  assign n54650 = ~n54648 & ~n54649;
  assign n54651 = ~i_hbusreq5 & ~n54650;
  assign n54652 = ~n54647 & ~n54651;
  assign n54653 = ~controllable_hgrant5 & ~n54652;
  assign n54654 = ~n44596 & ~n54653;
  assign n54655 = controllable_hmaster2 & ~n54654;
  assign n54656 = i_hbusreq5 & ~n54424;
  assign n54657 = n8426 & ~n14153;
  assign n54658 = ~n8426 & ~n18965;
  assign n54659 = ~n54657 & ~n54658;
  assign n54660 = ~i_hbusreq9 & ~n54659;
  assign n54661 = ~n49592 & ~n54660;
  assign n54662 = i_hlock4 & ~n54661;
  assign n54663 = ~n8426 & ~n18979;
  assign n54664 = ~n54657 & ~n54663;
  assign n54665 = ~i_hbusreq9 & ~n54664;
  assign n54666 = ~n49599 & ~n54665;
  assign n54667 = ~i_hlock4 & ~n54666;
  assign n54668 = ~n54662 & ~n54667;
  assign n54669 = ~i_hbusreq4 & ~n54668;
  assign n54670 = ~n49591 & ~n54669;
  assign n54671 = controllable_hgrant4 & ~n54670;
  assign n54672 = ~n44663 & ~n54671;
  assign n54673 = ~i_hbusreq5 & ~n54672;
  assign n54674 = ~n54656 & ~n54673;
  assign n54675 = ~controllable_hgrant5 & ~n54674;
  assign n54676 = ~n44612 & ~n54675;
  assign n54677 = ~controllable_hmaster2 & ~n54676;
  assign n54678 = ~n54655 & ~n54677;
  assign n54679 = ~controllable_hmaster1 & ~n54678;
  assign n54680 = ~n54646 & ~n54679;
  assign n54681 = ~i_hbusreq6 & ~n54680;
  assign n54682 = ~n54621 & ~n54681;
  assign n54683 = ~controllable_hgrant6 & ~n54682;
  assign n54684 = ~n44527 & ~n54683;
  assign n54685 = controllable_hmaster0 & ~n54684;
  assign n54686 = i_hbusreq6 & ~n54442;
  assign n54687 = ~n15481 & ~n44680;
  assign n54688 = n8217 & ~n54687;
  assign n54689 = ~n22965 & ~n44684;
  assign n54690 = ~n8217 & ~n54689;
  assign n54691 = ~n54688 & ~n54690;
  assign n54692 = i_hlock6 & ~n54691;
  assign n54693 = ~n15481 & ~n44690;
  assign n54694 = n8217 & ~n54693;
  assign n54695 = ~n22965 & ~n44694;
  assign n54696 = ~n8217 & ~n54695;
  assign n54697 = ~n54694 & ~n54696;
  assign n54698 = ~i_hlock6 & ~n54697;
  assign n54699 = ~n54692 & ~n54698;
  assign n54700 = ~i_hbusreq6 & ~n54699;
  assign n54701 = ~n54686 & ~n54700;
  assign n54702 = controllable_hgrant6 & ~n54701;
  assign n54703 = i_hbusreq6 & ~n54474;
  assign n54704 = i_hbusreq5 & ~n54444;
  assign n54705 = n8426 & ~n14192;
  assign n54706 = ~n8426 & ~n19015;
  assign n54707 = ~n54705 & ~n54706;
  assign n54708 = ~i_hbusreq9 & ~n54707;
  assign n54709 = ~n49707 & ~n54708;
  assign n54710 = i_hlock4 & ~n54709;
  assign n54711 = ~n8426 & ~n19027;
  assign n54712 = ~n54705 & ~n54711;
  assign n54713 = ~i_hbusreq9 & ~n54712;
  assign n54714 = ~n49714 & ~n54713;
  assign n54715 = ~i_hlock4 & ~n54714;
  assign n54716 = ~n54710 & ~n54715;
  assign n54717 = ~i_hbusreq4 & ~n54716;
  assign n54718 = ~n49706 & ~n54717;
  assign n54719 = controllable_hgrant4 & ~n54718;
  assign n54720 = ~n44770 & ~n54719;
  assign n54721 = ~i_hbusreq5 & ~n54720;
  assign n54722 = ~n54704 & ~n54721;
  assign n54723 = ~controllable_hgrant5 & ~n54722;
  assign n54724 = ~n44710 & ~n54723;
  assign n54725 = ~controllable_hmaster2 & ~n54724;
  assign n54726 = ~n54622 & ~n54725;
  assign n54727 = controllable_hmaster1 & ~n54726;
  assign n54728 = i_hbusreq5 & ~n54451;
  assign n54729 = n8378 & ~n15474;
  assign n54730 = ~n8378 & ~n22958;
  assign n54731 = ~n54729 & ~n54730;
  assign n54732 = ~i_hbusreq5 & ~n54731;
  assign n54733 = ~n54728 & ~n54732;
  assign n54734 = controllable_hgrant5 & ~n54733;
  assign n54735 = i_hbusreq5 & ~n54457;
  assign n54736 = i_hbusreq4 & ~n54455;
  assign n54737 = i_hlock4 & ~n45244;
  assign n54738 = ~i_hlock4 & ~n45290;
  assign n54739 = ~n54737 & ~n54738;
  assign n54740 = ~i_hbusreq4 & ~n54739;
  assign n54741 = ~n54736 & ~n54740;
  assign n54742 = ~controllable_hgrant4 & ~n54741;
  assign n54743 = ~n49828 & ~n54742;
  assign n54744 = ~i_hbusreq5 & ~n54743;
  assign n54745 = ~n54735 & ~n54744;
  assign n54746 = ~controllable_hgrant5 & ~n54745;
  assign n54747 = ~n54734 & ~n54746;
  assign n54748 = controllable_hmaster2 & ~n54747;
  assign n54749 = i_hbusreq5 & ~n54461;
  assign n54750 = n8426 & ~n14264;
  assign n54751 = ~n8426 & ~n19096;
  assign n54752 = ~n54750 & ~n54751;
  assign n54753 = ~i_hbusreq9 & ~n54752;
  assign n54754 = ~n49856 & ~n54753;
  assign n54755 = i_hlock4 & ~n54754;
  assign n54756 = ~n8426 & ~n19116;
  assign n54757 = ~n54750 & ~n54756;
  assign n54758 = ~i_hbusreq9 & ~n54757;
  assign n54759 = ~n49863 & ~n54758;
  assign n54760 = ~i_hlock4 & ~n54759;
  assign n54761 = ~n54755 & ~n54760;
  assign n54762 = ~i_hbusreq4 & ~n54761;
  assign n54763 = ~n49855 & ~n54762;
  assign n54764 = controllable_hgrant4 & ~n54763;
  assign n54765 = ~n44885 & ~n54764;
  assign n54766 = ~i_hbusreq5 & ~n54765;
  assign n54767 = ~n54749 & ~n54766;
  assign n54768 = ~controllable_hgrant5 & ~n54767;
  assign n54769 = ~n44825 & ~n54768;
  assign n54770 = ~controllable_hmaster2 & ~n54769;
  assign n54771 = ~n54748 & ~n54770;
  assign n54772 = ~controllable_hmaster1 & ~n54771;
  assign n54773 = ~n54727 & ~n54772;
  assign n54774 = i_hlock6 & ~n54773;
  assign n54775 = controllable_hmaster2 & ~n54604;
  assign n54776 = ~n54725 & ~n54775;
  assign n54777 = controllable_hmaster1 & ~n54776;
  assign n54778 = ~n54772 & ~n54777;
  assign n54779 = ~i_hlock6 & ~n54778;
  assign n54780 = ~n54774 & ~n54779;
  assign n54781 = ~i_hbusreq6 & ~n54780;
  assign n54782 = ~n54703 & ~n54781;
  assign n54783 = ~controllable_hgrant6 & ~n54782;
  assign n54784 = ~n54702 & ~n54783;
  assign n54785 = ~controllable_hmaster0 & ~n54784;
  assign n54786 = ~n54685 & ~n54785;
  assign n54787 = ~i_hbusreq8 & ~n54786;
  assign n54788 = ~n54620 & ~n54787;
  assign n54789 = ~controllable_hmaster3 & ~n54788;
  assign n54790 = ~n54619 & ~n54789;
  assign n54791 = i_hlock7 & ~n54790;
  assign n54792 = i_hbusreq8 & ~n54488;
  assign n54793 = i_hbusreq6 & ~n54484;
  assign n54794 = ~n54644 & ~n54775;
  assign n54795 = controllable_hmaster1 & ~n54794;
  assign n54796 = ~n54679 & ~n54795;
  assign n54797 = ~i_hbusreq6 & ~n54796;
  assign n54798 = ~n54793 & ~n54797;
  assign n54799 = ~controllable_hgrant6 & ~n54798;
  assign n54800 = ~n44920 & ~n54799;
  assign n54801 = controllable_hmaster0 & ~n54800;
  assign n54802 = ~n54785 & ~n54801;
  assign n54803 = ~i_hbusreq8 & ~n54802;
  assign n54804 = ~n54792 & ~n54803;
  assign n54805 = ~controllable_hmaster3 & ~n54804;
  assign n54806 = ~n54619 & ~n54805;
  assign n54807 = ~i_hlock7 & ~n54806;
  assign n54808 = ~n54791 & ~n54807;
  assign n54809 = ~i_hbusreq7 & ~n54808;
  assign n54810 = ~n54493 & ~n54809;
  assign n54811 = n7924 & ~n54810;
  assign n54812 = ~n54369 & ~n54811;
  assign n54813 = n8214 & ~n54812;
  assign n54814 = ~n54023 & ~n54813;
  assign n54815 = ~n8202 & ~n54814;
  assign n54816 = ~n42732 & ~n48014;
  assign n54817 = ~controllable_hgrant4 & ~n54816;
  assign n54818 = ~n42713 & ~n54817;
  assign n54819 = ~controllable_hgrant5 & ~n54818;
  assign n54820 = ~n42709 & ~n54819;
  assign n54821 = controllable_hmaster1 & ~n54820;
  assign n54822 = controllable_hmaster2 & ~n54820;
  assign n54823 = ~n40210 & ~n42766;
  assign n54824 = i_hlock9 & ~n54823;
  assign n54825 = ~n40240 & ~n42799;
  assign n54826 = ~i_hlock9 & ~n54825;
  assign n54827 = ~n54824 & ~n54826;
  assign n54828 = ~controllable_hgrant4 & ~n54827;
  assign n54829 = ~n44951 & ~n54828;
  assign n54830 = ~controllable_hgrant5 & ~n54829;
  assign n54831 = ~n44947 & ~n54830;
  assign n54832 = ~controllable_hmaster2 & ~n54831;
  assign n54833 = ~n54822 & ~n54832;
  assign n54834 = ~controllable_hmaster1 & ~n54833;
  assign n54835 = ~n54821 & ~n54834;
  assign n54836 = ~controllable_hgrant6 & ~n54835;
  assign n54837 = ~n44944 & ~n54836;
  assign n54838 = controllable_hmaster0 & ~n54837;
  assign n54839 = ~controllable_hgrant4 & ~n54823;
  assign n54840 = ~n42754 & ~n54839;
  assign n54841 = ~controllable_hgrant5 & ~n54840;
  assign n54842 = ~n42751 & ~n54841;
  assign n54843 = ~controllable_hmaster2 & ~n54842;
  assign n54844 = ~n54822 & ~n54843;
  assign n54845 = ~controllable_hmaster1 & ~n54844;
  assign n54846 = ~n54821 & ~n54845;
  assign n54847 = ~controllable_hgrant6 & ~n54846;
  assign n54848 = ~n42748 & ~n54847;
  assign n54849 = ~controllable_hmaster0 & ~n54848;
  assign n54850 = ~n54838 & ~n54849;
  assign n54851 = i_hlock8 & ~n54850;
  assign n54852 = ~controllable_hgrant4 & ~n54825;
  assign n54853 = ~n42789 & ~n54852;
  assign n54854 = ~controllable_hgrant5 & ~n54853;
  assign n54855 = ~n42786 & ~n54854;
  assign n54856 = ~controllable_hmaster2 & ~n54855;
  assign n54857 = ~n54822 & ~n54856;
  assign n54858 = ~controllable_hmaster1 & ~n54857;
  assign n54859 = ~n54821 & ~n54858;
  assign n54860 = ~controllable_hgrant6 & ~n54859;
  assign n54861 = ~n42783 & ~n54860;
  assign n54862 = ~controllable_hmaster0 & ~n54861;
  assign n54863 = ~n54838 & ~n54862;
  assign n54864 = ~i_hlock8 & ~n54863;
  assign n54865 = ~n54851 & ~n54864;
  assign n54866 = controllable_hmaster3 & ~n54865;
  assign n54867 = ~n8217 & ~n22999;
  assign n54868 = ~n42816 & ~n54867;
  assign n54869 = controllable_hgrant6 & ~n54868;
  assign n54870 = controllable_hmaster2 & ~n54842;
  assign n54871 = ~n48081 & ~n54870;
  assign n54872 = controllable_hmaster1 & ~n54871;
  assign n54873 = i_hlock5 & ~n54840;
  assign n54874 = ~i_hlock5 & ~n54853;
  assign n54875 = ~n54873 & ~n54874;
  assign n54876 = ~controllable_hgrant5 & ~n54875;
  assign n54877 = ~n42860 & ~n54876;
  assign n54878 = controllable_hmaster2 & ~n54877;
  assign n54879 = ~n42894 & ~n48106;
  assign n54880 = ~controllable_hgrant4 & ~n54879;
  assign n54881 = ~n42874 & ~n54880;
  assign n54882 = ~controllable_hgrant5 & ~n54881;
  assign n54883 = ~n42870 & ~n54882;
  assign n54884 = ~controllable_hmaster2 & ~n54883;
  assign n54885 = ~n54878 & ~n54884;
  assign n54886 = ~controllable_hmaster1 & ~n54885;
  assign n54887 = ~n54872 & ~n54886;
  assign n54888 = ~controllable_hgrant6 & ~n54887;
  assign n54889 = ~n54869 & ~n54888;
  assign n54890 = controllable_hmaster0 & ~n54889;
  assign n54891 = ~n42978 & ~n48141;
  assign n54892 = ~controllable_hgrant4 & ~n54891;
  assign n54893 = ~n42936 & ~n54892;
  assign n54894 = ~controllable_hgrant5 & ~n54893;
  assign n54895 = ~n42932 & ~n54894;
  assign n54896 = ~controllable_hmaster2 & ~n54895;
  assign n54897 = ~n54870 & ~n54896;
  assign n54898 = controllable_hmaster1 & ~n54897;
  assign n54899 = i_hlock4 & ~n54823;
  assign n54900 = ~i_hlock4 & ~n54825;
  assign n54901 = ~n54899 & ~n54900;
  assign n54902 = ~controllable_hgrant4 & ~n54901;
  assign n54903 = ~n43000 & ~n54902;
  assign n54904 = ~controllable_hgrant5 & ~n54903;
  assign n54905 = ~n42990 & ~n54904;
  assign n54906 = controllable_hmaster2 & ~n54905;
  assign n54907 = ~n43028 & ~n48194;
  assign n54908 = ~controllable_hgrant4 & ~n54907;
  assign n54909 = ~n43016 & ~n54908;
  assign n54910 = ~controllable_hgrant5 & ~n54909;
  assign n54911 = ~n43012 & ~n54910;
  assign n54912 = ~controllable_hmaster2 & ~n54911;
  assign n54913 = ~n54906 & ~n54912;
  assign n54914 = ~controllable_hmaster1 & ~n54913;
  assign n54915 = ~n54898 & ~n54914;
  assign n54916 = i_hlock6 & ~n54915;
  assign n54917 = controllable_hmaster2 & ~n54855;
  assign n54918 = ~n54896 & ~n54917;
  assign n54919 = controllable_hmaster1 & ~n54918;
  assign n54920 = ~n54914 & ~n54919;
  assign n54921 = ~i_hlock6 & ~n54920;
  assign n54922 = ~n54916 & ~n54921;
  assign n54923 = ~controllable_hgrant6 & ~n54922;
  assign n54924 = ~n42928 & ~n54923;
  assign n54925 = ~controllable_hmaster0 & ~n54924;
  assign n54926 = ~n54890 & ~n54925;
  assign n54927 = ~controllable_hmaster3 & ~n54926;
  assign n54928 = ~n54866 & ~n54927;
  assign n54929 = i_hlock7 & ~n54928;
  assign n54930 = ~n8217 & ~n23009;
  assign n54931 = ~n43052 & ~n54930;
  assign n54932 = controllable_hgrant6 & ~n54931;
  assign n54933 = ~n48081 & ~n54917;
  assign n54934 = controllable_hmaster1 & ~n54933;
  assign n54935 = ~n54886 & ~n54934;
  assign n54936 = ~controllable_hgrant6 & ~n54935;
  assign n54937 = ~n54932 & ~n54936;
  assign n54938 = controllable_hmaster0 & ~n54937;
  assign n54939 = ~n54925 & ~n54938;
  assign n54940 = ~controllable_hmaster3 & ~n54939;
  assign n54941 = ~n54866 & ~n54940;
  assign n54942 = ~i_hlock7 & ~n54941;
  assign n54943 = ~n54929 & ~n54942;
  assign n54944 = i_hbusreq7 & ~n54943;
  assign n54945 = i_hbusreq8 & ~n54865;
  assign n54946 = i_hbusreq6 & ~n54835;
  assign n54947 = i_hbusreq5 & ~n54818;
  assign n54948 = i_hbusreq4 & ~n54816;
  assign n54949 = i_hbusreq9 & ~n54816;
  assign n54950 = ~n8365 & ~n18232;
  assign n54951 = ~n43098 & ~n54950;
  assign n54952 = ~i_hbusreq3 & ~n54951;
  assign n54953 = ~n48264 & ~n54952;
  assign n54954 = controllable_hgrant3 & ~n54953;
  assign n54955 = ~n43134 & ~n54954;
  assign n54956 = ~i_hbusreq9 & ~n54955;
  assign n54957 = ~n54949 & ~n54956;
  assign n54958 = ~i_hbusreq4 & ~n54957;
  assign n54959 = ~n54948 & ~n54958;
  assign n54960 = ~controllable_hgrant4 & ~n54959;
  assign n54961 = ~n43094 & ~n54960;
  assign n54962 = ~i_hbusreq5 & ~n54961;
  assign n54963 = ~n54947 & ~n54962;
  assign n54964 = ~controllable_hgrant5 & ~n54963;
  assign n54965 = ~n43083 & ~n54964;
  assign n54966 = controllable_hmaster1 & ~n54965;
  assign n54967 = controllable_hmaster2 & ~n54965;
  assign n54968 = i_hbusreq5 & ~n54829;
  assign n54969 = i_hbusreq4 & ~n54827;
  assign n54970 = i_hbusreq9 & ~n54827;
  assign n54971 = ~n8365 & ~n18264;
  assign n54972 = ~n43185 & ~n54971;
  assign n54973 = ~i_hbusreq3 & ~n54972;
  assign n54974 = ~n40302 & ~n54973;
  assign n54975 = controllable_hgrant3 & ~n54974;
  assign n54976 = ~n43209 & ~n54975;
  assign n54977 = i_hlock9 & ~n54976;
  assign n54978 = ~n8365 & ~n18295;
  assign n54979 = ~n43261 & ~n54978;
  assign n54980 = ~i_hbusreq3 & ~n54979;
  assign n54981 = ~n40370 & ~n54980;
  assign n54982 = controllable_hgrant3 & ~n54981;
  assign n54983 = ~n43283 & ~n54982;
  assign n54984 = ~i_hlock9 & ~n54983;
  assign n54985 = ~n54977 & ~n54984;
  assign n54986 = ~i_hbusreq9 & ~n54985;
  assign n54987 = ~n54970 & ~n54986;
  assign n54988 = ~i_hbusreq4 & ~n54987;
  assign n54989 = ~n54969 & ~n54988;
  assign n54990 = ~controllable_hgrant4 & ~n54989;
  assign n54991 = ~n45022 & ~n54990;
  assign n54992 = ~i_hbusreq5 & ~n54991;
  assign n54993 = ~n54968 & ~n54992;
  assign n54994 = ~controllable_hgrant5 & ~n54993;
  assign n54995 = ~n45011 & ~n54994;
  assign n54996 = ~controllable_hmaster2 & ~n54995;
  assign n54997 = ~n54967 & ~n54996;
  assign n54998 = ~controllable_hmaster1 & ~n54997;
  assign n54999 = ~n54966 & ~n54998;
  assign n55000 = ~i_hbusreq6 & ~n54999;
  assign n55001 = ~n54946 & ~n55000;
  assign n55002 = ~controllable_hgrant6 & ~n55001;
  assign n55003 = ~n45003 & ~n55002;
  assign n55004 = controllable_hmaster0 & ~n55003;
  assign n55005 = i_hbusreq6 & ~n54846;
  assign n55006 = i_hbusreq5 & ~n54840;
  assign n55007 = i_hbusreq4 & ~n54823;
  assign n55008 = i_hbusreq9 & ~n54823;
  assign n55009 = ~i_hbusreq9 & ~n54976;
  assign n55010 = ~n55008 & ~n55009;
  assign n55011 = ~i_hbusreq4 & ~n55010;
  assign n55012 = ~n55007 & ~n55011;
  assign n55013 = ~controllable_hgrant4 & ~n55012;
  assign n55014 = ~n43181 & ~n55013;
  assign n55015 = ~i_hbusreq5 & ~n55014;
  assign n55016 = ~n55006 & ~n55015;
  assign n55017 = ~controllable_hgrant5 & ~n55016;
  assign n55018 = ~n43170 & ~n55017;
  assign n55019 = ~controllable_hmaster2 & ~n55018;
  assign n55020 = ~n54967 & ~n55019;
  assign n55021 = ~controllable_hmaster1 & ~n55020;
  assign n55022 = ~n54966 & ~n55021;
  assign n55023 = ~i_hbusreq6 & ~n55022;
  assign n55024 = ~n55005 & ~n55023;
  assign n55025 = ~controllable_hgrant6 & ~n55024;
  assign n55026 = ~n43162 & ~n55025;
  assign n55027 = ~controllable_hmaster0 & ~n55026;
  assign n55028 = ~n55004 & ~n55027;
  assign n55029 = i_hlock8 & ~n55028;
  assign n55030 = i_hbusreq6 & ~n54859;
  assign n55031 = i_hbusreq5 & ~n54853;
  assign n55032 = i_hbusreq4 & ~n54825;
  assign n55033 = i_hbusreq9 & ~n54825;
  assign n55034 = ~i_hbusreq9 & ~n54983;
  assign n55035 = ~n55033 & ~n55034;
  assign n55036 = ~i_hbusreq4 & ~n55035;
  assign n55037 = ~n55032 & ~n55036;
  assign n55038 = ~controllable_hgrant4 & ~n55037;
  assign n55039 = ~n43257 & ~n55038;
  assign n55040 = ~i_hbusreq5 & ~n55039;
  assign n55041 = ~n55031 & ~n55040;
  assign n55042 = ~controllable_hgrant5 & ~n55041;
  assign n55043 = ~n43246 & ~n55042;
  assign n55044 = ~controllable_hmaster2 & ~n55043;
  assign n55045 = ~n54967 & ~n55044;
  assign n55046 = ~controllable_hmaster1 & ~n55045;
  assign n55047 = ~n54966 & ~n55046;
  assign n55048 = ~i_hbusreq6 & ~n55047;
  assign n55049 = ~n55030 & ~n55048;
  assign n55050 = ~controllable_hgrant6 & ~n55049;
  assign n55051 = ~n43238 & ~n55050;
  assign n55052 = ~controllable_hmaster0 & ~n55051;
  assign n55053 = ~n55004 & ~n55052;
  assign n55054 = ~i_hlock8 & ~n55053;
  assign n55055 = ~n55029 & ~n55054;
  assign n55056 = ~i_hbusreq8 & ~n55055;
  assign n55057 = ~n54945 & ~n55056;
  assign n55058 = controllable_hmaster3 & ~n55057;
  assign n55059 = i_hbusreq8 & ~n54926;
  assign n55060 = i_hbusreq6 & ~n54868;
  assign n55061 = n8217 & ~n10217;
  assign n55062 = ~n8217 & ~n23023;
  assign n55063 = ~n55061 & ~n55062;
  assign n55064 = ~i_hbusreq6 & ~n55063;
  assign n55065 = ~n55060 & ~n55064;
  assign n55066 = controllable_hgrant6 & ~n55065;
  assign n55067 = i_hbusreq6 & ~n54887;
  assign n55068 = controllable_hmaster2 & ~n55018;
  assign n55069 = ~n48408 & ~n55068;
  assign n55070 = controllable_hmaster1 & ~n55069;
  assign n55071 = i_hbusreq5 & ~n54875;
  assign n55072 = i_hlock5 & ~n55014;
  assign n55073 = ~i_hlock5 & ~n55039;
  assign n55074 = ~n55072 & ~n55073;
  assign n55075 = ~i_hbusreq5 & ~n55074;
  assign n55076 = ~n55071 & ~n55075;
  assign n55077 = ~controllable_hgrant5 & ~n55076;
  assign n55078 = ~n43386 & ~n55077;
  assign n55079 = controllable_hmaster2 & ~n55078;
  assign n55080 = i_hbusreq5 & ~n54881;
  assign n55081 = i_hbusreq4 & ~n54879;
  assign n55082 = i_hbusreq9 & ~n54879;
  assign n55083 = ~n8365 & ~n18372;
  assign n55084 = ~n43417 & ~n55083;
  assign n55085 = ~i_hbusreq3 & ~n55084;
  assign n55086 = ~n48453 & ~n55085;
  assign n55087 = controllable_hgrant3 & ~n55086;
  assign n55088 = ~n43447 & ~n55087;
  assign n55089 = ~i_hbusreq9 & ~n55088;
  assign n55090 = ~n55082 & ~n55089;
  assign n55091 = ~i_hbusreq4 & ~n55090;
  assign n55092 = ~n55081 & ~n55091;
  assign n55093 = ~controllable_hgrant4 & ~n55092;
  assign n55094 = ~n43413 & ~n55093;
  assign n55095 = ~i_hbusreq5 & ~n55094;
  assign n55096 = ~n55080 & ~n55095;
  assign n55097 = ~controllable_hgrant5 & ~n55096;
  assign n55098 = ~n43402 & ~n55097;
  assign n55099 = ~controllable_hmaster2 & ~n55098;
  assign n55100 = ~n55079 & ~n55099;
  assign n55101 = ~controllable_hmaster1 & ~n55100;
  assign n55102 = ~n55070 & ~n55101;
  assign n55103 = ~i_hbusreq6 & ~n55102;
  assign n55104 = ~n55067 & ~n55103;
  assign n55105 = ~controllable_hgrant6 & ~n55104;
  assign n55106 = ~n55066 & ~n55105;
  assign n55107 = controllable_hmaster0 & ~n55106;
  assign n55108 = i_hbusreq6 & ~n54922;
  assign n55109 = i_hbusreq5 & ~n54893;
  assign n55110 = i_hbusreq4 & ~n54891;
  assign n55111 = i_hbusreq9 & ~n54891;
  assign n55112 = ~n8365 & ~n18406;
  assign n55113 = ~n43515 & ~n55112;
  assign n55114 = ~i_hbusreq3 & ~n55113;
  assign n55115 = ~n48550 & ~n55114;
  assign n55116 = controllable_hgrant3 & ~n55115;
  assign n55117 = ~n43568 & ~n55116;
  assign n55118 = ~i_hbusreq9 & ~n55117;
  assign n55119 = ~n55111 & ~n55118;
  assign n55120 = ~i_hbusreq4 & ~n55119;
  assign n55121 = ~n55110 & ~n55120;
  assign n55122 = ~controllable_hgrant4 & ~n55121;
  assign n55123 = ~n43511 & ~n55122;
  assign n55124 = ~i_hbusreq5 & ~n55123;
  assign n55125 = ~n55109 & ~n55124;
  assign n55126 = ~controllable_hgrant5 & ~n55125;
  assign n55127 = ~n43500 & ~n55126;
  assign n55128 = ~controllable_hmaster2 & ~n55127;
  assign n55129 = ~n55068 & ~n55128;
  assign n55130 = controllable_hmaster1 & ~n55129;
  assign n55131 = i_hbusreq5 & ~n54903;
  assign n55132 = i_hbusreq4 & ~n54901;
  assign n55133 = i_hlock4 & ~n55010;
  assign n55134 = ~i_hlock4 & ~n55035;
  assign n55135 = ~n55133 & ~n55134;
  assign n55136 = ~i_hbusreq4 & ~n55135;
  assign n55137 = ~n55132 & ~n55136;
  assign n55138 = ~controllable_hgrant4 & ~n55137;
  assign n55139 = ~n43609 & ~n55138;
  assign n55140 = ~i_hbusreq5 & ~n55139;
  assign n55141 = ~n55131 & ~n55140;
  assign n55142 = ~controllable_hgrant5 & ~n55141;
  assign n55143 = ~n43589 & ~n55142;
  assign n55144 = controllable_hmaster2 & ~n55143;
  assign n55145 = i_hbusreq5 & ~n54909;
  assign n55146 = i_hbusreq4 & ~n54907;
  assign n55147 = i_hbusreq9 & ~n54907;
  assign n55148 = ~n8365 & ~n18473;
  assign n55149 = ~n43644 & ~n55148;
  assign n55150 = ~i_hbusreq3 & ~n55149;
  assign n55151 = ~n48669 & ~n55150;
  assign n55152 = controllable_hgrant3 & ~n55151;
  assign n55153 = ~n43679 & ~n55152;
  assign n55154 = ~i_hbusreq9 & ~n55153;
  assign n55155 = ~n55147 & ~n55154;
  assign n55156 = ~i_hbusreq4 & ~n55155;
  assign n55157 = ~n55146 & ~n55156;
  assign n55158 = ~controllable_hgrant4 & ~n55157;
  assign n55159 = ~n43640 & ~n55158;
  assign n55160 = ~i_hbusreq5 & ~n55159;
  assign n55161 = ~n55145 & ~n55160;
  assign n55162 = ~controllable_hgrant5 & ~n55161;
  assign n55163 = ~n43629 & ~n55162;
  assign n55164 = ~controllable_hmaster2 & ~n55163;
  assign n55165 = ~n55144 & ~n55164;
  assign n55166 = ~controllable_hmaster1 & ~n55165;
  assign n55167 = ~n55130 & ~n55166;
  assign n55168 = i_hlock6 & ~n55167;
  assign n55169 = controllable_hmaster2 & ~n55043;
  assign n55170 = ~n55128 & ~n55169;
  assign n55171 = controllable_hmaster1 & ~n55170;
  assign n55172 = ~n55166 & ~n55171;
  assign n55173 = ~i_hlock6 & ~n55172;
  assign n55174 = ~n55168 & ~n55173;
  assign n55175 = ~i_hbusreq6 & ~n55174;
  assign n55176 = ~n55108 & ~n55175;
  assign n55177 = ~controllable_hgrant6 & ~n55176;
  assign n55178 = ~n43492 & ~n55177;
  assign n55179 = ~controllable_hmaster0 & ~n55178;
  assign n55180 = ~n55107 & ~n55179;
  assign n55181 = ~i_hbusreq8 & ~n55180;
  assign n55182 = ~n55059 & ~n55181;
  assign n55183 = ~controllable_hmaster3 & ~n55182;
  assign n55184 = ~n55058 & ~n55183;
  assign n55185 = i_hlock7 & ~n55184;
  assign n55186 = i_hbusreq8 & ~n54939;
  assign n55187 = i_hbusreq6 & ~n54931;
  assign n55188 = n8217 & ~n10229;
  assign n55189 = ~n8217 & ~n23039;
  assign n55190 = ~n55188 & ~n55189;
  assign n55191 = ~i_hbusreq6 & ~n55190;
  assign n55192 = ~n55187 & ~n55191;
  assign n55193 = controllable_hgrant6 & ~n55192;
  assign n55194 = i_hbusreq6 & ~n54935;
  assign n55195 = ~n48408 & ~n55169;
  assign n55196 = controllable_hmaster1 & ~n55195;
  assign n55197 = ~n55101 & ~n55196;
  assign n55198 = ~i_hbusreq6 & ~n55197;
  assign n55199 = ~n55194 & ~n55198;
  assign n55200 = ~controllable_hgrant6 & ~n55199;
  assign n55201 = ~n55193 & ~n55200;
  assign n55202 = controllable_hmaster0 & ~n55201;
  assign n55203 = ~n55179 & ~n55202;
  assign n55204 = ~i_hbusreq8 & ~n55203;
  assign n55205 = ~n55186 & ~n55204;
  assign n55206 = ~controllable_hmaster3 & ~n55205;
  assign n55207 = ~n55058 & ~n55206;
  assign n55208 = ~i_hlock7 & ~n55207;
  assign n55209 = ~n55185 & ~n55208;
  assign n55210 = ~i_hbusreq7 & ~n55209;
  assign n55211 = ~n54944 & ~n55210;
  assign n55212 = ~n7924 & ~n55211;
  assign n55213 = ~n43770 & ~n48785;
  assign n55214 = ~controllable_hgrant4 & ~n55213;
  assign n55215 = ~n43750 & ~n55214;
  assign n55216 = ~controllable_hgrant5 & ~n55215;
  assign n55217 = ~n43746 & ~n55216;
  assign n55218 = controllable_hmaster1 & ~n55217;
  assign n55219 = controllable_hmaster2 & ~n55217;
  assign n55220 = ~n43855 & ~n46038;
  assign n55221 = i_hlock9 & ~n55220;
  assign n55222 = ~n43888 & ~n46077;
  assign n55223 = ~i_hlock9 & ~n55222;
  assign n55224 = ~n55221 & ~n55223;
  assign n55225 = ~controllable_hgrant4 & ~n55224;
  assign n55226 = ~n45104 & ~n55225;
  assign n55227 = ~controllable_hgrant5 & ~n55226;
  assign n55228 = ~n45100 & ~n55227;
  assign n55229 = ~controllable_hmaster2 & ~n55228;
  assign n55230 = ~n55219 & ~n55229;
  assign n55231 = ~controllable_hmaster1 & ~n55230;
  assign n55232 = ~n55218 & ~n55231;
  assign n55233 = ~controllable_hgrant6 & ~n55232;
  assign n55234 = ~n45097 & ~n55233;
  assign n55235 = controllable_hmaster0 & ~n55234;
  assign n55236 = ~controllable_hgrant4 & ~n55220;
  assign n55237 = ~n43839 & ~n55236;
  assign n55238 = ~controllable_hgrant5 & ~n55237;
  assign n55239 = ~n43836 & ~n55238;
  assign n55240 = ~controllable_hmaster2 & ~n55239;
  assign n55241 = ~n55219 & ~n55240;
  assign n55242 = ~controllable_hmaster1 & ~n55241;
  assign n55243 = ~n55218 & ~n55242;
  assign n55244 = ~controllable_hgrant6 & ~n55243;
  assign n55245 = ~n43833 & ~n55244;
  assign n55246 = ~controllable_hmaster0 & ~n55245;
  assign n55247 = ~n55235 & ~n55246;
  assign n55248 = i_hlock8 & ~n55247;
  assign n55249 = ~controllable_hgrant4 & ~n55222;
  assign n55250 = ~n43878 & ~n55249;
  assign n55251 = ~controllable_hgrant5 & ~n55250;
  assign n55252 = ~n43875 & ~n55251;
  assign n55253 = ~controllable_hmaster2 & ~n55252;
  assign n55254 = ~n55219 & ~n55253;
  assign n55255 = ~controllable_hmaster1 & ~n55254;
  assign n55256 = ~n55218 & ~n55255;
  assign n55257 = ~controllable_hgrant6 & ~n55256;
  assign n55258 = ~n43872 & ~n55257;
  assign n55259 = ~controllable_hmaster0 & ~n55258;
  assign n55260 = ~n55235 & ~n55259;
  assign n55261 = ~i_hlock8 & ~n55260;
  assign n55262 = ~n55248 & ~n55261;
  assign n55263 = controllable_hmaster3 & ~n55262;
  assign n55264 = ~n8217 & ~n23067;
  assign n55265 = ~n43905 & ~n55264;
  assign n55266 = controllable_hgrant6 & ~n55265;
  assign n55267 = controllable_hmaster2 & ~n55239;
  assign n55268 = ~n8378 & ~n23061;
  assign n55269 = ~n43910 & ~n55268;
  assign n55270 = controllable_hgrant5 & ~n55269;
  assign n55271 = ~n8426 & ~n23059;
  assign n55272 = ~n43914 & ~n55271;
  assign n55273 = controllable_hgrant4 & ~n55272;
  assign n55274 = i_hlock3 & ~n43803;
  assign n55275 = ~i_hlock3 & ~n43815;
  assign n55276 = ~n55274 & ~n55275;
  assign n55277 = ~controllable_hgrant3 & ~n55276;
  assign n55278 = ~n48859 & ~n55277;
  assign n55279 = ~controllable_hgrant4 & ~n55278;
  assign n55280 = ~n55273 & ~n55279;
  assign n55281 = ~controllable_hgrant5 & ~n55280;
  assign n55282 = ~n55270 & ~n55281;
  assign n55283 = ~controllable_hmaster2 & ~n55282;
  assign n55284 = ~n55267 & ~n55283;
  assign n55285 = controllable_hmaster1 & ~n55284;
  assign n55286 = i_hlock5 & ~n55237;
  assign n55287 = ~i_hlock5 & ~n55250;
  assign n55288 = ~n55286 & ~n55287;
  assign n55289 = ~controllable_hgrant5 & ~n55288;
  assign n55290 = ~n43949 & ~n55289;
  assign n55291 = controllable_hmaster2 & ~n55290;
  assign n55292 = ~n43983 & ~n48909;
  assign n55293 = ~controllable_hgrant4 & ~n55292;
  assign n55294 = ~n43963 & ~n55293;
  assign n55295 = ~controllable_hgrant5 & ~n55294;
  assign n55296 = ~n43959 & ~n55295;
  assign n55297 = ~controllable_hmaster2 & ~n55296;
  assign n55298 = ~n55291 & ~n55297;
  assign n55299 = ~controllable_hmaster1 & ~n55298;
  assign n55300 = ~n55285 & ~n55299;
  assign n55301 = ~controllable_hgrant6 & ~n55300;
  assign n55302 = ~n55266 & ~n55301;
  assign n55303 = controllable_hmaster0 & ~n55302;
  assign n55304 = ~n44045 & ~n48959;
  assign n55305 = ~controllable_hgrant4 & ~n55304;
  assign n55306 = ~n44025 & ~n55305;
  assign n55307 = ~controllable_hgrant5 & ~n55306;
  assign n55308 = ~n44021 & ~n55307;
  assign n55309 = ~controllable_hmaster2 & ~n55308;
  assign n55310 = ~n55267 & ~n55309;
  assign n55311 = controllable_hmaster1 & ~n55310;
  assign n55312 = i_hlock4 & ~n55220;
  assign n55313 = ~i_hlock4 & ~n55222;
  assign n55314 = ~n55312 & ~n55313;
  assign n55315 = ~controllable_hgrant4 & ~n55314;
  assign n55316 = ~n44067 & ~n55315;
  assign n55317 = ~controllable_hgrant5 & ~n55316;
  assign n55318 = ~n44057 & ~n55317;
  assign n55319 = controllable_hmaster2 & ~n55318;
  assign n55320 = ~n44095 & ~n49041;
  assign n55321 = ~controllable_hgrant4 & ~n55320;
  assign n55322 = ~n44083 & ~n55321;
  assign n55323 = ~controllable_hgrant5 & ~n55322;
  assign n55324 = ~n44079 & ~n55323;
  assign n55325 = ~controllable_hmaster2 & ~n55324;
  assign n55326 = ~n55319 & ~n55325;
  assign n55327 = ~controllable_hmaster1 & ~n55326;
  assign n55328 = ~n55311 & ~n55327;
  assign n55329 = i_hlock6 & ~n55328;
  assign n55330 = controllable_hmaster2 & ~n55252;
  assign n55331 = ~n55309 & ~n55330;
  assign n55332 = controllable_hmaster1 & ~n55331;
  assign n55333 = ~n55327 & ~n55332;
  assign n55334 = ~i_hlock6 & ~n55333;
  assign n55335 = ~n55329 & ~n55334;
  assign n55336 = ~controllable_hgrant6 & ~n55335;
  assign n55337 = ~n44017 & ~n55336;
  assign n55338 = ~controllable_hmaster0 & ~n55337;
  assign n55339 = ~n55303 & ~n55338;
  assign n55340 = ~controllable_hmaster3 & ~n55339;
  assign n55341 = ~n55263 & ~n55340;
  assign n55342 = i_hlock7 & ~n55341;
  assign n55343 = ~n8217 & ~n23077;
  assign n55344 = ~n44119 & ~n55343;
  assign n55345 = controllable_hgrant6 & ~n55344;
  assign n55346 = ~n55283 & ~n55330;
  assign n55347 = controllable_hmaster1 & ~n55346;
  assign n55348 = ~n55299 & ~n55347;
  assign n55349 = ~controllable_hgrant6 & ~n55348;
  assign n55350 = ~n55345 & ~n55349;
  assign n55351 = controllable_hmaster0 & ~n55350;
  assign n55352 = ~n55338 & ~n55351;
  assign n55353 = ~controllable_hmaster3 & ~n55352;
  assign n55354 = ~n55263 & ~n55353;
  assign n55355 = ~i_hlock7 & ~n55354;
  assign n55356 = ~n55342 & ~n55355;
  assign n55357 = i_hbusreq7 & ~n55356;
  assign n55358 = i_hbusreq8 & ~n55262;
  assign n55359 = i_hbusreq6 & ~n55232;
  assign n55360 = i_hbusreq5 & ~n55215;
  assign n55361 = i_hbusreq4 & ~n55213;
  assign n55362 = i_hbusreq9 & ~n55213;
  assign n55363 = n8365 & ~n13994;
  assign n55364 = ~n8365 & ~n18741;
  assign n55365 = ~n55363 & ~n55364;
  assign n55366 = i_hlock3 & ~n55365;
  assign n55367 = ~n8365 & ~n18759;
  assign n55368 = ~n55363 & ~n55367;
  assign n55369 = ~i_hlock3 & ~n55368;
  assign n55370 = ~n55366 & ~n55369;
  assign n55371 = ~i_hbusreq3 & ~n55370;
  assign n55372 = ~n49134 & ~n55371;
  assign n55373 = controllable_hgrant3 & ~n55372;
  assign n55374 = ~n44211 & ~n55373;
  assign n55375 = ~i_hbusreq9 & ~n55374;
  assign n55376 = ~n55362 & ~n55375;
  assign n55377 = ~i_hbusreq4 & ~n55376;
  assign n55378 = ~n55361 & ~n55377;
  assign n55379 = ~controllable_hgrant4 & ~n55378;
  assign n55380 = ~n44161 & ~n55379;
  assign n55381 = ~i_hbusreq5 & ~n55380;
  assign n55382 = ~n55360 & ~n55381;
  assign n55383 = ~controllable_hgrant5 & ~n55382;
  assign n55384 = ~n44150 & ~n55383;
  assign n55385 = controllable_hmaster1 & ~n55384;
  assign n55386 = controllable_hmaster2 & ~n55384;
  assign n55387 = i_hbusreq5 & ~n55226;
  assign n55388 = i_hbusreq4 & ~n55224;
  assign n55389 = i_hbusreq9 & ~n55224;
  assign n55390 = n8365 & ~n14028;
  assign n55391 = ~n8365 & ~n18807;
  assign n55392 = ~n55390 & ~n55391;
  assign n55393 = i_hlock3 & ~n55392;
  assign n55394 = ~n8365 & ~n18821;
  assign n55395 = ~n55390 & ~n55394;
  assign n55396 = ~i_hlock3 & ~n55395;
  assign n55397 = ~n55393 & ~n55396;
  assign n55398 = ~i_hbusreq3 & ~n55397;
  assign n55399 = ~n46664 & ~n55398;
  assign n55400 = controllable_hgrant3 & ~n55399;
  assign n55401 = ~n44419 & ~n55400;
  assign n55402 = i_hlock9 & ~n55401;
  assign n55403 = n8365 & ~n14063;
  assign n55404 = ~n8365 & ~n18859;
  assign n55405 = ~n55403 & ~n55404;
  assign n55406 = i_hlock3 & ~n55405;
  assign n55407 = ~n8365 & ~n18871;
  assign n55408 = ~n55403 & ~n55407;
  assign n55409 = ~i_hlock3 & ~n55408;
  assign n55410 = ~n55406 & ~n55409;
  assign n55411 = ~i_hbusreq3 & ~n55410;
  assign n55412 = ~n46728 & ~n55411;
  assign n55413 = controllable_hgrant3 & ~n55412;
  assign n55414 = ~n44493 & ~n55413;
  assign n55415 = ~i_hlock9 & ~n55414;
  assign n55416 = ~n55402 & ~n55415;
  assign n55417 = ~i_hbusreq9 & ~n55416;
  assign n55418 = ~n55389 & ~n55417;
  assign n55419 = ~i_hbusreq4 & ~n55418;
  assign n55420 = ~n55388 & ~n55419;
  assign n55421 = ~controllable_hgrant4 & ~n55420;
  assign n55422 = ~n45193 & ~n55421;
  assign n55423 = ~i_hbusreq5 & ~n55422;
  assign n55424 = ~n55387 & ~n55423;
  assign n55425 = ~controllable_hgrant5 & ~n55424;
  assign n55426 = ~n45182 & ~n55425;
  assign n55427 = ~controllable_hmaster2 & ~n55426;
  assign n55428 = ~n55386 & ~n55427;
  assign n55429 = ~controllable_hmaster1 & ~n55428;
  assign n55430 = ~n55385 & ~n55429;
  assign n55431 = ~i_hbusreq6 & ~n55430;
  assign n55432 = ~n55359 & ~n55431;
  assign n55433 = ~controllable_hgrant6 & ~n55432;
  assign n55434 = ~n45174 & ~n55433;
  assign n55435 = controllable_hmaster0 & ~n55434;
  assign n55436 = i_hbusreq6 & ~n55243;
  assign n55437 = i_hbusreq5 & ~n55237;
  assign n55438 = i_hbusreq4 & ~n55220;
  assign n55439 = i_hbusreq9 & ~n55220;
  assign n55440 = ~i_hbusreq9 & ~n55401;
  assign n55441 = ~n55439 & ~n55440;
  assign n55442 = ~i_hbusreq4 & ~n55441;
  assign n55443 = ~n55438 & ~n55442;
  assign n55444 = ~controllable_hgrant4 & ~n55443;
  assign n55445 = ~n44387 & ~n55444;
  assign n55446 = ~i_hbusreq5 & ~n55445;
  assign n55447 = ~n55437 & ~n55446;
  assign n55448 = ~controllable_hgrant5 & ~n55447;
  assign n55449 = ~n44376 & ~n55448;
  assign n55450 = ~controllable_hmaster2 & ~n55449;
  assign n55451 = ~n55386 & ~n55450;
  assign n55452 = ~controllable_hmaster1 & ~n55451;
  assign n55453 = ~n55385 & ~n55452;
  assign n55454 = ~i_hbusreq6 & ~n55453;
  assign n55455 = ~n55436 & ~n55454;
  assign n55456 = ~controllable_hgrant6 & ~n55455;
  assign n55457 = ~n44368 & ~n55456;
  assign n55458 = ~controllable_hmaster0 & ~n55457;
  assign n55459 = ~n55435 & ~n55458;
  assign n55460 = i_hlock8 & ~n55459;
  assign n55461 = i_hbusreq6 & ~n55256;
  assign n55462 = i_hbusreq5 & ~n55250;
  assign n55463 = i_hbusreq4 & ~n55222;
  assign n55464 = i_hbusreq9 & ~n55222;
  assign n55465 = ~i_hbusreq9 & ~n55414;
  assign n55466 = ~n55464 & ~n55465;
  assign n55467 = ~i_hbusreq4 & ~n55466;
  assign n55468 = ~n55463 & ~n55467;
  assign n55469 = ~controllable_hgrant4 & ~n55468;
  assign n55470 = ~n44467 & ~n55469;
  assign n55471 = ~i_hbusreq5 & ~n55470;
  assign n55472 = ~n55462 & ~n55471;
  assign n55473 = ~controllable_hgrant5 & ~n55472;
  assign n55474 = ~n44456 & ~n55473;
  assign n55475 = ~controllable_hmaster2 & ~n55474;
  assign n55476 = ~n55386 & ~n55475;
  assign n55477 = ~controllable_hmaster1 & ~n55476;
  assign n55478 = ~n55385 & ~n55477;
  assign n55479 = ~i_hbusreq6 & ~n55478;
  assign n55480 = ~n55461 & ~n55479;
  assign n55481 = ~controllable_hgrant6 & ~n55480;
  assign n55482 = ~n44448 & ~n55481;
  assign n55483 = ~controllable_hmaster0 & ~n55482;
  assign n55484 = ~n55435 & ~n55483;
  assign n55485 = ~i_hlock8 & ~n55484;
  assign n55486 = ~n55460 & ~n55485;
  assign n55487 = ~i_hbusreq8 & ~n55486;
  assign n55488 = ~n55358 & ~n55487;
  assign n55489 = controllable_hmaster3 & ~n55488;
  assign n55490 = i_hbusreq8 & ~n55339;
  assign n55491 = i_hbusreq6 & ~n55265;
  assign n55492 = n8217 & ~n15541;
  assign n55493 = ~n8217 & ~n23113;
  assign n55494 = ~n55492 & ~n55493;
  assign n55495 = ~i_hbusreq6 & ~n55494;
  assign n55496 = ~n55491 & ~n55495;
  assign n55497 = controllable_hgrant6 & ~n55496;
  assign n55498 = i_hbusreq6 & ~n55300;
  assign n55499 = controllable_hmaster2 & ~n55449;
  assign n55500 = i_hbusreq5 & ~n55269;
  assign n55501 = n8378 & ~n15533;
  assign n55502 = ~n8378 & ~n23105;
  assign n55503 = ~n55501 & ~n55502;
  assign n55504 = ~i_hbusreq5 & ~n55503;
  assign n55505 = ~n55500 & ~n55504;
  assign n55506 = controllable_hgrant5 & ~n55505;
  assign n55507 = i_hbusreq5 & ~n55280;
  assign n55508 = i_hbusreq4 & ~n55272;
  assign n55509 = i_hbusreq9 & ~n55272;
  assign n55510 = n8426 & ~n15527;
  assign n55511 = ~n8426 & ~n23099;
  assign n55512 = ~n55510 & ~n55511;
  assign n55513 = ~i_hbusreq9 & ~n55512;
  assign n55514 = ~n55509 & ~n55513;
  assign n55515 = ~i_hbusreq4 & ~n55514;
  assign n55516 = ~n55508 & ~n55515;
  assign n55517 = controllable_hgrant4 & ~n55516;
  assign n55518 = i_hbusreq4 & ~n55278;
  assign n55519 = i_hbusreq9 & ~n55278;
  assign n55520 = i_hbusreq3 & ~n55276;
  assign n55521 = i_hlock3 & ~n44310;
  assign n55522 = ~i_hlock3 & ~n44336;
  assign n55523 = ~n55521 & ~n55522;
  assign n55524 = ~i_hbusreq3 & ~n55523;
  assign n55525 = ~n55520 & ~n55524;
  assign n55526 = ~controllable_hgrant3 & ~n55525;
  assign n55527 = ~n49534 & ~n55526;
  assign n55528 = ~i_hbusreq9 & ~n55527;
  assign n55529 = ~n55519 & ~n55528;
  assign n55530 = ~i_hbusreq4 & ~n55529;
  assign n55531 = ~n55518 & ~n55530;
  assign n55532 = ~controllable_hgrant4 & ~n55531;
  assign n55533 = ~n55517 & ~n55532;
  assign n55534 = ~i_hbusreq5 & ~n55533;
  assign n55535 = ~n55507 & ~n55534;
  assign n55536 = ~controllable_hgrant5 & ~n55535;
  assign n55537 = ~n55506 & ~n55536;
  assign n55538 = ~controllable_hmaster2 & ~n55537;
  assign n55539 = ~n55499 & ~n55538;
  assign n55540 = controllable_hmaster1 & ~n55539;
  assign n55541 = i_hbusreq5 & ~n55288;
  assign n55542 = i_hlock5 & ~n55445;
  assign n55543 = ~i_hlock5 & ~n55470;
  assign n55544 = ~n55542 & ~n55543;
  assign n55545 = ~i_hbusreq5 & ~n55544;
  assign n55546 = ~n55541 & ~n55545;
  assign n55547 = ~controllable_hgrant5 & ~n55546;
  assign n55548 = ~n44596 & ~n55547;
  assign n55549 = controllable_hmaster2 & ~n55548;
  assign n55550 = i_hbusreq5 & ~n55294;
  assign n55551 = i_hbusreq4 & ~n55292;
  assign n55552 = i_hbusreq9 & ~n55292;
  assign n55553 = n8365 & ~n14149;
  assign n55554 = ~n8365 & ~n18961;
  assign n55555 = ~n55553 & ~n55554;
  assign n55556 = i_hlock3 & ~n55555;
  assign n55557 = ~n8365 & ~n18975;
  assign n55558 = ~n55553 & ~n55557;
  assign n55559 = ~i_hlock3 & ~n55558;
  assign n55560 = ~n55556 & ~n55559;
  assign n55561 = ~i_hbusreq3 & ~n55560;
  assign n55562 = ~n49611 & ~n55561;
  assign n55563 = controllable_hgrant3 & ~n55562;
  assign n55564 = ~n44657 & ~n55563;
  assign n55565 = ~i_hbusreq9 & ~n55564;
  assign n55566 = ~n55552 & ~n55565;
  assign n55567 = ~i_hbusreq4 & ~n55566;
  assign n55568 = ~n55551 & ~n55567;
  assign n55569 = ~controllable_hgrant4 & ~n55568;
  assign n55570 = ~n44623 & ~n55569;
  assign n55571 = ~i_hbusreq5 & ~n55570;
  assign n55572 = ~n55550 & ~n55571;
  assign n55573 = ~controllable_hgrant5 & ~n55572;
  assign n55574 = ~n44612 & ~n55573;
  assign n55575 = ~controllable_hmaster2 & ~n55574;
  assign n55576 = ~n55549 & ~n55575;
  assign n55577 = ~controllable_hmaster1 & ~n55576;
  assign n55578 = ~n55540 & ~n55577;
  assign n55579 = ~i_hbusreq6 & ~n55578;
  assign n55580 = ~n55498 & ~n55579;
  assign n55581 = ~controllable_hgrant6 & ~n55580;
  assign n55582 = ~n55497 & ~n55581;
  assign n55583 = controllable_hmaster0 & ~n55582;
  assign n55584 = i_hbusreq6 & ~n55335;
  assign n55585 = i_hbusreq5 & ~n55306;
  assign n55586 = i_hbusreq4 & ~n55304;
  assign n55587 = i_hbusreq9 & ~n55304;
  assign n55588 = n8365 & ~n14188;
  assign n55589 = ~n8365 & ~n19011;
  assign n55590 = ~n55588 & ~n55589;
  assign n55591 = i_hlock3 & ~n55590;
  assign n55592 = ~n8365 & ~n19023;
  assign n55593 = ~n55588 & ~n55592;
  assign n55594 = ~i_hlock3 & ~n55593;
  assign n55595 = ~n55591 & ~n55594;
  assign n55596 = ~i_hbusreq3 & ~n55595;
  assign n55597 = ~n49726 & ~n55596;
  assign n55598 = controllable_hgrant3 & ~n55597;
  assign n55599 = ~n44764 & ~n55598;
  assign n55600 = ~i_hbusreq9 & ~n55599;
  assign n55601 = ~n55587 & ~n55600;
  assign n55602 = ~i_hbusreq4 & ~n55601;
  assign n55603 = ~n55586 & ~n55602;
  assign n55604 = ~controllable_hgrant4 & ~n55603;
  assign n55605 = ~n44721 & ~n55604;
  assign n55606 = ~i_hbusreq5 & ~n55605;
  assign n55607 = ~n55585 & ~n55606;
  assign n55608 = ~controllable_hgrant5 & ~n55607;
  assign n55609 = ~n44710 & ~n55608;
  assign n55610 = ~controllable_hmaster2 & ~n55609;
  assign n55611 = ~n55499 & ~n55610;
  assign n55612 = controllable_hmaster1 & ~n55611;
  assign n55613 = i_hbusreq5 & ~n55316;
  assign n55614 = i_hbusreq4 & ~n55314;
  assign n55615 = i_hlock4 & ~n55441;
  assign n55616 = ~i_hlock4 & ~n55466;
  assign n55617 = ~n55615 & ~n55616;
  assign n55618 = ~i_hbusreq4 & ~n55617;
  assign n55619 = ~n55614 & ~n55618;
  assign n55620 = ~controllable_hgrant4 & ~n55619;
  assign n55621 = ~n44805 & ~n55620;
  assign n55622 = ~i_hbusreq5 & ~n55621;
  assign n55623 = ~n55613 & ~n55622;
  assign n55624 = ~controllable_hgrant5 & ~n55623;
  assign n55625 = ~n44785 & ~n55624;
  assign n55626 = controllable_hmaster2 & ~n55625;
  assign n55627 = i_hbusreq5 & ~n55322;
  assign n55628 = i_hbusreq4 & ~n55320;
  assign n55629 = i_hbusreq9 & ~n55320;
  assign n55630 = n8365 & ~n14260;
  assign n55631 = ~n8365 & ~n19092;
  assign n55632 = ~n55630 & ~n55631;
  assign n55633 = i_hlock3 & ~n55632;
  assign n55634 = ~n8365 & ~n19112;
  assign n55635 = ~n55630 & ~n55634;
  assign n55636 = ~i_hlock3 & ~n55635;
  assign n55637 = ~n55633 & ~n55636;
  assign n55638 = ~i_hbusreq3 & ~n55637;
  assign n55639 = ~n49875 & ~n55638;
  assign n55640 = controllable_hgrant3 & ~n55639;
  assign n55641 = ~n44879 & ~n55640;
  assign n55642 = ~i_hbusreq9 & ~n55641;
  assign n55643 = ~n55629 & ~n55642;
  assign n55644 = ~i_hbusreq4 & ~n55643;
  assign n55645 = ~n55628 & ~n55644;
  assign n55646 = ~controllable_hgrant4 & ~n55645;
  assign n55647 = ~n44836 & ~n55646;
  assign n55648 = ~i_hbusreq5 & ~n55647;
  assign n55649 = ~n55627 & ~n55648;
  assign n55650 = ~controllable_hgrant5 & ~n55649;
  assign n55651 = ~n44825 & ~n55650;
  assign n55652 = ~controllable_hmaster2 & ~n55651;
  assign n55653 = ~n55626 & ~n55652;
  assign n55654 = ~controllable_hmaster1 & ~n55653;
  assign n55655 = ~n55612 & ~n55654;
  assign n55656 = i_hlock6 & ~n55655;
  assign n55657 = controllable_hmaster2 & ~n55474;
  assign n55658 = ~n55610 & ~n55657;
  assign n55659 = controllable_hmaster1 & ~n55658;
  assign n55660 = ~n55654 & ~n55659;
  assign n55661 = ~i_hlock6 & ~n55660;
  assign n55662 = ~n55656 & ~n55661;
  assign n55663 = ~i_hbusreq6 & ~n55662;
  assign n55664 = ~n55584 & ~n55663;
  assign n55665 = ~controllable_hgrant6 & ~n55664;
  assign n55666 = ~n44702 & ~n55665;
  assign n55667 = ~controllable_hmaster0 & ~n55666;
  assign n55668 = ~n55583 & ~n55667;
  assign n55669 = ~i_hbusreq8 & ~n55668;
  assign n55670 = ~n55490 & ~n55669;
  assign n55671 = ~controllable_hmaster3 & ~n55670;
  assign n55672 = ~n55489 & ~n55671;
  assign n55673 = i_hlock7 & ~n55672;
  assign n55674 = i_hbusreq8 & ~n55352;
  assign n55675 = i_hbusreq6 & ~n55344;
  assign n55676 = n8217 & ~n15556;
  assign n55677 = ~n8217 & ~n23129;
  assign n55678 = ~n55676 & ~n55677;
  assign n55679 = ~i_hbusreq6 & ~n55678;
  assign n55680 = ~n55675 & ~n55679;
  assign n55681 = controllable_hgrant6 & ~n55680;
  assign n55682 = i_hbusreq6 & ~n55348;
  assign n55683 = ~n55538 & ~n55657;
  assign n55684 = controllable_hmaster1 & ~n55683;
  assign n55685 = ~n55577 & ~n55684;
  assign n55686 = ~i_hbusreq6 & ~n55685;
  assign n55687 = ~n55682 & ~n55686;
  assign n55688 = ~controllable_hgrant6 & ~n55687;
  assign n55689 = ~n55681 & ~n55688;
  assign n55690 = controllable_hmaster0 & ~n55689;
  assign n55691 = ~n55667 & ~n55690;
  assign n55692 = ~i_hbusreq8 & ~n55691;
  assign n55693 = ~n55674 & ~n55692;
  assign n55694 = ~controllable_hmaster3 & ~n55693;
  assign n55695 = ~n55489 & ~n55694;
  assign n55696 = ~i_hlock7 & ~n55695;
  assign n55697 = ~n55673 & ~n55696;
  assign n55698 = ~i_hbusreq7 & ~n55697;
  assign n55699 = ~n55357 & ~n55698;
  assign n55700 = n7924 & ~n55699;
  assign n55701 = ~n55212 & ~n55700;
  assign n55702 = ~n8214 & ~n55701;
  assign n55703 = ~n16349 & ~n48018;
  assign n55704 = ~n7733 & ~n55703;
  assign n55705 = ~n16349 & ~n40226;
  assign n55706 = n7733 & ~n55705;
  assign n55707 = ~n55704 & ~n55706;
  assign n55708 = ~n7928 & ~n55707;
  assign n55709 = ~n48020 & ~n55706;
  assign n55710 = n7928 & ~n55709;
  assign n55711 = ~n55708 & ~n55710;
  assign n55712 = ~controllable_hgrant1 & ~n55711;
  assign n55713 = ~n42721 & ~n55712;
  assign n55714 = ~controllable_hgrant3 & ~n55713;
  assign n55715 = ~n42717 & ~n55714;
  assign n55716 = ~controllable_hgrant4 & ~n55715;
  assign n55717 = ~n42713 & ~n55716;
  assign n55718 = ~controllable_hgrant5 & ~n55717;
  assign n55719 = ~n42709 & ~n55718;
  assign n55720 = controllable_hmaster1 & ~n55719;
  assign n55721 = controllable_hmaster2 & ~n55719;
  assign n55722 = ~n7733 & ~n42761;
  assign n55723 = ~n16724 & ~n40226;
  assign n55724 = n7733 & ~n55723;
  assign n55725 = ~n55722 & ~n55724;
  assign n55726 = n7928 & ~n55725;
  assign n55727 = ~n8221 & ~n55726;
  assign n55728 = ~controllable_hgrant1 & ~n55727;
  assign n55729 = ~n42760 & ~n55728;
  assign n55730 = ~controllable_hgrant3 & ~n55729;
  assign n55731 = ~n42757 & ~n55730;
  assign n55732 = i_hlock9 & ~n55731;
  assign n55733 = ~n8235 & ~n55726;
  assign n55734 = ~controllable_hgrant1 & ~n55733;
  assign n55735 = ~n42795 & ~n55734;
  assign n55736 = ~controllable_hgrant3 & ~n55735;
  assign n55737 = ~n42792 & ~n55736;
  assign n55738 = ~i_hlock9 & ~n55737;
  assign n55739 = ~n55732 & ~n55738;
  assign n55740 = ~controllable_hgrant4 & ~n55739;
  assign n55741 = ~n44951 & ~n55740;
  assign n55742 = ~controllable_hgrant5 & ~n55741;
  assign n55743 = ~n44947 & ~n55742;
  assign n55744 = ~controllable_hmaster2 & ~n55743;
  assign n55745 = ~n55721 & ~n55744;
  assign n55746 = ~controllable_hmaster1 & ~n55745;
  assign n55747 = ~n55720 & ~n55746;
  assign n55748 = ~controllable_hgrant6 & ~n55747;
  assign n55749 = ~n44944 & ~n55748;
  assign n55750 = controllable_hmaster0 & ~n55749;
  assign n55751 = ~controllable_hgrant4 & ~n55731;
  assign n55752 = ~n42754 & ~n55751;
  assign n55753 = ~controllable_hgrant5 & ~n55752;
  assign n55754 = ~n42751 & ~n55753;
  assign n55755 = ~controllable_hmaster2 & ~n55754;
  assign n55756 = ~n55721 & ~n55755;
  assign n55757 = ~controllable_hmaster1 & ~n55756;
  assign n55758 = ~n55720 & ~n55757;
  assign n55759 = ~controllable_hgrant6 & ~n55758;
  assign n55760 = ~n42748 & ~n55759;
  assign n55761 = ~controllable_hmaster0 & ~n55760;
  assign n55762 = ~n55750 & ~n55761;
  assign n55763 = i_hlock8 & ~n55762;
  assign n55764 = ~controllable_hgrant4 & ~n55737;
  assign n55765 = ~n42789 & ~n55764;
  assign n55766 = ~controllable_hgrant5 & ~n55765;
  assign n55767 = ~n42786 & ~n55766;
  assign n55768 = ~controllable_hmaster2 & ~n55767;
  assign n55769 = ~n55721 & ~n55768;
  assign n55770 = ~controllable_hmaster1 & ~n55769;
  assign n55771 = ~n55720 & ~n55770;
  assign n55772 = ~controllable_hgrant6 & ~n55771;
  assign n55773 = ~n42783 & ~n55772;
  assign n55774 = ~controllable_hmaster0 & ~n55773;
  assign n55775 = ~n55750 & ~n55774;
  assign n55776 = ~i_hlock8 & ~n55775;
  assign n55777 = ~n55763 & ~n55776;
  assign n55778 = controllable_hmaster3 & ~n55777;
  assign n55779 = controllable_hmaster2 & ~n55754;
  assign n55780 = i_hlock3 & ~n55729;
  assign n55781 = ~i_hlock3 & ~n55735;
  assign n55782 = ~n55780 & ~n55781;
  assign n55783 = ~controllable_hgrant3 & ~n55782;
  assign n55784 = ~n42838 & ~n55783;
  assign n55785 = ~controllable_hgrant4 & ~n55784;
  assign n55786 = ~n42828 & ~n55785;
  assign n55787 = ~controllable_hgrant5 & ~n55786;
  assign n55788 = ~n42824 & ~n55787;
  assign n55789 = ~controllable_hmaster2 & ~n55788;
  assign n55790 = ~n55779 & ~n55789;
  assign n55791 = controllable_hmaster1 & ~n55790;
  assign n55792 = i_hlock5 & ~n55752;
  assign n55793 = ~i_hlock5 & ~n55765;
  assign n55794 = ~n55792 & ~n55793;
  assign n55795 = ~controllable_hgrant5 & ~n55794;
  assign n55796 = ~n42860 & ~n55795;
  assign n55797 = controllable_hmaster2 & ~n55796;
  assign n55798 = i_hlock1 & ~n55727;
  assign n55799 = ~i_hlock1 & ~n55733;
  assign n55800 = ~n55798 & ~n55799;
  assign n55801 = ~controllable_hgrant1 & ~n55800;
  assign n55802 = ~n42888 & ~n55801;
  assign n55803 = ~controllable_hgrant3 & ~n55802;
  assign n55804 = ~n42878 & ~n55803;
  assign n55805 = ~controllable_hgrant4 & ~n55804;
  assign n55806 = ~n42874 & ~n55805;
  assign n55807 = ~controllable_hgrant5 & ~n55806;
  assign n55808 = ~n42870 & ~n55807;
  assign n55809 = ~controllable_hmaster2 & ~n55808;
  assign n55810 = ~n55797 & ~n55809;
  assign n55811 = ~controllable_hmaster1 & ~n55810;
  assign n55812 = ~n55791 & ~n55811;
  assign n55813 = ~controllable_hgrant6 & ~n55812;
  assign n55814 = ~n42819 & ~n55813;
  assign n55815 = controllable_hmaster0 & ~n55814;
  assign n55816 = ~n18159 & ~n29735;
  assign n55817 = controllable_hmaster1 & ~n55816;
  assign n55818 = ~n19311 & ~n55817;
  assign n55819 = ~n8217 & ~n55818;
  assign n55820 = ~n42910 & ~n55819;
  assign n55821 = i_hlock6 & ~n55820;
  assign n55822 = ~n18159 & ~n29750;
  assign n55823 = controllable_hmaster1 & ~n55822;
  assign n55824 = ~n19311 & ~n55823;
  assign n55825 = ~n8217 & ~n55824;
  assign n55826 = ~n42920 & ~n55825;
  assign n55827 = ~i_hlock6 & ~n55826;
  assign n55828 = ~n55821 & ~n55827;
  assign n55829 = controllable_hgrant6 & ~n55828;
  assign n55830 = ~n48164 & ~n55779;
  assign n55831 = controllable_hmaster1 & ~n55830;
  assign n55832 = i_hlock4 & ~n55731;
  assign n55833 = ~i_hlock4 & ~n55737;
  assign n55834 = ~n55832 & ~n55833;
  assign n55835 = ~controllable_hgrant4 & ~n55834;
  assign n55836 = ~n43000 & ~n55835;
  assign n55837 = ~controllable_hgrant5 & ~n55836;
  assign n55838 = ~n42990 & ~n55837;
  assign n55839 = controllable_hmaster2 & ~n55838;
  assign n55840 = ~n8440 & ~n55726;
  assign n55841 = ~controllable_hgrant1 & ~n55840;
  assign n55842 = ~n43024 & ~n55841;
  assign n55843 = ~controllable_hgrant3 & ~n55842;
  assign n55844 = ~n43020 & ~n55843;
  assign n55845 = ~controllable_hgrant4 & ~n55844;
  assign n55846 = ~n43016 & ~n55845;
  assign n55847 = ~controllable_hgrant5 & ~n55846;
  assign n55848 = ~n43012 & ~n55847;
  assign n55849 = ~controllable_hmaster2 & ~n55848;
  assign n55850 = ~n55839 & ~n55849;
  assign n55851 = ~controllable_hmaster1 & ~n55850;
  assign n55852 = ~n55831 & ~n55851;
  assign n55853 = i_hlock6 & ~n55852;
  assign n55854 = controllable_hmaster2 & ~n55767;
  assign n55855 = ~n48164 & ~n55854;
  assign n55856 = controllable_hmaster1 & ~n55855;
  assign n55857 = ~n55851 & ~n55856;
  assign n55858 = ~i_hlock6 & ~n55857;
  assign n55859 = ~n55853 & ~n55858;
  assign n55860 = ~controllable_hgrant6 & ~n55859;
  assign n55861 = ~n55829 & ~n55860;
  assign n55862 = ~controllable_hmaster0 & ~n55861;
  assign n55863 = ~n55815 & ~n55862;
  assign n55864 = ~controllable_hmaster3 & ~n55863;
  assign n55865 = ~n55778 & ~n55864;
  assign n55866 = i_hlock7 & ~n55865;
  assign n55867 = ~n55789 & ~n55854;
  assign n55868 = controllable_hmaster1 & ~n55867;
  assign n55869 = ~n55811 & ~n55868;
  assign n55870 = ~controllable_hgrant6 & ~n55869;
  assign n55871 = ~n43055 & ~n55870;
  assign n55872 = controllable_hmaster0 & ~n55871;
  assign n55873 = ~n55862 & ~n55872;
  assign n55874 = ~controllable_hmaster3 & ~n55873;
  assign n55875 = ~n55778 & ~n55874;
  assign n55876 = ~i_hlock7 & ~n55875;
  assign n55877 = ~n55866 & ~n55876;
  assign n55878 = i_hbusreq7 & ~n55877;
  assign n55879 = i_hbusreq8 & ~n55777;
  assign n55880 = i_hbusreq6 & ~n55747;
  assign n55881 = i_hbusreq5 & ~n55717;
  assign n55882 = i_hbusreq4 & ~n55715;
  assign n55883 = i_hbusreq9 & ~n55715;
  assign n55884 = i_hbusreq3 & ~n55713;
  assign n55885 = i_hbusreq1 & ~n55711;
  assign n55886 = i_hlock0 & ~n40320;
  assign n55887 = ~i_hlock0 & ~n40216;
  assign n55888 = ~n55886 & ~n55887;
  assign n55889 = ~i_hbusreq0 & ~n55888;
  assign n55890 = ~n51393 & ~n55889;
  assign n55891 = ~i_hbusreq2 & ~n55890;
  assign n55892 = ~n51392 & ~n55891;
  assign n55893 = controllable_hgrant2 & ~n55892;
  assign n55894 = ~n16400 & ~n55893;
  assign n55895 = ~n7733 & ~n55894;
  assign n55896 = i_hlock0 & ~n52901;
  assign n55897 = ~n40342 & ~n55896;
  assign n55898 = ~i_hbusreq0 & ~n55897;
  assign n55899 = ~n40334 & ~n55898;
  assign n55900 = ~i_hbusreq2 & ~n55899;
  assign n55901 = ~n40333 & ~n55900;
  assign n55902 = controllable_hgrant2 & ~n55901;
  assign n55903 = ~n16400 & ~n55902;
  assign n55904 = n7733 & ~n55903;
  assign n55905 = ~n55895 & ~n55904;
  assign n55906 = ~n7928 & ~n55905;
  assign n55907 = ~n43121 & ~n55893;
  assign n55908 = ~n7733 & ~n55907;
  assign n55909 = ~n55904 & ~n55908;
  assign n55910 = n7928 & ~n55909;
  assign n55911 = ~n55906 & ~n55910;
  assign n55912 = ~i_hbusreq1 & ~n55911;
  assign n55913 = ~n55885 & ~n55912;
  assign n55914 = ~controllable_hgrant1 & ~n55913;
  assign n55915 = ~n43111 & ~n55914;
  assign n55916 = ~i_hbusreq3 & ~n55915;
  assign n55917 = ~n55884 & ~n55916;
  assign n55918 = ~controllable_hgrant3 & ~n55917;
  assign n55919 = ~n43103 & ~n55918;
  assign n55920 = ~i_hbusreq9 & ~n55919;
  assign n55921 = ~n55883 & ~n55920;
  assign n55922 = ~i_hbusreq4 & ~n55921;
  assign n55923 = ~n55882 & ~n55922;
  assign n55924 = ~controllable_hgrant4 & ~n55923;
  assign n55925 = ~n43094 & ~n55924;
  assign n55926 = ~i_hbusreq5 & ~n55925;
  assign n55927 = ~n55881 & ~n55926;
  assign n55928 = ~controllable_hgrant5 & ~n55927;
  assign n55929 = ~n43083 & ~n55928;
  assign n55930 = controllable_hmaster1 & ~n55929;
  assign n55931 = controllable_hmaster2 & ~n55929;
  assign n55932 = i_hbusreq5 & ~n55741;
  assign n55933 = i_hbusreq4 & ~n55739;
  assign n55934 = i_hbusreq9 & ~n55739;
  assign n55935 = i_hbusreq3 & ~n55729;
  assign n55936 = i_hbusreq1 & ~n55727;
  assign n55937 = ~n7733 & ~n43200;
  assign n55938 = ~n16796 & ~n55902;
  assign n55939 = n7733 & ~n55938;
  assign n55940 = ~n55937 & ~n55939;
  assign n55941 = n7928 & ~n55940;
  assign n55942 = ~n8265 & ~n55941;
  assign n55943 = ~i_hbusreq1 & ~n55942;
  assign n55944 = ~n55936 & ~n55943;
  assign n55945 = ~controllable_hgrant1 & ~n55944;
  assign n55946 = ~n43198 & ~n55945;
  assign n55947 = ~i_hbusreq3 & ~n55946;
  assign n55948 = ~n55935 & ~n55947;
  assign n55949 = ~controllable_hgrant3 & ~n55948;
  assign n55950 = ~n43190 & ~n55949;
  assign n55951 = i_hlock9 & ~n55950;
  assign n55952 = i_hbusreq3 & ~n55735;
  assign n55953 = i_hbusreq1 & ~n55733;
  assign n55954 = ~n8297 & ~n55941;
  assign n55955 = ~i_hbusreq1 & ~n55954;
  assign n55956 = ~n55953 & ~n55955;
  assign n55957 = ~controllable_hgrant1 & ~n55956;
  assign n55958 = ~n43274 & ~n55957;
  assign n55959 = ~i_hbusreq3 & ~n55958;
  assign n55960 = ~n55952 & ~n55959;
  assign n55961 = ~controllable_hgrant3 & ~n55960;
  assign n55962 = ~n43266 & ~n55961;
  assign n55963 = ~i_hlock9 & ~n55962;
  assign n55964 = ~n55951 & ~n55963;
  assign n55965 = ~i_hbusreq9 & ~n55964;
  assign n55966 = ~n55934 & ~n55965;
  assign n55967 = ~i_hbusreq4 & ~n55966;
  assign n55968 = ~n55933 & ~n55967;
  assign n55969 = ~controllable_hgrant4 & ~n55968;
  assign n55970 = ~n45022 & ~n55969;
  assign n55971 = ~i_hbusreq5 & ~n55970;
  assign n55972 = ~n55932 & ~n55971;
  assign n55973 = ~controllable_hgrant5 & ~n55972;
  assign n55974 = ~n45011 & ~n55973;
  assign n55975 = ~controllable_hmaster2 & ~n55974;
  assign n55976 = ~n55931 & ~n55975;
  assign n55977 = ~controllable_hmaster1 & ~n55976;
  assign n55978 = ~n55930 & ~n55977;
  assign n55979 = ~i_hbusreq6 & ~n55978;
  assign n55980 = ~n55880 & ~n55979;
  assign n55981 = ~controllable_hgrant6 & ~n55980;
  assign n55982 = ~n45003 & ~n55981;
  assign n55983 = controllable_hmaster0 & ~n55982;
  assign n55984 = i_hbusreq6 & ~n55758;
  assign n55985 = i_hbusreq5 & ~n55752;
  assign n55986 = i_hbusreq4 & ~n55731;
  assign n55987 = i_hbusreq9 & ~n55731;
  assign n55988 = ~i_hbusreq9 & ~n55950;
  assign n55989 = ~n55987 & ~n55988;
  assign n55990 = ~i_hbusreq4 & ~n55989;
  assign n55991 = ~n55986 & ~n55990;
  assign n55992 = ~controllable_hgrant4 & ~n55991;
  assign n55993 = ~n43181 & ~n55992;
  assign n55994 = ~i_hbusreq5 & ~n55993;
  assign n55995 = ~n55985 & ~n55994;
  assign n55996 = ~controllable_hgrant5 & ~n55995;
  assign n55997 = ~n43170 & ~n55996;
  assign n55998 = ~controllable_hmaster2 & ~n55997;
  assign n55999 = ~n55931 & ~n55998;
  assign n56000 = ~controllable_hmaster1 & ~n55999;
  assign n56001 = ~n55930 & ~n56000;
  assign n56002 = ~i_hbusreq6 & ~n56001;
  assign n56003 = ~n55984 & ~n56002;
  assign n56004 = ~controllable_hgrant6 & ~n56003;
  assign n56005 = ~n43162 & ~n56004;
  assign n56006 = ~controllable_hmaster0 & ~n56005;
  assign n56007 = ~n55983 & ~n56006;
  assign n56008 = i_hlock8 & ~n56007;
  assign n56009 = i_hbusreq6 & ~n55771;
  assign n56010 = i_hbusreq5 & ~n55765;
  assign n56011 = i_hbusreq4 & ~n55737;
  assign n56012 = i_hbusreq9 & ~n55737;
  assign n56013 = ~i_hbusreq9 & ~n55962;
  assign n56014 = ~n56012 & ~n56013;
  assign n56015 = ~i_hbusreq4 & ~n56014;
  assign n56016 = ~n56011 & ~n56015;
  assign n56017 = ~controllable_hgrant4 & ~n56016;
  assign n56018 = ~n43257 & ~n56017;
  assign n56019 = ~i_hbusreq5 & ~n56018;
  assign n56020 = ~n56010 & ~n56019;
  assign n56021 = ~controllable_hgrant5 & ~n56020;
  assign n56022 = ~n43246 & ~n56021;
  assign n56023 = ~controllable_hmaster2 & ~n56022;
  assign n56024 = ~n55931 & ~n56023;
  assign n56025 = ~controllable_hmaster1 & ~n56024;
  assign n56026 = ~n55930 & ~n56025;
  assign n56027 = ~i_hbusreq6 & ~n56026;
  assign n56028 = ~n56009 & ~n56027;
  assign n56029 = ~controllable_hgrant6 & ~n56028;
  assign n56030 = ~n43238 & ~n56029;
  assign n56031 = ~controllable_hmaster0 & ~n56030;
  assign n56032 = ~n55983 & ~n56031;
  assign n56033 = ~i_hlock8 & ~n56032;
  assign n56034 = ~n56008 & ~n56033;
  assign n56035 = ~i_hbusreq8 & ~n56034;
  assign n56036 = ~n55879 & ~n56035;
  assign n56037 = controllable_hmaster3 & ~n56036;
  assign n56038 = i_hbusreq8 & ~n55863;
  assign n56039 = i_hbusreq6 & ~n55812;
  assign n56040 = controllable_hmaster2 & ~n55997;
  assign n56041 = i_hbusreq5 & ~n55786;
  assign n56042 = i_hbusreq4 & ~n55784;
  assign n56043 = i_hbusreq9 & ~n55784;
  assign n56044 = i_hbusreq3 & ~n55782;
  assign n56045 = i_hlock3 & ~n55946;
  assign n56046 = ~i_hlock3 & ~n55958;
  assign n56047 = ~n56045 & ~n56046;
  assign n56048 = ~i_hbusreq3 & ~n56047;
  assign n56049 = ~n56044 & ~n56048;
  assign n56050 = ~controllable_hgrant3 & ~n56049;
  assign n56051 = ~n43352 & ~n56050;
  assign n56052 = ~i_hbusreq9 & ~n56051;
  assign n56053 = ~n56043 & ~n56052;
  assign n56054 = ~i_hbusreq4 & ~n56053;
  assign n56055 = ~n56042 & ~n56054;
  assign n56056 = ~controllable_hgrant4 & ~n56055;
  assign n56057 = ~n43337 & ~n56056;
  assign n56058 = ~i_hbusreq5 & ~n56057;
  assign n56059 = ~n56041 & ~n56058;
  assign n56060 = ~controllable_hgrant5 & ~n56059;
  assign n56061 = ~n43326 & ~n56060;
  assign n56062 = ~controllable_hmaster2 & ~n56061;
  assign n56063 = ~n56040 & ~n56062;
  assign n56064 = controllable_hmaster1 & ~n56063;
  assign n56065 = i_hbusreq5 & ~n55794;
  assign n56066 = i_hlock5 & ~n55993;
  assign n56067 = ~i_hlock5 & ~n56018;
  assign n56068 = ~n56066 & ~n56067;
  assign n56069 = ~i_hbusreq5 & ~n56068;
  assign n56070 = ~n56065 & ~n56069;
  assign n56071 = ~controllable_hgrant5 & ~n56070;
  assign n56072 = ~n43386 & ~n56071;
  assign n56073 = controllable_hmaster2 & ~n56072;
  assign n56074 = i_hbusreq5 & ~n55806;
  assign n56075 = i_hbusreq4 & ~n55804;
  assign n56076 = i_hbusreq9 & ~n55804;
  assign n56077 = i_hbusreq3 & ~n55802;
  assign n56078 = i_hbusreq1 & ~n55800;
  assign n56079 = i_hlock1 & ~n55942;
  assign n56080 = ~i_hlock1 & ~n55954;
  assign n56081 = ~n56079 & ~n56080;
  assign n56082 = ~i_hbusreq1 & ~n56081;
  assign n56083 = ~n56078 & ~n56082;
  assign n56084 = ~controllable_hgrant1 & ~n56083;
  assign n56085 = ~n43436 & ~n56084;
  assign n56086 = ~i_hbusreq3 & ~n56085;
  assign n56087 = ~n56077 & ~n56086;
  assign n56088 = ~controllable_hgrant3 & ~n56087;
  assign n56089 = ~n43422 & ~n56088;
  assign n56090 = ~i_hbusreq9 & ~n56089;
  assign n56091 = ~n56076 & ~n56090;
  assign n56092 = ~i_hbusreq4 & ~n56091;
  assign n56093 = ~n56075 & ~n56092;
  assign n56094 = ~controllable_hgrant4 & ~n56093;
  assign n56095 = ~n43413 & ~n56094;
  assign n56096 = ~i_hbusreq5 & ~n56095;
  assign n56097 = ~n56074 & ~n56096;
  assign n56098 = ~controllable_hgrant5 & ~n56097;
  assign n56099 = ~n43402 & ~n56098;
  assign n56100 = ~controllable_hmaster2 & ~n56099;
  assign n56101 = ~n56073 & ~n56100;
  assign n56102 = ~controllable_hmaster1 & ~n56101;
  assign n56103 = ~n56064 & ~n56102;
  assign n56104 = ~i_hbusreq6 & ~n56103;
  assign n56105 = ~n56039 & ~n56104;
  assign n56106 = ~controllable_hgrant6 & ~n56105;
  assign n56107 = ~n43317 & ~n56106;
  assign n56108 = controllable_hmaster0 & ~n56107;
  assign n56109 = i_hbusreq6 & ~n55828;
  assign n56110 = ~n9678 & ~n27226;
  assign n56111 = controllable_hmaster1 & ~n56110;
  assign n56112 = ~n9428 & ~n56111;
  assign n56113 = n8217 & ~n56112;
  assign n56114 = ~n21759 & ~n29796;
  assign n56115 = controllable_hmaster1 & ~n56114;
  assign n56116 = ~n19626 & ~n56115;
  assign n56117 = ~n8217 & ~n56116;
  assign n56118 = ~n56113 & ~n56117;
  assign n56119 = i_hlock6 & ~n56118;
  assign n56120 = ~n9678 & ~n27253;
  assign n56121 = controllable_hmaster1 & ~n56120;
  assign n56122 = ~n9428 & ~n56121;
  assign n56123 = n8217 & ~n56122;
  assign n56124 = ~n21759 & ~n29826;
  assign n56125 = controllable_hmaster1 & ~n56124;
  assign n56126 = ~n19626 & ~n56125;
  assign n56127 = ~n8217 & ~n56126;
  assign n56128 = ~n56123 & ~n56127;
  assign n56129 = ~i_hlock6 & ~n56128;
  assign n56130 = ~n56119 & ~n56129;
  assign n56131 = ~i_hbusreq6 & ~n56130;
  assign n56132 = ~n56109 & ~n56131;
  assign n56133 = controllable_hgrant6 & ~n56132;
  assign n56134 = i_hbusreq6 & ~n55859;
  assign n56135 = ~n48606 & ~n56040;
  assign n56136 = controllable_hmaster1 & ~n56135;
  assign n56137 = i_hbusreq5 & ~n55836;
  assign n56138 = i_hbusreq4 & ~n55834;
  assign n56139 = i_hlock4 & ~n55989;
  assign n56140 = ~i_hlock4 & ~n56014;
  assign n56141 = ~n56139 & ~n56140;
  assign n56142 = ~i_hbusreq4 & ~n56141;
  assign n56143 = ~n56138 & ~n56142;
  assign n56144 = ~controllable_hgrant4 & ~n56143;
  assign n56145 = ~n43609 & ~n56144;
  assign n56146 = ~i_hbusreq5 & ~n56145;
  assign n56147 = ~n56137 & ~n56146;
  assign n56148 = ~controllable_hgrant5 & ~n56147;
  assign n56149 = ~n43589 & ~n56148;
  assign n56150 = controllable_hmaster2 & ~n56149;
  assign n56151 = i_hbusreq5 & ~n55846;
  assign n56152 = i_hbusreq4 & ~n55844;
  assign n56153 = i_hbusreq9 & ~n55844;
  assign n56154 = i_hbusreq3 & ~n55842;
  assign n56155 = i_hbusreq1 & ~n55840;
  assign n56156 = ~n7733 & ~n43670;
  assign n56157 = ~n7818 & ~n43659;
  assign n56158 = controllable_locked & ~n56157;
  assign n56159 = ~n43661 & ~n56158;
  assign n56160 = i_hlock0 & ~n56159;
  assign n56161 = ~n40342 & ~n56160;
  assign n56162 = ~i_hbusreq0 & ~n56161;
  assign n56163 = ~n40334 & ~n56162;
  assign n56164 = ~i_hbusreq2 & ~n56163;
  assign n56165 = ~n40333 & ~n56164;
  assign n56166 = controllable_hgrant2 & ~n56165;
  assign n56167 = ~n18452 & ~n56166;
  assign n56168 = n7733 & ~n56167;
  assign n56169 = ~n56156 & ~n56168;
  assign n56170 = n7928 & ~n56169;
  assign n56171 = ~n8440 & ~n56170;
  assign n56172 = ~i_hbusreq1 & ~n56171;
  assign n56173 = ~n56155 & ~n56172;
  assign n56174 = ~controllable_hgrant1 & ~n56173;
  assign n56175 = ~n43657 & ~n56174;
  assign n56176 = ~i_hbusreq3 & ~n56175;
  assign n56177 = ~n56154 & ~n56176;
  assign n56178 = ~controllable_hgrant3 & ~n56177;
  assign n56179 = ~n43649 & ~n56178;
  assign n56180 = ~i_hbusreq9 & ~n56179;
  assign n56181 = ~n56153 & ~n56180;
  assign n56182 = ~i_hbusreq4 & ~n56181;
  assign n56183 = ~n56152 & ~n56182;
  assign n56184 = ~controllable_hgrant4 & ~n56183;
  assign n56185 = ~n43640 & ~n56184;
  assign n56186 = ~i_hbusreq5 & ~n56185;
  assign n56187 = ~n56151 & ~n56186;
  assign n56188 = ~controllable_hgrant5 & ~n56187;
  assign n56189 = ~n43629 & ~n56188;
  assign n56190 = ~controllable_hmaster2 & ~n56189;
  assign n56191 = ~n56150 & ~n56190;
  assign n56192 = ~controllable_hmaster1 & ~n56191;
  assign n56193 = ~n56136 & ~n56192;
  assign n56194 = i_hlock6 & ~n56193;
  assign n56195 = controllable_hmaster2 & ~n56022;
  assign n56196 = ~n48606 & ~n56195;
  assign n56197 = controllable_hmaster1 & ~n56196;
  assign n56198 = ~n56192 & ~n56197;
  assign n56199 = ~i_hlock6 & ~n56198;
  assign n56200 = ~n56194 & ~n56199;
  assign n56201 = ~i_hbusreq6 & ~n56200;
  assign n56202 = ~n56134 & ~n56201;
  assign n56203 = ~controllable_hgrant6 & ~n56202;
  assign n56204 = ~n56133 & ~n56203;
  assign n56205 = ~controllable_hmaster0 & ~n56204;
  assign n56206 = ~n56108 & ~n56205;
  assign n56207 = ~i_hbusreq8 & ~n56206;
  assign n56208 = ~n56038 & ~n56207;
  assign n56209 = ~controllable_hmaster3 & ~n56208;
  assign n56210 = ~n56037 & ~n56209;
  assign n56211 = i_hlock7 & ~n56210;
  assign n56212 = i_hbusreq8 & ~n55873;
  assign n56213 = i_hbusreq6 & ~n55869;
  assign n56214 = ~n56062 & ~n56195;
  assign n56215 = controllable_hmaster1 & ~n56214;
  assign n56216 = ~n56102 & ~n56215;
  assign n56217 = ~i_hbusreq6 & ~n56216;
  assign n56218 = ~n56213 & ~n56217;
  assign n56219 = ~controllable_hgrant6 & ~n56218;
  assign n56220 = ~n43720 & ~n56219;
  assign n56221 = controllable_hmaster0 & ~n56220;
  assign n56222 = ~n56205 & ~n56221;
  assign n56223 = ~i_hbusreq8 & ~n56222;
  assign n56224 = ~n56212 & ~n56223;
  assign n56225 = ~controllable_hmaster3 & ~n56224;
  assign n56226 = ~n56037 & ~n56225;
  assign n56227 = ~i_hlock7 & ~n56226;
  assign n56228 = ~n56211 & ~n56227;
  assign n56229 = ~i_hbusreq7 & ~n56228;
  assign n56230 = ~n55878 & ~n56229;
  assign n56231 = ~n7924 & ~n56230;
  assign n56232 = ~n16505 & ~n46060;
  assign n56233 = n7733 & ~n56232;
  assign n56234 = ~n48798 & ~n56233;
  assign n56235 = n7928 & ~n56234;
  assign n56236 = ~n55708 & ~n56235;
  assign n56237 = ~controllable_hgrant1 & ~n56236;
  assign n56238 = ~n43758 & ~n56237;
  assign n56239 = ~controllable_hgrant3 & ~n56238;
  assign n56240 = ~n43754 & ~n56239;
  assign n56241 = ~controllable_hgrant4 & ~n56240;
  assign n56242 = ~n43750 & ~n56241;
  assign n56243 = ~controllable_hgrant5 & ~n56242;
  assign n56244 = ~n43746 & ~n56243;
  assign n56245 = controllable_hmaster1 & ~n56244;
  assign n56246 = controllable_hmaster2 & ~n56244;
  assign n56247 = ~n17505 & ~n46060;
  assign n56248 = n7733 & ~n56247;
  assign n56249 = ~n43847 & ~n56248;
  assign n56250 = n7928 & ~n56249;
  assign n56251 = ~n8221 & ~n56250;
  assign n56252 = ~controllable_hgrant1 & ~n56251;
  assign n56253 = ~n43845 & ~n56252;
  assign n56254 = ~controllable_hgrant3 & ~n56253;
  assign n56255 = ~n43842 & ~n56254;
  assign n56256 = i_hlock9 & ~n56255;
  assign n56257 = ~n8235 & ~n56250;
  assign n56258 = ~controllable_hgrant1 & ~n56257;
  assign n56259 = ~n43884 & ~n56258;
  assign n56260 = ~controllable_hgrant3 & ~n56259;
  assign n56261 = ~n43881 & ~n56260;
  assign n56262 = ~i_hlock9 & ~n56261;
  assign n56263 = ~n56256 & ~n56262;
  assign n56264 = ~controllable_hgrant4 & ~n56263;
  assign n56265 = ~n45104 & ~n56264;
  assign n56266 = ~controllable_hgrant5 & ~n56265;
  assign n56267 = ~n45100 & ~n56266;
  assign n56268 = ~controllable_hmaster2 & ~n56267;
  assign n56269 = ~n56246 & ~n56268;
  assign n56270 = ~controllable_hmaster1 & ~n56269;
  assign n56271 = ~n56245 & ~n56270;
  assign n56272 = ~controllable_hgrant6 & ~n56271;
  assign n56273 = ~n45097 & ~n56272;
  assign n56274 = controllable_hmaster0 & ~n56273;
  assign n56275 = ~controllable_hgrant4 & ~n56255;
  assign n56276 = ~n43839 & ~n56275;
  assign n56277 = ~controllable_hgrant5 & ~n56276;
  assign n56278 = ~n43836 & ~n56277;
  assign n56279 = ~controllable_hmaster2 & ~n56278;
  assign n56280 = ~n56246 & ~n56279;
  assign n56281 = ~controllable_hmaster1 & ~n56280;
  assign n56282 = ~n56245 & ~n56281;
  assign n56283 = ~controllable_hgrant6 & ~n56282;
  assign n56284 = ~n43833 & ~n56283;
  assign n56285 = ~controllable_hmaster0 & ~n56284;
  assign n56286 = ~n56274 & ~n56285;
  assign n56287 = i_hlock8 & ~n56286;
  assign n56288 = ~controllable_hgrant4 & ~n56261;
  assign n56289 = ~n43878 & ~n56288;
  assign n56290 = ~controllable_hgrant5 & ~n56289;
  assign n56291 = ~n43875 & ~n56290;
  assign n56292 = ~controllable_hmaster2 & ~n56291;
  assign n56293 = ~n56246 & ~n56292;
  assign n56294 = ~controllable_hmaster1 & ~n56293;
  assign n56295 = ~n56245 & ~n56294;
  assign n56296 = ~controllable_hgrant6 & ~n56295;
  assign n56297 = ~n43872 & ~n56296;
  assign n56298 = ~controllable_hmaster0 & ~n56297;
  assign n56299 = ~n56274 & ~n56298;
  assign n56300 = ~i_hlock8 & ~n56299;
  assign n56301 = ~n56287 & ~n56300;
  assign n56302 = controllable_hmaster3 & ~n56301;
  assign n56303 = controllable_hmaster2 & ~n56278;
  assign n56304 = i_hlock3 & ~n56253;
  assign n56305 = ~i_hlock3 & ~n56259;
  assign n56306 = ~n56304 & ~n56305;
  assign n56307 = ~controllable_hgrant3 & ~n56306;
  assign n56308 = ~n43927 & ~n56307;
  assign n56309 = ~controllable_hgrant4 & ~n56308;
  assign n56310 = ~n43917 & ~n56309;
  assign n56311 = ~controllable_hgrant5 & ~n56310;
  assign n56312 = ~n43913 & ~n56311;
  assign n56313 = ~controllable_hmaster2 & ~n56312;
  assign n56314 = ~n56303 & ~n56313;
  assign n56315 = controllable_hmaster1 & ~n56314;
  assign n56316 = i_hlock5 & ~n56276;
  assign n56317 = ~i_hlock5 & ~n56289;
  assign n56318 = ~n56316 & ~n56317;
  assign n56319 = ~controllable_hgrant5 & ~n56318;
  assign n56320 = ~n43949 & ~n56319;
  assign n56321 = controllable_hmaster2 & ~n56320;
  assign n56322 = i_hlock1 & ~n56251;
  assign n56323 = ~i_hlock1 & ~n56257;
  assign n56324 = ~n56322 & ~n56323;
  assign n56325 = ~controllable_hgrant1 & ~n56324;
  assign n56326 = ~n43977 & ~n56325;
  assign n56327 = ~controllable_hgrant3 & ~n56326;
  assign n56328 = ~n43967 & ~n56327;
  assign n56329 = ~controllable_hgrant4 & ~n56328;
  assign n56330 = ~n43963 & ~n56329;
  assign n56331 = ~controllable_hgrant5 & ~n56330;
  assign n56332 = ~n43959 & ~n56331;
  assign n56333 = ~controllable_hmaster2 & ~n56332;
  assign n56334 = ~n56321 & ~n56333;
  assign n56335 = ~controllable_hmaster1 & ~n56334;
  assign n56336 = ~n56315 & ~n56335;
  assign n56337 = ~controllable_hgrant6 & ~n56336;
  assign n56338 = ~n43908 & ~n56337;
  assign n56339 = controllable_hmaster0 & ~n56338;
  assign n56340 = ~n23211 & ~n29869;
  assign n56341 = controllable_hmaster1 & ~n56340;
  assign n56342 = ~n19836 & ~n56341;
  assign n56343 = ~n8217 & ~n56342;
  assign n56344 = ~n43999 & ~n56343;
  assign n56345 = i_hlock6 & ~n56344;
  assign n56346 = ~n23211 & ~n29884;
  assign n56347 = controllable_hmaster1 & ~n56346;
  assign n56348 = ~n19836 & ~n56347;
  assign n56349 = ~n8217 & ~n56348;
  assign n56350 = ~n44009 & ~n56349;
  assign n56351 = ~i_hlock6 & ~n56350;
  assign n56352 = ~n56345 & ~n56351;
  assign n56353 = controllable_hgrant6 & ~n56352;
  assign n56354 = ~n8378 & ~n23208;
  assign n56355 = ~n44018 & ~n56354;
  assign n56356 = controllable_hgrant5 & ~n56355;
  assign n56357 = ~n8426 & ~n23206;
  assign n56358 = ~n44022 & ~n56357;
  assign n56359 = controllable_hgrant4 & ~n56358;
  assign n56360 = ~n8365 & ~n23204;
  assign n56361 = ~n44026 & ~n56360;
  assign n56362 = controllable_hgrant3 & ~n56361;
  assign n56363 = ~n8389 & ~n23202;
  assign n56364 = ~n44030 & ~n56363;
  assign n56365 = controllable_hgrant1 & ~n56364;
  assign n56366 = ~n17090 & ~n48978;
  assign n56367 = n7733 & ~n56366;
  assign n56368 = ~n48968 & ~n56367;
  assign n56369 = n7928 & ~n56368;
  assign n56370 = ~n42965 & ~n56369;
  assign n56371 = ~controllable_hgrant1 & ~n56370;
  assign n56372 = ~n56365 & ~n56371;
  assign n56373 = ~controllable_hgrant3 & ~n56372;
  assign n56374 = ~n56362 & ~n56373;
  assign n56375 = ~controllable_hgrant4 & ~n56374;
  assign n56376 = ~n56359 & ~n56375;
  assign n56377 = ~controllable_hgrant5 & ~n56376;
  assign n56378 = ~n56356 & ~n56377;
  assign n56379 = ~controllable_hmaster2 & ~n56378;
  assign n56380 = ~n56303 & ~n56379;
  assign n56381 = controllable_hmaster1 & ~n56380;
  assign n56382 = i_hlock4 & ~n56255;
  assign n56383 = ~i_hlock4 & ~n56261;
  assign n56384 = ~n56382 & ~n56383;
  assign n56385 = ~controllable_hgrant4 & ~n56384;
  assign n56386 = ~n44067 & ~n56385;
  assign n56387 = ~controllable_hgrant5 & ~n56386;
  assign n56388 = ~n44057 & ~n56387;
  assign n56389 = controllable_hmaster2 & ~n56388;
  assign n56390 = ~n8440 & ~n56250;
  assign n56391 = ~controllable_hgrant1 & ~n56390;
  assign n56392 = ~n44091 & ~n56391;
  assign n56393 = ~controllable_hgrant3 & ~n56392;
  assign n56394 = ~n44087 & ~n56393;
  assign n56395 = ~controllable_hgrant4 & ~n56394;
  assign n56396 = ~n44083 & ~n56395;
  assign n56397 = ~controllable_hgrant5 & ~n56396;
  assign n56398 = ~n44079 & ~n56397;
  assign n56399 = ~controllable_hmaster2 & ~n56398;
  assign n56400 = ~n56389 & ~n56399;
  assign n56401 = ~controllable_hmaster1 & ~n56400;
  assign n56402 = ~n56381 & ~n56401;
  assign n56403 = i_hlock6 & ~n56402;
  assign n56404 = controllable_hmaster2 & ~n56291;
  assign n56405 = ~n56379 & ~n56404;
  assign n56406 = controllable_hmaster1 & ~n56405;
  assign n56407 = ~n56401 & ~n56406;
  assign n56408 = ~i_hlock6 & ~n56407;
  assign n56409 = ~n56403 & ~n56408;
  assign n56410 = ~controllable_hgrant6 & ~n56409;
  assign n56411 = ~n56353 & ~n56410;
  assign n56412 = ~controllable_hmaster0 & ~n56411;
  assign n56413 = ~n56339 & ~n56412;
  assign n56414 = ~controllable_hmaster3 & ~n56413;
  assign n56415 = ~n56302 & ~n56414;
  assign n56416 = i_hlock7 & ~n56415;
  assign n56417 = ~n56313 & ~n56404;
  assign n56418 = controllable_hmaster1 & ~n56417;
  assign n56419 = ~n56335 & ~n56418;
  assign n56420 = ~controllable_hgrant6 & ~n56419;
  assign n56421 = ~n44122 & ~n56420;
  assign n56422 = controllable_hmaster0 & ~n56421;
  assign n56423 = ~n56412 & ~n56422;
  assign n56424 = ~controllable_hmaster3 & ~n56423;
  assign n56425 = ~n56302 & ~n56424;
  assign n56426 = ~i_hlock7 & ~n56425;
  assign n56427 = ~n56416 & ~n56426;
  assign n56428 = i_hbusreq7 & ~n56427;
  assign n56429 = i_hbusreq8 & ~n56301;
  assign n56430 = i_hbusreq6 & ~n56271;
  assign n56431 = i_hbusreq5 & ~n56242;
  assign n56432 = i_hbusreq4 & ~n56240;
  assign n56433 = i_hbusreq9 & ~n56240;
  assign n56434 = i_hbusreq3 & ~n56238;
  assign n56435 = i_hbusreq1 & ~n56236;
  assign n56436 = ~n49166 & ~n51511;
  assign n56437 = ~i_hbusreq0 & ~n56436;
  assign n56438 = ~n49162 & ~n56437;
  assign n56439 = ~i_hbusreq2 & ~n56438;
  assign n56440 = ~n49161 & ~n56439;
  assign n56441 = controllable_hgrant2 & ~n56440;
  assign n56442 = ~n44197 & ~n56441;
  assign n56443 = ~n7733 & ~n56442;
  assign n56444 = i_hlock0 & ~n53192;
  assign n56445 = ~n46695 & ~n56444;
  assign n56446 = ~i_hbusreq0 & ~n56445;
  assign n56447 = ~n46689 & ~n56446;
  assign n56448 = i_hlock2 & ~n56447;
  assign n56449 = ~n46700 & ~n56446;
  assign n56450 = ~i_hlock2 & ~n56449;
  assign n56451 = ~n56448 & ~n56450;
  assign n56452 = ~i_hbusreq2 & ~n56451;
  assign n56453 = ~n46688 & ~n56452;
  assign n56454 = controllable_hgrant2 & ~n56453;
  assign n56455 = ~n16633 & ~n56454;
  assign n56456 = n7733 & ~n56455;
  assign n56457 = ~n56443 & ~n56456;
  assign n56458 = n7928 & ~n56457;
  assign n56459 = ~n55906 & ~n56458;
  assign n56460 = ~i_hbusreq1 & ~n56459;
  assign n56461 = ~n56435 & ~n56460;
  assign n56462 = ~controllable_hgrant1 & ~n56461;
  assign n56463 = ~n44178 & ~n56462;
  assign n56464 = ~i_hbusreq3 & ~n56463;
  assign n56465 = ~n56434 & ~n56464;
  assign n56466 = ~controllable_hgrant3 & ~n56465;
  assign n56467 = ~n44170 & ~n56466;
  assign n56468 = ~i_hbusreq9 & ~n56467;
  assign n56469 = ~n56433 & ~n56468;
  assign n56470 = ~i_hbusreq4 & ~n56469;
  assign n56471 = ~n56432 & ~n56470;
  assign n56472 = ~controllable_hgrant4 & ~n56471;
  assign n56473 = ~n44161 & ~n56472;
  assign n56474 = ~i_hbusreq5 & ~n56473;
  assign n56475 = ~n56431 & ~n56474;
  assign n56476 = ~controllable_hgrant5 & ~n56475;
  assign n56477 = ~n44150 & ~n56476;
  assign n56478 = controllable_hmaster1 & ~n56477;
  assign n56479 = controllable_hmaster2 & ~n56477;
  assign n56480 = i_hbusreq5 & ~n56265;
  assign n56481 = i_hbusreq4 & ~n56263;
  assign n56482 = i_hbusreq9 & ~n56263;
  assign n56483 = i_hbusreq3 & ~n56253;
  assign n56484 = i_hbusreq1 & ~n56251;
  assign n56485 = ~n18798 & ~n56454;
  assign n56486 = n7733 & ~n56485;
  assign n56487 = ~n44407 & ~n56486;
  assign n56488 = n7928 & ~n56487;
  assign n56489 = ~n8265 & ~n56488;
  assign n56490 = ~i_hbusreq1 & ~n56489;
  assign n56491 = ~n56484 & ~n56490;
  assign n56492 = ~controllable_hgrant1 & ~n56491;
  assign n56493 = ~n44404 & ~n56492;
  assign n56494 = ~i_hbusreq3 & ~n56493;
  assign n56495 = ~n56483 & ~n56494;
  assign n56496 = ~controllable_hgrant3 & ~n56495;
  assign n56497 = ~n44396 & ~n56496;
  assign n56498 = i_hlock9 & ~n56497;
  assign n56499 = i_hbusreq3 & ~n56259;
  assign n56500 = i_hbusreq1 & ~n56257;
  assign n56501 = ~n8297 & ~n56488;
  assign n56502 = ~i_hbusreq1 & ~n56501;
  assign n56503 = ~n56500 & ~n56502;
  assign n56504 = ~controllable_hgrant1 & ~n56503;
  assign n56505 = ~n44484 & ~n56504;
  assign n56506 = ~i_hbusreq3 & ~n56505;
  assign n56507 = ~n56499 & ~n56506;
  assign n56508 = ~controllable_hgrant3 & ~n56507;
  assign n56509 = ~n44476 & ~n56508;
  assign n56510 = ~i_hlock9 & ~n56509;
  assign n56511 = ~n56498 & ~n56510;
  assign n56512 = ~i_hbusreq9 & ~n56511;
  assign n56513 = ~n56482 & ~n56512;
  assign n56514 = ~i_hbusreq4 & ~n56513;
  assign n56515 = ~n56481 & ~n56514;
  assign n56516 = ~controllable_hgrant4 & ~n56515;
  assign n56517 = ~n45193 & ~n56516;
  assign n56518 = ~i_hbusreq5 & ~n56517;
  assign n56519 = ~n56480 & ~n56518;
  assign n56520 = ~controllable_hgrant5 & ~n56519;
  assign n56521 = ~n45182 & ~n56520;
  assign n56522 = ~controllable_hmaster2 & ~n56521;
  assign n56523 = ~n56479 & ~n56522;
  assign n56524 = ~controllable_hmaster1 & ~n56523;
  assign n56525 = ~n56478 & ~n56524;
  assign n56526 = ~i_hbusreq6 & ~n56525;
  assign n56527 = ~n56430 & ~n56526;
  assign n56528 = ~controllable_hgrant6 & ~n56527;
  assign n56529 = ~n45174 & ~n56528;
  assign n56530 = controllable_hmaster0 & ~n56529;
  assign n56531 = i_hbusreq6 & ~n56282;
  assign n56532 = i_hbusreq5 & ~n56276;
  assign n56533 = i_hbusreq4 & ~n56255;
  assign n56534 = i_hbusreq9 & ~n56255;
  assign n56535 = ~i_hbusreq9 & ~n56497;
  assign n56536 = ~n56534 & ~n56535;
  assign n56537 = ~i_hbusreq4 & ~n56536;
  assign n56538 = ~n56533 & ~n56537;
  assign n56539 = ~controllable_hgrant4 & ~n56538;
  assign n56540 = ~n44387 & ~n56539;
  assign n56541 = ~i_hbusreq5 & ~n56540;
  assign n56542 = ~n56532 & ~n56541;
  assign n56543 = ~controllable_hgrant5 & ~n56542;
  assign n56544 = ~n44376 & ~n56543;
  assign n56545 = ~controllable_hmaster2 & ~n56544;
  assign n56546 = ~n56479 & ~n56545;
  assign n56547 = ~controllable_hmaster1 & ~n56546;
  assign n56548 = ~n56478 & ~n56547;
  assign n56549 = ~i_hbusreq6 & ~n56548;
  assign n56550 = ~n56531 & ~n56549;
  assign n56551 = ~controllable_hgrant6 & ~n56550;
  assign n56552 = ~n44368 & ~n56551;
  assign n56553 = ~controllable_hmaster0 & ~n56552;
  assign n56554 = ~n56530 & ~n56553;
  assign n56555 = i_hlock8 & ~n56554;
  assign n56556 = i_hbusreq6 & ~n56295;
  assign n56557 = i_hbusreq5 & ~n56289;
  assign n56558 = i_hbusreq4 & ~n56261;
  assign n56559 = i_hbusreq9 & ~n56261;
  assign n56560 = ~i_hbusreq9 & ~n56509;
  assign n56561 = ~n56559 & ~n56560;
  assign n56562 = ~i_hbusreq4 & ~n56561;
  assign n56563 = ~n56558 & ~n56562;
  assign n56564 = ~controllable_hgrant4 & ~n56563;
  assign n56565 = ~n44467 & ~n56564;
  assign n56566 = ~i_hbusreq5 & ~n56565;
  assign n56567 = ~n56557 & ~n56566;
  assign n56568 = ~controllable_hgrant5 & ~n56567;
  assign n56569 = ~n44456 & ~n56568;
  assign n56570 = ~controllable_hmaster2 & ~n56569;
  assign n56571 = ~n56479 & ~n56570;
  assign n56572 = ~controllable_hmaster1 & ~n56571;
  assign n56573 = ~n56478 & ~n56572;
  assign n56574 = ~i_hbusreq6 & ~n56573;
  assign n56575 = ~n56556 & ~n56574;
  assign n56576 = ~controllable_hgrant6 & ~n56575;
  assign n56577 = ~n44448 & ~n56576;
  assign n56578 = ~controllable_hmaster0 & ~n56577;
  assign n56579 = ~n56530 & ~n56578;
  assign n56580 = ~i_hlock8 & ~n56579;
  assign n56581 = ~n56555 & ~n56580;
  assign n56582 = ~i_hbusreq8 & ~n56581;
  assign n56583 = ~n56429 & ~n56582;
  assign n56584 = controllable_hmaster3 & ~n56583;
  assign n56585 = i_hbusreq8 & ~n56413;
  assign n56586 = i_hbusreq6 & ~n56336;
  assign n56587 = controllable_hmaster2 & ~n56544;
  assign n56588 = i_hbusreq5 & ~n56310;
  assign n56589 = i_hbusreq4 & ~n56308;
  assign n56590 = i_hbusreq9 & ~n56308;
  assign n56591 = i_hbusreq3 & ~n56306;
  assign n56592 = i_hlock3 & ~n56493;
  assign n56593 = ~i_hlock3 & ~n56505;
  assign n56594 = ~n56592 & ~n56593;
  assign n56595 = ~i_hbusreq3 & ~n56594;
  assign n56596 = ~n56591 & ~n56595;
  assign n56597 = ~controllable_hgrant3 & ~n56596;
  assign n56598 = ~n44562 & ~n56597;
  assign n56599 = ~i_hbusreq9 & ~n56598;
  assign n56600 = ~n56590 & ~n56599;
  assign n56601 = ~i_hbusreq4 & ~n56600;
  assign n56602 = ~n56589 & ~n56601;
  assign n56603 = ~controllable_hgrant4 & ~n56602;
  assign n56604 = ~n44547 & ~n56603;
  assign n56605 = ~i_hbusreq5 & ~n56604;
  assign n56606 = ~n56588 & ~n56605;
  assign n56607 = ~controllable_hgrant5 & ~n56606;
  assign n56608 = ~n44536 & ~n56607;
  assign n56609 = ~controllable_hmaster2 & ~n56608;
  assign n56610 = ~n56587 & ~n56609;
  assign n56611 = controllable_hmaster1 & ~n56610;
  assign n56612 = i_hbusreq5 & ~n56318;
  assign n56613 = i_hlock5 & ~n56540;
  assign n56614 = ~i_hlock5 & ~n56565;
  assign n56615 = ~n56613 & ~n56614;
  assign n56616 = ~i_hbusreq5 & ~n56615;
  assign n56617 = ~n56612 & ~n56616;
  assign n56618 = ~controllable_hgrant5 & ~n56617;
  assign n56619 = ~n44596 & ~n56618;
  assign n56620 = controllable_hmaster2 & ~n56619;
  assign n56621 = i_hbusreq5 & ~n56330;
  assign n56622 = i_hbusreq4 & ~n56328;
  assign n56623 = i_hbusreq9 & ~n56328;
  assign n56624 = i_hbusreq3 & ~n56326;
  assign n56625 = i_hbusreq1 & ~n56324;
  assign n56626 = i_hlock1 & ~n56489;
  assign n56627 = ~i_hlock1 & ~n56501;
  assign n56628 = ~n56626 & ~n56627;
  assign n56629 = ~i_hbusreq1 & ~n56628;
  assign n56630 = ~n56625 & ~n56629;
  assign n56631 = ~controllable_hgrant1 & ~n56630;
  assign n56632 = ~n44646 & ~n56631;
  assign n56633 = ~i_hbusreq3 & ~n56632;
  assign n56634 = ~n56624 & ~n56633;
  assign n56635 = ~controllable_hgrant3 & ~n56634;
  assign n56636 = ~n44632 & ~n56635;
  assign n56637 = ~i_hbusreq9 & ~n56636;
  assign n56638 = ~n56623 & ~n56637;
  assign n56639 = ~i_hbusreq4 & ~n56638;
  assign n56640 = ~n56622 & ~n56639;
  assign n56641 = ~controllable_hgrant4 & ~n56640;
  assign n56642 = ~n44623 & ~n56641;
  assign n56643 = ~i_hbusreq5 & ~n56642;
  assign n56644 = ~n56621 & ~n56643;
  assign n56645 = ~controllable_hgrant5 & ~n56644;
  assign n56646 = ~n44612 & ~n56645;
  assign n56647 = ~controllable_hmaster2 & ~n56646;
  assign n56648 = ~n56620 & ~n56647;
  assign n56649 = ~controllable_hmaster1 & ~n56648;
  assign n56650 = ~n56611 & ~n56649;
  assign n56651 = ~i_hbusreq6 & ~n56650;
  assign n56652 = ~n56586 & ~n56651;
  assign n56653 = ~controllable_hgrant6 & ~n56652;
  assign n56654 = ~n44527 & ~n56653;
  assign n56655 = controllable_hmaster0 & ~n56654;
  assign n56656 = i_hbusreq6 & ~n56352;
  assign n56657 = ~n15602 & ~n27343;
  assign n56658 = controllable_hmaster1 & ~n56657;
  assign n56659 = ~n14668 & ~n56658;
  assign n56660 = n8217 & ~n56659;
  assign n56661 = ~n23260 & ~n29947;
  assign n56662 = controllable_hmaster1 & ~n56661;
  assign n56663 = ~n20219 & ~n56662;
  assign n56664 = ~n8217 & ~n56663;
  assign n56665 = ~n56660 & ~n56664;
  assign n56666 = i_hlock6 & ~n56665;
  assign n56667 = ~n15602 & ~n27370;
  assign n56668 = controllable_hmaster1 & ~n56667;
  assign n56669 = ~n14668 & ~n56668;
  assign n56670 = n8217 & ~n56669;
  assign n56671 = ~n23260 & ~n29977;
  assign n56672 = controllable_hmaster1 & ~n56671;
  assign n56673 = ~n20219 & ~n56672;
  assign n56674 = ~n8217 & ~n56673;
  assign n56675 = ~n56670 & ~n56674;
  assign n56676 = ~i_hlock6 & ~n56675;
  assign n56677 = ~n56666 & ~n56676;
  assign n56678 = ~i_hbusreq6 & ~n56677;
  assign n56679 = ~n56656 & ~n56678;
  assign n56680 = controllable_hgrant6 & ~n56679;
  assign n56681 = i_hbusreq6 & ~n56409;
  assign n56682 = i_hbusreq5 & ~n56355;
  assign n56683 = n8378 & ~n15597;
  assign n56684 = ~n8378 & ~n23255;
  assign n56685 = ~n56683 & ~n56684;
  assign n56686 = ~i_hbusreq5 & ~n56685;
  assign n56687 = ~n56682 & ~n56686;
  assign n56688 = controllable_hgrant5 & ~n56687;
  assign n56689 = i_hbusreq5 & ~n56376;
  assign n56690 = i_hbusreq4 & ~n56358;
  assign n56691 = i_hbusreq9 & ~n56358;
  assign n56692 = n8426 & ~n15591;
  assign n56693 = ~n8426 & ~n23249;
  assign n56694 = ~n56692 & ~n56693;
  assign n56695 = ~i_hbusreq9 & ~n56694;
  assign n56696 = ~n56691 & ~n56695;
  assign n56697 = ~i_hbusreq4 & ~n56696;
  assign n56698 = ~n56690 & ~n56697;
  assign n56699 = controllable_hgrant4 & ~n56698;
  assign n56700 = i_hbusreq4 & ~n56374;
  assign n56701 = i_hbusreq9 & ~n56374;
  assign n56702 = i_hbusreq3 & ~n56361;
  assign n56703 = n8365 & ~n15587;
  assign n56704 = ~n8365 & ~n23245;
  assign n56705 = ~n56703 & ~n56704;
  assign n56706 = ~i_hbusreq3 & ~n56705;
  assign n56707 = ~n56702 & ~n56706;
  assign n56708 = controllable_hgrant3 & ~n56707;
  assign n56709 = i_hbusreq3 & ~n56372;
  assign n56710 = i_hbusreq1 & ~n56364;
  assign n56711 = n8389 & ~n15583;
  assign n56712 = ~n8389 & ~n23241;
  assign n56713 = ~n56711 & ~n56712;
  assign n56714 = ~i_hbusreq1 & ~n56713;
  assign n56715 = ~n56710 & ~n56714;
  assign n56716 = controllable_hgrant1 & ~n56715;
  assign n56717 = i_hbusreq1 & ~n56370;
  assign n56718 = ~n44275 & ~n44750;
  assign n56719 = ~n7733 & ~n56718;
  assign n56720 = ~n44301 & ~n49770;
  assign n56721 = n7733 & ~n56720;
  assign n56722 = ~n56719 & ~n56721;
  assign n56723 = n7928 & ~n56722;
  assign n56724 = ~n43545 & ~n56723;
  assign n56725 = ~i_hbusreq1 & ~n56724;
  assign n56726 = ~n56717 & ~n56725;
  assign n56727 = ~controllable_hgrant1 & ~n56726;
  assign n56728 = ~n56716 & ~n56727;
  assign n56729 = ~i_hbusreq3 & ~n56728;
  assign n56730 = ~n56709 & ~n56729;
  assign n56731 = ~controllable_hgrant3 & ~n56730;
  assign n56732 = ~n56708 & ~n56731;
  assign n56733 = ~i_hbusreq9 & ~n56732;
  assign n56734 = ~n56701 & ~n56733;
  assign n56735 = ~i_hbusreq4 & ~n56734;
  assign n56736 = ~n56700 & ~n56735;
  assign n56737 = ~controllable_hgrant4 & ~n56736;
  assign n56738 = ~n56699 & ~n56737;
  assign n56739 = ~i_hbusreq5 & ~n56738;
  assign n56740 = ~n56689 & ~n56739;
  assign n56741 = ~controllable_hgrant5 & ~n56740;
  assign n56742 = ~n56688 & ~n56741;
  assign n56743 = ~controllable_hmaster2 & ~n56742;
  assign n56744 = ~n56587 & ~n56743;
  assign n56745 = controllable_hmaster1 & ~n56744;
  assign n56746 = i_hbusreq5 & ~n56386;
  assign n56747 = i_hbusreq4 & ~n56384;
  assign n56748 = i_hlock4 & ~n56536;
  assign n56749 = ~i_hlock4 & ~n56561;
  assign n56750 = ~n56748 & ~n56749;
  assign n56751 = ~i_hbusreq4 & ~n56750;
  assign n56752 = ~n56747 & ~n56751;
  assign n56753 = ~controllable_hgrant4 & ~n56752;
  assign n56754 = ~n44805 & ~n56753;
  assign n56755 = ~i_hbusreq5 & ~n56754;
  assign n56756 = ~n56746 & ~n56755;
  assign n56757 = ~controllable_hgrant5 & ~n56756;
  assign n56758 = ~n44785 & ~n56757;
  assign n56759 = controllable_hmaster2 & ~n56758;
  assign n56760 = i_hbusreq5 & ~n56396;
  assign n56761 = i_hbusreq4 & ~n56394;
  assign n56762 = i_hbusreq9 & ~n56394;
  assign n56763 = i_hbusreq3 & ~n56392;
  assign n56764 = i_hbusreq1 & ~n56390;
  assign n56765 = ~n39848 & ~n46054;
  assign n56766 = controllable_locked & ~n56765;
  assign n56767 = ~controllable_hmastlock & ~n49180;
  assign n56768 = ~n42945 & ~n56767;
  assign n56769 = ~controllable_locked & ~n56768;
  assign n56770 = ~n56766 & ~n56769;
  assign n56771 = i_hlock0 & ~n56770;
  assign n56772 = ~n46695 & ~n56771;
  assign n56773 = ~i_hbusreq0 & ~n56772;
  assign n56774 = ~n46689 & ~n56773;
  assign n56775 = i_hlock2 & ~n56774;
  assign n56776 = ~n46700 & ~n56773;
  assign n56777 = ~i_hlock2 & ~n56776;
  assign n56778 = ~n56775 & ~n56777;
  assign n56779 = ~i_hbusreq2 & ~n56778;
  assign n56780 = ~n46688 & ~n56779;
  assign n56781 = controllable_hgrant2 & ~n56780;
  assign n56782 = ~n19070 & ~n56781;
  assign n56783 = n7733 & ~n56782;
  assign n56784 = ~n44867 & ~n56783;
  assign n56785 = n7928 & ~n56784;
  assign n56786 = ~n8440 & ~n56785;
  assign n56787 = ~i_hbusreq1 & ~n56786;
  assign n56788 = ~n56764 & ~n56787;
  assign n56789 = ~controllable_hgrant1 & ~n56788;
  assign n56790 = ~n44853 & ~n56789;
  assign n56791 = ~i_hbusreq3 & ~n56790;
  assign n56792 = ~n56763 & ~n56791;
  assign n56793 = ~controllable_hgrant3 & ~n56792;
  assign n56794 = ~n44845 & ~n56793;
  assign n56795 = ~i_hbusreq9 & ~n56794;
  assign n56796 = ~n56762 & ~n56795;
  assign n56797 = ~i_hbusreq4 & ~n56796;
  assign n56798 = ~n56761 & ~n56797;
  assign n56799 = ~controllable_hgrant4 & ~n56798;
  assign n56800 = ~n44836 & ~n56799;
  assign n56801 = ~i_hbusreq5 & ~n56800;
  assign n56802 = ~n56760 & ~n56801;
  assign n56803 = ~controllable_hgrant5 & ~n56802;
  assign n56804 = ~n44825 & ~n56803;
  assign n56805 = ~controllable_hmaster2 & ~n56804;
  assign n56806 = ~n56759 & ~n56805;
  assign n56807 = ~controllable_hmaster1 & ~n56806;
  assign n56808 = ~n56745 & ~n56807;
  assign n56809 = i_hlock6 & ~n56808;
  assign n56810 = controllable_hmaster2 & ~n56569;
  assign n56811 = ~n56743 & ~n56810;
  assign n56812 = controllable_hmaster1 & ~n56811;
  assign n56813 = ~n56807 & ~n56812;
  assign n56814 = ~i_hlock6 & ~n56813;
  assign n56815 = ~n56809 & ~n56814;
  assign n56816 = ~i_hbusreq6 & ~n56815;
  assign n56817 = ~n56681 & ~n56816;
  assign n56818 = ~controllable_hgrant6 & ~n56817;
  assign n56819 = ~n56680 & ~n56818;
  assign n56820 = ~controllable_hmaster0 & ~n56819;
  assign n56821 = ~n56655 & ~n56820;
  assign n56822 = ~i_hbusreq8 & ~n56821;
  assign n56823 = ~n56585 & ~n56822;
  assign n56824 = ~controllable_hmaster3 & ~n56823;
  assign n56825 = ~n56584 & ~n56824;
  assign n56826 = i_hlock7 & ~n56825;
  assign n56827 = i_hbusreq8 & ~n56423;
  assign n56828 = i_hbusreq6 & ~n56419;
  assign n56829 = ~n56609 & ~n56810;
  assign n56830 = controllable_hmaster1 & ~n56829;
  assign n56831 = ~n56649 & ~n56830;
  assign n56832 = ~i_hbusreq6 & ~n56831;
  assign n56833 = ~n56828 & ~n56832;
  assign n56834 = ~controllable_hgrant6 & ~n56833;
  assign n56835 = ~n44920 & ~n56834;
  assign n56836 = controllable_hmaster0 & ~n56835;
  assign n56837 = ~n56820 & ~n56836;
  assign n56838 = ~i_hbusreq8 & ~n56837;
  assign n56839 = ~n56827 & ~n56838;
  assign n56840 = ~controllable_hmaster3 & ~n56839;
  assign n56841 = ~n56584 & ~n56840;
  assign n56842 = ~i_hlock7 & ~n56841;
  assign n56843 = ~n56826 & ~n56842;
  assign n56844 = ~i_hbusreq7 & ~n56843;
  assign n56845 = ~n56428 & ~n56844;
  assign n56846 = n7924 & ~n56845;
  assign n56847 = ~n56231 & ~n56846;
  assign n56848 = n8214 & ~n56847;
  assign n56849 = ~n55702 & ~n56848;
  assign n56850 = n8202 & ~n56849;
  assign n56851 = ~n54815 & ~n56850;
  assign n56852 = n7920 & ~n56851;
  assign n56853 = ~n50812 & ~n56852;
  assign n56854 = ~n7728 & ~n56853;
  assign n56855 = ~n53432 & ~n56854;
  assign n56856 = n7723 & ~n56855;
  assign n56857 = ~n7723 & ~n56853;
  assign n56858 = ~n56856 & ~n56857;
  assign n56859 = n7714 & ~n56858;
  assign n56860 = n7723 & ~n56853;
  assign n56861 = ~n46001 & ~n48769;
  assign n56862 = controllable_hmaster1 & ~n56861;
  assign n56863 = controllable_hmaster2 & ~n56861;
  assign n56864 = ~n46012 & ~n47504;
  assign n56865 = ~controllable_hmaster2 & ~n56864;
  assign n56866 = ~n56863 & ~n56865;
  assign n56867 = ~controllable_hmaster1 & ~n56866;
  assign n56868 = ~n56862 & ~n56867;
  assign n56869 = ~controllable_hgrant6 & ~n56868;
  assign n56870 = ~n47480 & ~n56869;
  assign n56871 = controllable_hmaster0 & ~n56870;
  assign n56872 = ~n46155 & ~n47528;
  assign n56873 = ~controllable_hmaster2 & ~n56872;
  assign n56874 = ~n56863 & ~n56873;
  assign n56875 = ~controllable_hmaster1 & ~n56874;
  assign n56876 = ~n56862 & ~n56875;
  assign n56877 = ~controllable_hgrant6 & ~n56876;
  assign n56878 = ~n46111 & ~n56877;
  assign n56879 = ~controllable_hmaster0 & ~n56878;
  assign n56880 = ~n56871 & ~n56879;
  assign n56881 = i_hlock8 & ~n56880;
  assign n56882 = ~n46213 & ~n47561;
  assign n56883 = ~controllable_hmaster2 & ~n56882;
  assign n56884 = ~n56863 & ~n56883;
  assign n56885 = ~controllable_hmaster1 & ~n56884;
  assign n56886 = ~n56862 & ~n56885;
  assign n56887 = ~controllable_hgrant6 & ~n56886;
  assign n56888 = ~n46173 & ~n56887;
  assign n56889 = ~controllable_hmaster0 & ~n56888;
  assign n56890 = ~n56871 & ~n56889;
  assign n56891 = ~i_hlock8 & ~n56890;
  assign n56892 = ~n56881 & ~n56891;
  assign n56893 = controllable_hmaster3 & ~n56892;
  assign n56894 = ~n8217 & ~n38078;
  assign n56895 = ~n43905 & ~n56894;
  assign n56896 = i_hlock6 & ~n56895;
  assign n56897 = ~n8217 & ~n38084;
  assign n56898 = ~n43905 & ~n56897;
  assign n56899 = ~i_hlock6 & ~n56898;
  assign n56900 = ~n56896 & ~n56899;
  assign n56901 = controllable_hgrant6 & ~n56900;
  assign n56902 = controllable_hmaster2 & ~n56872;
  assign n56903 = ~n46266 & ~n48843;
  assign n56904 = ~controllable_hmaster2 & ~n56903;
  assign n56905 = ~n56902 & ~n56904;
  assign n56906 = controllable_hmaster1 & ~n56905;
  assign n56907 = ~n46326 & ~n48893;
  assign n56908 = ~controllable_hmaster2 & ~n56907;
  assign n56909 = ~n48885 & ~n56908;
  assign n56910 = ~controllable_hmaster1 & ~n56909;
  assign n56911 = ~n56906 & ~n56910;
  assign n56912 = ~controllable_hgrant6 & ~n56911;
  assign n56913 = ~n56901 & ~n56912;
  assign n56914 = controllable_hmaster0 & ~n56913;
  assign n56915 = ~n46404 & ~n48943;
  assign n56916 = ~controllable_hmaster2 & ~n56915;
  assign n56917 = ~n56902 & ~n56916;
  assign n56918 = controllable_hmaster1 & ~n56917;
  assign n56919 = ~n46430 & ~n49001;
  assign n56920 = controllable_hmaster2 & ~n56919;
  assign n56921 = ~n46472 & ~n49025;
  assign n56922 = ~controllable_hmaster2 & ~n56921;
  assign n56923 = ~n56920 & ~n56922;
  assign n56924 = ~controllable_hmaster1 & ~n56923;
  assign n56925 = ~n56918 & ~n56924;
  assign n56926 = i_hlock6 & ~n56925;
  assign n56927 = controllable_hmaster2 & ~n56882;
  assign n56928 = ~n56916 & ~n56927;
  assign n56929 = controllable_hmaster1 & ~n56928;
  assign n56930 = ~n56924 & ~n56929;
  assign n56931 = ~i_hlock6 & ~n56930;
  assign n56932 = ~n56926 & ~n56931;
  assign n56933 = ~controllable_hgrant6 & ~n56932;
  assign n56934 = ~n46348 & ~n56933;
  assign n56935 = ~controllable_hmaster0 & ~n56934;
  assign n56936 = ~n56914 & ~n56935;
  assign n56937 = ~controllable_hmaster3 & ~n56936;
  assign n56938 = ~n56893 & ~n56937;
  assign n56939 = i_hlock7 & ~n56938;
  assign n56940 = ~n8217 & ~n38094;
  assign n56941 = ~n44119 & ~n56940;
  assign n56942 = i_hlock6 & ~n56941;
  assign n56943 = ~n8217 & ~n38100;
  assign n56944 = ~n44119 & ~n56943;
  assign n56945 = ~i_hlock6 & ~n56944;
  assign n56946 = ~n56942 & ~n56945;
  assign n56947 = controllable_hgrant6 & ~n56946;
  assign n56948 = ~n56904 & ~n56927;
  assign n56949 = controllable_hmaster1 & ~n56948;
  assign n56950 = ~n56910 & ~n56949;
  assign n56951 = ~controllable_hgrant6 & ~n56950;
  assign n56952 = ~n56947 & ~n56951;
  assign n56953 = controllable_hmaster0 & ~n56952;
  assign n56954 = ~n56935 & ~n56953;
  assign n56955 = ~controllable_hmaster3 & ~n56954;
  assign n56956 = ~n56893 & ~n56955;
  assign n56957 = ~i_hlock7 & ~n56956;
  assign n56958 = ~n56939 & ~n56957;
  assign n56959 = i_hbusreq7 & ~n56958;
  assign n56960 = i_hbusreq8 & ~n56892;
  assign n56961 = i_hbusreq6 & ~n56868;
  assign n56962 = ~n46619 & ~n53800;
  assign n56963 = controllable_hmaster1 & ~n56962;
  assign n56964 = controllable_hmaster2 & ~n56962;
  assign n56965 = ~n47644 & ~n53814;
  assign n56966 = ~controllable_hmaster2 & ~n56965;
  assign n56967 = ~n56964 & ~n56966;
  assign n56968 = ~controllable_hmaster1 & ~n56967;
  assign n56969 = ~n56963 & ~n56968;
  assign n56970 = ~i_hbusreq6 & ~n56969;
  assign n56971 = ~n56961 & ~n56970;
  assign n56972 = ~controllable_hgrant6 & ~n56971;
  assign n56973 = ~n47598 & ~n56972;
  assign n56974 = controllable_hmaster0 & ~n56973;
  assign n56975 = i_hbusreq6 & ~n56876;
  assign n56976 = ~n46870 & ~n53836;
  assign n56977 = ~controllable_hmaster2 & ~n56976;
  assign n56978 = ~n56964 & ~n56977;
  assign n56979 = ~controllable_hmaster1 & ~n56978;
  assign n56980 = ~n56963 & ~n56979;
  assign n56981 = ~i_hbusreq6 & ~n56980;
  assign n56982 = ~n56975 & ~n56981;
  assign n56983 = ~controllable_hgrant6 & ~n56982;
  assign n56984 = ~n46792 & ~n56983;
  assign n56985 = ~controllable_hmaster0 & ~n56984;
  assign n56986 = ~n56974 & ~n56985;
  assign n56987 = i_hlock8 & ~n56986;
  assign n56988 = i_hbusreq6 & ~n56886;
  assign n56989 = ~n46967 & ~n53860;
  assign n56990 = ~controllable_hmaster2 & ~n56989;
  assign n56991 = ~n56964 & ~n56990;
  assign n56992 = ~controllable_hmaster1 & ~n56991;
  assign n56993 = ~n56963 & ~n56992;
  assign n56994 = ~i_hbusreq6 & ~n56993;
  assign n56995 = ~n56988 & ~n56994;
  assign n56996 = ~controllable_hgrant6 & ~n56995;
  assign n56997 = ~n46893 & ~n56996;
  assign n56998 = ~controllable_hmaster0 & ~n56997;
  assign n56999 = ~n56974 & ~n56998;
  assign n57000 = ~i_hlock8 & ~n56999;
  assign n57001 = ~n56987 & ~n57000;
  assign n57002 = ~i_hbusreq8 & ~n57001;
  assign n57003 = ~n56960 & ~n57002;
  assign n57004 = controllable_hmaster3 & ~n57003;
  assign n57005 = i_hbusreq8 & ~n56936;
  assign n57006 = i_hbusreq6 & ~n56900;
  assign n57007 = ~n8217 & ~n38114;
  assign n57008 = ~n53879 & ~n57007;
  assign n57009 = i_hlock6 & ~n57008;
  assign n57010 = ~n8217 & ~n38123;
  assign n57011 = ~n53879 & ~n57010;
  assign n57012 = ~i_hlock6 & ~n57011;
  assign n57013 = ~n57009 & ~n57012;
  assign n57014 = ~i_hbusreq6 & ~n57013;
  assign n57015 = ~n57006 & ~n57014;
  assign n57016 = controllable_hgrant6 & ~n57015;
  assign n57017 = i_hbusreq6 & ~n56911;
  assign n57018 = controllable_hmaster2 & ~n56976;
  assign n57019 = ~n47056 & ~n53897;
  assign n57020 = ~controllable_hmaster2 & ~n57019;
  assign n57021 = ~n57018 & ~n57020;
  assign n57022 = controllable_hmaster1 & ~n57021;
  assign n57023 = i_hlock5 & ~n47699;
  assign n57024 = ~i_hlock5 & ~n47759;
  assign n57025 = ~n57023 & ~n57024;
  assign n57026 = ~i_hbusreq5 & ~n57025;
  assign n57027 = ~n49569 & ~n57026;
  assign n57028 = ~controllable_hgrant5 & ~n57027;
  assign n57029 = ~n49568 & ~n57028;
  assign n57030 = controllable_hmaster2 & ~n57029;
  assign n57031 = ~n47155 & ~n53921;
  assign n57032 = ~controllable_hmaster2 & ~n57031;
  assign n57033 = ~n57030 & ~n57032;
  assign n57034 = ~controllable_hmaster1 & ~n57033;
  assign n57035 = ~n57022 & ~n57034;
  assign n57036 = ~i_hbusreq6 & ~n57035;
  assign n57037 = ~n57017 & ~n57036;
  assign n57038 = ~controllable_hgrant6 & ~n57037;
  assign n57039 = ~n57016 & ~n57038;
  assign n57040 = controllable_hmaster0 & ~n57039;
  assign n57041 = i_hbusreq6 & ~n56932;
  assign n57042 = ~n47279 & ~n53943;
  assign n57043 = ~controllable_hmaster2 & ~n57042;
  assign n57044 = ~n57018 & ~n57043;
  assign n57045 = controllable_hmaster1 & ~n57044;
  assign n57046 = ~n47323 & ~n53958;
  assign n57047 = controllable_hmaster2 & ~n57046;
  assign n57048 = ~n47416 & ~n53971;
  assign n57049 = ~controllable_hmaster2 & ~n57048;
  assign n57050 = ~n57047 & ~n57049;
  assign n57051 = ~controllable_hmaster1 & ~n57050;
  assign n57052 = ~n57045 & ~n57051;
  assign n57053 = i_hlock6 & ~n57052;
  assign n57054 = controllable_hmaster2 & ~n56989;
  assign n57055 = ~n57043 & ~n57054;
  assign n57056 = controllable_hmaster1 & ~n57055;
  assign n57057 = ~n57051 & ~n57056;
  assign n57058 = ~i_hlock6 & ~n57057;
  assign n57059 = ~n57053 & ~n57058;
  assign n57060 = ~i_hbusreq6 & ~n57059;
  assign n57061 = ~n57041 & ~n57060;
  assign n57062 = ~controllable_hgrant6 & ~n57061;
  assign n57063 = ~n47182 & ~n57062;
  assign n57064 = ~controllable_hmaster0 & ~n57063;
  assign n57065 = ~n57040 & ~n57064;
  assign n57066 = ~i_hbusreq8 & ~n57065;
  assign n57067 = ~n57005 & ~n57066;
  assign n57068 = ~controllable_hmaster3 & ~n57067;
  assign n57069 = ~n57004 & ~n57068;
  assign n57070 = i_hlock7 & ~n57069;
  assign n57071 = i_hbusreq8 & ~n56954;
  assign n57072 = i_hbusreq6 & ~n56946;
  assign n57073 = ~n8217 & ~n38139;
  assign n57074 = ~n53997 & ~n57073;
  assign n57075 = i_hlock6 & ~n57074;
  assign n57076 = ~n8217 & ~n38148;
  assign n57077 = ~n53997 & ~n57076;
  assign n57078 = ~i_hlock6 & ~n57077;
  assign n57079 = ~n57075 & ~n57078;
  assign n57080 = ~i_hbusreq6 & ~n57079;
  assign n57081 = ~n57072 & ~n57080;
  assign n57082 = controllable_hgrant6 & ~n57081;
  assign n57083 = i_hbusreq6 & ~n56950;
  assign n57084 = ~n57020 & ~n57054;
  assign n57085 = controllable_hmaster1 & ~n57084;
  assign n57086 = ~n57034 & ~n57085;
  assign n57087 = ~i_hbusreq6 & ~n57086;
  assign n57088 = ~n57083 & ~n57087;
  assign n57089 = ~controllable_hgrant6 & ~n57088;
  assign n57090 = ~n57082 & ~n57089;
  assign n57091 = controllable_hmaster0 & ~n57090;
  assign n57092 = ~n57064 & ~n57091;
  assign n57093 = ~i_hbusreq8 & ~n57092;
  assign n57094 = ~n57071 & ~n57093;
  assign n57095 = ~controllable_hmaster3 & ~n57094;
  assign n57096 = ~n57004 & ~n57095;
  assign n57097 = ~i_hlock7 & ~n57096;
  assign n57098 = ~n57070 & ~n57097;
  assign n57099 = ~i_hbusreq7 & ~n57098;
  assign n57100 = ~n56959 & ~n57099;
  assign n57101 = n7924 & ~n57100;
  assign n57102 = ~n53692 & ~n57101;
  assign n57103 = ~n8214 & ~n57102;
  assign n57104 = ~n45999 & ~n48777;
  assign n57105 = ~controllable_hgrant5 & ~n57104;
  assign n57106 = ~n45950 & ~n57105;
  assign n57107 = controllable_hmaster1 & ~n57106;
  assign n57108 = controllable_hmaster2 & ~n57106;
  assign n57109 = ~n46030 & ~n47502;
  assign n57110 = ~controllable_hgrant5 & ~n57109;
  assign n57111 = ~n47488 & ~n57110;
  assign n57112 = ~controllable_hmaster2 & ~n57111;
  assign n57113 = ~n57108 & ~n57112;
  assign n57114 = ~controllable_hmaster1 & ~n57113;
  assign n57115 = ~n57107 & ~n57114;
  assign n57116 = ~controllable_hgrant6 & ~n57115;
  assign n57117 = ~n47480 & ~n57116;
  assign n57118 = controllable_hmaster0 & ~n57117;
  assign n57119 = ~n46153 & ~n47532;
  assign n57120 = ~controllable_hgrant5 & ~n57119;
  assign n57121 = ~n46119 & ~n57120;
  assign n57122 = ~controllable_hmaster2 & ~n57121;
  assign n57123 = ~n57108 & ~n57122;
  assign n57124 = ~controllable_hmaster1 & ~n57123;
  assign n57125 = ~n57107 & ~n57124;
  assign n57126 = ~controllable_hgrant6 & ~n57125;
  assign n57127 = ~n46111 & ~n57126;
  assign n57128 = ~controllable_hmaster0 & ~n57127;
  assign n57129 = ~n57118 & ~n57128;
  assign n57130 = i_hlock8 & ~n57129;
  assign n57131 = ~n46211 & ~n47565;
  assign n57132 = ~controllable_hgrant5 & ~n57131;
  assign n57133 = ~n46181 & ~n57132;
  assign n57134 = ~controllable_hmaster2 & ~n57133;
  assign n57135 = ~n57108 & ~n57134;
  assign n57136 = ~controllable_hmaster1 & ~n57135;
  assign n57137 = ~n57107 & ~n57136;
  assign n57138 = ~controllable_hgrant6 & ~n57137;
  assign n57139 = ~n46173 & ~n57138;
  assign n57140 = ~controllable_hmaster0 & ~n57139;
  assign n57141 = ~n57118 & ~n57140;
  assign n57142 = ~i_hlock8 & ~n57141;
  assign n57143 = ~n57130 & ~n57142;
  assign n57144 = controllable_hmaster3 & ~n57143;
  assign n57145 = controllable_hmaster2 & ~n57121;
  assign n57146 = ~n46264 & ~n48851;
  assign n57147 = ~controllable_hgrant5 & ~n57146;
  assign n57148 = ~n46242 & ~n57147;
  assign n57149 = ~controllable_hmaster2 & ~n57148;
  assign n57150 = ~n57145 & ~n57149;
  assign n57151 = controllable_hmaster1 & ~n57150;
  assign n57152 = i_hlock5 & ~n57119;
  assign n57153 = ~i_hlock5 & ~n57131;
  assign n57154 = ~n57152 & ~n57153;
  assign n57155 = ~controllable_hgrant5 & ~n57154;
  assign n57156 = ~n46278 & ~n57155;
  assign n57157 = controllable_hmaster2 & ~n57156;
  assign n57158 = ~n46324 & ~n48901;
  assign n57159 = ~controllable_hgrant5 & ~n57158;
  assign n57160 = ~n46292 & ~n57159;
  assign n57161 = ~controllable_hmaster2 & ~n57160;
  assign n57162 = ~n57157 & ~n57161;
  assign n57163 = ~controllable_hmaster1 & ~n57162;
  assign n57164 = ~n57151 & ~n57163;
  assign n57165 = ~controllable_hgrant6 & ~n57164;
  assign n57166 = ~n46233 & ~n57165;
  assign n57167 = controllable_hmaster0 & ~n57166;
  assign n57168 = ~n33019 & ~n46336;
  assign n57169 = ~n8217 & ~n57168;
  assign n57170 = ~n43999 & ~n57169;
  assign n57171 = i_hlock6 & ~n57170;
  assign n57172 = ~n33033 & ~n46342;
  assign n57173 = ~n8217 & ~n57172;
  assign n57174 = ~n44009 & ~n57173;
  assign n57175 = ~i_hlock6 & ~n57174;
  assign n57176 = ~n57171 & ~n57175;
  assign n57177 = controllable_hgrant6 & ~n57176;
  assign n57178 = ~n46402 & ~n48951;
  assign n57179 = ~controllable_hgrant5 & ~n57178;
  assign n57180 = ~n46356 & ~n57179;
  assign n57181 = ~controllable_hmaster2 & ~n57180;
  assign n57182 = ~n57145 & ~n57181;
  assign n57183 = controllable_hmaster1 & ~n57182;
  assign n57184 = ~n46470 & ~n49033;
  assign n57185 = ~controllable_hgrant5 & ~n57184;
  assign n57186 = ~n46440 & ~n57185;
  assign n57187 = ~controllable_hmaster2 & ~n57186;
  assign n57188 = ~n49017 & ~n57187;
  assign n57189 = ~controllable_hmaster1 & ~n57188;
  assign n57190 = ~n57183 & ~n57189;
  assign n57191 = i_hlock6 & ~n57190;
  assign n57192 = controllable_hmaster2 & ~n57133;
  assign n57193 = ~n57181 & ~n57192;
  assign n57194 = controllable_hmaster1 & ~n57193;
  assign n57195 = ~n57189 & ~n57194;
  assign n57196 = ~i_hlock6 & ~n57195;
  assign n57197 = ~n57191 & ~n57196;
  assign n57198 = ~controllable_hgrant6 & ~n57197;
  assign n57199 = ~n57177 & ~n57198;
  assign n57200 = ~controllable_hmaster0 & ~n57199;
  assign n57201 = ~n57167 & ~n57200;
  assign n57202 = ~controllable_hmaster3 & ~n57201;
  assign n57203 = ~n57144 & ~n57202;
  assign n57204 = i_hlock7 & ~n57203;
  assign n57205 = ~n57149 & ~n57192;
  assign n57206 = controllable_hmaster1 & ~n57205;
  assign n57207 = ~n57163 & ~n57206;
  assign n57208 = ~controllable_hgrant6 & ~n57207;
  assign n57209 = ~n46499 & ~n57208;
  assign n57210 = controllable_hmaster0 & ~n57209;
  assign n57211 = ~n57200 & ~n57210;
  assign n57212 = ~controllable_hmaster3 & ~n57211;
  assign n57213 = ~n57144 & ~n57212;
  assign n57214 = ~i_hlock7 & ~n57213;
  assign n57215 = ~n57204 & ~n57214;
  assign n57216 = i_hbusreq7 & ~n57215;
  assign n57217 = i_hbusreq8 & ~n57143;
  assign n57218 = i_hbusreq6 & ~n57115;
  assign n57219 = i_hbusreq5 & ~n57104;
  assign n57220 = ~n46615 & ~n54511;
  assign n57221 = ~i_hbusreq5 & ~n57220;
  assign n57222 = ~n57219 & ~n57221;
  assign n57223 = ~controllable_hgrant5 & ~n57222;
  assign n57224 = ~n46535 & ~n57223;
  assign n57225 = controllable_hmaster1 & ~n57224;
  assign n57226 = controllable_hmaster2 & ~n57224;
  assign n57227 = i_hbusreq5 & ~n57109;
  assign n57228 = ~n47640 & ~n54545;
  assign n57229 = ~i_hbusreq5 & ~n57228;
  assign n57230 = ~n57227 & ~n57229;
  assign n57231 = ~controllable_hgrant5 & ~n57230;
  assign n57232 = ~n47610 & ~n57231;
  assign n57233 = ~controllable_hmaster2 & ~n57232;
  assign n57234 = ~n57226 & ~n57233;
  assign n57235 = ~controllable_hmaster1 & ~n57234;
  assign n57236 = ~n57225 & ~n57235;
  assign n57237 = ~i_hbusreq6 & ~n57236;
  assign n57238 = ~n57218 & ~n57237;
  assign n57239 = ~controllable_hgrant6 & ~n57238;
  assign n57240 = ~n47598 & ~n57239;
  assign n57241 = controllable_hmaster0 & ~n57240;
  assign n57242 = i_hbusreq6 & ~n57125;
  assign n57243 = i_hbusreq5 & ~n57119;
  assign n57244 = ~n46866 & ~n54571;
  assign n57245 = ~i_hbusreq5 & ~n57244;
  assign n57246 = ~n57243 & ~n57245;
  assign n57247 = ~controllable_hgrant5 & ~n57246;
  assign n57248 = ~n46804 & ~n57247;
  assign n57249 = ~controllable_hmaster2 & ~n57248;
  assign n57250 = ~n57226 & ~n57249;
  assign n57251 = ~controllable_hmaster1 & ~n57250;
  assign n57252 = ~n57225 & ~n57251;
  assign n57253 = ~i_hbusreq6 & ~n57252;
  assign n57254 = ~n57242 & ~n57253;
  assign n57255 = ~controllable_hgrant6 & ~n57254;
  assign n57256 = ~n46792 & ~n57255;
  assign n57257 = ~controllable_hmaster0 & ~n57256;
  assign n57258 = ~n57241 & ~n57257;
  assign n57259 = i_hlock8 & ~n57258;
  assign n57260 = i_hbusreq6 & ~n57137;
  assign n57261 = i_hbusreq5 & ~n57131;
  assign n57262 = ~n46963 & ~n54599;
  assign n57263 = ~i_hbusreq5 & ~n57262;
  assign n57264 = ~n57261 & ~n57263;
  assign n57265 = ~controllable_hgrant5 & ~n57264;
  assign n57266 = ~n46905 & ~n57265;
  assign n57267 = ~controllable_hmaster2 & ~n57266;
  assign n57268 = ~n57226 & ~n57267;
  assign n57269 = ~controllable_hmaster1 & ~n57268;
  assign n57270 = ~n57225 & ~n57269;
  assign n57271 = ~i_hbusreq6 & ~n57270;
  assign n57272 = ~n57260 & ~n57271;
  assign n57273 = ~controllable_hgrant6 & ~n57272;
  assign n57274 = ~n46893 & ~n57273;
  assign n57275 = ~controllable_hmaster0 & ~n57274;
  assign n57276 = ~n57241 & ~n57275;
  assign n57277 = ~i_hlock8 & ~n57276;
  assign n57278 = ~n57259 & ~n57277;
  assign n57279 = ~i_hbusreq8 & ~n57278;
  assign n57280 = ~n57217 & ~n57279;
  assign n57281 = controllable_hmaster3 & ~n57280;
  assign n57282 = i_hbusreq8 & ~n57201;
  assign n57283 = i_hbusreq6 & ~n57164;
  assign n57284 = controllable_hmaster2 & ~n57248;
  assign n57285 = i_hbusreq5 & ~n57146;
  assign n57286 = ~n47052 & ~n54638;
  assign n57287 = ~i_hbusreq5 & ~n57286;
  assign n57288 = ~n57285 & ~n57287;
  assign n57289 = ~controllable_hgrant5 & ~n57288;
  assign n57290 = ~n47008 & ~n57289;
  assign n57291 = ~controllable_hmaster2 & ~n57290;
  assign n57292 = ~n57284 & ~n57291;
  assign n57293 = controllable_hmaster1 & ~n57292;
  assign n57294 = i_hbusreq5 & ~n57154;
  assign n57295 = i_hlock5 & ~n57244;
  assign n57296 = ~i_hlock5 & ~n57262;
  assign n57297 = ~n57295 & ~n57296;
  assign n57298 = ~i_hbusreq5 & ~n57297;
  assign n57299 = ~n57294 & ~n57298;
  assign n57300 = ~controllable_hgrant5 & ~n57299;
  assign n57301 = ~n47071 & ~n57300;
  assign n57302 = controllable_hmaster2 & ~n57301;
  assign n57303 = i_hbusreq5 & ~n57158;
  assign n57304 = ~n47151 & ~n54671;
  assign n57305 = ~i_hbusreq5 & ~n57304;
  assign n57306 = ~n57303 & ~n57305;
  assign n57307 = ~controllable_hgrant5 & ~n57306;
  assign n57308 = ~n47091 & ~n57307;
  assign n57309 = ~controllable_hmaster2 & ~n57308;
  assign n57310 = ~n57302 & ~n57309;
  assign n57311 = ~controllable_hmaster1 & ~n57310;
  assign n57312 = ~n57293 & ~n57311;
  assign n57313 = ~i_hbusreq6 & ~n57312;
  assign n57314 = ~n57283 & ~n57313;
  assign n57315 = ~controllable_hgrant6 & ~n57314;
  assign n57316 = ~n46995 & ~n57315;
  assign n57317 = controllable_hmaster0 & ~n57316;
  assign n57318 = i_hbusreq6 & ~n57176;
  assign n57319 = ~n33063 & ~n47168;
  assign n57320 = ~n8217 & ~n57319;
  assign n57321 = ~n54688 & ~n57320;
  assign n57322 = i_hlock6 & ~n57321;
  assign n57323 = ~n33095 & ~n47174;
  assign n57324 = ~n8217 & ~n57323;
  assign n57325 = ~n54694 & ~n57324;
  assign n57326 = ~i_hlock6 & ~n57325;
  assign n57327 = ~n57322 & ~n57326;
  assign n57328 = ~i_hbusreq6 & ~n57327;
  assign n57329 = ~n57318 & ~n57328;
  assign n57330 = controllable_hgrant6 & ~n57329;
  assign n57331 = i_hbusreq6 & ~n57197;
  assign n57332 = i_hbusreq5 & ~n57178;
  assign n57333 = ~n47275 & ~n54719;
  assign n57334 = ~i_hbusreq5 & ~n57333;
  assign n57335 = ~n57332 & ~n57334;
  assign n57336 = ~controllable_hgrant5 & ~n57335;
  assign n57337 = ~n47194 & ~n57336;
  assign n57338 = ~controllable_hmaster2 & ~n57337;
  assign n57339 = ~n57284 & ~n57338;
  assign n57340 = controllable_hmaster1 & ~n57339;
  assign n57341 = ~n8378 & ~n33056;
  assign n57342 = ~n54729 & ~n57341;
  assign n57343 = i_hlock5 & ~n57342;
  assign n57344 = ~n8378 & ~n33088;
  assign n57345 = ~n54729 & ~n57344;
  assign n57346 = ~i_hlock5 & ~n57345;
  assign n57347 = ~n57343 & ~n57346;
  assign n57348 = ~i_hbusreq5 & ~n57347;
  assign n57349 = ~n49797 & ~n57348;
  assign n57350 = controllable_hgrant5 & ~n57349;
  assign n57351 = i_hlock4 & ~n47695;
  assign n57352 = ~i_hlock4 & ~n47755;
  assign n57353 = ~n57351 & ~n57352;
  assign n57354 = ~i_hbusreq4 & ~n57353;
  assign n57355 = ~n49829 & ~n57354;
  assign n57356 = ~controllable_hgrant4 & ~n57355;
  assign n57357 = ~n49828 & ~n57356;
  assign n57358 = ~i_hbusreq5 & ~n57357;
  assign n57359 = ~n49809 & ~n57358;
  assign n57360 = ~controllable_hgrant5 & ~n57359;
  assign n57361 = ~n57350 & ~n57360;
  assign n57362 = controllable_hmaster2 & ~n57361;
  assign n57363 = i_hbusreq5 & ~n57184;
  assign n57364 = ~n47412 & ~n54764;
  assign n57365 = ~i_hbusreq5 & ~n57364;
  assign n57366 = ~n57363 & ~n57365;
  assign n57367 = ~controllable_hgrant5 & ~n57366;
  assign n57368 = ~n47336 & ~n57367;
  assign n57369 = ~controllable_hmaster2 & ~n57368;
  assign n57370 = ~n57362 & ~n57369;
  assign n57371 = ~controllable_hmaster1 & ~n57370;
  assign n57372 = ~n57340 & ~n57371;
  assign n57373 = i_hlock6 & ~n57372;
  assign n57374 = controllable_hmaster2 & ~n57266;
  assign n57375 = ~n57338 & ~n57374;
  assign n57376 = controllable_hmaster1 & ~n57375;
  assign n57377 = ~n57371 & ~n57376;
  assign n57378 = ~i_hlock6 & ~n57377;
  assign n57379 = ~n57373 & ~n57378;
  assign n57380 = ~i_hbusreq6 & ~n57379;
  assign n57381 = ~n57331 & ~n57380;
  assign n57382 = ~controllable_hgrant6 & ~n57381;
  assign n57383 = ~n57330 & ~n57382;
  assign n57384 = ~controllable_hmaster0 & ~n57383;
  assign n57385 = ~n57317 & ~n57384;
  assign n57386 = ~i_hbusreq8 & ~n57385;
  assign n57387 = ~n57282 & ~n57386;
  assign n57388 = ~controllable_hmaster3 & ~n57387;
  assign n57389 = ~n57281 & ~n57388;
  assign n57390 = i_hlock7 & ~n57389;
  assign n57391 = i_hbusreq8 & ~n57211;
  assign n57392 = i_hbusreq6 & ~n57207;
  assign n57393 = ~n57291 & ~n57374;
  assign n57394 = controllable_hmaster1 & ~n57393;
  assign n57395 = ~n57311 & ~n57394;
  assign n57396 = ~i_hbusreq6 & ~n57395;
  assign n57397 = ~n57392 & ~n57396;
  assign n57398 = ~controllable_hgrant6 & ~n57397;
  assign n57399 = ~n47451 & ~n57398;
  assign n57400 = controllable_hmaster0 & ~n57399;
  assign n57401 = ~n57384 & ~n57400;
  assign n57402 = ~i_hbusreq8 & ~n57401;
  assign n57403 = ~n57391 & ~n57402;
  assign n57404 = ~controllable_hmaster3 & ~n57403;
  assign n57405 = ~n57281 & ~n57404;
  assign n57406 = ~i_hlock7 & ~n57405;
  assign n57407 = ~n57390 & ~n57406;
  assign n57408 = ~i_hbusreq7 & ~n57407;
  assign n57409 = ~n57216 & ~n57408;
  assign n57410 = n7924 & ~n57409;
  assign n57411 = ~n54369 & ~n57410;
  assign n57412 = n8214 & ~n57411;
  assign n57413 = ~n57103 & ~n57412;
  assign n57414 = ~n8202 & ~n57413;
  assign n57415 = ~n45997 & ~n48785;
  assign n57416 = ~controllable_hgrant4 & ~n57415;
  assign n57417 = ~n45958 & ~n57416;
  assign n57418 = ~controllable_hgrant5 & ~n57417;
  assign n57419 = ~n45950 & ~n57418;
  assign n57420 = controllable_hmaster1 & ~n57419;
  assign n57421 = controllable_hmaster2 & ~n57419;
  assign n57422 = ~n46038 & ~n46151;
  assign n57423 = i_hlock9 & ~n57422;
  assign n57424 = ~n46077 & ~n46209;
  assign n57425 = ~i_hlock9 & ~n57424;
  assign n57426 = ~n57423 & ~n57425;
  assign n57427 = ~controllable_hgrant4 & ~n57426;
  assign n57428 = ~n47498 & ~n57427;
  assign n57429 = ~controllable_hgrant5 & ~n57428;
  assign n57430 = ~n47488 & ~n57429;
  assign n57431 = ~controllable_hmaster2 & ~n57430;
  assign n57432 = ~n57421 & ~n57431;
  assign n57433 = ~controllable_hmaster1 & ~n57432;
  assign n57434 = ~n57420 & ~n57433;
  assign n57435 = ~controllable_hgrant6 & ~n57434;
  assign n57436 = ~n47480 & ~n57435;
  assign n57437 = controllable_hmaster0 & ~n57436;
  assign n57438 = ~controllable_hgrant4 & ~n57422;
  assign n57439 = ~n46127 & ~n57438;
  assign n57440 = ~controllable_hgrant5 & ~n57439;
  assign n57441 = ~n46119 & ~n57440;
  assign n57442 = ~controllable_hmaster2 & ~n57441;
  assign n57443 = ~n57421 & ~n57442;
  assign n57444 = ~controllable_hmaster1 & ~n57443;
  assign n57445 = ~n57420 & ~n57444;
  assign n57446 = ~controllable_hgrant6 & ~n57445;
  assign n57447 = ~n46111 & ~n57446;
  assign n57448 = ~controllable_hmaster0 & ~n57447;
  assign n57449 = ~n57437 & ~n57448;
  assign n57450 = i_hlock8 & ~n57449;
  assign n57451 = ~controllable_hgrant4 & ~n57424;
  assign n57452 = ~n46189 & ~n57451;
  assign n57453 = ~controllable_hgrant5 & ~n57452;
  assign n57454 = ~n46181 & ~n57453;
  assign n57455 = ~controllable_hmaster2 & ~n57454;
  assign n57456 = ~n57421 & ~n57455;
  assign n57457 = ~controllable_hmaster1 & ~n57456;
  assign n57458 = ~n57420 & ~n57457;
  assign n57459 = ~controllable_hgrant6 & ~n57458;
  assign n57460 = ~n46173 & ~n57459;
  assign n57461 = ~controllable_hmaster0 & ~n57460;
  assign n57462 = ~n57437 & ~n57461;
  assign n57463 = ~i_hlock8 & ~n57462;
  assign n57464 = ~n57450 & ~n57463;
  assign n57465 = controllable_hmaster3 & ~n57464;
  assign n57466 = ~n8217 & ~n38218;
  assign n57467 = ~n43905 & ~n57466;
  assign n57468 = i_hlock6 & ~n57467;
  assign n57469 = ~n8217 & ~n38226;
  assign n57470 = ~n43905 & ~n57469;
  assign n57471 = ~i_hlock6 & ~n57470;
  assign n57472 = ~n57468 & ~n57471;
  assign n57473 = controllable_hgrant6 & ~n57472;
  assign n57474 = controllable_hmaster2 & ~n57441;
  assign n57475 = ~n48869 & ~n57474;
  assign n57476 = controllable_hmaster1 & ~n57475;
  assign n57477 = i_hlock5 & ~n57439;
  assign n57478 = ~i_hlock5 & ~n57452;
  assign n57479 = ~n57477 & ~n57478;
  assign n57480 = ~controllable_hgrant5 & ~n57479;
  assign n57481 = ~n46278 & ~n57480;
  assign n57482 = controllable_hmaster2 & ~n57481;
  assign n57483 = ~n46322 & ~n48909;
  assign n57484 = ~controllable_hgrant4 & ~n57483;
  assign n57485 = ~n46300 & ~n57484;
  assign n57486 = ~controllable_hgrant5 & ~n57485;
  assign n57487 = ~n46292 & ~n57486;
  assign n57488 = ~controllable_hmaster2 & ~n57487;
  assign n57489 = ~n57482 & ~n57488;
  assign n57490 = ~controllable_hmaster1 & ~n57489;
  assign n57491 = ~n57476 & ~n57490;
  assign n57492 = ~controllable_hgrant6 & ~n57491;
  assign n57493 = ~n57473 & ~n57492;
  assign n57494 = controllable_hmaster0 & ~n57493;
  assign n57495 = ~n46400 & ~n48959;
  assign n57496 = ~controllable_hgrant4 & ~n57495;
  assign n57497 = ~n46364 & ~n57496;
  assign n57498 = ~controllable_hgrant5 & ~n57497;
  assign n57499 = ~n46356 & ~n57498;
  assign n57500 = ~controllable_hmaster2 & ~n57499;
  assign n57501 = ~n57474 & ~n57500;
  assign n57502 = controllable_hmaster1 & ~n57501;
  assign n57503 = i_hlock4 & ~n57422;
  assign n57504 = ~i_hlock4 & ~n57424;
  assign n57505 = ~n57503 & ~n57504;
  assign n57506 = ~controllable_hgrant4 & ~n57505;
  assign n57507 = ~n46424 & ~n57506;
  assign n57508 = ~controllable_hgrant5 & ~n57507;
  assign n57509 = ~n46416 & ~n57508;
  assign n57510 = controllable_hmaster2 & ~n57509;
  assign n57511 = ~n46468 & ~n49041;
  assign n57512 = ~controllable_hgrant4 & ~n57511;
  assign n57513 = ~n46448 & ~n57512;
  assign n57514 = ~controllable_hgrant5 & ~n57513;
  assign n57515 = ~n46440 & ~n57514;
  assign n57516 = ~controllable_hmaster2 & ~n57515;
  assign n57517 = ~n57510 & ~n57516;
  assign n57518 = ~controllable_hmaster1 & ~n57517;
  assign n57519 = ~n57502 & ~n57518;
  assign n57520 = i_hlock6 & ~n57519;
  assign n57521 = controllable_hmaster2 & ~n57454;
  assign n57522 = ~n57500 & ~n57521;
  assign n57523 = controllable_hmaster1 & ~n57522;
  assign n57524 = ~n57518 & ~n57523;
  assign n57525 = ~i_hlock6 & ~n57524;
  assign n57526 = ~n57520 & ~n57525;
  assign n57527 = ~controllable_hgrant6 & ~n57526;
  assign n57528 = ~n46348 & ~n57527;
  assign n57529 = ~controllable_hmaster0 & ~n57528;
  assign n57530 = ~n57494 & ~n57529;
  assign n57531 = ~controllable_hmaster3 & ~n57530;
  assign n57532 = ~n57465 & ~n57531;
  assign n57533 = i_hlock7 & ~n57532;
  assign n57534 = ~n8217 & ~n38238;
  assign n57535 = ~n44119 & ~n57534;
  assign n57536 = i_hlock6 & ~n57535;
  assign n57537 = ~n8217 & ~n38246;
  assign n57538 = ~n44119 & ~n57537;
  assign n57539 = ~i_hlock6 & ~n57538;
  assign n57540 = ~n57536 & ~n57539;
  assign n57541 = controllable_hgrant6 & ~n57540;
  assign n57542 = ~n48869 & ~n57521;
  assign n57543 = controllable_hmaster1 & ~n57542;
  assign n57544 = ~n57490 & ~n57543;
  assign n57545 = ~controllable_hgrant6 & ~n57544;
  assign n57546 = ~n57541 & ~n57545;
  assign n57547 = controllable_hmaster0 & ~n57546;
  assign n57548 = ~n57529 & ~n57547;
  assign n57549 = ~controllable_hmaster3 & ~n57548;
  assign n57550 = ~n57465 & ~n57549;
  assign n57551 = ~i_hlock7 & ~n57550;
  assign n57552 = ~n57533 & ~n57551;
  assign n57553 = i_hbusreq7 & ~n57552;
  assign n57554 = i_hbusreq8 & ~n57464;
  assign n57555 = i_hbusreq6 & ~n57434;
  assign n57556 = i_hbusreq5 & ~n57417;
  assign n57557 = i_hbusreq4 & ~n57415;
  assign n57558 = i_hbusreq9 & ~n57415;
  assign n57559 = ~n46609 & ~n55373;
  assign n57560 = ~i_hbusreq9 & ~n57559;
  assign n57561 = ~n57558 & ~n57560;
  assign n57562 = ~i_hbusreq4 & ~n57561;
  assign n57563 = ~n57557 & ~n57562;
  assign n57564 = ~controllable_hgrant4 & ~n57563;
  assign n57565 = ~n46553 & ~n57564;
  assign n57566 = ~i_hbusreq5 & ~n57565;
  assign n57567 = ~n57556 & ~n57566;
  assign n57568 = ~controllable_hgrant5 & ~n57567;
  assign n57569 = ~n46535 & ~n57568;
  assign n57570 = controllable_hmaster1 & ~n57569;
  assign n57571 = controllable_hmaster2 & ~n57569;
  assign n57572 = i_hbusreq5 & ~n57428;
  assign n57573 = i_hbusreq4 & ~n57426;
  assign n57574 = i_hbusreq9 & ~n57426;
  assign n57575 = ~n46860 & ~n55400;
  assign n57576 = i_hlock9 & ~n57575;
  assign n57577 = ~n46957 & ~n55413;
  assign n57578 = ~i_hlock9 & ~n57577;
  assign n57579 = ~n57576 & ~n57578;
  assign n57580 = ~i_hbusreq9 & ~n57579;
  assign n57581 = ~n57574 & ~n57580;
  assign n57582 = ~i_hbusreq4 & ~n57581;
  assign n57583 = ~n57573 & ~n57582;
  assign n57584 = ~controllable_hgrant4 & ~n57583;
  assign n57585 = ~n47630 & ~n57584;
  assign n57586 = ~i_hbusreq5 & ~n57585;
  assign n57587 = ~n57572 & ~n57586;
  assign n57588 = ~controllable_hgrant5 & ~n57587;
  assign n57589 = ~n47610 & ~n57588;
  assign n57590 = ~controllable_hmaster2 & ~n57589;
  assign n57591 = ~n57571 & ~n57590;
  assign n57592 = ~controllable_hmaster1 & ~n57591;
  assign n57593 = ~n57570 & ~n57592;
  assign n57594 = ~i_hbusreq6 & ~n57593;
  assign n57595 = ~n57555 & ~n57594;
  assign n57596 = ~controllable_hgrant6 & ~n57595;
  assign n57597 = ~n47598 & ~n57596;
  assign n57598 = controllable_hmaster0 & ~n57597;
  assign n57599 = i_hbusreq6 & ~n57445;
  assign n57600 = i_hbusreq5 & ~n57439;
  assign n57601 = i_hbusreq4 & ~n57422;
  assign n57602 = i_hbusreq9 & ~n57422;
  assign n57603 = ~i_hbusreq9 & ~n57575;
  assign n57604 = ~n57602 & ~n57603;
  assign n57605 = ~i_hbusreq4 & ~n57604;
  assign n57606 = ~n57601 & ~n57605;
  assign n57607 = ~controllable_hgrant4 & ~n57606;
  assign n57608 = ~n46822 & ~n57607;
  assign n57609 = ~i_hbusreq5 & ~n57608;
  assign n57610 = ~n57600 & ~n57609;
  assign n57611 = ~controllable_hgrant5 & ~n57610;
  assign n57612 = ~n46804 & ~n57611;
  assign n57613 = ~controllable_hmaster2 & ~n57612;
  assign n57614 = ~n57571 & ~n57613;
  assign n57615 = ~controllable_hmaster1 & ~n57614;
  assign n57616 = ~n57570 & ~n57615;
  assign n57617 = ~i_hbusreq6 & ~n57616;
  assign n57618 = ~n57599 & ~n57617;
  assign n57619 = ~controllable_hgrant6 & ~n57618;
  assign n57620 = ~n46792 & ~n57619;
  assign n57621 = ~controllable_hmaster0 & ~n57620;
  assign n57622 = ~n57598 & ~n57621;
  assign n57623 = i_hlock8 & ~n57622;
  assign n57624 = i_hbusreq6 & ~n57458;
  assign n57625 = i_hbusreq5 & ~n57452;
  assign n57626 = i_hbusreq4 & ~n57424;
  assign n57627 = i_hbusreq9 & ~n57424;
  assign n57628 = ~i_hbusreq9 & ~n57577;
  assign n57629 = ~n57627 & ~n57628;
  assign n57630 = ~i_hbusreq4 & ~n57629;
  assign n57631 = ~n57626 & ~n57630;
  assign n57632 = ~controllable_hgrant4 & ~n57631;
  assign n57633 = ~n46923 & ~n57632;
  assign n57634 = ~i_hbusreq5 & ~n57633;
  assign n57635 = ~n57625 & ~n57634;
  assign n57636 = ~controllable_hgrant5 & ~n57635;
  assign n57637 = ~n46905 & ~n57636;
  assign n57638 = ~controllable_hmaster2 & ~n57637;
  assign n57639 = ~n57571 & ~n57638;
  assign n57640 = ~controllable_hmaster1 & ~n57639;
  assign n57641 = ~n57570 & ~n57640;
  assign n57642 = ~i_hbusreq6 & ~n57641;
  assign n57643 = ~n57624 & ~n57642;
  assign n57644 = ~controllable_hgrant6 & ~n57643;
  assign n57645 = ~n46893 & ~n57644;
  assign n57646 = ~controllable_hmaster0 & ~n57645;
  assign n57647 = ~n57598 & ~n57646;
  assign n57648 = ~i_hlock8 & ~n57647;
  assign n57649 = ~n57623 & ~n57648;
  assign n57650 = ~i_hbusreq8 & ~n57649;
  assign n57651 = ~n57554 & ~n57650;
  assign n57652 = controllable_hmaster3 & ~n57651;
  assign n57653 = i_hbusreq8 & ~n57530;
  assign n57654 = i_hbusreq6 & ~n57472;
  assign n57655 = ~n8217 & ~n38262;
  assign n57656 = ~n55492 & ~n57655;
  assign n57657 = i_hlock6 & ~n57656;
  assign n57658 = ~n8217 & ~n38273;
  assign n57659 = ~n55492 & ~n57658;
  assign n57660 = ~i_hlock6 & ~n57659;
  assign n57661 = ~n57657 & ~n57660;
  assign n57662 = ~i_hbusreq6 & ~n57661;
  assign n57663 = ~n57654 & ~n57662;
  assign n57664 = controllable_hgrant6 & ~n57663;
  assign n57665 = i_hbusreq6 & ~n57491;
  assign n57666 = controllable_hmaster2 & ~n57612;
  assign n57667 = ~n8378 & ~n33149;
  assign n57668 = ~n55501 & ~n57667;
  assign n57669 = i_hlock5 & ~n57668;
  assign n57670 = ~n8378 & ~n33176;
  assign n57671 = ~n55501 & ~n57670;
  assign n57672 = ~i_hlock5 & ~n57671;
  assign n57673 = ~n57669 & ~n57672;
  assign n57674 = ~i_hbusreq5 & ~n57673;
  assign n57675 = ~n49489 & ~n57674;
  assign n57676 = controllable_hgrant5 & ~n57675;
  assign n57677 = ~n8426 & ~n23467;
  assign n57678 = ~n55510 & ~n57677;
  assign n57679 = ~i_hbusreq9 & ~n57678;
  assign n57680 = ~n49503 & ~n57679;
  assign n57681 = i_hlock4 & ~n57680;
  assign n57682 = ~n8426 & ~n23475;
  assign n57683 = ~n55510 & ~n57682;
  assign n57684 = ~i_hbusreq9 & ~n57683;
  assign n57685 = ~n49510 & ~n57684;
  assign n57686 = ~i_hlock4 & ~n57685;
  assign n57687 = ~n57681 & ~n57686;
  assign n57688 = ~i_hbusreq4 & ~n57687;
  assign n57689 = ~n49502 & ~n57688;
  assign n57690 = controllable_hgrant4 & ~n57689;
  assign n57691 = i_hlock3 & ~n46722;
  assign n57692 = ~i_hlock3 & ~n46756;
  assign n57693 = ~n57691 & ~n57692;
  assign n57694 = ~i_hbusreq3 & ~n57693;
  assign n57695 = ~n49535 & ~n57694;
  assign n57696 = ~controllable_hgrant3 & ~n57695;
  assign n57697 = ~n49534 & ~n57696;
  assign n57698 = ~i_hbusreq9 & ~n57697;
  assign n57699 = ~n49521 & ~n57698;
  assign n57700 = ~i_hbusreq4 & ~n57699;
  assign n57701 = ~n49520 & ~n57700;
  assign n57702 = ~controllable_hgrant4 & ~n57701;
  assign n57703 = ~n57690 & ~n57702;
  assign n57704 = ~i_hbusreq5 & ~n57703;
  assign n57705 = ~n49501 & ~n57704;
  assign n57706 = ~controllable_hgrant5 & ~n57705;
  assign n57707 = ~n57676 & ~n57706;
  assign n57708 = ~controllable_hmaster2 & ~n57707;
  assign n57709 = ~n57666 & ~n57708;
  assign n57710 = controllable_hmaster1 & ~n57709;
  assign n57711 = i_hbusreq5 & ~n57479;
  assign n57712 = i_hlock5 & ~n57608;
  assign n57713 = ~i_hlock5 & ~n57633;
  assign n57714 = ~n57712 & ~n57713;
  assign n57715 = ~i_hbusreq5 & ~n57714;
  assign n57716 = ~n57711 & ~n57715;
  assign n57717 = ~controllable_hgrant5 & ~n57716;
  assign n57718 = ~n47071 & ~n57717;
  assign n57719 = controllable_hmaster2 & ~n57718;
  assign n57720 = i_hbusreq5 & ~n57485;
  assign n57721 = i_hbusreq4 & ~n57483;
  assign n57722 = i_hbusreq9 & ~n57483;
  assign n57723 = ~n47145 & ~n55563;
  assign n57724 = ~i_hbusreq9 & ~n57723;
  assign n57725 = ~n57722 & ~n57724;
  assign n57726 = ~i_hbusreq4 & ~n57725;
  assign n57727 = ~n57721 & ~n57726;
  assign n57728 = ~controllable_hgrant4 & ~n57727;
  assign n57729 = ~n47109 & ~n57728;
  assign n57730 = ~i_hbusreq5 & ~n57729;
  assign n57731 = ~n57720 & ~n57730;
  assign n57732 = ~controllable_hgrant5 & ~n57731;
  assign n57733 = ~n47091 & ~n57732;
  assign n57734 = ~controllable_hmaster2 & ~n57733;
  assign n57735 = ~n57719 & ~n57734;
  assign n57736 = ~controllable_hmaster1 & ~n57735;
  assign n57737 = ~n57710 & ~n57736;
  assign n57738 = ~i_hbusreq6 & ~n57737;
  assign n57739 = ~n57665 & ~n57738;
  assign n57740 = ~controllable_hgrant6 & ~n57739;
  assign n57741 = ~n57664 & ~n57740;
  assign n57742 = controllable_hmaster0 & ~n57741;
  assign n57743 = i_hbusreq6 & ~n57526;
  assign n57744 = i_hbusreq5 & ~n57497;
  assign n57745 = i_hbusreq4 & ~n57495;
  assign n57746 = i_hbusreq9 & ~n57495;
  assign n57747 = ~n47269 & ~n55598;
  assign n57748 = ~i_hbusreq9 & ~n57747;
  assign n57749 = ~n57746 & ~n57748;
  assign n57750 = ~i_hbusreq4 & ~n57749;
  assign n57751 = ~n57745 & ~n57750;
  assign n57752 = ~controllable_hgrant4 & ~n57751;
  assign n57753 = ~n47212 & ~n57752;
  assign n57754 = ~i_hbusreq5 & ~n57753;
  assign n57755 = ~n57744 & ~n57754;
  assign n57756 = ~controllable_hgrant5 & ~n57755;
  assign n57757 = ~n47194 & ~n57756;
  assign n57758 = ~controllable_hmaster2 & ~n57757;
  assign n57759 = ~n57666 & ~n57758;
  assign n57760 = controllable_hmaster1 & ~n57759;
  assign n57761 = i_hbusreq5 & ~n57507;
  assign n57762 = i_hbusreq4 & ~n57505;
  assign n57763 = i_hlock4 & ~n57604;
  assign n57764 = ~i_hlock4 & ~n57629;
  assign n57765 = ~n57763 & ~n57764;
  assign n57766 = ~i_hbusreq4 & ~n57765;
  assign n57767 = ~n57762 & ~n57766;
  assign n57768 = ~controllable_hgrant4 & ~n57767;
  assign n57769 = ~n47312 & ~n57768;
  assign n57770 = ~i_hbusreq5 & ~n57769;
  assign n57771 = ~n57761 & ~n57770;
  assign n57772 = ~controllable_hgrant5 & ~n57771;
  assign n57773 = ~n47294 & ~n57772;
  assign n57774 = controllable_hmaster2 & ~n57773;
  assign n57775 = i_hbusreq5 & ~n57513;
  assign n57776 = i_hbusreq4 & ~n57511;
  assign n57777 = i_hbusreq9 & ~n57511;
  assign n57778 = ~n47406 & ~n55640;
  assign n57779 = ~i_hbusreq9 & ~n57778;
  assign n57780 = ~n57777 & ~n57779;
  assign n57781 = ~i_hbusreq4 & ~n57780;
  assign n57782 = ~n57776 & ~n57781;
  assign n57783 = ~controllable_hgrant4 & ~n57782;
  assign n57784 = ~n47354 & ~n57783;
  assign n57785 = ~i_hbusreq5 & ~n57784;
  assign n57786 = ~n57775 & ~n57785;
  assign n57787 = ~controllable_hgrant5 & ~n57786;
  assign n57788 = ~n47336 & ~n57787;
  assign n57789 = ~controllable_hmaster2 & ~n57788;
  assign n57790 = ~n57774 & ~n57789;
  assign n57791 = ~controllable_hmaster1 & ~n57790;
  assign n57792 = ~n57760 & ~n57791;
  assign n57793 = i_hlock6 & ~n57792;
  assign n57794 = controllable_hmaster2 & ~n57637;
  assign n57795 = ~n57758 & ~n57794;
  assign n57796 = controllable_hmaster1 & ~n57795;
  assign n57797 = ~n57791 & ~n57796;
  assign n57798 = ~i_hlock6 & ~n57797;
  assign n57799 = ~n57793 & ~n57798;
  assign n57800 = ~i_hbusreq6 & ~n57799;
  assign n57801 = ~n57743 & ~n57800;
  assign n57802 = ~controllable_hgrant6 & ~n57801;
  assign n57803 = ~n47182 & ~n57802;
  assign n57804 = ~controllable_hmaster0 & ~n57803;
  assign n57805 = ~n57742 & ~n57804;
  assign n57806 = ~i_hbusreq8 & ~n57805;
  assign n57807 = ~n57653 & ~n57806;
  assign n57808 = ~controllable_hmaster3 & ~n57807;
  assign n57809 = ~n57652 & ~n57808;
  assign n57810 = i_hlock7 & ~n57809;
  assign n57811 = i_hbusreq8 & ~n57548;
  assign n57812 = i_hbusreq6 & ~n57540;
  assign n57813 = ~n8217 & ~n38291;
  assign n57814 = ~n55676 & ~n57813;
  assign n57815 = i_hlock6 & ~n57814;
  assign n57816 = ~n8217 & ~n38302;
  assign n57817 = ~n55676 & ~n57816;
  assign n57818 = ~i_hlock6 & ~n57817;
  assign n57819 = ~n57815 & ~n57818;
  assign n57820 = ~i_hbusreq6 & ~n57819;
  assign n57821 = ~n57812 & ~n57820;
  assign n57822 = controllable_hgrant6 & ~n57821;
  assign n57823 = i_hbusreq6 & ~n57544;
  assign n57824 = ~n57708 & ~n57794;
  assign n57825 = controllable_hmaster1 & ~n57824;
  assign n57826 = ~n57736 & ~n57825;
  assign n57827 = ~i_hbusreq6 & ~n57826;
  assign n57828 = ~n57823 & ~n57827;
  assign n57829 = ~controllable_hgrant6 & ~n57828;
  assign n57830 = ~n57822 & ~n57829;
  assign n57831 = controllable_hmaster0 & ~n57830;
  assign n57832 = ~n57804 & ~n57831;
  assign n57833 = ~i_hbusreq8 & ~n57832;
  assign n57834 = ~n57811 & ~n57833;
  assign n57835 = ~controllable_hmaster3 & ~n57834;
  assign n57836 = ~n57652 & ~n57835;
  assign n57837 = ~i_hlock7 & ~n57836;
  assign n57838 = ~n57810 & ~n57837;
  assign n57839 = ~i_hbusreq7 & ~n57838;
  assign n57840 = ~n57553 & ~n57839;
  assign n57841 = n7924 & ~n57840;
  assign n57842 = ~n55212 & ~n57841;
  assign n57843 = ~n8214 & ~n57842;
  assign n57844 = ~n20645 & ~n46060;
  assign n57845 = n7733 & ~n57844;
  assign n57846 = ~n48798 & ~n57845;
  assign n57847 = n7928 & ~n57846;
  assign n57848 = ~n55708 & ~n57847;
  assign n57849 = ~controllable_hgrant1 & ~n57848;
  assign n57850 = ~n45974 & ~n57849;
  assign n57851 = ~controllable_hgrant3 & ~n57850;
  assign n57852 = ~n45966 & ~n57851;
  assign n57853 = ~controllable_hgrant4 & ~n57852;
  assign n57854 = ~n45958 & ~n57853;
  assign n57855 = ~controllable_hgrant5 & ~n57854;
  assign n57856 = ~n45950 & ~n57855;
  assign n57857 = controllable_hmaster1 & ~n57856;
  assign n57858 = controllable_hmaster2 & ~n57856;
  assign n57859 = ~n20613 & ~n46060;
  assign n57860 = n7733 & ~n57859;
  assign n57861 = ~n43847 & ~n57860;
  assign n57862 = n7928 & ~n57861;
  assign n57863 = ~n8221 & ~n57862;
  assign n57864 = ~controllable_hgrant1 & ~n57863;
  assign n57865 = ~n46143 & ~n57864;
  assign n57866 = ~controllable_hgrant3 & ~n57865;
  assign n57867 = ~n46135 & ~n57866;
  assign n57868 = i_hlock9 & ~n57867;
  assign n57869 = ~n8235 & ~n57862;
  assign n57870 = ~controllable_hgrant1 & ~n57869;
  assign n57871 = ~n46205 & ~n57870;
  assign n57872 = ~controllable_hgrant3 & ~n57871;
  assign n57873 = ~n46197 & ~n57872;
  assign n57874 = ~i_hlock9 & ~n57873;
  assign n57875 = ~n57868 & ~n57874;
  assign n57876 = ~controllable_hgrant4 & ~n57875;
  assign n57877 = ~n47498 & ~n57876;
  assign n57878 = ~controllable_hgrant5 & ~n57877;
  assign n57879 = ~n47488 & ~n57878;
  assign n57880 = ~controllable_hmaster2 & ~n57879;
  assign n57881 = ~n57858 & ~n57880;
  assign n57882 = ~controllable_hmaster1 & ~n57881;
  assign n57883 = ~n57857 & ~n57882;
  assign n57884 = ~controllable_hgrant6 & ~n57883;
  assign n57885 = ~n47480 & ~n57884;
  assign n57886 = controllable_hmaster0 & ~n57885;
  assign n57887 = ~controllable_hgrant4 & ~n57867;
  assign n57888 = ~n46127 & ~n57887;
  assign n57889 = ~controllable_hgrant5 & ~n57888;
  assign n57890 = ~n46119 & ~n57889;
  assign n57891 = ~controllable_hmaster2 & ~n57890;
  assign n57892 = ~n57858 & ~n57891;
  assign n57893 = ~controllable_hmaster1 & ~n57892;
  assign n57894 = ~n57857 & ~n57893;
  assign n57895 = ~controllable_hgrant6 & ~n57894;
  assign n57896 = ~n46111 & ~n57895;
  assign n57897 = ~controllable_hmaster0 & ~n57896;
  assign n57898 = ~n57886 & ~n57897;
  assign n57899 = i_hlock8 & ~n57898;
  assign n57900 = ~controllable_hgrant4 & ~n57873;
  assign n57901 = ~n46189 & ~n57900;
  assign n57902 = ~controllable_hgrant5 & ~n57901;
  assign n57903 = ~n46181 & ~n57902;
  assign n57904 = ~controllable_hmaster2 & ~n57903;
  assign n57905 = ~n57858 & ~n57904;
  assign n57906 = ~controllable_hmaster1 & ~n57905;
  assign n57907 = ~n57857 & ~n57906;
  assign n57908 = ~controllable_hgrant6 & ~n57907;
  assign n57909 = ~n46173 & ~n57908;
  assign n57910 = ~controllable_hmaster0 & ~n57909;
  assign n57911 = ~n57886 & ~n57910;
  assign n57912 = ~i_hlock8 & ~n57911;
  assign n57913 = ~n57899 & ~n57912;
  assign n57914 = controllable_hmaster3 & ~n57913;
  assign n57915 = controllable_hmaster2 & ~n57890;
  assign n57916 = i_hlock3 & ~n57865;
  assign n57917 = ~i_hlock3 & ~n57871;
  assign n57918 = ~n57916 & ~n57917;
  assign n57919 = ~controllable_hgrant3 & ~n57918;
  assign n57920 = ~n46258 & ~n57919;
  assign n57921 = ~controllable_hgrant4 & ~n57920;
  assign n57922 = ~n46250 & ~n57921;
  assign n57923 = ~controllable_hgrant5 & ~n57922;
  assign n57924 = ~n46242 & ~n57923;
  assign n57925 = ~controllable_hmaster2 & ~n57924;
  assign n57926 = ~n57915 & ~n57925;
  assign n57927 = controllable_hmaster1 & ~n57926;
  assign n57928 = i_hlock5 & ~n57888;
  assign n57929 = ~i_hlock5 & ~n57901;
  assign n57930 = ~n57928 & ~n57929;
  assign n57931 = ~controllable_hgrant5 & ~n57930;
  assign n57932 = ~n46278 & ~n57931;
  assign n57933 = controllable_hmaster2 & ~n57932;
  assign n57934 = i_hlock1 & ~n57863;
  assign n57935 = ~i_hlock1 & ~n57869;
  assign n57936 = ~n57934 & ~n57935;
  assign n57937 = ~controllable_hgrant1 & ~n57936;
  assign n57938 = ~n46316 & ~n57937;
  assign n57939 = ~controllable_hgrant3 & ~n57938;
  assign n57940 = ~n46308 & ~n57939;
  assign n57941 = ~controllable_hgrant4 & ~n57940;
  assign n57942 = ~n46300 & ~n57941;
  assign n57943 = ~controllable_hgrant5 & ~n57942;
  assign n57944 = ~n46292 & ~n57943;
  assign n57945 = ~controllable_hmaster2 & ~n57944;
  assign n57946 = ~n57933 & ~n57945;
  assign n57947 = ~controllable_hmaster1 & ~n57946;
  assign n57948 = ~n57927 & ~n57947;
  assign n57949 = ~controllable_hgrant6 & ~n57948;
  assign n57950 = ~n46233 & ~n57949;
  assign n57951 = controllable_hmaster0 & ~n57950;
  assign n57952 = ~n30312 & ~n31016;
  assign n57953 = controllable_hmaster1 & ~n57952;
  assign n57954 = ~n31063 & ~n57953;
  assign n57955 = ~n8217 & ~n57954;
  assign n57956 = ~n43999 & ~n57955;
  assign n57957 = i_hlock6 & ~n57956;
  assign n57958 = ~n30415 & ~n31123;
  assign n57959 = controllable_hmaster1 & ~n57958;
  assign n57960 = ~n31170 & ~n57959;
  assign n57961 = ~n8217 & ~n57960;
  assign n57962 = ~n44009 & ~n57961;
  assign n57963 = ~i_hlock6 & ~n57962;
  assign n57964 = ~n57957 & ~n57963;
  assign n57965 = controllable_hgrant6 & ~n57964;
  assign n57966 = ~n48991 & ~n57915;
  assign n57967 = controllable_hmaster1 & ~n57966;
  assign n57968 = i_hlock4 & ~n57867;
  assign n57969 = ~i_hlock4 & ~n57873;
  assign n57970 = ~n57968 & ~n57969;
  assign n57971 = ~controllable_hgrant4 & ~n57970;
  assign n57972 = ~n46424 & ~n57971;
  assign n57973 = ~controllable_hgrant5 & ~n57972;
  assign n57974 = ~n46416 & ~n57973;
  assign n57975 = controllable_hmaster2 & ~n57974;
  assign n57976 = ~n8440 & ~n57862;
  assign n57977 = ~controllable_hgrant1 & ~n57976;
  assign n57978 = ~n46464 & ~n57977;
  assign n57979 = ~controllable_hgrant3 & ~n57978;
  assign n57980 = ~n46456 & ~n57979;
  assign n57981 = ~controllable_hgrant4 & ~n57980;
  assign n57982 = ~n46448 & ~n57981;
  assign n57983 = ~controllable_hgrant5 & ~n57982;
  assign n57984 = ~n46440 & ~n57983;
  assign n57985 = ~controllable_hmaster2 & ~n57984;
  assign n57986 = ~n57975 & ~n57985;
  assign n57987 = ~controllable_hmaster1 & ~n57986;
  assign n57988 = ~n57967 & ~n57987;
  assign n57989 = i_hlock6 & ~n57988;
  assign n57990 = controllable_hmaster2 & ~n57903;
  assign n57991 = ~n48991 & ~n57990;
  assign n57992 = controllable_hmaster1 & ~n57991;
  assign n57993 = ~n57987 & ~n57992;
  assign n57994 = ~i_hlock6 & ~n57993;
  assign n57995 = ~n57989 & ~n57994;
  assign n57996 = ~controllable_hgrant6 & ~n57995;
  assign n57997 = ~n57965 & ~n57996;
  assign n57998 = ~controllable_hmaster0 & ~n57997;
  assign n57999 = ~n57951 & ~n57998;
  assign n58000 = ~controllable_hmaster3 & ~n57999;
  assign n58001 = ~n57914 & ~n58000;
  assign n58002 = i_hlock7 & ~n58001;
  assign n58003 = ~n57925 & ~n57990;
  assign n58004 = controllable_hmaster1 & ~n58003;
  assign n58005 = ~n57947 & ~n58004;
  assign n58006 = ~controllable_hgrant6 & ~n58005;
  assign n58007 = ~n46499 & ~n58006;
  assign n58008 = controllable_hmaster0 & ~n58007;
  assign n58009 = ~n57998 & ~n58008;
  assign n58010 = ~controllable_hmaster3 & ~n58009;
  assign n58011 = ~n57914 & ~n58010;
  assign n58012 = ~i_hlock7 & ~n58011;
  assign n58013 = ~n58002 & ~n58012;
  assign n58014 = i_hbusreq7 & ~n58013;
  assign n58015 = i_hbusreq8 & ~n57913;
  assign n58016 = i_hbusreq6 & ~n57883;
  assign n58017 = i_hbusreq5 & ~n57854;
  assign n58018 = i_hbusreq4 & ~n57852;
  assign n58019 = i_hbusreq9 & ~n57852;
  assign n58020 = i_hbusreq3 & ~n57850;
  assign n58021 = i_hbusreq1 & ~n57848;
  assign n58022 = ~n20950 & ~n56454;
  assign n58023 = n7733 & ~n58022;
  assign n58024 = ~n56443 & ~n58023;
  assign n58025 = n7928 & ~n58024;
  assign n58026 = ~n55906 & ~n58025;
  assign n58027 = ~i_hbusreq1 & ~n58026;
  assign n58028 = ~n58021 & ~n58027;
  assign n58029 = ~controllable_hgrant1 & ~n58028;
  assign n58030 = ~n46578 & ~n58029;
  assign n58031 = ~i_hbusreq3 & ~n58030;
  assign n58032 = ~n58020 & ~n58031;
  assign n58033 = ~controllable_hgrant3 & ~n58032;
  assign n58034 = ~n46566 & ~n58033;
  assign n58035 = ~i_hbusreq9 & ~n58034;
  assign n58036 = ~n58019 & ~n58035;
  assign n58037 = ~i_hbusreq4 & ~n58036;
  assign n58038 = ~n58018 & ~n58037;
  assign n58039 = ~controllable_hgrant4 & ~n58038;
  assign n58040 = ~n46553 & ~n58039;
  assign n58041 = ~i_hbusreq5 & ~n58040;
  assign n58042 = ~n58017 & ~n58041;
  assign n58043 = ~controllable_hgrant5 & ~n58042;
  assign n58044 = ~n46535 & ~n58043;
  assign n58045 = controllable_hmaster1 & ~n58044;
  assign n58046 = controllable_hmaster2 & ~n58044;
  assign n58047 = i_hbusreq5 & ~n57877;
  assign n58048 = i_hbusreq4 & ~n57875;
  assign n58049 = i_hbusreq9 & ~n57875;
  assign n58050 = i_hbusreq3 & ~n57865;
  assign n58051 = i_hbusreq1 & ~n57863;
  assign n58052 = ~n20882 & ~n56454;
  assign n58053 = n7733 & ~n58052;
  assign n58054 = ~n44407 & ~n58053;
  assign n58055 = n7928 & ~n58054;
  assign n58056 = ~n8265 & ~n58055;
  assign n58057 = ~i_hbusreq1 & ~n58056;
  assign n58058 = ~n58051 & ~n58057;
  assign n58059 = ~controllable_hgrant1 & ~n58058;
  assign n58060 = ~n46847 & ~n58059;
  assign n58061 = ~i_hbusreq3 & ~n58060;
  assign n58062 = ~n58050 & ~n58061;
  assign n58063 = ~controllable_hgrant3 & ~n58062;
  assign n58064 = ~n46835 & ~n58063;
  assign n58065 = i_hlock9 & ~n58064;
  assign n58066 = i_hbusreq3 & ~n57871;
  assign n58067 = i_hbusreq1 & ~n57869;
  assign n58068 = ~n8297 & ~n58055;
  assign n58069 = ~i_hbusreq1 & ~n58068;
  assign n58070 = ~n58067 & ~n58069;
  assign n58071 = ~controllable_hgrant1 & ~n58070;
  assign n58072 = ~n46948 & ~n58071;
  assign n58073 = ~i_hbusreq3 & ~n58072;
  assign n58074 = ~n58066 & ~n58073;
  assign n58075 = ~controllable_hgrant3 & ~n58074;
  assign n58076 = ~n46936 & ~n58075;
  assign n58077 = ~i_hlock9 & ~n58076;
  assign n58078 = ~n58065 & ~n58077;
  assign n58079 = ~i_hbusreq9 & ~n58078;
  assign n58080 = ~n58049 & ~n58079;
  assign n58081 = ~i_hbusreq4 & ~n58080;
  assign n58082 = ~n58048 & ~n58081;
  assign n58083 = ~controllable_hgrant4 & ~n58082;
  assign n58084 = ~n47630 & ~n58083;
  assign n58085 = ~i_hbusreq5 & ~n58084;
  assign n58086 = ~n58047 & ~n58085;
  assign n58087 = ~controllable_hgrant5 & ~n58086;
  assign n58088 = ~n47610 & ~n58087;
  assign n58089 = ~controllable_hmaster2 & ~n58088;
  assign n58090 = ~n58046 & ~n58089;
  assign n58091 = ~controllable_hmaster1 & ~n58090;
  assign n58092 = ~n58045 & ~n58091;
  assign n58093 = ~i_hbusreq6 & ~n58092;
  assign n58094 = ~n58016 & ~n58093;
  assign n58095 = ~controllable_hgrant6 & ~n58094;
  assign n58096 = ~n47598 & ~n58095;
  assign n58097 = controllable_hmaster0 & ~n58096;
  assign n58098 = i_hbusreq6 & ~n57894;
  assign n58099 = i_hbusreq5 & ~n57888;
  assign n58100 = i_hbusreq4 & ~n57867;
  assign n58101 = i_hbusreq9 & ~n57867;
  assign n58102 = ~i_hbusreq9 & ~n58064;
  assign n58103 = ~n58101 & ~n58102;
  assign n58104 = ~i_hbusreq4 & ~n58103;
  assign n58105 = ~n58100 & ~n58104;
  assign n58106 = ~controllable_hgrant4 & ~n58105;
  assign n58107 = ~n46822 & ~n58106;
  assign n58108 = ~i_hbusreq5 & ~n58107;
  assign n58109 = ~n58099 & ~n58108;
  assign n58110 = ~controllable_hgrant5 & ~n58109;
  assign n58111 = ~n46804 & ~n58110;
  assign n58112 = ~controllable_hmaster2 & ~n58111;
  assign n58113 = ~n58046 & ~n58112;
  assign n58114 = ~controllable_hmaster1 & ~n58113;
  assign n58115 = ~n58045 & ~n58114;
  assign n58116 = ~i_hbusreq6 & ~n58115;
  assign n58117 = ~n58098 & ~n58116;
  assign n58118 = ~controllable_hgrant6 & ~n58117;
  assign n58119 = ~n46792 & ~n58118;
  assign n58120 = ~controllable_hmaster0 & ~n58119;
  assign n58121 = ~n58097 & ~n58120;
  assign n58122 = i_hlock8 & ~n58121;
  assign n58123 = i_hbusreq6 & ~n57907;
  assign n58124 = i_hbusreq5 & ~n57901;
  assign n58125 = i_hbusreq4 & ~n57873;
  assign n58126 = i_hbusreq9 & ~n57873;
  assign n58127 = ~i_hbusreq9 & ~n58076;
  assign n58128 = ~n58126 & ~n58127;
  assign n58129 = ~i_hbusreq4 & ~n58128;
  assign n58130 = ~n58125 & ~n58129;
  assign n58131 = ~controllable_hgrant4 & ~n58130;
  assign n58132 = ~n46923 & ~n58131;
  assign n58133 = ~i_hbusreq5 & ~n58132;
  assign n58134 = ~n58124 & ~n58133;
  assign n58135 = ~controllable_hgrant5 & ~n58134;
  assign n58136 = ~n46905 & ~n58135;
  assign n58137 = ~controllable_hmaster2 & ~n58136;
  assign n58138 = ~n58046 & ~n58137;
  assign n58139 = ~controllable_hmaster1 & ~n58138;
  assign n58140 = ~n58045 & ~n58139;
  assign n58141 = ~i_hbusreq6 & ~n58140;
  assign n58142 = ~n58123 & ~n58141;
  assign n58143 = ~controllable_hgrant6 & ~n58142;
  assign n58144 = ~n46893 & ~n58143;
  assign n58145 = ~controllable_hmaster0 & ~n58144;
  assign n58146 = ~n58097 & ~n58145;
  assign n58147 = ~i_hlock8 & ~n58146;
  assign n58148 = ~n58122 & ~n58147;
  assign n58149 = ~i_hbusreq8 & ~n58148;
  assign n58150 = ~n58015 & ~n58149;
  assign n58151 = controllable_hmaster3 & ~n58150;
  assign n58152 = i_hbusreq8 & ~n57999;
  assign n58153 = i_hbusreq6 & ~n57948;
  assign n58154 = controllable_hmaster2 & ~n58111;
  assign n58155 = i_hbusreq5 & ~n57922;
  assign n58156 = i_hbusreq4 & ~n57920;
  assign n58157 = i_hbusreq9 & ~n57920;
  assign n58158 = i_hbusreq3 & ~n57918;
  assign n58159 = i_hlock3 & ~n58060;
  assign n58160 = ~i_hlock3 & ~n58072;
  assign n58161 = ~n58159 & ~n58160;
  assign n58162 = ~i_hbusreq3 & ~n58161;
  assign n58163 = ~n58158 & ~n58162;
  assign n58164 = ~controllable_hgrant3 & ~n58163;
  assign n58165 = ~n47039 & ~n58164;
  assign n58166 = ~i_hbusreq9 & ~n58165;
  assign n58167 = ~n58157 & ~n58166;
  assign n58168 = ~i_hbusreq4 & ~n58167;
  assign n58169 = ~n58156 & ~n58168;
  assign n58170 = ~controllable_hgrant4 & ~n58169;
  assign n58171 = ~n47026 & ~n58170;
  assign n58172 = ~i_hbusreq5 & ~n58171;
  assign n58173 = ~n58155 & ~n58172;
  assign n58174 = ~controllable_hgrant5 & ~n58173;
  assign n58175 = ~n47008 & ~n58174;
  assign n58176 = ~controllable_hmaster2 & ~n58175;
  assign n58177 = ~n58154 & ~n58176;
  assign n58178 = controllable_hmaster1 & ~n58177;
  assign n58179 = i_hbusreq5 & ~n57930;
  assign n58180 = i_hlock5 & ~n58107;
  assign n58181 = ~i_hlock5 & ~n58132;
  assign n58182 = ~n58180 & ~n58181;
  assign n58183 = ~i_hbusreq5 & ~n58182;
  assign n58184 = ~n58179 & ~n58183;
  assign n58185 = ~controllable_hgrant5 & ~n58184;
  assign n58186 = ~n47071 & ~n58185;
  assign n58187 = controllable_hmaster2 & ~n58186;
  assign n58188 = i_hbusreq5 & ~n57942;
  assign n58189 = i_hbusreq4 & ~n57940;
  assign n58190 = i_hbusreq9 & ~n57940;
  assign n58191 = i_hbusreq3 & ~n57938;
  assign n58192 = i_hbusreq1 & ~n57936;
  assign n58193 = i_hlock1 & ~n58056;
  assign n58194 = ~i_hlock1 & ~n58068;
  assign n58195 = ~n58193 & ~n58194;
  assign n58196 = ~i_hbusreq1 & ~n58195;
  assign n58197 = ~n58192 & ~n58196;
  assign n58198 = ~controllable_hgrant1 & ~n58197;
  assign n58199 = ~n47134 & ~n58198;
  assign n58200 = ~i_hbusreq3 & ~n58199;
  assign n58201 = ~n58191 & ~n58200;
  assign n58202 = ~controllable_hgrant3 & ~n58201;
  assign n58203 = ~n47122 & ~n58202;
  assign n58204 = ~i_hbusreq9 & ~n58203;
  assign n58205 = ~n58190 & ~n58204;
  assign n58206 = ~i_hbusreq4 & ~n58205;
  assign n58207 = ~n58189 & ~n58206;
  assign n58208 = ~controllable_hgrant4 & ~n58207;
  assign n58209 = ~n47109 & ~n58208;
  assign n58210 = ~i_hbusreq5 & ~n58209;
  assign n58211 = ~n58188 & ~n58210;
  assign n58212 = ~controllable_hgrant5 & ~n58211;
  assign n58213 = ~n47091 & ~n58212;
  assign n58214 = ~controllable_hmaster2 & ~n58213;
  assign n58215 = ~n58187 & ~n58214;
  assign n58216 = ~controllable_hmaster1 & ~n58215;
  assign n58217 = ~n58178 & ~n58216;
  assign n58218 = ~i_hbusreq6 & ~n58217;
  assign n58219 = ~n58153 & ~n58218;
  assign n58220 = ~controllable_hgrant6 & ~n58219;
  assign n58221 = ~n46995 & ~n58220;
  assign n58222 = controllable_hmaster0 & ~n58221;
  assign n58223 = i_hbusreq6 & ~n57964;
  assign n58224 = ~n31295 & ~n33248;
  assign n58225 = controllable_hmaster1 & ~n58224;
  assign n58226 = ~n31390 & ~n58225;
  assign n58227 = ~n8217 & ~n58226;
  assign n58228 = ~n56660 & ~n58227;
  assign n58229 = i_hlock6 & ~n58228;
  assign n58230 = ~n31517 & ~n33281;
  assign n58231 = controllable_hmaster1 & ~n58230;
  assign n58232 = ~n31612 & ~n58231;
  assign n58233 = ~n8217 & ~n58232;
  assign n58234 = ~n56670 & ~n58233;
  assign n58235 = ~i_hlock6 & ~n58234;
  assign n58236 = ~n58229 & ~n58235;
  assign n58237 = ~i_hbusreq6 & ~n58236;
  assign n58238 = ~n58223 & ~n58237;
  assign n58239 = controllable_hgrant6 & ~n58238;
  assign n58240 = i_hbusreq6 & ~n57995;
  assign n58241 = ~n8378 & ~n33243;
  assign n58242 = ~n56683 & ~n58241;
  assign n58243 = i_hlock5 & ~n58242;
  assign n58244 = ~n8378 & ~n33276;
  assign n58245 = ~n56683 & ~n58244;
  assign n58246 = ~i_hlock5 & ~n58245;
  assign n58247 = ~n58243 & ~n58246;
  assign n58248 = ~i_hbusreq5 & ~n58247;
  assign n58249 = ~n49693 & ~n58248;
  assign n58250 = controllable_hgrant5 & ~n58249;
  assign n58251 = ~n8426 & ~n23557;
  assign n58252 = ~n56692 & ~n58251;
  assign n58253 = ~i_hbusreq9 & ~n58252;
  assign n58254 = ~n49707 & ~n58253;
  assign n58255 = i_hlock4 & ~n58254;
  assign n58256 = ~n8426 & ~n23567;
  assign n58257 = ~n56692 & ~n58256;
  assign n58258 = ~i_hbusreq9 & ~n58257;
  assign n58259 = ~n49714 & ~n58258;
  assign n58260 = ~i_hlock4 & ~n58259;
  assign n58261 = ~n58255 & ~n58260;
  assign n58262 = ~i_hbusreq4 & ~n58261;
  assign n58263 = ~n49706 & ~n58262;
  assign n58264 = controllable_hgrant4 & ~n58263;
  assign n58265 = ~n8365 & ~n23553;
  assign n58266 = ~n56703 & ~n58265;
  assign n58267 = i_hlock3 & ~n58266;
  assign n58268 = ~n8365 & ~n23563;
  assign n58269 = ~n56703 & ~n58268;
  assign n58270 = ~i_hlock3 & ~n58269;
  assign n58271 = ~n58267 & ~n58270;
  assign n58272 = ~i_hbusreq3 & ~n58271;
  assign n58273 = ~n49726 & ~n58272;
  assign n58274 = controllable_hgrant3 & ~n58273;
  assign n58275 = ~n8389 & ~n23549;
  assign n58276 = ~n56711 & ~n58275;
  assign n58277 = i_hlock1 & ~n58276;
  assign n58278 = ~n8389 & ~n23559;
  assign n58279 = ~n56711 & ~n58278;
  assign n58280 = ~i_hlock1 & ~n58279;
  assign n58281 = ~n58277 & ~n58280;
  assign n58282 = ~i_hbusreq1 & ~n58281;
  assign n58283 = ~n49739 & ~n58282;
  assign n58284 = controllable_hgrant1 & ~n58283;
  assign n58285 = ~n46713 & ~n49770;
  assign n58286 = n7733 & ~n58285;
  assign n58287 = ~n56719 & ~n58286;
  assign n58288 = n7928 & ~n58287;
  assign n58289 = ~n43545 & ~n58288;
  assign n58290 = ~i_hbusreq1 & ~n58289;
  assign n58291 = ~n49751 & ~n58290;
  assign n58292 = ~controllable_hgrant1 & ~n58291;
  assign n58293 = ~n58284 & ~n58292;
  assign n58294 = ~i_hbusreq3 & ~n58293;
  assign n58295 = ~n49738 & ~n58294;
  assign n58296 = ~controllable_hgrant3 & ~n58295;
  assign n58297 = ~n58274 & ~n58296;
  assign n58298 = ~i_hbusreq9 & ~n58297;
  assign n58299 = ~n49725 & ~n58298;
  assign n58300 = ~i_hbusreq4 & ~n58299;
  assign n58301 = ~n49724 & ~n58300;
  assign n58302 = ~controllable_hgrant4 & ~n58301;
  assign n58303 = ~n58264 & ~n58302;
  assign n58304 = ~i_hbusreq5 & ~n58303;
  assign n58305 = ~n49705 & ~n58304;
  assign n58306 = ~controllable_hgrant5 & ~n58305;
  assign n58307 = ~n58250 & ~n58306;
  assign n58308 = ~controllable_hmaster2 & ~n58307;
  assign n58309 = ~n58154 & ~n58308;
  assign n58310 = controllable_hmaster1 & ~n58309;
  assign n58311 = i_hbusreq5 & ~n57972;
  assign n58312 = i_hbusreq4 & ~n57970;
  assign n58313 = i_hlock4 & ~n58103;
  assign n58314 = ~i_hlock4 & ~n58128;
  assign n58315 = ~n58313 & ~n58314;
  assign n58316 = ~i_hbusreq4 & ~n58315;
  assign n58317 = ~n58312 & ~n58316;
  assign n58318 = ~controllable_hgrant4 & ~n58317;
  assign n58319 = ~n47312 & ~n58318;
  assign n58320 = ~i_hbusreq5 & ~n58319;
  assign n58321 = ~n58311 & ~n58320;
  assign n58322 = ~controllable_hgrant5 & ~n58321;
  assign n58323 = ~n47294 & ~n58322;
  assign n58324 = controllable_hmaster2 & ~n58323;
  assign n58325 = i_hbusreq5 & ~n57982;
  assign n58326 = i_hbusreq4 & ~n57980;
  assign n58327 = i_hbusreq9 & ~n57980;
  assign n58328 = i_hbusreq3 & ~n57978;
  assign n58329 = i_hbusreq1 & ~n57976;
  assign n58330 = ~n21358 & ~n56781;
  assign n58331 = n7733 & ~n58330;
  assign n58332 = ~n44867 & ~n58331;
  assign n58333 = n7928 & ~n58332;
  assign n58334 = ~n8440 & ~n58333;
  assign n58335 = ~i_hbusreq1 & ~n58334;
  assign n58336 = ~n58329 & ~n58335;
  assign n58337 = ~controllable_hgrant1 & ~n58336;
  assign n58338 = ~n47379 & ~n58337;
  assign n58339 = ~i_hbusreq3 & ~n58338;
  assign n58340 = ~n58328 & ~n58339;
  assign n58341 = ~controllable_hgrant3 & ~n58340;
  assign n58342 = ~n47367 & ~n58341;
  assign n58343 = ~i_hbusreq9 & ~n58342;
  assign n58344 = ~n58327 & ~n58343;
  assign n58345 = ~i_hbusreq4 & ~n58344;
  assign n58346 = ~n58326 & ~n58345;
  assign n58347 = ~controllable_hgrant4 & ~n58346;
  assign n58348 = ~n47354 & ~n58347;
  assign n58349 = ~i_hbusreq5 & ~n58348;
  assign n58350 = ~n58325 & ~n58349;
  assign n58351 = ~controllable_hgrant5 & ~n58350;
  assign n58352 = ~n47336 & ~n58351;
  assign n58353 = ~controllable_hmaster2 & ~n58352;
  assign n58354 = ~n58324 & ~n58353;
  assign n58355 = ~controllable_hmaster1 & ~n58354;
  assign n58356 = ~n58310 & ~n58355;
  assign n58357 = i_hlock6 & ~n58356;
  assign n58358 = controllable_hmaster2 & ~n58136;
  assign n58359 = ~n58308 & ~n58358;
  assign n58360 = controllable_hmaster1 & ~n58359;
  assign n58361 = ~n58355 & ~n58360;
  assign n58362 = ~i_hlock6 & ~n58361;
  assign n58363 = ~n58357 & ~n58362;
  assign n58364 = ~i_hbusreq6 & ~n58363;
  assign n58365 = ~n58240 & ~n58364;
  assign n58366 = ~controllable_hgrant6 & ~n58365;
  assign n58367 = ~n58239 & ~n58366;
  assign n58368 = ~controllable_hmaster0 & ~n58367;
  assign n58369 = ~n58222 & ~n58368;
  assign n58370 = ~i_hbusreq8 & ~n58369;
  assign n58371 = ~n58152 & ~n58370;
  assign n58372 = ~controllable_hmaster3 & ~n58371;
  assign n58373 = ~n58151 & ~n58372;
  assign n58374 = i_hlock7 & ~n58373;
  assign n58375 = i_hbusreq8 & ~n58009;
  assign n58376 = i_hbusreq6 & ~n58005;
  assign n58377 = ~n58176 & ~n58358;
  assign n58378 = controllable_hmaster1 & ~n58377;
  assign n58379 = ~n58216 & ~n58378;
  assign n58380 = ~i_hbusreq6 & ~n58379;
  assign n58381 = ~n58376 & ~n58380;
  assign n58382 = ~controllable_hgrant6 & ~n58381;
  assign n58383 = ~n47451 & ~n58382;
  assign n58384 = controllable_hmaster0 & ~n58383;
  assign n58385 = ~n58368 & ~n58384;
  assign n58386 = ~i_hbusreq8 & ~n58385;
  assign n58387 = ~n58375 & ~n58386;
  assign n58388 = ~controllable_hmaster3 & ~n58387;
  assign n58389 = ~n58151 & ~n58388;
  assign n58390 = ~i_hlock7 & ~n58389;
  assign n58391 = ~n58374 & ~n58390;
  assign n58392 = ~i_hbusreq7 & ~n58391;
  assign n58393 = ~n58014 & ~n58392;
  assign n58394 = n7924 & ~n58393;
  assign n58395 = ~n56231 & ~n58394;
  assign n58396 = n8214 & ~n58395;
  assign n58397 = ~n57843 & ~n58396;
  assign n58398 = n8202 & ~n58397;
  assign n58399 = ~n57414 & ~n58398;
  assign n58400 = n7920 & ~n58399;
  assign n58401 = ~n40177 & ~n58400;
  assign n58402 = n7728 & ~n58401;
  assign n58403 = ~n50003 & ~n58402;
  assign n58404 = ~n7723 & ~n58403;
  assign n58405 = ~n56860 & ~n58404;
  assign n58406 = ~n7714 & ~n58405;
  assign n58407 = ~n56859 & ~n58406;
  assign n58408 = ~n7705 & ~n58407;
  assign n58409 = ~n51653 & ~n58408;
  assign n58410 = n7808 & ~n58409;
  assign n58411 = ~n50195 & ~n58410;
  assign n58412 = ~n8195 & ~n58411;
  assign n58413 = controllable_hgrant6 & ~n10297;
  assign n58414 = ~controllable_hmaster2 & ~n39818;
  assign n58415 = ~controllable_hmaster1 & ~n58414;
  assign n58416 = ~controllable_hmaster1 & ~n58415;
  assign n58417 = ~controllable_hgrant6 & ~n58416;
  assign n58418 = ~n58413 & ~n58417;
  assign n58419 = controllable_hmaster0 & ~n58418;
  assign n58420 = controllable_hmaster0 & ~n58419;
  assign n58421 = ~controllable_hmaster3 & ~n58420;
  assign n58422 = ~controllable_hmaster3 & ~n58421;
  assign n58423 = i_hbusreq7 & ~n58422;
  assign n58424 = i_hbusreq8 & ~n58420;
  assign n58425 = controllable_hgrant6 & ~n10309;
  assign n58426 = i_hbusreq6 & ~n58416;
  assign n58427 = ~controllable_hmaster2 & ~n40039;
  assign n58428 = ~controllable_hmaster1 & ~n58427;
  assign n58429 = ~controllable_hmaster1 & ~n58428;
  assign n58430 = ~i_hbusreq6 & ~n58429;
  assign n58431 = ~n58426 & ~n58430;
  assign n58432 = ~controllable_hgrant6 & ~n58431;
  assign n58433 = ~n58425 & ~n58432;
  assign n58434 = controllable_hmaster0 & ~n58433;
  assign n58435 = controllable_hmaster0 & ~n58434;
  assign n58436 = ~i_hbusreq8 & ~n58435;
  assign n58437 = ~n58424 & ~n58436;
  assign n58438 = ~controllable_hmaster3 & ~n58437;
  assign n58439 = ~controllable_hmaster3 & ~n58438;
  assign n58440 = ~i_hbusreq7 & ~n58439;
  assign n58441 = ~n58423 & ~n58440;
  assign n58442 = n7924 & ~n58441;
  assign n58443 = n7924 & ~n58442;
  assign n58444 = ~n8214 & ~n58443;
  assign n58445 = ~n10330 & ~n58444;
  assign n58446 = ~n8202 & ~n58445;
  assign n58447 = controllable_hgrant6 & ~n10339;
  assign n58448 = controllable_hgrant5 & ~n10334;
  assign n58449 = controllable_hgrant4 & ~n10334;
  assign n58450 = controllable_hgrant3 & ~n10334;
  assign n58451 = controllable_hgrant1 & ~n10334;
  assign n58452 = ~n7824 & n7928;
  assign n58453 = n7928 & ~n58452;
  assign n58454 = ~controllable_hgrant1 & ~n58453;
  assign n58455 = ~n58451 & ~n58454;
  assign n58456 = ~controllable_hgrant3 & ~n58455;
  assign n58457 = ~n58450 & ~n58456;
  assign n58458 = ~controllable_hgrant4 & ~n58457;
  assign n58459 = ~n58449 & ~n58458;
  assign n58460 = ~controllable_hgrant5 & ~n58459;
  assign n58461 = ~n58448 & ~n58460;
  assign n58462 = controllable_hmaster1 & ~n58461;
  assign n58463 = controllable_hmaster2 & ~n58461;
  assign n58464 = controllable_hmaster2 & ~n58463;
  assign n58465 = ~controllable_hmaster1 & ~n58464;
  assign n58466 = ~n58462 & ~n58465;
  assign n58467 = ~controllable_hgrant6 & ~n58466;
  assign n58468 = ~n58447 & ~n58467;
  assign n58469 = controllable_hmaster3 & ~n58468;
  assign n58470 = controllable_hmaster3 & ~n58469;
  assign n58471 = i_hbusreq7 & ~n58470;
  assign n58472 = i_hbusreq8 & ~n58468;
  assign n58473 = controllable_hgrant6 & ~n10368;
  assign n58474 = i_hbusreq6 & ~n58466;
  assign n58475 = controllable_hgrant5 & ~n10361;
  assign n58476 = i_hbusreq5 & ~n58459;
  assign n58477 = controllable_hgrant4 & ~n10359;
  assign n58478 = i_hbusreq4 & ~n58457;
  assign n58479 = i_hbusreq9 & ~n58457;
  assign n58480 = controllable_hgrant3 & ~n10355;
  assign n58481 = i_hbusreq3 & ~n58455;
  assign n58482 = controllable_hgrant1 & ~n10353;
  assign n58483 = i_hbusreq1 & ~n58453;
  assign n58484 = ~n7871 & n7928;
  assign n58485 = n7928 & ~n58484;
  assign n58486 = ~i_hbusreq1 & ~n58485;
  assign n58487 = ~n58483 & ~n58486;
  assign n58488 = ~controllable_hgrant1 & ~n58487;
  assign n58489 = ~n58482 & ~n58488;
  assign n58490 = ~i_hbusreq3 & ~n58489;
  assign n58491 = ~n58481 & ~n58490;
  assign n58492 = ~controllable_hgrant3 & ~n58491;
  assign n58493 = ~n58480 & ~n58492;
  assign n58494 = ~i_hbusreq9 & ~n58493;
  assign n58495 = ~n58479 & ~n58494;
  assign n58496 = ~i_hbusreq4 & ~n58495;
  assign n58497 = ~n58478 & ~n58496;
  assign n58498 = ~controllable_hgrant4 & ~n58497;
  assign n58499 = ~n58477 & ~n58498;
  assign n58500 = ~i_hbusreq5 & ~n58499;
  assign n58501 = ~n58476 & ~n58500;
  assign n58502 = ~controllable_hgrant5 & ~n58501;
  assign n58503 = ~n58475 & ~n58502;
  assign n58504 = controllable_hmaster1 & ~n58503;
  assign n58505 = controllable_hmaster2 & ~n58503;
  assign n58506 = controllable_hmaster2 & ~n58505;
  assign n58507 = ~controllable_hmaster1 & ~n58506;
  assign n58508 = ~n58504 & ~n58507;
  assign n58509 = ~i_hbusreq6 & ~n58508;
  assign n58510 = ~n58474 & ~n58509;
  assign n58511 = ~controllable_hgrant6 & ~n58510;
  assign n58512 = ~n58473 & ~n58511;
  assign n58513 = ~i_hbusreq8 & ~n58512;
  assign n58514 = ~n58472 & ~n58513;
  assign n58515 = controllable_hmaster3 & ~n58514;
  assign n58516 = controllable_hmaster3 & ~n58515;
  assign n58517 = ~i_hbusreq7 & ~n58516;
  assign n58518 = ~n58471 & ~n58517;
  assign n58519 = ~n7924 & ~n58518;
  assign n58520 = controllable_hgrant6 & ~n10378;
  assign n58521 = ~n7822 & n7928;
  assign n58522 = n7928 & ~n58521;
  assign n58523 = ~controllable_hgrant1 & ~n58522;
  assign n58524 = ~n13179 & ~n58523;
  assign n58525 = ~controllable_hgrant3 & ~n58524;
  assign n58526 = ~n13178 & ~n58525;
  assign n58527 = ~controllable_hgrant4 & ~n58526;
  assign n58528 = ~n13177 & ~n58527;
  assign n58529 = ~controllable_hgrant5 & ~n58528;
  assign n58530 = ~n13176 & ~n58529;
  assign n58531 = controllable_hmaster1 & ~n58530;
  assign n58532 = controllable_hmaster2 & ~n58530;
  assign n58533 = controllable_hmaster2 & ~n58532;
  assign n58534 = ~controllable_hmaster1 & ~n58533;
  assign n58535 = ~n58531 & ~n58534;
  assign n58536 = ~controllable_hgrant6 & ~n58535;
  assign n58537 = ~n58520 & ~n58536;
  assign n58538 = controllable_hmaster3 & ~n58537;
  assign n58539 = controllable_hgrant6 & ~n10410;
  assign n58540 = controllable_hgrant5 & ~n10388;
  assign n58541 = controllable_hgrant4 & ~n10388;
  assign n58542 = ~n8365 & ~n23637;
  assign n58543 = ~n8365 & ~n58542;
  assign n58544 = i_hlock3 & ~n58543;
  assign n58545 = ~n8365 & ~n23645;
  assign n58546 = ~n8365 & ~n58545;
  assign n58547 = ~i_hlock3 & ~n58546;
  assign n58548 = ~n58544 & ~n58547;
  assign n58549 = controllable_hgrant3 & ~n58548;
  assign n58550 = ~controllable_hgrant3 & ~n10388;
  assign n58551 = ~n58549 & ~n58550;
  assign n58552 = ~controllable_hgrant4 & ~n58551;
  assign n58553 = ~n58541 & ~n58552;
  assign n58554 = ~controllable_hgrant5 & ~n58553;
  assign n58555 = ~n58540 & ~n58554;
  assign n58556 = ~controllable_hmaster2 & ~n58555;
  assign n58557 = ~controllable_hmaster2 & ~n58556;
  assign n58558 = controllable_hmaster1 & ~n58557;
  assign n58559 = ~n8378 & ~n33328;
  assign n58560 = ~n8378 & ~n58559;
  assign n58561 = i_hlock5 & ~n58560;
  assign n58562 = ~n8378 & ~n33346;
  assign n58563 = ~n8378 & ~n58562;
  assign n58564 = ~i_hlock5 & ~n58563;
  assign n58565 = ~n58561 & ~n58564;
  assign n58566 = controllable_hgrant5 & ~n58565;
  assign n58567 = ~controllable_hgrant5 & ~n10398;
  assign n58568 = ~n58566 & ~n58567;
  assign n58569 = controllable_hmaster2 & ~n58568;
  assign n58570 = controllable_hgrant5 & ~n10406;
  assign n58571 = controllable_hgrant4 & ~n10406;
  assign n58572 = controllable_hgrant3 & ~n10406;
  assign n58573 = ~n8389 & ~n23635;
  assign n58574 = ~n8389 & ~n58573;
  assign n58575 = i_hlock1 & ~n58574;
  assign n58576 = ~n8389 & ~n23643;
  assign n58577 = ~n8389 & ~n58576;
  assign n58578 = ~i_hlock1 & ~n58577;
  assign n58579 = ~n58575 & ~n58578;
  assign n58580 = controllable_hgrant1 & ~n58579;
  assign n58581 = ~controllable_hgrant1 & ~n10406;
  assign n58582 = ~n58580 & ~n58581;
  assign n58583 = ~controllable_hgrant3 & ~n58582;
  assign n58584 = ~n58572 & ~n58583;
  assign n58585 = ~controllable_hgrant4 & ~n58584;
  assign n58586 = ~n58571 & ~n58585;
  assign n58587 = ~controllable_hgrant5 & ~n58586;
  assign n58588 = ~n58570 & ~n58587;
  assign n58589 = ~controllable_hmaster2 & ~n58588;
  assign n58590 = ~n58569 & ~n58589;
  assign n58591 = ~controllable_hmaster1 & ~n58590;
  assign n58592 = ~n58558 & ~n58591;
  assign n58593 = ~controllable_hgrant6 & ~n58592;
  assign n58594 = ~n58539 & ~n58593;
  assign n58595 = controllable_hmaster0 & ~n58594;
  assign n58596 = ~n10413 & ~n33331;
  assign n58597 = controllable_hmaster1 & ~n58596;
  assign n58598 = ~n10427 & ~n58597;
  assign n58599 = ~n8217 & ~n58598;
  assign n58600 = ~n10429 & ~n58599;
  assign n58601 = i_hlock6 & ~n58600;
  assign n58602 = ~n10413 & ~n33349;
  assign n58603 = controllable_hmaster1 & ~n58602;
  assign n58604 = ~n10427 & ~n58603;
  assign n58605 = ~n8217 & ~n58604;
  assign n58606 = ~n10429 & ~n58605;
  assign n58607 = ~i_hlock6 & ~n58606;
  assign n58608 = ~n58601 & ~n58607;
  assign n58609 = controllable_hgrant6 & ~n58608;
  assign n58610 = controllable_hgrant5 & ~n10412;
  assign n58611 = controllable_hgrant4 & ~n10412;
  assign n58612 = controllable_hgrant3 & ~n10412;
  assign n58613 = controllable_hgrant1 & ~n10412;
  assign n58614 = n7928 & ~n39868;
  assign n58615 = ~controllable_hgrant1 & ~n58614;
  assign n58616 = ~n58613 & ~n58615;
  assign n58617 = ~controllable_hgrant3 & ~n58616;
  assign n58618 = ~n58612 & ~n58617;
  assign n58619 = ~controllable_hgrant4 & ~n58618;
  assign n58620 = ~n58611 & ~n58619;
  assign n58621 = ~controllable_hgrant5 & ~n58620;
  assign n58622 = ~n58610 & ~n58621;
  assign n58623 = ~controllable_hmaster2 & ~n58622;
  assign n58624 = ~controllable_hmaster2 & ~n58623;
  assign n58625 = controllable_hmaster1 & ~n58624;
  assign n58626 = controllable_hgrant5 & ~n10422;
  assign n58627 = ~n8426 & ~n23639;
  assign n58628 = ~n8426 & ~n58627;
  assign n58629 = i_hlock4 & ~n58628;
  assign n58630 = ~n8426 & ~n23647;
  assign n58631 = ~n8426 & ~n58630;
  assign n58632 = ~i_hlock4 & ~n58631;
  assign n58633 = ~n58629 & ~n58632;
  assign n58634 = controllable_hgrant4 & ~n58633;
  assign n58635 = ~controllable_hgrant4 & ~n10422;
  assign n58636 = ~n58634 & ~n58635;
  assign n58637 = ~controllable_hgrant5 & ~n58636;
  assign n58638 = ~n58626 & ~n58637;
  assign n58639 = controllable_hmaster2 & ~n58638;
  assign n58640 = ~n10425 & ~n58639;
  assign n58641 = ~controllable_hmaster1 & ~n58640;
  assign n58642 = ~n58625 & ~n58641;
  assign n58643 = n8217 & ~n58642;
  assign n58644 = ~n10430 & ~n58623;
  assign n58645 = controllable_hmaster1 & ~n58644;
  assign n58646 = ~n58641 & ~n58645;
  assign n58647 = ~n8217 & ~n58646;
  assign n58648 = ~n58643 & ~n58647;
  assign n58649 = i_hlock6 & ~n58648;
  assign n58650 = ~n10437 & ~n58623;
  assign n58651 = controllable_hmaster1 & ~n58650;
  assign n58652 = ~n58641 & ~n58651;
  assign n58653 = ~n8217 & ~n58652;
  assign n58654 = ~n58643 & ~n58653;
  assign n58655 = ~i_hlock6 & ~n58654;
  assign n58656 = ~n58649 & ~n58655;
  assign n58657 = ~controllable_hgrant6 & ~n58656;
  assign n58658 = ~n58609 & ~n58657;
  assign n58659 = ~controllable_hmaster0 & ~n58658;
  assign n58660 = ~n58595 & ~n58659;
  assign n58661 = ~controllable_hmaster3 & ~n58660;
  assign n58662 = ~n58538 & ~n58661;
  assign n58663 = i_hbusreq7 & ~n58662;
  assign n58664 = i_hbusreq8 & ~n58537;
  assign n58665 = controllable_hgrant6 & ~n10456;
  assign n58666 = i_hbusreq6 & ~n58535;
  assign n58667 = i_hbusreq5 & ~n58528;
  assign n58668 = i_hbusreq4 & ~n58526;
  assign n58669 = i_hbusreq9 & ~n58526;
  assign n58670 = i_hbusreq3 & ~n58524;
  assign n58671 = i_hbusreq1 & ~n58522;
  assign n58672 = ~n7869 & n7928;
  assign n58673 = n7928 & ~n58672;
  assign n58674 = ~i_hbusreq1 & ~n58673;
  assign n58675 = ~n58671 & ~n58674;
  assign n58676 = ~controllable_hgrant1 & ~n58675;
  assign n58677 = ~n13263 & ~n58676;
  assign n58678 = ~i_hbusreq3 & ~n58677;
  assign n58679 = ~n58670 & ~n58678;
  assign n58680 = ~controllable_hgrant3 & ~n58679;
  assign n58681 = ~n13261 & ~n58680;
  assign n58682 = ~i_hbusreq9 & ~n58681;
  assign n58683 = ~n58669 & ~n58682;
  assign n58684 = ~i_hbusreq4 & ~n58683;
  assign n58685 = ~n58668 & ~n58684;
  assign n58686 = ~controllable_hgrant4 & ~n58685;
  assign n58687 = ~n13258 & ~n58686;
  assign n58688 = ~i_hbusreq5 & ~n58687;
  assign n58689 = ~n58667 & ~n58688;
  assign n58690 = ~controllable_hgrant5 & ~n58689;
  assign n58691 = ~n13256 & ~n58690;
  assign n58692 = controllable_hmaster1 & ~n58691;
  assign n58693 = controllable_hmaster2 & ~n58691;
  assign n58694 = controllable_hmaster2 & ~n58693;
  assign n58695 = ~controllable_hmaster1 & ~n58694;
  assign n58696 = ~n58692 & ~n58695;
  assign n58697 = ~i_hbusreq6 & ~n58696;
  assign n58698 = ~n58666 & ~n58697;
  assign n58699 = ~controllable_hgrant6 & ~n58698;
  assign n58700 = ~n58665 & ~n58699;
  assign n58701 = ~i_hbusreq8 & ~n58700;
  assign n58702 = ~n58664 & ~n58701;
  assign n58703 = controllable_hmaster3 & ~n58702;
  assign n58704 = i_hbusreq8 & ~n58660;
  assign n58705 = controllable_hgrant6 & ~n10548;
  assign n58706 = i_hbusreq6 & ~n58592;
  assign n58707 = controllable_hgrant5 & ~n10488;
  assign n58708 = i_hbusreq5 & ~n58553;
  assign n58709 = controllable_hgrant4 & ~n10486;
  assign n58710 = i_hbusreq4 & ~n58551;
  assign n58711 = i_hbusreq9 & ~n58551;
  assign n58712 = i_hbusreq3 & ~n58548;
  assign n58713 = ~n8365 & ~n23681;
  assign n58714 = ~n8365 & ~n58713;
  assign n58715 = i_hlock3 & ~n58714;
  assign n58716 = ~n8365 & ~n23695;
  assign n58717 = ~n8365 & ~n58716;
  assign n58718 = ~i_hlock3 & ~n58717;
  assign n58719 = ~n58715 & ~n58718;
  assign n58720 = ~i_hbusreq3 & ~n58719;
  assign n58721 = ~n58712 & ~n58720;
  assign n58722 = controllable_hgrant3 & ~n58721;
  assign n58723 = ~controllable_hgrant3 & ~n10482;
  assign n58724 = ~n58722 & ~n58723;
  assign n58725 = ~i_hbusreq9 & ~n58724;
  assign n58726 = ~n58711 & ~n58725;
  assign n58727 = ~i_hbusreq4 & ~n58726;
  assign n58728 = ~n58710 & ~n58727;
  assign n58729 = ~controllable_hgrant4 & ~n58728;
  assign n58730 = ~n58709 & ~n58729;
  assign n58731 = ~i_hbusreq5 & ~n58730;
  assign n58732 = ~n58708 & ~n58731;
  assign n58733 = ~controllable_hgrant5 & ~n58732;
  assign n58734 = ~n58707 & ~n58733;
  assign n58735 = ~controllable_hmaster2 & ~n58734;
  assign n58736 = ~controllable_hmaster2 & ~n58735;
  assign n58737 = controllable_hmaster1 & ~n58736;
  assign n58738 = i_hbusreq5 & ~n58565;
  assign n58739 = ~n8378 & ~n33375;
  assign n58740 = ~n8378 & ~n58739;
  assign n58741 = i_hlock5 & ~n58740;
  assign n58742 = ~n8378 & ~n33408;
  assign n58743 = ~n8378 & ~n58742;
  assign n58744 = ~i_hlock5 & ~n58743;
  assign n58745 = ~n58741 & ~n58744;
  assign n58746 = ~i_hbusreq5 & ~n58745;
  assign n58747 = ~n58738 & ~n58746;
  assign n58748 = controllable_hgrant5 & ~n58747;
  assign n58749 = ~controllable_hgrant5 & ~n10519;
  assign n58750 = ~n58748 & ~n58749;
  assign n58751 = controllable_hmaster2 & ~n58750;
  assign n58752 = controllable_hgrant5 & ~n10542;
  assign n58753 = i_hbusreq5 & ~n58586;
  assign n58754 = controllable_hgrant4 & ~n10540;
  assign n58755 = i_hbusreq4 & ~n58584;
  assign n58756 = i_hbusreq9 & ~n58584;
  assign n58757 = controllable_hgrant3 & ~n10536;
  assign n58758 = i_hbusreq3 & ~n58582;
  assign n58759 = i_hbusreq1 & ~n58579;
  assign n58760 = ~n8389 & ~n23677;
  assign n58761 = ~n8389 & ~n58760;
  assign n58762 = i_hlock1 & ~n58761;
  assign n58763 = ~n8389 & ~n23691;
  assign n58764 = ~n8389 & ~n58763;
  assign n58765 = ~i_hlock1 & ~n58764;
  assign n58766 = ~n58762 & ~n58765;
  assign n58767 = ~i_hbusreq1 & ~n58766;
  assign n58768 = ~n58759 & ~n58767;
  assign n58769 = controllable_hgrant1 & ~n58768;
  assign n58770 = ~controllable_hgrant1 & ~n10534;
  assign n58771 = ~n58769 & ~n58770;
  assign n58772 = ~i_hbusreq3 & ~n58771;
  assign n58773 = ~n58758 & ~n58772;
  assign n58774 = ~controllable_hgrant3 & ~n58773;
  assign n58775 = ~n58757 & ~n58774;
  assign n58776 = ~i_hbusreq9 & ~n58775;
  assign n58777 = ~n58756 & ~n58776;
  assign n58778 = ~i_hbusreq4 & ~n58777;
  assign n58779 = ~n58755 & ~n58778;
  assign n58780 = ~controllable_hgrant4 & ~n58779;
  assign n58781 = ~n58754 & ~n58780;
  assign n58782 = ~i_hbusreq5 & ~n58781;
  assign n58783 = ~n58753 & ~n58782;
  assign n58784 = ~controllable_hgrant5 & ~n58783;
  assign n58785 = ~n58752 & ~n58784;
  assign n58786 = ~controllable_hmaster2 & ~n58785;
  assign n58787 = ~n58751 & ~n58786;
  assign n58788 = ~controllable_hmaster1 & ~n58787;
  assign n58789 = ~n58737 & ~n58788;
  assign n58790 = ~i_hbusreq6 & ~n58789;
  assign n58791 = ~n58706 & ~n58790;
  assign n58792 = ~controllable_hgrant6 & ~n58791;
  assign n58793 = ~n58705 & ~n58792;
  assign n58794 = controllable_hmaster0 & ~n58793;
  assign n58795 = i_hbusreq6 & ~n58608;
  assign n58796 = ~n10567 & ~n33380;
  assign n58797 = controllable_hmaster1 & ~n58796;
  assign n58798 = ~n10591 & ~n58797;
  assign n58799 = ~n8217 & ~n58798;
  assign n58800 = ~n10593 & ~n58799;
  assign n58801 = i_hlock6 & ~n58800;
  assign n58802 = ~n10567 & ~n33413;
  assign n58803 = controllable_hmaster1 & ~n58802;
  assign n58804 = ~n10591 & ~n58803;
  assign n58805 = ~n8217 & ~n58804;
  assign n58806 = ~n10593 & ~n58805;
  assign n58807 = ~i_hlock6 & ~n58806;
  assign n58808 = ~n58801 & ~n58807;
  assign n58809 = ~i_hbusreq6 & ~n58808;
  assign n58810 = ~n58795 & ~n58809;
  assign n58811 = controllable_hgrant6 & ~n58810;
  assign n58812 = i_hbusreq6 & ~n58656;
  assign n58813 = controllable_hgrant5 & ~n10566;
  assign n58814 = i_hbusreq5 & ~n58620;
  assign n58815 = controllable_hgrant4 & ~n10564;
  assign n58816 = i_hbusreq4 & ~n58618;
  assign n58817 = i_hbusreq9 & ~n58618;
  assign n58818 = controllable_hgrant3 & ~n10560;
  assign n58819 = i_hbusreq3 & ~n58616;
  assign n58820 = controllable_hgrant1 & ~n10558;
  assign n58821 = i_hbusreq1 & ~n58614;
  assign n58822 = n7928 & ~n40097;
  assign n58823 = ~i_hbusreq1 & ~n58822;
  assign n58824 = ~n58821 & ~n58823;
  assign n58825 = ~controllable_hgrant1 & ~n58824;
  assign n58826 = ~n58820 & ~n58825;
  assign n58827 = ~i_hbusreq3 & ~n58826;
  assign n58828 = ~n58819 & ~n58827;
  assign n58829 = ~controllable_hgrant3 & ~n58828;
  assign n58830 = ~n58818 & ~n58829;
  assign n58831 = ~i_hbusreq9 & ~n58830;
  assign n58832 = ~n58817 & ~n58831;
  assign n58833 = ~i_hbusreq4 & ~n58832;
  assign n58834 = ~n58816 & ~n58833;
  assign n58835 = ~controllable_hgrant4 & ~n58834;
  assign n58836 = ~n58815 & ~n58835;
  assign n58837 = ~i_hbusreq5 & ~n58836;
  assign n58838 = ~n58814 & ~n58837;
  assign n58839 = ~controllable_hgrant5 & ~n58838;
  assign n58840 = ~n58813 & ~n58839;
  assign n58841 = ~controllable_hmaster2 & ~n58840;
  assign n58842 = ~controllable_hmaster2 & ~n58841;
  assign n58843 = controllable_hmaster1 & ~n58842;
  assign n58844 = controllable_hgrant5 & ~n10588;
  assign n58845 = i_hbusreq5 & ~n58636;
  assign n58846 = i_hbusreq4 & ~n58633;
  assign n58847 = i_hbusreq9 & ~n58628;
  assign n58848 = ~n8426 & ~n23685;
  assign n58849 = ~n8426 & ~n58848;
  assign n58850 = ~i_hbusreq9 & ~n58849;
  assign n58851 = ~n58847 & ~n58850;
  assign n58852 = i_hlock4 & ~n58851;
  assign n58853 = i_hbusreq9 & ~n58631;
  assign n58854 = ~n8426 & ~n23699;
  assign n58855 = ~n8426 & ~n58854;
  assign n58856 = ~i_hbusreq9 & ~n58855;
  assign n58857 = ~n58853 & ~n58856;
  assign n58858 = ~i_hlock4 & ~n58857;
  assign n58859 = ~n58852 & ~n58858;
  assign n58860 = ~i_hbusreq4 & ~n58859;
  assign n58861 = ~n58846 & ~n58860;
  assign n58862 = controllable_hgrant4 & ~n58861;
  assign n58863 = ~controllable_hgrant4 & ~n10586;
  assign n58864 = ~n58862 & ~n58863;
  assign n58865 = ~i_hbusreq5 & ~n58864;
  assign n58866 = ~n58845 & ~n58865;
  assign n58867 = ~controllable_hgrant5 & ~n58866;
  assign n58868 = ~n58844 & ~n58867;
  assign n58869 = controllable_hmaster2 & ~n58868;
  assign n58870 = ~n10425 & ~n58869;
  assign n58871 = ~controllable_hmaster1 & ~n58870;
  assign n58872 = ~n58843 & ~n58871;
  assign n58873 = n8217 & ~n58872;
  assign n58874 = ~n10597 & ~n58841;
  assign n58875 = controllable_hmaster1 & ~n58874;
  assign n58876 = ~n58871 & ~n58875;
  assign n58877 = ~n8217 & ~n58876;
  assign n58878 = ~n58873 & ~n58877;
  assign n58879 = i_hlock6 & ~n58878;
  assign n58880 = ~n10607 & ~n58841;
  assign n58881 = controllable_hmaster1 & ~n58880;
  assign n58882 = ~n58871 & ~n58881;
  assign n58883 = ~n8217 & ~n58882;
  assign n58884 = ~n58873 & ~n58883;
  assign n58885 = ~i_hlock6 & ~n58884;
  assign n58886 = ~n58879 & ~n58885;
  assign n58887 = ~i_hbusreq6 & ~n58886;
  assign n58888 = ~n58812 & ~n58887;
  assign n58889 = ~controllable_hgrant6 & ~n58888;
  assign n58890 = ~n58811 & ~n58889;
  assign n58891 = ~controllable_hmaster0 & ~n58890;
  assign n58892 = ~n58794 & ~n58891;
  assign n58893 = ~i_hbusreq8 & ~n58892;
  assign n58894 = ~n58704 & ~n58893;
  assign n58895 = ~controllable_hmaster3 & ~n58894;
  assign n58896 = ~n58703 & ~n58895;
  assign n58897 = ~i_hbusreq7 & ~n58896;
  assign n58898 = ~n58663 & ~n58897;
  assign n58899 = n7924 & ~n58898;
  assign n58900 = ~n58519 & ~n58899;
  assign n58901 = n8214 & ~n58900;
  assign n58902 = n8214 & ~n58901;
  assign n58903 = n8202 & ~n58902;
  assign n58904 = ~n58446 & ~n58903;
  assign n58905 = n7728 & ~n58904;
  assign n58906 = ~n7840 & ~n58421;
  assign n58907 = i_hbusreq7 & ~n58906;
  assign n58908 = ~n7901 & ~n58438;
  assign n58909 = ~i_hbusreq7 & ~n58908;
  assign n58910 = ~n58907 & ~n58909;
  assign n58911 = n7924 & ~n58910;
  assign n58912 = ~n39731 & ~n58911;
  assign n58913 = ~n8214 & ~n58912;
  assign n58914 = ~n7840 & ~n10326;
  assign n58915 = i_hbusreq7 & ~n58914;
  assign n58916 = ~n7901 & ~n10326;
  assign n58917 = ~i_hbusreq7 & ~n58916;
  assign n58918 = ~n58915 & ~n58917;
  assign n58919 = n7924 & ~n58918;
  assign n58920 = ~n39731 & ~n58919;
  assign n58921 = n8214 & ~n58920;
  assign n58922 = ~n58913 & ~n58921;
  assign n58923 = ~n8202 & ~n58922;
  assign n58924 = n8214 & ~n40176;
  assign n58925 = ~n39730 & ~n58924;
  assign n58926 = n8202 & ~n58925;
  assign n58927 = ~n58923 & ~n58926;
  assign n58928 = ~n7728 & ~n58927;
  assign n58929 = ~n58905 & ~n58928;
  assign n58930 = ~n7723 & ~n58929;
  assign n58931 = ~n7723 & ~n58930;
  assign n58932 = ~n7714 & ~n58931;
  assign n58933 = ~n7714 & ~n58932;
  assign n58934 = n7705 & ~n58933;
  assign n58935 = n7723 & ~n58927;
  assign n58936 = n7920 & ~n58927;
  assign n58937 = ~n40177 & ~n58936;
  assign n58938 = ~n7723 & ~n58937;
  assign n58939 = ~n58935 & ~n58938;
  assign n58940 = n7714 & ~n58939;
  assign n58941 = ~n40183 & ~n58940;
  assign n58942 = ~n7705 & ~n58941;
  assign n58943 = ~n58934 & ~n58942;
  assign n58944 = ~n7808 & ~n58943;
  assign n58945 = ~n7920 & ~n58904;
  assign n58946 = n8217 & ~n10674;
  assign n58947 = ~n8217 & ~n23760;
  assign n58948 = ~n58946 & ~n58947;
  assign n58949 = controllable_hgrant6 & ~n58948;
  assign n58950 = ~controllable_hmaster2 & ~n48126;
  assign n58951 = ~controllable_hmaster1 & ~n58950;
  assign n58952 = ~controllable_hmaster1 & ~n58951;
  assign n58953 = ~controllable_hgrant6 & ~n58952;
  assign n58954 = ~n58949 & ~n58953;
  assign n58955 = controllable_hmaster0 & ~n58954;
  assign n58956 = controllable_hmaster0 & ~n58955;
  assign n58957 = ~controllable_hmaster3 & ~n58956;
  assign n58958 = ~controllable_hmaster3 & ~n58957;
  assign n58959 = i_hbusreq7 & ~n58958;
  assign n58960 = i_hbusreq8 & ~n58956;
  assign n58961 = i_hbusreq6 & ~n58948;
  assign n58962 = n8217 & ~n10684;
  assign n58963 = ~n8217 & ~n23773;
  assign n58964 = ~n58962 & ~n58963;
  assign n58965 = ~i_hbusreq6 & ~n58964;
  assign n58966 = ~n58961 & ~n58965;
  assign n58967 = controllable_hgrant6 & ~n58966;
  assign n58968 = i_hbusreq6 & ~n58952;
  assign n58969 = ~controllable_hmaster2 & ~n48496;
  assign n58970 = ~controllable_hmaster1 & ~n58969;
  assign n58971 = ~controllable_hmaster1 & ~n58970;
  assign n58972 = ~i_hbusreq6 & ~n58971;
  assign n58973 = ~n58968 & ~n58972;
  assign n58974 = ~controllable_hgrant6 & ~n58973;
  assign n58975 = ~n58967 & ~n58974;
  assign n58976 = controllable_hmaster0 & ~n58975;
  assign n58977 = controllable_hmaster0 & ~n58976;
  assign n58978 = ~i_hbusreq8 & ~n58977;
  assign n58979 = ~n58960 & ~n58978;
  assign n58980 = ~controllable_hmaster3 & ~n58979;
  assign n58981 = ~controllable_hmaster3 & ~n58980;
  assign n58982 = ~i_hbusreq7 & ~n58981;
  assign n58983 = ~n58959 & ~n58982;
  assign n58984 = ~n7924 & ~n58983;
  assign n58985 = n8389 & ~n12788;
  assign n58986 = ~n8389 & ~n16477;
  assign n58987 = ~n58985 & ~n58986;
  assign n58988 = i_hlock1 & ~n58987;
  assign n58989 = ~n8389 & ~n16491;
  assign n58990 = ~n58985 & ~n58989;
  assign n58991 = ~i_hlock1 & ~n58990;
  assign n58992 = ~n58988 & ~n58991;
  assign n58993 = controllable_hgrant1 & ~n58992;
  assign n58994 = controllable_hgrant1 & ~n58993;
  assign n58995 = ~controllable_hgrant3 & ~n58994;
  assign n58996 = ~controllable_hgrant3 & ~n58995;
  assign n58997 = ~controllable_hgrant4 & ~n58996;
  assign n58998 = ~controllable_hgrant4 & ~n58997;
  assign n58999 = ~controllable_hgrant5 & ~n58998;
  assign n59000 = ~controllable_hgrant5 & ~n58999;
  assign n59001 = ~controllable_hgrant6 & ~n59000;
  assign n59002 = ~controllable_hgrant6 & ~n59001;
  assign n59003 = controllable_hmaster3 & ~n59002;
  assign n59004 = controllable_hmaster1 & ~n59000;
  assign n59005 = controllable_hmaster2 & ~n59000;
  assign n59006 = ~n48118 & ~n48917;
  assign n59007 = ~controllable_hgrant3 & ~n59006;
  assign n59008 = ~n48106 & ~n59007;
  assign n59009 = ~controllable_hgrant4 & ~n59008;
  assign n59010 = ~n48103 & ~n59009;
  assign n59011 = ~controllable_hgrant5 & ~n59010;
  assign n59012 = ~n48100 & ~n59011;
  assign n59013 = ~controllable_hmaster2 & ~n59012;
  assign n59014 = ~n59005 & ~n59013;
  assign n59015 = ~controllable_hmaster1 & ~n59014;
  assign n59016 = ~n59004 & ~n59015;
  assign n59017 = ~controllable_hgrant6 & ~n59016;
  assign n59018 = ~n58949 & ~n59017;
  assign n59019 = controllable_hmaster0 & ~n59018;
  assign n59020 = ~controllable_hmaster0 & ~n59002;
  assign n59021 = ~n59019 & ~n59020;
  assign n59022 = ~controllable_hmaster3 & ~n59021;
  assign n59023 = ~n59003 & ~n59022;
  assign n59024 = i_hbusreq7 & ~n59023;
  assign n59025 = i_hbusreq8 & ~n59002;
  assign n59026 = i_hbusreq6 & ~n59000;
  assign n59027 = i_hbusreq5 & ~n58998;
  assign n59028 = i_hbusreq4 & ~n58996;
  assign n59029 = i_hbusreq9 & ~n58996;
  assign n59030 = i_hbusreq3 & ~n58994;
  assign n59031 = i_hbusreq1 & ~n58992;
  assign n59032 = n8389 & ~n12857;
  assign n59033 = ~n8389 & ~n16581;
  assign n59034 = ~n59032 & ~n59033;
  assign n59035 = i_hlock1 & ~n59034;
  assign n59036 = ~n8389 & ~n16595;
  assign n59037 = ~n59032 & ~n59036;
  assign n59038 = ~i_hlock1 & ~n59037;
  assign n59039 = ~n59035 & ~n59038;
  assign n59040 = ~i_hbusreq1 & ~n59039;
  assign n59041 = ~n59031 & ~n59040;
  assign n59042 = controllable_hgrant1 & ~n59041;
  assign n59043 = controllable_hgrant1 & ~n59042;
  assign n59044 = ~i_hbusreq3 & ~n59043;
  assign n59045 = ~n59030 & ~n59044;
  assign n59046 = ~controllable_hgrant3 & ~n59045;
  assign n59047 = ~controllable_hgrant3 & ~n59046;
  assign n59048 = ~i_hbusreq9 & ~n59047;
  assign n59049 = ~n59029 & ~n59048;
  assign n59050 = ~i_hbusreq4 & ~n59049;
  assign n59051 = ~n59028 & ~n59050;
  assign n59052 = ~controllable_hgrant4 & ~n59051;
  assign n59053 = ~controllable_hgrant4 & ~n59052;
  assign n59054 = ~i_hbusreq5 & ~n59053;
  assign n59055 = ~n59027 & ~n59054;
  assign n59056 = ~controllable_hgrant5 & ~n59055;
  assign n59057 = ~controllable_hgrant5 & ~n59056;
  assign n59058 = ~i_hbusreq6 & ~n59057;
  assign n59059 = ~n59026 & ~n59058;
  assign n59060 = ~controllable_hgrant6 & ~n59059;
  assign n59061 = ~controllable_hgrant6 & ~n59060;
  assign n59062 = ~i_hbusreq8 & ~n59061;
  assign n59063 = ~n59025 & ~n59062;
  assign n59064 = controllable_hmaster3 & ~n59063;
  assign n59065 = i_hbusreq8 & ~n59021;
  assign n59066 = i_hbusreq6 & ~n59016;
  assign n59067 = controllable_hmaster1 & ~n59057;
  assign n59068 = controllable_hmaster2 & ~n59057;
  assign n59069 = i_hbusreq5 & ~n59010;
  assign n59070 = i_hbusreq4 & ~n59008;
  assign n59071 = i_hbusreq9 & ~n59008;
  assign n59072 = i_hbusreq3 & ~n59006;
  assign n59073 = ~n48480 & ~n49636;
  assign n59074 = ~i_hbusreq3 & ~n59073;
  assign n59075 = ~n59072 & ~n59074;
  assign n59076 = ~controllable_hgrant3 & ~n59075;
  assign n59077 = ~n48459 & ~n59076;
  assign n59078 = ~i_hbusreq9 & ~n59077;
  assign n59079 = ~n59071 & ~n59078;
  assign n59080 = ~i_hbusreq4 & ~n59079;
  assign n59081 = ~n59070 & ~n59080;
  assign n59082 = ~controllable_hgrant4 & ~n59081;
  assign n59083 = ~n48450 & ~n59082;
  assign n59084 = ~i_hbusreq5 & ~n59083;
  assign n59085 = ~n59069 & ~n59084;
  assign n59086 = ~controllable_hgrant5 & ~n59085;
  assign n59087 = ~n48439 & ~n59086;
  assign n59088 = ~controllable_hmaster2 & ~n59087;
  assign n59089 = ~n59068 & ~n59088;
  assign n59090 = ~controllable_hmaster1 & ~n59089;
  assign n59091 = ~n59067 & ~n59090;
  assign n59092 = ~i_hbusreq6 & ~n59091;
  assign n59093 = ~n59066 & ~n59092;
  assign n59094 = ~controllable_hgrant6 & ~n59093;
  assign n59095 = ~n58967 & ~n59094;
  assign n59096 = controllable_hmaster0 & ~n59095;
  assign n59097 = ~controllable_hmaster0 & ~n59061;
  assign n59098 = ~n59096 & ~n59097;
  assign n59099 = ~i_hbusreq8 & ~n59098;
  assign n59100 = ~n59065 & ~n59099;
  assign n59101 = ~controllable_hmaster3 & ~n59100;
  assign n59102 = ~n59064 & ~n59101;
  assign n59103 = ~i_hbusreq7 & ~n59102;
  assign n59104 = ~n59024 & ~n59103;
  assign n59105 = n7924 & ~n59104;
  assign n59106 = ~n58984 & ~n59105;
  assign n59107 = ~n8214 & ~n59106;
  assign n59108 = n8217 & ~n10698;
  assign n59109 = ~n8217 & ~n23790;
  assign n59110 = ~n59108 & ~n59109;
  assign n59111 = controllable_hgrant6 & ~n59110;
  assign n59112 = ~controllable_hmaster2 & ~n48207;
  assign n59113 = ~controllable_hmaster1 & ~n59112;
  assign n59114 = ~controllable_hmaster1 & ~n59113;
  assign n59115 = ~controllable_hgrant6 & ~n59114;
  assign n59116 = ~n59111 & ~n59115;
  assign n59117 = ~controllable_hmaster0 & ~n59116;
  assign n59118 = ~controllable_hmaster0 & ~n59117;
  assign n59119 = ~controllable_hmaster3 & ~n59118;
  assign n59120 = ~controllable_hmaster3 & ~n59119;
  assign n59121 = i_hbusreq7 & ~n59120;
  assign n59122 = i_hbusreq8 & ~n59118;
  assign n59123 = i_hbusreq6 & ~n59110;
  assign n59124 = n8217 & ~n10708;
  assign n59125 = ~n8217 & ~n23803;
  assign n59126 = ~n59124 & ~n59125;
  assign n59127 = ~i_hbusreq6 & ~n59126;
  assign n59128 = ~n59123 & ~n59127;
  assign n59129 = controllable_hgrant6 & ~n59128;
  assign n59130 = i_hbusreq6 & ~n59114;
  assign n59131 = ~controllable_hmaster2 & ~n48715;
  assign n59132 = ~controllable_hmaster1 & ~n59131;
  assign n59133 = ~controllable_hmaster1 & ~n59132;
  assign n59134 = ~i_hbusreq6 & ~n59133;
  assign n59135 = ~n59130 & ~n59134;
  assign n59136 = ~controllable_hgrant6 & ~n59135;
  assign n59137 = ~n59129 & ~n59136;
  assign n59138 = ~controllable_hmaster0 & ~n59137;
  assign n59139 = ~controllable_hmaster0 & ~n59138;
  assign n59140 = ~i_hbusreq8 & ~n59139;
  assign n59141 = ~n59122 & ~n59140;
  assign n59142 = ~controllable_hmaster3 & ~n59141;
  assign n59143 = ~controllable_hmaster3 & ~n59142;
  assign n59144 = ~i_hbusreq7 & ~n59143;
  assign n59145 = ~n59121 & ~n59144;
  assign n59146 = n8214 & ~n59145;
  assign n59147 = ~n59107 & ~n59146;
  assign n59148 = ~n8202 & ~n59147;
  assign n59149 = n7924 & ~n49999;
  assign n59150 = ~n8214 & ~n59149;
  assign n59151 = ~n8217 & ~n23851;
  assign n59152 = ~n42489 & ~n59151;
  assign n59153 = controllable_hgrant6 & ~n59152;
  assign n59154 = ~n8378 & ~n23828;
  assign n59155 = ~n51657 & ~n59154;
  assign n59156 = controllable_hgrant5 & ~n59155;
  assign n59157 = ~n8426 & ~n23826;
  assign n59158 = ~n51941 & ~n59157;
  assign n59159 = controllable_hgrant4 & ~n59158;
  assign n59160 = ~n8365 & ~n23824;
  assign n59161 = ~n52337 & ~n59160;
  assign n59162 = controllable_hgrant3 & ~n59161;
  assign n59163 = n8389 & ~n8987;
  assign n59164 = ~n8389 & ~n23822;
  assign n59165 = ~n59163 & ~n59164;
  assign n59166 = controllable_hgrant1 & ~n59165;
  assign n59167 = n7928 & ~n48023;
  assign n59168 = n7928 & ~n59167;
  assign n59169 = ~controllable_hgrant1 & ~n59168;
  assign n59170 = ~n59166 & ~n59169;
  assign n59171 = ~controllable_hgrant3 & ~n59170;
  assign n59172 = ~n59162 & ~n59171;
  assign n59173 = ~controllable_hgrant4 & ~n59172;
  assign n59174 = ~n59159 & ~n59173;
  assign n59175 = ~controllable_hgrant5 & ~n59174;
  assign n59176 = ~n59156 & ~n59175;
  assign n59177 = controllable_hmaster1 & ~n59176;
  assign n59178 = controllable_hmaster2 & ~n59176;
  assign n59179 = ~n8389 & ~n17331;
  assign n59180 = ~n59163 & ~n59179;
  assign n59181 = controllable_hgrant1 & ~n59180;
  assign n59182 = n7928 & ~n40230;
  assign n59183 = ~controllable_hgrant1 & ~n59182;
  assign n59184 = ~n59181 & ~n59183;
  assign n59185 = ~controllable_hgrant3 & ~n59184;
  assign n59186 = ~n52340 & ~n59185;
  assign n59187 = ~controllable_hgrant4 & ~n59186;
  assign n59188 = ~n51944 & ~n59187;
  assign n59189 = ~controllable_hgrant5 & ~n59188;
  assign n59190 = ~n51660 & ~n59189;
  assign n59191 = ~controllable_hmaster2 & ~n59190;
  assign n59192 = ~n59178 & ~n59191;
  assign n59193 = ~controllable_hmaster1 & ~n59192;
  assign n59194 = ~n59177 & ~n59193;
  assign n59195 = ~controllable_hgrant6 & ~n59194;
  assign n59196 = ~n59153 & ~n59195;
  assign n59197 = controllable_hmaster3 & ~n59196;
  assign n59198 = controllable_hmaster2 & ~n59190;
  assign n59199 = n8365 & ~n13315;
  assign n59200 = ~n8365 & ~n23835;
  assign n59201 = ~n59199 & ~n59200;
  assign n59202 = controllable_hgrant3 & ~n59201;
  assign n59203 = ~n59185 & ~n59202;
  assign n59204 = ~controllable_hgrant4 & ~n59203;
  assign n59205 = ~n51944 & ~n59204;
  assign n59206 = ~controllable_hgrant5 & ~n59205;
  assign n59207 = ~n51660 & ~n59206;
  assign n59208 = ~controllable_hmaster2 & ~n59207;
  assign n59209 = ~n59198 & ~n59208;
  assign n59210 = controllable_hmaster1 & ~n59209;
  assign n59211 = n8378 & ~n13319;
  assign n59212 = ~n8378 & ~n23839;
  assign n59213 = ~n59211 & ~n59212;
  assign n59214 = controllable_hgrant5 & ~n59213;
  assign n59215 = ~n59189 & ~n59214;
  assign n59216 = controllable_hmaster2 & ~n59215;
  assign n59217 = n8389 & ~n13313;
  assign n59218 = ~n8389 & ~n23833;
  assign n59219 = ~n59217 & ~n59218;
  assign n59220 = controllable_hgrant1 & ~n59219;
  assign n59221 = ~n59183 & ~n59220;
  assign n59222 = ~controllable_hgrant3 & ~n59221;
  assign n59223 = ~n52340 & ~n59222;
  assign n59224 = ~controllable_hgrant4 & ~n59223;
  assign n59225 = ~n51944 & ~n59224;
  assign n59226 = ~controllable_hgrant5 & ~n59225;
  assign n59227 = ~n51660 & ~n59226;
  assign n59228 = ~controllable_hmaster2 & ~n59227;
  assign n59229 = ~n59216 & ~n59228;
  assign n59230 = ~controllable_hmaster1 & ~n59229;
  assign n59231 = ~n59210 & ~n59230;
  assign n59232 = ~controllable_hgrant6 & ~n59231;
  assign n59233 = ~n42492 & ~n59232;
  assign n59234 = controllable_hmaster0 & ~n59233;
  assign n59235 = n8217 & ~n26891;
  assign n59236 = ~n8217 & ~n33466;
  assign n59237 = ~n59235 & ~n59236;
  assign n59238 = controllable_hgrant6 & ~n59237;
  assign n59239 = n7928 & ~n48154;
  assign n59240 = ~controllable_hgrant1 & ~n59239;
  assign n59241 = ~n59181 & ~n59240;
  assign n59242 = ~controllable_hgrant3 & ~n59241;
  assign n59243 = ~n52340 & ~n59242;
  assign n59244 = ~controllable_hgrant4 & ~n59243;
  assign n59245 = ~n51944 & ~n59244;
  assign n59246 = ~controllable_hgrant5 & ~n59245;
  assign n59247 = ~n51660 & ~n59246;
  assign n59248 = ~controllable_hmaster2 & ~n59247;
  assign n59249 = ~n59198 & ~n59248;
  assign n59250 = controllable_hmaster1 & ~n59249;
  assign n59251 = n8426 & ~n13317;
  assign n59252 = ~n8426 & ~n23837;
  assign n59253 = ~n59251 & ~n59252;
  assign n59254 = controllable_hgrant4 & ~n59253;
  assign n59255 = ~n59187 & ~n59254;
  assign n59256 = ~controllable_hgrant5 & ~n59255;
  assign n59257 = ~n51660 & ~n59256;
  assign n59258 = controllable_hmaster2 & ~n59257;
  assign n59259 = ~n59191 & ~n59258;
  assign n59260 = ~controllable_hmaster1 & ~n59259;
  assign n59261 = ~n59250 & ~n59260;
  assign n59262 = ~controllable_hgrant6 & ~n59261;
  assign n59263 = ~n59238 & ~n59262;
  assign n59264 = ~controllable_hmaster0 & ~n59263;
  assign n59265 = ~n59234 & ~n59264;
  assign n59266 = ~controllable_hmaster3 & ~n59265;
  assign n59267 = ~n59197 & ~n59266;
  assign n59268 = i_hbusreq7 & ~n59267;
  assign n59269 = i_hbusreq8 & ~n59196;
  assign n59270 = i_hbusreq6 & ~n59152;
  assign n59271 = n8217 & ~n10754;
  assign n59272 = ~n8217 & ~n23944;
  assign n59273 = ~n59271 & ~n59272;
  assign n59274 = ~i_hbusreq6 & ~n59273;
  assign n59275 = ~n59270 & ~n59274;
  assign n59276 = controllable_hgrant6 & ~n59275;
  assign n59277 = i_hbusreq6 & ~n59194;
  assign n59278 = i_hbusreq5 & ~n59155;
  assign n59279 = n8378 & ~n10735;
  assign n59280 = ~n8378 & ~n23881;
  assign n59281 = ~n59279 & ~n59280;
  assign n59282 = ~i_hbusreq5 & ~n59281;
  assign n59283 = ~n59278 & ~n59282;
  assign n59284 = controllable_hgrant5 & ~n59283;
  assign n59285 = i_hbusreq5 & ~n59174;
  assign n59286 = i_hbusreq4 & ~n59158;
  assign n59287 = i_hbusreq9 & ~n59158;
  assign n59288 = n8426 & ~n10731;
  assign n59289 = ~n8426 & ~n23875;
  assign n59290 = ~n59288 & ~n59289;
  assign n59291 = ~i_hbusreq9 & ~n59290;
  assign n59292 = ~n59287 & ~n59291;
  assign n59293 = ~i_hbusreq4 & ~n59292;
  assign n59294 = ~n59286 & ~n59293;
  assign n59295 = controllable_hgrant4 & ~n59294;
  assign n59296 = i_hbusreq4 & ~n59172;
  assign n59297 = i_hbusreq9 & ~n59172;
  assign n59298 = i_hbusreq3 & ~n59161;
  assign n59299 = n8365 & ~n10729;
  assign n59300 = ~n8365 & ~n23871;
  assign n59301 = ~n59299 & ~n59300;
  assign n59302 = ~i_hbusreq3 & ~n59301;
  assign n59303 = ~n59298 & ~n59302;
  assign n59304 = controllable_hgrant3 & ~n59303;
  assign n59305 = i_hbusreq3 & ~n59170;
  assign n59306 = i_hbusreq1 & ~n59165;
  assign n59307 = n8389 & ~n10727;
  assign n59308 = ~n8389 & ~n23867;
  assign n59309 = ~n59307 & ~n59308;
  assign n59310 = ~i_hbusreq1 & ~n59309;
  assign n59311 = ~n59306 & ~n59310;
  assign n59312 = controllable_hgrant1 & ~n59311;
  assign n59313 = i_hbusreq1 & ~n59168;
  assign n59314 = n7928 & ~n48282;
  assign n59315 = n7928 & ~n59314;
  assign n59316 = ~i_hbusreq1 & ~n59315;
  assign n59317 = ~n59313 & ~n59316;
  assign n59318 = ~controllable_hgrant1 & ~n59317;
  assign n59319 = ~n59312 & ~n59318;
  assign n59320 = ~i_hbusreq3 & ~n59319;
  assign n59321 = ~n59305 & ~n59320;
  assign n59322 = ~controllable_hgrant3 & ~n59321;
  assign n59323 = ~n59304 & ~n59322;
  assign n59324 = ~i_hbusreq9 & ~n59323;
  assign n59325 = ~n59297 & ~n59324;
  assign n59326 = ~i_hbusreq4 & ~n59325;
  assign n59327 = ~n59296 & ~n59326;
  assign n59328 = ~controllable_hgrant4 & ~n59327;
  assign n59329 = ~n59295 & ~n59328;
  assign n59330 = ~i_hbusreq5 & ~n59329;
  assign n59331 = ~n59285 & ~n59330;
  assign n59332 = ~controllable_hgrant5 & ~n59331;
  assign n59333 = ~n59284 & ~n59332;
  assign n59334 = controllable_hmaster1 & ~n59333;
  assign n59335 = controllable_hmaster2 & ~n59333;
  assign n59336 = n8378 & ~n10748;
  assign n59337 = ~n8378 & ~n23936;
  assign n59338 = ~n59336 & ~n59337;
  assign n59339 = ~i_hbusreq5 & ~n59338;
  assign n59340 = ~n51713 & ~n59339;
  assign n59341 = controllable_hgrant5 & ~n59340;
  assign n59342 = i_hbusreq5 & ~n59188;
  assign n59343 = n8426 & ~n10744;
  assign n59344 = ~n8426 & ~n23930;
  assign n59345 = ~n59343 & ~n59344;
  assign n59346 = ~i_hbusreq9 & ~n59345;
  assign n59347 = ~n52016 & ~n59346;
  assign n59348 = ~i_hbusreq4 & ~n59347;
  assign n59349 = ~n52015 & ~n59348;
  assign n59350 = controllable_hgrant4 & ~n59349;
  assign n59351 = i_hbusreq4 & ~n59186;
  assign n59352 = i_hbusreq9 & ~n59186;
  assign n59353 = n8365 & ~n10742;
  assign n59354 = ~n8365 & ~n23926;
  assign n59355 = ~n59353 & ~n59354;
  assign n59356 = ~i_hbusreq3 & ~n59355;
  assign n59357 = ~n52423 & ~n59356;
  assign n59358 = controllable_hgrant3 & ~n59357;
  assign n59359 = i_hbusreq3 & ~n59184;
  assign n59360 = i_hbusreq1 & ~n59180;
  assign n59361 = n8389 & ~n10740;
  assign n59362 = ~n8389 & ~n23922;
  assign n59363 = ~n59361 & ~n59362;
  assign n59364 = ~i_hbusreq1 & ~n59363;
  assign n59365 = ~n59360 & ~n59364;
  assign n59366 = controllable_hgrant1 & ~n59365;
  assign n59367 = i_hbusreq1 & ~n59182;
  assign n59368 = n7928 & ~n40359;
  assign n59369 = ~i_hbusreq1 & ~n59368;
  assign n59370 = ~n59367 & ~n59369;
  assign n59371 = ~controllable_hgrant1 & ~n59370;
  assign n59372 = ~n59366 & ~n59371;
  assign n59373 = ~i_hbusreq3 & ~n59372;
  assign n59374 = ~n59359 & ~n59373;
  assign n59375 = ~controllable_hgrant3 & ~n59374;
  assign n59376 = ~n59358 & ~n59375;
  assign n59377 = ~i_hbusreq9 & ~n59376;
  assign n59378 = ~n59352 & ~n59377;
  assign n59379 = ~i_hbusreq4 & ~n59378;
  assign n59380 = ~n59351 & ~n59379;
  assign n59381 = ~controllable_hgrant4 & ~n59380;
  assign n59382 = ~n59350 & ~n59381;
  assign n59383 = ~i_hbusreq5 & ~n59382;
  assign n59384 = ~n59342 & ~n59383;
  assign n59385 = ~controllable_hgrant5 & ~n59384;
  assign n59386 = ~n59341 & ~n59385;
  assign n59387 = ~controllable_hmaster2 & ~n59386;
  assign n59388 = ~n59335 & ~n59387;
  assign n59389 = ~controllable_hmaster1 & ~n59388;
  assign n59390 = ~n59334 & ~n59389;
  assign n59391 = ~i_hbusreq6 & ~n59390;
  assign n59392 = ~n59277 & ~n59391;
  assign n59393 = ~controllable_hgrant6 & ~n59392;
  assign n59394 = ~n59276 & ~n59393;
  assign n59395 = ~i_hbusreq8 & ~n59394;
  assign n59396 = ~n59269 & ~n59395;
  assign n59397 = controllable_hmaster3 & ~n59396;
  assign n59398 = i_hbusreq8 & ~n59265;
  assign n59399 = n8217 & ~n10750;
  assign n59400 = ~n8217 & ~n23940;
  assign n59401 = ~n59399 & ~n59400;
  assign n59402 = ~i_hbusreq6 & ~n59401;
  assign n59403 = ~n42534 & ~n59402;
  assign n59404 = controllable_hgrant6 & ~n59403;
  assign n59405 = i_hbusreq6 & ~n59231;
  assign n59406 = controllable_hmaster2 & ~n59386;
  assign n59407 = i_hbusreq5 & ~n59205;
  assign n59408 = i_hbusreq4 & ~n59203;
  assign n59409 = i_hbusreq9 & ~n59203;
  assign n59410 = i_hbusreq3 & ~n59201;
  assign n59411 = n8365 & ~n15682;
  assign n59412 = ~n8365 & ~n23897;
  assign n59413 = ~n59411 & ~n59412;
  assign n59414 = ~i_hbusreq3 & ~n59413;
  assign n59415 = ~n59410 & ~n59414;
  assign n59416 = controllable_hgrant3 & ~n59415;
  assign n59417 = ~n59375 & ~n59416;
  assign n59418 = ~i_hbusreq9 & ~n59417;
  assign n59419 = ~n59409 & ~n59418;
  assign n59420 = ~i_hbusreq4 & ~n59419;
  assign n59421 = ~n59408 & ~n59420;
  assign n59422 = ~controllable_hgrant4 & ~n59421;
  assign n59423 = ~n59350 & ~n59422;
  assign n59424 = ~i_hbusreq5 & ~n59423;
  assign n59425 = ~n59407 & ~n59424;
  assign n59426 = ~controllable_hgrant5 & ~n59425;
  assign n59427 = ~n59341 & ~n59426;
  assign n59428 = ~controllable_hmaster2 & ~n59427;
  assign n59429 = ~n59406 & ~n59428;
  assign n59430 = controllable_hmaster1 & ~n59429;
  assign n59431 = i_hbusreq5 & ~n59213;
  assign n59432 = n8378 & ~n15692;
  assign n59433 = ~n8378 & ~n23907;
  assign n59434 = ~n59432 & ~n59433;
  assign n59435 = ~i_hbusreq5 & ~n59434;
  assign n59436 = ~n59431 & ~n59435;
  assign n59437 = controllable_hgrant5 & ~n59436;
  assign n59438 = ~n59385 & ~n59437;
  assign n59439 = controllable_hmaster2 & ~n59438;
  assign n59440 = i_hbusreq5 & ~n59225;
  assign n59441 = i_hbusreq4 & ~n59223;
  assign n59442 = i_hbusreq9 & ~n59223;
  assign n59443 = i_hbusreq3 & ~n59221;
  assign n59444 = i_hbusreq1 & ~n59219;
  assign n59445 = n8389 & ~n15678;
  assign n59446 = ~n8389 & ~n23893;
  assign n59447 = ~n59445 & ~n59446;
  assign n59448 = ~i_hbusreq1 & ~n59447;
  assign n59449 = ~n59444 & ~n59448;
  assign n59450 = controllable_hgrant1 & ~n59449;
  assign n59451 = ~n59371 & ~n59450;
  assign n59452 = ~i_hbusreq3 & ~n59451;
  assign n59453 = ~n59443 & ~n59452;
  assign n59454 = ~controllable_hgrant3 & ~n59453;
  assign n59455 = ~n59358 & ~n59454;
  assign n59456 = ~i_hbusreq9 & ~n59455;
  assign n59457 = ~n59442 & ~n59456;
  assign n59458 = ~i_hbusreq4 & ~n59457;
  assign n59459 = ~n59441 & ~n59458;
  assign n59460 = ~controllable_hgrant4 & ~n59459;
  assign n59461 = ~n59350 & ~n59460;
  assign n59462 = ~i_hbusreq5 & ~n59461;
  assign n59463 = ~n59440 & ~n59462;
  assign n59464 = ~controllable_hgrant5 & ~n59463;
  assign n59465 = ~n59341 & ~n59464;
  assign n59466 = ~controllable_hmaster2 & ~n59465;
  assign n59467 = ~n59439 & ~n59466;
  assign n59468 = ~controllable_hmaster1 & ~n59467;
  assign n59469 = ~n59430 & ~n59468;
  assign n59470 = ~i_hbusreq6 & ~n59469;
  assign n59471 = ~n59405 & ~n59470;
  assign n59472 = ~controllable_hgrant6 & ~n59471;
  assign n59473 = ~n59404 & ~n59472;
  assign n59474 = controllable_hmaster0 & ~n59473;
  assign n59475 = i_hbusreq6 & ~n59237;
  assign n59476 = ~n10778 & ~n28100;
  assign n59477 = n8217 & ~n59476;
  assign n59478 = ~n23982 & ~n33482;
  assign n59479 = ~n8217 & ~n59478;
  assign n59480 = ~n59477 & ~n59479;
  assign n59481 = ~i_hbusreq6 & ~n59480;
  assign n59482 = ~n59475 & ~n59481;
  assign n59483 = controllable_hgrant6 & ~n59482;
  assign n59484 = i_hbusreq6 & ~n59261;
  assign n59485 = i_hbusreq5 & ~n59245;
  assign n59486 = i_hbusreq4 & ~n59243;
  assign n59487 = i_hbusreq9 & ~n59243;
  assign n59488 = i_hbusreq3 & ~n59241;
  assign n59489 = i_hbusreq1 & ~n59239;
  assign n59490 = n7928 & ~n48586;
  assign n59491 = ~i_hbusreq1 & ~n59490;
  assign n59492 = ~n59489 & ~n59491;
  assign n59493 = ~controllable_hgrant1 & ~n59492;
  assign n59494 = ~n59366 & ~n59493;
  assign n59495 = ~i_hbusreq3 & ~n59494;
  assign n59496 = ~n59488 & ~n59495;
  assign n59497 = ~controllable_hgrant3 & ~n59496;
  assign n59498 = ~n59358 & ~n59497;
  assign n59499 = ~i_hbusreq9 & ~n59498;
  assign n59500 = ~n59487 & ~n59499;
  assign n59501 = ~i_hbusreq4 & ~n59500;
  assign n59502 = ~n59486 & ~n59501;
  assign n59503 = ~controllable_hgrant4 & ~n59502;
  assign n59504 = ~n59350 & ~n59503;
  assign n59505 = ~i_hbusreq5 & ~n59504;
  assign n59506 = ~n59485 & ~n59505;
  assign n59507 = ~controllable_hgrant5 & ~n59506;
  assign n59508 = ~n59341 & ~n59507;
  assign n59509 = ~controllable_hmaster2 & ~n59508;
  assign n59510 = ~n59406 & ~n59509;
  assign n59511 = controllable_hmaster1 & ~n59510;
  assign n59512 = i_hbusreq5 & ~n59255;
  assign n59513 = i_hbusreq4 & ~n59253;
  assign n59514 = i_hbusreq9 & ~n59253;
  assign n59515 = n8426 & ~n15686;
  assign n59516 = ~n8426 & ~n23901;
  assign n59517 = ~n59515 & ~n59516;
  assign n59518 = ~i_hbusreq9 & ~n59517;
  assign n59519 = ~n59514 & ~n59518;
  assign n59520 = ~i_hbusreq4 & ~n59519;
  assign n59521 = ~n59513 & ~n59520;
  assign n59522 = controllable_hgrant4 & ~n59521;
  assign n59523 = ~n59381 & ~n59522;
  assign n59524 = ~i_hbusreq5 & ~n59523;
  assign n59525 = ~n59512 & ~n59524;
  assign n59526 = ~controllable_hgrant5 & ~n59525;
  assign n59527 = ~n59341 & ~n59526;
  assign n59528 = controllable_hmaster2 & ~n59527;
  assign n59529 = n8378 & ~n10773;
  assign n59530 = ~n8378 & ~n23975;
  assign n59531 = ~n59529 & ~n59530;
  assign n59532 = ~i_hbusreq5 & ~n59531;
  assign n59533 = ~n51713 & ~n59532;
  assign n59534 = controllable_hgrant5 & ~n59533;
  assign n59535 = n8426 & ~n10769;
  assign n59536 = ~n8426 & ~n23969;
  assign n59537 = ~n59535 & ~n59536;
  assign n59538 = ~i_hbusreq9 & ~n59537;
  assign n59539 = ~n52016 & ~n59538;
  assign n59540 = ~i_hbusreq4 & ~n59539;
  assign n59541 = ~n52015 & ~n59540;
  assign n59542 = controllable_hgrant4 & ~n59541;
  assign n59543 = n8365 & ~n10767;
  assign n59544 = ~n8365 & ~n23965;
  assign n59545 = ~n59543 & ~n59544;
  assign n59546 = ~i_hbusreq3 & ~n59545;
  assign n59547 = ~n52423 & ~n59546;
  assign n59548 = controllable_hgrant3 & ~n59547;
  assign n59549 = n8389 & ~n10765;
  assign n59550 = ~n8389 & ~n23961;
  assign n59551 = ~n59549 & ~n59550;
  assign n59552 = ~i_hbusreq1 & ~n59551;
  assign n59553 = ~n59360 & ~n59552;
  assign n59554 = controllable_hgrant1 & ~n59553;
  assign n59555 = n7928 & ~n48695;
  assign n59556 = ~i_hbusreq1 & ~n59555;
  assign n59557 = ~n59367 & ~n59556;
  assign n59558 = ~controllable_hgrant1 & ~n59557;
  assign n59559 = ~n59554 & ~n59558;
  assign n59560 = ~i_hbusreq3 & ~n59559;
  assign n59561 = ~n59359 & ~n59560;
  assign n59562 = ~controllable_hgrant3 & ~n59561;
  assign n59563 = ~n59548 & ~n59562;
  assign n59564 = ~i_hbusreq9 & ~n59563;
  assign n59565 = ~n59352 & ~n59564;
  assign n59566 = ~i_hbusreq4 & ~n59565;
  assign n59567 = ~n59351 & ~n59566;
  assign n59568 = ~controllable_hgrant4 & ~n59567;
  assign n59569 = ~n59542 & ~n59568;
  assign n59570 = ~i_hbusreq5 & ~n59569;
  assign n59571 = ~n59342 & ~n59570;
  assign n59572 = ~controllable_hgrant5 & ~n59571;
  assign n59573 = ~n59534 & ~n59572;
  assign n59574 = ~controllable_hmaster2 & ~n59573;
  assign n59575 = ~n59528 & ~n59574;
  assign n59576 = ~controllable_hmaster1 & ~n59575;
  assign n59577 = ~n59511 & ~n59576;
  assign n59578 = ~i_hbusreq6 & ~n59577;
  assign n59579 = ~n59484 & ~n59578;
  assign n59580 = ~controllable_hgrant6 & ~n59579;
  assign n59581 = ~n59483 & ~n59580;
  assign n59582 = ~controllable_hmaster0 & ~n59581;
  assign n59583 = ~n59474 & ~n59582;
  assign n59584 = ~i_hbusreq8 & ~n59583;
  assign n59585 = ~n59398 & ~n59584;
  assign n59586 = ~controllable_hmaster3 & ~n59585;
  assign n59587 = ~n59397 & ~n59586;
  assign n59588 = ~i_hbusreq7 & ~n59587;
  assign n59589 = ~n59268 & ~n59588;
  assign n59590 = ~n7924 & ~n59589;
  assign n59591 = ~n8217 & ~n33506;
  assign n59592 = ~n42590 & ~n59591;
  assign n59593 = i_hlock6 & ~n59592;
  assign n59594 = ~n8217 & ~n33533;
  assign n59595 = ~n42590 & ~n59594;
  assign n59596 = ~i_hlock6 & ~n59595;
  assign n59597 = ~n59593 & ~n59596;
  assign n59598 = controllable_hgrant6 & ~n59597;
  assign n59599 = ~n8378 & ~n33499;
  assign n59600 = ~n51782 & ~n59599;
  assign n59601 = i_hlock5 & ~n59600;
  assign n59602 = ~n8378 & ~n33526;
  assign n59603 = ~n51782 & ~n59602;
  assign n59604 = ~i_hlock5 & ~n59603;
  assign n59605 = ~n59601 & ~n59604;
  assign n59606 = controllable_hgrant5 & ~n59605;
  assign n59607 = ~n8426 & ~n24001;
  assign n59608 = ~n52110 & ~n59607;
  assign n59609 = i_hlock4 & ~n59608;
  assign n59610 = ~n8426 & ~n24007;
  assign n59611 = ~n52110 & ~n59610;
  assign n59612 = ~i_hlock4 & ~n59611;
  assign n59613 = ~n59609 & ~n59612;
  assign n59614 = controllable_hgrant4 & ~n59613;
  assign n59615 = ~n8365 & ~n23999;
  assign n59616 = ~n52537 & ~n59615;
  assign n59617 = i_hlock3 & ~n59616;
  assign n59618 = ~n8365 & ~n24005;
  assign n59619 = ~n52537 & ~n59618;
  assign n59620 = ~i_hlock3 & ~n59619;
  assign n59621 = ~n59617 & ~n59620;
  assign n59622 = controllable_hgrant3 & ~n59621;
  assign n59623 = n8389 & ~n13180;
  assign n59624 = ~n8389 & ~n23997;
  assign n59625 = ~n59623 & ~n59624;
  assign n59626 = i_hlock1 & ~n59625;
  assign n59627 = ~n8389 & ~n24003;
  assign n59628 = ~n59623 & ~n59627;
  assign n59629 = ~i_hlock1 & ~n59628;
  assign n59630 = ~n59626 & ~n59629;
  assign n59631 = controllable_hgrant1 & ~n59630;
  assign n59632 = n7928 & ~n48800;
  assign n59633 = ~controllable_hgrant1 & ~n59632;
  assign n59634 = ~n59631 & ~n59633;
  assign n59635 = ~controllable_hgrant3 & ~n59634;
  assign n59636 = ~n59622 & ~n59635;
  assign n59637 = ~controllable_hgrant4 & ~n59636;
  assign n59638 = ~n59614 & ~n59637;
  assign n59639 = ~controllable_hgrant5 & ~n59638;
  assign n59640 = ~n59606 & ~n59639;
  assign n59641 = controllable_hmaster1 & ~n59640;
  assign n59642 = controllable_hmaster2 & ~n59640;
  assign n59643 = ~n8389 & ~n17510;
  assign n59644 = ~n59623 & ~n59643;
  assign n59645 = i_hlock1 & ~n59644;
  assign n59646 = ~n8389 & ~n17518;
  assign n59647 = ~n59623 & ~n59646;
  assign n59648 = ~i_hlock1 & ~n59647;
  assign n59649 = ~n59645 & ~n59648;
  assign n59650 = controllable_hgrant1 & ~n59649;
  assign n59651 = n7928 & ~n46063;
  assign n59652 = ~controllable_hgrant1 & ~n59651;
  assign n59653 = ~n59650 & ~n59652;
  assign n59654 = ~controllable_hgrant3 & ~n59653;
  assign n59655 = ~n52545 & ~n59654;
  assign n59656 = ~controllable_hgrant4 & ~n59655;
  assign n59657 = ~n52118 & ~n59656;
  assign n59658 = ~controllable_hgrant5 & ~n59657;
  assign n59659 = ~n51790 & ~n59658;
  assign n59660 = ~controllable_hmaster2 & ~n59659;
  assign n59661 = ~n59642 & ~n59660;
  assign n59662 = ~controllable_hmaster1 & ~n59661;
  assign n59663 = ~n59641 & ~n59662;
  assign n59664 = ~controllable_hgrant6 & ~n59663;
  assign n59665 = ~n59598 & ~n59664;
  assign n59666 = controllable_hmaster3 & ~n59665;
  assign n59667 = controllable_hmaster2 & ~n59659;
  assign n59668 = n8365 & ~n13392;
  assign n59669 = ~n8365 & ~n24018;
  assign n59670 = ~n59668 & ~n59669;
  assign n59671 = i_hlock3 & ~n59670;
  assign n59672 = ~n8365 & ~n24024;
  assign n59673 = ~n59668 & ~n59672;
  assign n59674 = ~i_hlock3 & ~n59673;
  assign n59675 = ~n59671 & ~n59674;
  assign n59676 = controllable_hgrant3 & ~n59675;
  assign n59677 = ~n59654 & ~n59676;
  assign n59678 = ~controllable_hgrant4 & ~n59677;
  assign n59679 = ~n52118 & ~n59678;
  assign n59680 = ~controllable_hgrant5 & ~n59679;
  assign n59681 = ~n51790 & ~n59680;
  assign n59682 = ~controllable_hmaster2 & ~n59681;
  assign n59683 = ~n59667 & ~n59682;
  assign n59684 = controllable_hmaster1 & ~n59683;
  assign n59685 = n8378 & ~n13396;
  assign n59686 = ~n8378 & ~n33511;
  assign n59687 = ~n59685 & ~n59686;
  assign n59688 = i_hlock5 & ~n59687;
  assign n59689 = ~n8378 & ~n33538;
  assign n59690 = ~n59685 & ~n59689;
  assign n59691 = ~i_hlock5 & ~n59690;
  assign n59692 = ~n59688 & ~n59691;
  assign n59693 = controllable_hgrant5 & ~n59692;
  assign n59694 = ~n59658 & ~n59693;
  assign n59695 = controllable_hmaster2 & ~n59694;
  assign n59696 = n8389 & ~n13390;
  assign n59697 = ~n8389 & ~n24016;
  assign n59698 = ~n59696 & ~n59697;
  assign n59699 = i_hlock1 & ~n59698;
  assign n59700 = ~n8389 & ~n24022;
  assign n59701 = ~n59696 & ~n59700;
  assign n59702 = ~i_hlock1 & ~n59701;
  assign n59703 = ~n59699 & ~n59702;
  assign n59704 = controllable_hgrant1 & ~n59703;
  assign n59705 = ~n59652 & ~n59704;
  assign n59706 = ~controllable_hgrant3 & ~n59705;
  assign n59707 = ~n52545 & ~n59706;
  assign n59708 = ~controllable_hgrant4 & ~n59707;
  assign n59709 = ~n52118 & ~n59708;
  assign n59710 = ~controllable_hgrant5 & ~n59709;
  assign n59711 = ~n51790 & ~n59710;
  assign n59712 = ~controllable_hmaster2 & ~n59711;
  assign n59713 = ~n59695 & ~n59712;
  assign n59714 = ~controllable_hmaster1 & ~n59713;
  assign n59715 = ~n59684 & ~n59714;
  assign n59716 = ~controllable_hgrant6 & ~n59715;
  assign n59717 = ~n42598 & ~n59716;
  assign n59718 = controllable_hmaster0 & ~n59717;
  assign n59719 = n8217 & ~n26937;
  assign n59720 = ~n8217 & ~n33517;
  assign n59721 = ~n59719 & ~n59720;
  assign n59722 = i_hlock6 & ~n59721;
  assign n59723 = ~n8217 & ~n33544;
  assign n59724 = ~n59719 & ~n59723;
  assign n59725 = ~i_hlock6 & ~n59724;
  assign n59726 = ~n59722 & ~n59725;
  assign n59727 = controllable_hgrant6 & ~n59726;
  assign n59728 = n7928 & ~n48981;
  assign n59729 = ~controllable_hgrant1 & ~n59728;
  assign n59730 = ~n59650 & ~n59729;
  assign n59731 = ~controllable_hgrant3 & ~n59730;
  assign n59732 = ~n52545 & ~n59731;
  assign n59733 = ~controllable_hgrant4 & ~n59732;
  assign n59734 = ~n52118 & ~n59733;
  assign n59735 = ~controllable_hgrant5 & ~n59734;
  assign n59736 = ~n51790 & ~n59735;
  assign n59737 = ~controllable_hmaster2 & ~n59736;
  assign n59738 = ~n59667 & ~n59737;
  assign n59739 = controllable_hmaster1 & ~n59738;
  assign n59740 = n8426 & ~n13394;
  assign n59741 = ~n8426 & ~n24020;
  assign n59742 = ~n59740 & ~n59741;
  assign n59743 = i_hlock4 & ~n59742;
  assign n59744 = ~n8426 & ~n24026;
  assign n59745 = ~n59740 & ~n59744;
  assign n59746 = ~i_hlock4 & ~n59745;
  assign n59747 = ~n59743 & ~n59746;
  assign n59748 = controllable_hgrant4 & ~n59747;
  assign n59749 = ~n59656 & ~n59748;
  assign n59750 = ~controllable_hgrant5 & ~n59749;
  assign n59751 = ~n51790 & ~n59750;
  assign n59752 = controllable_hmaster2 & ~n59751;
  assign n59753 = ~n59660 & ~n59752;
  assign n59754 = ~controllable_hmaster1 & ~n59753;
  assign n59755 = ~n59739 & ~n59754;
  assign n59756 = ~controllable_hgrant6 & ~n59755;
  assign n59757 = ~n59727 & ~n59756;
  assign n59758 = ~controllable_hmaster0 & ~n59757;
  assign n59759 = ~n59718 & ~n59758;
  assign n59760 = ~controllable_hmaster3 & ~n59759;
  assign n59761 = ~n59666 & ~n59760;
  assign n59762 = i_hbusreq7 & ~n59761;
  assign n59763 = i_hbusreq8 & ~n59665;
  assign n59764 = i_hbusreq6 & ~n59597;
  assign n59765 = n8217 & ~n15802;
  assign n59766 = ~n8217 & ~n33584;
  assign n59767 = ~n59765 & ~n59766;
  assign n59768 = i_hlock6 & ~n59767;
  assign n59769 = ~n8217 & ~n33674;
  assign n59770 = ~n59765 & ~n59769;
  assign n59771 = ~i_hlock6 & ~n59770;
  assign n59772 = ~n59768 & ~n59771;
  assign n59773 = ~i_hbusreq6 & ~n59772;
  assign n59774 = ~n59764 & ~n59773;
  assign n59775 = controllable_hgrant6 & ~n59774;
  assign n59776 = i_hbusreq6 & ~n59663;
  assign n59777 = i_hbusreq5 & ~n59605;
  assign n59778 = n8378 & ~n15745;
  assign n59779 = ~n8378 & ~n33564;
  assign n59780 = ~n59778 & ~n59779;
  assign n59781 = i_hlock5 & ~n59780;
  assign n59782 = ~n8378 & ~n33654;
  assign n59783 = ~n59778 & ~n59782;
  assign n59784 = ~i_hlock5 & ~n59783;
  assign n59785 = ~n59781 & ~n59784;
  assign n59786 = ~i_hbusreq5 & ~n59785;
  assign n59787 = ~n59777 & ~n59786;
  assign n59788 = controllable_hgrant5 & ~n59787;
  assign n59789 = i_hbusreq5 & ~n59638;
  assign n59790 = i_hbusreq4 & ~n59613;
  assign n59791 = i_hbusreq9 & ~n59608;
  assign n59792 = n8426 & ~n15739;
  assign n59793 = ~n8426 & ~n24065;
  assign n59794 = ~n59792 & ~n59793;
  assign n59795 = ~i_hbusreq9 & ~n59794;
  assign n59796 = ~n59791 & ~n59795;
  assign n59797 = i_hlock4 & ~n59796;
  assign n59798 = i_hbusreq9 & ~n59611;
  assign n59799 = ~n8426 & ~n24077;
  assign n59800 = ~n59792 & ~n59799;
  assign n59801 = ~i_hbusreq9 & ~n59800;
  assign n59802 = ~n59798 & ~n59801;
  assign n59803 = ~i_hlock4 & ~n59802;
  assign n59804 = ~n59797 & ~n59803;
  assign n59805 = ~i_hbusreq4 & ~n59804;
  assign n59806 = ~n59790 & ~n59805;
  assign n59807 = controllable_hgrant4 & ~n59806;
  assign n59808 = i_hbusreq4 & ~n59636;
  assign n59809 = i_hbusreq9 & ~n59636;
  assign n59810 = i_hbusreq3 & ~n59621;
  assign n59811 = n8365 & ~n15735;
  assign n59812 = ~n8365 & ~n24061;
  assign n59813 = ~n59811 & ~n59812;
  assign n59814 = i_hlock3 & ~n59813;
  assign n59815 = ~n8365 & ~n24073;
  assign n59816 = ~n59811 & ~n59815;
  assign n59817 = ~i_hlock3 & ~n59816;
  assign n59818 = ~n59814 & ~n59817;
  assign n59819 = ~i_hbusreq3 & ~n59818;
  assign n59820 = ~n59810 & ~n59819;
  assign n59821 = controllable_hgrant3 & ~n59820;
  assign n59822 = i_hbusreq3 & ~n59634;
  assign n59823 = i_hbusreq1 & ~n59630;
  assign n59824 = n8389 & ~n15731;
  assign n59825 = ~n8389 & ~n24057;
  assign n59826 = ~n59824 & ~n59825;
  assign n59827 = i_hlock1 & ~n59826;
  assign n59828 = ~n8389 & ~n24069;
  assign n59829 = ~n59824 & ~n59828;
  assign n59830 = ~i_hlock1 & ~n59829;
  assign n59831 = ~n59827 & ~n59830;
  assign n59832 = ~i_hbusreq1 & ~n59831;
  assign n59833 = ~n59823 & ~n59832;
  assign n59834 = controllable_hgrant1 & ~n59833;
  assign n59835 = i_hbusreq1 & ~n59632;
  assign n59836 = n7928 & ~n49199;
  assign n59837 = ~i_hbusreq1 & ~n59836;
  assign n59838 = ~n59835 & ~n59837;
  assign n59839 = ~controllable_hgrant1 & ~n59838;
  assign n59840 = ~n59834 & ~n59839;
  assign n59841 = ~i_hbusreq3 & ~n59840;
  assign n59842 = ~n59822 & ~n59841;
  assign n59843 = ~controllable_hgrant3 & ~n59842;
  assign n59844 = ~n59821 & ~n59843;
  assign n59845 = ~i_hbusreq9 & ~n59844;
  assign n59846 = ~n59809 & ~n59845;
  assign n59847 = ~i_hbusreq4 & ~n59846;
  assign n59848 = ~n59808 & ~n59847;
  assign n59849 = ~controllable_hgrant4 & ~n59848;
  assign n59850 = ~n59807 & ~n59849;
  assign n59851 = ~i_hbusreq5 & ~n59850;
  assign n59852 = ~n59789 & ~n59851;
  assign n59853 = ~controllable_hgrant5 & ~n59852;
  assign n59854 = ~n59788 & ~n59853;
  assign n59855 = controllable_hmaster1 & ~n59854;
  assign n59856 = controllable_hmaster2 & ~n59854;
  assign n59857 = n8378 & ~n15794;
  assign n59858 = ~n8378 & ~n33576;
  assign n59859 = ~n59857 & ~n59858;
  assign n59860 = i_hlock5 & ~n59859;
  assign n59861 = ~n8378 & ~n33666;
  assign n59862 = ~n59857 & ~n59861;
  assign n59863 = ~i_hlock5 & ~n59862;
  assign n59864 = ~n59860 & ~n59863;
  assign n59865 = ~i_hbusreq5 & ~n59864;
  assign n59866 = ~n51854 & ~n59865;
  assign n59867 = controllable_hgrant5 & ~n59866;
  assign n59868 = i_hbusreq5 & ~n59657;
  assign n59869 = n8426 & ~n15788;
  assign n59870 = ~n8426 & ~n24148;
  assign n59871 = ~n59869 & ~n59870;
  assign n59872 = ~i_hbusreq9 & ~n59871;
  assign n59873 = ~n52208 & ~n59872;
  assign n59874 = i_hlock4 & ~n59873;
  assign n59875 = ~n8426 & ~n24158;
  assign n59876 = ~n59869 & ~n59875;
  assign n59877 = ~i_hbusreq9 & ~n59876;
  assign n59878 = ~n52215 & ~n59877;
  assign n59879 = ~i_hlock4 & ~n59878;
  assign n59880 = ~n59874 & ~n59879;
  assign n59881 = ~i_hbusreq4 & ~n59880;
  assign n59882 = ~n52207 & ~n59881;
  assign n59883 = controllable_hgrant4 & ~n59882;
  assign n59884 = i_hbusreq4 & ~n59655;
  assign n59885 = i_hbusreq9 & ~n59655;
  assign n59886 = n8365 & ~n15784;
  assign n59887 = ~n8365 & ~n24144;
  assign n59888 = ~n59886 & ~n59887;
  assign n59889 = i_hlock3 & ~n59888;
  assign n59890 = ~n8365 & ~n24154;
  assign n59891 = ~n59886 & ~n59890;
  assign n59892 = ~i_hlock3 & ~n59891;
  assign n59893 = ~n59889 & ~n59892;
  assign n59894 = ~i_hbusreq3 & ~n59893;
  assign n59895 = ~n52649 & ~n59894;
  assign n59896 = controllable_hgrant3 & ~n59895;
  assign n59897 = i_hbusreq3 & ~n59653;
  assign n59898 = i_hbusreq1 & ~n59649;
  assign n59899 = n8389 & ~n15780;
  assign n59900 = ~n8389 & ~n24140;
  assign n59901 = ~n59899 & ~n59900;
  assign n59902 = i_hlock1 & ~n59901;
  assign n59903 = ~n8389 & ~n24150;
  assign n59904 = ~n59899 & ~n59903;
  assign n59905 = ~i_hlock1 & ~n59904;
  assign n59906 = ~n59902 & ~n59905;
  assign n59907 = ~i_hbusreq1 & ~n59906;
  assign n59908 = ~n59898 & ~n59907;
  assign n59909 = controllable_hgrant1 & ~n59908;
  assign n59910 = i_hbusreq1 & ~n59651;
  assign n59911 = n7928 & ~n49300;
  assign n59912 = ~i_hbusreq1 & ~n59911;
  assign n59913 = ~n59910 & ~n59912;
  assign n59914 = ~controllable_hgrant1 & ~n59913;
  assign n59915 = ~n59909 & ~n59914;
  assign n59916 = ~i_hbusreq3 & ~n59915;
  assign n59917 = ~n59897 & ~n59916;
  assign n59918 = ~controllable_hgrant3 & ~n59917;
  assign n59919 = ~n59896 & ~n59918;
  assign n59920 = ~i_hbusreq9 & ~n59919;
  assign n59921 = ~n59885 & ~n59920;
  assign n59922 = ~i_hbusreq4 & ~n59921;
  assign n59923 = ~n59884 & ~n59922;
  assign n59924 = ~controllable_hgrant4 & ~n59923;
  assign n59925 = ~n59883 & ~n59924;
  assign n59926 = ~i_hbusreq5 & ~n59925;
  assign n59927 = ~n59868 & ~n59926;
  assign n59928 = ~controllable_hgrant5 & ~n59927;
  assign n59929 = ~n59867 & ~n59928;
  assign n59930 = ~controllable_hmaster2 & ~n59929;
  assign n59931 = ~n59856 & ~n59930;
  assign n59932 = ~controllable_hmaster1 & ~n59931;
  assign n59933 = ~n59855 & ~n59932;
  assign n59934 = ~i_hbusreq6 & ~n59933;
  assign n59935 = ~n59776 & ~n59934;
  assign n59936 = ~controllable_hgrant6 & ~n59935;
  assign n59937 = ~n59775 & ~n59936;
  assign n59938 = ~i_hbusreq8 & ~n59937;
  assign n59939 = ~n59763 & ~n59938;
  assign n59940 = controllable_hmaster3 & ~n59939;
  assign n59941 = i_hbusreq8 & ~n59759;
  assign n59942 = n8217 & ~n15798;
  assign n59943 = ~n8217 & ~n33580;
  assign n59944 = ~n59942 & ~n59943;
  assign n59945 = i_hlock6 & ~n59944;
  assign n59946 = ~n8217 & ~n33670;
  assign n59947 = ~n59942 & ~n59946;
  assign n59948 = ~i_hlock6 & ~n59947;
  assign n59949 = ~n59945 & ~n59948;
  assign n59950 = ~i_hbusreq6 & ~n59949;
  assign n59951 = ~n42645 & ~n59950;
  assign n59952 = controllable_hgrant6 & ~n59951;
  assign n59953 = i_hbusreq6 & ~n59715;
  assign n59954 = controllable_hmaster2 & ~n59929;
  assign n59955 = i_hbusreq5 & ~n59679;
  assign n59956 = i_hbusreq4 & ~n59677;
  assign n59957 = i_hbusreq9 & ~n59677;
  assign n59958 = i_hbusreq3 & ~n59675;
  assign n59959 = n8365 & ~n15756;
  assign n59960 = ~n8365 & ~n24101;
  assign n59961 = ~n59959 & ~n59960;
  assign n59962 = i_hlock3 & ~n59961;
  assign n59963 = ~n8365 & ~n24113;
  assign n59964 = ~n59959 & ~n59963;
  assign n59965 = ~i_hlock3 & ~n59964;
  assign n59966 = ~n59962 & ~n59965;
  assign n59967 = ~i_hbusreq3 & ~n59966;
  assign n59968 = ~n59958 & ~n59967;
  assign n59969 = controllable_hgrant3 & ~n59968;
  assign n59970 = ~n59918 & ~n59969;
  assign n59971 = ~i_hbusreq9 & ~n59970;
  assign n59972 = ~n59957 & ~n59971;
  assign n59973 = ~i_hbusreq4 & ~n59972;
  assign n59974 = ~n59956 & ~n59973;
  assign n59975 = ~controllable_hgrant4 & ~n59974;
  assign n59976 = ~n59883 & ~n59975;
  assign n59977 = ~i_hbusreq5 & ~n59976;
  assign n59978 = ~n59955 & ~n59977;
  assign n59979 = ~controllable_hgrant5 & ~n59978;
  assign n59980 = ~n59867 & ~n59979;
  assign n59981 = ~controllable_hmaster2 & ~n59980;
  assign n59982 = ~n59954 & ~n59981;
  assign n59983 = controllable_hmaster1 & ~n59982;
  assign n59984 = i_hbusreq5 & ~n59692;
  assign n59985 = n8378 & ~n15766;
  assign n59986 = ~n8378 & ~n33602;
  assign n59987 = ~n59985 & ~n59986;
  assign n59988 = i_hlock5 & ~n59987;
  assign n59989 = ~n8378 & ~n33692;
  assign n59990 = ~n59985 & ~n59989;
  assign n59991 = ~i_hlock5 & ~n59990;
  assign n59992 = ~n59988 & ~n59991;
  assign n59993 = ~i_hbusreq5 & ~n59992;
  assign n59994 = ~n59984 & ~n59993;
  assign n59995 = controllable_hgrant5 & ~n59994;
  assign n59996 = ~n59928 & ~n59995;
  assign n59997 = controllable_hmaster2 & ~n59996;
  assign n59998 = i_hbusreq5 & ~n59709;
  assign n59999 = i_hbusreq4 & ~n59707;
  assign n60000 = i_hbusreq9 & ~n59707;
  assign n60001 = i_hbusreq3 & ~n59705;
  assign n60002 = i_hbusreq1 & ~n59703;
  assign n60003 = n8389 & ~n15752;
  assign n60004 = ~n8389 & ~n24097;
  assign n60005 = ~n60003 & ~n60004;
  assign n60006 = i_hlock1 & ~n60005;
  assign n60007 = ~n8389 & ~n24109;
  assign n60008 = ~n60003 & ~n60007;
  assign n60009 = ~i_hlock1 & ~n60008;
  assign n60010 = ~n60006 & ~n60009;
  assign n60011 = ~i_hbusreq1 & ~n60010;
  assign n60012 = ~n60002 & ~n60011;
  assign n60013 = controllable_hgrant1 & ~n60012;
  assign n60014 = ~n59914 & ~n60013;
  assign n60015 = ~i_hbusreq3 & ~n60014;
  assign n60016 = ~n60001 & ~n60015;
  assign n60017 = ~controllable_hgrant3 & ~n60016;
  assign n60018 = ~n59896 & ~n60017;
  assign n60019 = ~i_hbusreq9 & ~n60018;
  assign n60020 = ~n60000 & ~n60019;
  assign n60021 = ~i_hbusreq4 & ~n60020;
  assign n60022 = ~n59999 & ~n60021;
  assign n60023 = ~controllable_hgrant4 & ~n60022;
  assign n60024 = ~n59883 & ~n60023;
  assign n60025 = ~i_hbusreq5 & ~n60024;
  assign n60026 = ~n59998 & ~n60025;
  assign n60027 = ~controllable_hgrant5 & ~n60026;
  assign n60028 = ~n59867 & ~n60027;
  assign n60029 = ~controllable_hmaster2 & ~n60028;
  assign n60030 = ~n59997 & ~n60029;
  assign n60031 = ~controllable_hmaster1 & ~n60030;
  assign n60032 = ~n59983 & ~n60031;
  assign n60033 = ~i_hbusreq6 & ~n60032;
  assign n60034 = ~n59953 & ~n60033;
  assign n60035 = ~controllable_hgrant6 & ~n60034;
  assign n60036 = ~n59952 & ~n60035;
  assign n60037 = controllable_hmaster0 & ~n60036;
  assign n60038 = i_hbusreq6 & ~n59726;
  assign n60039 = ~n15846 & ~n28124;
  assign n60040 = n8217 & ~n60039;
  assign n60041 = ~n33609 & ~n33631;
  assign n60042 = ~n8217 & ~n60041;
  assign n60043 = ~n60040 & ~n60042;
  assign n60044 = i_hlock6 & ~n60043;
  assign n60045 = ~n33699 & ~n33721;
  assign n60046 = ~n8217 & ~n60045;
  assign n60047 = ~n60040 & ~n60046;
  assign n60048 = ~i_hlock6 & ~n60047;
  assign n60049 = ~n60044 & ~n60048;
  assign n60050 = ~i_hbusreq6 & ~n60049;
  assign n60051 = ~n60038 & ~n60050;
  assign n60052 = controllable_hgrant6 & ~n60051;
  assign n60053 = i_hbusreq6 & ~n59755;
  assign n60054 = i_hbusreq5 & ~n59734;
  assign n60055 = i_hbusreq4 & ~n59732;
  assign n60056 = i_hbusreq9 & ~n59732;
  assign n60057 = i_hbusreq3 & ~n59730;
  assign n60058 = i_hbusreq1 & ~n59728;
  assign n60059 = n7928 & ~n49774;
  assign n60060 = ~i_hbusreq1 & ~n60059;
  assign n60061 = ~n60058 & ~n60060;
  assign n60062 = ~controllable_hgrant1 & ~n60061;
  assign n60063 = ~n59909 & ~n60062;
  assign n60064 = ~i_hbusreq3 & ~n60063;
  assign n60065 = ~n60057 & ~n60064;
  assign n60066 = ~controllable_hgrant3 & ~n60065;
  assign n60067 = ~n59896 & ~n60066;
  assign n60068 = ~i_hbusreq9 & ~n60067;
  assign n60069 = ~n60056 & ~n60068;
  assign n60070 = ~i_hbusreq4 & ~n60069;
  assign n60071 = ~n60055 & ~n60070;
  assign n60072 = ~controllable_hgrant4 & ~n60071;
  assign n60073 = ~n59883 & ~n60072;
  assign n60074 = ~i_hbusreq5 & ~n60073;
  assign n60075 = ~n60054 & ~n60074;
  assign n60076 = ~controllable_hgrant5 & ~n60075;
  assign n60077 = ~n59867 & ~n60076;
  assign n60078 = ~controllable_hmaster2 & ~n60077;
  assign n60079 = ~n59954 & ~n60078;
  assign n60080 = controllable_hmaster1 & ~n60079;
  assign n60081 = i_hbusreq5 & ~n59749;
  assign n60082 = i_hbusreq4 & ~n59747;
  assign n60083 = i_hbusreq9 & ~n59742;
  assign n60084 = n8426 & ~n15760;
  assign n60085 = ~n8426 & ~n24105;
  assign n60086 = ~n60084 & ~n60085;
  assign n60087 = ~i_hbusreq9 & ~n60086;
  assign n60088 = ~n60083 & ~n60087;
  assign n60089 = i_hlock4 & ~n60088;
  assign n60090 = i_hbusreq9 & ~n59745;
  assign n60091 = ~n8426 & ~n24117;
  assign n60092 = ~n60084 & ~n60091;
  assign n60093 = ~i_hbusreq9 & ~n60092;
  assign n60094 = ~n60090 & ~n60093;
  assign n60095 = ~i_hlock4 & ~n60094;
  assign n60096 = ~n60089 & ~n60095;
  assign n60097 = ~i_hbusreq4 & ~n60096;
  assign n60098 = ~n60082 & ~n60097;
  assign n60099 = controllable_hgrant4 & ~n60098;
  assign n60100 = ~n59924 & ~n60099;
  assign n60101 = ~i_hbusreq5 & ~n60100;
  assign n60102 = ~n60081 & ~n60101;
  assign n60103 = ~controllable_hgrant5 & ~n60102;
  assign n60104 = ~n59867 & ~n60103;
  assign n60105 = controllable_hmaster2 & ~n60104;
  assign n60106 = n8378 & ~n15839;
  assign n60107 = ~n8378 & ~n33624;
  assign n60108 = ~n60106 & ~n60107;
  assign n60109 = i_hlock5 & ~n60108;
  assign n60110 = ~n8378 & ~n33714;
  assign n60111 = ~n60106 & ~n60110;
  assign n60112 = ~i_hlock5 & ~n60111;
  assign n60113 = ~n60109 & ~n60112;
  assign n60114 = ~i_hbusreq5 & ~n60113;
  assign n60115 = ~n51854 & ~n60114;
  assign n60116 = controllable_hgrant5 & ~n60115;
  assign n60117 = n8426 & ~n15833;
  assign n60118 = ~n8426 & ~n24199;
  assign n60119 = ~n60117 & ~n60118;
  assign n60120 = ~i_hbusreq9 & ~n60119;
  assign n60121 = ~n52208 & ~n60120;
  assign n60122 = i_hlock4 & ~n60121;
  assign n60123 = ~n8426 & ~n24209;
  assign n60124 = ~n60117 & ~n60123;
  assign n60125 = ~i_hbusreq9 & ~n60124;
  assign n60126 = ~n52215 & ~n60125;
  assign n60127 = ~i_hlock4 & ~n60126;
  assign n60128 = ~n60122 & ~n60127;
  assign n60129 = ~i_hbusreq4 & ~n60128;
  assign n60130 = ~n52207 & ~n60129;
  assign n60131 = controllable_hgrant4 & ~n60130;
  assign n60132 = n8365 & ~n15829;
  assign n60133 = ~n8365 & ~n24195;
  assign n60134 = ~n60132 & ~n60133;
  assign n60135 = i_hlock3 & ~n60134;
  assign n60136 = ~n8365 & ~n24205;
  assign n60137 = ~n60132 & ~n60136;
  assign n60138 = ~i_hlock3 & ~n60137;
  assign n60139 = ~n60135 & ~n60138;
  assign n60140 = ~i_hbusreq3 & ~n60139;
  assign n60141 = ~n52649 & ~n60140;
  assign n60142 = controllable_hgrant3 & ~n60141;
  assign n60143 = n8389 & ~n15825;
  assign n60144 = ~n8389 & ~n24191;
  assign n60145 = ~n60143 & ~n60144;
  assign n60146 = i_hlock1 & ~n60145;
  assign n60147 = ~n8389 & ~n24201;
  assign n60148 = ~n60143 & ~n60147;
  assign n60149 = ~i_hlock1 & ~n60148;
  assign n60150 = ~n60146 & ~n60149;
  assign n60151 = ~i_hbusreq1 & ~n60150;
  assign n60152 = ~n59898 & ~n60151;
  assign n60153 = controllable_hgrant1 & ~n60152;
  assign n60154 = n7928 & ~n49927;
  assign n60155 = ~i_hbusreq1 & ~n60154;
  assign n60156 = ~n59910 & ~n60155;
  assign n60157 = ~controllable_hgrant1 & ~n60156;
  assign n60158 = ~n60153 & ~n60157;
  assign n60159 = ~i_hbusreq3 & ~n60158;
  assign n60160 = ~n59897 & ~n60159;
  assign n60161 = ~controllable_hgrant3 & ~n60160;
  assign n60162 = ~n60142 & ~n60161;
  assign n60163 = ~i_hbusreq9 & ~n60162;
  assign n60164 = ~n59885 & ~n60163;
  assign n60165 = ~i_hbusreq4 & ~n60164;
  assign n60166 = ~n59884 & ~n60165;
  assign n60167 = ~controllable_hgrant4 & ~n60166;
  assign n60168 = ~n60131 & ~n60167;
  assign n60169 = ~i_hbusreq5 & ~n60168;
  assign n60170 = ~n59868 & ~n60169;
  assign n60171 = ~controllable_hgrant5 & ~n60170;
  assign n60172 = ~n60116 & ~n60171;
  assign n60173 = ~controllable_hmaster2 & ~n60172;
  assign n60174 = ~n60105 & ~n60173;
  assign n60175 = ~controllable_hmaster1 & ~n60174;
  assign n60176 = ~n60080 & ~n60175;
  assign n60177 = ~i_hbusreq6 & ~n60176;
  assign n60178 = ~n60053 & ~n60177;
  assign n60179 = ~controllable_hgrant6 & ~n60178;
  assign n60180 = ~n60052 & ~n60179;
  assign n60181 = ~controllable_hmaster0 & ~n60180;
  assign n60182 = ~n60037 & ~n60181;
  assign n60183 = ~i_hbusreq8 & ~n60182;
  assign n60184 = ~n59941 & ~n60183;
  assign n60185 = ~controllable_hmaster3 & ~n60184;
  assign n60186 = ~n59940 & ~n60185;
  assign n60187 = ~i_hbusreq7 & ~n60186;
  assign n60188 = ~n59762 & ~n60187;
  assign n60189 = n7924 & ~n60188;
  assign n60190 = ~n59590 & ~n60189;
  assign n60191 = n8214 & ~n60190;
  assign n60192 = ~n59150 & ~n60191;
  assign n60193 = n8202 & ~n60192;
  assign n60194 = ~n59148 & ~n60193;
  assign n60195 = n7920 & ~n60194;
  assign n60196 = ~n58945 & ~n60195;
  assign n60197 = n7728 & ~n60196;
  assign n60198 = ~n7920 & ~n58927;
  assign n60199 = ~n7737 & n8389;
  assign n60200 = ~n8389 & ~n17001;
  assign n60201 = ~n60199 & ~n60200;
  assign n60202 = controllable_hgrant1 & ~n60201;
  assign n60203 = ~n7942 & ~n60202;
  assign n60204 = ~controllable_hgrant3 & ~n60203;
  assign n60205 = ~n7812 & ~n60204;
  assign n60206 = ~controllable_hgrant4 & ~n60205;
  assign n60207 = ~n7811 & ~n60206;
  assign n60208 = ~controllable_hgrant5 & ~n60207;
  assign n60209 = ~n7810 & ~n60208;
  assign n60210 = controllable_hmaster1 & ~n60209;
  assign n60211 = controllable_hmaster2 & ~n60209;
  assign n60212 = controllable_hmaster2 & ~n60211;
  assign n60213 = ~controllable_hmaster1 & ~n60212;
  assign n60214 = ~n60210 & ~n60213;
  assign n60215 = ~controllable_hgrant6 & ~n60214;
  assign n60216 = ~n7809 & ~n60215;
  assign n60217 = controllable_hmaster3 & ~n60216;
  assign n60218 = ~n58957 & ~n60217;
  assign n60219 = i_hbusreq7 & ~n60218;
  assign n60220 = i_hbusreq8 & ~n60216;
  assign n60221 = i_hbusreq6 & ~n60214;
  assign n60222 = i_hbusreq5 & ~n60207;
  assign n60223 = i_hbusreq4 & ~n60205;
  assign n60224 = i_hbusreq9 & ~n60205;
  assign n60225 = i_hbusreq3 & ~n60203;
  assign n60226 = i_hbusreq1 & ~n60201;
  assign n60227 = ~n7759 & n8389;
  assign n60228 = ~n8389 & ~n17042;
  assign n60229 = ~n60227 & ~n60228;
  assign n60230 = ~i_hbusreq1 & ~n60229;
  assign n60231 = ~n60226 & ~n60230;
  assign n60232 = controllable_hgrant1 & ~n60231;
  assign n60233 = ~n7991 & ~n60232;
  assign n60234 = ~i_hbusreq3 & ~n60233;
  assign n60235 = ~n60225 & ~n60234;
  assign n60236 = ~controllable_hgrant3 & ~n60235;
  assign n60237 = ~n7851 & ~n60236;
  assign n60238 = ~i_hbusreq9 & ~n60237;
  assign n60239 = ~n60224 & ~n60238;
  assign n60240 = ~i_hbusreq4 & ~n60239;
  assign n60241 = ~n60223 & ~n60240;
  assign n60242 = ~controllable_hgrant4 & ~n60241;
  assign n60243 = ~n7848 & ~n60242;
  assign n60244 = ~i_hbusreq5 & ~n60243;
  assign n60245 = ~n60222 & ~n60244;
  assign n60246 = ~controllable_hgrant5 & ~n60245;
  assign n60247 = ~n7846 & ~n60246;
  assign n60248 = controllable_hmaster1 & ~n60247;
  assign n60249 = controllable_hmaster2 & ~n60247;
  assign n60250 = controllable_hmaster2 & ~n60249;
  assign n60251 = ~controllable_hmaster1 & ~n60250;
  assign n60252 = ~n60248 & ~n60251;
  assign n60253 = ~i_hbusreq6 & ~n60252;
  assign n60254 = ~n60221 & ~n60253;
  assign n60255 = ~controllable_hgrant6 & ~n60254;
  assign n60256 = ~n7844 & ~n60255;
  assign n60257 = ~i_hbusreq8 & ~n60256;
  assign n60258 = ~n60220 & ~n60257;
  assign n60259 = controllable_hmaster3 & ~n60258;
  assign n60260 = ~n58980 & ~n60259;
  assign n60261 = ~i_hbusreq7 & ~n60260;
  assign n60262 = ~n60219 & ~n60261;
  assign n60263 = ~n7924 & ~n60262;
  assign n60264 = n8389 & ~n13015;
  assign n60265 = ~n8389 & ~n17095;
  assign n60266 = ~n60264 & ~n60265;
  assign n60267 = i_hlock1 & ~n60266;
  assign n60268 = ~n8389 & ~n17103;
  assign n60269 = ~n60264 & ~n60268;
  assign n60270 = ~i_hlock1 & ~n60269;
  assign n60271 = ~n60267 & ~n60270;
  assign n60272 = controllable_hgrant1 & ~n60271;
  assign n60273 = ~n8027 & ~n60272;
  assign n60274 = ~controllable_hgrant3 & ~n60273;
  assign n60275 = ~n7812 & ~n60274;
  assign n60276 = ~controllable_hgrant4 & ~n60275;
  assign n60277 = ~n7811 & ~n60276;
  assign n60278 = ~controllable_hgrant5 & ~n60277;
  assign n60279 = ~n7810 & ~n60278;
  assign n60280 = controllable_hmaster1 & ~n60279;
  assign n60281 = controllable_hmaster2 & ~n60279;
  assign n60282 = ~n8043 & ~n58993;
  assign n60283 = ~controllable_hgrant3 & ~n60282;
  assign n60284 = ~controllable_hgrant3 & ~n60283;
  assign n60285 = ~controllable_hgrant4 & ~n60284;
  assign n60286 = ~controllable_hgrant4 & ~n60285;
  assign n60287 = ~controllable_hgrant5 & ~n60286;
  assign n60288 = ~controllable_hgrant5 & ~n60287;
  assign n60289 = ~controllable_hmaster2 & ~n60288;
  assign n60290 = ~n60281 & ~n60289;
  assign n60291 = ~controllable_hmaster1 & ~n60290;
  assign n60292 = ~n60280 & ~n60291;
  assign n60293 = ~controllable_hgrant6 & ~n60292;
  assign n60294 = ~n7809 & ~n60293;
  assign n60295 = controllable_hmaster3 & ~n60294;
  assign n60296 = controllable_hmaster1 & ~n60288;
  assign n60297 = controllable_hmaster2 & ~n60288;
  assign n60298 = i_hlock1 & ~n40833;
  assign n60299 = ~i_hlock1 & ~n40839;
  assign n60300 = ~n60298 & ~n60299;
  assign n60301 = ~controllable_hgrant1 & ~n60300;
  assign n60302 = ~n48917 & ~n60301;
  assign n60303 = ~controllable_hgrant3 & ~n60302;
  assign n60304 = ~n48106 & ~n60303;
  assign n60305 = ~controllable_hgrant4 & ~n60304;
  assign n60306 = ~n48103 & ~n60305;
  assign n60307 = ~controllable_hgrant5 & ~n60306;
  assign n60308 = ~n48100 & ~n60307;
  assign n60309 = ~controllable_hmaster2 & ~n60308;
  assign n60310 = ~n60297 & ~n60309;
  assign n60311 = ~controllable_hmaster1 & ~n60310;
  assign n60312 = ~n60296 & ~n60311;
  assign n60313 = ~controllable_hgrant6 & ~n60312;
  assign n60314 = ~n58949 & ~n60313;
  assign n60315 = controllable_hmaster0 & ~n60314;
  assign n60316 = ~controllable_hgrant6 & ~n60288;
  assign n60317 = ~controllable_hgrant6 & ~n60316;
  assign n60318 = ~controllable_hmaster0 & ~n60317;
  assign n60319 = ~n60315 & ~n60318;
  assign n60320 = ~controllable_hmaster3 & ~n60319;
  assign n60321 = ~n60295 & ~n60320;
  assign n60322 = i_hbusreq7 & ~n60321;
  assign n60323 = i_hbusreq8 & ~n60294;
  assign n60324 = i_hbusreq6 & ~n60292;
  assign n60325 = i_hbusreq5 & ~n60277;
  assign n60326 = i_hbusreq4 & ~n60275;
  assign n60327 = i_hbusreq9 & ~n60275;
  assign n60328 = i_hbusreq3 & ~n60273;
  assign n60329 = i_hbusreq1 & ~n60271;
  assign n60330 = n8389 & ~n13061;
  assign n60331 = ~n8389 & ~n17160;
  assign n60332 = ~n60330 & ~n60331;
  assign n60333 = i_hlock1 & ~n60332;
  assign n60334 = ~n8389 & ~n17174;
  assign n60335 = ~n60330 & ~n60334;
  assign n60336 = ~i_hlock1 & ~n60335;
  assign n60337 = ~n60333 & ~n60336;
  assign n60338 = ~i_hbusreq1 & ~n60337;
  assign n60339 = ~n60329 & ~n60338;
  assign n60340 = controllable_hgrant1 & ~n60339;
  assign n60341 = ~n8082 & ~n60340;
  assign n60342 = ~i_hbusreq3 & ~n60341;
  assign n60343 = ~n60328 & ~n60342;
  assign n60344 = ~controllable_hgrant3 & ~n60343;
  assign n60345 = ~n7851 & ~n60344;
  assign n60346 = ~i_hbusreq9 & ~n60345;
  assign n60347 = ~n60327 & ~n60346;
  assign n60348 = ~i_hbusreq4 & ~n60347;
  assign n60349 = ~n60326 & ~n60348;
  assign n60350 = ~controllable_hgrant4 & ~n60349;
  assign n60351 = ~n7848 & ~n60350;
  assign n60352 = ~i_hbusreq5 & ~n60351;
  assign n60353 = ~n60325 & ~n60352;
  assign n60354 = ~controllable_hgrant5 & ~n60353;
  assign n60355 = ~n7846 & ~n60354;
  assign n60356 = controllable_hmaster1 & ~n60355;
  assign n60357 = controllable_hmaster2 & ~n60355;
  assign n60358 = i_hbusreq5 & ~n60286;
  assign n60359 = i_hbusreq4 & ~n60284;
  assign n60360 = i_hbusreq9 & ~n60284;
  assign n60361 = i_hbusreq3 & ~n60282;
  assign n60362 = ~n8119 & ~n59042;
  assign n60363 = ~i_hbusreq3 & ~n60362;
  assign n60364 = ~n60361 & ~n60363;
  assign n60365 = ~controllable_hgrant3 & ~n60364;
  assign n60366 = ~controllable_hgrant3 & ~n60365;
  assign n60367 = ~i_hbusreq9 & ~n60366;
  assign n60368 = ~n60360 & ~n60367;
  assign n60369 = ~i_hbusreq4 & ~n60368;
  assign n60370 = ~n60359 & ~n60369;
  assign n60371 = ~controllable_hgrant4 & ~n60370;
  assign n60372 = ~controllable_hgrant4 & ~n60371;
  assign n60373 = ~i_hbusreq5 & ~n60372;
  assign n60374 = ~n60358 & ~n60373;
  assign n60375 = ~controllable_hgrant5 & ~n60374;
  assign n60376 = ~controllable_hgrant5 & ~n60375;
  assign n60377 = ~controllable_hmaster2 & ~n60376;
  assign n60378 = ~n60357 & ~n60377;
  assign n60379 = ~controllable_hmaster1 & ~n60378;
  assign n60380 = ~n60356 & ~n60379;
  assign n60381 = ~i_hbusreq6 & ~n60380;
  assign n60382 = ~n60324 & ~n60381;
  assign n60383 = ~controllable_hgrant6 & ~n60382;
  assign n60384 = ~n7844 & ~n60383;
  assign n60385 = ~i_hbusreq8 & ~n60384;
  assign n60386 = ~n60323 & ~n60385;
  assign n60387 = controllable_hmaster3 & ~n60386;
  assign n60388 = i_hbusreq8 & ~n60319;
  assign n60389 = i_hbusreq6 & ~n60312;
  assign n60390 = controllable_hmaster1 & ~n60376;
  assign n60391 = controllable_hmaster2 & ~n60376;
  assign n60392 = i_hbusreq5 & ~n60306;
  assign n60393 = i_hbusreq4 & ~n60304;
  assign n60394 = i_hbusreq9 & ~n60304;
  assign n60395 = i_hbusreq3 & ~n60302;
  assign n60396 = i_hbusreq1 & ~n60300;
  assign n60397 = i_hlock1 & ~n40881;
  assign n60398 = ~i_hlock1 & ~n40893;
  assign n60399 = ~n60397 & ~n60398;
  assign n60400 = ~i_hbusreq1 & ~n60399;
  assign n60401 = ~n60396 & ~n60400;
  assign n60402 = ~controllable_hgrant1 & ~n60401;
  assign n60403 = ~n49636 & ~n60402;
  assign n60404 = ~i_hbusreq3 & ~n60403;
  assign n60405 = ~n60395 & ~n60404;
  assign n60406 = ~controllable_hgrant3 & ~n60405;
  assign n60407 = ~n48459 & ~n60406;
  assign n60408 = ~i_hbusreq9 & ~n60407;
  assign n60409 = ~n60394 & ~n60408;
  assign n60410 = ~i_hbusreq4 & ~n60409;
  assign n60411 = ~n60393 & ~n60410;
  assign n60412 = ~controllable_hgrant4 & ~n60411;
  assign n60413 = ~n48450 & ~n60412;
  assign n60414 = ~i_hbusreq5 & ~n60413;
  assign n60415 = ~n60392 & ~n60414;
  assign n60416 = ~controllable_hgrant5 & ~n60415;
  assign n60417 = ~n48439 & ~n60416;
  assign n60418 = ~controllable_hmaster2 & ~n60417;
  assign n60419 = ~n60391 & ~n60418;
  assign n60420 = ~controllable_hmaster1 & ~n60419;
  assign n60421 = ~n60390 & ~n60420;
  assign n60422 = ~i_hbusreq6 & ~n60421;
  assign n60423 = ~n60389 & ~n60422;
  assign n60424 = ~controllable_hgrant6 & ~n60423;
  assign n60425 = ~n58967 & ~n60424;
  assign n60426 = controllable_hmaster0 & ~n60425;
  assign n60427 = i_hbusreq6 & ~n60288;
  assign n60428 = ~i_hbusreq6 & ~n60376;
  assign n60429 = ~n60427 & ~n60428;
  assign n60430 = ~controllable_hgrant6 & ~n60429;
  assign n60431 = ~controllable_hgrant6 & ~n60430;
  assign n60432 = ~controllable_hmaster0 & ~n60431;
  assign n60433 = ~n60426 & ~n60432;
  assign n60434 = ~i_hbusreq8 & ~n60433;
  assign n60435 = ~n60388 & ~n60434;
  assign n60436 = ~controllable_hmaster3 & ~n60435;
  assign n60437 = ~n60387 & ~n60436;
  assign n60438 = ~i_hbusreq7 & ~n60437;
  assign n60439 = ~n60322 & ~n60438;
  assign n60440 = n7924 & ~n60439;
  assign n60441 = ~n60263 & ~n60440;
  assign n60442 = ~n8214 & ~n60441;
  assign n60443 = ~n7957 & ~n59119;
  assign n60444 = i_hbusreq7 & ~n60443;
  assign n60445 = ~n7957 & ~n59142;
  assign n60446 = ~i_hbusreq7 & ~n60445;
  assign n60447 = ~n60444 & ~n60446;
  assign n60448 = ~n7924 & ~n60447;
  assign n60449 = controllable_hmaster0 & ~n8059;
  assign n60450 = controllable_hmaster1 & ~n8050;
  assign n60451 = controllable_hmaster2 & ~n8050;
  assign n60452 = ~n8440 & ~n40832;
  assign n60453 = ~controllable_hgrant1 & ~n60452;
  assign n60454 = ~n48197 & ~n60453;
  assign n60455 = ~controllable_hgrant3 & ~n60454;
  assign n60456 = ~n48194 & ~n60455;
  assign n60457 = ~controllable_hgrant4 & ~n60456;
  assign n60458 = ~n48191 & ~n60457;
  assign n60459 = ~controllable_hgrant5 & ~n60458;
  assign n60460 = ~n48188 & ~n60459;
  assign n60461 = ~controllable_hmaster2 & ~n60460;
  assign n60462 = ~n60451 & ~n60461;
  assign n60463 = ~controllable_hmaster1 & ~n60462;
  assign n60464 = ~n60450 & ~n60463;
  assign n60465 = ~controllable_hgrant6 & ~n60464;
  assign n60466 = ~n59111 & ~n60465;
  assign n60467 = ~controllable_hmaster0 & ~n60466;
  assign n60468 = ~n60449 & ~n60467;
  assign n60469 = ~controllable_hmaster3 & ~n60468;
  assign n60470 = ~n8057 & ~n60469;
  assign n60471 = i_hbusreq7 & ~n60470;
  assign n60472 = ~n7814 & ~n49177;
  assign n60473 = ~n7733 & ~n60472;
  assign n60474 = ~n7733 & ~n60473;
  assign n60475 = n7928 & ~n60474;
  assign n60476 = ~n7929 & ~n60475;
  assign n60477 = ~i_hbusreq1 & ~n60476;
  assign n60478 = ~n8069 & ~n60477;
  assign n60479 = ~controllable_hgrant1 & ~n60478;
  assign n60480 = ~n7813 & ~n60479;
  assign n60481 = ~i_hbusreq3 & ~n60480;
  assign n60482 = ~n8068 & ~n60481;
  assign n60483 = ~controllable_hgrant3 & ~n60482;
  assign n60484 = ~n7812 & ~n60483;
  assign n60485 = ~i_hbusreq9 & ~n60484;
  assign n60486 = ~n8067 & ~n60485;
  assign n60487 = ~i_hbusreq4 & ~n60486;
  assign n60488 = ~n8066 & ~n60487;
  assign n60489 = ~controllable_hgrant4 & ~n60488;
  assign n60490 = ~n7811 & ~n60489;
  assign n60491 = ~i_hbusreq5 & ~n60490;
  assign n60492 = ~n8065 & ~n60491;
  assign n60493 = ~controllable_hgrant5 & ~n60492;
  assign n60494 = ~n7810 & ~n60493;
  assign n60495 = controllable_hmaster1 & ~n60494;
  assign n60496 = controllable_hmaster2 & ~n60494;
  assign n60497 = ~n7733 & ~n16577;
  assign n60498 = ~n7733 & ~n60497;
  assign n60499 = n7928 & ~n60498;
  assign n60500 = n7928 & ~n60499;
  assign n60501 = ~i_hbusreq1 & ~n60500;
  assign n60502 = ~n8104 & ~n60501;
  assign n60503 = ~controllable_hgrant1 & ~n60502;
  assign n60504 = ~controllable_hgrant1 & ~n60503;
  assign n60505 = ~i_hbusreq3 & ~n60504;
  assign n60506 = ~n8103 & ~n60505;
  assign n60507 = ~controllable_hgrant3 & ~n60506;
  assign n60508 = ~controllable_hgrant3 & ~n60507;
  assign n60509 = ~i_hbusreq9 & ~n60508;
  assign n60510 = ~n8102 & ~n60509;
  assign n60511 = ~i_hbusreq4 & ~n60510;
  assign n60512 = ~n8101 & ~n60511;
  assign n60513 = ~controllable_hgrant4 & ~n60512;
  assign n60514 = ~controllable_hgrant4 & ~n60513;
  assign n60515 = ~i_hbusreq5 & ~n60514;
  assign n60516 = ~n8100 & ~n60515;
  assign n60517 = ~controllable_hgrant5 & ~n60516;
  assign n60518 = ~controllable_hgrant5 & ~n60517;
  assign n60519 = ~controllable_hmaster2 & ~n60518;
  assign n60520 = ~n60496 & ~n60519;
  assign n60521 = ~controllable_hmaster1 & ~n60520;
  assign n60522 = ~n60495 & ~n60521;
  assign n60523 = ~i_hbusreq6 & ~n60522;
  assign n60524 = ~n8064 & ~n60523;
  assign n60525 = ~controllable_hgrant6 & ~n60524;
  assign n60526 = ~n7809 & ~n60525;
  assign n60527 = ~i_hbusreq8 & ~n60526;
  assign n60528 = ~n8063 & ~n60527;
  assign n60529 = controllable_hmaster3 & ~n60528;
  assign n60530 = i_hbusreq8 & ~n60468;
  assign n60531 = ~i_hbusreq6 & ~n60518;
  assign n60532 = ~n8147 & ~n60531;
  assign n60533 = ~controllable_hgrant6 & ~n60532;
  assign n60534 = ~controllable_hgrant6 & ~n60533;
  assign n60535 = controllable_hmaster0 & ~n60534;
  assign n60536 = i_hbusreq6 & ~n60464;
  assign n60537 = controllable_hmaster1 & ~n60518;
  assign n60538 = controllable_hmaster2 & ~n60518;
  assign n60539 = i_hbusreq5 & ~n60458;
  assign n60540 = i_hbusreq4 & ~n60456;
  assign n60541 = i_hbusreq9 & ~n60456;
  assign n60542 = i_hbusreq3 & ~n60454;
  assign n60543 = i_hbusreq1 & ~n60452;
  assign n60544 = ~n43669 & ~n49909;
  assign n60545 = ~n7733 & ~n60544;
  assign n60546 = ~n40228 & ~n60545;
  assign n60547 = n7928 & ~n60546;
  assign n60548 = ~n8440 & ~n60547;
  assign n60549 = ~i_hbusreq1 & ~n60548;
  assign n60550 = ~n60543 & ~n60549;
  assign n60551 = ~controllable_hgrant1 & ~n60550;
  assign n60552 = ~n48683 & ~n60551;
  assign n60553 = ~i_hbusreq3 & ~n60552;
  assign n60554 = ~n60542 & ~n60553;
  assign n60555 = ~controllable_hgrant3 & ~n60554;
  assign n60556 = ~n48675 & ~n60555;
  assign n60557 = ~i_hbusreq9 & ~n60556;
  assign n60558 = ~n60541 & ~n60557;
  assign n60559 = ~i_hbusreq4 & ~n60558;
  assign n60560 = ~n60540 & ~n60559;
  assign n60561 = ~controllable_hgrant4 & ~n60560;
  assign n60562 = ~n48666 & ~n60561;
  assign n60563 = ~i_hbusreq5 & ~n60562;
  assign n60564 = ~n60539 & ~n60563;
  assign n60565 = ~controllable_hgrant5 & ~n60564;
  assign n60566 = ~n48655 & ~n60565;
  assign n60567 = ~controllable_hmaster2 & ~n60566;
  assign n60568 = ~n60538 & ~n60567;
  assign n60569 = ~controllable_hmaster1 & ~n60568;
  assign n60570 = ~n60537 & ~n60569;
  assign n60571 = ~i_hbusreq6 & ~n60570;
  assign n60572 = ~n60536 & ~n60571;
  assign n60573 = ~controllable_hgrant6 & ~n60572;
  assign n60574 = ~n59129 & ~n60573;
  assign n60575 = ~controllable_hmaster0 & ~n60574;
  assign n60576 = ~n60535 & ~n60575;
  assign n60577 = ~i_hbusreq8 & ~n60576;
  assign n60578 = ~n60530 & ~n60577;
  assign n60579 = ~controllable_hmaster3 & ~n60578;
  assign n60580 = ~n60529 & ~n60579;
  assign n60581 = ~i_hbusreq7 & ~n60580;
  assign n60582 = ~n60471 & ~n60581;
  assign n60583 = n7924 & ~n60582;
  assign n60584 = ~n60448 & ~n60583;
  assign n60585 = n8214 & ~n60584;
  assign n60586 = ~n60442 & ~n60585;
  assign n60587 = ~n8202 & ~n60586;
  assign n60588 = ~controllable_hgrant1 & ~n51364;
  assign n60589 = ~n60202 & ~n60588;
  assign n60590 = ~controllable_hgrant3 & ~n60589;
  assign n60591 = ~n51147 & ~n60590;
  assign n60592 = ~controllable_hgrant4 & ~n60591;
  assign n60593 = ~n50962 & ~n60592;
  assign n60594 = ~controllable_hgrant5 & ~n60593;
  assign n60595 = ~n50816 & ~n60594;
  assign n60596 = controllable_hmaster1 & ~n60595;
  assign n60597 = controllable_hmaster2 & ~n60595;
  assign n60598 = controllable_hmaster2 & ~n60597;
  assign n60599 = ~controllable_hmaster1 & ~n60598;
  assign n60600 = ~n60596 & ~n60599;
  assign n60601 = ~controllable_hgrant6 & ~n60600;
  assign n60602 = ~n41189 & ~n60601;
  assign n60603 = controllable_hmaster3 & ~n60602;
  assign n60604 = controllable_hmaster3 & ~n60603;
  assign n60605 = ~n7924 & ~n60604;
  assign n60606 = ~n49999 & ~n60605;
  assign n60607 = ~n8214 & ~n60606;
  assign n60608 = n8214 & ~n50000;
  assign n60609 = ~n60607 & ~n60608;
  assign n60610 = n8202 & ~n60609;
  assign n60611 = ~n60587 & ~n60610;
  assign n60612 = n7920 & ~n60611;
  assign n60613 = ~n60198 & ~n60612;
  assign n60614 = ~n7728 & ~n60613;
  assign n60615 = ~n60197 & ~n60614;
  assign n60616 = ~n7723 & ~n60615;
  assign n60617 = ~n7723 & ~n60616;
  assign n60618 = ~n7714 & ~n60617;
  assign n60619 = ~n7714 & ~n60618;
  assign n60620 = n7705 & ~n60619;
  assign n60621 = ~n41294 & ~n48017;
  assign n60622 = ~controllable_hgrant3 & ~n60621;
  assign n60623 = ~n13154 & ~n60622;
  assign n60624 = ~controllable_hgrant4 & ~n60623;
  assign n60625 = ~n13153 & ~n60624;
  assign n60626 = ~controllable_hgrant5 & ~n60625;
  assign n60627 = ~n13152 & ~n60626;
  assign n60628 = controllable_hmaster1 & ~n60627;
  assign n60629 = controllable_hmaster2 & ~n60627;
  assign n60630 = ~n41333 & ~n59181;
  assign n60631 = ~controllable_hgrant3 & ~n60630;
  assign n60632 = ~n13178 & ~n60631;
  assign n60633 = ~controllable_hgrant4 & ~n60632;
  assign n60634 = ~n13177 & ~n60633;
  assign n60635 = ~controllable_hgrant5 & ~n60634;
  assign n60636 = ~n13176 & ~n60635;
  assign n60637 = ~controllable_hmaster2 & ~n60636;
  assign n60638 = ~n60629 & ~n60637;
  assign n60639 = ~controllable_hmaster1 & ~n60638;
  assign n60640 = ~n60628 & ~n60639;
  assign n60641 = ~controllable_hgrant6 & ~n60640;
  assign n60642 = ~n13175 & ~n60641;
  assign n60643 = controllable_hmaster3 & ~n60642;
  assign n60644 = n8217 & ~n10830;
  assign n60645 = ~n8217 & ~n24282;
  assign n60646 = ~n60644 & ~n60645;
  assign n60647 = controllable_hgrant6 & ~n60646;
  assign n60648 = controllable_hmaster2 & ~n60636;
  assign n60649 = ~n41318 & ~n60631;
  assign n60650 = ~controllable_hgrant4 & ~n60649;
  assign n60651 = ~n13177 & ~n60650;
  assign n60652 = ~controllable_hgrant5 & ~n60651;
  assign n60653 = ~n13176 & ~n60652;
  assign n60654 = ~controllable_hmaster2 & ~n60653;
  assign n60655 = ~n60648 & ~n60654;
  assign n60656 = controllable_hmaster1 & ~n60655;
  assign n60657 = ~n41328 & ~n60635;
  assign n60658 = controllable_hmaster2 & ~n60657;
  assign n60659 = ~n48126 & ~n60658;
  assign n60660 = ~controllable_hmaster1 & ~n60659;
  assign n60661 = ~n60656 & ~n60660;
  assign n60662 = ~controllable_hgrant6 & ~n60661;
  assign n60663 = ~n60647 & ~n60662;
  assign n60664 = controllable_hmaster0 & ~n60663;
  assign n60665 = ~n41354 & ~n59181;
  assign n60666 = ~controllable_hgrant3 & ~n60665;
  assign n60667 = ~n13178 & ~n60666;
  assign n60668 = ~controllable_hgrant4 & ~n60667;
  assign n60669 = ~n13177 & ~n60668;
  assign n60670 = ~controllable_hgrant5 & ~n60669;
  assign n60671 = ~n13176 & ~n60670;
  assign n60672 = ~controllable_hmaster2 & ~n60671;
  assign n60673 = ~n60648 & ~n60672;
  assign n60674 = controllable_hmaster1 & ~n60673;
  assign n60675 = ~n41365 & ~n60633;
  assign n60676 = ~controllable_hgrant5 & ~n60675;
  assign n60677 = ~n13176 & ~n60676;
  assign n60678 = controllable_hmaster2 & ~n60677;
  assign n60679 = ~n60637 & ~n60678;
  assign n60680 = ~controllable_hmaster1 & ~n60679;
  assign n60681 = ~n60674 & ~n60680;
  assign n60682 = ~controllable_hgrant6 & ~n60681;
  assign n60683 = ~n41348 & ~n60682;
  assign n60684 = ~controllable_hmaster0 & ~n60683;
  assign n60685 = ~n60664 & ~n60684;
  assign n60686 = ~controllable_hmaster3 & ~n60685;
  assign n60687 = ~n60643 & ~n60686;
  assign n60688 = i_hbusreq7 & ~n60687;
  assign n60689 = i_hbusreq8 & ~n60642;
  assign n60690 = i_hbusreq6 & ~n60640;
  assign n60691 = i_hbusreq5 & ~n60625;
  assign n60692 = i_hbusreq4 & ~n60623;
  assign n60693 = i_hbusreq9 & ~n60623;
  assign n60694 = i_hbusreq3 & ~n60621;
  assign n60695 = ~n7757 & n8389;
  assign n60696 = ~n8389 & ~n17372;
  assign n60697 = ~n60695 & ~n60696;
  assign n60698 = ~i_hbusreq1 & ~n60697;
  assign n60699 = ~n48272 & ~n60698;
  assign n60700 = controllable_hgrant1 & ~n60699;
  assign n60701 = ~n41403 & ~n60700;
  assign n60702 = ~i_hbusreq3 & ~n60701;
  assign n60703 = ~n60694 & ~n60702;
  assign n60704 = ~controllable_hgrant3 & ~n60703;
  assign n60705 = ~n13211 & ~n60704;
  assign n60706 = ~i_hbusreq9 & ~n60705;
  assign n60707 = ~n60693 & ~n60706;
  assign n60708 = ~i_hbusreq4 & ~n60707;
  assign n60709 = ~n60692 & ~n60708;
  assign n60710 = ~controllable_hgrant4 & ~n60709;
  assign n60711 = ~n13208 & ~n60710;
  assign n60712 = ~i_hbusreq5 & ~n60711;
  assign n60713 = ~n60691 & ~n60712;
  assign n60714 = ~controllable_hgrant5 & ~n60713;
  assign n60715 = ~n13206 & ~n60714;
  assign n60716 = controllable_hmaster1 & ~n60715;
  assign n60717 = controllable_hmaster2 & ~n60715;
  assign n60718 = i_hbusreq5 & ~n60634;
  assign n60719 = i_hbusreq4 & ~n60632;
  assign n60720 = i_hbusreq9 & ~n60632;
  assign n60721 = i_hbusreq3 & ~n60630;
  assign n60722 = n8389 & ~n9013;
  assign n60723 = ~n8389 & ~n17416;
  assign n60724 = ~n60722 & ~n60723;
  assign n60725 = ~i_hbusreq1 & ~n60724;
  assign n60726 = ~n59360 & ~n60725;
  assign n60727 = controllable_hgrant1 & ~n60726;
  assign n60728 = ~n41472 & ~n60727;
  assign n60729 = ~i_hbusreq3 & ~n60728;
  assign n60730 = ~n60721 & ~n60729;
  assign n60731 = ~controllable_hgrant3 & ~n60730;
  assign n60732 = ~n13261 & ~n60731;
  assign n60733 = ~i_hbusreq9 & ~n60732;
  assign n60734 = ~n60720 & ~n60733;
  assign n60735 = ~i_hbusreq4 & ~n60734;
  assign n60736 = ~n60719 & ~n60735;
  assign n60737 = ~controllable_hgrant4 & ~n60736;
  assign n60738 = ~n13258 & ~n60737;
  assign n60739 = ~i_hbusreq5 & ~n60738;
  assign n60740 = ~n60718 & ~n60739;
  assign n60741 = ~controllable_hgrant5 & ~n60740;
  assign n60742 = ~n13256 & ~n60741;
  assign n60743 = ~controllable_hmaster2 & ~n60742;
  assign n60744 = ~n60717 & ~n60743;
  assign n60745 = ~controllable_hmaster1 & ~n60744;
  assign n60746 = ~n60716 & ~n60745;
  assign n60747 = ~i_hbusreq6 & ~n60746;
  assign n60748 = ~n60690 & ~n60747;
  assign n60749 = ~controllable_hgrant6 & ~n60748;
  assign n60750 = ~n13254 & ~n60749;
  assign n60751 = ~i_hbusreq8 & ~n60750;
  assign n60752 = ~n60689 & ~n60751;
  assign n60753 = controllable_hmaster3 & ~n60752;
  assign n60754 = i_hbusreq8 & ~n60685;
  assign n60755 = i_hbusreq6 & ~n60646;
  assign n60756 = n8217 & ~n10840;
  assign n60757 = ~n8217 & ~n24294;
  assign n60758 = ~n60756 & ~n60757;
  assign n60759 = ~i_hbusreq6 & ~n60758;
  assign n60760 = ~n60755 & ~n60759;
  assign n60761 = controllable_hgrant6 & ~n60760;
  assign n60762 = i_hbusreq6 & ~n60661;
  assign n60763 = controllable_hmaster2 & ~n60742;
  assign n60764 = i_hbusreq5 & ~n60651;
  assign n60765 = i_hbusreq4 & ~n60649;
  assign n60766 = i_hbusreq9 & ~n60649;
  assign n60767 = ~n41447 & ~n60731;
  assign n60768 = ~i_hbusreq9 & ~n60767;
  assign n60769 = ~n60766 & ~n60768;
  assign n60770 = ~i_hbusreq4 & ~n60769;
  assign n60771 = ~n60765 & ~n60770;
  assign n60772 = ~controllable_hgrant4 & ~n60771;
  assign n60773 = ~n13258 & ~n60772;
  assign n60774 = ~i_hbusreq5 & ~n60773;
  assign n60775 = ~n60764 & ~n60774;
  assign n60776 = ~controllable_hgrant5 & ~n60775;
  assign n60777 = ~n13256 & ~n60776;
  assign n60778 = ~controllable_hmaster2 & ~n60777;
  assign n60779 = ~n60763 & ~n60778;
  assign n60780 = controllable_hmaster1 & ~n60779;
  assign n60781 = ~n41463 & ~n60741;
  assign n60782 = controllable_hmaster2 & ~n60781;
  assign n60783 = ~n48496 & ~n60782;
  assign n60784 = ~controllable_hmaster1 & ~n60783;
  assign n60785 = ~n60780 & ~n60784;
  assign n60786 = ~i_hbusreq6 & ~n60785;
  assign n60787 = ~n60762 & ~n60786;
  assign n60788 = ~controllable_hgrant6 & ~n60787;
  assign n60789 = ~n60761 & ~n60788;
  assign n60790 = controllable_hmaster0 & ~n60789;
  assign n60791 = i_hbusreq6 & ~n60681;
  assign n60792 = i_hbusreq5 & ~n60669;
  assign n60793 = i_hbusreq4 & ~n60667;
  assign n60794 = i_hbusreq9 & ~n60667;
  assign n60795 = i_hbusreq3 & ~n60665;
  assign n60796 = ~n41511 & ~n60727;
  assign n60797 = ~i_hbusreq3 & ~n60796;
  assign n60798 = ~n60795 & ~n60797;
  assign n60799 = ~controllable_hgrant3 & ~n60798;
  assign n60800 = ~n13261 & ~n60799;
  assign n60801 = ~i_hbusreq9 & ~n60800;
  assign n60802 = ~n60794 & ~n60801;
  assign n60803 = ~i_hbusreq4 & ~n60802;
  assign n60804 = ~n60793 & ~n60803;
  assign n60805 = ~controllable_hgrant4 & ~n60804;
  assign n60806 = ~n13258 & ~n60805;
  assign n60807 = ~i_hbusreq5 & ~n60806;
  assign n60808 = ~n60792 & ~n60807;
  assign n60809 = ~controllable_hgrant5 & ~n60808;
  assign n60810 = ~n13256 & ~n60809;
  assign n60811 = ~controllable_hmaster2 & ~n60810;
  assign n60812 = ~n60763 & ~n60811;
  assign n60813 = controllable_hmaster1 & ~n60812;
  assign n60814 = i_hbusreq5 & ~n60675;
  assign n60815 = ~n41531 & ~n60737;
  assign n60816 = ~i_hbusreq5 & ~n60815;
  assign n60817 = ~n60814 & ~n60816;
  assign n60818 = ~controllable_hgrant5 & ~n60817;
  assign n60819 = ~n13256 & ~n60818;
  assign n60820 = controllable_hmaster2 & ~n60819;
  assign n60821 = ~n60743 & ~n60820;
  assign n60822 = ~controllable_hmaster1 & ~n60821;
  assign n60823 = ~n60813 & ~n60822;
  assign n60824 = ~i_hbusreq6 & ~n60823;
  assign n60825 = ~n60791 & ~n60824;
  assign n60826 = ~controllable_hgrant6 & ~n60825;
  assign n60827 = ~n41497 & ~n60826;
  assign n60828 = ~controllable_hmaster0 & ~n60827;
  assign n60829 = ~n60790 & ~n60828;
  assign n60830 = ~i_hbusreq8 & ~n60829;
  assign n60831 = ~n60754 & ~n60830;
  assign n60832 = ~controllable_hmaster3 & ~n60831;
  assign n60833 = ~n60753 & ~n60832;
  assign n60834 = ~i_hbusreq7 & ~n60833;
  assign n60835 = ~n60688 & ~n60834;
  assign n60836 = ~n7924 & ~n60835;
  assign n60837 = ~n41570 & ~n48793;
  assign n60838 = ~controllable_hgrant3 & ~n60837;
  assign n60839 = ~n41561 & ~n60838;
  assign n60840 = ~controllable_hgrant4 & ~n60839;
  assign n60841 = ~n41560 & ~n60840;
  assign n60842 = ~controllable_hgrant5 & ~n60841;
  assign n60843 = ~n41559 & ~n60842;
  assign n60844 = controllable_hmaster1 & ~n60843;
  assign n60845 = controllable_hmaster2 & ~n60843;
  assign n60846 = ~n41658 & ~n59650;
  assign n60847 = ~controllable_hgrant3 & ~n60846;
  assign n60848 = ~n41649 & ~n60847;
  assign n60849 = ~controllable_hgrant4 & ~n60848;
  assign n60850 = ~n41648 & ~n60849;
  assign n60851 = ~controllable_hgrant5 & ~n60850;
  assign n60852 = ~n41647 & ~n60851;
  assign n60853 = ~controllable_hmaster2 & ~n60852;
  assign n60854 = ~n60845 & ~n60853;
  assign n60855 = ~controllable_hmaster1 & ~n60854;
  assign n60856 = ~n60844 & ~n60855;
  assign n60857 = ~controllable_hgrant6 & ~n60856;
  assign n60858 = ~n41646 & ~n60857;
  assign n60859 = controllable_hmaster3 & ~n60858;
  assign n60860 = n8217 & ~n15893;
  assign n60861 = ~n8217 & ~n24322;
  assign n60862 = ~n60860 & ~n60861;
  assign n60863 = controllable_hgrant6 & ~n60862;
  assign n60864 = controllable_hmaster2 & ~n60852;
  assign n60865 = ~n41677 & ~n60847;
  assign n60866 = ~controllable_hgrant4 & ~n60865;
  assign n60867 = ~n41648 & ~n60866;
  assign n60868 = ~controllable_hgrant5 & ~n60867;
  assign n60869 = ~n41647 & ~n60868;
  assign n60870 = ~controllable_hmaster2 & ~n60869;
  assign n60871 = ~n60864 & ~n60870;
  assign n60872 = controllable_hmaster1 & ~n60871;
  assign n60873 = ~n41686 & ~n60851;
  assign n60874 = controllable_hmaster2 & ~n60873;
  assign n60875 = ~n8378 & ~n24316;
  assign n60876 = ~n43956 & ~n60875;
  assign n60877 = controllable_hgrant5 & ~n60876;
  assign n60878 = ~n8426 & ~n24314;
  assign n60879 = ~n43960 & ~n60878;
  assign n60880 = controllable_hgrant4 & ~n60879;
  assign n60881 = ~n8365 & ~n24312;
  assign n60882 = ~n43964 & ~n60881;
  assign n60883 = controllable_hgrant3 & ~n60882;
  assign n60884 = i_hlock1 & ~n41614;
  assign n60885 = ~i_hlock1 & ~n41628;
  assign n60886 = ~n60884 & ~n60885;
  assign n60887 = ~controllable_hgrant1 & ~n60886;
  assign n60888 = ~n48917 & ~n60887;
  assign n60889 = ~controllable_hgrant3 & ~n60888;
  assign n60890 = ~n60883 & ~n60889;
  assign n60891 = ~controllable_hgrant4 & ~n60890;
  assign n60892 = ~n60880 & ~n60891;
  assign n60893 = ~controllable_hgrant5 & ~n60892;
  assign n60894 = ~n60877 & ~n60893;
  assign n60895 = ~controllable_hmaster2 & ~n60894;
  assign n60896 = ~n60874 & ~n60895;
  assign n60897 = ~controllable_hmaster1 & ~n60896;
  assign n60898 = ~n60872 & ~n60897;
  assign n60899 = ~controllable_hgrant6 & ~n60898;
  assign n60900 = ~n60863 & ~n60899;
  assign n60901 = controllable_hmaster0 & ~n60900;
  assign n60902 = ~n41713 & ~n59650;
  assign n60903 = ~controllable_hgrant3 & ~n60902;
  assign n60904 = ~n41649 & ~n60903;
  assign n60905 = ~controllable_hgrant4 & ~n60904;
  assign n60906 = ~n41648 & ~n60905;
  assign n60907 = ~controllable_hgrant5 & ~n60906;
  assign n60908 = ~n41647 & ~n60907;
  assign n60909 = ~controllable_hmaster2 & ~n60908;
  assign n60910 = ~n60864 & ~n60909;
  assign n60911 = controllable_hmaster1 & ~n60910;
  assign n60912 = ~n41724 & ~n60849;
  assign n60913 = ~controllable_hgrant5 & ~n60912;
  assign n60914 = ~n41647 & ~n60913;
  assign n60915 = controllable_hmaster2 & ~n60914;
  assign n60916 = ~n60853 & ~n60915;
  assign n60917 = ~controllable_hmaster1 & ~n60916;
  assign n60918 = ~n60911 & ~n60917;
  assign n60919 = ~controllable_hgrant6 & ~n60918;
  assign n60920 = ~n41704 & ~n60919;
  assign n60921 = ~controllable_hmaster0 & ~n60920;
  assign n60922 = ~n60901 & ~n60921;
  assign n60923 = ~controllable_hmaster3 & ~n60922;
  assign n60924 = ~n60859 & ~n60923;
  assign n60925 = i_hbusreq7 & ~n60924;
  assign n60926 = i_hbusreq8 & ~n60858;
  assign n60927 = i_hbusreq6 & ~n60856;
  assign n60928 = i_hbusreq5 & ~n60841;
  assign n60929 = i_hbusreq4 & ~n60839;
  assign n60930 = i_hbusreq9 & ~n60839;
  assign n60931 = i_hbusreq3 & ~n60837;
  assign n60932 = n8389 & ~n13225;
  assign n60933 = ~n8389 & ~n17567;
  assign n60934 = ~n60932 & ~n60933;
  assign n60935 = i_hlock1 & ~n60934;
  assign n60936 = ~n8389 & ~n17589;
  assign n60937 = ~n60932 & ~n60936;
  assign n60938 = ~i_hlock1 & ~n60937;
  assign n60939 = ~n60935 & ~n60938;
  assign n60940 = ~i_hbusreq1 & ~n60939;
  assign n60941 = ~n49147 & ~n60940;
  assign n60942 = controllable_hgrant1 & ~n60941;
  assign n60943 = ~n41767 & ~n60942;
  assign n60944 = ~i_hbusreq3 & ~n60943;
  assign n60945 = ~n60931 & ~n60944;
  assign n60946 = ~controllable_hgrant3 & ~n60945;
  assign n60947 = ~n41753 & ~n60946;
  assign n60948 = ~i_hbusreq9 & ~n60947;
  assign n60949 = ~n60930 & ~n60948;
  assign n60950 = ~i_hbusreq4 & ~n60949;
  assign n60951 = ~n60929 & ~n60950;
  assign n60952 = ~controllable_hgrant4 & ~n60951;
  assign n60953 = ~n41750 & ~n60952;
  assign n60954 = ~i_hbusreq5 & ~n60953;
  assign n60955 = ~n60928 & ~n60954;
  assign n60956 = ~controllable_hgrant5 & ~n60955;
  assign n60957 = ~n41748 & ~n60956;
  assign n60958 = controllable_hmaster1 & ~n60957;
  assign n60959 = controllable_hmaster2 & ~n60957;
  assign n60960 = i_hbusreq5 & ~n60850;
  assign n60961 = i_hbusreq4 & ~n60848;
  assign n60962 = i_hbusreq9 & ~n60848;
  assign n60963 = i_hbusreq3 & ~n60846;
  assign n60964 = n8389 & ~n13265;
  assign n60965 = ~n8389 & ~n17642;
  assign n60966 = ~n60964 & ~n60965;
  assign n60967 = i_hlock1 & ~n60966;
  assign n60968 = ~n8389 & ~n17656;
  assign n60969 = ~n60964 & ~n60968;
  assign n60970 = ~i_hlock1 & ~n60969;
  assign n60971 = ~n60967 & ~n60970;
  assign n60972 = ~i_hbusreq1 & ~n60971;
  assign n60973 = ~n59898 & ~n60972;
  assign n60974 = controllable_hgrant1 & ~n60973;
  assign n60975 = ~n41932 & ~n60974;
  assign n60976 = ~i_hbusreq3 & ~n60975;
  assign n60977 = ~n60963 & ~n60976;
  assign n60978 = ~controllable_hgrant3 & ~n60977;
  assign n60979 = ~n41914 & ~n60978;
  assign n60980 = ~i_hbusreq9 & ~n60979;
  assign n60981 = ~n60962 & ~n60980;
  assign n60982 = ~i_hbusreq4 & ~n60981;
  assign n60983 = ~n60961 & ~n60982;
  assign n60984 = ~controllable_hgrant4 & ~n60983;
  assign n60985 = ~n41911 & ~n60984;
  assign n60986 = ~i_hbusreq5 & ~n60985;
  assign n60987 = ~n60960 & ~n60986;
  assign n60988 = ~controllable_hgrant5 & ~n60987;
  assign n60989 = ~n41909 & ~n60988;
  assign n60990 = ~controllable_hmaster2 & ~n60989;
  assign n60991 = ~n60959 & ~n60990;
  assign n60992 = ~controllable_hmaster1 & ~n60991;
  assign n60993 = ~n60958 & ~n60992;
  assign n60994 = ~i_hbusreq6 & ~n60993;
  assign n60995 = ~n60927 & ~n60994;
  assign n60996 = ~controllable_hgrant6 & ~n60995;
  assign n60997 = ~n41907 & ~n60996;
  assign n60998 = ~i_hbusreq8 & ~n60997;
  assign n60999 = ~n60926 & ~n60998;
  assign n61000 = controllable_hmaster3 & ~n60999;
  assign n61001 = i_hbusreq8 & ~n60922;
  assign n61002 = i_hbusreq6 & ~n60862;
  assign n61003 = n8217 & ~n15928;
  assign n61004 = ~n8217 & ~n24361;
  assign n61005 = ~n61003 & ~n61004;
  assign n61006 = ~i_hbusreq6 & ~n61005;
  assign n61007 = ~n61002 & ~n61006;
  assign n61008 = controllable_hgrant6 & ~n61007;
  assign n61009 = i_hbusreq6 & ~n60898;
  assign n61010 = controllable_hmaster2 & ~n60989;
  assign n61011 = i_hbusreq5 & ~n60867;
  assign n61012 = i_hbusreq4 & ~n60865;
  assign n61013 = i_hbusreq9 & ~n60865;
  assign n61014 = ~n41968 & ~n60978;
  assign n61015 = ~i_hbusreq9 & ~n61014;
  assign n61016 = ~n61013 & ~n61015;
  assign n61017 = ~i_hbusreq4 & ~n61016;
  assign n61018 = ~n61012 & ~n61017;
  assign n61019 = ~controllable_hgrant4 & ~n61018;
  assign n61020 = ~n41911 & ~n61019;
  assign n61021 = ~i_hbusreq5 & ~n61020;
  assign n61022 = ~n61011 & ~n61021;
  assign n61023 = ~controllable_hgrant5 & ~n61022;
  assign n61024 = ~n41909 & ~n61023;
  assign n61025 = ~controllable_hmaster2 & ~n61024;
  assign n61026 = ~n61010 & ~n61025;
  assign n61027 = controllable_hmaster1 & ~n61026;
  assign n61028 = ~n41983 & ~n60988;
  assign n61029 = controllable_hmaster2 & ~n61028;
  assign n61030 = i_hbusreq5 & ~n60876;
  assign n61031 = n8378 & ~n15920;
  assign n61032 = ~n8378 & ~n24353;
  assign n61033 = ~n61031 & ~n61032;
  assign n61034 = ~i_hbusreq5 & ~n61033;
  assign n61035 = ~n61030 & ~n61034;
  assign n61036 = controllable_hgrant5 & ~n61035;
  assign n61037 = i_hbusreq5 & ~n60892;
  assign n61038 = i_hbusreq4 & ~n60879;
  assign n61039 = i_hbusreq9 & ~n60879;
  assign n61040 = n8426 & ~n15914;
  assign n61041 = ~n8426 & ~n24347;
  assign n61042 = ~n61040 & ~n61041;
  assign n61043 = ~i_hbusreq9 & ~n61042;
  assign n61044 = ~n61039 & ~n61043;
  assign n61045 = ~i_hbusreq4 & ~n61044;
  assign n61046 = ~n61038 & ~n61045;
  assign n61047 = controllable_hgrant4 & ~n61046;
  assign n61048 = i_hbusreq4 & ~n60890;
  assign n61049 = i_hbusreq9 & ~n60890;
  assign n61050 = i_hbusreq3 & ~n60882;
  assign n61051 = n8365 & ~n15910;
  assign n61052 = ~n8365 & ~n24343;
  assign n61053 = ~n61051 & ~n61052;
  assign n61054 = ~i_hbusreq3 & ~n61053;
  assign n61055 = ~n61050 & ~n61054;
  assign n61056 = controllable_hgrant3 & ~n61055;
  assign n61057 = i_hbusreq3 & ~n60888;
  assign n61058 = i_hbusreq1 & ~n60886;
  assign n61059 = i_hlock1 & ~n41851;
  assign n61060 = ~i_hlock1 & ~n41877;
  assign n61061 = ~n61059 & ~n61060;
  assign n61062 = ~i_hbusreq1 & ~n61061;
  assign n61063 = ~n61058 & ~n61062;
  assign n61064 = ~controllable_hgrant1 & ~n61063;
  assign n61065 = ~n49636 & ~n61064;
  assign n61066 = ~i_hbusreq3 & ~n61065;
  assign n61067 = ~n61057 & ~n61066;
  assign n61068 = ~controllable_hgrant3 & ~n61067;
  assign n61069 = ~n61056 & ~n61068;
  assign n61070 = ~i_hbusreq9 & ~n61069;
  assign n61071 = ~n61049 & ~n61070;
  assign n61072 = ~i_hbusreq4 & ~n61071;
  assign n61073 = ~n61048 & ~n61072;
  assign n61074 = ~controllable_hgrant4 & ~n61073;
  assign n61075 = ~n61047 & ~n61074;
  assign n61076 = ~i_hbusreq5 & ~n61075;
  assign n61077 = ~n61037 & ~n61076;
  assign n61078 = ~controllable_hgrant5 & ~n61077;
  assign n61079 = ~n61036 & ~n61078;
  assign n61080 = ~controllable_hmaster2 & ~n61079;
  assign n61081 = ~n61029 & ~n61080;
  assign n61082 = ~controllable_hmaster1 & ~n61081;
  assign n61083 = ~n61027 & ~n61082;
  assign n61084 = ~i_hbusreq6 & ~n61083;
  assign n61085 = ~n61009 & ~n61084;
  assign n61086 = ~controllable_hgrant6 & ~n61085;
  assign n61087 = ~n61008 & ~n61086;
  assign n61088 = controllable_hmaster0 & ~n61087;
  assign n61089 = i_hbusreq6 & ~n60918;
  assign n61090 = i_hbusreq5 & ~n60906;
  assign n61091 = i_hbusreq4 & ~n60904;
  assign n61092 = i_hbusreq9 & ~n60904;
  assign n61093 = i_hbusreq3 & ~n60902;
  assign n61094 = ~n42032 & ~n60974;
  assign n61095 = ~i_hbusreq3 & ~n61094;
  assign n61096 = ~n61093 & ~n61095;
  assign n61097 = ~controllable_hgrant3 & ~n61096;
  assign n61098 = ~n41914 & ~n61097;
  assign n61099 = ~i_hbusreq9 & ~n61098;
  assign n61100 = ~n61092 & ~n61099;
  assign n61101 = ~i_hbusreq4 & ~n61100;
  assign n61102 = ~n61091 & ~n61101;
  assign n61103 = ~controllable_hgrant4 & ~n61102;
  assign n61104 = ~n41911 & ~n61103;
  assign n61105 = ~i_hbusreq5 & ~n61104;
  assign n61106 = ~n61090 & ~n61105;
  assign n61107 = ~controllable_hgrant5 & ~n61106;
  assign n61108 = ~n41909 & ~n61107;
  assign n61109 = ~controllable_hmaster2 & ~n61108;
  assign n61110 = ~n61010 & ~n61109;
  assign n61111 = controllable_hmaster1 & ~n61110;
  assign n61112 = i_hbusreq5 & ~n60912;
  assign n61113 = ~n42052 & ~n60984;
  assign n61114 = ~i_hbusreq5 & ~n61113;
  assign n61115 = ~n61112 & ~n61114;
  assign n61116 = ~controllable_hgrant5 & ~n61115;
  assign n61117 = ~n41909 & ~n61116;
  assign n61118 = controllable_hmaster2 & ~n61117;
  assign n61119 = ~n60990 & ~n61118;
  assign n61120 = ~controllable_hmaster1 & ~n61119;
  assign n61121 = ~n61111 & ~n61120;
  assign n61122 = ~i_hbusreq6 & ~n61121;
  assign n61123 = ~n61089 & ~n61122;
  assign n61124 = ~controllable_hgrant6 & ~n61123;
  assign n61125 = ~n42015 & ~n61124;
  assign n61126 = ~controllable_hmaster0 & ~n61125;
  assign n61127 = ~n61088 & ~n61126;
  assign n61128 = ~i_hbusreq8 & ~n61127;
  assign n61129 = ~n61001 & ~n61128;
  assign n61130 = ~controllable_hmaster3 & ~n61129;
  assign n61131 = ~n61000 & ~n61130;
  assign n61132 = ~i_hbusreq7 & ~n61131;
  assign n61133 = ~n60925 & ~n61132;
  assign n61134 = n7924 & ~n61133;
  assign n61135 = ~n60836 & ~n61134;
  assign n61136 = ~n8214 & ~n61135;
  assign n61137 = ~n10853 & ~n26890;
  assign n61138 = n8217 & ~n61137;
  assign n61139 = ~n24378 & ~n26890;
  assign n61140 = ~n8217 & ~n61139;
  assign n61141 = ~n61138 & ~n61140;
  assign n61142 = controllable_hgrant6 & ~n61141;
  assign n61143 = ~n41370 & ~n48207;
  assign n61144 = ~controllable_hmaster1 & ~n61143;
  assign n61145 = ~n41364 & ~n61144;
  assign n61146 = ~controllable_hgrant6 & ~n61145;
  assign n61147 = ~n61142 & ~n61146;
  assign n61148 = ~controllable_hmaster0 & ~n61147;
  assign n61149 = ~n41347 & ~n61148;
  assign n61150 = ~controllable_hmaster3 & ~n61149;
  assign n61151 = ~n42307 & ~n61150;
  assign n61152 = i_hbusreq7 & ~n61151;
  assign n61153 = ~n7823 & ~n12715;
  assign n61154 = ~n7928 & ~n61153;
  assign n61155 = ~n7938 & ~n12715;
  assign n61156 = n7928 & ~n61155;
  assign n61157 = ~n61154 & ~n61156;
  assign n61158 = ~i_hbusreq1 & ~n61157;
  assign n61159 = ~n41394 & ~n61158;
  assign n61160 = ~controllable_hgrant1 & ~n61159;
  assign n61161 = ~n14877 & ~n61160;
  assign n61162 = ~i_hbusreq3 & ~n61161;
  assign n61163 = ~n41393 & ~n61162;
  assign n61164 = ~controllable_hgrant3 & ~n61163;
  assign n61165 = ~n14876 & ~n61164;
  assign n61166 = ~i_hbusreq9 & ~n61165;
  assign n61167 = ~n41392 & ~n61166;
  assign n61168 = ~i_hbusreq4 & ~n61167;
  assign n61169 = ~n41391 & ~n61168;
  assign n61170 = ~controllable_hgrant4 & ~n61169;
  assign n61171 = ~n14875 & ~n61170;
  assign n61172 = ~i_hbusreq5 & ~n61171;
  assign n61173 = ~n41390 & ~n61172;
  assign n61174 = ~controllable_hgrant5 & ~n61173;
  assign n61175 = ~n14874 & ~n61174;
  assign n61176 = controllable_hmaster1 & ~n61175;
  assign n61177 = controllable_hmaster2 & ~n61175;
  assign n61178 = ~n10751 & ~n61177;
  assign n61179 = ~controllable_hmaster1 & ~n61178;
  assign n61180 = ~n61176 & ~n61179;
  assign n61181 = ~i_hbusreq6 & ~n61180;
  assign n61182 = ~n41429 & ~n61181;
  assign n61183 = ~controllable_hgrant6 & ~n61182;
  assign n61184 = ~n15946 & ~n61183;
  assign n61185 = ~i_hbusreq8 & ~n61184;
  assign n61186 = ~n42338 & ~n61185;
  assign n61187 = controllable_hmaster3 & ~n61186;
  assign n61188 = i_hbusreq8 & ~n61149;
  assign n61189 = controllable_hgrant3 & ~n15684;
  assign n61190 = ~controllable_hgrant3 & ~n10744;
  assign n61191 = ~n61189 & ~n61190;
  assign n61192 = ~i_hbusreq9 & ~n61191;
  assign n61193 = ~n41446 & ~n61192;
  assign n61194 = ~i_hbusreq4 & ~n61193;
  assign n61195 = ~n41445 & ~n61194;
  assign n61196 = ~controllable_hgrant4 & ~n61195;
  assign n61197 = ~n15675 & ~n61196;
  assign n61198 = ~i_hbusreq5 & ~n61197;
  assign n61199 = ~n41444 & ~n61198;
  assign n61200 = ~controllable_hgrant5 & ~n61199;
  assign n61201 = ~n15674 & ~n61200;
  assign n61202 = ~controllable_hmaster2 & ~n61201;
  assign n61203 = ~n10764 & ~n61202;
  assign n61204 = controllable_hmaster1 & ~n61203;
  assign n61205 = controllable_hgrant5 & ~n15694;
  assign n61206 = ~controllable_hgrant5 & ~n10750;
  assign n61207 = ~n61205 & ~n61206;
  assign n61208 = controllable_hmaster2 & ~n61207;
  assign n61209 = controllable_hgrant1 & ~n15680;
  assign n61210 = ~controllable_hgrant1 & ~n10742;
  assign n61211 = ~n61209 & ~n61210;
  assign n61212 = ~i_hbusreq3 & ~n61211;
  assign n61213 = ~n41470 & ~n61212;
  assign n61214 = ~controllable_hgrant3 & ~n61213;
  assign n61215 = ~n15676 & ~n61214;
  assign n61216 = ~i_hbusreq9 & ~n61215;
  assign n61217 = ~n41469 & ~n61216;
  assign n61218 = ~i_hbusreq4 & ~n61217;
  assign n61219 = ~n41468 & ~n61218;
  assign n61220 = ~controllable_hgrant4 & ~n61219;
  assign n61221 = ~n15675 & ~n61220;
  assign n61222 = ~i_hbusreq5 & ~n61221;
  assign n61223 = ~n41467 & ~n61222;
  assign n61224 = ~controllable_hgrant5 & ~n61223;
  assign n61225 = ~n15674 & ~n61224;
  assign n61226 = ~controllable_hmaster2 & ~n61225;
  assign n61227 = ~n61208 & ~n61226;
  assign n61228 = ~controllable_hmaster1 & ~n61227;
  assign n61229 = ~n61204 & ~n61228;
  assign n61230 = ~i_hbusreq6 & ~n61229;
  assign n61231 = ~n41443 & ~n61230;
  assign n61232 = ~controllable_hgrant6 & ~n61231;
  assign n61233 = ~n15812 & ~n61232;
  assign n61234 = controllable_hmaster0 & ~n61233;
  assign n61235 = i_hbusreq6 & ~n61141;
  assign n61236 = ~n10871 & ~n28100;
  assign n61237 = n8217 & ~n61236;
  assign n61238 = ~n24390 & ~n28100;
  assign n61239 = ~n8217 & ~n61238;
  assign n61240 = ~n61237 & ~n61239;
  assign n61241 = ~i_hbusreq6 & ~n61240;
  assign n61242 = ~n61235 & ~n61241;
  assign n61243 = controllable_hgrant6 & ~n61242;
  assign n61244 = i_hbusreq6 & ~n61145;
  assign n61245 = controllable_hgrant2 & ~n12702;
  assign n61246 = ~controllable_hgrant2 & ~n8679;
  assign n61247 = ~n61245 & ~n61246;
  assign n61248 = ~n7733 & ~n61247;
  assign n61249 = controllable_hgrant2 & ~n12712;
  assign n61250 = ~controllable_hgrant2 & ~n8686;
  assign n61251 = ~n61249 & ~n61250;
  assign n61252 = n7733 & ~n61251;
  assign n61253 = ~n61248 & ~n61252;
  assign n61254 = n7928 & ~n61253;
  assign n61255 = n7928 & ~n61254;
  assign n61256 = ~i_hbusreq1 & ~n61255;
  assign n61257 = ~n41503 & ~n61256;
  assign n61258 = ~controllable_hgrant1 & ~n61257;
  assign n61259 = ~n15677 & ~n61258;
  assign n61260 = ~i_hbusreq3 & ~n61259;
  assign n61261 = ~n41502 & ~n61260;
  assign n61262 = ~controllable_hgrant3 & ~n61261;
  assign n61263 = ~n15676 & ~n61262;
  assign n61264 = ~i_hbusreq9 & ~n61263;
  assign n61265 = ~n41501 & ~n61264;
  assign n61266 = ~i_hbusreq4 & ~n61265;
  assign n61267 = ~n41500 & ~n61266;
  assign n61268 = ~controllable_hgrant4 & ~n61267;
  assign n61269 = ~n15675 & ~n61268;
  assign n61270 = ~i_hbusreq5 & ~n61269;
  assign n61271 = ~n41499 & ~n61270;
  assign n61272 = ~controllable_hgrant5 & ~n61271;
  assign n61273 = ~n15674 & ~n61272;
  assign n61274 = ~controllable_hmaster2 & ~n61273;
  assign n61275 = ~n10764 & ~n61274;
  assign n61276 = controllable_hmaster1 & ~n61275;
  assign n61277 = controllable_hgrant4 & ~n15690;
  assign n61278 = ~controllable_hgrant4 & ~n10748;
  assign n61279 = ~n61277 & ~n61278;
  assign n61280 = ~i_hbusreq5 & ~n61279;
  assign n61281 = ~n41530 & ~n61280;
  assign n61282 = ~controllable_hgrant5 & ~n61281;
  assign n61283 = ~n15674 & ~n61282;
  assign n61284 = controllable_hmaster2 & ~n61283;
  assign n61285 = ~n48715 & ~n61284;
  assign n61286 = ~controllable_hmaster1 & ~n61285;
  assign n61287 = ~n61276 & ~n61286;
  assign n61288 = ~i_hbusreq6 & ~n61287;
  assign n61289 = ~n61244 & ~n61288;
  assign n61290 = ~controllable_hgrant6 & ~n61289;
  assign n61291 = ~n61243 & ~n61290;
  assign n61292 = ~controllable_hmaster0 & ~n61291;
  assign n61293 = ~n61234 & ~n61292;
  assign n61294 = ~i_hbusreq8 & ~n61293;
  assign n61295 = ~n61188 & ~n61294;
  assign n61296 = ~controllable_hmaster3 & ~n61295;
  assign n61297 = ~n61187 & ~n61296;
  assign n61298 = ~i_hbusreq7 & ~n61297;
  assign n61299 = ~n61152 & ~n61298;
  assign n61300 = ~n7924 & ~n61299;
  assign n61301 = ~n15966 & ~n26936;
  assign n61302 = n8217 & ~n61301;
  assign n61303 = ~n24416 & ~n26936;
  assign n61304 = ~n8217 & ~n61303;
  assign n61305 = ~n61302 & ~n61304;
  assign n61306 = controllable_hgrant6 & ~n61305;
  assign n61307 = ~n8378 & ~n24411;
  assign n61308 = ~n44076 & ~n61307;
  assign n61309 = controllable_hgrant5 & ~n61308;
  assign n61310 = ~n8426 & ~n24409;
  assign n61311 = ~n44080 & ~n61310;
  assign n61312 = controllable_hgrant4 & ~n61311;
  assign n61313 = ~n8365 & ~n24407;
  assign n61314 = ~n44084 & ~n61313;
  assign n61315 = controllable_hgrant3 & ~n61314;
  assign n61316 = ~n8389 & ~n24405;
  assign n61317 = ~n44088 & ~n61316;
  assign n61318 = controllable_hgrant1 & ~n61317;
  assign n61319 = ~n8440 & ~n41613;
  assign n61320 = ~controllable_hgrant1 & ~n61319;
  assign n61321 = ~n61318 & ~n61320;
  assign n61322 = ~controllable_hgrant3 & ~n61321;
  assign n61323 = ~n61315 & ~n61322;
  assign n61324 = ~controllable_hgrant4 & ~n61323;
  assign n61325 = ~n61312 & ~n61324;
  assign n61326 = ~controllable_hgrant5 & ~n61325;
  assign n61327 = ~n61309 & ~n61326;
  assign n61328 = ~controllable_hmaster2 & ~n61327;
  assign n61329 = ~n41728 & ~n61328;
  assign n61330 = ~controllable_hmaster1 & ~n61329;
  assign n61331 = ~n41723 & ~n61330;
  assign n61332 = ~controllable_hgrant6 & ~n61331;
  assign n61333 = ~n61306 & ~n61332;
  assign n61334 = ~controllable_hmaster0 & ~n61333;
  assign n61335 = ~n41703 & ~n61334;
  assign n61336 = ~controllable_hmaster3 & ~n61335;
  assign n61337 = ~n42392 & ~n61336;
  assign n61338 = i_hbusreq7 & ~n61337;
  assign n61339 = controllable_hgrant6 & ~n15987;
  assign n61340 = controllable_hgrant5 & ~n14914;
  assign n61341 = controllable_hgrant4 & ~n14910;
  assign n61342 = controllable_hgrant3 & ~n14904;
  assign n61343 = controllable_hgrant1 & ~n14900;
  assign n61344 = controllable_hgrant2 & ~n14884;
  assign n61345 = ~n49177 & ~n61344;
  assign n61346 = ~n7733 & ~n61345;
  assign n61347 = controllable_hgrant2 & ~n14892;
  assign n61348 = ~n12904 & ~n61347;
  assign n61349 = n7733 & ~n61348;
  assign n61350 = ~n61346 & ~n61349;
  assign n61351 = n7928 & ~n61350;
  assign n61352 = ~n61154 & ~n61351;
  assign n61353 = ~i_hbusreq1 & ~n61352;
  assign n61354 = ~n41756 & ~n61353;
  assign n61355 = ~controllable_hgrant1 & ~n61354;
  assign n61356 = ~n61343 & ~n61355;
  assign n61357 = ~i_hbusreq3 & ~n61356;
  assign n61358 = ~n41754 & ~n61357;
  assign n61359 = ~controllable_hgrant3 & ~n61358;
  assign n61360 = ~n61342 & ~n61359;
  assign n61361 = ~i_hbusreq9 & ~n61360;
  assign n61362 = ~n41752 & ~n61361;
  assign n61363 = ~i_hbusreq4 & ~n61362;
  assign n61364 = ~n41751 & ~n61363;
  assign n61365 = ~controllable_hgrant4 & ~n61364;
  assign n61366 = ~n61341 & ~n61365;
  assign n61367 = ~i_hbusreq5 & ~n61366;
  assign n61368 = ~n41749 & ~n61367;
  assign n61369 = ~controllable_hgrant5 & ~n61368;
  assign n61370 = ~n61340 & ~n61369;
  assign n61371 = controllable_hmaster1 & ~n61370;
  assign n61372 = controllable_hmaster2 & ~n61370;
  assign n61373 = controllable_hgrant5 & ~n15796;
  assign n61374 = controllable_hgrant4 & ~n15792;
  assign n61375 = controllable_hgrant3 & ~n15786;
  assign n61376 = controllable_hgrant1 & ~n15782;
  assign n61377 = controllable_hgrant2 & ~n13975;
  assign n61378 = i_hlock0 & ~n16485;
  assign n61379 = ~n16787 & ~n20624;
  assign n61380 = ~i_hlock0 & ~n61379;
  assign n61381 = ~n61378 & ~n61380;
  assign n61382 = ~i_hbusreq0 & ~n61381;
  assign n61383 = ~n41919 & ~n61382;
  assign n61384 = ~i_hbusreq2 & ~n61383;
  assign n61385 = ~n41918 & ~n61384;
  assign n61386 = ~controllable_hgrant2 & n61385;
  assign n61387 = ~n61377 & ~n61386;
  assign n61388 = ~n7733 & ~n61387;
  assign n61389 = n7733 & ~n14892;
  assign n61390 = ~n61388 & ~n61389;
  assign n61391 = n7928 & ~n61390;
  assign n61392 = n7928 & ~n61391;
  assign n61393 = ~i_hbusreq1 & ~n61392;
  assign n61394 = ~n41917 & ~n61393;
  assign n61395 = ~controllable_hgrant1 & ~n61394;
  assign n61396 = ~n61376 & ~n61395;
  assign n61397 = ~i_hbusreq3 & ~n61396;
  assign n61398 = ~n41915 & ~n61397;
  assign n61399 = ~controllable_hgrant3 & ~n61398;
  assign n61400 = ~n61375 & ~n61399;
  assign n61401 = ~i_hbusreq9 & ~n61400;
  assign n61402 = ~n41913 & ~n61401;
  assign n61403 = ~i_hbusreq4 & ~n61402;
  assign n61404 = ~n41912 & ~n61403;
  assign n61405 = ~controllable_hgrant4 & ~n61404;
  assign n61406 = ~n61374 & ~n61405;
  assign n61407 = ~i_hbusreq5 & ~n61406;
  assign n61408 = ~n41910 & ~n61407;
  assign n61409 = ~controllable_hgrant5 & ~n61408;
  assign n61410 = ~n61373 & ~n61409;
  assign n61411 = ~controllable_hmaster2 & ~n61410;
  assign n61412 = ~n61372 & ~n61411;
  assign n61413 = ~controllable_hmaster1 & ~n61412;
  assign n61414 = ~n61371 & ~n61413;
  assign n61415 = ~i_hbusreq6 & ~n61414;
  assign n61416 = ~n41908 & ~n61415;
  assign n61417 = ~controllable_hgrant6 & ~n61416;
  assign n61418 = ~n61339 & ~n61417;
  assign n61419 = ~i_hbusreq8 & ~n61418;
  assign n61420 = ~n42425 & ~n61419;
  assign n61421 = controllable_hmaster3 & ~n61420;
  assign n61422 = i_hbusreq8 & ~n61335;
  assign n61423 = controllable_hgrant6 & ~n15814;
  assign n61424 = controllable_hmaster2 & ~n61410;
  assign n61425 = controllable_hgrant3 & ~n15758;
  assign n61426 = ~n61399 & ~n61425;
  assign n61427 = ~i_hbusreq9 & ~n61426;
  assign n61428 = ~n41967 & ~n61427;
  assign n61429 = ~i_hbusreq4 & ~n61428;
  assign n61430 = ~n41966 & ~n61429;
  assign n61431 = ~controllable_hgrant4 & ~n61430;
  assign n61432 = ~n61374 & ~n61431;
  assign n61433 = ~i_hbusreq5 & ~n61432;
  assign n61434 = ~n41965 & ~n61433;
  assign n61435 = ~controllable_hgrant5 & ~n61434;
  assign n61436 = ~n61373 & ~n61435;
  assign n61437 = ~controllable_hmaster2 & ~n61436;
  assign n61438 = ~n61424 & ~n61437;
  assign n61439 = controllable_hmaster1 & ~n61438;
  assign n61440 = controllable_hgrant5 & ~n15768;
  assign n61441 = ~n61409 & ~n61440;
  assign n61442 = controllable_hmaster2 & ~n61441;
  assign n61443 = controllable_hgrant1 & ~n15754;
  assign n61444 = ~n61395 & ~n61443;
  assign n61445 = ~i_hbusreq3 & ~n61444;
  assign n61446 = ~n41989 & ~n61445;
  assign n61447 = ~controllable_hgrant3 & ~n61446;
  assign n61448 = ~n61375 & ~n61447;
  assign n61449 = ~i_hbusreq9 & ~n61448;
  assign n61450 = ~n41988 & ~n61449;
  assign n61451 = ~i_hbusreq4 & ~n61450;
  assign n61452 = ~n41987 & ~n61451;
  assign n61453 = ~controllable_hgrant4 & ~n61452;
  assign n61454 = ~n61374 & ~n61453;
  assign n61455 = ~i_hbusreq5 & ~n61454;
  assign n61456 = ~n41986 & ~n61455;
  assign n61457 = ~controllable_hgrant5 & ~n61456;
  assign n61458 = ~n61373 & ~n61457;
  assign n61459 = ~controllable_hmaster2 & ~n61458;
  assign n61460 = ~n61442 & ~n61459;
  assign n61461 = ~controllable_hmaster1 & ~n61460;
  assign n61462 = ~n61439 & ~n61461;
  assign n61463 = ~i_hbusreq6 & ~n61462;
  assign n61464 = ~n41963 & ~n61463;
  assign n61465 = ~controllable_hgrant6 & ~n61464;
  assign n61466 = ~n61423 & ~n61465;
  assign n61467 = controllable_hmaster0 & ~n61466;
  assign n61468 = i_hbusreq6 & ~n61305;
  assign n61469 = ~n15999 & ~n28124;
  assign n61470 = n8217 & ~n61469;
  assign n61471 = ~n24464 & ~n28124;
  assign n61472 = ~n8217 & ~n61471;
  assign n61473 = ~n61470 & ~n61472;
  assign n61474 = ~i_hbusreq6 & ~n61473;
  assign n61475 = ~n61468 & ~n61474;
  assign n61476 = controllable_hgrant6 & ~n61475;
  assign n61477 = i_hbusreq6 & ~n61331;
  assign n61478 = controllable_hgrant2 & ~n12890;
  assign n61479 = ~n61386 & ~n61478;
  assign n61480 = ~n7733 & ~n61479;
  assign n61481 = controllable_hgrant2 & ~n12903;
  assign n61482 = ~n14893 & ~n61481;
  assign n61483 = n7733 & ~n61482;
  assign n61484 = ~n61480 & ~n61483;
  assign n61485 = n7928 & ~n61484;
  assign n61486 = n7928 & ~n61485;
  assign n61487 = ~i_hbusreq1 & ~n61486;
  assign n61488 = ~n42021 & ~n61487;
  assign n61489 = ~controllable_hgrant1 & ~n61488;
  assign n61490 = ~n61376 & ~n61489;
  assign n61491 = ~i_hbusreq3 & ~n61490;
  assign n61492 = ~n42020 & ~n61491;
  assign n61493 = ~controllable_hgrant3 & ~n61492;
  assign n61494 = ~n61375 & ~n61493;
  assign n61495 = ~i_hbusreq9 & ~n61494;
  assign n61496 = ~n42019 & ~n61495;
  assign n61497 = ~i_hbusreq4 & ~n61496;
  assign n61498 = ~n42018 & ~n61497;
  assign n61499 = ~controllable_hgrant4 & ~n61498;
  assign n61500 = ~n61374 & ~n61499;
  assign n61501 = ~i_hbusreq5 & ~n61500;
  assign n61502 = ~n42017 & ~n61501;
  assign n61503 = ~controllable_hgrant5 & ~n61502;
  assign n61504 = ~n61373 & ~n61503;
  assign n61505 = ~controllable_hmaster2 & ~n61504;
  assign n61506 = ~n61424 & ~n61505;
  assign n61507 = controllable_hmaster1 & ~n61506;
  assign n61508 = controllable_hgrant4 & ~n15764;
  assign n61509 = ~n61405 & ~n61508;
  assign n61510 = ~i_hbusreq5 & ~n61509;
  assign n61511 = ~n42051 & ~n61510;
  assign n61512 = ~controllable_hgrant5 & ~n61511;
  assign n61513 = ~n61373 & ~n61512;
  assign n61514 = controllable_hmaster2 & ~n61513;
  assign n61515 = i_hbusreq5 & ~n61308;
  assign n61516 = ~n8378 & ~n24457;
  assign n61517 = ~n49843 & ~n61516;
  assign n61518 = ~i_hbusreq5 & ~n61517;
  assign n61519 = ~n61515 & ~n61518;
  assign n61520 = controllable_hgrant5 & ~n61519;
  assign n61521 = i_hbusreq5 & ~n61325;
  assign n61522 = i_hbusreq4 & ~n61311;
  assign n61523 = i_hbusreq9 & ~n61311;
  assign n61524 = ~n8426 & ~n24451;
  assign n61525 = ~n49857 & ~n61524;
  assign n61526 = ~i_hbusreq9 & ~n61525;
  assign n61527 = ~n61523 & ~n61526;
  assign n61528 = ~i_hbusreq4 & ~n61527;
  assign n61529 = ~n61522 & ~n61528;
  assign n61530 = controllable_hgrant4 & ~n61529;
  assign n61531 = i_hbusreq4 & ~n61323;
  assign n61532 = i_hbusreq9 & ~n61323;
  assign n61533 = i_hbusreq3 & ~n61314;
  assign n61534 = ~n8365 & ~n24447;
  assign n61535 = ~n49876 & ~n61534;
  assign n61536 = ~i_hbusreq3 & ~n61535;
  assign n61537 = ~n61533 & ~n61536;
  assign n61538 = controllable_hgrant3 & ~n61537;
  assign n61539 = i_hbusreq3 & ~n61321;
  assign n61540 = i_hbusreq1 & ~n61317;
  assign n61541 = ~n8389 & ~n24443;
  assign n61542 = ~n49889 & ~n61541;
  assign n61543 = ~i_hbusreq1 & ~n61542;
  assign n61544 = ~n61540 & ~n61543;
  assign n61545 = controllable_hgrant1 & ~n61544;
  assign n61546 = i_hbusreq1 & ~n61319;
  assign n61547 = ~i_hlock0 & ~n41603;
  assign n61548 = ~n43663 & ~n61547;
  assign n61549 = ~i_hbusreq0 & ~n61548;
  assign n61550 = ~n41828 & ~n61549;
  assign n61551 = ~i_hbusreq2 & ~n61550;
  assign n61552 = ~n41827 & ~n61551;
  assign n61553 = controllable_hgrant2 & ~n61552;
  assign n61554 = ~n49909 & ~n61553;
  assign n61555 = ~n7733 & ~n61554;
  assign n61556 = ~n41611 & ~n61555;
  assign n61557 = n7928 & ~n61556;
  assign n61558 = ~n8440 & ~n61557;
  assign n61559 = ~i_hbusreq1 & ~n61558;
  assign n61560 = ~n61546 & ~n61559;
  assign n61561 = ~controllable_hgrant1 & ~n61560;
  assign n61562 = ~n61545 & ~n61561;
  assign n61563 = ~i_hbusreq3 & ~n61562;
  assign n61564 = ~n61539 & ~n61563;
  assign n61565 = ~controllable_hgrant3 & ~n61564;
  assign n61566 = ~n61538 & ~n61565;
  assign n61567 = ~i_hbusreq9 & ~n61566;
  assign n61568 = ~n61532 & ~n61567;
  assign n61569 = ~i_hbusreq4 & ~n61568;
  assign n61570 = ~n61531 & ~n61569;
  assign n61571 = ~controllable_hgrant4 & ~n61570;
  assign n61572 = ~n61530 & ~n61571;
  assign n61573 = ~i_hbusreq5 & ~n61572;
  assign n61574 = ~n61521 & ~n61573;
  assign n61575 = ~controllable_hgrant5 & ~n61574;
  assign n61576 = ~n61520 & ~n61575;
  assign n61577 = ~controllable_hmaster2 & ~n61576;
  assign n61578 = ~n61514 & ~n61577;
  assign n61579 = ~controllable_hmaster1 & ~n61578;
  assign n61580 = ~n61507 & ~n61579;
  assign n61581 = ~i_hbusreq6 & ~n61580;
  assign n61582 = ~n61477 & ~n61581;
  assign n61583 = ~controllable_hgrant6 & ~n61582;
  assign n61584 = ~n61476 & ~n61583;
  assign n61585 = ~controllable_hmaster0 & ~n61584;
  assign n61586 = ~n61467 & ~n61585;
  assign n61587 = ~i_hbusreq8 & ~n61586;
  assign n61588 = ~n61422 & ~n61587;
  assign n61589 = ~controllable_hmaster3 & ~n61588;
  assign n61590 = ~n61421 & ~n61589;
  assign n61591 = ~i_hbusreq7 & ~n61590;
  assign n61592 = ~n61338 & ~n61591;
  assign n61593 = n7924 & ~n61592;
  assign n61594 = ~n61300 & ~n61593;
  assign n61595 = n8214 & ~n61594;
  assign n61596 = ~n61136 & ~n61595;
  assign n61597 = ~n8202 & ~n61596;
  assign n61598 = n8202 & ~n50000;
  assign n61599 = ~n61597 & ~n61598;
  assign n61600 = n7920 & ~n61599;
  assign n61601 = ~n60198 & ~n61600;
  assign n61602 = n7728 & ~n61601;
  assign n61603 = ~n42730 & ~n48017;
  assign n61604 = ~controllable_hgrant3 & ~n61603;
  assign n61605 = ~n42717 & ~n61604;
  assign n61606 = ~controllable_hgrant4 & ~n61605;
  assign n61607 = ~n42713 & ~n61606;
  assign n61608 = ~controllable_hgrant5 & ~n61607;
  assign n61609 = ~n42709 & ~n61608;
  assign n61610 = controllable_hmaster1 & ~n61609;
  assign n61611 = controllable_hmaster2 & ~n61609;
  assign n61612 = ~n40214 & ~n42764;
  assign n61613 = ~controllable_hgrant3 & ~n61612;
  assign n61614 = ~n42757 & ~n61613;
  assign n61615 = i_hlock9 & ~n61614;
  assign n61616 = ~n40244 & ~n42797;
  assign n61617 = ~controllable_hgrant3 & ~n61616;
  assign n61618 = ~n42792 & ~n61617;
  assign n61619 = ~i_hlock9 & ~n61618;
  assign n61620 = ~n61615 & ~n61619;
  assign n61621 = ~controllable_hgrant4 & ~n61620;
  assign n61622 = ~n44951 & ~n61621;
  assign n61623 = ~controllable_hgrant5 & ~n61622;
  assign n61624 = ~n44947 & ~n61623;
  assign n61625 = ~controllable_hmaster2 & ~n61624;
  assign n61626 = ~n61611 & ~n61625;
  assign n61627 = ~controllable_hmaster1 & ~n61626;
  assign n61628 = ~n61610 & ~n61627;
  assign n61629 = ~controllable_hgrant6 & ~n61628;
  assign n61630 = ~n44944 & ~n61629;
  assign n61631 = controllable_hmaster0 & ~n61630;
  assign n61632 = ~controllable_hgrant4 & ~n61614;
  assign n61633 = ~n42754 & ~n61632;
  assign n61634 = ~controllable_hgrant5 & ~n61633;
  assign n61635 = ~n42751 & ~n61634;
  assign n61636 = ~controllable_hmaster2 & ~n61635;
  assign n61637 = ~n61611 & ~n61636;
  assign n61638 = ~controllable_hmaster1 & ~n61637;
  assign n61639 = ~n61610 & ~n61638;
  assign n61640 = ~controllable_hgrant6 & ~n61639;
  assign n61641 = ~n42748 & ~n61640;
  assign n61642 = ~controllable_hmaster0 & ~n61641;
  assign n61643 = ~n61631 & ~n61642;
  assign n61644 = i_hlock8 & ~n61643;
  assign n61645 = ~controllable_hgrant4 & ~n61618;
  assign n61646 = ~n42789 & ~n61645;
  assign n61647 = ~controllable_hgrant5 & ~n61646;
  assign n61648 = ~n42786 & ~n61647;
  assign n61649 = ~controllable_hmaster2 & ~n61648;
  assign n61650 = ~n61611 & ~n61649;
  assign n61651 = ~controllable_hmaster1 & ~n61650;
  assign n61652 = ~n61610 & ~n61651;
  assign n61653 = ~controllable_hgrant6 & ~n61652;
  assign n61654 = ~n42783 & ~n61653;
  assign n61655 = ~controllable_hmaster0 & ~n61654;
  assign n61656 = ~n61631 & ~n61655;
  assign n61657 = ~i_hlock8 & ~n61656;
  assign n61658 = ~n61644 & ~n61657;
  assign n61659 = controllable_hmaster3 & ~n61658;
  assign n61660 = ~n8217 & ~n24490;
  assign n61661 = ~n42816 & ~n61660;
  assign n61662 = controllable_hgrant6 & ~n61661;
  assign n61663 = controllable_hmaster2 & ~n61635;
  assign n61664 = i_hlock3 & ~n61612;
  assign n61665 = ~i_hlock3 & ~n61616;
  assign n61666 = ~n61664 & ~n61665;
  assign n61667 = ~controllable_hgrant3 & ~n61666;
  assign n61668 = ~n42838 & ~n61667;
  assign n61669 = ~controllable_hgrant4 & ~n61668;
  assign n61670 = ~n42828 & ~n61669;
  assign n61671 = ~controllable_hgrant5 & ~n61670;
  assign n61672 = ~n42824 & ~n61671;
  assign n61673 = ~controllable_hmaster2 & ~n61672;
  assign n61674 = ~n61663 & ~n61673;
  assign n61675 = controllable_hmaster1 & ~n61674;
  assign n61676 = i_hlock5 & ~n61633;
  assign n61677 = ~i_hlock5 & ~n61646;
  assign n61678 = ~n61676 & ~n61677;
  assign n61679 = ~controllable_hgrant5 & ~n61678;
  assign n61680 = ~n42860 & ~n61679;
  assign n61681 = controllable_hmaster2 & ~n61680;
  assign n61682 = ~n48126 & ~n61681;
  assign n61683 = ~controllable_hmaster1 & ~n61682;
  assign n61684 = ~n61675 & ~n61683;
  assign n61685 = ~controllable_hgrant6 & ~n61684;
  assign n61686 = ~n61662 & ~n61685;
  assign n61687 = controllable_hmaster0 & ~n61686;
  assign n61688 = ~n42976 & ~n48144;
  assign n61689 = ~controllable_hgrant3 & ~n61688;
  assign n61690 = ~n42940 & ~n61689;
  assign n61691 = ~controllable_hgrant4 & ~n61690;
  assign n61692 = ~n42936 & ~n61691;
  assign n61693 = ~controllable_hgrant5 & ~n61692;
  assign n61694 = ~n42932 & ~n61693;
  assign n61695 = ~controllable_hmaster2 & ~n61694;
  assign n61696 = ~n61663 & ~n61695;
  assign n61697 = controllable_hmaster1 & ~n61696;
  assign n61698 = i_hlock4 & ~n61614;
  assign n61699 = ~i_hlock4 & ~n61618;
  assign n61700 = ~n61698 & ~n61699;
  assign n61701 = ~controllable_hgrant4 & ~n61700;
  assign n61702 = ~n43000 & ~n61701;
  assign n61703 = ~controllable_hgrant5 & ~n61702;
  assign n61704 = ~n42990 & ~n61703;
  assign n61705 = controllable_hmaster2 & ~n61704;
  assign n61706 = ~n43026 & ~n48197;
  assign n61707 = ~controllable_hgrant3 & ~n61706;
  assign n61708 = ~n43020 & ~n61707;
  assign n61709 = ~controllable_hgrant4 & ~n61708;
  assign n61710 = ~n43016 & ~n61709;
  assign n61711 = ~controllable_hgrant5 & ~n61710;
  assign n61712 = ~n43012 & ~n61711;
  assign n61713 = ~controllable_hmaster2 & ~n61712;
  assign n61714 = ~n61705 & ~n61713;
  assign n61715 = ~controllable_hmaster1 & ~n61714;
  assign n61716 = ~n61697 & ~n61715;
  assign n61717 = i_hlock6 & ~n61716;
  assign n61718 = controllable_hmaster2 & ~n61648;
  assign n61719 = ~n61695 & ~n61718;
  assign n61720 = controllable_hmaster1 & ~n61719;
  assign n61721 = ~n61715 & ~n61720;
  assign n61722 = ~i_hlock6 & ~n61721;
  assign n61723 = ~n61717 & ~n61722;
  assign n61724 = ~controllable_hgrant6 & ~n61723;
  assign n61725 = ~n42928 & ~n61724;
  assign n61726 = ~controllable_hmaster0 & ~n61725;
  assign n61727 = ~n61687 & ~n61726;
  assign n61728 = ~controllable_hmaster3 & ~n61727;
  assign n61729 = ~n61659 & ~n61728;
  assign n61730 = i_hlock7 & ~n61729;
  assign n61731 = ~n8217 & ~n24498;
  assign n61732 = ~n43052 & ~n61731;
  assign n61733 = controllable_hgrant6 & ~n61732;
  assign n61734 = ~n61673 & ~n61718;
  assign n61735 = controllable_hmaster1 & ~n61734;
  assign n61736 = ~n61683 & ~n61735;
  assign n61737 = ~controllable_hgrant6 & ~n61736;
  assign n61738 = ~n61733 & ~n61737;
  assign n61739 = controllable_hmaster0 & ~n61738;
  assign n61740 = ~n61726 & ~n61739;
  assign n61741 = ~controllable_hmaster3 & ~n61740;
  assign n61742 = ~n61659 & ~n61741;
  assign n61743 = ~i_hlock7 & ~n61742;
  assign n61744 = ~n61730 & ~n61743;
  assign n61745 = i_hbusreq7 & ~n61744;
  assign n61746 = i_hbusreq8 & ~n61658;
  assign n61747 = i_hbusreq6 & ~n61628;
  assign n61748 = i_hbusreq5 & ~n61607;
  assign n61749 = i_hbusreq4 & ~n61605;
  assign n61750 = i_hbusreq9 & ~n61605;
  assign n61751 = i_hbusreq3 & ~n61603;
  assign n61752 = ~n8389 & ~n18228;
  assign n61753 = ~n43106 & ~n61752;
  assign n61754 = ~i_hbusreq1 & ~n61753;
  assign n61755 = ~n48272 & ~n61754;
  assign n61756 = controllable_hgrant1 & ~n61755;
  assign n61757 = ~n43130 & ~n61756;
  assign n61758 = ~i_hbusreq3 & ~n61757;
  assign n61759 = ~n61751 & ~n61758;
  assign n61760 = ~controllable_hgrant3 & ~n61759;
  assign n61761 = ~n43103 & ~n61760;
  assign n61762 = ~i_hbusreq9 & ~n61761;
  assign n61763 = ~n61750 & ~n61762;
  assign n61764 = ~i_hbusreq4 & ~n61763;
  assign n61765 = ~n61749 & ~n61764;
  assign n61766 = ~controllable_hgrant4 & ~n61765;
  assign n61767 = ~n43094 & ~n61766;
  assign n61768 = ~i_hbusreq5 & ~n61767;
  assign n61769 = ~n61748 & ~n61768;
  assign n61770 = ~controllable_hgrant5 & ~n61769;
  assign n61771 = ~n43083 & ~n61770;
  assign n61772 = controllable_hmaster1 & ~n61771;
  assign n61773 = controllable_hmaster2 & ~n61771;
  assign n61774 = i_hbusreq5 & ~n61622;
  assign n61775 = i_hbusreq4 & ~n61620;
  assign n61776 = i_hbusreq9 & ~n61620;
  assign n61777 = i_hbusreq3 & ~n61612;
  assign n61778 = ~n8389 & ~n18260;
  assign n61779 = ~n43193 & ~n61778;
  assign n61780 = ~i_hbusreq1 & ~n61779;
  assign n61781 = ~n40310 & ~n61780;
  assign n61782 = controllable_hgrant1 & ~n61781;
  assign n61783 = ~n43205 & ~n61782;
  assign n61784 = ~i_hbusreq3 & ~n61783;
  assign n61785 = ~n61777 & ~n61784;
  assign n61786 = ~controllable_hgrant3 & ~n61785;
  assign n61787 = ~n43190 & ~n61786;
  assign n61788 = i_hlock9 & ~n61787;
  assign n61789 = i_hbusreq3 & ~n61616;
  assign n61790 = ~n8389 & ~n18291;
  assign n61791 = ~n43269 & ~n61790;
  assign n61792 = ~i_hbusreq1 & ~n61791;
  assign n61793 = ~n40378 & ~n61792;
  assign n61794 = controllable_hgrant1 & ~n61793;
  assign n61795 = ~n43279 & ~n61794;
  assign n61796 = ~i_hbusreq3 & ~n61795;
  assign n61797 = ~n61789 & ~n61796;
  assign n61798 = ~controllable_hgrant3 & ~n61797;
  assign n61799 = ~n43266 & ~n61798;
  assign n61800 = ~i_hlock9 & ~n61799;
  assign n61801 = ~n61788 & ~n61800;
  assign n61802 = ~i_hbusreq9 & ~n61801;
  assign n61803 = ~n61776 & ~n61802;
  assign n61804 = ~i_hbusreq4 & ~n61803;
  assign n61805 = ~n61775 & ~n61804;
  assign n61806 = ~controllable_hgrant4 & ~n61805;
  assign n61807 = ~n45022 & ~n61806;
  assign n61808 = ~i_hbusreq5 & ~n61807;
  assign n61809 = ~n61774 & ~n61808;
  assign n61810 = ~controllable_hgrant5 & ~n61809;
  assign n61811 = ~n45011 & ~n61810;
  assign n61812 = ~controllable_hmaster2 & ~n61811;
  assign n61813 = ~n61773 & ~n61812;
  assign n61814 = ~controllable_hmaster1 & ~n61813;
  assign n61815 = ~n61772 & ~n61814;
  assign n61816 = ~i_hbusreq6 & ~n61815;
  assign n61817 = ~n61747 & ~n61816;
  assign n61818 = ~controllable_hgrant6 & ~n61817;
  assign n61819 = ~n45003 & ~n61818;
  assign n61820 = controllable_hmaster0 & ~n61819;
  assign n61821 = i_hbusreq6 & ~n61639;
  assign n61822 = i_hbusreq5 & ~n61633;
  assign n61823 = i_hbusreq4 & ~n61614;
  assign n61824 = i_hbusreq9 & ~n61614;
  assign n61825 = ~i_hbusreq9 & ~n61787;
  assign n61826 = ~n61824 & ~n61825;
  assign n61827 = ~i_hbusreq4 & ~n61826;
  assign n61828 = ~n61823 & ~n61827;
  assign n61829 = ~controllable_hgrant4 & ~n61828;
  assign n61830 = ~n43181 & ~n61829;
  assign n61831 = ~i_hbusreq5 & ~n61830;
  assign n61832 = ~n61822 & ~n61831;
  assign n61833 = ~controllable_hgrant5 & ~n61832;
  assign n61834 = ~n43170 & ~n61833;
  assign n61835 = ~controllable_hmaster2 & ~n61834;
  assign n61836 = ~n61773 & ~n61835;
  assign n61837 = ~controllable_hmaster1 & ~n61836;
  assign n61838 = ~n61772 & ~n61837;
  assign n61839 = ~i_hbusreq6 & ~n61838;
  assign n61840 = ~n61821 & ~n61839;
  assign n61841 = ~controllable_hgrant6 & ~n61840;
  assign n61842 = ~n43162 & ~n61841;
  assign n61843 = ~controllable_hmaster0 & ~n61842;
  assign n61844 = ~n61820 & ~n61843;
  assign n61845 = i_hlock8 & ~n61844;
  assign n61846 = i_hbusreq6 & ~n61652;
  assign n61847 = i_hbusreq5 & ~n61646;
  assign n61848 = i_hbusreq4 & ~n61618;
  assign n61849 = i_hbusreq9 & ~n61618;
  assign n61850 = ~i_hbusreq9 & ~n61799;
  assign n61851 = ~n61849 & ~n61850;
  assign n61852 = ~i_hbusreq4 & ~n61851;
  assign n61853 = ~n61848 & ~n61852;
  assign n61854 = ~controllable_hgrant4 & ~n61853;
  assign n61855 = ~n43257 & ~n61854;
  assign n61856 = ~i_hbusreq5 & ~n61855;
  assign n61857 = ~n61847 & ~n61856;
  assign n61858 = ~controllable_hgrant5 & ~n61857;
  assign n61859 = ~n43246 & ~n61858;
  assign n61860 = ~controllable_hmaster2 & ~n61859;
  assign n61861 = ~n61773 & ~n61860;
  assign n61862 = ~controllable_hmaster1 & ~n61861;
  assign n61863 = ~n61772 & ~n61862;
  assign n61864 = ~i_hbusreq6 & ~n61863;
  assign n61865 = ~n61846 & ~n61864;
  assign n61866 = ~controllable_hgrant6 & ~n61865;
  assign n61867 = ~n43238 & ~n61866;
  assign n61868 = ~controllable_hmaster0 & ~n61867;
  assign n61869 = ~n61820 & ~n61868;
  assign n61870 = ~i_hlock8 & ~n61869;
  assign n61871 = ~n61845 & ~n61870;
  assign n61872 = ~i_hbusreq8 & ~n61871;
  assign n61873 = ~n61746 & ~n61872;
  assign n61874 = controllable_hmaster3 & ~n61873;
  assign n61875 = i_hbusreq8 & ~n61727;
  assign n61876 = i_hbusreq6 & ~n61661;
  assign n61877 = n8217 & ~n10893;
  assign n61878 = ~n8217 & ~n24512;
  assign n61879 = ~n61877 & ~n61878;
  assign n61880 = ~i_hbusreq6 & ~n61879;
  assign n61881 = ~n61876 & ~n61880;
  assign n61882 = controllable_hgrant6 & ~n61881;
  assign n61883 = i_hbusreq6 & ~n61684;
  assign n61884 = controllable_hmaster2 & ~n61834;
  assign n61885 = i_hbusreq5 & ~n61670;
  assign n61886 = i_hbusreq4 & ~n61668;
  assign n61887 = i_hbusreq9 & ~n61668;
  assign n61888 = i_hbusreq3 & ~n61666;
  assign n61889 = i_hlock3 & ~n61783;
  assign n61890 = ~i_hlock3 & ~n61795;
  assign n61891 = ~n61889 & ~n61890;
  assign n61892 = ~i_hbusreq3 & ~n61891;
  assign n61893 = ~n61888 & ~n61892;
  assign n61894 = ~controllable_hgrant3 & ~n61893;
  assign n61895 = ~n43352 & ~n61894;
  assign n61896 = ~i_hbusreq9 & ~n61895;
  assign n61897 = ~n61887 & ~n61896;
  assign n61898 = ~i_hbusreq4 & ~n61897;
  assign n61899 = ~n61886 & ~n61898;
  assign n61900 = ~controllable_hgrant4 & ~n61899;
  assign n61901 = ~n43337 & ~n61900;
  assign n61902 = ~i_hbusreq5 & ~n61901;
  assign n61903 = ~n61885 & ~n61902;
  assign n61904 = ~controllable_hgrant5 & ~n61903;
  assign n61905 = ~n43326 & ~n61904;
  assign n61906 = ~controllable_hmaster2 & ~n61905;
  assign n61907 = ~n61884 & ~n61906;
  assign n61908 = controllable_hmaster1 & ~n61907;
  assign n61909 = i_hbusreq5 & ~n61678;
  assign n61910 = i_hlock5 & ~n61830;
  assign n61911 = ~i_hlock5 & ~n61855;
  assign n61912 = ~n61910 & ~n61911;
  assign n61913 = ~i_hbusreq5 & ~n61912;
  assign n61914 = ~n61909 & ~n61913;
  assign n61915 = ~controllable_hgrant5 & ~n61914;
  assign n61916 = ~n43386 & ~n61915;
  assign n61917 = controllable_hmaster2 & ~n61916;
  assign n61918 = ~n48496 & ~n61917;
  assign n61919 = ~controllable_hmaster1 & ~n61918;
  assign n61920 = ~n61908 & ~n61919;
  assign n61921 = ~i_hbusreq6 & ~n61920;
  assign n61922 = ~n61883 & ~n61921;
  assign n61923 = ~controllable_hgrant6 & ~n61922;
  assign n61924 = ~n61882 & ~n61923;
  assign n61925 = controllable_hmaster0 & ~n61924;
  assign n61926 = i_hbusreq6 & ~n61723;
  assign n61927 = i_hbusreq5 & ~n61692;
  assign n61928 = i_hbusreq4 & ~n61690;
  assign n61929 = i_hbusreq9 & ~n61690;
  assign n61930 = i_hbusreq3 & ~n61688;
  assign n61931 = ~n8389 & ~n18402;
  assign n61932 = ~n43523 & ~n61931;
  assign n61933 = ~i_hbusreq1 & ~n61932;
  assign n61934 = ~n48558 & ~n61933;
  assign n61935 = controllable_hgrant1 & ~n61934;
  assign n61936 = ~n43564 & ~n61935;
  assign n61937 = ~i_hbusreq3 & ~n61936;
  assign n61938 = ~n61930 & ~n61937;
  assign n61939 = ~controllable_hgrant3 & ~n61938;
  assign n61940 = ~n43520 & ~n61939;
  assign n61941 = ~i_hbusreq9 & ~n61940;
  assign n61942 = ~n61929 & ~n61941;
  assign n61943 = ~i_hbusreq4 & ~n61942;
  assign n61944 = ~n61928 & ~n61943;
  assign n61945 = ~controllable_hgrant4 & ~n61944;
  assign n61946 = ~n43511 & ~n61945;
  assign n61947 = ~i_hbusreq5 & ~n61946;
  assign n61948 = ~n61927 & ~n61947;
  assign n61949 = ~controllable_hgrant5 & ~n61948;
  assign n61950 = ~n43500 & ~n61949;
  assign n61951 = ~controllable_hmaster2 & ~n61950;
  assign n61952 = ~n61884 & ~n61951;
  assign n61953 = controllable_hmaster1 & ~n61952;
  assign n61954 = i_hbusreq5 & ~n61702;
  assign n61955 = i_hbusreq4 & ~n61700;
  assign n61956 = i_hlock4 & ~n61826;
  assign n61957 = ~i_hlock4 & ~n61851;
  assign n61958 = ~n61956 & ~n61957;
  assign n61959 = ~i_hbusreq4 & ~n61958;
  assign n61960 = ~n61955 & ~n61959;
  assign n61961 = ~controllable_hgrant4 & ~n61960;
  assign n61962 = ~n43609 & ~n61961;
  assign n61963 = ~i_hbusreq5 & ~n61962;
  assign n61964 = ~n61954 & ~n61963;
  assign n61965 = ~controllable_hgrant5 & ~n61964;
  assign n61966 = ~n43589 & ~n61965;
  assign n61967 = controllable_hmaster2 & ~n61966;
  assign n61968 = i_hbusreq5 & ~n61710;
  assign n61969 = i_hbusreq4 & ~n61708;
  assign n61970 = i_hbusreq9 & ~n61708;
  assign n61971 = i_hbusreq3 & ~n61706;
  assign n61972 = ~n8389 & ~n18469;
  assign n61973 = ~n43652 & ~n61972;
  assign n61974 = ~i_hbusreq1 & ~n61973;
  assign n61975 = ~n48677 & ~n61974;
  assign n61976 = controllable_hgrant1 & ~n61975;
  assign n61977 = ~n43675 & ~n61976;
  assign n61978 = ~i_hbusreq3 & ~n61977;
  assign n61979 = ~n61971 & ~n61978;
  assign n61980 = ~controllable_hgrant3 & ~n61979;
  assign n61981 = ~n43649 & ~n61980;
  assign n61982 = ~i_hbusreq9 & ~n61981;
  assign n61983 = ~n61970 & ~n61982;
  assign n61984 = ~i_hbusreq4 & ~n61983;
  assign n61985 = ~n61969 & ~n61984;
  assign n61986 = ~controllable_hgrant4 & ~n61985;
  assign n61987 = ~n43640 & ~n61986;
  assign n61988 = ~i_hbusreq5 & ~n61987;
  assign n61989 = ~n61968 & ~n61988;
  assign n61990 = ~controllable_hgrant5 & ~n61989;
  assign n61991 = ~n43629 & ~n61990;
  assign n61992 = ~controllable_hmaster2 & ~n61991;
  assign n61993 = ~n61967 & ~n61992;
  assign n61994 = ~controllable_hmaster1 & ~n61993;
  assign n61995 = ~n61953 & ~n61994;
  assign n61996 = i_hlock6 & ~n61995;
  assign n61997 = controllable_hmaster2 & ~n61859;
  assign n61998 = ~n61951 & ~n61997;
  assign n61999 = controllable_hmaster1 & ~n61998;
  assign n62000 = ~n61994 & ~n61999;
  assign n62001 = ~i_hlock6 & ~n62000;
  assign n62002 = ~n61996 & ~n62001;
  assign n62003 = ~i_hbusreq6 & ~n62002;
  assign n62004 = ~n61926 & ~n62003;
  assign n62005 = ~controllable_hgrant6 & ~n62004;
  assign n62006 = ~n43492 & ~n62005;
  assign n62007 = ~controllable_hmaster0 & ~n62006;
  assign n62008 = ~n61925 & ~n62007;
  assign n62009 = ~i_hbusreq8 & ~n62008;
  assign n62010 = ~n61875 & ~n62009;
  assign n62011 = ~controllable_hmaster3 & ~n62010;
  assign n62012 = ~n61874 & ~n62011;
  assign n62013 = i_hlock7 & ~n62012;
  assign n62014 = i_hbusreq8 & ~n61740;
  assign n62015 = i_hbusreq6 & ~n61732;
  assign n62016 = n8217 & ~n10903;
  assign n62017 = ~n8217 & ~n24526;
  assign n62018 = ~n62016 & ~n62017;
  assign n62019 = ~i_hbusreq6 & ~n62018;
  assign n62020 = ~n62015 & ~n62019;
  assign n62021 = controllable_hgrant6 & ~n62020;
  assign n62022 = i_hbusreq6 & ~n61736;
  assign n62023 = ~n61906 & ~n61997;
  assign n62024 = controllable_hmaster1 & ~n62023;
  assign n62025 = ~n61919 & ~n62024;
  assign n62026 = ~i_hbusreq6 & ~n62025;
  assign n62027 = ~n62022 & ~n62026;
  assign n62028 = ~controllable_hgrant6 & ~n62027;
  assign n62029 = ~n62021 & ~n62028;
  assign n62030 = controllable_hmaster0 & ~n62029;
  assign n62031 = ~n62007 & ~n62030;
  assign n62032 = ~i_hbusreq8 & ~n62031;
  assign n62033 = ~n62014 & ~n62032;
  assign n62034 = ~controllable_hmaster3 & ~n62033;
  assign n62035 = ~n61874 & ~n62034;
  assign n62036 = ~i_hlock7 & ~n62035;
  assign n62037 = ~n62013 & ~n62036;
  assign n62038 = ~i_hbusreq7 & ~n62037;
  assign n62039 = ~n61745 & ~n62038;
  assign n62040 = ~n7924 & ~n62039;
  assign n62041 = ~n43768 & ~n48793;
  assign n62042 = ~controllable_hgrant3 & ~n62041;
  assign n62043 = ~n43754 & ~n62042;
  assign n62044 = ~controllable_hgrant4 & ~n62043;
  assign n62045 = ~n43750 & ~n62044;
  assign n62046 = ~controllable_hgrant5 & ~n62045;
  assign n62047 = ~n43746 & ~n62046;
  assign n62048 = controllable_hmaster1 & ~n62047;
  assign n62049 = controllable_hmaster2 & ~n62047;
  assign n62050 = ~n43853 & ~n46046;
  assign n62051 = ~controllable_hgrant3 & ~n62050;
  assign n62052 = ~n43842 & ~n62051;
  assign n62053 = i_hlock9 & ~n62052;
  assign n62054 = ~n43886 & ~n46085;
  assign n62055 = ~controllable_hgrant3 & ~n62054;
  assign n62056 = ~n43881 & ~n62055;
  assign n62057 = ~i_hlock9 & ~n62056;
  assign n62058 = ~n62053 & ~n62057;
  assign n62059 = ~controllable_hgrant4 & ~n62058;
  assign n62060 = ~n45104 & ~n62059;
  assign n62061 = ~controllable_hgrant5 & ~n62060;
  assign n62062 = ~n45100 & ~n62061;
  assign n62063 = ~controllable_hmaster2 & ~n62062;
  assign n62064 = ~n62049 & ~n62063;
  assign n62065 = ~controllable_hmaster1 & ~n62064;
  assign n62066 = ~n62048 & ~n62065;
  assign n62067 = ~controllable_hgrant6 & ~n62066;
  assign n62068 = ~n45097 & ~n62067;
  assign n62069 = controllable_hmaster0 & ~n62068;
  assign n62070 = ~controllable_hgrant4 & ~n62052;
  assign n62071 = ~n43839 & ~n62070;
  assign n62072 = ~controllable_hgrant5 & ~n62071;
  assign n62073 = ~n43836 & ~n62072;
  assign n62074 = ~controllable_hmaster2 & ~n62073;
  assign n62075 = ~n62049 & ~n62074;
  assign n62076 = ~controllable_hmaster1 & ~n62075;
  assign n62077 = ~n62048 & ~n62076;
  assign n62078 = ~controllable_hgrant6 & ~n62077;
  assign n62079 = ~n43833 & ~n62078;
  assign n62080 = ~controllable_hmaster0 & ~n62079;
  assign n62081 = ~n62069 & ~n62080;
  assign n62082 = i_hlock8 & ~n62081;
  assign n62083 = ~controllable_hgrant4 & ~n62056;
  assign n62084 = ~n43878 & ~n62083;
  assign n62085 = ~controllable_hgrant5 & ~n62084;
  assign n62086 = ~n43875 & ~n62085;
  assign n62087 = ~controllable_hmaster2 & ~n62086;
  assign n62088 = ~n62049 & ~n62087;
  assign n62089 = ~controllable_hmaster1 & ~n62088;
  assign n62090 = ~n62048 & ~n62089;
  assign n62091 = ~controllable_hgrant6 & ~n62090;
  assign n62092 = ~n43872 & ~n62091;
  assign n62093 = ~controllable_hmaster0 & ~n62092;
  assign n62094 = ~n62069 & ~n62093;
  assign n62095 = ~i_hlock8 & ~n62094;
  assign n62096 = ~n62082 & ~n62095;
  assign n62097 = controllable_hmaster3 & ~n62096;
  assign n62098 = ~n8217 & ~n24556;
  assign n62099 = ~n43905 & ~n62098;
  assign n62100 = controllable_hgrant6 & ~n62099;
  assign n62101 = controllable_hmaster2 & ~n62073;
  assign n62102 = i_hlock3 & ~n62050;
  assign n62103 = ~i_hlock3 & ~n62054;
  assign n62104 = ~n62102 & ~n62103;
  assign n62105 = ~controllable_hgrant3 & ~n62104;
  assign n62106 = ~n43927 & ~n62105;
  assign n62107 = ~controllable_hgrant4 & ~n62106;
  assign n62108 = ~n43917 & ~n62107;
  assign n62109 = ~controllable_hgrant5 & ~n62108;
  assign n62110 = ~n43913 & ~n62109;
  assign n62111 = ~controllable_hmaster2 & ~n62110;
  assign n62112 = ~n62101 & ~n62111;
  assign n62113 = controllable_hmaster1 & ~n62112;
  assign n62114 = i_hlock5 & ~n62071;
  assign n62115 = ~i_hlock5 & ~n62084;
  assign n62116 = ~n62114 & ~n62115;
  assign n62117 = ~controllable_hgrant5 & ~n62116;
  assign n62118 = ~n43949 & ~n62117;
  assign n62119 = controllable_hmaster2 & ~n62118;
  assign n62120 = ~n8378 & ~n24550;
  assign n62121 = ~n43956 & ~n62120;
  assign n62122 = controllable_hgrant5 & ~n62121;
  assign n62123 = ~n8426 & ~n24548;
  assign n62124 = ~n43960 & ~n62123;
  assign n62125 = controllable_hgrant4 & ~n62124;
  assign n62126 = ~n8365 & ~n24546;
  assign n62127 = ~n43964 & ~n62126;
  assign n62128 = controllable_hgrant3 & ~n62127;
  assign n62129 = i_hlock1 & ~n43801;
  assign n62130 = ~i_hlock1 & ~n43813;
  assign n62131 = ~n62129 & ~n62130;
  assign n62132 = ~controllable_hgrant1 & ~n62131;
  assign n62133 = ~n48917 & ~n62132;
  assign n62134 = ~controllable_hgrant3 & ~n62133;
  assign n62135 = ~n62128 & ~n62134;
  assign n62136 = ~controllable_hgrant4 & ~n62135;
  assign n62137 = ~n62125 & ~n62136;
  assign n62138 = ~controllable_hgrant5 & ~n62137;
  assign n62139 = ~n62122 & ~n62138;
  assign n62140 = ~controllable_hmaster2 & ~n62139;
  assign n62141 = ~n62119 & ~n62140;
  assign n62142 = ~controllable_hmaster1 & ~n62141;
  assign n62143 = ~n62113 & ~n62142;
  assign n62144 = ~controllable_hgrant6 & ~n62143;
  assign n62145 = ~n62100 & ~n62144;
  assign n62146 = controllable_hmaster0 & ~n62145;
  assign n62147 = ~n44043 & ~n48967;
  assign n62148 = ~controllable_hgrant3 & ~n62147;
  assign n62149 = ~n44029 & ~n62148;
  assign n62150 = ~controllable_hgrant4 & ~n62149;
  assign n62151 = ~n44025 & ~n62150;
  assign n62152 = ~controllable_hgrant5 & ~n62151;
  assign n62153 = ~n44021 & ~n62152;
  assign n62154 = ~controllable_hmaster2 & ~n62153;
  assign n62155 = ~n62101 & ~n62154;
  assign n62156 = controllable_hmaster1 & ~n62155;
  assign n62157 = i_hlock4 & ~n62052;
  assign n62158 = ~i_hlock4 & ~n62056;
  assign n62159 = ~n62157 & ~n62158;
  assign n62160 = ~controllable_hgrant4 & ~n62159;
  assign n62161 = ~n44067 & ~n62160;
  assign n62162 = ~controllable_hgrant5 & ~n62161;
  assign n62163 = ~n44057 & ~n62162;
  assign n62164 = controllable_hmaster2 & ~n62163;
  assign n62165 = ~n44093 & ~n49049;
  assign n62166 = ~controllable_hgrant3 & ~n62165;
  assign n62167 = ~n44087 & ~n62166;
  assign n62168 = ~controllable_hgrant4 & ~n62167;
  assign n62169 = ~n44083 & ~n62168;
  assign n62170 = ~controllable_hgrant5 & ~n62169;
  assign n62171 = ~n44079 & ~n62170;
  assign n62172 = ~controllable_hmaster2 & ~n62171;
  assign n62173 = ~n62164 & ~n62172;
  assign n62174 = ~controllable_hmaster1 & ~n62173;
  assign n62175 = ~n62156 & ~n62174;
  assign n62176 = i_hlock6 & ~n62175;
  assign n62177 = controllable_hmaster2 & ~n62086;
  assign n62178 = ~n62154 & ~n62177;
  assign n62179 = controllable_hmaster1 & ~n62178;
  assign n62180 = ~n62174 & ~n62179;
  assign n62181 = ~i_hlock6 & ~n62180;
  assign n62182 = ~n62176 & ~n62181;
  assign n62183 = ~controllable_hgrant6 & ~n62182;
  assign n62184 = ~n44017 & ~n62183;
  assign n62185 = ~controllable_hmaster0 & ~n62184;
  assign n62186 = ~n62146 & ~n62185;
  assign n62187 = ~controllable_hmaster3 & ~n62186;
  assign n62188 = ~n62097 & ~n62187;
  assign n62189 = i_hlock7 & ~n62188;
  assign n62190 = ~n8217 & ~n24564;
  assign n62191 = ~n44119 & ~n62190;
  assign n62192 = controllable_hgrant6 & ~n62191;
  assign n62193 = ~n62111 & ~n62177;
  assign n62194 = controllable_hmaster1 & ~n62193;
  assign n62195 = ~n62142 & ~n62194;
  assign n62196 = ~controllable_hgrant6 & ~n62195;
  assign n62197 = ~n62192 & ~n62196;
  assign n62198 = controllable_hmaster0 & ~n62197;
  assign n62199 = ~n62185 & ~n62198;
  assign n62200 = ~controllable_hmaster3 & ~n62199;
  assign n62201 = ~n62097 & ~n62200;
  assign n62202 = ~i_hlock7 & ~n62201;
  assign n62203 = ~n62189 & ~n62202;
  assign n62204 = i_hbusreq7 & ~n62203;
  assign n62205 = i_hbusreq8 & ~n62096;
  assign n62206 = i_hbusreq6 & ~n62066;
  assign n62207 = i_hbusreq5 & ~n62045;
  assign n62208 = i_hbusreq4 & ~n62043;
  assign n62209 = i_hbusreq9 & ~n62043;
  assign n62210 = i_hbusreq3 & ~n62041;
  assign n62211 = n8389 & ~n13990;
  assign n62212 = ~n8389 & ~n18737;
  assign n62213 = ~n62211 & ~n62212;
  assign n62214 = i_hlock1 & ~n62213;
  assign n62215 = ~n8389 & ~n18755;
  assign n62216 = ~n62211 & ~n62215;
  assign n62217 = ~i_hlock1 & ~n62216;
  assign n62218 = ~n62214 & ~n62217;
  assign n62219 = ~i_hbusreq1 & ~n62218;
  assign n62220 = ~n49147 & ~n62219;
  assign n62221 = controllable_hgrant1 & ~n62220;
  assign n62222 = ~n44207 & ~n62221;
  assign n62223 = ~i_hbusreq3 & ~n62222;
  assign n62224 = ~n62210 & ~n62223;
  assign n62225 = ~controllable_hgrant3 & ~n62224;
  assign n62226 = ~n44170 & ~n62225;
  assign n62227 = ~i_hbusreq9 & ~n62226;
  assign n62228 = ~n62209 & ~n62227;
  assign n62229 = ~i_hbusreq4 & ~n62228;
  assign n62230 = ~n62208 & ~n62229;
  assign n62231 = ~controllable_hgrant4 & ~n62230;
  assign n62232 = ~n44161 & ~n62231;
  assign n62233 = ~i_hbusreq5 & ~n62232;
  assign n62234 = ~n62207 & ~n62233;
  assign n62235 = ~controllable_hgrant5 & ~n62234;
  assign n62236 = ~n44150 & ~n62235;
  assign n62237 = controllable_hmaster1 & ~n62236;
  assign n62238 = controllable_hmaster2 & ~n62236;
  assign n62239 = i_hbusreq5 & ~n62060;
  assign n62240 = i_hbusreq4 & ~n62058;
  assign n62241 = i_hbusreq9 & ~n62058;
  assign n62242 = i_hbusreq3 & ~n62050;
  assign n62243 = n8389 & ~n14024;
  assign n62244 = ~n8389 & ~n18803;
  assign n62245 = ~n62243 & ~n62244;
  assign n62246 = i_hlock1 & ~n62245;
  assign n62247 = ~n8389 & ~n18817;
  assign n62248 = ~n62243 & ~n62247;
  assign n62249 = ~i_hlock1 & ~n62248;
  assign n62250 = ~n62246 & ~n62249;
  assign n62251 = ~i_hbusreq1 & ~n62250;
  assign n62252 = ~n46676 & ~n62251;
  assign n62253 = controllable_hgrant1 & ~n62252;
  assign n62254 = ~n44415 & ~n62253;
  assign n62255 = ~i_hbusreq3 & ~n62254;
  assign n62256 = ~n62242 & ~n62255;
  assign n62257 = ~controllable_hgrant3 & ~n62256;
  assign n62258 = ~n44396 & ~n62257;
  assign n62259 = i_hlock9 & ~n62258;
  assign n62260 = i_hbusreq3 & ~n62054;
  assign n62261 = n8389 & ~n14059;
  assign n62262 = ~n8389 & ~n18855;
  assign n62263 = ~n62261 & ~n62262;
  assign n62264 = i_hlock1 & ~n62263;
  assign n62265 = ~n8389 & ~n18867;
  assign n62266 = ~n62261 & ~n62265;
  assign n62267 = ~i_hlock1 & ~n62266;
  assign n62268 = ~n62264 & ~n62267;
  assign n62269 = ~i_hbusreq1 & ~n62268;
  assign n62270 = ~n46740 & ~n62269;
  assign n62271 = controllable_hgrant1 & ~n62270;
  assign n62272 = ~n44489 & ~n62271;
  assign n62273 = ~i_hbusreq3 & ~n62272;
  assign n62274 = ~n62260 & ~n62273;
  assign n62275 = ~controllable_hgrant3 & ~n62274;
  assign n62276 = ~n44476 & ~n62275;
  assign n62277 = ~i_hlock9 & ~n62276;
  assign n62278 = ~n62259 & ~n62277;
  assign n62279 = ~i_hbusreq9 & ~n62278;
  assign n62280 = ~n62241 & ~n62279;
  assign n62281 = ~i_hbusreq4 & ~n62280;
  assign n62282 = ~n62240 & ~n62281;
  assign n62283 = ~controllable_hgrant4 & ~n62282;
  assign n62284 = ~n45193 & ~n62283;
  assign n62285 = ~i_hbusreq5 & ~n62284;
  assign n62286 = ~n62239 & ~n62285;
  assign n62287 = ~controllable_hgrant5 & ~n62286;
  assign n62288 = ~n45182 & ~n62287;
  assign n62289 = ~controllable_hmaster2 & ~n62288;
  assign n62290 = ~n62238 & ~n62289;
  assign n62291 = ~controllable_hmaster1 & ~n62290;
  assign n62292 = ~n62237 & ~n62291;
  assign n62293 = ~i_hbusreq6 & ~n62292;
  assign n62294 = ~n62206 & ~n62293;
  assign n62295 = ~controllable_hgrant6 & ~n62294;
  assign n62296 = ~n45174 & ~n62295;
  assign n62297 = controllable_hmaster0 & ~n62296;
  assign n62298 = i_hbusreq6 & ~n62077;
  assign n62299 = i_hbusreq5 & ~n62071;
  assign n62300 = i_hbusreq4 & ~n62052;
  assign n62301 = i_hbusreq9 & ~n62052;
  assign n62302 = ~i_hbusreq9 & ~n62258;
  assign n62303 = ~n62301 & ~n62302;
  assign n62304 = ~i_hbusreq4 & ~n62303;
  assign n62305 = ~n62300 & ~n62304;
  assign n62306 = ~controllable_hgrant4 & ~n62305;
  assign n62307 = ~n44387 & ~n62306;
  assign n62308 = ~i_hbusreq5 & ~n62307;
  assign n62309 = ~n62299 & ~n62308;
  assign n62310 = ~controllable_hgrant5 & ~n62309;
  assign n62311 = ~n44376 & ~n62310;
  assign n62312 = ~controllable_hmaster2 & ~n62311;
  assign n62313 = ~n62238 & ~n62312;
  assign n62314 = ~controllable_hmaster1 & ~n62313;
  assign n62315 = ~n62237 & ~n62314;
  assign n62316 = ~i_hbusreq6 & ~n62315;
  assign n62317 = ~n62298 & ~n62316;
  assign n62318 = ~controllable_hgrant6 & ~n62317;
  assign n62319 = ~n44368 & ~n62318;
  assign n62320 = ~controllable_hmaster0 & ~n62319;
  assign n62321 = ~n62297 & ~n62320;
  assign n62322 = i_hlock8 & ~n62321;
  assign n62323 = i_hbusreq6 & ~n62090;
  assign n62324 = i_hbusreq5 & ~n62084;
  assign n62325 = i_hbusreq4 & ~n62056;
  assign n62326 = i_hbusreq9 & ~n62056;
  assign n62327 = ~i_hbusreq9 & ~n62276;
  assign n62328 = ~n62326 & ~n62327;
  assign n62329 = ~i_hbusreq4 & ~n62328;
  assign n62330 = ~n62325 & ~n62329;
  assign n62331 = ~controllable_hgrant4 & ~n62330;
  assign n62332 = ~n44467 & ~n62331;
  assign n62333 = ~i_hbusreq5 & ~n62332;
  assign n62334 = ~n62324 & ~n62333;
  assign n62335 = ~controllable_hgrant5 & ~n62334;
  assign n62336 = ~n44456 & ~n62335;
  assign n62337 = ~controllable_hmaster2 & ~n62336;
  assign n62338 = ~n62238 & ~n62337;
  assign n62339 = ~controllable_hmaster1 & ~n62338;
  assign n62340 = ~n62237 & ~n62339;
  assign n62341 = ~i_hbusreq6 & ~n62340;
  assign n62342 = ~n62323 & ~n62341;
  assign n62343 = ~controllable_hgrant6 & ~n62342;
  assign n62344 = ~n44448 & ~n62343;
  assign n62345 = ~controllable_hmaster0 & ~n62344;
  assign n62346 = ~n62297 & ~n62345;
  assign n62347 = ~i_hlock8 & ~n62346;
  assign n62348 = ~n62322 & ~n62347;
  assign n62349 = ~i_hbusreq8 & ~n62348;
  assign n62350 = ~n62205 & ~n62349;
  assign n62351 = controllable_hmaster3 & ~n62350;
  assign n62352 = i_hbusreq8 & ~n62186;
  assign n62353 = i_hbusreq6 & ~n62099;
  assign n62354 = n8217 & ~n16056;
  assign n62355 = ~n8217 & ~n24605;
  assign n62356 = ~n62354 & ~n62355;
  assign n62357 = ~i_hbusreq6 & ~n62356;
  assign n62358 = ~n62353 & ~n62357;
  assign n62359 = controllable_hgrant6 & ~n62358;
  assign n62360 = i_hbusreq6 & ~n62143;
  assign n62361 = controllable_hmaster2 & ~n62311;
  assign n62362 = i_hbusreq5 & ~n62108;
  assign n62363 = i_hbusreq4 & ~n62106;
  assign n62364 = i_hbusreq9 & ~n62106;
  assign n62365 = i_hbusreq3 & ~n62104;
  assign n62366 = i_hlock3 & ~n62254;
  assign n62367 = ~i_hlock3 & ~n62272;
  assign n62368 = ~n62366 & ~n62367;
  assign n62369 = ~i_hbusreq3 & ~n62368;
  assign n62370 = ~n62365 & ~n62369;
  assign n62371 = ~controllable_hgrant3 & ~n62370;
  assign n62372 = ~n44562 & ~n62371;
  assign n62373 = ~i_hbusreq9 & ~n62372;
  assign n62374 = ~n62364 & ~n62373;
  assign n62375 = ~i_hbusreq4 & ~n62374;
  assign n62376 = ~n62363 & ~n62375;
  assign n62377 = ~controllable_hgrant4 & ~n62376;
  assign n62378 = ~n44547 & ~n62377;
  assign n62379 = ~i_hbusreq5 & ~n62378;
  assign n62380 = ~n62362 & ~n62379;
  assign n62381 = ~controllable_hgrant5 & ~n62380;
  assign n62382 = ~n44536 & ~n62381;
  assign n62383 = ~controllable_hmaster2 & ~n62382;
  assign n62384 = ~n62361 & ~n62383;
  assign n62385 = controllable_hmaster1 & ~n62384;
  assign n62386 = i_hbusreq5 & ~n62116;
  assign n62387 = i_hlock5 & ~n62307;
  assign n62388 = ~i_hlock5 & ~n62332;
  assign n62389 = ~n62387 & ~n62388;
  assign n62390 = ~i_hbusreq5 & ~n62389;
  assign n62391 = ~n62386 & ~n62390;
  assign n62392 = ~controllable_hgrant5 & ~n62391;
  assign n62393 = ~n44596 & ~n62392;
  assign n62394 = controllable_hmaster2 & ~n62393;
  assign n62395 = i_hbusreq5 & ~n62121;
  assign n62396 = n8378 & ~n16048;
  assign n62397 = ~n8378 & ~n24597;
  assign n62398 = ~n62396 & ~n62397;
  assign n62399 = ~i_hbusreq5 & ~n62398;
  assign n62400 = ~n62395 & ~n62399;
  assign n62401 = controllable_hgrant5 & ~n62400;
  assign n62402 = i_hbusreq5 & ~n62137;
  assign n62403 = i_hbusreq4 & ~n62124;
  assign n62404 = i_hbusreq9 & ~n62124;
  assign n62405 = n8426 & ~n16042;
  assign n62406 = ~n8426 & ~n24591;
  assign n62407 = ~n62405 & ~n62406;
  assign n62408 = ~i_hbusreq9 & ~n62407;
  assign n62409 = ~n62404 & ~n62408;
  assign n62410 = ~i_hbusreq4 & ~n62409;
  assign n62411 = ~n62403 & ~n62410;
  assign n62412 = controllable_hgrant4 & ~n62411;
  assign n62413 = i_hbusreq4 & ~n62135;
  assign n62414 = i_hbusreq9 & ~n62135;
  assign n62415 = i_hbusreq3 & ~n62127;
  assign n62416 = n8365 & ~n16038;
  assign n62417 = ~n8365 & ~n24587;
  assign n62418 = ~n62416 & ~n62417;
  assign n62419 = ~i_hbusreq3 & ~n62418;
  assign n62420 = ~n62415 & ~n62419;
  assign n62421 = controllable_hgrant3 & ~n62420;
  assign n62422 = i_hbusreq3 & ~n62133;
  assign n62423 = i_hbusreq1 & ~n62131;
  assign n62424 = i_hlock1 & ~n44306;
  assign n62425 = ~i_hlock1 & ~n44332;
  assign n62426 = ~n62424 & ~n62425;
  assign n62427 = ~i_hbusreq1 & ~n62426;
  assign n62428 = ~n62423 & ~n62427;
  assign n62429 = ~controllable_hgrant1 & ~n62428;
  assign n62430 = ~n49636 & ~n62429;
  assign n62431 = ~i_hbusreq3 & ~n62430;
  assign n62432 = ~n62422 & ~n62431;
  assign n62433 = ~controllable_hgrant3 & ~n62432;
  assign n62434 = ~n62421 & ~n62433;
  assign n62435 = ~i_hbusreq9 & ~n62434;
  assign n62436 = ~n62414 & ~n62435;
  assign n62437 = ~i_hbusreq4 & ~n62436;
  assign n62438 = ~n62413 & ~n62437;
  assign n62439 = ~controllable_hgrant4 & ~n62438;
  assign n62440 = ~n62412 & ~n62439;
  assign n62441 = ~i_hbusreq5 & ~n62440;
  assign n62442 = ~n62402 & ~n62441;
  assign n62443 = ~controllable_hgrant5 & ~n62442;
  assign n62444 = ~n62401 & ~n62443;
  assign n62445 = ~controllable_hmaster2 & ~n62444;
  assign n62446 = ~n62394 & ~n62445;
  assign n62447 = ~controllable_hmaster1 & ~n62446;
  assign n62448 = ~n62385 & ~n62447;
  assign n62449 = ~i_hbusreq6 & ~n62448;
  assign n62450 = ~n62360 & ~n62449;
  assign n62451 = ~controllable_hgrant6 & ~n62450;
  assign n62452 = ~n62359 & ~n62451;
  assign n62453 = controllable_hmaster0 & ~n62452;
  assign n62454 = i_hbusreq6 & ~n62182;
  assign n62455 = i_hbusreq5 & ~n62151;
  assign n62456 = i_hbusreq4 & ~n62149;
  assign n62457 = i_hbusreq9 & ~n62149;
  assign n62458 = i_hbusreq3 & ~n62147;
  assign n62459 = n8389 & ~n14184;
  assign n62460 = ~n8389 & ~n19007;
  assign n62461 = ~n62459 & ~n62460;
  assign n62462 = i_hlock1 & ~n62461;
  assign n62463 = ~n8389 & ~n19019;
  assign n62464 = ~n62459 & ~n62463;
  assign n62465 = ~i_hlock1 & ~n62464;
  assign n62466 = ~n62462 & ~n62465;
  assign n62467 = ~i_hbusreq1 & ~n62466;
  assign n62468 = ~n49739 & ~n62467;
  assign n62469 = controllable_hgrant1 & ~n62468;
  assign n62470 = ~n44760 & ~n62469;
  assign n62471 = ~i_hbusreq3 & ~n62470;
  assign n62472 = ~n62458 & ~n62471;
  assign n62473 = ~controllable_hgrant3 & ~n62472;
  assign n62474 = ~n44730 & ~n62473;
  assign n62475 = ~i_hbusreq9 & ~n62474;
  assign n62476 = ~n62457 & ~n62475;
  assign n62477 = ~i_hbusreq4 & ~n62476;
  assign n62478 = ~n62456 & ~n62477;
  assign n62479 = ~controllable_hgrant4 & ~n62478;
  assign n62480 = ~n44721 & ~n62479;
  assign n62481 = ~i_hbusreq5 & ~n62480;
  assign n62482 = ~n62455 & ~n62481;
  assign n62483 = ~controllable_hgrant5 & ~n62482;
  assign n62484 = ~n44710 & ~n62483;
  assign n62485 = ~controllable_hmaster2 & ~n62484;
  assign n62486 = ~n62361 & ~n62485;
  assign n62487 = controllable_hmaster1 & ~n62486;
  assign n62488 = i_hbusreq5 & ~n62161;
  assign n62489 = i_hbusreq4 & ~n62159;
  assign n62490 = i_hlock4 & ~n62303;
  assign n62491 = ~i_hlock4 & ~n62328;
  assign n62492 = ~n62490 & ~n62491;
  assign n62493 = ~i_hbusreq4 & ~n62492;
  assign n62494 = ~n62489 & ~n62493;
  assign n62495 = ~controllable_hgrant4 & ~n62494;
  assign n62496 = ~n44805 & ~n62495;
  assign n62497 = ~i_hbusreq5 & ~n62496;
  assign n62498 = ~n62488 & ~n62497;
  assign n62499 = ~controllable_hgrant5 & ~n62498;
  assign n62500 = ~n44785 & ~n62499;
  assign n62501 = controllable_hmaster2 & ~n62500;
  assign n62502 = i_hbusreq5 & ~n62169;
  assign n62503 = i_hbusreq4 & ~n62167;
  assign n62504 = i_hbusreq9 & ~n62167;
  assign n62505 = i_hbusreq3 & ~n62165;
  assign n62506 = n8389 & ~n14256;
  assign n62507 = ~n8389 & ~n19088;
  assign n62508 = ~n62506 & ~n62507;
  assign n62509 = i_hlock1 & ~n62508;
  assign n62510 = ~n8389 & ~n19108;
  assign n62511 = ~n62506 & ~n62510;
  assign n62512 = ~i_hlock1 & ~n62511;
  assign n62513 = ~n62509 & ~n62512;
  assign n62514 = ~i_hbusreq1 & ~n62513;
  assign n62515 = ~n49888 & ~n62514;
  assign n62516 = controllable_hgrant1 & ~n62515;
  assign n62517 = ~n44875 & ~n62516;
  assign n62518 = ~i_hbusreq3 & ~n62517;
  assign n62519 = ~n62505 & ~n62518;
  assign n62520 = ~controllable_hgrant3 & ~n62519;
  assign n62521 = ~n44845 & ~n62520;
  assign n62522 = ~i_hbusreq9 & ~n62521;
  assign n62523 = ~n62504 & ~n62522;
  assign n62524 = ~i_hbusreq4 & ~n62523;
  assign n62525 = ~n62503 & ~n62524;
  assign n62526 = ~controllable_hgrant4 & ~n62525;
  assign n62527 = ~n44836 & ~n62526;
  assign n62528 = ~i_hbusreq5 & ~n62527;
  assign n62529 = ~n62502 & ~n62528;
  assign n62530 = ~controllable_hgrant5 & ~n62529;
  assign n62531 = ~n44825 & ~n62530;
  assign n62532 = ~controllable_hmaster2 & ~n62531;
  assign n62533 = ~n62501 & ~n62532;
  assign n62534 = ~controllable_hmaster1 & ~n62533;
  assign n62535 = ~n62487 & ~n62534;
  assign n62536 = i_hlock6 & ~n62535;
  assign n62537 = controllable_hmaster2 & ~n62336;
  assign n62538 = ~n62485 & ~n62537;
  assign n62539 = controllable_hmaster1 & ~n62538;
  assign n62540 = ~n62534 & ~n62539;
  assign n62541 = ~i_hlock6 & ~n62540;
  assign n62542 = ~n62536 & ~n62541;
  assign n62543 = ~i_hbusreq6 & ~n62542;
  assign n62544 = ~n62454 & ~n62543;
  assign n62545 = ~controllable_hgrant6 & ~n62544;
  assign n62546 = ~n44702 & ~n62545;
  assign n62547 = ~controllable_hmaster0 & ~n62546;
  assign n62548 = ~n62453 & ~n62547;
  assign n62549 = ~i_hbusreq8 & ~n62548;
  assign n62550 = ~n62352 & ~n62549;
  assign n62551 = ~controllable_hmaster3 & ~n62550;
  assign n62552 = ~n62351 & ~n62551;
  assign n62553 = i_hlock7 & ~n62552;
  assign n62554 = i_hbusreq8 & ~n62199;
  assign n62555 = i_hbusreq6 & ~n62191;
  assign n62556 = n8217 & ~n16069;
  assign n62557 = ~n8217 & ~n24619;
  assign n62558 = ~n62556 & ~n62557;
  assign n62559 = ~i_hbusreq6 & ~n62558;
  assign n62560 = ~n62555 & ~n62559;
  assign n62561 = controllable_hgrant6 & ~n62560;
  assign n62562 = i_hbusreq6 & ~n62195;
  assign n62563 = ~n62383 & ~n62537;
  assign n62564 = controllable_hmaster1 & ~n62563;
  assign n62565 = ~n62447 & ~n62564;
  assign n62566 = ~i_hbusreq6 & ~n62565;
  assign n62567 = ~n62562 & ~n62566;
  assign n62568 = ~controllable_hgrant6 & ~n62567;
  assign n62569 = ~n62561 & ~n62568;
  assign n62570 = controllable_hmaster0 & ~n62569;
  assign n62571 = ~n62547 & ~n62570;
  assign n62572 = ~i_hbusreq8 & ~n62571;
  assign n62573 = ~n62554 & ~n62572;
  assign n62574 = ~controllable_hmaster3 & ~n62573;
  assign n62575 = ~n62351 & ~n62574;
  assign n62576 = ~i_hlock7 & ~n62575;
  assign n62577 = ~n62553 & ~n62576;
  assign n62578 = ~i_hbusreq7 & ~n62577;
  assign n62579 = ~n62204 & ~n62578;
  assign n62580 = n7924 & ~n62579;
  assign n62581 = ~n62040 & ~n62580;
  assign n62582 = ~n8214 & ~n62581;
  assign n62583 = ~n24638 & ~n42912;
  assign n62584 = ~n8217 & ~n62583;
  assign n62585 = ~n42910 & ~n62584;
  assign n62586 = i_hlock6 & ~n62585;
  assign n62587 = ~n24638 & ~n42922;
  assign n62588 = ~n8217 & ~n62587;
  assign n62589 = ~n42920 & ~n62588;
  assign n62590 = ~i_hlock6 & ~n62589;
  assign n62591 = ~n62586 & ~n62590;
  assign n62592 = controllable_hgrant6 & ~n62591;
  assign n62593 = ~n43008 & ~n48207;
  assign n62594 = ~controllable_hmaster1 & ~n62593;
  assign n62595 = ~n42986 & ~n62594;
  assign n62596 = i_hlock6 & ~n62595;
  assign n62597 = ~n43041 & ~n62594;
  assign n62598 = ~i_hlock6 & ~n62597;
  assign n62599 = ~n62596 & ~n62598;
  assign n62600 = ~controllable_hgrant6 & ~n62599;
  assign n62601 = ~n62592 & ~n62600;
  assign n62602 = ~controllable_hmaster0 & ~n62601;
  assign n62603 = ~n42906 & ~n62602;
  assign n62604 = ~controllable_hmaster3 & ~n62603;
  assign n62605 = ~n45331 & ~n62604;
  assign n62606 = i_hlock7 & ~n62605;
  assign n62607 = ~n43061 & ~n62602;
  assign n62608 = ~controllable_hmaster3 & ~n62607;
  assign n62609 = ~n45331 & ~n62608;
  assign n62610 = ~i_hlock7 & ~n62609;
  assign n62611 = ~n62606 & ~n62610;
  assign n62612 = i_hbusreq7 & ~n62611;
  assign n62613 = ~n8217 & ~n33975;
  assign n62614 = ~n48237 & ~n62613;
  assign n62615 = ~i_hbusreq6 & ~n62614;
  assign n62616 = ~n44997 & ~n62615;
  assign n62617 = controllable_hgrant6 & ~n62616;
  assign n62618 = ~n8378 & ~n24681;
  assign n62619 = ~n48245 & ~n62618;
  assign n62620 = ~i_hbusreq5 & ~n62619;
  assign n62621 = ~n43077 & ~n62620;
  assign n62622 = controllable_hgrant5 & ~n62621;
  assign n62623 = ~n8426 & ~n24675;
  assign n62624 = ~n48254 & ~n62623;
  assign n62625 = ~i_hbusreq9 & ~n62624;
  assign n62626 = ~n43086 & ~n62625;
  assign n62627 = ~i_hbusreq4 & ~n62626;
  assign n62628 = ~n43085 & ~n62627;
  assign n62629 = controllable_hgrant4 & ~n62628;
  assign n62630 = ~n8365 & ~n24671;
  assign n62631 = ~n48265 & ~n62630;
  assign n62632 = ~i_hbusreq3 & ~n62631;
  assign n62633 = ~n43097 & ~n62632;
  assign n62634 = controllable_hgrant3 & ~n62633;
  assign n62635 = ~n8389 & ~n24667;
  assign n62636 = ~n48273 & ~n62635;
  assign n62637 = ~i_hbusreq1 & ~n62636;
  assign n62638 = ~n43105 & ~n62637;
  assign n62639 = controllable_hgrant1 & ~n62638;
  assign n62640 = ~n7733 & ~n42722;
  assign n62641 = ~n12640 & ~n40339;
  assign n62642 = i_hlock0 & ~n62641;
  assign n62643 = ~n40324 & ~n62642;
  assign n62644 = ~i_hbusreq0 & ~n62643;
  assign n62645 = ~n40319 & ~n62644;
  assign n62646 = ~i_hbusreq2 & ~n62645;
  assign n62647 = ~n40318 & ~n62646;
  assign n62648 = controllable_hgrant2 & ~n62647;
  assign n62649 = ~n24695 & ~n62648;
  assign n62650 = n7733 & ~n62649;
  assign n62651 = ~n62640 & ~n62650;
  assign n62652 = ~n7928 & ~n62651;
  assign n62653 = ~n42725 & ~n62650;
  assign n62654 = n7928 & ~n62653;
  assign n62655 = ~n62652 & ~n62654;
  assign n62656 = ~i_hbusreq1 & ~n62655;
  assign n62657 = ~n43112 & ~n62656;
  assign n62658 = ~controllable_hgrant1 & ~n62657;
  assign n62659 = ~n62639 & ~n62658;
  assign n62660 = ~i_hbusreq3 & ~n62659;
  assign n62661 = ~n43104 & ~n62660;
  assign n62662 = ~controllable_hgrant3 & ~n62661;
  assign n62663 = ~n62634 & ~n62662;
  assign n62664 = ~i_hbusreq9 & ~n62663;
  assign n62665 = ~n43096 & ~n62664;
  assign n62666 = ~i_hbusreq4 & ~n62665;
  assign n62667 = ~n43095 & ~n62666;
  assign n62668 = ~controllable_hgrant4 & ~n62667;
  assign n62669 = ~n62629 & ~n62668;
  assign n62670 = ~i_hbusreq5 & ~n62669;
  assign n62671 = ~n43084 & ~n62670;
  assign n62672 = ~controllable_hgrant5 & ~n62671;
  assign n62673 = ~n62622 & ~n62672;
  assign n62674 = controllable_hmaster1 & ~n62673;
  assign n62675 = controllable_hmaster2 & ~n62673;
  assign n62676 = ~n8378 & ~n33967;
  assign n62677 = ~n40277 & ~n62676;
  assign n62678 = ~i_hbusreq5 & ~n62677;
  assign n62679 = ~n45005 & ~n62678;
  assign n62680 = controllable_hgrant5 & ~n62679;
  assign n62681 = ~n8426 & ~n24750;
  assign n62682 = ~n40286 & ~n62681;
  assign n62683 = i_hlock9 & ~n62682;
  assign n62684 = ~n8426 & ~n24780;
  assign n62685 = ~n40290 & ~n62684;
  assign n62686 = ~i_hlock9 & ~n62685;
  assign n62687 = ~n62683 & ~n62686;
  assign n62688 = ~i_hbusreq9 & ~n62687;
  assign n62689 = ~n45014 & ~n62688;
  assign n62690 = ~i_hbusreq4 & ~n62689;
  assign n62691 = ~n45013 & ~n62690;
  assign n62692 = controllable_hgrant4 & ~n62691;
  assign n62693 = ~n8365 & ~n24746;
  assign n62694 = ~n40303 & ~n62693;
  assign n62695 = ~i_hbusreq3 & ~n62694;
  assign n62696 = ~n43184 & ~n62695;
  assign n62697 = controllable_hgrant3 & ~n62696;
  assign n62698 = ~n8389 & ~n24742;
  assign n62699 = ~n40311 & ~n62698;
  assign n62700 = ~i_hbusreq1 & ~n62699;
  assign n62701 = ~n43192 & ~n62700;
  assign n62702 = controllable_hgrant1 & ~n62701;
  assign n62703 = ~n24664 & ~n62648;
  assign n62704 = n7733 & ~n62703;
  assign n62705 = ~n55937 & ~n62704;
  assign n62706 = n7928 & ~n62705;
  assign n62707 = ~n8265 & ~n62706;
  assign n62708 = ~i_hbusreq1 & ~n62707;
  assign n62709 = ~n43199 & ~n62708;
  assign n62710 = ~controllable_hgrant1 & ~n62709;
  assign n62711 = ~n62702 & ~n62710;
  assign n62712 = ~i_hbusreq3 & ~n62711;
  assign n62713 = ~n43191 & ~n62712;
  assign n62714 = ~controllable_hgrant3 & ~n62713;
  assign n62715 = ~n62697 & ~n62714;
  assign n62716 = i_hlock9 & ~n62715;
  assign n62717 = ~n8365 & ~n24776;
  assign n62718 = ~n40371 & ~n62717;
  assign n62719 = ~i_hbusreq3 & ~n62718;
  assign n62720 = ~n43260 & ~n62719;
  assign n62721 = controllable_hgrant3 & ~n62720;
  assign n62722 = ~n8389 & ~n24772;
  assign n62723 = ~n40379 & ~n62722;
  assign n62724 = ~i_hbusreq1 & ~n62723;
  assign n62725 = ~n43268 & ~n62724;
  assign n62726 = controllable_hgrant1 & ~n62725;
  assign n62727 = ~n8297 & ~n62706;
  assign n62728 = ~i_hbusreq1 & ~n62727;
  assign n62729 = ~n43275 & ~n62728;
  assign n62730 = ~controllable_hgrant1 & ~n62729;
  assign n62731 = ~n62726 & ~n62730;
  assign n62732 = ~i_hbusreq3 & ~n62731;
  assign n62733 = ~n43267 & ~n62732;
  assign n62734 = ~controllable_hgrant3 & ~n62733;
  assign n62735 = ~n62721 & ~n62734;
  assign n62736 = ~i_hlock9 & ~n62735;
  assign n62737 = ~n62716 & ~n62736;
  assign n62738 = ~i_hbusreq9 & ~n62737;
  assign n62739 = ~n45024 & ~n62738;
  assign n62740 = ~i_hbusreq4 & ~n62739;
  assign n62741 = ~n45023 & ~n62740;
  assign n62742 = ~controllable_hgrant4 & ~n62741;
  assign n62743 = ~n62692 & ~n62742;
  assign n62744 = ~i_hbusreq5 & ~n62743;
  assign n62745 = ~n45012 & ~n62744;
  assign n62746 = ~controllable_hgrant5 & ~n62745;
  assign n62747 = ~n62680 & ~n62746;
  assign n62748 = ~controllable_hmaster2 & ~n62747;
  assign n62749 = ~n62675 & ~n62748;
  assign n62750 = ~controllable_hmaster1 & ~n62749;
  assign n62751 = ~n62674 & ~n62750;
  assign n62752 = ~i_hbusreq6 & ~n62751;
  assign n62753 = ~n45004 & ~n62752;
  assign n62754 = ~controllable_hgrant6 & ~n62753;
  assign n62755 = ~n62617 & ~n62754;
  assign n62756 = controllable_hmaster0 & ~n62755;
  assign n62757 = ~n8217 & ~n24764;
  assign n62758 = ~n48311 & ~n62757;
  assign n62759 = ~i_hbusreq6 & ~n62758;
  assign n62760 = ~n43156 & ~n62759;
  assign n62761 = controllable_hgrant6 & ~n62760;
  assign n62762 = ~n8378 & ~n24756;
  assign n62763 = ~n40482 & ~n62762;
  assign n62764 = ~i_hbusreq5 & ~n62763;
  assign n62765 = ~n43164 & ~n62764;
  assign n62766 = controllable_hgrant5 & ~n62765;
  assign n62767 = ~i_hbusreq9 & ~n62682;
  assign n62768 = ~n43173 & ~n62767;
  assign n62769 = ~i_hbusreq4 & ~n62768;
  assign n62770 = ~n43172 & ~n62769;
  assign n62771 = controllable_hgrant4 & ~n62770;
  assign n62772 = ~i_hbusreq9 & ~n62715;
  assign n62773 = ~n43183 & ~n62772;
  assign n62774 = ~i_hbusreq4 & ~n62773;
  assign n62775 = ~n43182 & ~n62774;
  assign n62776 = ~controllable_hgrant4 & ~n62775;
  assign n62777 = ~n62771 & ~n62776;
  assign n62778 = ~i_hbusreq5 & ~n62777;
  assign n62779 = ~n43171 & ~n62778;
  assign n62780 = ~controllable_hgrant5 & ~n62779;
  assign n62781 = ~n62766 & ~n62780;
  assign n62782 = ~controllable_hmaster2 & ~n62781;
  assign n62783 = ~n62675 & ~n62782;
  assign n62784 = ~controllable_hmaster1 & ~n62783;
  assign n62785 = ~n62674 & ~n62784;
  assign n62786 = ~i_hbusreq6 & ~n62785;
  assign n62787 = ~n43163 & ~n62786;
  assign n62788 = ~controllable_hgrant6 & ~n62787;
  assign n62789 = ~n62761 & ~n62788;
  assign n62790 = ~controllable_hmaster0 & ~n62789;
  assign n62791 = ~n62756 & ~n62790;
  assign n62792 = i_hlock8 & ~n62791;
  assign n62793 = ~n8217 & ~n24794;
  assign n62794 = ~n48328 & ~n62793;
  assign n62795 = ~i_hbusreq6 & ~n62794;
  assign n62796 = ~n43232 & ~n62795;
  assign n62797 = controllable_hgrant6 & ~n62796;
  assign n62798 = ~n8378 & ~n24786;
  assign n62799 = ~n40528 & ~n62798;
  assign n62800 = ~i_hbusreq5 & ~n62799;
  assign n62801 = ~n43240 & ~n62800;
  assign n62802 = controllable_hgrant5 & ~n62801;
  assign n62803 = ~i_hbusreq9 & ~n62685;
  assign n62804 = ~n43249 & ~n62803;
  assign n62805 = ~i_hbusreq4 & ~n62804;
  assign n62806 = ~n43248 & ~n62805;
  assign n62807 = controllable_hgrant4 & ~n62806;
  assign n62808 = ~i_hbusreq9 & ~n62735;
  assign n62809 = ~n43259 & ~n62808;
  assign n62810 = ~i_hbusreq4 & ~n62809;
  assign n62811 = ~n43258 & ~n62810;
  assign n62812 = ~controllable_hgrant4 & ~n62811;
  assign n62813 = ~n62807 & ~n62812;
  assign n62814 = ~i_hbusreq5 & ~n62813;
  assign n62815 = ~n43247 & ~n62814;
  assign n62816 = ~controllable_hgrant5 & ~n62815;
  assign n62817 = ~n62802 & ~n62816;
  assign n62818 = ~controllable_hmaster2 & ~n62817;
  assign n62819 = ~n62675 & ~n62818;
  assign n62820 = ~controllable_hmaster1 & ~n62819;
  assign n62821 = ~n62674 & ~n62820;
  assign n62822 = ~i_hbusreq6 & ~n62821;
  assign n62823 = ~n43239 & ~n62822;
  assign n62824 = ~controllable_hgrant6 & ~n62823;
  assign n62825 = ~n62797 & ~n62824;
  assign n62826 = ~controllable_hmaster0 & ~n62825;
  assign n62827 = ~n62756 & ~n62826;
  assign n62828 = ~i_hlock8 & ~n62827;
  assign n62829 = ~n62792 & ~n62828;
  assign n62830 = ~i_hbusreq8 & ~n62829;
  assign n62831 = ~n45360 & ~n62830;
  assign n62832 = controllable_hmaster3 & ~n62831;
  assign n62833 = i_hbusreq8 & ~n62603;
  assign n62834 = ~n8217 & ~n24860;
  assign n62835 = ~n48350 & ~n62834;
  assign n62836 = ~i_hbusreq6 & ~n62835;
  assign n62837 = ~n43311 & ~n62836;
  assign n62838 = controllable_hgrant6 & ~n62837;
  assign n62839 = controllable_hmaster2 & ~n62781;
  assign n62840 = ~n8378 & ~n24820;
  assign n62841 = ~n48358 & ~n62840;
  assign n62842 = ~i_hbusreq5 & ~n62841;
  assign n62843 = ~n43320 & ~n62842;
  assign n62844 = controllable_hgrant5 & ~n62843;
  assign n62845 = ~n8426 & ~n24814;
  assign n62846 = ~n48367 & ~n62845;
  assign n62847 = ~i_hbusreq9 & ~n62846;
  assign n62848 = ~n43329 & ~n62847;
  assign n62849 = ~i_hbusreq4 & ~n62848;
  assign n62850 = ~n43328 & ~n62849;
  assign n62851 = controllable_hgrant4 & ~n62850;
  assign n62852 = ~n8365 & ~n24704;
  assign n62853 = ~n48378 & ~n62852;
  assign n62854 = i_hlock3 & ~n62853;
  assign n62855 = ~n8365 & ~n24714;
  assign n62856 = ~n48382 & ~n62855;
  assign n62857 = ~i_hlock3 & ~n62856;
  assign n62858 = ~n62854 & ~n62857;
  assign n62859 = ~i_hbusreq3 & ~n62858;
  assign n62860 = ~n43340 & ~n62859;
  assign n62861 = controllable_hgrant3 & ~n62860;
  assign n62862 = i_hlock3 & ~n62711;
  assign n62863 = ~i_hlock3 & ~n62731;
  assign n62864 = ~n62862 & ~n62863;
  assign n62865 = ~i_hbusreq3 & ~n62864;
  assign n62866 = ~n43353 & ~n62865;
  assign n62867 = ~controllable_hgrant3 & ~n62866;
  assign n62868 = ~n62861 & ~n62867;
  assign n62869 = ~i_hbusreq9 & ~n62868;
  assign n62870 = ~n43339 & ~n62869;
  assign n62871 = ~i_hbusreq4 & ~n62870;
  assign n62872 = ~n43338 & ~n62871;
  assign n62873 = ~controllable_hgrant4 & ~n62872;
  assign n62874 = ~n62851 & ~n62873;
  assign n62875 = ~i_hbusreq5 & ~n62874;
  assign n62876 = ~n43327 & ~n62875;
  assign n62877 = ~controllable_hgrant5 & ~n62876;
  assign n62878 = ~n62844 & ~n62877;
  assign n62879 = ~controllable_hmaster2 & ~n62878;
  assign n62880 = ~n62839 & ~n62879;
  assign n62881 = controllable_hmaster1 & ~n62880;
  assign n62882 = ~n8378 & ~n33995;
  assign n62883 = ~n48412 & ~n62882;
  assign n62884 = i_hlock5 & ~n62883;
  assign n62885 = ~n8378 & ~n34021;
  assign n62886 = ~n48416 & ~n62885;
  assign n62887 = ~i_hlock5 & ~n62886;
  assign n62888 = ~n62884 & ~n62887;
  assign n62889 = ~i_hbusreq5 & ~n62888;
  assign n62890 = ~n43374 & ~n62889;
  assign n62891 = controllable_hgrant5 & ~n62890;
  assign n62892 = i_hlock5 & ~n62777;
  assign n62893 = ~i_hlock5 & ~n62813;
  assign n62894 = ~n62892 & ~n62893;
  assign n62895 = ~i_hbusreq5 & ~n62894;
  assign n62896 = ~n43387 & ~n62895;
  assign n62897 = ~controllable_hgrant5 & ~n62896;
  assign n62898 = ~n62891 & ~n62897;
  assign n62899 = controllable_hmaster2 & ~n62898;
  assign n62900 = ~n8378 & ~n24852;
  assign n62901 = ~n48434 & ~n62900;
  assign n62902 = ~i_hbusreq5 & ~n62901;
  assign n62903 = ~n43396 & ~n62902;
  assign n62904 = controllable_hgrant5 & ~n62903;
  assign n62905 = ~n8426 & ~n24846;
  assign n62906 = ~n48443 & ~n62905;
  assign n62907 = ~i_hbusreq9 & ~n62906;
  assign n62908 = ~n43405 & ~n62907;
  assign n62909 = ~i_hbusreq4 & ~n62908;
  assign n62910 = ~n43404 & ~n62909;
  assign n62911 = controllable_hgrant4 & ~n62910;
  assign n62912 = ~n8365 & ~n24842;
  assign n62913 = ~n48454 & ~n62912;
  assign n62914 = ~i_hbusreq3 & ~n62913;
  assign n62915 = ~n43416 & ~n62914;
  assign n62916 = controllable_hgrant3 & ~n62915;
  assign n62917 = ~n8389 & ~n24700;
  assign n62918 = ~n48462 & ~n62917;
  assign n62919 = i_hlock1 & ~n62918;
  assign n62920 = ~n8389 & ~n24710;
  assign n62921 = ~n48466 & ~n62920;
  assign n62922 = ~i_hlock1 & ~n62921;
  assign n62923 = ~n62919 & ~n62922;
  assign n62924 = ~i_hbusreq1 & ~n62923;
  assign n62925 = ~n43424 & ~n62924;
  assign n62926 = controllable_hgrant1 & ~n62925;
  assign n62927 = i_hlock1 & ~n62707;
  assign n62928 = ~i_hlock1 & ~n62727;
  assign n62929 = ~n62927 & ~n62928;
  assign n62930 = ~i_hbusreq1 & ~n62929;
  assign n62931 = ~n43437 & ~n62930;
  assign n62932 = ~controllable_hgrant1 & ~n62931;
  assign n62933 = ~n62926 & ~n62932;
  assign n62934 = ~i_hbusreq3 & ~n62933;
  assign n62935 = ~n43423 & ~n62934;
  assign n62936 = ~controllable_hgrant3 & ~n62935;
  assign n62937 = ~n62916 & ~n62936;
  assign n62938 = ~i_hbusreq9 & ~n62937;
  assign n62939 = ~n43415 & ~n62938;
  assign n62940 = ~i_hbusreq4 & ~n62939;
  assign n62941 = ~n43414 & ~n62940;
  assign n62942 = ~controllable_hgrant4 & ~n62941;
  assign n62943 = ~n62911 & ~n62942;
  assign n62944 = ~i_hbusreq5 & ~n62943;
  assign n62945 = ~n43403 & ~n62944;
  assign n62946 = ~controllable_hgrant5 & ~n62945;
  assign n62947 = ~n62904 & ~n62946;
  assign n62948 = ~controllable_hmaster2 & ~n62947;
  assign n62949 = ~n62899 & ~n62948;
  assign n62950 = ~controllable_hmaster1 & ~n62949;
  assign n62951 = ~n62881 & ~n62950;
  assign n62952 = ~i_hbusreq6 & ~n62951;
  assign n62953 = ~n43318 & ~n62952;
  assign n62954 = ~controllable_hgrant6 & ~n62953;
  assign n62955 = ~n62838 & ~n62954;
  assign n62956 = controllable_hmaster0 & ~n62955;
  assign n62957 = i_hbusreq6 & ~n62591;
  assign n62958 = ~n24886 & ~n34000;
  assign n62959 = controllable_hmaster1 & ~n62958;
  assign n62960 = ~n24902 & ~n62959;
  assign n62961 = ~n8217 & ~n62960;
  assign n62962 = ~n48508 & ~n62961;
  assign n62963 = i_hlock6 & ~n62962;
  assign n62964 = ~n24886 & ~n34026;
  assign n62965 = controllable_hmaster1 & ~n62964;
  assign n62966 = ~n24902 & ~n62965;
  assign n62967 = ~n8217 & ~n62966;
  assign n62968 = ~n48518 & ~n62967;
  assign n62969 = ~i_hlock6 & ~n62968;
  assign n62970 = ~n62963 & ~n62969;
  assign n62971 = ~i_hbusreq6 & ~n62970;
  assign n62972 = ~n62957 & ~n62971;
  assign n62973 = controllable_hgrant6 & ~n62972;
  assign n62974 = i_hbusreq6 & ~n62599;
  assign n62975 = ~n8378 & ~n24881;
  assign n62976 = ~n48531 & ~n62975;
  assign n62977 = ~i_hbusreq5 & ~n62976;
  assign n62978 = ~n43494 & ~n62977;
  assign n62979 = controllable_hgrant5 & ~n62978;
  assign n62980 = ~n8426 & ~n24875;
  assign n62981 = ~n48540 & ~n62980;
  assign n62982 = ~i_hbusreq9 & ~n62981;
  assign n62983 = ~n43503 & ~n62982;
  assign n62984 = ~i_hbusreq4 & ~n62983;
  assign n62985 = ~n43502 & ~n62984;
  assign n62986 = controllable_hgrant4 & ~n62985;
  assign n62987 = ~n8365 & ~n24871;
  assign n62988 = ~n48551 & ~n62987;
  assign n62989 = ~i_hbusreq3 & ~n62988;
  assign n62990 = ~n43514 & ~n62989;
  assign n62991 = controllable_hgrant3 & ~n62990;
  assign n62992 = ~n8389 & ~n24867;
  assign n62993 = ~n48559 & ~n62992;
  assign n62994 = ~i_hbusreq1 & ~n62993;
  assign n62995 = ~n43522 & ~n62994;
  assign n62996 = controllable_hgrant1 & ~n62995;
  assign n62997 = ~n7733 & ~n43559;
  assign n62998 = ~n42953 & ~n48573;
  assign n62999 = i_hlock0 & ~n62998;
  assign n63000 = ~n43552 & ~n62999;
  assign n63001 = ~i_hbusreq0 & ~n63000;
  assign n63002 = ~n43547 & ~n63001;
  assign n63003 = ~i_hbusreq2 & ~n63002;
  assign n63004 = ~n43546 & ~n63003;
  assign n63005 = controllable_hgrant2 & ~n63004;
  assign n63006 = ~n24664 & ~n63005;
  assign n63007 = n7733 & ~n63006;
  assign n63008 = ~n62997 & ~n63007;
  assign n63009 = n7928 & ~n63008;
  assign n63010 = ~n43545 & ~n63009;
  assign n63011 = ~i_hbusreq1 & ~n63010;
  assign n63012 = ~n43529 & ~n63011;
  assign n63013 = ~controllable_hgrant1 & ~n63012;
  assign n63014 = ~n62996 & ~n63013;
  assign n63015 = ~i_hbusreq3 & ~n63014;
  assign n63016 = ~n43521 & ~n63015;
  assign n63017 = ~controllable_hgrant3 & ~n63016;
  assign n63018 = ~n62991 & ~n63017;
  assign n63019 = ~i_hbusreq9 & ~n63018;
  assign n63020 = ~n43513 & ~n63019;
  assign n63021 = ~i_hbusreq4 & ~n63020;
  assign n63022 = ~n43512 & ~n63021;
  assign n63023 = ~controllable_hgrant4 & ~n63022;
  assign n63024 = ~n62986 & ~n63023;
  assign n63025 = ~i_hbusreq5 & ~n63024;
  assign n63026 = ~n43501 & ~n63025;
  assign n63027 = ~controllable_hgrant5 & ~n63026;
  assign n63028 = ~n62979 & ~n63027;
  assign n63029 = ~controllable_hmaster2 & ~n63028;
  assign n63030 = ~n62839 & ~n63029;
  assign n63031 = controllable_hmaster1 & ~n63030;
  assign n63032 = ~n8378 & ~n24895;
  assign n63033 = ~n48610 & ~n63032;
  assign n63034 = ~i_hbusreq5 & ~n63033;
  assign n63035 = ~n43583 & ~n63034;
  assign n63036 = controllable_hgrant5 & ~n63035;
  assign n63037 = ~n8426 & ~n24708;
  assign n63038 = ~n48619 & ~n63037;
  assign n63039 = ~i_hbusreq9 & ~n63038;
  assign n63040 = ~n43592 & ~n63039;
  assign n63041 = i_hlock4 & ~n63040;
  assign n63042 = ~n8426 & ~n24718;
  assign n63043 = ~n48626 & ~n63042;
  assign n63044 = ~i_hbusreq9 & ~n63043;
  assign n63045 = ~n43599 & ~n63044;
  assign n63046 = ~i_hlock4 & ~n63045;
  assign n63047 = ~n63041 & ~n63046;
  assign n63048 = ~i_hbusreq4 & ~n63047;
  assign n63049 = ~n43591 & ~n63048;
  assign n63050 = controllable_hgrant4 & ~n63049;
  assign n63051 = i_hlock4 & ~n62773;
  assign n63052 = ~i_hlock4 & ~n62809;
  assign n63053 = ~n63051 & ~n63052;
  assign n63054 = ~i_hbusreq4 & ~n63053;
  assign n63055 = ~n43610 & ~n63054;
  assign n63056 = ~controllable_hgrant4 & ~n63055;
  assign n63057 = ~n63050 & ~n63056;
  assign n63058 = ~i_hbusreq5 & ~n63057;
  assign n63059 = ~n43590 & ~n63058;
  assign n63060 = ~controllable_hgrant5 & ~n63059;
  assign n63061 = ~n63036 & ~n63060;
  assign n63062 = controllable_hmaster2 & ~n63061;
  assign n63063 = ~n48715 & ~n63062;
  assign n63064 = ~controllable_hmaster1 & ~n63063;
  assign n63065 = ~n63031 & ~n63064;
  assign n63066 = i_hlock6 & ~n63065;
  assign n63067 = controllable_hmaster2 & ~n62817;
  assign n63068 = ~n63029 & ~n63067;
  assign n63069 = controllable_hmaster1 & ~n63068;
  assign n63070 = ~n63064 & ~n63069;
  assign n63071 = ~i_hlock6 & ~n63070;
  assign n63072 = ~n63066 & ~n63071;
  assign n63073 = ~i_hbusreq6 & ~n63072;
  assign n63074 = ~n62974 & ~n63073;
  assign n63075 = ~controllable_hgrant6 & ~n63074;
  assign n63076 = ~n62973 & ~n63075;
  assign n63077 = ~controllable_hmaster0 & ~n63076;
  assign n63078 = ~n62956 & ~n63077;
  assign n63079 = ~i_hbusreq8 & ~n63078;
  assign n63080 = ~n62833 & ~n63079;
  assign n63081 = ~controllable_hmaster3 & ~n63080;
  assign n63082 = ~n62832 & ~n63081;
  assign n63083 = i_hlock7 & ~n63082;
  assign n63084 = i_hbusreq8 & ~n62607;
  assign n63085 = ~n8217 & ~n24925;
  assign n63086 = ~n48737 & ~n63085;
  assign n63087 = ~i_hbusreq6 & ~n63086;
  assign n63088 = ~n43714 & ~n63087;
  assign n63089 = controllable_hgrant6 & ~n63088;
  assign n63090 = ~n62879 & ~n63067;
  assign n63091 = controllable_hmaster1 & ~n63090;
  assign n63092 = ~n62950 & ~n63091;
  assign n63093 = ~i_hbusreq6 & ~n63092;
  assign n63094 = ~n43721 & ~n63093;
  assign n63095 = ~controllable_hgrant6 & ~n63094;
  assign n63096 = ~n63089 & ~n63095;
  assign n63097 = controllable_hmaster0 & ~n63096;
  assign n63098 = ~n63077 & ~n63097;
  assign n63099 = ~i_hbusreq8 & ~n63098;
  assign n63100 = ~n63084 & ~n63099;
  assign n63101 = ~controllable_hmaster3 & ~n63100;
  assign n63102 = ~n62832 & ~n63101;
  assign n63103 = ~i_hlock7 & ~n63102;
  assign n63104 = ~n63083 & ~n63103;
  assign n63105 = ~i_hbusreq7 & ~n63104;
  assign n63106 = ~n62612 & ~n63105;
  assign n63107 = ~n7924 & ~n63106;
  assign n63108 = ~n24952 & ~n44001;
  assign n63109 = ~n8217 & ~n63108;
  assign n63110 = ~n43999 & ~n63109;
  assign n63111 = i_hlock6 & ~n63110;
  assign n63112 = ~n24952 & ~n44011;
  assign n63113 = ~n8217 & ~n63112;
  assign n63114 = ~n44009 & ~n63113;
  assign n63115 = ~i_hlock6 & ~n63114;
  assign n63116 = ~n63111 & ~n63115;
  assign n63117 = controllable_hgrant6 & ~n63116;
  assign n63118 = ~n8378 & ~n24947;
  assign n63119 = ~n44076 & ~n63118;
  assign n63120 = controllable_hgrant5 & ~n63119;
  assign n63121 = ~n8426 & ~n24945;
  assign n63122 = ~n44080 & ~n63121;
  assign n63123 = controllable_hgrant4 & ~n63122;
  assign n63124 = ~n8365 & ~n24943;
  assign n63125 = ~n44084 & ~n63124;
  assign n63126 = controllable_hgrant3 & ~n63125;
  assign n63127 = ~n8389 & ~n24941;
  assign n63128 = ~n44088 & ~n63127;
  assign n63129 = controllable_hgrant1 & ~n63128;
  assign n63130 = ~n8440 & ~n43800;
  assign n63131 = ~controllable_hgrant1 & ~n63130;
  assign n63132 = ~n63129 & ~n63131;
  assign n63133 = ~controllable_hgrant3 & ~n63132;
  assign n63134 = ~n63126 & ~n63133;
  assign n63135 = ~controllable_hgrant4 & ~n63134;
  assign n63136 = ~n63123 & ~n63135;
  assign n63137 = ~controllable_hgrant5 & ~n63136;
  assign n63138 = ~n63120 & ~n63137;
  assign n63139 = ~controllable_hmaster2 & ~n63138;
  assign n63140 = ~n44075 & ~n63139;
  assign n63141 = ~controllable_hmaster1 & ~n63140;
  assign n63142 = ~n44053 & ~n63141;
  assign n63143 = i_hlock6 & ~n63142;
  assign n63144 = ~n44108 & ~n63141;
  assign n63145 = ~i_hlock6 & ~n63144;
  assign n63146 = ~n63143 & ~n63145;
  assign n63147 = ~controllable_hgrant6 & ~n63146;
  assign n63148 = ~n63117 & ~n63147;
  assign n63149 = ~controllable_hmaster0 & ~n63148;
  assign n63150 = ~n43995 & ~n63149;
  assign n63151 = ~controllable_hmaster3 & ~n63150;
  assign n63152 = ~n45424 & ~n63151;
  assign n63153 = i_hlock7 & ~n63152;
  assign n63154 = ~n44128 & ~n63149;
  assign n63155 = ~controllable_hmaster3 & ~n63154;
  assign n63156 = ~n45424 & ~n63155;
  assign n63157 = ~i_hlock7 & ~n63156;
  assign n63158 = ~n63153 & ~n63157;
  assign n63159 = i_hbusreq7 & ~n63158;
  assign n63160 = ~n8217 & ~n34071;
  assign n63161 = ~n49089 & ~n63160;
  assign n63162 = ~i_hbusreq6 & ~n63161;
  assign n63163 = ~n45168 & ~n63162;
  assign n63164 = controllable_hgrant6 & ~n63163;
  assign n63165 = ~n8378 & ~n25009;
  assign n63166 = ~n49102 & ~n63165;
  assign n63167 = ~i_hbusreq5 & ~n63166;
  assign n63168 = ~n44144 & ~n63167;
  assign n63169 = controllable_hgrant5 & ~n63168;
  assign n63170 = ~n8426 & ~n25003;
  assign n63171 = ~n49116 & ~n63170;
  assign n63172 = ~i_hbusreq9 & ~n63171;
  assign n63173 = ~n44153 & ~n63172;
  assign n63174 = ~i_hbusreq4 & ~n63173;
  assign n63175 = ~n44152 & ~n63174;
  assign n63176 = controllable_hgrant4 & ~n63175;
  assign n63177 = ~n8365 & ~n24999;
  assign n63178 = ~n49135 & ~n63177;
  assign n63179 = ~i_hbusreq3 & ~n63178;
  assign n63180 = ~n44164 & ~n63179;
  assign n63181 = controllable_hgrant3 & ~n63180;
  assign n63182 = ~n8389 & ~n24995;
  assign n63183 = ~n49148 & ~n63182;
  assign n63184 = ~i_hbusreq1 & ~n63183;
  assign n63185 = ~n44172 & ~n63184;
  assign n63186 = controllable_hgrant1 & ~n63185;
  assign n63187 = ~n13008 & ~n49163;
  assign n63188 = i_hlock0 & ~n63187;
  assign n63189 = ~n44185 & ~n63188;
  assign n63190 = ~i_hbusreq0 & ~n63189;
  assign n63191 = ~n44181 & ~n63190;
  assign n63192 = ~i_hbusreq2 & ~n63191;
  assign n63193 = ~n44180 & ~n63192;
  assign n63194 = controllable_hgrant2 & ~n63193;
  assign n63195 = ~n49177 & ~n63194;
  assign n63196 = ~n7733 & ~n63195;
  assign n63197 = ~n12640 & ~n49183;
  assign n63198 = i_hlock0 & ~n63197;
  assign n63199 = ~n44185 & ~n63198;
  assign n63200 = ~i_hbusreq0 & ~n63199;
  assign n63201 = ~n44181 & ~n63200;
  assign n63202 = ~i_hbusreq2 & ~n63201;
  assign n63203 = ~n44180 & ~n63202;
  assign n63204 = controllable_hgrant2 & ~n63203;
  assign n63205 = ~n25023 & ~n63204;
  assign n63206 = n7733 & ~n63205;
  assign n63207 = ~n63196 & ~n63206;
  assign n63208 = n7928 & ~n63207;
  assign n63209 = ~n62652 & ~n63208;
  assign n63210 = ~i_hbusreq1 & ~n63209;
  assign n63211 = ~n44179 & ~n63210;
  assign n63212 = ~controllable_hgrant1 & ~n63211;
  assign n63213 = ~n63186 & ~n63212;
  assign n63214 = ~i_hbusreq3 & ~n63213;
  assign n63215 = ~n44171 & ~n63214;
  assign n63216 = ~controllable_hgrant3 & ~n63215;
  assign n63217 = ~n63181 & ~n63216;
  assign n63218 = ~i_hbusreq9 & ~n63217;
  assign n63219 = ~n44163 & ~n63218;
  assign n63220 = ~i_hbusreq4 & ~n63219;
  assign n63221 = ~n44162 & ~n63220;
  assign n63222 = ~controllable_hgrant4 & ~n63221;
  assign n63223 = ~n63176 & ~n63222;
  assign n63224 = ~i_hbusreq5 & ~n63223;
  assign n63225 = ~n44151 & ~n63224;
  assign n63226 = ~controllable_hgrant5 & ~n63225;
  assign n63227 = ~n63169 & ~n63226;
  assign n63228 = controllable_hmaster1 & ~n63227;
  assign n63229 = controllable_hmaster2 & ~n63227;
  assign n63230 = ~n8378 & ~n34063;
  assign n63231 = ~n49221 & ~n63230;
  assign n63232 = ~i_hbusreq5 & ~n63231;
  assign n63233 = ~n45176 & ~n63232;
  assign n63234 = controllable_hgrant5 & ~n63233;
  assign n63235 = ~n8426 & ~n25078;
  assign n63236 = ~n49232 & ~n63235;
  assign n63237 = i_hlock9 & ~n63236;
  assign n63238 = ~n8426 & ~n25108;
  assign n63239 = ~n49236 & ~n63238;
  assign n63240 = ~i_hlock9 & ~n63239;
  assign n63241 = ~n63237 & ~n63240;
  assign n63242 = ~i_hbusreq9 & ~n63241;
  assign n63243 = ~n45185 & ~n63242;
  assign n63244 = ~i_hbusreq4 & ~n63243;
  assign n63245 = ~n45184 & ~n63244;
  assign n63246 = controllable_hgrant4 & ~n63245;
  assign n63247 = ~n8365 & ~n25074;
  assign n63248 = ~n49258 & ~n63247;
  assign n63249 = ~i_hbusreq3 & ~n63248;
  assign n63250 = ~n44390 & ~n63249;
  assign n63251 = controllable_hgrant3 & ~n63250;
  assign n63252 = ~n8389 & ~n25070;
  assign n63253 = ~n49269 & ~n63252;
  assign n63254 = ~i_hbusreq1 & ~n63253;
  assign n63255 = ~n44398 & ~n63254;
  assign n63256 = controllable_hgrant1 & ~n63255;
  assign n63257 = ~n16483 & ~n17556;
  assign n63258 = i_hlock0 & ~n63257;
  assign n63259 = ~n20876 & ~n63258;
  assign n63260 = ~i_hbusreq0 & ~n63259;
  assign n63261 = ~n20873 & ~n63260;
  assign n63262 = ~i_hbusreq2 & ~n63261;
  assign n63263 = ~n20872 & ~n63262;
  assign n63264 = ~controllable_hgrant2 & n63263;
  assign n63265 = ~n44191 & ~n63264;
  assign n63266 = ~n7733 & ~n63265;
  assign n63267 = ~n24990 & ~n63204;
  assign n63268 = n7733 & ~n63267;
  assign n63269 = ~n63266 & ~n63268;
  assign n63270 = n7928 & ~n63269;
  assign n63271 = ~n8265 & ~n63270;
  assign n63272 = ~i_hbusreq1 & ~n63271;
  assign n63273 = ~n44405 & ~n63272;
  assign n63274 = ~controllable_hgrant1 & ~n63273;
  assign n63275 = ~n63256 & ~n63274;
  assign n63276 = ~i_hbusreq3 & ~n63275;
  assign n63277 = ~n44397 & ~n63276;
  assign n63278 = ~controllable_hgrant3 & ~n63277;
  assign n63279 = ~n63251 & ~n63278;
  assign n63280 = i_hlock9 & ~n63279;
  assign n63281 = ~n8365 & ~n25104;
  assign n63282 = ~n49311 & ~n63281;
  assign n63283 = ~i_hbusreq3 & ~n63282;
  assign n63284 = ~n44470 & ~n63283;
  assign n63285 = controllable_hgrant3 & ~n63284;
  assign n63286 = ~n8389 & ~n25100;
  assign n63287 = ~n49322 & ~n63286;
  assign n63288 = ~i_hbusreq1 & ~n63287;
  assign n63289 = ~n44478 & ~n63288;
  assign n63290 = controllable_hgrant1 & ~n63289;
  assign n63291 = ~n8297 & ~n63270;
  assign n63292 = ~i_hbusreq1 & ~n63291;
  assign n63293 = ~n44485 & ~n63292;
  assign n63294 = ~controllable_hgrant1 & ~n63293;
  assign n63295 = ~n63290 & ~n63294;
  assign n63296 = ~i_hbusreq3 & ~n63295;
  assign n63297 = ~n44477 & ~n63296;
  assign n63298 = ~controllable_hgrant3 & ~n63297;
  assign n63299 = ~n63285 & ~n63298;
  assign n63300 = ~i_hlock9 & ~n63299;
  assign n63301 = ~n63280 & ~n63300;
  assign n63302 = ~i_hbusreq9 & ~n63301;
  assign n63303 = ~n45195 & ~n63302;
  assign n63304 = ~i_hbusreq4 & ~n63303;
  assign n63305 = ~n45194 & ~n63304;
  assign n63306 = ~controllable_hgrant4 & ~n63305;
  assign n63307 = ~n63246 & ~n63306;
  assign n63308 = ~i_hbusreq5 & ~n63307;
  assign n63309 = ~n45183 & ~n63308;
  assign n63310 = ~controllable_hgrant5 & ~n63309;
  assign n63311 = ~n63234 & ~n63310;
  assign n63312 = ~controllable_hmaster2 & ~n63311;
  assign n63313 = ~n63229 & ~n63312;
  assign n63314 = ~controllable_hmaster1 & ~n63313;
  assign n63315 = ~n63228 & ~n63314;
  assign n63316 = ~i_hbusreq6 & ~n63315;
  assign n63317 = ~n45175 & ~n63316;
  assign n63318 = ~controllable_hgrant6 & ~n63317;
  assign n63319 = ~n63164 & ~n63318;
  assign n63320 = controllable_hmaster0 & ~n63319;
  assign n63321 = ~n8217 & ~n25092;
  assign n63322 = ~n49363 & ~n63321;
  assign n63323 = ~i_hbusreq6 & ~n63322;
  assign n63324 = ~n44362 & ~n63323;
  assign n63325 = controllable_hgrant6 & ~n63324;
  assign n63326 = ~n8378 & ~n25084;
  assign n63327 = ~n49375 & ~n63326;
  assign n63328 = ~i_hbusreq5 & ~n63327;
  assign n63329 = ~n44370 & ~n63328;
  assign n63330 = controllable_hgrant5 & ~n63329;
  assign n63331 = ~i_hbusreq9 & ~n63236;
  assign n63332 = ~n44379 & ~n63331;
  assign n63333 = ~i_hbusreq4 & ~n63332;
  assign n63334 = ~n44378 & ~n63333;
  assign n63335 = controllable_hgrant4 & ~n63334;
  assign n63336 = ~i_hbusreq9 & ~n63279;
  assign n63337 = ~n44389 & ~n63336;
  assign n63338 = ~i_hbusreq4 & ~n63337;
  assign n63339 = ~n44388 & ~n63338;
  assign n63340 = ~controllable_hgrant4 & ~n63339;
  assign n63341 = ~n63335 & ~n63340;
  assign n63342 = ~i_hbusreq5 & ~n63341;
  assign n63343 = ~n44377 & ~n63342;
  assign n63344 = ~controllable_hgrant5 & ~n63343;
  assign n63345 = ~n63330 & ~n63344;
  assign n63346 = ~controllable_hmaster2 & ~n63345;
  assign n63347 = ~n63229 & ~n63346;
  assign n63348 = ~controllable_hmaster1 & ~n63347;
  assign n63349 = ~n63228 & ~n63348;
  assign n63350 = ~i_hbusreq6 & ~n63349;
  assign n63351 = ~n44369 & ~n63350;
  assign n63352 = ~controllable_hgrant6 & ~n63351;
  assign n63353 = ~n63325 & ~n63352;
  assign n63354 = ~controllable_hmaster0 & ~n63353;
  assign n63355 = ~n63320 & ~n63354;
  assign n63356 = i_hlock8 & ~n63355;
  assign n63357 = ~n8217 & ~n25122;
  assign n63358 = ~n49417 & ~n63357;
  assign n63359 = ~i_hbusreq6 & ~n63358;
  assign n63360 = ~n44442 & ~n63359;
  assign n63361 = controllable_hgrant6 & ~n63360;
  assign n63362 = ~n8378 & ~n25114;
  assign n63363 = ~n49429 & ~n63362;
  assign n63364 = ~i_hbusreq5 & ~n63363;
  assign n63365 = ~n44450 & ~n63364;
  assign n63366 = controllable_hgrant5 & ~n63365;
  assign n63367 = ~i_hbusreq9 & ~n63239;
  assign n63368 = ~n44459 & ~n63367;
  assign n63369 = ~i_hbusreq4 & ~n63368;
  assign n63370 = ~n44458 & ~n63369;
  assign n63371 = controllable_hgrant4 & ~n63370;
  assign n63372 = ~i_hbusreq9 & ~n63299;
  assign n63373 = ~n44469 & ~n63372;
  assign n63374 = ~i_hbusreq4 & ~n63373;
  assign n63375 = ~n44468 & ~n63374;
  assign n63376 = ~controllable_hgrant4 & ~n63375;
  assign n63377 = ~n63371 & ~n63376;
  assign n63378 = ~i_hbusreq5 & ~n63377;
  assign n63379 = ~n44457 & ~n63378;
  assign n63380 = ~controllable_hgrant5 & ~n63379;
  assign n63381 = ~n63366 & ~n63380;
  assign n63382 = ~controllable_hmaster2 & ~n63381;
  assign n63383 = ~n63229 & ~n63382;
  assign n63384 = ~controllable_hmaster1 & ~n63383;
  assign n63385 = ~n63228 & ~n63384;
  assign n63386 = ~i_hbusreq6 & ~n63385;
  assign n63387 = ~n44449 & ~n63386;
  assign n63388 = ~controllable_hgrant6 & ~n63387;
  assign n63389 = ~n63361 & ~n63388;
  assign n63390 = ~controllable_hmaster0 & ~n63389;
  assign n63391 = ~n63320 & ~n63390;
  assign n63392 = ~i_hlock8 & ~n63391;
  assign n63393 = ~n63356 & ~n63392;
  assign n63394 = ~i_hbusreq8 & ~n63393;
  assign n63395 = ~n45455 & ~n63394;
  assign n63396 = controllable_hmaster3 & ~n63395;
  assign n63397 = i_hbusreq8 & ~n63150;
  assign n63398 = ~n8217 & ~n25188;
  assign n63399 = ~n49476 & ~n63398;
  assign n63400 = ~i_hbusreq6 & ~n63399;
  assign n63401 = ~n44521 & ~n63400;
  assign n63402 = controllable_hgrant6 & ~n63401;
  assign n63403 = controllable_hmaster2 & ~n63345;
  assign n63404 = ~n8378 & ~n25148;
  assign n63405 = ~n49490 & ~n63404;
  assign n63406 = ~i_hbusreq5 & ~n63405;
  assign n63407 = ~n44530 & ~n63406;
  assign n63408 = controllable_hgrant5 & ~n63407;
  assign n63409 = ~n8426 & ~n25142;
  assign n63410 = ~n49504 & ~n63409;
  assign n63411 = ~i_hbusreq9 & ~n63410;
  assign n63412 = ~n44539 & ~n63411;
  assign n63413 = ~i_hbusreq4 & ~n63412;
  assign n63414 = ~n44538 & ~n63413;
  assign n63415 = controllable_hgrant4 & ~n63414;
  assign n63416 = ~n8365 & ~n25032;
  assign n63417 = ~n49523 & ~n63416;
  assign n63418 = i_hlock3 & ~n63417;
  assign n63419 = ~n8365 & ~n25042;
  assign n63420 = ~n49527 & ~n63419;
  assign n63421 = ~i_hlock3 & ~n63420;
  assign n63422 = ~n63418 & ~n63421;
  assign n63423 = ~i_hbusreq3 & ~n63422;
  assign n63424 = ~n44550 & ~n63423;
  assign n63425 = controllable_hgrant3 & ~n63424;
  assign n63426 = i_hlock3 & ~n63275;
  assign n63427 = ~i_hlock3 & ~n63295;
  assign n63428 = ~n63426 & ~n63427;
  assign n63429 = ~i_hbusreq3 & ~n63428;
  assign n63430 = ~n44563 & ~n63429;
  assign n63431 = ~controllable_hgrant3 & ~n63430;
  assign n63432 = ~n63425 & ~n63431;
  assign n63433 = ~i_hbusreq9 & ~n63432;
  assign n63434 = ~n44549 & ~n63433;
  assign n63435 = ~i_hbusreq4 & ~n63434;
  assign n63436 = ~n44548 & ~n63435;
  assign n63437 = ~controllable_hgrant4 & ~n63436;
  assign n63438 = ~n63415 & ~n63437;
  assign n63439 = ~i_hbusreq5 & ~n63438;
  assign n63440 = ~n44537 & ~n63439;
  assign n63441 = ~controllable_hgrant5 & ~n63440;
  assign n63442 = ~n63408 & ~n63441;
  assign n63443 = ~controllable_hmaster2 & ~n63442;
  assign n63444 = ~n63403 & ~n63443;
  assign n63445 = controllable_hmaster1 & ~n63444;
  assign n63446 = ~n8378 & ~n34091;
  assign n63447 = ~n49557 & ~n63446;
  assign n63448 = i_hlock5 & ~n63447;
  assign n63449 = ~n8378 & ~n34117;
  assign n63450 = ~n49561 & ~n63449;
  assign n63451 = ~i_hlock5 & ~n63450;
  assign n63452 = ~n63448 & ~n63451;
  assign n63453 = ~i_hbusreq5 & ~n63452;
  assign n63454 = ~n44584 & ~n63453;
  assign n63455 = controllable_hgrant5 & ~n63454;
  assign n63456 = i_hlock5 & ~n63341;
  assign n63457 = ~i_hlock5 & ~n63377;
  assign n63458 = ~n63456 & ~n63457;
  assign n63459 = ~i_hbusreq5 & ~n63458;
  assign n63460 = ~n44597 & ~n63459;
  assign n63461 = ~controllable_hgrant5 & ~n63460;
  assign n63462 = ~n63455 & ~n63461;
  assign n63463 = controllable_hmaster2 & ~n63462;
  assign n63464 = ~n8378 & ~n25180;
  assign n63465 = ~n49579 & ~n63464;
  assign n63466 = ~i_hbusreq5 & ~n63465;
  assign n63467 = ~n44606 & ~n63466;
  assign n63468 = controllable_hgrant5 & ~n63467;
  assign n63469 = ~n8426 & ~n25174;
  assign n63470 = ~n49593 & ~n63469;
  assign n63471 = ~i_hbusreq9 & ~n63470;
  assign n63472 = ~n44615 & ~n63471;
  assign n63473 = ~i_hbusreq4 & ~n63472;
  assign n63474 = ~n44614 & ~n63473;
  assign n63475 = controllable_hgrant4 & ~n63474;
  assign n63476 = ~n8365 & ~n25170;
  assign n63477 = ~n49612 & ~n63476;
  assign n63478 = ~i_hbusreq3 & ~n63477;
  assign n63479 = ~n44626 & ~n63478;
  assign n63480 = controllable_hgrant3 & ~n63479;
  assign n63481 = ~n8389 & ~n25028;
  assign n63482 = ~n49625 & ~n63481;
  assign n63483 = i_hlock1 & ~n63482;
  assign n63484 = ~n8389 & ~n25038;
  assign n63485 = ~n49629 & ~n63484;
  assign n63486 = ~i_hlock1 & ~n63485;
  assign n63487 = ~n63483 & ~n63486;
  assign n63488 = ~i_hbusreq1 & ~n63487;
  assign n63489 = ~n44634 & ~n63488;
  assign n63490 = controllable_hgrant1 & ~n63489;
  assign n63491 = i_hlock1 & ~n63271;
  assign n63492 = ~i_hlock1 & ~n63291;
  assign n63493 = ~n63491 & ~n63492;
  assign n63494 = ~i_hbusreq1 & ~n63493;
  assign n63495 = ~n44647 & ~n63494;
  assign n63496 = ~controllable_hgrant1 & ~n63495;
  assign n63497 = ~n63490 & ~n63496;
  assign n63498 = ~i_hbusreq3 & ~n63497;
  assign n63499 = ~n44633 & ~n63498;
  assign n63500 = ~controllable_hgrant3 & ~n63499;
  assign n63501 = ~n63480 & ~n63500;
  assign n63502 = ~i_hbusreq9 & ~n63501;
  assign n63503 = ~n44625 & ~n63502;
  assign n63504 = ~i_hbusreq4 & ~n63503;
  assign n63505 = ~n44624 & ~n63504;
  assign n63506 = ~controllable_hgrant4 & ~n63505;
  assign n63507 = ~n63475 & ~n63506;
  assign n63508 = ~i_hbusreq5 & ~n63507;
  assign n63509 = ~n44613 & ~n63508;
  assign n63510 = ~controllable_hgrant5 & ~n63509;
  assign n63511 = ~n63468 & ~n63510;
  assign n63512 = ~controllable_hmaster2 & ~n63511;
  assign n63513 = ~n63463 & ~n63512;
  assign n63514 = ~controllable_hmaster1 & ~n63513;
  assign n63515 = ~n63445 & ~n63514;
  assign n63516 = ~i_hbusreq6 & ~n63515;
  assign n63517 = ~n44528 & ~n63516;
  assign n63518 = ~controllable_hgrant6 & ~n63517;
  assign n63519 = ~n63402 & ~n63518;
  assign n63520 = controllable_hmaster0 & ~n63519;
  assign n63521 = i_hbusreq6 & ~n63116;
  assign n63522 = ~n25214 & ~n34096;
  assign n63523 = controllable_hmaster1 & ~n63522;
  assign n63524 = ~n25257 & ~n63523;
  assign n63525 = ~n8217 & ~n63524;
  assign n63526 = ~n49671 & ~n63525;
  assign n63527 = i_hlock6 & ~n63526;
  assign n63528 = ~n25214 & ~n34122;
  assign n63529 = controllable_hmaster1 & ~n63528;
  assign n63530 = ~n25257 & ~n63529;
  assign n63531 = ~n8217 & ~n63530;
  assign n63532 = ~n49681 & ~n63531;
  assign n63533 = ~i_hlock6 & ~n63532;
  assign n63534 = ~n63527 & ~n63533;
  assign n63535 = ~i_hbusreq6 & ~n63534;
  assign n63536 = ~n63521 & ~n63535;
  assign n63537 = controllable_hgrant6 & ~n63536;
  assign n63538 = i_hbusreq6 & ~n63146;
  assign n63539 = ~n8378 & ~n25209;
  assign n63540 = ~n49694 & ~n63539;
  assign n63541 = ~i_hbusreq5 & ~n63540;
  assign n63542 = ~n44704 & ~n63541;
  assign n63543 = controllable_hgrant5 & ~n63542;
  assign n63544 = ~n8426 & ~n25203;
  assign n63545 = ~n49708 & ~n63544;
  assign n63546 = ~i_hbusreq9 & ~n63545;
  assign n63547 = ~n44713 & ~n63546;
  assign n63548 = ~i_hbusreq4 & ~n63547;
  assign n63549 = ~n44712 & ~n63548;
  assign n63550 = controllable_hgrant4 & ~n63549;
  assign n63551 = ~n8365 & ~n25199;
  assign n63552 = ~n49727 & ~n63551;
  assign n63553 = ~i_hbusreq3 & ~n63552;
  assign n63554 = ~n44724 & ~n63553;
  assign n63555 = controllable_hgrant3 & ~n63554;
  assign n63556 = ~n8389 & ~n25195;
  assign n63557 = ~n49740 & ~n63556;
  assign n63558 = ~i_hbusreq1 & ~n63557;
  assign n63559 = ~n44732 & ~n63558;
  assign n63560 = controllable_hgrant1 & ~n63559;
  assign n63561 = ~n44750 & ~n63264;
  assign n63562 = ~n7733 & ~n63561;
  assign n63563 = ~n42953 & ~n49183;
  assign n63564 = i_hlock0 & ~n63563;
  assign n63565 = ~n44744 & ~n63564;
  assign n63566 = ~i_hbusreq0 & ~n63565;
  assign n63567 = ~n44741 & ~n63566;
  assign n63568 = ~i_hbusreq2 & ~n63567;
  assign n63569 = ~n44740 & ~n63568;
  assign n63570 = controllable_hgrant2 & ~n63569;
  assign n63571 = ~n24990 & ~n63570;
  assign n63572 = n7733 & ~n63571;
  assign n63573 = ~n63562 & ~n63572;
  assign n63574 = n7928 & ~n63573;
  assign n63575 = ~n43545 & ~n63574;
  assign n63576 = ~i_hbusreq1 & ~n63575;
  assign n63577 = ~n44739 & ~n63576;
  assign n63578 = ~controllable_hgrant1 & ~n63577;
  assign n63579 = ~n63560 & ~n63578;
  assign n63580 = ~i_hbusreq3 & ~n63579;
  assign n63581 = ~n44731 & ~n63580;
  assign n63582 = ~controllable_hgrant3 & ~n63581;
  assign n63583 = ~n63555 & ~n63582;
  assign n63584 = ~i_hbusreq9 & ~n63583;
  assign n63585 = ~n44723 & ~n63584;
  assign n63586 = ~i_hbusreq4 & ~n63585;
  assign n63587 = ~n44722 & ~n63586;
  assign n63588 = ~controllable_hgrant4 & ~n63587;
  assign n63589 = ~n63550 & ~n63588;
  assign n63590 = ~i_hbusreq5 & ~n63589;
  assign n63591 = ~n44711 & ~n63590;
  assign n63592 = ~controllable_hgrant5 & ~n63591;
  assign n63593 = ~n63543 & ~n63592;
  assign n63594 = ~controllable_hmaster2 & ~n63593;
  assign n63595 = ~n63403 & ~n63594;
  assign n63596 = controllable_hmaster1 & ~n63595;
  assign n63597 = ~n8378 & ~n25223;
  assign n63598 = ~n49798 & ~n63597;
  assign n63599 = ~i_hbusreq5 & ~n63598;
  assign n63600 = ~n44779 & ~n63599;
  assign n63601 = controllable_hgrant5 & ~n63600;
  assign n63602 = ~n8426 & ~n25036;
  assign n63603 = ~n49812 & ~n63602;
  assign n63604 = ~i_hbusreq9 & ~n63603;
  assign n63605 = ~n44788 & ~n63604;
  assign n63606 = i_hlock4 & ~n63605;
  assign n63607 = ~n8426 & ~n25046;
  assign n63608 = ~n49819 & ~n63607;
  assign n63609 = ~i_hbusreq9 & ~n63608;
  assign n63610 = ~n44795 & ~n63609;
  assign n63611 = ~i_hlock4 & ~n63610;
  assign n63612 = ~n63606 & ~n63611;
  assign n63613 = ~i_hbusreq4 & ~n63612;
  assign n63614 = ~n44787 & ~n63613;
  assign n63615 = controllable_hgrant4 & ~n63614;
  assign n63616 = i_hlock4 & ~n63337;
  assign n63617 = ~i_hlock4 & ~n63373;
  assign n63618 = ~n63616 & ~n63617;
  assign n63619 = ~i_hbusreq4 & ~n63618;
  assign n63620 = ~n44806 & ~n63619;
  assign n63621 = ~controllable_hgrant4 & ~n63620;
  assign n63622 = ~n63615 & ~n63621;
  assign n63623 = ~i_hbusreq5 & ~n63622;
  assign n63624 = ~n44786 & ~n63623;
  assign n63625 = ~controllable_hgrant5 & ~n63624;
  assign n63626 = ~n63601 & ~n63625;
  assign n63627 = controllable_hmaster2 & ~n63626;
  assign n63628 = i_hbusreq5 & ~n63119;
  assign n63629 = ~n8378 & ~n25250;
  assign n63630 = ~n49843 & ~n63629;
  assign n63631 = ~i_hbusreq5 & ~n63630;
  assign n63632 = ~n63628 & ~n63631;
  assign n63633 = controllable_hgrant5 & ~n63632;
  assign n63634 = i_hbusreq5 & ~n63136;
  assign n63635 = i_hbusreq4 & ~n63122;
  assign n63636 = i_hbusreq9 & ~n63122;
  assign n63637 = ~n8426 & ~n25244;
  assign n63638 = ~n49857 & ~n63637;
  assign n63639 = ~i_hbusreq9 & ~n63638;
  assign n63640 = ~n63636 & ~n63639;
  assign n63641 = ~i_hbusreq4 & ~n63640;
  assign n63642 = ~n63635 & ~n63641;
  assign n63643 = controllable_hgrant4 & ~n63642;
  assign n63644 = i_hbusreq4 & ~n63134;
  assign n63645 = i_hbusreq9 & ~n63134;
  assign n63646 = i_hbusreq3 & ~n63125;
  assign n63647 = ~n8365 & ~n25240;
  assign n63648 = ~n49876 & ~n63647;
  assign n63649 = ~i_hbusreq3 & ~n63648;
  assign n63650 = ~n63646 & ~n63649;
  assign n63651 = controllable_hgrant3 & ~n63650;
  assign n63652 = i_hbusreq3 & ~n63132;
  assign n63653 = i_hbusreq1 & ~n63128;
  assign n63654 = ~n8389 & ~n25236;
  assign n63655 = ~n49889 & ~n63654;
  assign n63656 = ~i_hbusreq1 & ~n63655;
  assign n63657 = ~n63653 & ~n63656;
  assign n63658 = controllable_hgrant1 & ~n63657;
  assign n63659 = i_hbusreq1 & ~n63130;
  assign n63660 = ~n43798 & ~n49911;
  assign n63661 = n7928 & ~n63660;
  assign n63662 = ~n8440 & ~n63661;
  assign n63663 = ~i_hbusreq1 & ~n63662;
  assign n63664 = ~n63659 & ~n63663;
  assign n63665 = ~controllable_hgrant1 & ~n63664;
  assign n63666 = ~n63658 & ~n63665;
  assign n63667 = ~i_hbusreq3 & ~n63666;
  assign n63668 = ~n63652 & ~n63667;
  assign n63669 = ~controllable_hgrant3 & ~n63668;
  assign n63670 = ~n63651 & ~n63669;
  assign n63671 = ~i_hbusreq9 & ~n63670;
  assign n63672 = ~n63645 & ~n63671;
  assign n63673 = ~i_hbusreq4 & ~n63672;
  assign n63674 = ~n63644 & ~n63673;
  assign n63675 = ~controllable_hgrant4 & ~n63674;
  assign n63676 = ~n63643 & ~n63675;
  assign n63677 = ~i_hbusreq5 & ~n63676;
  assign n63678 = ~n63634 & ~n63677;
  assign n63679 = ~controllable_hgrant5 & ~n63678;
  assign n63680 = ~n63633 & ~n63679;
  assign n63681 = ~controllable_hmaster2 & ~n63680;
  assign n63682 = ~n63627 & ~n63681;
  assign n63683 = ~controllable_hmaster1 & ~n63682;
  assign n63684 = ~n63596 & ~n63683;
  assign n63685 = i_hlock6 & ~n63684;
  assign n63686 = controllable_hmaster2 & ~n63381;
  assign n63687 = ~n63594 & ~n63686;
  assign n63688 = controllable_hmaster1 & ~n63687;
  assign n63689 = ~n63683 & ~n63688;
  assign n63690 = ~i_hlock6 & ~n63689;
  assign n63691 = ~n63685 & ~n63690;
  assign n63692 = ~i_hbusreq6 & ~n63691;
  assign n63693 = ~n63538 & ~n63692;
  assign n63694 = ~controllable_hgrant6 & ~n63693;
  assign n63695 = ~n63537 & ~n63694;
  assign n63696 = ~controllable_hmaster0 & ~n63695;
  assign n63697 = ~n63520 & ~n63696;
  assign n63698 = ~i_hbusreq8 & ~n63697;
  assign n63699 = ~n63397 & ~n63698;
  assign n63700 = ~controllable_hmaster3 & ~n63699;
  assign n63701 = ~n63396 & ~n63700;
  assign n63702 = i_hlock7 & ~n63701;
  assign n63703 = i_hbusreq8 & ~n63154;
  assign n63704 = ~n8217 & ~n25280;
  assign n63705 = ~n49970 & ~n63704;
  assign n63706 = ~i_hbusreq6 & ~n63705;
  assign n63707 = ~n44914 & ~n63706;
  assign n63708 = controllable_hgrant6 & ~n63707;
  assign n63709 = ~n63443 & ~n63686;
  assign n63710 = controllable_hmaster1 & ~n63709;
  assign n63711 = ~n63514 & ~n63710;
  assign n63712 = ~i_hbusreq6 & ~n63711;
  assign n63713 = ~n44921 & ~n63712;
  assign n63714 = ~controllable_hgrant6 & ~n63713;
  assign n63715 = ~n63708 & ~n63714;
  assign n63716 = controllable_hmaster0 & ~n63715;
  assign n63717 = ~n63696 & ~n63716;
  assign n63718 = ~i_hbusreq8 & ~n63717;
  assign n63719 = ~n63703 & ~n63718;
  assign n63720 = ~controllable_hmaster3 & ~n63719;
  assign n63721 = ~n63396 & ~n63720;
  assign n63722 = ~i_hlock7 & ~n63721;
  assign n63723 = ~n63702 & ~n63722;
  assign n63724 = ~i_hbusreq7 & ~n63723;
  assign n63725 = ~n63159 & ~n63724;
  assign n63726 = n7924 & ~n63725;
  assign n63727 = ~n63107 & ~n63726;
  assign n63728 = n8214 & ~n63727;
  assign n63729 = ~n62582 & ~n63728;
  assign n63730 = ~n8202 & ~n63729;
  assign n63731 = ~n61598 & ~n63730;
  assign n63732 = n7920 & ~n63731;
  assign n63733 = ~n60198 & ~n63732;
  assign n63734 = ~n7728 & ~n63733;
  assign n63735 = ~n61602 & ~n63734;
  assign n63736 = n7723 & ~n63735;
  assign n63737 = ~n7723 & ~n63733;
  assign n63738 = ~n63736 & ~n63737;
  assign n63739 = n7714 & ~n63738;
  assign n63740 = n7723 & ~n63733;
  assign n63741 = ~n45995 & ~n48793;
  assign n63742 = ~controllable_hgrant3 & ~n63741;
  assign n63743 = ~n45966 & ~n63742;
  assign n63744 = ~controllable_hgrant4 & ~n63743;
  assign n63745 = ~n45958 & ~n63744;
  assign n63746 = ~controllable_hgrant5 & ~n63745;
  assign n63747 = ~n45950 & ~n63746;
  assign n63748 = controllable_hmaster1 & ~n63747;
  assign n63749 = controllable_hmaster2 & ~n63747;
  assign n63750 = ~n46046 & ~n46149;
  assign n63751 = ~controllable_hgrant3 & ~n63750;
  assign n63752 = ~n46135 & ~n63751;
  assign n63753 = i_hlock9 & ~n63752;
  assign n63754 = ~n46085 & ~n46207;
  assign n63755 = ~controllable_hgrant3 & ~n63754;
  assign n63756 = ~n46197 & ~n63755;
  assign n63757 = ~i_hlock9 & ~n63756;
  assign n63758 = ~n63753 & ~n63757;
  assign n63759 = ~controllable_hgrant4 & ~n63758;
  assign n63760 = ~n47498 & ~n63759;
  assign n63761 = ~controllable_hgrant5 & ~n63760;
  assign n63762 = ~n47488 & ~n63761;
  assign n63763 = ~controllable_hmaster2 & ~n63762;
  assign n63764 = ~n63749 & ~n63763;
  assign n63765 = ~controllable_hmaster1 & ~n63764;
  assign n63766 = ~n63748 & ~n63765;
  assign n63767 = ~controllable_hgrant6 & ~n63766;
  assign n63768 = ~n47480 & ~n63767;
  assign n63769 = controllable_hmaster0 & ~n63768;
  assign n63770 = ~controllable_hgrant4 & ~n63752;
  assign n63771 = ~n46127 & ~n63770;
  assign n63772 = ~controllable_hgrant5 & ~n63771;
  assign n63773 = ~n46119 & ~n63772;
  assign n63774 = ~controllable_hmaster2 & ~n63773;
  assign n63775 = ~n63749 & ~n63774;
  assign n63776 = ~controllable_hmaster1 & ~n63775;
  assign n63777 = ~n63748 & ~n63776;
  assign n63778 = ~controllable_hgrant6 & ~n63777;
  assign n63779 = ~n46111 & ~n63778;
  assign n63780 = ~controllable_hmaster0 & ~n63779;
  assign n63781 = ~n63769 & ~n63780;
  assign n63782 = i_hlock8 & ~n63781;
  assign n63783 = ~controllable_hgrant4 & ~n63756;
  assign n63784 = ~n46189 & ~n63783;
  assign n63785 = ~controllable_hgrant5 & ~n63784;
  assign n63786 = ~n46181 & ~n63785;
  assign n63787 = ~controllable_hmaster2 & ~n63786;
  assign n63788 = ~n63749 & ~n63787;
  assign n63789 = ~controllable_hmaster1 & ~n63788;
  assign n63790 = ~n63748 & ~n63789;
  assign n63791 = ~controllable_hgrant6 & ~n63790;
  assign n63792 = ~n46173 & ~n63791;
  assign n63793 = ~controllable_hmaster0 & ~n63792;
  assign n63794 = ~n63769 & ~n63793;
  assign n63795 = ~i_hlock8 & ~n63794;
  assign n63796 = ~n63782 & ~n63795;
  assign n63797 = controllable_hmaster3 & ~n63796;
  assign n63798 = ~n8217 & ~n38750;
  assign n63799 = ~n43905 & ~n63798;
  assign n63800 = i_hlock6 & ~n63799;
  assign n63801 = ~n8217 & ~n38756;
  assign n63802 = ~n43905 & ~n63801;
  assign n63803 = ~i_hlock6 & ~n63802;
  assign n63804 = ~n63800 & ~n63803;
  assign n63805 = controllable_hgrant6 & ~n63804;
  assign n63806 = controllable_hmaster2 & ~n63773;
  assign n63807 = i_hlock3 & ~n63750;
  assign n63808 = ~i_hlock3 & ~n63754;
  assign n63809 = ~n63807 & ~n63808;
  assign n63810 = ~controllable_hgrant3 & ~n63809;
  assign n63811 = ~n46258 & ~n63810;
  assign n63812 = ~controllable_hgrant4 & ~n63811;
  assign n63813 = ~n46250 & ~n63812;
  assign n63814 = ~controllable_hgrant5 & ~n63813;
  assign n63815 = ~n46242 & ~n63814;
  assign n63816 = ~controllable_hmaster2 & ~n63815;
  assign n63817 = ~n63806 & ~n63816;
  assign n63818 = controllable_hmaster1 & ~n63817;
  assign n63819 = i_hlock5 & ~n63771;
  assign n63820 = ~i_hlock5 & ~n63784;
  assign n63821 = ~n63819 & ~n63820;
  assign n63822 = ~controllable_hgrant5 & ~n63821;
  assign n63823 = ~n46278 & ~n63822;
  assign n63824 = controllable_hmaster2 & ~n63823;
  assign n63825 = ~n48929 & ~n63824;
  assign n63826 = ~controllable_hmaster1 & ~n63825;
  assign n63827 = ~n63818 & ~n63826;
  assign n63828 = ~controllable_hgrant6 & ~n63827;
  assign n63829 = ~n63805 & ~n63828;
  assign n63830 = controllable_hmaster0 & ~n63829;
  assign n63831 = ~n46398 & ~n48967;
  assign n63832 = ~controllable_hgrant3 & ~n63831;
  assign n63833 = ~n46372 & ~n63832;
  assign n63834 = ~controllable_hgrant4 & ~n63833;
  assign n63835 = ~n46364 & ~n63834;
  assign n63836 = ~controllable_hgrant5 & ~n63835;
  assign n63837 = ~n46356 & ~n63836;
  assign n63838 = ~controllable_hmaster2 & ~n63837;
  assign n63839 = ~n63806 & ~n63838;
  assign n63840 = controllable_hmaster1 & ~n63839;
  assign n63841 = i_hlock4 & ~n63752;
  assign n63842 = ~i_hlock4 & ~n63756;
  assign n63843 = ~n63841 & ~n63842;
  assign n63844 = ~controllable_hgrant4 & ~n63843;
  assign n63845 = ~n46424 & ~n63844;
  assign n63846 = ~controllable_hgrant5 & ~n63845;
  assign n63847 = ~n46416 & ~n63846;
  assign n63848 = controllable_hmaster2 & ~n63847;
  assign n63849 = ~n46466 & ~n49049;
  assign n63850 = ~controllable_hgrant3 & ~n63849;
  assign n63851 = ~n46456 & ~n63850;
  assign n63852 = ~controllable_hgrant4 & ~n63851;
  assign n63853 = ~n46448 & ~n63852;
  assign n63854 = ~controllable_hgrant5 & ~n63853;
  assign n63855 = ~n46440 & ~n63854;
  assign n63856 = ~controllable_hmaster2 & ~n63855;
  assign n63857 = ~n63848 & ~n63856;
  assign n63858 = ~controllable_hmaster1 & ~n63857;
  assign n63859 = ~n63840 & ~n63858;
  assign n63860 = i_hlock6 & ~n63859;
  assign n63861 = controllable_hmaster2 & ~n63786;
  assign n63862 = ~n63838 & ~n63861;
  assign n63863 = controllable_hmaster1 & ~n63862;
  assign n63864 = ~n63858 & ~n63863;
  assign n63865 = ~i_hlock6 & ~n63864;
  assign n63866 = ~n63860 & ~n63865;
  assign n63867 = ~controllable_hgrant6 & ~n63866;
  assign n63868 = ~n46348 & ~n63867;
  assign n63869 = ~controllable_hmaster0 & ~n63868;
  assign n63870 = ~n63830 & ~n63869;
  assign n63871 = ~controllable_hmaster3 & ~n63870;
  assign n63872 = ~n63797 & ~n63871;
  assign n63873 = i_hlock7 & ~n63872;
  assign n63874 = ~n8217 & ~n38766;
  assign n63875 = ~n44119 & ~n63874;
  assign n63876 = i_hlock6 & ~n63875;
  assign n63877 = ~n8217 & ~n38772;
  assign n63878 = ~n44119 & ~n63877;
  assign n63879 = ~i_hlock6 & ~n63878;
  assign n63880 = ~n63876 & ~n63879;
  assign n63881 = controllable_hgrant6 & ~n63880;
  assign n63882 = ~n63816 & ~n63861;
  assign n63883 = controllable_hmaster1 & ~n63882;
  assign n63884 = ~n63826 & ~n63883;
  assign n63885 = ~controllable_hgrant6 & ~n63884;
  assign n63886 = ~n63881 & ~n63885;
  assign n63887 = controllable_hmaster0 & ~n63886;
  assign n63888 = ~n63869 & ~n63887;
  assign n63889 = ~controllable_hmaster3 & ~n63888;
  assign n63890 = ~n63797 & ~n63889;
  assign n63891 = ~i_hlock7 & ~n63890;
  assign n63892 = ~n63873 & ~n63891;
  assign n63893 = i_hbusreq7 & ~n63892;
  assign n63894 = i_hbusreq8 & ~n63796;
  assign n63895 = i_hbusreq6 & ~n63766;
  assign n63896 = i_hbusreq5 & ~n63745;
  assign n63897 = i_hbusreq4 & ~n63743;
  assign n63898 = i_hbusreq9 & ~n63743;
  assign n63899 = i_hbusreq3 & ~n63741;
  assign n63900 = ~n46605 & ~n62221;
  assign n63901 = ~i_hbusreq3 & ~n63900;
  assign n63902 = ~n63899 & ~n63901;
  assign n63903 = ~controllable_hgrant3 & ~n63902;
  assign n63904 = ~n46566 & ~n63903;
  assign n63905 = ~i_hbusreq9 & ~n63904;
  assign n63906 = ~n63898 & ~n63905;
  assign n63907 = ~i_hbusreq4 & ~n63906;
  assign n63908 = ~n63897 & ~n63907;
  assign n63909 = ~controllable_hgrant4 & ~n63908;
  assign n63910 = ~n46553 & ~n63909;
  assign n63911 = ~i_hbusreq5 & ~n63910;
  assign n63912 = ~n63896 & ~n63911;
  assign n63913 = ~controllable_hgrant5 & ~n63912;
  assign n63914 = ~n46535 & ~n63913;
  assign n63915 = controllable_hmaster1 & ~n63914;
  assign n63916 = controllable_hmaster2 & ~n63914;
  assign n63917 = i_hbusreq5 & ~n63760;
  assign n63918 = i_hbusreq4 & ~n63758;
  assign n63919 = i_hbusreq9 & ~n63758;
  assign n63920 = i_hbusreq3 & ~n63750;
  assign n63921 = ~n46856 & ~n62253;
  assign n63922 = ~i_hbusreq3 & ~n63921;
  assign n63923 = ~n63920 & ~n63922;
  assign n63924 = ~controllable_hgrant3 & ~n63923;
  assign n63925 = ~n46835 & ~n63924;
  assign n63926 = i_hlock9 & ~n63925;
  assign n63927 = i_hbusreq3 & ~n63754;
  assign n63928 = ~n46953 & ~n62271;
  assign n63929 = ~i_hbusreq3 & ~n63928;
  assign n63930 = ~n63927 & ~n63929;
  assign n63931 = ~controllable_hgrant3 & ~n63930;
  assign n63932 = ~n46936 & ~n63931;
  assign n63933 = ~i_hlock9 & ~n63932;
  assign n63934 = ~n63926 & ~n63933;
  assign n63935 = ~i_hbusreq9 & ~n63934;
  assign n63936 = ~n63919 & ~n63935;
  assign n63937 = ~i_hbusreq4 & ~n63936;
  assign n63938 = ~n63918 & ~n63937;
  assign n63939 = ~controllable_hgrant4 & ~n63938;
  assign n63940 = ~n47630 & ~n63939;
  assign n63941 = ~i_hbusreq5 & ~n63940;
  assign n63942 = ~n63917 & ~n63941;
  assign n63943 = ~controllable_hgrant5 & ~n63942;
  assign n63944 = ~n47610 & ~n63943;
  assign n63945 = ~controllable_hmaster2 & ~n63944;
  assign n63946 = ~n63916 & ~n63945;
  assign n63947 = ~controllable_hmaster1 & ~n63946;
  assign n63948 = ~n63915 & ~n63947;
  assign n63949 = ~i_hbusreq6 & ~n63948;
  assign n63950 = ~n63895 & ~n63949;
  assign n63951 = ~controllable_hgrant6 & ~n63950;
  assign n63952 = ~n47598 & ~n63951;
  assign n63953 = controllable_hmaster0 & ~n63952;
  assign n63954 = i_hbusreq6 & ~n63777;
  assign n63955 = i_hbusreq5 & ~n63771;
  assign n63956 = i_hbusreq4 & ~n63752;
  assign n63957 = i_hbusreq9 & ~n63752;
  assign n63958 = ~i_hbusreq9 & ~n63925;
  assign n63959 = ~n63957 & ~n63958;
  assign n63960 = ~i_hbusreq4 & ~n63959;
  assign n63961 = ~n63956 & ~n63960;
  assign n63962 = ~controllable_hgrant4 & ~n63961;
  assign n63963 = ~n46822 & ~n63962;
  assign n63964 = ~i_hbusreq5 & ~n63963;
  assign n63965 = ~n63955 & ~n63964;
  assign n63966 = ~controllable_hgrant5 & ~n63965;
  assign n63967 = ~n46804 & ~n63966;
  assign n63968 = ~controllable_hmaster2 & ~n63967;
  assign n63969 = ~n63916 & ~n63968;
  assign n63970 = ~controllable_hmaster1 & ~n63969;
  assign n63971 = ~n63915 & ~n63970;
  assign n63972 = ~i_hbusreq6 & ~n63971;
  assign n63973 = ~n63954 & ~n63972;
  assign n63974 = ~controllable_hgrant6 & ~n63973;
  assign n63975 = ~n46792 & ~n63974;
  assign n63976 = ~controllable_hmaster0 & ~n63975;
  assign n63977 = ~n63953 & ~n63976;
  assign n63978 = i_hlock8 & ~n63977;
  assign n63979 = i_hbusreq6 & ~n63790;
  assign n63980 = i_hbusreq5 & ~n63784;
  assign n63981 = i_hbusreq4 & ~n63756;
  assign n63982 = i_hbusreq9 & ~n63756;
  assign n63983 = ~i_hbusreq9 & ~n63932;
  assign n63984 = ~n63982 & ~n63983;
  assign n63985 = ~i_hbusreq4 & ~n63984;
  assign n63986 = ~n63981 & ~n63985;
  assign n63987 = ~controllable_hgrant4 & ~n63986;
  assign n63988 = ~n46923 & ~n63987;
  assign n63989 = ~i_hbusreq5 & ~n63988;
  assign n63990 = ~n63980 & ~n63989;
  assign n63991 = ~controllable_hgrant5 & ~n63990;
  assign n63992 = ~n46905 & ~n63991;
  assign n63993 = ~controllable_hmaster2 & ~n63992;
  assign n63994 = ~n63916 & ~n63993;
  assign n63995 = ~controllable_hmaster1 & ~n63994;
  assign n63996 = ~n63915 & ~n63995;
  assign n63997 = ~i_hbusreq6 & ~n63996;
  assign n63998 = ~n63979 & ~n63997;
  assign n63999 = ~controllable_hgrant6 & ~n63998;
  assign n64000 = ~n46893 & ~n63999;
  assign n64001 = ~controllable_hmaster0 & ~n64000;
  assign n64002 = ~n63953 & ~n64001;
  assign n64003 = ~i_hlock8 & ~n64002;
  assign n64004 = ~n63978 & ~n64003;
  assign n64005 = ~i_hbusreq8 & ~n64004;
  assign n64006 = ~n63894 & ~n64005;
  assign n64007 = controllable_hmaster3 & ~n64006;
  assign n64008 = i_hbusreq8 & ~n63870;
  assign n64009 = i_hbusreq6 & ~n63804;
  assign n64010 = ~n8217 & ~n38786;
  assign n64011 = ~n62354 & ~n64010;
  assign n64012 = i_hlock6 & ~n64011;
  assign n64013 = ~n8217 & ~n38795;
  assign n64014 = ~n62354 & ~n64013;
  assign n64015 = ~i_hlock6 & ~n64014;
  assign n64016 = ~n64012 & ~n64015;
  assign n64017 = ~i_hbusreq6 & ~n64016;
  assign n64018 = ~n64009 & ~n64017;
  assign n64019 = controllable_hgrant6 & ~n64018;
  assign n64020 = i_hbusreq6 & ~n63827;
  assign n64021 = controllable_hmaster2 & ~n63967;
  assign n64022 = i_hbusreq5 & ~n63813;
  assign n64023 = i_hbusreq4 & ~n63811;
  assign n64024 = i_hbusreq9 & ~n63811;
  assign n64025 = i_hbusreq3 & ~n63809;
  assign n64026 = i_hlock3 & ~n63921;
  assign n64027 = ~i_hlock3 & ~n63928;
  assign n64028 = ~n64026 & ~n64027;
  assign n64029 = ~i_hbusreq3 & ~n64028;
  assign n64030 = ~n64025 & ~n64029;
  assign n64031 = ~controllable_hgrant3 & ~n64030;
  assign n64032 = ~n47039 & ~n64031;
  assign n64033 = ~i_hbusreq9 & ~n64032;
  assign n64034 = ~n64024 & ~n64033;
  assign n64035 = ~i_hbusreq4 & ~n64034;
  assign n64036 = ~n64023 & ~n64035;
  assign n64037 = ~controllable_hgrant4 & ~n64036;
  assign n64038 = ~n47026 & ~n64037;
  assign n64039 = ~i_hbusreq5 & ~n64038;
  assign n64040 = ~n64022 & ~n64039;
  assign n64041 = ~controllable_hgrant5 & ~n64040;
  assign n64042 = ~n47008 & ~n64041;
  assign n64043 = ~controllable_hmaster2 & ~n64042;
  assign n64044 = ~n64021 & ~n64043;
  assign n64045 = controllable_hmaster1 & ~n64044;
  assign n64046 = i_hbusreq5 & ~n63821;
  assign n64047 = i_hlock5 & ~n63963;
  assign n64048 = ~i_hlock5 & ~n63988;
  assign n64049 = ~n64047 & ~n64048;
  assign n64050 = ~i_hbusreq5 & ~n64049;
  assign n64051 = ~n64046 & ~n64050;
  assign n64052 = ~controllable_hgrant5 & ~n64051;
  assign n64053 = ~n47071 & ~n64052;
  assign n64054 = controllable_hmaster2 & ~n64053;
  assign n64055 = ~n8378 & ~n34184;
  assign n64056 = ~n62396 & ~n64055;
  assign n64057 = i_hlock5 & ~n64056;
  assign n64058 = ~n8378 & ~n34211;
  assign n64059 = ~n62396 & ~n64058;
  assign n64060 = ~i_hlock5 & ~n64059;
  assign n64061 = ~n64057 & ~n64060;
  assign n64062 = ~i_hbusreq5 & ~n64061;
  assign n64063 = ~n49578 & ~n64062;
  assign n64064 = controllable_hgrant5 & ~n64063;
  assign n64065 = ~n8426 & ~n25342;
  assign n64066 = ~n62405 & ~n64065;
  assign n64067 = ~i_hbusreq9 & ~n64066;
  assign n64068 = ~n49592 & ~n64067;
  assign n64069 = i_hlock4 & ~n64068;
  assign n64070 = ~n8426 & ~n25354;
  assign n64071 = ~n62405 & ~n64070;
  assign n64072 = ~i_hbusreq9 & ~n64071;
  assign n64073 = ~n49599 & ~n64072;
  assign n64074 = ~i_hlock4 & ~n64073;
  assign n64075 = ~n64069 & ~n64074;
  assign n64076 = ~i_hbusreq4 & ~n64075;
  assign n64077 = ~n49591 & ~n64076;
  assign n64078 = controllable_hgrant4 & ~n64077;
  assign n64079 = ~n8365 & ~n25338;
  assign n64080 = ~n62416 & ~n64079;
  assign n64081 = i_hlock3 & ~n64080;
  assign n64082 = ~n8365 & ~n25350;
  assign n64083 = ~n62416 & ~n64082;
  assign n64084 = ~i_hlock3 & ~n64083;
  assign n64085 = ~n64081 & ~n64084;
  assign n64086 = ~i_hbusreq3 & ~n64085;
  assign n64087 = ~n49611 & ~n64086;
  assign n64088 = controllable_hgrant3 & ~n64087;
  assign n64089 = i_hlock1 & ~n46718;
  assign n64090 = ~i_hlock1 & ~n46752;
  assign n64091 = ~n64089 & ~n64090;
  assign n64092 = ~i_hbusreq1 & ~n64091;
  assign n64093 = ~n49637 & ~n64092;
  assign n64094 = ~controllable_hgrant1 & ~n64093;
  assign n64095 = ~n49636 & ~n64094;
  assign n64096 = ~i_hbusreq3 & ~n64095;
  assign n64097 = ~n49623 & ~n64096;
  assign n64098 = ~controllable_hgrant3 & ~n64097;
  assign n64099 = ~n64088 & ~n64098;
  assign n64100 = ~i_hbusreq9 & ~n64099;
  assign n64101 = ~n49610 & ~n64100;
  assign n64102 = ~i_hbusreq4 & ~n64101;
  assign n64103 = ~n49609 & ~n64102;
  assign n64104 = ~controllable_hgrant4 & ~n64103;
  assign n64105 = ~n64078 & ~n64104;
  assign n64106 = ~i_hbusreq5 & ~n64105;
  assign n64107 = ~n49590 & ~n64106;
  assign n64108 = ~controllable_hgrant5 & ~n64107;
  assign n64109 = ~n64064 & ~n64108;
  assign n64110 = ~controllable_hmaster2 & ~n64109;
  assign n64111 = ~n64054 & ~n64110;
  assign n64112 = ~controllable_hmaster1 & ~n64111;
  assign n64113 = ~n64045 & ~n64112;
  assign n64114 = ~i_hbusreq6 & ~n64113;
  assign n64115 = ~n64020 & ~n64114;
  assign n64116 = ~controllable_hgrant6 & ~n64115;
  assign n64117 = ~n64019 & ~n64116;
  assign n64118 = controllable_hmaster0 & ~n64117;
  assign n64119 = i_hbusreq6 & ~n63866;
  assign n64120 = i_hbusreq5 & ~n63835;
  assign n64121 = i_hbusreq4 & ~n63833;
  assign n64122 = i_hbusreq9 & ~n63833;
  assign n64123 = i_hbusreq3 & ~n63831;
  assign n64124 = ~n47265 & ~n62469;
  assign n64125 = ~i_hbusreq3 & ~n64124;
  assign n64126 = ~n64123 & ~n64125;
  assign n64127 = ~controllable_hgrant3 & ~n64126;
  assign n64128 = ~n47225 & ~n64127;
  assign n64129 = ~i_hbusreq9 & ~n64128;
  assign n64130 = ~n64122 & ~n64129;
  assign n64131 = ~i_hbusreq4 & ~n64130;
  assign n64132 = ~n64121 & ~n64131;
  assign n64133 = ~controllable_hgrant4 & ~n64132;
  assign n64134 = ~n47212 & ~n64133;
  assign n64135 = ~i_hbusreq5 & ~n64134;
  assign n64136 = ~n64120 & ~n64135;
  assign n64137 = ~controllable_hgrant5 & ~n64136;
  assign n64138 = ~n47194 & ~n64137;
  assign n64139 = ~controllable_hmaster2 & ~n64138;
  assign n64140 = ~n64021 & ~n64139;
  assign n64141 = controllable_hmaster1 & ~n64140;
  assign n64142 = i_hbusreq5 & ~n63845;
  assign n64143 = i_hbusreq4 & ~n63843;
  assign n64144 = i_hlock4 & ~n63959;
  assign n64145 = ~i_hlock4 & ~n63984;
  assign n64146 = ~n64144 & ~n64145;
  assign n64147 = ~i_hbusreq4 & ~n64146;
  assign n64148 = ~n64143 & ~n64147;
  assign n64149 = ~controllable_hgrant4 & ~n64148;
  assign n64150 = ~n47312 & ~n64149;
  assign n64151 = ~i_hbusreq5 & ~n64150;
  assign n64152 = ~n64142 & ~n64151;
  assign n64153 = ~controllable_hgrant5 & ~n64152;
  assign n64154 = ~n47294 & ~n64153;
  assign n64155 = controllable_hmaster2 & ~n64154;
  assign n64156 = i_hbusreq5 & ~n63853;
  assign n64157 = i_hbusreq4 & ~n63851;
  assign n64158 = i_hbusreq9 & ~n63851;
  assign n64159 = i_hbusreq3 & ~n63849;
  assign n64160 = ~n47402 & ~n62516;
  assign n64161 = ~i_hbusreq3 & ~n64160;
  assign n64162 = ~n64159 & ~n64161;
  assign n64163 = ~controllable_hgrant3 & ~n64162;
  assign n64164 = ~n47367 & ~n64163;
  assign n64165 = ~i_hbusreq9 & ~n64164;
  assign n64166 = ~n64158 & ~n64165;
  assign n64167 = ~i_hbusreq4 & ~n64166;
  assign n64168 = ~n64157 & ~n64167;
  assign n64169 = ~controllable_hgrant4 & ~n64168;
  assign n64170 = ~n47354 & ~n64169;
  assign n64171 = ~i_hbusreq5 & ~n64170;
  assign n64172 = ~n64156 & ~n64171;
  assign n64173 = ~controllable_hgrant5 & ~n64172;
  assign n64174 = ~n47336 & ~n64173;
  assign n64175 = ~controllable_hmaster2 & ~n64174;
  assign n64176 = ~n64155 & ~n64175;
  assign n64177 = ~controllable_hmaster1 & ~n64176;
  assign n64178 = ~n64141 & ~n64177;
  assign n64179 = i_hlock6 & ~n64178;
  assign n64180 = controllable_hmaster2 & ~n63992;
  assign n64181 = ~n64139 & ~n64180;
  assign n64182 = controllable_hmaster1 & ~n64181;
  assign n64183 = ~n64177 & ~n64182;
  assign n64184 = ~i_hlock6 & ~n64183;
  assign n64185 = ~n64179 & ~n64184;
  assign n64186 = ~i_hbusreq6 & ~n64185;
  assign n64187 = ~n64119 & ~n64186;
  assign n64188 = ~controllable_hgrant6 & ~n64187;
  assign n64189 = ~n47182 & ~n64188;
  assign n64190 = ~controllable_hmaster0 & ~n64189;
  assign n64191 = ~n64118 & ~n64190;
  assign n64192 = ~i_hbusreq8 & ~n64191;
  assign n64193 = ~n64008 & ~n64192;
  assign n64194 = ~controllable_hmaster3 & ~n64193;
  assign n64195 = ~n64007 & ~n64194;
  assign n64196 = i_hlock7 & ~n64195;
  assign n64197 = i_hbusreq8 & ~n63888;
  assign n64198 = i_hbusreq6 & ~n63880;
  assign n64199 = ~n8217 & ~n38811;
  assign n64200 = ~n62556 & ~n64199;
  assign n64201 = i_hlock6 & ~n64200;
  assign n64202 = ~n8217 & ~n38820;
  assign n64203 = ~n62556 & ~n64202;
  assign n64204 = ~i_hlock6 & ~n64203;
  assign n64205 = ~n64201 & ~n64204;
  assign n64206 = ~i_hbusreq6 & ~n64205;
  assign n64207 = ~n64198 & ~n64206;
  assign n64208 = controllable_hgrant6 & ~n64207;
  assign n64209 = i_hbusreq6 & ~n63884;
  assign n64210 = ~n64043 & ~n64180;
  assign n64211 = controllable_hmaster1 & ~n64210;
  assign n64212 = ~n64112 & ~n64211;
  assign n64213 = ~i_hbusreq6 & ~n64212;
  assign n64214 = ~n64209 & ~n64213;
  assign n64215 = ~controllable_hgrant6 & ~n64214;
  assign n64216 = ~n64208 & ~n64215;
  assign n64217 = controllable_hmaster0 & ~n64216;
  assign n64218 = ~n64190 & ~n64217;
  assign n64219 = ~i_hbusreq8 & ~n64218;
  assign n64220 = ~n64197 & ~n64219;
  assign n64221 = ~controllable_hmaster3 & ~n64220;
  assign n64222 = ~n64007 & ~n64221;
  assign n64223 = ~i_hlock7 & ~n64222;
  assign n64224 = ~n64196 & ~n64223;
  assign n64225 = ~i_hbusreq7 & ~n64224;
  assign n64226 = ~n63893 & ~n64225;
  assign n64227 = n7924 & ~n64226;
  assign n64228 = ~n62040 & ~n64227;
  assign n64229 = ~n8214 & ~n64228;
  assign n64230 = ~n34238 & ~n46336;
  assign n64231 = ~n8217 & ~n64230;
  assign n64232 = ~n43999 & ~n64231;
  assign n64233 = i_hlock6 & ~n64232;
  assign n64234 = ~n34252 & ~n46342;
  assign n64235 = ~n8217 & ~n64234;
  assign n64236 = ~n44009 & ~n64235;
  assign n64237 = ~i_hlock6 & ~n64236;
  assign n64238 = ~n64233 & ~n64237;
  assign n64239 = controllable_hgrant6 & ~n64238;
  assign n64240 = ~n46432 & ~n49059;
  assign n64241 = ~controllable_hmaster1 & ~n64240;
  assign n64242 = ~n46408 & ~n64241;
  assign n64243 = i_hlock6 & ~n64242;
  assign n64244 = ~n46481 & ~n64241;
  assign n64245 = ~i_hlock6 & ~n64244;
  assign n64246 = ~n64243 & ~n64245;
  assign n64247 = ~controllable_hgrant6 & ~n64246;
  assign n64248 = ~n64239 & ~n64247;
  assign n64249 = ~controllable_hmaster0 & ~n64248;
  assign n64250 = ~n46334 & ~n64249;
  assign n64251 = ~controllable_hmaster3 & ~n64250;
  assign n64252 = ~n47796 & ~n64251;
  assign n64253 = i_hlock7 & ~n64252;
  assign n64254 = ~n46505 & ~n64249;
  assign n64255 = ~controllable_hmaster3 & ~n64254;
  assign n64256 = ~n47796 & ~n64255;
  assign n64257 = ~i_hlock7 & ~n64256;
  assign n64258 = ~n64253 & ~n64257;
  assign n64259 = i_hbusreq7 & ~n64258;
  assign n64260 = ~n8217 & ~n34294;
  assign n64261 = ~n49089 & ~n64260;
  assign n64262 = i_hlock6 & ~n64261;
  assign n64263 = ~n8217 & ~n34473;
  assign n64264 = ~n49089 & ~n64263;
  assign n64265 = ~i_hlock6 & ~n64264;
  assign n64266 = ~n64262 & ~n64265;
  assign n64267 = ~i_hbusreq6 & ~n64266;
  assign n64268 = ~n47588 & ~n64267;
  assign n64269 = controllable_hgrant6 & ~n64268;
  assign n64270 = ~n8378 & ~n34272;
  assign n64271 = ~n49102 & ~n64270;
  assign n64272 = i_hlock5 & ~n64271;
  assign n64273 = ~n8378 & ~n34451;
  assign n64274 = ~n49102 & ~n64273;
  assign n64275 = ~i_hlock5 & ~n64274;
  assign n64276 = ~n64272 & ~n64275;
  assign n64277 = ~i_hbusreq5 & ~n64276;
  assign n64278 = ~n46525 & ~n64277;
  assign n64279 = controllable_hgrant5 & ~n64278;
  assign n64280 = ~n8426 & ~n25444;
  assign n64281 = ~n49116 & ~n64280;
  assign n64282 = ~i_hbusreq9 & ~n64281;
  assign n64283 = ~n46538 & ~n64282;
  assign n64284 = i_hlock4 & ~n64283;
  assign n64285 = ~n8426 & ~n25462;
  assign n64286 = ~n49116 & ~n64285;
  assign n64287 = ~i_hbusreq9 & ~n64286;
  assign n64288 = ~n46544 & ~n64287;
  assign n64289 = ~i_hlock4 & ~n64288;
  assign n64290 = ~n64284 & ~n64289;
  assign n64291 = ~i_hbusreq4 & ~n64290;
  assign n64292 = ~n46537 & ~n64291;
  assign n64293 = controllable_hgrant4 & ~n64292;
  assign n64294 = ~n8365 & ~n25440;
  assign n64295 = ~n49135 & ~n64294;
  assign n64296 = i_hlock3 & ~n64295;
  assign n64297 = ~n8365 & ~n25458;
  assign n64298 = ~n49135 & ~n64297;
  assign n64299 = ~i_hlock3 & ~n64298;
  assign n64300 = ~n64296 & ~n64299;
  assign n64301 = ~i_hbusreq3 & ~n64300;
  assign n64302 = ~n46556 & ~n64301;
  assign n64303 = controllable_hgrant3 & ~n64302;
  assign n64304 = ~n8389 & ~n25436;
  assign n64305 = ~n49148 & ~n64304;
  assign n64306 = i_hlock1 & ~n64305;
  assign n64307 = ~n8389 & ~n25454;
  assign n64308 = ~n49148 & ~n64307;
  assign n64309 = ~i_hlock1 & ~n64308;
  assign n64310 = ~n64306 & ~n64309;
  assign n64311 = ~i_hbusreq1 & ~n64310;
  assign n64312 = ~n46568 & ~n64311;
  assign n64313 = controllable_hgrant1 & ~n64312;
  assign n64314 = ~n46386 & ~n46690;
  assign n64315 = controllable_locked & ~n64314;
  assign n64316 = ~n49183 & ~n64315;
  assign n64317 = i_hlock0 & ~n64316;
  assign n64318 = ~n46586 & ~n64317;
  assign n64319 = ~i_hbusreq0 & ~n64318;
  assign n64320 = ~n46581 & ~n64319;
  assign n64321 = i_hlock2 & ~n64320;
  assign n64322 = ~n46591 & ~n64319;
  assign n64323 = ~i_hlock2 & ~n64322;
  assign n64324 = ~n64321 & ~n64323;
  assign n64325 = ~i_hbusreq2 & ~n64324;
  assign n64326 = ~n46580 & ~n64325;
  assign n64327 = controllable_hgrant2 & ~n64326;
  assign n64328 = ~n25486 & ~n64327;
  assign n64329 = n7733 & ~n64328;
  assign n64330 = ~n63196 & ~n64329;
  assign n64331 = n7928 & ~n64330;
  assign n64332 = ~n62652 & ~n64331;
  assign n64333 = ~i_hbusreq1 & ~n64332;
  assign n64334 = ~n46579 & ~n64333;
  assign n64335 = ~controllable_hgrant1 & ~n64334;
  assign n64336 = ~n64313 & ~n64335;
  assign n64337 = ~i_hbusreq3 & ~n64336;
  assign n64338 = ~n46567 & ~n64337;
  assign n64339 = ~controllable_hgrant3 & ~n64338;
  assign n64340 = ~n64303 & ~n64339;
  assign n64341 = ~i_hbusreq9 & ~n64340;
  assign n64342 = ~n46555 & ~n64341;
  assign n64343 = ~i_hbusreq4 & ~n64342;
  assign n64344 = ~n46554 & ~n64343;
  assign n64345 = ~controllable_hgrant4 & ~n64344;
  assign n64346 = ~n64293 & ~n64345;
  assign n64347 = ~i_hbusreq5 & ~n64346;
  assign n64348 = ~n46536 & ~n64347;
  assign n64349 = ~controllable_hgrant5 & ~n64348;
  assign n64350 = ~n64279 & ~n64349;
  assign n64351 = controllable_hmaster1 & ~n64350;
  assign n64352 = controllable_hmaster2 & ~n64350;
  assign n64353 = ~n8378 & ~n34286;
  assign n64354 = ~n49221 & ~n64353;
  assign n64355 = i_hlock5 & ~n64354;
  assign n64356 = ~n8378 & ~n34465;
  assign n64357 = ~n49221 & ~n64356;
  assign n64358 = ~i_hlock5 & ~n64357;
  assign n64359 = ~n64355 & ~n64358;
  assign n64360 = ~i_hbusreq5 & ~n64359;
  assign n64361 = ~n47600 & ~n64360;
  assign n64362 = controllable_hgrant5 & ~n64361;
  assign n64363 = ~n8426 & ~n25549;
  assign n64364 = ~n49232 & ~n64363;
  assign n64365 = i_hlock9 & ~n64364;
  assign n64366 = ~n8426 & ~n25593;
  assign n64367 = ~n49236 & ~n64366;
  assign n64368 = ~i_hlock9 & ~n64367;
  assign n64369 = ~n64365 & ~n64368;
  assign n64370 = ~i_hbusreq9 & ~n64369;
  assign n64371 = ~n47613 & ~n64370;
  assign n64372 = i_hlock4 & ~n64371;
  assign n64373 = ~n8426 & ~n25561;
  assign n64374 = ~n49232 & ~n64373;
  assign n64375 = i_hlock9 & ~n64374;
  assign n64376 = ~n8426 & ~n25603;
  assign n64377 = ~n49236 & ~n64376;
  assign n64378 = ~i_hlock9 & ~n64377;
  assign n64379 = ~n64375 & ~n64378;
  assign n64380 = ~i_hbusreq9 & ~n64379;
  assign n64381 = ~n47620 & ~n64380;
  assign n64382 = ~i_hlock4 & ~n64381;
  assign n64383 = ~n64372 & ~n64382;
  assign n64384 = ~i_hbusreq4 & ~n64383;
  assign n64385 = ~n47612 & ~n64384;
  assign n64386 = controllable_hgrant4 & ~n64385;
  assign n64387 = ~n8365 & ~n25545;
  assign n64388 = ~n49258 & ~n64387;
  assign n64389 = i_hlock3 & ~n64388;
  assign n64390 = ~n8365 & ~n25557;
  assign n64391 = ~n49258 & ~n64390;
  assign n64392 = ~i_hlock3 & ~n64391;
  assign n64393 = ~n64389 & ~n64392;
  assign n64394 = ~i_hbusreq3 & ~n64393;
  assign n64395 = ~n46825 & ~n64394;
  assign n64396 = controllable_hgrant3 & ~n64395;
  assign n64397 = ~n8389 & ~n25541;
  assign n64398 = ~n49269 & ~n64397;
  assign n64399 = i_hlock1 & ~n64398;
  assign n64400 = ~n8389 & ~n25553;
  assign n64401 = ~n49269 & ~n64400;
  assign n64402 = ~i_hlock1 & ~n64401;
  assign n64403 = ~n64399 & ~n64402;
  assign n64404 = ~i_hbusreq1 & ~n64403;
  assign n64405 = ~n46837 & ~n64404;
  assign n64406 = controllable_hgrant1 & ~n64405;
  assign n64407 = ~n25431 & ~n64327;
  assign n64408 = n7733 & ~n64407;
  assign n64409 = ~n63266 & ~n64408;
  assign n64410 = n7928 & ~n64409;
  assign n64411 = ~n8265 & ~n64410;
  assign n64412 = ~i_hbusreq1 & ~n64411;
  assign n64413 = ~n46848 & ~n64412;
  assign n64414 = ~controllable_hgrant1 & ~n64413;
  assign n64415 = ~n64406 & ~n64414;
  assign n64416 = ~i_hbusreq3 & ~n64415;
  assign n64417 = ~n46836 & ~n64416;
  assign n64418 = ~controllable_hgrant3 & ~n64417;
  assign n64419 = ~n64396 & ~n64418;
  assign n64420 = i_hlock9 & ~n64419;
  assign n64421 = ~n8365 & ~n25589;
  assign n64422 = ~n49311 & ~n64421;
  assign n64423 = i_hlock3 & ~n64422;
  assign n64424 = ~n8365 & ~n25599;
  assign n64425 = ~n49311 & ~n64424;
  assign n64426 = ~i_hlock3 & ~n64425;
  assign n64427 = ~n64423 & ~n64426;
  assign n64428 = ~i_hbusreq3 & ~n64427;
  assign n64429 = ~n46926 & ~n64428;
  assign n64430 = controllable_hgrant3 & ~n64429;
  assign n64431 = ~n8389 & ~n25585;
  assign n64432 = ~n49322 & ~n64431;
  assign n64433 = i_hlock1 & ~n64432;
  assign n64434 = ~n8389 & ~n25595;
  assign n64435 = ~n49322 & ~n64434;
  assign n64436 = ~i_hlock1 & ~n64435;
  assign n64437 = ~n64433 & ~n64436;
  assign n64438 = ~i_hbusreq1 & ~n64437;
  assign n64439 = ~n46938 & ~n64438;
  assign n64440 = controllable_hgrant1 & ~n64439;
  assign n64441 = ~n8297 & ~n64410;
  assign n64442 = ~i_hbusreq1 & ~n64441;
  assign n64443 = ~n46949 & ~n64442;
  assign n64444 = ~controllable_hgrant1 & ~n64443;
  assign n64445 = ~n64440 & ~n64444;
  assign n64446 = ~i_hbusreq3 & ~n64445;
  assign n64447 = ~n46937 & ~n64446;
  assign n64448 = ~controllable_hgrant3 & ~n64447;
  assign n64449 = ~n64430 & ~n64448;
  assign n64450 = ~i_hlock9 & ~n64449;
  assign n64451 = ~n64420 & ~n64450;
  assign n64452 = ~i_hbusreq9 & ~n64451;
  assign n64453 = ~n47632 & ~n64452;
  assign n64454 = ~i_hbusreq4 & ~n64453;
  assign n64455 = ~n47631 & ~n64454;
  assign n64456 = ~controllable_hgrant4 & ~n64455;
  assign n64457 = ~n64386 & ~n64456;
  assign n64458 = ~i_hbusreq5 & ~n64457;
  assign n64459 = ~n47611 & ~n64458;
  assign n64460 = ~controllable_hgrant5 & ~n64459;
  assign n64461 = ~n64362 & ~n64460;
  assign n64462 = ~controllable_hmaster2 & ~n64461;
  assign n64463 = ~n64352 & ~n64462;
  assign n64464 = ~controllable_hmaster1 & ~n64463;
  assign n64465 = ~n64351 & ~n64464;
  assign n64466 = ~i_hbusreq6 & ~n64465;
  assign n64467 = ~n47599 & ~n64466;
  assign n64468 = ~controllable_hgrant6 & ~n64467;
  assign n64469 = ~n64269 & ~n64468;
  assign n64470 = controllable_hmaster0 & ~n64469;
  assign n64471 = ~n8217 & ~n34313;
  assign n64472 = ~n49363 & ~n64471;
  assign n64473 = i_hlock6 & ~n64472;
  assign n64474 = ~n8217 & ~n34492;
  assign n64475 = ~n49363 & ~n64474;
  assign n64476 = ~i_hlock6 & ~n64475;
  assign n64477 = ~n64473 & ~n64476;
  assign n64478 = ~i_hbusreq6 & ~n64477;
  assign n64479 = ~n46782 & ~n64478;
  assign n64480 = controllable_hgrant6 & ~n64479;
  assign n64481 = ~n8378 & ~n34305;
  assign n64482 = ~n49375 & ~n64481;
  assign n64483 = i_hlock5 & ~n64482;
  assign n64484 = ~n8378 & ~n34484;
  assign n64485 = ~n49375 & ~n64484;
  assign n64486 = ~i_hlock5 & ~n64485;
  assign n64487 = ~n64483 & ~n64486;
  assign n64488 = ~i_hbusreq5 & ~n64487;
  assign n64489 = ~n46794 & ~n64488;
  assign n64490 = controllable_hgrant5 & ~n64489;
  assign n64491 = ~i_hbusreq9 & ~n64364;
  assign n64492 = ~n46807 & ~n64491;
  assign n64493 = i_hlock4 & ~n64492;
  assign n64494 = ~i_hbusreq9 & ~n64374;
  assign n64495 = ~n46813 & ~n64494;
  assign n64496 = ~i_hlock4 & ~n64495;
  assign n64497 = ~n64493 & ~n64496;
  assign n64498 = ~i_hbusreq4 & ~n64497;
  assign n64499 = ~n46806 & ~n64498;
  assign n64500 = controllable_hgrant4 & ~n64499;
  assign n64501 = ~i_hbusreq9 & ~n64419;
  assign n64502 = ~n46824 & ~n64501;
  assign n64503 = ~i_hbusreq4 & ~n64502;
  assign n64504 = ~n46823 & ~n64503;
  assign n64505 = ~controllable_hgrant4 & ~n64504;
  assign n64506 = ~n64500 & ~n64505;
  assign n64507 = ~i_hbusreq5 & ~n64506;
  assign n64508 = ~n46805 & ~n64507;
  assign n64509 = ~controllable_hgrant5 & ~n64508;
  assign n64510 = ~n64490 & ~n64509;
  assign n64511 = ~controllable_hmaster2 & ~n64510;
  assign n64512 = ~n64352 & ~n64511;
  assign n64513 = ~controllable_hmaster1 & ~n64512;
  assign n64514 = ~n64351 & ~n64513;
  assign n64515 = ~i_hbusreq6 & ~n64514;
  assign n64516 = ~n46793 & ~n64515;
  assign n64517 = ~controllable_hgrant6 & ~n64516;
  assign n64518 = ~n64480 & ~n64517;
  assign n64519 = ~controllable_hmaster0 & ~n64518;
  assign n64520 = ~n64470 & ~n64519;
  assign n64521 = i_hlock8 & ~n64520;
  assign n64522 = ~n8217 & ~n34334;
  assign n64523 = ~n49417 & ~n64522;
  assign n64524 = i_hlock6 & ~n64523;
  assign n64525 = ~n8217 & ~n34513;
  assign n64526 = ~n49417 & ~n64525;
  assign n64527 = ~i_hlock6 & ~n64526;
  assign n64528 = ~n64524 & ~n64527;
  assign n64529 = ~i_hbusreq6 & ~n64528;
  assign n64530 = ~n46883 & ~n64529;
  assign n64531 = controllable_hgrant6 & ~n64530;
  assign n64532 = ~n8378 & ~n34326;
  assign n64533 = ~n49429 & ~n64532;
  assign n64534 = i_hlock5 & ~n64533;
  assign n64535 = ~n8378 & ~n34505;
  assign n64536 = ~n49429 & ~n64535;
  assign n64537 = ~i_hlock5 & ~n64536;
  assign n64538 = ~n64534 & ~n64537;
  assign n64539 = ~i_hbusreq5 & ~n64538;
  assign n64540 = ~n46895 & ~n64539;
  assign n64541 = controllable_hgrant5 & ~n64540;
  assign n64542 = ~i_hbusreq9 & ~n64367;
  assign n64543 = ~n46908 & ~n64542;
  assign n64544 = i_hlock4 & ~n64543;
  assign n64545 = ~i_hbusreq9 & ~n64377;
  assign n64546 = ~n46914 & ~n64545;
  assign n64547 = ~i_hlock4 & ~n64546;
  assign n64548 = ~n64544 & ~n64547;
  assign n64549 = ~i_hbusreq4 & ~n64548;
  assign n64550 = ~n46907 & ~n64549;
  assign n64551 = controllable_hgrant4 & ~n64550;
  assign n64552 = ~i_hbusreq9 & ~n64449;
  assign n64553 = ~n46925 & ~n64552;
  assign n64554 = ~i_hbusreq4 & ~n64553;
  assign n64555 = ~n46924 & ~n64554;
  assign n64556 = ~controllable_hgrant4 & ~n64555;
  assign n64557 = ~n64551 & ~n64556;
  assign n64558 = ~i_hbusreq5 & ~n64557;
  assign n64559 = ~n46906 & ~n64558;
  assign n64560 = ~controllable_hgrant5 & ~n64559;
  assign n64561 = ~n64541 & ~n64560;
  assign n64562 = ~controllable_hmaster2 & ~n64561;
  assign n64563 = ~n64352 & ~n64562;
  assign n64564 = ~controllable_hmaster1 & ~n64563;
  assign n64565 = ~n64351 & ~n64564;
  assign n64566 = ~i_hbusreq6 & ~n64565;
  assign n64567 = ~n46894 & ~n64566;
  assign n64568 = ~controllable_hgrant6 & ~n64567;
  assign n64569 = ~n64531 & ~n64568;
  assign n64570 = ~controllable_hmaster0 & ~n64569;
  assign n64571 = ~n64470 & ~n64570;
  assign n64572 = ~i_hlock8 & ~n64571;
  assign n64573 = ~n64521 & ~n64572;
  assign n64574 = ~i_hbusreq8 & ~n64573;
  assign n64575 = ~n47837 & ~n64574;
  assign n64576 = controllable_hmaster3 & ~n64575;
  assign n64577 = i_hbusreq8 & ~n64250;
  assign n64578 = ~n8217 & ~n38887;
  assign n64579 = ~n49476 & ~n64578;
  assign n64580 = i_hlock6 & ~n64579;
  assign n64581 = ~n8217 & ~n38897;
  assign n64582 = ~n49476 & ~n64581;
  assign n64583 = ~i_hlock6 & ~n64582;
  assign n64584 = ~n64580 & ~n64583;
  assign n64585 = ~i_hbusreq6 & ~n64584;
  assign n64586 = ~n46985 & ~n64585;
  assign n64587 = controllable_hgrant6 & ~n64586;
  assign n64588 = controllable_hmaster2 & ~n64510;
  assign n64589 = ~n8378 & ~n34363;
  assign n64590 = ~n49490 & ~n64589;
  assign n64591 = i_hlock5 & ~n64590;
  assign n64592 = ~n8378 & ~n34542;
  assign n64593 = ~n49490 & ~n64592;
  assign n64594 = ~i_hlock5 & ~n64593;
  assign n64595 = ~n64591 & ~n64594;
  assign n64596 = ~i_hbusreq5 & ~n64595;
  assign n64597 = ~n46998 & ~n64596;
  assign n64598 = controllable_hgrant5 & ~n64597;
  assign n64599 = ~n8426 & ~n25639;
  assign n64600 = ~n49504 & ~n64599;
  assign n64601 = ~i_hbusreq9 & ~n64600;
  assign n64602 = ~n47011 & ~n64601;
  assign n64603 = i_hlock4 & ~n64602;
  assign n64604 = ~n8426 & ~n25647;
  assign n64605 = ~n49504 & ~n64604;
  assign n64606 = ~i_hbusreq9 & ~n64605;
  assign n64607 = ~n47017 & ~n64606;
  assign n64608 = ~i_hlock4 & ~n64607;
  assign n64609 = ~n64603 & ~n64608;
  assign n64610 = ~i_hbusreq4 & ~n64609;
  assign n64611 = ~n47010 & ~n64610;
  assign n64612 = controllable_hgrant4 & ~n64611;
  assign n64613 = ~n8365 & ~n25495;
  assign n64614 = ~n49523 & ~n64613;
  assign n64615 = i_hlock3 & ~n64614;
  assign n64616 = ~n8365 & ~n25513;
  assign n64617 = ~n49527 & ~n64616;
  assign n64618 = ~i_hlock3 & ~n64617;
  assign n64619 = ~n64615 & ~n64618;
  assign n64620 = ~i_hbusreq3 & ~n64619;
  assign n64621 = ~n47029 & ~n64620;
  assign n64622 = controllable_hgrant3 & ~n64621;
  assign n64623 = i_hlock3 & ~n64415;
  assign n64624 = ~i_hlock3 & ~n64445;
  assign n64625 = ~n64623 & ~n64624;
  assign n64626 = ~i_hbusreq3 & ~n64625;
  assign n64627 = ~n47040 & ~n64626;
  assign n64628 = ~controllable_hgrant3 & ~n64627;
  assign n64629 = ~n64622 & ~n64628;
  assign n64630 = ~i_hbusreq9 & ~n64629;
  assign n64631 = ~n47028 & ~n64630;
  assign n64632 = ~i_hbusreq4 & ~n64631;
  assign n64633 = ~n47027 & ~n64632;
  assign n64634 = ~controllable_hgrant4 & ~n64633;
  assign n64635 = ~n64612 & ~n64634;
  assign n64636 = ~i_hbusreq5 & ~n64635;
  assign n64637 = ~n47009 & ~n64636;
  assign n64638 = ~controllable_hgrant5 & ~n64637;
  assign n64639 = ~n64598 & ~n64638;
  assign n64640 = ~controllable_hmaster2 & ~n64639;
  assign n64641 = ~n64588 & ~n64640;
  assign n64642 = controllable_hmaster1 & ~n64641;
  assign n64643 = ~n8378 & ~n34352;
  assign n64644 = ~n49557 & ~n64643;
  assign n64645 = i_hlock5 & ~n64644;
  assign n64646 = ~n8378 & ~n34531;
  assign n64647 = ~n49561 & ~n64646;
  assign n64648 = ~i_hlock5 & ~n64647;
  assign n64649 = ~n64645 & ~n64648;
  assign n64650 = ~i_hbusreq5 & ~n64649;
  assign n64651 = ~n47061 & ~n64650;
  assign n64652 = controllable_hgrant5 & ~n64651;
  assign n64653 = i_hlock5 & ~n64506;
  assign n64654 = ~i_hlock5 & ~n64557;
  assign n64655 = ~n64653 & ~n64654;
  assign n64656 = ~i_hbusreq5 & ~n64655;
  assign n64657 = ~n47072 & ~n64656;
  assign n64658 = ~controllable_hgrant5 & ~n64657;
  assign n64659 = ~n64652 & ~n64658;
  assign n64660 = controllable_hmaster2 & ~n64659;
  assign n64661 = ~n8378 & ~n34384;
  assign n64662 = ~n49579 & ~n64661;
  assign n64663 = i_hlock5 & ~n64662;
  assign n64664 = ~n8378 & ~n34563;
  assign n64665 = ~n49579 & ~n64664;
  assign n64666 = ~i_hlock5 & ~n64665;
  assign n64667 = ~n64663 & ~n64666;
  assign n64668 = ~i_hbusreq5 & ~n64667;
  assign n64669 = ~n47081 & ~n64668;
  assign n64670 = controllable_hgrant5 & ~n64669;
  assign n64671 = ~n8426 & ~n25681;
  assign n64672 = ~n49593 & ~n64671;
  assign n64673 = ~i_hbusreq9 & ~n64672;
  assign n64674 = ~n47094 & ~n64673;
  assign n64675 = i_hlock4 & ~n64674;
  assign n64676 = ~n8426 & ~n25693;
  assign n64677 = ~n49593 & ~n64676;
  assign n64678 = ~i_hbusreq9 & ~n64677;
  assign n64679 = ~n47100 & ~n64678;
  assign n64680 = ~i_hlock4 & ~n64679;
  assign n64681 = ~n64675 & ~n64680;
  assign n64682 = ~i_hbusreq4 & ~n64681;
  assign n64683 = ~n47093 & ~n64682;
  assign n64684 = controllable_hgrant4 & ~n64683;
  assign n64685 = ~n8365 & ~n25677;
  assign n64686 = ~n49612 & ~n64685;
  assign n64687 = i_hlock3 & ~n64686;
  assign n64688 = ~n8365 & ~n25689;
  assign n64689 = ~n49612 & ~n64688;
  assign n64690 = ~i_hlock3 & ~n64689;
  assign n64691 = ~n64687 & ~n64690;
  assign n64692 = ~i_hbusreq3 & ~n64691;
  assign n64693 = ~n47112 & ~n64692;
  assign n64694 = controllable_hgrant3 & ~n64693;
  assign n64695 = ~n8389 & ~n25491;
  assign n64696 = ~n49625 & ~n64695;
  assign n64697 = i_hlock1 & ~n64696;
  assign n64698 = ~n8389 & ~n25509;
  assign n64699 = ~n49629 & ~n64698;
  assign n64700 = ~i_hlock1 & ~n64699;
  assign n64701 = ~n64697 & ~n64700;
  assign n64702 = ~i_hbusreq1 & ~n64701;
  assign n64703 = ~n47124 & ~n64702;
  assign n64704 = controllable_hgrant1 & ~n64703;
  assign n64705 = i_hlock1 & ~n64411;
  assign n64706 = ~i_hlock1 & ~n64441;
  assign n64707 = ~n64705 & ~n64706;
  assign n64708 = ~i_hbusreq1 & ~n64707;
  assign n64709 = ~n47135 & ~n64708;
  assign n64710 = ~controllable_hgrant1 & ~n64709;
  assign n64711 = ~n64704 & ~n64710;
  assign n64712 = ~i_hbusreq3 & ~n64711;
  assign n64713 = ~n47123 & ~n64712;
  assign n64714 = ~controllable_hgrant3 & ~n64713;
  assign n64715 = ~n64694 & ~n64714;
  assign n64716 = ~i_hbusreq9 & ~n64715;
  assign n64717 = ~n47111 & ~n64716;
  assign n64718 = ~i_hbusreq4 & ~n64717;
  assign n64719 = ~n47110 & ~n64718;
  assign n64720 = ~controllable_hgrant4 & ~n64719;
  assign n64721 = ~n64684 & ~n64720;
  assign n64722 = ~i_hbusreq5 & ~n64721;
  assign n64723 = ~n47092 & ~n64722;
  assign n64724 = ~controllable_hgrant5 & ~n64723;
  assign n64725 = ~n64670 & ~n64724;
  assign n64726 = ~controllable_hmaster2 & ~n64725;
  assign n64727 = ~n64660 & ~n64726;
  assign n64728 = ~controllable_hmaster1 & ~n64727;
  assign n64729 = ~n64642 & ~n64728;
  assign n64730 = ~i_hbusreq6 & ~n64729;
  assign n64731 = ~n46996 & ~n64730;
  assign n64732 = ~controllable_hgrant6 & ~n64731;
  assign n64733 = ~n64587 & ~n64732;
  assign n64734 = controllable_hmaster0 & ~n64733;
  assign n64735 = i_hbusreq6 & ~n64238;
  assign n64736 = ~n34357 & ~n34410;
  assign n64737 = controllable_hmaster1 & ~n64736;
  assign n64738 = ~n34426 & ~n64737;
  assign n64739 = ~n8217 & ~n64738;
  assign n64740 = ~n49671 & ~n64739;
  assign n64741 = i_hlock6 & ~n64740;
  assign n64742 = ~n34536 & ~n34589;
  assign n64743 = controllable_hmaster1 & ~n64742;
  assign n64744 = ~n34605 & ~n64743;
  assign n64745 = ~n8217 & ~n64744;
  assign n64746 = ~n49681 & ~n64745;
  assign n64747 = ~i_hlock6 & ~n64746;
  assign n64748 = ~n64741 & ~n64747;
  assign n64749 = ~i_hbusreq6 & ~n64748;
  assign n64750 = ~n64735 & ~n64749;
  assign n64751 = controllable_hgrant6 & ~n64750;
  assign n64752 = i_hbusreq6 & ~n64246;
  assign n64753 = ~n8378 & ~n34405;
  assign n64754 = ~n49694 & ~n64753;
  assign n64755 = i_hlock5 & ~n64754;
  assign n64756 = ~n8378 & ~n34584;
  assign n64757 = ~n49694 & ~n64756;
  assign n64758 = ~i_hlock5 & ~n64757;
  assign n64759 = ~n64755 & ~n64758;
  assign n64760 = ~i_hbusreq5 & ~n64759;
  assign n64761 = ~n47184 & ~n64760;
  assign n64762 = controllable_hgrant5 & ~n64761;
  assign n64763 = ~n8426 & ~n25724;
  assign n64764 = ~n49708 & ~n64763;
  assign n64765 = ~i_hbusreq9 & ~n64764;
  assign n64766 = ~n47197 & ~n64765;
  assign n64767 = i_hlock4 & ~n64766;
  assign n64768 = ~n8426 & ~n25734;
  assign n64769 = ~n49708 & ~n64768;
  assign n64770 = ~i_hbusreq9 & ~n64769;
  assign n64771 = ~n47203 & ~n64770;
  assign n64772 = ~i_hlock4 & ~n64771;
  assign n64773 = ~n64767 & ~n64772;
  assign n64774 = ~i_hbusreq4 & ~n64773;
  assign n64775 = ~n47196 & ~n64774;
  assign n64776 = controllable_hgrant4 & ~n64775;
  assign n64777 = ~n8365 & ~n25720;
  assign n64778 = ~n49727 & ~n64777;
  assign n64779 = i_hlock3 & ~n64778;
  assign n64780 = ~n8365 & ~n25730;
  assign n64781 = ~n49727 & ~n64780;
  assign n64782 = ~i_hlock3 & ~n64781;
  assign n64783 = ~n64779 & ~n64782;
  assign n64784 = ~i_hbusreq3 & ~n64783;
  assign n64785 = ~n47215 & ~n64784;
  assign n64786 = controllable_hgrant3 & ~n64785;
  assign n64787 = ~n8389 & ~n25716;
  assign n64788 = ~n49740 & ~n64787;
  assign n64789 = i_hlock1 & ~n64788;
  assign n64790 = ~n8389 & ~n25726;
  assign n64791 = ~n49740 & ~n64790;
  assign n64792 = ~i_hlock1 & ~n64791;
  assign n64793 = ~n64789 & ~n64792;
  assign n64794 = ~i_hbusreq1 & ~n64793;
  assign n64795 = ~n47227 & ~n64794;
  assign n64796 = controllable_hgrant1 & ~n64795;
  assign n64797 = ~n39853 & ~n46386;
  assign n64798 = controllable_locked & ~n64797;
  assign n64799 = ~n49183 & ~n64798;
  assign n64800 = i_hlock0 & ~n64799;
  assign n64801 = ~n47246 & ~n64800;
  assign n64802 = ~i_hbusreq0 & ~n64801;
  assign n64803 = ~n47240 & ~n64802;
  assign n64804 = i_hlock2 & ~n64803;
  assign n64805 = ~n47251 & ~n64802;
  assign n64806 = ~i_hlock2 & ~n64805;
  assign n64807 = ~n64804 & ~n64806;
  assign n64808 = ~i_hbusreq2 & ~n64807;
  assign n64809 = ~n47239 & ~n64808;
  assign n64810 = controllable_hgrant2 & ~n64809;
  assign n64811 = ~n25431 & ~n64810;
  assign n64812 = n7733 & ~n64811;
  assign n64813 = ~n63562 & ~n64812;
  assign n64814 = n7928 & ~n64813;
  assign n64815 = ~n43545 & ~n64814;
  assign n64816 = ~i_hbusreq1 & ~n64815;
  assign n64817 = ~n47238 & ~n64816;
  assign n64818 = ~controllable_hgrant1 & ~n64817;
  assign n64819 = ~n64796 & ~n64818;
  assign n64820 = ~i_hbusreq3 & ~n64819;
  assign n64821 = ~n47226 & ~n64820;
  assign n64822 = ~controllable_hgrant3 & ~n64821;
  assign n64823 = ~n64786 & ~n64822;
  assign n64824 = ~i_hbusreq9 & ~n64823;
  assign n64825 = ~n47214 & ~n64824;
  assign n64826 = ~i_hbusreq4 & ~n64825;
  assign n64827 = ~n47213 & ~n64826;
  assign n64828 = ~controllable_hgrant4 & ~n64827;
  assign n64829 = ~n64776 & ~n64828;
  assign n64830 = ~i_hbusreq5 & ~n64829;
  assign n64831 = ~n47195 & ~n64830;
  assign n64832 = ~controllable_hgrant5 & ~n64831;
  assign n64833 = ~n64762 & ~n64832;
  assign n64834 = ~controllable_hmaster2 & ~n64833;
  assign n64835 = ~n64588 & ~n64834;
  assign n64836 = controllable_hmaster1 & ~n64835;
  assign n64837 = ~n8378 & ~n34419;
  assign n64838 = ~n49798 & ~n64837;
  assign n64839 = i_hlock5 & ~n64838;
  assign n64840 = ~n8378 & ~n34598;
  assign n64841 = ~n49798 & ~n64840;
  assign n64842 = ~i_hlock5 & ~n64841;
  assign n64843 = ~n64839 & ~n64842;
  assign n64844 = ~i_hbusreq5 & ~n64843;
  assign n64845 = ~n47284 & ~n64844;
  assign n64846 = controllable_hgrant5 & ~n64845;
  assign n64847 = ~n8426 & ~n25499;
  assign n64848 = ~n49812 & ~n64847;
  assign n64849 = ~i_hbusreq9 & ~n64848;
  assign n64850 = ~n47297 & ~n64849;
  assign n64851 = i_hlock4 & ~n64850;
  assign n64852 = ~n8426 & ~n25517;
  assign n64853 = ~n49819 & ~n64852;
  assign n64854 = ~i_hbusreq9 & ~n64853;
  assign n64855 = ~n47303 & ~n64854;
  assign n64856 = ~i_hlock4 & ~n64855;
  assign n64857 = ~n64851 & ~n64856;
  assign n64858 = ~i_hbusreq4 & ~n64857;
  assign n64859 = ~n47296 & ~n64858;
  assign n64860 = controllable_hgrant4 & ~n64859;
  assign n64861 = i_hlock4 & ~n64502;
  assign n64862 = ~i_hlock4 & ~n64553;
  assign n64863 = ~n64861 & ~n64862;
  assign n64864 = ~i_hbusreq4 & ~n64863;
  assign n64865 = ~n47313 & ~n64864;
  assign n64866 = ~controllable_hgrant4 & ~n64865;
  assign n64867 = ~n64860 & ~n64866;
  assign n64868 = ~i_hbusreq5 & ~n64867;
  assign n64869 = ~n47295 & ~n64868;
  assign n64870 = ~controllable_hgrant5 & ~n64869;
  assign n64871 = ~n64846 & ~n64870;
  assign n64872 = controllable_hmaster2 & ~n64871;
  assign n64873 = ~n49947 & ~n64872;
  assign n64874 = ~controllable_hmaster1 & ~n64873;
  assign n64875 = ~n64836 & ~n64874;
  assign n64876 = i_hlock6 & ~n64875;
  assign n64877 = controllable_hmaster2 & ~n64561;
  assign n64878 = ~n64834 & ~n64877;
  assign n64879 = controllable_hmaster1 & ~n64878;
  assign n64880 = ~n64874 & ~n64879;
  assign n64881 = ~i_hlock6 & ~n64880;
  assign n64882 = ~n64876 & ~n64881;
  assign n64883 = ~i_hbusreq6 & ~n64882;
  assign n64884 = ~n64752 & ~n64883;
  assign n64885 = ~controllable_hgrant6 & ~n64884;
  assign n64886 = ~n64751 & ~n64885;
  assign n64887 = ~controllable_hmaster0 & ~n64886;
  assign n64888 = ~n64734 & ~n64887;
  assign n64889 = ~i_hbusreq8 & ~n64888;
  assign n64890 = ~n64577 & ~n64889;
  assign n64891 = ~controllable_hmaster3 & ~n64890;
  assign n64892 = ~n64576 & ~n64891;
  assign n64893 = i_hlock7 & ~n64892;
  assign n64894 = i_hbusreq8 & ~n64254;
  assign n64895 = ~n8217 & ~n38914;
  assign n64896 = ~n49970 & ~n64895;
  assign n64897 = i_hlock6 & ~n64896;
  assign n64898 = ~n8217 & ~n38924;
  assign n64899 = ~n49970 & ~n64898;
  assign n64900 = ~i_hlock6 & ~n64899;
  assign n64901 = ~n64897 & ~n64900;
  assign n64902 = ~i_hbusreq6 & ~n64901;
  assign n64903 = ~n47441 & ~n64902;
  assign n64904 = controllable_hgrant6 & ~n64903;
  assign n64905 = ~n64640 & ~n64877;
  assign n64906 = controllable_hmaster1 & ~n64905;
  assign n64907 = ~n64728 & ~n64906;
  assign n64908 = ~i_hbusreq6 & ~n64907;
  assign n64909 = ~n47452 & ~n64908;
  assign n64910 = ~controllable_hgrant6 & ~n64909;
  assign n64911 = ~n64904 & ~n64910;
  assign n64912 = controllable_hmaster0 & ~n64911;
  assign n64913 = ~n64887 & ~n64912;
  assign n64914 = ~i_hbusreq8 & ~n64913;
  assign n64915 = ~n64894 & ~n64914;
  assign n64916 = ~controllable_hmaster3 & ~n64915;
  assign n64917 = ~n64576 & ~n64916;
  assign n64918 = ~i_hlock7 & ~n64917;
  assign n64919 = ~n64893 & ~n64918;
  assign n64920 = ~i_hbusreq7 & ~n64919;
  assign n64921 = ~n64259 & ~n64920;
  assign n64922 = n7924 & ~n64921;
  assign n64923 = ~n63107 & ~n64922;
  assign n64924 = n8214 & ~n64923;
  assign n64925 = ~n64229 & ~n64924;
  assign n64926 = ~n8202 & ~n64925;
  assign n64927 = ~n61598 & ~n64926;
  assign n64928 = n7920 & ~n64927;
  assign n64929 = ~n40177 & ~n64928;
  assign n64930 = n7728 & ~n64929;
  assign n64931 = ~n50003 & ~n64930;
  assign n64932 = ~n7723 & ~n64931;
  assign n64933 = ~n63740 & ~n64932;
  assign n64934 = ~n7714 & ~n64933;
  assign n64935 = ~n63739 & ~n64934;
  assign n64936 = ~n7705 & ~n64935;
  assign n64937 = ~n60620 & ~n64936;
  assign n64938 = n7808 & ~n64937;
  assign n64939 = ~n58944 & ~n64938;
  assign n64940 = n8195 & ~n64939;
  assign n64941 = ~n58412 & ~n64940;
  assign n64942 = n8193 & ~n64941;
  assign n64943 = ~n50015 & ~n64942;
  assign n64944 = n8191 & ~n64943;
  assign n64945 = ~n10989 & ~n39726;
  assign n64946 = n7728 & ~n64945;
  assign n64947 = ~n7834 & ~n10948;
  assign n64948 = ~controllable_hmaster1 & ~n64947;
  assign n64949 = ~n7833 & ~n64948;
  assign n64950 = ~controllable_hgrant6 & ~n64949;
  assign n64951 = ~n16262 & ~n64950;
  assign n64952 = controllable_hmaster0 & ~n64951;
  assign n64953 = ~controllable_hmaster0 & ~n7839;
  assign n64954 = ~n64952 & ~n64953;
  assign n64955 = controllable_hmaster3 & ~n64954;
  assign n64956 = controllable_hmaster3 & ~n64955;
  assign n64957 = i_hbusreq7 & ~n64956;
  assign n64958 = i_hbusreq8 & ~n64954;
  assign n64959 = i_hbusreq6 & ~n64949;
  assign n64960 = ~n7891 & ~n10971;
  assign n64961 = ~controllable_hmaster1 & ~n64960;
  assign n64962 = ~n7890 & ~n64961;
  assign n64963 = ~i_hbusreq6 & ~n64962;
  assign n64964 = ~n64959 & ~n64963;
  assign n64965 = ~controllable_hgrant6 & ~n64964;
  assign n64966 = ~n16274 & ~n64965;
  assign n64967 = controllable_hmaster0 & ~n64966;
  assign n64968 = ~controllable_hmaster0 & ~n7898;
  assign n64969 = ~n64967 & ~n64968;
  assign n64970 = ~i_hbusreq8 & ~n64969;
  assign n64971 = ~n64958 & ~n64970;
  assign n64972 = controllable_hmaster3 & ~n64971;
  assign n64973 = controllable_hmaster3 & ~n64972;
  assign n64974 = ~i_hbusreq7 & ~n64973;
  assign n64975 = ~n64957 & ~n64974;
  assign n64976 = n7924 & ~n64975;
  assign n64977 = ~n39731 & ~n64976;
  assign n64978 = ~n8214 & ~n64977;
  assign n64979 = ~n7904 & n8214;
  assign n64980 = ~n64978 & ~n64979;
  assign n64981 = ~n8202 & ~n64980;
  assign n64982 = ~n39741 & ~n64981;
  assign n64983 = ~n7728 & ~n64982;
  assign n64984 = ~n64946 & ~n64983;
  assign n64985 = ~n7723 & ~n64984;
  assign n64986 = ~n7723 & ~n64985;
  assign n64987 = ~n7714 & ~n64986;
  assign n64988 = ~n7714 & ~n64987;
  assign n64989 = n7705 & ~n64988;
  assign n64990 = n7723 & ~n64982;
  assign n64991 = ~n10948 & ~n39761;
  assign n64992 = ~controllable_hmaster1 & ~n64991;
  assign n64993 = ~n39760 & ~n64992;
  assign n64994 = ~controllable_hgrant6 & ~n64993;
  assign n64995 = ~n16305 & ~n64994;
  assign n64996 = controllable_hmaster0 & ~n64995;
  assign n64997 = ~controllable_hmaster0 & ~n39766;
  assign n64998 = ~n64996 & ~n64997;
  assign n64999 = controllable_hmaster3 & ~n64998;
  assign n65000 = ~n39916 & ~n64999;
  assign n65001 = i_hbusreq7 & ~n65000;
  assign n65002 = i_hbusreq8 & ~n64998;
  assign n65003 = i_hbusreq6 & ~n64993;
  assign n65004 = ~n10971 & ~n39946;
  assign n65005 = ~controllable_hmaster1 & ~n65004;
  assign n65006 = ~n39945 & ~n65005;
  assign n65007 = ~i_hbusreq6 & ~n65006;
  assign n65008 = ~n65003 & ~n65007;
  assign n65009 = ~controllable_hgrant6 & ~n65008;
  assign n65010 = ~n16317 & ~n65009;
  assign n65011 = controllable_hmaster0 & ~n65010;
  assign n65012 = ~controllable_hmaster0 & ~n39953;
  assign n65013 = ~n65011 & ~n65012;
  assign n65014 = ~i_hbusreq8 & ~n65013;
  assign n65015 = ~n65002 & ~n65014;
  assign n65016 = controllable_hmaster3 & ~n65015;
  assign n65017 = ~n40171 & ~n65016;
  assign n65018 = ~i_hbusreq7 & ~n65017;
  assign n65019 = ~n65001 & ~n65018;
  assign n65020 = n7924 & ~n65019;
  assign n65021 = ~n39731 & ~n65020;
  assign n65022 = ~n7920 & ~n65021;
  assign n65023 = n7920 & ~n64982;
  assign n65024 = ~n65022 & ~n65023;
  assign n65025 = ~n7723 & ~n65024;
  assign n65026 = ~n64990 & ~n65025;
  assign n65027 = n7714 & ~n65026;
  assign n65028 = ~n7714 & ~n65021;
  assign n65029 = ~n65027 & ~n65028;
  assign n65030 = ~n7705 & ~n65029;
  assign n65031 = ~n64989 & ~n65030;
  assign n65032 = ~n7808 & ~n65031;
  assign n65033 = ~n7920 & ~n64945;
  assign n65034 = ~n40785 & ~n65033;
  assign n65035 = n7728 & ~n65034;
  assign n65036 = ~n7920 & ~n64982;
  assign n65037 = ~n41275 & ~n65036;
  assign n65038 = ~n7728 & ~n65037;
  assign n65039 = ~n65035 & ~n65038;
  assign n65040 = ~n7723 & ~n65039;
  assign n65041 = ~n7723 & ~n65040;
  assign n65042 = ~n7714 & ~n65041;
  assign n65043 = ~n7714 & ~n65042;
  assign n65044 = n7705 & ~n65043;
  assign n65045 = ~n42700 & ~n65036;
  assign n65046 = n7728 & ~n65045;
  assign n65047 = ~n45926 & ~n65036;
  assign n65048 = ~n7728 & ~n65047;
  assign n65049 = ~n65046 & ~n65048;
  assign n65050 = n7723 & ~n65049;
  assign n65051 = ~n7723 & ~n65047;
  assign n65052 = ~n65050 & ~n65051;
  assign n65053 = n7714 & ~n65052;
  assign n65054 = n7723 & ~n65047;
  assign n65055 = ~n48003 & ~n65022;
  assign n65056 = n7728 & ~n65055;
  assign n65057 = ~n50001 & ~n65022;
  assign n65058 = ~n7728 & ~n65057;
  assign n65059 = ~n65056 & ~n65058;
  assign n65060 = ~n7723 & ~n65059;
  assign n65061 = ~n65054 & ~n65060;
  assign n65062 = ~n7714 & ~n65061;
  assign n65063 = ~n65053 & ~n65062;
  assign n65064 = ~n7705 & ~n65063;
  assign n65065 = ~n65044 & ~n65064;
  assign n65066 = n7808 & ~n65065;
  assign n65067 = ~n65032 & ~n65066;
  assign n65068 = n8195 & ~n65067;
  assign n65069 = ~n39684 & ~n65068;
  assign n65070 = ~n8193 & ~n65069;
  assign n65071 = ~n50187 & ~n65022;
  assign n65072 = ~n7723 & ~n65071;
  assign n65073 = ~n50186 & ~n65072;
  assign n65074 = n7714 & ~n65073;
  assign n65075 = ~n65028 & ~n65074;
  assign n65076 = ~n7705 & ~n65075;
  assign n65077 = ~n50185 & ~n65076;
  assign n65078 = ~n7808 & ~n65077;
  assign n65079 = ~n58400 & ~n65022;
  assign n65080 = n7728 & ~n65079;
  assign n65081 = ~n65058 & ~n65080;
  assign n65082 = ~n7723 & ~n65081;
  assign n65083 = ~n56860 & ~n65082;
  assign n65084 = ~n7714 & ~n65083;
  assign n65085 = ~n56859 & ~n65084;
  assign n65086 = ~n7705 & ~n65085;
  assign n65087 = ~n51653 & ~n65086;
  assign n65088 = n7808 & ~n65087;
  assign n65089 = ~n65078 & ~n65088;
  assign n65090 = ~n8195 & ~n65089;
  assign n65091 = ~n11129 & ~n58532;
  assign n65092 = ~controllable_hmaster1 & ~n65091;
  assign n65093 = ~n58531 & ~n65092;
  assign n65094 = ~controllable_hgrant6 & ~n65093;
  assign n65095 = ~n23630 & ~n65094;
  assign n65096 = controllable_hmaster0 & ~n65095;
  assign n65097 = ~controllable_hmaster0 & ~n58537;
  assign n65098 = ~n65096 & ~n65097;
  assign n65099 = controllable_hmaster3 & ~n65098;
  assign n65100 = ~n58661 & ~n65099;
  assign n65101 = i_hbusreq7 & ~n65100;
  assign n65102 = i_hbusreq8 & ~n65098;
  assign n65103 = i_hbusreq6 & ~n65093;
  assign n65104 = ~n11153 & ~n58693;
  assign n65105 = ~controllable_hmaster1 & ~n65104;
  assign n65106 = ~n58692 & ~n65105;
  assign n65107 = ~i_hbusreq6 & ~n65106;
  assign n65108 = ~n65103 & ~n65107;
  assign n65109 = ~controllable_hgrant6 & ~n65108;
  assign n65110 = ~n23666 & ~n65109;
  assign n65111 = controllable_hmaster0 & ~n65110;
  assign n65112 = ~controllable_hmaster0 & ~n58700;
  assign n65113 = ~n65111 & ~n65112;
  assign n65114 = ~i_hbusreq8 & ~n65113;
  assign n65115 = ~n65102 & ~n65114;
  assign n65116 = controllable_hmaster3 & ~n65115;
  assign n65117 = ~n58895 & ~n65116;
  assign n65118 = ~i_hbusreq7 & ~n65117;
  assign n65119 = ~n65101 & ~n65118;
  assign n65120 = n7924 & ~n65119;
  assign n65121 = ~n58519 & ~n65120;
  assign n65122 = n8214 & ~n65121;
  assign n65123 = n8214 & ~n65122;
  assign n65124 = n8202 & ~n65123;
  assign n65125 = ~n58446 & ~n65124;
  assign n65126 = n7728 & ~n65125;
  assign n65127 = n8214 & ~n65021;
  assign n65128 = ~n39730 & ~n65127;
  assign n65129 = n8202 & ~n65128;
  assign n65130 = ~n58923 & ~n65129;
  assign n65131 = ~n7728 & ~n65130;
  assign n65132 = ~n65126 & ~n65131;
  assign n65133 = ~n7723 & ~n65132;
  assign n65134 = ~n7723 & ~n65133;
  assign n65135 = ~n7714 & ~n65134;
  assign n65136 = ~n7714 & ~n65135;
  assign n65137 = n7705 & ~n65136;
  assign n65138 = n7723 & ~n65130;
  assign n65139 = n7920 & ~n65130;
  assign n65140 = ~n65022 & ~n65139;
  assign n65141 = ~n7723 & ~n65140;
  assign n65142 = ~n65138 & ~n65141;
  assign n65143 = n7714 & ~n65142;
  assign n65144 = ~n65028 & ~n65143;
  assign n65145 = ~n7705 & ~n65144;
  assign n65146 = ~n65137 & ~n65145;
  assign n65147 = ~n7808 & ~n65146;
  assign n65148 = ~n7920 & ~n65125;
  assign n65149 = ~n60195 & ~n65148;
  assign n65150 = n7728 & ~n65149;
  assign n65151 = ~n7920 & ~n65130;
  assign n65152 = ~n60612 & ~n65151;
  assign n65153 = ~n7728 & ~n65152;
  assign n65154 = ~n65150 & ~n65153;
  assign n65155 = ~n7723 & ~n65154;
  assign n65156 = ~n7723 & ~n65155;
  assign n65157 = ~n7714 & ~n65156;
  assign n65158 = ~n7714 & ~n65157;
  assign n65159 = n7705 & ~n65158;
  assign n65160 = ~n61600 & ~n65151;
  assign n65161 = n7728 & ~n65160;
  assign n65162 = ~n63732 & ~n65151;
  assign n65163 = ~n7728 & ~n65162;
  assign n65164 = ~n65161 & ~n65163;
  assign n65165 = n7723 & ~n65164;
  assign n65166 = ~n7723 & ~n65162;
  assign n65167 = ~n65165 & ~n65166;
  assign n65168 = n7714 & ~n65167;
  assign n65169 = n7723 & ~n65162;
  assign n65170 = ~n64928 & ~n65022;
  assign n65171 = n7728 & ~n65170;
  assign n65172 = ~n65058 & ~n65171;
  assign n65173 = ~n7723 & ~n65172;
  assign n65174 = ~n65169 & ~n65173;
  assign n65175 = ~n7714 & ~n65174;
  assign n65176 = ~n65168 & ~n65175;
  assign n65177 = ~n7705 & ~n65176;
  assign n65178 = ~n65159 & ~n65177;
  assign n65179 = n7808 & ~n65178;
  assign n65180 = ~n65147 & ~n65179;
  assign n65181 = n8195 & ~n65180;
  assign n65182 = ~n65090 & ~n65181;
  assign n65183 = n8193 & ~n65182;
  assign n65184 = ~n65070 & ~n65183;
  assign n65185 = ~n8191 & ~n65184;
  assign n65186 = ~n64944 & ~n65185;
  assign n65187 = n8188 & ~n65186;
  assign n65188 = ~n11286 & ~n39726;
  assign n65189 = n7728 & ~n65188;
  assign n65190 = controllable_hmaster0 & ~n7839;
  assign n65191 = ~n7834 & ~n11236;
  assign n65192 = ~controllable_hmaster1 & ~n65191;
  assign n65193 = ~n7833 & ~n65192;
  assign n65194 = ~controllable_hgrant6 & ~n65193;
  assign n65195 = ~n36399 & ~n65194;
  assign n65196 = ~controllable_hmaster0 & ~n65195;
  assign n65197 = ~n65190 & ~n65196;
  assign n65198 = i_hlock8 & ~n65197;
  assign n65199 = ~n7834 & ~n11243;
  assign n65200 = ~controllable_hmaster1 & ~n65199;
  assign n65201 = ~n7833 & ~n65200;
  assign n65202 = ~controllable_hgrant6 & ~n65201;
  assign n65203 = ~n36408 & ~n65202;
  assign n65204 = ~controllable_hmaster0 & ~n65203;
  assign n65205 = ~n65190 & ~n65204;
  assign n65206 = ~i_hlock8 & ~n65205;
  assign n65207 = ~n65198 & ~n65206;
  assign n65208 = controllable_hmaster3 & ~n65207;
  assign n65209 = controllable_hmaster3 & ~n65208;
  assign n65210 = i_hbusreq7 & ~n65209;
  assign n65211 = i_hbusreq8 & ~n65207;
  assign n65212 = controllable_hmaster0 & ~n7898;
  assign n65213 = i_hbusreq6 & ~n65193;
  assign n65214 = ~n7891 & ~n11256;
  assign n65215 = ~controllable_hmaster1 & ~n65214;
  assign n65216 = ~n7890 & ~n65215;
  assign n65217 = ~i_hbusreq6 & ~n65216;
  assign n65218 = ~n65213 & ~n65217;
  assign n65219 = ~controllable_hgrant6 & ~n65218;
  assign n65220 = ~n36422 & ~n65219;
  assign n65221 = ~controllable_hmaster0 & ~n65220;
  assign n65222 = ~n65212 & ~n65221;
  assign n65223 = i_hlock8 & ~n65222;
  assign n65224 = i_hbusreq6 & ~n65201;
  assign n65225 = ~n7891 & ~n11266;
  assign n65226 = ~controllable_hmaster1 & ~n65225;
  assign n65227 = ~n7890 & ~n65226;
  assign n65228 = ~i_hbusreq6 & ~n65227;
  assign n65229 = ~n65224 & ~n65228;
  assign n65230 = ~controllable_hgrant6 & ~n65229;
  assign n65231 = ~n36434 & ~n65230;
  assign n65232 = ~controllable_hmaster0 & ~n65231;
  assign n65233 = ~n65212 & ~n65232;
  assign n65234 = ~i_hlock8 & ~n65233;
  assign n65235 = ~n65223 & ~n65234;
  assign n65236 = ~i_hbusreq8 & ~n65235;
  assign n65237 = ~n65211 & ~n65236;
  assign n65238 = controllable_hmaster3 & ~n65237;
  assign n65239 = controllable_hmaster3 & ~n65238;
  assign n65240 = ~i_hbusreq7 & ~n65239;
  assign n65241 = ~n65210 & ~n65240;
  assign n65242 = n7924 & ~n65241;
  assign n65243 = ~n39731 & ~n65242;
  assign n65244 = n8214 & ~n65243;
  assign n65245 = ~n39730 & ~n65244;
  assign n65246 = ~n8202 & ~n65245;
  assign n65247 = ~n39741 & ~n65246;
  assign n65248 = ~n7728 & ~n65247;
  assign n65249 = ~n65189 & ~n65248;
  assign n65250 = ~n7723 & ~n65249;
  assign n65251 = ~n7723 & ~n65250;
  assign n65252 = ~n7714 & ~n65251;
  assign n65253 = ~n7714 & ~n65252;
  assign n65254 = n7705 & ~n65253;
  assign n65255 = n7723 & ~n65247;
  assign n65256 = controllable_hmaster0 & ~n39766;
  assign n65257 = ~n11236 & ~n39761;
  assign n65258 = ~controllable_hmaster1 & ~n65257;
  assign n65259 = ~n39760 & ~n65258;
  assign n65260 = ~controllable_hgrant6 & ~n65259;
  assign n65261 = ~n36467 & ~n65260;
  assign n65262 = ~controllable_hmaster0 & ~n65261;
  assign n65263 = ~n65256 & ~n65262;
  assign n65264 = i_hlock8 & ~n65263;
  assign n65265 = ~n11243 & ~n39761;
  assign n65266 = ~controllable_hmaster1 & ~n65265;
  assign n65267 = ~n39760 & ~n65266;
  assign n65268 = ~controllable_hgrant6 & ~n65267;
  assign n65269 = ~n36476 & ~n65268;
  assign n65270 = ~controllable_hmaster0 & ~n65269;
  assign n65271 = ~n65256 & ~n65270;
  assign n65272 = ~i_hlock8 & ~n65271;
  assign n65273 = ~n65264 & ~n65272;
  assign n65274 = controllable_hmaster3 & ~n65273;
  assign n65275 = ~n39916 & ~n65274;
  assign n65276 = i_hbusreq7 & ~n65275;
  assign n65277 = i_hbusreq8 & ~n65273;
  assign n65278 = controllable_hmaster0 & ~n39953;
  assign n65279 = i_hbusreq6 & ~n65259;
  assign n65280 = ~n11256 & ~n39946;
  assign n65281 = ~controllable_hmaster1 & ~n65280;
  assign n65282 = ~n39945 & ~n65281;
  assign n65283 = ~i_hbusreq6 & ~n65282;
  assign n65284 = ~n65279 & ~n65283;
  assign n65285 = ~controllable_hgrant6 & ~n65284;
  assign n65286 = ~n36490 & ~n65285;
  assign n65287 = ~controllable_hmaster0 & ~n65286;
  assign n65288 = ~n65278 & ~n65287;
  assign n65289 = i_hlock8 & ~n65288;
  assign n65290 = i_hbusreq6 & ~n65267;
  assign n65291 = ~n11266 & ~n39946;
  assign n65292 = ~controllable_hmaster1 & ~n65291;
  assign n65293 = ~n39945 & ~n65292;
  assign n65294 = ~i_hbusreq6 & ~n65293;
  assign n65295 = ~n65290 & ~n65294;
  assign n65296 = ~controllable_hgrant6 & ~n65295;
  assign n65297 = ~n36502 & ~n65296;
  assign n65298 = ~controllable_hmaster0 & ~n65297;
  assign n65299 = ~n65278 & ~n65298;
  assign n65300 = ~i_hlock8 & ~n65299;
  assign n65301 = ~n65289 & ~n65300;
  assign n65302 = ~i_hbusreq8 & ~n65301;
  assign n65303 = ~n65277 & ~n65302;
  assign n65304 = controllable_hmaster3 & ~n65303;
  assign n65305 = ~n40171 & ~n65304;
  assign n65306 = ~i_hbusreq7 & ~n65305;
  assign n65307 = ~n65276 & ~n65306;
  assign n65308 = n7924 & ~n65307;
  assign n65309 = ~n39731 & ~n65308;
  assign n65310 = ~n7920 & ~n65309;
  assign n65311 = n7920 & ~n65247;
  assign n65312 = ~n65310 & ~n65311;
  assign n65313 = ~n7723 & ~n65312;
  assign n65314 = ~n65255 & ~n65313;
  assign n65315 = n7714 & ~n65314;
  assign n65316 = ~n7714 & ~n65309;
  assign n65317 = ~n65315 & ~n65316;
  assign n65318 = ~n7705 & ~n65317;
  assign n65319 = ~n65254 & ~n65318;
  assign n65320 = ~n7808 & ~n65319;
  assign n65321 = ~n7920 & ~n65188;
  assign n65322 = ~n40785 & ~n65321;
  assign n65323 = n7728 & ~n65322;
  assign n65324 = ~n7920 & ~n65247;
  assign n65325 = ~n41275 & ~n65324;
  assign n65326 = ~n7728 & ~n65325;
  assign n65327 = ~n65323 & ~n65326;
  assign n65328 = ~n7723 & ~n65327;
  assign n65329 = ~n7723 & ~n65328;
  assign n65330 = ~n7714 & ~n65329;
  assign n65331 = ~n7714 & ~n65330;
  assign n65332 = n7705 & ~n65331;
  assign n65333 = ~n42700 & ~n65324;
  assign n65334 = n7728 & ~n65333;
  assign n65335 = ~n45926 & ~n65324;
  assign n65336 = ~n7728 & ~n65335;
  assign n65337 = ~n65334 & ~n65336;
  assign n65338 = n7723 & ~n65337;
  assign n65339 = ~n7723 & ~n65335;
  assign n65340 = ~n65338 & ~n65339;
  assign n65341 = n7714 & ~n65340;
  assign n65342 = n7723 & ~n65335;
  assign n65343 = ~n48003 & ~n65310;
  assign n65344 = n7728 & ~n65343;
  assign n65345 = ~n50001 & ~n65310;
  assign n65346 = ~n7728 & ~n65345;
  assign n65347 = ~n65344 & ~n65346;
  assign n65348 = ~n7723 & ~n65347;
  assign n65349 = ~n65342 & ~n65348;
  assign n65350 = ~n7714 & ~n65349;
  assign n65351 = ~n65341 & ~n65350;
  assign n65352 = ~n7705 & ~n65351;
  assign n65353 = ~n65332 & ~n65352;
  assign n65354 = n7808 & ~n65353;
  assign n65355 = ~n65320 & ~n65354;
  assign n65356 = n8195 & ~n65355;
  assign n65357 = ~n39684 & ~n65356;
  assign n65358 = ~n8193 & ~n65357;
  assign n65359 = ~n50187 & ~n65310;
  assign n65360 = ~n7723 & ~n65359;
  assign n65361 = ~n50186 & ~n65360;
  assign n65362 = n7714 & ~n65361;
  assign n65363 = ~n65316 & ~n65362;
  assign n65364 = ~n7705 & ~n65363;
  assign n65365 = ~n50185 & ~n65364;
  assign n65366 = ~n7808 & ~n65365;
  assign n65367 = ~n58400 & ~n65310;
  assign n65368 = n7728 & ~n65367;
  assign n65369 = ~n65346 & ~n65368;
  assign n65370 = ~n7723 & ~n65369;
  assign n65371 = ~n56860 & ~n65370;
  assign n65372 = ~n7714 & ~n65371;
  assign n65373 = ~n56859 & ~n65372;
  assign n65374 = ~n7705 & ~n65373;
  assign n65375 = ~n51653 & ~n65374;
  assign n65376 = n7808 & ~n65375;
  assign n65377 = ~n65366 & ~n65376;
  assign n65378 = ~n8195 & ~n65377;
  assign n65379 = controllable_hmaster0 & ~n58537;
  assign n65380 = ~n11461 & ~n58532;
  assign n65381 = ~controllable_hmaster1 & ~n65380;
  assign n65382 = ~n58531 & ~n65381;
  assign n65383 = ~controllable_hgrant6 & ~n65382;
  assign n65384 = ~n38384 & ~n65383;
  assign n65385 = ~controllable_hmaster0 & ~n65384;
  assign n65386 = ~n65379 & ~n65385;
  assign n65387 = i_hlock8 & ~n65386;
  assign n65388 = ~n11468 & ~n58532;
  assign n65389 = ~controllable_hmaster1 & ~n65388;
  assign n65390 = ~n58531 & ~n65389;
  assign n65391 = ~controllable_hgrant6 & ~n65390;
  assign n65392 = ~n38394 & ~n65391;
  assign n65393 = ~controllable_hmaster0 & ~n65392;
  assign n65394 = ~n65379 & ~n65393;
  assign n65395 = ~i_hlock8 & ~n65394;
  assign n65396 = ~n65387 & ~n65395;
  assign n65397 = controllable_hmaster3 & ~n65396;
  assign n65398 = ~n58661 & ~n65397;
  assign n65399 = i_hbusreq7 & ~n65398;
  assign n65400 = i_hbusreq8 & ~n65396;
  assign n65401 = controllable_hmaster0 & ~n58700;
  assign n65402 = i_hbusreq6 & ~n65382;
  assign n65403 = ~n11482 & ~n58693;
  assign n65404 = ~controllable_hmaster1 & ~n65403;
  assign n65405 = ~n58692 & ~n65404;
  assign n65406 = ~i_hbusreq6 & ~n65405;
  assign n65407 = ~n65402 & ~n65406;
  assign n65408 = ~controllable_hgrant6 & ~n65407;
  assign n65409 = ~n38409 & ~n65408;
  assign n65410 = ~controllable_hmaster0 & ~n65409;
  assign n65411 = ~n65401 & ~n65410;
  assign n65412 = i_hlock8 & ~n65411;
  assign n65413 = i_hbusreq6 & ~n65390;
  assign n65414 = ~n11492 & ~n58693;
  assign n65415 = ~controllable_hmaster1 & ~n65414;
  assign n65416 = ~n58692 & ~n65415;
  assign n65417 = ~i_hbusreq6 & ~n65416;
  assign n65418 = ~n65413 & ~n65417;
  assign n65419 = ~controllable_hgrant6 & ~n65418;
  assign n65420 = ~n38422 & ~n65419;
  assign n65421 = ~controllable_hmaster0 & ~n65420;
  assign n65422 = ~n65401 & ~n65421;
  assign n65423 = ~i_hlock8 & ~n65422;
  assign n65424 = ~n65412 & ~n65423;
  assign n65425 = ~i_hbusreq8 & ~n65424;
  assign n65426 = ~n65400 & ~n65425;
  assign n65427 = controllable_hmaster3 & ~n65426;
  assign n65428 = ~n58895 & ~n65427;
  assign n65429 = ~i_hbusreq7 & ~n65428;
  assign n65430 = ~n65399 & ~n65429;
  assign n65431 = n7924 & ~n65430;
  assign n65432 = ~n58519 & ~n65431;
  assign n65433 = n8214 & ~n65432;
  assign n65434 = n8214 & ~n65433;
  assign n65435 = n8202 & ~n65434;
  assign n65436 = ~n58446 & ~n65435;
  assign n65437 = n7728 & ~n65436;
  assign n65438 = n8214 & ~n65309;
  assign n65439 = ~n39730 & ~n65438;
  assign n65440 = n8202 & ~n65439;
  assign n65441 = ~n58923 & ~n65440;
  assign n65442 = ~n7728 & ~n65441;
  assign n65443 = ~n65437 & ~n65442;
  assign n65444 = ~n7723 & ~n65443;
  assign n65445 = ~n7723 & ~n65444;
  assign n65446 = ~n7714 & ~n65445;
  assign n65447 = ~n7714 & ~n65446;
  assign n65448 = n7705 & ~n65447;
  assign n65449 = n7723 & ~n65441;
  assign n65450 = n7920 & ~n65441;
  assign n65451 = ~n65310 & ~n65450;
  assign n65452 = ~n7723 & ~n65451;
  assign n65453 = ~n65449 & ~n65452;
  assign n65454 = n7714 & ~n65453;
  assign n65455 = ~n65316 & ~n65454;
  assign n65456 = ~n7705 & ~n65455;
  assign n65457 = ~n65448 & ~n65456;
  assign n65458 = ~n7808 & ~n65457;
  assign n65459 = ~n7920 & ~n65436;
  assign n65460 = ~n60195 & ~n65459;
  assign n65461 = n7728 & ~n65460;
  assign n65462 = ~n7920 & ~n65441;
  assign n65463 = ~n60612 & ~n65462;
  assign n65464 = ~n7728 & ~n65463;
  assign n65465 = ~n65461 & ~n65464;
  assign n65466 = ~n7723 & ~n65465;
  assign n65467 = ~n7723 & ~n65466;
  assign n65468 = ~n7714 & ~n65467;
  assign n65469 = ~n7714 & ~n65468;
  assign n65470 = n7705 & ~n65469;
  assign n65471 = ~n61600 & ~n65462;
  assign n65472 = n7728 & ~n65471;
  assign n65473 = ~n63732 & ~n65462;
  assign n65474 = ~n7728 & ~n65473;
  assign n65475 = ~n65472 & ~n65474;
  assign n65476 = n7723 & ~n65475;
  assign n65477 = ~n7723 & ~n65473;
  assign n65478 = ~n65476 & ~n65477;
  assign n65479 = n7714 & ~n65478;
  assign n65480 = n7723 & ~n65473;
  assign n65481 = ~n64928 & ~n65310;
  assign n65482 = n7728 & ~n65481;
  assign n65483 = ~n65346 & ~n65482;
  assign n65484 = ~n7723 & ~n65483;
  assign n65485 = ~n65480 & ~n65484;
  assign n65486 = ~n7714 & ~n65485;
  assign n65487 = ~n65479 & ~n65486;
  assign n65488 = ~n7705 & ~n65487;
  assign n65489 = ~n65470 & ~n65488;
  assign n65490 = n7808 & ~n65489;
  assign n65491 = ~n65458 & ~n65490;
  assign n65492 = n8195 & ~n65491;
  assign n65493 = ~n65378 & ~n65492;
  assign n65494 = n8193 & ~n65493;
  assign n65495 = ~n65358 & ~n65494;
  assign n65496 = n8191 & ~n65495;
  assign n65497 = ~n11575 & ~n39726;
  assign n65498 = n7728 & ~n65497;
  assign n65499 = ~n64978 & ~n65244;
  assign n65500 = ~n8202 & ~n65499;
  assign n65501 = ~n39741 & ~n65500;
  assign n65502 = ~n7728 & ~n65501;
  assign n65503 = ~n65498 & ~n65502;
  assign n65504 = ~n7723 & ~n65503;
  assign n65505 = ~n7723 & ~n65504;
  assign n65506 = ~n7714 & ~n65505;
  assign n65507 = ~n7714 & ~n65506;
  assign n65508 = n7705 & ~n65507;
  assign n65509 = n7723 & ~n65501;
  assign n65510 = ~n64996 & ~n65262;
  assign n65511 = i_hlock8 & ~n65510;
  assign n65512 = ~n64996 & ~n65270;
  assign n65513 = ~i_hlock8 & ~n65512;
  assign n65514 = ~n65511 & ~n65513;
  assign n65515 = controllable_hmaster3 & ~n65514;
  assign n65516 = ~n39916 & ~n65515;
  assign n65517 = i_hbusreq7 & ~n65516;
  assign n65518 = i_hbusreq8 & ~n65514;
  assign n65519 = ~n65011 & ~n65287;
  assign n65520 = i_hlock8 & ~n65519;
  assign n65521 = ~n65011 & ~n65298;
  assign n65522 = ~i_hlock8 & ~n65521;
  assign n65523 = ~n65520 & ~n65522;
  assign n65524 = ~i_hbusreq8 & ~n65523;
  assign n65525 = ~n65518 & ~n65524;
  assign n65526 = controllable_hmaster3 & ~n65525;
  assign n65527 = ~n40171 & ~n65526;
  assign n65528 = ~i_hbusreq7 & ~n65527;
  assign n65529 = ~n65517 & ~n65528;
  assign n65530 = n7924 & ~n65529;
  assign n65531 = ~n39731 & ~n65530;
  assign n65532 = ~n7920 & ~n65531;
  assign n65533 = n7920 & ~n65501;
  assign n65534 = ~n65532 & ~n65533;
  assign n65535 = ~n7723 & ~n65534;
  assign n65536 = ~n65509 & ~n65535;
  assign n65537 = n7714 & ~n65536;
  assign n65538 = ~n7714 & ~n65531;
  assign n65539 = ~n65537 & ~n65538;
  assign n65540 = ~n7705 & ~n65539;
  assign n65541 = ~n65508 & ~n65540;
  assign n65542 = ~n7808 & ~n65541;
  assign n65543 = ~n7920 & ~n65497;
  assign n65544 = ~n40785 & ~n65543;
  assign n65545 = n7728 & ~n65544;
  assign n65546 = ~n7920 & ~n65501;
  assign n65547 = ~n41275 & ~n65546;
  assign n65548 = ~n7728 & ~n65547;
  assign n65549 = ~n65545 & ~n65548;
  assign n65550 = ~n7723 & ~n65549;
  assign n65551 = ~n7723 & ~n65550;
  assign n65552 = ~n7714 & ~n65551;
  assign n65553 = ~n7714 & ~n65552;
  assign n65554 = n7705 & ~n65553;
  assign n65555 = ~n42700 & ~n65546;
  assign n65556 = n7728 & ~n65555;
  assign n65557 = ~n45926 & ~n65546;
  assign n65558 = ~n7728 & ~n65557;
  assign n65559 = ~n65556 & ~n65558;
  assign n65560 = n7723 & ~n65559;
  assign n65561 = ~n7723 & ~n65557;
  assign n65562 = ~n65560 & ~n65561;
  assign n65563 = n7714 & ~n65562;
  assign n65564 = n7723 & ~n65557;
  assign n65565 = ~n48003 & ~n65532;
  assign n65566 = n7728 & ~n65565;
  assign n65567 = ~n50001 & ~n65532;
  assign n65568 = ~n7728 & ~n65567;
  assign n65569 = ~n65566 & ~n65568;
  assign n65570 = ~n7723 & ~n65569;
  assign n65571 = ~n65564 & ~n65570;
  assign n65572 = ~n7714 & ~n65571;
  assign n65573 = ~n65563 & ~n65572;
  assign n65574 = ~n7705 & ~n65573;
  assign n65575 = ~n65554 & ~n65574;
  assign n65576 = n7808 & ~n65575;
  assign n65577 = ~n65542 & ~n65576;
  assign n65578 = n8195 & ~n65577;
  assign n65579 = ~n39684 & ~n65578;
  assign n65580 = ~n8193 & ~n65579;
  assign n65581 = ~n50187 & ~n65532;
  assign n65582 = ~n7723 & ~n65581;
  assign n65583 = ~n50186 & ~n65582;
  assign n65584 = n7714 & ~n65583;
  assign n65585 = ~n65538 & ~n65584;
  assign n65586 = ~n7705 & ~n65585;
  assign n65587 = ~n50185 & ~n65586;
  assign n65588 = ~n7808 & ~n65587;
  assign n65589 = ~n58400 & ~n65532;
  assign n65590 = n7728 & ~n65589;
  assign n65591 = ~n65568 & ~n65590;
  assign n65592 = ~n7723 & ~n65591;
  assign n65593 = ~n56860 & ~n65592;
  assign n65594 = ~n7714 & ~n65593;
  assign n65595 = ~n56859 & ~n65594;
  assign n65596 = ~n7705 & ~n65595;
  assign n65597 = ~n51653 & ~n65596;
  assign n65598 = n7808 & ~n65597;
  assign n65599 = ~n65588 & ~n65598;
  assign n65600 = ~n8195 & ~n65599;
  assign n65601 = ~n65096 & ~n65385;
  assign n65602 = i_hlock8 & ~n65601;
  assign n65603 = ~n65096 & ~n65393;
  assign n65604 = ~i_hlock8 & ~n65603;
  assign n65605 = ~n65602 & ~n65604;
  assign n65606 = controllable_hmaster3 & ~n65605;
  assign n65607 = ~n58661 & ~n65606;
  assign n65608 = i_hbusreq7 & ~n65607;
  assign n65609 = i_hbusreq8 & ~n65605;
  assign n65610 = ~n65111 & ~n65410;
  assign n65611 = i_hlock8 & ~n65610;
  assign n65612 = ~n65111 & ~n65421;
  assign n65613 = ~i_hlock8 & ~n65612;
  assign n65614 = ~n65611 & ~n65613;
  assign n65615 = ~i_hbusreq8 & ~n65614;
  assign n65616 = ~n65609 & ~n65615;
  assign n65617 = controllable_hmaster3 & ~n65616;
  assign n65618 = ~n58895 & ~n65617;
  assign n65619 = ~i_hbusreq7 & ~n65618;
  assign n65620 = ~n65608 & ~n65619;
  assign n65621 = n7924 & ~n65620;
  assign n65622 = ~n58519 & ~n65621;
  assign n65623 = n8214 & ~n65622;
  assign n65624 = n8214 & ~n65623;
  assign n65625 = n8202 & ~n65624;
  assign n65626 = ~n58446 & ~n65625;
  assign n65627 = n7728 & ~n65626;
  assign n65628 = n8214 & ~n65531;
  assign n65629 = ~n39730 & ~n65628;
  assign n65630 = n8202 & ~n65629;
  assign n65631 = ~n58923 & ~n65630;
  assign n65632 = ~n7728 & ~n65631;
  assign n65633 = ~n65627 & ~n65632;
  assign n65634 = ~n7723 & ~n65633;
  assign n65635 = ~n7723 & ~n65634;
  assign n65636 = ~n7714 & ~n65635;
  assign n65637 = ~n7714 & ~n65636;
  assign n65638 = n7705 & ~n65637;
  assign n65639 = n7723 & ~n65631;
  assign n65640 = n7920 & ~n65631;
  assign n65641 = ~n65532 & ~n65640;
  assign n65642 = ~n7723 & ~n65641;
  assign n65643 = ~n65639 & ~n65642;
  assign n65644 = n7714 & ~n65643;
  assign n65645 = ~n65538 & ~n65644;
  assign n65646 = ~n7705 & ~n65645;
  assign n65647 = ~n65638 & ~n65646;
  assign n65648 = ~n7808 & ~n65647;
  assign n65649 = ~n7920 & ~n65626;
  assign n65650 = ~n60195 & ~n65649;
  assign n65651 = n7728 & ~n65650;
  assign n65652 = ~n7920 & ~n65631;
  assign n65653 = ~n60612 & ~n65652;
  assign n65654 = ~n7728 & ~n65653;
  assign n65655 = ~n65651 & ~n65654;
  assign n65656 = ~n7723 & ~n65655;
  assign n65657 = ~n7723 & ~n65656;
  assign n65658 = ~n7714 & ~n65657;
  assign n65659 = ~n7714 & ~n65658;
  assign n65660 = n7705 & ~n65659;
  assign n65661 = ~n61600 & ~n65652;
  assign n65662 = n7728 & ~n65661;
  assign n65663 = ~n63732 & ~n65652;
  assign n65664 = ~n7728 & ~n65663;
  assign n65665 = ~n65662 & ~n65664;
  assign n65666 = n7723 & ~n65665;
  assign n65667 = ~n7723 & ~n65663;
  assign n65668 = ~n65666 & ~n65667;
  assign n65669 = n7714 & ~n65668;
  assign n65670 = n7723 & ~n65663;
  assign n65671 = ~n64928 & ~n65532;
  assign n65672 = n7728 & ~n65671;
  assign n65673 = ~n65568 & ~n65672;
  assign n65674 = ~n7723 & ~n65673;
  assign n65675 = ~n65670 & ~n65674;
  assign n65676 = ~n7714 & ~n65675;
  assign n65677 = ~n65669 & ~n65676;
  assign n65678 = ~n7705 & ~n65677;
  assign n65679 = ~n65660 & ~n65678;
  assign n65680 = n7808 & ~n65679;
  assign n65681 = ~n65648 & ~n65680;
  assign n65682 = n8195 & ~n65681;
  assign n65683 = ~n65600 & ~n65682;
  assign n65684 = n8193 & ~n65683;
  assign n65685 = ~n65580 & ~n65684;
  assign n65686 = ~n8191 & ~n65685;
  assign n65687 = ~n65496 & ~n65686;
  assign n65688 = ~n8188 & ~n65687;
  assign n65689 = ~n65187 & ~n65688;
  assign n65690 = n8185 & ~n65689;
  assign n65691 = ~n11809 & ~n39724;
  assign n65692 = n8202 & ~n65691;
  assign n65693 = n8202 & ~n65692;
  assign n65694 = n7728 & ~n65693;
  assign n65695 = ~n7840 & ~n11772;
  assign n65696 = i_hlock7 & ~n65695;
  assign n65697 = ~n7840 & ~n11777;
  assign n65698 = ~i_hlock7 & ~n65697;
  assign n65699 = ~n65696 & ~n65698;
  assign n65700 = i_hbusreq7 & ~n65699;
  assign n65701 = ~n7901 & ~n11790;
  assign n65702 = i_hlock7 & ~n65701;
  assign n65703 = ~n7901 & ~n11801;
  assign n65704 = ~i_hlock7 & ~n65703;
  assign n65705 = ~n65702 & ~n65704;
  assign n65706 = ~i_hbusreq7 & ~n65705;
  assign n65707 = ~n65700 & ~n65706;
  assign n65708 = n7924 & ~n65707;
  assign n65709 = ~n39731 & ~n65708;
  assign n65710 = ~n8214 & ~n65709;
  assign n65711 = ~n39739 & ~n65710;
  assign n65712 = n8202 & ~n65711;
  assign n65713 = ~n39729 & ~n65712;
  assign n65714 = ~n7728 & ~n65713;
  assign n65715 = ~n65694 & ~n65714;
  assign n65716 = ~n7723 & ~n65715;
  assign n65717 = ~n7723 & ~n65716;
  assign n65718 = ~n7714 & ~n65717;
  assign n65719 = ~n7714 & ~n65718;
  assign n65720 = n7705 & ~n65719;
  assign n65721 = n7723 & ~n65713;
  assign n65722 = ~n8224 & ~n39785;
  assign n65723 = controllable_hmaster1 & ~n65722;
  assign n65724 = ~n39820 & ~n65723;
  assign n65725 = ~controllable_hgrant6 & ~n65724;
  assign n65726 = ~n28736 & ~n65725;
  assign n65727 = controllable_hmaster0 & ~n65726;
  assign n65728 = ~n39914 & ~n65727;
  assign n65729 = ~controllable_hmaster3 & ~n65728;
  assign n65730 = ~n39767 & ~n65729;
  assign n65731 = i_hlock7 & ~n65730;
  assign n65732 = ~n8238 & ~n39785;
  assign n65733 = controllable_hmaster1 & ~n65732;
  assign n65734 = ~n39820 & ~n65733;
  assign n65735 = ~controllable_hgrant6 & ~n65734;
  assign n65736 = ~n28747 & ~n65735;
  assign n65737 = controllable_hmaster0 & ~n65736;
  assign n65738 = ~n39914 & ~n65737;
  assign n65739 = ~controllable_hmaster3 & ~n65738;
  assign n65740 = ~n39767 & ~n65739;
  assign n65741 = ~i_hlock7 & ~n65740;
  assign n65742 = ~n65731 & ~n65741;
  assign n65743 = i_hbusreq7 & ~n65742;
  assign n65744 = i_hbusreq8 & ~n65728;
  assign n65745 = i_hbusreq6 & ~n65724;
  assign n65746 = ~n8278 & ~n39988;
  assign n65747 = controllable_hmaster1 & ~n65746;
  assign n65748 = ~n40041 & ~n65747;
  assign n65749 = ~i_hbusreq6 & ~n65748;
  assign n65750 = ~n65745 & ~n65749;
  assign n65751 = ~controllable_hgrant6 & ~n65750;
  assign n65752 = ~n28761 & ~n65751;
  assign n65753 = controllable_hmaster0 & ~n65752;
  assign n65754 = ~n40167 & ~n65753;
  assign n65755 = ~i_hbusreq8 & ~n65754;
  assign n65756 = ~n65744 & ~n65755;
  assign n65757 = ~controllable_hmaster3 & ~n65756;
  assign n65758 = ~n39956 & ~n65757;
  assign n65759 = i_hlock7 & ~n65758;
  assign n65760 = i_hbusreq8 & ~n65738;
  assign n65761 = i_hbusreq6 & ~n65734;
  assign n65762 = ~n8310 & ~n39988;
  assign n65763 = controllable_hmaster1 & ~n65762;
  assign n65764 = ~n40041 & ~n65763;
  assign n65765 = ~i_hbusreq6 & ~n65764;
  assign n65766 = ~n65761 & ~n65765;
  assign n65767 = ~controllable_hgrant6 & ~n65766;
  assign n65768 = ~n28778 & ~n65767;
  assign n65769 = controllable_hmaster0 & ~n65768;
  assign n65770 = ~n40167 & ~n65769;
  assign n65771 = ~i_hbusreq8 & ~n65770;
  assign n65772 = ~n65760 & ~n65771;
  assign n65773 = ~controllable_hmaster3 & ~n65772;
  assign n65774 = ~n39956 & ~n65773;
  assign n65775 = ~i_hlock7 & ~n65774;
  assign n65776 = ~n65759 & ~n65775;
  assign n65777 = ~i_hbusreq7 & ~n65776;
  assign n65778 = ~n65743 & ~n65777;
  assign n65779 = n7924 & ~n65778;
  assign n65780 = ~n39731 & ~n65779;
  assign n65781 = ~n7920 & ~n65780;
  assign n65782 = n7920 & ~n65713;
  assign n65783 = ~n65781 & ~n65782;
  assign n65784 = ~n7723 & ~n65783;
  assign n65785 = ~n65721 & ~n65784;
  assign n65786 = n7714 & ~n65785;
  assign n65787 = ~n7714 & ~n65780;
  assign n65788 = ~n65786 & ~n65787;
  assign n65789 = ~n7705 & ~n65788;
  assign n65790 = ~n65720 & ~n65789;
  assign n65791 = ~n7808 & ~n65790;
  assign n65792 = ~n7920 & ~n65693;
  assign n65793 = ~n40785 & ~n65792;
  assign n65794 = n7728 & ~n65793;
  assign n65795 = ~n7920 & ~n65713;
  assign n65796 = ~n41275 & ~n65795;
  assign n65797 = ~n7728 & ~n65796;
  assign n65798 = ~n65794 & ~n65797;
  assign n65799 = ~n7723 & ~n65798;
  assign n65800 = ~n7723 & ~n65799;
  assign n65801 = ~n7714 & ~n65800;
  assign n65802 = ~n7714 & ~n65801;
  assign n65803 = n7705 & ~n65802;
  assign n65804 = ~n42700 & ~n65795;
  assign n65805 = n7728 & ~n65804;
  assign n65806 = ~n45926 & ~n65795;
  assign n65807 = ~n7728 & ~n65806;
  assign n65808 = ~n65805 & ~n65807;
  assign n65809 = n7723 & ~n65808;
  assign n65810 = ~n7723 & ~n65806;
  assign n65811 = ~n65809 & ~n65810;
  assign n65812 = n7714 & ~n65811;
  assign n65813 = n7723 & ~n65806;
  assign n65814 = ~n48003 & ~n65781;
  assign n65815 = n7728 & ~n65814;
  assign n65816 = ~n50001 & ~n65781;
  assign n65817 = ~n7728 & ~n65816;
  assign n65818 = ~n65815 & ~n65817;
  assign n65819 = ~n7723 & ~n65818;
  assign n65820 = ~n65813 & ~n65819;
  assign n65821 = ~n7714 & ~n65820;
  assign n65822 = ~n65812 & ~n65821;
  assign n65823 = ~n7705 & ~n65822;
  assign n65824 = ~n65803 & ~n65823;
  assign n65825 = n7808 & ~n65824;
  assign n65826 = ~n65791 & ~n65825;
  assign n65827 = n8195 & ~n65826;
  assign n65828 = ~n39684 & ~n65827;
  assign n65829 = ~n8193 & ~n65828;
  assign n65830 = ~n50187 & ~n65781;
  assign n65831 = ~n7723 & ~n65830;
  assign n65832 = ~n50186 & ~n65831;
  assign n65833 = n7714 & ~n65832;
  assign n65834 = ~n65787 & ~n65833;
  assign n65835 = ~n7705 & ~n65834;
  assign n65836 = ~n50185 & ~n65835;
  assign n65837 = ~n7808 & ~n65836;
  assign n65838 = ~n58400 & ~n65781;
  assign n65839 = n7728 & ~n65838;
  assign n65840 = ~n65817 & ~n65839;
  assign n65841 = ~n7723 & ~n65840;
  assign n65842 = ~n56860 & ~n65841;
  assign n65843 = ~n7714 & ~n65842;
  assign n65844 = ~n56859 & ~n65843;
  assign n65845 = ~n7705 & ~n65844;
  assign n65846 = ~n51653 & ~n65845;
  assign n65847 = n7808 & ~n65846;
  assign n65848 = ~n65837 & ~n65847;
  assign n65849 = ~n8195 & ~n65848;
  assign n65850 = ~n10430 & ~n58556;
  assign n65851 = controllable_hmaster1 & ~n65850;
  assign n65852 = ~n58591 & ~n65851;
  assign n65853 = ~controllable_hgrant6 & ~n65852;
  assign n65854 = ~n33324 & ~n65853;
  assign n65855 = controllable_hmaster0 & ~n65854;
  assign n65856 = ~n58659 & ~n65855;
  assign n65857 = ~controllable_hmaster3 & ~n65856;
  assign n65858 = ~n58538 & ~n65857;
  assign n65859 = i_hlock7 & ~n65858;
  assign n65860 = ~n10437 & ~n58556;
  assign n65861 = controllable_hmaster1 & ~n65860;
  assign n65862 = ~n58591 & ~n65861;
  assign n65863 = ~controllable_hgrant6 & ~n65862;
  assign n65864 = ~n33342 & ~n65863;
  assign n65865 = controllable_hmaster0 & ~n65864;
  assign n65866 = ~n58659 & ~n65865;
  assign n65867 = ~controllable_hmaster3 & ~n65866;
  assign n65868 = ~n58538 & ~n65867;
  assign n65869 = ~i_hlock7 & ~n65868;
  assign n65870 = ~n65859 & ~n65869;
  assign n65871 = i_hbusreq7 & ~n65870;
  assign n65872 = i_hbusreq8 & ~n65856;
  assign n65873 = i_hbusreq6 & ~n65852;
  assign n65874 = ~n10597 & ~n58735;
  assign n65875 = controllable_hmaster1 & ~n65874;
  assign n65876 = ~n58788 & ~n65875;
  assign n65877 = ~i_hbusreq6 & ~n65876;
  assign n65878 = ~n65873 & ~n65877;
  assign n65879 = ~controllable_hgrant6 & ~n65878;
  assign n65880 = ~n33363 & ~n65879;
  assign n65881 = controllable_hmaster0 & ~n65880;
  assign n65882 = ~n58891 & ~n65881;
  assign n65883 = ~i_hbusreq8 & ~n65882;
  assign n65884 = ~n65872 & ~n65883;
  assign n65885 = ~controllable_hmaster3 & ~n65884;
  assign n65886 = ~n58703 & ~n65885;
  assign n65887 = i_hlock7 & ~n65886;
  assign n65888 = i_hbusreq8 & ~n65866;
  assign n65889 = i_hbusreq6 & ~n65862;
  assign n65890 = ~n10607 & ~n58735;
  assign n65891 = controllable_hmaster1 & ~n65890;
  assign n65892 = ~n58788 & ~n65891;
  assign n65893 = ~i_hbusreq6 & ~n65892;
  assign n65894 = ~n65889 & ~n65893;
  assign n65895 = ~controllable_hgrant6 & ~n65894;
  assign n65896 = ~n33396 & ~n65895;
  assign n65897 = controllable_hmaster0 & ~n65896;
  assign n65898 = ~n58891 & ~n65897;
  assign n65899 = ~i_hbusreq8 & ~n65898;
  assign n65900 = ~n65888 & ~n65899;
  assign n65901 = ~controllable_hmaster3 & ~n65900;
  assign n65902 = ~n58703 & ~n65901;
  assign n65903 = ~i_hlock7 & ~n65902;
  assign n65904 = ~n65887 & ~n65903;
  assign n65905 = ~i_hbusreq7 & ~n65904;
  assign n65906 = ~n65871 & ~n65905;
  assign n65907 = n7924 & ~n65906;
  assign n65908 = ~n58519 & ~n65907;
  assign n65909 = n8214 & ~n65908;
  assign n65910 = n8214 & ~n65909;
  assign n65911 = n8202 & ~n65910;
  assign n65912 = ~n58446 & ~n65911;
  assign n65913 = n7728 & ~n65912;
  assign n65914 = n8214 & ~n65780;
  assign n65915 = ~n39730 & ~n65914;
  assign n65916 = n8202 & ~n65915;
  assign n65917 = ~n58923 & ~n65916;
  assign n65918 = ~n7728 & ~n65917;
  assign n65919 = ~n65913 & ~n65918;
  assign n65920 = ~n7723 & ~n65919;
  assign n65921 = ~n7723 & ~n65920;
  assign n65922 = ~n7714 & ~n65921;
  assign n65923 = ~n7714 & ~n65922;
  assign n65924 = n7705 & ~n65923;
  assign n65925 = n7723 & ~n65917;
  assign n65926 = n7920 & ~n65917;
  assign n65927 = ~n65781 & ~n65926;
  assign n65928 = ~n7723 & ~n65927;
  assign n65929 = ~n65925 & ~n65928;
  assign n65930 = n7714 & ~n65929;
  assign n65931 = ~n65787 & ~n65930;
  assign n65932 = ~n7705 & ~n65931;
  assign n65933 = ~n65924 & ~n65932;
  assign n65934 = ~n7808 & ~n65933;
  assign n65935 = ~n7920 & ~n65912;
  assign n65936 = ~n60195 & ~n65935;
  assign n65937 = n7728 & ~n65936;
  assign n65938 = ~n7920 & ~n65917;
  assign n65939 = ~n60612 & ~n65938;
  assign n65940 = ~n7728 & ~n65939;
  assign n65941 = ~n65937 & ~n65940;
  assign n65942 = ~n7723 & ~n65941;
  assign n65943 = ~n7723 & ~n65942;
  assign n65944 = ~n7714 & ~n65943;
  assign n65945 = ~n7714 & ~n65944;
  assign n65946 = n7705 & ~n65945;
  assign n65947 = ~n61600 & ~n65938;
  assign n65948 = n7728 & ~n65947;
  assign n65949 = ~n63732 & ~n65938;
  assign n65950 = ~n7728 & ~n65949;
  assign n65951 = ~n65948 & ~n65950;
  assign n65952 = n7723 & ~n65951;
  assign n65953 = ~n7723 & ~n65949;
  assign n65954 = ~n65952 & ~n65953;
  assign n65955 = n7714 & ~n65954;
  assign n65956 = n7723 & ~n65949;
  assign n65957 = ~n64928 & ~n65781;
  assign n65958 = n7728 & ~n65957;
  assign n65959 = ~n65817 & ~n65958;
  assign n65960 = ~n7723 & ~n65959;
  assign n65961 = ~n65956 & ~n65960;
  assign n65962 = ~n7714 & ~n65961;
  assign n65963 = ~n65955 & ~n65962;
  assign n65964 = ~n7705 & ~n65963;
  assign n65965 = ~n65946 & ~n65964;
  assign n65966 = n7808 & ~n65965;
  assign n65967 = ~n65934 & ~n65966;
  assign n65968 = n8195 & ~n65967;
  assign n65969 = ~n65849 & ~n65968;
  assign n65970 = n8193 & ~n65969;
  assign n65971 = ~n65829 & ~n65970;
  assign n65972 = n8191 & ~n65971;
  assign n65973 = ~n10989 & ~n65692;
  assign n65974 = n7728 & ~n65973;
  assign n65975 = ~n64981 & ~n65712;
  assign n65976 = ~n7728 & ~n65975;
  assign n65977 = ~n65974 & ~n65976;
  assign n65978 = ~n7723 & ~n65977;
  assign n65979 = ~n7723 & ~n65978;
  assign n65980 = ~n7714 & ~n65979;
  assign n65981 = ~n7714 & ~n65980;
  assign n65982 = n7705 & ~n65981;
  assign n65983 = n7723 & ~n65975;
  assign n65984 = ~n64999 & ~n65729;
  assign n65985 = i_hlock7 & ~n65984;
  assign n65986 = ~n64999 & ~n65739;
  assign n65987 = ~i_hlock7 & ~n65986;
  assign n65988 = ~n65985 & ~n65987;
  assign n65989 = i_hbusreq7 & ~n65988;
  assign n65990 = ~n65016 & ~n65757;
  assign n65991 = i_hlock7 & ~n65990;
  assign n65992 = ~n65016 & ~n65773;
  assign n65993 = ~i_hlock7 & ~n65992;
  assign n65994 = ~n65991 & ~n65993;
  assign n65995 = ~i_hbusreq7 & ~n65994;
  assign n65996 = ~n65989 & ~n65995;
  assign n65997 = n7924 & ~n65996;
  assign n65998 = ~n39731 & ~n65997;
  assign n65999 = ~n7920 & ~n65998;
  assign n66000 = n7920 & ~n65975;
  assign n66001 = ~n65999 & ~n66000;
  assign n66002 = ~n7723 & ~n66001;
  assign n66003 = ~n65983 & ~n66002;
  assign n66004 = n7714 & ~n66003;
  assign n66005 = ~n7714 & ~n65998;
  assign n66006 = ~n66004 & ~n66005;
  assign n66007 = ~n7705 & ~n66006;
  assign n66008 = ~n65982 & ~n66007;
  assign n66009 = ~n7808 & ~n66008;
  assign n66010 = ~n7920 & ~n65973;
  assign n66011 = ~n40785 & ~n66010;
  assign n66012 = n7728 & ~n66011;
  assign n66013 = ~n7920 & ~n65975;
  assign n66014 = ~n41275 & ~n66013;
  assign n66015 = ~n7728 & ~n66014;
  assign n66016 = ~n66012 & ~n66015;
  assign n66017 = ~n7723 & ~n66016;
  assign n66018 = ~n7723 & ~n66017;
  assign n66019 = ~n7714 & ~n66018;
  assign n66020 = ~n7714 & ~n66019;
  assign n66021 = n7705 & ~n66020;
  assign n66022 = ~n42700 & ~n66013;
  assign n66023 = n7728 & ~n66022;
  assign n66024 = ~n45926 & ~n66013;
  assign n66025 = ~n7728 & ~n66024;
  assign n66026 = ~n66023 & ~n66025;
  assign n66027 = n7723 & ~n66026;
  assign n66028 = ~n7723 & ~n66024;
  assign n66029 = ~n66027 & ~n66028;
  assign n66030 = n7714 & ~n66029;
  assign n66031 = n7723 & ~n66024;
  assign n66032 = ~n48003 & ~n65999;
  assign n66033 = n7728 & ~n66032;
  assign n66034 = ~n50001 & ~n65999;
  assign n66035 = ~n7728 & ~n66034;
  assign n66036 = ~n66033 & ~n66035;
  assign n66037 = ~n7723 & ~n66036;
  assign n66038 = ~n66031 & ~n66037;
  assign n66039 = ~n7714 & ~n66038;
  assign n66040 = ~n66030 & ~n66039;
  assign n66041 = ~n7705 & ~n66040;
  assign n66042 = ~n66021 & ~n66041;
  assign n66043 = n7808 & ~n66042;
  assign n66044 = ~n66009 & ~n66043;
  assign n66045 = n8195 & ~n66044;
  assign n66046 = ~n39684 & ~n66045;
  assign n66047 = ~n8193 & ~n66046;
  assign n66048 = ~n50187 & ~n65999;
  assign n66049 = ~n7723 & ~n66048;
  assign n66050 = ~n50186 & ~n66049;
  assign n66051 = n7714 & ~n66050;
  assign n66052 = ~n66005 & ~n66051;
  assign n66053 = ~n7705 & ~n66052;
  assign n66054 = ~n50185 & ~n66053;
  assign n66055 = ~n7808 & ~n66054;
  assign n66056 = ~n58400 & ~n65999;
  assign n66057 = n7728 & ~n66056;
  assign n66058 = ~n66035 & ~n66057;
  assign n66059 = ~n7723 & ~n66058;
  assign n66060 = ~n56860 & ~n66059;
  assign n66061 = ~n7714 & ~n66060;
  assign n66062 = ~n56859 & ~n66061;
  assign n66063 = ~n7705 & ~n66062;
  assign n66064 = ~n51653 & ~n66063;
  assign n66065 = n7808 & ~n66064;
  assign n66066 = ~n66055 & ~n66065;
  assign n66067 = ~n8195 & ~n66066;
  assign n66068 = ~n65099 & ~n65857;
  assign n66069 = i_hlock7 & ~n66068;
  assign n66070 = ~n65099 & ~n65867;
  assign n66071 = ~i_hlock7 & ~n66070;
  assign n66072 = ~n66069 & ~n66071;
  assign n66073 = i_hbusreq7 & ~n66072;
  assign n66074 = ~n65116 & ~n65885;
  assign n66075 = i_hlock7 & ~n66074;
  assign n66076 = ~n65116 & ~n65901;
  assign n66077 = ~i_hlock7 & ~n66076;
  assign n66078 = ~n66075 & ~n66077;
  assign n66079 = ~i_hbusreq7 & ~n66078;
  assign n66080 = ~n66073 & ~n66079;
  assign n66081 = n7924 & ~n66080;
  assign n66082 = ~n58519 & ~n66081;
  assign n66083 = n8214 & ~n66082;
  assign n66084 = n8214 & ~n66083;
  assign n66085 = n8202 & ~n66084;
  assign n66086 = ~n58446 & ~n66085;
  assign n66087 = n7728 & ~n66086;
  assign n66088 = n8214 & ~n65998;
  assign n66089 = ~n39730 & ~n66088;
  assign n66090 = n8202 & ~n66089;
  assign n66091 = ~n58923 & ~n66090;
  assign n66092 = ~n7728 & ~n66091;
  assign n66093 = ~n66087 & ~n66092;
  assign n66094 = ~n7723 & ~n66093;
  assign n66095 = ~n7723 & ~n66094;
  assign n66096 = ~n7714 & ~n66095;
  assign n66097 = ~n7714 & ~n66096;
  assign n66098 = n7705 & ~n66097;
  assign n66099 = n7723 & ~n66091;
  assign n66100 = n7920 & ~n66091;
  assign n66101 = ~n65999 & ~n66100;
  assign n66102 = ~n7723 & ~n66101;
  assign n66103 = ~n66099 & ~n66102;
  assign n66104 = n7714 & ~n66103;
  assign n66105 = ~n66005 & ~n66104;
  assign n66106 = ~n7705 & ~n66105;
  assign n66107 = ~n66098 & ~n66106;
  assign n66108 = ~n7808 & ~n66107;
  assign n66109 = ~n7920 & ~n66086;
  assign n66110 = ~n60195 & ~n66109;
  assign n66111 = n7728 & ~n66110;
  assign n66112 = ~n7920 & ~n66091;
  assign n66113 = ~n60612 & ~n66112;
  assign n66114 = ~n7728 & ~n66113;
  assign n66115 = ~n66111 & ~n66114;
  assign n66116 = ~n7723 & ~n66115;
  assign n66117 = ~n7723 & ~n66116;
  assign n66118 = ~n7714 & ~n66117;
  assign n66119 = ~n7714 & ~n66118;
  assign n66120 = n7705 & ~n66119;
  assign n66121 = ~n61600 & ~n66112;
  assign n66122 = n7728 & ~n66121;
  assign n66123 = ~n63732 & ~n66112;
  assign n66124 = ~n7728 & ~n66123;
  assign n66125 = ~n66122 & ~n66124;
  assign n66126 = n7723 & ~n66125;
  assign n66127 = ~n7723 & ~n66123;
  assign n66128 = ~n66126 & ~n66127;
  assign n66129 = n7714 & ~n66128;
  assign n66130 = n7723 & ~n66123;
  assign n66131 = ~n64928 & ~n65999;
  assign n66132 = n7728 & ~n66131;
  assign n66133 = ~n66035 & ~n66132;
  assign n66134 = ~n7723 & ~n66133;
  assign n66135 = ~n66130 & ~n66134;
  assign n66136 = ~n7714 & ~n66135;
  assign n66137 = ~n66129 & ~n66136;
  assign n66138 = ~n7705 & ~n66137;
  assign n66139 = ~n66120 & ~n66138;
  assign n66140 = n7808 & ~n66139;
  assign n66141 = ~n66108 & ~n66140;
  assign n66142 = n8195 & ~n66141;
  assign n66143 = ~n66067 & ~n66142;
  assign n66144 = n8193 & ~n66143;
  assign n66145 = ~n66047 & ~n66144;
  assign n66146 = ~n8191 & ~n66145;
  assign n66147 = ~n65972 & ~n66146;
  assign n66148 = n8188 & ~n66147;
  assign n66149 = ~n11286 & ~n65692;
  assign n66150 = n7728 & ~n66149;
  assign n66151 = ~n65246 & ~n65712;
  assign n66152 = ~n7728 & ~n66151;
  assign n66153 = ~n66150 & ~n66152;
  assign n66154 = ~n7723 & ~n66153;
  assign n66155 = ~n7723 & ~n66154;
  assign n66156 = ~n7714 & ~n66155;
  assign n66157 = ~n7714 & ~n66156;
  assign n66158 = n7705 & ~n66157;
  assign n66159 = n7723 & ~n66151;
  assign n66160 = ~n65274 & ~n65729;
  assign n66161 = i_hlock7 & ~n66160;
  assign n66162 = ~n65274 & ~n65739;
  assign n66163 = ~i_hlock7 & ~n66162;
  assign n66164 = ~n66161 & ~n66163;
  assign n66165 = i_hbusreq7 & ~n66164;
  assign n66166 = ~n65304 & ~n65757;
  assign n66167 = i_hlock7 & ~n66166;
  assign n66168 = ~n65304 & ~n65773;
  assign n66169 = ~i_hlock7 & ~n66168;
  assign n66170 = ~n66167 & ~n66169;
  assign n66171 = ~i_hbusreq7 & ~n66170;
  assign n66172 = ~n66165 & ~n66171;
  assign n66173 = n7924 & ~n66172;
  assign n66174 = ~n39731 & ~n66173;
  assign n66175 = ~n7920 & ~n66174;
  assign n66176 = n7920 & ~n66151;
  assign n66177 = ~n66175 & ~n66176;
  assign n66178 = ~n7723 & ~n66177;
  assign n66179 = ~n66159 & ~n66178;
  assign n66180 = n7714 & ~n66179;
  assign n66181 = ~n7714 & ~n66174;
  assign n66182 = ~n66180 & ~n66181;
  assign n66183 = ~n7705 & ~n66182;
  assign n66184 = ~n66158 & ~n66183;
  assign n66185 = ~n7808 & ~n66184;
  assign n66186 = ~n7920 & ~n66149;
  assign n66187 = ~n40785 & ~n66186;
  assign n66188 = n7728 & ~n66187;
  assign n66189 = ~n7920 & ~n66151;
  assign n66190 = ~n41275 & ~n66189;
  assign n66191 = ~n7728 & ~n66190;
  assign n66192 = ~n66188 & ~n66191;
  assign n66193 = ~n7723 & ~n66192;
  assign n66194 = ~n7723 & ~n66193;
  assign n66195 = ~n7714 & ~n66194;
  assign n66196 = ~n7714 & ~n66195;
  assign n66197 = n7705 & ~n66196;
  assign n66198 = ~n42700 & ~n66189;
  assign n66199 = n7728 & ~n66198;
  assign n66200 = ~n45926 & ~n66189;
  assign n66201 = ~n7728 & ~n66200;
  assign n66202 = ~n66199 & ~n66201;
  assign n66203 = n7723 & ~n66202;
  assign n66204 = ~n7723 & ~n66200;
  assign n66205 = ~n66203 & ~n66204;
  assign n66206 = n7714 & ~n66205;
  assign n66207 = n7723 & ~n66200;
  assign n66208 = ~n48003 & ~n66175;
  assign n66209 = n7728 & ~n66208;
  assign n66210 = ~n50001 & ~n66175;
  assign n66211 = ~n7728 & ~n66210;
  assign n66212 = ~n66209 & ~n66211;
  assign n66213 = ~n7723 & ~n66212;
  assign n66214 = ~n66207 & ~n66213;
  assign n66215 = ~n7714 & ~n66214;
  assign n66216 = ~n66206 & ~n66215;
  assign n66217 = ~n7705 & ~n66216;
  assign n66218 = ~n66197 & ~n66217;
  assign n66219 = n7808 & ~n66218;
  assign n66220 = ~n66185 & ~n66219;
  assign n66221 = n8195 & ~n66220;
  assign n66222 = ~n39684 & ~n66221;
  assign n66223 = ~n8193 & ~n66222;
  assign n66224 = ~n50187 & ~n66175;
  assign n66225 = ~n7723 & ~n66224;
  assign n66226 = ~n50186 & ~n66225;
  assign n66227 = n7714 & ~n66226;
  assign n66228 = ~n66181 & ~n66227;
  assign n66229 = ~n7705 & ~n66228;
  assign n66230 = ~n50185 & ~n66229;
  assign n66231 = ~n7808 & ~n66230;
  assign n66232 = ~n58400 & ~n66175;
  assign n66233 = n7728 & ~n66232;
  assign n66234 = ~n66211 & ~n66233;
  assign n66235 = ~n7723 & ~n66234;
  assign n66236 = ~n56860 & ~n66235;
  assign n66237 = ~n7714 & ~n66236;
  assign n66238 = ~n56859 & ~n66237;
  assign n66239 = ~n7705 & ~n66238;
  assign n66240 = ~n51653 & ~n66239;
  assign n66241 = n7808 & ~n66240;
  assign n66242 = ~n66231 & ~n66241;
  assign n66243 = ~n8195 & ~n66242;
  assign n66244 = ~n65397 & ~n65857;
  assign n66245 = i_hlock7 & ~n66244;
  assign n66246 = ~n65397 & ~n65867;
  assign n66247 = ~i_hlock7 & ~n66246;
  assign n66248 = ~n66245 & ~n66247;
  assign n66249 = i_hbusreq7 & ~n66248;
  assign n66250 = ~n65427 & ~n65885;
  assign n66251 = i_hlock7 & ~n66250;
  assign n66252 = ~n65427 & ~n65901;
  assign n66253 = ~i_hlock7 & ~n66252;
  assign n66254 = ~n66251 & ~n66253;
  assign n66255 = ~i_hbusreq7 & ~n66254;
  assign n66256 = ~n66249 & ~n66255;
  assign n66257 = n7924 & ~n66256;
  assign n66258 = ~n58519 & ~n66257;
  assign n66259 = n8214 & ~n66258;
  assign n66260 = n8214 & ~n66259;
  assign n66261 = n8202 & ~n66260;
  assign n66262 = ~n58446 & ~n66261;
  assign n66263 = n7728 & ~n66262;
  assign n66264 = n8214 & ~n66174;
  assign n66265 = ~n39730 & ~n66264;
  assign n66266 = n8202 & ~n66265;
  assign n66267 = ~n58923 & ~n66266;
  assign n66268 = ~n7728 & ~n66267;
  assign n66269 = ~n66263 & ~n66268;
  assign n66270 = ~n7723 & ~n66269;
  assign n66271 = ~n7723 & ~n66270;
  assign n66272 = ~n7714 & ~n66271;
  assign n66273 = ~n7714 & ~n66272;
  assign n66274 = n7705 & ~n66273;
  assign n66275 = n7723 & ~n66267;
  assign n66276 = n7920 & ~n66267;
  assign n66277 = ~n66175 & ~n66276;
  assign n66278 = ~n7723 & ~n66277;
  assign n66279 = ~n66275 & ~n66278;
  assign n66280 = n7714 & ~n66279;
  assign n66281 = ~n66181 & ~n66280;
  assign n66282 = ~n7705 & ~n66281;
  assign n66283 = ~n66274 & ~n66282;
  assign n66284 = ~n7808 & ~n66283;
  assign n66285 = ~n7920 & ~n66262;
  assign n66286 = ~n60195 & ~n66285;
  assign n66287 = n7728 & ~n66286;
  assign n66288 = ~n7920 & ~n66267;
  assign n66289 = ~n60612 & ~n66288;
  assign n66290 = ~n7728 & ~n66289;
  assign n66291 = ~n66287 & ~n66290;
  assign n66292 = ~n7723 & ~n66291;
  assign n66293 = ~n7723 & ~n66292;
  assign n66294 = ~n7714 & ~n66293;
  assign n66295 = ~n7714 & ~n66294;
  assign n66296 = n7705 & ~n66295;
  assign n66297 = ~n61600 & ~n66288;
  assign n66298 = n7728 & ~n66297;
  assign n66299 = ~n63732 & ~n66288;
  assign n66300 = ~n7728 & ~n66299;
  assign n66301 = ~n66298 & ~n66300;
  assign n66302 = n7723 & ~n66301;
  assign n66303 = ~n7723 & ~n66299;
  assign n66304 = ~n66302 & ~n66303;
  assign n66305 = n7714 & ~n66304;
  assign n66306 = n7723 & ~n66299;
  assign n66307 = ~n64928 & ~n66175;
  assign n66308 = n7728 & ~n66307;
  assign n66309 = ~n66211 & ~n66308;
  assign n66310 = ~n7723 & ~n66309;
  assign n66311 = ~n66306 & ~n66310;
  assign n66312 = ~n7714 & ~n66311;
  assign n66313 = ~n66305 & ~n66312;
  assign n66314 = ~n7705 & ~n66313;
  assign n66315 = ~n66296 & ~n66314;
  assign n66316 = n7808 & ~n66315;
  assign n66317 = ~n66284 & ~n66316;
  assign n66318 = n8195 & ~n66317;
  assign n66319 = ~n66243 & ~n66318;
  assign n66320 = n8193 & ~n66319;
  assign n66321 = ~n66223 & ~n66320;
  assign n66322 = n8191 & ~n66321;
  assign n66323 = ~n11575 & ~n65692;
  assign n66324 = n7728 & ~n66323;
  assign n66325 = ~n65500 & ~n65712;
  assign n66326 = ~n7728 & ~n66325;
  assign n66327 = ~n66324 & ~n66326;
  assign n66328 = ~n7723 & ~n66327;
  assign n66329 = ~n7723 & ~n66328;
  assign n66330 = ~n7714 & ~n66329;
  assign n66331 = ~n7714 & ~n66330;
  assign n66332 = n7705 & ~n66331;
  assign n66333 = n7723 & ~n66325;
  assign n66334 = ~n65515 & ~n65729;
  assign n66335 = i_hlock7 & ~n66334;
  assign n66336 = ~n65515 & ~n65739;
  assign n66337 = ~i_hlock7 & ~n66336;
  assign n66338 = ~n66335 & ~n66337;
  assign n66339 = i_hbusreq7 & ~n66338;
  assign n66340 = ~n65526 & ~n65757;
  assign n66341 = i_hlock7 & ~n66340;
  assign n66342 = ~n65526 & ~n65773;
  assign n66343 = ~i_hlock7 & ~n66342;
  assign n66344 = ~n66341 & ~n66343;
  assign n66345 = ~i_hbusreq7 & ~n66344;
  assign n66346 = ~n66339 & ~n66345;
  assign n66347 = n7924 & ~n66346;
  assign n66348 = ~n39731 & ~n66347;
  assign n66349 = ~n7920 & ~n66348;
  assign n66350 = n7920 & ~n66325;
  assign n66351 = ~n66349 & ~n66350;
  assign n66352 = ~n7723 & ~n66351;
  assign n66353 = ~n66333 & ~n66352;
  assign n66354 = n7714 & ~n66353;
  assign n66355 = ~n7714 & ~n66348;
  assign n66356 = ~n66354 & ~n66355;
  assign n66357 = ~n7705 & ~n66356;
  assign n66358 = ~n66332 & ~n66357;
  assign n66359 = ~n7808 & ~n66358;
  assign n66360 = ~n7920 & ~n66323;
  assign n66361 = ~n40785 & ~n66360;
  assign n66362 = n7728 & ~n66361;
  assign n66363 = ~n7920 & ~n66325;
  assign n66364 = ~n41275 & ~n66363;
  assign n66365 = ~n7728 & ~n66364;
  assign n66366 = ~n66362 & ~n66365;
  assign n66367 = ~n7723 & ~n66366;
  assign n66368 = ~n7723 & ~n66367;
  assign n66369 = ~n7714 & ~n66368;
  assign n66370 = ~n7714 & ~n66369;
  assign n66371 = n7705 & ~n66370;
  assign n66372 = ~n42700 & ~n66363;
  assign n66373 = n7728 & ~n66372;
  assign n66374 = ~n45926 & ~n66363;
  assign n66375 = ~n7728 & ~n66374;
  assign n66376 = ~n66373 & ~n66375;
  assign n66377 = n7723 & ~n66376;
  assign n66378 = ~n7723 & ~n66374;
  assign n66379 = ~n66377 & ~n66378;
  assign n66380 = n7714 & ~n66379;
  assign n66381 = n7723 & ~n66374;
  assign n66382 = ~n48003 & ~n66349;
  assign n66383 = n7728 & ~n66382;
  assign n66384 = ~n50001 & ~n66349;
  assign n66385 = ~n7728 & ~n66384;
  assign n66386 = ~n66383 & ~n66385;
  assign n66387 = ~n7723 & ~n66386;
  assign n66388 = ~n66381 & ~n66387;
  assign n66389 = ~n7714 & ~n66388;
  assign n66390 = ~n66380 & ~n66389;
  assign n66391 = ~n7705 & ~n66390;
  assign n66392 = ~n66371 & ~n66391;
  assign n66393 = n7808 & ~n66392;
  assign n66394 = ~n66359 & ~n66393;
  assign n66395 = n8195 & ~n66394;
  assign n66396 = ~n39684 & ~n66395;
  assign n66397 = ~n8193 & ~n66396;
  assign n66398 = ~n50187 & ~n66349;
  assign n66399 = ~n7723 & ~n66398;
  assign n66400 = ~n50186 & ~n66399;
  assign n66401 = n7714 & ~n66400;
  assign n66402 = ~n66355 & ~n66401;
  assign n66403 = ~n7705 & ~n66402;
  assign n66404 = ~n50185 & ~n66403;
  assign n66405 = ~n7808 & ~n66404;
  assign n66406 = ~n58400 & ~n66349;
  assign n66407 = n7728 & ~n66406;
  assign n66408 = ~n66385 & ~n66407;
  assign n66409 = ~n7723 & ~n66408;
  assign n66410 = ~n56860 & ~n66409;
  assign n66411 = ~n7714 & ~n66410;
  assign n66412 = ~n56859 & ~n66411;
  assign n66413 = ~n7705 & ~n66412;
  assign n66414 = ~n51653 & ~n66413;
  assign n66415 = n7808 & ~n66414;
  assign n66416 = ~n66405 & ~n66415;
  assign n66417 = ~n8195 & ~n66416;
  assign n66418 = ~n65606 & ~n65857;
  assign n66419 = i_hlock7 & ~n66418;
  assign n66420 = ~n65606 & ~n65867;
  assign n66421 = ~i_hlock7 & ~n66420;
  assign n66422 = ~n66419 & ~n66421;
  assign n66423 = i_hbusreq7 & ~n66422;
  assign n66424 = ~n65617 & ~n65885;
  assign n66425 = i_hlock7 & ~n66424;
  assign n66426 = ~n65617 & ~n65901;
  assign n66427 = ~i_hlock7 & ~n66426;
  assign n66428 = ~n66425 & ~n66427;
  assign n66429 = ~i_hbusreq7 & ~n66428;
  assign n66430 = ~n66423 & ~n66429;
  assign n66431 = n7924 & ~n66430;
  assign n66432 = ~n58519 & ~n66431;
  assign n66433 = n8214 & ~n66432;
  assign n66434 = n8214 & ~n66433;
  assign n66435 = n8202 & ~n66434;
  assign n66436 = ~n58446 & ~n66435;
  assign n66437 = n7728 & ~n66436;
  assign n66438 = n8214 & ~n66348;
  assign n66439 = ~n39730 & ~n66438;
  assign n66440 = n8202 & ~n66439;
  assign n66441 = ~n58923 & ~n66440;
  assign n66442 = ~n7728 & ~n66441;
  assign n66443 = ~n66437 & ~n66442;
  assign n66444 = ~n7723 & ~n66443;
  assign n66445 = ~n7723 & ~n66444;
  assign n66446 = ~n7714 & ~n66445;
  assign n66447 = ~n7714 & ~n66446;
  assign n66448 = n7705 & ~n66447;
  assign n66449 = n7723 & ~n66441;
  assign n66450 = n7920 & ~n66441;
  assign n66451 = ~n66349 & ~n66450;
  assign n66452 = ~n7723 & ~n66451;
  assign n66453 = ~n66449 & ~n66452;
  assign n66454 = n7714 & ~n66453;
  assign n66455 = ~n66355 & ~n66454;
  assign n66456 = ~n7705 & ~n66455;
  assign n66457 = ~n66448 & ~n66456;
  assign n66458 = ~n7808 & ~n66457;
  assign n66459 = ~n7920 & ~n66436;
  assign n66460 = ~n60195 & ~n66459;
  assign n66461 = n7728 & ~n66460;
  assign n66462 = ~n7920 & ~n66441;
  assign n66463 = ~n60612 & ~n66462;
  assign n66464 = ~n7728 & ~n66463;
  assign n66465 = ~n66461 & ~n66464;
  assign n66466 = ~n7723 & ~n66465;
  assign n66467 = ~n7723 & ~n66466;
  assign n66468 = ~n7714 & ~n66467;
  assign n66469 = ~n7714 & ~n66468;
  assign n66470 = n7705 & ~n66469;
  assign n66471 = ~n61600 & ~n66462;
  assign n66472 = n7728 & ~n66471;
  assign n66473 = ~n63732 & ~n66462;
  assign n66474 = ~n7728 & ~n66473;
  assign n66475 = ~n66472 & ~n66474;
  assign n66476 = n7723 & ~n66475;
  assign n66477 = ~n7723 & ~n66473;
  assign n66478 = ~n66476 & ~n66477;
  assign n66479 = n7714 & ~n66478;
  assign n66480 = n7723 & ~n66473;
  assign n66481 = ~n64928 & ~n66349;
  assign n66482 = n7728 & ~n66481;
  assign n66483 = ~n66385 & ~n66482;
  assign n66484 = ~n7723 & ~n66483;
  assign n66485 = ~n66480 & ~n66484;
  assign n66486 = ~n7714 & ~n66485;
  assign n66487 = ~n66479 & ~n66486;
  assign n66488 = ~n7705 & ~n66487;
  assign n66489 = ~n66470 & ~n66488;
  assign n66490 = n7808 & ~n66489;
  assign n66491 = ~n66458 & ~n66490;
  assign n66492 = n8195 & ~n66491;
  assign n66493 = ~n66417 & ~n66492;
  assign n66494 = n8193 & ~n66493;
  assign n66495 = ~n66397 & ~n66494;
  assign n66496 = ~n8191 & ~n66495;
  assign n66497 = ~n66322 & ~n66496;
  assign n66498 = ~n8188 & ~n66497;
  assign n66499 = ~n66148 & ~n66498;
  assign n66500 = ~n8185 & ~n66499;
  assign n66501 = ~n65690 & ~n66500;
  assign n66502 = ~controllable_hgrant8 & ~n66501;
  assign n66503 = ~n39683 & ~n66502;
  assign n66504 = controllable_nhgrant0 & ~n66503;
  assign n66505 = controllable_hgrant6 & ~n8460;
  assign n66506 = controllable_hgrant5 & ~n8442;
  assign n66507 = controllable_hgrant4 & ~n8442;
  assign n66508 = controllable_hgrant3 & ~n8442;
  assign n66509 = controllable_hgrant1 & ~n8442;
  assign n66510 = controllable_hgrant2 & ~n8437;
  assign n66511 = i_hlock0 & ~n16123;
  assign n66512 = ~i_hlock0 & ~n16141;
  assign n66513 = ~n66511 & ~n66512;
  assign n66514 = ~controllable_hgrant2 & n66513;
  assign n66515 = ~n66510 & ~n66514;
  assign n66516 = ~n7733 & ~n66515;
  assign n66517 = ~n7733 & ~n66516;
  assign n66518 = ~n7928 & ~n66517;
  assign n66519 = n7928 & ~n66515;
  assign n66520 = ~n66518 & ~n66519;
  assign n66521 = ~controllable_hgrant1 & ~n66520;
  assign n66522 = ~n66509 & ~n66521;
  assign n66523 = ~controllable_hgrant3 & ~n66522;
  assign n66524 = ~n66508 & ~n66523;
  assign n66525 = ~controllable_hgrant4 & ~n66524;
  assign n66526 = ~n66507 & ~n66525;
  assign n66527 = ~controllable_hgrant5 & ~n66526;
  assign n66528 = ~n66506 & ~n66527;
  assign n66529 = ~controllable_hmaster2 & ~n66528;
  assign n66530 = ~n8434 & ~n66529;
  assign n66531 = ~controllable_hmaster1 & ~n66530;
  assign n66532 = ~n8423 & ~n66531;
  assign n66533 = n8217 & ~n66532;
  assign n66534 = ~n8449 & ~n66531;
  assign n66535 = ~n8217 & ~n66534;
  assign n66536 = ~n66533 & ~n66535;
  assign n66537 = i_hlock6 & ~n66536;
  assign n66538 = ~n8455 & ~n66531;
  assign n66539 = ~n8217 & ~n66538;
  assign n66540 = ~n66533 & ~n66539;
  assign n66541 = ~i_hlock6 & ~n66540;
  assign n66542 = ~n66537 & ~n66541;
  assign n66543 = ~controllable_hgrant6 & ~n66542;
  assign n66544 = ~n66505 & ~n66543;
  assign n66545 = ~controllable_hmaster0 & ~n66544;
  assign n66546 = ~n8401 & ~n66545;
  assign n66547 = ~controllable_hmaster3 & ~n66546;
  assign n66548 = ~n8362 & ~n66547;
  assign n66549 = i_hbusreq7 & ~n66548;
  assign n66550 = i_hbusreq8 & ~n66546;
  assign n66551 = controllable_hgrant6 & ~n8629;
  assign n66552 = i_hbusreq6 & ~n66542;
  assign n66553 = ~n8610 & ~n66529;
  assign n66554 = ~controllable_hmaster1 & ~n66553;
  assign n66555 = ~n8590 & ~n66554;
  assign n66556 = n8217 & ~n66555;
  assign n66557 = ~n8616 & ~n66554;
  assign n66558 = ~n8217 & ~n66557;
  assign n66559 = ~n66556 & ~n66558;
  assign n66560 = i_hlock6 & ~n66559;
  assign n66561 = ~n8622 & ~n66554;
  assign n66562 = ~n8217 & ~n66561;
  assign n66563 = ~n66556 & ~n66562;
  assign n66564 = ~i_hlock6 & ~n66563;
  assign n66565 = ~n66560 & ~n66564;
  assign n66566 = ~i_hbusreq6 & ~n66565;
  assign n66567 = ~n66552 & ~n66566;
  assign n66568 = ~controllable_hgrant6 & ~n66567;
  assign n66569 = ~n66551 & ~n66568;
  assign n66570 = ~controllable_hmaster0 & ~n66569;
  assign n66571 = ~n8556 & ~n66570;
  assign n66572 = ~i_hbusreq8 & ~n66571;
  assign n66573 = ~n66550 & ~n66572;
  assign n66574 = ~controllable_hmaster3 & ~n66573;
  assign n66575 = ~n8492 & ~n66574;
  assign n66576 = ~i_hbusreq7 & ~n66575;
  assign n66577 = ~n66549 & ~n66576;
  assign n66578 = n7924 & ~n66577;
  assign n66579 = ~n8337 & ~n66578;
  assign n66580 = ~n7920 & ~n66579;
  assign n66581 = ~n8641 & ~n66580;
  assign n66582 = ~n7723 & ~n66581;
  assign n66583 = ~n8356 & ~n66582;
  assign n66584 = n7714 & ~n66583;
  assign n66585 = ~n7714 & ~n66579;
  assign n66586 = ~n66584 & ~n66585;
  assign n66587 = ~n7705 & ~n66586;
  assign n66588 = ~n8355 & ~n66587;
  assign n66589 = ~n7808 & ~n66588;
  assign n66590 = ~n16992 & ~n28865;
  assign n66591 = n7920 & ~n66590;
  assign n66592 = ~n8651 & ~n66591;
  assign n66593 = n7728 & ~n66592;
  assign n66594 = ~n17303 & ~n29166;
  assign n66595 = n7920 & ~n66594;
  assign n66596 = ~n8877 & ~n66595;
  assign n66597 = ~n7728 & ~n66596;
  assign n66598 = ~n66593 & ~n66597;
  assign n66599 = ~n7723 & ~n66598;
  assign n66600 = ~n7723 & ~n66599;
  assign n66601 = ~n7714 & ~n66600;
  assign n66602 = ~n7714 & ~n66601;
  assign n66603 = n7705 & ~n66602;
  assign n66604 = ~controllable_hmaster3 & ~n36101;
  assign n66605 = ~n29298 & ~n66604;
  assign n66606 = i_hbusreq7 & ~n66605;
  assign n66607 = ~n10116 & ~n13369;
  assign n66608 = ~controllable_hmaster1 & ~n66607;
  assign n66609 = ~n10064 & ~n66608;
  assign n66610 = ~i_hbusreq6 & ~n66609;
  assign n66611 = ~n15673 & ~n66610;
  assign n66612 = ~controllable_hgrant6 & ~n66611;
  assign n66613 = ~n13298 & ~n66612;
  assign n66614 = ~controllable_hmaster0 & ~n66613;
  assign n66615 = ~n9162 & ~n66614;
  assign n66616 = ~i_hbusreq8 & ~n66615;
  assign n66617 = ~n36105 & ~n66616;
  assign n66618 = ~controllable_hmaster3 & ~n66617;
  assign n66619 = ~n29314 & ~n66618;
  assign n66620 = ~i_hbusreq7 & ~n66619;
  assign n66621 = ~n66606 & ~n66620;
  assign n66622 = ~n7924 & ~n66621;
  assign n66623 = ~controllable_hmaster3 & ~n36117;
  assign n66624 = ~n29334 & ~n66623;
  assign n66625 = i_hbusreq7 & ~n66624;
  assign n66626 = ~n13511 & ~n15308;
  assign n66627 = ~controllable_hmaster1 & ~n66626;
  assign n66628 = ~n15208 & ~n66627;
  assign n66629 = ~i_hbusreq6 & ~n66628;
  assign n66630 = ~n15726 & ~n66629;
  assign n66631 = ~controllable_hgrant6 & ~n66630;
  assign n66632 = ~n13298 & ~n66631;
  assign n66633 = ~controllable_hmaster0 & ~n66632;
  assign n66634 = ~n13778 & ~n66633;
  assign n66635 = ~i_hbusreq8 & ~n66634;
  assign n66636 = ~n36121 & ~n66635;
  assign n66637 = ~controllable_hmaster3 & ~n66636;
  assign n66638 = ~n29367 & ~n66637;
  assign n66639 = ~i_hbusreq7 & ~n66638;
  assign n66640 = ~n66625 & ~n66639;
  assign n66641 = n7924 & ~n66640;
  assign n66642 = ~n66622 & ~n66641;
  assign n66643 = ~n8214 & ~n66642;
  assign n66644 = ~n29379 & ~n66604;
  assign n66645 = i_hbusreq7 & ~n66644;
  assign n66646 = ~n29390 & ~n66618;
  assign n66647 = ~i_hbusreq7 & ~n66646;
  assign n66648 = ~n66645 & ~n66647;
  assign n66649 = ~n7924 & ~n66648;
  assign n66650 = ~n29400 & ~n66623;
  assign n66651 = i_hbusreq7 & ~n66650;
  assign n66652 = ~n29411 & ~n66637;
  assign n66653 = ~i_hbusreq7 & ~n66652;
  assign n66654 = ~n66651 & ~n66653;
  assign n66655 = n7924 & ~n66654;
  assign n66656 = ~n66649 & ~n66655;
  assign n66657 = n8214 & ~n66656;
  assign n66658 = ~n66643 & ~n66657;
  assign n66659 = ~n8202 & ~n66658;
  assign n66660 = ~n17915 & ~n36100;
  assign n66661 = ~controllable_hmaster3 & ~n66660;
  assign n66662 = ~n9093 & ~n66661;
  assign n66663 = i_hlock7 & ~n66662;
  assign n66664 = ~n17925 & ~n36100;
  assign n66665 = ~controllable_hmaster3 & ~n66664;
  assign n66666 = ~n9093 & ~n66665;
  assign n66667 = ~i_hlock7 & ~n66666;
  assign n66668 = ~n66663 & ~n66667;
  assign n66669 = i_hbusreq7 & ~n66668;
  assign n66670 = i_hbusreq8 & ~n66660;
  assign n66671 = ~n17941 & ~n66614;
  assign n66672 = ~i_hbusreq8 & ~n66671;
  assign n66673 = ~n66670 & ~n66672;
  assign n66674 = ~controllable_hmaster3 & ~n66673;
  assign n66675 = ~n9117 & ~n66674;
  assign n66676 = i_hlock7 & ~n66675;
  assign n66677 = i_hbusreq8 & ~n66664;
  assign n66678 = ~n17957 & ~n66614;
  assign n66679 = ~i_hbusreq8 & ~n66678;
  assign n66680 = ~n66677 & ~n66679;
  assign n66681 = ~controllable_hmaster3 & ~n66680;
  assign n66682 = ~n9117 & ~n66681;
  assign n66683 = ~i_hlock7 & ~n66682;
  assign n66684 = ~n66676 & ~n66683;
  assign n66685 = ~i_hbusreq7 & ~n66684;
  assign n66686 = ~n66669 & ~n66685;
  assign n66687 = ~n7924 & ~n66686;
  assign n66688 = ~n17974 & ~n36116;
  assign n66689 = ~controllable_hmaster3 & ~n66688;
  assign n66690 = ~n27088 & ~n66689;
  assign n66691 = i_hlock7 & ~n66690;
  assign n66692 = ~n17985 & ~n36116;
  assign n66693 = ~controllable_hmaster3 & ~n66692;
  assign n66694 = ~n27088 & ~n66693;
  assign n66695 = ~i_hlock7 & ~n66694;
  assign n66696 = ~n66691 & ~n66695;
  assign n66697 = i_hbusreq7 & ~n66696;
  assign n66698 = i_hbusreq8 & ~n66688;
  assign n66699 = ~n18002 & ~n66633;
  assign n66700 = ~i_hbusreq8 & ~n66699;
  assign n66701 = ~n66698 & ~n66700;
  assign n66702 = ~controllable_hmaster3 & ~n66701;
  assign n66703 = ~n27174 & ~n66702;
  assign n66704 = i_hlock7 & ~n66703;
  assign n66705 = i_hbusreq8 & ~n66692;
  assign n66706 = ~n18019 & ~n66633;
  assign n66707 = ~i_hbusreq8 & ~n66706;
  assign n66708 = ~n66705 & ~n66707;
  assign n66709 = ~controllable_hmaster3 & ~n66708;
  assign n66710 = ~n27174 & ~n66709;
  assign n66711 = ~i_hlock7 & ~n66710;
  assign n66712 = ~n66704 & ~n66711;
  assign n66713 = ~i_hbusreq7 & ~n66712;
  assign n66714 = ~n66697 & ~n66713;
  assign n66715 = n7924 & ~n66714;
  assign n66716 = ~n66687 & ~n66715;
  assign n66717 = ~n8214 & ~n66716;
  assign n66718 = ~n15662 & ~n17911;
  assign n66719 = i_hlock6 & ~n66718;
  assign n66720 = ~n15662 & ~n17921;
  assign n66721 = ~i_hlock6 & ~n66720;
  assign n66722 = ~n66719 & ~n66721;
  assign n66723 = ~controllable_hgrant6 & ~n66722;
  assign n66724 = ~n13766 & ~n66723;
  assign n66725 = ~controllable_hmaster0 & ~n66724;
  assign n66726 = ~n9152 & ~n66725;
  assign n66727 = ~controllable_hmaster3 & ~n66726;
  assign n66728 = ~n9093 & ~n66727;
  assign n66729 = i_hbusreq7 & ~n66728;
  assign n66730 = i_hbusreq8 & ~n66726;
  assign n66731 = i_hbusreq6 & ~n66722;
  assign n66732 = ~n17935 & ~n66608;
  assign n66733 = i_hlock6 & ~n66732;
  assign n66734 = ~n17951 & ~n66608;
  assign n66735 = ~i_hlock6 & ~n66734;
  assign n66736 = ~n66733 & ~n66735;
  assign n66737 = ~i_hbusreq6 & ~n66736;
  assign n66738 = ~n66731 & ~n66737;
  assign n66739 = ~controllable_hgrant6 & ~n66738;
  assign n66740 = ~n13779 & ~n66739;
  assign n66741 = ~controllable_hmaster0 & ~n66740;
  assign n66742 = ~n9162 & ~n66741;
  assign n66743 = ~i_hbusreq8 & ~n66742;
  assign n66744 = ~n66730 & ~n66743;
  assign n66745 = ~controllable_hmaster3 & ~n66744;
  assign n66746 = ~n9117 & ~n66745;
  assign n66747 = ~i_hbusreq7 & ~n66746;
  assign n66748 = ~n66729 & ~n66747;
  assign n66749 = ~n7924 & ~n66748;
  assign n66750 = ~n15716 & ~n17970;
  assign n66751 = i_hlock6 & ~n66750;
  assign n66752 = ~n15716 & ~n17981;
  assign n66753 = ~i_hlock6 & ~n66752;
  assign n66754 = ~n66751 & ~n66753;
  assign n66755 = ~controllable_hgrant6 & ~n66754;
  assign n66756 = ~n13766 & ~n66755;
  assign n66757 = ~controllable_hmaster0 & ~n66756;
  assign n66758 = ~n13765 & ~n66757;
  assign n66759 = ~controllable_hmaster3 & ~n66758;
  assign n66760 = ~n27088 & ~n66759;
  assign n66761 = i_hbusreq7 & ~n66760;
  assign n66762 = i_hbusreq8 & ~n66758;
  assign n66763 = i_hbusreq6 & ~n66754;
  assign n66764 = ~n17996 & ~n66627;
  assign n66765 = i_hlock6 & ~n66764;
  assign n66766 = ~n18013 & ~n66627;
  assign n66767 = ~i_hlock6 & ~n66766;
  assign n66768 = ~n66765 & ~n66767;
  assign n66769 = ~i_hbusreq6 & ~n66768;
  assign n66770 = ~n66763 & ~n66769;
  assign n66771 = ~controllable_hgrant6 & ~n66770;
  assign n66772 = ~n13779 & ~n66771;
  assign n66773 = ~controllable_hmaster0 & ~n66772;
  assign n66774 = ~n13778 & ~n66773;
  assign n66775 = ~i_hbusreq8 & ~n66774;
  assign n66776 = ~n66762 & ~n66775;
  assign n66777 = ~controllable_hmaster3 & ~n66776;
  assign n66778 = ~n27174 & ~n66777;
  assign n66779 = ~i_hbusreq7 & ~n66778;
  assign n66780 = ~n66761 & ~n66779;
  assign n66781 = n7924 & ~n66780;
  assign n66782 = ~n66749 & ~n66781;
  assign n66783 = n8214 & ~n66782;
  assign n66784 = ~n66717 & ~n66783;
  assign n66785 = n8202 & ~n66784;
  assign n66786 = ~n66659 & ~n66785;
  assign n66787 = n7920 & ~n66786;
  assign n66788 = ~n8877 & ~n66787;
  assign n66789 = n7728 & ~n66788;
  assign n66790 = ~n19183 & ~n66518;
  assign n66791 = ~controllable_hgrant1 & ~n66790;
  assign n66792 = ~n13924 & ~n66791;
  assign n66793 = ~controllable_hgrant3 & ~n66792;
  assign n66794 = ~n13923 & ~n66793;
  assign n66795 = ~controllable_hgrant4 & ~n66794;
  assign n66796 = ~n13922 & ~n66795;
  assign n66797 = ~controllable_hgrant5 & ~n66796;
  assign n66798 = ~n13921 & ~n66797;
  assign n66799 = ~controllable_hmaster2 & ~n66798;
  assign n66800 = ~n19299 & ~n66799;
  assign n66801 = ~controllable_hmaster1 & ~n66800;
  assign n66802 = ~n19291 & ~n66801;
  assign n66803 = i_hlock6 & ~n66802;
  assign n66804 = ~n19318 & ~n66801;
  assign n66805 = ~i_hlock6 & ~n66804;
  assign n66806 = ~n66803 & ~n66805;
  assign n66807 = ~controllable_hgrant6 & ~n66806;
  assign n66808 = ~n13894 & ~n66807;
  assign n66809 = ~controllable_hmaster0 & ~n66808;
  assign n66810 = ~n19279 & ~n66809;
  assign n66811 = ~controllable_hmaster3 & ~n66810;
  assign n66812 = ~n29730 & ~n66811;
  assign n66813 = i_hlock7 & ~n66812;
  assign n66814 = ~n19334 & ~n66809;
  assign n66815 = ~controllable_hmaster3 & ~n66814;
  assign n66816 = ~n29730 & ~n66815;
  assign n66817 = ~i_hlock7 & ~n66816;
  assign n66818 = ~n66813 & ~n66817;
  assign n66819 = i_hbusreq7 & ~n66818;
  assign n66820 = i_hbusreq8 & ~n66810;
  assign n66821 = i_hbusreq6 & ~n66806;
  assign n66822 = i_hbusreq5 & ~n66796;
  assign n66823 = i_hbusreq4 & ~n66794;
  assign n66824 = i_hbusreq9 & ~n66794;
  assign n66825 = i_hbusreq3 & ~n66792;
  assign n66826 = i_hbusreq1 & ~n66790;
  assign n66827 = ~n7860 & ~n7933;
  assign n66828 = ~controllable_locked & n66827;
  assign n66829 = ~n16120 & ~n66828;
  assign n66830 = i_hlock0 & ~n66829;
  assign n66831 = ~n16394 & ~n66830;
  assign n66832 = ~i_hbusreq0 & ~n66831;
  assign n66833 = ~n16391 & ~n66832;
  assign n66834 = ~i_hbusreq2 & ~n66833;
  assign n66835 = ~n16390 & ~n66834;
  assign n66836 = ~controllable_hgrant2 & n66835;
  assign n66837 = ~n14231 & ~n66836;
  assign n66838 = n7928 & ~n66837;
  assign n66839 = ~n66518 & ~n66838;
  assign n66840 = ~i_hbusreq1 & ~n66839;
  assign n66841 = ~n66826 & ~n66840;
  assign n66842 = ~controllable_hgrant1 & ~n66841;
  assign n66843 = ~n14229 & ~n66842;
  assign n66844 = ~i_hbusreq3 & ~n66843;
  assign n66845 = ~n66825 & ~n66844;
  assign n66846 = ~controllable_hgrant3 & ~n66845;
  assign n66847 = ~n14227 & ~n66846;
  assign n66848 = ~i_hbusreq9 & ~n66847;
  assign n66849 = ~n66824 & ~n66848;
  assign n66850 = ~i_hbusreq4 & ~n66849;
  assign n66851 = ~n66823 & ~n66850;
  assign n66852 = ~controllable_hgrant4 & ~n66851;
  assign n66853 = ~n14224 & ~n66852;
  assign n66854 = ~i_hbusreq5 & ~n66853;
  assign n66855 = ~n66822 & ~n66854;
  assign n66856 = ~controllable_hgrant5 & ~n66855;
  assign n66857 = ~n14222 & ~n66856;
  assign n66858 = ~controllable_hmaster2 & ~n66857;
  assign n66859 = ~n19598 & ~n66858;
  assign n66860 = ~controllable_hmaster1 & ~n66859;
  assign n66861 = ~n19584 & ~n66860;
  assign n66862 = i_hlock6 & ~n66861;
  assign n66863 = ~n19636 & ~n66860;
  assign n66864 = ~i_hlock6 & ~n66863;
  assign n66865 = ~n66862 & ~n66864;
  assign n66866 = ~i_hbusreq6 & ~n66865;
  assign n66867 = ~n66821 & ~n66866;
  assign n66868 = ~controllable_hgrant6 & ~n66867;
  assign n66869 = ~n14173 & ~n66868;
  assign n66870 = ~controllable_hmaster0 & ~n66869;
  assign n66871 = ~n19556 & ~n66870;
  assign n66872 = ~i_hbusreq8 & ~n66871;
  assign n66873 = ~n66820 & ~n66872;
  assign n66874 = ~controllable_hmaster3 & ~n66873;
  assign n66875 = ~n29780 & ~n66874;
  assign n66876 = i_hlock7 & ~n66875;
  assign n66877 = i_hbusreq8 & ~n66814;
  assign n66878 = ~n19660 & ~n66870;
  assign n66879 = ~i_hbusreq8 & ~n66878;
  assign n66880 = ~n66877 & ~n66879;
  assign n66881 = ~controllable_hmaster3 & ~n66880;
  assign n66882 = ~n29780 & ~n66881;
  assign n66883 = ~i_hlock7 & ~n66882;
  assign n66884 = ~n66876 & ~n66883;
  assign n66885 = ~i_hbusreq7 & ~n66884;
  assign n66886 = ~n66819 & ~n66885;
  assign n66887 = ~n7924 & ~n66886;
  assign n66888 = ~n19684 & ~n66518;
  assign n66889 = ~controllable_hgrant1 & ~n66888;
  assign n66890 = ~n13924 & ~n66889;
  assign n66891 = ~controllable_hgrant3 & ~n66890;
  assign n66892 = ~n13923 & ~n66891;
  assign n66893 = ~controllable_hgrant4 & ~n66892;
  assign n66894 = ~n13922 & ~n66893;
  assign n66895 = ~controllable_hgrant5 & ~n66894;
  assign n66896 = ~n13921 & ~n66895;
  assign n66897 = ~controllable_hmaster2 & ~n66896;
  assign n66898 = ~n19824 & ~n66897;
  assign n66899 = ~controllable_hmaster1 & ~n66898;
  assign n66900 = ~n19816 & ~n66899;
  assign n66901 = i_hlock6 & ~n66900;
  assign n66902 = ~n19843 & ~n66899;
  assign n66903 = ~i_hlock6 & ~n66902;
  assign n66904 = ~n66901 & ~n66903;
  assign n66905 = ~controllable_hgrant6 & ~n66904;
  assign n66906 = ~n13894 & ~n66905;
  assign n66907 = ~controllable_hmaster0 & ~n66906;
  assign n66908 = ~n19804 & ~n66907;
  assign n66909 = ~controllable_hmaster3 & ~n66908;
  assign n66910 = ~n29864 & ~n66909;
  assign n66911 = i_hlock7 & ~n66910;
  assign n66912 = ~n19859 & ~n66907;
  assign n66913 = ~controllable_hmaster3 & ~n66912;
  assign n66914 = ~n29864 & ~n66913;
  assign n66915 = ~i_hlock7 & ~n66914;
  assign n66916 = ~n66911 & ~n66915;
  assign n66917 = i_hbusreq7 & ~n66916;
  assign n66918 = i_hbusreq8 & ~n66908;
  assign n66919 = i_hbusreq6 & ~n66904;
  assign n66920 = i_hbusreq5 & ~n66894;
  assign n66921 = i_hbusreq4 & ~n66892;
  assign n66922 = i_hbusreq9 & ~n66892;
  assign n66923 = i_hbusreq3 & ~n66890;
  assign n66924 = i_hbusreq1 & ~n66888;
  assign n66925 = ~n12896 & ~n16120;
  assign n66926 = i_hlock0 & ~n66925;
  assign n66927 = ~n16627 & ~n66926;
  assign n66928 = ~i_hbusreq0 & ~n66927;
  assign n66929 = ~n16624 & ~n66928;
  assign n66930 = ~i_hbusreq2 & ~n66929;
  assign n66931 = ~n16623 & ~n66930;
  assign n66932 = ~controllable_hgrant2 & n66931;
  assign n66933 = ~n14231 & ~n66932;
  assign n66934 = n7928 & ~n66933;
  assign n66935 = ~n66518 & ~n66934;
  assign n66936 = ~i_hbusreq1 & ~n66935;
  assign n66937 = ~n66924 & ~n66936;
  assign n66938 = ~controllable_hgrant1 & ~n66937;
  assign n66939 = ~n14229 & ~n66938;
  assign n66940 = ~i_hbusreq3 & ~n66939;
  assign n66941 = ~n66923 & ~n66940;
  assign n66942 = ~controllable_hgrant3 & ~n66941;
  assign n66943 = ~n14227 & ~n66942;
  assign n66944 = ~i_hbusreq9 & ~n66943;
  assign n66945 = ~n66922 & ~n66944;
  assign n66946 = ~i_hbusreq4 & ~n66945;
  assign n66947 = ~n66921 & ~n66946;
  assign n66948 = ~controllable_hgrant4 & ~n66947;
  assign n66949 = ~n14224 & ~n66948;
  assign n66950 = ~i_hbusreq5 & ~n66949;
  assign n66951 = ~n66920 & ~n66950;
  assign n66952 = ~controllable_hgrant5 & ~n66951;
  assign n66953 = ~n14222 & ~n66952;
  assign n66954 = ~controllable_hmaster2 & ~n66953;
  assign n66955 = ~n20191 & ~n66954;
  assign n66956 = ~controllable_hmaster1 & ~n66955;
  assign n66957 = ~n20177 & ~n66956;
  assign n66958 = i_hlock6 & ~n66957;
  assign n66959 = ~n20229 & ~n66956;
  assign n66960 = ~i_hlock6 & ~n66959;
  assign n66961 = ~n66958 & ~n66960;
  assign n66962 = ~i_hbusreq6 & ~n66961;
  assign n66963 = ~n66919 & ~n66962;
  assign n66964 = ~controllable_hgrant6 & ~n66963;
  assign n66965 = ~n14173 & ~n66964;
  assign n66966 = ~controllable_hmaster0 & ~n66965;
  assign n66967 = ~n20149 & ~n66966;
  assign n66968 = ~i_hbusreq8 & ~n66967;
  assign n66969 = ~n66918 & ~n66968;
  assign n66970 = ~controllable_hmaster3 & ~n66969;
  assign n66971 = ~n29931 & ~n66970;
  assign n66972 = i_hlock7 & ~n66971;
  assign n66973 = i_hbusreq8 & ~n66912;
  assign n66974 = ~n20253 & ~n66966;
  assign n66975 = ~i_hbusreq8 & ~n66974;
  assign n66976 = ~n66973 & ~n66975;
  assign n66977 = ~controllable_hmaster3 & ~n66976;
  assign n66978 = ~n29931 & ~n66977;
  assign n66979 = ~i_hlock7 & ~n66978;
  assign n66980 = ~n66972 & ~n66979;
  assign n66981 = ~i_hbusreq7 & ~n66980;
  assign n66982 = ~n66917 & ~n66981;
  assign n66983 = n7924 & ~n66982;
  assign n66984 = ~n66887 & ~n66983;
  assign n66985 = ~n8214 & ~n66984;
  assign n66986 = ~n30017 & ~n66811;
  assign n66987 = i_hlock7 & ~n66986;
  assign n66988 = ~n30017 & ~n66815;
  assign n66989 = ~i_hlock7 & ~n66988;
  assign n66990 = ~n66987 & ~n66989;
  assign n66991 = i_hbusreq7 & ~n66990;
  assign n66992 = ~n30058 & ~n66874;
  assign n66993 = i_hlock7 & ~n66992;
  assign n66994 = ~n30058 & ~n66881;
  assign n66995 = ~i_hlock7 & ~n66994;
  assign n66996 = ~n66993 & ~n66995;
  assign n66997 = ~i_hbusreq7 & ~n66996;
  assign n66998 = ~n66991 & ~n66997;
  assign n66999 = ~n7924 & ~n66998;
  assign n67000 = ~n30086 & ~n66909;
  assign n67001 = i_hlock7 & ~n67000;
  assign n67002 = ~n30086 & ~n66913;
  assign n67003 = ~i_hlock7 & ~n67002;
  assign n67004 = ~n67001 & ~n67003;
  assign n67005 = i_hbusreq7 & ~n67004;
  assign n67006 = ~n30127 & ~n66970;
  assign n67007 = i_hlock7 & ~n67006;
  assign n67008 = ~n30127 & ~n66977;
  assign n67009 = ~i_hlock7 & ~n67008;
  assign n67010 = ~n67007 & ~n67009;
  assign n67011 = ~i_hbusreq7 & ~n67010;
  assign n67012 = ~n67005 & ~n67011;
  assign n67013 = n7924 & ~n67012;
  assign n67014 = ~n66999 & ~n67013;
  assign n67015 = n8214 & ~n67014;
  assign n67016 = ~n66985 & ~n67015;
  assign n67017 = ~n8202 & ~n67016;
  assign n67018 = ~n20293 & ~n66809;
  assign n67019 = ~controllable_hmaster3 & ~n67018;
  assign n67020 = ~n30877 & ~n67019;
  assign n67021 = i_hlock7 & ~n67020;
  assign n67022 = ~n20303 & ~n66809;
  assign n67023 = ~controllable_hmaster3 & ~n67022;
  assign n67024 = ~n30877 & ~n67023;
  assign n67025 = ~i_hlock7 & ~n67024;
  assign n67026 = ~n67021 & ~n67025;
  assign n67027 = i_hbusreq7 & ~n67026;
  assign n67028 = i_hbusreq8 & ~n67018;
  assign n67029 = ~n20348 & ~n66870;
  assign n67030 = ~i_hbusreq8 & ~n67029;
  assign n67031 = ~n67028 & ~n67030;
  assign n67032 = ~controllable_hmaster3 & ~n67031;
  assign n67033 = ~n30896 & ~n67032;
  assign n67034 = i_hlock7 & ~n67033;
  assign n67035 = i_hbusreq8 & ~n67022;
  assign n67036 = ~n20364 & ~n66870;
  assign n67037 = ~i_hbusreq8 & ~n67036;
  assign n67038 = ~n67035 & ~n67037;
  assign n67039 = ~controllable_hmaster3 & ~n67038;
  assign n67040 = ~n30896 & ~n67039;
  assign n67041 = ~i_hlock7 & ~n67040;
  assign n67042 = ~n67034 & ~n67041;
  assign n67043 = ~i_hbusreq7 & ~n67042;
  assign n67044 = ~n67027 & ~n67043;
  assign n67045 = ~n7924 & ~n67044;
  assign n67046 = ~n20401 & ~n66907;
  assign n67047 = ~controllable_hmaster3 & ~n67046;
  assign n67048 = ~n30920 & ~n67047;
  assign n67049 = i_hlock7 & ~n67048;
  assign n67050 = ~n20412 & ~n66907;
  assign n67051 = ~controllable_hmaster3 & ~n67050;
  assign n67052 = ~n30920 & ~n67051;
  assign n67053 = ~i_hlock7 & ~n67052;
  assign n67054 = ~n67049 & ~n67053;
  assign n67055 = i_hbusreq7 & ~n67054;
  assign n67056 = i_hbusreq8 & ~n67046;
  assign n67057 = ~n20458 & ~n66966;
  assign n67058 = ~i_hbusreq8 & ~n67057;
  assign n67059 = ~n67056 & ~n67058;
  assign n67060 = ~controllable_hmaster3 & ~n67059;
  assign n67061 = ~n30939 & ~n67060;
  assign n67062 = i_hlock7 & ~n67061;
  assign n67063 = i_hbusreq8 & ~n67050;
  assign n67064 = ~n20475 & ~n66966;
  assign n67065 = ~i_hbusreq8 & ~n67064;
  assign n67066 = ~n67063 & ~n67065;
  assign n67067 = ~controllable_hmaster3 & ~n67066;
  assign n67068 = ~n30939 & ~n67067;
  assign n67069 = ~i_hlock7 & ~n67068;
  assign n67070 = ~n67062 & ~n67069;
  assign n67071 = ~i_hbusreq7 & ~n67070;
  assign n67072 = ~n67055 & ~n67071;
  assign n67073 = n7924 & ~n67072;
  assign n67074 = ~n67045 & ~n67073;
  assign n67075 = ~n8214 & ~n67074;
  assign n67076 = ~n20489 & ~n66801;
  assign n67077 = i_hlock6 & ~n67076;
  assign n67078 = ~n20493 & ~n66801;
  assign n67079 = ~i_hlock6 & ~n67078;
  assign n67080 = ~n67077 & ~n67079;
  assign n67081 = ~controllable_hgrant6 & ~n67080;
  assign n67082 = ~n13894 & ~n67081;
  assign n67083 = ~controllable_hmaster0 & ~n67082;
  assign n67084 = ~n19279 & ~n67083;
  assign n67085 = ~controllable_hmaster3 & ~n67084;
  assign n67086 = ~n30877 & ~n67085;
  assign n67087 = i_hlock7 & ~n67086;
  assign n67088 = ~n19334 & ~n67083;
  assign n67089 = ~controllable_hmaster3 & ~n67088;
  assign n67090 = ~n30877 & ~n67089;
  assign n67091 = ~i_hlock7 & ~n67090;
  assign n67092 = ~n67087 & ~n67091;
  assign n67093 = i_hbusreq7 & ~n67092;
  assign n67094 = i_hbusreq8 & ~n67084;
  assign n67095 = i_hbusreq6 & ~n67080;
  assign n67096 = ~n20513 & ~n66860;
  assign n67097 = i_hlock6 & ~n67096;
  assign n67098 = ~n20517 & ~n66860;
  assign n67099 = ~i_hlock6 & ~n67098;
  assign n67100 = ~n67097 & ~n67099;
  assign n67101 = ~i_hbusreq6 & ~n67100;
  assign n67102 = ~n67095 & ~n67101;
  assign n67103 = ~controllable_hgrant6 & ~n67102;
  assign n67104 = ~n14802 & ~n67103;
  assign n67105 = ~controllable_hmaster0 & ~n67104;
  assign n67106 = ~n19556 & ~n67105;
  assign n67107 = ~i_hbusreq8 & ~n67106;
  assign n67108 = ~n67094 & ~n67107;
  assign n67109 = ~controllable_hmaster3 & ~n67108;
  assign n67110 = ~n30896 & ~n67109;
  assign n67111 = i_hlock7 & ~n67110;
  assign n67112 = i_hbusreq8 & ~n67088;
  assign n67113 = ~n19660 & ~n67105;
  assign n67114 = ~i_hbusreq8 & ~n67113;
  assign n67115 = ~n67112 & ~n67114;
  assign n67116 = ~controllable_hmaster3 & ~n67115;
  assign n67117 = ~n30896 & ~n67116;
  assign n67118 = ~i_hlock7 & ~n67117;
  assign n67119 = ~n67111 & ~n67118;
  assign n67120 = ~i_hbusreq7 & ~n67119;
  assign n67121 = ~n67093 & ~n67120;
  assign n67122 = ~n7924 & ~n67121;
  assign n67123 = ~n20544 & ~n66899;
  assign n67124 = i_hlock6 & ~n67123;
  assign n67125 = ~n20548 & ~n66899;
  assign n67126 = ~i_hlock6 & ~n67125;
  assign n67127 = ~n67124 & ~n67126;
  assign n67128 = ~controllable_hgrant6 & ~n67127;
  assign n67129 = ~n13894 & ~n67128;
  assign n67130 = ~controllable_hmaster0 & ~n67129;
  assign n67131 = ~n19804 & ~n67130;
  assign n67132 = ~controllable_hmaster3 & ~n67131;
  assign n67133 = ~n30920 & ~n67132;
  assign n67134 = i_hlock7 & ~n67133;
  assign n67135 = ~n19859 & ~n67130;
  assign n67136 = ~controllable_hmaster3 & ~n67135;
  assign n67137 = ~n30920 & ~n67136;
  assign n67138 = ~i_hlock7 & ~n67137;
  assign n67139 = ~n67134 & ~n67138;
  assign n67140 = i_hbusreq7 & ~n67139;
  assign n67141 = i_hbusreq8 & ~n67131;
  assign n67142 = i_hbusreq6 & ~n67127;
  assign n67143 = ~n20568 & ~n66956;
  assign n67144 = i_hlock6 & ~n67143;
  assign n67145 = ~n20572 & ~n66956;
  assign n67146 = ~i_hlock6 & ~n67145;
  assign n67147 = ~n67144 & ~n67146;
  assign n67148 = ~i_hbusreq6 & ~n67147;
  assign n67149 = ~n67142 & ~n67148;
  assign n67150 = ~controllable_hgrant6 & ~n67149;
  assign n67151 = ~n14802 & ~n67150;
  assign n67152 = ~controllable_hmaster0 & ~n67151;
  assign n67153 = ~n20149 & ~n67152;
  assign n67154 = ~i_hbusreq8 & ~n67153;
  assign n67155 = ~n67141 & ~n67154;
  assign n67156 = ~controllable_hmaster3 & ~n67155;
  assign n67157 = ~n30939 & ~n67156;
  assign n67158 = i_hlock7 & ~n67157;
  assign n67159 = i_hbusreq8 & ~n67135;
  assign n67160 = ~n20253 & ~n67152;
  assign n67161 = ~i_hbusreq8 & ~n67160;
  assign n67162 = ~n67159 & ~n67161;
  assign n67163 = ~controllable_hmaster3 & ~n67162;
  assign n67164 = ~n30939 & ~n67163;
  assign n67165 = ~i_hlock7 & ~n67164;
  assign n67166 = ~n67158 & ~n67165;
  assign n67167 = ~i_hbusreq7 & ~n67166;
  assign n67168 = ~n67140 & ~n67167;
  assign n67169 = n7924 & ~n67168;
  assign n67170 = ~n67122 & ~n67169;
  assign n67171 = n8214 & ~n67170;
  assign n67172 = ~n67075 & ~n67171;
  assign n67173 = n8202 & ~n67172;
  assign n67174 = ~n67017 & ~n67173;
  assign n67175 = n7920 & ~n67174;
  assign n67176 = ~n8877 & ~n67175;
  assign n67177 = ~n7728 & ~n67176;
  assign n67178 = ~n66789 & ~n67177;
  assign n67179 = n7723 & ~n67178;
  assign n67180 = ~n7723 & ~n67176;
  assign n67181 = ~n67179 & ~n67180;
  assign n67182 = n7714 & ~n67181;
  assign n67183 = n7723 & ~n67176;
  assign n67184 = i_hlock0 & ~n20612;
  assign n67185 = ~n20876 & ~n67184;
  assign n67186 = ~controllable_hgrant2 & n67185;
  assign n67187 = ~n7814 & ~n67186;
  assign n67188 = n7733 & ~n67187;
  assign n67189 = ~n17507 & ~n67188;
  assign n67190 = n7928 & ~n67189;
  assign n67191 = ~n19671 & ~n67190;
  assign n67192 = ~controllable_hgrant1 & ~n67191;
  assign n67193 = ~n13155 & ~n67192;
  assign n67194 = ~controllable_hgrant3 & ~n67193;
  assign n67195 = ~n13154 & ~n67194;
  assign n67196 = ~controllable_hgrant4 & ~n67195;
  assign n67197 = ~n13153 & ~n67196;
  assign n67198 = ~controllable_hgrant5 & ~n67197;
  assign n67199 = ~n13152 & ~n67198;
  assign n67200 = controllable_hmaster1 & ~n67199;
  assign n67201 = controllable_hmaster2 & ~n67199;
  assign n67202 = i_hlock0 & ~n17464;
  assign n67203 = ~n18726 & ~n67202;
  assign n67204 = ~controllable_hgrant2 & n67203;
  assign n67205 = ~n7814 & ~n67204;
  assign n67206 = n7733 & ~n67205;
  assign n67207 = ~n17507 & ~n67206;
  assign n67208 = n7928 & ~n67207;
  assign n67209 = ~n8221 & ~n67208;
  assign n67210 = ~controllable_hgrant1 & ~n67209;
  assign n67211 = ~n12611 & ~n67210;
  assign n67212 = ~controllable_hgrant3 & ~n67211;
  assign n67213 = ~n12610 & ~n67212;
  assign n67214 = i_hlock9 & ~n67213;
  assign n67215 = ~n8235 & ~n67208;
  assign n67216 = ~controllable_hgrant1 & ~n67215;
  assign n67217 = ~n12638 & ~n67216;
  assign n67218 = ~controllable_hgrant3 & ~n67217;
  assign n67219 = ~n12637 & ~n67218;
  assign n67220 = ~i_hlock9 & ~n67219;
  assign n67221 = ~n67214 & ~n67220;
  assign n67222 = ~controllable_hgrant4 & ~n67221;
  assign n67223 = ~n12609 & ~n67222;
  assign n67224 = ~controllable_hgrant5 & ~n67223;
  assign n67225 = ~n12608 & ~n67224;
  assign n67226 = ~controllable_hmaster2 & ~n67225;
  assign n67227 = ~n67201 & ~n67226;
  assign n67228 = ~controllable_hmaster1 & ~n67227;
  assign n67229 = ~n67200 & ~n67228;
  assign n67230 = ~controllable_hgrant6 & ~n67229;
  assign n67231 = ~n13122 & ~n67230;
  assign n67232 = controllable_hmaster0 & ~n67231;
  assign n67233 = ~n8221 & ~n67190;
  assign n67234 = ~controllable_hgrant1 & ~n67233;
  assign n67235 = ~n12611 & ~n67234;
  assign n67236 = ~controllable_hgrant3 & ~n67235;
  assign n67237 = ~n12610 & ~n67236;
  assign n67238 = ~controllable_hgrant4 & ~n67237;
  assign n67239 = ~n13408 & ~n67238;
  assign n67240 = ~controllable_hgrant5 & ~n67239;
  assign n67241 = ~n13407 & ~n67240;
  assign n67242 = ~controllable_hmaster2 & ~n67241;
  assign n67243 = ~n67201 & ~n67242;
  assign n67244 = ~controllable_hmaster1 & ~n67243;
  assign n67245 = ~n67200 & ~n67244;
  assign n67246 = ~controllable_hgrant6 & ~n67245;
  assign n67247 = ~n13406 & ~n67246;
  assign n67248 = ~controllable_hmaster0 & ~n67247;
  assign n67249 = ~n67232 & ~n67248;
  assign n67250 = i_hlock8 & ~n67249;
  assign n67251 = ~n8235 & ~n67190;
  assign n67252 = ~controllable_hgrant1 & ~n67251;
  assign n67253 = ~n12638 & ~n67252;
  assign n67254 = ~controllable_hgrant3 & ~n67253;
  assign n67255 = ~n12637 & ~n67254;
  assign n67256 = ~controllable_hgrant4 & ~n67255;
  assign n67257 = ~n13429 & ~n67256;
  assign n67258 = ~controllable_hgrant5 & ~n67257;
  assign n67259 = ~n13428 & ~n67258;
  assign n67260 = ~controllable_hmaster2 & ~n67259;
  assign n67261 = ~n67201 & ~n67260;
  assign n67262 = ~controllable_hmaster1 & ~n67261;
  assign n67263 = ~n67200 & ~n67262;
  assign n67264 = ~controllable_hgrant6 & ~n67263;
  assign n67265 = ~n13427 & ~n67264;
  assign n67266 = ~controllable_hmaster0 & ~n67265;
  assign n67267 = ~n67232 & ~n67266;
  assign n67268 = ~i_hlock8 & ~n67267;
  assign n67269 = ~n67250 & ~n67268;
  assign n67270 = controllable_hmaster3 & ~n67269;
  assign n67271 = controllable_hmaster2 & ~n67241;
  assign n67272 = i_hlock3 & ~n67235;
  assign n67273 = ~i_hlock3 & ~n67253;
  assign n67274 = ~n67272 & ~n67273;
  assign n67275 = ~controllable_hgrant3 & ~n67274;
  assign n67276 = ~n13852 & ~n67275;
  assign n67277 = ~controllable_hgrant4 & ~n67276;
  assign n67278 = ~n13851 & ~n67277;
  assign n67279 = ~controllable_hgrant5 & ~n67278;
  assign n67280 = ~n13850 & ~n67279;
  assign n67281 = ~controllable_hmaster2 & ~n67280;
  assign n67282 = ~n67271 & ~n67281;
  assign n67283 = controllable_hmaster1 & ~n67282;
  assign n67284 = i_hlock5 & ~n67239;
  assign n67285 = ~i_hlock5 & ~n67257;
  assign n67286 = ~n67284 & ~n67285;
  assign n67287 = ~controllable_hgrant5 & ~n67286;
  assign n67288 = ~n13865 & ~n67287;
  assign n67289 = controllable_hmaster2 & ~n67288;
  assign n67290 = i_hlock1 & ~n67233;
  assign n67291 = ~i_hlock1 & ~n67251;
  assign n67292 = ~n67290 & ~n67291;
  assign n67293 = ~controllable_hgrant1 & ~n67292;
  assign n67294 = ~n13875 & ~n67293;
  assign n67295 = ~controllable_hgrant3 & ~n67294;
  assign n67296 = ~n13874 & ~n67295;
  assign n67297 = ~controllable_hgrant4 & ~n67296;
  assign n67298 = ~n13873 & ~n67297;
  assign n67299 = ~controllable_hgrant5 & ~n67298;
  assign n67300 = ~n13872 & ~n67299;
  assign n67301 = ~controllable_hmaster2 & ~n67300;
  assign n67302 = ~n67289 & ~n67301;
  assign n67303 = ~controllable_hmaster1 & ~n67302;
  assign n67304 = ~n67283 & ~n67303;
  assign n67305 = ~controllable_hgrant6 & ~n67304;
  assign n67306 = ~n13849 & ~n67305;
  assign n67307 = controllable_hmaster0 & ~n67306;
  assign n67308 = ~n9213 & ~n67190;
  assign n67309 = ~controllable_hgrant1 & ~n67308;
  assign n67310 = ~n13898 & ~n67309;
  assign n67311 = ~controllable_hgrant3 & ~n67310;
  assign n67312 = ~n13897 & ~n67311;
  assign n67313 = ~controllable_hgrant4 & ~n67312;
  assign n67314 = ~n13896 & ~n67313;
  assign n67315 = ~controllable_hgrant5 & ~n67314;
  assign n67316 = ~n13895 & ~n67315;
  assign n67317 = ~controllable_hmaster2 & ~n67316;
  assign n67318 = ~n67271 & ~n67317;
  assign n67319 = controllable_hmaster1 & ~n67318;
  assign n67320 = i_hlock4 & ~n67237;
  assign n67321 = ~i_hlock4 & ~n67255;
  assign n67322 = ~n67320 & ~n67321;
  assign n67323 = ~controllable_hgrant4 & ~n67322;
  assign n67324 = ~n13912 & ~n67323;
  assign n67325 = ~controllable_hgrant5 & ~n67324;
  assign n67326 = ~n13911 & ~n67325;
  assign n67327 = controllable_hmaster2 & ~n67326;
  assign n67328 = i_hlock0 & ~n20644;
  assign n67329 = ~n20944 & ~n67328;
  assign n67330 = ~controllable_hgrant2 & n67329;
  assign n67331 = ~n7814 & ~n67330;
  assign n67332 = n7733 & ~n67331;
  assign n67333 = ~n16507 & ~n67332;
  assign n67334 = n7928 & ~n67333;
  assign n67335 = ~n66518 & ~n67334;
  assign n67336 = ~controllable_hgrant1 & ~n67335;
  assign n67337 = ~n13924 & ~n67336;
  assign n67338 = ~controllable_hgrant3 & ~n67337;
  assign n67339 = ~n13923 & ~n67338;
  assign n67340 = ~controllable_hgrant4 & ~n67339;
  assign n67341 = ~n13922 & ~n67340;
  assign n67342 = ~controllable_hgrant5 & ~n67341;
  assign n67343 = ~n13921 & ~n67342;
  assign n67344 = ~controllable_hmaster2 & ~n67343;
  assign n67345 = ~n67327 & ~n67344;
  assign n67346 = ~controllable_hmaster1 & ~n67345;
  assign n67347 = ~n67319 & ~n67346;
  assign n67348 = i_hlock6 & ~n67347;
  assign n67349 = controllable_hmaster2 & ~n67259;
  assign n67350 = ~n67317 & ~n67349;
  assign n67351 = controllable_hmaster1 & ~n67350;
  assign n67352 = ~n67346 & ~n67351;
  assign n67353 = ~i_hlock6 & ~n67352;
  assign n67354 = ~n67348 & ~n67353;
  assign n67355 = ~controllable_hgrant6 & ~n67354;
  assign n67356 = ~n13894 & ~n67355;
  assign n67357 = ~controllable_hmaster0 & ~n67356;
  assign n67358 = ~n67307 & ~n67357;
  assign n67359 = ~controllable_hmaster3 & ~n67358;
  assign n67360 = ~n67270 & ~n67359;
  assign n67361 = i_hlock7 & ~n67360;
  assign n67362 = ~n67281 & ~n67349;
  assign n67363 = controllable_hmaster1 & ~n67362;
  assign n67364 = ~n67303 & ~n67363;
  assign n67365 = ~controllable_hgrant6 & ~n67364;
  assign n67366 = ~n13951 & ~n67365;
  assign n67367 = controllable_hmaster0 & ~n67366;
  assign n67368 = ~n67357 & ~n67367;
  assign n67369 = ~controllable_hmaster3 & ~n67368;
  assign n67370 = ~n67270 & ~n67369;
  assign n67371 = ~i_hlock7 & ~n67370;
  assign n67372 = ~n67361 & ~n67371;
  assign n67373 = i_hbusreq7 & ~n67372;
  assign n67374 = i_hbusreq8 & ~n67269;
  assign n67375 = i_hbusreq6 & ~n67229;
  assign n67376 = i_hbusreq5 & ~n67197;
  assign n67377 = i_hbusreq4 & ~n67195;
  assign n67378 = i_hbusreq9 & ~n67195;
  assign n67379 = i_hbusreq3 & ~n67193;
  assign n67380 = i_hbusreq1 & ~n67191;
  assign n67381 = i_hbusreq2 & ~n67185;
  assign n67382 = i_hbusreq0 & ~n67185;
  assign n67383 = ~n12799 & ~n17089;
  assign n67384 = i_hlock0 & ~n67383;
  assign n67385 = ~n20876 & ~n67384;
  assign n67386 = ~i_hbusreq0 & ~n67385;
  assign n67387 = ~n67382 & ~n67386;
  assign n67388 = ~i_hbusreq2 & ~n67387;
  assign n67389 = ~n67381 & ~n67388;
  assign n67390 = ~controllable_hgrant2 & n67389;
  assign n67391 = ~n12694 & ~n67390;
  assign n67392 = n7733 & ~n67391;
  assign n67393 = ~n18800 & ~n67392;
  assign n67394 = n7928 & ~n67393;
  assign n67395 = ~n19873 & ~n67394;
  assign n67396 = ~i_hbusreq1 & ~n67395;
  assign n67397 = ~n67380 & ~n67396;
  assign n67398 = ~controllable_hgrant1 & ~n67397;
  assign n67399 = ~n13968 & ~n67398;
  assign n67400 = ~i_hbusreq3 & ~n67399;
  assign n67401 = ~n67379 & ~n67400;
  assign n67402 = ~controllable_hgrant3 & ~n67401;
  assign n67403 = ~n13967 & ~n67402;
  assign n67404 = ~i_hbusreq9 & ~n67403;
  assign n67405 = ~n67378 & ~n67404;
  assign n67406 = ~i_hbusreq4 & ~n67405;
  assign n67407 = ~n67377 & ~n67406;
  assign n67408 = ~controllable_hgrant4 & ~n67407;
  assign n67409 = ~n13966 & ~n67408;
  assign n67410 = ~i_hbusreq5 & ~n67409;
  assign n67411 = ~n67376 & ~n67410;
  assign n67412 = ~controllable_hgrant5 & ~n67411;
  assign n67413 = ~n13965 & ~n67412;
  assign n67414 = controllable_hmaster1 & ~n67413;
  assign n67415 = controllable_hmaster2 & ~n67413;
  assign n67416 = i_hbusreq5 & ~n67223;
  assign n67417 = i_hbusreq4 & ~n67221;
  assign n67418 = i_hbusreq9 & ~n67221;
  assign n67419 = i_hbusreq3 & ~n67211;
  assign n67420 = i_hbusreq1 & ~n67209;
  assign n67421 = i_hbusreq2 & ~n67203;
  assign n67422 = i_hbusreq0 & ~n67203;
  assign n67423 = controllable_hmastlock & ~n7933;
  assign n67424 = controllable_locked & ~n67423;
  assign n67425 = ~n14243 & ~n67424;
  assign n67426 = i_hlock0 & ~n67425;
  assign n67427 = ~n18726 & ~n67426;
  assign n67428 = ~i_hbusreq0 & ~n67427;
  assign n67429 = ~n67422 & ~n67428;
  assign n67430 = ~i_hbusreq2 & ~n67429;
  assign n67431 = ~n67421 & ~n67430;
  assign n67432 = ~controllable_hgrant2 & n67431;
  assign n67433 = ~n12706 & ~n67432;
  assign n67434 = n7733 & ~n67433;
  assign n67435 = ~n18800 & ~n67434;
  assign n67436 = n7928 & ~n67435;
  assign n67437 = ~n8265 & ~n67436;
  assign n67438 = ~i_hbusreq1 & ~n67437;
  assign n67439 = ~n67420 & ~n67438;
  assign n67440 = ~controllable_hgrant1 & ~n67439;
  assign n67441 = ~n12681 & ~n67440;
  assign n67442 = ~i_hbusreq3 & ~n67441;
  assign n67443 = ~n67419 & ~n67442;
  assign n67444 = ~controllable_hgrant3 & ~n67443;
  assign n67445 = ~n12679 & ~n67444;
  assign n67446 = i_hlock9 & ~n67445;
  assign n67447 = i_hbusreq3 & ~n67217;
  assign n67448 = i_hbusreq1 & ~n67215;
  assign n67449 = ~n8297 & ~n67436;
  assign n67450 = ~i_hbusreq1 & ~n67449;
  assign n67451 = ~n67448 & ~n67450;
  assign n67452 = ~controllable_hgrant1 & ~n67451;
  assign n67453 = ~n12730 & ~n67452;
  assign n67454 = ~i_hbusreq3 & ~n67453;
  assign n67455 = ~n67447 & ~n67454;
  assign n67456 = ~controllable_hgrant3 & ~n67455;
  assign n67457 = ~n12728 & ~n67456;
  assign n67458 = ~i_hlock9 & ~n67457;
  assign n67459 = ~n67446 & ~n67458;
  assign n67460 = ~i_hbusreq9 & ~n67459;
  assign n67461 = ~n67418 & ~n67460;
  assign n67462 = ~i_hbusreq4 & ~n67461;
  assign n67463 = ~n67417 & ~n67462;
  assign n67464 = ~controllable_hgrant4 & ~n67463;
  assign n67465 = ~n12676 & ~n67464;
  assign n67466 = ~i_hbusreq5 & ~n67465;
  assign n67467 = ~n67416 & ~n67466;
  assign n67468 = ~controllable_hgrant5 & ~n67467;
  assign n67469 = ~n12674 & ~n67468;
  assign n67470 = ~controllable_hmaster2 & ~n67469;
  assign n67471 = ~n67415 & ~n67470;
  assign n67472 = ~controllable_hmaster1 & ~n67471;
  assign n67473 = ~n67414 & ~n67472;
  assign n67474 = ~i_hbusreq6 & ~n67473;
  assign n67475 = ~n67375 & ~n67474;
  assign n67476 = ~controllable_hgrant6 & ~n67475;
  assign n67477 = ~n13818 & ~n67476;
  assign n67478 = controllable_hmaster0 & ~n67477;
  assign n67479 = i_hbusreq6 & ~n67245;
  assign n67480 = i_hbusreq5 & ~n67239;
  assign n67481 = i_hbusreq4 & ~n67237;
  assign n67482 = i_hbusreq9 & ~n67237;
  assign n67483 = i_hbusreq3 & ~n67235;
  assign n67484 = i_hbusreq1 & ~n67233;
  assign n67485 = ~n8265 & ~n67394;
  assign n67486 = ~i_hbusreq1 & ~n67485;
  assign n67487 = ~n67484 & ~n67486;
  assign n67488 = ~controllable_hgrant1 & ~n67487;
  assign n67489 = ~n14023 & ~n67488;
  assign n67490 = ~i_hbusreq3 & ~n67489;
  assign n67491 = ~n67483 & ~n67490;
  assign n67492 = ~controllable_hgrant3 & ~n67491;
  assign n67493 = ~n14022 & ~n67492;
  assign n67494 = ~i_hbusreq9 & ~n67493;
  assign n67495 = ~n67482 & ~n67494;
  assign n67496 = ~i_hbusreq4 & ~n67495;
  assign n67497 = ~n67481 & ~n67496;
  assign n67498 = ~controllable_hgrant4 & ~n67497;
  assign n67499 = ~n14021 & ~n67498;
  assign n67500 = ~i_hbusreq5 & ~n67499;
  assign n67501 = ~n67480 & ~n67500;
  assign n67502 = ~controllable_hgrant5 & ~n67501;
  assign n67503 = ~n14020 & ~n67502;
  assign n67504 = ~controllable_hmaster2 & ~n67503;
  assign n67505 = ~n67415 & ~n67504;
  assign n67506 = ~controllable_hmaster1 & ~n67505;
  assign n67507 = ~n67414 & ~n67506;
  assign n67508 = ~i_hbusreq6 & ~n67507;
  assign n67509 = ~n67479 & ~n67508;
  assign n67510 = ~controllable_hgrant6 & ~n67509;
  assign n67511 = ~n14019 & ~n67510;
  assign n67512 = ~controllable_hmaster0 & ~n67511;
  assign n67513 = ~n67478 & ~n67512;
  assign n67514 = i_hlock8 & ~n67513;
  assign n67515 = i_hbusreq6 & ~n67263;
  assign n67516 = i_hbusreq5 & ~n67257;
  assign n67517 = i_hbusreq4 & ~n67255;
  assign n67518 = i_hbusreq9 & ~n67255;
  assign n67519 = i_hbusreq3 & ~n67253;
  assign n67520 = i_hbusreq1 & ~n67251;
  assign n67521 = ~n8297 & ~n67394;
  assign n67522 = ~i_hbusreq1 & ~n67521;
  assign n67523 = ~n67520 & ~n67522;
  assign n67524 = ~controllable_hgrant1 & ~n67523;
  assign n67525 = ~n14058 & ~n67524;
  assign n67526 = ~i_hbusreq3 & ~n67525;
  assign n67527 = ~n67519 & ~n67526;
  assign n67528 = ~controllable_hgrant3 & ~n67527;
  assign n67529 = ~n14057 & ~n67528;
  assign n67530 = ~i_hbusreq9 & ~n67529;
  assign n67531 = ~n67518 & ~n67530;
  assign n67532 = ~i_hbusreq4 & ~n67531;
  assign n67533 = ~n67517 & ~n67532;
  assign n67534 = ~controllable_hgrant4 & ~n67533;
  assign n67535 = ~n14056 & ~n67534;
  assign n67536 = ~i_hbusreq5 & ~n67535;
  assign n67537 = ~n67516 & ~n67536;
  assign n67538 = ~controllable_hgrant5 & ~n67537;
  assign n67539 = ~n14055 & ~n67538;
  assign n67540 = ~controllable_hmaster2 & ~n67539;
  assign n67541 = ~n67415 & ~n67540;
  assign n67542 = ~controllable_hmaster1 & ~n67541;
  assign n67543 = ~n67414 & ~n67542;
  assign n67544 = ~i_hbusreq6 & ~n67543;
  assign n67545 = ~n67515 & ~n67544;
  assign n67546 = ~controllable_hgrant6 & ~n67545;
  assign n67547 = ~n14054 & ~n67546;
  assign n67548 = ~controllable_hmaster0 & ~n67547;
  assign n67549 = ~n67478 & ~n67548;
  assign n67550 = ~i_hlock8 & ~n67549;
  assign n67551 = ~n67514 & ~n67550;
  assign n67552 = ~i_hbusreq8 & ~n67551;
  assign n67553 = ~n67374 & ~n67552;
  assign n67554 = controllable_hmaster3 & ~n67553;
  assign n67555 = i_hbusreq8 & ~n67358;
  assign n67556 = i_hbusreq6 & ~n67304;
  assign n67557 = controllable_hmaster2 & ~n67503;
  assign n67558 = i_hbusreq5 & ~n67278;
  assign n67559 = i_hbusreq4 & ~n67276;
  assign n67560 = i_hbusreq9 & ~n67276;
  assign n67561 = i_hbusreq3 & ~n67274;
  assign n67562 = i_hlock3 & ~n67489;
  assign n67563 = ~i_hlock3 & ~n67525;
  assign n67564 = ~n67562 & ~n67563;
  assign n67565 = ~i_hbusreq3 & ~n67564;
  assign n67566 = ~n67561 & ~n67565;
  assign n67567 = ~controllable_hgrant3 & ~n67566;
  assign n67568 = ~n14102 & ~n67567;
  assign n67569 = ~i_hbusreq9 & ~n67568;
  assign n67570 = ~n67560 & ~n67569;
  assign n67571 = ~i_hbusreq4 & ~n67570;
  assign n67572 = ~n67559 & ~n67571;
  assign n67573 = ~controllable_hgrant4 & ~n67572;
  assign n67574 = ~n14099 & ~n67573;
  assign n67575 = ~i_hbusreq5 & ~n67574;
  assign n67576 = ~n67558 & ~n67575;
  assign n67577 = ~controllable_hgrant5 & ~n67576;
  assign n67578 = ~n14097 & ~n67577;
  assign n67579 = ~controllable_hmaster2 & ~n67578;
  assign n67580 = ~n67557 & ~n67579;
  assign n67581 = controllable_hmaster1 & ~n67580;
  assign n67582 = i_hbusreq5 & ~n67286;
  assign n67583 = i_hlock5 & ~n67499;
  assign n67584 = ~i_hlock5 & ~n67535;
  assign n67585 = ~n67583 & ~n67584;
  assign n67586 = ~i_hbusreq5 & ~n67585;
  assign n67587 = ~n67582 & ~n67586;
  assign n67588 = ~controllable_hgrant5 & ~n67587;
  assign n67589 = ~n14124 & ~n67588;
  assign n67590 = controllable_hmaster2 & ~n67589;
  assign n67591 = i_hbusreq5 & ~n67298;
  assign n67592 = i_hbusreq4 & ~n67296;
  assign n67593 = i_hbusreq9 & ~n67296;
  assign n67594 = i_hbusreq3 & ~n67294;
  assign n67595 = i_hbusreq1 & ~n67292;
  assign n67596 = i_hlock1 & ~n67485;
  assign n67597 = ~i_hlock1 & ~n67521;
  assign n67598 = ~n67596 & ~n67597;
  assign n67599 = ~i_hbusreq1 & ~n67598;
  assign n67600 = ~n67595 & ~n67599;
  assign n67601 = ~controllable_hgrant1 & ~n67600;
  assign n67602 = ~n14141 & ~n67601;
  assign n67603 = ~i_hbusreq3 & ~n67602;
  assign n67604 = ~n67594 & ~n67603;
  assign n67605 = ~controllable_hgrant3 & ~n67604;
  assign n67606 = ~n14139 & ~n67605;
  assign n67607 = ~i_hbusreq9 & ~n67606;
  assign n67608 = ~n67593 & ~n67607;
  assign n67609 = ~i_hbusreq4 & ~n67608;
  assign n67610 = ~n67592 & ~n67609;
  assign n67611 = ~controllable_hgrant4 & ~n67610;
  assign n67612 = ~n14136 & ~n67611;
  assign n67613 = ~i_hbusreq5 & ~n67612;
  assign n67614 = ~n67591 & ~n67613;
  assign n67615 = ~controllable_hgrant5 & ~n67614;
  assign n67616 = ~n14134 & ~n67615;
  assign n67617 = ~controllable_hmaster2 & ~n67616;
  assign n67618 = ~n67590 & ~n67617;
  assign n67619 = ~controllable_hmaster1 & ~n67618;
  assign n67620 = ~n67581 & ~n67619;
  assign n67621 = ~i_hbusreq6 & ~n67620;
  assign n67622 = ~n67556 & ~n67621;
  assign n67623 = ~controllable_hgrant6 & ~n67622;
  assign n67624 = ~n14094 & ~n67623;
  assign n67625 = controllable_hmaster0 & ~n67624;
  assign n67626 = i_hbusreq6 & ~n67354;
  assign n67627 = i_hbusreq5 & ~n67314;
  assign n67628 = i_hbusreq4 & ~n67312;
  assign n67629 = i_hbusreq9 & ~n67312;
  assign n67630 = i_hbusreq3 & ~n67310;
  assign n67631 = i_hbusreq1 & ~n67308;
  assign n67632 = ~n9379 & ~n67394;
  assign n67633 = ~i_hbusreq1 & ~n67632;
  assign n67634 = ~n67631 & ~n67633;
  assign n67635 = ~controllable_hgrant1 & ~n67634;
  assign n67636 = ~n14182 & ~n67635;
  assign n67637 = ~i_hbusreq3 & ~n67636;
  assign n67638 = ~n67630 & ~n67637;
  assign n67639 = ~controllable_hgrant3 & ~n67638;
  assign n67640 = ~n14180 & ~n67639;
  assign n67641 = ~i_hbusreq9 & ~n67640;
  assign n67642 = ~n67629 & ~n67641;
  assign n67643 = ~i_hbusreq4 & ~n67642;
  assign n67644 = ~n67628 & ~n67643;
  assign n67645 = ~controllable_hgrant4 & ~n67644;
  assign n67646 = ~n14177 & ~n67645;
  assign n67647 = ~i_hbusreq5 & ~n67646;
  assign n67648 = ~n67627 & ~n67647;
  assign n67649 = ~controllable_hgrant5 & ~n67648;
  assign n67650 = ~n14175 & ~n67649;
  assign n67651 = ~controllable_hmaster2 & ~n67650;
  assign n67652 = ~n67557 & ~n67651;
  assign n67653 = controllable_hmaster1 & ~n67652;
  assign n67654 = i_hbusreq5 & ~n67324;
  assign n67655 = i_hbusreq4 & ~n67322;
  assign n67656 = i_hlock4 & ~n67495;
  assign n67657 = ~i_hlock4 & ~n67531;
  assign n67658 = ~n67656 & ~n67657;
  assign n67659 = ~i_hbusreq4 & ~n67658;
  assign n67660 = ~n67655 & ~n67659;
  assign n67661 = ~controllable_hgrant4 & ~n67660;
  assign n67662 = ~n14208 & ~n67661;
  assign n67663 = ~i_hbusreq5 & ~n67662;
  assign n67664 = ~n67654 & ~n67663;
  assign n67665 = ~controllable_hgrant5 & ~n67664;
  assign n67666 = ~n14206 & ~n67665;
  assign n67667 = controllable_hmaster2 & ~n67666;
  assign n67668 = i_hbusreq5 & ~n67341;
  assign n67669 = i_hbusreq4 & ~n67339;
  assign n67670 = i_hbusreq9 & ~n67339;
  assign n67671 = i_hbusreq3 & ~n67337;
  assign n67672 = i_hbusreq1 & ~n67335;
  assign n67673 = ~n7733 & ~n66933;
  assign n67674 = i_hbusreq2 & ~n67329;
  assign n67675 = i_hbusreq0 & ~n67329;
  assign n67676 = ~n12896 & ~n16802;
  assign n67677 = i_hlock0 & ~n67676;
  assign n67678 = ~n20944 & ~n67677;
  assign n67679 = ~i_hbusreq0 & ~n67678;
  assign n67680 = ~n67675 & ~n67679;
  assign n67681 = ~i_hbusreq2 & ~n67680;
  assign n67682 = ~n67674 & ~n67681;
  assign n67683 = ~controllable_hgrant2 & n67682;
  assign n67684 = ~n14231 & ~n67683;
  assign n67685 = n7733 & ~n67684;
  assign n67686 = ~n67673 & ~n67685;
  assign n67687 = n7928 & ~n67686;
  assign n67688 = ~n66518 & ~n67687;
  assign n67689 = ~i_hbusreq1 & ~n67688;
  assign n67690 = ~n67672 & ~n67689;
  assign n67691 = ~controllable_hgrant1 & ~n67690;
  assign n67692 = ~n14229 & ~n67691;
  assign n67693 = ~i_hbusreq3 & ~n67692;
  assign n67694 = ~n67671 & ~n67693;
  assign n67695 = ~controllable_hgrant3 & ~n67694;
  assign n67696 = ~n14227 & ~n67695;
  assign n67697 = ~i_hbusreq9 & ~n67696;
  assign n67698 = ~n67670 & ~n67697;
  assign n67699 = ~i_hbusreq4 & ~n67698;
  assign n67700 = ~n67669 & ~n67699;
  assign n67701 = ~controllable_hgrant4 & ~n67700;
  assign n67702 = ~n14224 & ~n67701;
  assign n67703 = ~i_hbusreq5 & ~n67702;
  assign n67704 = ~n67668 & ~n67703;
  assign n67705 = ~controllable_hgrant5 & ~n67704;
  assign n67706 = ~n14222 & ~n67705;
  assign n67707 = ~controllable_hmaster2 & ~n67706;
  assign n67708 = ~n67667 & ~n67707;
  assign n67709 = ~controllable_hmaster1 & ~n67708;
  assign n67710 = ~n67653 & ~n67709;
  assign n67711 = i_hlock6 & ~n67710;
  assign n67712 = controllable_hmaster2 & ~n67539;
  assign n67713 = ~n67651 & ~n67712;
  assign n67714 = controllable_hmaster1 & ~n67713;
  assign n67715 = ~n67709 & ~n67714;
  assign n67716 = ~i_hlock6 & ~n67715;
  assign n67717 = ~n67711 & ~n67716;
  assign n67718 = ~i_hbusreq6 & ~n67717;
  assign n67719 = ~n67626 & ~n67718;
  assign n67720 = ~controllable_hgrant6 & ~n67719;
  assign n67721 = ~n14173 & ~n67720;
  assign n67722 = ~controllable_hmaster0 & ~n67721;
  assign n67723 = ~n67625 & ~n67722;
  assign n67724 = ~i_hbusreq8 & ~n67723;
  assign n67725 = ~n67555 & ~n67724;
  assign n67726 = ~controllable_hmaster3 & ~n67725;
  assign n67727 = ~n67554 & ~n67726;
  assign n67728 = i_hlock7 & ~n67727;
  assign n67729 = i_hbusreq8 & ~n67368;
  assign n67730 = i_hbusreq6 & ~n67364;
  assign n67731 = ~n67579 & ~n67712;
  assign n67732 = controllable_hmaster1 & ~n67731;
  assign n67733 = ~n67619 & ~n67732;
  assign n67734 = ~i_hbusreq6 & ~n67733;
  assign n67735 = ~n67730 & ~n67734;
  assign n67736 = ~controllable_hgrant6 & ~n67735;
  assign n67737 = ~n14298 & ~n67736;
  assign n67738 = controllable_hmaster0 & ~n67737;
  assign n67739 = ~n67722 & ~n67738;
  assign n67740 = ~i_hbusreq8 & ~n67739;
  assign n67741 = ~n67729 & ~n67740;
  assign n67742 = ~controllable_hmaster3 & ~n67741;
  assign n67743 = ~n67554 & ~n67742;
  assign n67744 = ~i_hlock7 & ~n67743;
  assign n67745 = ~n67728 & ~n67744;
  assign n67746 = ~i_hbusreq7 & ~n67745;
  assign n67747 = ~n67373 & ~n67746;
  assign n67748 = n7924 & ~n67747;
  assign n67749 = ~n66887 & ~n67748;
  assign n67750 = ~n8214 & ~n67749;
  assign n67751 = i_hlock9 & ~n67237;
  assign n67752 = ~i_hlock9 & ~n67255;
  assign n67753 = ~n67751 & ~n67752;
  assign n67754 = ~controllable_hgrant4 & ~n67753;
  assign n67755 = ~n12609 & ~n67754;
  assign n67756 = ~controllable_hgrant5 & ~n67755;
  assign n67757 = ~n12608 & ~n67756;
  assign n67758 = ~controllable_hmaster2 & ~n67757;
  assign n67759 = ~n67201 & ~n67758;
  assign n67760 = ~controllable_hmaster1 & ~n67759;
  assign n67761 = ~n67200 & ~n67760;
  assign n67762 = ~controllable_hgrant6 & ~n67761;
  assign n67763 = ~n13122 & ~n67762;
  assign n67764 = controllable_hmaster0 & ~n67763;
  assign n67765 = ~controllable_hgrant4 & ~n67213;
  assign n67766 = ~n13408 & ~n67765;
  assign n67767 = ~controllable_hgrant5 & ~n67766;
  assign n67768 = ~n13407 & ~n67767;
  assign n67769 = ~controllable_hmaster2 & ~n67768;
  assign n67770 = ~n67201 & ~n67769;
  assign n67771 = ~controllable_hmaster1 & ~n67770;
  assign n67772 = ~n67200 & ~n67771;
  assign n67773 = ~controllable_hgrant6 & ~n67772;
  assign n67774 = ~n13406 & ~n67773;
  assign n67775 = ~controllable_hmaster0 & ~n67774;
  assign n67776 = ~n67764 & ~n67775;
  assign n67777 = i_hlock8 & ~n67776;
  assign n67778 = ~controllable_hgrant4 & ~n67219;
  assign n67779 = ~n13429 & ~n67778;
  assign n67780 = ~controllable_hgrant5 & ~n67779;
  assign n67781 = ~n13428 & ~n67780;
  assign n67782 = ~controllable_hmaster2 & ~n67781;
  assign n67783 = ~n67201 & ~n67782;
  assign n67784 = ~controllable_hmaster1 & ~n67783;
  assign n67785 = ~n67200 & ~n67784;
  assign n67786 = ~controllable_hgrant6 & ~n67785;
  assign n67787 = ~n13427 & ~n67786;
  assign n67788 = ~controllable_hmaster0 & ~n67787;
  assign n67789 = ~n67764 & ~n67788;
  assign n67790 = ~i_hlock8 & ~n67789;
  assign n67791 = ~n67777 & ~n67790;
  assign n67792 = controllable_hmaster3 & ~n67791;
  assign n67793 = ~n67359 & ~n67792;
  assign n67794 = i_hlock7 & ~n67793;
  assign n67795 = ~n67369 & ~n67792;
  assign n67796 = ~i_hlock7 & ~n67795;
  assign n67797 = ~n67794 & ~n67796;
  assign n67798 = i_hbusreq7 & ~n67797;
  assign n67799 = i_hbusreq8 & ~n67791;
  assign n67800 = i_hbusreq6 & ~n67761;
  assign n67801 = i_hbusreq5 & ~n67755;
  assign n67802 = i_hbusreq4 & ~n67753;
  assign n67803 = i_hbusreq9 & ~n67753;
  assign n67804 = i_hlock9 & ~n67493;
  assign n67805 = ~i_hlock9 & ~n67529;
  assign n67806 = ~n67804 & ~n67805;
  assign n67807 = ~i_hbusreq9 & ~n67806;
  assign n67808 = ~n67803 & ~n67807;
  assign n67809 = ~i_hbusreq4 & ~n67808;
  assign n67810 = ~n67802 & ~n67809;
  assign n67811 = ~controllable_hgrant4 & ~n67810;
  assign n67812 = ~n14322 & ~n67811;
  assign n67813 = ~i_hbusreq5 & ~n67812;
  assign n67814 = ~n67801 & ~n67813;
  assign n67815 = ~controllable_hgrant5 & ~n67814;
  assign n67816 = ~n14321 & ~n67815;
  assign n67817 = ~controllable_hmaster2 & ~n67816;
  assign n67818 = ~n67415 & ~n67817;
  assign n67819 = ~controllable_hmaster1 & ~n67818;
  assign n67820 = ~n67414 & ~n67819;
  assign n67821 = ~i_hbusreq6 & ~n67820;
  assign n67822 = ~n67800 & ~n67821;
  assign n67823 = ~controllable_hgrant6 & ~n67822;
  assign n67824 = ~n14320 & ~n67823;
  assign n67825 = controllable_hmaster0 & ~n67824;
  assign n67826 = i_hbusreq6 & ~n67772;
  assign n67827 = i_hbusreq5 & ~n67766;
  assign n67828 = i_hbusreq4 & ~n67213;
  assign n67829 = i_hbusreq9 & ~n67213;
  assign n67830 = ~i_hbusreq9 & ~n67445;
  assign n67831 = ~n67829 & ~n67830;
  assign n67832 = ~i_hbusreq4 & ~n67831;
  assign n67833 = ~n67828 & ~n67832;
  assign n67834 = ~controllable_hgrant4 & ~n67833;
  assign n67835 = ~n13524 & ~n67834;
  assign n67836 = ~i_hbusreq5 & ~n67835;
  assign n67837 = ~n67827 & ~n67836;
  assign n67838 = ~controllable_hgrant5 & ~n67837;
  assign n67839 = ~n13522 & ~n67838;
  assign n67840 = ~controllable_hmaster2 & ~n67839;
  assign n67841 = ~n67415 & ~n67840;
  assign n67842 = ~controllable_hmaster1 & ~n67841;
  assign n67843 = ~n67414 & ~n67842;
  assign n67844 = ~i_hbusreq6 & ~n67843;
  assign n67845 = ~n67826 & ~n67844;
  assign n67846 = ~controllable_hgrant6 & ~n67845;
  assign n67847 = ~n14443 & ~n67846;
  assign n67848 = ~controllable_hmaster0 & ~n67847;
  assign n67849 = ~n67825 & ~n67848;
  assign n67850 = i_hlock8 & ~n67849;
  assign n67851 = i_hbusreq6 & ~n67785;
  assign n67852 = i_hbusreq5 & ~n67779;
  assign n67853 = i_hbusreq4 & ~n67219;
  assign n67854 = i_hbusreq9 & ~n67219;
  assign n67855 = ~i_hbusreq9 & ~n67457;
  assign n67856 = ~n67854 & ~n67855;
  assign n67857 = ~i_hbusreq4 & ~n67856;
  assign n67858 = ~n67853 & ~n67857;
  assign n67859 = ~controllable_hgrant4 & ~n67858;
  assign n67860 = ~n13577 & ~n67859;
  assign n67861 = ~i_hbusreq5 & ~n67860;
  assign n67862 = ~n67852 & ~n67861;
  assign n67863 = ~controllable_hgrant5 & ~n67862;
  assign n67864 = ~n13575 & ~n67863;
  assign n67865 = ~controllable_hmaster2 & ~n67864;
  assign n67866 = ~n67415 & ~n67865;
  assign n67867 = ~controllable_hmaster1 & ~n67866;
  assign n67868 = ~n67414 & ~n67867;
  assign n67869 = ~i_hbusreq6 & ~n67868;
  assign n67870 = ~n67851 & ~n67869;
  assign n67871 = ~controllable_hgrant6 & ~n67870;
  assign n67872 = ~n14484 & ~n67871;
  assign n67873 = ~controllable_hmaster0 & ~n67872;
  assign n67874 = ~n67825 & ~n67873;
  assign n67875 = ~i_hlock8 & ~n67874;
  assign n67876 = ~n67850 & ~n67875;
  assign n67877 = ~i_hbusreq8 & ~n67876;
  assign n67878 = ~n67799 & ~n67877;
  assign n67879 = controllable_hmaster3 & ~n67878;
  assign n67880 = ~n67726 & ~n67879;
  assign n67881 = i_hlock7 & ~n67880;
  assign n67882 = ~n67742 & ~n67879;
  assign n67883 = ~i_hlock7 & ~n67882;
  assign n67884 = ~n67881 & ~n67883;
  assign n67885 = ~i_hbusreq7 & ~n67884;
  assign n67886 = ~n67798 & ~n67885;
  assign n67887 = n7924 & ~n67886;
  assign n67888 = ~n66999 & ~n67887;
  assign n67889 = n8214 & ~n67888;
  assign n67890 = ~n67750 & ~n67889;
  assign n67891 = ~n8202 & ~n67890;
  assign n67892 = ~n67248 & ~n67764;
  assign n67893 = i_hlock8 & ~n67892;
  assign n67894 = ~n67266 & ~n67764;
  assign n67895 = ~i_hlock8 & ~n67894;
  assign n67896 = ~n67893 & ~n67895;
  assign n67897 = controllable_hmaster3 & ~n67896;
  assign n67898 = controllable_hmaster2 & ~n67768;
  assign n67899 = ~n67281 & ~n67898;
  assign n67900 = controllable_hmaster1 & ~n67899;
  assign n67901 = ~n67303 & ~n67900;
  assign n67902 = ~controllable_hgrant6 & ~n67901;
  assign n67903 = ~n13849 & ~n67902;
  assign n67904 = controllable_hmaster0 & ~n67903;
  assign n67905 = ~n67357 & ~n67904;
  assign n67906 = ~controllable_hmaster3 & ~n67905;
  assign n67907 = ~n67897 & ~n67906;
  assign n67908 = i_hlock7 & ~n67907;
  assign n67909 = controllable_hmaster2 & ~n67781;
  assign n67910 = ~n67281 & ~n67909;
  assign n67911 = controllable_hmaster1 & ~n67910;
  assign n67912 = ~n67303 & ~n67911;
  assign n67913 = ~controllable_hgrant6 & ~n67912;
  assign n67914 = ~n13951 & ~n67913;
  assign n67915 = controllable_hmaster0 & ~n67914;
  assign n67916 = ~n67357 & ~n67915;
  assign n67917 = ~controllable_hmaster3 & ~n67916;
  assign n67918 = ~n67897 & ~n67917;
  assign n67919 = ~i_hlock7 & ~n67918;
  assign n67920 = ~n67908 & ~n67919;
  assign n67921 = i_hbusreq7 & ~n67920;
  assign n67922 = i_hbusreq8 & ~n67896;
  assign n67923 = ~n67512 & ~n67825;
  assign n67924 = i_hlock8 & ~n67923;
  assign n67925 = ~n67548 & ~n67825;
  assign n67926 = ~i_hlock8 & ~n67925;
  assign n67927 = ~n67924 & ~n67926;
  assign n67928 = ~i_hbusreq8 & ~n67927;
  assign n67929 = ~n67922 & ~n67928;
  assign n67930 = controllable_hmaster3 & ~n67929;
  assign n67931 = i_hbusreq8 & ~n67905;
  assign n67932 = i_hbusreq6 & ~n67901;
  assign n67933 = controllable_hmaster2 & ~n67839;
  assign n67934 = ~n67579 & ~n67933;
  assign n67935 = controllable_hmaster1 & ~n67934;
  assign n67936 = ~n67619 & ~n67935;
  assign n67937 = ~i_hbusreq6 & ~n67936;
  assign n67938 = ~n67932 & ~n67937;
  assign n67939 = ~controllable_hgrant6 & ~n67938;
  assign n67940 = ~n14756 & ~n67939;
  assign n67941 = controllable_hmaster0 & ~n67940;
  assign n67942 = ~n67722 & ~n67941;
  assign n67943 = ~i_hbusreq8 & ~n67942;
  assign n67944 = ~n67931 & ~n67943;
  assign n67945 = ~controllable_hmaster3 & ~n67944;
  assign n67946 = ~n67930 & ~n67945;
  assign n67947 = i_hlock7 & ~n67946;
  assign n67948 = i_hbusreq8 & ~n67916;
  assign n67949 = i_hbusreq6 & ~n67912;
  assign n67950 = controllable_hmaster2 & ~n67864;
  assign n67951 = ~n67579 & ~n67950;
  assign n67952 = controllable_hmaster1 & ~n67951;
  assign n67953 = ~n67619 & ~n67952;
  assign n67954 = ~i_hbusreq6 & ~n67953;
  assign n67955 = ~n67949 & ~n67954;
  assign n67956 = ~controllable_hgrant6 & ~n67955;
  assign n67957 = ~n14772 & ~n67956;
  assign n67958 = controllable_hmaster0 & ~n67957;
  assign n67959 = ~n67722 & ~n67958;
  assign n67960 = ~i_hbusreq8 & ~n67959;
  assign n67961 = ~n67948 & ~n67960;
  assign n67962 = ~controllable_hmaster3 & ~n67961;
  assign n67963 = ~n67930 & ~n67962;
  assign n67964 = ~i_hlock7 & ~n67963;
  assign n67965 = ~n67947 & ~n67964;
  assign n67966 = ~i_hbusreq7 & ~n67965;
  assign n67967 = ~n67921 & ~n67966;
  assign n67968 = n7924 & ~n67967;
  assign n67969 = ~n67045 & ~n67968;
  assign n67970 = ~n8214 & ~n67969;
  assign n67971 = ~n67317 & ~n67898;
  assign n67972 = controllable_hmaster1 & ~n67971;
  assign n67973 = ~n67346 & ~n67972;
  assign n67974 = i_hlock6 & ~n67973;
  assign n67975 = ~n67317 & ~n67909;
  assign n67976 = controllable_hmaster1 & ~n67975;
  assign n67977 = ~n67346 & ~n67976;
  assign n67978 = ~i_hlock6 & ~n67977;
  assign n67979 = ~n67974 & ~n67978;
  assign n67980 = ~controllable_hgrant6 & ~n67979;
  assign n67981 = ~n13894 & ~n67980;
  assign n67982 = ~controllable_hmaster0 & ~n67981;
  assign n67983 = ~n67307 & ~n67982;
  assign n67984 = ~controllable_hmaster3 & ~n67983;
  assign n67985 = ~n67897 & ~n67984;
  assign n67986 = i_hlock7 & ~n67985;
  assign n67987 = ~n67367 & ~n67982;
  assign n67988 = ~controllable_hmaster3 & ~n67987;
  assign n67989 = ~n67897 & ~n67988;
  assign n67990 = ~i_hlock7 & ~n67989;
  assign n67991 = ~n67986 & ~n67990;
  assign n67992 = i_hbusreq7 & ~n67991;
  assign n67993 = i_hbusreq8 & ~n67983;
  assign n67994 = i_hbusreq6 & ~n67979;
  assign n67995 = ~n67651 & ~n67933;
  assign n67996 = controllable_hmaster1 & ~n67995;
  assign n67997 = ~n67709 & ~n67996;
  assign n67998 = i_hlock6 & ~n67997;
  assign n67999 = ~n67651 & ~n67950;
  assign n68000 = controllable_hmaster1 & ~n67999;
  assign n68001 = ~n67709 & ~n68000;
  assign n68002 = ~i_hlock6 & ~n68001;
  assign n68003 = ~n67998 & ~n68002;
  assign n68004 = ~i_hbusreq6 & ~n68003;
  assign n68005 = ~n67994 & ~n68004;
  assign n68006 = ~controllable_hgrant6 & ~n68005;
  assign n68007 = ~n14802 & ~n68006;
  assign n68008 = ~controllable_hmaster0 & ~n68007;
  assign n68009 = ~n67625 & ~n68008;
  assign n68010 = ~i_hbusreq8 & ~n68009;
  assign n68011 = ~n67993 & ~n68010;
  assign n68012 = ~controllable_hmaster3 & ~n68011;
  assign n68013 = ~n67930 & ~n68012;
  assign n68014 = i_hlock7 & ~n68013;
  assign n68015 = i_hbusreq8 & ~n67987;
  assign n68016 = ~n67738 & ~n68008;
  assign n68017 = ~i_hbusreq8 & ~n68016;
  assign n68018 = ~n68015 & ~n68017;
  assign n68019 = ~controllable_hmaster3 & ~n68018;
  assign n68020 = ~n67930 & ~n68019;
  assign n68021 = ~i_hlock7 & ~n68020;
  assign n68022 = ~n68014 & ~n68021;
  assign n68023 = ~i_hbusreq7 & ~n68022;
  assign n68024 = ~n67992 & ~n68023;
  assign n68025 = n7924 & ~n68024;
  assign n68026 = ~n67122 & ~n68025;
  assign n68027 = n8214 & ~n68026;
  assign n68028 = ~n67970 & ~n68027;
  assign n68029 = n8202 & ~n68028;
  assign n68030 = ~n67891 & ~n68029;
  assign n68031 = n7920 & ~n68030;
  assign n68032 = ~n66580 & ~n68031;
  assign n68033 = n7728 & ~n68032;
  assign n68034 = ~n16354 & ~n66518;
  assign n68035 = ~controllable_hgrant1 & ~n68034;
  assign n68036 = ~n13924 & ~n68035;
  assign n68037 = ~controllable_hgrant3 & ~n68036;
  assign n68038 = ~n13923 & ~n68037;
  assign n68039 = ~controllable_hgrant4 & ~n68038;
  assign n68040 = ~n13922 & ~n68039;
  assign n68041 = ~controllable_hgrant5 & ~n68040;
  assign n68042 = ~n13921 & ~n68041;
  assign n68043 = ~controllable_hmaster2 & ~n68042;
  assign n68044 = ~n18169 & ~n68043;
  assign n68045 = ~controllable_hmaster1 & ~n68044;
  assign n68046 = ~n18161 & ~n68045;
  assign n68047 = i_hlock6 & ~n68046;
  assign n68048 = ~n18185 & ~n68045;
  assign n68049 = ~i_hlock6 & ~n68048;
  assign n68050 = ~n68047 & ~n68049;
  assign n68051 = ~controllable_hgrant6 & ~n68050;
  assign n68052 = ~n13894 & ~n68051;
  assign n68053 = ~controllable_hmaster0 & ~n68052;
  assign n68054 = ~n18149 & ~n68053;
  assign n68055 = ~controllable_hmaster3 & ~n68054;
  assign n68056 = ~n30151 & ~n68055;
  assign n68057 = i_hlock7 & ~n68056;
  assign n68058 = ~n18201 & ~n68053;
  assign n68059 = ~controllable_hmaster3 & ~n68058;
  assign n68060 = ~n30151 & ~n68059;
  assign n68061 = ~i_hlock7 & ~n68060;
  assign n68062 = ~n68057 & ~n68061;
  assign n68063 = i_hbusreq7 & ~n68062;
  assign n68064 = i_hbusreq8 & ~n68054;
  assign n68065 = i_hbusreq6 & ~n68050;
  assign n68066 = i_hbusreq5 & ~n68040;
  assign n68067 = i_hbusreq4 & ~n68038;
  assign n68068 = i_hbusreq9 & ~n68038;
  assign n68069 = i_hbusreq3 & ~n68036;
  assign n68070 = i_hbusreq1 & ~n68034;
  assign n68071 = ~n7733 & ~n66837;
  assign n68072 = ~n16352 & ~n68071;
  assign n68073 = n7928 & ~n68072;
  assign n68074 = ~n66518 & ~n68073;
  assign n68075 = ~i_hbusreq1 & ~n68074;
  assign n68076 = ~n68070 & ~n68075;
  assign n68077 = ~controllable_hgrant1 & ~n68076;
  assign n68078 = ~n15107 & ~n68077;
  assign n68079 = ~i_hbusreq3 & ~n68078;
  assign n68080 = ~n68069 & ~n68079;
  assign n68081 = ~controllable_hgrant3 & ~n68080;
  assign n68082 = ~n15106 & ~n68081;
  assign n68083 = ~i_hbusreq9 & ~n68082;
  assign n68084 = ~n68068 & ~n68083;
  assign n68085 = ~i_hbusreq4 & ~n68084;
  assign n68086 = ~n68067 & ~n68085;
  assign n68087 = ~controllable_hgrant4 & ~n68086;
  assign n68088 = ~n15105 & ~n68087;
  assign n68089 = ~i_hbusreq5 & ~n68088;
  assign n68090 = ~n68066 & ~n68089;
  assign n68091 = ~controllable_hgrant5 & ~n68090;
  assign n68092 = ~n15104 & ~n68091;
  assign n68093 = ~controllable_hmaster2 & ~n68092;
  assign n68094 = ~n21773 & ~n68093;
  assign n68095 = ~controllable_hmaster1 & ~n68094;
  assign n68096 = ~n21761 & ~n68095;
  assign n68097 = i_hlock6 & ~n68096;
  assign n68098 = ~n21801 & ~n68095;
  assign n68099 = ~i_hlock6 & ~n68098;
  assign n68100 = ~n68097 & ~n68099;
  assign n68101 = ~i_hbusreq6 & ~n68100;
  assign n68102 = ~n68065 & ~n68101;
  assign n68103 = ~controllable_hgrant6 & ~n68102;
  assign n68104 = ~n15063 & ~n68103;
  assign n68105 = ~controllable_hmaster0 & ~n68104;
  assign n68106 = ~n21739 & ~n68105;
  assign n68107 = ~i_hbusreq8 & ~n68106;
  assign n68108 = ~n68064 & ~n68107;
  assign n68109 = ~controllable_hmaster3 & ~n68108;
  assign n68110 = ~n32005 & ~n68109;
  assign n68111 = i_hlock7 & ~n68110;
  assign n68112 = i_hbusreq8 & ~n68058;
  assign n68113 = ~n21823 & ~n68105;
  assign n68114 = ~i_hbusreq8 & ~n68113;
  assign n68115 = ~n68112 & ~n68114;
  assign n68116 = ~controllable_hmaster3 & ~n68115;
  assign n68117 = ~n32005 & ~n68116;
  assign n68118 = ~i_hlock7 & ~n68117;
  assign n68119 = ~n68111 & ~n68118;
  assign n68120 = ~i_hbusreq7 & ~n68119;
  assign n68121 = ~n68063 & ~n68120;
  assign n68122 = ~n7924 & ~n68121;
  assign n68123 = ~n17092 & ~n67206;
  assign n68124 = n7928 & ~n68123;
  assign n68125 = ~n17461 & ~n68124;
  assign n68126 = ~controllable_hgrant1 & ~n68125;
  assign n68127 = ~n13155 & ~n68126;
  assign n68128 = ~controllable_hgrant3 & ~n68127;
  assign n68129 = ~n13154 & ~n68128;
  assign n68130 = ~controllable_hgrant4 & ~n68129;
  assign n68131 = ~n13153 & ~n68130;
  assign n68132 = ~controllable_hgrant5 & ~n68131;
  assign n68133 = ~n13152 & ~n68132;
  assign n68134 = controllable_hmaster1 & ~n68133;
  assign n68135 = controllable_hmaster2 & ~n68133;
  assign n68136 = ~n67226 & ~n68135;
  assign n68137 = ~controllable_hmaster1 & ~n68136;
  assign n68138 = ~n68134 & ~n68137;
  assign n68139 = ~controllable_hgrant6 & ~n68138;
  assign n68140 = ~n13122 & ~n68139;
  assign n68141 = controllable_hmaster0 & ~n68140;
  assign n68142 = ~n67769 & ~n68135;
  assign n68143 = ~controllable_hmaster1 & ~n68142;
  assign n68144 = ~n68134 & ~n68143;
  assign n68145 = ~controllable_hgrant6 & ~n68144;
  assign n68146 = ~n13406 & ~n68145;
  assign n68147 = ~controllable_hmaster0 & ~n68146;
  assign n68148 = ~n68141 & ~n68147;
  assign n68149 = i_hlock8 & ~n68148;
  assign n68150 = ~n67782 & ~n68135;
  assign n68151 = ~controllable_hmaster1 & ~n68150;
  assign n68152 = ~n68134 & ~n68151;
  assign n68153 = ~controllable_hgrant6 & ~n68152;
  assign n68154 = ~n13427 & ~n68153;
  assign n68155 = ~controllable_hmaster0 & ~n68154;
  assign n68156 = ~n68141 & ~n68155;
  assign n68157 = ~i_hlock8 & ~n68156;
  assign n68158 = ~n68149 & ~n68157;
  assign n68159 = controllable_hmaster3 & ~n68158;
  assign n68160 = i_hlock3 & ~n67211;
  assign n68161 = ~i_hlock3 & ~n67217;
  assign n68162 = ~n68160 & ~n68161;
  assign n68163 = ~controllable_hgrant3 & ~n68162;
  assign n68164 = ~n13852 & ~n68163;
  assign n68165 = ~controllable_hgrant4 & ~n68164;
  assign n68166 = ~n13851 & ~n68165;
  assign n68167 = ~controllable_hgrant5 & ~n68166;
  assign n68168 = ~n13850 & ~n68167;
  assign n68169 = ~controllable_hmaster2 & ~n68168;
  assign n68170 = ~n67898 & ~n68169;
  assign n68171 = controllable_hmaster1 & ~n68170;
  assign n68172 = i_hlock5 & ~n67766;
  assign n68173 = ~i_hlock5 & ~n67779;
  assign n68174 = ~n68172 & ~n68173;
  assign n68175 = ~controllable_hgrant5 & ~n68174;
  assign n68176 = ~n13865 & ~n68175;
  assign n68177 = controllable_hmaster2 & ~n68176;
  assign n68178 = i_hlock1 & ~n67209;
  assign n68179 = ~i_hlock1 & ~n67215;
  assign n68180 = ~n68178 & ~n68179;
  assign n68181 = ~controllable_hgrant1 & ~n68180;
  assign n68182 = ~n13875 & ~n68181;
  assign n68183 = ~controllable_hgrant3 & ~n68182;
  assign n68184 = ~n13874 & ~n68183;
  assign n68185 = ~controllable_hgrant4 & ~n68184;
  assign n68186 = ~n13873 & ~n68185;
  assign n68187 = ~controllable_hgrant5 & ~n68186;
  assign n68188 = ~n13872 & ~n68187;
  assign n68189 = ~controllable_hmaster2 & ~n68188;
  assign n68190 = ~n68177 & ~n68189;
  assign n68191 = ~controllable_hmaster1 & ~n68190;
  assign n68192 = ~n68171 & ~n68191;
  assign n68193 = ~controllable_hgrant6 & ~n68192;
  assign n68194 = ~n13849 & ~n68193;
  assign n68195 = controllable_hmaster0 & ~n68194;
  assign n68196 = ~n9213 & ~n67208;
  assign n68197 = ~controllable_hgrant1 & ~n68196;
  assign n68198 = ~n13898 & ~n68197;
  assign n68199 = ~controllable_hgrant3 & ~n68198;
  assign n68200 = ~n13897 & ~n68199;
  assign n68201 = ~controllable_hgrant4 & ~n68200;
  assign n68202 = ~n13896 & ~n68201;
  assign n68203 = ~controllable_hgrant5 & ~n68202;
  assign n68204 = ~n13895 & ~n68203;
  assign n68205 = ~controllable_hmaster2 & ~n68204;
  assign n68206 = ~n67898 & ~n68205;
  assign n68207 = controllable_hmaster1 & ~n68206;
  assign n68208 = i_hlock4 & ~n67213;
  assign n68209 = ~i_hlock4 & ~n67219;
  assign n68210 = ~n68208 & ~n68209;
  assign n68211 = ~controllable_hgrant4 & ~n68210;
  assign n68212 = ~n13912 & ~n68211;
  assign n68213 = ~controllable_hgrant5 & ~n68212;
  assign n68214 = ~n13911 & ~n68213;
  assign n68215 = controllable_hmaster2 & ~n68214;
  assign n68216 = ~i_hlock0 & ~n16639;
  assign n68217 = ~controllable_hgrant2 & n68216;
  assign n68218 = ~n7814 & ~n68217;
  assign n68219 = n7733 & ~n68218;
  assign n68220 = ~n16507 & ~n68219;
  assign n68221 = n7928 & ~n68220;
  assign n68222 = ~n66518 & ~n68221;
  assign n68223 = ~controllable_hgrant1 & ~n68222;
  assign n68224 = ~n13924 & ~n68223;
  assign n68225 = ~controllable_hgrant3 & ~n68224;
  assign n68226 = ~n13923 & ~n68225;
  assign n68227 = ~controllable_hgrant4 & ~n68226;
  assign n68228 = ~n13922 & ~n68227;
  assign n68229 = ~controllable_hgrant5 & ~n68228;
  assign n68230 = ~n13921 & ~n68229;
  assign n68231 = ~controllable_hmaster2 & ~n68230;
  assign n68232 = ~n68215 & ~n68231;
  assign n68233 = ~controllable_hmaster1 & ~n68232;
  assign n68234 = ~n68207 & ~n68233;
  assign n68235 = i_hlock6 & ~n68234;
  assign n68236 = ~n67909 & ~n68205;
  assign n68237 = controllable_hmaster1 & ~n68236;
  assign n68238 = ~n68233 & ~n68237;
  assign n68239 = ~i_hlock6 & ~n68238;
  assign n68240 = ~n68235 & ~n68239;
  assign n68241 = ~controllable_hgrant6 & ~n68240;
  assign n68242 = ~n13894 & ~n68241;
  assign n68243 = ~controllable_hmaster0 & ~n68242;
  assign n68244 = ~n68195 & ~n68243;
  assign n68245 = ~controllable_hmaster3 & ~n68244;
  assign n68246 = ~n68159 & ~n68245;
  assign n68247 = i_hlock7 & ~n68246;
  assign n68248 = ~n67909 & ~n68169;
  assign n68249 = controllable_hmaster1 & ~n68248;
  assign n68250 = ~n68191 & ~n68249;
  assign n68251 = ~controllable_hgrant6 & ~n68250;
  assign n68252 = ~n13951 & ~n68251;
  assign n68253 = controllable_hmaster0 & ~n68252;
  assign n68254 = ~n68243 & ~n68253;
  assign n68255 = ~controllable_hmaster3 & ~n68254;
  assign n68256 = ~n68159 & ~n68255;
  assign n68257 = ~i_hlock7 & ~n68256;
  assign n68258 = ~n68247 & ~n68257;
  assign n68259 = i_hbusreq7 & ~n68258;
  assign n68260 = i_hbusreq8 & ~n68158;
  assign n68261 = i_hbusreq6 & ~n68138;
  assign n68262 = i_hbusreq5 & ~n68131;
  assign n68263 = i_hbusreq4 & ~n68129;
  assign n68264 = i_hbusreq9 & ~n68129;
  assign n68265 = i_hbusreq3 & ~n68127;
  assign n68266 = i_hbusreq1 & ~n68125;
  assign n68267 = ~n12615 & ~n67424;
  assign n68268 = i_hlock0 & ~n68267;
  assign n68269 = ~n18726 & ~n68268;
  assign n68270 = ~i_hbusreq0 & ~n68269;
  assign n68271 = ~n67422 & ~n68270;
  assign n68272 = ~i_hbusreq2 & ~n68271;
  assign n68273 = ~n67421 & ~n68272;
  assign n68274 = ~controllable_hgrant2 & n68273;
  assign n68275 = ~n12706 & ~n68274;
  assign n68276 = n7733 & ~n68275;
  assign n68277 = ~n21845 & ~n68276;
  assign n68278 = n7928 & ~n68277;
  assign n68279 = ~n21834 & ~n68278;
  assign n68280 = ~i_hbusreq1 & ~n68279;
  assign n68281 = ~n68266 & ~n68280;
  assign n68282 = ~controllable_hgrant1 & ~n68281;
  assign n68283 = ~n14877 & ~n68282;
  assign n68284 = ~i_hbusreq3 & ~n68283;
  assign n68285 = ~n68265 & ~n68284;
  assign n68286 = ~controllable_hgrant3 & ~n68285;
  assign n68287 = ~n14876 & ~n68286;
  assign n68288 = ~i_hbusreq9 & ~n68287;
  assign n68289 = ~n68264 & ~n68288;
  assign n68290 = ~i_hbusreq4 & ~n68289;
  assign n68291 = ~n68263 & ~n68290;
  assign n68292 = ~controllable_hgrant4 & ~n68291;
  assign n68293 = ~n14875 & ~n68292;
  assign n68294 = ~i_hbusreq5 & ~n68293;
  assign n68295 = ~n68262 & ~n68294;
  assign n68296 = ~controllable_hgrant5 & ~n68295;
  assign n68297 = ~n14874 & ~n68296;
  assign n68298 = controllable_hmaster1 & ~n68297;
  assign n68299 = controllable_hmaster2 & ~n68297;
  assign n68300 = ~n18800 & ~n68276;
  assign n68301 = n7928 & ~n68300;
  assign n68302 = ~n8265 & ~n68301;
  assign n68303 = ~i_hbusreq1 & ~n68302;
  assign n68304 = ~n67420 & ~n68303;
  assign n68305 = ~controllable_hgrant1 & ~n68304;
  assign n68306 = ~n12681 & ~n68305;
  assign n68307 = ~i_hbusreq3 & ~n68306;
  assign n68308 = ~n67419 & ~n68307;
  assign n68309 = ~controllable_hgrant3 & ~n68308;
  assign n68310 = ~n12679 & ~n68309;
  assign n68311 = i_hlock9 & ~n68310;
  assign n68312 = ~n8297 & ~n68301;
  assign n68313 = ~i_hbusreq1 & ~n68312;
  assign n68314 = ~n67448 & ~n68313;
  assign n68315 = ~controllable_hgrant1 & ~n68314;
  assign n68316 = ~n12730 & ~n68315;
  assign n68317 = ~i_hbusreq3 & ~n68316;
  assign n68318 = ~n67447 & ~n68317;
  assign n68319 = ~controllable_hgrant3 & ~n68318;
  assign n68320 = ~n12728 & ~n68319;
  assign n68321 = ~i_hlock9 & ~n68320;
  assign n68322 = ~n68311 & ~n68321;
  assign n68323 = ~i_hbusreq9 & ~n68322;
  assign n68324 = ~n67418 & ~n68323;
  assign n68325 = ~i_hbusreq4 & ~n68324;
  assign n68326 = ~n67417 & ~n68325;
  assign n68327 = ~controllable_hgrant4 & ~n68326;
  assign n68328 = ~n12676 & ~n68327;
  assign n68329 = ~i_hbusreq5 & ~n68328;
  assign n68330 = ~n67416 & ~n68329;
  assign n68331 = ~controllable_hgrant5 & ~n68330;
  assign n68332 = ~n12674 & ~n68331;
  assign n68333 = ~controllable_hmaster2 & ~n68332;
  assign n68334 = ~n68299 & ~n68333;
  assign n68335 = ~controllable_hmaster1 & ~n68334;
  assign n68336 = ~n68298 & ~n68335;
  assign n68337 = ~i_hbusreq6 & ~n68336;
  assign n68338 = ~n68261 & ~n68337;
  assign n68339 = ~controllable_hgrant6 & ~n68338;
  assign n68340 = ~n14849 & ~n68339;
  assign n68341 = controllable_hmaster0 & ~n68340;
  assign n68342 = i_hbusreq6 & ~n68144;
  assign n68343 = ~i_hbusreq9 & ~n68310;
  assign n68344 = ~n67829 & ~n68343;
  assign n68345 = ~i_hbusreq4 & ~n68344;
  assign n68346 = ~n67828 & ~n68345;
  assign n68347 = ~controllable_hgrant4 & ~n68346;
  assign n68348 = ~n13524 & ~n68347;
  assign n68349 = ~i_hbusreq5 & ~n68348;
  assign n68350 = ~n67827 & ~n68349;
  assign n68351 = ~controllable_hgrant5 & ~n68350;
  assign n68352 = ~n13522 & ~n68351;
  assign n68353 = ~controllable_hmaster2 & ~n68352;
  assign n68354 = ~n68299 & ~n68353;
  assign n68355 = ~controllable_hmaster1 & ~n68354;
  assign n68356 = ~n68298 & ~n68355;
  assign n68357 = ~i_hbusreq6 & ~n68356;
  assign n68358 = ~n68342 & ~n68357;
  assign n68359 = ~controllable_hgrant6 & ~n68358;
  assign n68360 = ~n14927 & ~n68359;
  assign n68361 = ~controllable_hmaster0 & ~n68360;
  assign n68362 = ~n68341 & ~n68361;
  assign n68363 = i_hlock8 & ~n68362;
  assign n68364 = i_hbusreq6 & ~n68152;
  assign n68365 = ~i_hbusreq9 & ~n68320;
  assign n68366 = ~n67854 & ~n68365;
  assign n68367 = ~i_hbusreq4 & ~n68366;
  assign n68368 = ~n67853 & ~n68367;
  assign n68369 = ~controllable_hgrant4 & ~n68368;
  assign n68370 = ~n13577 & ~n68369;
  assign n68371 = ~i_hbusreq5 & ~n68370;
  assign n68372 = ~n67852 & ~n68371;
  assign n68373 = ~controllable_hgrant5 & ~n68372;
  assign n68374 = ~n13575 & ~n68373;
  assign n68375 = ~controllable_hmaster2 & ~n68374;
  assign n68376 = ~n68299 & ~n68375;
  assign n68377 = ~controllable_hmaster1 & ~n68376;
  assign n68378 = ~n68298 & ~n68377;
  assign n68379 = ~i_hbusreq6 & ~n68378;
  assign n68380 = ~n68364 & ~n68379;
  assign n68381 = ~controllable_hgrant6 & ~n68380;
  assign n68382 = ~n14960 & ~n68381;
  assign n68383 = ~controllable_hmaster0 & ~n68382;
  assign n68384 = ~n68341 & ~n68383;
  assign n68385 = ~i_hlock8 & ~n68384;
  assign n68386 = ~n68363 & ~n68385;
  assign n68387 = ~i_hbusreq8 & ~n68386;
  assign n68388 = ~n68260 & ~n68387;
  assign n68389 = controllable_hmaster3 & ~n68388;
  assign n68390 = i_hbusreq8 & ~n68244;
  assign n68391 = i_hbusreq6 & ~n68192;
  assign n68392 = controllable_hmaster2 & ~n68352;
  assign n68393 = i_hbusreq5 & ~n68166;
  assign n68394 = i_hbusreq4 & ~n68164;
  assign n68395 = i_hbusreq9 & ~n68164;
  assign n68396 = i_hbusreq3 & ~n68162;
  assign n68397 = i_hlock3 & ~n68306;
  assign n68398 = ~i_hlock3 & ~n68316;
  assign n68399 = ~n68397 & ~n68398;
  assign n68400 = ~i_hbusreq3 & ~n68399;
  assign n68401 = ~n68396 & ~n68400;
  assign n68402 = ~controllable_hgrant3 & ~n68401;
  assign n68403 = ~n14999 & ~n68402;
  assign n68404 = ~i_hbusreq9 & ~n68403;
  assign n68405 = ~n68395 & ~n68404;
  assign n68406 = ~i_hbusreq4 & ~n68405;
  assign n68407 = ~n68394 & ~n68406;
  assign n68408 = ~controllable_hgrant4 & ~n68407;
  assign n68409 = ~n14998 & ~n68408;
  assign n68410 = ~i_hbusreq5 & ~n68409;
  assign n68411 = ~n68393 & ~n68410;
  assign n68412 = ~controllable_hgrant5 & ~n68411;
  assign n68413 = ~n14997 & ~n68412;
  assign n68414 = ~controllable_hmaster2 & ~n68413;
  assign n68415 = ~n68392 & ~n68414;
  assign n68416 = controllable_hmaster1 & ~n68415;
  assign n68417 = i_hbusreq5 & ~n68174;
  assign n68418 = i_hlock5 & ~n68348;
  assign n68419 = ~i_hlock5 & ~n68370;
  assign n68420 = ~n68418 & ~n68419;
  assign n68421 = ~i_hbusreq5 & ~n68420;
  assign n68422 = ~n68417 & ~n68421;
  assign n68423 = ~controllable_hgrant5 & ~n68422;
  assign n68424 = ~n15020 & ~n68423;
  assign n68425 = controllable_hmaster2 & ~n68424;
  assign n68426 = i_hbusreq5 & ~n68186;
  assign n68427 = i_hbusreq4 & ~n68184;
  assign n68428 = i_hbusreq9 & ~n68184;
  assign n68429 = i_hbusreq3 & ~n68182;
  assign n68430 = i_hbusreq1 & ~n68180;
  assign n68431 = i_hlock1 & ~n68302;
  assign n68432 = ~i_hlock1 & ~n68312;
  assign n68433 = ~n68431 & ~n68432;
  assign n68434 = ~i_hbusreq1 & ~n68433;
  assign n68435 = ~n68430 & ~n68434;
  assign n68436 = ~controllable_hgrant1 & ~n68435;
  assign n68437 = ~n15032 & ~n68436;
  assign n68438 = ~i_hbusreq3 & ~n68437;
  assign n68439 = ~n68429 & ~n68438;
  assign n68440 = ~controllable_hgrant3 & ~n68439;
  assign n68441 = ~n15031 & ~n68440;
  assign n68442 = ~i_hbusreq9 & ~n68441;
  assign n68443 = ~n68428 & ~n68442;
  assign n68444 = ~i_hbusreq4 & ~n68443;
  assign n68445 = ~n68427 & ~n68444;
  assign n68446 = ~controllable_hgrant4 & ~n68445;
  assign n68447 = ~n15030 & ~n68446;
  assign n68448 = ~i_hbusreq5 & ~n68447;
  assign n68449 = ~n68426 & ~n68448;
  assign n68450 = ~controllable_hgrant5 & ~n68449;
  assign n68451 = ~n15029 & ~n68450;
  assign n68452 = ~controllable_hmaster2 & ~n68451;
  assign n68453 = ~n68425 & ~n68452;
  assign n68454 = ~controllable_hmaster1 & ~n68453;
  assign n68455 = ~n68416 & ~n68454;
  assign n68456 = ~i_hbusreq6 & ~n68455;
  assign n68457 = ~n68391 & ~n68456;
  assign n68458 = ~controllable_hgrant6 & ~n68457;
  assign n68459 = ~n14995 & ~n68458;
  assign n68460 = controllable_hmaster0 & ~n68459;
  assign n68461 = i_hbusreq6 & ~n68240;
  assign n68462 = i_hbusreq5 & ~n68202;
  assign n68463 = i_hbusreq4 & ~n68200;
  assign n68464 = i_hbusreq9 & ~n68200;
  assign n68465 = i_hbusreq3 & ~n68198;
  assign n68466 = i_hbusreq1 & ~n68196;
  assign n68467 = ~n9379 & ~n68301;
  assign n68468 = ~i_hbusreq1 & ~n68467;
  assign n68469 = ~n68466 & ~n68468;
  assign n68470 = ~controllable_hgrant1 & ~n68469;
  assign n68471 = ~n15067 & ~n68470;
  assign n68472 = ~i_hbusreq3 & ~n68471;
  assign n68473 = ~n68465 & ~n68472;
  assign n68474 = ~controllable_hgrant3 & ~n68473;
  assign n68475 = ~n15066 & ~n68474;
  assign n68476 = ~i_hbusreq9 & ~n68475;
  assign n68477 = ~n68464 & ~n68476;
  assign n68478 = ~i_hbusreq4 & ~n68477;
  assign n68479 = ~n68463 & ~n68478;
  assign n68480 = ~controllable_hgrant4 & ~n68479;
  assign n68481 = ~n15065 & ~n68480;
  assign n68482 = ~i_hbusreq5 & ~n68481;
  assign n68483 = ~n68462 & ~n68482;
  assign n68484 = ~controllable_hgrant5 & ~n68483;
  assign n68485 = ~n15064 & ~n68484;
  assign n68486 = ~controllable_hmaster2 & ~n68485;
  assign n68487 = ~n68392 & ~n68486;
  assign n68488 = controllable_hmaster1 & ~n68487;
  assign n68489 = i_hbusreq5 & ~n68212;
  assign n68490 = i_hbusreq4 & ~n68210;
  assign n68491 = i_hlock4 & ~n68344;
  assign n68492 = ~i_hlock4 & ~n68366;
  assign n68493 = ~n68491 & ~n68492;
  assign n68494 = ~i_hbusreq4 & ~n68493;
  assign n68495 = ~n68490 & ~n68494;
  assign n68496 = ~controllable_hgrant4 & ~n68495;
  assign n68497 = ~n15091 & ~n68496;
  assign n68498 = ~i_hbusreq5 & ~n68497;
  assign n68499 = ~n68489 & ~n68498;
  assign n68500 = ~controllable_hgrant5 & ~n68499;
  assign n68501 = ~n15090 & ~n68500;
  assign n68502 = controllable_hmaster2 & ~n68501;
  assign n68503 = i_hbusreq5 & ~n68228;
  assign n68504 = i_hbusreq4 & ~n68226;
  assign n68505 = i_hbusreq9 & ~n68226;
  assign n68506 = i_hbusreq3 & ~n68224;
  assign n68507 = i_hbusreq1 & ~n68222;
  assign n68508 = ~n67673 & ~n68219;
  assign n68509 = n7928 & ~n68508;
  assign n68510 = ~n66518 & ~n68509;
  assign n68511 = ~i_hbusreq1 & ~n68510;
  assign n68512 = ~n68507 & ~n68511;
  assign n68513 = ~controllable_hgrant1 & ~n68512;
  assign n68514 = ~n15107 & ~n68513;
  assign n68515 = ~i_hbusreq3 & ~n68514;
  assign n68516 = ~n68506 & ~n68515;
  assign n68517 = ~controllable_hgrant3 & ~n68516;
  assign n68518 = ~n15106 & ~n68517;
  assign n68519 = ~i_hbusreq9 & ~n68518;
  assign n68520 = ~n68505 & ~n68519;
  assign n68521 = ~i_hbusreq4 & ~n68520;
  assign n68522 = ~n68504 & ~n68521;
  assign n68523 = ~controllable_hgrant4 & ~n68522;
  assign n68524 = ~n15105 & ~n68523;
  assign n68525 = ~i_hbusreq5 & ~n68524;
  assign n68526 = ~n68503 & ~n68525;
  assign n68527 = ~controllable_hgrant5 & ~n68526;
  assign n68528 = ~n15104 & ~n68527;
  assign n68529 = ~controllable_hmaster2 & ~n68528;
  assign n68530 = ~n68502 & ~n68529;
  assign n68531 = ~controllable_hmaster1 & ~n68530;
  assign n68532 = ~n68488 & ~n68531;
  assign n68533 = i_hlock6 & ~n68532;
  assign n68534 = controllable_hmaster2 & ~n68374;
  assign n68535 = ~n68486 & ~n68534;
  assign n68536 = controllable_hmaster1 & ~n68535;
  assign n68537 = ~n68531 & ~n68536;
  assign n68538 = ~i_hlock6 & ~n68537;
  assign n68539 = ~n68533 & ~n68538;
  assign n68540 = ~i_hbusreq6 & ~n68539;
  assign n68541 = ~n68461 & ~n68540;
  assign n68542 = ~controllable_hgrant6 & ~n68541;
  assign n68543 = ~n15063 & ~n68542;
  assign n68544 = ~controllable_hmaster0 & ~n68543;
  assign n68545 = ~n68460 & ~n68544;
  assign n68546 = ~i_hbusreq8 & ~n68545;
  assign n68547 = ~n68390 & ~n68546;
  assign n68548 = ~controllable_hmaster3 & ~n68547;
  assign n68549 = ~n68389 & ~n68548;
  assign n68550 = i_hlock7 & ~n68549;
  assign n68551 = i_hbusreq8 & ~n68254;
  assign n68552 = i_hbusreq6 & ~n68250;
  assign n68553 = ~n68414 & ~n68534;
  assign n68554 = controllable_hmaster1 & ~n68553;
  assign n68555 = ~n68454 & ~n68554;
  assign n68556 = ~i_hbusreq6 & ~n68555;
  assign n68557 = ~n68552 & ~n68556;
  assign n68558 = ~controllable_hgrant6 & ~n68557;
  assign n68559 = ~n15152 & ~n68558;
  assign n68560 = controllable_hmaster0 & ~n68559;
  assign n68561 = ~n68544 & ~n68560;
  assign n68562 = ~i_hbusreq8 & ~n68561;
  assign n68563 = ~n68551 & ~n68562;
  assign n68564 = ~controllable_hmaster3 & ~n68563;
  assign n68565 = ~n68389 & ~n68564;
  assign n68566 = ~i_hlock7 & ~n68565;
  assign n68567 = ~n68550 & ~n68566;
  assign n68568 = ~i_hbusreq7 & ~n68567;
  assign n68569 = ~n68259 & ~n68568;
  assign n68570 = n7924 & ~n68569;
  assign n68571 = ~n68122 & ~n68570;
  assign n68572 = n7920 & ~n68571;
  assign n68573 = ~n66580 & ~n68572;
  assign n68574 = ~n7728 & ~n68573;
  assign n68575 = ~n68033 & ~n68574;
  assign n68576 = ~n7723 & ~n68575;
  assign n68577 = ~n67183 & ~n68576;
  assign n68578 = ~n7714 & ~n68577;
  assign n68579 = ~n67182 & ~n68578;
  assign n68580 = ~n7705 & ~n68579;
  assign n68581 = ~n66603 & ~n68580;
  assign n68582 = n7808 & ~n68581;
  assign n68583 = ~n66589 & ~n68582;
  assign n68584 = n8195 & ~n68583;
  assign n68585 = ~n8196 & ~n68584;
  assign n68586 = ~n8193 & ~n68585;
  assign n68587 = ~n9900 & ~n66580;
  assign n68588 = ~n7723 & ~n68587;
  assign n68589 = ~n9899 & ~n68588;
  assign n68590 = n7714 & ~n68589;
  assign n68591 = ~n66585 & ~n68590;
  assign n68592 = ~n7705 & ~n68591;
  assign n68593 = ~n9898 & ~n68592;
  assign n68594 = ~n7808 & ~n68593;
  assign n68595 = ~n22405 & ~n36100;
  assign n68596 = ~controllable_hmaster3 & ~n68595;
  assign n68597 = ~n9093 & ~n68596;
  assign n68598 = i_hbusreq7 & ~n68597;
  assign n68599 = i_hbusreq8 & ~n68595;
  assign n68600 = ~n22419 & ~n66614;
  assign n68601 = ~i_hbusreq8 & ~n68600;
  assign n68602 = ~n68599 & ~n68601;
  assign n68603 = ~controllable_hmaster3 & ~n68602;
  assign n68604 = ~n9117 & ~n68603;
  assign n68605 = ~i_hbusreq7 & ~n68604;
  assign n68606 = ~n68598 & ~n68605;
  assign n68607 = ~n7924 & ~n68606;
  assign n68608 = ~n22439 & ~n36116;
  assign n68609 = ~controllable_hmaster3 & ~n68608;
  assign n68610 = ~n27088 & ~n68609;
  assign n68611 = i_hbusreq7 & ~n68610;
  assign n68612 = i_hbusreq8 & ~n68608;
  assign n68613 = ~n22462 & ~n66633;
  assign n68614 = ~i_hbusreq8 & ~n68613;
  assign n68615 = ~n68612 & ~n68614;
  assign n68616 = ~controllable_hmaster3 & ~n68615;
  assign n68617 = ~n27174 & ~n68616;
  assign n68618 = ~i_hbusreq7 & ~n68617;
  assign n68619 = ~n68611 & ~n68618;
  assign n68620 = n7924 & ~n68619;
  assign n68621 = ~n68607 & ~n68620;
  assign n68622 = ~n8214 & ~n68621;
  assign n68623 = ~n13322 & ~n18169;
  assign n68624 = ~controllable_hmaster1 & ~n68623;
  assign n68625 = ~n10053 & ~n68624;
  assign n68626 = ~controllable_hgrant6 & ~n68625;
  assign n68627 = ~n15241 & ~n68626;
  assign n68628 = ~controllable_hmaster0 & ~n68627;
  assign n68629 = ~n9152 & ~n68628;
  assign n68630 = ~controllable_hmaster3 & ~n68629;
  assign n68631 = ~n9093 & ~n68630;
  assign n68632 = i_hbusreq7 & ~n68631;
  assign n68633 = i_hbusreq8 & ~n68629;
  assign n68634 = i_hbusreq6 & ~n68625;
  assign n68635 = ~n13369 & ~n21773;
  assign n68636 = ~controllable_hmaster1 & ~n68635;
  assign n68637 = ~n10064 & ~n68636;
  assign n68638 = ~i_hbusreq6 & ~n68637;
  assign n68639 = ~n68634 & ~n68638;
  assign n68640 = ~controllable_hgrant6 & ~n68639;
  assign n68641 = ~n15253 & ~n68640;
  assign n68642 = ~controllable_hmaster0 & ~n68641;
  assign n68643 = ~n9162 & ~n68642;
  assign n68644 = ~i_hbusreq8 & ~n68643;
  assign n68645 = ~n68633 & ~n68644;
  assign n68646 = ~controllable_hmaster3 & ~n68645;
  assign n68647 = ~n9117 & ~n68646;
  assign n68648 = ~i_hbusreq7 & ~n68647;
  assign n68649 = ~n68632 & ~n68648;
  assign n68650 = ~n7924 & ~n68649;
  assign n68651 = ~n13399 & ~n22508;
  assign n68652 = ~controllable_hmaster1 & ~n68651;
  assign n68653 = ~n15194 & ~n68652;
  assign n68654 = ~controllable_hgrant6 & ~n68653;
  assign n68655 = ~n15241 & ~n68654;
  assign n68656 = ~controllable_hmaster0 & ~n68655;
  assign n68657 = ~n13765 & ~n68656;
  assign n68658 = ~controllable_hmaster3 & ~n68657;
  assign n68659 = ~n27088 & ~n68658;
  assign n68660 = i_hbusreq7 & ~n68659;
  assign n68661 = i_hbusreq8 & ~n68657;
  assign n68662 = i_hbusreq6 & ~n68653;
  assign n68663 = ~n13511 & ~n22534;
  assign n68664 = ~controllable_hmaster1 & ~n68663;
  assign n68665 = ~n15208 & ~n68664;
  assign n68666 = ~i_hbusreq6 & ~n68665;
  assign n68667 = ~n68662 & ~n68666;
  assign n68668 = ~controllable_hgrant6 & ~n68667;
  assign n68669 = ~n15253 & ~n68668;
  assign n68670 = ~controllable_hmaster0 & ~n68669;
  assign n68671 = ~n13778 & ~n68670;
  assign n68672 = ~i_hbusreq8 & ~n68671;
  assign n68673 = ~n68661 & ~n68672;
  assign n68674 = ~controllable_hmaster3 & ~n68673;
  assign n68675 = ~n27174 & ~n68674;
  assign n68676 = ~i_hbusreq7 & ~n68675;
  assign n68677 = ~n68660 & ~n68676;
  assign n68678 = n7924 & ~n68677;
  assign n68679 = ~n68650 & ~n68678;
  assign n68680 = n8214 & ~n68679;
  assign n68681 = ~n68622 & ~n68680;
  assign n68682 = ~n8202 & ~n68681;
  assign n68683 = ~n22560 & ~n36100;
  assign n68684 = ~controllable_hmaster3 & ~n68683;
  assign n68685 = ~n9093 & ~n68684;
  assign n68686 = i_hbusreq7 & ~n68685;
  assign n68687 = i_hbusreq8 & ~n68683;
  assign n68688 = ~n22574 & ~n66614;
  assign n68689 = ~i_hbusreq8 & ~n68688;
  assign n68690 = ~n68687 & ~n68689;
  assign n68691 = ~controllable_hmaster3 & ~n68690;
  assign n68692 = ~n9117 & ~n68691;
  assign n68693 = ~i_hbusreq7 & ~n68692;
  assign n68694 = ~n68686 & ~n68693;
  assign n68695 = ~n7924 & ~n68694;
  assign n68696 = ~n22598 & ~n36116;
  assign n68697 = ~controllable_hmaster3 & ~n68696;
  assign n68698 = ~n27088 & ~n68697;
  assign n68699 = i_hbusreq7 & ~n68698;
  assign n68700 = i_hbusreq8 & ~n68696;
  assign n68701 = ~n22634 & ~n66633;
  assign n68702 = ~i_hbusreq8 & ~n68701;
  assign n68703 = ~n68700 & ~n68702;
  assign n68704 = ~controllable_hmaster3 & ~n68703;
  assign n68705 = ~n27174 & ~n68704;
  assign n68706 = ~i_hbusreq7 & ~n68705;
  assign n68707 = ~n68699 & ~n68706;
  assign n68708 = n7924 & ~n68707;
  assign n68709 = ~n68695 & ~n68708;
  assign n68710 = ~n8214 & ~n68709;
  assign n68711 = ~n15662 & ~n22646;
  assign n68712 = ~controllable_hgrant6 & ~n68711;
  assign n68713 = ~n15351 & ~n68712;
  assign n68714 = ~controllable_hmaster0 & ~n68713;
  assign n68715 = ~n9152 & ~n68714;
  assign n68716 = ~controllable_hmaster3 & ~n68715;
  assign n68717 = ~n9093 & ~n68716;
  assign n68718 = i_hbusreq7 & ~n68717;
  assign n68719 = i_hbusreq8 & ~n68715;
  assign n68720 = i_hbusreq6 & ~n68711;
  assign n68721 = ~n22658 & ~n66608;
  assign n68722 = ~i_hbusreq6 & ~n68721;
  assign n68723 = ~n68720 & ~n68722;
  assign n68724 = ~controllable_hgrant6 & ~n68723;
  assign n68725 = ~n15363 & ~n68724;
  assign n68726 = ~controllable_hmaster0 & ~n68725;
  assign n68727 = ~n9162 & ~n68726;
  assign n68728 = ~i_hbusreq8 & ~n68727;
  assign n68729 = ~n68719 & ~n68728;
  assign n68730 = ~controllable_hmaster3 & ~n68729;
  assign n68731 = ~n9117 & ~n68730;
  assign n68732 = ~i_hbusreq7 & ~n68731;
  assign n68733 = ~n68718 & ~n68732;
  assign n68734 = ~n7924 & ~n68733;
  assign n68735 = ~n15716 & ~n22684;
  assign n68736 = ~controllable_hgrant6 & ~n68735;
  assign n68737 = ~n15351 & ~n68736;
  assign n68738 = ~controllable_hmaster0 & ~n68737;
  assign n68739 = ~n13765 & ~n68738;
  assign n68740 = ~controllable_hmaster3 & ~n68739;
  assign n68741 = ~n27088 & ~n68740;
  assign n68742 = i_hbusreq7 & ~n68741;
  assign n68743 = i_hbusreq8 & ~n68739;
  assign n68744 = i_hbusreq6 & ~n68735;
  assign n68745 = ~n22721 & ~n66627;
  assign n68746 = ~i_hbusreq6 & ~n68745;
  assign n68747 = ~n68744 & ~n68746;
  assign n68748 = ~controllable_hgrant6 & ~n68747;
  assign n68749 = ~n15363 & ~n68748;
  assign n68750 = ~controllable_hmaster0 & ~n68749;
  assign n68751 = ~n13778 & ~n68750;
  assign n68752 = ~i_hbusreq8 & ~n68751;
  assign n68753 = ~n68743 & ~n68752;
  assign n68754 = ~controllable_hmaster3 & ~n68753;
  assign n68755 = ~n27174 & ~n68754;
  assign n68756 = ~i_hbusreq7 & ~n68755;
  assign n68757 = ~n68742 & ~n68756;
  assign n68758 = n7924 & ~n68757;
  assign n68759 = ~n68734 & ~n68758;
  assign n68760 = n8214 & ~n68759;
  assign n68761 = ~n68710 & ~n68760;
  assign n68762 = n8202 & ~n68761;
  assign n68763 = ~n68682 & ~n68762;
  assign n68764 = n7920 & ~n68763;
  assign n68765 = ~n10014 & ~n68764;
  assign n68766 = n7728 & ~n68765;
  assign n68767 = ~n22749 & ~n66809;
  assign n68768 = ~controllable_hmaster3 & ~n68767;
  assign n68769 = ~n30877 & ~n68768;
  assign n68770 = i_hlock7 & ~n68769;
  assign n68771 = ~n22757 & ~n66809;
  assign n68772 = ~controllable_hmaster3 & ~n68771;
  assign n68773 = ~n30877 & ~n68772;
  assign n68774 = ~i_hlock7 & ~n68773;
  assign n68775 = ~n68770 & ~n68774;
  assign n68776 = i_hbusreq7 & ~n68775;
  assign n68777 = i_hbusreq8 & ~n68767;
  assign n68778 = ~n22773 & ~n66870;
  assign n68779 = ~i_hbusreq8 & ~n68778;
  assign n68780 = ~n68777 & ~n68779;
  assign n68781 = ~controllable_hmaster3 & ~n68780;
  assign n68782 = ~n30896 & ~n68781;
  assign n68783 = i_hlock7 & ~n68782;
  assign n68784 = i_hbusreq8 & ~n68771;
  assign n68785 = ~n22787 & ~n66870;
  assign n68786 = ~i_hbusreq8 & ~n68785;
  assign n68787 = ~n68784 & ~n68786;
  assign n68788 = ~controllable_hmaster3 & ~n68787;
  assign n68789 = ~n30896 & ~n68788;
  assign n68790 = ~i_hlock7 & ~n68789;
  assign n68791 = ~n68783 & ~n68790;
  assign n68792 = ~i_hbusreq7 & ~n68791;
  assign n68793 = ~n68776 & ~n68792;
  assign n68794 = ~n7924 & ~n68793;
  assign n68795 = ~n22809 & ~n66907;
  assign n68796 = ~controllable_hmaster3 & ~n68795;
  assign n68797 = ~n30920 & ~n68796;
  assign n68798 = i_hlock7 & ~n68797;
  assign n68799 = ~n22817 & ~n66907;
  assign n68800 = ~controllable_hmaster3 & ~n68799;
  assign n68801 = ~n30920 & ~n68800;
  assign n68802 = ~i_hlock7 & ~n68801;
  assign n68803 = ~n68798 & ~n68802;
  assign n68804 = i_hbusreq7 & ~n68803;
  assign n68805 = i_hbusreq8 & ~n68795;
  assign n68806 = ~n22842 & ~n66966;
  assign n68807 = ~i_hbusreq8 & ~n68806;
  assign n68808 = ~n68805 & ~n68807;
  assign n68809 = ~controllable_hmaster3 & ~n68808;
  assign n68810 = ~n30939 & ~n68809;
  assign n68811 = i_hlock7 & ~n68810;
  assign n68812 = i_hbusreq8 & ~n68799;
  assign n68813 = ~n22856 & ~n66966;
  assign n68814 = ~i_hbusreq8 & ~n68813;
  assign n68815 = ~n68812 & ~n68814;
  assign n68816 = ~controllable_hmaster3 & ~n68815;
  assign n68817 = ~n30939 & ~n68816;
  assign n68818 = ~i_hlock7 & ~n68817;
  assign n68819 = ~n68811 & ~n68818;
  assign n68820 = ~i_hbusreq7 & ~n68819;
  assign n68821 = ~n68804 & ~n68820;
  assign n68822 = n7924 & ~n68821;
  assign n68823 = ~n68794 & ~n68822;
  assign n68824 = ~n8214 & ~n68823;
  assign n68825 = ~n18169 & ~n66799;
  assign n68826 = ~controllable_hmaster1 & ~n68825;
  assign n68827 = ~n19291 & ~n68826;
  assign n68828 = i_hlock6 & ~n68827;
  assign n68829 = ~n19318 & ~n68826;
  assign n68830 = ~i_hlock6 & ~n68829;
  assign n68831 = ~n68828 & ~n68830;
  assign n68832 = ~controllable_hgrant6 & ~n68831;
  assign n68833 = ~n13894 & ~n68832;
  assign n68834 = ~controllable_hmaster0 & ~n68833;
  assign n68835 = ~n19279 & ~n68834;
  assign n68836 = ~controllable_hmaster3 & ~n68835;
  assign n68837 = ~n30877 & ~n68836;
  assign n68838 = i_hlock7 & ~n68837;
  assign n68839 = ~n19334 & ~n68834;
  assign n68840 = ~controllable_hmaster3 & ~n68839;
  assign n68841 = ~n30877 & ~n68840;
  assign n68842 = ~i_hlock7 & ~n68841;
  assign n68843 = ~n68838 & ~n68842;
  assign n68844 = i_hbusreq7 & ~n68843;
  assign n68845 = i_hbusreq8 & ~n68835;
  assign n68846 = i_hbusreq6 & ~n68831;
  assign n68847 = ~n21773 & ~n66858;
  assign n68848 = ~controllable_hmaster1 & ~n68847;
  assign n68849 = ~n19584 & ~n68848;
  assign n68850 = i_hlock6 & ~n68849;
  assign n68851 = ~n19636 & ~n68848;
  assign n68852 = ~i_hlock6 & ~n68851;
  assign n68853 = ~n68850 & ~n68852;
  assign n68854 = ~i_hbusreq6 & ~n68853;
  assign n68855 = ~n68846 & ~n68854;
  assign n68856 = ~controllable_hgrant6 & ~n68855;
  assign n68857 = ~n15467 & ~n68856;
  assign n68858 = ~controllable_hmaster0 & ~n68857;
  assign n68859 = ~n19556 & ~n68858;
  assign n68860 = ~i_hbusreq8 & ~n68859;
  assign n68861 = ~n68845 & ~n68860;
  assign n68862 = ~controllable_hmaster3 & ~n68861;
  assign n68863 = ~n30896 & ~n68862;
  assign n68864 = i_hlock7 & ~n68863;
  assign n68865 = i_hbusreq8 & ~n68839;
  assign n68866 = ~n19660 & ~n68858;
  assign n68867 = ~i_hbusreq8 & ~n68866;
  assign n68868 = ~n68865 & ~n68867;
  assign n68869 = ~controllable_hmaster3 & ~n68868;
  assign n68870 = ~n30896 & ~n68869;
  assign n68871 = ~i_hlock7 & ~n68870;
  assign n68872 = ~n68864 & ~n68871;
  assign n68873 = ~i_hbusreq7 & ~n68872;
  assign n68874 = ~n68844 & ~n68873;
  assign n68875 = ~n7924 & ~n68874;
  assign n68876 = ~n22927 & ~n66897;
  assign n68877 = ~controllable_hmaster1 & ~n68876;
  assign n68878 = ~n19816 & ~n68877;
  assign n68879 = i_hlock6 & ~n68878;
  assign n68880 = ~n19843 & ~n68877;
  assign n68881 = ~i_hlock6 & ~n68880;
  assign n68882 = ~n68879 & ~n68881;
  assign n68883 = ~controllable_hgrant6 & ~n68882;
  assign n68884 = ~n13894 & ~n68883;
  assign n68885 = ~controllable_hmaster0 & ~n68884;
  assign n68886 = ~n19804 & ~n68885;
  assign n68887 = ~controllable_hmaster3 & ~n68886;
  assign n68888 = ~n30920 & ~n68887;
  assign n68889 = i_hlock7 & ~n68888;
  assign n68890 = ~n19859 & ~n68885;
  assign n68891 = ~controllable_hmaster3 & ~n68890;
  assign n68892 = ~n30920 & ~n68891;
  assign n68893 = ~i_hlock7 & ~n68892;
  assign n68894 = ~n68889 & ~n68893;
  assign n68895 = i_hbusreq7 & ~n68894;
  assign n68896 = i_hbusreq8 & ~n68886;
  assign n68897 = i_hbusreq6 & ~n68882;
  assign n68898 = ~n22963 & ~n66954;
  assign n68899 = ~controllable_hmaster1 & ~n68898;
  assign n68900 = ~n20177 & ~n68899;
  assign n68901 = i_hlock6 & ~n68900;
  assign n68902 = ~n20229 & ~n68899;
  assign n68903 = ~i_hlock6 & ~n68902;
  assign n68904 = ~n68901 & ~n68903;
  assign n68905 = ~i_hbusreq6 & ~n68904;
  assign n68906 = ~n68897 & ~n68905;
  assign n68907 = ~controllable_hgrant6 & ~n68906;
  assign n68908 = ~n15467 & ~n68907;
  assign n68909 = ~controllable_hmaster0 & ~n68908;
  assign n68910 = ~n20149 & ~n68909;
  assign n68911 = ~i_hbusreq8 & ~n68910;
  assign n68912 = ~n68896 & ~n68911;
  assign n68913 = ~controllable_hmaster3 & ~n68912;
  assign n68914 = ~n30939 & ~n68913;
  assign n68915 = i_hlock7 & ~n68914;
  assign n68916 = i_hbusreq8 & ~n68890;
  assign n68917 = ~n20253 & ~n68909;
  assign n68918 = ~i_hbusreq8 & ~n68917;
  assign n68919 = ~n68916 & ~n68918;
  assign n68920 = ~controllable_hmaster3 & ~n68919;
  assign n68921 = ~n30939 & ~n68920;
  assign n68922 = ~i_hlock7 & ~n68921;
  assign n68923 = ~n68915 & ~n68922;
  assign n68924 = ~i_hbusreq7 & ~n68923;
  assign n68925 = ~n68895 & ~n68924;
  assign n68926 = n7924 & ~n68925;
  assign n68927 = ~n68875 & ~n68926;
  assign n68928 = n8214 & ~n68927;
  assign n68929 = ~n68824 & ~n68928;
  assign n68930 = ~n8202 & ~n68929;
  assign n68931 = ~n23002 & ~n66809;
  assign n68932 = ~controllable_hmaster3 & ~n68931;
  assign n68933 = ~n30877 & ~n68932;
  assign n68934 = i_hlock7 & ~n68933;
  assign n68935 = ~n23012 & ~n66809;
  assign n68936 = ~controllable_hmaster3 & ~n68935;
  assign n68937 = ~n30877 & ~n68936;
  assign n68938 = ~i_hlock7 & ~n68937;
  assign n68939 = ~n68934 & ~n68938;
  assign n68940 = i_hbusreq7 & ~n68939;
  assign n68941 = i_hbusreq8 & ~n68931;
  assign n68942 = ~n23028 & ~n66870;
  assign n68943 = ~i_hbusreq8 & ~n68942;
  assign n68944 = ~n68941 & ~n68943;
  assign n68945 = ~controllable_hmaster3 & ~n68944;
  assign n68946 = ~n30896 & ~n68945;
  assign n68947 = i_hlock7 & ~n68946;
  assign n68948 = i_hbusreq8 & ~n68935;
  assign n68949 = ~n23044 & ~n66870;
  assign n68950 = ~i_hbusreq8 & ~n68949;
  assign n68951 = ~n68948 & ~n68950;
  assign n68952 = ~controllable_hmaster3 & ~n68951;
  assign n68953 = ~n30896 & ~n68952;
  assign n68954 = ~i_hlock7 & ~n68953;
  assign n68955 = ~n68947 & ~n68954;
  assign n68956 = ~i_hbusreq7 & ~n68955;
  assign n68957 = ~n68940 & ~n68956;
  assign n68958 = ~n7924 & ~n68957;
  assign n68959 = ~n23070 & ~n66907;
  assign n68960 = ~controllable_hmaster3 & ~n68959;
  assign n68961 = ~n30920 & ~n68960;
  assign n68962 = i_hlock7 & ~n68961;
  assign n68963 = ~n23080 & ~n66907;
  assign n68964 = ~controllable_hmaster3 & ~n68963;
  assign n68965 = ~n30920 & ~n68964;
  assign n68966 = ~i_hlock7 & ~n68965;
  assign n68967 = ~n68962 & ~n68966;
  assign n68968 = i_hbusreq7 & ~n68967;
  assign n68969 = i_hbusreq8 & ~n68959;
  assign n68970 = ~n23118 & ~n66966;
  assign n68971 = ~i_hbusreq8 & ~n68970;
  assign n68972 = ~n68969 & ~n68971;
  assign n68973 = ~controllable_hmaster3 & ~n68972;
  assign n68974 = ~n30939 & ~n68973;
  assign n68975 = i_hlock7 & ~n68974;
  assign n68976 = i_hbusreq8 & ~n68963;
  assign n68977 = ~n23134 & ~n66966;
  assign n68978 = ~i_hbusreq8 & ~n68977;
  assign n68979 = ~n68976 & ~n68978;
  assign n68980 = ~controllable_hmaster3 & ~n68979;
  assign n68981 = ~n30939 & ~n68980;
  assign n68982 = ~i_hlock7 & ~n68981;
  assign n68983 = ~n68975 & ~n68982;
  assign n68984 = ~i_hbusreq7 & ~n68983;
  assign n68985 = ~n68968 & ~n68984;
  assign n68986 = n7924 & ~n68985;
  assign n68987 = ~n68958 & ~n68986;
  assign n68988 = ~n8214 & ~n68987;
  assign n68989 = ~n23148 & ~n66801;
  assign n68990 = i_hlock6 & ~n68989;
  assign n68991 = ~n23152 & ~n66801;
  assign n68992 = ~i_hlock6 & ~n68991;
  assign n68993 = ~n68990 & ~n68992;
  assign n68994 = ~controllable_hgrant6 & ~n68993;
  assign n68995 = ~n13894 & ~n68994;
  assign n68996 = ~controllable_hmaster0 & ~n68995;
  assign n68997 = ~n19279 & ~n68996;
  assign n68998 = ~controllable_hmaster3 & ~n68997;
  assign n68999 = ~n30877 & ~n68998;
  assign n69000 = i_hlock7 & ~n68999;
  assign n69001 = ~n19334 & ~n68996;
  assign n69002 = ~controllable_hmaster3 & ~n69001;
  assign n69003 = ~n30877 & ~n69002;
  assign n69004 = ~i_hlock7 & ~n69003;
  assign n69005 = ~n69000 & ~n69004;
  assign n69006 = i_hbusreq7 & ~n69005;
  assign n69007 = i_hbusreq8 & ~n68997;
  assign n69008 = i_hbusreq6 & ~n68993;
  assign n69009 = ~n23172 & ~n66860;
  assign n69010 = i_hlock6 & ~n69009;
  assign n69011 = ~n23176 & ~n66860;
  assign n69012 = ~i_hlock6 & ~n69011;
  assign n69013 = ~n69010 & ~n69012;
  assign n69014 = ~i_hbusreq6 & ~n69013;
  assign n69015 = ~n69008 & ~n69014;
  assign n69016 = ~controllable_hgrant6 & ~n69015;
  assign n69017 = ~n15582 & ~n69016;
  assign n69018 = ~controllable_hmaster0 & ~n69017;
  assign n69019 = ~n19556 & ~n69018;
  assign n69020 = ~i_hbusreq8 & ~n69019;
  assign n69021 = ~n69007 & ~n69020;
  assign n69022 = ~controllable_hmaster3 & ~n69021;
  assign n69023 = ~n30896 & ~n69022;
  assign n69024 = i_hlock7 & ~n69023;
  assign n69025 = i_hbusreq8 & ~n69001;
  assign n69026 = ~n19660 & ~n69018;
  assign n69027 = ~i_hbusreq8 & ~n69026;
  assign n69028 = ~n69025 & ~n69027;
  assign n69029 = ~controllable_hmaster3 & ~n69028;
  assign n69030 = ~n30896 & ~n69029;
  assign n69031 = ~i_hlock7 & ~n69030;
  assign n69032 = ~n69024 & ~n69031;
  assign n69033 = ~i_hbusreq7 & ~n69032;
  assign n69034 = ~n69006 & ~n69033;
  assign n69035 = ~n7924 & ~n69034;
  assign n69036 = ~n23213 & ~n66899;
  assign n69037 = i_hlock6 & ~n69036;
  assign n69038 = ~n23217 & ~n66899;
  assign n69039 = ~i_hlock6 & ~n69038;
  assign n69040 = ~n69037 & ~n69039;
  assign n69041 = ~controllable_hgrant6 & ~n69040;
  assign n69042 = ~n13894 & ~n69041;
  assign n69043 = ~controllable_hmaster0 & ~n69042;
  assign n69044 = ~n19804 & ~n69043;
  assign n69045 = ~controllable_hmaster3 & ~n69044;
  assign n69046 = ~n30920 & ~n69045;
  assign n69047 = i_hlock7 & ~n69046;
  assign n69048 = ~n19859 & ~n69043;
  assign n69049 = ~controllable_hmaster3 & ~n69048;
  assign n69050 = ~n30920 & ~n69049;
  assign n69051 = ~i_hlock7 & ~n69050;
  assign n69052 = ~n69047 & ~n69051;
  assign n69053 = i_hbusreq7 & ~n69052;
  assign n69054 = i_hbusreq8 & ~n69044;
  assign n69055 = i_hbusreq6 & ~n69040;
  assign n69056 = ~n23262 & ~n66956;
  assign n69057 = i_hlock6 & ~n69056;
  assign n69058 = ~n23266 & ~n66956;
  assign n69059 = ~i_hlock6 & ~n69058;
  assign n69060 = ~n69057 & ~n69059;
  assign n69061 = ~i_hbusreq6 & ~n69060;
  assign n69062 = ~n69055 & ~n69061;
  assign n69063 = ~controllable_hgrant6 & ~n69062;
  assign n69064 = ~n15582 & ~n69063;
  assign n69065 = ~controllable_hmaster0 & ~n69064;
  assign n69066 = ~n20149 & ~n69065;
  assign n69067 = ~i_hbusreq8 & ~n69066;
  assign n69068 = ~n69054 & ~n69067;
  assign n69069 = ~controllable_hmaster3 & ~n69068;
  assign n69070 = ~n30939 & ~n69069;
  assign n69071 = i_hlock7 & ~n69070;
  assign n69072 = i_hbusreq8 & ~n69048;
  assign n69073 = ~n20253 & ~n69065;
  assign n69074 = ~i_hbusreq8 & ~n69073;
  assign n69075 = ~n69072 & ~n69074;
  assign n69076 = ~controllable_hmaster3 & ~n69075;
  assign n69077 = ~n30939 & ~n69076;
  assign n69078 = ~i_hlock7 & ~n69077;
  assign n69079 = ~n69071 & ~n69078;
  assign n69080 = ~i_hbusreq7 & ~n69079;
  assign n69081 = ~n69053 & ~n69080;
  assign n69082 = n7924 & ~n69081;
  assign n69083 = ~n69035 & ~n69082;
  assign n69084 = n8214 & ~n69083;
  assign n69085 = ~n68988 & ~n69084;
  assign n69086 = n8202 & ~n69085;
  assign n69087 = ~n68930 & ~n69086;
  assign n69088 = n7920 & ~n69087;
  assign n69089 = ~n10014 & ~n69088;
  assign n69090 = ~n7728 & ~n69089;
  assign n69091 = ~n68766 & ~n69090;
  assign n69092 = n7723 & ~n69091;
  assign n69093 = ~n7723 & ~n69089;
  assign n69094 = ~n69092 & ~n69093;
  assign n69095 = n7714 & ~n69094;
  assign n69096 = n7723 & ~n69089;
  assign n69097 = ~n67301 & ~n68177;
  assign n69098 = ~controllable_hmaster1 & ~n69097;
  assign n69099 = ~n67283 & ~n69098;
  assign n69100 = ~controllable_hgrant6 & ~n69099;
  assign n69101 = ~n13849 & ~n69100;
  assign n69102 = controllable_hmaster0 & ~n69101;
  assign n69103 = ~n67357 & ~n69102;
  assign n69104 = ~controllable_hmaster3 & ~n69103;
  assign n69105 = ~n67897 & ~n69104;
  assign n69106 = i_hlock7 & ~n69105;
  assign n69107 = ~n67363 & ~n69098;
  assign n69108 = ~controllable_hgrant6 & ~n69107;
  assign n69109 = ~n13951 & ~n69108;
  assign n69110 = controllable_hmaster0 & ~n69109;
  assign n69111 = ~n67357 & ~n69110;
  assign n69112 = ~controllable_hmaster3 & ~n69111;
  assign n69113 = ~n67897 & ~n69112;
  assign n69114 = ~i_hlock7 & ~n69113;
  assign n69115 = ~n69106 & ~n69114;
  assign n69116 = i_hbusreq7 & ~n69115;
  assign n69117 = i_hbusreq8 & ~n69103;
  assign n69118 = i_hbusreq6 & ~n69099;
  assign n69119 = i_hlock5 & ~n67835;
  assign n69120 = ~i_hlock5 & ~n67860;
  assign n69121 = ~n69119 & ~n69120;
  assign n69122 = ~i_hbusreq5 & ~n69121;
  assign n69123 = ~n68417 & ~n69122;
  assign n69124 = ~controllable_hgrant5 & ~n69123;
  assign n69125 = ~n15020 & ~n69124;
  assign n69126 = controllable_hmaster2 & ~n69125;
  assign n69127 = ~n67617 & ~n69126;
  assign n69128 = ~controllable_hmaster1 & ~n69127;
  assign n69129 = ~n67581 & ~n69128;
  assign n69130 = ~i_hbusreq6 & ~n69129;
  assign n69131 = ~n69118 & ~n69130;
  assign n69132 = ~controllable_hgrant6 & ~n69131;
  assign n69133 = ~n15417 & ~n69132;
  assign n69134 = controllable_hmaster0 & ~n69133;
  assign n69135 = ~n67722 & ~n69134;
  assign n69136 = ~i_hbusreq8 & ~n69135;
  assign n69137 = ~n69117 & ~n69136;
  assign n69138 = ~controllable_hmaster3 & ~n69137;
  assign n69139 = ~n67930 & ~n69138;
  assign n69140 = i_hlock7 & ~n69139;
  assign n69141 = i_hbusreq8 & ~n69111;
  assign n69142 = i_hbusreq6 & ~n69107;
  assign n69143 = ~n67732 & ~n69128;
  assign n69144 = ~i_hbusreq6 & ~n69143;
  assign n69145 = ~n69142 & ~n69144;
  assign n69146 = ~controllable_hgrant6 & ~n69145;
  assign n69147 = ~n15440 & ~n69146;
  assign n69148 = controllable_hmaster0 & ~n69147;
  assign n69149 = ~n67722 & ~n69148;
  assign n69150 = ~i_hbusreq8 & ~n69149;
  assign n69151 = ~n69141 & ~n69150;
  assign n69152 = ~controllable_hmaster3 & ~n69151;
  assign n69153 = ~n67930 & ~n69152;
  assign n69154 = ~i_hlock7 & ~n69153;
  assign n69155 = ~n69140 & ~n69154;
  assign n69156 = ~i_hbusreq7 & ~n69155;
  assign n69157 = ~n69116 & ~n69156;
  assign n69158 = n7924 & ~n69157;
  assign n69159 = ~n68794 & ~n69158;
  assign n69160 = ~n8214 & ~n69159;
  assign n69161 = ~n67344 & ~n68215;
  assign n69162 = ~controllable_hmaster1 & ~n69161;
  assign n69163 = ~n67319 & ~n69162;
  assign n69164 = i_hlock6 & ~n69163;
  assign n69165 = ~n67351 & ~n69162;
  assign n69166 = ~i_hlock6 & ~n69165;
  assign n69167 = ~n69164 & ~n69166;
  assign n69168 = ~controllable_hgrant6 & ~n69167;
  assign n69169 = ~n13894 & ~n69168;
  assign n69170 = ~controllable_hmaster0 & ~n69169;
  assign n69171 = ~n67307 & ~n69170;
  assign n69172 = ~controllable_hmaster3 & ~n69171;
  assign n69173 = ~n67897 & ~n69172;
  assign n69174 = i_hlock7 & ~n69173;
  assign n69175 = ~n67367 & ~n69170;
  assign n69176 = ~controllable_hmaster3 & ~n69175;
  assign n69177 = ~n67897 & ~n69176;
  assign n69178 = ~i_hlock7 & ~n69177;
  assign n69179 = ~n69174 & ~n69178;
  assign n69180 = i_hbusreq7 & ~n69179;
  assign n69181 = i_hbusreq8 & ~n69171;
  assign n69182 = i_hbusreq6 & ~n69167;
  assign n69183 = i_hlock4 & ~n67831;
  assign n69184 = ~i_hlock4 & ~n67856;
  assign n69185 = ~n69183 & ~n69184;
  assign n69186 = ~i_hbusreq4 & ~n69185;
  assign n69187 = ~n68490 & ~n69186;
  assign n69188 = ~controllable_hgrant4 & ~n69187;
  assign n69189 = ~n15091 & ~n69188;
  assign n69190 = ~i_hbusreq5 & ~n69189;
  assign n69191 = ~n68489 & ~n69190;
  assign n69192 = ~controllable_hgrant5 & ~n69191;
  assign n69193 = ~n15090 & ~n69192;
  assign n69194 = controllable_hmaster2 & ~n69193;
  assign n69195 = ~n67707 & ~n69194;
  assign n69196 = ~controllable_hmaster1 & ~n69195;
  assign n69197 = ~n67653 & ~n69196;
  assign n69198 = i_hlock6 & ~n69197;
  assign n69199 = ~n67714 & ~n69196;
  assign n69200 = ~i_hlock6 & ~n69199;
  assign n69201 = ~n69198 & ~n69200;
  assign n69202 = ~i_hbusreq6 & ~n69201;
  assign n69203 = ~n69182 & ~n69202;
  assign n69204 = ~controllable_hgrant6 & ~n69203;
  assign n69205 = ~n15467 & ~n69204;
  assign n69206 = ~controllable_hmaster0 & ~n69205;
  assign n69207 = ~n67625 & ~n69206;
  assign n69208 = ~i_hbusreq8 & ~n69207;
  assign n69209 = ~n69181 & ~n69208;
  assign n69210 = ~controllable_hmaster3 & ~n69209;
  assign n69211 = ~n67930 & ~n69210;
  assign n69212 = i_hlock7 & ~n69211;
  assign n69213 = i_hbusreq8 & ~n69175;
  assign n69214 = ~n67738 & ~n69206;
  assign n69215 = ~i_hbusreq8 & ~n69214;
  assign n69216 = ~n69213 & ~n69215;
  assign n69217 = ~controllable_hmaster3 & ~n69216;
  assign n69218 = ~n67930 & ~n69217;
  assign n69219 = ~i_hlock7 & ~n69218;
  assign n69220 = ~n69212 & ~n69219;
  assign n69221 = ~i_hbusreq7 & ~n69220;
  assign n69222 = ~n69180 & ~n69221;
  assign n69223 = n7924 & ~n69222;
  assign n69224 = ~n68875 & ~n69223;
  assign n69225 = n8214 & ~n69224;
  assign n69226 = ~n69160 & ~n69225;
  assign n69227 = ~n8202 & ~n69226;
  assign n69228 = ~n67271 & ~n68169;
  assign n69229 = controllable_hmaster1 & ~n69228;
  assign n69230 = ~n67303 & ~n69229;
  assign n69231 = ~controllable_hgrant6 & ~n69230;
  assign n69232 = ~n13849 & ~n69231;
  assign n69233 = controllable_hmaster0 & ~n69232;
  assign n69234 = ~n67357 & ~n69233;
  assign n69235 = ~controllable_hmaster3 & ~n69234;
  assign n69236 = ~n67897 & ~n69235;
  assign n69237 = i_hlock7 & ~n69236;
  assign n69238 = ~n67349 & ~n68169;
  assign n69239 = controllable_hmaster1 & ~n69238;
  assign n69240 = ~n67303 & ~n69239;
  assign n69241 = ~controllable_hgrant6 & ~n69240;
  assign n69242 = ~n13951 & ~n69241;
  assign n69243 = controllable_hmaster0 & ~n69242;
  assign n69244 = ~n67357 & ~n69243;
  assign n69245 = ~controllable_hmaster3 & ~n69244;
  assign n69246 = ~n67897 & ~n69245;
  assign n69247 = ~i_hlock7 & ~n69246;
  assign n69248 = ~n69237 & ~n69247;
  assign n69249 = i_hbusreq7 & ~n69248;
  assign n69250 = i_hbusreq8 & ~n69234;
  assign n69251 = i_hbusreq6 & ~n69230;
  assign n69252 = i_hlock3 & ~n67441;
  assign n69253 = ~i_hlock3 & ~n67453;
  assign n69254 = ~n69252 & ~n69253;
  assign n69255 = ~i_hbusreq3 & ~n69254;
  assign n69256 = ~n68396 & ~n69255;
  assign n69257 = ~controllable_hgrant3 & ~n69256;
  assign n69258 = ~n14999 & ~n69257;
  assign n69259 = ~i_hbusreq9 & ~n69258;
  assign n69260 = ~n68395 & ~n69259;
  assign n69261 = ~i_hbusreq4 & ~n69260;
  assign n69262 = ~n68394 & ~n69261;
  assign n69263 = ~controllable_hgrant4 & ~n69262;
  assign n69264 = ~n14998 & ~n69263;
  assign n69265 = ~i_hbusreq5 & ~n69264;
  assign n69266 = ~n68393 & ~n69265;
  assign n69267 = ~controllable_hgrant5 & ~n69266;
  assign n69268 = ~n14997 & ~n69267;
  assign n69269 = ~controllable_hmaster2 & ~n69268;
  assign n69270 = ~n67557 & ~n69269;
  assign n69271 = controllable_hmaster1 & ~n69270;
  assign n69272 = ~n67619 & ~n69271;
  assign n69273 = ~i_hbusreq6 & ~n69272;
  assign n69274 = ~n69251 & ~n69273;
  assign n69275 = ~controllable_hgrant6 & ~n69274;
  assign n69276 = ~n15520 & ~n69275;
  assign n69277 = controllable_hmaster0 & ~n69276;
  assign n69278 = ~n67722 & ~n69277;
  assign n69279 = ~i_hbusreq8 & ~n69278;
  assign n69280 = ~n69250 & ~n69279;
  assign n69281 = ~controllable_hmaster3 & ~n69280;
  assign n69282 = ~n67930 & ~n69281;
  assign n69283 = i_hlock7 & ~n69282;
  assign n69284 = i_hbusreq8 & ~n69244;
  assign n69285 = i_hbusreq6 & ~n69240;
  assign n69286 = ~n67712 & ~n69269;
  assign n69287 = controllable_hmaster1 & ~n69286;
  assign n69288 = ~n67619 & ~n69287;
  assign n69289 = ~i_hbusreq6 & ~n69288;
  assign n69290 = ~n69285 & ~n69289;
  assign n69291 = ~controllable_hgrant6 & ~n69290;
  assign n69292 = ~n15553 & ~n69291;
  assign n69293 = controllable_hmaster0 & ~n69292;
  assign n69294 = ~n67722 & ~n69293;
  assign n69295 = ~i_hbusreq8 & ~n69294;
  assign n69296 = ~n69284 & ~n69295;
  assign n69297 = ~controllable_hmaster3 & ~n69296;
  assign n69298 = ~n67930 & ~n69297;
  assign n69299 = ~i_hlock7 & ~n69298;
  assign n69300 = ~n69283 & ~n69299;
  assign n69301 = ~i_hbusreq7 & ~n69300;
  assign n69302 = ~n69249 & ~n69301;
  assign n69303 = n7924 & ~n69302;
  assign n69304 = ~n68958 & ~n69303;
  assign n69305 = ~n8214 & ~n69304;
  assign n69306 = ~n67271 & ~n68205;
  assign n69307 = controllable_hmaster1 & ~n69306;
  assign n69308 = ~n67346 & ~n69307;
  assign n69309 = i_hlock6 & ~n69308;
  assign n69310 = ~n67349 & ~n68205;
  assign n69311 = controllable_hmaster1 & ~n69310;
  assign n69312 = ~n67346 & ~n69311;
  assign n69313 = ~i_hlock6 & ~n69312;
  assign n69314 = ~n69309 & ~n69313;
  assign n69315 = ~controllable_hgrant6 & ~n69314;
  assign n69316 = ~n13894 & ~n69315;
  assign n69317 = ~controllable_hmaster0 & ~n69316;
  assign n69318 = ~n67307 & ~n69317;
  assign n69319 = ~controllable_hmaster3 & ~n69318;
  assign n69320 = ~n67897 & ~n69319;
  assign n69321 = i_hlock7 & ~n69320;
  assign n69322 = ~n67367 & ~n69317;
  assign n69323 = ~controllable_hmaster3 & ~n69322;
  assign n69324 = ~n67897 & ~n69323;
  assign n69325 = ~i_hlock7 & ~n69324;
  assign n69326 = ~n69321 & ~n69325;
  assign n69327 = i_hbusreq7 & ~n69326;
  assign n69328 = i_hbusreq8 & ~n69318;
  assign n69329 = i_hbusreq6 & ~n69314;
  assign n69330 = ~n9379 & ~n67436;
  assign n69331 = ~i_hbusreq1 & ~n69330;
  assign n69332 = ~n68466 & ~n69331;
  assign n69333 = ~controllable_hgrant1 & ~n69332;
  assign n69334 = ~n15067 & ~n69333;
  assign n69335 = ~i_hbusreq3 & ~n69334;
  assign n69336 = ~n68465 & ~n69335;
  assign n69337 = ~controllable_hgrant3 & ~n69336;
  assign n69338 = ~n15066 & ~n69337;
  assign n69339 = ~i_hbusreq9 & ~n69338;
  assign n69340 = ~n68464 & ~n69339;
  assign n69341 = ~i_hbusreq4 & ~n69340;
  assign n69342 = ~n68463 & ~n69341;
  assign n69343 = ~controllable_hgrant4 & ~n69342;
  assign n69344 = ~n15065 & ~n69343;
  assign n69345 = ~i_hbusreq5 & ~n69344;
  assign n69346 = ~n68462 & ~n69345;
  assign n69347 = ~controllable_hgrant5 & ~n69346;
  assign n69348 = ~n15064 & ~n69347;
  assign n69349 = ~controllable_hmaster2 & ~n69348;
  assign n69350 = ~n67557 & ~n69349;
  assign n69351 = controllable_hmaster1 & ~n69350;
  assign n69352 = ~n67709 & ~n69351;
  assign n69353 = i_hlock6 & ~n69352;
  assign n69354 = ~n67712 & ~n69349;
  assign n69355 = controllable_hmaster1 & ~n69354;
  assign n69356 = ~n67709 & ~n69355;
  assign n69357 = ~i_hlock6 & ~n69356;
  assign n69358 = ~n69353 & ~n69357;
  assign n69359 = ~i_hbusreq6 & ~n69358;
  assign n69360 = ~n69329 & ~n69359;
  assign n69361 = ~controllable_hgrant6 & ~n69360;
  assign n69362 = ~n15582 & ~n69361;
  assign n69363 = ~controllable_hmaster0 & ~n69362;
  assign n69364 = ~n67625 & ~n69363;
  assign n69365 = ~i_hbusreq8 & ~n69364;
  assign n69366 = ~n69328 & ~n69365;
  assign n69367 = ~controllable_hmaster3 & ~n69366;
  assign n69368 = ~n67930 & ~n69367;
  assign n69369 = i_hlock7 & ~n69368;
  assign n69370 = i_hbusreq8 & ~n69322;
  assign n69371 = ~n67738 & ~n69363;
  assign n69372 = ~i_hbusreq8 & ~n69371;
  assign n69373 = ~n69370 & ~n69372;
  assign n69374 = ~controllable_hmaster3 & ~n69373;
  assign n69375 = ~n67930 & ~n69374;
  assign n69376 = ~i_hlock7 & ~n69375;
  assign n69377 = ~n69369 & ~n69376;
  assign n69378 = ~i_hbusreq7 & ~n69377;
  assign n69379 = ~n69327 & ~n69378;
  assign n69380 = n7924 & ~n69379;
  assign n69381 = ~n69035 & ~n69380;
  assign n69382 = n8214 & ~n69381;
  assign n69383 = ~n69305 & ~n69382;
  assign n69384 = n8202 & ~n69383;
  assign n69385 = ~n69227 & ~n69384;
  assign n69386 = n7920 & ~n69385;
  assign n69387 = ~n66580 & ~n69386;
  assign n69388 = n7728 & ~n69387;
  assign n69389 = ~n68574 & ~n69388;
  assign n69390 = ~n7723 & ~n69389;
  assign n69391 = ~n69096 & ~n69390;
  assign n69392 = ~n7714 & ~n69391;
  assign n69393 = ~n69095 & ~n69392;
  assign n69394 = ~n7705 & ~n69393;
  assign n69395 = ~n22399 & ~n69394;
  assign n69396 = n7808 & ~n69395;
  assign n69397 = ~n68594 & ~n69396;
  assign n69398 = ~n8195 & ~n69397;
  assign n69399 = controllable_hgrant6 & ~n10323;
  assign n69400 = ~controllable_hmaster2 & ~n66529;
  assign n69401 = ~controllable_hmaster1 & ~n69400;
  assign n69402 = ~controllable_hmaster1 & ~n69401;
  assign n69403 = ~controllable_hgrant6 & ~n69402;
  assign n69404 = ~n69399 & ~n69403;
  assign n69405 = ~controllable_hmaster0 & ~n69404;
  assign n69406 = ~controllable_hmaster0 & ~n69405;
  assign n69407 = ~controllable_hmaster3 & ~n69406;
  assign n69408 = ~controllable_hmaster3 & ~n69407;
  assign n69409 = n7924 & ~n69408;
  assign n69410 = n7924 & ~n69409;
  assign n69411 = n8214 & ~n69410;
  assign n69412 = ~n10320 & ~n69411;
  assign n69413 = ~n8202 & ~n69412;
  assign n69414 = controllable_hgrant6 & ~n10444;
  assign n69415 = controllable_hgrant5 & ~n10424;
  assign n69416 = controllable_hgrant4 & ~n10424;
  assign n69417 = controllable_hgrant3 & ~n10424;
  assign n69418 = controllable_hgrant1 & ~n10424;
  assign n69419 = n7928 & ~n66519;
  assign n69420 = ~controllable_hgrant1 & ~n69419;
  assign n69421 = ~n69418 & ~n69420;
  assign n69422 = ~controllable_hgrant3 & ~n69421;
  assign n69423 = ~n69417 & ~n69422;
  assign n69424 = ~controllable_hgrant4 & ~n69423;
  assign n69425 = ~n69416 & ~n69424;
  assign n69426 = ~controllable_hgrant5 & ~n69425;
  assign n69427 = ~n69415 & ~n69426;
  assign n69428 = ~controllable_hmaster2 & ~n69427;
  assign n69429 = ~n10423 & ~n69428;
  assign n69430 = ~controllable_hmaster1 & ~n69429;
  assign n69431 = ~n10415 & ~n69430;
  assign n69432 = n8217 & ~n69431;
  assign n69433 = ~n10432 & ~n69430;
  assign n69434 = ~n8217 & ~n69433;
  assign n69435 = ~n69432 & ~n69434;
  assign n69436 = i_hlock6 & ~n69435;
  assign n69437 = ~n10439 & ~n69430;
  assign n69438 = ~n8217 & ~n69437;
  assign n69439 = ~n69432 & ~n69438;
  assign n69440 = ~i_hlock6 & ~n69439;
  assign n69441 = ~n69436 & ~n69440;
  assign n69442 = ~controllable_hgrant6 & ~n69441;
  assign n69443 = ~n69414 & ~n69442;
  assign n69444 = ~controllable_hmaster0 & ~n69443;
  assign n69445 = ~n10411 & ~n69444;
  assign n69446 = ~controllable_hmaster3 & ~n69445;
  assign n69447 = ~n10379 & ~n69446;
  assign n69448 = i_hbusreq7 & ~n69447;
  assign n69449 = i_hbusreq8 & ~n69445;
  assign n69450 = controllable_hgrant6 & ~n10616;
  assign n69451 = i_hbusreq6 & ~n69441;
  assign n69452 = ~n10589 & ~n69428;
  assign n69453 = ~controllable_hmaster1 & ~n69452;
  assign n69454 = ~n10569 & ~n69453;
  assign n69455 = n8217 & ~n69454;
  assign n69456 = ~n10599 & ~n69453;
  assign n69457 = ~n8217 & ~n69456;
  assign n69458 = ~n69455 & ~n69457;
  assign n69459 = i_hlock6 & ~n69458;
  assign n69460 = ~n10609 & ~n69453;
  assign n69461 = ~n8217 & ~n69460;
  assign n69462 = ~n69455 & ~n69461;
  assign n69463 = ~i_hlock6 & ~n69462;
  assign n69464 = ~n69459 & ~n69463;
  assign n69465 = ~i_hbusreq6 & ~n69464;
  assign n69466 = ~n69451 & ~n69465;
  assign n69467 = ~controllable_hgrant6 & ~n69466;
  assign n69468 = ~n69450 & ~n69467;
  assign n69469 = ~controllable_hmaster0 & ~n69468;
  assign n69470 = ~n10549 & ~n69469;
  assign n69471 = ~i_hbusreq8 & ~n69470;
  assign n69472 = ~n69449 & ~n69471;
  assign n69473 = ~controllable_hmaster3 & ~n69472;
  assign n69474 = ~n10459 & ~n69473;
  assign n69475 = ~i_hbusreq7 & ~n69474;
  assign n69476 = ~n69448 & ~n69475;
  assign n69477 = n7924 & ~n69476;
  assign n69478 = ~n10375 & ~n69477;
  assign n69479 = n8214 & ~n69478;
  assign n69480 = n8214 & ~n69479;
  assign n69481 = n8202 & ~n69480;
  assign n69482 = ~n69413 & ~n69481;
  assign n69483 = n7728 & ~n69482;
  assign n69484 = ~n7743 & ~n69407;
  assign n69485 = i_hbusreq7 & ~n69484;
  assign n69486 = ~n7779 & ~n69407;
  assign n69487 = ~i_hbusreq7 & ~n69486;
  assign n69488 = ~n69485 & ~n69487;
  assign n69489 = n7924 & ~n69488;
  assign n69490 = ~n8337 & ~n69489;
  assign n69491 = n8214 & ~n69490;
  assign n69492 = ~n10639 & ~n69491;
  assign n69493 = ~n8202 & ~n69492;
  assign n69494 = n8214 & ~n66579;
  assign n69495 = ~n8336 & ~n69494;
  assign n69496 = n8202 & ~n69495;
  assign n69497 = ~n69493 & ~n69496;
  assign n69498 = ~n7728 & ~n69497;
  assign n69499 = ~n69483 & ~n69498;
  assign n69500 = ~n7723 & ~n69499;
  assign n69501 = ~n7723 & ~n69500;
  assign n69502 = ~n7714 & ~n69501;
  assign n69503 = ~n7714 & ~n69502;
  assign n69504 = n7705 & ~n69503;
  assign n69505 = n7723 & ~n69497;
  assign n69506 = n7920 & ~n69497;
  assign n69507 = ~n66580 & ~n69506;
  assign n69508 = ~n7723 & ~n69507;
  assign n69509 = ~n69505 & ~n69508;
  assign n69510 = n7714 & ~n69509;
  assign n69511 = ~n66585 & ~n69510;
  assign n69512 = ~n7705 & ~n69511;
  assign n69513 = ~n69504 & ~n69512;
  assign n69514 = ~n7808 & ~n69513;
  assign n69515 = ~n7920 & ~n69482;
  assign n69516 = ~controllable_hmaster2 & ~n68043;
  assign n69517 = ~controllable_hmaster1 & ~n69516;
  assign n69518 = ~controllable_hmaster1 & ~n69517;
  assign n69519 = ~controllable_hgrant6 & ~n69518;
  assign n69520 = ~n23787 & ~n69519;
  assign n69521 = ~controllable_hmaster0 & ~n69520;
  assign n69522 = ~controllable_hmaster0 & ~n69521;
  assign n69523 = ~controllable_hmaster3 & ~n69522;
  assign n69524 = ~controllable_hmaster3 & ~n69523;
  assign n69525 = i_hbusreq7 & ~n69524;
  assign n69526 = i_hbusreq8 & ~n69522;
  assign n69527 = i_hbusreq6 & ~n69518;
  assign n69528 = ~controllable_hmaster2 & ~n68093;
  assign n69529 = ~controllable_hmaster1 & ~n69528;
  assign n69530 = ~controllable_hmaster1 & ~n69529;
  assign n69531 = ~i_hbusreq6 & ~n69530;
  assign n69532 = ~n69527 & ~n69531;
  assign n69533 = ~controllable_hgrant6 & ~n69532;
  assign n69534 = ~n23799 & ~n69533;
  assign n69535 = ~controllable_hmaster0 & ~n69534;
  assign n69536 = ~controllable_hmaster0 & ~n69535;
  assign n69537 = ~i_hbusreq8 & ~n69536;
  assign n69538 = ~n69526 & ~n69537;
  assign n69539 = ~controllable_hmaster3 & ~n69538;
  assign n69540 = ~controllable_hmaster3 & ~n69539;
  assign n69541 = ~i_hbusreq7 & ~n69540;
  assign n69542 = ~n69525 & ~n69541;
  assign n69543 = ~n7924 & ~n69542;
  assign n69544 = i_hlock0 & i_hready;
  assign n69545 = ~i_hlock0 & ~n16485;
  assign n69546 = ~n69544 & ~n69545;
  assign n69547 = ~controllable_hgrant2 & n69546;
  assign n69548 = ~controllable_hgrant2 & ~n69547;
  assign n69549 = n7733 & ~n69548;
  assign n69550 = ~n16473 & ~n69549;
  assign n69551 = n7928 & ~n69550;
  assign n69552 = n7928 & ~n69551;
  assign n69553 = ~controllable_hgrant1 & ~n69552;
  assign n69554 = ~controllable_hgrant1 & ~n69553;
  assign n69555 = ~controllable_hgrant3 & ~n69554;
  assign n69556 = ~controllable_hgrant3 & ~n69555;
  assign n69557 = ~controllable_hgrant4 & ~n69556;
  assign n69558 = ~controllable_hgrant4 & ~n69557;
  assign n69559 = ~controllable_hgrant5 & ~n69558;
  assign n69560 = ~controllable_hgrant5 & ~n69559;
  assign n69561 = ~controllable_hgrant6 & ~n69560;
  assign n69562 = ~controllable_hgrant6 & ~n69561;
  assign n69563 = controllable_hmaster3 & ~n69562;
  assign n69564 = controllable_hmaster0 & ~n69562;
  assign n69565 = controllable_hmaster1 & ~n69560;
  assign n69566 = controllable_hmaster2 & ~n69560;
  assign n69567 = ~n68231 & ~n69566;
  assign n69568 = ~controllable_hmaster1 & ~n69567;
  assign n69569 = ~n69565 & ~n69568;
  assign n69570 = ~controllable_hgrant6 & ~n69569;
  assign n69571 = ~n23787 & ~n69570;
  assign n69572 = ~controllable_hmaster0 & ~n69571;
  assign n69573 = ~n69564 & ~n69572;
  assign n69574 = ~controllable_hmaster3 & ~n69573;
  assign n69575 = ~n69563 & ~n69574;
  assign n69576 = i_hbusreq7 & ~n69575;
  assign n69577 = i_hbusreq8 & ~n69562;
  assign n69578 = i_hbusreq6 & ~n69560;
  assign n69579 = i_hbusreq5 & ~n69558;
  assign n69580 = i_hbusreq4 & ~n69556;
  assign n69581 = i_hbusreq9 & ~n69556;
  assign n69582 = i_hbusreq3 & ~n69554;
  assign n69583 = i_hbusreq1 & ~n69552;
  assign n69584 = ~n16571 & ~n69549;
  assign n69585 = n7928 & ~n69584;
  assign n69586 = n7928 & ~n69585;
  assign n69587 = ~i_hbusreq1 & ~n69586;
  assign n69588 = ~n69583 & ~n69587;
  assign n69589 = ~controllable_hgrant1 & ~n69588;
  assign n69590 = ~controllable_hgrant1 & ~n69589;
  assign n69591 = ~i_hbusreq3 & ~n69590;
  assign n69592 = ~n69582 & ~n69591;
  assign n69593 = ~controllable_hgrant3 & ~n69592;
  assign n69594 = ~controllable_hgrant3 & ~n69593;
  assign n69595 = ~i_hbusreq9 & ~n69594;
  assign n69596 = ~n69581 & ~n69595;
  assign n69597 = ~i_hbusreq4 & ~n69596;
  assign n69598 = ~n69580 & ~n69597;
  assign n69599 = ~controllable_hgrant4 & ~n69598;
  assign n69600 = ~controllable_hgrant4 & ~n69599;
  assign n69601 = ~i_hbusreq5 & ~n69600;
  assign n69602 = ~n69579 & ~n69601;
  assign n69603 = ~controllable_hgrant5 & ~n69602;
  assign n69604 = ~controllable_hgrant5 & ~n69603;
  assign n69605 = ~i_hbusreq6 & ~n69604;
  assign n69606 = ~n69578 & ~n69605;
  assign n69607 = ~controllable_hgrant6 & ~n69606;
  assign n69608 = ~controllable_hgrant6 & ~n69607;
  assign n69609 = ~i_hbusreq8 & ~n69608;
  assign n69610 = ~n69577 & ~n69609;
  assign n69611 = controllable_hmaster3 & ~n69610;
  assign n69612 = i_hbusreq8 & ~n69573;
  assign n69613 = controllable_hmaster0 & ~n69608;
  assign n69614 = i_hbusreq6 & ~n69569;
  assign n69615 = controllable_hmaster1 & ~n69604;
  assign n69616 = controllable_hmaster2 & ~n69604;
  assign n69617 = ~n68529 & ~n69616;
  assign n69618 = ~controllable_hmaster1 & ~n69617;
  assign n69619 = ~n69615 & ~n69618;
  assign n69620 = ~i_hbusreq6 & ~n69619;
  assign n69621 = ~n69614 & ~n69620;
  assign n69622 = ~controllable_hgrant6 & ~n69621;
  assign n69623 = ~n23799 & ~n69622;
  assign n69624 = ~controllable_hmaster0 & ~n69623;
  assign n69625 = ~n69613 & ~n69624;
  assign n69626 = ~i_hbusreq8 & ~n69625;
  assign n69627 = ~n69612 & ~n69626;
  assign n69628 = ~controllable_hmaster3 & ~n69627;
  assign n69629 = ~n69611 & ~n69628;
  assign n69630 = ~i_hbusreq7 & ~n69629;
  assign n69631 = ~n69576 & ~n69630;
  assign n69632 = n7924 & ~n69631;
  assign n69633 = ~n69543 & ~n69632;
  assign n69634 = n8214 & ~n69633;
  assign n69635 = ~n23786 & ~n69634;
  assign n69636 = ~n8202 & ~n69635;
  assign n69637 = n7924 & ~n68570;
  assign n69638 = ~n8214 & ~n69637;
  assign n69639 = controllable_hmaster0 & ~n17350;
  assign n69640 = controllable_hmaster1 & ~n17339;
  assign n69641 = controllable_hmaster2 & ~n17339;
  assign n69642 = ~n23842 & ~n69641;
  assign n69643 = ~controllable_hmaster1 & ~n69642;
  assign n69644 = ~n69640 & ~n69643;
  assign n69645 = ~controllable_hgrant6 & ~n69644;
  assign n69646 = ~n13198 & ~n69645;
  assign n69647 = ~controllable_hmaster0 & ~n69646;
  assign n69648 = ~n69639 & ~n69647;
  assign n69649 = ~controllable_hmaster3 & ~n69648;
  assign n69650 = ~n33462 & ~n69649;
  assign n69651 = i_hbusreq7 & ~n69650;
  assign n69652 = i_hbusreq8 & ~n69648;
  assign n69653 = i_hbusreq6 & ~n69644;
  assign n69654 = n7928 & ~n68073;
  assign n69655 = ~i_hbusreq1 & ~n69654;
  assign n69656 = ~n23892 & ~n69655;
  assign n69657 = ~controllable_hgrant1 & ~n69656;
  assign n69658 = ~n15824 & ~n69657;
  assign n69659 = ~i_hbusreq3 & ~n69658;
  assign n69660 = ~n23891 & ~n69659;
  assign n69661 = ~controllable_hgrant3 & ~n69660;
  assign n69662 = ~n15823 & ~n69661;
  assign n69663 = ~i_hbusreq9 & ~n69662;
  assign n69664 = ~n23890 & ~n69663;
  assign n69665 = ~i_hbusreq4 & ~n69664;
  assign n69666 = ~n23889 & ~n69665;
  assign n69667 = ~controllable_hgrant4 & ~n69666;
  assign n69668 = ~n15822 & ~n69667;
  assign n69669 = ~i_hbusreq5 & ~n69668;
  assign n69670 = ~n23888 & ~n69669;
  assign n69671 = ~controllable_hgrant5 & ~n69670;
  assign n69672 = ~n15821 & ~n69671;
  assign n69673 = ~controllable_hmaster2 & ~n69672;
  assign n69674 = ~n23960 & ~n69673;
  assign n69675 = ~controllable_hmaster1 & ~n69674;
  assign n69676 = ~n23959 & ~n69675;
  assign n69677 = ~i_hbusreq6 & ~n69676;
  assign n69678 = ~n69653 & ~n69677;
  assign n69679 = ~controllable_hgrant6 & ~n69678;
  assign n69680 = ~n15818 & ~n69679;
  assign n69681 = ~controllable_hmaster0 & ~n69680;
  assign n69682 = ~n23958 & ~n69681;
  assign n69683 = ~i_hbusreq8 & ~n69682;
  assign n69684 = ~n69652 & ~n69683;
  assign n69685 = ~controllable_hmaster3 & ~n69684;
  assign n69686 = ~n33477 & ~n69685;
  assign n69687 = ~i_hbusreq7 & ~n69686;
  assign n69688 = ~n69651 & ~n69687;
  assign n69689 = ~n7924 & ~n69688;
  assign n69690 = n7928 & ~n68124;
  assign n69691 = ~controllable_hgrant1 & ~n69690;
  assign n69692 = ~n13179 & ~n69691;
  assign n69693 = ~controllable_hgrant3 & ~n69692;
  assign n69694 = ~n13178 & ~n69693;
  assign n69695 = ~controllable_hgrant4 & ~n69694;
  assign n69696 = ~n13177 & ~n69695;
  assign n69697 = ~controllable_hgrant5 & ~n69696;
  assign n69698 = ~n13176 & ~n69697;
  assign n69699 = controllable_hmaster1 & ~n69698;
  assign n69700 = controllable_hmaster2 & ~n69698;
  assign n69701 = n7928 & ~n67208;
  assign n69702 = ~controllable_hgrant1 & ~n69701;
  assign n69703 = ~n13179 & ~n69702;
  assign n69704 = ~controllable_hgrant3 & ~n69703;
  assign n69705 = ~n13178 & ~n69704;
  assign n69706 = ~controllable_hgrant4 & ~n69705;
  assign n69707 = ~n13177 & ~n69706;
  assign n69708 = ~controllable_hgrant5 & ~n69707;
  assign n69709 = ~n13176 & ~n69708;
  assign n69710 = ~controllable_hmaster2 & ~n69709;
  assign n69711 = ~n69700 & ~n69710;
  assign n69712 = ~controllable_hmaster1 & ~n69711;
  assign n69713 = ~n69699 & ~n69712;
  assign n69714 = ~controllable_hgrant6 & ~n69713;
  assign n69715 = ~n13198 & ~n69714;
  assign n69716 = controllable_hmaster3 & ~n69715;
  assign n69717 = ~controllable_hgrant6 & ~n69709;
  assign n69718 = ~n13198 & ~n69717;
  assign n69719 = controllable_hmaster0 & ~n69718;
  assign n69720 = controllable_hmaster1 & ~n69709;
  assign n69721 = controllable_hmaster2 & ~n69709;
  assign n69722 = n7928 & ~n68221;
  assign n69723 = ~controllable_hgrant1 & ~n69722;
  assign n69724 = ~n13179 & ~n69723;
  assign n69725 = ~controllable_hgrant3 & ~n69724;
  assign n69726 = ~n13178 & ~n69725;
  assign n69727 = ~controllable_hgrant4 & ~n69726;
  assign n69728 = ~n13177 & ~n69727;
  assign n69729 = ~controllable_hgrant5 & ~n69728;
  assign n69730 = ~n13176 & ~n69729;
  assign n69731 = ~controllable_hmaster2 & ~n69730;
  assign n69732 = ~n69721 & ~n69731;
  assign n69733 = ~controllable_hmaster1 & ~n69732;
  assign n69734 = ~n69720 & ~n69733;
  assign n69735 = ~controllable_hgrant6 & ~n69734;
  assign n69736 = ~n13198 & ~n69735;
  assign n69737 = ~controllable_hmaster0 & ~n69736;
  assign n69738 = ~n69719 & ~n69737;
  assign n69739 = ~controllable_hmaster3 & ~n69738;
  assign n69740 = ~n69716 & ~n69739;
  assign n69741 = i_hbusreq7 & ~n69740;
  assign n69742 = i_hbusreq8 & ~n69715;
  assign n69743 = i_hbusreq6 & ~n69713;
  assign n69744 = i_hbusreq5 & ~n69696;
  assign n69745 = i_hbusreq4 & ~n69694;
  assign n69746 = i_hbusreq9 & ~n69694;
  assign n69747 = i_hbusreq3 & ~n69692;
  assign n69748 = i_hbusreq1 & ~n69690;
  assign n69749 = n7928 & ~n68278;
  assign n69750 = ~i_hbusreq1 & ~n69749;
  assign n69751 = ~n69748 & ~n69750;
  assign n69752 = ~controllable_hgrant1 & ~n69751;
  assign n69753 = ~n15730 & ~n69752;
  assign n69754 = ~i_hbusreq3 & ~n69753;
  assign n69755 = ~n69747 & ~n69754;
  assign n69756 = ~controllable_hgrant3 & ~n69755;
  assign n69757 = ~n15729 & ~n69756;
  assign n69758 = ~i_hbusreq9 & ~n69757;
  assign n69759 = ~n69746 & ~n69758;
  assign n69760 = ~i_hbusreq4 & ~n69759;
  assign n69761 = ~n69745 & ~n69760;
  assign n69762 = ~controllable_hgrant4 & ~n69761;
  assign n69763 = ~n15728 & ~n69762;
  assign n69764 = ~i_hbusreq5 & ~n69763;
  assign n69765 = ~n69744 & ~n69764;
  assign n69766 = ~controllable_hgrant5 & ~n69765;
  assign n69767 = ~n15727 & ~n69766;
  assign n69768 = controllable_hmaster1 & ~n69767;
  assign n69769 = controllable_hmaster2 & ~n69767;
  assign n69770 = i_hbusreq5 & ~n69707;
  assign n69771 = i_hbusreq4 & ~n69705;
  assign n69772 = i_hbusreq9 & ~n69705;
  assign n69773 = i_hbusreq3 & ~n69703;
  assign n69774 = i_hbusreq1 & ~n69701;
  assign n69775 = n7928 & ~n68301;
  assign n69776 = ~i_hbusreq1 & ~n69775;
  assign n69777 = ~n69774 & ~n69776;
  assign n69778 = ~controllable_hgrant1 & ~n69777;
  assign n69779 = ~n15677 & ~n69778;
  assign n69780 = ~i_hbusreq3 & ~n69779;
  assign n69781 = ~n69773 & ~n69780;
  assign n69782 = ~controllable_hgrant3 & ~n69781;
  assign n69783 = ~n15676 & ~n69782;
  assign n69784 = ~i_hbusreq9 & ~n69783;
  assign n69785 = ~n69772 & ~n69784;
  assign n69786 = ~i_hbusreq4 & ~n69785;
  assign n69787 = ~n69771 & ~n69786;
  assign n69788 = ~controllable_hgrant4 & ~n69787;
  assign n69789 = ~n15675 & ~n69788;
  assign n69790 = ~i_hbusreq5 & ~n69789;
  assign n69791 = ~n69770 & ~n69790;
  assign n69792 = ~controllable_hgrant5 & ~n69791;
  assign n69793 = ~n15674 & ~n69792;
  assign n69794 = ~controllable_hmaster2 & ~n69793;
  assign n69795 = ~n69769 & ~n69794;
  assign n69796 = ~controllable_hmaster1 & ~n69795;
  assign n69797 = ~n69768 & ~n69796;
  assign n69798 = ~i_hbusreq6 & ~n69797;
  assign n69799 = ~n69743 & ~n69798;
  assign n69800 = ~controllable_hgrant6 & ~n69799;
  assign n69801 = ~n15672 & ~n69800;
  assign n69802 = ~i_hbusreq8 & ~n69801;
  assign n69803 = ~n69742 & ~n69802;
  assign n69804 = controllable_hmaster3 & ~n69803;
  assign n69805 = i_hbusreq8 & ~n69738;
  assign n69806 = i_hbusreq6 & ~n69709;
  assign n69807 = ~i_hbusreq6 & ~n69793;
  assign n69808 = ~n69806 & ~n69807;
  assign n69809 = ~controllable_hgrant6 & ~n69808;
  assign n69810 = ~n15812 & ~n69809;
  assign n69811 = controllable_hmaster0 & ~n69810;
  assign n69812 = i_hbusreq6 & ~n69734;
  assign n69813 = controllable_hmaster1 & ~n69793;
  assign n69814 = controllable_hmaster2 & ~n69793;
  assign n69815 = i_hbusreq5 & ~n69728;
  assign n69816 = i_hbusreq4 & ~n69726;
  assign n69817 = i_hbusreq9 & ~n69726;
  assign n69818 = i_hbusreq3 & ~n69724;
  assign n69819 = i_hbusreq1 & ~n69722;
  assign n69820 = n7928 & ~n68509;
  assign n69821 = ~i_hbusreq1 & ~n69820;
  assign n69822 = ~n69819 & ~n69821;
  assign n69823 = ~controllable_hgrant1 & ~n69822;
  assign n69824 = ~n15824 & ~n69823;
  assign n69825 = ~i_hbusreq3 & ~n69824;
  assign n69826 = ~n69818 & ~n69825;
  assign n69827 = ~controllable_hgrant3 & ~n69826;
  assign n69828 = ~n15823 & ~n69827;
  assign n69829 = ~i_hbusreq9 & ~n69828;
  assign n69830 = ~n69817 & ~n69829;
  assign n69831 = ~i_hbusreq4 & ~n69830;
  assign n69832 = ~n69816 & ~n69831;
  assign n69833 = ~controllable_hgrant4 & ~n69832;
  assign n69834 = ~n15822 & ~n69833;
  assign n69835 = ~i_hbusreq5 & ~n69834;
  assign n69836 = ~n69815 & ~n69835;
  assign n69837 = ~controllable_hgrant5 & ~n69836;
  assign n69838 = ~n15821 & ~n69837;
  assign n69839 = ~controllable_hmaster2 & ~n69838;
  assign n69840 = ~n69814 & ~n69839;
  assign n69841 = ~controllable_hmaster1 & ~n69840;
  assign n69842 = ~n69813 & ~n69841;
  assign n69843 = ~i_hbusreq6 & ~n69842;
  assign n69844 = ~n69812 & ~n69843;
  assign n69845 = ~controllable_hgrant6 & ~n69844;
  assign n69846 = ~n15818 & ~n69845;
  assign n69847 = ~controllable_hmaster0 & ~n69846;
  assign n69848 = ~n69811 & ~n69847;
  assign n69849 = ~i_hbusreq8 & ~n69848;
  assign n69850 = ~n69805 & ~n69849;
  assign n69851 = ~controllable_hmaster3 & ~n69850;
  assign n69852 = ~n69804 & ~n69851;
  assign n69853 = ~i_hbusreq7 & ~n69852;
  assign n69854 = ~n69741 & ~n69853;
  assign n69855 = n7924 & ~n69854;
  assign n69856 = ~n69689 & ~n69855;
  assign n69857 = n8214 & ~n69856;
  assign n69858 = ~n69638 & ~n69857;
  assign n69859 = n8202 & ~n69858;
  assign n69860 = ~n69636 & ~n69859;
  assign n69861 = n7920 & ~n69860;
  assign n69862 = ~n69515 & ~n69861;
  assign n69863 = n7728 & ~n69862;
  assign n69864 = ~n7920 & ~n69497;
  assign n69865 = ~n24262 & ~n69523;
  assign n69866 = i_hbusreq7 & ~n69865;
  assign n69867 = ~n24262 & ~n69539;
  assign n69868 = ~i_hbusreq7 & ~n69867;
  assign n69869 = ~n69866 & ~n69868;
  assign n69870 = ~n7924 & ~n69869;
  assign n69871 = ~n17092 & ~n69549;
  assign n69872 = n7928 & ~n69871;
  assign n69873 = ~n17088 & ~n69872;
  assign n69874 = ~controllable_hgrant1 & ~n69873;
  assign n69875 = ~n7813 & ~n69874;
  assign n69876 = ~controllable_hgrant3 & ~n69875;
  assign n69877 = ~n7812 & ~n69876;
  assign n69878 = ~controllable_hgrant4 & ~n69877;
  assign n69879 = ~n7811 & ~n69878;
  assign n69880 = ~controllable_hgrant5 & ~n69879;
  assign n69881 = ~n7810 & ~n69880;
  assign n69882 = controllable_hmaster1 & ~n69881;
  assign n69883 = controllable_hmaster2 & ~n69881;
  assign n69884 = ~controllable_hmaster2 & ~n69560;
  assign n69885 = ~n69883 & ~n69884;
  assign n69886 = ~controllable_hmaster1 & ~n69885;
  assign n69887 = ~n69882 & ~n69886;
  assign n69888 = ~controllable_hgrant6 & ~n69887;
  assign n69889 = ~n7809 & ~n69888;
  assign n69890 = controllable_hmaster3 & ~n69889;
  assign n69891 = ~n69574 & ~n69890;
  assign n69892 = i_hbusreq7 & ~n69891;
  assign n69893 = i_hbusreq8 & ~n69889;
  assign n69894 = i_hbusreq6 & ~n69887;
  assign n69895 = i_hbusreq5 & ~n69879;
  assign n69896 = i_hbusreq4 & ~n69877;
  assign n69897 = i_hbusreq9 & ~n69877;
  assign n69898 = i_hbusreq3 & ~n69875;
  assign n69899 = i_hbusreq1 & ~n69873;
  assign n69900 = ~n21845 & ~n69549;
  assign n69901 = n7928 & ~n69900;
  assign n69902 = ~n17088 & ~n69901;
  assign n69903 = ~i_hbusreq1 & ~n69902;
  assign n69904 = ~n69899 & ~n69903;
  assign n69905 = ~controllable_hgrant1 & ~n69904;
  assign n69906 = ~n7813 & ~n69905;
  assign n69907 = ~i_hbusreq3 & ~n69906;
  assign n69908 = ~n69898 & ~n69907;
  assign n69909 = ~controllable_hgrant3 & ~n69908;
  assign n69910 = ~n7812 & ~n69909;
  assign n69911 = ~i_hbusreq9 & ~n69910;
  assign n69912 = ~n69897 & ~n69911;
  assign n69913 = ~i_hbusreq4 & ~n69912;
  assign n69914 = ~n69896 & ~n69913;
  assign n69915 = ~controllable_hgrant4 & ~n69914;
  assign n69916 = ~n7811 & ~n69915;
  assign n69917 = ~i_hbusreq5 & ~n69916;
  assign n69918 = ~n69895 & ~n69917;
  assign n69919 = ~controllable_hgrant5 & ~n69918;
  assign n69920 = ~n7810 & ~n69919;
  assign n69921 = controllable_hmaster1 & ~n69920;
  assign n69922 = controllable_hmaster2 & ~n69920;
  assign n69923 = ~controllable_hmaster2 & ~n69604;
  assign n69924 = ~n69922 & ~n69923;
  assign n69925 = ~controllable_hmaster1 & ~n69924;
  assign n69926 = ~n69921 & ~n69925;
  assign n69927 = ~i_hbusreq6 & ~n69926;
  assign n69928 = ~n69894 & ~n69927;
  assign n69929 = ~controllable_hgrant6 & ~n69928;
  assign n69930 = ~n7809 & ~n69929;
  assign n69931 = ~i_hbusreq8 & ~n69930;
  assign n69932 = ~n69893 & ~n69931;
  assign n69933 = controllable_hmaster3 & ~n69932;
  assign n69934 = ~n69628 & ~n69933;
  assign n69935 = ~i_hbusreq7 & ~n69934;
  assign n69936 = ~n69892 & ~n69935;
  assign n69937 = n7924 & ~n69936;
  assign n69938 = ~n69870 & ~n69937;
  assign n69939 = n8214 & ~n69938;
  assign n69940 = ~n24253 & ~n69939;
  assign n69941 = ~n8202 & ~n69940;
  assign n69942 = ~n24264 & ~n68570;
  assign n69943 = ~n8214 & ~n69942;
  assign n69944 = n8214 & ~n68571;
  assign n69945 = ~n69943 & ~n69944;
  assign n69946 = n8202 & ~n69945;
  assign n69947 = ~n69941 & ~n69946;
  assign n69948 = n7920 & ~n69947;
  assign n69949 = ~n69864 & ~n69948;
  assign n69950 = ~n7728 & ~n69949;
  assign n69951 = ~n69863 & ~n69950;
  assign n69952 = ~n7723 & ~n69951;
  assign n69953 = ~n7723 & ~n69952;
  assign n69954 = ~n7714 & ~n69953;
  assign n69955 = ~n7714 & ~n69954;
  assign n69956 = n7705 & ~n69955;
  assign n69957 = ~n24285 & ~n36100;
  assign n69958 = ~controllable_hmaster3 & ~n69957;
  assign n69959 = ~n9093 & ~n69958;
  assign n69960 = i_hbusreq7 & ~n69959;
  assign n69961 = i_hbusreq8 & ~n69957;
  assign n69962 = ~n24299 & ~n66614;
  assign n69963 = ~i_hbusreq8 & ~n69962;
  assign n69964 = ~n69961 & ~n69963;
  assign n69965 = ~controllable_hmaster3 & ~n69964;
  assign n69966 = ~n9117 & ~n69965;
  assign n69967 = ~i_hbusreq7 & ~n69966;
  assign n69968 = ~n69960 & ~n69967;
  assign n69969 = ~n7924 & ~n69968;
  assign n69970 = ~n24325 & ~n36116;
  assign n69971 = ~controllable_hmaster3 & ~n69970;
  assign n69972 = ~n27088 & ~n69971;
  assign n69973 = i_hbusreq7 & ~n69972;
  assign n69974 = i_hbusreq8 & ~n69970;
  assign n69975 = ~n24366 & ~n66633;
  assign n69976 = ~i_hbusreq8 & ~n69975;
  assign n69977 = ~n69974 & ~n69976;
  assign n69978 = ~controllable_hmaster3 & ~n69977;
  assign n69979 = ~n27174 & ~n69978;
  assign n69980 = ~i_hbusreq7 & ~n69979;
  assign n69981 = ~n69973 & ~n69980;
  assign n69982 = n7924 & ~n69981;
  assign n69983 = ~n69969 & ~n69982;
  assign n69984 = ~n8214 & ~n69983;
  assign n69985 = ~n68043 & ~n69641;
  assign n69986 = ~controllable_hmaster1 & ~n69985;
  assign n69987 = ~n69640 & ~n69986;
  assign n69988 = ~controllable_hgrant6 & ~n69987;
  assign n69989 = ~n15964 & ~n69988;
  assign n69990 = ~controllable_hmaster0 & ~n69989;
  assign n69991 = ~n69639 & ~n69990;
  assign n69992 = ~controllable_hmaster3 & ~n69991;
  assign n69993 = ~n29420 & ~n69992;
  assign n69994 = i_hbusreq7 & ~n69993;
  assign n69995 = ~n21649 & ~n23941;
  assign n69996 = ~controllable_hmaster1 & ~n69995;
  assign n69997 = ~n21648 & ~n69996;
  assign n69998 = ~i_hbusreq6 & ~n69997;
  assign n69999 = ~n17401 & ~n69998;
  assign n70000 = ~controllable_hgrant6 & ~n69999;
  assign n70001 = ~n15946 & ~n70000;
  assign n70002 = ~i_hbusreq8 & ~n70001;
  assign n70003 = ~n29445 & ~n70002;
  assign n70004 = controllable_hmaster3 & ~n70003;
  assign n70005 = i_hbusreq8 & ~n69991;
  assign n70006 = i_hbusreq6 & ~n69987;
  assign n70007 = ~n23960 & ~n68093;
  assign n70008 = ~controllable_hmaster1 & ~n70007;
  assign n70009 = ~n23959 & ~n70008;
  assign n70010 = ~i_hbusreq6 & ~n70009;
  assign n70011 = ~n70006 & ~n70010;
  assign n70012 = ~controllable_hgrant6 & ~n70011;
  assign n70013 = ~n15996 & ~n70012;
  assign n70014 = ~controllable_hmaster0 & ~n70013;
  assign n70015 = ~n23958 & ~n70014;
  assign n70016 = ~i_hbusreq8 & ~n70015;
  assign n70017 = ~n70005 & ~n70016;
  assign n70018 = ~controllable_hmaster3 & ~n70017;
  assign n70019 = ~n70004 & ~n70018;
  assign n70020 = ~i_hbusreq7 & ~n70019;
  assign n70021 = ~n69994 & ~n70020;
  assign n70022 = ~n7924 & ~n70021;
  assign n70023 = ~n68135 & ~n69710;
  assign n70024 = ~controllable_hmaster1 & ~n70023;
  assign n70025 = ~n68134 & ~n70024;
  assign n70026 = ~controllable_hgrant6 & ~n70025;
  assign n70027 = ~n13175 & ~n70026;
  assign n70028 = controllable_hmaster3 & ~n70027;
  assign n70029 = ~n68231 & ~n69721;
  assign n70030 = ~controllable_hmaster1 & ~n70029;
  assign n70031 = ~n69720 & ~n70030;
  assign n70032 = ~controllable_hgrant6 & ~n70031;
  assign n70033 = ~n15964 & ~n70032;
  assign n70034 = ~controllable_hmaster0 & ~n70033;
  assign n70035 = ~n69719 & ~n70034;
  assign n70036 = ~controllable_hmaster3 & ~n70035;
  assign n70037 = ~n70028 & ~n70036;
  assign n70038 = i_hbusreq7 & ~n70037;
  assign n70039 = i_hbusreq8 & ~n70027;
  assign n70040 = i_hbusreq6 & ~n70025;
  assign n70041 = ~n68299 & ~n69794;
  assign n70042 = ~controllable_hmaster1 & ~n70041;
  assign n70043 = ~n68298 & ~n70042;
  assign n70044 = ~i_hbusreq6 & ~n70043;
  assign n70045 = ~n70040 & ~n70044;
  assign n70046 = ~controllable_hgrant6 & ~n70045;
  assign n70047 = ~n15946 & ~n70046;
  assign n70048 = ~i_hbusreq8 & ~n70047;
  assign n70049 = ~n70039 & ~n70048;
  assign n70050 = controllable_hmaster3 & ~n70049;
  assign n70051 = i_hbusreq8 & ~n70035;
  assign n70052 = i_hbusreq6 & ~n70031;
  assign n70053 = ~n68529 & ~n69814;
  assign n70054 = ~controllable_hmaster1 & ~n70053;
  assign n70055 = ~n69813 & ~n70054;
  assign n70056 = ~i_hbusreq6 & ~n70055;
  assign n70057 = ~n70052 & ~n70056;
  assign n70058 = ~controllable_hgrant6 & ~n70057;
  assign n70059 = ~n15996 & ~n70058;
  assign n70060 = ~controllable_hmaster0 & ~n70059;
  assign n70061 = ~n69811 & ~n70060;
  assign n70062 = ~i_hbusreq8 & ~n70061;
  assign n70063 = ~n70051 & ~n70062;
  assign n70064 = ~controllable_hmaster3 & ~n70063;
  assign n70065 = ~n70050 & ~n70064;
  assign n70066 = ~i_hbusreq7 & ~n70065;
  assign n70067 = ~n70038 & ~n70066;
  assign n70068 = n7924 & ~n70067;
  assign n70069 = ~n70022 & ~n70068;
  assign n70070 = n8214 & ~n70069;
  assign n70071 = ~n69984 & ~n70070;
  assign n70072 = ~n8202 & ~n70071;
  assign n70073 = n8202 & ~n68571;
  assign n70074 = ~n70072 & ~n70073;
  assign n70075 = n7920 & ~n70074;
  assign n70076 = ~n69864 & ~n70075;
  assign n70077 = n7728 & ~n70076;
  assign n70078 = ~n24493 & ~n66809;
  assign n70079 = ~controllable_hmaster3 & ~n70078;
  assign n70080 = ~n30877 & ~n70079;
  assign n70081 = i_hlock7 & ~n70080;
  assign n70082 = ~n24501 & ~n66809;
  assign n70083 = ~controllable_hmaster3 & ~n70082;
  assign n70084 = ~n30877 & ~n70083;
  assign n70085 = ~i_hlock7 & ~n70084;
  assign n70086 = ~n70081 & ~n70085;
  assign n70087 = i_hbusreq7 & ~n70086;
  assign n70088 = i_hbusreq8 & ~n70078;
  assign n70089 = ~n24517 & ~n66870;
  assign n70090 = ~i_hbusreq8 & ~n70089;
  assign n70091 = ~n70088 & ~n70090;
  assign n70092 = ~controllable_hmaster3 & ~n70091;
  assign n70093 = ~n30896 & ~n70092;
  assign n70094 = i_hlock7 & ~n70093;
  assign n70095 = i_hbusreq8 & ~n70082;
  assign n70096 = ~n24531 & ~n66870;
  assign n70097 = ~i_hbusreq8 & ~n70096;
  assign n70098 = ~n70095 & ~n70097;
  assign n70099 = ~controllable_hmaster3 & ~n70098;
  assign n70100 = ~n30896 & ~n70099;
  assign n70101 = ~i_hlock7 & ~n70100;
  assign n70102 = ~n70094 & ~n70101;
  assign n70103 = ~i_hbusreq7 & ~n70102;
  assign n70104 = ~n70087 & ~n70103;
  assign n70105 = ~n7924 & ~n70104;
  assign n70106 = ~n24559 & ~n66907;
  assign n70107 = ~controllable_hmaster3 & ~n70106;
  assign n70108 = ~n30920 & ~n70107;
  assign n70109 = i_hlock7 & ~n70108;
  assign n70110 = ~n24567 & ~n66907;
  assign n70111 = ~controllable_hmaster3 & ~n70110;
  assign n70112 = ~n30920 & ~n70111;
  assign n70113 = ~i_hlock7 & ~n70112;
  assign n70114 = ~n70109 & ~n70113;
  assign n70115 = i_hbusreq7 & ~n70114;
  assign n70116 = i_hbusreq8 & ~n70106;
  assign n70117 = ~n24610 & ~n66966;
  assign n70118 = ~i_hbusreq8 & ~n70117;
  assign n70119 = ~n70116 & ~n70118;
  assign n70120 = ~controllable_hmaster3 & ~n70119;
  assign n70121 = ~n30939 & ~n70120;
  assign n70122 = i_hlock7 & ~n70121;
  assign n70123 = i_hbusreq8 & ~n70110;
  assign n70124 = ~n24624 & ~n66966;
  assign n70125 = ~i_hbusreq8 & ~n70124;
  assign n70126 = ~n70123 & ~n70125;
  assign n70127 = ~controllable_hmaster3 & ~n70126;
  assign n70128 = ~n30939 & ~n70127;
  assign n70129 = ~i_hlock7 & ~n70128;
  assign n70130 = ~n70122 & ~n70129;
  assign n70131 = ~i_hbusreq7 & ~n70130;
  assign n70132 = ~n70115 & ~n70131;
  assign n70133 = n7924 & ~n70132;
  assign n70134 = ~n70105 & ~n70133;
  assign n70135 = ~n8214 & ~n70134;
  assign n70136 = ~n69944 & ~n70135;
  assign n70137 = ~n8202 & ~n70136;
  assign n70138 = ~n70073 & ~n70137;
  assign n70139 = n7920 & ~n70138;
  assign n70140 = ~n69864 & ~n70139;
  assign n70141 = ~n7728 & ~n70140;
  assign n70142 = ~n70077 & ~n70141;
  assign n70143 = n7723 & ~n70142;
  assign n70144 = ~n7723 & ~n70140;
  assign n70145 = ~n70143 & ~n70144;
  assign n70146 = n7714 & ~n70145;
  assign n70147 = n7723 & ~n70140;
  assign n70148 = ~n67289 & ~n68189;
  assign n70149 = ~controllable_hmaster1 & ~n70148;
  assign n70150 = ~n67283 & ~n70149;
  assign n70151 = ~controllable_hgrant6 & ~n70150;
  assign n70152 = ~n13849 & ~n70151;
  assign n70153 = controllable_hmaster0 & ~n70152;
  assign n70154 = ~n67357 & ~n70153;
  assign n70155 = ~controllable_hmaster3 & ~n70154;
  assign n70156 = ~n67897 & ~n70155;
  assign n70157 = i_hlock7 & ~n70156;
  assign n70158 = ~n67363 & ~n70149;
  assign n70159 = ~controllable_hgrant6 & ~n70158;
  assign n70160 = ~n13951 & ~n70159;
  assign n70161 = controllable_hmaster0 & ~n70160;
  assign n70162 = ~n67357 & ~n70161;
  assign n70163 = ~controllable_hmaster3 & ~n70162;
  assign n70164 = ~n67897 & ~n70163;
  assign n70165 = ~i_hlock7 & ~n70164;
  assign n70166 = ~n70157 & ~n70165;
  assign n70167 = i_hbusreq7 & ~n70166;
  assign n70168 = i_hbusreq8 & ~n70154;
  assign n70169 = i_hbusreq6 & ~n70150;
  assign n70170 = i_hlock1 & ~n67437;
  assign n70171 = ~i_hlock1 & ~n67449;
  assign n70172 = ~n70170 & ~n70171;
  assign n70173 = ~i_hbusreq1 & ~n70172;
  assign n70174 = ~n68430 & ~n70173;
  assign n70175 = ~controllable_hgrant1 & ~n70174;
  assign n70176 = ~n15032 & ~n70175;
  assign n70177 = ~i_hbusreq3 & ~n70176;
  assign n70178 = ~n68429 & ~n70177;
  assign n70179 = ~controllable_hgrant3 & ~n70178;
  assign n70180 = ~n15031 & ~n70179;
  assign n70181 = ~i_hbusreq9 & ~n70180;
  assign n70182 = ~n68428 & ~n70181;
  assign n70183 = ~i_hbusreq4 & ~n70182;
  assign n70184 = ~n68427 & ~n70183;
  assign n70185 = ~controllable_hgrant4 & ~n70184;
  assign n70186 = ~n15030 & ~n70185;
  assign n70187 = ~i_hbusreq5 & ~n70186;
  assign n70188 = ~n68426 & ~n70187;
  assign n70189 = ~controllable_hgrant5 & ~n70188;
  assign n70190 = ~n15029 & ~n70189;
  assign n70191 = ~controllable_hmaster2 & ~n70190;
  assign n70192 = ~n67590 & ~n70191;
  assign n70193 = ~controllable_hmaster1 & ~n70192;
  assign n70194 = ~n67581 & ~n70193;
  assign n70195 = ~i_hbusreq6 & ~n70194;
  assign n70196 = ~n70169 & ~n70195;
  assign n70197 = ~controllable_hgrant6 & ~n70196;
  assign n70198 = ~n16031 & ~n70197;
  assign n70199 = controllable_hmaster0 & ~n70198;
  assign n70200 = ~n67722 & ~n70199;
  assign n70201 = ~i_hbusreq8 & ~n70200;
  assign n70202 = ~n70168 & ~n70201;
  assign n70203 = ~controllable_hmaster3 & ~n70202;
  assign n70204 = ~n67930 & ~n70203;
  assign n70205 = i_hlock7 & ~n70204;
  assign n70206 = i_hbusreq8 & ~n70162;
  assign n70207 = i_hbusreq6 & ~n70158;
  assign n70208 = ~n67732 & ~n70193;
  assign n70209 = ~i_hbusreq6 & ~n70208;
  assign n70210 = ~n70207 & ~n70209;
  assign n70211 = ~controllable_hgrant6 & ~n70210;
  assign n70212 = ~n16068 & ~n70211;
  assign n70213 = controllable_hmaster0 & ~n70212;
  assign n70214 = ~n67722 & ~n70213;
  assign n70215 = ~i_hbusreq8 & ~n70214;
  assign n70216 = ~n70206 & ~n70215;
  assign n70217 = ~controllable_hmaster3 & ~n70216;
  assign n70218 = ~n67930 & ~n70217;
  assign n70219 = ~i_hlock7 & ~n70218;
  assign n70220 = ~n70205 & ~n70219;
  assign n70221 = ~i_hbusreq7 & ~n70220;
  assign n70222 = ~n70167 & ~n70221;
  assign n70223 = n7924 & ~n70222;
  assign n70224 = ~n70105 & ~n70223;
  assign n70225 = ~n8214 & ~n70224;
  assign n70226 = ~n69944 & ~n70225;
  assign n70227 = ~n8202 & ~n70226;
  assign n70228 = ~n70073 & ~n70227;
  assign n70229 = n7920 & ~n70228;
  assign n70230 = ~n66580 & ~n70229;
  assign n70231 = n7728 & ~n70230;
  assign n70232 = ~n68574 & ~n70231;
  assign n70233 = ~n7723 & ~n70232;
  assign n70234 = ~n70147 & ~n70233;
  assign n70235 = ~n7714 & ~n70234;
  assign n70236 = ~n70146 & ~n70235;
  assign n70237 = ~n7705 & ~n70236;
  assign n70238 = ~n69956 & ~n70237;
  assign n70239 = n7808 & ~n70238;
  assign n70240 = ~n69514 & ~n70239;
  assign n70241 = n8195 & ~n70240;
  assign n70242 = ~n69398 & ~n70241;
  assign n70243 = n8193 & ~n70242;
  assign n70244 = ~n68586 & ~n70243;
  assign n70245 = n8191 & ~n70244;
  assign n70246 = ~n11036 & ~n66547;
  assign n70247 = i_hbusreq7 & ~n70246;
  assign n70248 = ~n11051 & ~n66574;
  assign n70249 = ~i_hbusreq7 & ~n70248;
  assign n70250 = ~n70247 & ~n70249;
  assign n70251 = n7924 & ~n70250;
  assign n70252 = ~n8337 & ~n70251;
  assign n70253 = ~n7920 & ~n70252;
  assign n70254 = ~n11058 & ~n70253;
  assign n70255 = ~n7723 & ~n70254;
  assign n70256 = ~n11029 & ~n70255;
  assign n70257 = n7714 & ~n70256;
  assign n70258 = ~n7714 & ~n70252;
  assign n70259 = ~n70257 & ~n70258;
  assign n70260 = ~n7705 & ~n70259;
  assign n70261 = ~n11028 & ~n70260;
  assign n70262 = ~n7808 & ~n70261;
  assign n70263 = ~n11068 & ~n66591;
  assign n70264 = n7728 & ~n70263;
  assign n70265 = ~n11071 & ~n66595;
  assign n70266 = ~n7728 & ~n70265;
  assign n70267 = ~n70264 & ~n70266;
  assign n70268 = ~n7723 & ~n70267;
  assign n70269 = ~n7723 & ~n70268;
  assign n70270 = ~n7714 & ~n70269;
  assign n70271 = ~n7714 & ~n70270;
  assign n70272 = n7705 & ~n70271;
  assign n70273 = ~n11071 & ~n66787;
  assign n70274 = n7728 & ~n70273;
  assign n70275 = ~n11071 & ~n67175;
  assign n70276 = ~n7728 & ~n70275;
  assign n70277 = ~n70274 & ~n70276;
  assign n70278 = n7723 & ~n70277;
  assign n70279 = ~n7723 & ~n70275;
  assign n70280 = ~n70278 & ~n70279;
  assign n70281 = n7714 & ~n70280;
  assign n70282 = n7723 & ~n70275;
  assign n70283 = ~n68031 & ~n70253;
  assign n70284 = n7728 & ~n70283;
  assign n70285 = ~n68572 & ~n70253;
  assign n70286 = ~n7728 & ~n70285;
  assign n70287 = ~n70284 & ~n70286;
  assign n70288 = ~n7723 & ~n70287;
  assign n70289 = ~n70282 & ~n70288;
  assign n70290 = ~n7714 & ~n70289;
  assign n70291 = ~n70281 & ~n70290;
  assign n70292 = ~n7705 & ~n70291;
  assign n70293 = ~n70272 & ~n70292;
  assign n70294 = n7808 & ~n70293;
  assign n70295 = ~n70262 & ~n70294;
  assign n70296 = n8195 & ~n70295;
  assign n70297 = ~n8196 & ~n70296;
  assign n70298 = ~n8193 & ~n70297;
  assign n70299 = ~n9900 & ~n70253;
  assign n70300 = ~n7723 & ~n70299;
  assign n70301 = ~n9899 & ~n70300;
  assign n70302 = n7714 & ~n70301;
  assign n70303 = ~n70258 & ~n70302;
  assign n70304 = ~n7705 & ~n70303;
  assign n70305 = ~n9898 & ~n70304;
  assign n70306 = ~n7808 & ~n70305;
  assign n70307 = ~n69386 & ~n70253;
  assign n70308 = n7728 & ~n70307;
  assign n70309 = ~n70286 & ~n70308;
  assign n70310 = ~n7723 & ~n70309;
  assign n70311 = ~n69096 & ~n70310;
  assign n70312 = ~n7714 & ~n70311;
  assign n70313 = ~n69095 & ~n70312;
  assign n70314 = ~n7705 & ~n70313;
  assign n70315 = ~n22399 & ~n70314;
  assign n70316 = n7808 & ~n70315;
  assign n70317 = ~n70306 & ~n70316;
  assign n70318 = ~n8195 & ~n70317;
  assign n70319 = ~n11136 & ~n69446;
  assign n70320 = i_hbusreq7 & ~n70319;
  assign n70321 = ~n11164 & ~n69473;
  assign n70322 = ~i_hbusreq7 & ~n70321;
  assign n70323 = ~n70320 & ~n70322;
  assign n70324 = n7924 & ~n70323;
  assign n70325 = ~n10375 & ~n70324;
  assign n70326 = n8214 & ~n70325;
  assign n70327 = n8214 & ~n70326;
  assign n70328 = n8202 & ~n70327;
  assign n70329 = ~n69413 & ~n70328;
  assign n70330 = n7728 & ~n70329;
  assign n70331 = n8214 & ~n70252;
  assign n70332 = ~n8336 & ~n70331;
  assign n70333 = n8202 & ~n70332;
  assign n70334 = ~n69493 & ~n70333;
  assign n70335 = ~n7728 & ~n70334;
  assign n70336 = ~n70330 & ~n70335;
  assign n70337 = ~n7723 & ~n70336;
  assign n70338 = ~n7723 & ~n70337;
  assign n70339 = ~n7714 & ~n70338;
  assign n70340 = ~n7714 & ~n70339;
  assign n70341 = n7705 & ~n70340;
  assign n70342 = n7723 & ~n70334;
  assign n70343 = n7920 & ~n70334;
  assign n70344 = ~n70253 & ~n70343;
  assign n70345 = ~n7723 & ~n70344;
  assign n70346 = ~n70342 & ~n70345;
  assign n70347 = n7714 & ~n70346;
  assign n70348 = ~n70258 & ~n70347;
  assign n70349 = ~n7705 & ~n70348;
  assign n70350 = ~n70341 & ~n70349;
  assign n70351 = ~n7808 & ~n70350;
  assign n70352 = ~n7920 & ~n70329;
  assign n70353 = ~n69861 & ~n70352;
  assign n70354 = n7728 & ~n70353;
  assign n70355 = ~n7920 & ~n70334;
  assign n70356 = ~n69948 & ~n70355;
  assign n70357 = ~n7728 & ~n70356;
  assign n70358 = ~n70354 & ~n70357;
  assign n70359 = ~n7723 & ~n70358;
  assign n70360 = ~n7723 & ~n70359;
  assign n70361 = ~n7714 & ~n70360;
  assign n70362 = ~n7714 & ~n70361;
  assign n70363 = n7705 & ~n70362;
  assign n70364 = ~n70075 & ~n70355;
  assign n70365 = n7728 & ~n70364;
  assign n70366 = ~n70139 & ~n70355;
  assign n70367 = ~n7728 & ~n70366;
  assign n70368 = ~n70365 & ~n70367;
  assign n70369 = n7723 & ~n70368;
  assign n70370 = ~n7723 & ~n70366;
  assign n70371 = ~n70369 & ~n70370;
  assign n70372 = n7714 & ~n70371;
  assign n70373 = n7723 & ~n70366;
  assign n70374 = ~n70229 & ~n70253;
  assign n70375 = n7728 & ~n70374;
  assign n70376 = ~n70286 & ~n70375;
  assign n70377 = ~n7723 & ~n70376;
  assign n70378 = ~n70373 & ~n70377;
  assign n70379 = ~n7714 & ~n70378;
  assign n70380 = ~n70372 & ~n70379;
  assign n70381 = ~n7705 & ~n70380;
  assign n70382 = ~n70363 & ~n70381;
  assign n70383 = n7808 & ~n70382;
  assign n70384 = ~n70351 & ~n70383;
  assign n70385 = n8195 & ~n70384;
  assign n70386 = ~n70318 & ~n70385;
  assign n70387 = n8193 & ~n70386;
  assign n70388 = ~n70298 & ~n70387;
  assign n70389 = ~n8191 & ~n70388;
  assign n70390 = ~n70245 & ~n70389;
  assign n70391 = n8188 & ~n70390;
  assign n70392 = ~n11359 & ~n66547;
  assign n70393 = i_hbusreq7 & ~n70392;
  assign n70394 = ~n11385 & ~n66574;
  assign n70395 = ~i_hbusreq7 & ~n70394;
  assign n70396 = ~n70393 & ~n70395;
  assign n70397 = n7924 & ~n70396;
  assign n70398 = ~n8337 & ~n70397;
  assign n70399 = ~n7920 & ~n70398;
  assign n70400 = ~n11392 & ~n70399;
  assign n70401 = ~n7723 & ~n70400;
  assign n70402 = ~n11344 & ~n70401;
  assign n70403 = n7714 & ~n70402;
  assign n70404 = ~n7714 & ~n70398;
  assign n70405 = ~n70403 & ~n70404;
  assign n70406 = ~n7705 & ~n70405;
  assign n70407 = ~n11343 & ~n70406;
  assign n70408 = ~n7808 & ~n70407;
  assign n70409 = ~n11402 & ~n66591;
  assign n70410 = n7728 & ~n70409;
  assign n70411 = ~n11405 & ~n66595;
  assign n70412 = ~n7728 & ~n70411;
  assign n70413 = ~n70410 & ~n70412;
  assign n70414 = ~n7723 & ~n70413;
  assign n70415 = ~n7723 & ~n70414;
  assign n70416 = ~n7714 & ~n70415;
  assign n70417 = ~n7714 & ~n70416;
  assign n70418 = n7705 & ~n70417;
  assign n70419 = ~n11405 & ~n66787;
  assign n70420 = n7728 & ~n70419;
  assign n70421 = ~n11405 & ~n67175;
  assign n70422 = ~n7728 & ~n70421;
  assign n70423 = ~n70420 & ~n70422;
  assign n70424 = n7723 & ~n70423;
  assign n70425 = ~n7723 & ~n70421;
  assign n70426 = ~n70424 & ~n70425;
  assign n70427 = n7714 & ~n70426;
  assign n70428 = n7723 & ~n70421;
  assign n70429 = ~n68031 & ~n70399;
  assign n70430 = n7728 & ~n70429;
  assign n70431 = ~n68572 & ~n70399;
  assign n70432 = ~n7728 & ~n70431;
  assign n70433 = ~n70430 & ~n70432;
  assign n70434 = ~n7723 & ~n70433;
  assign n70435 = ~n70428 & ~n70434;
  assign n70436 = ~n7714 & ~n70435;
  assign n70437 = ~n70427 & ~n70436;
  assign n70438 = ~n7705 & ~n70437;
  assign n70439 = ~n70418 & ~n70438;
  assign n70440 = n7808 & ~n70439;
  assign n70441 = ~n70408 & ~n70440;
  assign n70442 = n8195 & ~n70441;
  assign n70443 = ~n8196 & ~n70442;
  assign n70444 = ~n8193 & ~n70443;
  assign n70445 = ~n9900 & ~n70399;
  assign n70446 = ~n7723 & ~n70445;
  assign n70447 = ~n9899 & ~n70446;
  assign n70448 = n7714 & ~n70447;
  assign n70449 = ~n70404 & ~n70448;
  assign n70450 = ~n7705 & ~n70449;
  assign n70451 = ~n9898 & ~n70450;
  assign n70452 = ~n7808 & ~n70451;
  assign n70453 = ~n69386 & ~n70399;
  assign n70454 = n7728 & ~n70453;
  assign n70455 = ~n70432 & ~n70454;
  assign n70456 = ~n7723 & ~n70455;
  assign n70457 = ~n69096 & ~n70456;
  assign n70458 = ~n7714 & ~n70457;
  assign n70459 = ~n69095 & ~n70458;
  assign n70460 = ~n7705 & ~n70459;
  assign n70461 = ~n22399 & ~n70460;
  assign n70462 = n7808 & ~n70461;
  assign n70463 = ~n70452 & ~n70462;
  assign n70464 = ~n8195 & ~n70463;
  assign n70465 = ~n11476 & ~n69446;
  assign n70466 = i_hbusreq7 & ~n70465;
  assign n70467 = ~n11504 & ~n69473;
  assign n70468 = ~i_hbusreq7 & ~n70467;
  assign n70469 = ~n70466 & ~n70468;
  assign n70470 = n7924 & ~n70469;
  assign n70471 = ~n10375 & ~n70470;
  assign n70472 = n8214 & ~n70471;
  assign n70473 = n8214 & ~n70472;
  assign n70474 = n8202 & ~n70473;
  assign n70475 = ~n69413 & ~n70474;
  assign n70476 = n7728 & ~n70475;
  assign n70477 = n8214 & ~n70398;
  assign n70478 = ~n8336 & ~n70477;
  assign n70479 = n8202 & ~n70478;
  assign n70480 = ~n69493 & ~n70479;
  assign n70481 = ~n7728 & ~n70480;
  assign n70482 = ~n70476 & ~n70481;
  assign n70483 = ~n7723 & ~n70482;
  assign n70484 = ~n7723 & ~n70483;
  assign n70485 = ~n7714 & ~n70484;
  assign n70486 = ~n7714 & ~n70485;
  assign n70487 = n7705 & ~n70486;
  assign n70488 = n7723 & ~n70480;
  assign n70489 = n7920 & ~n70480;
  assign n70490 = ~n70399 & ~n70489;
  assign n70491 = ~n7723 & ~n70490;
  assign n70492 = ~n70488 & ~n70491;
  assign n70493 = n7714 & ~n70492;
  assign n70494 = ~n70404 & ~n70493;
  assign n70495 = ~n7705 & ~n70494;
  assign n70496 = ~n70487 & ~n70495;
  assign n70497 = ~n7808 & ~n70496;
  assign n70498 = ~n7920 & ~n70475;
  assign n70499 = ~n69861 & ~n70498;
  assign n70500 = n7728 & ~n70499;
  assign n70501 = ~n7920 & ~n70480;
  assign n70502 = ~n69948 & ~n70501;
  assign n70503 = ~n7728 & ~n70502;
  assign n70504 = ~n70500 & ~n70503;
  assign n70505 = ~n7723 & ~n70504;
  assign n70506 = ~n7723 & ~n70505;
  assign n70507 = ~n7714 & ~n70506;
  assign n70508 = ~n7714 & ~n70507;
  assign n70509 = n7705 & ~n70508;
  assign n70510 = ~n70075 & ~n70501;
  assign n70511 = n7728 & ~n70510;
  assign n70512 = ~n70139 & ~n70501;
  assign n70513 = ~n7728 & ~n70512;
  assign n70514 = ~n70511 & ~n70513;
  assign n70515 = n7723 & ~n70514;
  assign n70516 = ~n7723 & ~n70512;
  assign n70517 = ~n70515 & ~n70516;
  assign n70518 = n7714 & ~n70517;
  assign n70519 = n7723 & ~n70512;
  assign n70520 = ~n70229 & ~n70399;
  assign n70521 = n7728 & ~n70520;
  assign n70522 = ~n70432 & ~n70521;
  assign n70523 = ~n7723 & ~n70522;
  assign n70524 = ~n70519 & ~n70523;
  assign n70525 = ~n7714 & ~n70524;
  assign n70526 = ~n70518 & ~n70525;
  assign n70527 = ~n7705 & ~n70526;
  assign n70528 = ~n70509 & ~n70527;
  assign n70529 = n7808 & ~n70528;
  assign n70530 = ~n70497 & ~n70529;
  assign n70531 = n8195 & ~n70530;
  assign n70532 = ~n70464 & ~n70531;
  assign n70533 = n8193 & ~n70532;
  assign n70534 = ~n70444 & ~n70533;
  assign n70535 = n8191 & ~n70534;
  assign n70536 = ~n11594 & ~n66547;
  assign n70537 = i_hbusreq7 & ~n70536;
  assign n70538 = ~n11605 & ~n66574;
  assign n70539 = ~i_hbusreq7 & ~n70538;
  assign n70540 = ~n70537 & ~n70539;
  assign n70541 = n7924 & ~n70540;
  assign n70542 = ~n8337 & ~n70541;
  assign n70543 = ~n7920 & ~n70542;
  assign n70544 = ~n11612 & ~n70543;
  assign n70545 = ~n7723 & ~n70544;
  assign n70546 = ~n11588 & ~n70545;
  assign n70547 = n7714 & ~n70546;
  assign n70548 = ~n7714 & ~n70542;
  assign n70549 = ~n70547 & ~n70548;
  assign n70550 = ~n7705 & ~n70549;
  assign n70551 = ~n11587 & ~n70550;
  assign n70552 = ~n7808 & ~n70551;
  assign n70553 = ~n11622 & ~n66591;
  assign n70554 = n7728 & ~n70553;
  assign n70555 = ~n11625 & ~n66595;
  assign n70556 = ~n7728 & ~n70555;
  assign n70557 = ~n70554 & ~n70556;
  assign n70558 = ~n7723 & ~n70557;
  assign n70559 = ~n7723 & ~n70558;
  assign n70560 = ~n7714 & ~n70559;
  assign n70561 = ~n7714 & ~n70560;
  assign n70562 = n7705 & ~n70561;
  assign n70563 = ~n11625 & ~n66787;
  assign n70564 = n7728 & ~n70563;
  assign n70565 = ~n11625 & ~n67175;
  assign n70566 = ~n7728 & ~n70565;
  assign n70567 = ~n70564 & ~n70566;
  assign n70568 = n7723 & ~n70567;
  assign n70569 = ~n7723 & ~n70565;
  assign n70570 = ~n70568 & ~n70569;
  assign n70571 = n7714 & ~n70570;
  assign n70572 = n7723 & ~n70565;
  assign n70573 = ~n68031 & ~n70543;
  assign n70574 = n7728 & ~n70573;
  assign n70575 = ~n68572 & ~n70543;
  assign n70576 = ~n7728 & ~n70575;
  assign n70577 = ~n70574 & ~n70576;
  assign n70578 = ~n7723 & ~n70577;
  assign n70579 = ~n70572 & ~n70578;
  assign n70580 = ~n7714 & ~n70579;
  assign n70581 = ~n70571 & ~n70580;
  assign n70582 = ~n7705 & ~n70581;
  assign n70583 = ~n70562 & ~n70582;
  assign n70584 = n7808 & ~n70583;
  assign n70585 = ~n70552 & ~n70584;
  assign n70586 = n8195 & ~n70585;
  assign n70587 = ~n8196 & ~n70586;
  assign n70588 = ~n8193 & ~n70587;
  assign n70589 = ~n9900 & ~n70543;
  assign n70590 = ~n7723 & ~n70589;
  assign n70591 = ~n9899 & ~n70590;
  assign n70592 = n7714 & ~n70591;
  assign n70593 = ~n70548 & ~n70592;
  assign n70594 = ~n7705 & ~n70593;
  assign n70595 = ~n9898 & ~n70594;
  assign n70596 = ~n7808 & ~n70595;
  assign n70597 = ~n69386 & ~n70543;
  assign n70598 = n7728 & ~n70597;
  assign n70599 = ~n70576 & ~n70598;
  assign n70600 = ~n7723 & ~n70599;
  assign n70601 = ~n69096 & ~n70600;
  assign n70602 = ~n7714 & ~n70601;
  assign n70603 = ~n69095 & ~n70602;
  assign n70604 = ~n7705 & ~n70603;
  assign n70605 = ~n22399 & ~n70604;
  assign n70606 = n7808 & ~n70605;
  assign n70607 = ~n70596 & ~n70606;
  assign n70608 = ~n8195 & ~n70607;
  assign n70609 = ~n11685 & ~n69446;
  assign n70610 = i_hbusreq7 & ~n70609;
  assign n70611 = ~n11696 & ~n69473;
  assign n70612 = ~i_hbusreq7 & ~n70611;
  assign n70613 = ~n70610 & ~n70612;
  assign n70614 = n7924 & ~n70613;
  assign n70615 = ~n10375 & ~n70614;
  assign n70616 = n8214 & ~n70615;
  assign n70617 = n8214 & ~n70616;
  assign n70618 = n8202 & ~n70617;
  assign n70619 = ~n69413 & ~n70618;
  assign n70620 = n7728 & ~n70619;
  assign n70621 = n8214 & ~n70542;
  assign n70622 = ~n8336 & ~n70621;
  assign n70623 = n8202 & ~n70622;
  assign n70624 = ~n69493 & ~n70623;
  assign n70625 = ~n7728 & ~n70624;
  assign n70626 = ~n70620 & ~n70625;
  assign n70627 = ~n7723 & ~n70626;
  assign n70628 = ~n7723 & ~n70627;
  assign n70629 = ~n7714 & ~n70628;
  assign n70630 = ~n7714 & ~n70629;
  assign n70631 = n7705 & ~n70630;
  assign n70632 = n7723 & ~n70624;
  assign n70633 = n7920 & ~n70624;
  assign n70634 = ~n70543 & ~n70633;
  assign n70635 = ~n7723 & ~n70634;
  assign n70636 = ~n70632 & ~n70635;
  assign n70637 = n7714 & ~n70636;
  assign n70638 = ~n70548 & ~n70637;
  assign n70639 = ~n7705 & ~n70638;
  assign n70640 = ~n70631 & ~n70639;
  assign n70641 = ~n7808 & ~n70640;
  assign n70642 = ~n7920 & ~n70619;
  assign n70643 = ~n69861 & ~n70642;
  assign n70644 = n7728 & ~n70643;
  assign n70645 = ~n7920 & ~n70624;
  assign n70646 = ~n69948 & ~n70645;
  assign n70647 = ~n7728 & ~n70646;
  assign n70648 = ~n70644 & ~n70647;
  assign n70649 = ~n7723 & ~n70648;
  assign n70650 = ~n7723 & ~n70649;
  assign n70651 = ~n7714 & ~n70650;
  assign n70652 = ~n7714 & ~n70651;
  assign n70653 = n7705 & ~n70652;
  assign n70654 = ~n70075 & ~n70645;
  assign n70655 = n7728 & ~n70654;
  assign n70656 = ~n70139 & ~n70645;
  assign n70657 = ~n7728 & ~n70656;
  assign n70658 = ~n70655 & ~n70657;
  assign n70659 = n7723 & ~n70658;
  assign n70660 = ~n7723 & ~n70656;
  assign n70661 = ~n70659 & ~n70660;
  assign n70662 = n7714 & ~n70661;
  assign n70663 = n7723 & ~n70656;
  assign n70664 = ~n70229 & ~n70543;
  assign n70665 = n7728 & ~n70664;
  assign n70666 = ~n70576 & ~n70665;
  assign n70667 = ~n7723 & ~n70666;
  assign n70668 = ~n70663 & ~n70667;
  assign n70669 = ~n7714 & ~n70668;
  assign n70670 = ~n70662 & ~n70669;
  assign n70671 = ~n7705 & ~n70670;
  assign n70672 = ~n70653 & ~n70671;
  assign n70673 = n7808 & ~n70672;
  assign n70674 = ~n70641 & ~n70673;
  assign n70675 = n8195 & ~n70674;
  assign n70676 = ~n70608 & ~n70675;
  assign n70677 = n8193 & ~n70676;
  assign n70678 = ~n70588 & ~n70677;
  assign n70679 = ~n8191 & ~n70678;
  assign n70680 = ~n70535 & ~n70679;
  assign n70681 = ~n8188 & ~n70680;
  assign n70682 = ~n70391 & ~n70681;
  assign n70683 = n8185 & ~n70682;
  assign n70684 = ~n11844 & ~n66545;
  assign n70685 = ~controllable_hmaster3 & ~n70684;
  assign n70686 = ~n8362 & ~n70685;
  assign n70687 = i_hlock7 & ~n70686;
  assign n70688 = ~n11852 & ~n66545;
  assign n70689 = ~controllable_hmaster3 & ~n70688;
  assign n70690 = ~n8362 & ~n70689;
  assign n70691 = ~i_hlock7 & ~n70690;
  assign n70692 = ~n70687 & ~n70691;
  assign n70693 = i_hbusreq7 & ~n70692;
  assign n70694 = i_hbusreq8 & ~n70684;
  assign n70695 = ~n11866 & ~n66570;
  assign n70696 = ~i_hbusreq8 & ~n70695;
  assign n70697 = ~n70694 & ~n70696;
  assign n70698 = ~controllable_hmaster3 & ~n70697;
  assign n70699 = ~n8492 & ~n70698;
  assign n70700 = i_hlock7 & ~n70699;
  assign n70701 = i_hbusreq8 & ~n70688;
  assign n70702 = ~n11880 & ~n66570;
  assign n70703 = ~i_hbusreq8 & ~n70702;
  assign n70704 = ~n70701 & ~n70703;
  assign n70705 = ~controllable_hmaster3 & ~n70704;
  assign n70706 = ~n8492 & ~n70705;
  assign n70707 = ~i_hlock7 & ~n70706;
  assign n70708 = ~n70700 & ~n70707;
  assign n70709 = ~i_hbusreq7 & ~n70708;
  assign n70710 = ~n70693 & ~n70709;
  assign n70711 = n7924 & ~n70710;
  assign n70712 = ~n8337 & ~n70711;
  assign n70713 = ~n7920 & ~n70712;
  assign n70714 = ~n11893 & ~n70713;
  assign n70715 = ~n7723 & ~n70714;
  assign n70716 = ~n11840 & ~n70715;
  assign n70717 = n7714 & ~n70716;
  assign n70718 = ~n7714 & ~n70712;
  assign n70719 = ~n70717 & ~n70718;
  assign n70720 = ~n7705 & ~n70719;
  assign n70721 = ~n11839 & ~n70720;
  assign n70722 = ~n7808 & ~n70721;
  assign n70723 = ~n11903 & ~n66591;
  assign n70724 = n7728 & ~n70723;
  assign n70725 = ~n11906 & ~n66595;
  assign n70726 = ~n7728 & ~n70725;
  assign n70727 = ~n70724 & ~n70726;
  assign n70728 = ~n7723 & ~n70727;
  assign n70729 = ~n7723 & ~n70728;
  assign n70730 = ~n7714 & ~n70729;
  assign n70731 = ~n7714 & ~n70730;
  assign n70732 = n7705 & ~n70731;
  assign n70733 = ~n11906 & ~n66787;
  assign n70734 = n7728 & ~n70733;
  assign n70735 = ~n11906 & ~n67175;
  assign n70736 = ~n7728 & ~n70735;
  assign n70737 = ~n70734 & ~n70736;
  assign n70738 = n7723 & ~n70737;
  assign n70739 = ~n7723 & ~n70735;
  assign n70740 = ~n70738 & ~n70739;
  assign n70741 = n7714 & ~n70740;
  assign n70742 = n7723 & ~n70735;
  assign n70743 = ~n68031 & ~n70713;
  assign n70744 = n7728 & ~n70743;
  assign n70745 = ~n68572 & ~n70713;
  assign n70746 = ~n7728 & ~n70745;
  assign n70747 = ~n70744 & ~n70746;
  assign n70748 = ~n7723 & ~n70747;
  assign n70749 = ~n70742 & ~n70748;
  assign n70750 = ~n7714 & ~n70749;
  assign n70751 = ~n70741 & ~n70750;
  assign n70752 = ~n7705 & ~n70751;
  assign n70753 = ~n70732 & ~n70752;
  assign n70754 = n7808 & ~n70753;
  assign n70755 = ~n70722 & ~n70754;
  assign n70756 = n8195 & ~n70755;
  assign n70757 = ~n8196 & ~n70756;
  assign n70758 = ~n8193 & ~n70757;
  assign n70759 = ~n9900 & ~n70713;
  assign n70760 = ~n7723 & ~n70759;
  assign n70761 = ~n9899 & ~n70760;
  assign n70762 = n7714 & ~n70761;
  assign n70763 = ~n70718 & ~n70762;
  assign n70764 = ~n7705 & ~n70763;
  assign n70765 = ~n9898 & ~n70764;
  assign n70766 = ~n7808 & ~n70765;
  assign n70767 = ~n69386 & ~n70713;
  assign n70768 = n7728 & ~n70767;
  assign n70769 = ~n70746 & ~n70768;
  assign n70770 = ~n7723 & ~n70769;
  assign n70771 = ~n69096 & ~n70770;
  assign n70772 = ~n7714 & ~n70771;
  assign n70773 = ~n69095 & ~n70772;
  assign n70774 = ~n7705 & ~n70773;
  assign n70775 = ~n22399 & ~n70774;
  assign n70776 = n7808 & ~n70775;
  assign n70777 = ~n70766 & ~n70776;
  assign n70778 = ~n8195 & ~n70777;
  assign n70779 = ~n11964 & ~n69444;
  assign n70780 = ~controllable_hmaster3 & ~n70779;
  assign n70781 = ~n10379 & ~n70780;
  assign n70782 = i_hlock7 & ~n70781;
  assign n70783 = ~n11972 & ~n69444;
  assign n70784 = ~controllable_hmaster3 & ~n70783;
  assign n70785 = ~n10379 & ~n70784;
  assign n70786 = ~i_hlock7 & ~n70785;
  assign n70787 = ~n70782 & ~n70786;
  assign n70788 = i_hbusreq7 & ~n70787;
  assign n70789 = i_hbusreq8 & ~n70779;
  assign n70790 = ~n11986 & ~n69469;
  assign n70791 = ~i_hbusreq8 & ~n70790;
  assign n70792 = ~n70789 & ~n70791;
  assign n70793 = ~controllable_hmaster3 & ~n70792;
  assign n70794 = ~n10459 & ~n70793;
  assign n70795 = i_hlock7 & ~n70794;
  assign n70796 = i_hbusreq8 & ~n70783;
  assign n70797 = ~n12000 & ~n69469;
  assign n70798 = ~i_hbusreq8 & ~n70797;
  assign n70799 = ~n70796 & ~n70798;
  assign n70800 = ~controllable_hmaster3 & ~n70799;
  assign n70801 = ~n10459 & ~n70800;
  assign n70802 = ~i_hlock7 & ~n70801;
  assign n70803 = ~n70795 & ~n70802;
  assign n70804 = ~i_hbusreq7 & ~n70803;
  assign n70805 = ~n70788 & ~n70804;
  assign n70806 = n7924 & ~n70805;
  assign n70807 = ~n10375 & ~n70806;
  assign n70808 = n8214 & ~n70807;
  assign n70809 = n8214 & ~n70808;
  assign n70810 = n8202 & ~n70809;
  assign n70811 = ~n69413 & ~n70810;
  assign n70812 = n7728 & ~n70811;
  assign n70813 = n8214 & ~n70712;
  assign n70814 = ~n8336 & ~n70813;
  assign n70815 = n8202 & ~n70814;
  assign n70816 = ~n69493 & ~n70815;
  assign n70817 = ~n7728 & ~n70816;
  assign n70818 = ~n70812 & ~n70817;
  assign n70819 = ~n7723 & ~n70818;
  assign n70820 = ~n7723 & ~n70819;
  assign n70821 = ~n7714 & ~n70820;
  assign n70822 = ~n7714 & ~n70821;
  assign n70823 = n7705 & ~n70822;
  assign n70824 = n7723 & ~n70816;
  assign n70825 = n7920 & ~n70816;
  assign n70826 = ~n70713 & ~n70825;
  assign n70827 = ~n7723 & ~n70826;
  assign n70828 = ~n70824 & ~n70827;
  assign n70829 = n7714 & ~n70828;
  assign n70830 = ~n70718 & ~n70829;
  assign n70831 = ~n7705 & ~n70830;
  assign n70832 = ~n70823 & ~n70831;
  assign n70833 = ~n7808 & ~n70832;
  assign n70834 = ~n7920 & ~n70811;
  assign n70835 = ~n69861 & ~n70834;
  assign n70836 = n7728 & ~n70835;
  assign n70837 = ~n7920 & ~n70816;
  assign n70838 = ~n69948 & ~n70837;
  assign n70839 = ~n7728 & ~n70838;
  assign n70840 = ~n70836 & ~n70839;
  assign n70841 = ~n7723 & ~n70840;
  assign n70842 = ~n7723 & ~n70841;
  assign n70843 = ~n7714 & ~n70842;
  assign n70844 = ~n7714 & ~n70843;
  assign n70845 = n7705 & ~n70844;
  assign n70846 = ~n70075 & ~n70837;
  assign n70847 = n7728 & ~n70846;
  assign n70848 = ~n70139 & ~n70837;
  assign n70849 = ~n7728 & ~n70848;
  assign n70850 = ~n70847 & ~n70849;
  assign n70851 = n7723 & ~n70850;
  assign n70852 = ~n7723 & ~n70848;
  assign n70853 = ~n70851 & ~n70852;
  assign n70854 = n7714 & ~n70853;
  assign n70855 = n7723 & ~n70848;
  assign n70856 = ~n70229 & ~n70713;
  assign n70857 = n7728 & ~n70856;
  assign n70858 = ~n70746 & ~n70857;
  assign n70859 = ~n7723 & ~n70858;
  assign n70860 = ~n70855 & ~n70859;
  assign n70861 = ~n7714 & ~n70860;
  assign n70862 = ~n70854 & ~n70861;
  assign n70863 = ~n7705 & ~n70862;
  assign n70864 = ~n70845 & ~n70863;
  assign n70865 = n7808 & ~n70864;
  assign n70866 = ~n70833 & ~n70865;
  assign n70867 = n8195 & ~n70866;
  assign n70868 = ~n70778 & ~n70867;
  assign n70869 = n8193 & ~n70868;
  assign n70870 = ~n70758 & ~n70869;
  assign n70871 = n8191 & ~n70870;
  assign n70872 = ~n11036 & ~n70685;
  assign n70873 = i_hlock7 & ~n70872;
  assign n70874 = ~n11036 & ~n70689;
  assign n70875 = ~i_hlock7 & ~n70874;
  assign n70876 = ~n70873 & ~n70875;
  assign n70877 = i_hbusreq7 & ~n70876;
  assign n70878 = ~n11051 & ~n70698;
  assign n70879 = i_hlock7 & ~n70878;
  assign n70880 = ~n11051 & ~n70705;
  assign n70881 = ~i_hlock7 & ~n70880;
  assign n70882 = ~n70879 & ~n70881;
  assign n70883 = ~i_hbusreq7 & ~n70882;
  assign n70884 = ~n70877 & ~n70883;
  assign n70885 = n7924 & ~n70884;
  assign n70886 = ~n8337 & ~n70885;
  assign n70887 = ~n7920 & ~n70886;
  assign n70888 = ~n12103 & ~n70887;
  assign n70889 = ~n7723 & ~n70888;
  assign n70890 = ~n12086 & ~n70889;
  assign n70891 = n7714 & ~n70890;
  assign n70892 = ~n7714 & ~n70886;
  assign n70893 = ~n70891 & ~n70892;
  assign n70894 = ~n7705 & ~n70893;
  assign n70895 = ~n12085 & ~n70894;
  assign n70896 = ~n7808 & ~n70895;
  assign n70897 = ~n12113 & ~n66591;
  assign n70898 = n7728 & ~n70897;
  assign n70899 = ~n12116 & ~n66595;
  assign n70900 = ~n7728 & ~n70899;
  assign n70901 = ~n70898 & ~n70900;
  assign n70902 = ~n7723 & ~n70901;
  assign n70903 = ~n7723 & ~n70902;
  assign n70904 = ~n7714 & ~n70903;
  assign n70905 = ~n7714 & ~n70904;
  assign n70906 = n7705 & ~n70905;
  assign n70907 = ~n12116 & ~n66787;
  assign n70908 = n7728 & ~n70907;
  assign n70909 = ~n12116 & ~n67175;
  assign n70910 = ~n7728 & ~n70909;
  assign n70911 = ~n70908 & ~n70910;
  assign n70912 = n7723 & ~n70911;
  assign n70913 = ~n7723 & ~n70909;
  assign n70914 = ~n70912 & ~n70913;
  assign n70915 = n7714 & ~n70914;
  assign n70916 = n7723 & ~n70909;
  assign n70917 = ~n68031 & ~n70887;
  assign n70918 = n7728 & ~n70917;
  assign n70919 = ~n68572 & ~n70887;
  assign n70920 = ~n7728 & ~n70919;
  assign n70921 = ~n70918 & ~n70920;
  assign n70922 = ~n7723 & ~n70921;
  assign n70923 = ~n70916 & ~n70922;
  assign n70924 = ~n7714 & ~n70923;
  assign n70925 = ~n70915 & ~n70924;
  assign n70926 = ~n7705 & ~n70925;
  assign n70927 = ~n70906 & ~n70926;
  assign n70928 = n7808 & ~n70927;
  assign n70929 = ~n70896 & ~n70928;
  assign n70930 = n8195 & ~n70929;
  assign n70931 = ~n8196 & ~n70930;
  assign n70932 = ~n8193 & ~n70931;
  assign n70933 = ~n9900 & ~n70887;
  assign n70934 = ~n7723 & ~n70933;
  assign n70935 = ~n9899 & ~n70934;
  assign n70936 = n7714 & ~n70935;
  assign n70937 = ~n70892 & ~n70936;
  assign n70938 = ~n7705 & ~n70937;
  assign n70939 = ~n9898 & ~n70938;
  assign n70940 = ~n7808 & ~n70939;
  assign n70941 = ~n69386 & ~n70887;
  assign n70942 = n7728 & ~n70941;
  assign n70943 = ~n70920 & ~n70942;
  assign n70944 = ~n7723 & ~n70943;
  assign n70945 = ~n69096 & ~n70944;
  assign n70946 = ~n7714 & ~n70945;
  assign n70947 = ~n69095 & ~n70946;
  assign n70948 = ~n7705 & ~n70947;
  assign n70949 = ~n22399 & ~n70948;
  assign n70950 = n7808 & ~n70949;
  assign n70951 = ~n70940 & ~n70950;
  assign n70952 = ~n8195 & ~n70951;
  assign n70953 = ~n11136 & ~n70780;
  assign n70954 = i_hlock7 & ~n70953;
  assign n70955 = ~n11136 & ~n70784;
  assign n70956 = ~i_hlock7 & ~n70955;
  assign n70957 = ~n70954 & ~n70956;
  assign n70958 = i_hbusreq7 & ~n70957;
  assign n70959 = ~n11164 & ~n70793;
  assign n70960 = i_hlock7 & ~n70959;
  assign n70961 = ~n11164 & ~n70800;
  assign n70962 = ~i_hlock7 & ~n70961;
  assign n70963 = ~n70960 & ~n70962;
  assign n70964 = ~i_hbusreq7 & ~n70963;
  assign n70965 = ~n70958 & ~n70964;
  assign n70966 = n7924 & ~n70965;
  assign n70967 = ~n10375 & ~n70966;
  assign n70968 = n8214 & ~n70967;
  assign n70969 = n8214 & ~n70968;
  assign n70970 = n8202 & ~n70969;
  assign n70971 = ~n69413 & ~n70970;
  assign n70972 = n7728 & ~n70971;
  assign n70973 = n8214 & ~n70886;
  assign n70974 = ~n8336 & ~n70973;
  assign n70975 = n8202 & ~n70974;
  assign n70976 = ~n69493 & ~n70975;
  assign n70977 = ~n7728 & ~n70976;
  assign n70978 = ~n70972 & ~n70977;
  assign n70979 = ~n7723 & ~n70978;
  assign n70980 = ~n7723 & ~n70979;
  assign n70981 = ~n7714 & ~n70980;
  assign n70982 = ~n7714 & ~n70981;
  assign n70983 = n7705 & ~n70982;
  assign n70984 = n7723 & ~n70976;
  assign n70985 = n7920 & ~n70976;
  assign n70986 = ~n70887 & ~n70985;
  assign n70987 = ~n7723 & ~n70986;
  assign n70988 = ~n70984 & ~n70987;
  assign n70989 = n7714 & ~n70988;
  assign n70990 = ~n70892 & ~n70989;
  assign n70991 = ~n7705 & ~n70990;
  assign n70992 = ~n70983 & ~n70991;
  assign n70993 = ~n7808 & ~n70992;
  assign n70994 = ~n7920 & ~n70971;
  assign n70995 = ~n69861 & ~n70994;
  assign n70996 = n7728 & ~n70995;
  assign n70997 = ~n7920 & ~n70976;
  assign n70998 = ~n69948 & ~n70997;
  assign n70999 = ~n7728 & ~n70998;
  assign n71000 = ~n70996 & ~n70999;
  assign n71001 = ~n7723 & ~n71000;
  assign n71002 = ~n7723 & ~n71001;
  assign n71003 = ~n7714 & ~n71002;
  assign n71004 = ~n7714 & ~n71003;
  assign n71005 = n7705 & ~n71004;
  assign n71006 = ~n70075 & ~n70997;
  assign n71007 = n7728 & ~n71006;
  assign n71008 = ~n70139 & ~n70997;
  assign n71009 = ~n7728 & ~n71008;
  assign n71010 = ~n71007 & ~n71009;
  assign n71011 = n7723 & ~n71010;
  assign n71012 = ~n7723 & ~n71008;
  assign n71013 = ~n71011 & ~n71012;
  assign n71014 = n7714 & ~n71013;
  assign n71015 = n7723 & ~n71008;
  assign n71016 = ~n70229 & ~n70887;
  assign n71017 = n7728 & ~n71016;
  assign n71018 = ~n70920 & ~n71017;
  assign n71019 = ~n7723 & ~n71018;
  assign n71020 = ~n71015 & ~n71019;
  assign n71021 = ~n7714 & ~n71020;
  assign n71022 = ~n71014 & ~n71021;
  assign n71023 = ~n7705 & ~n71022;
  assign n71024 = ~n71005 & ~n71023;
  assign n71025 = n7808 & ~n71024;
  assign n71026 = ~n70993 & ~n71025;
  assign n71027 = n8195 & ~n71026;
  assign n71028 = ~n70952 & ~n71027;
  assign n71029 = n8193 & ~n71028;
  assign n71030 = ~n70932 & ~n71029;
  assign n71031 = ~n8191 & ~n71030;
  assign n71032 = ~n70871 & ~n71031;
  assign n71033 = n8188 & ~n71032;
  assign n71034 = ~n11359 & ~n70685;
  assign n71035 = i_hlock7 & ~n71034;
  assign n71036 = ~n11359 & ~n70689;
  assign n71037 = ~i_hlock7 & ~n71036;
  assign n71038 = ~n71035 & ~n71037;
  assign n71039 = i_hbusreq7 & ~n71038;
  assign n71040 = ~n11385 & ~n70698;
  assign n71041 = i_hlock7 & ~n71040;
  assign n71042 = ~n11385 & ~n70705;
  assign n71043 = ~i_hlock7 & ~n71042;
  assign n71044 = ~n71041 & ~n71043;
  assign n71045 = ~i_hbusreq7 & ~n71044;
  assign n71046 = ~n71039 & ~n71045;
  assign n71047 = n7924 & ~n71046;
  assign n71048 = ~n8337 & ~n71047;
  assign n71049 = ~n7920 & ~n71048;
  assign n71050 = ~n12279 & ~n71049;
  assign n71051 = ~n7723 & ~n71050;
  assign n71052 = ~n12262 & ~n71051;
  assign n71053 = n7714 & ~n71052;
  assign n71054 = ~n7714 & ~n71048;
  assign n71055 = ~n71053 & ~n71054;
  assign n71056 = ~n7705 & ~n71055;
  assign n71057 = ~n12261 & ~n71056;
  assign n71058 = ~n7808 & ~n71057;
  assign n71059 = ~n12289 & ~n66591;
  assign n71060 = n7728 & ~n71059;
  assign n71061 = ~n12292 & ~n66595;
  assign n71062 = ~n7728 & ~n71061;
  assign n71063 = ~n71060 & ~n71062;
  assign n71064 = ~n7723 & ~n71063;
  assign n71065 = ~n7723 & ~n71064;
  assign n71066 = ~n7714 & ~n71065;
  assign n71067 = ~n7714 & ~n71066;
  assign n71068 = n7705 & ~n71067;
  assign n71069 = ~n12292 & ~n66787;
  assign n71070 = n7728 & ~n71069;
  assign n71071 = ~n12292 & ~n67175;
  assign n71072 = ~n7728 & ~n71071;
  assign n71073 = ~n71070 & ~n71072;
  assign n71074 = n7723 & ~n71073;
  assign n71075 = ~n7723 & ~n71071;
  assign n71076 = ~n71074 & ~n71075;
  assign n71077 = n7714 & ~n71076;
  assign n71078 = n7723 & ~n71071;
  assign n71079 = ~n68031 & ~n71049;
  assign n71080 = n7728 & ~n71079;
  assign n71081 = ~n68572 & ~n71049;
  assign n71082 = ~n7728 & ~n71081;
  assign n71083 = ~n71080 & ~n71082;
  assign n71084 = ~n7723 & ~n71083;
  assign n71085 = ~n71078 & ~n71084;
  assign n71086 = ~n7714 & ~n71085;
  assign n71087 = ~n71077 & ~n71086;
  assign n71088 = ~n7705 & ~n71087;
  assign n71089 = ~n71068 & ~n71088;
  assign n71090 = n7808 & ~n71089;
  assign n71091 = ~n71058 & ~n71090;
  assign n71092 = n8195 & ~n71091;
  assign n71093 = ~n8196 & ~n71092;
  assign n71094 = ~n8193 & ~n71093;
  assign n71095 = ~n9900 & ~n71049;
  assign n71096 = ~n7723 & ~n71095;
  assign n71097 = ~n9899 & ~n71096;
  assign n71098 = n7714 & ~n71097;
  assign n71099 = ~n71054 & ~n71098;
  assign n71100 = ~n7705 & ~n71099;
  assign n71101 = ~n9898 & ~n71100;
  assign n71102 = ~n7808 & ~n71101;
  assign n71103 = ~n69386 & ~n71049;
  assign n71104 = n7728 & ~n71103;
  assign n71105 = ~n71082 & ~n71104;
  assign n71106 = ~n7723 & ~n71105;
  assign n71107 = ~n69096 & ~n71106;
  assign n71108 = ~n7714 & ~n71107;
  assign n71109 = ~n69095 & ~n71108;
  assign n71110 = ~n7705 & ~n71109;
  assign n71111 = ~n22399 & ~n71110;
  assign n71112 = n7808 & ~n71111;
  assign n71113 = ~n71102 & ~n71112;
  assign n71114 = ~n8195 & ~n71113;
  assign n71115 = ~n11476 & ~n70780;
  assign n71116 = i_hlock7 & ~n71115;
  assign n71117 = ~n11476 & ~n70784;
  assign n71118 = ~i_hlock7 & ~n71117;
  assign n71119 = ~n71116 & ~n71118;
  assign n71120 = i_hbusreq7 & ~n71119;
  assign n71121 = ~n11504 & ~n70793;
  assign n71122 = i_hlock7 & ~n71121;
  assign n71123 = ~n11504 & ~n70800;
  assign n71124 = ~i_hlock7 & ~n71123;
  assign n71125 = ~n71122 & ~n71124;
  assign n71126 = ~i_hbusreq7 & ~n71125;
  assign n71127 = ~n71120 & ~n71126;
  assign n71128 = n7924 & ~n71127;
  assign n71129 = ~n10375 & ~n71128;
  assign n71130 = n8214 & ~n71129;
  assign n71131 = n8214 & ~n71130;
  assign n71132 = n8202 & ~n71131;
  assign n71133 = ~n69413 & ~n71132;
  assign n71134 = n7728 & ~n71133;
  assign n71135 = n8214 & ~n71048;
  assign n71136 = ~n8336 & ~n71135;
  assign n71137 = n8202 & ~n71136;
  assign n71138 = ~n69493 & ~n71137;
  assign n71139 = ~n7728 & ~n71138;
  assign n71140 = ~n71134 & ~n71139;
  assign n71141 = ~n7723 & ~n71140;
  assign n71142 = ~n7723 & ~n71141;
  assign n71143 = ~n7714 & ~n71142;
  assign n71144 = ~n7714 & ~n71143;
  assign n71145 = n7705 & ~n71144;
  assign n71146 = n7723 & ~n71138;
  assign n71147 = n7920 & ~n71138;
  assign n71148 = ~n71049 & ~n71147;
  assign n71149 = ~n7723 & ~n71148;
  assign n71150 = ~n71146 & ~n71149;
  assign n71151 = n7714 & ~n71150;
  assign n71152 = ~n71054 & ~n71151;
  assign n71153 = ~n7705 & ~n71152;
  assign n71154 = ~n71145 & ~n71153;
  assign n71155 = ~n7808 & ~n71154;
  assign n71156 = ~n7920 & ~n71133;
  assign n71157 = ~n69861 & ~n71156;
  assign n71158 = n7728 & ~n71157;
  assign n71159 = ~n7920 & ~n71138;
  assign n71160 = ~n69948 & ~n71159;
  assign n71161 = ~n7728 & ~n71160;
  assign n71162 = ~n71158 & ~n71161;
  assign n71163 = ~n7723 & ~n71162;
  assign n71164 = ~n7723 & ~n71163;
  assign n71165 = ~n7714 & ~n71164;
  assign n71166 = ~n7714 & ~n71165;
  assign n71167 = n7705 & ~n71166;
  assign n71168 = ~n70075 & ~n71159;
  assign n71169 = n7728 & ~n71168;
  assign n71170 = ~n70139 & ~n71159;
  assign n71171 = ~n7728 & ~n71170;
  assign n71172 = ~n71169 & ~n71171;
  assign n71173 = n7723 & ~n71172;
  assign n71174 = ~n7723 & ~n71170;
  assign n71175 = ~n71173 & ~n71174;
  assign n71176 = n7714 & ~n71175;
  assign n71177 = n7723 & ~n71170;
  assign n71178 = ~n70229 & ~n71049;
  assign n71179 = n7728 & ~n71178;
  assign n71180 = ~n71082 & ~n71179;
  assign n71181 = ~n7723 & ~n71180;
  assign n71182 = ~n71177 & ~n71181;
  assign n71183 = ~n7714 & ~n71182;
  assign n71184 = ~n71176 & ~n71183;
  assign n71185 = ~n7705 & ~n71184;
  assign n71186 = ~n71167 & ~n71185;
  assign n71187 = n7808 & ~n71186;
  assign n71188 = ~n71155 & ~n71187;
  assign n71189 = n8195 & ~n71188;
  assign n71190 = ~n71114 & ~n71189;
  assign n71191 = n8193 & ~n71190;
  assign n71192 = ~n71094 & ~n71191;
  assign n71193 = n8191 & ~n71192;
  assign n71194 = ~n11594 & ~n70685;
  assign n71195 = i_hlock7 & ~n71194;
  assign n71196 = ~n11594 & ~n70689;
  assign n71197 = ~i_hlock7 & ~n71196;
  assign n71198 = ~n71195 & ~n71197;
  assign n71199 = i_hbusreq7 & ~n71198;
  assign n71200 = ~n11605 & ~n70698;
  assign n71201 = i_hlock7 & ~n71200;
  assign n71202 = ~n11605 & ~n70705;
  assign n71203 = ~i_hlock7 & ~n71202;
  assign n71204 = ~n71201 & ~n71203;
  assign n71205 = ~i_hbusreq7 & ~n71204;
  assign n71206 = ~n71199 & ~n71205;
  assign n71207 = n7924 & ~n71206;
  assign n71208 = ~n8337 & ~n71207;
  assign n71209 = ~n7920 & ~n71208;
  assign n71210 = ~n12453 & ~n71209;
  assign n71211 = ~n7723 & ~n71210;
  assign n71212 = ~n12436 & ~n71211;
  assign n71213 = n7714 & ~n71212;
  assign n71214 = ~n7714 & ~n71208;
  assign n71215 = ~n71213 & ~n71214;
  assign n71216 = ~n7705 & ~n71215;
  assign n71217 = ~n12435 & ~n71216;
  assign n71218 = ~n7808 & ~n71217;
  assign n71219 = ~n12463 & ~n66591;
  assign n71220 = n7728 & ~n71219;
  assign n71221 = ~n12466 & ~n66595;
  assign n71222 = ~n7728 & ~n71221;
  assign n71223 = ~n71220 & ~n71222;
  assign n71224 = ~n7723 & ~n71223;
  assign n71225 = ~n7723 & ~n71224;
  assign n71226 = ~n7714 & ~n71225;
  assign n71227 = ~n7714 & ~n71226;
  assign n71228 = n7705 & ~n71227;
  assign n71229 = ~n12466 & ~n66787;
  assign n71230 = n7728 & ~n71229;
  assign n71231 = ~n12466 & ~n67175;
  assign n71232 = ~n7728 & ~n71231;
  assign n71233 = ~n71230 & ~n71232;
  assign n71234 = n7723 & ~n71233;
  assign n71235 = ~n7723 & ~n71231;
  assign n71236 = ~n71234 & ~n71235;
  assign n71237 = n7714 & ~n71236;
  assign n71238 = n7723 & ~n71231;
  assign n71239 = ~n68031 & ~n71209;
  assign n71240 = n7728 & ~n71239;
  assign n71241 = ~n68572 & ~n71209;
  assign n71242 = ~n7728 & ~n71241;
  assign n71243 = ~n71240 & ~n71242;
  assign n71244 = ~n7723 & ~n71243;
  assign n71245 = ~n71238 & ~n71244;
  assign n71246 = ~n7714 & ~n71245;
  assign n71247 = ~n71237 & ~n71246;
  assign n71248 = ~n7705 & ~n71247;
  assign n71249 = ~n71228 & ~n71248;
  assign n71250 = n7808 & ~n71249;
  assign n71251 = ~n71218 & ~n71250;
  assign n71252 = n8195 & ~n71251;
  assign n71253 = ~n8196 & ~n71252;
  assign n71254 = ~n8193 & ~n71253;
  assign n71255 = ~n9900 & ~n71209;
  assign n71256 = ~n7723 & ~n71255;
  assign n71257 = ~n9899 & ~n71256;
  assign n71258 = n7714 & ~n71257;
  assign n71259 = ~n71214 & ~n71258;
  assign n71260 = ~n7705 & ~n71259;
  assign n71261 = ~n9898 & ~n71260;
  assign n71262 = ~n7808 & ~n71261;
  assign n71263 = ~n69386 & ~n71209;
  assign n71264 = n7728 & ~n71263;
  assign n71265 = ~n71242 & ~n71264;
  assign n71266 = ~n7723 & ~n71265;
  assign n71267 = ~n69096 & ~n71266;
  assign n71268 = ~n7714 & ~n71267;
  assign n71269 = ~n69095 & ~n71268;
  assign n71270 = ~n7705 & ~n71269;
  assign n71271 = ~n22399 & ~n71270;
  assign n71272 = n7808 & ~n71271;
  assign n71273 = ~n71262 & ~n71272;
  assign n71274 = ~n8195 & ~n71273;
  assign n71275 = ~n11685 & ~n70780;
  assign n71276 = i_hlock7 & ~n71275;
  assign n71277 = ~n11685 & ~n70784;
  assign n71278 = ~i_hlock7 & ~n71277;
  assign n71279 = ~n71276 & ~n71278;
  assign n71280 = i_hbusreq7 & ~n71279;
  assign n71281 = ~n11696 & ~n70793;
  assign n71282 = i_hlock7 & ~n71281;
  assign n71283 = ~n11696 & ~n70800;
  assign n71284 = ~i_hlock7 & ~n71283;
  assign n71285 = ~n71282 & ~n71284;
  assign n71286 = ~i_hbusreq7 & ~n71285;
  assign n71287 = ~n71280 & ~n71286;
  assign n71288 = n7924 & ~n71287;
  assign n71289 = ~n10375 & ~n71288;
  assign n71290 = n8214 & ~n71289;
  assign n71291 = n8214 & ~n71290;
  assign n71292 = n8202 & ~n71291;
  assign n71293 = ~n69413 & ~n71292;
  assign n71294 = n7728 & ~n71293;
  assign n71295 = n8214 & ~n71208;
  assign n71296 = ~n8336 & ~n71295;
  assign n71297 = n8202 & ~n71296;
  assign n71298 = ~n69493 & ~n71297;
  assign n71299 = ~n7728 & ~n71298;
  assign n71300 = ~n71294 & ~n71299;
  assign n71301 = ~n7723 & ~n71300;
  assign n71302 = ~n7723 & ~n71301;
  assign n71303 = ~n7714 & ~n71302;
  assign n71304 = ~n7714 & ~n71303;
  assign n71305 = n7705 & ~n71304;
  assign n71306 = n7723 & ~n71298;
  assign n71307 = n7920 & ~n71298;
  assign n71308 = ~n71209 & ~n71307;
  assign n71309 = ~n7723 & ~n71308;
  assign n71310 = ~n71306 & ~n71309;
  assign n71311 = n7714 & ~n71310;
  assign n71312 = ~n71214 & ~n71311;
  assign n71313 = ~n7705 & ~n71312;
  assign n71314 = ~n71305 & ~n71313;
  assign n71315 = ~n7808 & ~n71314;
  assign n71316 = ~n7920 & ~n71293;
  assign n71317 = ~n69861 & ~n71316;
  assign n71318 = n7728 & ~n71317;
  assign n71319 = ~n7920 & ~n71298;
  assign n71320 = ~n69948 & ~n71319;
  assign n71321 = ~n7728 & ~n71320;
  assign n71322 = ~n71318 & ~n71321;
  assign n71323 = ~n7723 & ~n71322;
  assign n71324 = ~n7723 & ~n71323;
  assign n71325 = ~n7714 & ~n71324;
  assign n71326 = ~n7714 & ~n71325;
  assign n71327 = n7705 & ~n71326;
  assign n71328 = ~n70075 & ~n71319;
  assign n71329 = n7728 & ~n71328;
  assign n71330 = ~n70139 & ~n71319;
  assign n71331 = ~n7728 & ~n71330;
  assign n71332 = ~n71329 & ~n71331;
  assign n71333 = n7723 & ~n71332;
  assign n71334 = ~n7723 & ~n71330;
  assign n71335 = ~n71333 & ~n71334;
  assign n71336 = n7714 & ~n71335;
  assign n71337 = n7723 & ~n71330;
  assign n71338 = ~n70229 & ~n71209;
  assign n71339 = n7728 & ~n71338;
  assign n71340 = ~n71242 & ~n71339;
  assign n71341 = ~n7723 & ~n71340;
  assign n71342 = ~n71337 & ~n71341;
  assign n71343 = ~n7714 & ~n71342;
  assign n71344 = ~n71336 & ~n71343;
  assign n71345 = ~n7705 & ~n71344;
  assign n71346 = ~n71327 & ~n71345;
  assign n71347 = n7808 & ~n71346;
  assign n71348 = ~n71315 & ~n71347;
  assign n71349 = n8195 & ~n71348;
  assign n71350 = ~n71274 & ~n71349;
  assign n71351 = n8193 & ~n71350;
  assign n71352 = ~n71254 & ~n71351;
  assign n71353 = ~n8191 & ~n71352;
  assign n71354 = ~n71193 & ~n71353;
  assign n71355 = ~n8188 & ~n71354;
  assign n71356 = ~n71033 & ~n71355;
  assign n71357 = ~n8185 & ~n71356;
  assign n71358 = ~n70683 & ~n71357;
  assign n71359 = ~controllable_hgrant8 & ~n71358;
  assign n71360 = ~n12606 & ~n71359;
  assign n71361 = ~controllable_nhgrant0 & ~n71360;
  assign n71362 = ~n66504 & ~n71361;
  assign n71363 = ~controllable_hgrant7 & ~n71362;
  assign n71364 = ~n35184 & ~n71363;
  assign n71365 = ~controllable_hgrant9 & ~n71364;
  assign n71366 = ~n26636 & ~n71365;
  assign n71367 = ~n7593 & ~n71366;
  assign n71368 = ~n8182 & ~n71367;
  assign n71369 = n7592 & n71368;
  assign n71370 = n7592 & ~n71369;
  assign inductivity_check  = ~n7571 & n71370;
endmodule


