// Benchmark "genbuf12b4y_cert" written by ABC on Sun Jul 30 11:41:47 2017

module genbuf12b4y_cert ( 
    n75, reg_i_StoB_REQ4_out, reg_controllable_SLC1_out, sys_fair8done_out,
    reg_i_RtoB_ACK1_out, reg_i_StoB_REQ3_out, reg_controllable_SLC2_out,
    sys_fair7done_out, reg_i_StoB_REQ2_out, reg_controllable_SLC3_out,
    sys_fair9done_out, reg_controllable_BtoS_ACK10_out, env_fair1done_out,
    reg_i_StoB_REQ1_out, reg_controllable_BtoS_ACK11_out,
    sys_fair10done_out, reg_i_StoB_REQ0_out, sys_fair6done_out,
    reg_controllable_BtoR_REQ0_out, reg_controllable_DEQ_out,
    sys_fair11done_out, sys_fair5done_out, reg_controllable_BtoR_REQ1_out,
    reg_controllable_ENQ_out, sys_fair12done_out, sys_fair4done_out,
    env_fair0done_out, reg_controllable_BtoS_ACK0_out, reg_nstateG7_1_out,
    reg_controllable_BtoS_ACK1_out, reg_controllable_BtoS_ACK2_out,
    sys_fair3done_out, reg_stateG7_0_out, fair_cnt<0>_out ,
    fair_cnt<1>_out , fair_cnt<2>_out , reg_controllable_BtoS_ACK3_out,
    sys_fair2done_out, reg_controllable_BtoS_ACK4_out,
    reg_controllable_BtoS_ACK5_out, reg_controllable_BtoS_ACK6_out,
    sys_fair1done_out, reg_controllable_BtoS_ACK7_out, reg_i_nEMPTY_out,
    reg_controllable_BtoS_ACK8_out, reg_stateG12_out, sys_fair0done_out,
    reg_controllable_BtoS_ACK9_out, reg_i_FULL_out, reg_i_StoB_REQ9_out,
    env_safe_err_happened_out, reg_i_StoB_REQ8_out, reg_i_StoB_REQ7_out,
    reg_i_StoB_REQ11_out, reg_i_StoB_REQ6_out, reg_i_StoB_REQ10_out,
    reg_i_RtoB_ACK0_out, reg_i_StoB_REQ5_out, reg_controllable_SLC0_out,
    i_StoB_REQ0, i_StoB_REQ1, i_FULL, i_StoB_REQ2, i_StoB_REQ3,
    i_StoB_REQ4, i_StoB_REQ5, i_StoB_REQ6, i_StoB_REQ7, i_StoB_REQ8,
    i_StoB_REQ9, i_StoB_REQ10, i_StoB_REQ11, i_nEMPTY, i_RtoB_ACK1,
    i_RtoB_ACK0, controllable_SLC2, controllable_SLC3, controllable_DEQ,
    controllable_BtoR_REQ0, controllable_BtoR_REQ1, controllable_BtoS_ACK0,
    controllable_BtoS_ACK1, controllable_BtoS_ACK2, controllable_BtoS_ACK3,
    controllable_BtoS_ACK4, controllable_BtoS_ACK5, controllable_BtoS_ACK6,
    controllable_BtoS_ACK7, controllable_BtoS_ACK8, controllable_BtoS_ACK9,
    controllable_BtoS_ACK10, controllable_ENQ, controllable_BtoS_ACK11,
    controllable_SLC0, controllable_SLC1,
    inductivity_check   );
  input  n75, reg_i_StoB_REQ4_out, reg_controllable_SLC1_out,
    sys_fair8done_out, reg_i_RtoB_ACK1_out, reg_i_StoB_REQ3_out,
    reg_controllable_SLC2_out, sys_fair7done_out, reg_i_StoB_REQ2_out,
    reg_controllable_SLC3_out, sys_fair9done_out,
    reg_controllable_BtoS_ACK10_out, env_fair1done_out,
    reg_i_StoB_REQ1_out, reg_controllable_BtoS_ACK11_out,
    sys_fair10done_out, reg_i_StoB_REQ0_out, sys_fair6done_out,
    reg_controllable_BtoR_REQ0_out, reg_controllable_DEQ_out,
    sys_fair11done_out, sys_fair5done_out, reg_controllable_BtoR_REQ1_out,
    reg_controllable_ENQ_out, sys_fair12done_out, sys_fair4done_out,
    env_fair0done_out, reg_controllable_BtoS_ACK0_out, reg_nstateG7_1_out,
    reg_controllable_BtoS_ACK1_out, reg_controllable_BtoS_ACK2_out,
    sys_fair3done_out, reg_stateG7_0_out, fair_cnt<0>_out ,
    fair_cnt<1>_out , fair_cnt<2>_out , reg_controllable_BtoS_ACK3_out,
    sys_fair2done_out, reg_controllable_BtoS_ACK4_out,
    reg_controllable_BtoS_ACK5_out, reg_controllable_BtoS_ACK6_out,
    sys_fair1done_out, reg_controllable_BtoS_ACK7_out, reg_i_nEMPTY_out,
    reg_controllable_BtoS_ACK8_out, reg_stateG12_out, sys_fair0done_out,
    reg_controllable_BtoS_ACK9_out, reg_i_FULL_out, reg_i_StoB_REQ9_out,
    env_safe_err_happened_out, reg_i_StoB_REQ8_out, reg_i_StoB_REQ7_out,
    reg_i_StoB_REQ11_out, reg_i_StoB_REQ6_out, reg_i_StoB_REQ10_out,
    reg_i_RtoB_ACK0_out, reg_i_StoB_REQ5_out, reg_controllable_SLC0_out,
    i_StoB_REQ0, i_StoB_REQ1, i_FULL, i_StoB_REQ2, i_StoB_REQ3,
    i_StoB_REQ4, i_StoB_REQ5, i_StoB_REQ6, i_StoB_REQ7, i_StoB_REQ8,
    i_StoB_REQ9, i_StoB_REQ10, i_StoB_REQ11, i_nEMPTY, i_RtoB_ACK1,
    i_RtoB_ACK0, controllable_SLC2, controllable_SLC3, controllable_DEQ,
    controllable_BtoR_REQ0, controllable_BtoR_REQ1, controllable_BtoS_ACK0,
    controllable_BtoS_ACK1, controllable_BtoS_ACK2, controllable_BtoS_ACK3,
    controllable_BtoS_ACK4, controllable_BtoS_ACK5, controllable_BtoS_ACK6,
    controllable_BtoS_ACK7, controllable_BtoS_ACK8, controllable_BtoS_ACK9,
    controllable_BtoS_ACK10, controllable_ENQ, controllable_BtoS_ACK11,
    controllable_SLC0, controllable_SLC1;
  output inductivity_check ;
  wire n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
    n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
    n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
    n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
    n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
    n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
    n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
    n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
    n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
    n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
    n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
    n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
    n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
    n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
    n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
    n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
    n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
    n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
    n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
    n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
    n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
    n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
    n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
    n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
    n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
    n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
    n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
    n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
    n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
    n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
    n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
    n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
    n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
    n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
    n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
    n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
    n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
    n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
    n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
    n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
    n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
    n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
    n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
    n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
    n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
    n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
    n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
    n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
    n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
    n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
    n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
    n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
    n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
    n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
    n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
    n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
    n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
    n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
    n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
    n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
    n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
    n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
    n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
    n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
    n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
    n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
    n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
    n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
    n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
    n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
    n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
    n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
    n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
    n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
    n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
    n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
    n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
    n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
    n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
    n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
    n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
    n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
    n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
    n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
    n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
    n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
    n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
    n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
    n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
    n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
    n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
    n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
    n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
    n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
    n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
    n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
    n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
    n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
    n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
    n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
    n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
    n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
    n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
    n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
    n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
    n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
    n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
    n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
    n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
    n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
    n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
    n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
    n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
    n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
    n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
    n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
    n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
    n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
    n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
    n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
    n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
    n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
    n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
    n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
    n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
    n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
    n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
    n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
    n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
    n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
    n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
    n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
    n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
    n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
    n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
    n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
    n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
    n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
    n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
    n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
    n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
    n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
    n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
    n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
    n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
    n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
    n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
    n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
    n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
    n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
    n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
    n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
    n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
    n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
    n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796,
    n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806,
    n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816,
    n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
    n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
    n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
    n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
    n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
    n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876,
    n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
    n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
    n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
    n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
    n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
    n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
    n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
    n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956,
    n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
    n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976,
    n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
    n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996,
    n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
    n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
    n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
    n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036,
    n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046,
    n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056,
    n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
    n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076,
    n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086,
    n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
    n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
    n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
    n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
    n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
    n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
    n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
    n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
    n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
    n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
    n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
    n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
    n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
    n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
    n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
    n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
    n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
    n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
    n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
    n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
    n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
    n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
    n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
    n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
    n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
    n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
    n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
    n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
    n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
    n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
    n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
    n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
    n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
    n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
    n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
    n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
    n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
    n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
    n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
    n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
    n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
    n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506,
    n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516,
    n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
    n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536,
    n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
    n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
    n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
    n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
    n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
    n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
    n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
    n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
    n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
    n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
    n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
    n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
    n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
    n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
    n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
    n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
    n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
    n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
    n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726,
    n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
    n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
    n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
    n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
    n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
    n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
    n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
    n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
    n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
    n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826,
    n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836,
    n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846,
    n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856,
    n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866,
    n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876,
    n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
    n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896,
    n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906,
    n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916,
    n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926,
    n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936,
    n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946,
    n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956,
    n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966,
    n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976,
    n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986,
    n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996,
    n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006,
    n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016,
    n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026,
    n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036,
    n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046,
    n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056,
    n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066,
    n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076,
    n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086,
    n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096,
    n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106,
    n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116,
    n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126,
    n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136,
    n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146,
    n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156,
    n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166,
    n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176,
    n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186,
    n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
    n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
    n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
    n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226,
    n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
    n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
    n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
    n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
    n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
    n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
    n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
    n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
    n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
    n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
    n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
    n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
    n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
    n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
    n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
    n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
    n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396,
    n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
    n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
    n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426,
    n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
    n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
    n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456,
    n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
    n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
    n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
    n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
    n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
    n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
    n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
    n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
    n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
    n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
    n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
    n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
    n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
    n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
    n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
    n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616,
    n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
    n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
    n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
    n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
    n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
    n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
    n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686,
    n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
    n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706,
    n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
    n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
    n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
    n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
    n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
    n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
    n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
    n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
    n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
    n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
    n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
    n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
    n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
    n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
    n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856,
    n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866,
    n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876,
    n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886,
    n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896,
    n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906,
    n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
    n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926,
    n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936,
    n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946,
    n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
    n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
    n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
    n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
    n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
    n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
    n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
    n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
    n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
    n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046,
    n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
    n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
    n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
    n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
    n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
    n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
    n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
    n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
    n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
    n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
    n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
    n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
    n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
    n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
    n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
    n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
    n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
    n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
    n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
    n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
    n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
    n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
    n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
    n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
    n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
    n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
    n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
    n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
    n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
    n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
    n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
    n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
    n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
    n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
    n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
    n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
    n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
    n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
    n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
    n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
    n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
    n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
    n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
    n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
    n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
    n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
    n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
    n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
    n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
    n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
    n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
    n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
    n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
    n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
    n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
    n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
    n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
    n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
    n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
    n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
    n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
    n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
    n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
    n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
    n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
    n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
    n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
    n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
    n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
    n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
    n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
    n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
    n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
    n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
    n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
    n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
    n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
    n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
    n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
    n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
    n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
    n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
    n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
    n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
    n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
    n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
    n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
    n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
    n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
    n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
    n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
    n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
    n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
    n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
    n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
    n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
    n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
    n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
    n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
    n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
    n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
    n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
    n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
    n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
    n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
    n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
    n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
    n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
    n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
    n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
    n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
    n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
    n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
    n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
    n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
    n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
    n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
    n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
    n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
    n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
    n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
    n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
    n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
    n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
    n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
    n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
    n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
    n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
    n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
    n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
    n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
    n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
    n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
    n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
    n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
    n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
    n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
    n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
    n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
    n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
    n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
    n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
    n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
    n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
    n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
    n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
    n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
    n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
    n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
    n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
    n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
    n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
    n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
    n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
    n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
    n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
    n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
    n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
    n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
    n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
    n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
    n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
    n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
    n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
    n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
    n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
    n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
    n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
    n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
    n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
    n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756,
    n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
    n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
    n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
    n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
    n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
    n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
    n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826,
    n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836,
    n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
    n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
    n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
    n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
    n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
    n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896,
    n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906,
    n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916,
    n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926,
    n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936,
    n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946,
    n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
    n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966,
    n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976,
    n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986,
    n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996,
    n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006,
    n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016,
    n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
    n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036,
    n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046,
    n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056,
    n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066,
    n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076,
    n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086,
    n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
    n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
    n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
    n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
    n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
    n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
    n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
    n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
    n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176,
    n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
    n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
    n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
    n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216,
    n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226,
    n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236,
    n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246,
    n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256,
    n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266,
    n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276,
    n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286,
    n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296,
    n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306,
    n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316,
    n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326,
    n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336,
    n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
    n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356,
    n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366,
    n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
    n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386,
    n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396,
    n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406,
    n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416,
    n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426,
    n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436,
    n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
    n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
    n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
    n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
    n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
    n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
    n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
    n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
    n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
    n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
    n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
    n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
    n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
    n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
    n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
    n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
    n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
    n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
    n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
    n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
    n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
    n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
    n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
    n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
    n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
    n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
    n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
    n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
    n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
    n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
    n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
    n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
    n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
    n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
    n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
    n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
    n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
    n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
    n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
    n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
    n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
    n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
    n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
    n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
    n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
    n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
    n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
    n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
    n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
    n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
    n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
    n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
    n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
    n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
    n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
    n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
    n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
    n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
    n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
    n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
    n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
    n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
    n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
    n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
    n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
    n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
    n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
    n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
    n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
    n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
    n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
    n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
    n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
    n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
    n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
    n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
    n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
    n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
    n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,
    n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
    n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
    n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
    n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,
    n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,
    n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
    n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,
    n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
    n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
    n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
    n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
    n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
    n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
    n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
    n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,
    n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
    n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
    n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406,
    n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416,
    n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426,
    n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436,
    n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446,
    n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456,
    n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466,
    n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476,
    n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486,
    n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496,
    n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506,
    n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516,
    n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
    n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536,
    n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546,
    n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556,
    n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566,
    n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576,
    n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586,
    n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596,
    n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606,
    n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616,
    n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626,
    n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636,
    n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646,
    n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656,
    n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666,
    n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676,
    n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686,
    n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696,
    n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706,
    n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716,
    n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726,
    n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736,
    n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746,
    n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756,
    n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766,
    n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776,
    n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786,
    n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796,
    n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806,
    n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816,
    n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826,
    n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836,
    n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846,
    n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856,
    n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866,
    n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876,
    n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886,
    n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896,
    n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906,
    n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916,
    n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926,
    n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936,
    n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946,
    n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956,
    n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966,
    n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976,
    n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986,
    n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996,
    n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006,
    n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016,
    n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026,
    n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036,
    n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046,
    n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056,
    n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066,
    n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076,
    n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086,
    n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096,
    n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106,
    n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116,
    n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126,
    n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136,
    n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146,
    n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156,
    n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166,
    n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176,
    n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186,
    n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196,
    n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206,
    n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216,
    n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226,
    n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236,
    n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246,
    n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256,
    n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266,
    n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276,
    n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286,
    n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296,
    n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306,
    n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316,
    n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326,
    n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336,
    n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346,
    n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356,
    n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366,
    n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376,
    n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386,
    n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396,
    n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406,
    n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416,
    n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426,
    n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436,
    n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446,
    n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456,
    n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466,
    n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476,
    n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486,
    n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496,
    n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506,
    n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516,
    n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526,
    n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536,
    n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546,
    n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556,
    n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566,
    n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576,
    n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586,
    n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596,
    n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606,
    n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616,
    n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626,
    n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636,
    n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646,
    n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656,
    n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666,
    n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676,
    n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686,
    n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696,
    n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706,
    n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716,
    n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726,
    n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736,
    n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746,
    n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756,
    n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766,
    n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776,
    n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786,
    n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796,
    n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806,
    n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816,
    n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826,
    n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836,
    n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846,
    n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856,
    n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866,
    n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876,
    n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886,
    n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896,
    n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906,
    n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916,
    n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926,
    n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936,
    n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946,
    n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956,
    n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966,
    n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976,
    n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986,
    n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996,
    n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006,
    n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016,
    n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026,
    n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036,
    n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046,
    n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056,
    n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066,
    n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076,
    n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086,
    n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096,
    n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106,
    n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116,
    n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126,
    n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136,
    n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146,
    n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156,
    n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166,
    n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176,
    n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186,
    n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196,
    n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206,
    n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216,
    n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226,
    n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236,
    n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246,
    n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256,
    n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266,
    n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276,
    n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286,
    n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296,
    n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306,
    n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316,
    n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326,
    n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336,
    n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346,
    n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356,
    n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366,
    n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376,
    n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386,
    n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396,
    n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406,
    n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416,
    n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426,
    n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436,
    n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446,
    n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456,
    n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466,
    n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476,
    n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486,
    n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496,
    n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506,
    n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516,
    n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526,
    n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536,
    n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546,
    n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556,
    n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566,
    n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576,
    n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586,
    n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596,
    n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606,
    n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616,
    n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626,
    n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636,
    n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646,
    n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656,
    n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
    n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
    n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
    n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
    n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
    n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
    n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
    n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
    n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
    n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
    n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
    n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
    n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
    n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
    n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
    n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
    n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
    n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
    n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
    n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
    n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
    n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
    n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
    n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
    n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
    n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
    n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
    n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
    n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
    n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
    n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
    n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
    n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
    n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
    n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
    n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014,
    n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
    n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
    n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
    n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
    n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
    n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068,
    n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
    n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086,
    n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
    n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
    n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
    n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
    n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
    n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140,
    n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
    n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158,
    n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
    n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
    n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
    n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
    n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
    n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212,
    n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221,
    n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230,
    n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
    n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
    n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
    n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
    n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
    n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284,
    n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293,
    n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302,
    n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
    n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
    n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
    n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
    n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347,
    n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356,
    n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365,
    n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374,
    n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
    n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
    n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
    n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
    n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419,
    n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428,
    n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437,
    n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446,
    n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
    n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
    n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
    n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
    n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491,
    n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500,
    n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509,
    n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518,
    n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
    n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
    n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
    n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
    n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563,
    n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572,
    n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581,
    n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590,
    n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
    n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
    n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
    n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626,
    n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635,
    n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644,
    n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653,
    n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662,
    n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
    n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
    n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
    n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698,
    n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707,
    n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716,
    n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725,
    n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734,
    n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
    n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
    n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
    n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770,
    n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779,
    n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788,
    n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797,
    n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806,
    n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
    n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
    n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
    n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842,
    n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851,
    n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860,
    n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869,
    n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878,
    n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
    n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
    n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
    n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914,
    n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923,
    n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932,
    n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941,
    n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950,
    n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
    n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
    n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
    n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986,
    n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995,
    n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004,
    n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013,
    n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022,
    n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
    n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
    n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
    n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058,
    n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067,
    n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076,
    n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085,
    n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094,
    n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
    n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
    n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
    n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130,
    n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139,
    n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148,
    n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157,
    n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166,
    n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
    n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
    n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
    n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202,
    n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211,
    n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220,
    n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229,
    n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238,
    n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
    n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
    n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
    n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274,
    n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283,
    n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292,
    n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301,
    n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310,
    n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
    n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
    n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
    n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346,
    n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355,
    n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364,
    n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373,
    n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382,
    n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
    n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
    n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
    n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418,
    n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427,
    n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436,
    n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445,
    n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454,
    n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
    n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
    n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
    n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490,
    n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499,
    n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508,
    n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517,
    n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526,
    n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
    n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
    n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
    n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562,
    n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571,
    n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580,
    n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589,
    n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598,
    n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
    n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
    n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
    n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634,
    n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643,
    n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652,
    n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661,
    n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670,
    n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
    n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
    n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
    n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706,
    n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715,
    n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724,
    n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733,
    n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742,
    n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
    n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
    n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
    n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778,
    n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787,
    n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796,
    n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805,
    n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814,
    n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
    n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
    n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
    n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850,
    n11851, n11852, n11853, n11854, n11855, n11856, n11857;
  assign n97 = reg_i_StoB_REQ0_out & reg_controllable_BtoS_ACK0_out;
  assign n98 = ~reg_controllable_BtoS_ACK1_out & n97;
  assign n99 = ~reg_controllable_BtoS_ACK1_out & ~n98;
  assign n100 = reg_i_StoB_REQ1_out & ~n99;
  assign n101 = ~reg_i_StoB_REQ1_out & n97;
  assign n102 = ~n100 & ~n101;
  assign n103 = sys_fair0done_out & ~n102;
  assign n104 = ~reg_i_StoB_REQ0_out & ~reg_controllable_BtoS_ACK0_out;
  assign n105 = ~reg_i_StoB_REQ0_out & ~n104;
  assign n106 = ~reg_controllable_BtoS_ACK1_out & ~n105;
  assign n107 = ~reg_controllable_BtoS_ACK1_out & ~n106;
  assign n108 = reg_i_StoB_REQ1_out & ~n107;
  assign n109 = ~reg_i_StoB_REQ1_out & ~n105;
  assign n110 = ~n108 & ~n109;
  assign n111 = ~sys_fair0done_out & ~n110;
  assign n112 = ~n103 & ~n111;
  assign n113 = sys_fair1done_out & ~n112;
  assign n114 = reg_controllable_BtoS_ACK1_out & n97;
  assign n115 = reg_controllable_BtoS_ACK1_out & ~n114;
  assign n116 = ~reg_i_StoB_REQ1_out & ~n115;
  assign n117 = ~reg_i_StoB_REQ1_out & ~n116;
  assign n118 = sys_fair0done_out & ~n117;
  assign n119 = ~n106 & ~n114;
  assign n120 = ~reg_i_StoB_REQ1_out & ~n119;
  assign n121 = ~n108 & ~n120;
  assign n122 = ~sys_fair0done_out & ~n121;
  assign n123 = ~n118 & ~n122;
  assign n124 = ~sys_fair1done_out & ~n123;
  assign n125 = ~n113 & ~n124;
  assign n126 = sys_fair12done_out & ~n125;
  assign n127 = ~sys_fair0done_out & ~n111;
  assign n128 = sys_fair1done_out & ~n127;
  assign n129 = ~n124 & ~n128;
  assign n130 = reg_stateG12_out & ~n129;
  assign n131 = ~reg_stateG12_out & ~n102;
  assign n132 = ~n130 & ~n131;
  assign n133 = ~sys_fair12done_out & ~n132;
  assign n134 = ~n126 & ~n133;
  assign n135 = sys_fair2done_out & ~n134;
  assign n136 = sys_fair12done_out & ~n129;
  assign n137 = ~n133 & ~n136;
  assign n138 = ~sys_fair2done_out & ~n137;
  assign n139 = ~n135 & ~n138;
  assign n140 = ~reg_controllable_BtoS_ACK2_out & ~n139;
  assign n141 = ~reg_controllable_BtoS_ACK2_out & ~n140;
  assign n142 = reg_i_StoB_REQ2_out & ~n141;
  assign n143 = ~sys_fair2done_out & ~n102;
  assign n144 = ~n135 & ~n143;
  assign n145 = reg_controllable_BtoS_ACK2_out & ~n144;
  assign n146 = ~n140 & ~n145;
  assign n147 = ~reg_i_StoB_REQ2_out & ~n146;
  assign n148 = ~n142 & ~n147;
  assign n149 = sys_fair3done_out & ~n148;
  assign n150 = ~reg_controllable_BtoS_ACK2_out & ~n137;
  assign n151 = ~reg_controllable_BtoS_ACK2_out & ~n150;
  assign n152 = reg_i_StoB_REQ2_out & ~n151;
  assign n153 = sys_fair2done_out & ~n137;
  assign n154 = ~n143 & ~n153;
  assign n155 = reg_controllable_BtoS_ACK2_out & ~n154;
  assign n156 = ~n150 & ~n155;
  assign n157 = ~reg_i_StoB_REQ2_out & ~n156;
  assign n158 = ~n152 & ~n157;
  assign n159 = ~sys_fair3done_out & ~n158;
  assign n160 = ~n149 & ~n159;
  assign n161 = ~reg_controllable_BtoS_ACK3_out & ~n160;
  assign n162 = ~reg_controllable_BtoS_ACK3_out & ~n161;
  assign n163 = reg_i_StoB_REQ3_out & ~n162;
  assign n164 = ~reg_controllable_BtoS_ACK2_out & ~n102;
  assign n165 = ~reg_controllable_BtoS_ACK2_out & ~n164;
  assign n166 = reg_i_StoB_REQ2_out & ~n165;
  assign n167 = ~reg_i_StoB_REQ2_out & ~n102;
  assign n168 = ~n166 & ~n167;
  assign n169 = ~sys_fair3done_out & ~n168;
  assign n170 = ~n149 & ~n169;
  assign n171 = reg_controllable_BtoS_ACK3_out & ~n170;
  assign n172 = ~n161 & ~n171;
  assign n173 = ~reg_i_StoB_REQ3_out & ~n172;
  assign n174 = ~n163 & ~n173;
  assign n175 = ~reg_controllable_BtoS_ACK4_out & ~n174;
  assign n176 = ~reg_controllable_BtoS_ACK4_out & ~n175;
  assign n177 = reg_i_StoB_REQ4_out & ~n176;
  assign n178 = ~reg_i_StoB_REQ4_out & ~n174;
  assign n179 = ~n177 & ~n178;
  assign n180 = sys_fair4done_out & ~n179;
  assign n181 = ~reg_controllable_BtoS_ACK3_out & ~n158;
  assign n182 = ~reg_controllable_BtoS_ACK3_out & ~n181;
  assign n183 = reg_i_StoB_REQ3_out & ~n182;
  assign n184 = sys_fair3done_out & ~n158;
  assign n185 = ~n169 & ~n184;
  assign n186 = reg_controllable_BtoS_ACK3_out & ~n185;
  assign n187 = ~n181 & ~n186;
  assign n188 = ~reg_i_StoB_REQ3_out & ~n187;
  assign n189 = ~n183 & ~n188;
  assign n190 = ~reg_controllable_BtoS_ACK4_out & ~n189;
  assign n191 = ~reg_controllable_BtoS_ACK4_out & ~n190;
  assign n192 = reg_i_StoB_REQ4_out & ~n191;
  assign n193 = ~reg_controllable_BtoS_ACK3_out & ~n168;
  assign n194 = ~reg_controllable_BtoS_ACK3_out & ~n193;
  assign n195 = reg_i_StoB_REQ3_out & ~n194;
  assign n196 = ~reg_i_StoB_REQ3_out & ~n168;
  assign n197 = ~n195 & ~n196;
  assign n198 = reg_controllable_BtoS_ACK4_out & ~n197;
  assign n199 = ~n190 & ~n198;
  assign n200 = ~reg_i_StoB_REQ4_out & ~n199;
  assign n201 = ~n192 & ~n200;
  assign n202 = ~sys_fair4done_out & ~n201;
  assign n203 = ~n180 & ~n202;
  assign n204 = ~reg_controllable_BtoS_ACK5_out & ~n203;
  assign n205 = ~reg_controllable_BtoS_ACK5_out & ~n204;
  assign n206 = reg_i_StoB_REQ5_out & ~n205;
  assign n207 = ~reg_i_StoB_REQ5_out & ~n203;
  assign n208 = ~n206 & ~n207;
  assign n209 = sys_fair5done_out & ~n208;
  assign n210 = ~reg_i_StoB_REQ4_out & ~n189;
  assign n211 = ~n192 & ~n210;
  assign n212 = sys_fair4done_out & ~n211;
  assign n213 = ~n202 & ~n212;
  assign n214 = ~reg_controllable_BtoS_ACK5_out & ~n213;
  assign n215 = ~reg_controllable_BtoS_ACK5_out & ~n214;
  assign n216 = reg_i_StoB_REQ5_out & ~n215;
  assign n217 = ~reg_controllable_BtoS_ACK4_out & ~n197;
  assign n218 = ~reg_controllable_BtoS_ACK4_out & ~n217;
  assign n219 = reg_i_StoB_REQ4_out & ~n218;
  assign n220 = ~reg_i_StoB_REQ4_out & ~n197;
  assign n221 = ~n219 & ~n220;
  assign n222 = reg_controllable_BtoS_ACK5_out & ~n221;
  assign n223 = ~n214 & ~n222;
  assign n224 = ~reg_i_StoB_REQ5_out & ~n223;
  assign n225 = ~n216 & ~n224;
  assign n226 = ~sys_fair5done_out & ~n225;
  assign n227 = ~n209 & ~n226;
  assign n228 = ~reg_controllable_BtoS_ACK6_out & ~n227;
  assign n229 = ~reg_controllable_BtoS_ACK6_out & ~n228;
  assign n230 = reg_i_StoB_REQ6_out & ~n229;
  assign n231 = ~reg_i_StoB_REQ6_out & ~n227;
  assign n232 = ~n230 & ~n231;
  assign n233 = sys_fair6done_out & ~n232;
  assign n234 = ~reg_i_StoB_REQ5_out & ~n213;
  assign n235 = ~n216 & ~n234;
  assign n236 = sys_fair5done_out & ~n235;
  assign n237 = ~n226 & ~n236;
  assign n238 = ~reg_controllable_BtoS_ACK6_out & ~n237;
  assign n239 = ~reg_controllable_BtoS_ACK6_out & ~n238;
  assign n240 = reg_i_StoB_REQ6_out & ~n239;
  assign n241 = ~reg_controllable_BtoS_ACK5_out & ~n221;
  assign n242 = ~reg_controllable_BtoS_ACK5_out & ~n241;
  assign n243 = reg_i_StoB_REQ5_out & ~n242;
  assign n244 = ~reg_i_StoB_REQ5_out & ~n221;
  assign n245 = ~n243 & ~n244;
  assign n246 = reg_controllable_BtoS_ACK6_out & ~n245;
  assign n247 = ~n238 & ~n246;
  assign n248 = ~reg_i_StoB_REQ6_out & ~n247;
  assign n249 = ~n240 & ~n248;
  assign n250 = ~sys_fair6done_out & ~n249;
  assign n251 = ~n233 & ~n250;
  assign n252 = ~reg_controllable_BtoS_ACK7_out & ~n251;
  assign n253 = ~reg_controllable_BtoS_ACK7_out & ~n252;
  assign n254 = reg_i_StoB_REQ7_out & ~n253;
  assign n255 = ~reg_i_StoB_REQ7_out & ~n251;
  assign n256 = ~n254 & ~n255;
  assign n257 = sys_fair7done_out & ~n256;
  assign n258 = ~reg_i_StoB_REQ6_out & ~n237;
  assign n259 = ~n240 & ~n258;
  assign n260 = sys_fair6done_out & ~n259;
  assign n261 = ~n250 & ~n260;
  assign n262 = ~reg_controllable_BtoS_ACK7_out & ~n261;
  assign n263 = ~reg_controllable_BtoS_ACK7_out & ~n262;
  assign n264 = reg_i_StoB_REQ7_out & ~n263;
  assign n265 = ~reg_controllable_BtoS_ACK6_out & ~n245;
  assign n266 = ~reg_controllable_BtoS_ACK6_out & ~n265;
  assign n267 = reg_i_StoB_REQ6_out & ~n266;
  assign n268 = ~reg_i_StoB_REQ6_out & ~n245;
  assign n269 = ~n267 & ~n268;
  assign n270 = reg_controllable_BtoS_ACK7_out & ~n269;
  assign n271 = ~n262 & ~n270;
  assign n272 = ~reg_i_StoB_REQ7_out & ~n271;
  assign n273 = ~n264 & ~n272;
  assign n274 = ~sys_fair7done_out & ~n273;
  assign n275 = ~n257 & ~n274;
  assign n276 = sys_fair8done_out & ~n275;
  assign n277 = ~reg_i_StoB_REQ7_out & ~n261;
  assign n278 = ~n264 & ~n277;
  assign n279 = sys_fair7done_out & ~n278;
  assign n280 = ~n274 & ~n279;
  assign n281 = ~sys_fair8done_out & ~n280;
  assign n282 = ~n276 & ~n281;
  assign n283 = ~reg_controllable_BtoS_ACK8_out & ~n282;
  assign n284 = ~reg_controllable_BtoS_ACK8_out & ~n283;
  assign n285 = reg_i_StoB_REQ8_out & ~n284;
  assign n286 = ~reg_controllable_BtoS_ACK7_out & ~n269;
  assign n287 = ~reg_controllable_BtoS_ACK7_out & ~n286;
  assign n288 = reg_i_StoB_REQ7_out & ~n287;
  assign n289 = ~reg_i_StoB_REQ7_out & ~n269;
  assign n290 = ~n288 & ~n289;
  assign n291 = ~sys_fair8done_out & ~n290;
  assign n292 = ~n276 & ~n291;
  assign n293 = reg_controllable_BtoS_ACK8_out & ~n292;
  assign n294 = ~n283 & ~n293;
  assign n295 = ~reg_i_StoB_REQ8_out & ~n294;
  assign n296 = ~n285 & ~n295;
  assign n297 = ~reg_controllable_BtoS_ACK10_out & ~n296;
  assign n298 = ~reg_controllable_BtoS_ACK10_out & ~n297;
  assign n299 = reg_i_StoB_REQ10_out & ~n298;
  assign n300 = ~reg_i_StoB_REQ10_out & ~n296;
  assign n301 = ~n299 & ~n300;
  assign n302 = sys_fair10done_out & ~n301;
  assign n303 = ~reg_controllable_BtoS_ACK8_out & ~n280;
  assign n304 = ~reg_controllable_BtoS_ACK8_out & ~n303;
  assign n305 = reg_i_StoB_REQ8_out & ~n304;
  assign n306 = sys_fair8done_out & ~n280;
  assign n307 = ~n291 & ~n306;
  assign n308 = reg_controllable_BtoS_ACK8_out & ~n307;
  assign n309 = ~n303 & ~n308;
  assign n310 = ~reg_i_StoB_REQ8_out & ~n309;
  assign n311 = ~n305 & ~n310;
  assign n312 = ~reg_controllable_BtoS_ACK10_out & ~n311;
  assign n313 = ~reg_controllable_BtoS_ACK10_out & ~n312;
  assign n314 = reg_i_StoB_REQ10_out & ~n313;
  assign n315 = ~reg_controllable_BtoS_ACK8_out & ~n290;
  assign n316 = ~reg_controllable_BtoS_ACK8_out & ~n315;
  assign n317 = reg_i_StoB_REQ8_out & ~n316;
  assign n318 = ~reg_i_StoB_REQ8_out & ~n290;
  assign n319 = ~n317 & ~n318;
  assign n320 = reg_controllable_BtoS_ACK10_out & ~n319;
  assign n321 = ~n312 & ~n320;
  assign n322 = ~reg_i_StoB_REQ10_out & ~n321;
  assign n323 = ~n314 & ~n322;
  assign n324 = ~sys_fair10done_out & ~n323;
  assign n325 = ~n302 & ~n324;
  assign n326 = sys_fair11done_out & ~n325;
  assign n327 = ~reg_i_StoB_REQ10_out & ~n311;
  assign n328 = ~n314 & ~n327;
  assign n329 = sys_fair10done_out & ~n328;
  assign n330 = ~n324 & ~n329;
  assign n331 = ~sys_fair11done_out & ~n330;
  assign n332 = ~n326 & ~n331;
  assign n333 = ~reg_controllable_BtoS_ACK11_out & ~n332;
  assign n334 = ~reg_controllable_BtoS_ACK11_out & ~n333;
  assign n335 = reg_i_StoB_REQ11_out & ~n334;
  assign n336 = ~reg_controllable_BtoS_ACK10_out & ~n319;
  assign n337 = ~reg_controllable_BtoS_ACK10_out & ~n336;
  assign n338 = reg_i_StoB_REQ10_out & ~n337;
  assign n339 = ~reg_i_StoB_REQ10_out & ~n319;
  assign n340 = ~n338 & ~n339;
  assign n341 = ~sys_fair11done_out & ~n340;
  assign n342 = ~n326 & ~n341;
  assign n343 = reg_controllable_BtoS_ACK11_out & ~n342;
  assign n344 = ~n333 & ~n343;
  assign n345 = ~reg_i_StoB_REQ11_out & ~n344;
  assign n346 = ~n335 & ~n345;
  assign n347 = sys_fair9done_out & ~n346;
  assign n348 = ~reg_controllable_BtoS_ACK11_out & ~n330;
  assign n349 = ~reg_controllable_BtoS_ACK11_out & ~n348;
  assign n350 = reg_i_StoB_REQ11_out & ~n349;
  assign n351 = sys_fair11done_out & ~n330;
  assign n352 = ~n341 & ~n351;
  assign n353 = reg_controllable_BtoS_ACK11_out & ~n352;
  assign n354 = ~n348 & ~n353;
  assign n355 = ~reg_i_StoB_REQ11_out & ~n354;
  assign n356 = ~n350 & ~n355;
  assign n357 = ~sys_fair9done_out & ~n356;
  assign n358 = ~n347 & ~n357;
  assign n359 = fair_cnt<1>_out  & ~n358;
  assign n360 = ~reg_controllable_BtoS_ACK11_out & ~n340;
  assign n361 = ~reg_controllable_BtoS_ACK11_out & ~n360;
  assign n362 = reg_i_StoB_REQ11_out & ~n361;
  assign n363 = ~reg_i_StoB_REQ11_out & ~n340;
  assign n364 = ~n362 & ~n363;
  assign n365 = ~fair_cnt<1>_out  & ~n364;
  assign n366 = ~n359 & ~n365;
  assign n367 = fair_cnt<0>_out  & ~n366;
  assign n368 = ~fair_cnt<0>_out  & ~n364;
  assign n369 = ~n367 & ~n368;
  assign n370 = ~reg_controllable_BtoR_REQ1_out & ~n369;
  assign n371 = ~reg_controllable_BtoR_REQ1_out & ~n370;
  assign n372 = ~reg_controllable_BtoR_REQ0_out & ~n371;
  assign n373 = ~reg_controllable_BtoR_REQ0_out & ~n372;
  assign n374 = reg_i_RtoB_ACK1_out & ~n373;
  assign n375 = env_fair1done_out & ~n369;
  assign n376 = sys_fair12done_out & ~n102;
  assign n377 = reg_i_StoB_REQ0_out & ~n97;
  assign n378 = ~reg_i_StoB_REQ1_out & ~n377;
  assign n379 = ~n100 & ~n378;
  assign n380 = sys_fair0done_out & ~n379;
  assign n381 = ~sys_fair0done_out & ~n102;
  assign n382 = ~n380 & ~n381;
  assign n383 = sys_fair1done_out & ~n382;
  assign n384 = ~sys_fair1done_out & ~n102;
  assign n385 = ~n383 & ~n384;
  assign n386 = reg_stateG12_out & ~n385;
  assign n387 = ~n131 & ~n386;
  assign n388 = ~sys_fair12done_out & ~n387;
  assign n389 = ~n376 & ~n388;
  assign n390 = sys_fair2done_out & ~n389;
  assign n391 = ~n143 & ~n390;
  assign n392 = ~reg_i_StoB_REQ2_out & ~n391;
  assign n393 = ~n166 & ~n392;
  assign n394 = sys_fair3done_out & ~n393;
  assign n395 = ~n169 & ~n394;
  assign n396 = ~reg_i_StoB_REQ3_out & ~n395;
  assign n397 = ~n195 & ~n396;
  assign n398 = ~reg_i_StoB_REQ4_out & ~n397;
  assign n399 = ~n219 & ~n398;
  assign n400 = sys_fair4done_out & ~n399;
  assign n401 = ~sys_fair4done_out & ~n221;
  assign n402 = ~n400 & ~n401;
  assign n403 = ~reg_i_StoB_REQ5_out & ~n402;
  assign n404 = ~n243 & ~n403;
  assign n405 = sys_fair5done_out & ~n404;
  assign n406 = ~sys_fair5done_out & ~n245;
  assign n407 = ~n405 & ~n406;
  assign n408 = ~reg_i_StoB_REQ6_out & ~n407;
  assign n409 = ~n267 & ~n408;
  assign n410 = sys_fair6done_out & ~n409;
  assign n411 = ~sys_fair6done_out & ~n269;
  assign n412 = ~n410 & ~n411;
  assign n413 = ~reg_i_StoB_REQ7_out & ~n412;
  assign n414 = ~n288 & ~n413;
  assign n415 = sys_fair7done_out & ~n414;
  assign n416 = ~sys_fair7done_out & ~n290;
  assign n417 = ~n415 & ~n416;
  assign n418 = sys_fair8done_out & ~n417;
  assign n419 = ~n291 & ~n418;
  assign n420 = ~reg_i_StoB_REQ8_out & ~n419;
  assign n421 = ~n317 & ~n420;
  assign n422 = ~reg_i_StoB_REQ10_out & ~n421;
  assign n423 = ~n338 & ~n422;
  assign n424 = sys_fair10done_out & ~n423;
  assign n425 = ~sys_fair10done_out & ~n340;
  assign n426 = ~n424 & ~n425;
  assign n427 = sys_fair11done_out & ~n426;
  assign n428 = ~n341 & ~n427;
  assign n429 = ~reg_i_StoB_REQ11_out & ~n428;
  assign n430 = ~n362 & ~n429;
  assign n431 = sys_fair9done_out & ~n430;
  assign n432 = sys_fair12done_out & ~n385;
  assign n433 = ~n388 & ~n432;
  assign n434 = sys_fair2done_out & ~n433;
  assign n435 = ~n143 & ~n434;
  assign n436 = ~reg_i_StoB_REQ2_out & ~n435;
  assign n437 = ~n166 & ~n436;
  assign n438 = sys_fair3done_out & ~n437;
  assign n439 = ~n169 & ~n438;
  assign n440 = ~reg_i_StoB_REQ3_out & ~n439;
  assign n441 = ~n195 & ~n440;
  assign n442 = ~reg_i_StoB_REQ4_out & ~n441;
  assign n443 = ~n219 & ~n442;
  assign n444 = sys_fair4done_out & ~n443;
  assign n445 = ~n401 & ~n444;
  assign n446 = ~reg_i_StoB_REQ5_out & ~n445;
  assign n447 = ~n243 & ~n446;
  assign n448 = sys_fair5done_out & ~n447;
  assign n449 = ~n406 & ~n448;
  assign n450 = ~reg_i_StoB_REQ6_out & ~n449;
  assign n451 = ~n267 & ~n450;
  assign n452 = sys_fair6done_out & ~n451;
  assign n453 = ~n411 & ~n452;
  assign n454 = ~reg_i_StoB_REQ7_out & ~n453;
  assign n455 = ~n288 & ~n454;
  assign n456 = sys_fair7done_out & ~n455;
  assign n457 = ~n416 & ~n456;
  assign n458 = sys_fair8done_out & ~n457;
  assign n459 = ~n291 & ~n458;
  assign n460 = ~reg_i_StoB_REQ8_out & ~n459;
  assign n461 = ~n317 & ~n460;
  assign n462 = ~reg_i_StoB_REQ10_out & ~n461;
  assign n463 = ~n338 & ~n462;
  assign n464 = sys_fair10done_out & ~n463;
  assign n465 = ~n425 & ~n464;
  assign n466 = sys_fair11done_out & ~n465;
  assign n467 = ~n341 & ~n466;
  assign n468 = ~reg_i_StoB_REQ11_out & ~n467;
  assign n469 = ~n362 & ~n468;
  assign n470 = ~sys_fair9done_out & ~n469;
  assign n471 = ~n431 & ~n470;
  assign n472 = fair_cnt<1>_out  & ~n471;
  assign n473 = ~n365 & ~n472;
  assign n474 = fair_cnt<0>_out  & ~n473;
  assign n475 = ~n368 & ~n474;
  assign n476 = ~env_fair1done_out & ~n475;
  assign n477 = ~n375 & ~n476;
  assign n478 = env_fair0done_out & ~n477;
  assign n479 = ~env_fair0done_out & ~n364;
  assign n480 = ~n478 & ~n479;
  assign n481 = ~reg_stateG7_0_out & ~n480;
  assign n482 = ~reg_stateG7_0_out & ~n481;
  assign n483 = reg_nstateG7_1_out & ~n482;
  assign n484 = ~reg_nstateG7_1_out & ~n480;
  assign n485 = ~n483 & ~n484;
  assign n486 = ~reg_controllable_BtoR_REQ1_out & ~n485;
  assign n487 = ~reg_controllable_BtoR_REQ1_out & ~n486;
  assign n488 = reg_controllable_BtoR_REQ0_out & ~n487;
  assign n489 = reg_i_StoB_REQ1_out & ~n108;
  assign n490 = ~sys_fair0done_out & ~n489;
  assign n491 = ~n380 & ~n490;
  assign n492 = sys_fair1done_out & ~n491;
  assign n493 = reg_controllable_BtoS_ACK1_out & ~n377;
  assign n494 = reg_controllable_BtoS_ACK1_out & ~n493;
  assign n495 = ~reg_i_StoB_REQ1_out & ~n494;
  assign n496 = ~reg_i_StoB_REQ1_out & ~n495;
  assign n497 = sys_fair0done_out & ~n496;
  assign n498 = ~n108 & ~n495;
  assign n499 = ~sys_fair0done_out & ~n498;
  assign n500 = ~n497 & ~n499;
  assign n501 = ~sys_fair1done_out & ~n500;
  assign n502 = ~n492 & ~n501;
  assign n503 = sys_fair12done_out & ~n502;
  assign n504 = ~sys_fair0done_out & ~n490;
  assign n505 = sys_fair1done_out & ~n504;
  assign n506 = ~n501 & ~n505;
  assign n507 = reg_stateG12_out & ~n506;
  assign n508 = ~reg_stateG12_out & ~n379;
  assign n509 = ~n507 & ~n508;
  assign n510 = ~sys_fair12done_out & ~n509;
  assign n511 = ~n503 & ~n510;
  assign n512 = sys_fair2done_out & ~n511;
  assign n513 = ~sys_fair2done_out & ~n379;
  assign n514 = ~n512 & ~n513;
  assign n515 = reg_controllable_BtoS_ACK2_out & ~n514;
  assign n516 = sys_fair12done_out & ~n506;
  assign n517 = ~n510 & ~n516;
  assign n518 = ~sys_fair2done_out & ~n517;
  assign n519 = ~n512 & ~n518;
  assign n520 = ~reg_controllable_BtoS_ACK2_out & ~n519;
  assign n521 = ~n515 & ~n520;
  assign n522 = ~reg_i_StoB_REQ2_out & ~n521;
  assign n523 = ~n142 & ~n522;
  assign n524 = sys_fair3done_out & ~n523;
  assign n525 = ~reg_i_StoB_REQ2_out & ~n379;
  assign n526 = ~n166 & ~n525;
  assign n527 = ~sys_fair3done_out & ~n526;
  assign n528 = ~n524 & ~n527;
  assign n529 = reg_controllable_BtoS_ACK3_out & ~n528;
  assign n530 = sys_fair2done_out & ~n517;
  assign n531 = ~n513 & ~n530;
  assign n532 = reg_controllable_BtoS_ACK2_out & ~n531;
  assign n533 = ~reg_controllable_BtoS_ACK2_out & ~n517;
  assign n534 = ~n532 & ~n533;
  assign n535 = ~reg_i_StoB_REQ2_out & ~n534;
  assign n536 = ~n152 & ~n535;
  assign n537 = ~sys_fair3done_out & ~n536;
  assign n538 = ~n524 & ~n537;
  assign n539 = ~reg_controllable_BtoS_ACK3_out & ~n538;
  assign n540 = ~n529 & ~n539;
  assign n541 = ~reg_i_StoB_REQ3_out & ~n540;
  assign n542 = ~n163 & ~n541;
  assign n543 = ~reg_i_StoB_REQ4_out & ~n542;
  assign n544 = ~n177 & ~n543;
  assign n545 = sys_fair4done_out & ~n544;
  assign n546 = ~reg_i_StoB_REQ3_out & ~n526;
  assign n547 = ~n195 & ~n546;
  assign n548 = reg_controllable_BtoS_ACK4_out & ~n547;
  assign n549 = sys_fair3done_out & ~n536;
  assign n550 = ~n527 & ~n549;
  assign n551 = reg_controllable_BtoS_ACK3_out & ~n550;
  assign n552 = ~reg_controllable_BtoS_ACK3_out & ~n536;
  assign n553 = ~n551 & ~n552;
  assign n554 = ~reg_i_StoB_REQ3_out & ~n553;
  assign n555 = ~n183 & ~n554;
  assign n556 = ~reg_controllable_BtoS_ACK4_out & ~n555;
  assign n557 = ~n548 & ~n556;
  assign n558 = ~reg_i_StoB_REQ4_out & ~n557;
  assign n559 = ~n192 & ~n558;
  assign n560 = ~sys_fair4done_out & ~n559;
  assign n561 = ~n545 & ~n560;
  assign n562 = ~reg_i_StoB_REQ5_out & ~n561;
  assign n563 = ~n206 & ~n562;
  assign n564 = sys_fair5done_out & ~n563;
  assign n565 = ~reg_i_StoB_REQ4_out & ~n547;
  assign n566 = ~n219 & ~n565;
  assign n567 = reg_controllable_BtoS_ACK5_out & ~n566;
  assign n568 = ~reg_i_StoB_REQ4_out & ~n555;
  assign n569 = ~n192 & ~n568;
  assign n570 = sys_fair4done_out & ~n569;
  assign n571 = ~n560 & ~n570;
  assign n572 = ~reg_controllable_BtoS_ACK5_out & ~n571;
  assign n573 = ~n567 & ~n572;
  assign n574 = ~reg_i_StoB_REQ5_out & ~n573;
  assign n575 = ~n216 & ~n574;
  assign n576 = ~sys_fair5done_out & ~n575;
  assign n577 = ~n564 & ~n576;
  assign n578 = ~reg_i_StoB_REQ6_out & ~n577;
  assign n579 = ~n230 & ~n578;
  assign n580 = sys_fair6done_out & ~n579;
  assign n581 = ~reg_i_StoB_REQ5_out & ~n566;
  assign n582 = ~n243 & ~n581;
  assign n583 = reg_controllable_BtoS_ACK6_out & ~n582;
  assign n584 = ~reg_i_StoB_REQ5_out & ~n571;
  assign n585 = ~n216 & ~n584;
  assign n586 = sys_fair5done_out & ~n585;
  assign n587 = ~n576 & ~n586;
  assign n588 = ~reg_controllable_BtoS_ACK6_out & ~n587;
  assign n589 = ~n583 & ~n588;
  assign n590 = ~reg_i_StoB_REQ6_out & ~n589;
  assign n591 = ~n240 & ~n590;
  assign n592 = ~sys_fair6done_out & ~n591;
  assign n593 = ~n580 & ~n592;
  assign n594 = ~reg_i_StoB_REQ7_out & ~n593;
  assign n595 = ~n254 & ~n594;
  assign n596 = sys_fair7done_out & ~n595;
  assign n597 = ~reg_i_StoB_REQ6_out & ~n582;
  assign n598 = ~n267 & ~n597;
  assign n599 = reg_controllable_BtoS_ACK7_out & ~n598;
  assign n600 = ~reg_i_StoB_REQ6_out & ~n587;
  assign n601 = ~n240 & ~n600;
  assign n602 = sys_fair6done_out & ~n601;
  assign n603 = ~n592 & ~n602;
  assign n604 = ~reg_controllable_BtoS_ACK7_out & ~n603;
  assign n605 = ~n599 & ~n604;
  assign n606 = ~reg_i_StoB_REQ7_out & ~n605;
  assign n607 = ~n264 & ~n606;
  assign n608 = ~sys_fair7done_out & ~n607;
  assign n609 = ~n596 & ~n608;
  assign n610 = sys_fair8done_out & ~n609;
  assign n611 = ~reg_i_StoB_REQ7_out & ~n598;
  assign n612 = ~n288 & ~n611;
  assign n613 = ~sys_fair8done_out & ~n612;
  assign n614 = ~n610 & ~n613;
  assign n615 = reg_controllable_BtoS_ACK8_out & ~n614;
  assign n616 = ~reg_i_StoB_REQ7_out & ~n603;
  assign n617 = ~n264 & ~n616;
  assign n618 = sys_fair7done_out & ~n617;
  assign n619 = ~n608 & ~n618;
  assign n620 = ~sys_fair8done_out & ~n619;
  assign n621 = ~n610 & ~n620;
  assign n622 = ~reg_controllable_BtoS_ACK8_out & ~n621;
  assign n623 = ~n615 & ~n622;
  assign n624 = ~reg_i_StoB_REQ8_out & ~n623;
  assign n625 = ~n285 & ~n624;
  assign n626 = ~reg_i_StoB_REQ10_out & ~n625;
  assign n627 = ~n299 & ~n626;
  assign n628 = sys_fair10done_out & ~n627;
  assign n629 = ~reg_i_StoB_REQ8_out & ~n612;
  assign n630 = ~n317 & ~n629;
  assign n631 = reg_controllable_BtoS_ACK10_out & ~n630;
  assign n632 = sys_fair8done_out & ~n619;
  assign n633 = ~n613 & ~n632;
  assign n634 = reg_controllable_BtoS_ACK8_out & ~n633;
  assign n635 = ~reg_controllable_BtoS_ACK8_out & ~n619;
  assign n636 = ~n634 & ~n635;
  assign n637 = ~reg_i_StoB_REQ8_out & ~n636;
  assign n638 = ~n305 & ~n637;
  assign n639 = ~reg_controllable_BtoS_ACK10_out & ~n638;
  assign n640 = ~n631 & ~n639;
  assign n641 = ~reg_i_StoB_REQ10_out & ~n640;
  assign n642 = ~n314 & ~n641;
  assign n643 = ~sys_fair10done_out & ~n642;
  assign n644 = ~n628 & ~n643;
  assign n645 = sys_fair11done_out & ~n644;
  assign n646 = ~reg_i_StoB_REQ10_out & ~n630;
  assign n647 = ~n338 & ~n646;
  assign n648 = ~sys_fair11done_out & ~n647;
  assign n649 = ~n645 & ~n648;
  assign n650 = reg_controllable_BtoS_ACK11_out & ~n649;
  assign n651 = ~reg_i_StoB_REQ10_out & ~n638;
  assign n652 = ~n314 & ~n651;
  assign n653 = sys_fair10done_out & ~n652;
  assign n654 = ~n643 & ~n653;
  assign n655 = ~sys_fair11done_out & ~n654;
  assign n656 = ~n645 & ~n655;
  assign n657 = ~reg_controllable_BtoS_ACK11_out & ~n656;
  assign n658 = ~n650 & ~n657;
  assign n659 = ~reg_i_StoB_REQ11_out & ~n658;
  assign n660 = ~n335 & ~n659;
  assign n661 = sys_fair9done_out & ~n660;
  assign n662 = sys_fair11done_out & ~n654;
  assign n663 = ~n648 & ~n662;
  assign n664 = reg_controllable_BtoS_ACK11_out & ~n663;
  assign n665 = ~reg_controllable_BtoS_ACK11_out & ~n654;
  assign n666 = ~n664 & ~n665;
  assign n667 = ~reg_i_StoB_REQ11_out & ~n666;
  assign n668 = ~n350 & ~n667;
  assign n669 = ~sys_fair9done_out & ~n668;
  assign n670 = ~n661 & ~n669;
  assign n671 = fair_cnt<1>_out  & ~n670;
  assign n672 = ~reg_i_StoB_REQ11_out & ~n647;
  assign n673 = ~n362 & ~n672;
  assign n674 = ~fair_cnt<1>_out  & ~n673;
  assign n675 = ~n671 & ~n674;
  assign n676 = fair_cnt<0>_out  & ~n675;
  assign n677 = ~fair_cnt<0>_out  & ~n673;
  assign n678 = ~n676 & ~n677;
  assign n679 = reg_nstateG7_1_out & ~n678;
  assign n680 = ~reg_stateG7_0_out & ~n678;
  assign n681 = ~reg_stateG7_0_out & ~n680;
  assign n682 = ~reg_nstateG7_1_out & ~n681;
  assign n683 = ~n679 & ~n682;
  assign n684 = reg_controllable_BtoR_REQ1_out & ~n683;
  assign n685 = reg_nstateG7_1_out & ~n477;
  assign n686 = ~reg_nstateG7_1_out & ~n369;
  assign n687 = ~n685 & ~n686;
  assign n688 = ~reg_controllable_BtoR_REQ1_out & ~n687;
  assign n689 = ~n684 & ~n688;
  assign n690 = ~reg_controllable_BtoR_REQ0_out & ~n689;
  assign n691 = ~n488 & ~n690;
  assign n692 = ~reg_i_RtoB_ACK1_out & ~n691;
  assign n693 = ~n374 & ~n692;
  assign n694 = reg_i_RtoB_ACK0_out & ~n693;
  assign n695 = reg_nstateG7_1_out & ~n681;
  assign n696 = ~reg_nstateG7_1_out & ~n678;
  assign n697 = ~n695 & ~n696;
  assign n698 = ~reg_controllable_BtoR_REQ1_out & ~n697;
  assign n699 = ~reg_controllable_BtoR_REQ1_out & ~n698;
  assign n700 = reg_controllable_BtoR_REQ0_out & ~n699;
  assign n701 = ~env_fair1done_out & ~n364;
  assign n702 = ~n375 & ~n701;
  assign n703 = env_fair0done_out & ~n702;
  assign n704 = env_fair1done_out & ~n475;
  assign n705 = ~n701 & ~n704;
  assign n706 = ~env_fair0done_out & ~n705;
  assign n707 = ~n703 & ~n706;
  assign n708 = reg_nstateG7_1_out & ~n707;
  assign n709 = ~reg_stateG7_0_out & ~n707;
  assign n710 = ~reg_stateG7_0_out & ~n709;
  assign n711 = ~reg_nstateG7_1_out & ~n710;
  assign n712 = ~n708 & ~n711;
  assign n713 = reg_controllable_BtoR_REQ1_out & ~n712;
  assign n714 = reg_nstateG7_1_out & ~n369;
  assign n715 = env_fair0done_out & ~n369;
  assign n716 = ~env_fair0done_out & ~n475;
  assign n717 = ~n715 & ~n716;
  assign n718 = ~reg_nstateG7_1_out & ~n717;
  assign n719 = ~n714 & ~n718;
  assign n720 = ~reg_controllable_BtoR_REQ1_out & ~n719;
  assign n721 = ~n713 & ~n720;
  assign n722 = ~reg_controllable_BtoR_REQ0_out & ~n721;
  assign n723 = ~n700 & ~n722;
  assign n724 = reg_i_RtoB_ACK1_out & ~n723;
  assign n725 = ~sys_fair12done_out & ~n102;
  assign n726 = ~n126 & ~n725;
  assign n727 = sys_fair2done_out & ~n726;
  assign n728 = ~n136 & ~n725;
  assign n729 = ~sys_fair2done_out & ~n728;
  assign n730 = ~n727 & ~n729;
  assign n731 = ~reg_controllable_BtoS_ACK2_out & ~n730;
  assign n732 = ~reg_controllable_BtoS_ACK2_out & ~n731;
  assign n733 = reg_i_StoB_REQ2_out & ~n732;
  assign n734 = ~n143 & ~n727;
  assign n735 = reg_controllable_BtoS_ACK2_out & ~n734;
  assign n736 = ~n731 & ~n735;
  assign n737 = ~reg_i_StoB_REQ2_out & ~n736;
  assign n738 = ~n733 & ~n737;
  assign n739 = sys_fair3done_out & ~n738;
  assign n740 = ~reg_controllable_BtoS_ACK2_out & ~n728;
  assign n741 = ~reg_controllable_BtoS_ACK2_out & ~n740;
  assign n742 = reg_i_StoB_REQ2_out & ~n741;
  assign n743 = sys_fair2done_out & ~n728;
  assign n744 = ~n143 & ~n743;
  assign n745 = reg_controllable_BtoS_ACK2_out & ~n744;
  assign n746 = ~n740 & ~n745;
  assign n747 = ~reg_i_StoB_REQ2_out & ~n746;
  assign n748 = ~n742 & ~n747;
  assign n749 = ~sys_fair3done_out & ~n748;
  assign n750 = ~n739 & ~n749;
  assign n751 = ~reg_controllable_BtoS_ACK3_out & ~n750;
  assign n752 = ~reg_controllable_BtoS_ACK3_out & ~n751;
  assign n753 = reg_i_StoB_REQ3_out & ~n752;
  assign n754 = ~n169 & ~n739;
  assign n755 = reg_controllable_BtoS_ACK3_out & ~n754;
  assign n756 = ~n751 & ~n755;
  assign n757 = ~reg_i_StoB_REQ3_out & ~n756;
  assign n758 = ~n753 & ~n757;
  assign n759 = ~reg_controllable_BtoS_ACK4_out & ~n758;
  assign n760 = ~reg_controllable_BtoS_ACK4_out & ~n759;
  assign n761 = reg_i_StoB_REQ4_out & ~n760;
  assign n762 = ~reg_i_StoB_REQ4_out & ~n758;
  assign n763 = ~n761 & ~n762;
  assign n764 = sys_fair4done_out & ~n763;
  assign n765 = ~reg_controllable_BtoS_ACK3_out & ~n748;
  assign n766 = ~reg_controllable_BtoS_ACK3_out & ~n765;
  assign n767 = reg_i_StoB_REQ3_out & ~n766;
  assign n768 = sys_fair3done_out & ~n748;
  assign n769 = ~n169 & ~n768;
  assign n770 = reg_controllable_BtoS_ACK3_out & ~n769;
  assign n771 = ~n765 & ~n770;
  assign n772 = ~reg_i_StoB_REQ3_out & ~n771;
  assign n773 = ~n767 & ~n772;
  assign n774 = ~reg_controllable_BtoS_ACK4_out & ~n773;
  assign n775 = ~reg_controllable_BtoS_ACK4_out & ~n774;
  assign n776 = reg_i_StoB_REQ4_out & ~n775;
  assign n777 = ~n198 & ~n774;
  assign n778 = ~reg_i_StoB_REQ4_out & ~n777;
  assign n779 = ~n776 & ~n778;
  assign n780 = ~sys_fair4done_out & ~n779;
  assign n781 = ~n764 & ~n780;
  assign n782 = ~reg_controllable_BtoS_ACK5_out & ~n781;
  assign n783 = ~reg_controllable_BtoS_ACK5_out & ~n782;
  assign n784 = reg_i_StoB_REQ5_out & ~n783;
  assign n785 = ~reg_i_StoB_REQ5_out & ~n781;
  assign n786 = ~n784 & ~n785;
  assign n787 = sys_fair5done_out & ~n786;
  assign n788 = ~reg_i_StoB_REQ4_out & ~n773;
  assign n789 = ~n776 & ~n788;
  assign n790 = sys_fair4done_out & ~n789;
  assign n791 = ~n780 & ~n790;
  assign n792 = ~reg_controllable_BtoS_ACK5_out & ~n791;
  assign n793 = ~reg_controllable_BtoS_ACK5_out & ~n792;
  assign n794 = reg_i_StoB_REQ5_out & ~n793;
  assign n795 = ~n222 & ~n792;
  assign n796 = ~reg_i_StoB_REQ5_out & ~n795;
  assign n797 = ~n794 & ~n796;
  assign n798 = ~sys_fair5done_out & ~n797;
  assign n799 = ~n787 & ~n798;
  assign n800 = ~reg_controllable_BtoS_ACK6_out & ~n799;
  assign n801 = ~reg_controllable_BtoS_ACK6_out & ~n800;
  assign n802 = reg_i_StoB_REQ6_out & ~n801;
  assign n803 = ~reg_i_StoB_REQ6_out & ~n799;
  assign n804 = ~n802 & ~n803;
  assign n805 = sys_fair6done_out & ~n804;
  assign n806 = ~reg_i_StoB_REQ5_out & ~n791;
  assign n807 = ~n794 & ~n806;
  assign n808 = sys_fair5done_out & ~n807;
  assign n809 = ~n798 & ~n808;
  assign n810 = ~reg_controllable_BtoS_ACK6_out & ~n809;
  assign n811 = ~reg_controllable_BtoS_ACK6_out & ~n810;
  assign n812 = reg_i_StoB_REQ6_out & ~n811;
  assign n813 = ~n246 & ~n810;
  assign n814 = ~reg_i_StoB_REQ6_out & ~n813;
  assign n815 = ~n812 & ~n814;
  assign n816 = ~sys_fair6done_out & ~n815;
  assign n817 = ~n805 & ~n816;
  assign n818 = ~reg_controllable_BtoS_ACK7_out & ~n817;
  assign n819 = ~reg_controllable_BtoS_ACK7_out & ~n818;
  assign n820 = reg_i_StoB_REQ7_out & ~n819;
  assign n821 = ~reg_i_StoB_REQ7_out & ~n817;
  assign n822 = ~n820 & ~n821;
  assign n823 = sys_fair7done_out & ~n822;
  assign n824 = ~reg_i_StoB_REQ6_out & ~n809;
  assign n825 = ~n812 & ~n824;
  assign n826 = sys_fair6done_out & ~n825;
  assign n827 = ~n816 & ~n826;
  assign n828 = ~reg_controllable_BtoS_ACK7_out & ~n827;
  assign n829 = ~reg_controllable_BtoS_ACK7_out & ~n828;
  assign n830 = reg_i_StoB_REQ7_out & ~n829;
  assign n831 = ~n270 & ~n828;
  assign n832 = ~reg_i_StoB_REQ7_out & ~n831;
  assign n833 = ~n830 & ~n832;
  assign n834 = ~sys_fair7done_out & ~n833;
  assign n835 = ~n823 & ~n834;
  assign n836 = sys_fair8done_out & ~n835;
  assign n837 = ~reg_i_StoB_REQ7_out & ~n827;
  assign n838 = ~n830 & ~n837;
  assign n839 = sys_fair7done_out & ~n838;
  assign n840 = ~n834 & ~n839;
  assign n841 = ~sys_fair8done_out & ~n840;
  assign n842 = ~n836 & ~n841;
  assign n843 = ~reg_controllable_BtoS_ACK8_out & ~n842;
  assign n844 = ~reg_controllable_BtoS_ACK8_out & ~n843;
  assign n845 = reg_i_StoB_REQ8_out & ~n844;
  assign n846 = ~n291 & ~n836;
  assign n847 = reg_controllable_BtoS_ACK8_out & ~n846;
  assign n848 = ~n843 & ~n847;
  assign n849 = ~reg_i_StoB_REQ8_out & ~n848;
  assign n850 = ~n845 & ~n849;
  assign n851 = ~reg_controllable_BtoS_ACK10_out & ~n850;
  assign n852 = ~reg_controllable_BtoS_ACK10_out & ~n851;
  assign n853 = reg_i_StoB_REQ10_out & ~n852;
  assign n854 = ~reg_i_StoB_REQ10_out & ~n850;
  assign n855 = ~n853 & ~n854;
  assign n856 = sys_fair10done_out & ~n855;
  assign n857 = ~reg_controllable_BtoS_ACK8_out & ~n840;
  assign n858 = ~reg_controllable_BtoS_ACK8_out & ~n857;
  assign n859 = reg_i_StoB_REQ8_out & ~n858;
  assign n860 = sys_fair8done_out & ~n840;
  assign n861 = ~n291 & ~n860;
  assign n862 = reg_controllable_BtoS_ACK8_out & ~n861;
  assign n863 = ~n857 & ~n862;
  assign n864 = ~reg_i_StoB_REQ8_out & ~n863;
  assign n865 = ~n859 & ~n864;
  assign n866 = ~reg_controllable_BtoS_ACK10_out & ~n865;
  assign n867 = ~reg_controllable_BtoS_ACK10_out & ~n866;
  assign n868 = reg_i_StoB_REQ10_out & ~n867;
  assign n869 = ~n320 & ~n866;
  assign n870 = ~reg_i_StoB_REQ10_out & ~n869;
  assign n871 = ~n868 & ~n870;
  assign n872 = ~sys_fair10done_out & ~n871;
  assign n873 = ~n856 & ~n872;
  assign n874 = sys_fair11done_out & ~n873;
  assign n875 = ~reg_i_StoB_REQ10_out & ~n865;
  assign n876 = ~n868 & ~n875;
  assign n877 = sys_fair10done_out & ~n876;
  assign n878 = ~n872 & ~n877;
  assign n879 = ~sys_fair11done_out & ~n878;
  assign n880 = ~n874 & ~n879;
  assign n881 = ~reg_controllable_BtoS_ACK11_out & ~n880;
  assign n882 = ~reg_controllable_BtoS_ACK11_out & ~n881;
  assign n883 = reg_i_StoB_REQ11_out & ~n882;
  assign n884 = ~n341 & ~n874;
  assign n885 = reg_controllable_BtoS_ACK11_out & ~n884;
  assign n886 = ~n881 & ~n885;
  assign n887 = ~reg_i_StoB_REQ11_out & ~n886;
  assign n888 = ~n883 & ~n887;
  assign n889 = sys_fair9done_out & ~n888;
  assign n890 = ~sys_fair9done_out & ~n364;
  assign n891 = ~n889 & ~n890;
  assign n892 = fair_cnt<1>_out  & ~n891;
  assign n893 = ~n365 & ~n892;
  assign n894 = ~fair_cnt<0>_out  & ~n893;
  assign n895 = ~n367 & ~n894;
  assign n896 = env_fair0done_out & ~n895;
  assign n897 = ~env_fair0done_out & ~n369;
  assign n898 = ~n896 & ~n897;
  assign n899 = ~reg_stateG7_0_out & ~n898;
  assign n900 = ~reg_stateG7_0_out & ~n899;
  assign n901 = reg_nstateG7_1_out & ~n900;
  assign n902 = ~reg_nstateG7_1_out & ~n898;
  assign n903 = ~n901 & ~n902;
  assign n904 = ~reg_controllable_BtoR_REQ1_out & ~n903;
  assign n905 = ~reg_controllable_BtoR_REQ1_out & ~n904;
  assign n906 = reg_controllable_BtoR_REQ0_out & ~n905;
  assign n907 = env_fair1done_out & ~n895;
  assign n908 = ~env_fair1done_out & ~n369;
  assign n909 = ~n907 & ~n908;
  assign n910 = reg_nstateG7_1_out & ~n909;
  assign n911 = ~reg_stateG7_0_out & ~n909;
  assign n912 = ~reg_stateG7_0_out & ~n911;
  assign n913 = ~reg_nstateG7_1_out & ~n912;
  assign n914 = ~n910 & ~n913;
  assign n915 = reg_controllable_BtoR_REQ1_out & ~n914;
  assign n916 = fair_cnt<0>_out  & ~n893;
  assign n917 = ~n368 & ~n916;
  assign n918 = ~env_fair1done_out & ~n917;
  assign n919 = ~n907 & ~n918;
  assign n920 = reg_nstateG7_1_out & ~n919;
  assign n921 = ~env_fair0done_out & ~n917;
  assign n922 = ~n896 & ~n921;
  assign n923 = ~reg_nstateG7_1_out & ~n922;
  assign n924 = ~n920 & ~n923;
  assign n925 = ~reg_controllable_BtoR_REQ1_out & ~n924;
  assign n926 = ~n915 & ~n925;
  assign n927 = ~reg_controllable_BtoR_REQ0_out & ~n926;
  assign n928 = ~n906 & ~n927;
  assign n929 = ~reg_i_RtoB_ACK1_out & ~n928;
  assign n930 = ~n724 & ~n929;
  assign n931 = ~reg_i_RtoB_ACK0_out & ~n930;
  assign n932 = ~n694 & ~n931;
  assign n933 = reg_i_StoB_REQ9_out & ~n932;
  assign n934 = ~n97 & ~n104;
  assign n935 = ~reg_controllable_BtoS_ACK1_out & ~n934;
  assign n936 = ~reg_controllable_BtoS_ACK1_out & ~n935;
  assign n937 = reg_i_StoB_REQ1_out & ~n936;
  assign n938 = ~reg_i_StoB_REQ1_out & ~n934;
  assign n939 = ~n937 & ~n938;
  assign n940 = ~sys_fair0done_out & ~n939;
  assign n941 = ~n103 & ~n940;
  assign n942 = sys_fair1done_out & ~n941;
  assign n943 = ~n100 & ~n116;
  assign n944 = sys_fair0done_out & ~n943;
  assign n945 = ~n114 & ~n935;
  assign n946 = ~reg_i_StoB_REQ1_out & ~n945;
  assign n947 = ~n100 & ~n946;
  assign n948 = ~sys_fair0done_out & ~n947;
  assign n949 = ~n944 & ~n948;
  assign n950 = ~sys_fair1done_out & ~n949;
  assign n951 = ~n942 & ~n950;
  assign n952 = sys_fair12done_out & ~n951;
  assign n953 = ~sys_fair0done_out & ~n940;
  assign n954 = sys_fair1done_out & ~n953;
  assign n955 = ~n950 & ~n954;
  assign n956 = reg_stateG12_out & ~n955;
  assign n957 = ~n131 & ~n956;
  assign n958 = ~sys_fair12done_out & ~n957;
  assign n959 = ~n952 & ~n958;
  assign n960 = sys_fair2done_out & ~n959;
  assign n961 = ~n143 & ~n960;
  assign n962 = ~reg_controllable_BtoS_ACK2_out & ~n961;
  assign n963 = ~reg_controllable_BtoS_ACK2_out & ~n962;
  assign n964 = reg_i_StoB_REQ2_out & ~n963;
  assign n965 = reg_controllable_BtoS_ACK2_out & ~n961;
  assign n966 = sys_fair12done_out & ~n955;
  assign n967 = ~n958 & ~n966;
  assign n968 = ~sys_fair2done_out & ~n967;
  assign n969 = ~n960 & ~n968;
  assign n970 = ~reg_controllable_BtoS_ACK2_out & ~n969;
  assign n971 = ~n965 & ~n970;
  assign n972 = ~reg_i_StoB_REQ2_out & ~n971;
  assign n973 = ~n964 & ~n972;
  assign n974 = sys_fair3done_out & ~n973;
  assign n975 = ~n169 & ~n974;
  assign n976 = ~reg_controllable_BtoS_ACK3_out & ~n975;
  assign n977 = ~reg_controllable_BtoS_ACK3_out & ~n976;
  assign n978 = reg_i_StoB_REQ3_out & ~n977;
  assign n979 = reg_controllable_BtoS_ACK3_out & ~n975;
  assign n980 = sys_fair2done_out & ~n967;
  assign n981 = ~n143 & ~n980;
  assign n982 = ~reg_controllable_BtoS_ACK2_out & ~n981;
  assign n983 = ~reg_controllable_BtoS_ACK2_out & ~n982;
  assign n984 = reg_i_StoB_REQ2_out & ~n983;
  assign n985 = reg_controllable_BtoS_ACK2_out & ~n981;
  assign n986 = ~reg_controllable_BtoS_ACK2_out & ~n967;
  assign n987 = ~n985 & ~n986;
  assign n988 = ~reg_i_StoB_REQ2_out & ~n987;
  assign n989 = ~n984 & ~n988;
  assign n990 = ~sys_fair3done_out & ~n989;
  assign n991 = ~n974 & ~n990;
  assign n992 = ~reg_controllable_BtoS_ACK3_out & ~n991;
  assign n993 = ~n979 & ~n992;
  assign n994 = ~reg_i_StoB_REQ3_out & ~n993;
  assign n995 = ~n978 & ~n994;
  assign n996 = ~reg_controllable_BtoS_ACK4_out & ~n995;
  assign n997 = ~reg_controllable_BtoS_ACK4_out & ~n996;
  assign n998 = reg_i_StoB_REQ4_out & ~n997;
  assign n999 = ~reg_i_StoB_REQ4_out & ~n995;
  assign n1000 = ~n998 & ~n999;
  assign n1001 = sys_fair4done_out & ~n1000;
  assign n1002 = sys_fair3done_out & ~n989;
  assign n1003 = ~n169 & ~n1002;
  assign n1004 = ~reg_controllable_BtoS_ACK3_out & ~n1003;
  assign n1005 = ~reg_controllable_BtoS_ACK3_out & ~n1004;
  assign n1006 = reg_i_StoB_REQ3_out & ~n1005;
  assign n1007 = reg_controllable_BtoS_ACK3_out & ~n1003;
  assign n1008 = ~reg_controllable_BtoS_ACK3_out & ~n989;
  assign n1009 = ~n1007 & ~n1008;
  assign n1010 = ~reg_i_StoB_REQ3_out & ~n1009;
  assign n1011 = ~n1006 & ~n1010;
  assign n1012 = ~reg_controllable_BtoS_ACK4_out & ~n1011;
  assign n1013 = ~n198 & ~n1012;
  assign n1014 = ~reg_i_StoB_REQ4_out & ~n1013;
  assign n1015 = ~n219 & ~n1014;
  assign n1016 = ~sys_fair4done_out & ~n1015;
  assign n1017 = ~n1001 & ~n1016;
  assign n1018 = ~reg_controllable_BtoS_ACK5_out & ~n1017;
  assign n1019 = ~reg_controllable_BtoS_ACK5_out & ~n1018;
  assign n1020 = reg_i_StoB_REQ5_out & ~n1019;
  assign n1021 = ~reg_i_StoB_REQ5_out & ~n1017;
  assign n1022 = ~n1020 & ~n1021;
  assign n1023 = sys_fair5done_out & ~n1022;
  assign n1024 = ~reg_controllable_BtoS_ACK4_out & ~n1012;
  assign n1025 = reg_i_StoB_REQ4_out & ~n1024;
  assign n1026 = ~reg_i_StoB_REQ4_out & ~n1011;
  assign n1027 = ~n1025 & ~n1026;
  assign n1028 = sys_fair4done_out & ~n1027;
  assign n1029 = ~n1016 & ~n1028;
  assign n1030 = ~reg_controllable_BtoS_ACK5_out & ~n1029;
  assign n1031 = ~n222 & ~n1030;
  assign n1032 = ~reg_i_StoB_REQ5_out & ~n1031;
  assign n1033 = ~n243 & ~n1032;
  assign n1034 = ~sys_fair5done_out & ~n1033;
  assign n1035 = ~n1023 & ~n1034;
  assign n1036 = ~reg_controllable_BtoS_ACK6_out & ~n1035;
  assign n1037 = ~reg_controllable_BtoS_ACK6_out & ~n1036;
  assign n1038 = reg_i_StoB_REQ6_out & ~n1037;
  assign n1039 = ~reg_i_StoB_REQ6_out & ~n1035;
  assign n1040 = ~n1038 & ~n1039;
  assign n1041 = sys_fair6done_out & ~n1040;
  assign n1042 = ~reg_controllable_BtoS_ACK5_out & ~n1030;
  assign n1043 = reg_i_StoB_REQ5_out & ~n1042;
  assign n1044 = ~reg_i_StoB_REQ5_out & ~n1029;
  assign n1045 = ~n1043 & ~n1044;
  assign n1046 = sys_fair5done_out & ~n1045;
  assign n1047 = ~n1034 & ~n1046;
  assign n1048 = ~reg_controllable_BtoS_ACK6_out & ~n1047;
  assign n1049 = ~n246 & ~n1048;
  assign n1050 = ~reg_i_StoB_REQ6_out & ~n1049;
  assign n1051 = ~n267 & ~n1050;
  assign n1052 = ~sys_fair6done_out & ~n1051;
  assign n1053 = ~n1041 & ~n1052;
  assign n1054 = ~reg_controllable_BtoS_ACK7_out & ~n1053;
  assign n1055 = ~reg_controllable_BtoS_ACK7_out & ~n1054;
  assign n1056 = reg_i_StoB_REQ7_out & ~n1055;
  assign n1057 = ~reg_i_StoB_REQ7_out & ~n1053;
  assign n1058 = ~n1056 & ~n1057;
  assign n1059 = sys_fair7done_out & ~n1058;
  assign n1060 = ~reg_controllable_BtoS_ACK6_out & ~n1048;
  assign n1061 = reg_i_StoB_REQ6_out & ~n1060;
  assign n1062 = ~reg_i_StoB_REQ6_out & ~n1047;
  assign n1063 = ~n1061 & ~n1062;
  assign n1064 = sys_fair6done_out & ~n1063;
  assign n1065 = ~n1052 & ~n1064;
  assign n1066 = ~reg_controllable_BtoS_ACK7_out & ~n1065;
  assign n1067 = ~n270 & ~n1066;
  assign n1068 = ~reg_i_StoB_REQ7_out & ~n1067;
  assign n1069 = ~n288 & ~n1068;
  assign n1070 = ~sys_fair7done_out & ~n1069;
  assign n1071 = ~n1059 & ~n1070;
  assign n1072 = sys_fair8done_out & ~n1071;
  assign n1073 = ~n291 & ~n1072;
  assign n1074 = ~reg_controllable_BtoS_ACK8_out & ~n1073;
  assign n1075 = ~reg_controllable_BtoS_ACK8_out & ~n1074;
  assign n1076 = reg_i_StoB_REQ8_out & ~n1075;
  assign n1077 = reg_controllable_BtoS_ACK8_out & ~n1073;
  assign n1078 = ~reg_controllable_BtoS_ACK7_out & ~n1066;
  assign n1079 = reg_i_StoB_REQ7_out & ~n1078;
  assign n1080 = ~reg_i_StoB_REQ7_out & ~n1065;
  assign n1081 = ~n1079 & ~n1080;
  assign n1082 = sys_fair7done_out & ~n1081;
  assign n1083 = ~n1070 & ~n1082;
  assign n1084 = ~sys_fair8done_out & ~n1083;
  assign n1085 = ~n1072 & ~n1084;
  assign n1086 = ~reg_controllable_BtoS_ACK8_out & ~n1085;
  assign n1087 = ~n1077 & ~n1086;
  assign n1088 = ~reg_i_StoB_REQ8_out & ~n1087;
  assign n1089 = ~n1076 & ~n1088;
  assign n1090 = ~reg_controllable_BtoS_ACK10_out & ~n1089;
  assign n1091 = ~reg_controllable_BtoS_ACK10_out & ~n1090;
  assign n1092 = reg_i_StoB_REQ10_out & ~n1091;
  assign n1093 = ~reg_i_StoB_REQ10_out & ~n1089;
  assign n1094 = ~n1092 & ~n1093;
  assign n1095 = sys_fair10done_out & ~n1094;
  assign n1096 = sys_fair8done_out & ~n1083;
  assign n1097 = ~n291 & ~n1096;
  assign n1098 = ~reg_controllable_BtoS_ACK8_out & ~n1097;
  assign n1099 = ~reg_controllable_BtoS_ACK8_out & ~n1098;
  assign n1100 = reg_i_StoB_REQ8_out & ~n1099;
  assign n1101 = reg_controllable_BtoS_ACK8_out & ~n1097;
  assign n1102 = ~reg_controllable_BtoS_ACK8_out & ~n1083;
  assign n1103 = ~n1101 & ~n1102;
  assign n1104 = ~reg_i_StoB_REQ8_out & ~n1103;
  assign n1105 = ~n1100 & ~n1104;
  assign n1106 = ~reg_controllable_BtoS_ACK10_out & ~n1105;
  assign n1107 = ~n320 & ~n1106;
  assign n1108 = ~reg_i_StoB_REQ10_out & ~n1107;
  assign n1109 = ~n338 & ~n1108;
  assign n1110 = ~sys_fair10done_out & ~n1109;
  assign n1111 = ~n1095 & ~n1110;
  assign n1112 = sys_fair11done_out & ~n1111;
  assign n1113 = ~n341 & ~n1112;
  assign n1114 = ~reg_controllable_BtoS_ACK11_out & ~n1113;
  assign n1115 = ~reg_controllable_BtoS_ACK11_out & ~n1114;
  assign n1116 = reg_i_StoB_REQ11_out & ~n1115;
  assign n1117 = ~n378 & ~n937;
  assign n1118 = ~sys_fair0done_out & ~n1117;
  assign n1119 = ~n380 & ~n1118;
  assign n1120 = sys_fair1done_out & ~n1119;
  assign n1121 = ~n100 & ~n495;
  assign n1122 = sys_fair0done_out & ~n1121;
  assign n1123 = ~sys_fair0done_out & ~n379;
  assign n1124 = ~n1122 & ~n1123;
  assign n1125 = ~sys_fair1done_out & ~n1124;
  assign n1126 = ~n1120 & ~n1125;
  assign n1127 = sys_fair12done_out & ~n1126;
  assign n1128 = ~sys_fair0done_out & ~n1118;
  assign n1129 = sys_fair1done_out & ~n1128;
  assign n1130 = ~n1125 & ~n1129;
  assign n1131 = reg_stateG12_out & ~n1130;
  assign n1132 = ~n508 & ~n1131;
  assign n1133 = ~sys_fair12done_out & ~n1132;
  assign n1134 = ~n1127 & ~n1133;
  assign n1135 = sys_fair2done_out & ~n1134;
  assign n1136 = ~n513 & ~n1135;
  assign n1137 = reg_controllable_BtoS_ACK2_out & ~n1136;
  assign n1138 = sys_fair12done_out & ~n1130;
  assign n1139 = ~n1133 & ~n1138;
  assign n1140 = ~sys_fair2done_out & ~n1139;
  assign n1141 = ~n1135 & ~n1140;
  assign n1142 = ~reg_controllable_BtoS_ACK2_out & ~n1141;
  assign n1143 = ~n1137 & ~n1142;
  assign n1144 = ~reg_i_StoB_REQ2_out & ~n1143;
  assign n1145 = ~n964 & ~n1144;
  assign n1146 = sys_fair3done_out & ~n1145;
  assign n1147 = ~n527 & ~n1146;
  assign n1148 = reg_controllable_BtoS_ACK3_out & ~n1147;
  assign n1149 = sys_fair2done_out & ~n1139;
  assign n1150 = ~n513 & ~n1149;
  assign n1151 = reg_controllable_BtoS_ACK2_out & ~n1150;
  assign n1152 = ~reg_controllable_BtoS_ACK2_out & ~n1139;
  assign n1153 = ~n1151 & ~n1152;
  assign n1154 = ~reg_i_StoB_REQ2_out & ~n1153;
  assign n1155 = ~n984 & ~n1154;
  assign n1156 = ~sys_fair3done_out & ~n1155;
  assign n1157 = ~n1146 & ~n1156;
  assign n1158 = ~reg_controllable_BtoS_ACK3_out & ~n1157;
  assign n1159 = ~n1148 & ~n1158;
  assign n1160 = ~reg_i_StoB_REQ3_out & ~n1159;
  assign n1161 = ~n978 & ~n1160;
  assign n1162 = ~reg_i_StoB_REQ4_out & ~n1161;
  assign n1163 = ~n998 & ~n1162;
  assign n1164 = sys_fair4done_out & ~n1163;
  assign n1165 = sys_fair3done_out & ~n1155;
  assign n1166 = ~n527 & ~n1165;
  assign n1167 = reg_controllable_BtoS_ACK3_out & ~n1166;
  assign n1168 = ~reg_controllable_BtoS_ACK3_out & ~n1155;
  assign n1169 = ~n1167 & ~n1168;
  assign n1170 = ~reg_i_StoB_REQ3_out & ~n1169;
  assign n1171 = ~n1006 & ~n1170;
  assign n1172 = ~reg_controllable_BtoS_ACK4_out & ~n1171;
  assign n1173 = ~n548 & ~n1172;
  assign n1174 = ~reg_i_StoB_REQ4_out & ~n1173;
  assign n1175 = ~n219 & ~n1174;
  assign n1176 = ~sys_fair4done_out & ~n1175;
  assign n1177 = ~n1164 & ~n1176;
  assign n1178 = ~reg_i_StoB_REQ5_out & ~n1177;
  assign n1179 = ~n1020 & ~n1178;
  assign n1180 = sys_fair5done_out & ~n1179;
  assign n1181 = ~reg_i_StoB_REQ4_out & ~n1171;
  assign n1182 = ~n1025 & ~n1181;
  assign n1183 = sys_fair4done_out & ~n1182;
  assign n1184 = ~n1176 & ~n1183;
  assign n1185 = ~reg_controllable_BtoS_ACK5_out & ~n1184;
  assign n1186 = ~n567 & ~n1185;
  assign n1187 = ~reg_i_StoB_REQ5_out & ~n1186;
  assign n1188 = ~n243 & ~n1187;
  assign n1189 = ~sys_fair5done_out & ~n1188;
  assign n1190 = ~n1180 & ~n1189;
  assign n1191 = ~reg_i_StoB_REQ6_out & ~n1190;
  assign n1192 = ~n1038 & ~n1191;
  assign n1193 = sys_fair6done_out & ~n1192;
  assign n1194 = ~reg_i_StoB_REQ5_out & ~n1184;
  assign n1195 = ~n1043 & ~n1194;
  assign n1196 = sys_fair5done_out & ~n1195;
  assign n1197 = ~n1189 & ~n1196;
  assign n1198 = ~reg_controllable_BtoS_ACK6_out & ~n1197;
  assign n1199 = ~n583 & ~n1198;
  assign n1200 = ~reg_i_StoB_REQ6_out & ~n1199;
  assign n1201 = ~n267 & ~n1200;
  assign n1202 = ~sys_fair6done_out & ~n1201;
  assign n1203 = ~n1193 & ~n1202;
  assign n1204 = ~reg_i_StoB_REQ7_out & ~n1203;
  assign n1205 = ~n1056 & ~n1204;
  assign n1206 = sys_fair7done_out & ~n1205;
  assign n1207 = ~reg_i_StoB_REQ6_out & ~n1197;
  assign n1208 = ~n1061 & ~n1207;
  assign n1209 = sys_fair6done_out & ~n1208;
  assign n1210 = ~n1202 & ~n1209;
  assign n1211 = ~reg_controllable_BtoS_ACK7_out & ~n1210;
  assign n1212 = ~n599 & ~n1211;
  assign n1213 = ~reg_i_StoB_REQ7_out & ~n1212;
  assign n1214 = ~n288 & ~n1213;
  assign n1215 = ~sys_fair7done_out & ~n1214;
  assign n1216 = ~n1206 & ~n1215;
  assign n1217 = sys_fair8done_out & ~n1216;
  assign n1218 = ~n613 & ~n1217;
  assign n1219 = reg_controllable_BtoS_ACK8_out & ~n1218;
  assign n1220 = ~reg_i_StoB_REQ7_out & ~n1210;
  assign n1221 = ~n1079 & ~n1220;
  assign n1222 = sys_fair7done_out & ~n1221;
  assign n1223 = ~n1215 & ~n1222;
  assign n1224 = ~sys_fair8done_out & ~n1223;
  assign n1225 = ~n1217 & ~n1224;
  assign n1226 = ~reg_controllable_BtoS_ACK8_out & ~n1225;
  assign n1227 = ~n1219 & ~n1226;
  assign n1228 = ~reg_i_StoB_REQ8_out & ~n1227;
  assign n1229 = ~n1076 & ~n1228;
  assign n1230 = ~reg_i_StoB_REQ10_out & ~n1229;
  assign n1231 = ~n1092 & ~n1230;
  assign n1232 = sys_fair10done_out & ~n1231;
  assign n1233 = sys_fair8done_out & ~n1223;
  assign n1234 = ~n613 & ~n1233;
  assign n1235 = reg_controllable_BtoS_ACK8_out & ~n1234;
  assign n1236 = ~reg_controllable_BtoS_ACK8_out & ~n1223;
  assign n1237 = ~n1235 & ~n1236;
  assign n1238 = ~reg_i_StoB_REQ8_out & ~n1237;
  assign n1239 = ~n1100 & ~n1238;
  assign n1240 = ~reg_controllable_BtoS_ACK10_out & ~n1239;
  assign n1241 = ~n631 & ~n1240;
  assign n1242 = ~reg_i_StoB_REQ10_out & ~n1241;
  assign n1243 = ~n338 & ~n1242;
  assign n1244 = ~sys_fair10done_out & ~n1243;
  assign n1245 = ~n1232 & ~n1244;
  assign n1246 = sys_fair11done_out & ~n1245;
  assign n1247 = ~n648 & ~n1246;
  assign n1248 = reg_controllable_BtoS_ACK11_out & ~n1247;
  assign n1249 = ~reg_controllable_BtoS_ACK10_out & ~n1106;
  assign n1250 = reg_i_StoB_REQ10_out & ~n1249;
  assign n1251 = ~reg_i_StoB_REQ10_out & ~n1239;
  assign n1252 = ~n1250 & ~n1251;
  assign n1253 = sys_fair10done_out & ~n1252;
  assign n1254 = ~n1244 & ~n1253;
  assign n1255 = ~sys_fair11done_out & ~n1254;
  assign n1256 = ~n1246 & ~n1255;
  assign n1257 = ~reg_controllable_BtoS_ACK11_out & ~n1256;
  assign n1258 = ~n1248 & ~n1257;
  assign n1259 = ~reg_i_StoB_REQ11_out & ~n1258;
  assign n1260 = ~n1116 & ~n1259;
  assign n1261 = sys_fair9done_out & ~n1260;
  assign n1262 = ~sys_fair9done_out & ~n673;
  assign n1263 = ~n1261 & ~n1262;
  assign n1264 = fair_cnt<1>_out  & ~n1263;
  assign n1265 = ~n674 & ~n1264;
  assign n1266 = fair_cnt<0>_out  & ~n1265;
  assign n1267 = ~n677 & ~n1266;
  assign n1268 = env_fair0done_out & ~n1267;
  assign n1269 = ~n725 & ~n952;
  assign n1270 = sys_fair2done_out & ~n1269;
  assign n1271 = ~n143 & ~n1270;
  assign n1272 = ~reg_controllable_BtoS_ACK2_out & ~n1271;
  assign n1273 = ~reg_controllable_BtoS_ACK2_out & ~n1272;
  assign n1274 = reg_i_StoB_REQ2_out & ~n1273;
  assign n1275 = reg_controllable_BtoS_ACK2_out & ~n1271;
  assign n1276 = ~n725 & ~n966;
  assign n1277 = ~sys_fair2done_out & ~n1276;
  assign n1278 = ~n1270 & ~n1277;
  assign n1279 = ~reg_controllable_BtoS_ACK2_out & ~n1278;
  assign n1280 = ~n1275 & ~n1279;
  assign n1281 = ~reg_i_StoB_REQ2_out & ~n1280;
  assign n1282 = ~n1274 & ~n1281;
  assign n1283 = sys_fair3done_out & ~n1282;
  assign n1284 = ~n169 & ~n1283;
  assign n1285 = ~reg_controllable_BtoS_ACK3_out & ~n1284;
  assign n1286 = ~reg_controllable_BtoS_ACK3_out & ~n1285;
  assign n1287 = reg_i_StoB_REQ3_out & ~n1286;
  assign n1288 = reg_controllable_BtoS_ACK3_out & ~n1284;
  assign n1289 = sys_fair2done_out & ~n1276;
  assign n1290 = ~n143 & ~n1289;
  assign n1291 = ~reg_controllable_BtoS_ACK2_out & ~n1290;
  assign n1292 = ~reg_controllable_BtoS_ACK2_out & ~n1291;
  assign n1293 = reg_i_StoB_REQ2_out & ~n1292;
  assign n1294 = reg_controllable_BtoS_ACK2_out & ~n1290;
  assign n1295 = ~reg_controllable_BtoS_ACK2_out & ~n1276;
  assign n1296 = ~n1294 & ~n1295;
  assign n1297 = ~reg_i_StoB_REQ2_out & ~n1296;
  assign n1298 = ~n1293 & ~n1297;
  assign n1299 = ~sys_fair3done_out & ~n1298;
  assign n1300 = ~n1283 & ~n1299;
  assign n1301 = ~reg_controllable_BtoS_ACK3_out & ~n1300;
  assign n1302 = ~n1288 & ~n1301;
  assign n1303 = ~reg_i_StoB_REQ3_out & ~n1302;
  assign n1304 = ~n1287 & ~n1303;
  assign n1305 = ~reg_controllable_BtoS_ACK4_out & ~n1304;
  assign n1306 = ~reg_controllable_BtoS_ACK4_out & ~n1305;
  assign n1307 = reg_i_StoB_REQ4_out & ~n1306;
  assign n1308 = ~reg_i_StoB_REQ4_out & ~n1304;
  assign n1309 = ~n1307 & ~n1308;
  assign n1310 = sys_fair4done_out & ~n1309;
  assign n1311 = sys_fair3done_out & ~n1298;
  assign n1312 = ~n169 & ~n1311;
  assign n1313 = ~reg_controllable_BtoS_ACK3_out & ~n1312;
  assign n1314 = ~reg_controllable_BtoS_ACK3_out & ~n1313;
  assign n1315 = reg_i_StoB_REQ3_out & ~n1314;
  assign n1316 = reg_controllable_BtoS_ACK3_out & ~n1312;
  assign n1317 = ~reg_controllable_BtoS_ACK3_out & ~n1298;
  assign n1318 = ~n1316 & ~n1317;
  assign n1319 = ~reg_i_StoB_REQ3_out & ~n1318;
  assign n1320 = ~n1315 & ~n1319;
  assign n1321 = ~reg_controllable_BtoS_ACK4_out & ~n1320;
  assign n1322 = ~n198 & ~n1321;
  assign n1323 = ~reg_i_StoB_REQ4_out & ~n1322;
  assign n1324 = ~n219 & ~n1323;
  assign n1325 = ~sys_fair4done_out & ~n1324;
  assign n1326 = ~n1310 & ~n1325;
  assign n1327 = ~reg_controllable_BtoS_ACK5_out & ~n1326;
  assign n1328 = ~reg_controllable_BtoS_ACK5_out & ~n1327;
  assign n1329 = reg_i_StoB_REQ5_out & ~n1328;
  assign n1330 = ~reg_i_StoB_REQ5_out & ~n1326;
  assign n1331 = ~n1329 & ~n1330;
  assign n1332 = sys_fair5done_out & ~n1331;
  assign n1333 = ~reg_controllable_BtoS_ACK4_out & ~n1321;
  assign n1334 = reg_i_StoB_REQ4_out & ~n1333;
  assign n1335 = ~reg_i_StoB_REQ4_out & ~n1320;
  assign n1336 = ~n1334 & ~n1335;
  assign n1337 = sys_fair4done_out & ~n1336;
  assign n1338 = ~n1325 & ~n1337;
  assign n1339 = ~reg_controllable_BtoS_ACK5_out & ~n1338;
  assign n1340 = ~n222 & ~n1339;
  assign n1341 = ~reg_i_StoB_REQ5_out & ~n1340;
  assign n1342 = ~n243 & ~n1341;
  assign n1343 = ~sys_fair5done_out & ~n1342;
  assign n1344 = ~n1332 & ~n1343;
  assign n1345 = ~reg_controllable_BtoS_ACK6_out & ~n1344;
  assign n1346 = ~reg_controllable_BtoS_ACK6_out & ~n1345;
  assign n1347 = reg_i_StoB_REQ6_out & ~n1346;
  assign n1348 = ~reg_i_StoB_REQ6_out & ~n1344;
  assign n1349 = ~n1347 & ~n1348;
  assign n1350 = sys_fair6done_out & ~n1349;
  assign n1351 = ~reg_controllable_BtoS_ACK5_out & ~n1339;
  assign n1352 = reg_i_StoB_REQ5_out & ~n1351;
  assign n1353 = ~reg_i_StoB_REQ5_out & ~n1338;
  assign n1354 = ~n1352 & ~n1353;
  assign n1355 = sys_fair5done_out & ~n1354;
  assign n1356 = ~n1343 & ~n1355;
  assign n1357 = ~reg_controllable_BtoS_ACK6_out & ~n1356;
  assign n1358 = ~n246 & ~n1357;
  assign n1359 = ~reg_i_StoB_REQ6_out & ~n1358;
  assign n1360 = ~n267 & ~n1359;
  assign n1361 = ~sys_fair6done_out & ~n1360;
  assign n1362 = ~n1350 & ~n1361;
  assign n1363 = ~reg_controllable_BtoS_ACK7_out & ~n1362;
  assign n1364 = ~reg_controllable_BtoS_ACK7_out & ~n1363;
  assign n1365 = reg_i_StoB_REQ7_out & ~n1364;
  assign n1366 = ~reg_i_StoB_REQ7_out & ~n1362;
  assign n1367 = ~n1365 & ~n1366;
  assign n1368 = sys_fair7done_out & ~n1367;
  assign n1369 = ~reg_controllable_BtoS_ACK6_out & ~n1357;
  assign n1370 = reg_i_StoB_REQ6_out & ~n1369;
  assign n1371 = ~reg_i_StoB_REQ6_out & ~n1356;
  assign n1372 = ~n1370 & ~n1371;
  assign n1373 = sys_fair6done_out & ~n1372;
  assign n1374 = ~n1361 & ~n1373;
  assign n1375 = ~reg_controllable_BtoS_ACK7_out & ~n1374;
  assign n1376 = ~n270 & ~n1375;
  assign n1377 = ~reg_i_StoB_REQ7_out & ~n1376;
  assign n1378 = ~n288 & ~n1377;
  assign n1379 = ~sys_fair7done_out & ~n1378;
  assign n1380 = ~n1368 & ~n1379;
  assign n1381 = sys_fair8done_out & ~n1380;
  assign n1382 = ~n291 & ~n1381;
  assign n1383 = ~reg_controllable_BtoS_ACK8_out & ~n1382;
  assign n1384 = ~reg_controllable_BtoS_ACK8_out & ~n1383;
  assign n1385 = reg_i_StoB_REQ8_out & ~n1384;
  assign n1386 = reg_controllable_BtoS_ACK8_out & ~n1382;
  assign n1387 = ~reg_controllable_BtoS_ACK7_out & ~n1375;
  assign n1388 = reg_i_StoB_REQ7_out & ~n1387;
  assign n1389 = ~reg_i_StoB_REQ7_out & ~n1374;
  assign n1390 = ~n1388 & ~n1389;
  assign n1391 = sys_fair7done_out & ~n1390;
  assign n1392 = ~n1379 & ~n1391;
  assign n1393 = ~sys_fair8done_out & ~n1392;
  assign n1394 = ~n1381 & ~n1393;
  assign n1395 = ~reg_controllable_BtoS_ACK8_out & ~n1394;
  assign n1396 = ~n1386 & ~n1395;
  assign n1397 = ~reg_i_StoB_REQ8_out & ~n1396;
  assign n1398 = ~n1385 & ~n1397;
  assign n1399 = ~reg_controllable_BtoS_ACK10_out & ~n1398;
  assign n1400 = ~reg_controllable_BtoS_ACK10_out & ~n1399;
  assign n1401 = reg_i_StoB_REQ10_out & ~n1400;
  assign n1402 = ~reg_i_StoB_REQ10_out & ~n1398;
  assign n1403 = ~n1401 & ~n1402;
  assign n1404 = sys_fair10done_out & ~n1403;
  assign n1405 = sys_fair8done_out & ~n1392;
  assign n1406 = ~n291 & ~n1405;
  assign n1407 = ~reg_controllable_BtoS_ACK8_out & ~n1406;
  assign n1408 = ~reg_controllable_BtoS_ACK8_out & ~n1407;
  assign n1409 = reg_i_StoB_REQ8_out & ~n1408;
  assign n1410 = reg_controllable_BtoS_ACK8_out & ~n1406;
  assign n1411 = ~reg_controllable_BtoS_ACK8_out & ~n1392;
  assign n1412 = ~n1410 & ~n1411;
  assign n1413 = ~reg_i_StoB_REQ8_out & ~n1412;
  assign n1414 = ~n1409 & ~n1413;
  assign n1415 = ~reg_controllable_BtoS_ACK10_out & ~n1414;
  assign n1416 = ~n320 & ~n1415;
  assign n1417 = ~reg_i_StoB_REQ10_out & ~n1416;
  assign n1418 = ~n338 & ~n1417;
  assign n1419 = ~sys_fair10done_out & ~n1418;
  assign n1420 = ~n1404 & ~n1419;
  assign n1421 = sys_fair11done_out & ~n1420;
  assign n1422 = ~n341 & ~n1421;
  assign n1423 = ~reg_controllable_BtoS_ACK11_out & ~n1422;
  assign n1424 = ~reg_controllable_BtoS_ACK11_out & ~n1423;
  assign n1425 = reg_i_StoB_REQ11_out & ~n1424;
  assign n1426 = ~sys_fair12done_out & ~n379;
  assign n1427 = ~n1127 & ~n1426;
  assign n1428 = sys_fair2done_out & ~n1427;
  assign n1429 = ~n513 & ~n1428;
  assign n1430 = reg_controllable_BtoS_ACK2_out & ~n1429;
  assign n1431 = ~n1138 & ~n1426;
  assign n1432 = ~sys_fair2done_out & ~n1431;
  assign n1433 = ~n1428 & ~n1432;
  assign n1434 = ~reg_controllable_BtoS_ACK2_out & ~n1433;
  assign n1435 = ~n1430 & ~n1434;
  assign n1436 = ~reg_i_StoB_REQ2_out & ~n1435;
  assign n1437 = ~n1274 & ~n1436;
  assign n1438 = sys_fair3done_out & ~n1437;
  assign n1439 = ~n527 & ~n1438;
  assign n1440 = reg_controllable_BtoS_ACK3_out & ~n1439;
  assign n1441 = sys_fair2done_out & ~n1431;
  assign n1442 = ~n513 & ~n1441;
  assign n1443 = reg_controllable_BtoS_ACK2_out & ~n1442;
  assign n1444 = ~reg_controllable_BtoS_ACK2_out & ~n1431;
  assign n1445 = ~n1443 & ~n1444;
  assign n1446 = ~reg_i_StoB_REQ2_out & ~n1445;
  assign n1447 = ~n1293 & ~n1446;
  assign n1448 = ~sys_fair3done_out & ~n1447;
  assign n1449 = ~n1438 & ~n1448;
  assign n1450 = ~reg_controllable_BtoS_ACK3_out & ~n1449;
  assign n1451 = ~n1440 & ~n1450;
  assign n1452 = ~reg_i_StoB_REQ3_out & ~n1451;
  assign n1453 = ~n1287 & ~n1452;
  assign n1454 = ~reg_i_StoB_REQ4_out & ~n1453;
  assign n1455 = ~n1307 & ~n1454;
  assign n1456 = sys_fair4done_out & ~n1455;
  assign n1457 = sys_fair3done_out & ~n1447;
  assign n1458 = ~n527 & ~n1457;
  assign n1459 = reg_controllable_BtoS_ACK3_out & ~n1458;
  assign n1460 = ~reg_controllable_BtoS_ACK3_out & ~n1447;
  assign n1461 = ~n1459 & ~n1460;
  assign n1462 = ~reg_i_StoB_REQ3_out & ~n1461;
  assign n1463 = ~n1315 & ~n1462;
  assign n1464 = ~reg_controllable_BtoS_ACK4_out & ~n1463;
  assign n1465 = ~n548 & ~n1464;
  assign n1466 = ~reg_i_StoB_REQ4_out & ~n1465;
  assign n1467 = ~n219 & ~n1466;
  assign n1468 = ~sys_fair4done_out & ~n1467;
  assign n1469 = ~n1456 & ~n1468;
  assign n1470 = ~reg_i_StoB_REQ5_out & ~n1469;
  assign n1471 = ~n1329 & ~n1470;
  assign n1472 = sys_fair5done_out & ~n1471;
  assign n1473 = ~reg_i_StoB_REQ4_out & ~n1463;
  assign n1474 = ~n1334 & ~n1473;
  assign n1475 = sys_fair4done_out & ~n1474;
  assign n1476 = ~n1468 & ~n1475;
  assign n1477 = ~reg_controllable_BtoS_ACK5_out & ~n1476;
  assign n1478 = ~n567 & ~n1477;
  assign n1479 = ~reg_i_StoB_REQ5_out & ~n1478;
  assign n1480 = ~n243 & ~n1479;
  assign n1481 = ~sys_fair5done_out & ~n1480;
  assign n1482 = ~n1472 & ~n1481;
  assign n1483 = ~reg_i_StoB_REQ6_out & ~n1482;
  assign n1484 = ~n1347 & ~n1483;
  assign n1485 = sys_fair6done_out & ~n1484;
  assign n1486 = ~reg_i_StoB_REQ5_out & ~n1476;
  assign n1487 = ~n1352 & ~n1486;
  assign n1488 = sys_fair5done_out & ~n1487;
  assign n1489 = ~n1481 & ~n1488;
  assign n1490 = ~reg_controllable_BtoS_ACK6_out & ~n1489;
  assign n1491 = ~n583 & ~n1490;
  assign n1492 = ~reg_i_StoB_REQ6_out & ~n1491;
  assign n1493 = ~n267 & ~n1492;
  assign n1494 = ~sys_fair6done_out & ~n1493;
  assign n1495 = ~n1485 & ~n1494;
  assign n1496 = ~reg_i_StoB_REQ7_out & ~n1495;
  assign n1497 = ~n1365 & ~n1496;
  assign n1498 = sys_fair7done_out & ~n1497;
  assign n1499 = ~reg_i_StoB_REQ6_out & ~n1489;
  assign n1500 = ~n1370 & ~n1499;
  assign n1501 = sys_fair6done_out & ~n1500;
  assign n1502 = ~n1494 & ~n1501;
  assign n1503 = ~reg_controllable_BtoS_ACK7_out & ~n1502;
  assign n1504 = ~n599 & ~n1503;
  assign n1505 = ~reg_i_StoB_REQ7_out & ~n1504;
  assign n1506 = ~n288 & ~n1505;
  assign n1507 = ~sys_fair7done_out & ~n1506;
  assign n1508 = ~n1498 & ~n1507;
  assign n1509 = sys_fair8done_out & ~n1508;
  assign n1510 = ~n613 & ~n1509;
  assign n1511 = reg_controllable_BtoS_ACK8_out & ~n1510;
  assign n1512 = ~reg_i_StoB_REQ7_out & ~n1502;
  assign n1513 = ~n1388 & ~n1512;
  assign n1514 = sys_fair7done_out & ~n1513;
  assign n1515 = ~n1507 & ~n1514;
  assign n1516 = ~sys_fair8done_out & ~n1515;
  assign n1517 = ~n1509 & ~n1516;
  assign n1518 = ~reg_controllable_BtoS_ACK8_out & ~n1517;
  assign n1519 = ~n1511 & ~n1518;
  assign n1520 = ~reg_i_StoB_REQ8_out & ~n1519;
  assign n1521 = ~n1385 & ~n1520;
  assign n1522 = ~reg_i_StoB_REQ10_out & ~n1521;
  assign n1523 = ~n1401 & ~n1522;
  assign n1524 = sys_fair10done_out & ~n1523;
  assign n1525 = sys_fair8done_out & ~n1515;
  assign n1526 = ~n613 & ~n1525;
  assign n1527 = reg_controllable_BtoS_ACK8_out & ~n1526;
  assign n1528 = ~reg_controllable_BtoS_ACK8_out & ~n1515;
  assign n1529 = ~n1527 & ~n1528;
  assign n1530 = ~reg_i_StoB_REQ8_out & ~n1529;
  assign n1531 = ~n1409 & ~n1530;
  assign n1532 = ~reg_controllable_BtoS_ACK10_out & ~n1531;
  assign n1533 = ~n631 & ~n1532;
  assign n1534 = ~reg_i_StoB_REQ10_out & ~n1533;
  assign n1535 = ~n338 & ~n1534;
  assign n1536 = ~sys_fair10done_out & ~n1535;
  assign n1537 = ~n1524 & ~n1536;
  assign n1538 = sys_fair11done_out & ~n1537;
  assign n1539 = ~n648 & ~n1538;
  assign n1540 = reg_controllable_BtoS_ACK11_out & ~n1539;
  assign n1541 = ~reg_controllable_BtoS_ACK10_out & ~n1415;
  assign n1542 = reg_i_StoB_REQ10_out & ~n1541;
  assign n1543 = ~reg_i_StoB_REQ10_out & ~n1531;
  assign n1544 = ~n1542 & ~n1543;
  assign n1545 = sys_fair10done_out & ~n1544;
  assign n1546 = ~n1536 & ~n1545;
  assign n1547 = ~sys_fair11done_out & ~n1546;
  assign n1548 = ~n1538 & ~n1547;
  assign n1549 = ~reg_controllable_BtoS_ACK11_out & ~n1548;
  assign n1550 = ~n1540 & ~n1549;
  assign n1551 = ~reg_i_StoB_REQ11_out & ~n1550;
  assign n1552 = ~n1425 & ~n1551;
  assign n1553 = sys_fair9done_out & ~n1552;
  assign n1554 = ~n1262 & ~n1553;
  assign n1555 = fair_cnt<1>_out  & ~n1554;
  assign n1556 = ~n674 & ~n1555;
  assign n1557 = fair_cnt<0>_out  & ~n1556;
  assign n1558 = ~n677 & ~n1557;
  assign n1559 = ~env_fair0done_out & ~n1558;
  assign n1560 = ~n1268 & ~n1559;
  assign n1561 = ~reg_stateG7_0_out & ~n1560;
  assign n1562 = ~reg_stateG7_0_out & ~n1561;
  assign n1563 = reg_nstateG7_1_out & ~n1562;
  assign n1564 = ~reg_nstateG7_1_out & ~n1560;
  assign n1565 = ~n1563 & ~n1564;
  assign n1566 = ~reg_controllable_BtoR_REQ1_out & ~n1565;
  assign n1567 = ~reg_controllable_BtoR_REQ1_out & ~n1566;
  assign n1568 = reg_controllable_BtoR_REQ0_out & ~n1567;
  assign n1569 = env_fair1done_out & ~n1267;
  assign n1570 = ~env_fair1done_out & ~n1558;
  assign n1571 = ~n1569 & ~n1570;
  assign n1572 = reg_nstateG7_1_out & ~n1571;
  assign n1573 = ~reg_stateG7_0_out & ~n1571;
  assign n1574 = ~reg_stateG7_0_out & ~n1573;
  assign n1575 = ~reg_nstateG7_1_out & ~n1574;
  assign n1576 = ~n1572 & ~n1575;
  assign n1577 = reg_controllable_BtoR_REQ1_out & ~n1576;
  assign n1578 = reg_controllable_BtoS_ACK11_out & ~n332;
  assign n1579 = reg_controllable_BtoS_ACK10_out & ~n296;
  assign n1580 = reg_controllable_BtoS_ACK8_out & ~n282;
  assign n1581 = reg_controllable_BtoS_ACK7_out & ~n251;
  assign n1582 = reg_controllable_BtoS_ACK6_out & ~n227;
  assign n1583 = reg_controllable_BtoS_ACK5_out & ~n203;
  assign n1584 = reg_controllable_BtoS_ACK4_out & ~n174;
  assign n1585 = reg_controllable_BtoS_ACK3_out & ~n160;
  assign n1586 = reg_controllable_BtoS_ACK2_out & ~n139;
  assign n1587 = reg_i_StoB_REQ1_out & n114;
  assign n1588 = sys_fair0done_out & n1587;
  assign n1589 = reg_controllable_BtoS_ACK1_out & ~n105;
  assign n1590 = ~n935 & ~n1589;
  assign n1591 = reg_i_StoB_REQ1_out & ~n1590;
  assign n1592 = ~n938 & ~n1591;
  assign n1593 = ~sys_fair0done_out & ~n1592;
  assign n1594 = ~n1588 & ~n1593;
  assign n1595 = sys_fair1done_out & ~n1594;
  assign n1596 = ~reg_i_StoB_REQ1_out & ~reg_controllable_BtoS_ACK1_out;
  assign n1597 = ~n100 & ~n1596;
  assign n1598 = sys_fair0done_out & ~n1597;
  assign n1599 = ~n98 & ~n1589;
  assign n1600 = reg_i_StoB_REQ1_out & ~n1599;
  assign n1601 = ~reg_controllable_BtoS_ACK1_out & n934;
  assign n1602 = ~reg_controllable_BtoS_ACK1_out & ~n1601;
  assign n1603 = ~reg_i_StoB_REQ1_out & n1602;
  assign n1604 = ~n1600 & ~n1603;
  assign n1605 = ~sys_fair0done_out & ~n1604;
  assign n1606 = ~n1598 & ~n1605;
  assign n1607 = ~sys_fair1done_out & ~n1606;
  assign n1608 = ~n1595 & ~n1607;
  assign n1609 = sys_fair12done_out & ~n1608;
  assign n1610 = ~sys_fair0done_out & ~n1593;
  assign n1611 = sys_fair1done_out & ~n1610;
  assign n1612 = ~n1607 & ~n1611;
  assign n1613 = reg_stateG12_out & ~n1612;
  assign n1614 = ~reg_stateG12_out & n1587;
  assign n1615 = ~n1613 & ~n1614;
  assign n1616 = ~sys_fair12done_out & ~n1615;
  assign n1617 = ~n1609 & ~n1616;
  assign n1618 = sys_fair2done_out & ~n1617;
  assign n1619 = ~n101 & ~n1600;
  assign n1620 = ~sys_fair0done_out & ~n1619;
  assign n1621 = ~n103 & ~n1620;
  assign n1622 = sys_fair1done_out & ~n1621;
  assign n1623 = ~reg_controllable_BtoS_ACK1_out & ~n97;
  assign n1624 = ~reg_controllable_BtoS_ACK1_out & ~n1623;
  assign n1625 = ~reg_i_StoB_REQ1_out & n1624;
  assign n1626 = ~n100 & ~n1625;
  assign n1627 = sys_fair0done_out & ~n1626;
  assign n1628 = ~n1600 & ~n1625;
  assign n1629 = ~sys_fair0done_out & ~n1628;
  assign n1630 = ~n1627 & ~n1629;
  assign n1631 = ~sys_fair1done_out & ~n1630;
  assign n1632 = ~n1622 & ~n1631;
  assign n1633 = sys_fair12done_out & ~n1632;
  assign n1634 = reg_stateG12_out & ~n1632;
  assign n1635 = ~n1614 & ~n1634;
  assign n1636 = ~sys_fair12done_out & ~n1635;
  assign n1637 = ~n1633 & ~n1636;
  assign n1638 = ~sys_fair2done_out & ~n1637;
  assign n1639 = ~n1618 & ~n1638;
  assign n1640 = ~reg_controllable_BtoS_ACK2_out & ~n1639;
  assign n1641 = ~n1586 & ~n1640;
  assign n1642 = reg_i_StoB_REQ2_out & ~n1641;
  assign n1643 = ~sys_fair2done_out & n1587;
  assign n1644 = ~n1618 & ~n1643;
  assign n1645 = reg_controllable_BtoS_ACK2_out & ~n1644;
  assign n1646 = sys_fair12done_out & ~n1612;
  assign n1647 = ~n1616 & ~n1646;
  assign n1648 = ~sys_fair2done_out & ~n1647;
  assign n1649 = ~n1618 & ~n1648;
  assign n1650 = ~reg_controllable_BtoS_ACK2_out & ~n1649;
  assign n1651 = ~n1645 & ~n1650;
  assign n1652 = ~reg_i_StoB_REQ2_out & ~n1651;
  assign n1653 = ~n1642 & ~n1652;
  assign n1654 = sys_fair3done_out & ~n1653;
  assign n1655 = reg_controllable_BtoS_ACK2_out & ~n137;
  assign n1656 = ~reg_controllable_BtoS_ACK2_out & ~n1637;
  assign n1657 = ~n1655 & ~n1656;
  assign n1658 = reg_i_StoB_REQ2_out & ~n1657;
  assign n1659 = sys_fair2done_out & ~n1637;
  assign n1660 = ~n1643 & ~n1659;
  assign n1661 = reg_controllable_BtoS_ACK2_out & ~n1660;
  assign n1662 = ~n1656 & ~n1661;
  assign n1663 = ~reg_i_StoB_REQ2_out & ~n1662;
  assign n1664 = ~n1658 & ~n1663;
  assign n1665 = ~sys_fair3done_out & ~n1664;
  assign n1666 = ~n1654 & ~n1665;
  assign n1667 = ~reg_controllable_BtoS_ACK3_out & ~n1666;
  assign n1668 = ~n1585 & ~n1667;
  assign n1669 = reg_i_StoB_REQ3_out & ~n1668;
  assign n1670 = reg_controllable_BtoS_ACK2_out & ~n102;
  assign n1671 = ~reg_controllable_BtoS_ACK2_out & n1587;
  assign n1672 = ~n1670 & ~n1671;
  assign n1673 = reg_i_StoB_REQ2_out & ~n1672;
  assign n1674 = ~reg_i_StoB_REQ2_out & n1587;
  assign n1675 = ~n1673 & ~n1674;
  assign n1676 = ~sys_fair3done_out & ~n1675;
  assign n1677 = ~n1654 & ~n1676;
  assign n1678 = reg_controllable_BtoS_ACK3_out & ~n1677;
  assign n1679 = sys_fair2done_out & ~n1647;
  assign n1680 = ~n1638 & ~n1679;
  assign n1681 = ~reg_controllable_BtoS_ACK2_out & ~n1680;
  assign n1682 = ~n1655 & ~n1681;
  assign n1683 = reg_i_StoB_REQ2_out & ~n1682;
  assign n1684 = ~n1643 & ~n1679;
  assign n1685 = reg_controllable_BtoS_ACK2_out & ~n1684;
  assign n1686 = ~reg_controllable_BtoS_ACK2_out & ~n1647;
  assign n1687 = ~n1685 & ~n1686;
  assign n1688 = ~reg_i_StoB_REQ2_out & ~n1687;
  assign n1689 = ~n1683 & ~n1688;
  assign n1690 = ~sys_fair3done_out & ~n1689;
  assign n1691 = ~n1654 & ~n1690;
  assign n1692 = ~reg_controllable_BtoS_ACK3_out & ~n1691;
  assign n1693 = ~n1678 & ~n1692;
  assign n1694 = ~reg_i_StoB_REQ3_out & ~n1693;
  assign n1695 = ~n1669 & ~n1694;
  assign n1696 = ~reg_controllable_BtoS_ACK4_out & ~n1695;
  assign n1697 = ~n1584 & ~n1696;
  assign n1698 = reg_i_StoB_REQ4_out & ~n1697;
  assign n1699 = ~reg_i_StoB_REQ4_out & ~n1695;
  assign n1700 = ~n1698 & ~n1699;
  assign n1701 = sys_fair4done_out & ~n1700;
  assign n1702 = reg_controllable_BtoS_ACK4_out & ~n189;
  assign n1703 = reg_controllable_BtoS_ACK3_out & ~n158;
  assign n1704 = ~reg_controllable_BtoS_ACK3_out & ~n1664;
  assign n1705 = ~n1703 & ~n1704;
  assign n1706 = reg_i_StoB_REQ3_out & ~n1705;
  assign n1707 = sys_fair3done_out & ~n1664;
  assign n1708 = ~n1676 & ~n1707;
  assign n1709 = reg_controllable_BtoS_ACK3_out & ~n1708;
  assign n1710 = ~n1704 & ~n1709;
  assign n1711 = ~reg_i_StoB_REQ3_out & ~n1710;
  assign n1712 = ~n1706 & ~n1711;
  assign n1713 = ~reg_controllable_BtoS_ACK4_out & ~n1712;
  assign n1714 = ~n1702 & ~n1713;
  assign n1715 = reg_i_StoB_REQ4_out & ~n1714;
  assign n1716 = reg_controllable_BtoS_ACK3_out & ~n168;
  assign n1717 = ~reg_controllable_BtoS_ACK3_out & ~n1675;
  assign n1718 = ~n1716 & ~n1717;
  assign n1719 = reg_i_StoB_REQ3_out & ~n1718;
  assign n1720 = ~reg_i_StoB_REQ3_out & ~n1675;
  assign n1721 = ~n1719 & ~n1720;
  assign n1722 = reg_controllable_BtoS_ACK4_out & ~n1721;
  assign n1723 = sys_fair3done_out & ~n1689;
  assign n1724 = ~n1665 & ~n1723;
  assign n1725 = ~reg_controllable_BtoS_ACK3_out & ~n1724;
  assign n1726 = ~n1703 & ~n1725;
  assign n1727 = reg_i_StoB_REQ3_out & ~n1726;
  assign n1728 = ~n1676 & ~n1723;
  assign n1729 = reg_controllable_BtoS_ACK3_out & ~n1728;
  assign n1730 = ~reg_controllable_BtoS_ACK3_out & ~n1689;
  assign n1731 = ~n1729 & ~n1730;
  assign n1732 = ~reg_i_StoB_REQ3_out & ~n1731;
  assign n1733 = ~n1727 & ~n1732;
  assign n1734 = ~reg_controllable_BtoS_ACK4_out & ~n1733;
  assign n1735 = ~n1722 & ~n1734;
  assign n1736 = ~reg_i_StoB_REQ4_out & ~n1735;
  assign n1737 = ~n1715 & ~n1736;
  assign n1738 = ~sys_fair4done_out & ~n1737;
  assign n1739 = ~n1701 & ~n1738;
  assign n1740 = ~reg_controllable_BtoS_ACK5_out & ~n1739;
  assign n1741 = ~n1583 & ~n1740;
  assign n1742 = reg_i_StoB_REQ5_out & ~n1741;
  assign n1743 = ~reg_i_StoB_REQ5_out & ~n1739;
  assign n1744 = ~n1742 & ~n1743;
  assign n1745 = sys_fair5done_out & ~n1744;
  assign n1746 = reg_controllable_BtoS_ACK5_out & ~n213;
  assign n1747 = ~reg_i_StoB_REQ4_out & ~n1712;
  assign n1748 = ~n1715 & ~n1747;
  assign n1749 = sys_fair4done_out & ~n1748;
  assign n1750 = ~n1713 & ~n1722;
  assign n1751 = ~reg_i_StoB_REQ4_out & ~n1750;
  assign n1752 = ~n1715 & ~n1751;
  assign n1753 = ~sys_fair4done_out & ~n1752;
  assign n1754 = ~n1749 & ~n1753;
  assign n1755 = ~reg_controllable_BtoS_ACK5_out & ~n1754;
  assign n1756 = ~n1746 & ~n1755;
  assign n1757 = reg_i_StoB_REQ5_out & ~n1756;
  assign n1758 = ~reg_controllable_BtoS_ACK4_out & ~n1721;
  assign n1759 = ~n198 & ~n1758;
  assign n1760 = reg_i_StoB_REQ4_out & ~n1759;
  assign n1761 = ~reg_i_StoB_REQ4_out & ~n1721;
  assign n1762 = ~n1760 & ~n1761;
  assign n1763 = reg_controllable_BtoS_ACK5_out & ~n1762;
  assign n1764 = ~n1702 & ~n1734;
  assign n1765 = reg_i_StoB_REQ4_out & ~n1764;
  assign n1766 = ~reg_i_StoB_REQ4_out & ~n1733;
  assign n1767 = ~n1765 & ~n1766;
  assign n1768 = sys_fair4done_out & ~n1767;
  assign n1769 = ~n1738 & ~n1768;
  assign n1770 = ~reg_controllable_BtoS_ACK5_out & ~n1769;
  assign n1771 = ~n1763 & ~n1770;
  assign n1772 = ~reg_i_StoB_REQ5_out & ~n1771;
  assign n1773 = ~n1757 & ~n1772;
  assign n1774 = ~sys_fair5done_out & ~n1773;
  assign n1775 = ~n1745 & ~n1774;
  assign n1776 = ~reg_controllable_BtoS_ACK6_out & ~n1775;
  assign n1777 = ~n1582 & ~n1776;
  assign n1778 = reg_i_StoB_REQ6_out & ~n1777;
  assign n1779 = ~reg_i_StoB_REQ6_out & ~n1775;
  assign n1780 = ~n1778 & ~n1779;
  assign n1781 = sys_fair6done_out & ~n1780;
  assign n1782 = reg_controllable_BtoS_ACK6_out & ~n237;
  assign n1783 = ~reg_i_StoB_REQ5_out & ~n1754;
  assign n1784 = ~n1757 & ~n1783;
  assign n1785 = sys_fair5done_out & ~n1784;
  assign n1786 = ~n1755 & ~n1763;
  assign n1787 = ~reg_i_StoB_REQ5_out & ~n1786;
  assign n1788 = ~n1757 & ~n1787;
  assign n1789 = ~sys_fair5done_out & ~n1788;
  assign n1790 = ~n1785 & ~n1789;
  assign n1791 = ~reg_controllable_BtoS_ACK6_out & ~n1790;
  assign n1792 = ~n1782 & ~n1791;
  assign n1793 = reg_i_StoB_REQ6_out & ~n1792;
  assign n1794 = ~reg_controllable_BtoS_ACK5_out & ~n1762;
  assign n1795 = ~n222 & ~n1794;
  assign n1796 = reg_i_StoB_REQ5_out & ~n1795;
  assign n1797 = ~reg_i_StoB_REQ5_out & ~n1762;
  assign n1798 = ~n1796 & ~n1797;
  assign n1799 = reg_controllable_BtoS_ACK6_out & ~n1798;
  assign n1800 = ~n1746 & ~n1770;
  assign n1801 = reg_i_StoB_REQ5_out & ~n1800;
  assign n1802 = ~reg_i_StoB_REQ5_out & ~n1769;
  assign n1803 = ~n1801 & ~n1802;
  assign n1804 = sys_fair5done_out & ~n1803;
  assign n1805 = ~n1774 & ~n1804;
  assign n1806 = ~reg_controllable_BtoS_ACK6_out & ~n1805;
  assign n1807 = ~n1799 & ~n1806;
  assign n1808 = ~reg_i_StoB_REQ6_out & ~n1807;
  assign n1809 = ~n1793 & ~n1808;
  assign n1810 = ~sys_fair6done_out & ~n1809;
  assign n1811 = ~n1781 & ~n1810;
  assign n1812 = ~reg_controllable_BtoS_ACK7_out & ~n1811;
  assign n1813 = ~n1581 & ~n1812;
  assign n1814 = reg_i_StoB_REQ7_out & ~n1813;
  assign n1815 = ~reg_i_StoB_REQ7_out & ~n1811;
  assign n1816 = ~n1814 & ~n1815;
  assign n1817 = sys_fair7done_out & ~n1816;
  assign n1818 = reg_controllable_BtoS_ACK7_out & ~n261;
  assign n1819 = ~reg_i_StoB_REQ6_out & ~n1790;
  assign n1820 = ~n1793 & ~n1819;
  assign n1821 = sys_fair6done_out & ~n1820;
  assign n1822 = ~n1791 & ~n1799;
  assign n1823 = ~reg_i_StoB_REQ6_out & ~n1822;
  assign n1824 = ~n1793 & ~n1823;
  assign n1825 = ~sys_fair6done_out & ~n1824;
  assign n1826 = ~n1821 & ~n1825;
  assign n1827 = ~reg_controllable_BtoS_ACK7_out & ~n1826;
  assign n1828 = ~n1818 & ~n1827;
  assign n1829 = reg_i_StoB_REQ7_out & ~n1828;
  assign n1830 = ~reg_controllable_BtoS_ACK6_out & ~n1798;
  assign n1831 = ~n246 & ~n1830;
  assign n1832 = reg_i_StoB_REQ6_out & ~n1831;
  assign n1833 = ~reg_i_StoB_REQ6_out & ~n1798;
  assign n1834 = ~n1832 & ~n1833;
  assign n1835 = reg_controllable_BtoS_ACK7_out & ~n1834;
  assign n1836 = ~n1782 & ~n1806;
  assign n1837 = reg_i_StoB_REQ6_out & ~n1836;
  assign n1838 = ~reg_i_StoB_REQ6_out & ~n1805;
  assign n1839 = ~n1837 & ~n1838;
  assign n1840 = sys_fair6done_out & ~n1839;
  assign n1841 = ~n1810 & ~n1840;
  assign n1842 = ~reg_controllable_BtoS_ACK7_out & ~n1841;
  assign n1843 = ~n1835 & ~n1842;
  assign n1844 = ~reg_i_StoB_REQ7_out & ~n1843;
  assign n1845 = ~n1829 & ~n1844;
  assign n1846 = ~sys_fair7done_out & ~n1845;
  assign n1847 = ~n1817 & ~n1846;
  assign n1848 = sys_fair8done_out & ~n1847;
  assign n1849 = ~reg_i_StoB_REQ7_out & ~n1826;
  assign n1850 = ~n1829 & ~n1849;
  assign n1851 = sys_fair7done_out & ~n1850;
  assign n1852 = ~n1827 & ~n1835;
  assign n1853 = ~reg_i_StoB_REQ7_out & ~n1852;
  assign n1854 = ~n1829 & ~n1853;
  assign n1855 = ~sys_fair7done_out & ~n1854;
  assign n1856 = ~n1851 & ~n1855;
  assign n1857 = ~sys_fair8done_out & ~n1856;
  assign n1858 = ~n1848 & ~n1857;
  assign n1859 = ~reg_controllable_BtoS_ACK8_out & ~n1858;
  assign n1860 = ~n1580 & ~n1859;
  assign n1861 = reg_i_StoB_REQ8_out & ~n1860;
  assign n1862 = ~reg_controllable_BtoS_ACK7_out & ~n1834;
  assign n1863 = ~n270 & ~n1862;
  assign n1864 = reg_i_StoB_REQ7_out & ~n1863;
  assign n1865 = ~reg_i_StoB_REQ7_out & ~n1834;
  assign n1866 = ~n1864 & ~n1865;
  assign n1867 = ~sys_fair8done_out & ~n1866;
  assign n1868 = ~n1848 & ~n1867;
  assign n1869 = reg_controllable_BtoS_ACK8_out & ~n1868;
  assign n1870 = ~n1818 & ~n1842;
  assign n1871 = reg_i_StoB_REQ7_out & ~n1870;
  assign n1872 = ~reg_i_StoB_REQ7_out & ~n1841;
  assign n1873 = ~n1871 & ~n1872;
  assign n1874 = sys_fair7done_out & ~n1873;
  assign n1875 = ~n1846 & ~n1874;
  assign n1876 = ~sys_fair8done_out & ~n1875;
  assign n1877 = ~n1848 & ~n1876;
  assign n1878 = ~reg_controllable_BtoS_ACK8_out & ~n1877;
  assign n1879 = ~n1869 & ~n1878;
  assign n1880 = ~reg_i_StoB_REQ8_out & ~n1879;
  assign n1881 = ~n1861 & ~n1880;
  assign n1882 = ~reg_controllable_BtoS_ACK10_out & ~n1881;
  assign n1883 = ~n1579 & ~n1882;
  assign n1884 = reg_i_StoB_REQ10_out & ~n1883;
  assign n1885 = ~reg_i_StoB_REQ10_out & ~n1881;
  assign n1886 = ~n1884 & ~n1885;
  assign n1887 = sys_fair10done_out & ~n1886;
  assign n1888 = reg_controllable_BtoS_ACK10_out & ~n311;
  assign n1889 = reg_controllable_BtoS_ACK8_out & ~n280;
  assign n1890 = ~reg_controllable_BtoS_ACK8_out & ~n1856;
  assign n1891 = ~n1889 & ~n1890;
  assign n1892 = reg_i_StoB_REQ8_out & ~n1891;
  assign n1893 = sys_fair8done_out & ~n1856;
  assign n1894 = ~n1867 & ~n1893;
  assign n1895 = reg_controllable_BtoS_ACK8_out & ~n1894;
  assign n1896 = ~n1890 & ~n1895;
  assign n1897 = ~reg_i_StoB_REQ8_out & ~n1896;
  assign n1898 = ~n1892 & ~n1897;
  assign n1899 = ~reg_controllable_BtoS_ACK10_out & ~n1898;
  assign n1900 = ~n1888 & ~n1899;
  assign n1901 = reg_i_StoB_REQ10_out & ~n1900;
  assign n1902 = reg_controllable_BtoS_ACK8_out & ~n290;
  assign n1903 = ~reg_controllable_BtoS_ACK8_out & ~n1866;
  assign n1904 = ~n1902 & ~n1903;
  assign n1905 = reg_i_StoB_REQ8_out & ~n1904;
  assign n1906 = ~reg_i_StoB_REQ8_out & ~n1866;
  assign n1907 = ~n1905 & ~n1906;
  assign n1908 = reg_controllable_BtoS_ACK10_out & ~n1907;
  assign n1909 = sys_fair8done_out & ~n1875;
  assign n1910 = ~n1857 & ~n1909;
  assign n1911 = ~reg_controllable_BtoS_ACK8_out & ~n1910;
  assign n1912 = ~n1889 & ~n1911;
  assign n1913 = reg_i_StoB_REQ8_out & ~n1912;
  assign n1914 = ~n1867 & ~n1909;
  assign n1915 = reg_controllable_BtoS_ACK8_out & ~n1914;
  assign n1916 = ~reg_controllable_BtoS_ACK8_out & ~n1875;
  assign n1917 = ~n1915 & ~n1916;
  assign n1918 = ~reg_i_StoB_REQ8_out & ~n1917;
  assign n1919 = ~n1913 & ~n1918;
  assign n1920 = ~reg_controllable_BtoS_ACK10_out & ~n1919;
  assign n1921 = ~n1908 & ~n1920;
  assign n1922 = ~reg_i_StoB_REQ10_out & ~n1921;
  assign n1923 = ~n1901 & ~n1922;
  assign n1924 = ~sys_fair10done_out & ~n1923;
  assign n1925 = ~n1887 & ~n1924;
  assign n1926 = sys_fair11done_out & ~n1925;
  assign n1927 = ~reg_i_StoB_REQ10_out & ~n1898;
  assign n1928 = ~n1901 & ~n1927;
  assign n1929 = sys_fair10done_out & ~n1928;
  assign n1930 = ~n1899 & ~n1908;
  assign n1931 = ~reg_i_StoB_REQ10_out & ~n1930;
  assign n1932 = ~n1901 & ~n1931;
  assign n1933 = ~sys_fair10done_out & ~n1932;
  assign n1934 = ~n1929 & ~n1933;
  assign n1935 = ~sys_fair11done_out & ~n1934;
  assign n1936 = ~n1926 & ~n1935;
  assign n1937 = ~reg_controllable_BtoS_ACK11_out & ~n1936;
  assign n1938 = ~n1578 & ~n1937;
  assign n1939 = reg_i_StoB_REQ11_out & ~n1938;
  assign n1940 = ~reg_controllable_BtoS_ACK10_out & ~n1907;
  assign n1941 = ~n320 & ~n1940;
  assign n1942 = reg_i_StoB_REQ10_out & ~n1941;
  assign n1943 = ~reg_i_StoB_REQ10_out & ~n1907;
  assign n1944 = ~n1942 & ~n1943;
  assign n1945 = ~sys_fair11done_out & ~n1944;
  assign n1946 = ~n1926 & ~n1945;
  assign n1947 = reg_controllable_BtoS_ACK11_out & ~n1946;
  assign n1948 = ~n1888 & ~n1920;
  assign n1949 = reg_i_StoB_REQ10_out & ~n1948;
  assign n1950 = ~reg_i_StoB_REQ10_out & ~n1919;
  assign n1951 = ~n1949 & ~n1950;
  assign n1952 = sys_fair10done_out & ~n1951;
  assign n1953 = ~n1924 & ~n1952;
  assign n1954 = ~sys_fair11done_out & ~n1953;
  assign n1955 = ~n1926 & ~n1954;
  assign n1956 = ~reg_controllable_BtoS_ACK11_out & ~n1955;
  assign n1957 = ~n1947 & ~n1956;
  assign n1958 = ~reg_i_StoB_REQ11_out & ~n1957;
  assign n1959 = ~n1939 & ~n1958;
  assign n1960 = sys_fair9done_out & ~n1959;
  assign n1961 = reg_controllable_BtoS_ACK11_out & ~n340;
  assign n1962 = ~reg_controllable_BtoS_ACK11_out & ~n1944;
  assign n1963 = ~n1961 & ~n1962;
  assign n1964 = reg_i_StoB_REQ11_out & ~n1963;
  assign n1965 = ~reg_i_StoB_REQ11_out & ~n1944;
  assign n1966 = ~n1964 & ~n1965;
  assign n1967 = ~sys_fair9done_out & ~n1966;
  assign n1968 = ~n1960 & ~n1967;
  assign n1969 = fair_cnt<1>_out  & ~n1968;
  assign n1970 = ~fair_cnt<1>_out  & ~n1966;
  assign n1971 = ~n1969 & ~n1970;
  assign n1972 = fair_cnt<0>_out  & ~n1971;
  assign n1973 = ~fair_cnt<0>_out  & ~n1966;
  assign n1974 = ~n1972 & ~n1973;
  assign n1975 = ~reg_controllable_BtoR_REQ1_out & ~n1974;
  assign n1976 = ~n1577 & ~n1975;
  assign n1977 = ~reg_controllable_BtoR_REQ0_out & ~n1976;
  assign n1978 = ~n1568 & ~n1977;
  assign n1979 = reg_i_RtoB_ACK1_out & ~n1978;
  assign n1980 = ~sys_fair0done_out & ~n105;
  assign n1981 = ~n1588 & ~n1980;
  assign n1982 = sys_fair1done_out & ~n1981;
  assign n1983 = ~reg_i_StoB_REQ1_out & ~n1596;
  assign n1984 = sys_fair0done_out & ~n1983;
  assign n1985 = reg_i_StoB_REQ1_out & ~n105;
  assign n1986 = ~reg_controllable_BtoS_ACK1_out & n105;
  assign n1987 = ~reg_controllable_BtoS_ACK1_out & ~n1986;
  assign n1988 = ~reg_i_StoB_REQ1_out & n1987;
  assign n1989 = ~n1985 & ~n1988;
  assign n1990 = ~sys_fair0done_out & ~n1989;
  assign n1991 = ~n1984 & ~n1990;
  assign n1992 = ~sys_fair1done_out & ~n1991;
  assign n1993 = ~n1982 & ~n1992;
  assign n1994 = sys_fair12done_out & ~n1993;
  assign n1995 = ~sys_fair0done_out & ~n1980;
  assign n1996 = sys_fair1done_out & ~n1995;
  assign n1997 = ~n1992 & ~n1996;
  assign n1998 = reg_stateG12_out & ~n1997;
  assign n1999 = ~n1614 & ~n1998;
  assign n2000 = ~sys_fair12done_out & ~n1999;
  assign n2001 = ~n1994 & ~n2000;
  assign n2002 = sys_fair2done_out & ~n2001;
  assign n2003 = sys_fair12done_out & ~n1997;
  assign n2004 = ~n2000 & ~n2003;
  assign n2005 = ~sys_fair2done_out & ~n2004;
  assign n2006 = ~n2002 & ~n2005;
  assign n2007 = ~reg_controllable_BtoS_ACK2_out & ~n2006;
  assign n2008 = ~n1586 & ~n2007;
  assign n2009 = reg_i_StoB_REQ2_out & ~n2008;
  assign n2010 = ~n1643 & ~n2002;
  assign n2011 = reg_controllable_BtoS_ACK2_out & ~n2010;
  assign n2012 = ~n2007 & ~n2011;
  assign n2013 = ~reg_i_StoB_REQ2_out & ~n2012;
  assign n2014 = ~n2009 & ~n2013;
  assign n2015 = sys_fair3done_out & ~n2014;
  assign n2016 = ~reg_controllable_BtoS_ACK2_out & ~n2004;
  assign n2017 = ~n1655 & ~n2016;
  assign n2018 = reg_i_StoB_REQ2_out & ~n2017;
  assign n2019 = sys_fair2done_out & ~n2004;
  assign n2020 = ~n1643 & ~n2019;
  assign n2021 = reg_controllable_BtoS_ACK2_out & ~n2020;
  assign n2022 = ~n2016 & ~n2021;
  assign n2023 = ~reg_i_StoB_REQ2_out & ~n2022;
  assign n2024 = ~n2018 & ~n2023;
  assign n2025 = ~sys_fair3done_out & ~n2024;
  assign n2026 = ~n2015 & ~n2025;
  assign n2027 = ~reg_controllable_BtoS_ACK3_out & ~n2026;
  assign n2028 = ~n1585 & ~n2027;
  assign n2029 = reg_i_StoB_REQ3_out & ~n2028;
  assign n2030 = ~n1676 & ~n2015;
  assign n2031 = reg_controllable_BtoS_ACK3_out & ~n2030;
  assign n2032 = ~n2027 & ~n2031;
  assign n2033 = ~reg_i_StoB_REQ3_out & ~n2032;
  assign n2034 = ~n2029 & ~n2033;
  assign n2035 = ~reg_controllable_BtoS_ACK4_out & ~n2034;
  assign n2036 = ~n1584 & ~n2035;
  assign n2037 = reg_i_StoB_REQ4_out & ~n2036;
  assign n2038 = ~reg_i_StoB_REQ4_out & ~n2034;
  assign n2039 = ~n2037 & ~n2038;
  assign n2040 = sys_fair4done_out & ~n2039;
  assign n2041 = ~reg_controllable_BtoS_ACK3_out & ~n2024;
  assign n2042 = ~n1703 & ~n2041;
  assign n2043 = reg_i_StoB_REQ3_out & ~n2042;
  assign n2044 = sys_fair3done_out & ~n2024;
  assign n2045 = ~n1676 & ~n2044;
  assign n2046 = reg_controllable_BtoS_ACK3_out & ~n2045;
  assign n2047 = ~n2041 & ~n2046;
  assign n2048 = ~reg_i_StoB_REQ3_out & ~n2047;
  assign n2049 = ~n2043 & ~n2048;
  assign n2050 = ~reg_controllable_BtoS_ACK4_out & ~n2049;
  assign n2051 = ~n1702 & ~n2050;
  assign n2052 = reg_i_StoB_REQ4_out & ~n2051;
  assign n2053 = ~n1722 & ~n2050;
  assign n2054 = ~reg_i_StoB_REQ4_out & ~n2053;
  assign n2055 = ~n2052 & ~n2054;
  assign n2056 = ~sys_fair4done_out & ~n2055;
  assign n2057 = ~n2040 & ~n2056;
  assign n2058 = ~reg_controllable_BtoS_ACK5_out & ~n2057;
  assign n2059 = ~n1583 & ~n2058;
  assign n2060 = reg_i_StoB_REQ5_out & ~n2059;
  assign n2061 = ~reg_i_StoB_REQ5_out & ~n2057;
  assign n2062 = ~n2060 & ~n2061;
  assign n2063 = sys_fair5done_out & ~n2062;
  assign n2064 = ~reg_i_StoB_REQ4_out & ~n2049;
  assign n2065 = ~n2052 & ~n2064;
  assign n2066 = sys_fair4done_out & ~n2065;
  assign n2067 = ~n2056 & ~n2066;
  assign n2068 = ~reg_controllable_BtoS_ACK5_out & ~n2067;
  assign n2069 = ~n1746 & ~n2068;
  assign n2070 = reg_i_StoB_REQ5_out & ~n2069;
  assign n2071 = ~n1763 & ~n2068;
  assign n2072 = ~reg_i_StoB_REQ5_out & ~n2071;
  assign n2073 = ~n2070 & ~n2072;
  assign n2074 = ~sys_fair5done_out & ~n2073;
  assign n2075 = ~n2063 & ~n2074;
  assign n2076 = ~reg_controllable_BtoS_ACK6_out & ~n2075;
  assign n2077 = ~n1582 & ~n2076;
  assign n2078 = reg_i_StoB_REQ6_out & ~n2077;
  assign n2079 = ~reg_i_StoB_REQ6_out & ~n2075;
  assign n2080 = ~n2078 & ~n2079;
  assign n2081 = sys_fair6done_out & ~n2080;
  assign n2082 = ~reg_i_StoB_REQ5_out & ~n2067;
  assign n2083 = ~n2070 & ~n2082;
  assign n2084 = sys_fair5done_out & ~n2083;
  assign n2085 = ~n2074 & ~n2084;
  assign n2086 = ~reg_controllable_BtoS_ACK6_out & ~n2085;
  assign n2087 = ~n1782 & ~n2086;
  assign n2088 = reg_i_StoB_REQ6_out & ~n2087;
  assign n2089 = ~n1799 & ~n2086;
  assign n2090 = ~reg_i_StoB_REQ6_out & ~n2089;
  assign n2091 = ~n2088 & ~n2090;
  assign n2092 = ~sys_fair6done_out & ~n2091;
  assign n2093 = ~n2081 & ~n2092;
  assign n2094 = ~reg_controllable_BtoS_ACK7_out & ~n2093;
  assign n2095 = ~n1581 & ~n2094;
  assign n2096 = reg_i_StoB_REQ7_out & ~n2095;
  assign n2097 = ~reg_i_StoB_REQ7_out & ~n2093;
  assign n2098 = ~n2096 & ~n2097;
  assign n2099 = sys_fair7done_out & ~n2098;
  assign n2100 = ~reg_i_StoB_REQ6_out & ~n2085;
  assign n2101 = ~n2088 & ~n2100;
  assign n2102 = sys_fair6done_out & ~n2101;
  assign n2103 = ~n2092 & ~n2102;
  assign n2104 = ~reg_controllable_BtoS_ACK7_out & ~n2103;
  assign n2105 = ~n1818 & ~n2104;
  assign n2106 = reg_i_StoB_REQ7_out & ~n2105;
  assign n2107 = ~n1835 & ~n2104;
  assign n2108 = ~reg_i_StoB_REQ7_out & ~n2107;
  assign n2109 = ~n2106 & ~n2108;
  assign n2110 = ~sys_fair7done_out & ~n2109;
  assign n2111 = ~n2099 & ~n2110;
  assign n2112 = sys_fair8done_out & ~n2111;
  assign n2113 = ~reg_i_StoB_REQ7_out & ~n2103;
  assign n2114 = ~n2106 & ~n2113;
  assign n2115 = sys_fair7done_out & ~n2114;
  assign n2116 = ~n2110 & ~n2115;
  assign n2117 = ~sys_fair8done_out & ~n2116;
  assign n2118 = ~n2112 & ~n2117;
  assign n2119 = ~reg_controllable_BtoS_ACK8_out & ~n2118;
  assign n2120 = ~n1580 & ~n2119;
  assign n2121 = reg_i_StoB_REQ8_out & ~n2120;
  assign n2122 = ~n1867 & ~n2112;
  assign n2123 = reg_controllable_BtoS_ACK8_out & ~n2122;
  assign n2124 = ~n2119 & ~n2123;
  assign n2125 = ~reg_i_StoB_REQ8_out & ~n2124;
  assign n2126 = ~n2121 & ~n2125;
  assign n2127 = ~reg_controllable_BtoS_ACK10_out & ~n2126;
  assign n2128 = ~n1579 & ~n2127;
  assign n2129 = reg_i_StoB_REQ10_out & ~n2128;
  assign n2130 = ~reg_i_StoB_REQ10_out & ~n2126;
  assign n2131 = ~n2129 & ~n2130;
  assign n2132 = sys_fair10done_out & ~n2131;
  assign n2133 = ~reg_controllable_BtoS_ACK8_out & ~n2116;
  assign n2134 = ~n1889 & ~n2133;
  assign n2135 = reg_i_StoB_REQ8_out & ~n2134;
  assign n2136 = sys_fair8done_out & ~n2116;
  assign n2137 = ~n1867 & ~n2136;
  assign n2138 = reg_controllable_BtoS_ACK8_out & ~n2137;
  assign n2139 = ~n2133 & ~n2138;
  assign n2140 = ~reg_i_StoB_REQ8_out & ~n2139;
  assign n2141 = ~n2135 & ~n2140;
  assign n2142 = ~reg_controllable_BtoS_ACK10_out & ~n2141;
  assign n2143 = ~n1888 & ~n2142;
  assign n2144 = reg_i_StoB_REQ10_out & ~n2143;
  assign n2145 = ~n1908 & ~n2142;
  assign n2146 = ~reg_i_StoB_REQ10_out & ~n2145;
  assign n2147 = ~n2144 & ~n2146;
  assign n2148 = ~sys_fair10done_out & ~n2147;
  assign n2149 = ~n2132 & ~n2148;
  assign n2150 = sys_fair11done_out & ~n2149;
  assign n2151 = ~reg_i_StoB_REQ10_out & ~n2141;
  assign n2152 = ~n2144 & ~n2151;
  assign n2153 = sys_fair10done_out & ~n2152;
  assign n2154 = ~n2148 & ~n2153;
  assign n2155 = ~sys_fair11done_out & ~n2154;
  assign n2156 = ~n2150 & ~n2155;
  assign n2157 = ~reg_controllable_BtoS_ACK11_out & ~n2156;
  assign n2158 = ~n1578 & ~n2157;
  assign n2159 = reg_i_StoB_REQ11_out & ~n2158;
  assign n2160 = ~n1945 & ~n2150;
  assign n2161 = reg_controllable_BtoS_ACK11_out & ~n2160;
  assign n2162 = ~n2157 & ~n2161;
  assign n2163 = ~reg_i_StoB_REQ11_out & ~n2162;
  assign n2164 = ~n2159 & ~n2163;
  assign n2165 = sys_fair9done_out & ~n2164;
  assign n2166 = ~n1967 & ~n2165;
  assign n2167 = fair_cnt<1>_out  & ~n2166;
  assign n2168 = ~n1970 & ~n2167;
  assign n2169 = fair_cnt<0>_out  & ~n2168;
  assign n2170 = ~n1973 & ~n2169;
  assign n2171 = env_fair1done_out & ~n2170;
  assign n2172 = ~sys_fair11done_out & ~n465;
  assign n2173 = ~n427 & ~n2172;
  assign n2174 = reg_controllable_BtoS_ACK11_out & ~n2173;
  assign n2175 = ~n1962 & ~n2174;
  assign n2176 = reg_i_StoB_REQ11_out & ~n2175;
  assign n2177 = reg_controllable_BtoS_ACK10_out & ~n421;
  assign n2178 = ~n1940 & ~n2177;
  assign n2179 = reg_i_StoB_REQ10_out & ~n2178;
  assign n2180 = ~sys_fair8done_out & ~n457;
  assign n2181 = ~n418 & ~n2180;
  assign n2182 = reg_controllable_BtoS_ACK8_out & ~n2181;
  assign n2183 = ~n1903 & ~n2182;
  assign n2184 = reg_i_StoB_REQ8_out & ~n2183;
  assign n2185 = reg_controllable_BtoS_ACK7_out & ~n412;
  assign n2186 = ~n1862 & ~n2185;
  assign n2187 = reg_i_StoB_REQ7_out & ~n2186;
  assign n2188 = reg_controllable_BtoS_ACK6_out & ~n407;
  assign n2189 = ~n1830 & ~n2188;
  assign n2190 = reg_i_StoB_REQ6_out & ~n2189;
  assign n2191 = reg_controllable_BtoS_ACK5_out & ~n402;
  assign n2192 = ~n1794 & ~n2191;
  assign n2193 = reg_i_StoB_REQ5_out & ~n2192;
  assign n2194 = reg_controllable_BtoS_ACK4_out & ~n397;
  assign n2195 = ~n1758 & ~n2194;
  assign n2196 = reg_i_StoB_REQ4_out & ~n2195;
  assign n2197 = ~sys_fair3done_out & ~n437;
  assign n2198 = ~n394 & ~n2197;
  assign n2199 = reg_controllable_BtoS_ACK3_out & ~n2198;
  assign n2200 = ~n1717 & ~n2199;
  assign n2201 = reg_i_StoB_REQ3_out & ~n2200;
  assign n2202 = ~sys_fair2done_out & ~n433;
  assign n2203 = ~n390 & ~n2202;
  assign n2204 = reg_controllable_BtoS_ACK2_out & ~n2203;
  assign n2205 = ~n1671 & ~n2204;
  assign n2206 = reg_i_StoB_REQ2_out & ~n2205;
  assign n2207 = ~n101 & ~n1587;
  assign n2208 = ~sys_fair0done_out & ~n2207;
  assign n2209 = ~n1588 & ~n2208;
  assign n2210 = sys_fair1done_out & ~n2209;
  assign n2211 = reg_i_StoB_REQ1_out & n493;
  assign n2212 = sys_fair0done_out & n2211;
  assign n2213 = ~sys_fair0done_out & n1587;
  assign n2214 = ~n2212 & ~n2213;
  assign n2215 = ~sys_fair1done_out & ~n2214;
  assign n2216 = ~n2210 & ~n2215;
  assign n2217 = sys_fair12done_out & ~n2216;
  assign n2218 = ~n378 & ~n2211;
  assign n2219 = sys_fair0done_out & ~n2218;
  assign n2220 = ~n2208 & ~n2219;
  assign n2221 = sys_fair1done_out & ~n2220;
  assign n2222 = ~n2215 & ~n2221;
  assign n2223 = reg_stateG12_out & ~n2222;
  assign n2224 = ~n1614 & ~n2223;
  assign n2225 = ~sys_fair12done_out & ~n2224;
  assign n2226 = ~n2217 & ~n2225;
  assign n2227 = sys_fair2done_out & ~n2226;
  assign n2228 = ~n1643 & ~n2227;
  assign n2229 = ~reg_i_StoB_REQ2_out & ~n2228;
  assign n2230 = ~n2206 & ~n2229;
  assign n2231 = sys_fair3done_out & ~n2230;
  assign n2232 = ~n1676 & ~n2231;
  assign n2233 = ~reg_i_StoB_REQ3_out & ~n2232;
  assign n2234 = ~n2201 & ~n2233;
  assign n2235 = ~reg_i_StoB_REQ4_out & ~n2234;
  assign n2236 = ~n2196 & ~n2235;
  assign n2237 = sys_fair4done_out & ~n2236;
  assign n2238 = reg_controllable_BtoS_ACK4_out & ~n441;
  assign n2239 = ~n1758 & ~n2238;
  assign n2240 = reg_i_StoB_REQ4_out & ~n2239;
  assign n2241 = ~n1761 & ~n2240;
  assign n2242 = ~sys_fair4done_out & ~n2241;
  assign n2243 = ~n2237 & ~n2242;
  assign n2244 = ~reg_i_StoB_REQ5_out & ~n2243;
  assign n2245 = ~n2193 & ~n2244;
  assign n2246 = sys_fair5done_out & ~n2245;
  assign n2247 = reg_controllable_BtoS_ACK5_out & ~n445;
  assign n2248 = ~n1794 & ~n2247;
  assign n2249 = reg_i_StoB_REQ5_out & ~n2248;
  assign n2250 = ~n1797 & ~n2249;
  assign n2251 = ~sys_fair5done_out & ~n2250;
  assign n2252 = ~n2246 & ~n2251;
  assign n2253 = ~reg_i_StoB_REQ6_out & ~n2252;
  assign n2254 = ~n2190 & ~n2253;
  assign n2255 = sys_fair6done_out & ~n2254;
  assign n2256 = reg_controllable_BtoS_ACK6_out & ~n449;
  assign n2257 = ~n1830 & ~n2256;
  assign n2258 = reg_i_StoB_REQ6_out & ~n2257;
  assign n2259 = ~n1833 & ~n2258;
  assign n2260 = ~sys_fair6done_out & ~n2259;
  assign n2261 = ~n2255 & ~n2260;
  assign n2262 = ~reg_i_StoB_REQ7_out & ~n2261;
  assign n2263 = ~n2187 & ~n2262;
  assign n2264 = sys_fair7done_out & ~n2263;
  assign n2265 = reg_controllable_BtoS_ACK7_out & ~n453;
  assign n2266 = ~n1862 & ~n2265;
  assign n2267 = reg_i_StoB_REQ7_out & ~n2266;
  assign n2268 = ~n1865 & ~n2267;
  assign n2269 = ~sys_fair7done_out & ~n2268;
  assign n2270 = ~n2264 & ~n2269;
  assign n2271 = sys_fair8done_out & ~n2270;
  assign n2272 = ~n1867 & ~n2271;
  assign n2273 = ~reg_i_StoB_REQ8_out & ~n2272;
  assign n2274 = ~n2184 & ~n2273;
  assign n2275 = ~reg_i_StoB_REQ10_out & ~n2274;
  assign n2276 = ~n2179 & ~n2275;
  assign n2277 = sys_fair10done_out & ~n2276;
  assign n2278 = reg_controllable_BtoS_ACK10_out & ~n461;
  assign n2279 = ~n1940 & ~n2278;
  assign n2280 = reg_i_StoB_REQ10_out & ~n2279;
  assign n2281 = ~n1943 & ~n2280;
  assign n2282 = ~sys_fair10done_out & ~n2281;
  assign n2283 = ~n2277 & ~n2282;
  assign n2284 = sys_fair11done_out & ~n2283;
  assign n2285 = ~n1945 & ~n2284;
  assign n2286 = ~reg_i_StoB_REQ11_out & ~n2285;
  assign n2287 = ~n2176 & ~n2286;
  assign n2288 = sys_fair9done_out & ~n2287;
  assign n2289 = ~n1967 & ~n2288;
  assign n2290 = fair_cnt<1>_out  & ~n2289;
  assign n2291 = ~n1970 & ~n2290;
  assign n2292 = fair_cnt<0>_out  & ~n2291;
  assign n2293 = ~n1973 & ~n2292;
  assign n2294 = ~env_fair1done_out & ~n2293;
  assign n2295 = ~n2171 & ~n2294;
  assign n2296 = env_fair0done_out & ~n2295;
  assign n2297 = ~env_fair0done_out & ~n1966;
  assign n2298 = ~n2296 & ~n2297;
  assign n2299 = ~reg_stateG7_0_out & ~n2298;
  assign n2300 = ~reg_stateG7_0_out & ~n2299;
  assign n2301 = reg_nstateG7_1_out & ~n2300;
  assign n2302 = ~reg_nstateG7_1_out & ~n2298;
  assign n2303 = ~n2301 & ~n2302;
  assign n2304 = ~reg_controllable_BtoR_REQ1_out & ~n2303;
  assign n2305 = ~reg_controllable_BtoR_REQ1_out & ~n2304;
  assign n2306 = reg_controllable_BtoR_REQ0_out & ~n2305;
  assign n2307 = reg_controllable_BtoS_ACK11_out & ~n656;
  assign n2308 = ~n1937 & ~n2307;
  assign n2309 = reg_i_StoB_REQ11_out & ~n2308;
  assign n2310 = reg_controllable_BtoS_ACK10_out & ~n625;
  assign n2311 = ~n1882 & ~n2310;
  assign n2312 = reg_i_StoB_REQ10_out & ~n2311;
  assign n2313 = reg_controllable_BtoS_ACK8_out & ~n621;
  assign n2314 = ~n1859 & ~n2313;
  assign n2315 = reg_i_StoB_REQ8_out & ~n2314;
  assign n2316 = reg_controllable_BtoS_ACK7_out & ~n593;
  assign n2317 = ~n1812 & ~n2316;
  assign n2318 = reg_i_StoB_REQ7_out & ~n2317;
  assign n2319 = reg_controllable_BtoS_ACK6_out & ~n577;
  assign n2320 = ~n1776 & ~n2319;
  assign n2321 = reg_i_StoB_REQ6_out & ~n2320;
  assign n2322 = reg_controllable_BtoS_ACK5_out & ~n561;
  assign n2323 = ~n1740 & ~n2322;
  assign n2324 = reg_i_StoB_REQ5_out & ~n2323;
  assign n2325 = reg_controllable_BtoS_ACK4_out & ~n542;
  assign n2326 = ~n1696 & ~n2325;
  assign n2327 = reg_i_StoB_REQ4_out & ~n2326;
  assign n2328 = reg_controllable_BtoS_ACK3_out & ~n538;
  assign n2329 = ~n1667 & ~n2328;
  assign n2330 = reg_i_StoB_REQ3_out & ~n2329;
  assign n2331 = reg_controllable_BtoS_ACK2_out & ~n519;
  assign n2332 = ~n1640 & ~n2331;
  assign n2333 = reg_i_StoB_REQ2_out & ~n2332;
  assign n2334 = ~n1118 & ~n2219;
  assign n2335 = sys_fair1done_out & ~n2334;
  assign n2336 = ~n1125 & ~n2335;
  assign n2337 = sys_fair12done_out & ~n2336;
  assign n2338 = ~reg_stateG12_out & ~n2218;
  assign n2339 = ~n1131 & ~n2338;
  assign n2340 = ~sys_fair12done_out & ~n2339;
  assign n2341 = ~n2337 & ~n2340;
  assign n2342 = sys_fair2done_out & ~n2341;
  assign n2343 = ~sys_fair2done_out & ~n2218;
  assign n2344 = ~n2342 & ~n2343;
  assign n2345 = reg_controllable_BtoS_ACK2_out & ~n2344;
  assign n2346 = ~n1138 & ~n2340;
  assign n2347 = ~sys_fair2done_out & ~n2346;
  assign n2348 = ~n2342 & ~n2347;
  assign n2349 = ~reg_controllable_BtoS_ACK2_out & ~n2348;
  assign n2350 = ~n2345 & ~n2349;
  assign n2351 = ~reg_i_StoB_REQ2_out & ~n2350;
  assign n2352 = ~n2333 & ~n2351;
  assign n2353 = sys_fair3done_out & ~n2352;
  assign n2354 = reg_controllable_BtoS_ACK2_out & ~n379;
  assign n2355 = ~n1671 & ~n2354;
  assign n2356 = reg_i_StoB_REQ2_out & ~n2355;
  assign n2357 = ~reg_i_StoB_REQ2_out & ~n2218;
  assign n2358 = ~n2356 & ~n2357;
  assign n2359 = ~sys_fair3done_out & ~n2358;
  assign n2360 = ~n2353 & ~n2359;
  assign n2361 = reg_controllable_BtoS_ACK3_out & ~n2360;
  assign n2362 = reg_controllable_BtoS_ACK2_out & ~n517;
  assign n2363 = ~n1681 & ~n2362;
  assign n2364 = reg_i_StoB_REQ2_out & ~n2363;
  assign n2365 = sys_fair2done_out & ~n2346;
  assign n2366 = ~n2343 & ~n2365;
  assign n2367 = reg_controllable_BtoS_ACK2_out & ~n2366;
  assign n2368 = ~reg_controllable_BtoS_ACK2_out & ~n2346;
  assign n2369 = ~n2367 & ~n2368;
  assign n2370 = ~reg_i_StoB_REQ2_out & ~n2369;
  assign n2371 = ~n2364 & ~n2370;
  assign n2372 = ~sys_fair3done_out & ~n2371;
  assign n2373 = ~n2353 & ~n2372;
  assign n2374 = ~reg_controllable_BtoS_ACK3_out & ~n2373;
  assign n2375 = ~n2361 & ~n2374;
  assign n2376 = ~reg_i_StoB_REQ3_out & ~n2375;
  assign n2377 = ~n2330 & ~n2376;
  assign n2378 = ~reg_i_StoB_REQ4_out & ~n2377;
  assign n2379 = ~n2327 & ~n2378;
  assign n2380 = sys_fair4done_out & ~n2379;
  assign n2381 = reg_controllable_BtoS_ACK4_out & ~n555;
  assign n2382 = ~n1713 & ~n2381;
  assign n2383 = reg_i_StoB_REQ4_out & ~n2382;
  assign n2384 = reg_controllable_BtoS_ACK3_out & ~n526;
  assign n2385 = ~n1717 & ~n2384;
  assign n2386 = reg_i_StoB_REQ3_out & ~n2385;
  assign n2387 = ~reg_i_StoB_REQ3_out & ~n2358;
  assign n2388 = ~n2386 & ~n2387;
  assign n2389 = reg_controllable_BtoS_ACK4_out & ~n2388;
  assign n2390 = reg_controllable_BtoS_ACK3_out & ~n536;
  assign n2391 = ~n1725 & ~n2390;
  assign n2392 = reg_i_StoB_REQ3_out & ~n2391;
  assign n2393 = sys_fair3done_out & ~n2371;
  assign n2394 = ~n2359 & ~n2393;
  assign n2395 = reg_controllable_BtoS_ACK3_out & ~n2394;
  assign n2396 = ~reg_controllable_BtoS_ACK3_out & ~n2371;
  assign n2397 = ~n2395 & ~n2396;
  assign n2398 = ~reg_i_StoB_REQ3_out & ~n2397;
  assign n2399 = ~n2392 & ~n2398;
  assign n2400 = ~reg_controllable_BtoS_ACK4_out & ~n2399;
  assign n2401 = ~n2389 & ~n2400;
  assign n2402 = ~reg_i_StoB_REQ4_out & ~n2401;
  assign n2403 = ~n2383 & ~n2402;
  assign n2404 = ~sys_fair4done_out & ~n2403;
  assign n2405 = ~n2380 & ~n2404;
  assign n2406 = ~reg_i_StoB_REQ5_out & ~n2405;
  assign n2407 = ~n2324 & ~n2406;
  assign n2408 = sys_fair5done_out & ~n2407;
  assign n2409 = reg_controllable_BtoS_ACK5_out & ~n571;
  assign n2410 = ~n1755 & ~n2409;
  assign n2411 = reg_i_StoB_REQ5_out & ~n2410;
  assign n2412 = ~n548 & ~n1758;
  assign n2413 = reg_i_StoB_REQ4_out & ~n2412;
  assign n2414 = ~reg_i_StoB_REQ4_out & ~n2388;
  assign n2415 = ~n2413 & ~n2414;
  assign n2416 = reg_controllable_BtoS_ACK5_out & ~n2415;
  assign n2417 = ~n1734 & ~n2381;
  assign n2418 = reg_i_StoB_REQ4_out & ~n2417;
  assign n2419 = ~reg_i_StoB_REQ4_out & ~n2399;
  assign n2420 = ~n2418 & ~n2419;
  assign n2421 = sys_fair4done_out & ~n2420;
  assign n2422 = ~n2404 & ~n2421;
  assign n2423 = ~reg_controllable_BtoS_ACK5_out & ~n2422;
  assign n2424 = ~n2416 & ~n2423;
  assign n2425 = ~reg_i_StoB_REQ5_out & ~n2424;
  assign n2426 = ~n2411 & ~n2425;
  assign n2427 = ~sys_fair5done_out & ~n2426;
  assign n2428 = ~n2408 & ~n2427;
  assign n2429 = ~reg_i_StoB_REQ6_out & ~n2428;
  assign n2430 = ~n2321 & ~n2429;
  assign n2431 = sys_fair6done_out & ~n2430;
  assign n2432 = reg_controllable_BtoS_ACK6_out & ~n587;
  assign n2433 = ~n1791 & ~n2432;
  assign n2434 = reg_i_StoB_REQ6_out & ~n2433;
  assign n2435 = ~n567 & ~n1794;
  assign n2436 = reg_i_StoB_REQ5_out & ~n2435;
  assign n2437 = ~reg_i_StoB_REQ5_out & ~n2415;
  assign n2438 = ~n2436 & ~n2437;
  assign n2439 = reg_controllable_BtoS_ACK6_out & ~n2438;
  assign n2440 = ~n1770 & ~n2409;
  assign n2441 = reg_i_StoB_REQ5_out & ~n2440;
  assign n2442 = ~reg_i_StoB_REQ5_out & ~n2422;
  assign n2443 = ~n2441 & ~n2442;
  assign n2444 = sys_fair5done_out & ~n2443;
  assign n2445 = ~n2427 & ~n2444;
  assign n2446 = ~reg_controllable_BtoS_ACK6_out & ~n2445;
  assign n2447 = ~n2439 & ~n2446;
  assign n2448 = ~reg_i_StoB_REQ6_out & ~n2447;
  assign n2449 = ~n2434 & ~n2448;
  assign n2450 = ~sys_fair6done_out & ~n2449;
  assign n2451 = ~n2431 & ~n2450;
  assign n2452 = ~reg_i_StoB_REQ7_out & ~n2451;
  assign n2453 = ~n2318 & ~n2452;
  assign n2454 = sys_fair7done_out & ~n2453;
  assign n2455 = reg_controllable_BtoS_ACK7_out & ~n603;
  assign n2456 = ~n1827 & ~n2455;
  assign n2457 = reg_i_StoB_REQ7_out & ~n2456;
  assign n2458 = ~n583 & ~n1830;
  assign n2459 = reg_i_StoB_REQ6_out & ~n2458;
  assign n2460 = ~reg_i_StoB_REQ6_out & ~n2438;
  assign n2461 = ~n2459 & ~n2460;
  assign n2462 = reg_controllable_BtoS_ACK7_out & ~n2461;
  assign n2463 = ~n1806 & ~n2432;
  assign n2464 = reg_i_StoB_REQ6_out & ~n2463;
  assign n2465 = ~reg_i_StoB_REQ6_out & ~n2445;
  assign n2466 = ~n2464 & ~n2465;
  assign n2467 = sys_fair6done_out & ~n2466;
  assign n2468 = ~n2450 & ~n2467;
  assign n2469 = ~reg_controllable_BtoS_ACK7_out & ~n2468;
  assign n2470 = ~n2462 & ~n2469;
  assign n2471 = ~reg_i_StoB_REQ7_out & ~n2470;
  assign n2472 = ~n2457 & ~n2471;
  assign n2473 = ~sys_fair7done_out & ~n2472;
  assign n2474 = ~n2454 & ~n2473;
  assign n2475 = sys_fair8done_out & ~n2474;
  assign n2476 = ~n599 & ~n1862;
  assign n2477 = reg_i_StoB_REQ7_out & ~n2476;
  assign n2478 = ~reg_i_StoB_REQ7_out & ~n2461;
  assign n2479 = ~n2477 & ~n2478;
  assign n2480 = ~sys_fair8done_out & ~n2479;
  assign n2481 = ~n2475 & ~n2480;
  assign n2482 = reg_controllable_BtoS_ACK8_out & ~n2481;
  assign n2483 = ~n1842 & ~n2455;
  assign n2484 = reg_i_StoB_REQ7_out & ~n2483;
  assign n2485 = ~reg_i_StoB_REQ7_out & ~n2468;
  assign n2486 = ~n2484 & ~n2485;
  assign n2487 = sys_fair7done_out & ~n2486;
  assign n2488 = ~n2473 & ~n2487;
  assign n2489 = ~sys_fair8done_out & ~n2488;
  assign n2490 = ~n2475 & ~n2489;
  assign n2491 = ~reg_controllable_BtoS_ACK8_out & ~n2490;
  assign n2492 = ~n2482 & ~n2491;
  assign n2493 = ~reg_i_StoB_REQ8_out & ~n2492;
  assign n2494 = ~n2315 & ~n2493;
  assign n2495 = ~reg_i_StoB_REQ10_out & ~n2494;
  assign n2496 = ~n2312 & ~n2495;
  assign n2497 = sys_fair10done_out & ~n2496;
  assign n2498 = reg_controllable_BtoS_ACK10_out & ~n638;
  assign n2499 = ~n1899 & ~n2498;
  assign n2500 = reg_i_StoB_REQ10_out & ~n2499;
  assign n2501 = reg_controllable_BtoS_ACK8_out & ~n612;
  assign n2502 = ~n1903 & ~n2501;
  assign n2503 = reg_i_StoB_REQ8_out & ~n2502;
  assign n2504 = ~reg_i_StoB_REQ8_out & ~n2479;
  assign n2505 = ~n2503 & ~n2504;
  assign n2506 = reg_controllable_BtoS_ACK10_out & ~n2505;
  assign n2507 = reg_controllable_BtoS_ACK8_out & ~n619;
  assign n2508 = ~n1911 & ~n2507;
  assign n2509 = reg_i_StoB_REQ8_out & ~n2508;
  assign n2510 = sys_fair8done_out & ~n2488;
  assign n2511 = ~n2480 & ~n2510;
  assign n2512 = reg_controllable_BtoS_ACK8_out & ~n2511;
  assign n2513 = ~reg_controllable_BtoS_ACK8_out & ~n2488;
  assign n2514 = ~n2512 & ~n2513;
  assign n2515 = ~reg_i_StoB_REQ8_out & ~n2514;
  assign n2516 = ~n2509 & ~n2515;
  assign n2517 = ~reg_controllable_BtoS_ACK10_out & ~n2516;
  assign n2518 = ~n2506 & ~n2517;
  assign n2519 = ~reg_i_StoB_REQ10_out & ~n2518;
  assign n2520 = ~n2500 & ~n2519;
  assign n2521 = ~sys_fair10done_out & ~n2520;
  assign n2522 = ~n2497 & ~n2521;
  assign n2523 = sys_fair11done_out & ~n2522;
  assign n2524 = ~n631 & ~n1940;
  assign n2525 = reg_i_StoB_REQ10_out & ~n2524;
  assign n2526 = ~reg_i_StoB_REQ10_out & ~n2505;
  assign n2527 = ~n2525 & ~n2526;
  assign n2528 = ~sys_fair11done_out & ~n2527;
  assign n2529 = ~n2523 & ~n2528;
  assign n2530 = reg_controllable_BtoS_ACK11_out & ~n2529;
  assign n2531 = ~n1920 & ~n2498;
  assign n2532 = reg_i_StoB_REQ10_out & ~n2531;
  assign n2533 = ~reg_i_StoB_REQ10_out & ~n2516;
  assign n2534 = ~n2532 & ~n2533;
  assign n2535 = sys_fair10done_out & ~n2534;
  assign n2536 = ~n2521 & ~n2535;
  assign n2537 = ~sys_fair11done_out & ~n2536;
  assign n2538 = ~n2523 & ~n2537;
  assign n2539 = ~reg_controllable_BtoS_ACK11_out & ~n2538;
  assign n2540 = ~n2530 & ~n2539;
  assign n2541 = ~reg_i_StoB_REQ11_out & ~n2540;
  assign n2542 = ~n2309 & ~n2541;
  assign n2543 = sys_fair9done_out & ~n2542;
  assign n2544 = reg_controllable_BtoS_ACK11_out & ~n647;
  assign n2545 = ~n1962 & ~n2544;
  assign n2546 = reg_i_StoB_REQ11_out & ~n2545;
  assign n2547 = ~reg_i_StoB_REQ11_out & ~n2527;
  assign n2548 = ~n2546 & ~n2547;
  assign n2549 = ~sys_fair9done_out & ~n2548;
  assign n2550 = ~n2543 & ~n2549;
  assign n2551 = fair_cnt<1>_out  & ~n2550;
  assign n2552 = ~fair_cnt<1>_out  & ~n2548;
  assign n2553 = ~n2551 & ~n2552;
  assign n2554 = fair_cnt<0>_out  & ~n2553;
  assign n2555 = ~fair_cnt<0>_out  & ~n2548;
  assign n2556 = ~n2554 & ~n2555;
  assign n2557 = reg_nstateG7_1_out & ~n2556;
  assign n2558 = ~reg_stateG7_0_out & ~n2556;
  assign n2559 = ~reg_stateG7_0_out & ~n2558;
  assign n2560 = ~reg_nstateG7_1_out & ~n2559;
  assign n2561 = ~n2557 & ~n2560;
  assign n2562 = reg_controllable_BtoR_REQ1_out & ~n2561;
  assign n2563 = env_fair1done_out & ~n1974;
  assign n2564 = ~n2294 & ~n2563;
  assign n2565 = reg_nstateG7_1_out & ~n2564;
  assign n2566 = ~reg_nstateG7_1_out & ~n1974;
  assign n2567 = ~n2565 & ~n2566;
  assign n2568 = ~reg_controllable_BtoR_REQ1_out & ~n2567;
  assign n2569 = ~n2562 & ~n2568;
  assign n2570 = ~reg_controllable_BtoR_REQ0_out & ~n2569;
  assign n2571 = ~n2306 & ~n2570;
  assign n2572 = ~reg_i_RtoB_ACK1_out & ~n2571;
  assign n2573 = ~n1979 & ~n2572;
  assign n2574 = reg_i_RtoB_ACK0_out & ~n2573;
  assign n2575 = reg_nstateG7_1_out & ~n2559;
  assign n2576 = ~reg_nstateG7_1_out & ~n2556;
  assign n2577 = ~n2575 & ~n2576;
  assign n2578 = ~reg_controllable_BtoR_REQ1_out & ~n2577;
  assign n2579 = ~reg_controllable_BtoR_REQ1_out & ~n2578;
  assign n2580 = reg_controllable_BtoR_REQ0_out & ~n2579;
  assign n2581 = ~env_fair1done_out & ~n1966;
  assign n2582 = ~n2171 & ~n2581;
  assign n2583 = env_fair0done_out & ~n2582;
  assign n2584 = env_fair1done_out & ~n2293;
  assign n2585 = ~n2581 & ~n2584;
  assign n2586 = ~env_fair0done_out & ~n2585;
  assign n2587 = ~n2583 & ~n2586;
  assign n2588 = reg_nstateG7_1_out & ~n2587;
  assign n2589 = ~reg_stateG7_0_out & ~n2587;
  assign n2590 = ~reg_stateG7_0_out & ~n2589;
  assign n2591 = ~reg_nstateG7_1_out & ~n2590;
  assign n2592 = ~n2588 & ~n2591;
  assign n2593 = reg_controllable_BtoR_REQ1_out & ~n2592;
  assign n2594 = reg_nstateG7_1_out & ~n1974;
  assign n2595 = env_fair0done_out & ~n1974;
  assign n2596 = ~env_fair0done_out & ~n2293;
  assign n2597 = ~n2595 & ~n2596;
  assign n2598 = ~reg_nstateG7_1_out & ~n2597;
  assign n2599 = ~n2594 & ~n2598;
  assign n2600 = ~reg_controllable_BtoR_REQ1_out & ~n2599;
  assign n2601 = ~n2593 & ~n2600;
  assign n2602 = ~reg_controllable_BtoR_REQ0_out & ~n2601;
  assign n2603 = ~n2580 & ~n2602;
  assign n2604 = reg_i_RtoB_ACK1_out & ~n2603;
  assign n2605 = reg_controllable_BtoS_ACK10_out & ~n850;
  assign n2606 = reg_controllable_BtoS_ACK7_out & ~n817;
  assign n2607 = reg_controllable_BtoS_ACK6_out & ~n799;
  assign n2608 = reg_controllable_BtoS_ACK5_out & ~n781;
  assign n2609 = reg_controllable_BtoS_ACK4_out & ~n758;
  assign n2610 = ~reg_controllable_BtoS_ACK0_out & ~reg_controllable_BtoS_ACK1_out;
  assign n2611 = ~n1589 & ~n2610;
  assign n2612 = reg_i_StoB_REQ1_out & ~n2611;
  assign n2613 = ~reg_i_StoB_REQ1_out & ~reg_controllable_BtoS_ACK0_out;
  assign n2614 = ~n2612 & ~n2613;
  assign n2615 = ~sys_fair0done_out & ~n2614;
  assign n2616 = ~n1588 & ~n2615;
  assign n2617 = sys_fair1done_out & ~n2616;
  assign n2618 = reg_i_StoB_REQ1_out & ~n115;
  assign n2619 = ~n1596 & ~n2618;
  assign n2620 = sys_fair0done_out & ~n2619;
  assign n2621 = ~n114 & ~n2610;
  assign n2622 = reg_i_StoB_REQ1_out & ~n2621;
  assign n2623 = reg_controllable_BtoS_ACK0_out & ~reg_controllable_BtoS_ACK1_out;
  assign n2624 = ~reg_controllable_BtoS_ACK1_out & ~n2623;
  assign n2625 = ~reg_i_StoB_REQ1_out & n2624;
  assign n2626 = ~n2622 & ~n2625;
  assign n2627 = ~sys_fair0done_out & ~n2626;
  assign n2628 = ~n2620 & ~n2627;
  assign n2629 = ~sys_fair1done_out & ~n2628;
  assign n2630 = ~n2617 & ~n2629;
  assign n2631 = sys_fair12done_out & ~n2630;
  assign n2632 = ~sys_fair12done_out & n1587;
  assign n2633 = ~n2631 & ~n2632;
  assign n2634 = sys_fair2done_out & ~n2633;
  assign n2635 = ~sys_fair0done_out & ~n2615;
  assign n2636 = sys_fair1done_out & ~n2635;
  assign n2637 = ~n2629 & ~n2636;
  assign n2638 = sys_fair12done_out & ~n2637;
  assign n2639 = ~n2632 & ~n2638;
  assign n2640 = ~sys_fair2done_out & ~n2639;
  assign n2641 = ~n2634 & ~n2640;
  assign n2642 = ~reg_controllable_BtoS_ACK2_out & ~n2641;
  assign n2643 = ~n735 & ~n2642;
  assign n2644 = reg_i_StoB_REQ2_out & ~n2643;
  assign n2645 = ~n1643 & ~n2634;
  assign n2646 = reg_controllable_BtoS_ACK2_out & ~n2645;
  assign n2647 = ~n2642 & ~n2646;
  assign n2648 = ~reg_i_StoB_REQ2_out & ~n2647;
  assign n2649 = ~n2644 & ~n2648;
  assign n2650 = sys_fair3done_out & ~n2649;
  assign n2651 = ~reg_controllable_BtoS_ACK2_out & ~n2639;
  assign n2652 = ~n745 & ~n2651;
  assign n2653 = reg_i_StoB_REQ2_out & ~n2652;
  assign n2654 = sys_fair2done_out & ~n2639;
  assign n2655 = ~n1643 & ~n2654;
  assign n2656 = reg_controllable_BtoS_ACK2_out & ~n2655;
  assign n2657 = ~n2651 & ~n2656;
  assign n2658 = ~reg_i_StoB_REQ2_out & ~n2657;
  assign n2659 = ~n2653 & ~n2658;
  assign n2660 = ~sys_fair3done_out & ~n2659;
  assign n2661 = ~n2650 & ~n2660;
  assign n2662 = ~reg_controllable_BtoS_ACK3_out & ~n2661;
  assign n2663 = ~n755 & ~n2662;
  assign n2664 = reg_i_StoB_REQ3_out & ~n2663;
  assign n2665 = ~n1676 & ~n2650;
  assign n2666 = reg_controllable_BtoS_ACK3_out & ~n2665;
  assign n2667 = ~n2662 & ~n2666;
  assign n2668 = ~reg_i_StoB_REQ3_out & ~n2667;
  assign n2669 = ~n2664 & ~n2668;
  assign n2670 = ~reg_controllable_BtoS_ACK4_out & ~n2669;
  assign n2671 = ~n2609 & ~n2670;
  assign n2672 = reg_i_StoB_REQ4_out & ~n2671;
  assign n2673 = ~reg_i_StoB_REQ4_out & ~n2669;
  assign n2674 = ~n2672 & ~n2673;
  assign n2675 = sys_fair4done_out & ~n2674;
  assign n2676 = ~reg_controllable_BtoS_ACK3_out & ~n2659;
  assign n2677 = ~n770 & ~n2676;
  assign n2678 = reg_i_StoB_REQ3_out & ~n2677;
  assign n2679 = sys_fair3done_out & ~n2659;
  assign n2680 = ~n1676 & ~n2679;
  assign n2681 = reg_controllable_BtoS_ACK3_out & ~n2680;
  assign n2682 = ~n2676 & ~n2681;
  assign n2683 = ~reg_i_StoB_REQ3_out & ~n2682;
  assign n2684 = ~n2678 & ~n2683;
  assign n2685 = ~reg_controllable_BtoS_ACK4_out & ~n2684;
  assign n2686 = ~n198 & ~n2685;
  assign n2687 = reg_i_StoB_REQ4_out & ~n2686;
  assign n2688 = ~n1722 & ~n2685;
  assign n2689 = ~reg_i_StoB_REQ4_out & ~n2688;
  assign n2690 = ~n2687 & ~n2689;
  assign n2691 = ~sys_fair4done_out & ~n2690;
  assign n2692 = ~n2675 & ~n2691;
  assign n2693 = ~reg_controllable_BtoS_ACK5_out & ~n2692;
  assign n2694 = ~n2608 & ~n2693;
  assign n2695 = reg_i_StoB_REQ5_out & ~n2694;
  assign n2696 = ~reg_i_StoB_REQ5_out & ~n2692;
  assign n2697 = ~n2695 & ~n2696;
  assign n2698 = sys_fair5done_out & ~n2697;
  assign n2699 = reg_controllable_BtoS_ACK4_out & ~n773;
  assign n2700 = ~n2685 & ~n2699;
  assign n2701 = reg_i_StoB_REQ4_out & ~n2700;
  assign n2702 = ~reg_i_StoB_REQ4_out & ~n2684;
  assign n2703 = ~n2701 & ~n2702;
  assign n2704 = sys_fair4done_out & ~n2703;
  assign n2705 = ~n2691 & ~n2704;
  assign n2706 = ~reg_controllable_BtoS_ACK5_out & ~n2705;
  assign n2707 = ~n222 & ~n2706;
  assign n2708 = reg_i_StoB_REQ5_out & ~n2707;
  assign n2709 = ~n1763 & ~n2706;
  assign n2710 = ~reg_i_StoB_REQ5_out & ~n2709;
  assign n2711 = ~n2708 & ~n2710;
  assign n2712 = ~sys_fair5done_out & ~n2711;
  assign n2713 = ~n2698 & ~n2712;
  assign n2714 = ~reg_controllable_BtoS_ACK6_out & ~n2713;
  assign n2715 = ~n2607 & ~n2714;
  assign n2716 = reg_i_StoB_REQ6_out & ~n2715;
  assign n2717 = ~reg_i_StoB_REQ6_out & ~n2713;
  assign n2718 = ~n2716 & ~n2717;
  assign n2719 = sys_fair6done_out & ~n2718;
  assign n2720 = reg_controllable_BtoS_ACK5_out & ~n791;
  assign n2721 = ~n2706 & ~n2720;
  assign n2722 = reg_i_StoB_REQ5_out & ~n2721;
  assign n2723 = ~reg_i_StoB_REQ5_out & ~n2705;
  assign n2724 = ~n2722 & ~n2723;
  assign n2725 = sys_fair5done_out & ~n2724;
  assign n2726 = ~n2712 & ~n2725;
  assign n2727 = ~reg_controllable_BtoS_ACK6_out & ~n2726;
  assign n2728 = ~n246 & ~n2727;
  assign n2729 = reg_i_StoB_REQ6_out & ~n2728;
  assign n2730 = ~n1799 & ~n2727;
  assign n2731 = ~reg_i_StoB_REQ6_out & ~n2730;
  assign n2732 = ~n2729 & ~n2731;
  assign n2733 = ~sys_fair6done_out & ~n2732;
  assign n2734 = ~n2719 & ~n2733;
  assign n2735 = ~reg_controllable_BtoS_ACK7_out & ~n2734;
  assign n2736 = ~n2606 & ~n2735;
  assign n2737 = reg_i_StoB_REQ7_out & ~n2736;
  assign n2738 = ~reg_i_StoB_REQ7_out & ~n2734;
  assign n2739 = ~n2737 & ~n2738;
  assign n2740 = sys_fair7done_out & ~n2739;
  assign n2741 = reg_controllable_BtoS_ACK6_out & ~n809;
  assign n2742 = ~n2727 & ~n2741;
  assign n2743 = reg_i_StoB_REQ6_out & ~n2742;
  assign n2744 = ~reg_i_StoB_REQ6_out & ~n2726;
  assign n2745 = ~n2743 & ~n2744;
  assign n2746 = sys_fair6done_out & ~n2745;
  assign n2747 = ~n2733 & ~n2746;
  assign n2748 = ~reg_controllable_BtoS_ACK7_out & ~n2747;
  assign n2749 = ~n270 & ~n2748;
  assign n2750 = reg_i_StoB_REQ7_out & ~n2749;
  assign n2751 = ~n1835 & ~n2748;
  assign n2752 = ~reg_i_StoB_REQ7_out & ~n2751;
  assign n2753 = ~n2750 & ~n2752;
  assign n2754 = ~sys_fair7done_out & ~n2753;
  assign n2755 = ~n2740 & ~n2754;
  assign n2756 = sys_fair8done_out & ~n2755;
  assign n2757 = reg_controllable_BtoS_ACK7_out & ~n827;
  assign n2758 = ~n2748 & ~n2757;
  assign n2759 = reg_i_StoB_REQ7_out & ~n2758;
  assign n2760 = ~reg_i_StoB_REQ7_out & ~n2747;
  assign n2761 = ~n2759 & ~n2760;
  assign n2762 = sys_fair7done_out & ~n2761;
  assign n2763 = ~n2754 & ~n2762;
  assign n2764 = ~sys_fair8done_out & ~n2763;
  assign n2765 = ~n2756 & ~n2764;
  assign n2766 = ~reg_controllable_BtoS_ACK8_out & ~n2765;
  assign n2767 = ~n847 & ~n2766;
  assign n2768 = reg_i_StoB_REQ8_out & ~n2767;
  assign n2769 = ~n1867 & ~n2756;
  assign n2770 = reg_controllable_BtoS_ACK8_out & ~n2769;
  assign n2771 = ~n2766 & ~n2770;
  assign n2772 = ~reg_i_StoB_REQ8_out & ~n2771;
  assign n2773 = ~n2768 & ~n2772;
  assign n2774 = ~reg_controllable_BtoS_ACK10_out & ~n2773;
  assign n2775 = ~n2605 & ~n2774;
  assign n2776 = reg_i_StoB_REQ10_out & ~n2775;
  assign n2777 = ~reg_i_StoB_REQ10_out & ~n2773;
  assign n2778 = ~n2776 & ~n2777;
  assign n2779 = sys_fair10done_out & ~n2778;
  assign n2780 = ~reg_controllable_BtoS_ACK8_out & ~n2763;
  assign n2781 = ~n862 & ~n2780;
  assign n2782 = reg_i_StoB_REQ8_out & ~n2781;
  assign n2783 = sys_fair8done_out & ~n2763;
  assign n2784 = ~n1867 & ~n2783;
  assign n2785 = reg_controllable_BtoS_ACK8_out & ~n2784;
  assign n2786 = ~n2780 & ~n2785;
  assign n2787 = ~reg_i_StoB_REQ8_out & ~n2786;
  assign n2788 = ~n2782 & ~n2787;
  assign n2789 = ~reg_controllable_BtoS_ACK10_out & ~n2788;
  assign n2790 = ~n320 & ~n2789;
  assign n2791 = reg_i_StoB_REQ10_out & ~n2790;
  assign n2792 = ~n1908 & ~n2789;
  assign n2793 = ~reg_i_StoB_REQ10_out & ~n2792;
  assign n2794 = ~n2791 & ~n2793;
  assign n2795 = ~sys_fair10done_out & ~n2794;
  assign n2796 = ~n2779 & ~n2795;
  assign n2797 = sys_fair11done_out & ~n2796;
  assign n2798 = reg_controllable_BtoS_ACK10_out & ~n865;
  assign n2799 = ~n2789 & ~n2798;
  assign n2800 = reg_i_StoB_REQ10_out & ~n2799;
  assign n2801 = ~reg_i_StoB_REQ10_out & ~n2788;
  assign n2802 = ~n2800 & ~n2801;
  assign n2803 = sys_fair10done_out & ~n2802;
  assign n2804 = ~n2795 & ~n2803;
  assign n2805 = ~sys_fair11done_out & ~n2804;
  assign n2806 = ~n2797 & ~n2805;
  assign n2807 = ~reg_controllable_BtoS_ACK11_out & ~n2806;
  assign n2808 = ~n885 & ~n2807;
  assign n2809 = reg_i_StoB_REQ11_out & ~n2808;
  assign n2810 = ~n1945 & ~n2797;
  assign n2811 = reg_controllable_BtoS_ACK11_out & ~n2810;
  assign n2812 = ~n2807 & ~n2811;
  assign n2813 = ~reg_i_StoB_REQ11_out & ~n2812;
  assign n2814 = ~n2809 & ~n2813;
  assign n2815 = sys_fair9done_out & ~n2814;
  assign n2816 = ~n1967 & ~n2815;
  assign n2817 = fair_cnt<1>_out  & ~n2816;
  assign n2818 = ~n1970 & ~n2817;
  assign n2819 = ~fair_cnt<0>_out  & ~n2818;
  assign n2820 = ~n2169 & ~n2819;
  assign n2821 = env_fair0done_out & ~n2820;
  assign n2822 = ~env_fair0done_out & ~n2170;
  assign n2823 = ~n2821 & ~n2822;
  assign n2824 = ~reg_stateG7_0_out & ~n2823;
  assign n2825 = ~reg_stateG7_0_out & ~n2824;
  assign n2826 = reg_nstateG7_1_out & ~n2825;
  assign n2827 = ~reg_nstateG7_1_out & ~n2823;
  assign n2828 = ~n2826 & ~n2827;
  assign n2829 = ~reg_controllable_BtoR_REQ1_out & ~n2828;
  assign n2830 = ~reg_controllable_BtoR_REQ1_out & ~n2829;
  assign n2831 = reg_controllable_BtoR_REQ0_out & ~n2830;
  assign n2832 = env_fair1done_out & ~n2820;
  assign n2833 = ~env_fair1done_out & ~n2170;
  assign n2834 = ~n2832 & ~n2833;
  assign n2835 = reg_nstateG7_1_out & ~n2834;
  assign n2836 = ~reg_stateG7_0_out & ~n2834;
  assign n2837 = ~reg_stateG7_0_out & ~n2836;
  assign n2838 = ~reg_nstateG7_1_out & ~n2837;
  assign n2839 = ~n2835 & ~n2838;
  assign n2840 = reg_controllable_BtoR_REQ1_out & ~n2839;
  assign n2841 = fair_cnt<0>_out  & ~n2818;
  assign n2842 = ~n1973 & ~n2841;
  assign n2843 = ~env_fair1done_out & ~n2842;
  assign n2844 = ~n2832 & ~n2843;
  assign n2845 = reg_nstateG7_1_out & ~n2844;
  assign n2846 = ~env_fair0done_out & ~n2842;
  assign n2847 = ~n2821 & ~n2846;
  assign n2848 = ~reg_nstateG7_1_out & ~n2847;
  assign n2849 = ~n2845 & ~n2848;
  assign n2850 = ~reg_controllable_BtoR_REQ1_out & ~n2849;
  assign n2851 = ~n2840 & ~n2850;
  assign n2852 = ~reg_controllable_BtoR_REQ0_out & ~n2851;
  assign n2853 = ~n2831 & ~n2852;
  assign n2854 = ~reg_i_RtoB_ACK1_out & ~n2853;
  assign n2855 = ~n2604 & ~n2854;
  assign n2856 = ~reg_i_RtoB_ACK0_out & ~n2855;
  assign n2857 = ~n2574 & ~n2856;
  assign n2858 = ~reg_i_StoB_REQ9_out & ~n2857;
  assign n2859 = ~n933 & ~n2858;
  assign n2860 = reg_controllable_BtoS_ACK9_out & ~n2859;
  assign n2861 = reg_controllable_BtoS_ACK11_out & ~n1113;
  assign n2862 = ~reg_i_StoB_REQ10_out & ~n1105;
  assign n2863 = ~n1250 & ~n2862;
  assign n2864 = sys_fair10done_out & ~n2863;
  assign n2865 = ~n1110 & ~n2864;
  assign n2866 = ~sys_fair11done_out & ~n2865;
  assign n2867 = ~n1112 & ~n2866;
  assign n2868 = ~reg_controllable_BtoS_ACK11_out & ~n2867;
  assign n2869 = ~n2861 & ~n2868;
  assign n2870 = ~reg_i_StoB_REQ11_out & ~n2869;
  assign n2871 = ~n1116 & ~n2870;
  assign n2872 = sys_fair9done_out & ~n2871;
  assign n2873 = ~n890 & ~n2872;
  assign n2874 = fair_cnt<1>_out  & ~n2873;
  assign n2875 = ~n365 & ~n2874;
  assign n2876 = fair_cnt<0>_out  & ~n2875;
  assign n2877 = ~n368 & ~n2876;
  assign n2878 = env_fair0done_out & ~n2877;
  assign n2879 = reg_controllable_BtoS_ACK11_out & ~n1422;
  assign n2880 = ~reg_i_StoB_REQ10_out & ~n1414;
  assign n2881 = ~n1542 & ~n2880;
  assign n2882 = sys_fair10done_out & ~n2881;
  assign n2883 = ~n1419 & ~n2882;
  assign n2884 = ~sys_fair11done_out & ~n2883;
  assign n2885 = ~n1421 & ~n2884;
  assign n2886 = ~reg_controllable_BtoS_ACK11_out & ~n2885;
  assign n2887 = ~n2879 & ~n2886;
  assign n2888 = ~reg_i_StoB_REQ11_out & ~n2887;
  assign n2889 = ~n1425 & ~n2888;
  assign n2890 = sys_fair9done_out & ~n2889;
  assign n2891 = ~n890 & ~n2890;
  assign n2892 = fair_cnt<1>_out  & ~n2891;
  assign n2893 = ~n365 & ~n2892;
  assign n2894 = fair_cnt<0>_out  & ~n2893;
  assign n2895 = ~n368 & ~n2894;
  assign n2896 = ~env_fair0done_out & ~n2895;
  assign n2897 = ~n2878 & ~n2896;
  assign n2898 = ~reg_stateG7_0_out & ~n2897;
  assign n2899 = ~reg_stateG7_0_out & ~n2898;
  assign n2900 = reg_nstateG7_1_out & ~n2899;
  assign n2901 = ~reg_nstateG7_1_out & ~n2897;
  assign n2902 = ~n2900 & ~n2901;
  assign n2903 = ~reg_controllable_BtoR_REQ1_out & ~n2902;
  assign n2904 = ~reg_controllable_BtoR_REQ1_out & ~n2903;
  assign n2905 = reg_controllable_BtoR_REQ0_out & ~n2904;
  assign n2906 = env_fair1done_out & ~n2877;
  assign n2907 = ~env_fair1done_out & ~n2895;
  assign n2908 = ~n2906 & ~n2907;
  assign n2909 = reg_nstateG7_1_out & ~n2908;
  assign n2910 = ~reg_stateG7_0_out & ~n2908;
  assign n2911 = ~reg_stateG7_0_out & ~n2910;
  assign n2912 = ~reg_nstateG7_1_out & ~n2911;
  assign n2913 = ~n2909 & ~n2912;
  assign n2914 = reg_controllable_BtoR_REQ1_out & ~n2913;
  assign n2915 = reg_controllable_BtoS_ACK11_out & ~n330;
  assign n2916 = ~reg_controllable_BtoS_ACK11_out & ~n1934;
  assign n2917 = ~n2915 & ~n2916;
  assign n2918 = reg_i_StoB_REQ11_out & ~n2917;
  assign n2919 = sys_fair11done_out & ~n1934;
  assign n2920 = ~n1945 & ~n2919;
  assign n2921 = reg_controllable_BtoS_ACK11_out & ~n2920;
  assign n2922 = ~n2916 & ~n2921;
  assign n2923 = ~reg_i_StoB_REQ11_out & ~n2922;
  assign n2924 = ~n2918 & ~n2923;
  assign n2925 = ~sys_fair9done_out & ~n2924;
  assign n2926 = ~n1960 & ~n2925;
  assign n2927 = fair_cnt<1>_out  & ~n2926;
  assign n2928 = ~n1970 & ~n2927;
  assign n2929 = fair_cnt<0>_out  & ~n2928;
  assign n2930 = ~n1973 & ~n2929;
  assign n2931 = ~reg_controllable_BtoR_REQ1_out & ~n2930;
  assign n2932 = ~n2914 & ~n2931;
  assign n2933 = ~reg_controllable_BtoR_REQ0_out & ~n2932;
  assign n2934 = ~n2905 & ~n2933;
  assign n2935 = reg_i_RtoB_ACK1_out & ~n2934;
  assign n2936 = ~reg_controllable_BtoS_ACK11_out & ~n2154;
  assign n2937 = ~n2915 & ~n2936;
  assign n2938 = reg_i_StoB_REQ11_out & ~n2937;
  assign n2939 = sys_fair11done_out & ~n2154;
  assign n2940 = ~n1945 & ~n2939;
  assign n2941 = reg_controllable_BtoS_ACK11_out & ~n2940;
  assign n2942 = ~n2936 & ~n2941;
  assign n2943 = ~reg_i_StoB_REQ11_out & ~n2942;
  assign n2944 = ~n2938 & ~n2943;
  assign n2945 = ~sys_fair9done_out & ~n2944;
  assign n2946 = ~n2165 & ~n2945;
  assign n2947 = fair_cnt<1>_out  & ~n2946;
  assign n2948 = ~n1970 & ~n2947;
  assign n2949 = fair_cnt<0>_out  & ~n2948;
  assign n2950 = ~n1973 & ~n2949;
  assign n2951 = env_fair1done_out & ~n2950;
  assign n2952 = ~n2581 & ~n2951;
  assign n2953 = env_fair0done_out & ~n2952;
  assign n2954 = ~n2297 & ~n2953;
  assign n2955 = ~reg_stateG7_0_out & ~n2954;
  assign n2956 = ~reg_stateG7_0_out & ~n2955;
  assign n2957 = reg_nstateG7_1_out & ~n2956;
  assign n2958 = ~reg_nstateG7_1_out & ~n2954;
  assign n2959 = ~n2957 & ~n2958;
  assign n2960 = ~reg_controllable_BtoR_REQ1_out & ~n2959;
  assign n2961 = ~reg_controllable_BtoR_REQ1_out & ~n2960;
  assign n2962 = reg_controllable_BtoR_REQ0_out & ~n2961;
  assign n2963 = reg_nstateG7_1_out & ~n2930;
  assign n2964 = ~reg_stateG7_0_out & ~n2930;
  assign n2965 = ~reg_stateG7_0_out & ~n2964;
  assign n2966 = ~reg_nstateG7_1_out & ~n2965;
  assign n2967 = ~n2963 & ~n2966;
  assign n2968 = reg_controllable_BtoR_REQ1_out & ~n2967;
  assign n2969 = env_fair1done_out & ~n2930;
  assign n2970 = ~n2581 & ~n2969;
  assign n2971 = reg_nstateG7_1_out & ~n2970;
  assign n2972 = ~reg_nstateG7_1_out & ~n2930;
  assign n2973 = ~n2971 & ~n2972;
  assign n2974 = ~reg_controllable_BtoR_REQ1_out & ~n2973;
  assign n2975 = ~n2968 & ~n2974;
  assign n2976 = ~reg_controllable_BtoR_REQ0_out & ~n2975;
  assign n2977 = ~n2962 & ~n2976;
  assign n2978 = ~reg_i_RtoB_ACK1_out & ~n2977;
  assign n2979 = ~n2935 & ~n2978;
  assign n2980 = reg_i_RtoB_ACK0_out & ~n2979;
  assign n2981 = reg_nstateG7_1_out & ~n2965;
  assign n2982 = ~n2972 & ~n2981;
  assign n2983 = ~reg_controllable_BtoR_REQ1_out & ~n2982;
  assign n2984 = ~reg_controllable_BtoR_REQ1_out & ~n2983;
  assign n2985 = reg_controllable_BtoR_REQ0_out & ~n2984;
  assign n2986 = reg_nstateG7_1_out & ~n2954;
  assign n2987 = ~reg_nstateG7_1_out & ~n2956;
  assign n2988 = ~n2986 & ~n2987;
  assign n2989 = reg_controllable_BtoR_REQ1_out & ~n2988;
  assign n2990 = env_fair0done_out & ~n2930;
  assign n2991 = ~n2297 & ~n2990;
  assign n2992 = ~reg_nstateG7_1_out & ~n2991;
  assign n2993 = ~n2963 & ~n2992;
  assign n2994 = ~reg_controllable_BtoR_REQ1_out & ~n2993;
  assign n2995 = ~n2989 & ~n2994;
  assign n2996 = ~reg_controllable_BtoR_REQ0_out & ~n2995;
  assign n2997 = ~n2985 & ~n2996;
  assign n2998 = reg_i_RtoB_ACK1_out & ~n2997;
  assign n2999 = sys_fair11done_out & ~n878;
  assign n3000 = ~n341 & ~n2999;
  assign n3001 = reg_controllable_BtoS_ACK11_out & ~n3000;
  assign n3002 = ~reg_controllable_BtoS_ACK11_out & ~n2804;
  assign n3003 = ~n3001 & ~n3002;
  assign n3004 = reg_i_StoB_REQ11_out & ~n3003;
  assign n3005 = sys_fair11done_out & ~n2804;
  assign n3006 = ~n1945 & ~n3005;
  assign n3007 = reg_controllable_BtoS_ACK11_out & ~n3006;
  assign n3008 = ~n3002 & ~n3007;
  assign n3009 = ~reg_i_StoB_REQ11_out & ~n3008;
  assign n3010 = ~n3004 & ~n3009;
  assign n3011 = ~sys_fair9done_out & ~n3010;
  assign n3012 = ~n2815 & ~n3011;
  assign n3013 = fair_cnt<1>_out  & ~n3012;
  assign n3014 = ~n1970 & ~n3013;
  assign n3015 = ~fair_cnt<0>_out  & ~n3014;
  assign n3016 = ~n2949 & ~n3015;
  assign n3017 = env_fair0done_out & ~n3016;
  assign n3018 = ~env_fair0done_out & ~n2950;
  assign n3019 = ~n3017 & ~n3018;
  assign n3020 = ~reg_stateG7_0_out & ~n3019;
  assign n3021 = ~reg_stateG7_0_out & ~n3020;
  assign n3022 = reg_nstateG7_1_out & ~n3021;
  assign n3023 = ~reg_nstateG7_1_out & ~n3019;
  assign n3024 = ~n3022 & ~n3023;
  assign n3025 = ~reg_controllable_BtoR_REQ1_out & ~n3024;
  assign n3026 = ~reg_controllable_BtoR_REQ1_out & ~n3025;
  assign n3027 = reg_controllable_BtoR_REQ0_out & ~n3026;
  assign n3028 = env_fair1done_out & ~n3016;
  assign n3029 = ~env_fair1done_out & ~n2950;
  assign n3030 = ~n3028 & ~n3029;
  assign n3031 = reg_nstateG7_1_out & ~n3030;
  assign n3032 = ~reg_stateG7_0_out & ~n3030;
  assign n3033 = ~reg_stateG7_0_out & ~n3032;
  assign n3034 = ~reg_nstateG7_1_out & ~n3033;
  assign n3035 = ~n3031 & ~n3034;
  assign n3036 = reg_controllable_BtoR_REQ1_out & ~n3035;
  assign n3037 = fair_cnt<0>_out  & ~n3014;
  assign n3038 = ~n1973 & ~n3037;
  assign n3039 = ~env_fair1done_out & ~n3038;
  assign n3040 = ~n3028 & ~n3039;
  assign n3041 = reg_nstateG7_1_out & ~n3040;
  assign n3042 = ~env_fair0done_out & ~n3038;
  assign n3043 = ~n3017 & ~n3042;
  assign n3044 = ~reg_nstateG7_1_out & ~n3043;
  assign n3045 = ~n3041 & ~n3044;
  assign n3046 = ~reg_controllable_BtoR_REQ1_out & ~n3045;
  assign n3047 = ~n3036 & ~n3046;
  assign n3048 = ~reg_controllable_BtoR_REQ0_out & ~n3047;
  assign n3049 = ~n3027 & ~n3048;
  assign n3050 = ~reg_i_RtoB_ACK1_out & ~n3049;
  assign n3051 = ~n2998 & ~n3050;
  assign n3052 = ~reg_i_RtoB_ACK0_out & ~n3051;
  assign n3053 = ~n2980 & ~n3052;
  assign n3054 = reg_i_StoB_REQ9_out & ~n3053;
  assign n3055 = sys_fair11done_out & ~n2865;
  assign n3056 = ~n341 & ~n3055;
  assign n3057 = ~reg_controllable_BtoS_ACK11_out & ~n3056;
  assign n3058 = ~reg_controllable_BtoS_ACK11_out & ~n3057;
  assign n3059 = reg_i_StoB_REQ11_out & ~n3058;
  assign n3060 = sys_fair11done_out & ~n1254;
  assign n3061 = ~n648 & ~n3060;
  assign n3062 = reg_controllable_BtoS_ACK11_out & ~n3061;
  assign n3063 = ~reg_controllable_BtoS_ACK11_out & ~n1254;
  assign n3064 = ~n3062 & ~n3063;
  assign n3065 = ~reg_i_StoB_REQ11_out & ~n3064;
  assign n3066 = ~n3059 & ~n3065;
  assign n3067 = ~sys_fair9done_out & ~n3066;
  assign n3068 = ~n1261 & ~n3067;
  assign n3069 = fair_cnt<1>_out  & ~n3068;
  assign n3070 = ~n674 & ~n3069;
  assign n3071 = fair_cnt<0>_out  & ~n3070;
  assign n3072 = ~n677 & ~n3071;
  assign n3073 = env_fair0done_out & ~n3072;
  assign n3074 = sys_fair11done_out & ~n2883;
  assign n3075 = ~n341 & ~n3074;
  assign n3076 = ~reg_controllable_BtoS_ACK11_out & ~n3075;
  assign n3077 = ~reg_controllable_BtoS_ACK11_out & ~n3076;
  assign n3078 = reg_i_StoB_REQ11_out & ~n3077;
  assign n3079 = sys_fair11done_out & ~n1546;
  assign n3080 = ~n648 & ~n3079;
  assign n3081 = reg_controllable_BtoS_ACK11_out & ~n3080;
  assign n3082 = ~reg_controllable_BtoS_ACK11_out & ~n1546;
  assign n3083 = ~n3081 & ~n3082;
  assign n3084 = ~reg_i_StoB_REQ11_out & ~n3083;
  assign n3085 = ~n3078 & ~n3084;
  assign n3086 = ~sys_fair9done_out & ~n3085;
  assign n3087 = ~n1553 & ~n3086;
  assign n3088 = fair_cnt<1>_out  & ~n3087;
  assign n3089 = ~n674 & ~n3088;
  assign n3090 = fair_cnt<0>_out  & ~n3089;
  assign n3091 = ~n677 & ~n3090;
  assign n3092 = ~env_fair0done_out & ~n3091;
  assign n3093 = ~n3073 & ~n3092;
  assign n3094 = ~reg_stateG7_0_out & ~n3093;
  assign n3095 = ~reg_stateG7_0_out & ~n3094;
  assign n3096 = reg_nstateG7_1_out & ~n3095;
  assign n3097 = ~reg_nstateG7_1_out & ~n3093;
  assign n3098 = ~n3096 & ~n3097;
  assign n3099 = ~reg_controllable_BtoR_REQ1_out & ~n3098;
  assign n3100 = ~reg_controllable_BtoR_REQ1_out & ~n3099;
  assign n3101 = reg_controllable_BtoR_REQ0_out & ~n3100;
  assign n3102 = env_fair1done_out & ~n3072;
  assign n3103 = ~env_fair1done_out & ~n3091;
  assign n3104 = ~n3102 & ~n3103;
  assign n3105 = reg_nstateG7_1_out & ~n3104;
  assign n3106 = ~reg_stateG7_0_out & ~n3104;
  assign n3107 = ~reg_stateG7_0_out & ~n3106;
  assign n3108 = ~reg_nstateG7_1_out & ~n3107;
  assign n3109 = ~n3105 & ~n3108;
  assign n3110 = reg_controllable_BtoR_REQ1_out & ~n3109;
  assign n3111 = sys_fair11done_out & ~n1953;
  assign n3112 = ~n1935 & ~n3111;
  assign n3113 = ~reg_controllable_BtoS_ACK11_out & ~n3112;
  assign n3114 = ~n2915 & ~n3113;
  assign n3115 = reg_i_StoB_REQ11_out & ~n3114;
  assign n3116 = ~n1945 & ~n3111;
  assign n3117 = reg_controllable_BtoS_ACK11_out & ~n3116;
  assign n3118 = ~reg_controllable_BtoS_ACK11_out & ~n1953;
  assign n3119 = ~n3117 & ~n3118;
  assign n3120 = ~reg_i_StoB_REQ11_out & ~n3119;
  assign n3121 = ~n3115 & ~n3120;
  assign n3122 = ~sys_fair9done_out & ~n3121;
  assign n3123 = ~n1960 & ~n3122;
  assign n3124 = fair_cnt<1>_out  & ~n3123;
  assign n3125 = ~n1970 & ~n3124;
  assign n3126 = fair_cnt<0>_out  & ~n3125;
  assign n3127 = ~n1973 & ~n3126;
  assign n3128 = ~reg_controllable_BtoR_REQ1_out & ~n3127;
  assign n3129 = ~n3110 & ~n3128;
  assign n3130 = ~reg_controllable_BtoR_REQ0_out & ~n3129;
  assign n3131 = ~n3101 & ~n3130;
  assign n3132 = reg_i_RtoB_ACK1_out & ~n3131;
  assign n3133 = ~n2294 & ~n2951;
  assign n3134 = env_fair0done_out & ~n3133;
  assign n3135 = ~n2297 & ~n3134;
  assign n3136 = ~reg_stateG7_0_out & ~n3135;
  assign n3137 = ~reg_stateG7_0_out & ~n3136;
  assign n3138 = reg_nstateG7_1_out & ~n3137;
  assign n3139 = ~reg_nstateG7_1_out & ~n3135;
  assign n3140 = ~n3138 & ~n3139;
  assign n3141 = ~reg_controllable_BtoR_REQ1_out & ~n3140;
  assign n3142 = ~reg_controllable_BtoR_REQ1_out & ~n3141;
  assign n3143 = reg_controllable_BtoR_REQ0_out & ~n3142;
  assign n3144 = reg_controllable_BtoS_ACK11_out & ~n654;
  assign n3145 = ~n3113 & ~n3144;
  assign n3146 = reg_i_StoB_REQ11_out & ~n3145;
  assign n3147 = sys_fair11done_out & ~n2536;
  assign n3148 = ~n2528 & ~n3147;
  assign n3149 = reg_controllable_BtoS_ACK11_out & ~n3148;
  assign n3150 = ~reg_controllable_BtoS_ACK11_out & ~n2536;
  assign n3151 = ~n3149 & ~n3150;
  assign n3152 = ~reg_i_StoB_REQ11_out & ~n3151;
  assign n3153 = ~n3146 & ~n3152;
  assign n3154 = ~sys_fair9done_out & ~n3153;
  assign n3155 = ~n2543 & ~n3154;
  assign n3156 = fair_cnt<1>_out  & ~n3155;
  assign n3157 = ~n2552 & ~n3156;
  assign n3158 = fair_cnt<0>_out  & ~n3157;
  assign n3159 = ~n2555 & ~n3158;
  assign n3160 = reg_nstateG7_1_out & ~n3159;
  assign n3161 = ~reg_stateG7_0_out & ~n3159;
  assign n3162 = ~reg_stateG7_0_out & ~n3161;
  assign n3163 = ~reg_nstateG7_1_out & ~n3162;
  assign n3164 = ~n3160 & ~n3163;
  assign n3165 = reg_controllable_BtoR_REQ1_out & ~n3164;
  assign n3166 = env_fair1done_out & ~n3127;
  assign n3167 = ~n2294 & ~n3166;
  assign n3168 = reg_nstateG7_1_out & ~n3167;
  assign n3169 = ~reg_nstateG7_1_out & ~n3127;
  assign n3170 = ~n3168 & ~n3169;
  assign n3171 = ~reg_controllable_BtoR_REQ1_out & ~n3170;
  assign n3172 = ~n3165 & ~n3171;
  assign n3173 = ~reg_controllable_BtoR_REQ0_out & ~n3172;
  assign n3174 = ~n3143 & ~n3173;
  assign n3175 = ~reg_i_RtoB_ACK1_out & ~n3174;
  assign n3176 = ~n3132 & ~n3175;
  assign n3177 = reg_i_RtoB_ACK0_out & ~n3176;
  assign n3178 = reg_nstateG7_1_out & ~n3162;
  assign n3179 = ~reg_nstateG7_1_out & ~n3159;
  assign n3180 = ~n3178 & ~n3179;
  assign n3181 = ~reg_controllable_BtoR_REQ1_out & ~n3180;
  assign n3182 = ~reg_controllable_BtoR_REQ1_out & ~n3181;
  assign n3183 = reg_controllable_BtoR_REQ0_out & ~n3182;
  assign n3184 = ~n2586 & ~n2953;
  assign n3185 = reg_nstateG7_1_out & ~n3184;
  assign n3186 = ~reg_stateG7_0_out & ~n3184;
  assign n3187 = ~reg_stateG7_0_out & ~n3186;
  assign n3188 = ~reg_nstateG7_1_out & ~n3187;
  assign n3189 = ~n3185 & ~n3188;
  assign n3190 = reg_controllable_BtoR_REQ1_out & ~n3189;
  assign n3191 = reg_nstateG7_1_out & ~n3127;
  assign n3192 = env_fair0done_out & ~n3127;
  assign n3193 = ~n2596 & ~n3192;
  assign n3194 = ~reg_nstateG7_1_out & ~n3193;
  assign n3195 = ~n3191 & ~n3194;
  assign n3196 = ~reg_controllable_BtoR_REQ1_out & ~n3195;
  assign n3197 = ~n3190 & ~n3196;
  assign n3198 = ~reg_controllable_BtoR_REQ0_out & ~n3197;
  assign n3199 = ~n3183 & ~n3198;
  assign n3200 = reg_i_RtoB_ACK1_out & ~n3199;
  assign n3201 = ~n3050 & ~n3200;
  assign n3202 = ~reg_i_RtoB_ACK0_out & ~n3201;
  assign n3203 = ~n3177 & ~n3202;
  assign n3204 = ~reg_i_StoB_REQ9_out & ~n3203;
  assign n3205 = ~n3054 & ~n3204;
  assign n3206 = ~reg_controllable_BtoS_ACK9_out & ~n3205;
  assign n3207 = ~n2860 & ~n3206;
  assign n3208 = reg_i_nEMPTY_out & ~n3207;
  assign n3209 = reg_i_nEMPTY_out & ~n3208;
  assign n3210 = reg_i_FULL_out & ~n3209;
  assign n3211 = ~reg_stateG7_0_out & ~n369;
  assign n3212 = ~reg_stateG7_0_out & ~n3211;
  assign n3213 = reg_nstateG7_1_out & ~n3212;
  assign n3214 = ~n686 & ~n3213;
  assign n3215 = ~reg_controllable_BtoR_REQ1_out & ~n3214;
  assign n3216 = ~reg_controllable_BtoR_REQ1_out & ~n3215;
  assign n3217 = reg_controllable_BtoR_REQ0_out & ~n3216;
  assign n3218 = ~reg_nstateG7_1_out & ~n3212;
  assign n3219 = ~n714 & ~n3218;
  assign n3220 = reg_controllable_BtoR_REQ1_out & ~n3219;
  assign n3221 = reg_nstateG7_1_out & ~n702;
  assign n3222 = ~n479 & ~n715;
  assign n3223 = ~reg_nstateG7_1_out & ~n3222;
  assign n3224 = ~n3221 & ~n3223;
  assign n3225 = ~reg_controllable_BtoR_REQ1_out & ~n3224;
  assign n3226 = ~n3220 & ~n3225;
  assign n3227 = ~reg_controllable_BtoR_REQ0_out & ~n3226;
  assign n3228 = ~n3217 & ~n3227;
  assign n3229 = ~reg_i_RtoB_ACK1_out & ~n3228;
  assign n3230 = ~n724 & ~n3229;
  assign n3231 = ~reg_i_RtoB_ACK0_out & ~n3230;
  assign n3232 = ~n694 & ~n3231;
  assign n3233 = reg_i_StoB_REQ9_out & ~n3232;
  assign n3234 = env_fair0done_out & ~n2564;
  assign n3235 = ~n2297 & ~n3234;
  assign n3236 = ~reg_stateG7_0_out & ~n3235;
  assign n3237 = ~reg_stateG7_0_out & ~n3236;
  assign n3238 = reg_nstateG7_1_out & ~n3237;
  assign n3239 = ~reg_nstateG7_1_out & ~n3235;
  assign n3240 = ~n3238 & ~n3239;
  assign n3241 = ~reg_controllable_BtoR_REQ1_out & ~n3240;
  assign n3242 = ~reg_controllable_BtoR_REQ1_out & ~n3241;
  assign n3243 = reg_controllable_BtoR_REQ0_out & ~n3242;
  assign n3244 = ~n2570 & ~n3243;
  assign n3245 = ~reg_i_RtoB_ACK1_out & ~n3244;
  assign n3246 = ~n1979 & ~n3245;
  assign n3247 = reg_i_RtoB_ACK0_out & ~n3246;
  assign n3248 = ~n2563 & ~n2581;
  assign n3249 = env_fair0done_out & ~n3248;
  assign n3250 = ~n2586 & ~n3249;
  assign n3251 = reg_nstateG7_1_out & ~n3250;
  assign n3252 = ~reg_stateG7_0_out & ~n3250;
  assign n3253 = ~reg_stateG7_0_out & ~n3252;
  assign n3254 = ~reg_nstateG7_1_out & ~n3253;
  assign n3255 = ~n3251 & ~n3254;
  assign n3256 = reg_controllable_BtoR_REQ1_out & ~n3255;
  assign n3257 = ~n2600 & ~n3256;
  assign n3258 = ~reg_controllable_BtoR_REQ0_out & ~n3257;
  assign n3259 = ~n2580 & ~n3258;
  assign n3260 = reg_i_RtoB_ACK1_out & ~n3259;
  assign n3261 = ~reg_stateG7_0_out & ~n1974;
  assign n3262 = ~reg_stateG7_0_out & ~n3261;
  assign n3263 = reg_nstateG7_1_out & ~n3262;
  assign n3264 = ~n2566 & ~n3263;
  assign n3265 = ~reg_controllable_BtoR_REQ1_out & ~n3264;
  assign n3266 = ~reg_controllable_BtoR_REQ1_out & ~n3265;
  assign n3267 = reg_controllable_BtoR_REQ0_out & ~n3266;
  assign n3268 = ~reg_nstateG7_1_out & ~n3262;
  assign n3269 = ~n2594 & ~n3268;
  assign n3270 = reg_controllable_BtoR_REQ1_out & ~n3269;
  assign n3271 = reg_nstateG7_1_out & ~n3248;
  assign n3272 = ~n2297 & ~n2595;
  assign n3273 = ~reg_nstateG7_1_out & ~n3272;
  assign n3274 = ~n3271 & ~n3273;
  assign n3275 = ~reg_controllable_BtoR_REQ1_out & ~n3274;
  assign n3276 = ~n3270 & ~n3275;
  assign n3277 = ~reg_controllable_BtoR_REQ0_out & ~n3276;
  assign n3278 = ~n3267 & ~n3277;
  assign n3279 = ~reg_i_RtoB_ACK1_out & ~n3278;
  assign n3280 = ~n3260 & ~n3279;
  assign n3281 = ~reg_i_RtoB_ACK0_out & ~n3280;
  assign n3282 = ~n3247 & ~n3281;
  assign n3283 = ~reg_i_StoB_REQ9_out & ~n3282;
  assign n3284 = ~n3233 & ~n3283;
  assign n3285 = reg_controllable_BtoS_ACK9_out & ~n3284;
  assign n3286 = env_fair0done_out & ~n2970;
  assign n3287 = ~n2297 & ~n3286;
  assign n3288 = ~reg_stateG7_0_out & ~n3287;
  assign n3289 = ~reg_stateG7_0_out & ~n3288;
  assign n3290 = reg_nstateG7_1_out & ~n3289;
  assign n3291 = ~reg_nstateG7_1_out & ~n3287;
  assign n3292 = ~n3290 & ~n3291;
  assign n3293 = ~reg_controllable_BtoR_REQ1_out & ~n3292;
  assign n3294 = ~reg_controllable_BtoR_REQ1_out & ~n3293;
  assign n3295 = reg_controllable_BtoR_REQ0_out & ~n3294;
  assign n3296 = ~n2976 & ~n3295;
  assign n3297 = ~reg_i_RtoB_ACK1_out & ~n3296;
  assign n3298 = ~n2935 & ~n3297;
  assign n3299 = reg_i_RtoB_ACK0_out & ~n3298;
  assign n3300 = reg_nstateG7_1_out & ~n3287;
  assign n3301 = ~reg_nstateG7_1_out & ~n3289;
  assign n3302 = ~n3300 & ~n3301;
  assign n3303 = reg_controllable_BtoR_REQ1_out & ~n3302;
  assign n3304 = ~n2994 & ~n3303;
  assign n3305 = ~reg_controllable_BtoR_REQ0_out & ~n3304;
  assign n3306 = ~n2985 & ~n3305;
  assign n3307 = reg_i_RtoB_ACK1_out & ~n3306;
  assign n3308 = ~n2971 & ~n2992;
  assign n3309 = ~reg_controllable_BtoR_REQ1_out & ~n3308;
  assign n3310 = ~n2968 & ~n3309;
  assign n3311 = ~reg_controllable_BtoR_REQ0_out & ~n3310;
  assign n3312 = ~n2985 & ~n3311;
  assign n3313 = ~reg_i_RtoB_ACK1_out & ~n3312;
  assign n3314 = ~n3307 & ~n3313;
  assign n3315 = ~reg_i_RtoB_ACK0_out & ~n3314;
  assign n3316 = ~n3299 & ~n3315;
  assign n3317 = reg_i_StoB_REQ9_out & ~n3316;
  assign n3318 = env_fair0done_out & ~n3167;
  assign n3319 = ~n2297 & ~n3318;
  assign n3320 = ~reg_stateG7_0_out & ~n3319;
  assign n3321 = ~reg_stateG7_0_out & ~n3320;
  assign n3322 = reg_nstateG7_1_out & ~n3321;
  assign n3323 = ~reg_nstateG7_1_out & ~n3319;
  assign n3324 = ~n3322 & ~n3323;
  assign n3325 = ~reg_controllable_BtoR_REQ1_out & ~n3324;
  assign n3326 = ~reg_controllable_BtoR_REQ1_out & ~n3325;
  assign n3327 = reg_controllable_BtoR_REQ0_out & ~n3326;
  assign n3328 = ~n3173 & ~n3327;
  assign n3329 = ~reg_i_RtoB_ACK1_out & ~n3328;
  assign n3330 = ~n3132 & ~n3329;
  assign n3331 = reg_i_RtoB_ACK0_out & ~n3330;
  assign n3332 = ~n2581 & ~n3166;
  assign n3333 = env_fair0done_out & ~n3332;
  assign n3334 = ~n2586 & ~n3333;
  assign n3335 = reg_nstateG7_1_out & ~n3334;
  assign n3336 = ~reg_stateG7_0_out & ~n3334;
  assign n3337 = ~reg_stateG7_0_out & ~n3336;
  assign n3338 = ~reg_nstateG7_1_out & ~n3337;
  assign n3339 = ~n3335 & ~n3338;
  assign n3340 = reg_controllable_BtoR_REQ1_out & ~n3339;
  assign n3341 = ~n3196 & ~n3340;
  assign n3342 = ~reg_controllable_BtoR_REQ0_out & ~n3341;
  assign n3343 = ~n3183 & ~n3342;
  assign n3344 = reg_i_RtoB_ACK1_out & ~n3343;
  assign n3345 = ~reg_stateG7_0_out & ~n3127;
  assign n3346 = ~reg_stateG7_0_out & ~n3345;
  assign n3347 = reg_nstateG7_1_out & ~n3346;
  assign n3348 = ~n3169 & ~n3347;
  assign n3349 = ~reg_controllable_BtoR_REQ1_out & ~n3348;
  assign n3350 = ~reg_controllable_BtoR_REQ1_out & ~n3349;
  assign n3351 = reg_controllable_BtoR_REQ0_out & ~n3350;
  assign n3352 = ~reg_nstateG7_1_out & ~n3346;
  assign n3353 = ~n3191 & ~n3352;
  assign n3354 = reg_controllable_BtoR_REQ1_out & ~n3353;
  assign n3355 = reg_nstateG7_1_out & ~n3332;
  assign n3356 = ~n2297 & ~n3192;
  assign n3357 = ~reg_nstateG7_1_out & ~n3356;
  assign n3358 = ~n3355 & ~n3357;
  assign n3359 = ~reg_controllable_BtoR_REQ1_out & ~n3358;
  assign n3360 = ~n3354 & ~n3359;
  assign n3361 = ~reg_controllable_BtoR_REQ0_out & ~n3360;
  assign n3362 = ~n3351 & ~n3361;
  assign n3363 = ~reg_i_RtoB_ACK1_out & ~n3362;
  assign n3364 = ~n3344 & ~n3363;
  assign n3365 = ~reg_i_RtoB_ACK0_out & ~n3364;
  assign n3366 = ~n3331 & ~n3365;
  assign n3367 = ~reg_i_StoB_REQ9_out & ~n3366;
  assign n3368 = ~n3317 & ~n3367;
  assign n3369 = ~reg_controllable_BtoS_ACK9_out & ~n3368;
  assign n3370 = ~n3285 & ~n3369;
  assign n3371 = reg_i_nEMPTY_out & ~n3370;
  assign n3372 = ~n685 & ~n718;
  assign n3373 = ~reg_controllable_BtoR_REQ1_out & ~n3372;
  assign n3374 = ~n684 & ~n3373;
  assign n3375 = ~reg_controllable_BtoR_REQ0_out & ~n3374;
  assign n3376 = ~n700 & ~n3375;
  assign n3377 = ~reg_i_RtoB_ACK1_out & ~n3376;
  assign n3378 = ~reg_i_RtoB_ACK1_out & ~n3377;
  assign n3379 = ~reg_i_RtoB_ACK0_out & ~n3378;
  assign n3380 = ~reg_i_RtoB_ACK0_out & ~n3379;
  assign n3381 = reg_i_StoB_REQ9_out & ~n3380;
  assign n3382 = ~n388 & ~n952;
  assign n3383 = sys_fair2done_out & ~n3382;
  assign n3384 = ~n143 & ~n3383;
  assign n3385 = reg_controllable_BtoS_ACK2_out & ~n3384;
  assign n3386 = ~n1277 & ~n3383;
  assign n3387 = ~reg_controllable_BtoS_ACK2_out & ~n3386;
  assign n3388 = ~n3385 & ~n3387;
  assign n3389 = ~reg_i_StoB_REQ2_out & ~n3388;
  assign n3390 = ~n1274 & ~n3389;
  assign n3391 = sys_fair3done_out & ~n3390;
  assign n3392 = ~n169 & ~n3391;
  assign n3393 = reg_controllable_BtoS_ACK3_out & ~n3392;
  assign n3394 = ~n1299 & ~n3391;
  assign n3395 = ~reg_controllable_BtoS_ACK3_out & ~n3394;
  assign n3396 = ~n3393 & ~n3395;
  assign n3397 = ~reg_i_StoB_REQ3_out & ~n3396;
  assign n3398 = ~n1287 & ~n3397;
  assign n3399 = ~reg_i_StoB_REQ4_out & ~n3398;
  assign n3400 = ~n1307 & ~n3399;
  assign n3401 = sys_fair4done_out & ~n3400;
  assign n3402 = ~n1325 & ~n3401;
  assign n3403 = ~reg_i_StoB_REQ5_out & ~n3402;
  assign n3404 = ~n1329 & ~n3403;
  assign n3405 = sys_fair5done_out & ~n3404;
  assign n3406 = ~n1343 & ~n3405;
  assign n3407 = ~reg_i_StoB_REQ6_out & ~n3406;
  assign n3408 = ~n1347 & ~n3407;
  assign n3409 = sys_fair6done_out & ~n3408;
  assign n3410 = ~n1361 & ~n3409;
  assign n3411 = ~reg_i_StoB_REQ7_out & ~n3410;
  assign n3412 = ~n1365 & ~n3411;
  assign n3413 = sys_fair7done_out & ~n3412;
  assign n3414 = ~n1379 & ~n3413;
  assign n3415 = sys_fair8done_out & ~n3414;
  assign n3416 = ~n291 & ~n3415;
  assign n3417 = reg_controllable_BtoS_ACK8_out & ~n3416;
  assign n3418 = ~n1393 & ~n3415;
  assign n3419 = ~reg_controllable_BtoS_ACK8_out & ~n3418;
  assign n3420 = ~n3417 & ~n3419;
  assign n3421 = ~reg_i_StoB_REQ8_out & ~n3420;
  assign n3422 = ~n1385 & ~n3421;
  assign n3423 = ~reg_i_StoB_REQ10_out & ~n3422;
  assign n3424 = ~n1401 & ~n3423;
  assign n3425 = sys_fair10done_out & ~n3424;
  assign n3426 = ~n1419 & ~n3425;
  assign n3427 = sys_fair11done_out & ~n3426;
  assign n3428 = ~n341 & ~n3427;
  assign n3429 = ~reg_controllable_BtoS_ACK11_out & ~n3428;
  assign n3430 = ~reg_controllable_BtoS_ACK11_out & ~n3429;
  assign n3431 = reg_i_StoB_REQ11_out & ~n3430;
  assign n3432 = ~reg_controllable_BtoS_ACK10_out & ~n3422;
  assign n3433 = ~reg_controllable_BtoS_ACK10_out & ~n3432;
  assign n3434 = reg_i_StoB_REQ10_out & ~n3433;
  assign n3435 = ~reg_controllable_BtoS_ACK8_out & ~n3416;
  assign n3436 = ~reg_controllable_BtoS_ACK8_out & ~n3435;
  assign n3437 = reg_i_StoB_REQ8_out & ~n3436;
  assign n3438 = ~reg_controllable_BtoS_ACK7_out & ~n3410;
  assign n3439 = ~reg_controllable_BtoS_ACK7_out & ~n3438;
  assign n3440 = reg_i_StoB_REQ7_out & ~n3439;
  assign n3441 = ~reg_controllable_BtoS_ACK6_out & ~n3406;
  assign n3442 = ~reg_controllable_BtoS_ACK6_out & ~n3441;
  assign n3443 = reg_i_StoB_REQ6_out & ~n3442;
  assign n3444 = ~reg_controllable_BtoS_ACK5_out & ~n3402;
  assign n3445 = ~reg_controllable_BtoS_ACK5_out & ~n3444;
  assign n3446 = reg_i_StoB_REQ5_out & ~n3445;
  assign n3447 = ~reg_controllable_BtoS_ACK4_out & ~n3398;
  assign n3448 = ~reg_controllable_BtoS_ACK4_out & ~n3447;
  assign n3449 = reg_i_StoB_REQ4_out & ~n3448;
  assign n3450 = ~reg_controllable_BtoS_ACK3_out & ~n3392;
  assign n3451 = ~reg_controllable_BtoS_ACK3_out & ~n3450;
  assign n3452 = reg_i_StoB_REQ3_out & ~n3451;
  assign n3453 = ~reg_controllable_BtoS_ACK2_out & ~n3384;
  assign n3454 = ~reg_controllable_BtoS_ACK2_out & ~n3453;
  assign n3455 = reg_i_StoB_REQ2_out & ~n3454;
  assign n3456 = ~reg_controllable_BtoS_ACK1_out & ~n377;
  assign n3457 = ~reg_controllable_BtoS_ACK1_out & ~n3456;
  assign n3458 = reg_i_StoB_REQ1_out & ~n3457;
  assign n3459 = reg_i_StoB_REQ1_out & ~n3458;
  assign n3460 = sys_fair0done_out & ~n3459;
  assign n3461 = ~n1123 & ~n3460;
  assign n3462 = sys_fair1done_out & ~n3461;
  assign n3463 = ~sys_fair1done_out & ~n379;
  assign n3464 = ~n3462 & ~n3463;
  assign n3465 = reg_stateG12_out & ~n3464;
  assign n3466 = ~n508 & ~n3465;
  assign n3467 = ~sys_fair12done_out & ~n3466;
  assign n3468 = ~n1127 & ~n3467;
  assign n3469 = sys_fair2done_out & ~n3468;
  assign n3470 = ~n513 & ~n3469;
  assign n3471 = reg_controllable_BtoS_ACK2_out & ~n3470;
  assign n3472 = ~n1432 & ~n3469;
  assign n3473 = ~reg_controllable_BtoS_ACK2_out & ~n3472;
  assign n3474 = ~n3471 & ~n3473;
  assign n3475 = ~reg_i_StoB_REQ2_out & ~n3474;
  assign n3476 = ~n3455 & ~n3475;
  assign n3477 = sys_fair3done_out & ~n3476;
  assign n3478 = ~n527 & ~n3477;
  assign n3479 = reg_controllable_BtoS_ACK3_out & ~n3478;
  assign n3480 = ~n1448 & ~n3477;
  assign n3481 = ~reg_controllable_BtoS_ACK3_out & ~n3480;
  assign n3482 = ~n3479 & ~n3481;
  assign n3483 = ~reg_i_StoB_REQ3_out & ~n3482;
  assign n3484 = ~n3452 & ~n3483;
  assign n3485 = ~reg_i_StoB_REQ4_out & ~n3484;
  assign n3486 = ~n3449 & ~n3485;
  assign n3487 = sys_fair4done_out & ~n3486;
  assign n3488 = ~n1468 & ~n3487;
  assign n3489 = ~reg_i_StoB_REQ5_out & ~n3488;
  assign n3490 = ~n3446 & ~n3489;
  assign n3491 = sys_fair5done_out & ~n3490;
  assign n3492 = ~n1481 & ~n3491;
  assign n3493 = ~reg_i_StoB_REQ6_out & ~n3492;
  assign n3494 = ~n3443 & ~n3493;
  assign n3495 = sys_fair6done_out & ~n3494;
  assign n3496 = ~n1494 & ~n3495;
  assign n3497 = ~reg_i_StoB_REQ7_out & ~n3496;
  assign n3498 = ~n3440 & ~n3497;
  assign n3499 = sys_fair7done_out & ~n3498;
  assign n3500 = ~n1507 & ~n3499;
  assign n3501 = sys_fair8done_out & ~n3500;
  assign n3502 = ~n613 & ~n3501;
  assign n3503 = reg_controllable_BtoS_ACK8_out & ~n3502;
  assign n3504 = ~n1516 & ~n3501;
  assign n3505 = ~reg_controllable_BtoS_ACK8_out & ~n3504;
  assign n3506 = ~n3503 & ~n3505;
  assign n3507 = ~reg_i_StoB_REQ8_out & ~n3506;
  assign n3508 = ~n3437 & ~n3507;
  assign n3509 = ~reg_i_StoB_REQ10_out & ~n3508;
  assign n3510 = ~n3434 & ~n3509;
  assign n3511 = sys_fair10done_out & ~n3510;
  assign n3512 = ~n1536 & ~n3511;
  assign n3513 = sys_fair11done_out & ~n3512;
  assign n3514 = ~n648 & ~n3513;
  assign n3515 = reg_controllable_BtoS_ACK11_out & ~n3514;
  assign n3516 = ~n1547 & ~n3513;
  assign n3517 = ~reg_controllable_BtoS_ACK11_out & ~n3516;
  assign n3518 = ~n3515 & ~n3517;
  assign n3519 = ~reg_i_StoB_REQ11_out & ~n3518;
  assign n3520 = ~n3431 & ~n3519;
  assign n3521 = sys_fair9done_out & ~n3520;
  assign n3522 = ~n1262 & ~n3521;
  assign n3523 = fair_cnt<1>_out  & ~n3522;
  assign n3524 = ~n674 & ~n3523;
  assign n3525 = fair_cnt<0>_out  & ~n3524;
  assign n3526 = ~n677 & ~n3525;
  assign n3527 = ~env_fair1done_out & ~n3526;
  assign n3528 = ~n1569 & ~n3527;
  assign n3529 = env_fair0done_out & ~n3528;
  assign n3530 = ~n1559 & ~n3529;
  assign n3531 = ~reg_stateG7_0_out & ~n3530;
  assign n3532 = ~reg_stateG7_0_out & ~n3531;
  assign n3533 = reg_nstateG7_1_out & ~n3532;
  assign n3534 = ~reg_nstateG7_1_out & ~n3530;
  assign n3535 = ~n3533 & ~n3534;
  assign n3536 = ~reg_controllable_BtoR_REQ1_out & ~n3535;
  assign n3537 = ~reg_controllable_BtoR_REQ1_out & ~n3536;
  assign n3538 = reg_controllable_BtoR_REQ0_out & ~n3537;
  assign n3539 = reg_controllable_BtoR_REQ0_out & ~n3538;
  assign n3540 = ~reg_i_RtoB_ACK1_out & ~n3539;
  assign n3541 = ~reg_i_RtoB_ACK1_out & ~n3540;
  assign n3542 = reg_i_RtoB_ACK0_out & ~n3541;
  assign n3543 = env_fair0done_out & ~n1571;
  assign n3544 = env_fair1done_out & ~n3526;
  assign n3545 = ~n1570 & ~n3544;
  assign n3546 = ~env_fair0done_out & ~n3545;
  assign n3547 = ~n3543 & ~n3546;
  assign n3548 = reg_nstateG7_1_out & ~n3547;
  assign n3549 = ~reg_stateG7_0_out & ~n3547;
  assign n3550 = ~reg_stateG7_0_out & ~n3549;
  assign n3551 = ~reg_nstateG7_1_out & ~n3550;
  assign n3552 = ~n3548 & ~n3551;
  assign n3553 = reg_controllable_BtoR_REQ1_out & ~n3552;
  assign n3554 = reg_controllable_BtoR_REQ1_out & ~n3553;
  assign n3555 = ~reg_controllable_BtoR_REQ0_out & ~n3554;
  assign n3556 = ~reg_controllable_BtoR_REQ0_out & ~n3555;
  assign n3557 = reg_i_RtoB_ACK1_out & ~n3556;
  assign n3558 = ~n2565 & ~n2598;
  assign n3559 = ~reg_controllable_BtoR_REQ1_out & ~n3558;
  assign n3560 = ~n2562 & ~n3559;
  assign n3561 = ~reg_controllable_BtoR_REQ0_out & ~n3560;
  assign n3562 = ~n2580 & ~n3561;
  assign n3563 = ~reg_i_RtoB_ACK1_out & ~n3562;
  assign n3564 = ~n3557 & ~n3563;
  assign n3565 = ~reg_i_RtoB_ACK0_out & ~n3564;
  assign n3566 = ~n3542 & ~n3565;
  assign n3567 = ~reg_i_StoB_REQ9_out & ~n3566;
  assign n3568 = ~n3381 & ~n3567;
  assign n3569 = reg_controllable_BtoS_ACK9_out & ~n3568;
  assign n3570 = reg_controllable_BtoS_ACK11_out & ~n3428;
  assign n3571 = ~n2884 & ~n3427;
  assign n3572 = ~reg_controllable_BtoS_ACK11_out & ~n3571;
  assign n3573 = ~n3570 & ~n3572;
  assign n3574 = ~reg_i_StoB_REQ11_out & ~n3573;
  assign n3575 = ~n1425 & ~n3574;
  assign n3576 = sys_fair9done_out & ~n3575;
  assign n3577 = ~n890 & ~n3576;
  assign n3578 = fair_cnt<1>_out  & ~n3577;
  assign n3579 = ~n365 & ~n3578;
  assign n3580 = fair_cnt<0>_out  & ~n3579;
  assign n3581 = ~n368 & ~n3580;
  assign n3582 = ~env_fair1done_out & ~n3581;
  assign n3583 = ~n2906 & ~n3582;
  assign n3584 = env_fair0done_out & ~n3583;
  assign n3585 = ~n2896 & ~n3584;
  assign n3586 = ~reg_stateG7_0_out & ~n3585;
  assign n3587 = ~reg_stateG7_0_out & ~n3586;
  assign n3588 = reg_nstateG7_1_out & ~n3587;
  assign n3589 = ~reg_nstateG7_1_out & ~n3585;
  assign n3590 = ~n3588 & ~n3589;
  assign n3591 = ~reg_controllable_BtoR_REQ1_out & ~n3590;
  assign n3592 = ~reg_controllable_BtoR_REQ1_out & ~n3591;
  assign n3593 = reg_controllable_BtoR_REQ0_out & ~n3592;
  assign n3594 = reg_controllable_BtoR_REQ0_out & ~n3593;
  assign n3595 = ~reg_i_RtoB_ACK1_out & ~n3594;
  assign n3596 = ~reg_i_RtoB_ACK1_out & ~n3595;
  assign n3597 = reg_i_RtoB_ACK0_out & ~n3596;
  assign n3598 = env_fair0done_out & ~n2908;
  assign n3599 = env_fair1done_out & ~n3581;
  assign n3600 = ~n2907 & ~n3599;
  assign n3601 = ~env_fair0done_out & ~n3600;
  assign n3602 = ~n3598 & ~n3601;
  assign n3603 = reg_nstateG7_1_out & ~n3602;
  assign n3604 = ~reg_stateG7_0_out & ~n3602;
  assign n3605 = ~reg_stateG7_0_out & ~n3604;
  assign n3606 = ~reg_nstateG7_1_out & ~n3605;
  assign n3607 = ~n3603 & ~n3606;
  assign n3608 = reg_controllable_BtoR_REQ1_out & ~n3607;
  assign n3609 = reg_controllable_BtoR_REQ1_out & ~n3608;
  assign n3610 = ~reg_controllable_BtoR_REQ0_out & ~n3609;
  assign n3611 = ~reg_controllable_BtoR_REQ0_out & ~n3610;
  assign n3612 = reg_i_RtoB_ACK1_out & ~n3611;
  assign n3613 = ~n3313 & ~n3612;
  assign n3614 = ~reg_i_RtoB_ACK0_out & ~n3613;
  assign n3615 = ~n3597 & ~n3614;
  assign n3616 = reg_i_StoB_REQ9_out & ~n3615;
  assign n3617 = ~n3086 & ~n3521;
  assign n3618 = fair_cnt<1>_out  & ~n3617;
  assign n3619 = ~n674 & ~n3618;
  assign n3620 = fair_cnt<0>_out  & ~n3619;
  assign n3621 = ~n677 & ~n3620;
  assign n3622 = ~env_fair1done_out & ~n3621;
  assign n3623 = ~n3102 & ~n3622;
  assign n3624 = env_fair0done_out & ~n3623;
  assign n3625 = ~n3092 & ~n3624;
  assign n3626 = ~reg_stateG7_0_out & ~n3625;
  assign n3627 = ~reg_stateG7_0_out & ~n3626;
  assign n3628 = reg_nstateG7_1_out & ~n3627;
  assign n3629 = ~reg_nstateG7_1_out & ~n3625;
  assign n3630 = ~n3628 & ~n3629;
  assign n3631 = ~reg_controllable_BtoR_REQ1_out & ~n3630;
  assign n3632 = ~reg_controllable_BtoR_REQ1_out & ~n3631;
  assign n3633 = reg_controllable_BtoR_REQ0_out & ~n3632;
  assign n3634 = reg_controllable_BtoR_REQ0_out & ~n3633;
  assign n3635 = ~reg_i_RtoB_ACK1_out & ~n3634;
  assign n3636 = ~reg_i_RtoB_ACK1_out & ~n3635;
  assign n3637 = reg_i_RtoB_ACK0_out & ~n3636;
  assign n3638 = env_fair0done_out & ~n3104;
  assign n3639 = env_fair1done_out & ~n3621;
  assign n3640 = ~n3103 & ~n3639;
  assign n3641 = ~env_fair0done_out & ~n3640;
  assign n3642 = ~n3638 & ~n3641;
  assign n3643 = reg_nstateG7_1_out & ~n3642;
  assign n3644 = ~reg_stateG7_0_out & ~n3642;
  assign n3645 = ~reg_stateG7_0_out & ~n3644;
  assign n3646 = ~reg_nstateG7_1_out & ~n3645;
  assign n3647 = ~n3643 & ~n3646;
  assign n3648 = reg_controllable_BtoR_REQ1_out & ~n3647;
  assign n3649 = reg_controllable_BtoR_REQ1_out & ~n3648;
  assign n3650 = ~reg_controllable_BtoR_REQ0_out & ~n3649;
  assign n3651 = ~reg_controllable_BtoR_REQ0_out & ~n3650;
  assign n3652 = reg_i_RtoB_ACK1_out & ~n3651;
  assign n3653 = ~n3168 & ~n3194;
  assign n3654 = ~reg_controllable_BtoR_REQ1_out & ~n3653;
  assign n3655 = ~n3165 & ~n3654;
  assign n3656 = ~reg_controllable_BtoR_REQ0_out & ~n3655;
  assign n3657 = ~n3183 & ~n3656;
  assign n3658 = ~reg_i_RtoB_ACK1_out & ~n3657;
  assign n3659 = ~n3652 & ~n3658;
  assign n3660 = ~reg_i_RtoB_ACK0_out & ~n3659;
  assign n3661 = ~n3637 & ~n3660;
  assign n3662 = ~reg_i_StoB_REQ9_out & ~n3661;
  assign n3663 = ~n3616 & ~n3662;
  assign n3664 = ~reg_controllable_BtoS_ACK9_out & ~n3663;
  assign n3665 = ~n3569 & ~n3664;
  assign n3666 = ~reg_i_nEMPTY_out & ~n3665;
  assign n3667 = ~n3371 & ~n3666;
  assign n3668 = ~reg_i_FULL_out & ~n3667;
  assign n3669 = ~n3210 & ~n3668;
  assign n3670 = reg_controllable_DEQ_out & ~n3669;
  assign n3671 = ~n431 & ~n890;
  assign n3672 = fair_cnt<1>_out  & ~n3671;
  assign n3673 = ~n365 & ~n3672;
  assign n3674 = ~fair_cnt<0>_out  & ~n3673;
  assign n3675 = ~n367 & ~n3674;
  assign n3676 = ~reg_controllable_BtoR_REQ1_out & ~n3675;
  assign n3677 = ~reg_controllable_BtoR_REQ1_out & ~n3676;
  assign n3678 = ~reg_controllable_BtoR_REQ0_out & ~n3677;
  assign n3679 = ~reg_controllable_BtoR_REQ0_out & ~n3678;
  assign n3680 = reg_i_RtoB_ACK1_out & ~n3679;
  assign n3681 = ~fair_cnt<1>_out  & ~n3671;
  assign n3682 = ~n359 & ~n3681;
  assign n3683 = fair_cnt<0>_out  & ~n3682;
  assign n3684 = ~sys_fair0done_out & ~n381;
  assign n3685 = sys_fair1done_out & ~n3684;
  assign n3686 = ~n384 & ~n3685;
  assign n3687 = reg_stateG12_out & ~n3686;
  assign n3688 = ~n131 & ~n3687;
  assign n3689 = ~sys_fair12done_out & ~n3688;
  assign n3690 = ~n376 & ~n3689;
  assign n3691 = sys_fair2done_out & ~n3690;
  assign n3692 = ~n143 & ~n3691;
  assign n3693 = ~reg_controllable_BtoS_ACK2_out & ~n3692;
  assign n3694 = ~reg_controllable_BtoS_ACK2_out & ~n3693;
  assign n3695 = reg_i_StoB_REQ2_out & ~n3694;
  assign n3696 = ~reg_i_StoB_REQ2_out & ~n3692;
  assign n3697 = ~n3695 & ~n3696;
  assign n3698 = sys_fair3done_out & ~n3697;
  assign n3699 = ~n169 & ~n3698;
  assign n3700 = ~reg_controllable_BtoS_ACK3_out & ~n3699;
  assign n3701 = ~reg_controllable_BtoS_ACK3_out & ~n3700;
  assign n3702 = reg_i_StoB_REQ3_out & ~n3701;
  assign n3703 = ~reg_i_StoB_REQ3_out & ~n3699;
  assign n3704 = ~n3702 & ~n3703;
  assign n3705 = ~reg_controllable_BtoS_ACK4_out & ~n3704;
  assign n3706 = ~reg_controllable_BtoS_ACK4_out & ~n3705;
  assign n3707 = reg_i_StoB_REQ4_out & ~n3706;
  assign n3708 = ~reg_i_StoB_REQ4_out & ~n3704;
  assign n3709 = ~n3707 & ~n3708;
  assign n3710 = sys_fair4done_out & ~n3709;
  assign n3711 = ~n401 & ~n3710;
  assign n3712 = ~reg_controllable_BtoS_ACK5_out & ~n3711;
  assign n3713 = ~reg_controllable_BtoS_ACK5_out & ~n3712;
  assign n3714 = reg_i_StoB_REQ5_out & ~n3713;
  assign n3715 = ~reg_i_StoB_REQ5_out & ~n3711;
  assign n3716 = ~n3714 & ~n3715;
  assign n3717 = sys_fair5done_out & ~n3716;
  assign n3718 = ~n406 & ~n3717;
  assign n3719 = ~reg_controllable_BtoS_ACK6_out & ~n3718;
  assign n3720 = ~reg_controllable_BtoS_ACK6_out & ~n3719;
  assign n3721 = reg_i_StoB_REQ6_out & ~n3720;
  assign n3722 = ~reg_i_StoB_REQ6_out & ~n3718;
  assign n3723 = ~n3721 & ~n3722;
  assign n3724 = sys_fair6done_out & ~n3723;
  assign n3725 = ~n411 & ~n3724;
  assign n3726 = ~reg_controllable_BtoS_ACK7_out & ~n3725;
  assign n3727 = ~reg_controllable_BtoS_ACK7_out & ~n3726;
  assign n3728 = reg_i_StoB_REQ7_out & ~n3727;
  assign n3729 = ~reg_i_StoB_REQ7_out & ~n3725;
  assign n3730 = ~n3728 & ~n3729;
  assign n3731 = sys_fair7done_out & ~n3730;
  assign n3732 = ~n416 & ~n3731;
  assign n3733 = sys_fair8done_out & ~n3732;
  assign n3734 = ~n291 & ~n3733;
  assign n3735 = ~reg_controllable_BtoS_ACK8_out & ~n3734;
  assign n3736 = ~reg_controllable_BtoS_ACK8_out & ~n3735;
  assign n3737 = reg_i_StoB_REQ8_out & ~n3736;
  assign n3738 = ~reg_i_StoB_REQ8_out & ~n3734;
  assign n3739 = ~n3737 & ~n3738;
  assign n3740 = ~reg_controllable_BtoS_ACK10_out & ~n3739;
  assign n3741 = ~reg_controllable_BtoS_ACK10_out & ~n3740;
  assign n3742 = reg_i_StoB_REQ10_out & ~n3741;
  assign n3743 = ~reg_i_StoB_REQ10_out & ~n3739;
  assign n3744 = ~n3742 & ~n3743;
  assign n3745 = sys_fair10done_out & ~n3744;
  assign n3746 = ~n425 & ~n3745;
  assign n3747 = sys_fair11done_out & ~n3746;
  assign n3748 = ~n341 & ~n3747;
  assign n3749 = ~reg_controllable_BtoS_ACK11_out & ~n3748;
  assign n3750 = ~reg_controllable_BtoS_ACK11_out & ~n3749;
  assign n3751 = reg_i_StoB_REQ11_out & ~n3750;
  assign n3752 = ~reg_i_StoB_REQ11_out & ~n3748;
  assign n3753 = ~n3751 & ~n3752;
  assign n3754 = sys_fair9done_out & ~n3753;
  assign n3755 = ~n890 & ~n3754;
  assign n3756 = fair_cnt<1>_out  & ~n3755;
  assign n3757 = ~n365 & ~n3756;
  assign n3758 = ~fair_cnt<0>_out  & ~n3757;
  assign n3759 = ~n3683 & ~n3758;
  assign n3760 = env_fair1done_out & ~n3759;
  assign n3761 = ~n470 & ~n3754;
  assign n3762 = fair_cnt<1>_out  & ~n3761;
  assign n3763 = ~n3681 & ~n3762;
  assign n3764 = fair_cnt<0>_out  & ~n3763;
  assign n3765 = ~n3674 & ~n3764;
  assign n3766 = ~env_fair1done_out & ~n3765;
  assign n3767 = ~n3760 & ~n3766;
  assign n3768 = env_fair0done_out & ~n3767;
  assign n3769 = fair_cnt<0>_out  & ~n3757;
  assign n3770 = ~n3674 & ~n3769;
  assign n3771 = ~env_fair0done_out & ~n3770;
  assign n3772 = ~n3768 & ~n3771;
  assign n3773 = ~reg_stateG7_0_out & ~n3772;
  assign n3774 = ~reg_stateG7_0_out & ~n3773;
  assign n3775 = reg_nstateG7_1_out & ~n3774;
  assign n3776 = ~reg_nstateG7_1_out & ~n3772;
  assign n3777 = ~n3775 & ~n3776;
  assign n3778 = ~reg_controllable_BtoR_REQ1_out & ~n3777;
  assign n3779 = ~reg_controllable_BtoR_REQ1_out & ~n3778;
  assign n3780 = reg_controllable_BtoR_REQ0_out & ~n3779;
  assign n3781 = sys_fair12done_out & ~n379;
  assign n3782 = ~sys_fair0done_out & ~n1123;
  assign n3783 = sys_fair1done_out & ~n3782;
  assign n3784 = ~n3463 & ~n3783;
  assign n3785 = reg_stateG12_out & ~n3784;
  assign n3786 = ~n508 & ~n3785;
  assign n3787 = ~sys_fair12done_out & ~n3786;
  assign n3788 = ~n3781 & ~n3787;
  assign n3789 = sys_fair2done_out & ~n3788;
  assign n3790 = ~n513 & ~n3789;
  assign n3791 = ~reg_i_StoB_REQ2_out & ~n3790;
  assign n3792 = ~n3695 & ~n3791;
  assign n3793 = sys_fair3done_out & ~n3792;
  assign n3794 = ~n527 & ~n3793;
  assign n3795 = ~reg_i_StoB_REQ3_out & ~n3794;
  assign n3796 = ~n3702 & ~n3795;
  assign n3797 = ~reg_i_StoB_REQ4_out & ~n3796;
  assign n3798 = ~n3707 & ~n3797;
  assign n3799 = sys_fair4done_out & ~n3798;
  assign n3800 = ~sys_fair4done_out & ~n566;
  assign n3801 = ~n3799 & ~n3800;
  assign n3802 = ~reg_i_StoB_REQ5_out & ~n3801;
  assign n3803 = ~n3714 & ~n3802;
  assign n3804 = sys_fair5done_out & ~n3803;
  assign n3805 = ~sys_fair5done_out & ~n582;
  assign n3806 = ~n3804 & ~n3805;
  assign n3807 = ~reg_i_StoB_REQ6_out & ~n3806;
  assign n3808 = ~n3721 & ~n3807;
  assign n3809 = sys_fair6done_out & ~n3808;
  assign n3810 = ~sys_fair6done_out & ~n598;
  assign n3811 = ~n3809 & ~n3810;
  assign n3812 = ~reg_i_StoB_REQ7_out & ~n3811;
  assign n3813 = ~n3728 & ~n3812;
  assign n3814 = sys_fair7done_out & ~n3813;
  assign n3815 = ~sys_fair7done_out & ~n612;
  assign n3816 = ~n3814 & ~n3815;
  assign n3817 = sys_fair8done_out & ~n3816;
  assign n3818 = ~n613 & ~n3817;
  assign n3819 = ~reg_i_StoB_REQ8_out & ~n3818;
  assign n3820 = ~n3737 & ~n3819;
  assign n3821 = ~reg_i_StoB_REQ10_out & ~n3820;
  assign n3822 = ~n3742 & ~n3821;
  assign n3823 = sys_fair10done_out & ~n3822;
  assign n3824 = ~sys_fair10done_out & ~n647;
  assign n3825 = ~n3823 & ~n3824;
  assign n3826 = sys_fair11done_out & ~n3825;
  assign n3827 = ~n648 & ~n3826;
  assign n3828 = ~reg_i_StoB_REQ11_out & ~n3827;
  assign n3829 = ~n3751 & ~n3828;
  assign n3830 = sys_fair9done_out & ~n3829;
  assign n3831 = ~n1262 & ~n3830;
  assign n3832 = fair_cnt<1>_out  & ~n3831;
  assign n3833 = ~n674 & ~n3832;
  assign n3834 = ~fair_cnt<0>_out  & ~n3833;
  assign n3835 = ~n676 & ~n3834;
  assign n3836 = env_fair1done_out & ~n3835;
  assign n3837 = ~env_fair1done_out & ~n678;
  assign n3838 = ~n3836 & ~n3837;
  assign n3839 = reg_nstateG7_1_out & ~n3838;
  assign n3840 = ~reg_stateG7_0_out & ~n3838;
  assign n3841 = ~reg_stateG7_0_out & ~n3840;
  assign n3842 = ~reg_nstateG7_1_out & ~n3841;
  assign n3843 = ~n3839 & ~n3842;
  assign n3844 = reg_controllable_BtoR_REQ1_out & ~n3843;
  assign n3845 = env_fair1done_out & ~n3675;
  assign n3846 = ~n365 & ~n3762;
  assign n3847 = fair_cnt<0>_out  & ~n3846;
  assign n3848 = ~n3674 & ~n3847;
  assign n3849 = ~env_fair1done_out & ~n3848;
  assign n3850 = ~n3845 & ~n3849;
  assign n3851 = reg_nstateG7_1_out & ~n3850;
  assign n3852 = ~reg_nstateG7_1_out & ~n3675;
  assign n3853 = ~n3851 & ~n3852;
  assign n3854 = ~reg_controllable_BtoR_REQ1_out & ~n3853;
  assign n3855 = ~n3844 & ~n3854;
  assign n3856 = ~reg_controllable_BtoR_REQ0_out & ~n3855;
  assign n3857 = ~n3780 & ~n3856;
  assign n3858 = ~reg_i_RtoB_ACK1_out & ~n3857;
  assign n3859 = ~n3680 & ~n3858;
  assign n3860 = reg_i_RtoB_ACK0_out & ~n3859;
  assign n3861 = env_fair0done_out & ~n3835;
  assign n3862 = ~env_fair0done_out & ~n678;
  assign n3863 = ~n3861 & ~n3862;
  assign n3864 = ~reg_stateG7_0_out & ~n3863;
  assign n3865 = ~reg_stateG7_0_out & ~n3864;
  assign n3866 = reg_nstateG7_1_out & ~n3865;
  assign n3867 = ~reg_nstateG7_1_out & ~n3863;
  assign n3868 = ~n3866 & ~n3867;
  assign n3869 = ~reg_controllable_BtoR_REQ1_out & ~n3868;
  assign n3870 = ~reg_controllable_BtoR_REQ1_out & ~n3869;
  assign n3871 = reg_controllable_BtoR_REQ0_out & ~n3870;
  assign n3872 = ~env_fair1done_out & ~n3770;
  assign n3873 = ~n3760 & ~n3872;
  assign n3874 = env_fair0done_out & ~n3873;
  assign n3875 = env_fair1done_out & ~n3765;
  assign n3876 = ~n3872 & ~n3875;
  assign n3877 = ~env_fair0done_out & ~n3876;
  assign n3878 = ~n3874 & ~n3877;
  assign n3879 = reg_nstateG7_1_out & ~n3878;
  assign n3880 = ~reg_stateG7_0_out & ~n3878;
  assign n3881 = ~reg_stateG7_0_out & ~n3880;
  assign n3882 = ~reg_nstateG7_1_out & ~n3881;
  assign n3883 = ~n3879 & ~n3882;
  assign n3884 = reg_controllable_BtoR_REQ1_out & ~n3883;
  assign n3885 = reg_nstateG7_1_out & ~n3675;
  assign n3886 = env_fair0done_out & ~n3675;
  assign n3887 = ~env_fair0done_out & ~n3848;
  assign n3888 = ~n3886 & ~n3887;
  assign n3889 = ~reg_nstateG7_1_out & ~n3888;
  assign n3890 = ~n3885 & ~n3889;
  assign n3891 = ~reg_controllable_BtoR_REQ1_out & ~n3890;
  assign n3892 = ~n3884 & ~n3891;
  assign n3893 = ~reg_controllable_BtoR_REQ0_out & ~n3892;
  assign n3894 = ~n3871 & ~n3893;
  assign n3895 = reg_i_RtoB_ACK1_out & ~n3894;
  assign n3896 = ~fair_cnt<1>_out  & ~n3755;
  assign n3897 = ~n359 & ~n3896;
  assign n3898 = fair_cnt<0>_out  & ~n3897;
  assign n3899 = ~n347 & ~n890;
  assign n3900 = fair_cnt<1>_out  & ~n3899;
  assign n3901 = ~n3681 & ~n3900;
  assign n3902 = ~fair_cnt<0>_out  & ~n3901;
  assign n3903 = ~n3898 & ~n3902;
  assign n3904 = env_fair0done_out & ~n3903;
  assign n3905 = ~env_fair0done_out & ~n3759;
  assign n3906 = ~n3904 & ~n3905;
  assign n3907 = ~reg_stateG7_0_out & ~n3906;
  assign n3908 = ~reg_stateG7_0_out & ~n3907;
  assign n3909 = reg_nstateG7_1_out & ~n3908;
  assign n3910 = ~reg_nstateG7_1_out & ~n3906;
  assign n3911 = ~n3909 & ~n3910;
  assign n3912 = ~reg_controllable_BtoR_REQ1_out & ~n3911;
  assign n3913 = ~reg_controllable_BtoR_REQ1_out & ~n3912;
  assign n3914 = reg_controllable_BtoR_REQ0_out & ~n3913;
  assign n3915 = env_fair1done_out & ~n3903;
  assign n3916 = ~env_fair1done_out & ~n3759;
  assign n3917 = ~n3915 & ~n3916;
  assign n3918 = reg_nstateG7_1_out & ~n3917;
  assign n3919 = ~reg_stateG7_0_out & ~n3917;
  assign n3920 = ~reg_stateG7_0_out & ~n3919;
  assign n3921 = ~reg_nstateG7_1_out & ~n3920;
  assign n3922 = ~n3918 & ~n3921;
  assign n3923 = reg_controllable_BtoR_REQ1_out & ~n3922;
  assign n3924 = fair_cnt<0>_out  & ~n3901;
  assign n3925 = ~n3758 & ~n3924;
  assign n3926 = ~env_fair1done_out & ~n3925;
  assign n3927 = ~n3915 & ~n3926;
  assign n3928 = reg_nstateG7_1_out & ~n3927;
  assign n3929 = ~env_fair0done_out & ~n3925;
  assign n3930 = ~n3904 & ~n3929;
  assign n3931 = ~reg_nstateG7_1_out & ~n3930;
  assign n3932 = ~n3928 & ~n3931;
  assign n3933 = ~reg_controllable_BtoR_REQ1_out & ~n3932;
  assign n3934 = ~n3923 & ~n3933;
  assign n3935 = ~reg_controllable_BtoR_REQ0_out & ~n3934;
  assign n3936 = ~n3914 & ~n3935;
  assign n3937 = ~reg_i_RtoB_ACK1_out & ~n3936;
  assign n3938 = ~n3895 & ~n3937;
  assign n3939 = ~reg_i_RtoB_ACK0_out & ~n3938;
  assign n3940 = ~n3860 & ~n3939;
  assign n3941 = reg_i_StoB_REQ9_out & ~n3940;
  assign n3942 = ~reg_controllable_BtoS_ACK11_out & ~n428;
  assign n3943 = ~reg_controllable_BtoS_ACK11_out & ~n3942;
  assign n3944 = reg_i_StoB_REQ11_out & ~n3943;
  assign n3945 = ~reg_controllable_BtoS_ACK10_out & ~n421;
  assign n3946 = ~reg_controllable_BtoS_ACK10_out & ~n3945;
  assign n3947 = reg_i_StoB_REQ10_out & ~n3946;
  assign n3948 = ~reg_controllable_BtoS_ACK8_out & ~n419;
  assign n3949 = ~reg_controllable_BtoS_ACK8_out & ~n3948;
  assign n3950 = reg_i_StoB_REQ8_out & ~n3949;
  assign n3951 = ~reg_controllable_BtoS_ACK7_out & ~n412;
  assign n3952 = ~reg_controllable_BtoS_ACK7_out & ~n3951;
  assign n3953 = reg_i_StoB_REQ7_out & ~n3952;
  assign n3954 = ~reg_controllable_BtoS_ACK6_out & ~n407;
  assign n3955 = ~reg_controllable_BtoS_ACK6_out & ~n3954;
  assign n3956 = reg_i_StoB_REQ6_out & ~n3955;
  assign n3957 = ~reg_controllable_BtoS_ACK5_out & ~n402;
  assign n3958 = ~reg_controllable_BtoS_ACK5_out & ~n3957;
  assign n3959 = reg_i_StoB_REQ5_out & ~n3958;
  assign n3960 = ~reg_controllable_BtoS_ACK4_out & ~n397;
  assign n3961 = ~reg_controllable_BtoS_ACK4_out & ~n3960;
  assign n3962 = reg_i_StoB_REQ4_out & ~n3961;
  assign n3963 = ~reg_controllable_BtoS_ACK3_out & ~n395;
  assign n3964 = ~reg_controllable_BtoS_ACK3_out & ~n3963;
  assign n3965 = reg_i_StoB_REQ3_out & ~n3964;
  assign n3966 = ~reg_controllable_BtoS_ACK2_out & ~n391;
  assign n3967 = ~reg_controllable_BtoS_ACK2_out & ~n3966;
  assign n3968 = reg_i_StoB_REQ2_out & ~n3967;
  assign n3969 = ~n3467 & ~n3781;
  assign n3970 = sys_fair2done_out & ~n3969;
  assign n3971 = ~n513 & ~n3970;
  assign n3972 = ~reg_i_StoB_REQ2_out & ~n3971;
  assign n3973 = ~n3968 & ~n3972;
  assign n3974 = sys_fair3done_out & ~n3973;
  assign n3975 = ~n527 & ~n3974;
  assign n3976 = ~reg_i_StoB_REQ3_out & ~n3975;
  assign n3977 = ~n3965 & ~n3976;
  assign n3978 = ~reg_i_StoB_REQ4_out & ~n3977;
  assign n3979 = ~n3962 & ~n3978;
  assign n3980 = sys_fair4done_out & ~n3979;
  assign n3981 = ~n3800 & ~n3980;
  assign n3982 = ~reg_i_StoB_REQ5_out & ~n3981;
  assign n3983 = ~n3959 & ~n3982;
  assign n3984 = sys_fair5done_out & ~n3983;
  assign n3985 = ~n3805 & ~n3984;
  assign n3986 = ~reg_i_StoB_REQ6_out & ~n3985;
  assign n3987 = ~n3956 & ~n3986;
  assign n3988 = sys_fair6done_out & ~n3987;
  assign n3989 = ~n3810 & ~n3988;
  assign n3990 = ~reg_i_StoB_REQ7_out & ~n3989;
  assign n3991 = ~n3953 & ~n3990;
  assign n3992 = sys_fair7done_out & ~n3991;
  assign n3993 = ~n3815 & ~n3992;
  assign n3994 = sys_fair8done_out & ~n3993;
  assign n3995 = ~n613 & ~n3994;
  assign n3996 = ~reg_i_StoB_REQ8_out & ~n3995;
  assign n3997 = ~n3950 & ~n3996;
  assign n3998 = ~reg_i_StoB_REQ10_out & ~n3997;
  assign n3999 = ~n3947 & ~n3998;
  assign n4000 = sys_fair10done_out & ~n3999;
  assign n4001 = ~n3824 & ~n4000;
  assign n4002 = sys_fair11done_out & ~n4001;
  assign n4003 = ~n648 & ~n4002;
  assign n4004 = ~reg_i_StoB_REQ11_out & ~n4003;
  assign n4005 = ~n3944 & ~n4004;
  assign n4006 = sys_fair9done_out & ~n4005;
  assign n4007 = ~n1262 & ~n4006;
  assign n4008 = fair_cnt<1>_out  & ~n4007;
  assign n4009 = ~n674 & ~n4008;
  assign n4010 = ~fair_cnt<0>_out  & ~n4009;
  assign n4011 = ~n1266 & ~n4010;
  assign n4012 = env_fair0done_out & ~n4011;
  assign n4013 = ~env_fair0done_out & ~n1267;
  assign n4014 = ~n4012 & ~n4013;
  assign n4015 = ~reg_stateG7_0_out & ~n4014;
  assign n4016 = ~reg_stateG7_0_out & ~n4015;
  assign n4017 = reg_nstateG7_1_out & ~n4016;
  assign n4018 = ~reg_nstateG7_1_out & ~n4014;
  assign n4019 = ~n4017 & ~n4018;
  assign n4020 = ~reg_controllable_BtoR_REQ1_out & ~n4019;
  assign n4021 = ~reg_controllable_BtoR_REQ1_out & ~n4020;
  assign n4022 = reg_controllable_BtoR_REQ0_out & ~n4021;
  assign n4023 = env_fair1done_out & ~n4011;
  assign n4024 = ~env_fair1done_out & ~n1267;
  assign n4025 = ~n4023 & ~n4024;
  assign n4026 = reg_nstateG7_1_out & ~n4025;
  assign n4027 = ~reg_stateG7_0_out & ~n4025;
  assign n4028 = ~reg_stateG7_0_out & ~n4027;
  assign n4029 = ~reg_nstateG7_1_out & ~n4028;
  assign n4030 = ~n4026 & ~n4029;
  assign n4031 = reg_controllable_BtoR_REQ1_out & ~n4030;
  assign n4032 = reg_controllable_BtoS_ACK11_out & ~n428;
  assign n4033 = ~n1962 & ~n4032;
  assign n4034 = reg_i_StoB_REQ11_out & ~n4033;
  assign n4035 = reg_controllable_BtoS_ACK8_out & ~n419;
  assign n4036 = ~n1903 & ~n4035;
  assign n4037 = reg_i_StoB_REQ8_out & ~n4036;
  assign n4038 = reg_controllable_BtoS_ACK3_out & ~n395;
  assign n4039 = ~n1717 & ~n4038;
  assign n4040 = reg_i_StoB_REQ3_out & ~n4039;
  assign n4041 = reg_controllable_BtoS_ACK2_out & ~n391;
  assign n4042 = ~n1671 & ~n4041;
  assign n4043 = reg_i_StoB_REQ2_out & ~n4042;
  assign n4044 = sys_fair12done_out & n1587;
  assign n4045 = ~n2213 & ~n2219;
  assign n4046 = sys_fair1done_out & ~n4045;
  assign n4047 = ~sys_fair1done_out & n1587;
  assign n4048 = ~n4046 & ~n4047;
  assign n4049 = reg_stateG12_out & ~n4048;
  assign n4050 = ~n1614 & ~n4049;
  assign n4051 = ~sys_fair12done_out & ~n4050;
  assign n4052 = ~n4044 & ~n4051;
  assign n4053 = sys_fair2done_out & ~n4052;
  assign n4054 = ~n1643 & ~n4053;
  assign n4055 = ~reg_i_StoB_REQ2_out & ~n4054;
  assign n4056 = ~n4043 & ~n4055;
  assign n4057 = sys_fair3done_out & ~n4056;
  assign n4058 = ~n1676 & ~n4057;
  assign n4059 = ~reg_i_StoB_REQ3_out & ~n4058;
  assign n4060 = ~n4040 & ~n4059;
  assign n4061 = ~reg_i_StoB_REQ4_out & ~n4060;
  assign n4062 = ~n2196 & ~n4061;
  assign n4063 = sys_fair4done_out & ~n4062;
  assign n4064 = ~sys_fair4done_out & ~n1762;
  assign n4065 = ~n4063 & ~n4064;
  assign n4066 = ~reg_i_StoB_REQ5_out & ~n4065;
  assign n4067 = ~n2193 & ~n4066;
  assign n4068 = sys_fair5done_out & ~n4067;
  assign n4069 = ~sys_fair5done_out & ~n1798;
  assign n4070 = ~n4068 & ~n4069;
  assign n4071 = ~reg_i_StoB_REQ6_out & ~n4070;
  assign n4072 = ~n2190 & ~n4071;
  assign n4073 = sys_fair6done_out & ~n4072;
  assign n4074 = ~sys_fair6done_out & ~n1834;
  assign n4075 = ~n4073 & ~n4074;
  assign n4076 = ~reg_i_StoB_REQ7_out & ~n4075;
  assign n4077 = ~n2187 & ~n4076;
  assign n4078 = sys_fair7done_out & ~n4077;
  assign n4079 = ~sys_fair7done_out & ~n1866;
  assign n4080 = ~n4078 & ~n4079;
  assign n4081 = sys_fair8done_out & ~n4080;
  assign n4082 = ~n1867 & ~n4081;
  assign n4083 = ~reg_i_StoB_REQ8_out & ~n4082;
  assign n4084 = ~n4037 & ~n4083;
  assign n4085 = ~reg_i_StoB_REQ10_out & ~n4084;
  assign n4086 = ~n2179 & ~n4085;
  assign n4087 = sys_fair10done_out & ~n4086;
  assign n4088 = ~sys_fair10done_out & ~n1944;
  assign n4089 = ~n4087 & ~n4088;
  assign n4090 = sys_fair11done_out & ~n4089;
  assign n4091 = ~n1945 & ~n4090;
  assign n4092 = ~reg_i_StoB_REQ11_out & ~n4091;
  assign n4093 = ~n4034 & ~n4092;
  assign n4094 = sys_fair9done_out & ~n4093;
  assign n4095 = ~n1967 & ~n4094;
  assign n4096 = fair_cnt<1>_out  & ~n4095;
  assign n4097 = ~n1970 & ~n4096;
  assign n4098 = ~fair_cnt<0>_out  & ~n4097;
  assign n4099 = ~n1972 & ~n4098;
  assign n4100 = ~reg_controllable_BtoR_REQ1_out & ~n4099;
  assign n4101 = ~n4031 & ~n4100;
  assign n4102 = ~reg_controllable_BtoR_REQ0_out & ~n4101;
  assign n4103 = ~n4022 & ~n4102;
  assign n4104 = reg_i_RtoB_ACK1_out & ~n4103;
  assign n4105 = ~fair_cnt<1>_out  & ~n4095;
  assign n4106 = ~n2167 & ~n4105;
  assign n4107 = fair_cnt<0>_out  & ~n4106;
  assign n4108 = reg_controllable_BtoS_ACK11_out & ~n3748;
  assign n4109 = reg_controllable_BtoS_ACK10_out & ~n3739;
  assign n4110 = reg_controllable_BtoS_ACK8_out & ~n3734;
  assign n4111 = reg_controllable_BtoS_ACK7_out & ~n3725;
  assign n4112 = reg_controllable_BtoS_ACK6_out & ~n3718;
  assign n4113 = reg_controllable_BtoS_ACK5_out & ~n3711;
  assign n4114 = reg_controllable_BtoS_ACK4_out & ~n3704;
  assign n4115 = reg_controllable_BtoS_ACK3_out & ~n3699;
  assign n4116 = reg_controllable_BtoS_ACK2_out & ~n3692;
  assign n4117 = ~sys_fair0done_out & ~n2213;
  assign n4118 = sys_fair1done_out & ~n4117;
  assign n4119 = ~n4047 & ~n4118;
  assign n4120 = reg_stateG12_out & ~n4119;
  assign n4121 = ~n1614 & ~n4120;
  assign n4122 = ~sys_fair12done_out & ~n4121;
  assign n4123 = ~n4044 & ~n4122;
  assign n4124 = sys_fair2done_out & ~n4123;
  assign n4125 = ~n1643 & ~n4124;
  assign n4126 = ~reg_controllable_BtoS_ACK2_out & ~n4125;
  assign n4127 = ~n4116 & ~n4126;
  assign n4128 = reg_i_StoB_REQ2_out & ~n4127;
  assign n4129 = ~reg_i_StoB_REQ2_out & ~n4125;
  assign n4130 = ~n4128 & ~n4129;
  assign n4131 = sys_fair3done_out & ~n4130;
  assign n4132 = ~n1676 & ~n4131;
  assign n4133 = ~reg_controllable_BtoS_ACK3_out & ~n4132;
  assign n4134 = ~n4115 & ~n4133;
  assign n4135 = reg_i_StoB_REQ3_out & ~n4134;
  assign n4136 = ~reg_i_StoB_REQ3_out & ~n4132;
  assign n4137 = ~n4135 & ~n4136;
  assign n4138 = ~reg_controllable_BtoS_ACK4_out & ~n4137;
  assign n4139 = ~n4114 & ~n4138;
  assign n4140 = reg_i_StoB_REQ4_out & ~n4139;
  assign n4141 = ~reg_i_StoB_REQ4_out & ~n4137;
  assign n4142 = ~n4140 & ~n4141;
  assign n4143 = sys_fair4done_out & ~n4142;
  assign n4144 = ~n4064 & ~n4143;
  assign n4145 = ~reg_controllable_BtoS_ACK5_out & ~n4144;
  assign n4146 = ~n4113 & ~n4145;
  assign n4147 = reg_i_StoB_REQ5_out & ~n4146;
  assign n4148 = ~reg_i_StoB_REQ5_out & ~n4144;
  assign n4149 = ~n4147 & ~n4148;
  assign n4150 = sys_fair5done_out & ~n4149;
  assign n4151 = ~n4069 & ~n4150;
  assign n4152 = ~reg_controllable_BtoS_ACK6_out & ~n4151;
  assign n4153 = ~n4112 & ~n4152;
  assign n4154 = reg_i_StoB_REQ6_out & ~n4153;
  assign n4155 = ~reg_i_StoB_REQ6_out & ~n4151;
  assign n4156 = ~n4154 & ~n4155;
  assign n4157 = sys_fair6done_out & ~n4156;
  assign n4158 = ~n4074 & ~n4157;
  assign n4159 = ~reg_controllable_BtoS_ACK7_out & ~n4158;
  assign n4160 = ~n4111 & ~n4159;
  assign n4161 = reg_i_StoB_REQ7_out & ~n4160;
  assign n4162 = ~reg_i_StoB_REQ7_out & ~n4158;
  assign n4163 = ~n4161 & ~n4162;
  assign n4164 = sys_fair7done_out & ~n4163;
  assign n4165 = ~n4079 & ~n4164;
  assign n4166 = sys_fair8done_out & ~n4165;
  assign n4167 = ~n1867 & ~n4166;
  assign n4168 = ~reg_controllable_BtoS_ACK8_out & ~n4167;
  assign n4169 = ~n4110 & ~n4168;
  assign n4170 = reg_i_StoB_REQ8_out & ~n4169;
  assign n4171 = ~reg_i_StoB_REQ8_out & ~n4167;
  assign n4172 = ~n4170 & ~n4171;
  assign n4173 = ~reg_controllable_BtoS_ACK10_out & ~n4172;
  assign n4174 = ~n4109 & ~n4173;
  assign n4175 = reg_i_StoB_REQ10_out & ~n4174;
  assign n4176 = ~reg_i_StoB_REQ10_out & ~n4172;
  assign n4177 = ~n4175 & ~n4176;
  assign n4178 = sys_fair10done_out & ~n4177;
  assign n4179 = ~n4088 & ~n4178;
  assign n4180 = sys_fair11done_out & ~n4179;
  assign n4181 = ~n1945 & ~n4180;
  assign n4182 = ~reg_controllable_BtoS_ACK11_out & ~n4181;
  assign n4183 = ~n4108 & ~n4182;
  assign n4184 = reg_i_StoB_REQ11_out & ~n4183;
  assign n4185 = ~reg_i_StoB_REQ11_out & ~n4181;
  assign n4186 = ~n4184 & ~n4185;
  assign n4187 = sys_fair9done_out & ~n4186;
  assign n4188 = ~n1967 & ~n4187;
  assign n4189 = fair_cnt<1>_out  & ~n4188;
  assign n4190 = ~n1970 & ~n4189;
  assign n4191 = ~fair_cnt<0>_out  & ~n4190;
  assign n4192 = ~n4107 & ~n4191;
  assign n4193 = env_fair1done_out & ~n4192;
  assign n4194 = ~n2172 & ~n3747;
  assign n4195 = reg_controllable_BtoS_ACK11_out & ~n4194;
  assign n4196 = ~n4182 & ~n4195;
  assign n4197 = reg_i_StoB_REQ11_out & ~n4196;
  assign n4198 = ~n2180 & ~n3733;
  assign n4199 = reg_controllable_BtoS_ACK8_out & ~n4198;
  assign n4200 = ~n4168 & ~n4199;
  assign n4201 = reg_i_StoB_REQ8_out & ~n4200;
  assign n4202 = ~n2197 & ~n3698;
  assign n4203 = reg_controllable_BtoS_ACK3_out & ~n4202;
  assign n4204 = ~n4133 & ~n4203;
  assign n4205 = reg_i_StoB_REQ3_out & ~n4204;
  assign n4206 = ~n2202 & ~n3691;
  assign n4207 = reg_controllable_BtoS_ACK2_out & ~n4206;
  assign n4208 = ~n4126 & ~n4207;
  assign n4209 = reg_i_StoB_REQ2_out & ~n4208;
  assign n4210 = ~sys_fair0done_out & ~n2208;
  assign n4211 = sys_fair1done_out & ~n4210;
  assign n4212 = ~n2215 & ~n4211;
  assign n4213 = reg_stateG12_out & ~n4212;
  assign n4214 = ~n1614 & ~n4213;
  assign n4215 = ~sys_fair12done_out & ~n4214;
  assign n4216 = ~n2217 & ~n4215;
  assign n4217 = sys_fair2done_out & ~n4216;
  assign n4218 = ~n1643 & ~n4217;
  assign n4219 = ~reg_i_StoB_REQ2_out & ~n4218;
  assign n4220 = ~n4209 & ~n4219;
  assign n4221 = sys_fair3done_out & ~n4220;
  assign n4222 = ~n1676 & ~n4221;
  assign n4223 = ~reg_i_StoB_REQ3_out & ~n4222;
  assign n4224 = ~n4205 & ~n4223;
  assign n4225 = ~reg_i_StoB_REQ4_out & ~n4224;
  assign n4226 = ~n4140 & ~n4225;
  assign n4227 = sys_fair4done_out & ~n4226;
  assign n4228 = ~n2242 & ~n4227;
  assign n4229 = ~reg_i_StoB_REQ5_out & ~n4228;
  assign n4230 = ~n4147 & ~n4229;
  assign n4231 = sys_fair5done_out & ~n4230;
  assign n4232 = ~n2251 & ~n4231;
  assign n4233 = ~reg_i_StoB_REQ6_out & ~n4232;
  assign n4234 = ~n4154 & ~n4233;
  assign n4235 = sys_fair6done_out & ~n4234;
  assign n4236 = ~n2260 & ~n4235;
  assign n4237 = ~reg_i_StoB_REQ7_out & ~n4236;
  assign n4238 = ~n4161 & ~n4237;
  assign n4239 = sys_fair7done_out & ~n4238;
  assign n4240 = ~n2269 & ~n4239;
  assign n4241 = sys_fair8done_out & ~n4240;
  assign n4242 = ~n1867 & ~n4241;
  assign n4243 = ~reg_i_StoB_REQ8_out & ~n4242;
  assign n4244 = ~n4201 & ~n4243;
  assign n4245 = ~reg_i_StoB_REQ10_out & ~n4244;
  assign n4246 = ~n4175 & ~n4245;
  assign n4247 = sys_fair10done_out & ~n4246;
  assign n4248 = ~n2282 & ~n4247;
  assign n4249 = sys_fair11done_out & ~n4248;
  assign n4250 = ~n1945 & ~n4249;
  assign n4251 = ~reg_i_StoB_REQ11_out & ~n4250;
  assign n4252 = ~n4197 & ~n4251;
  assign n4253 = sys_fair9done_out & ~n4252;
  assign n4254 = ~n1967 & ~n4253;
  assign n4255 = fair_cnt<1>_out  & ~n4254;
  assign n4256 = ~n4105 & ~n4255;
  assign n4257 = fair_cnt<0>_out  & ~n4256;
  assign n4258 = ~n4098 & ~n4257;
  assign n4259 = ~env_fair1done_out & ~n4258;
  assign n4260 = ~n4193 & ~n4259;
  assign n4261 = env_fair0done_out & ~n4260;
  assign n4262 = fair_cnt<0>_out  & ~n4190;
  assign n4263 = ~n4098 & ~n4262;
  assign n4264 = ~env_fair0done_out & ~n4263;
  assign n4265 = ~n4261 & ~n4264;
  assign n4266 = ~reg_stateG7_0_out & ~n4265;
  assign n4267 = ~reg_stateG7_0_out & ~n4266;
  assign n4268 = reg_nstateG7_1_out & ~n4267;
  assign n4269 = ~reg_nstateG7_1_out & ~n4265;
  assign n4270 = ~n4268 & ~n4269;
  assign n4271 = ~reg_controllable_BtoR_REQ1_out & ~n4270;
  assign n4272 = ~reg_controllable_BtoR_REQ1_out & ~n4271;
  assign n4273 = reg_controllable_BtoR_REQ0_out & ~n4272;
  assign n4274 = reg_controllable_BtoS_ACK11_out & ~n3827;
  assign n4275 = ~n4182 & ~n4274;
  assign n4276 = reg_i_StoB_REQ11_out & ~n4275;
  assign n4277 = reg_controllable_BtoS_ACK10_out & ~n3820;
  assign n4278 = ~n4173 & ~n4277;
  assign n4279 = reg_i_StoB_REQ10_out & ~n4278;
  assign n4280 = reg_controllable_BtoS_ACK8_out & ~n3818;
  assign n4281 = ~n4168 & ~n4280;
  assign n4282 = reg_i_StoB_REQ8_out & ~n4281;
  assign n4283 = reg_controllable_BtoS_ACK7_out & ~n3811;
  assign n4284 = ~n4159 & ~n4283;
  assign n4285 = reg_i_StoB_REQ7_out & ~n4284;
  assign n4286 = reg_controllable_BtoS_ACK6_out & ~n3806;
  assign n4287 = ~n4152 & ~n4286;
  assign n4288 = reg_i_StoB_REQ6_out & ~n4287;
  assign n4289 = reg_controllable_BtoS_ACK5_out & ~n3801;
  assign n4290 = ~n4145 & ~n4289;
  assign n4291 = reg_i_StoB_REQ5_out & ~n4290;
  assign n4292 = reg_controllable_BtoS_ACK4_out & ~n3796;
  assign n4293 = ~n4138 & ~n4292;
  assign n4294 = reg_i_StoB_REQ4_out & ~n4293;
  assign n4295 = reg_controllable_BtoS_ACK3_out & ~n3794;
  assign n4296 = ~n4133 & ~n4295;
  assign n4297 = reg_i_StoB_REQ3_out & ~n4296;
  assign n4298 = reg_controllable_BtoS_ACK2_out & ~n3790;
  assign n4299 = ~n4126 & ~n4298;
  assign n4300 = reg_i_StoB_REQ2_out & ~n4299;
  assign n4301 = sys_fair12done_out & ~n2218;
  assign n4302 = ~sys_fair0done_out & ~n2218;
  assign n4303 = ~sys_fair0done_out & ~n4302;
  assign n4304 = sys_fair1done_out & ~n4303;
  assign n4305 = ~sys_fair1done_out & ~n2218;
  assign n4306 = ~n4304 & ~n4305;
  assign n4307 = reg_stateG12_out & ~n4306;
  assign n4308 = ~n2338 & ~n4307;
  assign n4309 = ~sys_fair12done_out & ~n4308;
  assign n4310 = ~n4301 & ~n4309;
  assign n4311 = sys_fair2done_out & ~n4310;
  assign n4312 = ~n2343 & ~n4311;
  assign n4313 = ~reg_i_StoB_REQ2_out & ~n4312;
  assign n4314 = ~n4300 & ~n4313;
  assign n4315 = sys_fair3done_out & ~n4314;
  assign n4316 = ~n2359 & ~n4315;
  assign n4317 = ~reg_i_StoB_REQ3_out & ~n4316;
  assign n4318 = ~n4297 & ~n4317;
  assign n4319 = ~reg_i_StoB_REQ4_out & ~n4318;
  assign n4320 = ~n4294 & ~n4319;
  assign n4321 = sys_fair4done_out & ~n4320;
  assign n4322 = ~sys_fair4done_out & ~n2415;
  assign n4323 = ~n4321 & ~n4322;
  assign n4324 = ~reg_i_StoB_REQ5_out & ~n4323;
  assign n4325 = ~n4291 & ~n4324;
  assign n4326 = sys_fair5done_out & ~n4325;
  assign n4327 = ~sys_fair5done_out & ~n2438;
  assign n4328 = ~n4326 & ~n4327;
  assign n4329 = ~reg_i_StoB_REQ6_out & ~n4328;
  assign n4330 = ~n4288 & ~n4329;
  assign n4331 = sys_fair6done_out & ~n4330;
  assign n4332 = ~sys_fair6done_out & ~n2461;
  assign n4333 = ~n4331 & ~n4332;
  assign n4334 = ~reg_i_StoB_REQ7_out & ~n4333;
  assign n4335 = ~n4285 & ~n4334;
  assign n4336 = sys_fair7done_out & ~n4335;
  assign n4337 = ~sys_fair7done_out & ~n2479;
  assign n4338 = ~n4336 & ~n4337;
  assign n4339 = sys_fair8done_out & ~n4338;
  assign n4340 = ~n2480 & ~n4339;
  assign n4341 = ~reg_i_StoB_REQ8_out & ~n4340;
  assign n4342 = ~n4282 & ~n4341;
  assign n4343 = ~reg_i_StoB_REQ10_out & ~n4342;
  assign n4344 = ~n4279 & ~n4343;
  assign n4345 = sys_fair10done_out & ~n4344;
  assign n4346 = ~sys_fair10done_out & ~n2527;
  assign n4347 = ~n4345 & ~n4346;
  assign n4348 = sys_fair11done_out & ~n4347;
  assign n4349 = ~n2528 & ~n4348;
  assign n4350 = ~reg_i_StoB_REQ11_out & ~n4349;
  assign n4351 = ~n4276 & ~n4350;
  assign n4352 = sys_fair9done_out & ~n4351;
  assign n4353 = ~n2549 & ~n4352;
  assign n4354 = fair_cnt<1>_out  & ~n4353;
  assign n4355 = ~n2552 & ~n4354;
  assign n4356 = ~fair_cnt<0>_out  & ~n4355;
  assign n4357 = ~n2554 & ~n4356;
  assign n4358 = env_fair1done_out & ~n4357;
  assign n4359 = ~env_fair1done_out & ~n2556;
  assign n4360 = ~n4358 & ~n4359;
  assign n4361 = reg_nstateG7_1_out & ~n4360;
  assign n4362 = ~reg_stateG7_0_out & ~n4360;
  assign n4363 = ~reg_stateG7_0_out & ~n4362;
  assign n4364 = ~reg_nstateG7_1_out & ~n4363;
  assign n4365 = ~n4361 & ~n4364;
  assign n4366 = reg_controllable_BtoR_REQ1_out & ~n4365;
  assign n4367 = env_fair1done_out & ~n4099;
  assign n4368 = ~n1970 & ~n4255;
  assign n4369 = fair_cnt<0>_out  & ~n4368;
  assign n4370 = ~n4098 & ~n4369;
  assign n4371 = ~env_fair1done_out & ~n4370;
  assign n4372 = ~n4367 & ~n4371;
  assign n4373 = reg_nstateG7_1_out & ~n4372;
  assign n4374 = ~reg_nstateG7_1_out & ~n4099;
  assign n4375 = ~n4373 & ~n4374;
  assign n4376 = ~reg_controllable_BtoR_REQ1_out & ~n4375;
  assign n4377 = ~n4366 & ~n4376;
  assign n4378 = ~reg_controllable_BtoR_REQ0_out & ~n4377;
  assign n4379 = ~n4273 & ~n4378;
  assign n4380 = ~reg_i_RtoB_ACK1_out & ~n4379;
  assign n4381 = ~n4104 & ~n4380;
  assign n4382 = reg_i_RtoB_ACK0_out & ~n4381;
  assign n4383 = env_fair0done_out & ~n4357;
  assign n4384 = ~env_fair0done_out & ~n2556;
  assign n4385 = ~n4383 & ~n4384;
  assign n4386 = ~reg_stateG7_0_out & ~n4385;
  assign n4387 = ~reg_stateG7_0_out & ~n4386;
  assign n4388 = reg_nstateG7_1_out & ~n4387;
  assign n4389 = ~reg_nstateG7_1_out & ~n4385;
  assign n4390 = ~n4388 & ~n4389;
  assign n4391 = ~reg_controllable_BtoR_REQ1_out & ~n4390;
  assign n4392 = ~reg_controllable_BtoR_REQ1_out & ~n4391;
  assign n4393 = reg_controllable_BtoR_REQ0_out & ~n4392;
  assign n4394 = ~env_fair1done_out & ~n4263;
  assign n4395 = ~n4193 & ~n4394;
  assign n4396 = env_fair0done_out & ~n4395;
  assign n4397 = env_fair1done_out & ~n4258;
  assign n4398 = ~n4394 & ~n4397;
  assign n4399 = ~env_fair0done_out & ~n4398;
  assign n4400 = ~n4396 & ~n4399;
  assign n4401 = reg_nstateG7_1_out & ~n4400;
  assign n4402 = ~reg_stateG7_0_out & ~n4400;
  assign n4403 = ~reg_stateG7_0_out & ~n4402;
  assign n4404 = ~reg_nstateG7_1_out & ~n4403;
  assign n4405 = ~n4401 & ~n4404;
  assign n4406 = reg_controllable_BtoR_REQ1_out & ~n4405;
  assign n4407 = reg_nstateG7_1_out & ~n4099;
  assign n4408 = env_fair0done_out & ~n4099;
  assign n4409 = ~env_fair0done_out & ~n4370;
  assign n4410 = ~n4408 & ~n4409;
  assign n4411 = ~reg_nstateG7_1_out & ~n4410;
  assign n4412 = ~n4407 & ~n4411;
  assign n4413 = ~reg_controllable_BtoR_REQ1_out & ~n4412;
  assign n4414 = ~n4406 & ~n4413;
  assign n4415 = ~reg_controllable_BtoR_REQ0_out & ~n4414;
  assign n4416 = ~n4393 & ~n4415;
  assign n4417 = reg_i_RtoB_ACK1_out & ~n4416;
  assign n4418 = ~fair_cnt<1>_out  & ~n4188;
  assign n4419 = ~n2167 & ~n4418;
  assign n4420 = fair_cnt<0>_out  & ~n4419;
  assign n4421 = reg_stateG12_out & ~n2637;
  assign n4422 = ~n1614 & ~n4421;
  assign n4423 = ~sys_fair12done_out & ~n4422;
  assign n4424 = ~n2631 & ~n4423;
  assign n4425 = sys_fair2done_out & ~n4424;
  assign n4426 = ~n2638 & ~n4423;
  assign n4427 = ~sys_fair2done_out & ~n4426;
  assign n4428 = ~n4425 & ~n4427;
  assign n4429 = ~reg_controllable_BtoS_ACK2_out & ~n4428;
  assign n4430 = ~n145 & ~n4429;
  assign n4431 = reg_i_StoB_REQ2_out & ~n4430;
  assign n4432 = ~n1643 & ~n4425;
  assign n4433 = reg_controllable_BtoS_ACK2_out & ~n4432;
  assign n4434 = ~n4429 & ~n4433;
  assign n4435 = ~reg_i_StoB_REQ2_out & ~n4434;
  assign n4436 = ~n4431 & ~n4435;
  assign n4437 = sys_fair3done_out & ~n4436;
  assign n4438 = ~reg_controllable_BtoS_ACK2_out & ~n4426;
  assign n4439 = ~n155 & ~n4438;
  assign n4440 = reg_i_StoB_REQ2_out & ~n4439;
  assign n4441 = sys_fair2done_out & ~n4426;
  assign n4442 = ~n1643 & ~n4441;
  assign n4443 = reg_controllable_BtoS_ACK2_out & ~n4442;
  assign n4444 = ~n4438 & ~n4443;
  assign n4445 = ~reg_i_StoB_REQ2_out & ~n4444;
  assign n4446 = ~n4440 & ~n4445;
  assign n4447 = ~sys_fair3done_out & ~n4446;
  assign n4448 = ~n4437 & ~n4447;
  assign n4449 = ~reg_controllable_BtoS_ACK3_out & ~n4448;
  assign n4450 = ~n171 & ~n4449;
  assign n4451 = reg_i_StoB_REQ3_out & ~n4450;
  assign n4452 = ~n1676 & ~n4437;
  assign n4453 = reg_controllable_BtoS_ACK3_out & ~n4452;
  assign n4454 = ~n4449 & ~n4453;
  assign n4455 = ~reg_i_StoB_REQ3_out & ~n4454;
  assign n4456 = ~n4451 & ~n4455;
  assign n4457 = ~reg_controllable_BtoS_ACK4_out & ~n4456;
  assign n4458 = ~n1584 & ~n4457;
  assign n4459 = reg_i_StoB_REQ4_out & ~n4458;
  assign n4460 = ~reg_i_StoB_REQ4_out & ~n4456;
  assign n4461 = ~n4459 & ~n4460;
  assign n4462 = sys_fair4done_out & ~n4461;
  assign n4463 = ~reg_controllable_BtoS_ACK3_out & ~n4446;
  assign n4464 = ~n186 & ~n4463;
  assign n4465 = reg_i_StoB_REQ3_out & ~n4464;
  assign n4466 = sys_fair3done_out & ~n4446;
  assign n4467 = ~n1676 & ~n4466;
  assign n4468 = reg_controllable_BtoS_ACK3_out & ~n4467;
  assign n4469 = ~n4463 & ~n4468;
  assign n4470 = ~reg_i_StoB_REQ3_out & ~n4469;
  assign n4471 = ~n4465 & ~n4470;
  assign n4472 = ~reg_controllable_BtoS_ACK4_out & ~n4471;
  assign n4473 = ~n198 & ~n4472;
  assign n4474 = reg_i_StoB_REQ4_out & ~n4473;
  assign n4475 = ~n1722 & ~n4472;
  assign n4476 = ~reg_i_StoB_REQ4_out & ~n4475;
  assign n4477 = ~n4474 & ~n4476;
  assign n4478 = ~sys_fair4done_out & ~n4477;
  assign n4479 = ~n4462 & ~n4478;
  assign n4480 = ~reg_controllable_BtoS_ACK5_out & ~n4479;
  assign n4481 = ~n1583 & ~n4480;
  assign n4482 = reg_i_StoB_REQ5_out & ~n4481;
  assign n4483 = ~reg_i_StoB_REQ5_out & ~n4479;
  assign n4484 = ~n4482 & ~n4483;
  assign n4485 = sys_fair5done_out & ~n4484;
  assign n4486 = ~n1702 & ~n4472;
  assign n4487 = reg_i_StoB_REQ4_out & ~n4486;
  assign n4488 = ~reg_i_StoB_REQ4_out & ~n4471;
  assign n4489 = ~n4487 & ~n4488;
  assign n4490 = sys_fair4done_out & ~n4489;
  assign n4491 = ~n4478 & ~n4490;
  assign n4492 = ~reg_controllable_BtoS_ACK5_out & ~n4491;
  assign n4493 = ~n222 & ~n4492;
  assign n4494 = reg_i_StoB_REQ5_out & ~n4493;
  assign n4495 = ~n1763 & ~n4492;
  assign n4496 = ~reg_i_StoB_REQ5_out & ~n4495;
  assign n4497 = ~n4494 & ~n4496;
  assign n4498 = ~sys_fair5done_out & ~n4497;
  assign n4499 = ~n4485 & ~n4498;
  assign n4500 = ~reg_controllable_BtoS_ACK6_out & ~n4499;
  assign n4501 = ~n1582 & ~n4500;
  assign n4502 = reg_i_StoB_REQ6_out & ~n4501;
  assign n4503 = ~reg_i_StoB_REQ6_out & ~n4499;
  assign n4504 = ~n4502 & ~n4503;
  assign n4505 = sys_fair6done_out & ~n4504;
  assign n4506 = ~n1746 & ~n4492;
  assign n4507 = reg_i_StoB_REQ5_out & ~n4506;
  assign n4508 = ~reg_i_StoB_REQ5_out & ~n4491;
  assign n4509 = ~n4507 & ~n4508;
  assign n4510 = sys_fair5done_out & ~n4509;
  assign n4511 = ~n4498 & ~n4510;
  assign n4512 = ~reg_controllable_BtoS_ACK6_out & ~n4511;
  assign n4513 = ~n246 & ~n4512;
  assign n4514 = reg_i_StoB_REQ6_out & ~n4513;
  assign n4515 = ~n1799 & ~n4512;
  assign n4516 = ~reg_i_StoB_REQ6_out & ~n4515;
  assign n4517 = ~n4514 & ~n4516;
  assign n4518 = ~sys_fair6done_out & ~n4517;
  assign n4519 = ~n4505 & ~n4518;
  assign n4520 = ~reg_controllable_BtoS_ACK7_out & ~n4519;
  assign n4521 = ~n1581 & ~n4520;
  assign n4522 = reg_i_StoB_REQ7_out & ~n4521;
  assign n4523 = ~reg_i_StoB_REQ7_out & ~n4519;
  assign n4524 = ~n4522 & ~n4523;
  assign n4525 = sys_fair7done_out & ~n4524;
  assign n4526 = ~n1782 & ~n4512;
  assign n4527 = reg_i_StoB_REQ6_out & ~n4526;
  assign n4528 = ~reg_i_StoB_REQ6_out & ~n4511;
  assign n4529 = ~n4527 & ~n4528;
  assign n4530 = sys_fair6done_out & ~n4529;
  assign n4531 = ~n4518 & ~n4530;
  assign n4532 = ~reg_controllable_BtoS_ACK7_out & ~n4531;
  assign n4533 = ~n270 & ~n4532;
  assign n4534 = reg_i_StoB_REQ7_out & ~n4533;
  assign n4535 = ~n1835 & ~n4532;
  assign n4536 = ~reg_i_StoB_REQ7_out & ~n4535;
  assign n4537 = ~n4534 & ~n4536;
  assign n4538 = ~sys_fair7done_out & ~n4537;
  assign n4539 = ~n4525 & ~n4538;
  assign n4540 = sys_fair8done_out & ~n4539;
  assign n4541 = ~n1818 & ~n4532;
  assign n4542 = reg_i_StoB_REQ7_out & ~n4541;
  assign n4543 = ~reg_i_StoB_REQ7_out & ~n4531;
  assign n4544 = ~n4542 & ~n4543;
  assign n4545 = sys_fair7done_out & ~n4544;
  assign n4546 = ~n4538 & ~n4545;
  assign n4547 = ~sys_fair8done_out & ~n4546;
  assign n4548 = ~n4540 & ~n4547;
  assign n4549 = ~reg_controllable_BtoS_ACK8_out & ~n4548;
  assign n4550 = ~n293 & ~n4549;
  assign n4551 = reg_i_StoB_REQ8_out & ~n4550;
  assign n4552 = ~n1867 & ~n4540;
  assign n4553 = reg_controllable_BtoS_ACK8_out & ~n4552;
  assign n4554 = ~n4549 & ~n4553;
  assign n4555 = ~reg_i_StoB_REQ8_out & ~n4554;
  assign n4556 = ~n4551 & ~n4555;
  assign n4557 = ~reg_controllable_BtoS_ACK10_out & ~n4556;
  assign n4558 = ~n1579 & ~n4557;
  assign n4559 = reg_i_StoB_REQ10_out & ~n4558;
  assign n4560 = ~reg_i_StoB_REQ10_out & ~n4556;
  assign n4561 = ~n4559 & ~n4560;
  assign n4562 = sys_fair10done_out & ~n4561;
  assign n4563 = ~reg_controllable_BtoS_ACK8_out & ~n4546;
  assign n4564 = ~n308 & ~n4563;
  assign n4565 = reg_i_StoB_REQ8_out & ~n4564;
  assign n4566 = sys_fair8done_out & ~n4546;
  assign n4567 = ~n1867 & ~n4566;
  assign n4568 = reg_controllable_BtoS_ACK8_out & ~n4567;
  assign n4569 = ~n4563 & ~n4568;
  assign n4570 = ~reg_i_StoB_REQ8_out & ~n4569;
  assign n4571 = ~n4565 & ~n4570;
  assign n4572 = ~reg_controllable_BtoS_ACK10_out & ~n4571;
  assign n4573 = ~n320 & ~n4572;
  assign n4574 = reg_i_StoB_REQ10_out & ~n4573;
  assign n4575 = ~n1908 & ~n4572;
  assign n4576 = ~reg_i_StoB_REQ10_out & ~n4575;
  assign n4577 = ~n4574 & ~n4576;
  assign n4578 = ~sys_fair10done_out & ~n4577;
  assign n4579 = ~n4562 & ~n4578;
  assign n4580 = sys_fair11done_out & ~n4579;
  assign n4581 = ~n1888 & ~n4572;
  assign n4582 = reg_i_StoB_REQ10_out & ~n4581;
  assign n4583 = ~reg_i_StoB_REQ10_out & ~n4571;
  assign n4584 = ~n4582 & ~n4583;
  assign n4585 = sys_fair10done_out & ~n4584;
  assign n4586 = ~n4578 & ~n4585;
  assign n4587 = ~sys_fair11done_out & ~n4586;
  assign n4588 = ~n4580 & ~n4587;
  assign n4589 = ~reg_controllable_BtoS_ACK11_out & ~n4588;
  assign n4590 = ~n343 & ~n4589;
  assign n4591 = reg_i_StoB_REQ11_out & ~n4590;
  assign n4592 = ~n1945 & ~n4580;
  assign n4593 = reg_controllable_BtoS_ACK11_out & ~n4592;
  assign n4594 = ~n4589 & ~n4593;
  assign n4595 = ~reg_i_StoB_REQ11_out & ~n4594;
  assign n4596 = ~n4591 & ~n4595;
  assign n4597 = sys_fair9done_out & ~n4596;
  assign n4598 = ~n1967 & ~n4597;
  assign n4599 = fair_cnt<1>_out  & ~n4598;
  assign n4600 = ~n4105 & ~n4599;
  assign n4601 = ~fair_cnt<0>_out  & ~n4600;
  assign n4602 = ~n4420 & ~n4601;
  assign n4603 = env_fair0done_out & ~n4602;
  assign n4604 = ~env_fair0done_out & ~n4192;
  assign n4605 = ~n4603 & ~n4604;
  assign n4606 = ~reg_stateG7_0_out & ~n4605;
  assign n4607 = ~reg_stateG7_0_out & ~n4606;
  assign n4608 = reg_nstateG7_1_out & ~n4607;
  assign n4609 = ~reg_nstateG7_1_out & ~n4605;
  assign n4610 = ~n4608 & ~n4609;
  assign n4611 = ~reg_controllable_BtoR_REQ1_out & ~n4610;
  assign n4612 = ~reg_controllable_BtoR_REQ1_out & ~n4611;
  assign n4613 = reg_controllable_BtoR_REQ0_out & ~n4612;
  assign n4614 = env_fair1done_out & ~n4602;
  assign n4615 = ~env_fair1done_out & ~n4192;
  assign n4616 = ~n4614 & ~n4615;
  assign n4617 = reg_nstateG7_1_out & ~n4616;
  assign n4618 = ~reg_stateG7_0_out & ~n4616;
  assign n4619 = ~reg_stateG7_0_out & ~n4618;
  assign n4620 = ~reg_nstateG7_1_out & ~n4619;
  assign n4621 = ~n4617 & ~n4620;
  assign n4622 = reg_controllable_BtoR_REQ1_out & ~n4621;
  assign n4623 = fair_cnt<0>_out  & ~n4600;
  assign n4624 = ~n4191 & ~n4623;
  assign n4625 = ~env_fair1done_out & ~n4624;
  assign n4626 = ~n4614 & ~n4625;
  assign n4627 = reg_nstateG7_1_out & ~n4626;
  assign n4628 = ~env_fair0done_out & ~n4624;
  assign n4629 = ~n4603 & ~n4628;
  assign n4630 = ~reg_nstateG7_1_out & ~n4629;
  assign n4631 = ~n4627 & ~n4630;
  assign n4632 = ~reg_controllable_BtoR_REQ1_out & ~n4631;
  assign n4633 = ~n4622 & ~n4632;
  assign n4634 = ~reg_controllable_BtoR_REQ0_out & ~n4633;
  assign n4635 = ~n4613 & ~n4634;
  assign n4636 = ~reg_i_RtoB_ACK1_out & ~n4635;
  assign n4637 = ~n4417 & ~n4636;
  assign n4638 = ~reg_i_RtoB_ACK0_out & ~n4637;
  assign n4639 = ~n4382 & ~n4638;
  assign n4640 = ~reg_i_StoB_REQ9_out & ~n4639;
  assign n4641 = ~n3941 & ~n4640;
  assign n4642 = reg_controllable_BtoS_ACK9_out & ~n4641;
  assign n4643 = ~n2876 & ~n3674;
  assign n4644 = env_fair0done_out & ~n4643;
  assign n4645 = ~env_fair0done_out & ~n2877;
  assign n4646 = ~n4644 & ~n4645;
  assign n4647 = ~reg_stateG7_0_out & ~n4646;
  assign n4648 = ~reg_stateG7_0_out & ~n4647;
  assign n4649 = reg_nstateG7_1_out & ~n4648;
  assign n4650 = ~reg_nstateG7_1_out & ~n4646;
  assign n4651 = ~n4649 & ~n4650;
  assign n4652 = ~reg_controllable_BtoR_REQ1_out & ~n4651;
  assign n4653 = ~reg_controllable_BtoR_REQ1_out & ~n4652;
  assign n4654 = reg_controllable_BtoR_REQ0_out & ~n4653;
  assign n4655 = env_fair1done_out & ~n4643;
  assign n4656 = ~env_fair1done_out & ~n2877;
  assign n4657 = ~n4655 & ~n4656;
  assign n4658 = reg_nstateG7_1_out & ~n4657;
  assign n4659 = ~reg_stateG7_0_out & ~n4657;
  assign n4660 = ~reg_stateG7_0_out & ~n4659;
  assign n4661 = ~reg_nstateG7_1_out & ~n4660;
  assign n4662 = ~n4658 & ~n4661;
  assign n4663 = reg_controllable_BtoR_REQ1_out & ~n4662;
  assign n4664 = ~n2931 & ~n4663;
  assign n4665 = ~reg_controllable_BtoR_REQ0_out & ~n4664;
  assign n4666 = ~n4654 & ~n4665;
  assign n4667 = reg_i_RtoB_ACK1_out & ~n4666;
  assign n4668 = ~n2949 & ~n4191;
  assign n4669 = env_fair1done_out & ~n4668;
  assign n4670 = ~n1973 & ~n4262;
  assign n4671 = ~env_fair1done_out & ~n4670;
  assign n4672 = ~n4669 & ~n4671;
  assign n4673 = env_fair0done_out & ~n4672;
  assign n4674 = ~env_fair0done_out & ~n4670;
  assign n4675 = ~n4673 & ~n4674;
  assign n4676 = ~reg_stateG7_0_out & ~n4675;
  assign n4677 = ~reg_stateG7_0_out & ~n4676;
  assign n4678 = reg_nstateG7_1_out & ~n4677;
  assign n4679 = ~reg_nstateG7_1_out & ~n4675;
  assign n4680 = ~n4678 & ~n4679;
  assign n4681 = ~reg_controllable_BtoR_REQ1_out & ~n4680;
  assign n4682 = ~reg_controllable_BtoR_REQ1_out & ~n4681;
  assign n4683 = reg_controllable_BtoR_REQ0_out & ~n4682;
  assign n4684 = ~n2929 & ~n4191;
  assign n4685 = env_fair1done_out & ~n4684;
  assign n4686 = ~env_fair1done_out & ~n2930;
  assign n4687 = ~n4685 & ~n4686;
  assign n4688 = reg_nstateG7_1_out & ~n4687;
  assign n4689 = ~reg_stateG7_0_out & ~n4687;
  assign n4690 = ~reg_stateG7_0_out & ~n4689;
  assign n4691 = ~reg_nstateG7_1_out & ~n4690;
  assign n4692 = ~n4688 & ~n4691;
  assign n4693 = reg_controllable_BtoR_REQ1_out & ~n4692;
  assign n4694 = ~n2969 & ~n4671;
  assign n4695 = reg_nstateG7_1_out & ~n4694;
  assign n4696 = ~n2972 & ~n4695;
  assign n4697 = ~reg_controllable_BtoR_REQ1_out & ~n4696;
  assign n4698 = ~n4693 & ~n4697;
  assign n4699 = ~reg_controllable_BtoR_REQ0_out & ~n4698;
  assign n4700 = ~n4683 & ~n4699;
  assign n4701 = ~reg_i_RtoB_ACK1_out & ~n4700;
  assign n4702 = ~n4667 & ~n4701;
  assign n4703 = reg_i_RtoB_ACK0_out & ~n4702;
  assign n4704 = env_fair0done_out & ~n4684;
  assign n4705 = ~env_fair0done_out & ~n2930;
  assign n4706 = ~n4704 & ~n4705;
  assign n4707 = ~reg_stateG7_0_out & ~n4706;
  assign n4708 = ~reg_stateG7_0_out & ~n4707;
  assign n4709 = reg_nstateG7_1_out & ~n4708;
  assign n4710 = ~reg_nstateG7_1_out & ~n4706;
  assign n4711 = ~n4709 & ~n4710;
  assign n4712 = ~reg_controllable_BtoR_REQ1_out & ~n4711;
  assign n4713 = ~reg_controllable_BtoR_REQ1_out & ~n4712;
  assign n4714 = reg_controllable_BtoR_REQ0_out & ~n4713;
  assign n4715 = reg_nstateG7_1_out & ~n4675;
  assign n4716 = ~reg_nstateG7_1_out & ~n4677;
  assign n4717 = ~n4715 & ~n4716;
  assign n4718 = reg_controllable_BtoR_REQ1_out & ~n4717;
  assign n4719 = ~n2990 & ~n4674;
  assign n4720 = ~reg_nstateG7_1_out & ~n4719;
  assign n4721 = ~n2963 & ~n4720;
  assign n4722 = ~reg_controllable_BtoR_REQ1_out & ~n4721;
  assign n4723 = ~n4718 & ~n4722;
  assign n4724 = ~reg_controllable_BtoR_REQ0_out & ~n4723;
  assign n4725 = ~n4714 & ~n4724;
  assign n4726 = reg_i_RtoB_ACK1_out & ~n4725;
  assign n4727 = ~n2947 & ~n4418;
  assign n4728 = fair_cnt<0>_out  & ~n4727;
  assign n4729 = ~reg_controllable_BtoS_ACK11_out & ~n4586;
  assign n4730 = ~n353 & ~n4729;
  assign n4731 = reg_i_StoB_REQ11_out & ~n4730;
  assign n4732 = sys_fair11done_out & ~n4586;
  assign n4733 = ~n1945 & ~n4732;
  assign n4734 = reg_controllable_BtoS_ACK11_out & ~n4733;
  assign n4735 = ~n4729 & ~n4734;
  assign n4736 = ~reg_i_StoB_REQ11_out & ~n4735;
  assign n4737 = ~n4731 & ~n4736;
  assign n4738 = ~sys_fair9done_out & ~n4737;
  assign n4739 = ~n4597 & ~n4738;
  assign n4740 = fair_cnt<1>_out  & ~n4739;
  assign n4741 = ~n1970 & ~n4740;
  assign n4742 = ~fair_cnt<0>_out  & ~n4741;
  assign n4743 = ~n4728 & ~n4742;
  assign n4744 = env_fair0done_out & ~n4743;
  assign n4745 = ~env_fair0done_out & ~n4668;
  assign n4746 = ~n4744 & ~n4745;
  assign n4747 = ~reg_stateG7_0_out & ~n4746;
  assign n4748 = ~reg_stateG7_0_out & ~n4747;
  assign n4749 = reg_nstateG7_1_out & ~n4748;
  assign n4750 = ~reg_nstateG7_1_out & ~n4746;
  assign n4751 = ~n4749 & ~n4750;
  assign n4752 = ~reg_controllable_BtoR_REQ1_out & ~n4751;
  assign n4753 = ~reg_controllable_BtoR_REQ1_out & ~n4752;
  assign n4754 = reg_controllable_BtoR_REQ0_out & ~n4753;
  assign n4755 = env_fair1done_out & ~n4743;
  assign n4756 = ~env_fair1done_out & ~n4668;
  assign n4757 = ~n4755 & ~n4756;
  assign n4758 = reg_nstateG7_1_out & ~n4757;
  assign n4759 = ~reg_stateG7_0_out & ~n4757;
  assign n4760 = ~reg_stateG7_0_out & ~n4759;
  assign n4761 = ~reg_nstateG7_1_out & ~n4760;
  assign n4762 = ~n4758 & ~n4761;
  assign n4763 = reg_controllable_BtoR_REQ1_out & ~n4762;
  assign n4764 = fair_cnt<0>_out  & ~n4741;
  assign n4765 = ~n4191 & ~n4764;
  assign n4766 = ~env_fair1done_out & ~n4765;
  assign n4767 = ~n4755 & ~n4766;
  assign n4768 = reg_nstateG7_1_out & ~n4767;
  assign n4769 = ~env_fair0done_out & ~n4765;
  assign n4770 = ~n4744 & ~n4769;
  assign n4771 = ~reg_nstateG7_1_out & ~n4770;
  assign n4772 = ~n4768 & ~n4771;
  assign n4773 = ~reg_controllable_BtoR_REQ1_out & ~n4772;
  assign n4774 = ~n4763 & ~n4773;
  assign n4775 = ~reg_controllable_BtoR_REQ0_out & ~n4774;
  assign n4776 = ~n4754 & ~n4775;
  assign n4777 = ~reg_i_RtoB_ACK1_out & ~n4776;
  assign n4778 = ~n4726 & ~n4777;
  assign n4779 = ~reg_i_RtoB_ACK0_out & ~n4778;
  assign n4780 = ~n4703 & ~n4779;
  assign n4781 = reg_i_StoB_REQ9_out & ~n4780;
  assign n4782 = ~n3071 & ~n4010;
  assign n4783 = env_fair0done_out & ~n4782;
  assign n4784 = ~env_fair0done_out & ~n3072;
  assign n4785 = ~n4783 & ~n4784;
  assign n4786 = ~reg_stateG7_0_out & ~n4785;
  assign n4787 = ~reg_stateG7_0_out & ~n4786;
  assign n4788 = reg_nstateG7_1_out & ~n4787;
  assign n4789 = ~reg_nstateG7_1_out & ~n4785;
  assign n4790 = ~n4788 & ~n4789;
  assign n4791 = ~reg_controllable_BtoR_REQ1_out & ~n4790;
  assign n4792 = ~reg_controllable_BtoR_REQ1_out & ~n4791;
  assign n4793 = reg_controllable_BtoR_REQ0_out & ~n4792;
  assign n4794 = env_fair1done_out & ~n4782;
  assign n4795 = ~env_fair1done_out & ~n3072;
  assign n4796 = ~n4794 & ~n4795;
  assign n4797 = reg_nstateG7_1_out & ~n4796;
  assign n4798 = ~reg_stateG7_0_out & ~n4796;
  assign n4799 = ~reg_stateG7_0_out & ~n4798;
  assign n4800 = ~reg_nstateG7_1_out & ~n4799;
  assign n4801 = ~n4797 & ~n4800;
  assign n4802 = reg_controllable_BtoR_REQ1_out & ~n4801;
  assign n4803 = ~n3126 & ~n4098;
  assign n4804 = ~reg_controllable_BtoR_REQ1_out & ~n4803;
  assign n4805 = ~n4802 & ~n4804;
  assign n4806 = ~reg_controllable_BtoR_REQ0_out & ~n4805;
  assign n4807 = ~n4793 & ~n4806;
  assign n4808 = reg_i_RtoB_ACK1_out & ~n4807;
  assign n4809 = ~n2947 & ~n4105;
  assign n4810 = fair_cnt<0>_out  & ~n4809;
  assign n4811 = ~n4191 & ~n4810;
  assign n4812 = env_fair1done_out & ~n4811;
  assign n4813 = ~n4259 & ~n4812;
  assign n4814 = env_fair0done_out & ~n4813;
  assign n4815 = ~n4264 & ~n4814;
  assign n4816 = ~reg_stateG7_0_out & ~n4815;
  assign n4817 = ~reg_stateG7_0_out & ~n4816;
  assign n4818 = reg_nstateG7_1_out & ~n4817;
  assign n4819 = ~reg_nstateG7_1_out & ~n4815;
  assign n4820 = ~n4818 & ~n4819;
  assign n4821 = ~reg_controllable_BtoR_REQ1_out & ~n4820;
  assign n4822 = ~reg_controllable_BtoR_REQ1_out & ~n4821;
  assign n4823 = reg_controllable_BtoR_REQ0_out & ~n4822;
  assign n4824 = ~n3158 & ~n4356;
  assign n4825 = env_fair1done_out & ~n4824;
  assign n4826 = ~env_fair1done_out & ~n3159;
  assign n4827 = ~n4825 & ~n4826;
  assign n4828 = reg_nstateG7_1_out & ~n4827;
  assign n4829 = ~reg_stateG7_0_out & ~n4827;
  assign n4830 = ~reg_stateG7_0_out & ~n4829;
  assign n4831 = ~reg_nstateG7_1_out & ~n4830;
  assign n4832 = ~n4828 & ~n4831;
  assign n4833 = reg_controllable_BtoR_REQ1_out & ~n4832;
  assign n4834 = env_fair1done_out & ~n4803;
  assign n4835 = ~n4371 & ~n4834;
  assign n4836 = reg_nstateG7_1_out & ~n4835;
  assign n4837 = ~reg_nstateG7_1_out & ~n4803;
  assign n4838 = ~n4836 & ~n4837;
  assign n4839 = ~reg_controllable_BtoR_REQ1_out & ~n4838;
  assign n4840 = ~n4833 & ~n4839;
  assign n4841 = ~reg_controllable_BtoR_REQ0_out & ~n4840;
  assign n4842 = ~n4823 & ~n4841;
  assign n4843 = ~reg_i_RtoB_ACK1_out & ~n4842;
  assign n4844 = ~n4808 & ~n4843;
  assign n4845 = reg_i_RtoB_ACK0_out & ~n4844;
  assign n4846 = env_fair0done_out & ~n4824;
  assign n4847 = ~env_fair0done_out & ~n3159;
  assign n4848 = ~n4846 & ~n4847;
  assign n4849 = ~reg_stateG7_0_out & ~n4848;
  assign n4850 = ~reg_stateG7_0_out & ~n4849;
  assign n4851 = reg_nstateG7_1_out & ~n4850;
  assign n4852 = ~reg_nstateG7_1_out & ~n4848;
  assign n4853 = ~n4851 & ~n4852;
  assign n4854 = ~reg_controllable_BtoR_REQ1_out & ~n4853;
  assign n4855 = ~reg_controllable_BtoR_REQ1_out & ~n4854;
  assign n4856 = reg_controllable_BtoR_REQ0_out & ~n4855;
  assign n4857 = ~n4394 & ~n4812;
  assign n4858 = env_fair0done_out & ~n4857;
  assign n4859 = ~n4399 & ~n4858;
  assign n4860 = reg_nstateG7_1_out & ~n4859;
  assign n4861 = ~reg_stateG7_0_out & ~n4859;
  assign n4862 = ~reg_stateG7_0_out & ~n4861;
  assign n4863 = ~reg_nstateG7_1_out & ~n4862;
  assign n4864 = ~n4860 & ~n4863;
  assign n4865 = reg_controllable_BtoR_REQ1_out & ~n4864;
  assign n4866 = reg_nstateG7_1_out & ~n4803;
  assign n4867 = env_fair0done_out & ~n4803;
  assign n4868 = ~n4409 & ~n4867;
  assign n4869 = ~reg_nstateG7_1_out & ~n4868;
  assign n4870 = ~n4866 & ~n4869;
  assign n4871 = ~reg_controllable_BtoR_REQ1_out & ~n4870;
  assign n4872 = ~n4865 & ~n4871;
  assign n4873 = ~reg_controllable_BtoR_REQ0_out & ~n4872;
  assign n4874 = ~n4856 & ~n4873;
  assign n4875 = reg_i_RtoB_ACK1_out & ~n4874;
  assign n4876 = ~n4105 & ~n4740;
  assign n4877 = ~fair_cnt<0>_out  & ~n4876;
  assign n4878 = ~n4728 & ~n4877;
  assign n4879 = env_fair0done_out & ~n4878;
  assign n4880 = ~env_fair0done_out & ~n4811;
  assign n4881 = ~n4879 & ~n4880;
  assign n4882 = ~reg_stateG7_0_out & ~n4881;
  assign n4883 = ~reg_stateG7_0_out & ~n4882;
  assign n4884 = reg_nstateG7_1_out & ~n4883;
  assign n4885 = ~reg_nstateG7_1_out & ~n4881;
  assign n4886 = ~n4884 & ~n4885;
  assign n4887 = ~reg_controllable_BtoR_REQ1_out & ~n4886;
  assign n4888 = ~reg_controllable_BtoR_REQ1_out & ~n4887;
  assign n4889 = reg_controllable_BtoR_REQ0_out & ~n4888;
  assign n4890 = env_fair1done_out & ~n4878;
  assign n4891 = ~env_fair1done_out & ~n4811;
  assign n4892 = ~n4890 & ~n4891;
  assign n4893 = reg_nstateG7_1_out & ~n4892;
  assign n4894 = ~reg_stateG7_0_out & ~n4892;
  assign n4895 = ~reg_stateG7_0_out & ~n4894;
  assign n4896 = ~reg_nstateG7_1_out & ~n4895;
  assign n4897 = ~n4893 & ~n4896;
  assign n4898 = reg_controllable_BtoR_REQ1_out & ~n4897;
  assign n4899 = fair_cnt<0>_out  & ~n4876;
  assign n4900 = ~n4191 & ~n4899;
  assign n4901 = ~env_fair1done_out & ~n4900;
  assign n4902 = ~n4890 & ~n4901;
  assign n4903 = reg_nstateG7_1_out & ~n4902;
  assign n4904 = ~env_fair0done_out & ~n4900;
  assign n4905 = ~n4879 & ~n4904;
  assign n4906 = ~reg_nstateG7_1_out & ~n4905;
  assign n4907 = ~n4903 & ~n4906;
  assign n4908 = ~reg_controllable_BtoR_REQ1_out & ~n4907;
  assign n4909 = ~n4898 & ~n4908;
  assign n4910 = ~reg_controllable_BtoR_REQ0_out & ~n4909;
  assign n4911 = ~n4889 & ~n4910;
  assign n4912 = ~reg_i_RtoB_ACK1_out & ~n4911;
  assign n4913 = ~n4875 & ~n4912;
  assign n4914 = ~reg_i_RtoB_ACK0_out & ~n4913;
  assign n4915 = ~n4845 & ~n4914;
  assign n4916 = ~reg_i_StoB_REQ9_out & ~n4915;
  assign n4917 = ~n4781 & ~n4916;
  assign n4918 = ~reg_controllable_BtoS_ACK9_out & ~n4917;
  assign n4919 = ~n4642 & ~n4918;
  assign n4920 = ~reg_controllable_DEQ_out & ~n4919;
  assign n4921 = ~n3670 & ~n4920;
  assign n4922 = reg_controllable_ENQ_out & ~n4921;
  assign n4923 = reg_controllable_DEQ_out & ~n3665;
  assign n4924 = reg_i_nEMPTY_out & ~n4919;
  assign n4925 = reg_i_nEMPTY_out & ~n4924;
  assign n4926 = reg_i_FULL_out & ~n4925;
  assign n4927 = ~n3681 & ~n3756;
  assign n4928 = ~fair_cnt<0>_out  & ~n4927;
  assign n4929 = ~n3898 & ~n4928;
  assign n4930 = env_fair0done_out & ~n4929;
  assign n4931 = ~n3905 & ~n4930;
  assign n4932 = ~reg_stateG7_0_out & ~n4931;
  assign n4933 = ~reg_stateG7_0_out & ~n4932;
  assign n4934 = reg_nstateG7_1_out & ~n4933;
  assign n4935 = ~reg_nstateG7_1_out & ~n4931;
  assign n4936 = ~n4934 & ~n4935;
  assign n4937 = ~reg_controllable_BtoR_REQ1_out & ~n4936;
  assign n4938 = ~reg_controllable_BtoR_REQ1_out & ~n4937;
  assign n4939 = reg_controllable_BtoR_REQ0_out & ~n4938;
  assign n4940 = env_fair1done_out & ~n4929;
  assign n4941 = ~n3916 & ~n4940;
  assign n4942 = reg_nstateG7_1_out & ~n4941;
  assign n4943 = ~reg_stateG7_0_out & ~n4941;
  assign n4944 = ~reg_stateG7_0_out & ~n4943;
  assign n4945 = ~reg_nstateG7_1_out & ~n4944;
  assign n4946 = ~n4942 & ~n4945;
  assign n4947 = reg_controllable_BtoR_REQ1_out & ~n4946;
  assign n4948 = fair_cnt<0>_out  & ~n4927;
  assign n4949 = ~n3758 & ~n4948;
  assign n4950 = ~env_fair1done_out & ~n4949;
  assign n4951 = ~n4940 & ~n4950;
  assign n4952 = reg_nstateG7_1_out & ~n4951;
  assign n4953 = ~env_fair0done_out & ~n4949;
  assign n4954 = ~n4930 & ~n4953;
  assign n4955 = ~reg_nstateG7_1_out & ~n4954;
  assign n4956 = ~n4952 & ~n4955;
  assign n4957 = ~reg_controllable_BtoR_REQ1_out & ~n4956;
  assign n4958 = ~n4947 & ~n4957;
  assign n4959 = ~reg_controllable_BtoR_REQ0_out & ~n4958;
  assign n4960 = ~n4939 & ~n4959;
  assign n4961 = ~reg_i_RtoB_ACK1_out & ~n4960;
  assign n4962 = ~n3895 & ~n4961;
  assign n4963 = ~reg_i_RtoB_ACK0_out & ~n4962;
  assign n4964 = ~n3860 & ~n4963;
  assign n4965 = reg_i_StoB_REQ9_out & ~n4964;
  assign n4966 = ~n1969 & ~n4105;
  assign n4967 = fair_cnt<0>_out  & ~n4966;
  assign n4968 = ~n4191 & ~n4967;
  assign n4969 = env_fair1done_out & ~n4968;
  assign n4970 = ~n4259 & ~n4969;
  assign n4971 = env_fair0done_out & ~n4970;
  assign n4972 = ~n4264 & ~n4971;
  assign n4973 = ~reg_stateG7_0_out & ~n4972;
  assign n4974 = ~reg_stateG7_0_out & ~n4973;
  assign n4975 = reg_nstateG7_1_out & ~n4974;
  assign n4976 = ~reg_nstateG7_1_out & ~n4972;
  assign n4977 = ~n4975 & ~n4976;
  assign n4978 = ~reg_controllable_BtoR_REQ1_out & ~n4977;
  assign n4979 = ~reg_controllable_BtoR_REQ1_out & ~n4978;
  assign n4980 = reg_controllable_BtoR_REQ0_out & ~n4979;
  assign n4981 = ~n4378 & ~n4980;
  assign n4982 = ~reg_i_RtoB_ACK1_out & ~n4981;
  assign n4983 = ~n4104 & ~n4982;
  assign n4984 = reg_i_RtoB_ACK0_out & ~n4983;
  assign n4985 = ~n4394 & ~n4969;
  assign n4986 = env_fair0done_out & ~n4985;
  assign n4987 = ~n4399 & ~n4986;
  assign n4988 = reg_nstateG7_1_out & ~n4987;
  assign n4989 = ~reg_stateG7_0_out & ~n4987;
  assign n4990 = ~reg_stateG7_0_out & ~n4989;
  assign n4991 = ~reg_nstateG7_1_out & ~n4990;
  assign n4992 = ~n4988 & ~n4991;
  assign n4993 = reg_controllable_BtoR_REQ1_out & ~n4992;
  assign n4994 = ~n4413 & ~n4993;
  assign n4995 = ~reg_controllable_BtoR_REQ0_out & ~n4994;
  assign n4996 = ~n4393 & ~n4995;
  assign n4997 = reg_i_RtoB_ACK1_out & ~n4996;
  assign n4998 = ~n1969 & ~n4418;
  assign n4999 = fair_cnt<0>_out  & ~n4998;
  assign n5000 = ~n4105 & ~n4189;
  assign n5001 = ~fair_cnt<0>_out  & ~n5000;
  assign n5002 = ~n4999 & ~n5001;
  assign n5003 = env_fair0done_out & ~n5002;
  assign n5004 = ~env_fair0done_out & ~n4968;
  assign n5005 = ~n5003 & ~n5004;
  assign n5006 = ~reg_stateG7_0_out & ~n5005;
  assign n5007 = ~reg_stateG7_0_out & ~n5006;
  assign n5008 = reg_nstateG7_1_out & ~n5007;
  assign n5009 = ~reg_nstateG7_1_out & ~n5005;
  assign n5010 = ~n5008 & ~n5009;
  assign n5011 = ~reg_controllable_BtoR_REQ1_out & ~n5010;
  assign n5012 = ~reg_controllable_BtoR_REQ1_out & ~n5011;
  assign n5013 = reg_controllable_BtoR_REQ0_out & ~n5012;
  assign n5014 = env_fair1done_out & ~n5002;
  assign n5015 = ~env_fair1done_out & ~n4968;
  assign n5016 = ~n5014 & ~n5015;
  assign n5017 = reg_nstateG7_1_out & ~n5016;
  assign n5018 = ~reg_stateG7_0_out & ~n5016;
  assign n5019 = ~reg_stateG7_0_out & ~n5018;
  assign n5020 = ~reg_nstateG7_1_out & ~n5019;
  assign n5021 = ~n5017 & ~n5020;
  assign n5022 = reg_controllable_BtoR_REQ1_out & ~n5021;
  assign n5023 = fair_cnt<0>_out  & ~n5000;
  assign n5024 = ~n4191 & ~n5023;
  assign n5025 = ~env_fair1done_out & ~n5024;
  assign n5026 = ~n5014 & ~n5025;
  assign n5027 = reg_nstateG7_1_out & ~n5026;
  assign n5028 = ~env_fair0done_out & ~n5024;
  assign n5029 = ~n5003 & ~n5028;
  assign n5030 = ~reg_nstateG7_1_out & ~n5029;
  assign n5031 = ~n5027 & ~n5030;
  assign n5032 = ~reg_controllable_BtoR_REQ1_out & ~n5031;
  assign n5033 = ~n5022 & ~n5032;
  assign n5034 = ~reg_controllable_BtoR_REQ0_out & ~n5033;
  assign n5035 = ~n5013 & ~n5034;
  assign n5036 = ~reg_i_RtoB_ACK1_out & ~n5035;
  assign n5037 = ~n4997 & ~n5036;
  assign n5038 = ~reg_i_RtoB_ACK0_out & ~n5037;
  assign n5039 = ~n4984 & ~n5038;
  assign n5040 = ~reg_i_StoB_REQ9_out & ~n5039;
  assign n5041 = ~n4965 & ~n5040;
  assign n5042 = reg_controllable_BtoS_ACK9_out & ~n5041;
  assign n5043 = ~n4671 & ~n4685;
  assign n5044 = env_fair0done_out & ~n5043;
  assign n5045 = ~n4674 & ~n5044;
  assign n5046 = ~reg_stateG7_0_out & ~n5045;
  assign n5047 = ~reg_stateG7_0_out & ~n5046;
  assign n5048 = reg_nstateG7_1_out & ~n5047;
  assign n5049 = ~reg_nstateG7_1_out & ~n5045;
  assign n5050 = ~n5048 & ~n5049;
  assign n5051 = ~reg_controllable_BtoR_REQ1_out & ~n5050;
  assign n5052 = ~reg_controllable_BtoR_REQ1_out & ~n5051;
  assign n5053 = reg_controllable_BtoR_REQ0_out & ~n5052;
  assign n5054 = ~n4699 & ~n5053;
  assign n5055 = ~reg_i_RtoB_ACK1_out & ~n5054;
  assign n5056 = ~n4667 & ~n5055;
  assign n5057 = reg_i_RtoB_ACK0_out & ~n5056;
  assign n5058 = reg_nstateG7_1_out & ~n5045;
  assign n5059 = ~reg_nstateG7_1_out & ~n5047;
  assign n5060 = ~n5058 & ~n5059;
  assign n5061 = reg_controllable_BtoR_REQ1_out & ~n5060;
  assign n5062 = ~n4722 & ~n5061;
  assign n5063 = ~reg_controllable_BtoR_REQ0_out & ~n5062;
  assign n5064 = ~n4714 & ~n5063;
  assign n5065 = reg_i_RtoB_ACK1_out & ~n5064;
  assign n5066 = ~n2927 & ~n4418;
  assign n5067 = fair_cnt<0>_out  & ~n5066;
  assign n5068 = ~n4191 & ~n5067;
  assign n5069 = env_fair0done_out & ~n5068;
  assign n5070 = ~env_fair0done_out & ~n4684;
  assign n5071 = ~n5069 & ~n5070;
  assign n5072 = ~reg_stateG7_0_out & ~n5071;
  assign n5073 = ~reg_stateG7_0_out & ~n5072;
  assign n5074 = reg_nstateG7_1_out & ~n5073;
  assign n5075 = ~reg_nstateG7_1_out & ~n5071;
  assign n5076 = ~n5074 & ~n5075;
  assign n5077 = ~reg_controllable_BtoR_REQ1_out & ~n5076;
  assign n5078 = ~reg_controllable_BtoR_REQ1_out & ~n5077;
  assign n5079 = reg_controllable_BtoR_REQ0_out & ~n5078;
  assign n5080 = env_fair1done_out & ~n5068;
  assign n5081 = ~env_fair1done_out & ~n4684;
  assign n5082 = ~n5080 & ~n5081;
  assign n5083 = reg_nstateG7_1_out & ~n5082;
  assign n5084 = ~reg_stateG7_0_out & ~n5082;
  assign n5085 = ~reg_stateG7_0_out & ~n5084;
  assign n5086 = ~reg_nstateG7_1_out & ~n5085;
  assign n5087 = ~n5083 & ~n5086;
  assign n5088 = reg_controllable_BtoR_REQ1_out & ~n5087;
  assign n5089 = ~env_fair1done_out & ~n4190;
  assign n5090 = ~n5080 & ~n5089;
  assign n5091 = reg_nstateG7_1_out & ~n5090;
  assign n5092 = ~env_fair0done_out & ~n4190;
  assign n5093 = ~n5069 & ~n5092;
  assign n5094 = ~reg_nstateG7_1_out & ~n5093;
  assign n5095 = ~n5091 & ~n5094;
  assign n5096 = ~reg_controllable_BtoR_REQ1_out & ~n5095;
  assign n5097 = ~n5088 & ~n5096;
  assign n5098 = ~reg_controllable_BtoR_REQ0_out & ~n5097;
  assign n5099 = ~n5079 & ~n5098;
  assign n5100 = ~reg_i_RtoB_ACK1_out & ~n5099;
  assign n5101 = ~n5065 & ~n5100;
  assign n5102 = ~reg_i_RtoB_ACK0_out & ~n5101;
  assign n5103 = ~n5057 & ~n5102;
  assign n5104 = reg_i_StoB_REQ9_out & ~n5103;
  assign n5105 = ~n3124 & ~n4105;
  assign n5106 = fair_cnt<0>_out  & ~n5105;
  assign n5107 = ~n4191 & ~n5106;
  assign n5108 = env_fair1done_out & ~n5107;
  assign n5109 = ~n4259 & ~n5108;
  assign n5110 = env_fair0done_out & ~n5109;
  assign n5111 = ~n4264 & ~n5110;
  assign n5112 = ~reg_stateG7_0_out & ~n5111;
  assign n5113 = ~reg_stateG7_0_out & ~n5112;
  assign n5114 = reg_nstateG7_1_out & ~n5113;
  assign n5115 = ~reg_nstateG7_1_out & ~n5111;
  assign n5116 = ~n5114 & ~n5115;
  assign n5117 = ~reg_controllable_BtoR_REQ1_out & ~n5116;
  assign n5118 = ~reg_controllable_BtoR_REQ1_out & ~n5117;
  assign n5119 = reg_controllable_BtoR_REQ0_out & ~n5118;
  assign n5120 = ~n4841 & ~n5119;
  assign n5121 = ~reg_i_RtoB_ACK1_out & ~n5120;
  assign n5122 = ~n4808 & ~n5121;
  assign n5123 = reg_i_RtoB_ACK0_out & ~n5122;
  assign n5124 = ~n4394 & ~n5108;
  assign n5125 = env_fair0done_out & ~n5124;
  assign n5126 = ~n4399 & ~n5125;
  assign n5127 = reg_nstateG7_1_out & ~n5126;
  assign n5128 = ~reg_stateG7_0_out & ~n5126;
  assign n5129 = ~reg_stateG7_0_out & ~n5128;
  assign n5130 = ~reg_nstateG7_1_out & ~n5129;
  assign n5131 = ~n5127 & ~n5130;
  assign n5132 = reg_controllable_BtoR_REQ1_out & ~n5131;
  assign n5133 = ~n4871 & ~n5132;
  assign n5134 = ~reg_controllable_BtoR_REQ0_out & ~n5133;
  assign n5135 = ~n4856 & ~n5134;
  assign n5136 = reg_i_RtoB_ACK1_out & ~n5135;
  assign n5137 = ~n3124 & ~n4418;
  assign n5138 = fair_cnt<0>_out  & ~n5137;
  assign n5139 = ~n5001 & ~n5138;
  assign n5140 = env_fair0done_out & ~n5139;
  assign n5141 = ~env_fair0done_out & ~n5107;
  assign n5142 = ~n5140 & ~n5141;
  assign n5143 = ~reg_stateG7_0_out & ~n5142;
  assign n5144 = ~reg_stateG7_0_out & ~n5143;
  assign n5145 = reg_nstateG7_1_out & ~n5144;
  assign n5146 = ~reg_nstateG7_1_out & ~n5142;
  assign n5147 = ~n5145 & ~n5146;
  assign n5148 = ~reg_controllable_BtoR_REQ1_out & ~n5147;
  assign n5149 = ~reg_controllable_BtoR_REQ1_out & ~n5148;
  assign n5150 = reg_controllable_BtoR_REQ0_out & ~n5149;
  assign n5151 = env_fair1done_out & ~n5139;
  assign n5152 = ~env_fair1done_out & ~n5107;
  assign n5153 = ~n5151 & ~n5152;
  assign n5154 = reg_nstateG7_1_out & ~n5153;
  assign n5155 = ~reg_stateG7_0_out & ~n5153;
  assign n5156 = ~reg_stateG7_0_out & ~n5155;
  assign n5157 = ~reg_nstateG7_1_out & ~n5156;
  assign n5158 = ~n5154 & ~n5157;
  assign n5159 = reg_controllable_BtoR_REQ1_out & ~n5158;
  assign n5160 = ~n5025 & ~n5151;
  assign n5161 = reg_nstateG7_1_out & ~n5160;
  assign n5162 = ~n5028 & ~n5140;
  assign n5163 = ~reg_nstateG7_1_out & ~n5162;
  assign n5164 = ~n5161 & ~n5163;
  assign n5165 = ~reg_controllable_BtoR_REQ1_out & ~n5164;
  assign n5166 = ~n5159 & ~n5165;
  assign n5167 = ~reg_controllable_BtoR_REQ0_out & ~n5166;
  assign n5168 = ~n5150 & ~n5167;
  assign n5169 = ~reg_i_RtoB_ACK1_out & ~n5168;
  assign n5170 = ~n5136 & ~n5169;
  assign n5171 = ~reg_i_RtoB_ACK0_out & ~n5170;
  assign n5172 = ~n5123 & ~n5171;
  assign n5173 = ~reg_i_StoB_REQ9_out & ~n5172;
  assign n5174 = ~n5104 & ~n5173;
  assign n5175 = ~reg_controllable_BtoS_ACK9_out & ~n5174;
  assign n5176 = ~n5042 & ~n5175;
  assign n5177 = reg_i_nEMPTY_out & ~n5176;
  assign n5178 = ~fair_cnt<1>_out  & ~n3831;
  assign n5179 = ~n671 & ~n5178;
  assign n5180 = fair_cnt<0>_out  & ~n5179;
  assign n5181 = ~fair_cnt<1>_out  & ~n4007;
  assign n5182 = ~n3832 & ~n5181;
  assign n5183 = ~fair_cnt<0>_out  & ~n5182;
  assign n5184 = ~n5180 & ~n5183;
  assign n5185 = env_fair0done_out & ~n5184;
  assign n5186 = ~n671 & ~n5181;
  assign n5187 = fair_cnt<0>_out  & ~n5186;
  assign n5188 = ~n3834 & ~n5187;
  assign n5189 = ~env_fair0done_out & ~n5188;
  assign n5190 = ~n5185 & ~n5189;
  assign n5191 = ~reg_stateG7_0_out & ~n5190;
  assign n5192 = ~reg_stateG7_0_out & ~n5191;
  assign n5193 = reg_nstateG7_1_out & ~n5192;
  assign n5194 = ~reg_nstateG7_1_out & ~n5190;
  assign n5195 = ~n5193 & ~n5194;
  assign n5196 = ~reg_controllable_BtoR_REQ1_out & ~n5195;
  assign n5197 = ~reg_controllable_BtoR_REQ1_out & ~n5196;
  assign n5198 = reg_controllable_BtoR_REQ0_out & ~n5197;
  assign n5199 = env_fair1done_out & ~n5184;
  assign n5200 = ~env_fair1done_out & ~n5188;
  assign n5201 = ~n5199 & ~n5200;
  assign n5202 = reg_nstateG7_1_out & ~n5201;
  assign n5203 = ~reg_stateG7_0_out & ~n5201;
  assign n5204 = ~reg_stateG7_0_out & ~n5203;
  assign n5205 = ~reg_nstateG7_1_out & ~n5204;
  assign n5206 = ~n5202 & ~n5205;
  assign n5207 = reg_controllable_BtoR_REQ1_out & ~n5206;
  assign n5208 = reg_stateG12_out & ~n502;
  assign n5209 = ~reg_stateG12_out & ~n125;
  assign n5210 = ~n5208 & ~n5209;
  assign n5211 = sys_fair12done_out & ~n5210;
  assign n5212 = ~n131 & ~n507;
  assign n5213 = ~sys_fair12done_out & ~n5212;
  assign n5214 = ~n5211 & ~n5213;
  assign n5215 = sys_fair2done_out & ~n5214;
  assign n5216 = reg_stateG12_out & ~n379;
  assign n5217 = ~n131 & ~n5216;
  assign n5218 = ~sys_fair2done_out & ~n5217;
  assign n5219 = ~n5215 & ~n5218;
  assign n5220 = reg_controllable_BtoS_ACK2_out & ~n5219;
  assign n5221 = ~reg_stateG12_out & ~n129;
  assign n5222 = ~n507 & ~n5221;
  assign n5223 = sys_fair12done_out & ~n5222;
  assign n5224 = ~n5213 & ~n5223;
  assign n5225 = ~sys_fair2done_out & ~n5224;
  assign n5226 = ~n5215 & ~n5225;
  assign n5227 = ~reg_controllable_BtoS_ACK2_out & ~n5226;
  assign n5228 = ~n5220 & ~n5227;
  assign n5229 = ~reg_i_StoB_REQ2_out & ~n5228;
  assign n5230 = ~n142 & ~n5229;
  assign n5231 = sys_fair3done_out & ~n5230;
  assign n5232 = ~reg_i_StoB_REQ2_out & ~n5217;
  assign n5233 = ~n166 & ~n5232;
  assign n5234 = ~sys_fair3done_out & ~n5233;
  assign n5235 = ~n5231 & ~n5234;
  assign n5236 = reg_controllable_BtoS_ACK3_out & ~n5235;
  assign n5237 = sys_fair2done_out & ~n5224;
  assign n5238 = ~n5218 & ~n5237;
  assign n5239 = reg_controllable_BtoS_ACK2_out & ~n5238;
  assign n5240 = ~reg_controllable_BtoS_ACK2_out & ~n5224;
  assign n5241 = ~n5239 & ~n5240;
  assign n5242 = ~reg_i_StoB_REQ2_out & ~n5241;
  assign n5243 = ~n152 & ~n5242;
  assign n5244 = ~sys_fair3done_out & ~n5243;
  assign n5245 = ~n5231 & ~n5244;
  assign n5246 = ~reg_controllable_BtoS_ACK3_out & ~n5245;
  assign n5247 = ~n5236 & ~n5246;
  assign n5248 = ~reg_i_StoB_REQ3_out & ~n5247;
  assign n5249 = ~n163 & ~n5248;
  assign n5250 = ~reg_i_StoB_REQ4_out & ~n5249;
  assign n5251 = ~n177 & ~n5250;
  assign n5252 = sys_fair4done_out & ~n5251;
  assign n5253 = ~reg_i_StoB_REQ3_out & ~n5233;
  assign n5254 = ~n195 & ~n5253;
  assign n5255 = reg_controllable_BtoS_ACK4_out & ~n5254;
  assign n5256 = sys_fair3done_out & ~n5243;
  assign n5257 = ~n5234 & ~n5256;
  assign n5258 = reg_controllable_BtoS_ACK3_out & ~n5257;
  assign n5259 = ~reg_controllable_BtoS_ACK3_out & ~n5243;
  assign n5260 = ~n5258 & ~n5259;
  assign n5261 = ~reg_i_StoB_REQ3_out & ~n5260;
  assign n5262 = ~n183 & ~n5261;
  assign n5263 = ~reg_controllable_BtoS_ACK4_out & ~n5262;
  assign n5264 = ~n5255 & ~n5263;
  assign n5265 = ~reg_i_StoB_REQ4_out & ~n5264;
  assign n5266 = ~n192 & ~n5265;
  assign n5267 = ~sys_fair4done_out & ~n5266;
  assign n5268 = ~n5252 & ~n5267;
  assign n5269 = ~reg_i_StoB_REQ5_out & ~n5268;
  assign n5270 = ~n206 & ~n5269;
  assign n5271 = sys_fair5done_out & ~n5270;
  assign n5272 = ~reg_i_StoB_REQ4_out & ~n5254;
  assign n5273 = ~n219 & ~n5272;
  assign n5274 = reg_controllable_BtoS_ACK5_out & ~n5273;
  assign n5275 = ~reg_i_StoB_REQ4_out & ~n5262;
  assign n5276 = ~n192 & ~n5275;
  assign n5277 = sys_fair4done_out & ~n5276;
  assign n5278 = ~n5267 & ~n5277;
  assign n5279 = ~reg_controllable_BtoS_ACK5_out & ~n5278;
  assign n5280 = ~n5274 & ~n5279;
  assign n5281 = ~reg_i_StoB_REQ5_out & ~n5280;
  assign n5282 = ~n216 & ~n5281;
  assign n5283 = ~sys_fair5done_out & ~n5282;
  assign n5284 = ~n5271 & ~n5283;
  assign n5285 = ~reg_i_StoB_REQ6_out & ~n5284;
  assign n5286 = ~n230 & ~n5285;
  assign n5287 = sys_fair6done_out & ~n5286;
  assign n5288 = ~reg_i_StoB_REQ5_out & ~n5273;
  assign n5289 = ~n243 & ~n5288;
  assign n5290 = reg_controllable_BtoS_ACK6_out & ~n5289;
  assign n5291 = ~reg_i_StoB_REQ5_out & ~n5278;
  assign n5292 = ~n216 & ~n5291;
  assign n5293 = sys_fair5done_out & ~n5292;
  assign n5294 = ~n5283 & ~n5293;
  assign n5295 = ~reg_controllable_BtoS_ACK6_out & ~n5294;
  assign n5296 = ~n5290 & ~n5295;
  assign n5297 = ~reg_i_StoB_REQ6_out & ~n5296;
  assign n5298 = ~n240 & ~n5297;
  assign n5299 = ~sys_fair6done_out & ~n5298;
  assign n5300 = ~n5287 & ~n5299;
  assign n5301 = ~reg_i_StoB_REQ7_out & ~n5300;
  assign n5302 = ~n254 & ~n5301;
  assign n5303 = sys_fair7done_out & ~n5302;
  assign n5304 = ~reg_i_StoB_REQ6_out & ~n5289;
  assign n5305 = ~n267 & ~n5304;
  assign n5306 = reg_controllable_BtoS_ACK7_out & ~n5305;
  assign n5307 = ~reg_i_StoB_REQ6_out & ~n5294;
  assign n5308 = ~n240 & ~n5307;
  assign n5309 = sys_fair6done_out & ~n5308;
  assign n5310 = ~n5299 & ~n5309;
  assign n5311 = ~reg_controllable_BtoS_ACK7_out & ~n5310;
  assign n5312 = ~n5306 & ~n5311;
  assign n5313 = ~reg_i_StoB_REQ7_out & ~n5312;
  assign n5314 = ~n264 & ~n5313;
  assign n5315 = ~sys_fair7done_out & ~n5314;
  assign n5316 = ~n5303 & ~n5315;
  assign n5317 = sys_fair8done_out & ~n5316;
  assign n5318 = ~reg_i_StoB_REQ7_out & ~n5305;
  assign n5319 = ~n288 & ~n5318;
  assign n5320 = ~sys_fair8done_out & ~n5319;
  assign n5321 = ~n5317 & ~n5320;
  assign n5322 = reg_controllable_BtoS_ACK8_out & ~n5321;
  assign n5323 = ~reg_i_StoB_REQ7_out & ~n5310;
  assign n5324 = ~n264 & ~n5323;
  assign n5325 = sys_fair7done_out & ~n5324;
  assign n5326 = ~n5315 & ~n5325;
  assign n5327 = ~sys_fair8done_out & ~n5326;
  assign n5328 = ~n5317 & ~n5327;
  assign n5329 = ~reg_controllable_BtoS_ACK8_out & ~n5328;
  assign n5330 = ~n5322 & ~n5329;
  assign n5331 = ~reg_i_StoB_REQ8_out & ~n5330;
  assign n5332 = ~n285 & ~n5331;
  assign n5333 = ~reg_i_StoB_REQ10_out & ~n5332;
  assign n5334 = ~n299 & ~n5333;
  assign n5335 = sys_fair10done_out & ~n5334;
  assign n5336 = ~reg_i_StoB_REQ8_out & ~n5319;
  assign n5337 = ~n317 & ~n5336;
  assign n5338 = reg_controllable_BtoS_ACK10_out & ~n5337;
  assign n5339 = sys_fair8done_out & ~n5326;
  assign n5340 = ~n5320 & ~n5339;
  assign n5341 = reg_controllable_BtoS_ACK8_out & ~n5340;
  assign n5342 = ~reg_controllable_BtoS_ACK8_out & ~n5326;
  assign n5343 = ~n5341 & ~n5342;
  assign n5344 = ~reg_i_StoB_REQ8_out & ~n5343;
  assign n5345 = ~n305 & ~n5344;
  assign n5346 = ~reg_controllable_BtoS_ACK10_out & ~n5345;
  assign n5347 = ~n5338 & ~n5346;
  assign n5348 = ~reg_i_StoB_REQ10_out & ~n5347;
  assign n5349 = ~n314 & ~n5348;
  assign n5350 = ~sys_fair10done_out & ~n5349;
  assign n5351 = ~n5335 & ~n5350;
  assign n5352 = sys_fair11done_out & ~n5351;
  assign n5353 = ~reg_i_StoB_REQ10_out & ~n5337;
  assign n5354 = ~n338 & ~n5353;
  assign n5355 = ~sys_fair11done_out & ~n5354;
  assign n5356 = ~n5352 & ~n5355;
  assign n5357 = reg_controllable_BtoS_ACK11_out & ~n5356;
  assign n5358 = ~reg_i_StoB_REQ10_out & ~n5345;
  assign n5359 = ~n314 & ~n5358;
  assign n5360 = sys_fair10done_out & ~n5359;
  assign n5361 = ~n5350 & ~n5360;
  assign n5362 = ~sys_fair11done_out & ~n5361;
  assign n5363 = ~n5352 & ~n5362;
  assign n5364 = ~reg_controllable_BtoS_ACK11_out & ~n5363;
  assign n5365 = ~n5357 & ~n5364;
  assign n5366 = ~reg_i_StoB_REQ11_out & ~n5365;
  assign n5367 = ~n335 & ~n5366;
  assign n5368 = sys_fair9done_out & ~n5367;
  assign n5369 = sys_fair11done_out & ~n5361;
  assign n5370 = ~n5355 & ~n5369;
  assign n5371 = reg_controllable_BtoS_ACK11_out & ~n5370;
  assign n5372 = ~reg_controllable_BtoS_ACK11_out & ~n5361;
  assign n5373 = ~n5371 & ~n5372;
  assign n5374 = ~reg_i_StoB_REQ11_out & ~n5373;
  assign n5375 = ~n350 & ~n5374;
  assign n5376 = ~sys_fair9done_out & ~n5375;
  assign n5377 = ~n5368 & ~n5376;
  assign n5378 = fair_cnt<1>_out  & ~n5377;
  assign n5379 = sys_fair12done_out & ~n5217;
  assign n5380 = ~n131 & ~n3785;
  assign n5381 = ~sys_fair12done_out & ~n5380;
  assign n5382 = ~n5379 & ~n5381;
  assign n5383 = sys_fair2done_out & ~n5382;
  assign n5384 = ~n5218 & ~n5383;
  assign n5385 = ~reg_i_StoB_REQ2_out & ~n5384;
  assign n5386 = ~n3695 & ~n5385;
  assign n5387 = sys_fair3done_out & ~n5386;
  assign n5388 = ~n5234 & ~n5387;
  assign n5389 = ~reg_i_StoB_REQ3_out & ~n5388;
  assign n5390 = ~n3702 & ~n5389;
  assign n5391 = ~reg_i_StoB_REQ4_out & ~n5390;
  assign n5392 = ~n3707 & ~n5391;
  assign n5393 = sys_fair4done_out & ~n5392;
  assign n5394 = ~sys_fair4done_out & ~n5273;
  assign n5395 = ~n5393 & ~n5394;
  assign n5396 = ~reg_i_StoB_REQ5_out & ~n5395;
  assign n5397 = ~n3714 & ~n5396;
  assign n5398 = sys_fair5done_out & ~n5397;
  assign n5399 = ~sys_fair5done_out & ~n5289;
  assign n5400 = ~n5398 & ~n5399;
  assign n5401 = ~reg_i_StoB_REQ6_out & ~n5400;
  assign n5402 = ~n3721 & ~n5401;
  assign n5403 = sys_fair6done_out & ~n5402;
  assign n5404 = ~sys_fair6done_out & ~n5305;
  assign n5405 = ~n5403 & ~n5404;
  assign n5406 = ~reg_i_StoB_REQ7_out & ~n5405;
  assign n5407 = ~n3728 & ~n5406;
  assign n5408 = sys_fair7done_out & ~n5407;
  assign n5409 = ~sys_fair7done_out & ~n5319;
  assign n5410 = ~n5408 & ~n5409;
  assign n5411 = sys_fair8done_out & ~n5410;
  assign n5412 = ~n5320 & ~n5411;
  assign n5413 = ~reg_i_StoB_REQ8_out & ~n5412;
  assign n5414 = ~n3737 & ~n5413;
  assign n5415 = ~reg_i_StoB_REQ10_out & ~n5414;
  assign n5416 = ~n3742 & ~n5415;
  assign n5417 = sys_fair10done_out & ~n5416;
  assign n5418 = ~sys_fair10done_out & ~n5354;
  assign n5419 = ~n5417 & ~n5418;
  assign n5420 = sys_fair11done_out & ~n5419;
  assign n5421 = ~n5355 & ~n5420;
  assign n5422 = ~reg_i_StoB_REQ11_out & ~n5421;
  assign n5423 = ~n3751 & ~n5422;
  assign n5424 = sys_fair9done_out & ~n5423;
  assign n5425 = ~reg_i_StoB_REQ11_out & ~n5354;
  assign n5426 = ~n362 & ~n5425;
  assign n5427 = ~sys_fair9done_out & ~n5426;
  assign n5428 = ~n5424 & ~n5427;
  assign n5429 = ~fair_cnt<1>_out  & ~n5428;
  assign n5430 = ~n5378 & ~n5429;
  assign n5431 = fair_cnt<0>_out  & ~n5430;
  assign n5432 = fair_cnt<1>_out  & ~n5428;
  assign n5433 = ~n131 & ~n3465;
  assign n5434 = ~sys_fair12done_out & ~n5433;
  assign n5435 = ~n5379 & ~n5434;
  assign n5436 = sys_fair2done_out & ~n5435;
  assign n5437 = ~n5218 & ~n5436;
  assign n5438 = ~reg_i_StoB_REQ2_out & ~n5437;
  assign n5439 = ~n3968 & ~n5438;
  assign n5440 = sys_fair3done_out & ~n5439;
  assign n5441 = ~n5234 & ~n5440;
  assign n5442 = ~reg_i_StoB_REQ3_out & ~n5441;
  assign n5443 = ~n3965 & ~n5442;
  assign n5444 = ~reg_i_StoB_REQ4_out & ~n5443;
  assign n5445 = ~n3962 & ~n5444;
  assign n5446 = sys_fair4done_out & ~n5445;
  assign n5447 = ~n5394 & ~n5446;
  assign n5448 = ~reg_i_StoB_REQ5_out & ~n5447;
  assign n5449 = ~n3959 & ~n5448;
  assign n5450 = sys_fair5done_out & ~n5449;
  assign n5451 = ~n5399 & ~n5450;
  assign n5452 = ~reg_i_StoB_REQ6_out & ~n5451;
  assign n5453 = ~n3956 & ~n5452;
  assign n5454 = sys_fair6done_out & ~n5453;
  assign n5455 = ~n5404 & ~n5454;
  assign n5456 = ~reg_i_StoB_REQ7_out & ~n5455;
  assign n5457 = ~n3953 & ~n5456;
  assign n5458 = sys_fair7done_out & ~n5457;
  assign n5459 = ~n5409 & ~n5458;
  assign n5460 = sys_fair8done_out & ~n5459;
  assign n5461 = ~n5320 & ~n5460;
  assign n5462 = ~reg_i_StoB_REQ8_out & ~n5461;
  assign n5463 = ~n3950 & ~n5462;
  assign n5464 = ~reg_i_StoB_REQ10_out & ~n5463;
  assign n5465 = ~n3947 & ~n5464;
  assign n5466 = sys_fair10done_out & ~n5465;
  assign n5467 = ~n5418 & ~n5466;
  assign n5468 = sys_fair11done_out & ~n5467;
  assign n5469 = ~n5355 & ~n5468;
  assign n5470 = ~reg_i_StoB_REQ11_out & ~n5469;
  assign n5471 = ~n3944 & ~n5470;
  assign n5472 = sys_fair9done_out & ~n5471;
  assign n5473 = ~n5427 & ~n5472;
  assign n5474 = ~fair_cnt<1>_out  & ~n5473;
  assign n5475 = ~n5432 & ~n5474;
  assign n5476 = ~fair_cnt<0>_out  & ~n5475;
  assign n5477 = ~n5431 & ~n5476;
  assign n5478 = env_fair1done_out & ~n5477;
  assign n5479 = ~reg_stateG12_out & ~n385;
  assign n5480 = ~n5216 & ~n5479;
  assign n5481 = sys_fair12done_out & ~n5480;
  assign n5482 = ~sys_fair12done_out & ~n5217;
  assign n5483 = ~n5481 & ~n5482;
  assign n5484 = sys_fair2done_out & ~n5483;
  assign n5485 = ~n5218 & ~n5484;
  assign n5486 = ~reg_i_StoB_REQ2_out & ~n5485;
  assign n5487 = ~n166 & ~n5486;
  assign n5488 = sys_fair3done_out & ~n5487;
  assign n5489 = ~n5234 & ~n5488;
  assign n5490 = ~reg_i_StoB_REQ3_out & ~n5489;
  assign n5491 = ~n195 & ~n5490;
  assign n5492 = ~reg_i_StoB_REQ4_out & ~n5491;
  assign n5493 = ~n219 & ~n5492;
  assign n5494 = sys_fair4done_out & ~n5493;
  assign n5495 = ~n5394 & ~n5494;
  assign n5496 = ~reg_i_StoB_REQ5_out & ~n5495;
  assign n5497 = ~n243 & ~n5496;
  assign n5498 = sys_fair5done_out & ~n5497;
  assign n5499 = ~n5399 & ~n5498;
  assign n5500 = ~reg_i_StoB_REQ6_out & ~n5499;
  assign n5501 = ~n267 & ~n5500;
  assign n5502 = sys_fair6done_out & ~n5501;
  assign n5503 = ~n5404 & ~n5502;
  assign n5504 = ~reg_i_StoB_REQ7_out & ~n5503;
  assign n5505 = ~n288 & ~n5504;
  assign n5506 = sys_fair7done_out & ~n5505;
  assign n5507 = ~n5409 & ~n5506;
  assign n5508 = sys_fair8done_out & ~n5507;
  assign n5509 = ~n5320 & ~n5508;
  assign n5510 = ~reg_i_StoB_REQ8_out & ~n5509;
  assign n5511 = ~n317 & ~n5510;
  assign n5512 = ~reg_i_StoB_REQ10_out & ~n5511;
  assign n5513 = ~n338 & ~n5512;
  assign n5514 = sys_fair10done_out & ~n5513;
  assign n5515 = ~n5418 & ~n5514;
  assign n5516 = sys_fair11done_out & ~n5515;
  assign n5517 = ~n5355 & ~n5516;
  assign n5518 = ~reg_i_StoB_REQ11_out & ~n5517;
  assign n5519 = ~n362 & ~n5518;
  assign n5520 = ~sys_fair9done_out & ~n5519;
  assign n5521 = ~n5424 & ~n5520;
  assign n5522 = fair_cnt<1>_out  & ~n5521;
  assign n5523 = ~n5474 & ~n5522;
  assign n5524 = fair_cnt<0>_out  & ~n5523;
  assign n5525 = ~fair_cnt<1>_out  & ~n5426;
  assign n5526 = ~n5432 & ~n5525;
  assign n5527 = ~fair_cnt<0>_out  & ~n5526;
  assign n5528 = ~n5524 & ~n5527;
  assign n5529 = ~env_fair1done_out & ~n5528;
  assign n5530 = ~n5478 & ~n5529;
  assign n5531 = reg_nstateG7_1_out & ~n5530;
  assign n5532 = env_fair0done_out & ~n5477;
  assign n5533 = ~env_fair0done_out & ~n5528;
  assign n5534 = ~n5532 & ~n5533;
  assign n5535 = ~reg_nstateG7_1_out & ~n5534;
  assign n5536 = ~n5531 & ~n5535;
  assign n5537 = ~reg_controllable_BtoR_REQ1_out & ~n5536;
  assign n5538 = ~n5207 & ~n5537;
  assign n5539 = ~reg_controllable_BtoR_REQ0_out & ~n5538;
  assign n5540 = ~n5198 & ~n5539;
  assign n5541 = ~reg_i_RtoB_ACK1_out & ~n5540;
  assign n5542 = ~reg_i_RtoB_ACK1_out & ~n5541;
  assign n5543 = ~reg_i_RtoB_ACK0_out & ~n5542;
  assign n5544 = ~reg_i_RtoB_ACK0_out & ~n5543;
  assign n5545 = reg_i_StoB_REQ9_out & ~n5544;
  assign n5546 = ~n1264 & ~n5181;
  assign n5547 = fair_cnt<0>_out  & ~n5546;
  assign n5548 = ~n3834 & ~n5547;
  assign n5549 = env_fair1done_out & ~n5548;
  assign n5550 = ~n4010 & ~n5547;
  assign n5551 = ~env_fair1done_out & ~n5550;
  assign n5552 = ~n5549 & ~n5551;
  assign n5553 = env_fair0done_out & ~n5552;
  assign n5554 = ~env_fair0done_out & ~n4011;
  assign n5555 = ~n5553 & ~n5554;
  assign n5556 = ~reg_stateG7_0_out & ~n5555;
  assign n5557 = ~reg_stateG7_0_out & ~n5556;
  assign n5558 = reg_nstateG7_1_out & ~n5557;
  assign n5559 = ~reg_nstateG7_1_out & ~n5555;
  assign n5560 = ~n5558 & ~n5559;
  assign n5561 = ~reg_controllable_BtoR_REQ1_out & ~n5560;
  assign n5562 = ~reg_controllable_BtoR_REQ1_out & ~n5561;
  assign n5563 = reg_controllable_BtoR_REQ0_out & ~n5562;
  assign n5564 = reg_controllable_BtoR_REQ0_out & ~n5563;
  assign n5565 = ~reg_i_RtoB_ACK1_out & ~n5564;
  assign n5566 = ~reg_i_RtoB_ACK1_out & ~n5565;
  assign n5567 = reg_i_RtoB_ACK0_out & ~n5566;
  assign n5568 = ~env_fair1done_out & ~n4011;
  assign n5569 = ~n5549 & ~n5568;
  assign n5570 = env_fair0done_out & ~n5569;
  assign n5571 = env_fair1done_out & ~n5550;
  assign n5572 = ~n5568 & ~n5571;
  assign n5573 = ~env_fair0done_out & ~n5572;
  assign n5574 = ~n5570 & ~n5573;
  assign n5575 = reg_nstateG7_1_out & ~n5574;
  assign n5576 = ~reg_stateG7_0_out & ~n5574;
  assign n5577 = ~reg_stateG7_0_out & ~n5576;
  assign n5578 = ~reg_nstateG7_1_out & ~n5577;
  assign n5579 = ~n5575 & ~n5578;
  assign n5580 = reg_controllable_BtoR_REQ1_out & ~n5579;
  assign n5581 = reg_controllable_BtoR_REQ1_out & ~n5580;
  assign n5582 = ~reg_controllable_BtoR_REQ0_out & ~n5581;
  assign n5583 = ~reg_controllable_BtoR_REQ0_out & ~n5582;
  assign n5584 = reg_i_RtoB_ACK1_out & ~n5583;
  assign n5585 = ~fair_cnt<1>_out  & ~n4353;
  assign n5586 = ~n2551 & ~n5585;
  assign n5587 = fair_cnt<0>_out  & ~n5586;
  assign n5588 = reg_controllable_BtoS_ACK11_out & ~n4003;
  assign n5589 = ~reg_controllable_BtoS_ACK11_out & ~n4091;
  assign n5590 = ~n5588 & ~n5589;
  assign n5591 = reg_i_StoB_REQ11_out & ~n5590;
  assign n5592 = reg_controllable_BtoS_ACK10_out & ~n3997;
  assign n5593 = ~reg_controllable_BtoS_ACK10_out & ~n4084;
  assign n5594 = ~n5592 & ~n5593;
  assign n5595 = reg_i_StoB_REQ10_out & ~n5594;
  assign n5596 = reg_controllable_BtoS_ACK8_out & ~n3995;
  assign n5597 = ~reg_controllable_BtoS_ACK8_out & ~n4082;
  assign n5598 = ~n5596 & ~n5597;
  assign n5599 = reg_i_StoB_REQ8_out & ~n5598;
  assign n5600 = reg_controllable_BtoS_ACK7_out & ~n3989;
  assign n5601 = ~reg_controllable_BtoS_ACK7_out & ~n4075;
  assign n5602 = ~n5600 & ~n5601;
  assign n5603 = reg_i_StoB_REQ7_out & ~n5602;
  assign n5604 = reg_controllable_BtoS_ACK6_out & ~n3985;
  assign n5605 = ~reg_controllable_BtoS_ACK6_out & ~n4070;
  assign n5606 = ~n5604 & ~n5605;
  assign n5607 = reg_i_StoB_REQ6_out & ~n5606;
  assign n5608 = reg_controllable_BtoS_ACK5_out & ~n3981;
  assign n5609 = ~reg_controllable_BtoS_ACK5_out & ~n4065;
  assign n5610 = ~n5608 & ~n5609;
  assign n5611 = reg_i_StoB_REQ5_out & ~n5610;
  assign n5612 = reg_controllable_BtoS_ACK4_out & ~n3977;
  assign n5613 = ~reg_controllable_BtoS_ACK4_out & ~n4060;
  assign n5614 = ~n5612 & ~n5613;
  assign n5615 = reg_i_StoB_REQ4_out & ~n5614;
  assign n5616 = reg_controllable_BtoS_ACK3_out & ~n3975;
  assign n5617 = ~reg_controllable_BtoS_ACK3_out & ~n4058;
  assign n5618 = ~n5616 & ~n5617;
  assign n5619 = reg_i_StoB_REQ3_out & ~n5618;
  assign n5620 = reg_controllable_BtoS_ACK2_out & ~n3971;
  assign n5621 = ~reg_controllable_BtoS_ACK2_out & ~n4054;
  assign n5622 = ~n5620 & ~n5621;
  assign n5623 = reg_i_StoB_REQ2_out & ~n5622;
  assign n5624 = ~n3460 & ~n4302;
  assign n5625 = sys_fair1done_out & ~n5624;
  assign n5626 = ~n4305 & ~n5625;
  assign n5627 = reg_stateG12_out & ~n5626;
  assign n5628 = ~n2338 & ~n5627;
  assign n5629 = ~sys_fair12done_out & ~n5628;
  assign n5630 = ~n4301 & ~n5629;
  assign n5631 = sys_fair2done_out & ~n5630;
  assign n5632 = ~n2343 & ~n5631;
  assign n5633 = ~reg_i_StoB_REQ2_out & ~n5632;
  assign n5634 = ~n5623 & ~n5633;
  assign n5635 = sys_fair3done_out & ~n5634;
  assign n5636 = ~n2359 & ~n5635;
  assign n5637 = ~reg_i_StoB_REQ3_out & ~n5636;
  assign n5638 = ~n5619 & ~n5637;
  assign n5639 = ~reg_i_StoB_REQ4_out & ~n5638;
  assign n5640 = ~n5615 & ~n5639;
  assign n5641 = sys_fair4done_out & ~n5640;
  assign n5642 = ~n4322 & ~n5641;
  assign n5643 = ~reg_i_StoB_REQ5_out & ~n5642;
  assign n5644 = ~n5611 & ~n5643;
  assign n5645 = sys_fair5done_out & ~n5644;
  assign n5646 = ~n4327 & ~n5645;
  assign n5647 = ~reg_i_StoB_REQ6_out & ~n5646;
  assign n5648 = ~n5607 & ~n5647;
  assign n5649 = sys_fair6done_out & ~n5648;
  assign n5650 = ~n4332 & ~n5649;
  assign n5651 = ~reg_i_StoB_REQ7_out & ~n5650;
  assign n5652 = ~n5603 & ~n5651;
  assign n5653 = sys_fair7done_out & ~n5652;
  assign n5654 = ~n4337 & ~n5653;
  assign n5655 = sys_fair8done_out & ~n5654;
  assign n5656 = ~n2480 & ~n5655;
  assign n5657 = ~reg_i_StoB_REQ8_out & ~n5656;
  assign n5658 = ~n5599 & ~n5657;
  assign n5659 = ~reg_i_StoB_REQ10_out & ~n5658;
  assign n5660 = ~n5595 & ~n5659;
  assign n5661 = sys_fair10done_out & ~n5660;
  assign n5662 = ~n4346 & ~n5661;
  assign n5663 = sys_fair11done_out & ~n5662;
  assign n5664 = ~n2528 & ~n5663;
  assign n5665 = ~reg_i_StoB_REQ11_out & ~n5664;
  assign n5666 = ~n5591 & ~n5665;
  assign n5667 = sys_fair9done_out & ~n5666;
  assign n5668 = ~n2549 & ~n5667;
  assign n5669 = ~fair_cnt<1>_out  & ~n5668;
  assign n5670 = ~n4354 & ~n5669;
  assign n5671 = ~fair_cnt<0>_out  & ~n5670;
  assign n5672 = ~n5587 & ~n5671;
  assign n5673 = env_fair0done_out & ~n5672;
  assign n5674 = ~n2551 & ~n5669;
  assign n5675 = fair_cnt<0>_out  & ~n5674;
  assign n5676 = ~n4356 & ~n5675;
  assign n5677 = ~env_fair0done_out & ~n5676;
  assign n5678 = ~n5673 & ~n5677;
  assign n5679 = ~reg_stateG7_0_out & ~n5678;
  assign n5680 = ~reg_stateG7_0_out & ~n5679;
  assign n5681 = reg_nstateG7_1_out & ~n5680;
  assign n5682 = ~reg_nstateG7_1_out & ~n5678;
  assign n5683 = ~n5681 & ~n5682;
  assign n5684 = ~reg_controllable_BtoR_REQ1_out & ~n5683;
  assign n5685 = ~reg_controllable_BtoR_REQ1_out & ~n5684;
  assign n5686 = reg_controllable_BtoR_REQ0_out & ~n5685;
  assign n5687 = env_fair1done_out & ~n5672;
  assign n5688 = ~env_fair1done_out & ~n5676;
  assign n5689 = ~n5687 & ~n5688;
  assign n5690 = reg_nstateG7_1_out & ~n5689;
  assign n5691 = ~reg_stateG7_0_out & ~n5689;
  assign n5692 = ~reg_stateG7_0_out & ~n5691;
  assign n5693 = ~reg_nstateG7_1_out & ~n5692;
  assign n5694 = ~n5690 & ~n5693;
  assign n5695 = reg_controllable_BtoR_REQ1_out & ~n5694;
  assign n5696 = reg_controllable_BtoS_ACK11_out & ~n5363;
  assign n5697 = ~n1937 & ~n5696;
  assign n5698 = reg_i_StoB_REQ11_out & ~n5697;
  assign n5699 = reg_controllable_BtoS_ACK10_out & ~n5332;
  assign n5700 = ~n1882 & ~n5699;
  assign n5701 = reg_i_StoB_REQ10_out & ~n5700;
  assign n5702 = reg_controllable_BtoS_ACK8_out & ~n5328;
  assign n5703 = ~n1859 & ~n5702;
  assign n5704 = reg_i_StoB_REQ8_out & ~n5703;
  assign n5705 = reg_controllable_BtoS_ACK7_out & ~n5300;
  assign n5706 = ~n1812 & ~n5705;
  assign n5707 = reg_i_StoB_REQ7_out & ~n5706;
  assign n5708 = reg_controllable_BtoS_ACK6_out & ~n5284;
  assign n5709 = ~n1776 & ~n5708;
  assign n5710 = reg_i_StoB_REQ6_out & ~n5709;
  assign n5711 = reg_controllable_BtoS_ACK5_out & ~n5268;
  assign n5712 = ~n1740 & ~n5711;
  assign n5713 = reg_i_StoB_REQ5_out & ~n5712;
  assign n5714 = reg_controllable_BtoS_ACK4_out & ~n5249;
  assign n5715 = ~n1696 & ~n5714;
  assign n5716 = reg_i_StoB_REQ4_out & ~n5715;
  assign n5717 = reg_controllable_BtoS_ACK3_out & ~n5245;
  assign n5718 = ~n1667 & ~n5717;
  assign n5719 = reg_i_StoB_REQ3_out & ~n5718;
  assign n5720 = reg_controllable_BtoS_ACK2_out & ~n5226;
  assign n5721 = ~n1640 & ~n5720;
  assign n5722 = reg_i_StoB_REQ2_out & ~n5721;
  assign n5723 = reg_stateG12_out & ~n2336;
  assign n5724 = ~reg_stateG12_out & ~n1608;
  assign n5725 = ~n5723 & ~n5724;
  assign n5726 = sys_fair12done_out & ~n5725;
  assign n5727 = ~n1131 & ~n1614;
  assign n5728 = ~sys_fair12done_out & ~n5727;
  assign n5729 = ~n5726 & ~n5728;
  assign n5730 = sys_fair2done_out & ~n5729;
  assign n5731 = reg_stateG12_out & ~n2218;
  assign n5732 = ~n1614 & ~n5731;
  assign n5733 = ~sys_fair2done_out & ~n5732;
  assign n5734 = ~n5730 & ~n5733;
  assign n5735 = reg_controllable_BtoS_ACK2_out & ~n5734;
  assign n5736 = ~reg_stateG12_out & ~n1612;
  assign n5737 = ~n1131 & ~n5736;
  assign n5738 = sys_fair12done_out & ~n5737;
  assign n5739 = ~n5728 & ~n5738;
  assign n5740 = ~sys_fair2done_out & ~n5739;
  assign n5741 = ~n5730 & ~n5740;
  assign n5742 = ~reg_controllable_BtoS_ACK2_out & ~n5741;
  assign n5743 = ~n5735 & ~n5742;
  assign n5744 = ~reg_i_StoB_REQ2_out & ~n5743;
  assign n5745 = ~n5722 & ~n5744;
  assign n5746 = sys_fair3done_out & ~n5745;
  assign n5747 = reg_controllable_BtoS_ACK2_out & ~n5217;
  assign n5748 = ~n1671 & ~n5747;
  assign n5749 = reg_i_StoB_REQ2_out & ~n5748;
  assign n5750 = ~reg_i_StoB_REQ2_out & ~n5732;
  assign n5751 = ~n5749 & ~n5750;
  assign n5752 = ~sys_fair3done_out & ~n5751;
  assign n5753 = ~n5746 & ~n5752;
  assign n5754 = reg_controllable_BtoS_ACK3_out & ~n5753;
  assign n5755 = reg_controllable_BtoS_ACK2_out & ~n5224;
  assign n5756 = ~n1681 & ~n5755;
  assign n5757 = reg_i_StoB_REQ2_out & ~n5756;
  assign n5758 = sys_fair2done_out & ~n5739;
  assign n5759 = ~n5733 & ~n5758;
  assign n5760 = reg_controllable_BtoS_ACK2_out & ~n5759;
  assign n5761 = ~reg_controllable_BtoS_ACK2_out & ~n5739;
  assign n5762 = ~n5760 & ~n5761;
  assign n5763 = ~reg_i_StoB_REQ2_out & ~n5762;
  assign n5764 = ~n5757 & ~n5763;
  assign n5765 = ~sys_fair3done_out & ~n5764;
  assign n5766 = ~n5746 & ~n5765;
  assign n5767 = ~reg_controllable_BtoS_ACK3_out & ~n5766;
  assign n5768 = ~n5754 & ~n5767;
  assign n5769 = ~reg_i_StoB_REQ3_out & ~n5768;
  assign n5770 = ~n5719 & ~n5769;
  assign n5771 = ~reg_i_StoB_REQ4_out & ~n5770;
  assign n5772 = ~n5716 & ~n5771;
  assign n5773 = sys_fair4done_out & ~n5772;
  assign n5774 = reg_controllable_BtoS_ACK4_out & ~n5262;
  assign n5775 = ~n1713 & ~n5774;
  assign n5776 = reg_i_StoB_REQ4_out & ~n5775;
  assign n5777 = reg_controllable_BtoS_ACK3_out & ~n5233;
  assign n5778 = ~n1717 & ~n5777;
  assign n5779 = reg_i_StoB_REQ3_out & ~n5778;
  assign n5780 = ~reg_i_StoB_REQ3_out & ~n5751;
  assign n5781 = ~n5779 & ~n5780;
  assign n5782 = reg_controllable_BtoS_ACK4_out & ~n5781;
  assign n5783 = reg_controllable_BtoS_ACK3_out & ~n5243;
  assign n5784 = ~n1725 & ~n5783;
  assign n5785 = reg_i_StoB_REQ3_out & ~n5784;
  assign n5786 = sys_fair3done_out & ~n5764;
  assign n5787 = ~n5752 & ~n5786;
  assign n5788 = reg_controllable_BtoS_ACK3_out & ~n5787;
  assign n5789 = ~reg_controllable_BtoS_ACK3_out & ~n5764;
  assign n5790 = ~n5788 & ~n5789;
  assign n5791 = ~reg_i_StoB_REQ3_out & ~n5790;
  assign n5792 = ~n5785 & ~n5791;
  assign n5793 = ~reg_controllable_BtoS_ACK4_out & ~n5792;
  assign n5794 = ~n5782 & ~n5793;
  assign n5795 = ~reg_i_StoB_REQ4_out & ~n5794;
  assign n5796 = ~n5776 & ~n5795;
  assign n5797 = ~sys_fair4done_out & ~n5796;
  assign n5798 = ~n5773 & ~n5797;
  assign n5799 = ~reg_i_StoB_REQ5_out & ~n5798;
  assign n5800 = ~n5713 & ~n5799;
  assign n5801 = sys_fair5done_out & ~n5800;
  assign n5802 = reg_controllable_BtoS_ACK5_out & ~n5278;
  assign n5803 = ~n1755 & ~n5802;
  assign n5804 = reg_i_StoB_REQ5_out & ~n5803;
  assign n5805 = ~n1758 & ~n5255;
  assign n5806 = reg_i_StoB_REQ4_out & ~n5805;
  assign n5807 = ~reg_i_StoB_REQ4_out & ~n5781;
  assign n5808 = ~n5806 & ~n5807;
  assign n5809 = reg_controllable_BtoS_ACK5_out & ~n5808;
  assign n5810 = ~n1734 & ~n5774;
  assign n5811 = reg_i_StoB_REQ4_out & ~n5810;
  assign n5812 = ~reg_i_StoB_REQ4_out & ~n5792;
  assign n5813 = ~n5811 & ~n5812;
  assign n5814 = sys_fair4done_out & ~n5813;
  assign n5815 = ~n5797 & ~n5814;
  assign n5816 = ~reg_controllable_BtoS_ACK5_out & ~n5815;
  assign n5817 = ~n5809 & ~n5816;
  assign n5818 = ~reg_i_StoB_REQ5_out & ~n5817;
  assign n5819 = ~n5804 & ~n5818;
  assign n5820 = ~sys_fair5done_out & ~n5819;
  assign n5821 = ~n5801 & ~n5820;
  assign n5822 = ~reg_i_StoB_REQ6_out & ~n5821;
  assign n5823 = ~n5710 & ~n5822;
  assign n5824 = sys_fair6done_out & ~n5823;
  assign n5825 = reg_controllable_BtoS_ACK6_out & ~n5294;
  assign n5826 = ~n1791 & ~n5825;
  assign n5827 = reg_i_StoB_REQ6_out & ~n5826;
  assign n5828 = ~n1794 & ~n5274;
  assign n5829 = reg_i_StoB_REQ5_out & ~n5828;
  assign n5830 = ~reg_i_StoB_REQ5_out & ~n5808;
  assign n5831 = ~n5829 & ~n5830;
  assign n5832 = reg_controllable_BtoS_ACK6_out & ~n5831;
  assign n5833 = ~n1770 & ~n5802;
  assign n5834 = reg_i_StoB_REQ5_out & ~n5833;
  assign n5835 = ~reg_i_StoB_REQ5_out & ~n5815;
  assign n5836 = ~n5834 & ~n5835;
  assign n5837 = sys_fair5done_out & ~n5836;
  assign n5838 = ~n5820 & ~n5837;
  assign n5839 = ~reg_controllable_BtoS_ACK6_out & ~n5838;
  assign n5840 = ~n5832 & ~n5839;
  assign n5841 = ~reg_i_StoB_REQ6_out & ~n5840;
  assign n5842 = ~n5827 & ~n5841;
  assign n5843 = ~sys_fair6done_out & ~n5842;
  assign n5844 = ~n5824 & ~n5843;
  assign n5845 = ~reg_i_StoB_REQ7_out & ~n5844;
  assign n5846 = ~n5707 & ~n5845;
  assign n5847 = sys_fair7done_out & ~n5846;
  assign n5848 = reg_controllable_BtoS_ACK7_out & ~n5310;
  assign n5849 = ~n1827 & ~n5848;
  assign n5850 = reg_i_StoB_REQ7_out & ~n5849;
  assign n5851 = ~n1830 & ~n5290;
  assign n5852 = reg_i_StoB_REQ6_out & ~n5851;
  assign n5853 = ~reg_i_StoB_REQ6_out & ~n5831;
  assign n5854 = ~n5852 & ~n5853;
  assign n5855 = reg_controllable_BtoS_ACK7_out & ~n5854;
  assign n5856 = ~n1806 & ~n5825;
  assign n5857 = reg_i_StoB_REQ6_out & ~n5856;
  assign n5858 = ~reg_i_StoB_REQ6_out & ~n5838;
  assign n5859 = ~n5857 & ~n5858;
  assign n5860 = sys_fair6done_out & ~n5859;
  assign n5861 = ~n5843 & ~n5860;
  assign n5862 = ~reg_controllable_BtoS_ACK7_out & ~n5861;
  assign n5863 = ~n5855 & ~n5862;
  assign n5864 = ~reg_i_StoB_REQ7_out & ~n5863;
  assign n5865 = ~n5850 & ~n5864;
  assign n5866 = ~sys_fair7done_out & ~n5865;
  assign n5867 = ~n5847 & ~n5866;
  assign n5868 = sys_fair8done_out & ~n5867;
  assign n5869 = ~n1862 & ~n5306;
  assign n5870 = reg_i_StoB_REQ7_out & ~n5869;
  assign n5871 = ~reg_i_StoB_REQ7_out & ~n5854;
  assign n5872 = ~n5870 & ~n5871;
  assign n5873 = ~sys_fair8done_out & ~n5872;
  assign n5874 = ~n5868 & ~n5873;
  assign n5875 = reg_controllable_BtoS_ACK8_out & ~n5874;
  assign n5876 = ~n1842 & ~n5848;
  assign n5877 = reg_i_StoB_REQ7_out & ~n5876;
  assign n5878 = ~reg_i_StoB_REQ7_out & ~n5861;
  assign n5879 = ~n5877 & ~n5878;
  assign n5880 = sys_fair7done_out & ~n5879;
  assign n5881 = ~n5866 & ~n5880;
  assign n5882 = ~sys_fair8done_out & ~n5881;
  assign n5883 = ~n5868 & ~n5882;
  assign n5884 = ~reg_controllable_BtoS_ACK8_out & ~n5883;
  assign n5885 = ~n5875 & ~n5884;
  assign n5886 = ~reg_i_StoB_REQ8_out & ~n5885;
  assign n5887 = ~n5704 & ~n5886;
  assign n5888 = ~reg_i_StoB_REQ10_out & ~n5887;
  assign n5889 = ~n5701 & ~n5888;
  assign n5890 = sys_fair10done_out & ~n5889;
  assign n5891 = reg_controllable_BtoS_ACK10_out & ~n5345;
  assign n5892 = ~n1899 & ~n5891;
  assign n5893 = reg_i_StoB_REQ10_out & ~n5892;
  assign n5894 = reg_controllable_BtoS_ACK8_out & ~n5319;
  assign n5895 = ~n1903 & ~n5894;
  assign n5896 = reg_i_StoB_REQ8_out & ~n5895;
  assign n5897 = ~reg_i_StoB_REQ8_out & ~n5872;
  assign n5898 = ~n5896 & ~n5897;
  assign n5899 = reg_controllable_BtoS_ACK10_out & ~n5898;
  assign n5900 = reg_controllable_BtoS_ACK8_out & ~n5326;
  assign n5901 = ~n1911 & ~n5900;
  assign n5902 = reg_i_StoB_REQ8_out & ~n5901;
  assign n5903 = sys_fair8done_out & ~n5881;
  assign n5904 = ~n5873 & ~n5903;
  assign n5905 = reg_controllable_BtoS_ACK8_out & ~n5904;
  assign n5906 = ~reg_controllable_BtoS_ACK8_out & ~n5881;
  assign n5907 = ~n5905 & ~n5906;
  assign n5908 = ~reg_i_StoB_REQ8_out & ~n5907;
  assign n5909 = ~n5902 & ~n5908;
  assign n5910 = ~reg_controllable_BtoS_ACK10_out & ~n5909;
  assign n5911 = ~n5899 & ~n5910;
  assign n5912 = ~reg_i_StoB_REQ10_out & ~n5911;
  assign n5913 = ~n5893 & ~n5912;
  assign n5914 = ~sys_fair10done_out & ~n5913;
  assign n5915 = ~n5890 & ~n5914;
  assign n5916 = sys_fair11done_out & ~n5915;
  assign n5917 = ~n1940 & ~n5338;
  assign n5918 = reg_i_StoB_REQ10_out & ~n5917;
  assign n5919 = ~reg_i_StoB_REQ10_out & ~n5898;
  assign n5920 = ~n5918 & ~n5919;
  assign n5921 = ~sys_fair11done_out & ~n5920;
  assign n5922 = ~n5916 & ~n5921;
  assign n5923 = reg_controllable_BtoS_ACK11_out & ~n5922;
  assign n5924 = ~n1920 & ~n5891;
  assign n5925 = reg_i_StoB_REQ10_out & ~n5924;
  assign n5926 = ~reg_i_StoB_REQ10_out & ~n5909;
  assign n5927 = ~n5925 & ~n5926;
  assign n5928 = sys_fair10done_out & ~n5927;
  assign n5929 = ~n5914 & ~n5928;
  assign n5930 = ~sys_fair11done_out & ~n5929;
  assign n5931 = ~n5916 & ~n5930;
  assign n5932 = ~reg_controllable_BtoS_ACK11_out & ~n5931;
  assign n5933 = ~n5923 & ~n5932;
  assign n5934 = ~reg_i_StoB_REQ11_out & ~n5933;
  assign n5935 = ~n5698 & ~n5934;
  assign n5936 = sys_fair9done_out & ~n5935;
  assign n5937 = reg_controllable_BtoS_ACK11_out & ~n5354;
  assign n5938 = ~n1962 & ~n5937;
  assign n5939 = reg_i_StoB_REQ11_out & ~n5938;
  assign n5940 = ~reg_i_StoB_REQ11_out & ~n5920;
  assign n5941 = ~n5939 & ~n5940;
  assign n5942 = ~sys_fair9done_out & ~n5941;
  assign n5943 = ~n5936 & ~n5942;
  assign n5944 = fair_cnt<1>_out  & ~n5943;
  assign n5945 = reg_controllable_BtoS_ACK11_out & ~n5421;
  assign n5946 = ~n4182 & ~n5945;
  assign n5947 = reg_i_StoB_REQ11_out & ~n5946;
  assign n5948 = reg_controllable_BtoS_ACK10_out & ~n5414;
  assign n5949 = ~n4173 & ~n5948;
  assign n5950 = reg_i_StoB_REQ10_out & ~n5949;
  assign n5951 = reg_controllable_BtoS_ACK8_out & ~n5412;
  assign n5952 = ~n4168 & ~n5951;
  assign n5953 = reg_i_StoB_REQ8_out & ~n5952;
  assign n5954 = reg_controllable_BtoS_ACK7_out & ~n5405;
  assign n5955 = ~n4159 & ~n5954;
  assign n5956 = reg_i_StoB_REQ7_out & ~n5955;
  assign n5957 = reg_controllable_BtoS_ACK6_out & ~n5400;
  assign n5958 = ~n4152 & ~n5957;
  assign n5959 = reg_i_StoB_REQ6_out & ~n5958;
  assign n5960 = reg_controllable_BtoS_ACK5_out & ~n5395;
  assign n5961 = ~n4145 & ~n5960;
  assign n5962 = reg_i_StoB_REQ5_out & ~n5961;
  assign n5963 = reg_controllable_BtoS_ACK4_out & ~n5390;
  assign n5964 = ~n4138 & ~n5963;
  assign n5965 = reg_i_StoB_REQ4_out & ~n5964;
  assign n5966 = reg_controllable_BtoS_ACK3_out & ~n5388;
  assign n5967 = ~n4133 & ~n5966;
  assign n5968 = reg_i_StoB_REQ3_out & ~n5967;
  assign n5969 = reg_controllable_BtoS_ACK2_out & ~n5384;
  assign n5970 = ~n4126 & ~n5969;
  assign n5971 = reg_i_StoB_REQ2_out & ~n5970;
  assign n5972 = sys_fair12done_out & ~n5732;
  assign n5973 = ~n1614 & ~n4307;
  assign n5974 = ~sys_fair12done_out & ~n5973;
  assign n5975 = ~n5972 & ~n5974;
  assign n5976 = sys_fair2done_out & ~n5975;
  assign n5977 = ~n5733 & ~n5976;
  assign n5978 = ~reg_i_StoB_REQ2_out & ~n5977;
  assign n5979 = ~n5971 & ~n5978;
  assign n5980 = sys_fair3done_out & ~n5979;
  assign n5981 = ~n5752 & ~n5980;
  assign n5982 = ~reg_i_StoB_REQ3_out & ~n5981;
  assign n5983 = ~n5968 & ~n5982;
  assign n5984 = ~reg_i_StoB_REQ4_out & ~n5983;
  assign n5985 = ~n5965 & ~n5984;
  assign n5986 = sys_fair4done_out & ~n5985;
  assign n5987 = ~sys_fair4done_out & ~n5808;
  assign n5988 = ~n5986 & ~n5987;
  assign n5989 = ~reg_i_StoB_REQ5_out & ~n5988;
  assign n5990 = ~n5962 & ~n5989;
  assign n5991 = sys_fair5done_out & ~n5990;
  assign n5992 = ~sys_fair5done_out & ~n5831;
  assign n5993 = ~n5991 & ~n5992;
  assign n5994 = ~reg_i_StoB_REQ6_out & ~n5993;
  assign n5995 = ~n5959 & ~n5994;
  assign n5996 = sys_fair6done_out & ~n5995;
  assign n5997 = ~sys_fair6done_out & ~n5854;
  assign n5998 = ~n5996 & ~n5997;
  assign n5999 = ~reg_i_StoB_REQ7_out & ~n5998;
  assign n6000 = ~n5956 & ~n5999;
  assign n6001 = sys_fair7done_out & ~n6000;
  assign n6002 = ~sys_fair7done_out & ~n5872;
  assign n6003 = ~n6001 & ~n6002;
  assign n6004 = sys_fair8done_out & ~n6003;
  assign n6005 = ~n5873 & ~n6004;
  assign n6006 = ~reg_i_StoB_REQ8_out & ~n6005;
  assign n6007 = ~n5953 & ~n6006;
  assign n6008 = ~reg_i_StoB_REQ10_out & ~n6007;
  assign n6009 = ~n5950 & ~n6008;
  assign n6010 = sys_fair10done_out & ~n6009;
  assign n6011 = ~sys_fair10done_out & ~n5920;
  assign n6012 = ~n6010 & ~n6011;
  assign n6013 = sys_fair11done_out & ~n6012;
  assign n6014 = ~n5921 & ~n6013;
  assign n6015 = ~reg_i_StoB_REQ11_out & ~n6014;
  assign n6016 = ~n5947 & ~n6015;
  assign n6017 = sys_fair9done_out & ~n6016;
  assign n6018 = ~n5942 & ~n6017;
  assign n6019 = ~fair_cnt<1>_out  & ~n6018;
  assign n6020 = ~n5944 & ~n6019;
  assign n6021 = fair_cnt<0>_out  & ~n6020;
  assign n6022 = fair_cnt<1>_out  & ~n6018;
  assign n6023 = reg_controllable_BtoS_ACK11_out & ~n5469;
  assign n6024 = ~n5589 & ~n6023;
  assign n6025 = reg_i_StoB_REQ11_out & ~n6024;
  assign n6026 = reg_controllable_BtoS_ACK10_out & ~n5463;
  assign n6027 = ~n5593 & ~n6026;
  assign n6028 = reg_i_StoB_REQ10_out & ~n6027;
  assign n6029 = reg_controllable_BtoS_ACK8_out & ~n5461;
  assign n6030 = ~n5597 & ~n6029;
  assign n6031 = reg_i_StoB_REQ8_out & ~n6030;
  assign n6032 = reg_controllable_BtoS_ACK7_out & ~n5455;
  assign n6033 = ~n5601 & ~n6032;
  assign n6034 = reg_i_StoB_REQ7_out & ~n6033;
  assign n6035 = reg_controllable_BtoS_ACK6_out & ~n5451;
  assign n6036 = ~n5605 & ~n6035;
  assign n6037 = reg_i_StoB_REQ6_out & ~n6036;
  assign n6038 = reg_controllable_BtoS_ACK5_out & ~n5447;
  assign n6039 = ~n5609 & ~n6038;
  assign n6040 = reg_i_StoB_REQ5_out & ~n6039;
  assign n6041 = reg_controllable_BtoS_ACK4_out & ~n5443;
  assign n6042 = ~n5613 & ~n6041;
  assign n6043 = reg_i_StoB_REQ4_out & ~n6042;
  assign n6044 = reg_controllable_BtoS_ACK3_out & ~n5441;
  assign n6045 = ~n5617 & ~n6044;
  assign n6046 = reg_i_StoB_REQ3_out & ~n6045;
  assign n6047 = reg_controllable_BtoS_ACK2_out & ~n5437;
  assign n6048 = ~n5621 & ~n6047;
  assign n6049 = reg_i_StoB_REQ2_out & ~n6048;
  assign n6050 = ~n1614 & ~n5627;
  assign n6051 = ~sys_fair12done_out & ~n6050;
  assign n6052 = ~n5972 & ~n6051;
  assign n6053 = sys_fair2done_out & ~n6052;
  assign n6054 = ~n5733 & ~n6053;
  assign n6055 = ~reg_i_StoB_REQ2_out & ~n6054;
  assign n6056 = ~n6049 & ~n6055;
  assign n6057 = sys_fair3done_out & ~n6056;
  assign n6058 = ~n5752 & ~n6057;
  assign n6059 = ~reg_i_StoB_REQ3_out & ~n6058;
  assign n6060 = ~n6046 & ~n6059;
  assign n6061 = ~reg_i_StoB_REQ4_out & ~n6060;
  assign n6062 = ~n6043 & ~n6061;
  assign n6063 = sys_fair4done_out & ~n6062;
  assign n6064 = ~n5987 & ~n6063;
  assign n6065 = ~reg_i_StoB_REQ5_out & ~n6064;
  assign n6066 = ~n6040 & ~n6065;
  assign n6067 = sys_fair5done_out & ~n6066;
  assign n6068 = ~n5992 & ~n6067;
  assign n6069 = ~reg_i_StoB_REQ6_out & ~n6068;
  assign n6070 = ~n6037 & ~n6069;
  assign n6071 = sys_fair6done_out & ~n6070;
  assign n6072 = ~n5997 & ~n6071;
  assign n6073 = ~reg_i_StoB_REQ7_out & ~n6072;
  assign n6074 = ~n6034 & ~n6073;
  assign n6075 = sys_fair7done_out & ~n6074;
  assign n6076 = ~n6002 & ~n6075;
  assign n6077 = sys_fair8done_out & ~n6076;
  assign n6078 = ~n5873 & ~n6077;
  assign n6079 = ~reg_i_StoB_REQ8_out & ~n6078;
  assign n6080 = ~n6031 & ~n6079;
  assign n6081 = ~reg_i_StoB_REQ10_out & ~n6080;
  assign n6082 = ~n6028 & ~n6081;
  assign n6083 = sys_fair10done_out & ~n6082;
  assign n6084 = ~n6011 & ~n6083;
  assign n6085 = sys_fair11done_out & ~n6084;
  assign n6086 = ~n5921 & ~n6085;
  assign n6087 = ~reg_i_StoB_REQ11_out & ~n6086;
  assign n6088 = ~n6025 & ~n6087;
  assign n6089 = sys_fair9done_out & ~n6088;
  assign n6090 = ~n5942 & ~n6089;
  assign n6091 = ~fair_cnt<1>_out  & ~n6090;
  assign n6092 = ~n6022 & ~n6091;
  assign n6093 = ~fair_cnt<0>_out  & ~n6092;
  assign n6094 = ~n6021 & ~n6093;
  assign n6095 = env_fair1done_out & ~n6094;
  assign n6096 = ~sys_fair11done_out & ~n5515;
  assign n6097 = ~n5420 & ~n6096;
  assign n6098 = reg_controllable_BtoS_ACK11_out & ~n6097;
  assign n6099 = ~n4182 & ~n6098;
  assign n6100 = reg_i_StoB_REQ11_out & ~n6099;
  assign n6101 = ~sys_fair8done_out & ~n5507;
  assign n6102 = ~n5411 & ~n6101;
  assign n6103 = reg_controllable_BtoS_ACK8_out & ~n6102;
  assign n6104 = ~n4168 & ~n6103;
  assign n6105 = reg_i_StoB_REQ8_out & ~n6104;
  assign n6106 = ~sys_fair3done_out & ~n5487;
  assign n6107 = ~n5387 & ~n6106;
  assign n6108 = reg_controllable_BtoS_ACK3_out & ~n6107;
  assign n6109 = ~n4133 & ~n6108;
  assign n6110 = reg_i_StoB_REQ3_out & ~n6109;
  assign n6111 = ~sys_fair2done_out & ~n5483;
  assign n6112 = ~n5383 & ~n6111;
  assign n6113 = reg_controllable_BtoS_ACK2_out & ~n6112;
  assign n6114 = ~n4126 & ~n6113;
  assign n6115 = reg_i_StoB_REQ2_out & ~n6114;
  assign n6116 = ~reg_stateG12_out & ~n2216;
  assign n6117 = ~n5731 & ~n6116;
  assign n6118 = sys_fair12done_out & ~n6117;
  assign n6119 = ~n5974 & ~n6118;
  assign n6120 = sys_fair2done_out & ~n6119;
  assign n6121 = ~n5733 & ~n6120;
  assign n6122 = ~reg_i_StoB_REQ2_out & ~n6121;
  assign n6123 = ~n6115 & ~n6122;
  assign n6124 = sys_fair3done_out & ~n6123;
  assign n6125 = ~n5752 & ~n6124;
  assign n6126 = ~reg_i_StoB_REQ3_out & ~n6125;
  assign n6127 = ~n6110 & ~n6126;
  assign n6128 = ~reg_i_StoB_REQ4_out & ~n6127;
  assign n6129 = ~n5965 & ~n6128;
  assign n6130 = sys_fair4done_out & ~n6129;
  assign n6131 = reg_controllable_BtoS_ACK4_out & ~n5491;
  assign n6132 = ~n1758 & ~n6131;
  assign n6133 = reg_i_StoB_REQ4_out & ~n6132;
  assign n6134 = ~n5807 & ~n6133;
  assign n6135 = ~sys_fair4done_out & ~n6134;
  assign n6136 = ~n6130 & ~n6135;
  assign n6137 = ~reg_i_StoB_REQ5_out & ~n6136;
  assign n6138 = ~n5962 & ~n6137;
  assign n6139 = sys_fair5done_out & ~n6138;
  assign n6140 = reg_controllable_BtoS_ACK5_out & ~n5495;
  assign n6141 = ~n1794 & ~n6140;
  assign n6142 = reg_i_StoB_REQ5_out & ~n6141;
  assign n6143 = ~n5830 & ~n6142;
  assign n6144 = ~sys_fair5done_out & ~n6143;
  assign n6145 = ~n6139 & ~n6144;
  assign n6146 = ~reg_i_StoB_REQ6_out & ~n6145;
  assign n6147 = ~n5959 & ~n6146;
  assign n6148 = sys_fair6done_out & ~n6147;
  assign n6149 = reg_controllable_BtoS_ACK6_out & ~n5499;
  assign n6150 = ~n1830 & ~n6149;
  assign n6151 = reg_i_StoB_REQ6_out & ~n6150;
  assign n6152 = ~n5853 & ~n6151;
  assign n6153 = ~sys_fair6done_out & ~n6152;
  assign n6154 = ~n6148 & ~n6153;
  assign n6155 = ~reg_i_StoB_REQ7_out & ~n6154;
  assign n6156 = ~n5956 & ~n6155;
  assign n6157 = sys_fair7done_out & ~n6156;
  assign n6158 = reg_controllable_BtoS_ACK7_out & ~n5503;
  assign n6159 = ~n1862 & ~n6158;
  assign n6160 = reg_i_StoB_REQ7_out & ~n6159;
  assign n6161 = ~n5871 & ~n6160;
  assign n6162 = ~sys_fair7done_out & ~n6161;
  assign n6163 = ~n6157 & ~n6162;
  assign n6164 = sys_fair8done_out & ~n6163;
  assign n6165 = ~n5873 & ~n6164;
  assign n6166 = ~reg_i_StoB_REQ8_out & ~n6165;
  assign n6167 = ~n6105 & ~n6166;
  assign n6168 = ~reg_i_StoB_REQ10_out & ~n6167;
  assign n6169 = ~n5950 & ~n6168;
  assign n6170 = sys_fair10done_out & ~n6169;
  assign n6171 = reg_controllable_BtoS_ACK10_out & ~n5511;
  assign n6172 = ~n1940 & ~n6171;
  assign n6173 = reg_i_StoB_REQ10_out & ~n6172;
  assign n6174 = ~n5919 & ~n6173;
  assign n6175 = ~sys_fair10done_out & ~n6174;
  assign n6176 = ~n6170 & ~n6175;
  assign n6177 = sys_fair11done_out & ~n6176;
  assign n6178 = ~n5921 & ~n6177;
  assign n6179 = ~reg_i_StoB_REQ11_out & ~n6178;
  assign n6180 = ~n6100 & ~n6179;
  assign n6181 = sys_fair9done_out & ~n6180;
  assign n6182 = ~n5942 & ~n6181;
  assign n6183 = fair_cnt<1>_out  & ~n6182;
  assign n6184 = ~n6091 & ~n6183;
  assign n6185 = fair_cnt<0>_out  & ~n6184;
  assign n6186 = ~fair_cnt<1>_out  & ~n5941;
  assign n6187 = ~n6022 & ~n6186;
  assign n6188 = ~fair_cnt<0>_out  & ~n6187;
  assign n6189 = ~n6185 & ~n6188;
  assign n6190 = ~env_fair1done_out & ~n6189;
  assign n6191 = ~n6095 & ~n6190;
  assign n6192 = reg_nstateG7_1_out & ~n6191;
  assign n6193 = env_fair0done_out & ~n6094;
  assign n6194 = ~env_fair0done_out & ~n6189;
  assign n6195 = ~n6193 & ~n6194;
  assign n6196 = ~reg_nstateG7_1_out & ~n6195;
  assign n6197 = ~n6192 & ~n6196;
  assign n6198 = ~reg_controllable_BtoR_REQ1_out & ~n6197;
  assign n6199 = ~n5695 & ~n6198;
  assign n6200 = ~reg_controllable_BtoR_REQ0_out & ~n6199;
  assign n6201 = ~n5686 & ~n6200;
  assign n6202 = ~reg_i_RtoB_ACK1_out & ~n6201;
  assign n6203 = ~n5584 & ~n6202;
  assign n6204 = ~reg_i_RtoB_ACK0_out & ~n6203;
  assign n6205 = ~n5567 & ~n6204;
  assign n6206 = ~reg_i_StoB_REQ9_out & ~n6205;
  assign n6207 = ~n5545 & ~n6206;
  assign n6208 = reg_controllable_BtoS_ACK9_out & ~n6207;
  assign n6209 = ~n2874 & ~n3681;
  assign n6210 = fair_cnt<0>_out  & ~n6209;
  assign n6211 = ~n3758 & ~n6210;
  assign n6212 = env_fair1done_out & ~n6211;
  assign n6213 = ~n3674 & ~n6210;
  assign n6214 = ~env_fair1done_out & ~n6213;
  assign n6215 = ~n6212 & ~n6214;
  assign n6216 = env_fair0done_out & ~n6215;
  assign n6217 = ~env_fair0done_out & ~n4643;
  assign n6218 = ~n6216 & ~n6217;
  assign n6219 = ~reg_stateG7_0_out & ~n6218;
  assign n6220 = ~reg_stateG7_0_out & ~n6219;
  assign n6221 = reg_nstateG7_1_out & ~n6220;
  assign n6222 = ~reg_nstateG7_1_out & ~n6218;
  assign n6223 = ~n6221 & ~n6222;
  assign n6224 = ~reg_controllable_BtoR_REQ1_out & ~n6223;
  assign n6225 = ~reg_controllable_BtoR_REQ1_out & ~n6224;
  assign n6226 = reg_controllable_BtoR_REQ0_out & ~n6225;
  assign n6227 = reg_controllable_BtoR_REQ0_out & ~n6226;
  assign n6228 = ~reg_i_RtoB_ACK1_out & ~n6227;
  assign n6229 = ~reg_i_RtoB_ACK1_out & ~n6228;
  assign n6230 = reg_i_RtoB_ACK0_out & ~n6229;
  assign n6231 = ~env_fair1done_out & ~n4643;
  assign n6232 = ~n6212 & ~n6231;
  assign n6233 = env_fair0done_out & ~n6232;
  assign n6234 = env_fair1done_out & ~n6213;
  assign n6235 = ~n6231 & ~n6234;
  assign n6236 = ~env_fair0done_out & ~n6235;
  assign n6237 = ~n6233 & ~n6236;
  assign n6238 = reg_nstateG7_1_out & ~n6237;
  assign n6239 = ~reg_stateG7_0_out & ~n6237;
  assign n6240 = ~reg_stateG7_0_out & ~n6239;
  assign n6241 = ~reg_nstateG7_1_out & ~n6240;
  assign n6242 = ~n6238 & ~n6241;
  assign n6243 = reg_controllable_BtoR_REQ1_out & ~n6242;
  assign n6244 = reg_controllable_BtoR_REQ1_out & ~n6243;
  assign n6245 = ~reg_controllable_BtoR_REQ0_out & ~n6244;
  assign n6246 = ~reg_controllable_BtoR_REQ0_out & ~n6245;
  assign n6247 = reg_i_RtoB_ACK1_out & ~n6246;
  assign n6248 = ~n5001 & ~n5067;
  assign n6249 = env_fair0done_out & ~n6248;
  assign n6250 = ~n2927 & ~n4105;
  assign n6251 = fair_cnt<0>_out  & ~n6250;
  assign n6252 = ~n4191 & ~n6251;
  assign n6253 = ~env_fair0done_out & ~n6252;
  assign n6254 = ~n6249 & ~n6253;
  assign n6255 = ~reg_stateG7_0_out & ~n6254;
  assign n6256 = ~reg_stateG7_0_out & ~n6255;
  assign n6257 = reg_nstateG7_1_out & ~n6256;
  assign n6258 = ~reg_nstateG7_1_out & ~n6254;
  assign n6259 = ~n6257 & ~n6258;
  assign n6260 = ~reg_controllable_BtoR_REQ1_out & ~n6259;
  assign n6261 = ~reg_controllable_BtoR_REQ1_out & ~n6260;
  assign n6262 = reg_controllable_BtoR_REQ0_out & ~n6261;
  assign n6263 = env_fair1done_out & ~n6248;
  assign n6264 = ~env_fair1done_out & ~n6252;
  assign n6265 = ~n6263 & ~n6264;
  assign n6266 = reg_nstateG7_1_out & ~n6265;
  assign n6267 = ~reg_stateG7_0_out & ~n6265;
  assign n6268 = ~reg_stateG7_0_out & ~n6267;
  assign n6269 = ~reg_nstateG7_1_out & ~n6268;
  assign n6270 = ~n6266 & ~n6269;
  assign n6271 = reg_controllable_BtoR_REQ1_out & ~n6270;
  assign n6272 = ~n5025 & ~n6263;
  assign n6273 = reg_nstateG7_1_out & ~n6272;
  assign n6274 = ~n5028 & ~n6249;
  assign n6275 = ~reg_nstateG7_1_out & ~n6274;
  assign n6276 = ~n6273 & ~n6275;
  assign n6277 = ~reg_controllable_BtoR_REQ1_out & ~n6276;
  assign n6278 = ~n6271 & ~n6277;
  assign n6279 = ~reg_controllable_BtoR_REQ0_out & ~n6278;
  assign n6280 = ~n6262 & ~n6279;
  assign n6281 = ~reg_i_RtoB_ACK1_out & ~n6280;
  assign n6282 = ~n6247 & ~n6281;
  assign n6283 = ~reg_i_RtoB_ACK0_out & ~n6282;
  assign n6284 = ~n6230 & ~n6283;
  assign n6285 = reg_i_StoB_REQ9_out & ~n6284;
  assign n6286 = ~n3069 & ~n5181;
  assign n6287 = fair_cnt<0>_out  & ~n6286;
  assign n6288 = ~n3834 & ~n6287;
  assign n6289 = env_fair1done_out & ~n6288;
  assign n6290 = ~n4010 & ~n6287;
  assign n6291 = ~env_fair1done_out & ~n6290;
  assign n6292 = ~n6289 & ~n6291;
  assign n6293 = env_fair0done_out & ~n6292;
  assign n6294 = ~env_fair0done_out & ~n4782;
  assign n6295 = ~n6293 & ~n6294;
  assign n6296 = ~reg_stateG7_0_out & ~n6295;
  assign n6297 = ~reg_stateG7_0_out & ~n6296;
  assign n6298 = reg_nstateG7_1_out & ~n6297;
  assign n6299 = ~reg_nstateG7_1_out & ~n6295;
  assign n6300 = ~n6298 & ~n6299;
  assign n6301 = ~reg_controllable_BtoR_REQ1_out & ~n6300;
  assign n6302 = ~reg_controllable_BtoR_REQ1_out & ~n6301;
  assign n6303 = reg_controllable_BtoR_REQ0_out & ~n6302;
  assign n6304 = reg_controllable_BtoR_REQ0_out & ~n6303;
  assign n6305 = ~reg_i_RtoB_ACK1_out & ~n6304;
  assign n6306 = ~reg_i_RtoB_ACK1_out & ~n6305;
  assign n6307 = reg_i_RtoB_ACK0_out & ~n6306;
  assign n6308 = ~env_fair1done_out & ~n4782;
  assign n6309 = ~n6289 & ~n6308;
  assign n6310 = env_fair0done_out & ~n6309;
  assign n6311 = env_fair1done_out & ~n6290;
  assign n6312 = ~n6308 & ~n6311;
  assign n6313 = ~env_fair0done_out & ~n6312;
  assign n6314 = ~n6310 & ~n6313;
  assign n6315 = reg_nstateG7_1_out & ~n6314;
  assign n6316 = ~reg_stateG7_0_out & ~n6314;
  assign n6317 = ~reg_stateG7_0_out & ~n6316;
  assign n6318 = ~reg_nstateG7_1_out & ~n6317;
  assign n6319 = ~n6315 & ~n6318;
  assign n6320 = reg_controllable_BtoR_REQ1_out & ~n6319;
  assign n6321 = reg_controllable_BtoR_REQ1_out & ~n6320;
  assign n6322 = ~reg_controllable_BtoR_REQ0_out & ~n6321;
  assign n6323 = ~reg_controllable_BtoR_REQ0_out & ~n6322;
  assign n6324 = reg_i_RtoB_ACK1_out & ~n6323;
  assign n6325 = ~n3156 & ~n5585;
  assign n6326 = fair_cnt<0>_out  & ~n6325;
  assign n6327 = ~n5671 & ~n6326;
  assign n6328 = env_fair0done_out & ~n6327;
  assign n6329 = ~n3156 & ~n5669;
  assign n6330 = fair_cnt<0>_out  & ~n6329;
  assign n6331 = ~n4356 & ~n6330;
  assign n6332 = ~env_fair0done_out & ~n6331;
  assign n6333 = ~n6328 & ~n6332;
  assign n6334 = ~reg_stateG7_0_out & ~n6333;
  assign n6335 = ~reg_stateG7_0_out & ~n6334;
  assign n6336 = reg_nstateG7_1_out & ~n6335;
  assign n6337 = ~reg_nstateG7_1_out & ~n6333;
  assign n6338 = ~n6336 & ~n6337;
  assign n6339 = ~reg_controllable_BtoR_REQ1_out & ~n6338;
  assign n6340 = ~reg_controllable_BtoR_REQ1_out & ~n6339;
  assign n6341 = reg_controllable_BtoR_REQ0_out & ~n6340;
  assign n6342 = env_fair1done_out & ~n6327;
  assign n6343 = ~env_fair1done_out & ~n6331;
  assign n6344 = ~n6342 & ~n6343;
  assign n6345 = reg_nstateG7_1_out & ~n6344;
  assign n6346 = ~reg_stateG7_0_out & ~n6344;
  assign n6347 = ~reg_stateG7_0_out & ~n6346;
  assign n6348 = ~reg_nstateG7_1_out & ~n6347;
  assign n6349 = ~n6345 & ~n6348;
  assign n6350 = reg_controllable_BtoR_REQ1_out & ~n6349;
  assign n6351 = reg_controllable_BtoS_ACK11_out & ~n5361;
  assign n6352 = ~n3113 & ~n6351;
  assign n6353 = reg_i_StoB_REQ11_out & ~n6352;
  assign n6354 = sys_fair11done_out & ~n5929;
  assign n6355 = ~n5921 & ~n6354;
  assign n6356 = reg_controllable_BtoS_ACK11_out & ~n6355;
  assign n6357 = ~reg_controllable_BtoS_ACK11_out & ~n5929;
  assign n6358 = ~n6356 & ~n6357;
  assign n6359 = ~reg_i_StoB_REQ11_out & ~n6358;
  assign n6360 = ~n6353 & ~n6359;
  assign n6361 = ~sys_fair9done_out & ~n6360;
  assign n6362 = ~n5936 & ~n6361;
  assign n6363 = fair_cnt<1>_out  & ~n6362;
  assign n6364 = ~n6019 & ~n6363;
  assign n6365 = fair_cnt<0>_out  & ~n6364;
  assign n6366 = ~n6093 & ~n6365;
  assign n6367 = env_fair1done_out & ~n6366;
  assign n6368 = ~n6190 & ~n6367;
  assign n6369 = reg_nstateG7_1_out & ~n6368;
  assign n6370 = env_fair0done_out & ~n6366;
  assign n6371 = ~n6194 & ~n6370;
  assign n6372 = ~reg_nstateG7_1_out & ~n6371;
  assign n6373 = ~n6369 & ~n6372;
  assign n6374 = ~reg_controllable_BtoR_REQ1_out & ~n6373;
  assign n6375 = ~n6350 & ~n6374;
  assign n6376 = ~reg_controllable_BtoR_REQ0_out & ~n6375;
  assign n6377 = ~n6341 & ~n6376;
  assign n6378 = ~reg_i_RtoB_ACK1_out & ~n6377;
  assign n6379 = ~n6324 & ~n6378;
  assign n6380 = ~reg_i_RtoB_ACK0_out & ~n6379;
  assign n6381 = ~n6307 & ~n6380;
  assign n6382 = ~reg_i_StoB_REQ9_out & ~n6381;
  assign n6383 = ~n6285 & ~n6382;
  assign n6384 = ~reg_controllable_BtoS_ACK9_out & ~n6383;
  assign n6385 = ~n6208 & ~n6384;
  assign n6386 = ~reg_i_nEMPTY_out & ~n6385;
  assign n6387 = ~n5177 & ~n6386;
  assign n6388 = ~reg_i_FULL_out & ~n6387;
  assign n6389 = ~n4926 & ~n6388;
  assign n6390 = ~reg_controllable_DEQ_out & ~n6389;
  assign n6391 = ~n4923 & ~n6390;
  assign n6392 = ~reg_controllable_ENQ_out & ~n6391;
  assign n6393 = ~n4922 & ~n6392;
  assign n6394 = ~fair_cnt<2>_out  & ~n6393;
  assign n6395 = ~fair_cnt<2>_out  & ~n6394;
  assign n6396 = ~env_safe_err_happened_out & n6395;
  assign n6397 = ~env_safe_err_happened_out & ~n6396;
  assign n6398 = n75 & ~n6397;
  assign n6399 = n75 & ~n6398;
  assign n6400 = n75 & reg_i_StoB_REQ1_out;
  assign n6401 = n75 & reg_controllable_BtoS_ACK1_out;
  assign n6402 = n6400 & ~n6401;
  assign n6403 = ~i_StoB_REQ1 & n6402;
  assign n6404 = n75 & reg_controllable_BtoS_ACK0_out;
  assign n6405 = ~i_StoB_REQ0 & n6404;
  assign n6406 = n75 & reg_i_StoB_REQ0_out;
  assign n6407 = ~i_StoB_REQ0 & n6406;
  assign n6408 = ~n6404 & ~n6407;
  assign n6409 = ~n6405 & ~n6408;
  assign n6410 = ~n6403 & ~n6409;
  assign n6411 = i_StoB_REQ1 & n6401;
  assign n6412 = n6410 & ~n6411;
  assign n6413 = n75 & reg_i_StoB_REQ2_out;
  assign n6414 = n75 & reg_controllable_BtoS_ACK2_out;
  assign n6415 = n6413 & ~n6414;
  assign n6416 = ~i_StoB_REQ2 & n6415;
  assign n6417 = n6412 & ~n6416;
  assign n6418 = i_StoB_REQ2 & n6414;
  assign n6419 = n6417 & ~n6418;
  assign n6420 = n75 & reg_i_StoB_REQ3_out;
  assign n6421 = n75 & reg_controllable_BtoS_ACK3_out;
  assign n6422 = n6420 & ~n6421;
  assign n6423 = ~i_StoB_REQ3 & n6422;
  assign n6424 = n6419 & ~n6423;
  assign n6425 = i_StoB_REQ3 & n6421;
  assign n6426 = n6424 & ~n6425;
  assign n6427 = n75 & reg_i_StoB_REQ4_out;
  assign n6428 = n75 & reg_controllable_BtoS_ACK4_out;
  assign n6429 = n6427 & ~n6428;
  assign n6430 = ~i_StoB_REQ4 & n6429;
  assign n6431 = n6426 & ~n6430;
  assign n6432 = i_StoB_REQ4 & n6428;
  assign n6433 = n6431 & ~n6432;
  assign n6434 = n75 & reg_i_StoB_REQ5_out;
  assign n6435 = n75 & reg_controllable_BtoS_ACK5_out;
  assign n6436 = n6434 & ~n6435;
  assign n6437 = ~i_StoB_REQ5 & n6436;
  assign n6438 = n6433 & ~n6437;
  assign n6439 = i_StoB_REQ5 & n6435;
  assign n6440 = n6438 & ~n6439;
  assign n6441 = n75 & reg_i_StoB_REQ6_out;
  assign n6442 = n75 & reg_controllable_BtoS_ACK6_out;
  assign n6443 = n6441 & ~n6442;
  assign n6444 = ~i_StoB_REQ6 & n6443;
  assign n6445 = n6440 & ~n6444;
  assign n6446 = i_StoB_REQ6 & n6442;
  assign n6447 = n6445 & ~n6446;
  assign n6448 = n75 & reg_i_StoB_REQ7_out;
  assign n6449 = n75 & reg_controllable_BtoS_ACK7_out;
  assign n6450 = n6448 & ~n6449;
  assign n6451 = ~i_StoB_REQ7 & n6450;
  assign n6452 = n6447 & ~n6451;
  assign n6453 = i_StoB_REQ7 & n6449;
  assign n6454 = n6452 & ~n6453;
  assign n6455 = n75 & reg_i_StoB_REQ8_out;
  assign n6456 = n75 & reg_controllable_BtoS_ACK8_out;
  assign n6457 = n6455 & ~n6456;
  assign n6458 = ~i_StoB_REQ8 & n6457;
  assign n6459 = n6454 & ~n6458;
  assign n6460 = i_StoB_REQ8 & n6456;
  assign n6461 = n6459 & ~n6460;
  assign n6462 = n75 & reg_i_StoB_REQ9_out;
  assign n6463 = n75 & reg_controllable_BtoS_ACK9_out;
  assign n6464 = n6462 & ~n6463;
  assign n6465 = ~i_StoB_REQ9 & n6464;
  assign n6466 = n6461 & ~n6465;
  assign n6467 = i_StoB_REQ9 & n6463;
  assign n6468 = n6466 & ~n6467;
  assign n6469 = n75 & reg_i_StoB_REQ10_out;
  assign n6470 = n75 & reg_controllable_BtoS_ACK10_out;
  assign n6471 = n6469 & ~n6470;
  assign n6472 = ~i_StoB_REQ10 & n6471;
  assign n6473 = n6468 & ~n6472;
  assign n6474 = i_StoB_REQ10 & n6470;
  assign n6475 = n6473 & ~n6474;
  assign n6476 = n75 & reg_i_StoB_REQ11_out;
  assign n6477 = n75 & reg_controllable_BtoS_ACK11_out;
  assign n6478 = n6476 & ~n6477;
  assign n6479 = ~i_StoB_REQ11 & n6478;
  assign n6480 = n6475 & ~n6479;
  assign n6481 = i_StoB_REQ11 & n6477;
  assign n6482 = n6480 & ~n6481;
  assign n6483 = n75 & reg_controllable_BtoR_REQ0_out;
  assign n6484 = i_RtoB_ACK0 & ~n6483;
  assign n6485 = n6482 & ~n6484;
  assign n6486 = n75 & reg_i_RtoB_ACK0_out;
  assign n6487 = ~i_RtoB_ACK0 & n6486;
  assign n6488 = n6483 & n6487;
  assign n6489 = n6485 & ~n6488;
  assign n6490 = n75 & reg_controllable_BtoR_REQ1_out;
  assign n6491 = i_RtoB_ACK1 & ~n6490;
  assign n6492 = n6489 & ~n6491;
  assign n6493 = n75 & reg_i_RtoB_ACK1_out;
  assign n6494 = ~i_RtoB_ACK1 & n6493;
  assign n6495 = n6490 & n6494;
  assign n6496 = n6492 & ~n6495;
  assign n6497 = n75 & reg_controllable_DEQ_out;
  assign n6498 = n75 & reg_controllable_ENQ_out;
  assign n6499 = ~n6497 & n6498;
  assign n6500 = ~i_nEMPTY & n6499;
  assign n6501 = n6496 & ~n6500;
  assign n6502 = n6497 & ~n6498;
  assign n6503 = i_FULL & n6502;
  assign n6504 = n6501 & ~n6503;
  assign n6505 = ~n6499 & ~n6502;
  assign n6506 = n75 & reg_i_FULL_out;
  assign n6507 = i_FULL & ~n6506;
  assign n6508 = ~i_FULL & n6506;
  assign n6509 = ~n6507 & ~n6508;
  assign n6510 = n75 & reg_i_nEMPTY_out;
  assign n6511 = i_nEMPTY & ~n6510;
  assign n6512 = ~i_nEMPTY & n6510;
  assign n6513 = ~n6511 & ~n6512;
  assign n6514 = n6509 & n6513;
  assign n6515 = n6505 & ~n6514;
  assign n6516 = n6504 & ~n6515;
  assign n6517 = n75 & env_safe_err_happened_out;
  assign n6518 = n6516 & ~n6517;
  assign n6519 = n75 & sys_fair8done_out;
  assign n6520 = ~i_StoB_REQ8 & controllable_BtoS_ACK8;
  assign n6521 = i_StoB_REQ8 & ~controllable_BtoS_ACK8;
  assign n6522 = ~n6520 & ~n6521;
  assign n6523 = ~n6519 & ~n6522;
  assign n6524 = ~i_StoB_REQ0 & controllable_BtoS_ACK0;
  assign n6525 = i_StoB_REQ0 & ~controllable_BtoS_ACK0;
  assign n6526 = ~n6524 & ~n6525;
  assign n6527 = n75 & sys_fair0done_out;
  assign n6528 = ~n6526 & ~n6527;
  assign n6529 = ~i_StoB_REQ1 & controllable_BtoS_ACK1;
  assign n6530 = i_StoB_REQ1 & ~controllable_BtoS_ACK1;
  assign n6531 = ~n6529 & ~n6530;
  assign n6532 = n75 & sys_fair1done_out;
  assign n6533 = ~n6531 & ~n6532;
  assign n6534 = ~n6528 & ~n6533;
  assign n6535 = ~i_StoB_REQ2 & controllable_BtoS_ACK2;
  assign n6536 = i_StoB_REQ2 & ~controllable_BtoS_ACK2;
  assign n6537 = ~n6535 & ~n6536;
  assign n6538 = n75 & sys_fair2done_out;
  assign n6539 = ~n6537 & ~n6538;
  assign n6540 = n6534 & ~n6539;
  assign n6541 = ~i_StoB_REQ3 & controllable_BtoS_ACK3;
  assign n6542 = i_StoB_REQ3 & ~controllable_BtoS_ACK3;
  assign n6543 = ~n6541 & ~n6542;
  assign n6544 = n75 & sys_fair3done_out;
  assign n6545 = ~n6543 & ~n6544;
  assign n6546 = n6540 & ~n6545;
  assign n6547 = ~i_StoB_REQ4 & controllable_BtoS_ACK4;
  assign n6548 = i_StoB_REQ4 & ~controllable_BtoS_ACK4;
  assign n6549 = ~n6547 & ~n6548;
  assign n6550 = n75 & sys_fair4done_out;
  assign n6551 = ~n6549 & ~n6550;
  assign n6552 = n6546 & ~n6551;
  assign n6553 = ~i_StoB_REQ5 & controllable_BtoS_ACK5;
  assign n6554 = i_StoB_REQ5 & ~controllable_BtoS_ACK5;
  assign n6555 = ~n6553 & ~n6554;
  assign n6556 = n75 & sys_fair5done_out;
  assign n6557 = ~n6555 & ~n6556;
  assign n6558 = n6552 & ~n6557;
  assign n6559 = ~i_StoB_REQ6 & controllable_BtoS_ACK6;
  assign n6560 = i_StoB_REQ6 & ~controllable_BtoS_ACK6;
  assign n6561 = ~n6559 & ~n6560;
  assign n6562 = n75 & sys_fair6done_out;
  assign n6563 = ~n6561 & ~n6562;
  assign n6564 = n6558 & ~n6563;
  assign n6565 = ~i_StoB_REQ7 & controllable_BtoS_ACK7;
  assign n6566 = i_StoB_REQ7 & ~controllable_BtoS_ACK7;
  assign n6567 = ~n6565 & ~n6566;
  assign n6568 = n75 & sys_fair7done_out;
  assign n6569 = ~n6567 & ~n6568;
  assign n6570 = n6564 & ~n6569;
  assign n6571 = ~n6523 & n6570;
  assign n6572 = ~i_StoB_REQ9 & controllable_BtoS_ACK9;
  assign n6573 = i_StoB_REQ9 & ~controllable_BtoS_ACK9;
  assign n6574 = ~n6572 & ~n6573;
  assign n6575 = n75 & sys_fair9done_out;
  assign n6576 = ~n6574 & ~n6575;
  assign n6577 = n6571 & ~n6576;
  assign n6578 = ~i_StoB_REQ10 & controllable_BtoS_ACK10;
  assign n6579 = i_StoB_REQ10 & ~controllable_BtoS_ACK10;
  assign n6580 = ~n6578 & ~n6579;
  assign n6581 = n75 & sys_fair10done_out;
  assign n6582 = ~n6580 & ~n6581;
  assign n6583 = n6577 & ~n6582;
  assign n6584 = ~i_StoB_REQ11 & controllable_BtoS_ACK11;
  assign n6585 = i_StoB_REQ11 & ~controllable_BtoS_ACK11;
  assign n6586 = ~n6584 & ~n6585;
  assign n6587 = n75 & sys_fair11done_out;
  assign n6588 = ~n6586 & ~n6587;
  assign n6589 = n6583 & ~n6588;
  assign n6590 = n75 & reg_stateG12_out;
  assign n6591 = n75 & sys_fair12done_out;
  assign n6592 = n6590 & ~n6591;
  assign n6593 = n6589 & ~n6592;
  assign n6594 = n6526 & ~n6527;
  assign n6595 = n6531 & ~n6532;
  assign n6596 = ~n6594 & ~n6595;
  assign n6597 = n6537 & ~n6538;
  assign n6598 = n6596 & ~n6597;
  assign n6599 = n6543 & ~n6544;
  assign n6600 = n6598 & ~n6599;
  assign n6601 = n6549 & ~n6550;
  assign n6602 = n6600 & ~n6601;
  assign n6603 = n6555 & ~n6556;
  assign n6604 = n6602 & ~n6603;
  assign n6605 = n6561 & ~n6562;
  assign n6606 = n6604 & ~n6605;
  assign n6607 = n6567 & ~n6568;
  assign n6608 = n6606 & ~n6607;
  assign n6609 = ~n6519 & n6522;
  assign n6610 = n6608 & ~n6609;
  assign n6611 = n6574 & ~n6575;
  assign n6612 = n6610 & ~n6611;
  assign n6613 = n6580 & ~n6581;
  assign n6614 = n6612 & ~n6613;
  assign n6615 = n6586 & ~n6587;
  assign n6616 = n6614 & ~n6615;
  assign n6617 = ~n6590 & ~n6591;
  assign n6618 = n6616 & ~n6617;
  assign n6619 = ~n6593 & n6618;
  assign n6620 = n75 & fair_cnt<2>_out ;
  assign n6621 = i_RtoB_ACK1 & ~controllable_BtoR_REQ1;
  assign n6622 = ~i_RtoB_ACK1 & controllable_BtoR_REQ1;
  assign n6623 = ~n6621 & ~n6622;
  assign n6624 = n75 & env_fair1done_out;
  assign n6625 = ~n6623 & ~n6624;
  assign n6626 = i_RtoB_ACK0 & ~controllable_BtoR_REQ0;
  assign n6627 = ~i_RtoB_ACK0 & controllable_BtoR_REQ0;
  assign n6628 = ~n6626 & ~n6627;
  assign n6629 = n75 & env_fair0done_out;
  assign n6630 = ~n6628 & ~n6629;
  assign n6631 = ~n6625 & ~n6630;
  assign n6632 = n75 & fair_cnt<0>_out ;
  assign n6633 = n6631 & n6632;
  assign n6634 = n75 & fair_cnt<1>_out ;
  assign n6635 = n6633 & n6634;
  assign n6636 = ~n6620 & ~n6635;
  assign n6637 = n6620 & n6635;
  assign n6638 = ~n6636 & ~n6637;
  assign n6639 = n6619 & n6638;
  assign n6640 = ~n6631 & ~n6632;
  assign n6641 = ~n6633 & ~n6640;
  assign n6642 = n6619 & n6641;
  assign n6643 = ~n6633 & n6634;
  assign n6644 = n6633 & ~n6634;
  assign n6645 = ~n6643 & ~n6644;
  assign n6646 = n6619 & ~n6645;
  assign n6647 = ~n6592 & ~n6593;
  assign n6648 = ~n6510 & ~n6590;
  assign n6649 = ~n6497 & ~n6648;
  assign n6650 = n6619 & ~n6631;
  assign n6651 = ~n6625 & n6650;
  assign n6652 = ~n6630 & n6650;
  assign n6653 = n75 & reg_nstateG7_1_out;
  assign n6654 = ~n6483 & n6653;
  assign n6655 = n6483 & ~n6653;
  assign n6656 = ~n6654 & ~n6655;
  assign n6657 = ~n6490 & ~n6656;
  assign n6658 = n6483 & n6653;
  assign n6659 = ~n6657 & ~n6658;
  assign n6660 = ~n6576 & ~n6593;
  assign n6661 = ~n6588 & ~n6593;
  assign n6662 = ~n6582 & ~n6593;
  assign n6663 = ~n6523 & ~n6593;
  assign n6664 = ~n6569 & ~n6593;
  assign n6665 = ~n6563 & ~n6593;
  assign n6666 = ~n6557 & ~n6593;
  assign n6667 = ~n6551 & ~n6593;
  assign n6668 = ~n6545 & ~n6593;
  assign n6669 = ~n6539 & ~n6593;
  assign n6670 = ~n6533 & ~n6593;
  assign n6671 = ~n6528 & ~n6593;
  assign n6672 = i_StoB_REQ0 & controllable_BtoS_ACK0;
  assign n6673 = ~i_StoB_REQ1 & n6672;
  assign n6674 = ~i_StoB_REQ1 & ~n6673;
  assign n6675 = controllable_BtoS_ACK1 & ~n6674;
  assign n6676 = ~controllable_BtoS_ACK1 & n6672;
  assign n6677 = ~n6675 & ~n6676;
  assign n6678 = n6671 & ~n6677;
  assign n6679 = ~i_StoB_REQ0 & ~controllable_BtoS_ACK0;
  assign n6680 = ~n6672 & ~n6679;
  assign n6681 = ~i_StoB_REQ1 & ~n6680;
  assign n6682 = ~i_StoB_REQ1 & ~n6681;
  assign n6683 = controllable_BtoS_ACK1 & ~n6682;
  assign n6684 = ~controllable_BtoS_ACK1 & ~n6680;
  assign n6685 = ~n6683 & ~n6684;
  assign n6686 = ~n6671 & ~n6685;
  assign n6687 = ~n6678 & ~n6686;
  assign n6688 = n6670 & ~n6687;
  assign n6689 = i_StoB_REQ1 & n6672;
  assign n6690 = i_StoB_REQ1 & ~n6689;
  assign n6691 = ~controllable_BtoS_ACK1 & ~n6690;
  assign n6692 = ~n6675 & ~n6691;
  assign n6693 = n6671 & ~n6692;
  assign n6694 = ~n6681 & ~n6689;
  assign n6695 = ~controllable_BtoS_ACK1 & ~n6694;
  assign n6696 = ~n6675 & ~n6695;
  assign n6697 = ~n6671 & ~n6696;
  assign n6698 = ~n6693 & ~n6697;
  assign n6699 = ~n6670 & ~n6698;
  assign n6700 = ~n6688 & ~n6699;
  assign n6701 = n6669 & ~n6700;
  assign n6702 = ~n6669 & ~n6677;
  assign n6703 = ~n6701 & ~n6702;
  assign n6704 = ~i_StoB_REQ2 & ~n6703;
  assign n6705 = ~i_StoB_REQ2 & ~n6704;
  assign n6706 = controllable_BtoS_ACK2 & ~n6705;
  assign n6707 = i_StoB_REQ2 & ~n6703;
  assign n6708 = ~n6671 & ~n6686;
  assign n6709 = n6670 & ~n6708;
  assign n6710 = ~n6699 & ~n6709;
  assign n6711 = ~n6669 & ~n6710;
  assign n6712 = ~n6701 & ~n6711;
  assign n6713 = ~i_StoB_REQ2 & ~n6712;
  assign n6714 = ~n6707 & ~n6713;
  assign n6715 = ~controllable_BtoS_ACK2 & ~n6714;
  assign n6716 = ~n6706 & ~n6715;
  assign n6717 = n6668 & ~n6716;
  assign n6718 = ~i_StoB_REQ2 & ~n6677;
  assign n6719 = ~i_StoB_REQ2 & ~n6718;
  assign n6720 = controllable_BtoS_ACK2 & ~n6719;
  assign n6721 = ~controllable_BtoS_ACK2 & ~n6677;
  assign n6722 = ~n6720 & ~n6721;
  assign n6723 = ~n6668 & ~n6722;
  assign n6724 = ~n6717 & ~n6723;
  assign n6725 = ~i_StoB_REQ3 & ~n6724;
  assign n6726 = ~i_StoB_REQ3 & ~n6725;
  assign n6727 = controllable_BtoS_ACK3 & ~n6726;
  assign n6728 = i_StoB_REQ3 & ~n6724;
  assign n6729 = n6669 & ~n6710;
  assign n6730 = ~n6702 & ~n6729;
  assign n6731 = ~i_StoB_REQ2 & ~n6730;
  assign n6732 = ~i_StoB_REQ2 & ~n6731;
  assign n6733 = controllable_BtoS_ACK2 & ~n6732;
  assign n6734 = i_StoB_REQ2 & ~n6730;
  assign n6735 = ~i_StoB_REQ2 & ~n6710;
  assign n6736 = ~n6734 & ~n6735;
  assign n6737 = ~controllable_BtoS_ACK2 & ~n6736;
  assign n6738 = ~n6733 & ~n6737;
  assign n6739 = ~n6668 & ~n6738;
  assign n6740 = ~n6717 & ~n6739;
  assign n6741 = ~i_StoB_REQ3 & ~n6740;
  assign n6742 = ~n6728 & ~n6741;
  assign n6743 = ~controllable_BtoS_ACK3 & ~n6742;
  assign n6744 = ~n6727 & ~n6743;
  assign n6745 = ~controllable_BtoS_ACK4 & ~n6744;
  assign n6746 = ~controllable_BtoS_ACK4 & ~n6745;
  assign n6747 = n6667 & ~n6746;
  assign n6748 = ~i_StoB_REQ3 & ~n6722;
  assign n6749 = ~i_StoB_REQ3 & ~n6748;
  assign n6750 = controllable_BtoS_ACK3 & ~n6749;
  assign n6751 = ~controllable_BtoS_ACK3 & ~n6722;
  assign n6752 = ~n6750 & ~n6751;
  assign n6753 = ~controllable_BtoS_ACK4 & ~n6752;
  assign n6754 = ~controllable_BtoS_ACK4 & ~n6753;
  assign n6755 = ~n6667 & ~n6754;
  assign n6756 = ~n6747 & ~n6755;
  assign n6757 = i_StoB_REQ4 & ~n6756;
  assign n6758 = n6667 & ~n6744;
  assign n6759 = controllable_BtoS_ACK4 & ~n6752;
  assign n6760 = n6668 & ~n6738;
  assign n6761 = ~n6723 & ~n6760;
  assign n6762 = ~i_StoB_REQ3 & ~n6761;
  assign n6763 = ~i_StoB_REQ3 & ~n6762;
  assign n6764 = controllable_BtoS_ACK3 & ~n6763;
  assign n6765 = i_StoB_REQ3 & ~n6761;
  assign n6766 = ~i_StoB_REQ3 & ~n6738;
  assign n6767 = ~n6765 & ~n6766;
  assign n6768 = ~controllable_BtoS_ACK3 & ~n6767;
  assign n6769 = ~n6764 & ~n6768;
  assign n6770 = ~controllable_BtoS_ACK4 & ~n6769;
  assign n6771 = ~n6759 & ~n6770;
  assign n6772 = ~n6667 & ~n6771;
  assign n6773 = ~n6758 & ~n6772;
  assign n6774 = ~i_StoB_REQ4 & ~n6773;
  assign n6775 = ~n6757 & ~n6774;
  assign n6776 = n6666 & ~n6775;
  assign n6777 = i_StoB_REQ4 & ~n6754;
  assign n6778 = ~i_StoB_REQ4 & ~n6752;
  assign n6779 = ~n6777 & ~n6778;
  assign n6780 = ~n6666 & ~n6779;
  assign n6781 = ~n6776 & ~n6780;
  assign n6782 = ~i_StoB_REQ5 & ~n6781;
  assign n6783 = ~i_StoB_REQ5 & ~n6782;
  assign n6784 = controllable_BtoS_ACK5 & ~n6783;
  assign n6785 = i_StoB_REQ5 & ~n6781;
  assign n6786 = ~controllable_BtoS_ACK4 & ~n6770;
  assign n6787 = n6667 & ~n6786;
  assign n6788 = ~n6755 & ~n6787;
  assign n6789 = i_StoB_REQ4 & ~n6788;
  assign n6790 = n6667 & ~n6769;
  assign n6791 = ~n6772 & ~n6790;
  assign n6792 = ~i_StoB_REQ4 & ~n6791;
  assign n6793 = ~n6789 & ~n6792;
  assign n6794 = ~n6666 & ~n6793;
  assign n6795 = ~n6776 & ~n6794;
  assign n6796 = ~i_StoB_REQ5 & ~n6795;
  assign n6797 = ~n6785 & ~n6796;
  assign n6798 = ~controllable_BtoS_ACK5 & ~n6797;
  assign n6799 = ~n6784 & ~n6798;
  assign n6800 = n6665 & ~n6799;
  assign n6801 = ~i_StoB_REQ5 & ~n6779;
  assign n6802 = ~i_StoB_REQ5 & ~n6801;
  assign n6803 = controllable_BtoS_ACK5 & ~n6802;
  assign n6804 = ~controllable_BtoS_ACK5 & ~n6779;
  assign n6805 = ~n6803 & ~n6804;
  assign n6806 = ~n6665 & ~n6805;
  assign n6807 = ~n6800 & ~n6806;
  assign n6808 = ~i_StoB_REQ6 & ~n6807;
  assign n6809 = ~i_StoB_REQ6 & ~n6808;
  assign n6810 = controllable_BtoS_ACK6 & ~n6809;
  assign n6811 = i_StoB_REQ6 & ~n6807;
  assign n6812 = n6666 & ~n6793;
  assign n6813 = ~n6780 & ~n6812;
  assign n6814 = ~i_StoB_REQ5 & ~n6813;
  assign n6815 = ~i_StoB_REQ5 & ~n6814;
  assign n6816 = controllable_BtoS_ACK5 & ~n6815;
  assign n6817 = i_StoB_REQ5 & ~n6813;
  assign n6818 = ~i_StoB_REQ5 & ~n6793;
  assign n6819 = ~n6817 & ~n6818;
  assign n6820 = ~controllable_BtoS_ACK5 & ~n6819;
  assign n6821 = ~n6816 & ~n6820;
  assign n6822 = ~n6665 & ~n6821;
  assign n6823 = ~n6800 & ~n6822;
  assign n6824 = ~i_StoB_REQ6 & ~n6823;
  assign n6825 = ~n6811 & ~n6824;
  assign n6826 = ~controllable_BtoS_ACK6 & ~n6825;
  assign n6827 = ~n6810 & ~n6826;
  assign n6828 = ~i_StoB_REQ7 & ~n6827;
  assign n6829 = ~i_StoB_REQ7 & ~n6828;
  assign n6830 = n6664 & ~n6829;
  assign n6831 = ~i_StoB_REQ6 & ~n6805;
  assign n6832 = ~i_StoB_REQ6 & ~n6831;
  assign n6833 = controllable_BtoS_ACK6 & ~n6832;
  assign n6834 = ~controllable_BtoS_ACK6 & ~n6805;
  assign n6835 = ~n6833 & ~n6834;
  assign n6836 = ~i_StoB_REQ7 & ~n6835;
  assign n6837 = ~i_StoB_REQ7 & ~n6836;
  assign n6838 = ~n6664 & ~n6837;
  assign n6839 = ~n6830 & ~n6838;
  assign n6840 = controllable_BtoS_ACK7 & ~n6839;
  assign n6841 = n6664 & ~n6827;
  assign n6842 = i_StoB_REQ7 & ~n6835;
  assign n6843 = n6665 & ~n6821;
  assign n6844 = ~n6806 & ~n6843;
  assign n6845 = ~i_StoB_REQ6 & ~n6844;
  assign n6846 = ~i_StoB_REQ6 & ~n6845;
  assign n6847 = controllable_BtoS_ACK6 & ~n6846;
  assign n6848 = i_StoB_REQ6 & ~n6844;
  assign n6849 = ~i_StoB_REQ6 & ~n6821;
  assign n6850 = ~n6848 & ~n6849;
  assign n6851 = ~controllable_BtoS_ACK6 & ~n6850;
  assign n6852 = ~n6847 & ~n6851;
  assign n6853 = ~i_StoB_REQ7 & ~n6852;
  assign n6854 = ~n6842 & ~n6853;
  assign n6855 = ~n6664 & ~n6854;
  assign n6856 = ~n6841 & ~n6855;
  assign n6857 = ~controllable_BtoS_ACK7 & ~n6856;
  assign n6858 = ~n6840 & ~n6857;
  assign n6859 = n6663 & ~n6858;
  assign n6860 = controllable_BtoS_ACK7 & ~n6837;
  assign n6861 = ~controllable_BtoS_ACK7 & ~n6835;
  assign n6862 = ~n6860 & ~n6861;
  assign n6863 = ~n6663 & ~n6862;
  assign n6864 = ~n6859 & ~n6863;
  assign n6865 = ~i_StoB_REQ8 & ~n6864;
  assign n6866 = ~i_StoB_REQ8 & ~n6865;
  assign n6867 = controllable_BtoS_ACK8 & ~n6866;
  assign n6868 = i_StoB_REQ8 & ~n6864;
  assign n6869 = ~i_StoB_REQ7 & ~n6853;
  assign n6870 = n6664 & ~n6869;
  assign n6871 = ~n6838 & ~n6870;
  assign n6872 = controllable_BtoS_ACK7 & ~n6871;
  assign n6873 = n6664 & ~n6852;
  assign n6874 = ~n6855 & ~n6873;
  assign n6875 = ~controllable_BtoS_ACK7 & ~n6874;
  assign n6876 = ~n6872 & ~n6875;
  assign n6877 = ~n6663 & ~n6876;
  assign n6878 = ~n6859 & ~n6877;
  assign n6879 = ~i_StoB_REQ8 & ~n6878;
  assign n6880 = ~n6868 & ~n6879;
  assign n6881 = ~controllable_BtoS_ACK8 & ~n6880;
  assign n6882 = ~n6867 & ~n6881;
  assign n6883 = n6662 & ~n6882;
  assign n6884 = ~i_StoB_REQ8 & ~n6862;
  assign n6885 = ~i_StoB_REQ8 & ~n6884;
  assign n6886 = controllable_BtoS_ACK8 & ~n6885;
  assign n6887 = ~controllable_BtoS_ACK8 & ~n6862;
  assign n6888 = ~n6886 & ~n6887;
  assign n6889 = ~n6662 & ~n6888;
  assign n6890 = ~n6883 & ~n6889;
  assign n6891 = ~i_StoB_REQ10 & ~n6890;
  assign n6892 = ~i_StoB_REQ10 & ~n6891;
  assign n6893 = controllable_BtoS_ACK10 & ~n6892;
  assign n6894 = i_StoB_REQ10 & ~n6890;
  assign n6895 = n6663 & ~n6876;
  assign n6896 = ~n6863 & ~n6895;
  assign n6897 = ~i_StoB_REQ8 & ~n6896;
  assign n6898 = ~i_StoB_REQ8 & ~n6897;
  assign n6899 = controllable_BtoS_ACK8 & ~n6898;
  assign n6900 = i_StoB_REQ8 & ~n6896;
  assign n6901 = ~i_StoB_REQ8 & ~n6876;
  assign n6902 = ~n6900 & ~n6901;
  assign n6903 = ~controllable_BtoS_ACK8 & ~n6902;
  assign n6904 = ~n6899 & ~n6903;
  assign n6905 = ~n6662 & ~n6904;
  assign n6906 = ~n6883 & ~n6905;
  assign n6907 = ~i_StoB_REQ10 & ~n6906;
  assign n6908 = ~n6894 & ~n6907;
  assign n6909 = ~controllable_BtoS_ACK10 & ~n6908;
  assign n6910 = ~n6893 & ~n6909;
  assign n6911 = ~controllable_BtoS_ACK11 & ~n6910;
  assign n6912 = ~controllable_BtoS_ACK11 & ~n6911;
  assign n6913 = n6661 & ~n6912;
  assign n6914 = ~i_StoB_REQ10 & ~n6888;
  assign n6915 = ~i_StoB_REQ10 & ~n6914;
  assign n6916 = controllable_BtoS_ACK10 & ~n6915;
  assign n6917 = ~controllable_BtoS_ACK10 & ~n6888;
  assign n6918 = ~n6916 & ~n6917;
  assign n6919 = ~controllable_BtoS_ACK11 & ~n6918;
  assign n6920 = ~controllable_BtoS_ACK11 & ~n6919;
  assign n6921 = ~n6661 & ~n6920;
  assign n6922 = ~n6913 & ~n6921;
  assign n6923 = i_StoB_REQ11 & ~n6922;
  assign n6924 = ~controllable_BtoS_ACK0 & ~n6679;
  assign n6925 = ~i_StoB_REQ1 & ~n6924;
  assign n6926 = ~i_StoB_REQ1 & ~n6925;
  assign n6927 = controllable_BtoS_ACK1 & ~n6926;
  assign n6928 = ~n6689 & ~n6925;
  assign n6929 = ~controllable_BtoS_ACK1 & ~n6928;
  assign n6930 = ~n6927 & ~n6929;
  assign n6931 = n6671 & ~n6930;
  assign n6932 = i_StoB_REQ1 & ~n6680;
  assign n6933 = ~n6925 & ~n6932;
  assign n6934 = ~controllable_BtoS_ACK1 & ~n6933;
  assign n6935 = ~n6927 & ~n6934;
  assign n6936 = ~n6671 & ~n6935;
  assign n6937 = ~n6931 & ~n6936;
  assign n6938 = n6670 & ~n6937;
  assign n6939 = ~n6691 & ~n6927;
  assign n6940 = n6671 & ~n6939;
  assign n6941 = ~n6671 & ~n6930;
  assign n6942 = ~n6940 & ~n6941;
  assign n6943 = ~n6670 & ~n6942;
  assign n6944 = ~n6938 & ~n6943;
  assign n6945 = n6669 & ~n6944;
  assign n6946 = ~n6669 & ~n6930;
  assign n6947 = ~n6945 & ~n6946;
  assign n6948 = ~i_StoB_REQ2 & ~n6947;
  assign n6949 = ~i_StoB_REQ2 & ~n6948;
  assign n6950 = controllable_BtoS_ACK2 & ~n6949;
  assign n6951 = ~n6671 & ~n6936;
  assign n6952 = n6670 & ~n6951;
  assign n6953 = ~n6943 & ~n6952;
  assign n6954 = ~n6669 & ~n6953;
  assign n6955 = ~n6945 & ~n6954;
  assign n6956 = ~i_StoB_REQ2 & ~n6955;
  assign n6957 = ~n6707 & ~n6956;
  assign n6958 = ~controllable_BtoS_ACK2 & ~n6957;
  assign n6959 = ~n6950 & ~n6958;
  assign n6960 = n6668 & ~n6959;
  assign n6961 = ~i_StoB_REQ2 & ~n6930;
  assign n6962 = ~i_StoB_REQ2 & ~n6961;
  assign n6963 = controllable_BtoS_ACK2 & ~n6962;
  assign n6964 = i_StoB_REQ2 & ~n6677;
  assign n6965 = ~n6961 & ~n6964;
  assign n6966 = ~controllable_BtoS_ACK2 & ~n6965;
  assign n6967 = ~n6963 & ~n6966;
  assign n6968 = ~n6668 & ~n6967;
  assign n6969 = ~n6960 & ~n6968;
  assign n6970 = ~i_StoB_REQ3 & ~n6969;
  assign n6971 = ~i_StoB_REQ3 & ~n6970;
  assign n6972 = controllable_BtoS_ACK3 & ~n6971;
  assign n6973 = n6669 & ~n6953;
  assign n6974 = ~n6946 & ~n6973;
  assign n6975 = ~i_StoB_REQ2 & ~n6974;
  assign n6976 = ~i_StoB_REQ2 & ~n6975;
  assign n6977 = controllable_BtoS_ACK2 & ~n6976;
  assign n6978 = ~i_StoB_REQ2 & ~n6953;
  assign n6979 = ~n6734 & ~n6978;
  assign n6980 = ~controllable_BtoS_ACK2 & ~n6979;
  assign n6981 = ~n6977 & ~n6980;
  assign n6982 = ~n6668 & ~n6981;
  assign n6983 = ~n6960 & ~n6982;
  assign n6984 = ~i_StoB_REQ3 & ~n6983;
  assign n6985 = ~n6728 & ~n6984;
  assign n6986 = ~controllable_BtoS_ACK3 & ~n6985;
  assign n6987 = ~n6972 & ~n6986;
  assign n6988 = n6667 & ~n6987;
  assign n6989 = ~i_StoB_REQ3 & ~n6967;
  assign n6990 = ~i_StoB_REQ3 & ~n6989;
  assign n6991 = controllable_BtoS_ACK3 & ~n6990;
  assign n6992 = i_StoB_REQ3 & ~n6722;
  assign n6993 = ~n6989 & ~n6992;
  assign n6994 = ~controllable_BtoS_ACK3 & ~n6993;
  assign n6995 = ~n6991 & ~n6994;
  assign n6996 = controllable_BtoS_ACK4 & ~n6995;
  assign n6997 = n6668 & ~n6981;
  assign n6998 = ~n6968 & ~n6997;
  assign n6999 = ~i_StoB_REQ3 & ~n6998;
  assign n7000 = ~i_StoB_REQ3 & ~n6999;
  assign n7001 = controllable_BtoS_ACK3 & ~n7000;
  assign n7002 = ~i_StoB_REQ3 & ~n6981;
  assign n7003 = ~n6765 & ~n7002;
  assign n7004 = ~controllable_BtoS_ACK3 & ~n7003;
  assign n7005 = ~n7001 & ~n7004;
  assign n7006 = ~controllable_BtoS_ACK4 & ~n7005;
  assign n7007 = ~n6996 & ~n7006;
  assign n7008 = ~n6667 & ~n7007;
  assign n7009 = ~n6988 & ~n7008;
  assign n7010 = ~i_StoB_REQ4 & ~n7009;
  assign n7011 = ~n6757 & ~n7010;
  assign n7012 = n6666 & ~n7011;
  assign n7013 = ~i_StoB_REQ4 & ~n6995;
  assign n7014 = ~n6777 & ~n7013;
  assign n7015 = ~n6666 & ~n7014;
  assign n7016 = ~n7012 & ~n7015;
  assign n7017 = ~i_StoB_REQ5 & ~n7016;
  assign n7018 = ~i_StoB_REQ5 & ~n7017;
  assign n7019 = controllable_BtoS_ACK5 & ~n7018;
  assign n7020 = n6667 & ~n7005;
  assign n7021 = ~n7008 & ~n7020;
  assign n7022 = ~i_StoB_REQ4 & ~n7021;
  assign n7023 = ~n6789 & ~n7022;
  assign n7024 = ~n6666 & ~n7023;
  assign n7025 = ~n7012 & ~n7024;
  assign n7026 = ~i_StoB_REQ5 & ~n7025;
  assign n7027 = ~n6785 & ~n7026;
  assign n7028 = ~controllable_BtoS_ACK5 & ~n7027;
  assign n7029 = ~n7019 & ~n7028;
  assign n7030 = n6665 & ~n7029;
  assign n7031 = ~i_StoB_REQ5 & ~n7014;
  assign n7032 = ~i_StoB_REQ5 & ~n7031;
  assign n7033 = controllable_BtoS_ACK5 & ~n7032;
  assign n7034 = i_StoB_REQ5 & ~n6779;
  assign n7035 = ~n7031 & ~n7034;
  assign n7036 = ~controllable_BtoS_ACK5 & ~n7035;
  assign n7037 = ~n7033 & ~n7036;
  assign n7038 = ~n6665 & ~n7037;
  assign n7039 = ~n7030 & ~n7038;
  assign n7040 = ~i_StoB_REQ6 & ~n7039;
  assign n7041 = ~i_StoB_REQ6 & ~n7040;
  assign n7042 = controllable_BtoS_ACK6 & ~n7041;
  assign n7043 = n6666 & ~n7023;
  assign n7044 = ~n7015 & ~n7043;
  assign n7045 = ~i_StoB_REQ5 & ~n7044;
  assign n7046 = ~i_StoB_REQ5 & ~n7045;
  assign n7047 = controllable_BtoS_ACK5 & ~n7046;
  assign n7048 = ~i_StoB_REQ5 & ~n7023;
  assign n7049 = ~n6817 & ~n7048;
  assign n7050 = ~controllable_BtoS_ACK5 & ~n7049;
  assign n7051 = ~n7047 & ~n7050;
  assign n7052 = ~n6665 & ~n7051;
  assign n7053 = ~n7030 & ~n7052;
  assign n7054 = ~i_StoB_REQ6 & ~n7053;
  assign n7055 = ~n6811 & ~n7054;
  assign n7056 = ~controllable_BtoS_ACK6 & ~n7055;
  assign n7057 = ~n7042 & ~n7056;
  assign n7058 = ~i_StoB_REQ7 & ~n7057;
  assign n7059 = ~i_StoB_REQ7 & ~n7058;
  assign n7060 = n6664 & ~n7059;
  assign n7061 = ~i_StoB_REQ6 & ~n7037;
  assign n7062 = ~i_StoB_REQ6 & ~n7061;
  assign n7063 = controllable_BtoS_ACK6 & ~n7062;
  assign n7064 = i_StoB_REQ6 & ~n6805;
  assign n7065 = ~n7061 & ~n7064;
  assign n7066 = ~controllable_BtoS_ACK6 & ~n7065;
  assign n7067 = ~n7063 & ~n7066;
  assign n7068 = ~i_StoB_REQ7 & ~n7067;
  assign n7069 = ~i_StoB_REQ7 & ~n7068;
  assign n7070 = ~n6664 & ~n7069;
  assign n7071 = ~n7060 & ~n7070;
  assign n7072 = controllable_BtoS_ACK7 & ~n7071;
  assign n7073 = i_StoB_REQ7 & ~n6827;
  assign n7074 = ~n7058 & ~n7073;
  assign n7075 = n6664 & ~n7074;
  assign n7076 = n6665 & ~n7051;
  assign n7077 = ~n7038 & ~n7076;
  assign n7078 = ~i_StoB_REQ6 & ~n7077;
  assign n7079 = ~i_StoB_REQ6 & ~n7078;
  assign n7080 = controllable_BtoS_ACK6 & ~n7079;
  assign n7081 = ~i_StoB_REQ6 & ~n7051;
  assign n7082 = ~n6848 & ~n7081;
  assign n7083 = ~controllable_BtoS_ACK6 & ~n7082;
  assign n7084 = ~n7080 & ~n7083;
  assign n7085 = ~i_StoB_REQ7 & ~n7084;
  assign n7086 = ~n6842 & ~n7085;
  assign n7087 = ~n6664 & ~n7086;
  assign n7088 = ~n7075 & ~n7087;
  assign n7089 = ~controllable_BtoS_ACK7 & ~n7088;
  assign n7090 = ~n7072 & ~n7089;
  assign n7091 = n6663 & ~n7090;
  assign n7092 = controllable_BtoS_ACK7 & ~n7069;
  assign n7093 = ~n6842 & ~n7068;
  assign n7094 = ~controllable_BtoS_ACK7 & ~n7093;
  assign n7095 = ~n7092 & ~n7094;
  assign n7096 = ~n6663 & ~n7095;
  assign n7097 = ~n7091 & ~n7096;
  assign n7098 = ~i_StoB_REQ8 & ~n7097;
  assign n7099 = ~i_StoB_REQ8 & ~n7098;
  assign n7100 = controllable_BtoS_ACK8 & ~n7099;
  assign n7101 = ~i_StoB_REQ7 & ~n7085;
  assign n7102 = n6664 & ~n7101;
  assign n7103 = ~n7070 & ~n7102;
  assign n7104 = controllable_BtoS_ACK7 & ~n7103;
  assign n7105 = i_StoB_REQ7 & ~n6852;
  assign n7106 = ~n7085 & ~n7105;
  assign n7107 = n6664 & ~n7106;
  assign n7108 = ~n7087 & ~n7107;
  assign n7109 = ~controllable_BtoS_ACK7 & ~n7108;
  assign n7110 = ~n7104 & ~n7109;
  assign n7111 = ~n6663 & ~n7110;
  assign n7112 = ~n7091 & ~n7111;
  assign n7113 = ~i_StoB_REQ8 & ~n7112;
  assign n7114 = ~n6868 & ~n7113;
  assign n7115 = ~controllable_BtoS_ACK8 & ~n7114;
  assign n7116 = ~n7100 & ~n7115;
  assign n7117 = n6662 & ~n7116;
  assign n7118 = ~i_StoB_REQ8 & ~n7095;
  assign n7119 = ~i_StoB_REQ8 & ~n7118;
  assign n7120 = controllable_BtoS_ACK8 & ~n7119;
  assign n7121 = i_StoB_REQ8 & ~n6862;
  assign n7122 = ~n7118 & ~n7121;
  assign n7123 = ~controllable_BtoS_ACK8 & ~n7122;
  assign n7124 = ~n7120 & ~n7123;
  assign n7125 = ~n6662 & ~n7124;
  assign n7126 = ~n7117 & ~n7125;
  assign n7127 = ~i_StoB_REQ10 & ~n7126;
  assign n7128 = ~i_StoB_REQ10 & ~n7127;
  assign n7129 = controllable_BtoS_ACK10 & ~n7128;
  assign n7130 = n6663 & ~n7110;
  assign n7131 = ~n7096 & ~n7130;
  assign n7132 = ~i_StoB_REQ8 & ~n7131;
  assign n7133 = ~i_StoB_REQ8 & ~n7132;
  assign n7134 = controllable_BtoS_ACK8 & ~n7133;
  assign n7135 = ~i_StoB_REQ8 & ~n7110;
  assign n7136 = ~n6900 & ~n7135;
  assign n7137 = ~controllable_BtoS_ACK8 & ~n7136;
  assign n7138 = ~n7134 & ~n7137;
  assign n7139 = ~n6662 & ~n7138;
  assign n7140 = ~n7117 & ~n7139;
  assign n7141 = ~i_StoB_REQ10 & ~n7140;
  assign n7142 = ~n6894 & ~n7141;
  assign n7143 = ~controllable_BtoS_ACK10 & ~n7142;
  assign n7144 = ~n7129 & ~n7143;
  assign n7145 = n6661 & ~n7144;
  assign n7146 = ~i_StoB_REQ10 & ~n7124;
  assign n7147 = ~i_StoB_REQ10 & ~n7146;
  assign n7148 = controllable_BtoS_ACK10 & ~n7147;
  assign n7149 = i_StoB_REQ10 & ~n6888;
  assign n7150 = ~n7146 & ~n7149;
  assign n7151 = ~controllable_BtoS_ACK10 & ~n7150;
  assign n7152 = ~n7148 & ~n7151;
  assign n7153 = controllable_BtoS_ACK11 & ~n7152;
  assign n7154 = n6662 & ~n7138;
  assign n7155 = ~n7125 & ~n7154;
  assign n7156 = ~i_StoB_REQ10 & ~n7155;
  assign n7157 = ~i_StoB_REQ10 & ~n7156;
  assign n7158 = controllable_BtoS_ACK10 & ~n7157;
  assign n7159 = n6662 & ~n6904;
  assign n7160 = ~n6889 & ~n7159;
  assign n7161 = i_StoB_REQ10 & ~n7160;
  assign n7162 = ~i_StoB_REQ10 & ~n7138;
  assign n7163 = ~n7161 & ~n7162;
  assign n7164 = ~controllable_BtoS_ACK10 & ~n7163;
  assign n7165 = ~n7158 & ~n7164;
  assign n7166 = ~controllable_BtoS_ACK11 & ~n7165;
  assign n7167 = ~n7153 & ~n7166;
  assign n7168 = ~n6661 & ~n7167;
  assign n7169 = ~n7145 & ~n7168;
  assign n7170 = ~i_StoB_REQ11 & ~n7169;
  assign n7171 = ~n6923 & ~n7170;
  assign n7172 = controllable_ENQ & ~n7171;
  assign n7173 = controllable_ENQ & ~n7172;
  assign n7174 = ~i_StoB_REQ9 & ~n7173;
  assign n7175 = ~i_StoB_REQ9 & ~n7174;
  assign n7176 = controllable_BtoS_ACK9 & ~n7175;
  assign n7177 = n6661 & ~n6910;
  assign n7178 = controllable_BtoS_ACK11 & ~n6918;
  assign n7179 = ~i_StoB_REQ10 & ~n7160;
  assign n7180 = ~i_StoB_REQ10 & ~n7179;
  assign n7181 = controllable_BtoS_ACK10 & ~n7180;
  assign n7182 = ~i_StoB_REQ10 & ~n6904;
  assign n7183 = ~n7161 & ~n7182;
  assign n7184 = ~controllable_BtoS_ACK10 & ~n7183;
  assign n7185 = ~n7181 & ~n7184;
  assign n7186 = ~controllable_BtoS_ACK11 & ~n7185;
  assign n7187 = ~n7178 & ~n7186;
  assign n7188 = ~n6661 & ~n7187;
  assign n7189 = ~n7177 & ~n7188;
  assign n7190 = ~i_StoB_REQ11 & ~n7189;
  assign n7191 = ~n6923 & ~n7190;
  assign n7192 = controllable_ENQ & ~n7191;
  assign n7193 = controllable_ENQ & ~n7192;
  assign n7194 = i_StoB_REQ9 & ~n7193;
  assign n7195 = ~n7174 & ~n7194;
  assign n7196 = ~controllable_BtoS_ACK9 & ~n7195;
  assign n7197 = ~n7176 & ~n7196;
  assign n7198 = controllable_DEQ & ~n7197;
  assign n7199 = ~i_StoB_REQ9 & ~n7171;
  assign n7200 = ~i_StoB_REQ9 & ~n7199;
  assign n7201 = controllable_BtoS_ACK9 & ~n7200;
  assign n7202 = i_StoB_REQ9 & ~n7191;
  assign n7203 = ~n7199 & ~n7202;
  assign n7204 = ~controllable_BtoS_ACK9 & ~n7203;
  assign n7205 = ~n7201 & ~n7204;
  assign n7206 = ~controllable_DEQ & ~n7205;
  assign n7207 = ~n7198 & ~n7206;
  assign n7208 = i_nEMPTY & ~n7207;
  assign n7209 = ~controllable_DEQ & ~n7197;
  assign n7210 = ~controllable_DEQ & ~n7209;
  assign n7211 = ~i_nEMPTY & ~n7210;
  assign n7212 = ~n7208 & ~n7211;
  assign n7213 = i_RtoB_ACK0 & ~n7212;
  assign n7214 = controllable_BtoS_ACK0 & ~n6672;
  assign n7215 = ~i_StoB_REQ1 & ~n7214;
  assign n7216 = ~i_StoB_REQ1 & ~n7215;
  assign n7217 = controllable_BtoS_ACK1 & ~n7216;
  assign n7218 = ~controllable_BtoS_ACK1 & ~n7214;
  assign n7219 = ~n7217 & ~n7218;
  assign n7220 = ~n6671 & ~n7219;
  assign n7221 = ~n6678 & ~n7220;
  assign n7222 = n6670 & ~n7221;
  assign n7223 = controllable_BtoS_ACK1 & ~n6675;
  assign n7224 = n6671 & ~n7223;
  assign n7225 = ~n6675 & ~n7218;
  assign n7226 = ~n6671 & ~n7225;
  assign n7227 = ~n7224 & ~n7226;
  assign n7228 = ~n6670 & ~n7227;
  assign n7229 = ~n7222 & ~n7228;
  assign n7230 = n6669 & ~n7229;
  assign n7231 = ~n6702 & ~n7230;
  assign n7232 = ~i_StoB_REQ2 & ~n7231;
  assign n7233 = ~i_StoB_REQ2 & ~n7232;
  assign n7234 = controllable_BtoS_ACK2 & ~n7233;
  assign n7235 = ~n6671 & ~n7220;
  assign n7236 = n6670 & ~n7235;
  assign n7237 = ~n7228 & ~n7236;
  assign n7238 = ~n6669 & ~n7237;
  assign n7239 = ~n7230 & ~n7238;
  assign n7240 = ~controllable_BtoS_ACK2 & ~n7239;
  assign n7241 = ~n7234 & ~n7240;
  assign n7242 = n6668 & ~n7241;
  assign n7243 = ~n6723 & ~n7242;
  assign n7244 = ~i_StoB_REQ3 & ~n7243;
  assign n7245 = ~i_StoB_REQ3 & ~n7244;
  assign n7246 = controllable_BtoS_ACK3 & ~n7245;
  assign n7247 = n6669 & ~n7237;
  assign n7248 = ~n6702 & ~n7247;
  assign n7249 = ~i_StoB_REQ2 & ~n7248;
  assign n7250 = ~i_StoB_REQ2 & ~n7249;
  assign n7251 = controllable_BtoS_ACK2 & ~n7250;
  assign n7252 = ~controllable_BtoS_ACK2 & ~n7237;
  assign n7253 = ~n7251 & ~n7252;
  assign n7254 = ~n6668 & ~n7253;
  assign n7255 = ~n7242 & ~n7254;
  assign n7256 = ~controllable_BtoS_ACK3 & ~n7255;
  assign n7257 = ~n7246 & ~n7256;
  assign n7258 = ~controllable_BtoS_ACK4 & ~n7257;
  assign n7259 = ~controllable_BtoS_ACK4 & ~n7258;
  assign n7260 = n6667 & ~n7259;
  assign n7261 = n6668 & ~n7253;
  assign n7262 = ~n6723 & ~n7261;
  assign n7263 = ~i_StoB_REQ3 & ~n7262;
  assign n7264 = ~i_StoB_REQ3 & ~n7263;
  assign n7265 = controllable_BtoS_ACK3 & ~n7264;
  assign n7266 = ~controllable_BtoS_ACK3 & ~n7253;
  assign n7267 = ~n7265 & ~n7266;
  assign n7268 = ~controllable_BtoS_ACK4 & ~n7267;
  assign n7269 = ~controllable_BtoS_ACK4 & ~n7268;
  assign n7270 = ~n6667 & ~n7269;
  assign n7271 = ~n7260 & ~n7270;
  assign n7272 = i_StoB_REQ4 & ~n7271;
  assign n7273 = n6667 & ~n7257;
  assign n7274 = ~n6759 & ~n7268;
  assign n7275 = ~n6667 & ~n7274;
  assign n7276 = ~n7273 & ~n7275;
  assign n7277 = ~i_StoB_REQ4 & ~n7276;
  assign n7278 = ~n7272 & ~n7277;
  assign n7279 = n6666 & ~n7278;
  assign n7280 = ~n6780 & ~n7279;
  assign n7281 = ~i_StoB_REQ5 & ~n7280;
  assign n7282 = ~i_StoB_REQ5 & ~n7281;
  assign n7283 = controllable_BtoS_ACK5 & ~n7282;
  assign n7284 = i_StoB_REQ4 & ~n7269;
  assign n7285 = n6667 & ~n7267;
  assign n7286 = ~n7275 & ~n7285;
  assign n7287 = ~i_StoB_REQ4 & ~n7286;
  assign n7288 = ~n7284 & ~n7287;
  assign n7289 = ~n6666 & ~n7288;
  assign n7290 = ~n7279 & ~n7289;
  assign n7291 = ~controllable_BtoS_ACK5 & ~n7290;
  assign n7292 = ~n7283 & ~n7291;
  assign n7293 = n6665 & ~n7292;
  assign n7294 = ~n6806 & ~n7293;
  assign n7295 = ~i_StoB_REQ6 & ~n7294;
  assign n7296 = ~i_StoB_REQ6 & ~n7295;
  assign n7297 = controllable_BtoS_ACK6 & ~n7296;
  assign n7298 = n6666 & ~n7288;
  assign n7299 = ~n6780 & ~n7298;
  assign n7300 = ~i_StoB_REQ5 & ~n7299;
  assign n7301 = ~i_StoB_REQ5 & ~n7300;
  assign n7302 = controllable_BtoS_ACK5 & ~n7301;
  assign n7303 = ~controllable_BtoS_ACK5 & ~n7288;
  assign n7304 = ~n7302 & ~n7303;
  assign n7305 = ~n6665 & ~n7304;
  assign n7306 = ~n7293 & ~n7305;
  assign n7307 = ~controllable_BtoS_ACK6 & ~n7306;
  assign n7308 = ~n7297 & ~n7307;
  assign n7309 = ~i_StoB_REQ7 & ~n7308;
  assign n7310 = ~i_StoB_REQ7 & ~n7309;
  assign n7311 = n6664 & ~n7310;
  assign n7312 = ~n6838 & ~n7311;
  assign n7313 = controllable_BtoS_ACK7 & ~n7312;
  assign n7314 = n6664 & ~n7308;
  assign n7315 = n6665 & ~n7304;
  assign n7316 = ~n6806 & ~n7315;
  assign n7317 = ~i_StoB_REQ6 & ~n7316;
  assign n7318 = ~i_StoB_REQ6 & ~n7317;
  assign n7319 = controllable_BtoS_ACK6 & ~n7318;
  assign n7320 = ~controllable_BtoS_ACK6 & ~n7304;
  assign n7321 = ~n7319 & ~n7320;
  assign n7322 = ~n6664 & ~n7321;
  assign n7323 = ~n7314 & ~n7322;
  assign n7324 = ~controllable_BtoS_ACK7 & ~n7323;
  assign n7325 = ~n7313 & ~n7324;
  assign n7326 = n6663 & ~n7325;
  assign n7327 = ~n6863 & ~n7326;
  assign n7328 = ~i_StoB_REQ8 & ~n7327;
  assign n7329 = ~i_StoB_REQ8 & ~n7328;
  assign n7330 = controllable_BtoS_ACK8 & ~n7329;
  assign n7331 = ~i_StoB_REQ7 & ~n7321;
  assign n7332 = ~i_StoB_REQ7 & ~n7331;
  assign n7333 = n6664 & ~n7332;
  assign n7334 = ~n6838 & ~n7333;
  assign n7335 = controllable_BtoS_ACK7 & ~n7334;
  assign n7336 = ~controllable_BtoS_ACK7 & ~n7321;
  assign n7337 = ~n7335 & ~n7336;
  assign n7338 = ~n6663 & ~n7337;
  assign n7339 = ~n7326 & ~n7338;
  assign n7340 = ~controllable_BtoS_ACK8 & ~n7339;
  assign n7341 = ~n7330 & ~n7340;
  assign n7342 = n6662 & ~n7341;
  assign n7343 = ~n6889 & ~n7342;
  assign n7344 = ~i_StoB_REQ10 & ~n7343;
  assign n7345 = ~i_StoB_REQ10 & ~n7344;
  assign n7346 = controllable_BtoS_ACK10 & ~n7345;
  assign n7347 = n6663 & ~n7337;
  assign n7348 = ~n6863 & ~n7347;
  assign n7349 = ~i_StoB_REQ8 & ~n7348;
  assign n7350 = ~i_StoB_REQ8 & ~n7349;
  assign n7351 = controllable_BtoS_ACK8 & ~n7350;
  assign n7352 = ~controllable_BtoS_ACK8 & ~n7337;
  assign n7353 = ~n7351 & ~n7352;
  assign n7354 = ~n6662 & ~n7353;
  assign n7355 = ~n7342 & ~n7354;
  assign n7356 = ~controllable_BtoS_ACK10 & ~n7355;
  assign n7357 = ~n7346 & ~n7356;
  assign n7358 = ~controllable_BtoS_ACK11 & ~n7357;
  assign n7359 = ~controllable_BtoS_ACK11 & ~n7358;
  assign n7360 = n6661 & ~n7359;
  assign n7361 = n6662 & ~n7353;
  assign n7362 = ~n6889 & ~n7361;
  assign n7363 = ~i_StoB_REQ10 & ~n7362;
  assign n7364 = ~i_StoB_REQ10 & ~n7363;
  assign n7365 = controllable_BtoS_ACK10 & ~n7364;
  assign n7366 = ~controllable_BtoS_ACK10 & ~n7353;
  assign n7367 = ~n7365 & ~n7366;
  assign n7368 = ~controllable_BtoS_ACK11 & ~n7367;
  assign n7369 = ~controllable_BtoS_ACK11 & ~n7368;
  assign n7370 = ~n6661 & ~n7369;
  assign n7371 = ~n7360 & ~n7370;
  assign n7372 = i_StoB_REQ11 & ~n7371;
  assign n7373 = n6661 & ~n7357;
  assign n7374 = ~n7178 & ~n7368;
  assign n7375 = ~n6661 & ~n7374;
  assign n7376 = ~n7373 & ~n7375;
  assign n7377 = ~i_StoB_REQ11 & ~n7376;
  assign n7378 = ~n7372 & ~n7377;
  assign n7379 = controllable_ENQ & ~n7378;
  assign n7380 = controllable_ENQ & ~n7379;
  assign n7381 = i_StoB_REQ9 & ~n7380;
  assign n7382 = controllable_BtoS_ACK11 & ~n7357;
  assign n7383 = i_StoB_REQ10 & ~n7355;
  assign n7384 = i_StoB_REQ8 & ~n7339;
  assign n7385 = i_StoB_REQ7 & ~n7308;
  assign n7386 = i_StoB_REQ6 & ~n7306;
  assign n7387 = i_StoB_REQ5 & ~n7290;
  assign n7388 = controllable_BtoS_ACK4 & ~n7257;
  assign n7389 = i_StoB_REQ3 & ~n7255;
  assign n7390 = i_StoB_REQ2 & ~n7239;
  assign n7391 = controllable_BtoS_ACK1 & n6689;
  assign n7392 = n6671 & n7391;
  assign n7393 = ~n6671 & ~n7214;
  assign n7394 = ~n7392 & ~n7393;
  assign n7395 = n6670 & ~n7394;
  assign n7396 = i_StoB_REQ1 & controllable_BtoS_ACK1;
  assign n7397 = controllable_BtoS_ACK1 & ~n7396;
  assign n7398 = n6671 & ~n7397;
  assign n7399 = i_StoB_REQ1 & ~n7214;
  assign n7400 = controllable_BtoS_ACK1 & n7399;
  assign n7401 = ~n7218 & ~n7400;
  assign n7402 = ~n6671 & ~n7401;
  assign n7403 = ~n7398 & ~n7402;
  assign n7404 = ~n6670 & ~n7403;
  assign n7405 = ~n7395 & ~n7404;
  assign n7406 = n6669 & ~n7405;
  assign n7407 = ~n6669 & n7391;
  assign n7408 = ~n7406 & ~n7407;
  assign n7409 = ~i_StoB_REQ2 & ~n7408;
  assign n7410 = ~n7390 & ~n7409;
  assign n7411 = controllable_BtoS_ACK2 & ~n7410;
  assign n7412 = ~n6671 & ~n7393;
  assign n7413 = n6670 & ~n7412;
  assign n7414 = ~n7404 & ~n7413;
  assign n7415 = ~n6669 & ~n7414;
  assign n7416 = ~n7406 & ~n7415;
  assign n7417 = ~controllable_BtoS_ACK2 & ~n7416;
  assign n7418 = ~n7411 & ~n7417;
  assign n7419 = n6668 & ~n7418;
  assign n7420 = ~i_StoB_REQ2 & n7391;
  assign n7421 = ~n6964 & ~n7420;
  assign n7422 = controllable_BtoS_ACK2 & ~n7421;
  assign n7423 = ~controllable_BtoS_ACK2 & n7391;
  assign n7424 = ~n7422 & ~n7423;
  assign n7425 = ~n6668 & ~n7424;
  assign n7426 = ~n7419 & ~n7425;
  assign n7427 = ~i_StoB_REQ3 & ~n7426;
  assign n7428 = ~n7389 & ~n7427;
  assign n7429 = controllable_BtoS_ACK3 & ~n7428;
  assign n7430 = i_StoB_REQ2 & ~n7237;
  assign n7431 = n6669 & ~n7414;
  assign n7432 = ~n7407 & ~n7431;
  assign n7433 = ~i_StoB_REQ2 & ~n7432;
  assign n7434 = ~n7430 & ~n7433;
  assign n7435 = controllable_BtoS_ACK2 & ~n7434;
  assign n7436 = ~controllable_BtoS_ACK2 & ~n7414;
  assign n7437 = ~n7435 & ~n7436;
  assign n7438 = ~n6668 & ~n7437;
  assign n7439 = ~n7419 & ~n7438;
  assign n7440 = ~controllable_BtoS_ACK3 & ~n7439;
  assign n7441 = ~n7429 & ~n7440;
  assign n7442 = ~controllable_BtoS_ACK4 & ~n7441;
  assign n7443 = ~n7388 & ~n7442;
  assign n7444 = n6667 & ~n7443;
  assign n7445 = controllable_BtoS_ACK4 & ~n7267;
  assign n7446 = i_StoB_REQ3 & ~n7253;
  assign n7447 = n6668 & ~n7437;
  assign n7448 = ~n7425 & ~n7447;
  assign n7449 = ~i_StoB_REQ3 & ~n7448;
  assign n7450 = ~n7446 & ~n7449;
  assign n7451 = controllable_BtoS_ACK3 & ~n7450;
  assign n7452 = ~controllable_BtoS_ACK3 & ~n7437;
  assign n7453 = ~n7451 & ~n7452;
  assign n7454 = ~controllable_BtoS_ACK4 & ~n7453;
  assign n7455 = ~n7445 & ~n7454;
  assign n7456 = ~n6667 & ~n7455;
  assign n7457 = ~n7444 & ~n7456;
  assign n7458 = i_StoB_REQ4 & ~n7457;
  assign n7459 = n6667 & ~n7441;
  assign n7460 = ~i_StoB_REQ3 & ~n7424;
  assign n7461 = ~n6992 & ~n7460;
  assign n7462 = controllable_BtoS_ACK3 & ~n7461;
  assign n7463 = ~controllable_BtoS_ACK3 & ~n7424;
  assign n7464 = ~n7462 & ~n7463;
  assign n7465 = controllable_BtoS_ACK4 & ~n7464;
  assign n7466 = ~n7454 & ~n7465;
  assign n7467 = ~n6667 & ~n7466;
  assign n7468 = ~n7459 & ~n7467;
  assign n7469 = ~i_StoB_REQ4 & ~n7468;
  assign n7470 = ~n7458 & ~n7469;
  assign n7471 = n6666 & ~n7470;
  assign n7472 = ~controllable_BtoS_ACK4 & ~n7464;
  assign n7473 = ~n6759 & ~n7472;
  assign n7474 = i_StoB_REQ4 & ~n7473;
  assign n7475 = ~i_StoB_REQ4 & ~n7464;
  assign n7476 = ~n7474 & ~n7475;
  assign n7477 = ~n6666 & ~n7476;
  assign n7478 = ~n7471 & ~n7477;
  assign n7479 = ~i_StoB_REQ5 & ~n7478;
  assign n7480 = ~n7387 & ~n7479;
  assign n7481 = controllable_BtoS_ACK5 & ~n7480;
  assign n7482 = i_StoB_REQ4 & ~n7455;
  assign n7483 = n6667 & ~n7453;
  assign n7484 = ~n7467 & ~n7483;
  assign n7485 = ~i_StoB_REQ4 & ~n7484;
  assign n7486 = ~n7482 & ~n7485;
  assign n7487 = ~n6666 & ~n7486;
  assign n7488 = ~n7471 & ~n7487;
  assign n7489 = ~controllable_BtoS_ACK5 & ~n7488;
  assign n7490 = ~n7481 & ~n7489;
  assign n7491 = n6665 & ~n7490;
  assign n7492 = ~i_StoB_REQ5 & ~n7476;
  assign n7493 = ~n7034 & ~n7492;
  assign n7494 = controllable_BtoS_ACK5 & ~n7493;
  assign n7495 = ~controllable_BtoS_ACK5 & ~n7476;
  assign n7496 = ~n7494 & ~n7495;
  assign n7497 = ~n6665 & ~n7496;
  assign n7498 = ~n7491 & ~n7497;
  assign n7499 = ~i_StoB_REQ6 & ~n7498;
  assign n7500 = ~n7386 & ~n7499;
  assign n7501 = controllable_BtoS_ACK6 & ~n7500;
  assign n7502 = i_StoB_REQ5 & ~n7288;
  assign n7503 = n6666 & ~n7486;
  assign n7504 = ~n7477 & ~n7503;
  assign n7505 = ~i_StoB_REQ5 & ~n7504;
  assign n7506 = ~n7502 & ~n7505;
  assign n7507 = controllable_BtoS_ACK5 & ~n7506;
  assign n7508 = ~controllable_BtoS_ACK5 & ~n7486;
  assign n7509 = ~n7507 & ~n7508;
  assign n7510 = ~n6665 & ~n7509;
  assign n7511 = ~n7491 & ~n7510;
  assign n7512 = ~controllable_BtoS_ACK6 & ~n7511;
  assign n7513 = ~n7501 & ~n7512;
  assign n7514 = ~i_StoB_REQ7 & ~n7513;
  assign n7515 = ~n7385 & ~n7514;
  assign n7516 = n6664 & ~n7515;
  assign n7517 = i_StoB_REQ7 & ~n7321;
  assign n7518 = ~i_StoB_REQ6 & ~n7496;
  assign n7519 = ~n7064 & ~n7518;
  assign n7520 = controllable_BtoS_ACK6 & ~n7519;
  assign n7521 = ~controllable_BtoS_ACK6 & ~n7496;
  assign n7522 = ~n7520 & ~n7521;
  assign n7523 = ~i_StoB_REQ7 & ~n7522;
  assign n7524 = ~n7517 & ~n7523;
  assign n7525 = ~n6664 & ~n7524;
  assign n7526 = ~n7516 & ~n7525;
  assign n7527 = controllable_BtoS_ACK7 & ~n7526;
  assign n7528 = n6664 & ~n7513;
  assign n7529 = i_StoB_REQ6 & ~n7304;
  assign n7530 = n6665 & ~n7509;
  assign n7531 = ~n7497 & ~n7530;
  assign n7532 = ~i_StoB_REQ6 & ~n7531;
  assign n7533 = ~n7529 & ~n7532;
  assign n7534 = controllable_BtoS_ACK6 & ~n7533;
  assign n7535 = ~controllable_BtoS_ACK6 & ~n7509;
  assign n7536 = ~n7534 & ~n7535;
  assign n7537 = ~n6664 & ~n7536;
  assign n7538 = ~n7528 & ~n7537;
  assign n7539 = ~controllable_BtoS_ACK7 & ~n7538;
  assign n7540 = ~n7527 & ~n7539;
  assign n7541 = n6663 & ~n7540;
  assign n7542 = ~n6842 & ~n7523;
  assign n7543 = controllable_BtoS_ACK7 & ~n7542;
  assign n7544 = ~controllable_BtoS_ACK7 & ~n7522;
  assign n7545 = ~n7543 & ~n7544;
  assign n7546 = ~n6663 & ~n7545;
  assign n7547 = ~n7541 & ~n7546;
  assign n7548 = ~i_StoB_REQ8 & ~n7547;
  assign n7549 = ~n7384 & ~n7548;
  assign n7550 = controllable_BtoS_ACK8 & ~n7549;
  assign n7551 = ~i_StoB_REQ7 & ~n7536;
  assign n7552 = ~n7517 & ~n7551;
  assign n7553 = n6664 & ~n7552;
  assign n7554 = ~n7525 & ~n7553;
  assign n7555 = controllable_BtoS_ACK7 & ~n7554;
  assign n7556 = ~controllable_BtoS_ACK7 & ~n7536;
  assign n7557 = ~n7555 & ~n7556;
  assign n7558 = ~n6663 & ~n7557;
  assign n7559 = ~n7541 & ~n7558;
  assign n7560 = ~controllable_BtoS_ACK8 & ~n7559;
  assign n7561 = ~n7550 & ~n7560;
  assign n7562 = n6662 & ~n7561;
  assign n7563 = ~i_StoB_REQ8 & ~n7545;
  assign n7564 = ~n7121 & ~n7563;
  assign n7565 = controllable_BtoS_ACK8 & ~n7564;
  assign n7566 = ~controllable_BtoS_ACK8 & ~n7545;
  assign n7567 = ~n7565 & ~n7566;
  assign n7568 = ~n6662 & ~n7567;
  assign n7569 = ~n7562 & ~n7568;
  assign n7570 = ~i_StoB_REQ10 & ~n7569;
  assign n7571 = ~n7383 & ~n7570;
  assign n7572 = controllable_BtoS_ACK10 & ~n7571;
  assign n7573 = i_StoB_REQ8 & ~n7337;
  assign n7574 = n6663 & ~n7557;
  assign n7575 = ~n7546 & ~n7574;
  assign n7576 = ~i_StoB_REQ8 & ~n7575;
  assign n7577 = ~n7573 & ~n7576;
  assign n7578 = controllable_BtoS_ACK8 & ~n7577;
  assign n7579 = ~controllable_BtoS_ACK8 & ~n7557;
  assign n7580 = ~n7578 & ~n7579;
  assign n7581 = ~n6662 & ~n7580;
  assign n7582 = ~n7562 & ~n7581;
  assign n7583 = ~controllable_BtoS_ACK10 & ~n7582;
  assign n7584 = ~n7572 & ~n7583;
  assign n7585 = ~controllable_BtoS_ACK11 & ~n7584;
  assign n7586 = ~n7382 & ~n7585;
  assign n7587 = n6661 & ~n7586;
  assign n7588 = controllable_BtoS_ACK11 & ~n7367;
  assign n7589 = i_StoB_REQ10 & ~n7353;
  assign n7590 = n6662 & ~n7580;
  assign n7591 = ~n7568 & ~n7590;
  assign n7592 = ~i_StoB_REQ10 & ~n7591;
  assign n7593 = ~n7589 & ~n7592;
  assign n7594 = controllable_BtoS_ACK10 & ~n7593;
  assign n7595 = ~controllable_BtoS_ACK10 & ~n7580;
  assign n7596 = ~n7594 & ~n7595;
  assign n7597 = ~controllable_BtoS_ACK11 & ~n7596;
  assign n7598 = ~n7588 & ~n7597;
  assign n7599 = ~n6661 & ~n7598;
  assign n7600 = ~n7587 & ~n7599;
  assign n7601 = i_StoB_REQ11 & ~n7600;
  assign n7602 = n6661 & ~n7584;
  assign n7603 = ~i_StoB_REQ10 & ~n7567;
  assign n7604 = ~n7149 & ~n7603;
  assign n7605 = controllable_BtoS_ACK10 & ~n7604;
  assign n7606 = ~controllable_BtoS_ACK10 & ~n7567;
  assign n7607 = ~n7605 & ~n7606;
  assign n7608 = controllable_BtoS_ACK11 & ~n7607;
  assign n7609 = ~n7597 & ~n7608;
  assign n7610 = ~n6661 & ~n7609;
  assign n7611 = ~n7602 & ~n7610;
  assign n7612 = ~i_StoB_REQ11 & ~n7611;
  assign n7613 = ~n7601 & ~n7612;
  assign n7614 = controllable_ENQ & ~n7613;
  assign n7615 = ~controllable_ENQ & ~n7171;
  assign n7616 = ~n7614 & ~n7615;
  assign n7617 = ~i_StoB_REQ9 & ~n7616;
  assign n7618 = ~n7381 & ~n7617;
  assign n7619 = controllable_BtoS_ACK9 & ~n7618;
  assign n7620 = ~controllable_ENQ & ~n7191;
  assign n7621 = ~n7614 & ~n7620;
  assign n7622 = i_StoB_REQ9 & ~n7621;
  assign n7623 = ~n7617 & ~n7622;
  assign n7624 = ~controllable_BtoS_ACK9 & ~n7623;
  assign n7625 = ~n7619 & ~n7624;
  assign n7626 = controllable_DEQ & ~n7625;
  assign n7627 = i_StoB_REQ9 & ~n7378;
  assign n7628 = ~i_StoB_REQ9 & ~n7613;
  assign n7629 = ~n7627 & ~n7628;
  assign n7630 = controllable_BtoS_ACK9 & ~n7629;
  assign n7631 = ~controllable_BtoS_ACK9 & ~n7613;
  assign n7632 = ~n7630 & ~n7631;
  assign n7633 = ~controllable_DEQ & ~n7632;
  assign n7634 = ~n7626 & ~n7633;
  assign n7635 = i_nEMPTY & ~n7634;
  assign n7636 = ~controllable_ENQ & ~n7615;
  assign n7637 = ~i_StoB_REQ9 & ~n7636;
  assign n7638 = ~i_StoB_REQ9 & ~n7637;
  assign n7639 = controllable_BtoS_ACK9 & ~n7638;
  assign n7640 = ~controllable_ENQ & ~n7620;
  assign n7641 = i_StoB_REQ9 & ~n7640;
  assign n7642 = ~n7637 & ~n7641;
  assign n7643 = ~controllable_BtoS_ACK9 & ~n7642;
  assign n7644 = ~n7639 & ~n7643;
  assign n7645 = controllable_DEQ & ~n7644;
  assign n7646 = controllable_ENQ & ~n7614;
  assign n7647 = ~i_StoB_REQ9 & ~n7646;
  assign n7648 = ~n7381 & ~n7647;
  assign n7649 = controllable_BtoS_ACK9 & ~n7648;
  assign n7650 = ~controllable_BtoS_ACK9 & ~n7646;
  assign n7651 = ~n7649 & ~n7650;
  assign n7652 = ~controllable_DEQ & ~n7651;
  assign n7653 = ~n7645 & ~n7652;
  assign n7654 = ~i_nEMPTY & ~n7653;
  assign n7655 = ~n7635 & ~n7654;
  assign n7656 = i_FULL & ~n7655;
  assign n7657 = ~n6681 & ~n7399;
  assign n7658 = controllable_BtoS_ACK1 & ~n7657;
  assign n7659 = ~n6684 & ~n7658;
  assign n7660 = ~n6671 & ~n7659;
  assign n7661 = ~n7392 & ~n7660;
  assign n7662 = n6670 & ~n7661;
  assign n7663 = ~n6691 & ~n7396;
  assign n7664 = n6671 & ~n7663;
  assign n7665 = ~n6695 & ~n7400;
  assign n7666 = ~n6671 & ~n7665;
  assign n7667 = ~n7664 & ~n7666;
  assign n7668 = ~n6670 & ~n7667;
  assign n7669 = ~n7662 & ~n7668;
  assign n7670 = n6669 & ~n7669;
  assign n7671 = ~n7407 & ~n7670;
  assign n7672 = ~i_StoB_REQ2 & ~n7671;
  assign n7673 = ~n7390 & ~n7672;
  assign n7674 = controllable_BtoS_ACK2 & ~n7673;
  assign n7675 = ~n6673 & ~n7399;
  assign n7676 = controllable_BtoS_ACK1 & ~n7675;
  assign n7677 = ~n6676 & ~n7676;
  assign n7678 = ~n6671 & ~n7677;
  assign n7679 = ~n6678 & ~n7678;
  assign n7680 = n6670 & ~n7679;
  assign n7681 = ~n6676 & ~n7396;
  assign n7682 = n6671 & ~n7681;
  assign n7683 = ~n6676 & ~n7400;
  assign n7684 = ~n6671 & ~n7683;
  assign n7685 = ~n7682 & ~n7684;
  assign n7686 = ~n6670 & ~n7685;
  assign n7687 = ~n7680 & ~n7686;
  assign n7688 = ~n6669 & ~n7687;
  assign n7689 = ~n7670 & ~n7688;
  assign n7690 = i_StoB_REQ2 & ~n7689;
  assign n7691 = ~n6671 & ~n7660;
  assign n7692 = n6670 & ~n7691;
  assign n7693 = ~n7668 & ~n7692;
  assign n7694 = ~n6669 & ~n7693;
  assign n7695 = ~n7670 & ~n7694;
  assign n7696 = ~i_StoB_REQ2 & ~n7695;
  assign n7697 = ~n7690 & ~n7696;
  assign n7698 = ~controllable_BtoS_ACK2 & ~n7697;
  assign n7699 = ~n7674 & ~n7698;
  assign n7700 = n6668 & ~n7699;
  assign n7701 = ~n7425 & ~n7700;
  assign n7702 = ~i_StoB_REQ3 & ~n7701;
  assign n7703 = ~n7389 & ~n7702;
  assign n7704 = controllable_BtoS_ACK3 & ~n7703;
  assign n7705 = n6669 & ~n7687;
  assign n7706 = ~n7407 & ~n7705;
  assign n7707 = ~i_StoB_REQ2 & ~n7706;
  assign n7708 = ~n7430 & ~n7707;
  assign n7709 = controllable_BtoS_ACK2 & ~n7708;
  assign n7710 = ~controllable_BtoS_ACK2 & ~n7687;
  assign n7711 = ~n7709 & ~n7710;
  assign n7712 = ~n6668 & ~n7711;
  assign n7713 = ~n7700 & ~n7712;
  assign n7714 = i_StoB_REQ3 & ~n7713;
  assign n7715 = n6669 & ~n7693;
  assign n7716 = ~n7407 & ~n7715;
  assign n7717 = ~i_StoB_REQ2 & ~n7716;
  assign n7718 = ~n7430 & ~n7717;
  assign n7719 = controllable_BtoS_ACK2 & ~n7718;
  assign n7720 = ~n7688 & ~n7715;
  assign n7721 = i_StoB_REQ2 & ~n7720;
  assign n7722 = ~i_StoB_REQ2 & ~n7693;
  assign n7723 = ~n7721 & ~n7722;
  assign n7724 = ~controllable_BtoS_ACK2 & ~n7723;
  assign n7725 = ~n7719 & ~n7724;
  assign n7726 = ~n6668 & ~n7725;
  assign n7727 = ~n7700 & ~n7726;
  assign n7728 = ~i_StoB_REQ3 & ~n7727;
  assign n7729 = ~n7714 & ~n7728;
  assign n7730 = ~controllable_BtoS_ACK3 & ~n7729;
  assign n7731 = ~n7704 & ~n7730;
  assign n7732 = ~controllable_BtoS_ACK4 & ~n7731;
  assign n7733 = ~n7388 & ~n7732;
  assign n7734 = n6667 & ~n7733;
  assign n7735 = n6668 & ~n7711;
  assign n7736 = ~n7425 & ~n7735;
  assign n7737 = ~i_StoB_REQ3 & ~n7736;
  assign n7738 = ~n7446 & ~n7737;
  assign n7739 = controllable_BtoS_ACK3 & ~n7738;
  assign n7740 = ~controllable_BtoS_ACK3 & ~n7711;
  assign n7741 = ~n7739 & ~n7740;
  assign n7742 = ~controllable_BtoS_ACK4 & ~n7741;
  assign n7743 = ~n7445 & ~n7742;
  assign n7744 = ~n6667 & ~n7743;
  assign n7745 = ~n7734 & ~n7744;
  assign n7746 = i_StoB_REQ4 & ~n7745;
  assign n7747 = n6667 & ~n7731;
  assign n7748 = n6668 & ~n7725;
  assign n7749 = ~n7425 & ~n7748;
  assign n7750 = ~i_StoB_REQ3 & ~n7749;
  assign n7751 = ~n7446 & ~n7750;
  assign n7752 = controllable_BtoS_ACK3 & ~n7751;
  assign n7753 = ~n7712 & ~n7748;
  assign n7754 = i_StoB_REQ3 & ~n7753;
  assign n7755 = ~i_StoB_REQ3 & ~n7725;
  assign n7756 = ~n7754 & ~n7755;
  assign n7757 = ~controllable_BtoS_ACK3 & ~n7756;
  assign n7758 = ~n7752 & ~n7757;
  assign n7759 = ~controllable_BtoS_ACK4 & ~n7758;
  assign n7760 = ~n7465 & ~n7759;
  assign n7761 = ~n6667 & ~n7760;
  assign n7762 = ~n7747 & ~n7761;
  assign n7763 = ~i_StoB_REQ4 & ~n7762;
  assign n7764 = ~n7746 & ~n7763;
  assign n7765 = n6666 & ~n7764;
  assign n7766 = ~n7477 & ~n7765;
  assign n7767 = ~i_StoB_REQ5 & ~n7766;
  assign n7768 = ~n7387 & ~n7767;
  assign n7769 = controllable_BtoS_ACK5 & ~n7768;
  assign n7770 = i_StoB_REQ4 & ~n7743;
  assign n7771 = n6667 & ~n7741;
  assign n7772 = ~n7465 & ~n7742;
  assign n7773 = ~n6667 & ~n7772;
  assign n7774 = ~n7771 & ~n7773;
  assign n7775 = ~i_StoB_REQ4 & ~n7774;
  assign n7776 = ~n7770 & ~n7775;
  assign n7777 = ~n6666 & ~n7776;
  assign n7778 = ~n7765 & ~n7777;
  assign n7779 = i_StoB_REQ5 & ~n7778;
  assign n7780 = ~n7445 & ~n7759;
  assign n7781 = n6667 & ~n7780;
  assign n7782 = ~n7744 & ~n7781;
  assign n7783 = i_StoB_REQ4 & ~n7782;
  assign n7784 = n6667 & ~n7758;
  assign n7785 = ~n7761 & ~n7784;
  assign n7786 = ~i_StoB_REQ4 & ~n7785;
  assign n7787 = ~n7783 & ~n7786;
  assign n7788 = ~n6666 & ~n7787;
  assign n7789 = ~n7765 & ~n7788;
  assign n7790 = ~i_StoB_REQ5 & ~n7789;
  assign n7791 = ~n7779 & ~n7790;
  assign n7792 = ~controllable_BtoS_ACK5 & ~n7791;
  assign n7793 = ~n7769 & ~n7792;
  assign n7794 = n6665 & ~n7793;
  assign n7795 = ~n7497 & ~n7794;
  assign n7796 = ~i_StoB_REQ6 & ~n7795;
  assign n7797 = ~n7386 & ~n7796;
  assign n7798 = controllable_BtoS_ACK6 & ~n7797;
  assign n7799 = n6666 & ~n7776;
  assign n7800 = ~n7477 & ~n7799;
  assign n7801 = ~i_StoB_REQ5 & ~n7800;
  assign n7802 = ~n7502 & ~n7801;
  assign n7803 = controllable_BtoS_ACK5 & ~n7802;
  assign n7804 = ~controllable_BtoS_ACK5 & ~n7776;
  assign n7805 = ~n7803 & ~n7804;
  assign n7806 = ~n6665 & ~n7805;
  assign n7807 = ~n7794 & ~n7806;
  assign n7808 = i_StoB_REQ6 & ~n7807;
  assign n7809 = n6666 & ~n7787;
  assign n7810 = ~n7477 & ~n7809;
  assign n7811 = ~i_StoB_REQ5 & ~n7810;
  assign n7812 = ~n7502 & ~n7811;
  assign n7813 = controllable_BtoS_ACK5 & ~n7812;
  assign n7814 = ~n7777 & ~n7809;
  assign n7815 = i_StoB_REQ5 & ~n7814;
  assign n7816 = ~i_StoB_REQ5 & ~n7787;
  assign n7817 = ~n7815 & ~n7816;
  assign n7818 = ~controllable_BtoS_ACK5 & ~n7817;
  assign n7819 = ~n7813 & ~n7818;
  assign n7820 = ~n6665 & ~n7819;
  assign n7821 = ~n7794 & ~n7820;
  assign n7822 = ~i_StoB_REQ6 & ~n7821;
  assign n7823 = ~n7808 & ~n7822;
  assign n7824 = ~controllable_BtoS_ACK6 & ~n7823;
  assign n7825 = ~n7798 & ~n7824;
  assign n7826 = ~i_StoB_REQ7 & ~n7825;
  assign n7827 = ~n7385 & ~n7826;
  assign n7828 = n6664 & ~n7827;
  assign n7829 = ~n7525 & ~n7828;
  assign n7830 = controllable_BtoS_ACK7 & ~n7829;
  assign n7831 = n6664 & ~n7825;
  assign n7832 = n6665 & ~n7805;
  assign n7833 = ~n7497 & ~n7832;
  assign n7834 = ~i_StoB_REQ6 & ~n7833;
  assign n7835 = ~n7529 & ~n7834;
  assign n7836 = controllable_BtoS_ACK6 & ~n7835;
  assign n7837 = ~controllable_BtoS_ACK6 & ~n7805;
  assign n7838 = ~n7836 & ~n7837;
  assign n7839 = i_StoB_REQ7 & ~n7838;
  assign n7840 = n6665 & ~n7819;
  assign n7841 = ~n7497 & ~n7840;
  assign n7842 = ~i_StoB_REQ6 & ~n7841;
  assign n7843 = ~n7529 & ~n7842;
  assign n7844 = controllable_BtoS_ACK6 & ~n7843;
  assign n7845 = ~n7806 & ~n7840;
  assign n7846 = i_StoB_REQ6 & ~n7845;
  assign n7847 = ~i_StoB_REQ6 & ~n7819;
  assign n7848 = ~n7846 & ~n7847;
  assign n7849 = ~controllable_BtoS_ACK6 & ~n7848;
  assign n7850 = ~n7844 & ~n7849;
  assign n7851 = ~i_StoB_REQ7 & ~n7850;
  assign n7852 = ~n7839 & ~n7851;
  assign n7853 = ~n6664 & ~n7852;
  assign n7854 = ~n7831 & ~n7853;
  assign n7855 = ~controllable_BtoS_ACK7 & ~n7854;
  assign n7856 = ~n7830 & ~n7855;
  assign n7857 = n6663 & ~n7856;
  assign n7858 = ~n7546 & ~n7857;
  assign n7859 = ~i_StoB_REQ8 & ~n7858;
  assign n7860 = ~n7384 & ~n7859;
  assign n7861 = controllable_BtoS_ACK8 & ~n7860;
  assign n7862 = ~i_StoB_REQ7 & ~n7838;
  assign n7863 = ~n7517 & ~n7862;
  assign n7864 = n6664 & ~n7863;
  assign n7865 = ~n7525 & ~n7864;
  assign n7866 = controllable_BtoS_ACK7 & ~n7865;
  assign n7867 = ~controllable_BtoS_ACK7 & ~n7838;
  assign n7868 = ~n7866 & ~n7867;
  assign n7869 = ~n6663 & ~n7868;
  assign n7870 = ~n7857 & ~n7869;
  assign n7871 = i_StoB_REQ8 & ~n7870;
  assign n7872 = ~n7517 & ~n7851;
  assign n7873 = n6664 & ~n7872;
  assign n7874 = ~n7525 & ~n7873;
  assign n7875 = controllable_BtoS_ACK7 & ~n7874;
  assign n7876 = n6664 & ~n7850;
  assign n7877 = ~n7853 & ~n7876;
  assign n7878 = ~controllable_BtoS_ACK7 & ~n7877;
  assign n7879 = ~n7875 & ~n7878;
  assign n7880 = ~n6663 & ~n7879;
  assign n7881 = ~n7857 & ~n7880;
  assign n7882 = ~i_StoB_REQ8 & ~n7881;
  assign n7883 = ~n7871 & ~n7882;
  assign n7884 = ~controllable_BtoS_ACK8 & ~n7883;
  assign n7885 = ~n7861 & ~n7884;
  assign n7886 = n6662 & ~n7885;
  assign n7887 = ~n7568 & ~n7886;
  assign n7888 = ~i_StoB_REQ10 & ~n7887;
  assign n7889 = ~n7383 & ~n7888;
  assign n7890 = controllable_BtoS_ACK10 & ~n7889;
  assign n7891 = n6663 & ~n7868;
  assign n7892 = ~n7546 & ~n7891;
  assign n7893 = ~i_StoB_REQ8 & ~n7892;
  assign n7894 = ~n7573 & ~n7893;
  assign n7895 = controllable_BtoS_ACK8 & ~n7894;
  assign n7896 = ~controllable_BtoS_ACK8 & ~n7868;
  assign n7897 = ~n7895 & ~n7896;
  assign n7898 = ~n6662 & ~n7897;
  assign n7899 = ~n7886 & ~n7898;
  assign n7900 = i_StoB_REQ10 & ~n7899;
  assign n7901 = n6663 & ~n7879;
  assign n7902 = ~n7546 & ~n7901;
  assign n7903 = ~i_StoB_REQ8 & ~n7902;
  assign n7904 = ~n7573 & ~n7903;
  assign n7905 = controllable_BtoS_ACK8 & ~n7904;
  assign n7906 = ~n7869 & ~n7901;
  assign n7907 = i_StoB_REQ8 & ~n7906;
  assign n7908 = ~i_StoB_REQ8 & ~n7879;
  assign n7909 = ~n7907 & ~n7908;
  assign n7910 = ~controllable_BtoS_ACK8 & ~n7909;
  assign n7911 = ~n7905 & ~n7910;
  assign n7912 = ~n6662 & ~n7911;
  assign n7913 = ~n7886 & ~n7912;
  assign n7914 = ~i_StoB_REQ10 & ~n7913;
  assign n7915 = ~n7900 & ~n7914;
  assign n7916 = ~controllable_BtoS_ACK10 & ~n7915;
  assign n7917 = ~n7890 & ~n7916;
  assign n7918 = ~controllable_BtoS_ACK11 & ~n7917;
  assign n7919 = ~n7382 & ~n7918;
  assign n7920 = n6661 & ~n7919;
  assign n7921 = n6662 & ~n7897;
  assign n7922 = ~n7568 & ~n7921;
  assign n7923 = ~i_StoB_REQ10 & ~n7922;
  assign n7924 = ~n7589 & ~n7923;
  assign n7925 = controllable_BtoS_ACK10 & ~n7924;
  assign n7926 = ~controllable_BtoS_ACK10 & ~n7897;
  assign n7927 = ~n7925 & ~n7926;
  assign n7928 = ~controllable_BtoS_ACK11 & ~n7927;
  assign n7929 = ~n7588 & ~n7928;
  assign n7930 = ~n6661 & ~n7929;
  assign n7931 = ~n7920 & ~n7930;
  assign n7932 = i_StoB_REQ11 & ~n7931;
  assign n7933 = n6661 & ~n7917;
  assign n7934 = n6662 & ~n7911;
  assign n7935 = ~n7568 & ~n7934;
  assign n7936 = ~i_StoB_REQ10 & ~n7935;
  assign n7937 = ~n7589 & ~n7936;
  assign n7938 = controllable_BtoS_ACK10 & ~n7937;
  assign n7939 = ~n7898 & ~n7934;
  assign n7940 = i_StoB_REQ10 & ~n7939;
  assign n7941 = ~i_StoB_REQ10 & ~n7911;
  assign n7942 = ~n7940 & ~n7941;
  assign n7943 = ~controllable_BtoS_ACK10 & ~n7942;
  assign n7944 = ~n7938 & ~n7943;
  assign n7945 = ~controllable_BtoS_ACK11 & ~n7944;
  assign n7946 = ~n7608 & ~n7945;
  assign n7947 = ~n6661 & ~n7946;
  assign n7948 = ~n7933 & ~n7947;
  assign n7949 = ~i_StoB_REQ11 & ~n7948;
  assign n7950 = ~n7932 & ~n7949;
  assign n7951 = controllable_ENQ & ~n7950;
  assign n7952 = ~n7615 & ~n7951;
  assign n7953 = ~i_StoB_REQ9 & ~n7952;
  assign n7954 = ~n7381 & ~n7953;
  assign n7955 = controllable_BtoS_ACK9 & ~n7954;
  assign n7956 = ~n7620 & ~n7951;
  assign n7957 = i_StoB_REQ9 & ~n7956;
  assign n7958 = ~n7953 & ~n7957;
  assign n7959 = ~controllable_BtoS_ACK9 & ~n7958;
  assign n7960 = ~n7955 & ~n7959;
  assign n7961 = controllable_DEQ & ~n7960;
  assign n7962 = ~controllable_ENQ & ~n7950;
  assign n7963 = ~n7614 & ~n7962;
  assign n7964 = ~i_StoB_REQ9 & ~n7963;
  assign n7965 = ~n7627 & ~n7964;
  assign n7966 = controllable_BtoS_ACK9 & ~n7965;
  assign n7967 = ~controllable_BtoS_ACK9 & ~n7963;
  assign n7968 = ~n7966 & ~n7967;
  assign n7969 = ~controllable_DEQ & ~n7968;
  assign n7970 = ~n7961 & ~n7969;
  assign n7971 = i_nEMPTY & ~n7970;
  assign n7972 = controllable_DEQ & ~n7205;
  assign n7973 = ~controllable_DEQ & ~n7625;
  assign n7974 = ~n7972 & ~n7973;
  assign n7975 = ~i_nEMPTY & ~n7974;
  assign n7976 = ~n7971 & ~n7975;
  assign n7977 = ~i_FULL & ~n7976;
  assign n7978 = ~n7656 & ~n7977;
  assign n7979 = ~i_RtoB_ACK0 & ~n7978;
  assign n7980 = ~n7213 & ~n7979;
  assign n7981 = n6660 & ~n7980;
  assign n7982 = i_StoB_REQ11 & ~n6920;
  assign n7983 = ~i_StoB_REQ11 & ~n7152;
  assign n7984 = ~n7982 & ~n7983;
  assign n7985 = controllable_ENQ & ~n7984;
  assign n7986 = controllable_ENQ & ~n7985;
  assign n7987 = ~i_StoB_REQ9 & ~n7986;
  assign n7988 = ~i_StoB_REQ9 & ~n7987;
  assign n7989 = controllable_BtoS_ACK9 & ~n7988;
  assign n7990 = ~i_StoB_REQ11 & ~n6918;
  assign n7991 = ~n7982 & ~n7990;
  assign n7992 = controllable_ENQ & ~n7991;
  assign n7993 = controllable_ENQ & ~n7992;
  assign n7994 = i_StoB_REQ9 & ~n7993;
  assign n7995 = ~controllable_BtoS_ACK11 & ~n7186;
  assign n7996 = n6661 & ~n7995;
  assign n7997 = ~n6921 & ~n7996;
  assign n7998 = i_StoB_REQ11 & ~n7997;
  assign n7999 = n6661 & ~n7165;
  assign n8000 = ~n7168 & ~n7999;
  assign n8001 = ~i_StoB_REQ11 & ~n8000;
  assign n8002 = ~n7998 & ~n8001;
  assign n8003 = controllable_ENQ & ~n8002;
  assign n8004 = controllable_ENQ & ~n8003;
  assign n8005 = ~i_StoB_REQ9 & ~n8004;
  assign n8006 = ~n7994 & ~n8005;
  assign n8007 = ~controllable_BtoS_ACK9 & ~n8006;
  assign n8008 = ~n7989 & ~n8007;
  assign n8009 = controllable_DEQ & ~n8008;
  assign n8010 = ~i_StoB_REQ9 & ~n7984;
  assign n8011 = ~i_StoB_REQ9 & ~n8010;
  assign n8012 = controllable_BtoS_ACK9 & ~n8011;
  assign n8013 = i_StoB_REQ9 & ~n7991;
  assign n8014 = ~i_StoB_REQ9 & ~n8002;
  assign n8015 = ~n8013 & ~n8014;
  assign n8016 = ~controllable_BtoS_ACK9 & ~n8015;
  assign n8017 = ~n8012 & ~n8016;
  assign n8018 = ~controllable_DEQ & ~n8017;
  assign n8019 = ~n8009 & ~n8018;
  assign n8020 = i_nEMPTY & ~n8019;
  assign n8021 = ~controllable_DEQ & ~n8008;
  assign n8022 = ~controllable_DEQ & ~n8021;
  assign n8023 = ~i_nEMPTY & ~n8022;
  assign n8024 = ~n8020 & ~n8023;
  assign n8025 = i_RtoB_ACK0 & ~n8024;
  assign n8026 = i_StoB_REQ11 & ~n7369;
  assign n8027 = n6661 & ~n7367;
  assign n8028 = ~n7375 & ~n8027;
  assign n8029 = ~i_StoB_REQ11 & ~n8028;
  assign n8030 = ~n8026 & ~n8029;
  assign n8031 = controllable_ENQ & ~n8030;
  assign n8032 = controllable_ENQ & ~n8031;
  assign n8033 = i_StoB_REQ9 & ~n8032;
  assign n8034 = ~controllable_BtoS_ACK11 & ~n7607;
  assign n8035 = ~n7178 & ~n8034;
  assign n8036 = i_StoB_REQ11 & ~n8035;
  assign n8037 = ~i_StoB_REQ11 & ~n7607;
  assign n8038 = ~n8036 & ~n8037;
  assign n8039 = controllable_ENQ & ~n8038;
  assign n8040 = ~controllable_ENQ & ~n7984;
  assign n8041 = ~n8039 & ~n8040;
  assign n8042 = ~i_StoB_REQ9 & ~n8041;
  assign n8043 = ~n8033 & ~n8042;
  assign n8044 = controllable_BtoS_ACK9 & ~n8043;
  assign n8045 = i_StoB_REQ11 & ~n7598;
  assign n8046 = n6661 & ~n7596;
  assign n8047 = ~n7610 & ~n8046;
  assign n8048 = ~i_StoB_REQ11 & ~n8047;
  assign n8049 = ~n8045 & ~n8048;
  assign n8050 = controllable_ENQ & ~n8049;
  assign n8051 = ~controllable_ENQ & ~n7991;
  assign n8052 = ~n8050 & ~n8051;
  assign n8053 = i_StoB_REQ9 & ~n8052;
  assign n8054 = ~controllable_ENQ & ~n8002;
  assign n8055 = ~n8050 & ~n8054;
  assign n8056 = ~i_StoB_REQ9 & ~n8055;
  assign n8057 = ~n8053 & ~n8056;
  assign n8058 = ~controllable_BtoS_ACK9 & ~n8057;
  assign n8059 = ~n8044 & ~n8058;
  assign n8060 = controllable_DEQ & ~n8059;
  assign n8061 = i_StoB_REQ9 & ~n8030;
  assign n8062 = ~i_StoB_REQ9 & ~n8038;
  assign n8063 = ~n8061 & ~n8062;
  assign n8064 = controllable_BtoS_ACK9 & ~n8063;
  assign n8065 = ~controllable_BtoS_ACK9 & ~n8049;
  assign n8066 = ~n8064 & ~n8065;
  assign n8067 = ~controllable_DEQ & ~n8066;
  assign n8068 = ~n8060 & ~n8067;
  assign n8069 = i_nEMPTY & ~n8068;
  assign n8070 = ~controllable_ENQ & ~n8040;
  assign n8071 = ~i_StoB_REQ9 & ~n8070;
  assign n8072 = ~i_StoB_REQ9 & ~n8071;
  assign n8073 = controllable_BtoS_ACK9 & ~n8072;
  assign n8074 = ~controllable_ENQ & ~n8051;
  assign n8075 = i_StoB_REQ9 & ~n8074;
  assign n8076 = ~controllable_ENQ & ~n8054;
  assign n8077 = ~i_StoB_REQ9 & ~n8076;
  assign n8078 = ~n8075 & ~n8077;
  assign n8079 = ~controllable_BtoS_ACK9 & ~n8078;
  assign n8080 = ~n8073 & ~n8079;
  assign n8081 = controllable_DEQ & ~n8080;
  assign n8082 = controllable_ENQ & ~n8039;
  assign n8083 = ~i_StoB_REQ9 & ~n8082;
  assign n8084 = ~n8033 & ~n8083;
  assign n8085 = controllable_BtoS_ACK9 & ~n8084;
  assign n8086 = controllable_ENQ & ~n8050;
  assign n8087 = ~controllable_BtoS_ACK9 & ~n8086;
  assign n8088 = ~n8085 & ~n8087;
  assign n8089 = ~controllable_DEQ & ~n8088;
  assign n8090 = ~n8081 & ~n8089;
  assign n8091 = ~i_nEMPTY & ~n8090;
  assign n8092 = ~n8069 & ~n8091;
  assign n8093 = i_FULL & ~n8092;
  assign n8094 = i_StoB_REQ11 & ~n7929;
  assign n8095 = n6661 & ~n7927;
  assign n8096 = ~n7608 & ~n7928;
  assign n8097 = ~n6661 & ~n8096;
  assign n8098 = ~n8095 & ~n8097;
  assign n8099 = ~i_StoB_REQ11 & ~n8098;
  assign n8100 = ~n8094 & ~n8099;
  assign n8101 = controllable_ENQ & ~n8100;
  assign n8102 = ~n8051 & ~n8101;
  assign n8103 = i_StoB_REQ9 & ~n8102;
  assign n8104 = ~n7588 & ~n7945;
  assign n8105 = n6661 & ~n8104;
  assign n8106 = ~n7930 & ~n8105;
  assign n8107 = i_StoB_REQ11 & ~n8106;
  assign n8108 = n6661 & ~n7944;
  assign n8109 = ~n7947 & ~n8108;
  assign n8110 = ~i_StoB_REQ11 & ~n8109;
  assign n8111 = ~n8107 & ~n8110;
  assign n8112 = controllable_ENQ & ~n8111;
  assign n8113 = ~n8054 & ~n8112;
  assign n8114 = ~i_StoB_REQ9 & ~n8113;
  assign n8115 = ~n8103 & ~n8114;
  assign n8116 = ~controllable_BtoS_ACK9 & ~n8115;
  assign n8117 = ~n8044 & ~n8116;
  assign n8118 = controllable_DEQ & ~n8117;
  assign n8119 = ~controllable_ENQ & ~n8100;
  assign n8120 = ~n8050 & ~n8119;
  assign n8121 = i_StoB_REQ9 & ~n8120;
  assign n8122 = ~controllable_ENQ & ~n8111;
  assign n8123 = ~n8050 & ~n8122;
  assign n8124 = ~i_StoB_REQ9 & ~n8123;
  assign n8125 = ~n8121 & ~n8124;
  assign n8126 = ~controllable_BtoS_ACK9 & ~n8125;
  assign n8127 = ~n8064 & ~n8126;
  assign n8128 = ~controllable_DEQ & ~n8127;
  assign n8129 = ~n8118 & ~n8128;
  assign n8130 = i_nEMPTY & ~n8129;
  assign n8131 = controllable_DEQ & ~n8017;
  assign n8132 = ~controllable_DEQ & ~n8059;
  assign n8133 = ~n8131 & ~n8132;
  assign n8134 = ~i_nEMPTY & ~n8133;
  assign n8135 = ~n8130 & ~n8134;
  assign n8136 = ~i_FULL & ~n8135;
  assign n8137 = ~n8093 & ~n8136;
  assign n8138 = ~i_RtoB_ACK0 & ~n8137;
  assign n8139 = ~n8025 & ~n8138;
  assign n8140 = ~n6660 & ~n8139;
  assign n8141 = ~n7981 & ~n8140;
  assign n8142 = ~n6659 & ~n8141;
  assign n8143 = n6490 & n6654;
  assign n8144 = ~n6490 & n6655;
  assign n8145 = ~n8143 & ~n8144;
  assign n8146 = n75 & reg_stateG7_0_out;
  assign n8147 = ~n6483 & ~n6490;
  assign n8148 = ~n8146 & ~n8147;
  assign n8149 = n8145 & ~n8148;
  assign n8150 = ~n8141 & ~n8149;
  assign n8151 = ~n8149 & ~n8150;
  assign n8152 = n6659 & ~n8151;
  assign n8153 = ~n8142 & ~n8152;
  assign n8154 = n6652 & ~n8153;
  assign n8155 = n6661 & ~n8035;
  assign n8156 = ~n6671 & ~n6677;
  assign n8157 = ~n6931 & ~n8156;
  assign n8158 = n6670 & ~n8157;
  assign n8159 = ~n6670 & ~n6677;
  assign n8160 = ~n8158 & ~n8159;
  assign n8161 = n6669 & ~n8160;
  assign n8162 = ~n6702 & ~n8161;
  assign n8163 = ~i_StoB_REQ2 & ~n8162;
  assign n8164 = ~i_StoB_REQ2 & ~n8163;
  assign n8165 = controllable_BtoS_ACK2 & ~n8164;
  assign n8166 = ~n6964 & ~n8163;
  assign n8167 = ~controllable_BtoS_ACK2 & ~n8166;
  assign n8168 = ~n8165 & ~n8167;
  assign n8169 = n6668 & ~n8168;
  assign n8170 = ~n6723 & ~n8169;
  assign n8171 = ~i_StoB_REQ3 & ~n8170;
  assign n8172 = ~i_StoB_REQ3 & ~n8171;
  assign n8173 = controllable_BtoS_ACK3 & ~n8172;
  assign n8174 = ~n6992 & ~n8171;
  assign n8175 = ~controllable_BtoS_ACK3 & ~n8174;
  assign n8176 = ~n8173 & ~n8175;
  assign n8177 = n6667 & ~n8176;
  assign n8178 = ~n6667 & ~n6752;
  assign n8179 = ~n8177 & ~n8178;
  assign n8180 = ~i_StoB_REQ4 & ~n8179;
  assign n8181 = ~n6777 & ~n8180;
  assign n8182 = n6666 & ~n8181;
  assign n8183 = ~n6780 & ~n8182;
  assign n8184 = ~i_StoB_REQ5 & ~n8183;
  assign n8185 = ~i_StoB_REQ5 & ~n8184;
  assign n8186 = controllable_BtoS_ACK5 & ~n8185;
  assign n8187 = ~n7034 & ~n8184;
  assign n8188 = ~controllable_BtoS_ACK5 & ~n8187;
  assign n8189 = ~n8186 & ~n8188;
  assign n8190 = n6665 & ~n8189;
  assign n8191 = ~n6806 & ~n8190;
  assign n8192 = ~i_StoB_REQ6 & ~n8191;
  assign n8193 = ~i_StoB_REQ6 & ~n8192;
  assign n8194 = controllable_BtoS_ACK6 & ~n8193;
  assign n8195 = ~n7064 & ~n8192;
  assign n8196 = ~controllable_BtoS_ACK6 & ~n8195;
  assign n8197 = ~n8194 & ~n8196;
  assign n8198 = ~i_StoB_REQ7 & ~n8197;
  assign n8199 = ~i_StoB_REQ7 & ~n8198;
  assign n8200 = n6664 & ~n8199;
  assign n8201 = ~n6838 & ~n8200;
  assign n8202 = controllable_BtoS_ACK7 & ~n8201;
  assign n8203 = ~n6842 & ~n8198;
  assign n8204 = n6664 & ~n8203;
  assign n8205 = ~n6664 & ~n6835;
  assign n8206 = ~n8204 & ~n8205;
  assign n8207 = ~controllable_BtoS_ACK7 & ~n8206;
  assign n8208 = ~n8202 & ~n8207;
  assign n8209 = n6663 & ~n8208;
  assign n8210 = ~n6863 & ~n8209;
  assign n8211 = ~i_StoB_REQ8 & ~n8210;
  assign n8212 = ~i_StoB_REQ8 & ~n8211;
  assign n8213 = controllable_BtoS_ACK8 & ~n8212;
  assign n8214 = ~n7121 & ~n8211;
  assign n8215 = ~controllable_BtoS_ACK8 & ~n8214;
  assign n8216 = ~n8213 & ~n8215;
  assign n8217 = n6662 & ~n8216;
  assign n8218 = ~n6889 & ~n8217;
  assign n8219 = ~i_StoB_REQ10 & ~n8218;
  assign n8220 = ~i_StoB_REQ10 & ~n8219;
  assign n8221 = controllable_BtoS_ACK10 & ~n8220;
  assign n8222 = ~n7149 & ~n8219;
  assign n8223 = ~controllable_BtoS_ACK10 & ~n8222;
  assign n8224 = ~n8221 & ~n8223;
  assign n8225 = controllable_BtoS_ACK11 & ~n8224;
  assign n8226 = ~n8034 & ~n8225;
  assign n8227 = ~n6661 & ~n8226;
  assign n8228 = ~n8155 & ~n8227;
  assign n8229 = i_StoB_REQ11 & ~n8228;
  assign n8230 = n6662 & ~n6888;
  assign n8231 = ~n6662 & ~n8216;
  assign n8232 = ~n8230 & ~n8231;
  assign n8233 = i_StoB_REQ10 & ~n8232;
  assign n8234 = n6663 & ~n6862;
  assign n8235 = ~n6663 & ~n8208;
  assign n8236 = ~n8234 & ~n8235;
  assign n8237 = i_StoB_REQ8 & ~n8236;
  assign n8238 = n6665 & ~n6805;
  assign n8239 = ~n6665 & ~n8189;
  assign n8240 = ~n8238 & ~n8239;
  assign n8241 = i_StoB_REQ6 & ~n8240;
  assign n8242 = n6666 & ~n6779;
  assign n8243 = ~n6666 & ~n8181;
  assign n8244 = ~n8242 & ~n8243;
  assign n8245 = i_StoB_REQ5 & ~n8244;
  assign n8246 = n6667 & ~n7473;
  assign n8247 = controllable_BtoS_ACK4 & ~n8176;
  assign n8248 = ~n7472 & ~n8247;
  assign n8249 = ~n6667 & ~n8248;
  assign n8250 = ~n8246 & ~n8249;
  assign n8251 = i_StoB_REQ4 & ~n8250;
  assign n8252 = n6668 & ~n6722;
  assign n8253 = ~n6668 & ~n8168;
  assign n8254 = ~n8252 & ~n8253;
  assign n8255 = i_StoB_REQ3 & ~n8254;
  assign n8256 = n6669 & ~n6677;
  assign n8257 = ~n6669 & ~n8160;
  assign n8258 = ~n8256 & ~n8257;
  assign n8259 = i_StoB_REQ2 & ~n8258;
  assign n8260 = controllable_BtoS_ACK1 & n6672;
  assign n8261 = ~i_StoB_REQ1 & ~n6672;
  assign n8262 = ~i_StoB_REQ1 & ~n8261;
  assign n8263 = ~controllable_BtoS_ACK1 & n8262;
  assign n8264 = ~n8260 & ~n8263;
  assign n8265 = ~n6671 & ~n8264;
  assign n8266 = ~n7392 & ~n8265;
  assign n8267 = n6670 & ~n8266;
  assign n8268 = i_StoB_REQ1 & ~n6924;
  assign n8269 = controllable_BtoS_ACK1 & n8268;
  assign n8270 = n6671 & n8269;
  assign n8271 = ~n6671 & n7391;
  assign n8272 = ~n8270 & ~n8271;
  assign n8273 = ~n6670 & ~n8272;
  assign n8274 = ~n8267 & ~n8273;
  assign n8275 = n6669 & ~n8274;
  assign n8276 = ~n7407 & ~n8275;
  assign n8277 = ~i_StoB_REQ2 & ~n8276;
  assign n8278 = ~n8259 & ~n8277;
  assign n8279 = controllable_BtoS_ACK2 & ~n8278;
  assign n8280 = i_StoB_REQ2 & n7391;
  assign n8281 = ~n8277 & ~n8280;
  assign n8282 = ~controllable_BtoS_ACK2 & ~n8281;
  assign n8283 = ~n8279 & ~n8282;
  assign n8284 = n6668 & ~n8283;
  assign n8285 = ~n7425 & ~n8284;
  assign n8286 = ~i_StoB_REQ3 & ~n8285;
  assign n8287 = ~n8255 & ~n8286;
  assign n8288 = controllable_BtoS_ACK3 & ~n8287;
  assign n8289 = i_StoB_REQ3 & ~n7424;
  assign n8290 = ~n8286 & ~n8289;
  assign n8291 = ~controllable_BtoS_ACK3 & ~n8290;
  assign n8292 = ~n8288 & ~n8291;
  assign n8293 = n6667 & ~n8292;
  assign n8294 = ~n6667 & ~n7464;
  assign n8295 = ~n8293 & ~n8294;
  assign n8296 = ~i_StoB_REQ4 & ~n8295;
  assign n8297 = ~n8251 & ~n8296;
  assign n8298 = n6666 & ~n8297;
  assign n8299 = ~n7477 & ~n8298;
  assign n8300 = ~i_StoB_REQ5 & ~n8299;
  assign n8301 = ~n8245 & ~n8300;
  assign n8302 = controllable_BtoS_ACK5 & ~n8301;
  assign n8303 = i_StoB_REQ5 & ~n7476;
  assign n8304 = ~n8300 & ~n8303;
  assign n8305 = ~controllable_BtoS_ACK5 & ~n8304;
  assign n8306 = ~n8302 & ~n8305;
  assign n8307 = n6665 & ~n8306;
  assign n8308 = ~n7497 & ~n8307;
  assign n8309 = ~i_StoB_REQ6 & ~n8308;
  assign n8310 = ~n8241 & ~n8309;
  assign n8311 = controllable_BtoS_ACK6 & ~n8310;
  assign n8312 = i_StoB_REQ6 & ~n7496;
  assign n8313 = ~n8309 & ~n8312;
  assign n8314 = ~controllable_BtoS_ACK6 & ~n8313;
  assign n8315 = ~n8311 & ~n8314;
  assign n8316 = ~i_StoB_REQ7 & ~n8315;
  assign n8317 = ~n6842 & ~n8316;
  assign n8318 = n6664 & ~n8317;
  assign n8319 = i_StoB_REQ7 & ~n8197;
  assign n8320 = ~n7523 & ~n8319;
  assign n8321 = ~n6664 & ~n8320;
  assign n8322 = ~n8318 & ~n8321;
  assign n8323 = controllable_BtoS_ACK7 & ~n8322;
  assign n8324 = i_StoB_REQ7 & ~n7522;
  assign n8325 = ~n8316 & ~n8324;
  assign n8326 = n6664 & ~n8325;
  assign n8327 = ~n6664 & ~n7522;
  assign n8328 = ~n8326 & ~n8327;
  assign n8329 = ~controllable_BtoS_ACK7 & ~n8328;
  assign n8330 = ~n8323 & ~n8329;
  assign n8331 = n6663 & ~n8330;
  assign n8332 = ~n7546 & ~n8331;
  assign n8333 = ~i_StoB_REQ8 & ~n8332;
  assign n8334 = ~n8237 & ~n8333;
  assign n8335 = controllable_BtoS_ACK8 & ~n8334;
  assign n8336 = i_StoB_REQ8 & ~n7545;
  assign n8337 = ~n8333 & ~n8336;
  assign n8338 = ~controllable_BtoS_ACK8 & ~n8337;
  assign n8339 = ~n8335 & ~n8338;
  assign n8340 = n6662 & ~n8339;
  assign n8341 = ~n7568 & ~n8340;
  assign n8342 = ~i_StoB_REQ10 & ~n8341;
  assign n8343 = ~n8233 & ~n8342;
  assign n8344 = controllable_BtoS_ACK10 & ~n8343;
  assign n8345 = i_StoB_REQ10 & ~n7567;
  assign n8346 = ~n8342 & ~n8345;
  assign n8347 = ~controllable_BtoS_ACK10 & ~n8346;
  assign n8348 = ~n8344 & ~n8347;
  assign n8349 = n6661 & ~n8348;
  assign n8350 = ~n6661 & ~n7607;
  assign n8351 = ~n8349 & ~n8350;
  assign n8352 = ~i_StoB_REQ11 & ~n8351;
  assign n8353 = ~n8229 & ~n8352;
  assign n8354 = controllable_ENQ & ~n8353;
  assign n8355 = ~n7615 & ~n8354;
  assign n8356 = ~i_StoB_REQ9 & ~n8355;
  assign n8357 = ~n7994 & ~n8356;
  assign n8358 = controllable_BtoS_ACK9 & ~n8357;
  assign n8359 = ~n7620 & ~n8039;
  assign n8360 = i_StoB_REQ9 & ~n8359;
  assign n8361 = ~n8356 & ~n8360;
  assign n8362 = ~controllable_BtoS_ACK9 & ~n8361;
  assign n8363 = ~n8358 & ~n8362;
  assign n8364 = controllable_DEQ & ~n8363;
  assign n8365 = ~i_StoB_REQ9 & ~n8353;
  assign n8366 = ~n8013 & ~n8365;
  assign n8367 = controllable_BtoS_ACK9 & ~n8366;
  assign n8368 = i_StoB_REQ9 & ~n8038;
  assign n8369 = ~n8365 & ~n8368;
  assign n8370 = ~controllable_BtoS_ACK9 & ~n8369;
  assign n8371 = ~n8367 & ~n8370;
  assign n8372 = ~controllable_DEQ & ~n8371;
  assign n8373 = ~n8364 & ~n8372;
  assign n8374 = i_nEMPTY & ~n8373;
  assign n8375 = controllable_ENQ & ~n8354;
  assign n8376 = ~i_StoB_REQ9 & ~n8375;
  assign n8377 = ~n7994 & ~n8376;
  assign n8378 = controllable_BtoS_ACK9 & ~n8377;
  assign n8379 = i_StoB_REQ9 & ~n8082;
  assign n8380 = ~n8376 & ~n8379;
  assign n8381 = ~controllable_BtoS_ACK9 & ~n8380;
  assign n8382 = ~n8378 & ~n8381;
  assign n8383 = ~controllable_DEQ & ~n8382;
  assign n8384 = ~n7645 & ~n8383;
  assign n8385 = ~i_nEMPTY & ~n8384;
  assign n8386 = ~n8374 & ~n8385;
  assign n8387 = i_FULL & ~n8386;
  assign n8388 = ~controllable_DEQ & ~n8363;
  assign n8389 = ~n7972 & ~n8388;
  assign n8390 = ~i_nEMPTY & ~n8389;
  assign n8391 = ~n8374 & ~n8390;
  assign n8392 = ~i_FULL & ~n8391;
  assign n8393 = ~n8387 & ~n8392;
  assign n8394 = ~i_RtoB_ACK0 & ~n8393;
  assign n8395 = ~n7213 & ~n8394;
  assign n8396 = n6660 & ~n8395;
  assign n8397 = n6661 & ~n8224;
  assign n8398 = ~n6661 & ~n6918;
  assign n8399 = ~n8397 & ~n8398;
  assign n8400 = ~i_StoB_REQ11 & ~n8399;
  assign n8401 = ~n7982 & ~n8400;
  assign n8402 = controllable_ENQ & ~n8401;
  assign n8403 = controllable_ENQ & ~n8402;
  assign n8404 = i_StoB_REQ9 & ~n8403;
  assign n8405 = ~n8042 & ~n8404;
  assign n8406 = controllable_BtoS_ACK9 & ~n8405;
  assign n8407 = ~n8039 & ~n8051;
  assign n8408 = i_StoB_REQ9 & ~n8407;
  assign n8409 = ~n8039 & ~n8054;
  assign n8410 = ~i_StoB_REQ9 & ~n8409;
  assign n8411 = ~n8408 & ~n8410;
  assign n8412 = ~controllable_BtoS_ACK9 & ~n8411;
  assign n8413 = ~n8406 & ~n8412;
  assign n8414 = controllable_DEQ & ~n8413;
  assign n8415 = i_StoB_REQ9 & ~n8401;
  assign n8416 = ~n8062 & ~n8415;
  assign n8417 = controllable_BtoS_ACK9 & ~n8416;
  assign n8418 = ~controllable_BtoS_ACK9 & ~n8038;
  assign n8419 = ~n8417 & ~n8418;
  assign n8420 = ~controllable_DEQ & ~n8419;
  assign n8421 = ~n8414 & ~n8420;
  assign n8422 = i_nEMPTY & ~n8421;
  assign n8423 = ~n8083 & ~n8404;
  assign n8424 = controllable_BtoS_ACK9 & ~n8423;
  assign n8425 = ~controllable_BtoS_ACK9 & ~n8082;
  assign n8426 = ~n8424 & ~n8425;
  assign n8427 = ~controllable_DEQ & ~n8426;
  assign n8428 = ~n8081 & ~n8427;
  assign n8429 = ~i_nEMPTY & ~n8428;
  assign n8430 = ~n8422 & ~n8429;
  assign n8431 = i_FULL & ~n8430;
  assign n8432 = ~controllable_DEQ & ~n8413;
  assign n8433 = ~n8131 & ~n8432;
  assign n8434 = ~i_nEMPTY & ~n8433;
  assign n8435 = ~n8422 & ~n8434;
  assign n8436 = ~i_FULL & ~n8435;
  assign n8437 = ~n8431 & ~n8436;
  assign n8438 = ~i_RtoB_ACK0 & ~n8437;
  assign n8439 = ~n8025 & ~n8438;
  assign n8440 = ~n6660 & ~n8439;
  assign n8441 = ~n8396 & ~n8440;
  assign n8442 = ~n6659 & ~n8441;
  assign n8443 = ~n8149 & ~n8441;
  assign n8444 = ~n8149 & ~n8443;
  assign n8445 = n6659 & ~n8444;
  assign n8446 = ~n8442 & ~n8445;
  assign n8447 = ~n6652 & ~n8446;
  assign n8448 = ~n8154 & ~n8447;
  assign n8449 = n6651 & ~n8448;
  assign n8450 = ~n7615 & ~n8039;
  assign n8451 = ~i_StoB_REQ9 & ~n8450;
  assign n8452 = ~n7994 & ~n8451;
  assign n8453 = controllable_BtoS_ACK9 & ~n8452;
  assign n8454 = ~n8360 & ~n8451;
  assign n8455 = ~controllable_BtoS_ACK9 & ~n8454;
  assign n8456 = ~n8453 & ~n8455;
  assign n8457 = controllable_DEQ & ~n8456;
  assign n8458 = ~n8013 & ~n8062;
  assign n8459 = controllable_BtoS_ACK9 & ~n8458;
  assign n8460 = ~n8418 & ~n8459;
  assign n8461 = ~controllable_DEQ & ~n8460;
  assign n8462 = ~n8457 & ~n8461;
  assign n8463 = i_nEMPTY & ~n8462;
  assign n8464 = ~n7994 & ~n8083;
  assign n8465 = controllable_BtoS_ACK9 & ~n8464;
  assign n8466 = ~n8425 & ~n8465;
  assign n8467 = ~controllable_DEQ & ~n8466;
  assign n8468 = ~n7645 & ~n8467;
  assign n8469 = ~i_nEMPTY & ~n8468;
  assign n8470 = ~n8463 & ~n8469;
  assign n8471 = i_FULL & ~n8470;
  assign n8472 = ~controllable_DEQ & ~n8456;
  assign n8473 = ~n7972 & ~n8472;
  assign n8474 = ~i_nEMPTY & ~n8473;
  assign n8475 = ~n8463 & ~n8474;
  assign n8476 = ~i_FULL & ~n8475;
  assign n8477 = ~n8471 & ~n8476;
  assign n8478 = ~i_RtoB_ACK0 & ~n8477;
  assign n8479 = ~n7213 & ~n8478;
  assign n8480 = n6660 & ~n8479;
  assign n8481 = ~n7994 & ~n8042;
  assign n8482 = controllable_BtoS_ACK9 & ~n8481;
  assign n8483 = ~n8412 & ~n8482;
  assign n8484 = controllable_DEQ & ~n8483;
  assign n8485 = ~n8461 & ~n8484;
  assign n8486 = i_nEMPTY & ~n8485;
  assign n8487 = ~n8081 & ~n8467;
  assign n8488 = ~i_nEMPTY & ~n8487;
  assign n8489 = ~n8486 & ~n8488;
  assign n8490 = i_FULL & ~n8489;
  assign n8491 = ~controllable_DEQ & ~n8483;
  assign n8492 = ~n8131 & ~n8491;
  assign n8493 = ~i_nEMPTY & ~n8492;
  assign n8494 = ~n8486 & ~n8493;
  assign n8495 = ~i_FULL & ~n8494;
  assign n8496 = ~n8490 & ~n8495;
  assign n8497 = ~i_RtoB_ACK0 & ~n8496;
  assign n8498 = ~n8025 & ~n8497;
  assign n8499 = ~n6660 & ~n8498;
  assign n8500 = ~n8480 & ~n8499;
  assign n8501 = ~n6659 & ~n8500;
  assign n8502 = ~n8149 & ~n8500;
  assign n8503 = ~n8149 & ~n8502;
  assign n8504 = n6659 & ~n8503;
  assign n8505 = ~n8501 & ~n8504;
  assign n8506 = ~n6651 & ~n8505;
  assign n8507 = ~n8449 & ~n8506;
  assign n8508 = ~controllable_BtoR_REQ0 & ~n8507;
  assign n8509 = ~controllable_BtoR_REQ0 & ~n8508;
  assign n8510 = i_RtoB_ACK1 & ~n8509;
  assign n8511 = i_StoB_REQ1 & ~n7399;
  assign n8512 = ~controllable_BtoS_ACK1 & ~n8511;
  assign n8513 = ~controllable_BtoS_ACK1 & ~n8512;
  assign n8514 = ~n6671 & ~n8513;
  assign n8515 = ~n6931 & ~n8514;
  assign n8516 = n6670 & ~n8515;
  assign n8517 = controllable_BtoS_ACK1 & ~n6927;
  assign n8518 = n6671 & ~n8517;
  assign n8519 = ~n6927 & ~n8512;
  assign n8520 = ~n6671 & ~n8519;
  assign n8521 = ~n8518 & ~n8520;
  assign n8522 = ~n6670 & ~n8521;
  assign n8523 = ~n8516 & ~n8522;
  assign n8524 = n6669 & ~n8523;
  assign n8525 = ~n6946 & ~n8524;
  assign n8526 = ~i_StoB_REQ2 & ~n8525;
  assign n8527 = ~i_StoB_REQ2 & ~n8526;
  assign n8528 = controllable_BtoS_ACK2 & ~n8527;
  assign n8529 = ~n6671 & ~n8514;
  assign n8530 = n6670 & ~n8529;
  assign n8531 = ~n8522 & ~n8530;
  assign n8532 = ~n6669 & ~n8531;
  assign n8533 = ~n8524 & ~n8532;
  assign n8534 = ~i_StoB_REQ2 & ~n8533;
  assign n8535 = ~n7390 & ~n8534;
  assign n8536 = ~controllable_BtoS_ACK2 & ~n8535;
  assign n8537 = ~n8528 & ~n8536;
  assign n8538 = n6668 & ~n8537;
  assign n8539 = ~n6968 & ~n8538;
  assign n8540 = ~i_StoB_REQ3 & ~n8539;
  assign n8541 = ~i_StoB_REQ3 & ~n8540;
  assign n8542 = controllable_BtoS_ACK3 & ~n8541;
  assign n8543 = n6669 & ~n8531;
  assign n8544 = ~n6946 & ~n8543;
  assign n8545 = ~i_StoB_REQ2 & ~n8544;
  assign n8546 = ~i_StoB_REQ2 & ~n8545;
  assign n8547 = controllable_BtoS_ACK2 & ~n8546;
  assign n8548 = ~i_StoB_REQ2 & ~n8531;
  assign n8549 = ~n7430 & ~n8548;
  assign n8550 = ~controllable_BtoS_ACK2 & ~n8549;
  assign n8551 = ~n8547 & ~n8550;
  assign n8552 = ~n6668 & ~n8551;
  assign n8553 = ~n8538 & ~n8552;
  assign n8554 = ~i_StoB_REQ3 & ~n8553;
  assign n8555 = ~n7389 & ~n8554;
  assign n8556 = ~controllable_BtoS_ACK3 & ~n8555;
  assign n8557 = ~n8542 & ~n8556;
  assign n8558 = n6667 & ~n8557;
  assign n8559 = n6668 & ~n8551;
  assign n8560 = ~n6968 & ~n8559;
  assign n8561 = ~i_StoB_REQ3 & ~n8560;
  assign n8562 = ~i_StoB_REQ3 & ~n8561;
  assign n8563 = controllable_BtoS_ACK3 & ~n8562;
  assign n8564 = ~i_StoB_REQ3 & ~n8551;
  assign n8565 = ~n7446 & ~n8564;
  assign n8566 = ~controllable_BtoS_ACK3 & ~n8565;
  assign n8567 = ~n8563 & ~n8566;
  assign n8568 = ~controllable_BtoS_ACK4 & ~n8567;
  assign n8569 = ~n6996 & ~n8568;
  assign n8570 = ~n6667 & ~n8569;
  assign n8571 = ~n8558 & ~n8570;
  assign n8572 = ~i_StoB_REQ4 & ~n8571;
  assign n8573 = ~n7272 & ~n8572;
  assign n8574 = n6666 & ~n8573;
  assign n8575 = ~n7015 & ~n8574;
  assign n8576 = ~i_StoB_REQ5 & ~n8575;
  assign n8577 = ~i_StoB_REQ5 & ~n8576;
  assign n8578 = controllable_BtoS_ACK5 & ~n8577;
  assign n8579 = n6667 & ~n8567;
  assign n8580 = ~n8570 & ~n8579;
  assign n8581 = ~i_StoB_REQ4 & ~n8580;
  assign n8582 = ~n7284 & ~n8581;
  assign n8583 = ~n6666 & ~n8582;
  assign n8584 = ~n8574 & ~n8583;
  assign n8585 = ~i_StoB_REQ5 & ~n8584;
  assign n8586 = ~n7387 & ~n8585;
  assign n8587 = ~controllable_BtoS_ACK5 & ~n8586;
  assign n8588 = ~n8578 & ~n8587;
  assign n8589 = n6665 & ~n8588;
  assign n8590 = ~n7038 & ~n8589;
  assign n8591 = ~i_StoB_REQ6 & ~n8590;
  assign n8592 = ~i_StoB_REQ6 & ~n8591;
  assign n8593 = controllable_BtoS_ACK6 & ~n8592;
  assign n8594 = n6666 & ~n8582;
  assign n8595 = ~n7015 & ~n8594;
  assign n8596 = ~i_StoB_REQ5 & ~n8595;
  assign n8597 = ~i_StoB_REQ5 & ~n8596;
  assign n8598 = controllable_BtoS_ACK5 & ~n8597;
  assign n8599 = ~i_StoB_REQ5 & ~n8582;
  assign n8600 = ~n7502 & ~n8599;
  assign n8601 = ~controllable_BtoS_ACK5 & ~n8600;
  assign n8602 = ~n8598 & ~n8601;
  assign n8603 = ~n6665 & ~n8602;
  assign n8604 = ~n8589 & ~n8603;
  assign n8605 = ~i_StoB_REQ6 & ~n8604;
  assign n8606 = ~n7386 & ~n8605;
  assign n8607 = ~controllable_BtoS_ACK6 & ~n8606;
  assign n8608 = ~n8593 & ~n8607;
  assign n8609 = ~i_StoB_REQ7 & ~n8608;
  assign n8610 = ~i_StoB_REQ7 & ~n8609;
  assign n8611 = n6664 & ~n8610;
  assign n8612 = ~n7070 & ~n8611;
  assign n8613 = controllable_BtoS_ACK7 & ~n8612;
  assign n8614 = ~n7385 & ~n8609;
  assign n8615 = n6664 & ~n8614;
  assign n8616 = n6665 & ~n8602;
  assign n8617 = ~n7038 & ~n8616;
  assign n8618 = ~i_StoB_REQ6 & ~n8617;
  assign n8619 = ~i_StoB_REQ6 & ~n8618;
  assign n8620 = controllable_BtoS_ACK6 & ~n8619;
  assign n8621 = ~i_StoB_REQ6 & ~n8602;
  assign n8622 = ~n7529 & ~n8621;
  assign n8623 = ~controllable_BtoS_ACK6 & ~n8622;
  assign n8624 = ~n8620 & ~n8623;
  assign n8625 = ~i_StoB_REQ7 & ~n8624;
  assign n8626 = ~n7517 & ~n8625;
  assign n8627 = ~n6664 & ~n8626;
  assign n8628 = ~n8615 & ~n8627;
  assign n8629 = ~controllable_BtoS_ACK7 & ~n8628;
  assign n8630 = ~n8613 & ~n8629;
  assign n8631 = n6663 & ~n8630;
  assign n8632 = ~n7096 & ~n8631;
  assign n8633 = ~i_StoB_REQ8 & ~n8632;
  assign n8634 = ~i_StoB_REQ8 & ~n8633;
  assign n8635 = controllable_BtoS_ACK8 & ~n8634;
  assign n8636 = ~i_StoB_REQ7 & ~n8625;
  assign n8637 = n6664 & ~n8636;
  assign n8638 = ~n7070 & ~n8637;
  assign n8639 = controllable_BtoS_ACK7 & ~n8638;
  assign n8640 = ~controllable_BtoS_ACK7 & ~n8626;
  assign n8641 = ~n8639 & ~n8640;
  assign n8642 = ~n6663 & ~n8641;
  assign n8643 = ~n8631 & ~n8642;
  assign n8644 = ~i_StoB_REQ8 & ~n8643;
  assign n8645 = ~n7384 & ~n8644;
  assign n8646 = ~controllable_BtoS_ACK8 & ~n8645;
  assign n8647 = ~n8635 & ~n8646;
  assign n8648 = n6662 & ~n8647;
  assign n8649 = ~n7125 & ~n8648;
  assign n8650 = ~i_StoB_REQ10 & ~n8649;
  assign n8651 = ~i_StoB_REQ10 & ~n8650;
  assign n8652 = controllable_BtoS_ACK10 & ~n8651;
  assign n8653 = n6663 & ~n8641;
  assign n8654 = ~n7096 & ~n8653;
  assign n8655 = ~i_StoB_REQ8 & ~n8654;
  assign n8656 = ~i_StoB_REQ8 & ~n8655;
  assign n8657 = controllable_BtoS_ACK8 & ~n8656;
  assign n8658 = ~i_StoB_REQ8 & ~n8641;
  assign n8659 = ~n7573 & ~n8658;
  assign n8660 = ~controllable_BtoS_ACK8 & ~n8659;
  assign n8661 = ~n8657 & ~n8660;
  assign n8662 = ~n6662 & ~n8661;
  assign n8663 = ~n8648 & ~n8662;
  assign n8664 = ~i_StoB_REQ10 & ~n8663;
  assign n8665 = ~n7383 & ~n8664;
  assign n8666 = ~controllable_BtoS_ACK10 & ~n8665;
  assign n8667 = ~n8652 & ~n8666;
  assign n8668 = n6661 & ~n8667;
  assign n8669 = n6662 & ~n8661;
  assign n8670 = ~n7125 & ~n8669;
  assign n8671 = ~i_StoB_REQ10 & ~n8670;
  assign n8672 = ~i_StoB_REQ10 & ~n8671;
  assign n8673 = controllable_BtoS_ACK10 & ~n8672;
  assign n8674 = ~i_StoB_REQ10 & ~n8661;
  assign n8675 = ~n7589 & ~n8674;
  assign n8676 = ~controllable_BtoS_ACK10 & ~n8675;
  assign n8677 = ~n8673 & ~n8676;
  assign n8678 = ~controllable_BtoS_ACK11 & ~n8677;
  assign n8679 = ~n7153 & ~n8678;
  assign n8680 = ~n6661 & ~n8679;
  assign n8681 = ~n8668 & ~n8680;
  assign n8682 = ~i_StoB_REQ11 & ~n8681;
  assign n8683 = ~n7372 & ~n8682;
  assign n8684 = controllable_ENQ & ~n8683;
  assign n8685 = controllable_ENQ & ~n8684;
  assign n8686 = i_StoB_REQ9 & ~n8685;
  assign n8687 = controllable_BtoS_ACK11 & ~n8667;
  assign n8688 = ~n7918 & ~n8687;
  assign n8689 = n6661 & ~n8688;
  assign n8690 = controllable_BtoS_ACK11 & ~n8677;
  assign n8691 = ~n7928 & ~n8690;
  assign n8692 = ~n6661 & ~n8691;
  assign n8693 = ~n8689 & ~n8692;
  assign n8694 = i_StoB_REQ11 & ~n8693;
  assign n8695 = i_StoB_REQ10 & ~n8663;
  assign n8696 = i_StoB_REQ8 & ~n8643;
  assign n8697 = i_StoB_REQ7 & ~n8608;
  assign n8698 = i_StoB_REQ6 & ~n8604;
  assign n8699 = i_StoB_REQ5 & ~n8584;
  assign n8700 = controllable_BtoS_ACK4 & ~n8557;
  assign n8701 = ~n7732 & ~n8700;
  assign n8702 = n6667 & ~n8701;
  assign n8703 = controllable_BtoS_ACK4 & ~n8567;
  assign n8704 = ~n7742 & ~n8703;
  assign n8705 = ~n6667 & ~n8704;
  assign n8706 = ~n8702 & ~n8705;
  assign n8707 = i_StoB_REQ4 & ~n8706;
  assign n8708 = i_StoB_REQ3 & ~n8553;
  assign n8709 = i_StoB_REQ2 & ~n8533;
  assign n8710 = controllable_BtoS_ACK1 & ~n6924;
  assign n8711 = ~i_StoB_REQ1 & n6924;
  assign n8712 = ~i_StoB_REQ1 & ~n8711;
  assign n8713 = ~controllable_BtoS_ACK1 & n8712;
  assign n8714 = ~n8710 & ~n8713;
  assign n8715 = n6671 & ~n8714;
  assign n8716 = ~n6936 & ~n8715;
  assign n8717 = n6670 & ~n8716;
  assign n8718 = ~n6943 & ~n8717;
  assign n8719 = n6669 & ~n8718;
  assign n8720 = ~n6669 & ~n8714;
  assign n8721 = ~n8719 & ~n8720;
  assign n8722 = ~i_StoB_REQ2 & ~n8721;
  assign n8723 = ~n8709 & ~n8722;
  assign n8724 = controllable_BtoS_ACK2 & ~n8723;
  assign n8725 = ~n6954 & ~n8719;
  assign n8726 = ~i_StoB_REQ2 & ~n8725;
  assign n8727 = ~n7690 & ~n8726;
  assign n8728 = ~controllable_BtoS_ACK2 & ~n8727;
  assign n8729 = ~n8724 & ~n8728;
  assign n8730 = n6668 & ~n8729;
  assign n8731 = i_StoB_REQ2 & ~n6930;
  assign n8732 = ~i_StoB_REQ2 & ~n8714;
  assign n8733 = ~n8731 & ~n8732;
  assign n8734 = controllable_BtoS_ACK2 & ~n8733;
  assign n8735 = ~n8280 & ~n8732;
  assign n8736 = ~controllable_BtoS_ACK2 & ~n8735;
  assign n8737 = ~n8734 & ~n8736;
  assign n8738 = ~n6668 & ~n8737;
  assign n8739 = ~n8730 & ~n8738;
  assign n8740 = ~i_StoB_REQ3 & ~n8739;
  assign n8741 = ~n8708 & ~n8740;
  assign n8742 = controllable_BtoS_ACK3 & ~n8741;
  assign n8743 = i_StoB_REQ2 & ~n8531;
  assign n8744 = ~n6973 & ~n8720;
  assign n8745 = ~i_StoB_REQ2 & ~n8744;
  assign n8746 = ~n8743 & ~n8745;
  assign n8747 = controllable_BtoS_ACK2 & ~n8746;
  assign n8748 = ~n6978 & ~n7721;
  assign n8749 = ~controllable_BtoS_ACK2 & ~n8748;
  assign n8750 = ~n8747 & ~n8749;
  assign n8751 = ~n6668 & ~n8750;
  assign n8752 = ~n8730 & ~n8751;
  assign n8753 = ~i_StoB_REQ3 & ~n8752;
  assign n8754 = ~n7714 & ~n8753;
  assign n8755 = ~controllable_BtoS_ACK3 & ~n8754;
  assign n8756 = ~n8742 & ~n8755;
  assign n8757 = n6667 & ~n8756;
  assign n8758 = i_StoB_REQ3 & ~n6967;
  assign n8759 = ~i_StoB_REQ3 & ~n8737;
  assign n8760 = ~n8758 & ~n8759;
  assign n8761 = controllable_BtoS_ACK3 & ~n8760;
  assign n8762 = ~n8289 & ~n8759;
  assign n8763 = ~controllable_BtoS_ACK3 & ~n8762;
  assign n8764 = ~n8761 & ~n8763;
  assign n8765 = controllable_BtoS_ACK4 & ~n8764;
  assign n8766 = i_StoB_REQ3 & ~n8551;
  assign n8767 = n6668 & ~n8750;
  assign n8768 = ~n8738 & ~n8767;
  assign n8769 = ~i_StoB_REQ3 & ~n8768;
  assign n8770 = ~n8766 & ~n8769;
  assign n8771 = controllable_BtoS_ACK3 & ~n8770;
  assign n8772 = ~i_StoB_REQ3 & ~n8750;
  assign n8773 = ~n7754 & ~n8772;
  assign n8774 = ~controllable_BtoS_ACK3 & ~n8773;
  assign n8775 = ~n8771 & ~n8774;
  assign n8776 = ~controllable_BtoS_ACK4 & ~n8775;
  assign n8777 = ~n8765 & ~n8776;
  assign n8778 = ~n6667 & ~n8777;
  assign n8779 = ~n8757 & ~n8778;
  assign n8780 = ~i_StoB_REQ4 & ~n8779;
  assign n8781 = ~n8707 & ~n8780;
  assign n8782 = n6666 & ~n8781;
  assign n8783 = ~n6996 & ~n7472;
  assign n8784 = i_StoB_REQ4 & ~n8783;
  assign n8785 = ~i_StoB_REQ4 & ~n8764;
  assign n8786 = ~n8784 & ~n8785;
  assign n8787 = ~n6666 & ~n8786;
  assign n8788 = ~n8782 & ~n8787;
  assign n8789 = ~i_StoB_REQ5 & ~n8788;
  assign n8790 = ~n8699 & ~n8789;
  assign n8791 = controllable_BtoS_ACK5 & ~n8790;
  assign n8792 = ~n7759 & ~n8703;
  assign n8793 = n6667 & ~n8792;
  assign n8794 = ~n8705 & ~n8793;
  assign n8795 = i_StoB_REQ4 & ~n8794;
  assign n8796 = n6667 & ~n8775;
  assign n8797 = ~n8778 & ~n8796;
  assign n8798 = ~i_StoB_REQ4 & ~n8797;
  assign n8799 = ~n8795 & ~n8798;
  assign n8800 = ~n6666 & ~n8799;
  assign n8801 = ~n8782 & ~n8800;
  assign n8802 = ~i_StoB_REQ5 & ~n8801;
  assign n8803 = ~n7779 & ~n8802;
  assign n8804 = ~controllable_BtoS_ACK5 & ~n8803;
  assign n8805 = ~n8791 & ~n8804;
  assign n8806 = n6665 & ~n8805;
  assign n8807 = i_StoB_REQ5 & ~n7014;
  assign n8808 = ~i_StoB_REQ5 & ~n8786;
  assign n8809 = ~n8807 & ~n8808;
  assign n8810 = controllable_BtoS_ACK5 & ~n8809;
  assign n8811 = ~n8303 & ~n8808;
  assign n8812 = ~controllable_BtoS_ACK5 & ~n8811;
  assign n8813 = ~n8810 & ~n8812;
  assign n8814 = ~n6665 & ~n8813;
  assign n8815 = ~n8806 & ~n8814;
  assign n8816 = ~i_StoB_REQ6 & ~n8815;
  assign n8817 = ~n8698 & ~n8816;
  assign n8818 = controllable_BtoS_ACK6 & ~n8817;
  assign n8819 = i_StoB_REQ5 & ~n8582;
  assign n8820 = n6666 & ~n8799;
  assign n8821 = ~n8787 & ~n8820;
  assign n8822 = ~i_StoB_REQ5 & ~n8821;
  assign n8823 = ~n8819 & ~n8822;
  assign n8824 = controllable_BtoS_ACK5 & ~n8823;
  assign n8825 = ~i_StoB_REQ5 & ~n8799;
  assign n8826 = ~n7815 & ~n8825;
  assign n8827 = ~controllable_BtoS_ACK5 & ~n8826;
  assign n8828 = ~n8824 & ~n8827;
  assign n8829 = ~n6665 & ~n8828;
  assign n8830 = ~n8806 & ~n8829;
  assign n8831 = ~i_StoB_REQ6 & ~n8830;
  assign n8832 = ~n7808 & ~n8831;
  assign n8833 = ~controllable_BtoS_ACK6 & ~n8832;
  assign n8834 = ~n8818 & ~n8833;
  assign n8835 = ~i_StoB_REQ7 & ~n8834;
  assign n8836 = ~n8697 & ~n8835;
  assign n8837 = n6664 & ~n8836;
  assign n8838 = i_StoB_REQ7 & ~n8624;
  assign n8839 = i_StoB_REQ6 & ~n7037;
  assign n8840 = ~i_StoB_REQ6 & ~n8813;
  assign n8841 = ~n8839 & ~n8840;
  assign n8842 = controllable_BtoS_ACK6 & ~n8841;
  assign n8843 = ~n8312 & ~n8840;
  assign n8844 = ~controllable_BtoS_ACK6 & ~n8843;
  assign n8845 = ~n8842 & ~n8844;
  assign n8846 = ~i_StoB_REQ7 & ~n8845;
  assign n8847 = ~n8838 & ~n8846;
  assign n8848 = ~n6664 & ~n8847;
  assign n8849 = ~n8837 & ~n8848;
  assign n8850 = controllable_BtoS_ACK7 & ~n8849;
  assign n8851 = i_StoB_REQ7 & ~n7825;
  assign n8852 = ~n8835 & ~n8851;
  assign n8853 = n6664 & ~n8852;
  assign n8854 = i_StoB_REQ6 & ~n8602;
  assign n8855 = n6665 & ~n8828;
  assign n8856 = ~n8814 & ~n8855;
  assign n8857 = ~i_StoB_REQ6 & ~n8856;
  assign n8858 = ~n8854 & ~n8857;
  assign n8859 = controllable_BtoS_ACK6 & ~n8858;
  assign n8860 = ~i_StoB_REQ6 & ~n8828;
  assign n8861 = ~n7846 & ~n8860;
  assign n8862 = ~controllable_BtoS_ACK6 & ~n8861;
  assign n8863 = ~n8859 & ~n8862;
  assign n8864 = ~i_StoB_REQ7 & ~n8863;
  assign n8865 = ~n7839 & ~n8864;
  assign n8866 = ~n6664 & ~n8865;
  assign n8867 = ~n8853 & ~n8866;
  assign n8868 = ~controllable_BtoS_ACK7 & ~n8867;
  assign n8869 = ~n8850 & ~n8868;
  assign n8870 = n6663 & ~n8869;
  assign n8871 = i_StoB_REQ7 & ~n7067;
  assign n8872 = ~n8846 & ~n8871;
  assign n8873 = controllable_BtoS_ACK7 & ~n8872;
  assign n8874 = ~n8324 & ~n8846;
  assign n8875 = ~controllable_BtoS_ACK7 & ~n8874;
  assign n8876 = ~n8873 & ~n8875;
  assign n8877 = ~n6663 & ~n8876;
  assign n8878 = ~n8870 & ~n8877;
  assign n8879 = ~i_StoB_REQ8 & ~n8878;
  assign n8880 = ~n8696 & ~n8879;
  assign n8881 = controllable_BtoS_ACK8 & ~n8880;
  assign n8882 = ~n8838 & ~n8864;
  assign n8883 = n6664 & ~n8882;
  assign n8884 = ~n8848 & ~n8883;
  assign n8885 = controllable_BtoS_ACK7 & ~n8884;
  assign n8886 = i_StoB_REQ7 & ~n7850;
  assign n8887 = ~n8864 & ~n8886;
  assign n8888 = n6664 & ~n8887;
  assign n8889 = ~n8866 & ~n8888;
  assign n8890 = ~controllable_BtoS_ACK7 & ~n8889;
  assign n8891 = ~n8885 & ~n8890;
  assign n8892 = ~n6663 & ~n8891;
  assign n8893 = ~n8870 & ~n8892;
  assign n8894 = ~i_StoB_REQ8 & ~n8893;
  assign n8895 = ~n7871 & ~n8894;
  assign n8896 = ~controllable_BtoS_ACK8 & ~n8895;
  assign n8897 = ~n8881 & ~n8896;
  assign n8898 = n6662 & ~n8897;
  assign n8899 = i_StoB_REQ8 & ~n7095;
  assign n8900 = ~i_StoB_REQ8 & ~n8876;
  assign n8901 = ~n8899 & ~n8900;
  assign n8902 = controllable_BtoS_ACK8 & ~n8901;
  assign n8903 = ~n8336 & ~n8900;
  assign n8904 = ~controllable_BtoS_ACK8 & ~n8903;
  assign n8905 = ~n8902 & ~n8904;
  assign n8906 = ~n6662 & ~n8905;
  assign n8907 = ~n8898 & ~n8906;
  assign n8908 = ~i_StoB_REQ10 & ~n8907;
  assign n8909 = ~n8695 & ~n8908;
  assign n8910 = controllable_BtoS_ACK10 & ~n8909;
  assign n8911 = i_StoB_REQ8 & ~n8641;
  assign n8912 = n6663 & ~n8891;
  assign n8913 = ~n8877 & ~n8912;
  assign n8914 = ~i_StoB_REQ8 & ~n8913;
  assign n8915 = ~n8911 & ~n8914;
  assign n8916 = controllable_BtoS_ACK8 & ~n8915;
  assign n8917 = ~i_StoB_REQ8 & ~n8891;
  assign n8918 = ~n7907 & ~n8917;
  assign n8919 = ~controllable_BtoS_ACK8 & ~n8918;
  assign n8920 = ~n8916 & ~n8919;
  assign n8921 = ~n6662 & ~n8920;
  assign n8922 = ~n8898 & ~n8921;
  assign n8923 = ~i_StoB_REQ10 & ~n8922;
  assign n8924 = ~n7900 & ~n8923;
  assign n8925 = ~controllable_BtoS_ACK10 & ~n8924;
  assign n8926 = ~n8910 & ~n8925;
  assign n8927 = n6661 & ~n8926;
  assign n8928 = i_StoB_REQ10 & ~n7124;
  assign n8929 = ~i_StoB_REQ10 & ~n8905;
  assign n8930 = ~n8928 & ~n8929;
  assign n8931 = controllable_BtoS_ACK10 & ~n8930;
  assign n8932 = ~n8345 & ~n8929;
  assign n8933 = ~controllable_BtoS_ACK10 & ~n8932;
  assign n8934 = ~n8931 & ~n8933;
  assign n8935 = controllable_BtoS_ACK11 & ~n8934;
  assign n8936 = i_StoB_REQ10 & ~n8661;
  assign n8937 = n6662 & ~n8920;
  assign n8938 = ~n8906 & ~n8937;
  assign n8939 = ~i_StoB_REQ10 & ~n8938;
  assign n8940 = ~n8936 & ~n8939;
  assign n8941 = controllable_BtoS_ACK10 & ~n8940;
  assign n8942 = ~i_StoB_REQ10 & ~n8920;
  assign n8943 = ~n7940 & ~n8942;
  assign n8944 = ~controllable_BtoS_ACK10 & ~n8943;
  assign n8945 = ~n8941 & ~n8944;
  assign n8946 = ~controllable_BtoS_ACK11 & ~n8945;
  assign n8947 = ~n8935 & ~n8946;
  assign n8948 = ~n6661 & ~n8947;
  assign n8949 = ~n8927 & ~n8948;
  assign n8950 = ~i_StoB_REQ11 & ~n8949;
  assign n8951 = ~n8694 & ~n8950;
  assign n8952 = controllable_ENQ & ~n8951;
  assign n8953 = controllable_ENQ & ~n8952;
  assign n8954 = ~i_StoB_REQ9 & ~n8953;
  assign n8955 = ~n8686 & ~n8954;
  assign n8956 = controllable_BtoS_ACK9 & ~n8955;
  assign n8957 = controllable_ENQ & ~n7951;
  assign n8958 = i_StoB_REQ9 & ~n8957;
  assign n8959 = ~n8954 & ~n8958;
  assign n8960 = ~controllable_BtoS_ACK9 & ~n8959;
  assign n8961 = ~n8956 & ~n8960;
  assign n8962 = controllable_DEQ & ~n8961;
  assign n8963 = i_StoB_REQ9 & ~n8683;
  assign n8964 = ~i_StoB_REQ9 & ~n8951;
  assign n8965 = ~n8963 & ~n8964;
  assign n8966 = controllable_BtoS_ACK9 & ~n8965;
  assign n8967 = i_StoB_REQ9 & ~n7950;
  assign n8968 = ~n8964 & ~n8967;
  assign n8969 = ~controllable_BtoS_ACK9 & ~n8968;
  assign n8970 = ~n8966 & ~n8969;
  assign n8971 = ~controllable_DEQ & ~n8970;
  assign n8972 = ~n8962 & ~n8971;
  assign n8973 = i_nEMPTY & ~n8972;
  assign n8974 = ~controllable_DEQ & ~n8961;
  assign n8975 = ~controllable_DEQ & ~n8974;
  assign n8976 = ~i_nEMPTY & ~n8975;
  assign n8977 = ~n8973 & ~n8976;
  assign n8978 = i_RtoB_ACK0 & ~n8977;
  assign n8979 = ~controllable_ENQ & ~n8683;
  assign n8980 = ~n7379 & ~n8979;
  assign n8981 = i_StoB_REQ9 & ~n8980;
  assign n8982 = ~controllable_ENQ & ~n8951;
  assign n8983 = ~n7614 & ~n8982;
  assign n8984 = ~i_StoB_REQ9 & ~n8983;
  assign n8985 = ~n8981 & ~n8984;
  assign n8986 = controllable_BtoS_ACK9 & ~n8985;
  assign n8987 = i_StoB_REQ9 & ~n7963;
  assign n8988 = ~n8984 & ~n8987;
  assign n8989 = ~controllable_BtoS_ACK9 & ~n8988;
  assign n8990 = ~n8986 & ~n8989;
  assign n8991 = controllable_DEQ & ~n8990;
  assign n8992 = ~n7633 & ~n8991;
  assign n8993 = i_nEMPTY & ~n8992;
  assign n8994 = ~controllable_ENQ & ~n8979;
  assign n8995 = i_StoB_REQ9 & ~n8994;
  assign n8996 = ~controllable_ENQ & ~n8982;
  assign n8997 = ~i_StoB_REQ9 & ~n8996;
  assign n8998 = ~n8995 & ~n8997;
  assign n8999 = controllable_BtoS_ACK9 & ~n8998;
  assign n9000 = ~controllable_ENQ & ~n7962;
  assign n9001 = i_StoB_REQ9 & ~n9000;
  assign n9002 = ~n8997 & ~n9001;
  assign n9003 = ~controllable_BtoS_ACK9 & ~n9002;
  assign n9004 = ~n8999 & ~n9003;
  assign n9005 = controllable_DEQ & ~n9004;
  assign n9006 = ~n7652 & ~n9005;
  assign n9007 = ~i_nEMPTY & ~n9006;
  assign n9008 = ~n8993 & ~n9007;
  assign n9009 = i_FULL & ~n9008;
  assign n9010 = ~n7951 & ~n8982;
  assign n9011 = ~i_StoB_REQ9 & ~n9010;
  assign n9012 = ~n8981 & ~n9011;
  assign n9013 = controllable_BtoS_ACK9 & ~n9012;
  assign n9014 = ~n8967 & ~n9011;
  assign n9015 = ~controllable_BtoS_ACK9 & ~n9014;
  assign n9016 = ~n9013 & ~n9015;
  assign n9017 = controllable_DEQ & ~n9016;
  assign n9018 = ~n7969 & ~n9017;
  assign n9019 = i_nEMPTY & ~n9018;
  assign n9020 = controllable_DEQ & ~n8970;
  assign n9021 = ~controllable_DEQ & ~n8990;
  assign n9022 = ~n9020 & ~n9021;
  assign n9023 = ~i_nEMPTY & ~n9022;
  assign n9024 = ~n9019 & ~n9023;
  assign n9025 = ~i_FULL & ~n9024;
  assign n9026 = ~n9009 & ~n9025;
  assign n9027 = ~i_RtoB_ACK0 & ~n9026;
  assign n9028 = ~n8978 & ~n9027;
  assign n9029 = n6660 & ~n9028;
  assign n9030 = n6661 & ~n8677;
  assign n9031 = ~n8680 & ~n9030;
  assign n9032 = ~i_StoB_REQ11 & ~n9031;
  assign n9033 = ~n8026 & ~n9032;
  assign n9034 = controllable_ENQ & ~n9033;
  assign n9035 = controllable_ENQ & ~n9034;
  assign n9036 = i_StoB_REQ9 & ~n9035;
  assign n9037 = ~n7153 & ~n8034;
  assign n9038 = i_StoB_REQ11 & ~n9037;
  assign n9039 = ~i_StoB_REQ11 & ~n8934;
  assign n9040 = ~n9038 & ~n9039;
  assign n9041 = controllable_ENQ & ~n9040;
  assign n9042 = controllable_ENQ & ~n9041;
  assign n9043 = ~i_StoB_REQ9 & ~n9042;
  assign n9044 = ~n9036 & ~n9043;
  assign n9045 = controllable_BtoS_ACK9 & ~n9044;
  assign n9046 = controllable_ENQ & ~n8101;
  assign n9047 = i_StoB_REQ9 & ~n9046;
  assign n9048 = ~n7945 & ~n8690;
  assign n9049 = n6661 & ~n9048;
  assign n9050 = ~n8692 & ~n9049;
  assign n9051 = i_StoB_REQ11 & ~n9050;
  assign n9052 = n6661 & ~n8945;
  assign n9053 = ~n8948 & ~n9052;
  assign n9054 = ~i_StoB_REQ11 & ~n9053;
  assign n9055 = ~n9051 & ~n9054;
  assign n9056 = controllable_ENQ & ~n9055;
  assign n9057 = controllable_ENQ & ~n9056;
  assign n9058 = ~i_StoB_REQ9 & ~n9057;
  assign n9059 = ~n9047 & ~n9058;
  assign n9060 = ~controllable_BtoS_ACK9 & ~n9059;
  assign n9061 = ~n9045 & ~n9060;
  assign n9062 = controllable_DEQ & ~n9061;
  assign n9063 = i_StoB_REQ9 & ~n9033;
  assign n9064 = ~i_StoB_REQ9 & ~n9040;
  assign n9065 = ~n9063 & ~n9064;
  assign n9066 = controllable_BtoS_ACK9 & ~n9065;
  assign n9067 = i_StoB_REQ9 & ~n8100;
  assign n9068 = ~i_StoB_REQ9 & ~n9055;
  assign n9069 = ~n9067 & ~n9068;
  assign n9070 = ~controllable_BtoS_ACK9 & ~n9069;
  assign n9071 = ~n9066 & ~n9070;
  assign n9072 = ~controllable_DEQ & ~n9071;
  assign n9073 = ~n9062 & ~n9072;
  assign n9074 = i_nEMPTY & ~n9073;
  assign n9075 = ~controllable_DEQ & ~n9061;
  assign n9076 = ~controllable_DEQ & ~n9075;
  assign n9077 = ~i_nEMPTY & ~n9076;
  assign n9078 = ~n9074 & ~n9077;
  assign n9079 = i_RtoB_ACK0 & ~n9078;
  assign n9080 = ~controllable_ENQ & ~n9033;
  assign n9081 = ~n8031 & ~n9080;
  assign n9082 = i_StoB_REQ9 & ~n9081;
  assign n9083 = ~controllable_ENQ & ~n9040;
  assign n9084 = ~n8039 & ~n9083;
  assign n9085 = ~i_StoB_REQ9 & ~n9084;
  assign n9086 = ~n9082 & ~n9085;
  assign n9087 = controllable_BtoS_ACK9 & ~n9086;
  assign n9088 = ~controllable_ENQ & ~n9055;
  assign n9089 = ~n8050 & ~n9088;
  assign n9090 = ~i_StoB_REQ9 & ~n9089;
  assign n9091 = ~n8121 & ~n9090;
  assign n9092 = ~controllable_BtoS_ACK9 & ~n9091;
  assign n9093 = ~n9087 & ~n9092;
  assign n9094 = controllable_DEQ & ~n9093;
  assign n9095 = ~n8067 & ~n9094;
  assign n9096 = i_nEMPTY & ~n9095;
  assign n9097 = ~controllable_ENQ & ~n9080;
  assign n9098 = i_StoB_REQ9 & ~n9097;
  assign n9099 = ~controllable_ENQ & ~n9083;
  assign n9100 = ~i_StoB_REQ9 & ~n9099;
  assign n9101 = ~n9098 & ~n9100;
  assign n9102 = controllable_BtoS_ACK9 & ~n9101;
  assign n9103 = ~controllable_ENQ & ~n8119;
  assign n9104 = i_StoB_REQ9 & ~n9103;
  assign n9105 = ~controllable_ENQ & ~n9088;
  assign n9106 = ~i_StoB_REQ9 & ~n9105;
  assign n9107 = ~n9104 & ~n9106;
  assign n9108 = ~controllable_BtoS_ACK9 & ~n9107;
  assign n9109 = ~n9102 & ~n9108;
  assign n9110 = controllable_DEQ & ~n9109;
  assign n9111 = ~n8089 & ~n9110;
  assign n9112 = ~i_nEMPTY & ~n9111;
  assign n9113 = ~n9096 & ~n9112;
  assign n9114 = i_FULL & ~n9113;
  assign n9115 = ~n8112 & ~n9088;
  assign n9116 = ~i_StoB_REQ9 & ~n9115;
  assign n9117 = ~n9067 & ~n9116;
  assign n9118 = ~controllable_BtoS_ACK9 & ~n9117;
  assign n9119 = ~n9087 & ~n9118;
  assign n9120 = controllable_DEQ & ~n9119;
  assign n9121 = ~n8128 & ~n9120;
  assign n9122 = i_nEMPTY & ~n9121;
  assign n9123 = controllable_DEQ & ~n9071;
  assign n9124 = ~controllable_DEQ & ~n9093;
  assign n9125 = ~n9123 & ~n9124;
  assign n9126 = ~i_nEMPTY & ~n9125;
  assign n9127 = ~n9122 & ~n9126;
  assign n9128 = ~i_FULL & ~n9127;
  assign n9129 = ~n9114 & ~n9128;
  assign n9130 = ~i_RtoB_ACK0 & ~n9129;
  assign n9131 = ~n9079 & ~n9130;
  assign n9132 = ~n6660 & ~n9131;
  assign n9133 = ~n9029 & ~n9132;
  assign n9134 = ~n6659 & ~n9133;
  assign n9135 = ~n8149 & ~n9133;
  assign n9136 = ~n8149 & ~n9135;
  assign n9137 = n6659 & ~n9136;
  assign n9138 = ~n9134 & ~n9137;
  assign n9139 = ~controllable_BtoR_REQ0 & ~n9138;
  assign n9140 = ~controllable_BtoR_REQ0 & ~n9139;
  assign n9141 = ~i_RtoB_ACK1 & ~n9140;
  assign n9142 = ~n8510 & ~n9141;
  assign n9143 = controllable_BtoR_REQ1 & ~n9142;
  assign n9144 = ~i_RtoB_ACK0 & ~n8977;
  assign n9145 = ~n7213 & ~n9144;
  assign n9146 = n6660 & ~n9145;
  assign n9147 = ~i_RtoB_ACK0 & ~n9078;
  assign n9148 = ~n8025 & ~n9147;
  assign n9149 = ~n6660 & ~n9148;
  assign n9150 = ~n9146 & ~n9149;
  assign n9151 = ~n8149 & ~n9150;
  assign n9152 = ~n8149 & ~n9151;
  assign n9153 = ~n6659 & ~n9152;
  assign n9154 = n6659 & ~n9150;
  assign n9155 = ~n9153 & ~n9154;
  assign n9156 = controllable_BtoR_REQ0 & ~n9155;
  assign n9157 = ~i_StoB_REQ9 & ~n8957;
  assign n9158 = ~n7381 & ~n9157;
  assign n9159 = controllable_BtoS_ACK9 & ~n9158;
  assign n9160 = ~controllable_BtoS_ACK9 & ~n8957;
  assign n9161 = ~n9159 & ~n9160;
  assign n9162 = controllable_DEQ & ~n9161;
  assign n9163 = ~i_StoB_REQ9 & ~n7950;
  assign n9164 = ~n7627 & ~n9163;
  assign n9165 = controllable_BtoS_ACK9 & ~n9164;
  assign n9166 = ~controllable_BtoS_ACK9 & ~n7950;
  assign n9167 = ~n9165 & ~n9166;
  assign n9168 = ~controllable_DEQ & ~n9167;
  assign n9169 = ~n9162 & ~n9168;
  assign n9170 = i_nEMPTY & ~n9169;
  assign n9171 = ~controllable_DEQ & ~n9161;
  assign n9172 = ~controllable_DEQ & ~n9171;
  assign n9173 = ~i_nEMPTY & ~n9172;
  assign n9174 = ~n9170 & ~n9173;
  assign n9175 = n6660 & ~n9174;
  assign n9176 = controllable_ENQ & ~n8112;
  assign n9177 = ~i_StoB_REQ9 & ~n9176;
  assign n9178 = ~n9047 & ~n9177;
  assign n9179 = ~controllable_BtoS_ACK9 & ~n9178;
  assign n9180 = ~n8085 & ~n9179;
  assign n9181 = controllable_DEQ & ~n9180;
  assign n9182 = ~i_StoB_REQ9 & ~n8111;
  assign n9183 = ~n9067 & ~n9182;
  assign n9184 = ~controllable_BtoS_ACK9 & ~n9183;
  assign n9185 = ~n8064 & ~n9184;
  assign n9186 = ~controllable_DEQ & ~n9185;
  assign n9187 = ~n9181 & ~n9186;
  assign n9188 = i_nEMPTY & ~n9187;
  assign n9189 = ~controllable_DEQ & ~n9180;
  assign n9190 = ~controllable_DEQ & ~n9189;
  assign n9191 = ~i_nEMPTY & ~n9190;
  assign n9192 = ~n9188 & ~n9191;
  assign n9193 = ~n6660 & ~n9192;
  assign n9194 = ~n9175 & ~n9193;
  assign n9195 = n6652 & ~n9194;
  assign n9196 = ~n6659 & ~n9194;
  assign n9197 = i_RtoB_ACK0 & ~n9174;
  assign n9198 = controllable_DEQ & ~n8382;
  assign n9199 = ~n8372 & ~n9198;
  assign n9200 = i_nEMPTY & ~n9199;
  assign n9201 = ~controllable_DEQ & ~n8383;
  assign n9202 = ~i_nEMPTY & ~n9201;
  assign n9203 = ~n9200 & ~n9202;
  assign n9204 = ~i_RtoB_ACK0 & ~n9203;
  assign n9205 = ~n9197 & ~n9204;
  assign n9206 = n6660 & ~n9205;
  assign n9207 = i_RtoB_ACK0 & ~n9192;
  assign n9208 = controllable_DEQ & ~n8426;
  assign n9209 = ~n8420 & ~n9208;
  assign n9210 = i_nEMPTY & ~n9209;
  assign n9211 = ~controllable_DEQ & ~n8427;
  assign n9212 = ~i_nEMPTY & ~n9211;
  assign n9213 = ~n9210 & ~n9212;
  assign n9214 = ~i_RtoB_ACK0 & ~n9213;
  assign n9215 = ~n9207 & ~n9214;
  assign n9216 = ~n6660 & ~n9215;
  assign n9217 = ~n9206 & ~n9216;
  assign n9218 = n6659 & ~n9217;
  assign n9219 = ~n9196 & ~n9218;
  assign n9220 = ~n6652 & ~n9219;
  assign n9221 = ~n9195 & ~n9220;
  assign n9222 = ~controllable_BtoR_REQ0 & ~n9221;
  assign n9223 = ~n9156 & ~n9222;
  assign n9224 = i_RtoB_ACK1 & ~n9223;
  assign n9225 = i_RtoB_ACK0 & ~n7978;
  assign n9226 = ~n9027 & ~n9225;
  assign n9227 = n6660 & ~n9226;
  assign n9228 = i_RtoB_ACK0 & ~n8137;
  assign n9229 = ~n9130 & ~n9228;
  assign n9230 = ~n6660 & ~n9229;
  assign n9231 = ~n9227 & ~n9230;
  assign n9232 = ~n8149 & ~n9231;
  assign n9233 = ~n8149 & ~n9232;
  assign n9234 = ~n6659 & ~n9233;
  assign n9235 = n6659 & ~n9231;
  assign n9236 = ~n9234 & ~n9235;
  assign n9237 = n6652 & ~n9236;
  assign n9238 = i_RtoB_ACK0 & ~n8477;
  assign n9239 = ~n9027 & ~n9238;
  assign n9240 = n6660 & ~n9239;
  assign n9241 = i_RtoB_ACK0 & ~n8496;
  assign n9242 = ~n9130 & ~n9241;
  assign n9243 = ~n6660 & ~n9242;
  assign n9244 = ~n9240 & ~n9243;
  assign n9245 = ~n8149 & ~n9244;
  assign n9246 = ~n8149 & ~n9245;
  assign n9247 = ~n6659 & ~n9246;
  assign n9248 = n6659 & ~n9244;
  assign n9249 = ~n9247 & ~n9248;
  assign n9250 = ~n6652 & ~n9249;
  assign n9251 = ~n9237 & ~n9250;
  assign n9252 = n6651 & ~n9251;
  assign n9253 = i_RtoB_ACK0 & ~n8393;
  assign n9254 = ~n9027 & ~n9253;
  assign n9255 = n6660 & ~n9254;
  assign n9256 = i_RtoB_ACK0 & ~n8437;
  assign n9257 = ~n9130 & ~n9256;
  assign n9258 = ~n6660 & ~n9257;
  assign n9259 = ~n9255 & ~n9258;
  assign n9260 = ~n8149 & ~n9259;
  assign n9261 = ~n8149 & ~n9260;
  assign n9262 = ~n6659 & ~n9261;
  assign n9263 = n6659 & ~n9259;
  assign n9264 = ~n9262 & ~n9263;
  assign n9265 = n6652 & ~n9264;
  assign n9266 = ~n9250 & ~n9265;
  assign n9267 = ~n6651 & ~n9266;
  assign n9268 = ~n9252 & ~n9267;
  assign n9269 = controllable_BtoR_REQ0 & ~n9268;
  assign n9270 = controllable_DEQ & ~n7968;
  assign n9271 = ~n7633 & ~n9270;
  assign n9272 = i_nEMPTY & ~n9271;
  assign n9273 = ~controllable_ENQ & ~n7378;
  assign n9274 = ~controllable_ENQ & ~n9273;
  assign n9275 = i_StoB_REQ9 & ~n9274;
  assign n9276 = ~i_StoB_REQ9 & ~n9000;
  assign n9277 = ~n9275 & ~n9276;
  assign n9278 = controllable_BtoS_ACK9 & ~n9277;
  assign n9279 = ~controllable_BtoS_ACK9 & ~n9000;
  assign n9280 = ~n9278 & ~n9279;
  assign n9281 = controllable_DEQ & ~n9280;
  assign n9282 = ~n7652 & ~n9281;
  assign n9283 = ~i_nEMPTY & ~n9282;
  assign n9284 = ~n9272 & ~n9283;
  assign n9285 = i_FULL & ~n9284;
  assign n9286 = controllable_DEQ & ~n9167;
  assign n9287 = ~n7969 & ~n9286;
  assign n9288 = i_nEMPTY & ~n9287;
  assign n9289 = ~n9021 & ~n9286;
  assign n9290 = ~i_nEMPTY & ~n9289;
  assign n9291 = ~n9288 & ~n9290;
  assign n9292 = ~i_FULL & ~n9291;
  assign n9293 = ~n9285 & ~n9292;
  assign n9294 = ~i_RtoB_ACK0 & ~n9293;
  assign n9295 = ~n9197 & ~n9294;
  assign n9296 = n6660 & ~n9295;
  assign n9297 = controllable_DEQ & ~n8127;
  assign n9298 = ~n8067 & ~n9297;
  assign n9299 = i_nEMPTY & ~n9298;
  assign n9300 = ~controllable_ENQ & ~n8030;
  assign n9301 = ~controllable_ENQ & ~n9300;
  assign n9302 = i_StoB_REQ9 & ~n9301;
  assign n9303 = ~controllable_ENQ & ~n8038;
  assign n9304 = ~controllable_ENQ & ~n9303;
  assign n9305 = ~i_StoB_REQ9 & ~n9304;
  assign n9306 = ~n9302 & ~n9305;
  assign n9307 = controllable_BtoS_ACK9 & ~n9306;
  assign n9308 = ~controllable_ENQ & ~n8122;
  assign n9309 = ~i_StoB_REQ9 & ~n9308;
  assign n9310 = ~n9104 & ~n9309;
  assign n9311 = ~controllable_BtoS_ACK9 & ~n9310;
  assign n9312 = ~n9307 & ~n9311;
  assign n9313 = controllable_DEQ & ~n9312;
  assign n9314 = ~n8089 & ~n9313;
  assign n9315 = ~i_nEMPTY & ~n9314;
  assign n9316 = ~n9299 & ~n9315;
  assign n9317 = i_FULL & ~n9316;
  assign n9318 = controllable_DEQ & ~n9185;
  assign n9319 = ~n8128 & ~n9318;
  assign n9320 = i_nEMPTY & ~n9319;
  assign n9321 = ~n9124 & ~n9318;
  assign n9322 = ~i_nEMPTY & ~n9321;
  assign n9323 = ~n9320 & ~n9322;
  assign n9324 = ~i_FULL & ~n9323;
  assign n9325 = ~n9317 & ~n9324;
  assign n9326 = ~i_RtoB_ACK0 & ~n9325;
  assign n9327 = ~n9207 & ~n9326;
  assign n9328 = ~n6660 & ~n9327;
  assign n9329 = ~n9296 & ~n9328;
  assign n9330 = n6652 & ~n9329;
  assign n9331 = ~n6659 & ~n9329;
  assign n9332 = ~n7379 & ~n8051;
  assign n9333 = i_StoB_REQ9 & ~n9332;
  assign n9334 = i_StoB_REQ10 & ~n7343;
  assign n9335 = i_StoB_REQ8 & ~n7327;
  assign n9336 = i_StoB_REQ6 & ~n7294;
  assign n9337 = i_StoB_REQ5 & ~n7280;
  assign n9338 = i_StoB_REQ3 & ~n7243;
  assign n9339 = i_StoB_REQ2 & ~n7231;
  assign n9340 = ~i_StoB_REQ1 & ~controllable_BtoS_ACK0;
  assign n9341 = ~n7399 & ~n9340;
  assign n9342 = controllable_BtoS_ACK1 & ~n9341;
  assign n9343 = ~controllable_BtoS_ACK0 & ~controllable_BtoS_ACK1;
  assign n9344 = ~n9342 & ~n9343;
  assign n9345 = ~n6671 & ~n9344;
  assign n9346 = ~n7392 & ~n9345;
  assign n9347 = n6670 & ~n9346;
  assign n9348 = controllable_BtoS_ACK1 & ~n7391;
  assign n9349 = n6671 & ~n9348;
  assign n9350 = ~n7391 & ~n9343;
  assign n9351 = ~n6671 & ~n9350;
  assign n9352 = ~n9349 & ~n9351;
  assign n9353 = ~n6670 & ~n9352;
  assign n9354 = ~n9347 & ~n9353;
  assign n9355 = n6669 & ~n9354;
  assign n9356 = ~n7407 & ~n9355;
  assign n9357 = ~i_StoB_REQ2 & ~n9356;
  assign n9358 = ~n9339 & ~n9357;
  assign n9359 = controllable_BtoS_ACK2 & ~n9358;
  assign n9360 = ~n6671 & ~n9345;
  assign n9361 = n6670 & ~n9360;
  assign n9362 = ~n9353 & ~n9361;
  assign n9363 = ~n6669 & ~n9362;
  assign n9364 = ~n9355 & ~n9363;
  assign n9365 = ~controllable_BtoS_ACK2 & ~n9364;
  assign n9366 = ~n9359 & ~n9365;
  assign n9367 = n6668 & ~n9366;
  assign n9368 = ~n7425 & ~n9367;
  assign n9369 = ~i_StoB_REQ3 & ~n9368;
  assign n9370 = ~n9338 & ~n9369;
  assign n9371 = controllable_BtoS_ACK3 & ~n9370;
  assign n9372 = i_StoB_REQ2 & ~n7248;
  assign n9373 = n6669 & ~n9362;
  assign n9374 = ~n7407 & ~n9373;
  assign n9375 = ~i_StoB_REQ2 & ~n9374;
  assign n9376 = ~n9372 & ~n9375;
  assign n9377 = controllable_BtoS_ACK2 & ~n9376;
  assign n9378 = ~controllable_BtoS_ACK2 & ~n9362;
  assign n9379 = ~n9377 & ~n9378;
  assign n9380 = ~n6668 & ~n9379;
  assign n9381 = ~n9367 & ~n9380;
  assign n9382 = ~controllable_BtoS_ACK3 & ~n9381;
  assign n9383 = ~n9371 & ~n9382;
  assign n9384 = ~controllable_BtoS_ACK4 & ~n9383;
  assign n9385 = ~n7388 & ~n9384;
  assign n9386 = n6667 & ~n9385;
  assign n9387 = i_StoB_REQ3 & ~n7262;
  assign n9388 = n6668 & ~n9379;
  assign n9389 = ~n7425 & ~n9388;
  assign n9390 = ~i_StoB_REQ3 & ~n9389;
  assign n9391 = ~n9387 & ~n9390;
  assign n9392 = controllable_BtoS_ACK3 & ~n9391;
  assign n9393 = ~controllable_BtoS_ACK3 & ~n9379;
  assign n9394 = ~n9392 & ~n9393;
  assign n9395 = ~controllable_BtoS_ACK4 & ~n9394;
  assign n9396 = ~n6759 & ~n9395;
  assign n9397 = ~n6667 & ~n9396;
  assign n9398 = ~n9386 & ~n9397;
  assign n9399 = i_StoB_REQ4 & ~n9398;
  assign n9400 = n6667 & ~n9383;
  assign n9401 = ~n7465 & ~n9395;
  assign n9402 = ~n6667 & ~n9401;
  assign n9403 = ~n9400 & ~n9402;
  assign n9404 = ~i_StoB_REQ4 & ~n9403;
  assign n9405 = ~n9399 & ~n9404;
  assign n9406 = n6666 & ~n9405;
  assign n9407 = ~n7477 & ~n9406;
  assign n9408 = ~i_StoB_REQ5 & ~n9407;
  assign n9409 = ~n9337 & ~n9408;
  assign n9410 = controllable_BtoS_ACK5 & ~n9409;
  assign n9411 = ~n7445 & ~n9395;
  assign n9412 = n6667 & ~n9411;
  assign n9413 = ~n9397 & ~n9412;
  assign n9414 = i_StoB_REQ4 & ~n9413;
  assign n9415 = n6667 & ~n9394;
  assign n9416 = ~n9402 & ~n9415;
  assign n9417 = ~i_StoB_REQ4 & ~n9416;
  assign n9418 = ~n9414 & ~n9417;
  assign n9419 = ~n6666 & ~n9418;
  assign n9420 = ~n9406 & ~n9419;
  assign n9421 = ~controllable_BtoS_ACK5 & ~n9420;
  assign n9422 = ~n9410 & ~n9421;
  assign n9423 = n6665 & ~n9422;
  assign n9424 = ~n7497 & ~n9423;
  assign n9425 = ~i_StoB_REQ6 & ~n9424;
  assign n9426 = ~n9336 & ~n9425;
  assign n9427 = controllable_BtoS_ACK6 & ~n9426;
  assign n9428 = i_StoB_REQ5 & ~n7299;
  assign n9429 = n6666 & ~n9418;
  assign n9430 = ~n7477 & ~n9429;
  assign n9431 = ~i_StoB_REQ5 & ~n9430;
  assign n9432 = ~n9428 & ~n9431;
  assign n9433 = controllable_BtoS_ACK5 & ~n9432;
  assign n9434 = ~controllable_BtoS_ACK5 & ~n9418;
  assign n9435 = ~n9433 & ~n9434;
  assign n9436 = ~n6665 & ~n9435;
  assign n9437 = ~n9423 & ~n9436;
  assign n9438 = ~controllable_BtoS_ACK6 & ~n9437;
  assign n9439 = ~n9427 & ~n9438;
  assign n9440 = ~i_StoB_REQ7 & ~n9439;
  assign n9441 = ~n7385 & ~n9440;
  assign n9442 = n6664 & ~n9441;
  assign n9443 = ~n6664 & ~n7542;
  assign n9444 = ~n9442 & ~n9443;
  assign n9445 = controllable_BtoS_ACK7 & ~n9444;
  assign n9446 = n6664 & ~n9439;
  assign n9447 = i_StoB_REQ6 & ~n7316;
  assign n9448 = n6665 & ~n9435;
  assign n9449 = ~n7497 & ~n9448;
  assign n9450 = ~i_StoB_REQ6 & ~n9449;
  assign n9451 = ~n9447 & ~n9450;
  assign n9452 = controllable_BtoS_ACK6 & ~n9451;
  assign n9453 = ~controllable_BtoS_ACK6 & ~n9435;
  assign n9454 = ~n9452 & ~n9453;
  assign n9455 = ~n6664 & ~n9454;
  assign n9456 = ~n9446 & ~n9455;
  assign n9457 = ~controllable_BtoS_ACK7 & ~n9456;
  assign n9458 = ~n9445 & ~n9457;
  assign n9459 = n6663 & ~n9458;
  assign n9460 = ~n7546 & ~n9459;
  assign n9461 = ~i_StoB_REQ8 & ~n9460;
  assign n9462 = ~n9335 & ~n9461;
  assign n9463 = controllable_BtoS_ACK8 & ~n9462;
  assign n9464 = ~i_StoB_REQ7 & ~n9454;
  assign n9465 = ~n7517 & ~n9464;
  assign n9466 = n6664 & ~n9465;
  assign n9467 = ~n9443 & ~n9466;
  assign n9468 = controllable_BtoS_ACK7 & ~n9467;
  assign n9469 = ~controllable_BtoS_ACK7 & ~n9454;
  assign n9470 = ~n9468 & ~n9469;
  assign n9471 = ~n6663 & ~n9470;
  assign n9472 = ~n9459 & ~n9471;
  assign n9473 = ~controllable_BtoS_ACK8 & ~n9472;
  assign n9474 = ~n9463 & ~n9473;
  assign n9475 = n6662 & ~n9474;
  assign n9476 = ~n7568 & ~n9475;
  assign n9477 = ~i_StoB_REQ10 & ~n9476;
  assign n9478 = ~n9334 & ~n9477;
  assign n9479 = controllable_BtoS_ACK10 & ~n9478;
  assign n9480 = i_StoB_REQ8 & ~n7348;
  assign n9481 = n6663 & ~n9470;
  assign n9482 = ~n7546 & ~n9481;
  assign n9483 = ~i_StoB_REQ8 & ~n9482;
  assign n9484 = ~n9480 & ~n9483;
  assign n9485 = controllable_BtoS_ACK8 & ~n9484;
  assign n9486 = ~controllable_BtoS_ACK8 & ~n9470;
  assign n9487 = ~n9485 & ~n9486;
  assign n9488 = ~n6662 & ~n9487;
  assign n9489 = ~n9475 & ~n9488;
  assign n9490 = ~controllable_BtoS_ACK10 & ~n9489;
  assign n9491 = ~n9479 & ~n9490;
  assign n9492 = ~controllable_BtoS_ACK11 & ~n9491;
  assign n9493 = ~n7382 & ~n9492;
  assign n9494 = n6661 & ~n9493;
  assign n9495 = i_StoB_REQ10 & ~n7362;
  assign n9496 = n6662 & ~n9487;
  assign n9497 = ~n7568 & ~n9496;
  assign n9498 = ~i_StoB_REQ10 & ~n9497;
  assign n9499 = ~n9495 & ~n9498;
  assign n9500 = controllable_BtoS_ACK10 & ~n9499;
  assign n9501 = ~controllable_BtoS_ACK10 & ~n9487;
  assign n9502 = ~n9500 & ~n9501;
  assign n9503 = ~controllable_BtoS_ACK11 & ~n9502;
  assign n9504 = ~n7178 & ~n9503;
  assign n9505 = ~n6661 & ~n9504;
  assign n9506 = ~n9494 & ~n9505;
  assign n9507 = i_StoB_REQ11 & ~n9506;
  assign n9508 = n6661 & ~n9491;
  assign n9509 = ~n7608 & ~n9503;
  assign n9510 = ~n6661 & ~n9509;
  assign n9511 = ~n9508 & ~n9510;
  assign n9512 = ~i_StoB_REQ11 & ~n9511;
  assign n9513 = ~n9507 & ~n9512;
  assign n9514 = controllable_ENQ & ~n9513;
  assign n9515 = ~controllable_ENQ & ~n8353;
  assign n9516 = ~n9514 & ~n9515;
  assign n9517 = ~i_StoB_REQ9 & ~n9516;
  assign n9518 = ~n9333 & ~n9517;
  assign n9519 = controllable_BtoS_ACK9 & ~n9518;
  assign n9520 = ~n9303 & ~n9514;
  assign n9521 = i_StoB_REQ9 & ~n9520;
  assign n9522 = ~n9517 & ~n9521;
  assign n9523 = ~controllable_BtoS_ACK9 & ~n9522;
  assign n9524 = ~n9519 & ~n9523;
  assign n9525 = controllable_DEQ & ~n9524;
  assign n9526 = ~i_StoB_REQ9 & ~n9513;
  assign n9527 = ~n7627 & ~n9526;
  assign n9528 = controllable_BtoS_ACK9 & ~n9527;
  assign n9529 = ~controllable_BtoS_ACK9 & ~n9513;
  assign n9530 = ~n9528 & ~n9529;
  assign n9531 = ~controllable_DEQ & ~n9530;
  assign n9532 = ~n9525 & ~n9531;
  assign n9533 = i_nEMPTY & ~n9532;
  assign n9534 = ~controllable_ENQ & ~n9515;
  assign n9535 = ~i_StoB_REQ9 & ~n9534;
  assign n9536 = ~n8075 & ~n9535;
  assign n9537 = controllable_BtoS_ACK9 & ~n9536;
  assign n9538 = i_StoB_REQ9 & ~n9304;
  assign n9539 = ~n9535 & ~n9538;
  assign n9540 = ~controllable_BtoS_ACK9 & ~n9539;
  assign n9541 = ~n9537 & ~n9540;
  assign n9542 = controllable_DEQ & ~n9541;
  assign n9543 = controllable_ENQ & ~n9514;
  assign n9544 = ~i_StoB_REQ9 & ~n9543;
  assign n9545 = ~n7381 & ~n9544;
  assign n9546 = controllable_BtoS_ACK9 & ~n9545;
  assign n9547 = ~controllable_BtoS_ACK9 & ~n9543;
  assign n9548 = ~n9546 & ~n9547;
  assign n9549 = ~controllable_DEQ & ~n9548;
  assign n9550 = ~n9542 & ~n9549;
  assign n9551 = ~i_nEMPTY & ~n9550;
  assign n9552 = ~n9533 & ~n9551;
  assign n9553 = i_FULL & ~n9552;
  assign n9554 = ~n8039 & ~n9515;
  assign n9555 = ~i_StoB_REQ9 & ~n9554;
  assign n9556 = ~n8013 & ~n9555;
  assign n9557 = controllable_BtoS_ACK9 & ~n9556;
  assign n9558 = ~n8368 & ~n9555;
  assign n9559 = ~controllable_BtoS_ACK9 & ~n9558;
  assign n9560 = ~n9557 & ~n9559;
  assign n9561 = controllable_DEQ & ~n9560;
  assign n9562 = ~i_StoB_REQ9 & ~n9520;
  assign n9563 = ~n9333 & ~n9562;
  assign n9564 = controllable_BtoS_ACK9 & ~n9563;
  assign n9565 = ~controllable_BtoS_ACK9 & ~n9520;
  assign n9566 = ~n9564 & ~n9565;
  assign n9567 = ~controllable_DEQ & ~n9566;
  assign n9568 = ~n9561 & ~n9567;
  assign n9569 = i_nEMPTY & ~n9568;
  assign n9570 = controllable_DEQ & ~n8371;
  assign n9571 = ~n7379 & ~n8040;
  assign n9572 = i_StoB_REQ9 & ~n9571;
  assign n9573 = ~n9083 & ~n9514;
  assign n9574 = ~i_StoB_REQ9 & ~n9573;
  assign n9575 = ~n9572 & ~n9574;
  assign n9576 = controllable_BtoS_ACK9 & ~n9575;
  assign n9577 = ~n9521 & ~n9574;
  assign n9578 = ~controllable_BtoS_ACK9 & ~n9577;
  assign n9579 = ~n9576 & ~n9578;
  assign n9580 = ~controllable_DEQ & ~n9579;
  assign n9581 = ~n9570 & ~n9580;
  assign n9582 = ~i_nEMPTY & ~n9581;
  assign n9583 = ~n9569 & ~n9582;
  assign n9584 = ~i_FULL & ~n9583;
  assign n9585 = ~n9553 & ~n9584;
  assign n9586 = ~i_RtoB_ACK0 & ~n9585;
  assign n9587 = ~n9197 & ~n9586;
  assign n9588 = n6660 & ~n9587;
  assign n9589 = ~controllable_ENQ & ~n8401;
  assign n9590 = ~n7992 & ~n9589;
  assign n9591 = i_StoB_REQ9 & ~n9590;
  assign n9592 = ~n8062 & ~n9591;
  assign n9593 = controllable_BtoS_ACK9 & ~n9592;
  assign n9594 = ~n7588 & ~n9503;
  assign n9595 = n6661 & ~n9594;
  assign n9596 = ~n9505 & ~n9595;
  assign n9597 = i_StoB_REQ11 & ~n9596;
  assign n9598 = n6661 & ~n9502;
  assign n9599 = ~n9510 & ~n9598;
  assign n9600 = ~i_StoB_REQ11 & ~n9599;
  assign n9601 = ~n9597 & ~n9600;
  assign n9602 = controllable_ENQ & ~n9601;
  assign n9603 = ~n9303 & ~n9602;
  assign n9604 = ~controllable_BtoS_ACK9 & ~n9603;
  assign n9605 = ~n9593 & ~n9604;
  assign n9606 = controllable_DEQ & ~n9605;
  assign n9607 = ~controllable_BtoS_ACK9 & ~n9601;
  assign n9608 = ~n8459 & ~n9607;
  assign n9609 = ~controllable_DEQ & ~n9608;
  assign n9610 = ~n9606 & ~n9609;
  assign n9611 = i_nEMPTY & ~n9610;
  assign n9612 = ~controllable_ENQ & ~n9589;
  assign n9613 = i_StoB_REQ9 & ~n9612;
  assign n9614 = ~n9305 & ~n9613;
  assign n9615 = controllable_BtoS_ACK9 & ~n9614;
  assign n9616 = ~controllable_BtoS_ACK9 & ~n9304;
  assign n9617 = ~n9615 & ~n9616;
  assign n9618 = controllable_DEQ & ~n9617;
  assign n9619 = controllable_ENQ & ~n9602;
  assign n9620 = ~controllable_BtoS_ACK9 & ~n9619;
  assign n9621 = ~n8465 & ~n9620;
  assign n9622 = ~controllable_DEQ & ~n9621;
  assign n9623 = ~n9618 & ~n9622;
  assign n9624 = ~i_nEMPTY & ~n9623;
  assign n9625 = ~n9611 & ~n9624;
  assign n9626 = i_FULL & ~n9625;
  assign n9627 = ~n8418 & ~n9593;
  assign n9628 = controllable_DEQ & ~n9627;
  assign n9629 = ~n8459 & ~n9604;
  assign n9630 = ~controllable_DEQ & ~n9629;
  assign n9631 = ~n9628 & ~n9630;
  assign n9632 = i_nEMPTY & ~n9631;
  assign n9633 = controllable_DEQ & ~n8419;
  assign n9634 = ~n7992 & ~n8040;
  assign n9635 = i_StoB_REQ9 & ~n9634;
  assign n9636 = ~n9085 & ~n9635;
  assign n9637 = controllable_BtoS_ACK9 & ~n9636;
  assign n9638 = i_StoB_REQ9 & ~n9603;
  assign n9639 = ~n9083 & ~n9602;
  assign n9640 = ~i_StoB_REQ9 & ~n9639;
  assign n9641 = ~n9638 & ~n9640;
  assign n9642 = ~controllable_BtoS_ACK9 & ~n9641;
  assign n9643 = ~n9637 & ~n9642;
  assign n9644 = ~controllable_DEQ & ~n9643;
  assign n9645 = ~n9633 & ~n9644;
  assign n9646 = ~i_nEMPTY & ~n9645;
  assign n9647 = ~n9632 & ~n9646;
  assign n9648 = ~i_FULL & ~n9647;
  assign n9649 = ~n9626 & ~n9648;
  assign n9650 = ~i_RtoB_ACK0 & ~n9649;
  assign n9651 = ~n9207 & ~n9650;
  assign n9652 = ~n6660 & ~n9651;
  assign n9653 = ~n9588 & ~n9652;
  assign n9654 = n6659 & ~n9653;
  assign n9655 = ~n9331 & ~n9654;
  assign n9656 = ~n6652 & ~n9655;
  assign n9657 = ~n9330 & ~n9656;
  assign n9658 = n6651 & ~n9657;
  assign n9659 = i_RtoB_ACK0 & ~n9203;
  assign n9660 = ~n9586 & ~n9659;
  assign n9661 = n6660 & ~n9660;
  assign n9662 = i_RtoB_ACK0 & ~n9213;
  assign n9663 = ~n9650 & ~n9662;
  assign n9664 = ~n6660 & ~n9663;
  assign n9665 = ~n9661 & ~n9664;
  assign n9666 = ~n6659 & ~n9665;
  assign n9667 = n6659 & ~n9329;
  assign n9668 = ~n9666 & ~n9667;
  assign n9669 = n6652 & ~n9668;
  assign n9670 = ~n9654 & ~n9666;
  assign n9671 = ~n6652 & ~n9670;
  assign n9672 = ~n9669 & ~n9671;
  assign n9673 = ~n6651 & ~n9672;
  assign n9674 = ~n9658 & ~n9673;
  assign n9675 = ~controllable_BtoR_REQ0 & ~n9674;
  assign n9676 = ~n9269 & ~n9675;
  assign n9677 = ~i_RtoB_ACK1 & ~n9676;
  assign n9678 = ~n9224 & ~n9677;
  assign n9679 = ~controllable_BtoR_REQ1 & ~n9678;
  assign n9680 = ~n9143 & ~n9679;
  assign n9681 = n6649 & ~n9680;
  assign n9682 = ~i_FULL & ~n9287;
  assign n9683 = ~n9285 & ~n9682;
  assign n9684 = ~i_RtoB_ACK0 & ~n9683;
  assign n9685 = ~n9197 & ~n9684;
  assign n9686 = n6660 & ~n9685;
  assign n9687 = ~i_FULL & ~n9319;
  assign n9688 = ~n9317 & ~n9687;
  assign n9689 = ~i_RtoB_ACK0 & ~n9688;
  assign n9690 = ~n9207 & ~n9689;
  assign n9691 = ~n6660 & ~n9690;
  assign n9692 = ~n9686 & ~n9691;
  assign n9693 = n6652 & ~n9692;
  assign n9694 = ~n6659 & ~n9692;
  assign n9695 = ~controllable_DEQ & ~n9524;
  assign n9696 = ~n9570 & ~n9695;
  assign n9697 = ~i_nEMPTY & ~n9696;
  assign n9698 = ~n9569 & ~n9697;
  assign n9699 = ~i_FULL & ~n9698;
  assign n9700 = ~n9553 & ~n9699;
  assign n9701 = ~i_RtoB_ACK0 & ~n9700;
  assign n9702 = ~n9197 & ~n9701;
  assign n9703 = n6660 & ~n9702;
  assign n9704 = ~controllable_DEQ & ~n9605;
  assign n9705 = ~n9633 & ~n9704;
  assign n9706 = ~i_nEMPTY & ~n9705;
  assign n9707 = ~n9632 & ~n9706;
  assign n9708 = ~i_FULL & ~n9707;
  assign n9709 = ~n9626 & ~n9708;
  assign n9710 = ~i_RtoB_ACK0 & ~n9709;
  assign n9711 = ~n9207 & ~n9710;
  assign n9712 = ~n6660 & ~n9711;
  assign n9713 = ~n9703 & ~n9712;
  assign n9714 = n6659 & ~n9713;
  assign n9715 = ~n9694 & ~n9714;
  assign n9716 = ~n6652 & ~n9715;
  assign n9717 = ~n9693 & ~n9716;
  assign n9718 = n6651 & ~n9717;
  assign n9719 = ~n9659 & ~n9701;
  assign n9720 = n6660 & ~n9719;
  assign n9721 = ~n9662 & ~n9710;
  assign n9722 = ~n6660 & ~n9721;
  assign n9723 = ~n9720 & ~n9722;
  assign n9724 = ~n6659 & ~n9723;
  assign n9725 = n6659 & ~n9692;
  assign n9726 = ~n9724 & ~n9725;
  assign n9727 = n6652 & ~n9726;
  assign n9728 = ~n9714 & ~n9724;
  assign n9729 = ~n6652 & ~n9728;
  assign n9730 = ~n9727 & ~n9729;
  assign n9731 = ~n6651 & ~n9730;
  assign n9732 = ~n9718 & ~n9731;
  assign n9733 = ~controllable_BtoR_REQ0 & ~n9732;
  assign n9734 = ~n9269 & ~n9733;
  assign n9735 = ~i_RtoB_ACK1 & ~n9734;
  assign n9736 = ~n9224 & ~n9735;
  assign n9737 = ~controllable_BtoR_REQ1 & ~n9736;
  assign n9738 = ~n9143 & ~n9737;
  assign n9739 = ~n6649 & ~n9738;
  assign n9740 = ~n9681 & ~n9739;
  assign n9741 = n6647 & ~n9740;
  assign n9742 = ~i_StoB_REQ9 & ~n8005;
  assign n9743 = controllable_BtoS_ACK9 & ~n9742;
  assign n9744 = n6661 & ~n7185;
  assign n9745 = ~n7188 & ~n9744;
  assign n9746 = ~i_StoB_REQ11 & ~n9745;
  assign n9747 = ~n7998 & ~n9746;
  assign n9748 = controllable_ENQ & ~n9747;
  assign n9749 = controllable_ENQ & ~n9748;
  assign n9750 = i_StoB_REQ9 & ~n9749;
  assign n9751 = ~n8005 & ~n9750;
  assign n9752 = ~controllable_BtoS_ACK9 & ~n9751;
  assign n9753 = ~n9743 & ~n9752;
  assign n9754 = controllable_DEQ & ~n9753;
  assign n9755 = ~i_StoB_REQ9 & ~n8014;
  assign n9756 = controllable_BtoS_ACK9 & ~n9755;
  assign n9757 = i_StoB_REQ9 & ~n9747;
  assign n9758 = ~n8014 & ~n9757;
  assign n9759 = ~controllable_BtoS_ACK9 & ~n9758;
  assign n9760 = ~n9756 & ~n9759;
  assign n9761 = ~controllable_DEQ & ~n9760;
  assign n9762 = ~n9754 & ~n9761;
  assign n9763 = i_nEMPTY & ~n9762;
  assign n9764 = ~controllable_DEQ & ~n9753;
  assign n9765 = ~controllable_DEQ & ~n9764;
  assign n9766 = ~i_nEMPTY & ~n9765;
  assign n9767 = ~n9763 & ~n9766;
  assign n9768 = i_RtoB_ACK0 & ~n9767;
  assign n9769 = ~n8033 & ~n8056;
  assign n9770 = controllable_BtoS_ACK9 & ~n9769;
  assign n9771 = ~controllable_ENQ & ~n9747;
  assign n9772 = ~n8050 & ~n9771;
  assign n9773 = i_StoB_REQ9 & ~n9772;
  assign n9774 = ~n8056 & ~n9773;
  assign n9775 = ~controllable_BtoS_ACK9 & ~n9774;
  assign n9776 = ~n9770 & ~n9775;
  assign n9777 = controllable_DEQ & ~n9776;
  assign n9778 = ~i_StoB_REQ9 & ~n8049;
  assign n9779 = ~n8061 & ~n9778;
  assign n9780 = controllable_BtoS_ACK9 & ~n9779;
  assign n9781 = ~n8065 & ~n9780;
  assign n9782 = ~controllable_DEQ & ~n9781;
  assign n9783 = ~n9777 & ~n9782;
  assign n9784 = i_nEMPTY & ~n9783;
  assign n9785 = ~i_StoB_REQ9 & ~n8077;
  assign n9786 = controllable_BtoS_ACK9 & ~n9785;
  assign n9787 = ~controllable_ENQ & ~n9771;
  assign n9788 = i_StoB_REQ9 & ~n9787;
  assign n9789 = ~n8077 & ~n9788;
  assign n9790 = ~controllable_BtoS_ACK9 & ~n9789;
  assign n9791 = ~n9786 & ~n9790;
  assign n9792 = controllable_DEQ & ~n9791;
  assign n9793 = ~i_StoB_REQ9 & ~n8086;
  assign n9794 = ~n8033 & ~n9793;
  assign n9795 = controllable_BtoS_ACK9 & ~n9794;
  assign n9796 = ~n8087 & ~n9795;
  assign n9797 = ~controllable_DEQ & ~n9796;
  assign n9798 = ~n9792 & ~n9797;
  assign n9799 = ~i_nEMPTY & ~n9798;
  assign n9800 = ~n9784 & ~n9799;
  assign n9801 = i_FULL & ~n9800;
  assign n9802 = ~n8033 & ~n8114;
  assign n9803 = controllable_BtoS_ACK9 & ~n9802;
  assign n9804 = ~n8112 & ~n9771;
  assign n9805 = i_StoB_REQ9 & ~n9804;
  assign n9806 = ~n8114 & ~n9805;
  assign n9807 = ~controllable_BtoS_ACK9 & ~n9806;
  assign n9808 = ~n9803 & ~n9807;
  assign n9809 = controllable_DEQ & ~n9808;
  assign n9810 = ~n8061 & ~n8124;
  assign n9811 = controllable_BtoS_ACK9 & ~n9810;
  assign n9812 = ~controllable_BtoS_ACK9 & ~n8123;
  assign n9813 = ~n9811 & ~n9812;
  assign n9814 = ~controllable_DEQ & ~n9813;
  assign n9815 = ~n9809 & ~n9814;
  assign n9816 = i_nEMPTY & ~n9815;
  assign n9817 = controllable_DEQ & ~n9760;
  assign n9818 = ~controllable_DEQ & ~n9776;
  assign n9819 = ~n9817 & ~n9818;
  assign n9820 = ~i_nEMPTY & ~n9819;
  assign n9821 = ~n9816 & ~n9820;
  assign n9822 = ~i_FULL & ~n9821;
  assign n9823 = ~n9801 & ~n9822;
  assign n9824 = ~i_RtoB_ACK0 & ~n9823;
  assign n9825 = ~n9768 & ~n9824;
  assign n9826 = n6660 & ~n9825;
  assign n9827 = ~n8140 & ~n9826;
  assign n9828 = ~n6659 & ~n9827;
  assign n9829 = ~n8149 & ~n9827;
  assign n9830 = ~n8149 & ~n9829;
  assign n9831 = n6659 & ~n9830;
  assign n9832 = ~n9828 & ~n9831;
  assign n9833 = n6652 & ~n9832;
  assign n9834 = i_StoB_REQ11 & ~n8226;
  assign n9835 = i_StoB_REQ10 & ~n8216;
  assign n9836 = i_StoB_REQ8 & ~n8208;
  assign n9837 = i_StoB_REQ6 & ~n8189;
  assign n9838 = i_StoB_REQ5 & ~n8181;
  assign n9839 = i_StoB_REQ4 & ~n8248;
  assign n9840 = i_StoB_REQ3 & ~n8168;
  assign n9841 = i_StoB_REQ2 & ~n8160;
  assign n9842 = ~n8265 & ~n8715;
  assign n9843 = n6670 & ~n9842;
  assign n9844 = ~n8273 & ~n9843;
  assign n9845 = n6669 & ~n9844;
  assign n9846 = ~n7407 & ~n9845;
  assign n9847 = ~i_StoB_REQ2 & ~n9846;
  assign n9848 = ~n9841 & ~n9847;
  assign n9849 = controllable_BtoS_ACK2 & ~n9848;
  assign n9850 = ~n8280 & ~n9847;
  assign n9851 = ~controllable_BtoS_ACK2 & ~n9850;
  assign n9852 = ~n9849 & ~n9851;
  assign n9853 = n6668 & ~n9852;
  assign n9854 = ~n7425 & ~n9853;
  assign n9855 = ~i_StoB_REQ3 & ~n9854;
  assign n9856 = ~n9840 & ~n9855;
  assign n9857 = controllable_BtoS_ACK3 & ~n9856;
  assign n9858 = ~n8289 & ~n9855;
  assign n9859 = ~controllable_BtoS_ACK3 & ~n9858;
  assign n9860 = ~n9857 & ~n9859;
  assign n9861 = n6667 & ~n9860;
  assign n9862 = ~n8294 & ~n9861;
  assign n9863 = ~i_StoB_REQ4 & ~n9862;
  assign n9864 = ~n9839 & ~n9863;
  assign n9865 = n6666 & ~n9864;
  assign n9866 = ~n7477 & ~n9865;
  assign n9867 = ~i_StoB_REQ5 & ~n9866;
  assign n9868 = ~n9838 & ~n9867;
  assign n9869 = controllable_BtoS_ACK5 & ~n9868;
  assign n9870 = ~n8303 & ~n9867;
  assign n9871 = ~controllable_BtoS_ACK5 & ~n9870;
  assign n9872 = ~n9869 & ~n9871;
  assign n9873 = n6665 & ~n9872;
  assign n9874 = ~n7497 & ~n9873;
  assign n9875 = ~i_StoB_REQ6 & ~n9874;
  assign n9876 = ~n9837 & ~n9875;
  assign n9877 = controllable_BtoS_ACK6 & ~n9876;
  assign n9878 = ~n8312 & ~n9875;
  assign n9879 = ~controllable_BtoS_ACK6 & ~n9878;
  assign n9880 = ~n9877 & ~n9879;
  assign n9881 = ~i_StoB_REQ7 & ~n9880;
  assign n9882 = ~n8319 & ~n9881;
  assign n9883 = n6664 & ~n9882;
  assign n9884 = ~n8321 & ~n9883;
  assign n9885 = controllable_BtoS_ACK7 & ~n9884;
  assign n9886 = ~n8324 & ~n9881;
  assign n9887 = n6664 & ~n9886;
  assign n9888 = ~n8327 & ~n9887;
  assign n9889 = ~controllable_BtoS_ACK7 & ~n9888;
  assign n9890 = ~n9885 & ~n9889;
  assign n9891 = n6663 & ~n9890;
  assign n9892 = ~n7546 & ~n9891;
  assign n9893 = ~i_StoB_REQ8 & ~n9892;
  assign n9894 = ~n9836 & ~n9893;
  assign n9895 = controllable_BtoS_ACK8 & ~n9894;
  assign n9896 = ~n8336 & ~n9893;
  assign n9897 = ~controllable_BtoS_ACK8 & ~n9896;
  assign n9898 = ~n9895 & ~n9897;
  assign n9899 = n6662 & ~n9898;
  assign n9900 = ~n7568 & ~n9899;
  assign n9901 = ~i_StoB_REQ10 & ~n9900;
  assign n9902 = ~n9835 & ~n9901;
  assign n9903 = controllable_BtoS_ACK10 & ~n9902;
  assign n9904 = ~n8345 & ~n9901;
  assign n9905 = ~controllable_BtoS_ACK10 & ~n9904;
  assign n9906 = ~n9903 & ~n9905;
  assign n9907 = n6661 & ~n9906;
  assign n9908 = ~n8350 & ~n9907;
  assign n9909 = ~i_StoB_REQ11 & ~n9908;
  assign n9910 = ~n9834 & ~n9909;
  assign n9911 = controllable_ENQ & ~n9910;
  assign n9912 = ~controllable_BtoS_ACK11 & ~n8224;
  assign n9913 = ~controllable_BtoS_ACK11 & ~n9912;
  assign n9914 = n6661 & ~n9913;
  assign n9915 = ~n6921 & ~n9914;
  assign n9916 = i_StoB_REQ11 & ~n9915;
  assign n9917 = ~controllable_BtoS_ACK4 & ~n8176;
  assign n9918 = ~controllable_BtoS_ACK4 & ~n9917;
  assign n9919 = n6667 & ~n9918;
  assign n9920 = ~n6755 & ~n9919;
  assign n9921 = i_StoB_REQ4 & ~n9920;
  assign n9922 = i_StoB_REQ1 & ~n8268;
  assign n9923 = ~controllable_BtoS_ACK1 & ~n9922;
  assign n9924 = ~controllable_BtoS_ACK1 & ~n9923;
  assign n9925 = n6671 & ~n9924;
  assign n9926 = ~n6941 & ~n9925;
  assign n9927 = n6670 & ~n9926;
  assign n9928 = ~n6670 & ~n6930;
  assign n9929 = ~n9927 & ~n9928;
  assign n9930 = n6669 & ~n9929;
  assign n9931 = ~n6946 & ~n9930;
  assign n9932 = ~i_StoB_REQ2 & ~n9931;
  assign n9933 = ~i_StoB_REQ2 & ~n9932;
  assign n9934 = controllable_BtoS_ACK2 & ~n9933;
  assign n9935 = i_StoB_REQ2 & ~n8162;
  assign n9936 = ~n9932 & ~n9935;
  assign n9937 = ~controllable_BtoS_ACK2 & ~n9936;
  assign n9938 = ~n9934 & ~n9937;
  assign n9939 = n6668 & ~n9938;
  assign n9940 = ~n6968 & ~n9939;
  assign n9941 = ~i_StoB_REQ3 & ~n9940;
  assign n9942 = ~i_StoB_REQ3 & ~n9941;
  assign n9943 = controllable_BtoS_ACK3 & ~n9942;
  assign n9944 = i_StoB_REQ3 & ~n8170;
  assign n9945 = ~n9941 & ~n9944;
  assign n9946 = ~controllable_BtoS_ACK3 & ~n9945;
  assign n9947 = ~n9943 & ~n9946;
  assign n9948 = n6667 & ~n9947;
  assign n9949 = ~n6667 & ~n6995;
  assign n9950 = ~n9948 & ~n9949;
  assign n9951 = ~i_StoB_REQ4 & ~n9950;
  assign n9952 = ~n9921 & ~n9951;
  assign n9953 = n6666 & ~n9952;
  assign n9954 = ~n7015 & ~n9953;
  assign n9955 = ~i_StoB_REQ5 & ~n9954;
  assign n9956 = ~i_StoB_REQ5 & ~n9955;
  assign n9957 = controllable_BtoS_ACK5 & ~n9956;
  assign n9958 = i_StoB_REQ5 & ~n8183;
  assign n9959 = ~n9955 & ~n9958;
  assign n9960 = ~controllable_BtoS_ACK5 & ~n9959;
  assign n9961 = ~n9957 & ~n9960;
  assign n9962 = n6665 & ~n9961;
  assign n9963 = ~n7038 & ~n9962;
  assign n9964 = ~i_StoB_REQ6 & ~n9963;
  assign n9965 = ~i_StoB_REQ6 & ~n9964;
  assign n9966 = controllable_BtoS_ACK6 & ~n9965;
  assign n9967 = i_StoB_REQ6 & ~n8191;
  assign n9968 = ~n9964 & ~n9967;
  assign n9969 = ~controllable_BtoS_ACK6 & ~n9968;
  assign n9970 = ~n9966 & ~n9969;
  assign n9971 = ~i_StoB_REQ7 & ~n9970;
  assign n9972 = ~i_StoB_REQ7 & ~n9971;
  assign n9973 = n6664 & ~n9972;
  assign n9974 = ~n7070 & ~n9973;
  assign n9975 = controllable_BtoS_ACK7 & ~n9974;
  assign n9976 = ~n8319 & ~n9971;
  assign n9977 = n6664 & ~n9976;
  assign n9978 = ~n6664 & ~n7093;
  assign n9979 = ~n9977 & ~n9978;
  assign n9980 = ~controllable_BtoS_ACK7 & ~n9979;
  assign n9981 = ~n9975 & ~n9980;
  assign n9982 = n6663 & ~n9981;
  assign n9983 = ~n7096 & ~n9982;
  assign n9984 = ~i_StoB_REQ8 & ~n9983;
  assign n9985 = ~i_StoB_REQ8 & ~n9984;
  assign n9986 = controllable_BtoS_ACK8 & ~n9985;
  assign n9987 = i_StoB_REQ8 & ~n8210;
  assign n9988 = ~n9984 & ~n9987;
  assign n9989 = ~controllable_BtoS_ACK8 & ~n9988;
  assign n9990 = ~n9986 & ~n9989;
  assign n9991 = n6662 & ~n9990;
  assign n9992 = ~n7125 & ~n9991;
  assign n9993 = ~i_StoB_REQ10 & ~n9992;
  assign n9994 = ~i_StoB_REQ10 & ~n9993;
  assign n9995 = controllable_BtoS_ACK10 & ~n9994;
  assign n9996 = i_StoB_REQ10 & ~n8218;
  assign n9997 = ~n9993 & ~n9996;
  assign n9998 = ~controllable_BtoS_ACK10 & ~n9997;
  assign n9999 = ~n9995 & ~n9998;
  assign n10000 = n6661 & ~n9999;
  assign n10001 = ~n6661 & ~n7152;
  assign n10002 = ~n10000 & ~n10001;
  assign n10003 = ~i_StoB_REQ11 & ~n10002;
  assign n10004 = ~n9916 & ~n10003;
  assign n10005 = ~controllable_ENQ & ~n10004;
  assign n10006 = ~n9911 & ~n10005;
  assign n10007 = ~i_StoB_REQ9 & ~n10006;
  assign n10008 = ~n8404 & ~n10007;
  assign n10009 = controllable_BtoS_ACK9 & ~n10008;
  assign n10010 = ~n8039 & ~n9589;
  assign n10011 = i_StoB_REQ9 & ~n10010;
  assign n10012 = ~n10007 & ~n10011;
  assign n10013 = ~controllable_BtoS_ACK9 & ~n10012;
  assign n10014 = ~n10009 & ~n10013;
  assign n10015 = controllable_DEQ & ~n10014;
  assign n10016 = ~n6671 & ~n8156;
  assign n10017 = n6670 & ~n10016;
  assign n10018 = ~n8159 & ~n10017;
  assign n10019 = n6669 & ~n10018;
  assign n10020 = ~n6702 & ~n10019;
  assign n10021 = ~i_StoB_REQ2 & ~n10020;
  assign n10022 = ~i_StoB_REQ2 & ~n10021;
  assign n10023 = controllable_BtoS_ACK2 & ~n10022;
  assign n10024 = ~controllable_BtoS_ACK2 & ~n10020;
  assign n10025 = ~n10023 & ~n10024;
  assign n10026 = n6668 & ~n10025;
  assign n10027 = ~n6723 & ~n10026;
  assign n10028 = ~i_StoB_REQ3 & ~n10027;
  assign n10029 = ~i_StoB_REQ3 & ~n10028;
  assign n10030 = controllable_BtoS_ACK3 & ~n10029;
  assign n10031 = ~controllable_BtoS_ACK3 & ~n10027;
  assign n10032 = ~n10030 & ~n10031;
  assign n10033 = ~controllable_BtoS_ACK4 & ~n10032;
  assign n10034 = ~controllable_BtoS_ACK4 & ~n10033;
  assign n10035 = n6667 & ~n10034;
  assign n10036 = ~n6755 & ~n10035;
  assign n10037 = i_StoB_REQ4 & ~n10036;
  assign n10038 = n6667 & ~n10032;
  assign n10039 = ~n8178 & ~n10038;
  assign n10040 = ~i_StoB_REQ4 & ~n10039;
  assign n10041 = ~n10037 & ~n10040;
  assign n10042 = n6666 & ~n10041;
  assign n10043 = ~n6780 & ~n10042;
  assign n10044 = ~i_StoB_REQ5 & ~n10043;
  assign n10045 = ~i_StoB_REQ5 & ~n10044;
  assign n10046 = controllable_BtoS_ACK5 & ~n10045;
  assign n10047 = ~controllable_BtoS_ACK5 & ~n10043;
  assign n10048 = ~n10046 & ~n10047;
  assign n10049 = n6665 & ~n10048;
  assign n10050 = ~n6806 & ~n10049;
  assign n10051 = ~i_StoB_REQ6 & ~n10050;
  assign n10052 = ~i_StoB_REQ6 & ~n10051;
  assign n10053 = controllable_BtoS_ACK6 & ~n10052;
  assign n10054 = ~controllable_BtoS_ACK6 & ~n10050;
  assign n10055 = ~n10053 & ~n10054;
  assign n10056 = ~i_StoB_REQ7 & ~n10055;
  assign n10057 = ~i_StoB_REQ7 & ~n10056;
  assign n10058 = n6664 & ~n10057;
  assign n10059 = ~n6838 & ~n10058;
  assign n10060 = controllable_BtoS_ACK7 & ~n10059;
  assign n10061 = n6664 & ~n10055;
  assign n10062 = ~n8205 & ~n10061;
  assign n10063 = ~controllable_BtoS_ACK7 & ~n10062;
  assign n10064 = ~n10060 & ~n10063;
  assign n10065 = n6663 & ~n10064;
  assign n10066 = ~n6863 & ~n10065;
  assign n10067 = ~i_StoB_REQ8 & ~n10066;
  assign n10068 = ~i_StoB_REQ8 & ~n10067;
  assign n10069 = controllable_BtoS_ACK8 & ~n10068;
  assign n10070 = ~controllable_BtoS_ACK8 & ~n10066;
  assign n10071 = ~n10069 & ~n10070;
  assign n10072 = n6662 & ~n10071;
  assign n10073 = ~n6889 & ~n10072;
  assign n10074 = ~i_StoB_REQ10 & ~n10073;
  assign n10075 = ~i_StoB_REQ10 & ~n10074;
  assign n10076 = controllable_BtoS_ACK10 & ~n10075;
  assign n10077 = ~controllable_BtoS_ACK10 & ~n10073;
  assign n10078 = ~n10076 & ~n10077;
  assign n10079 = ~controllable_BtoS_ACK11 & ~n10078;
  assign n10080 = ~controllable_BtoS_ACK11 & ~n10079;
  assign n10081 = n6661 & ~n10080;
  assign n10082 = ~n6921 & ~n10081;
  assign n10083 = i_StoB_REQ11 & ~n10082;
  assign n10084 = n6661 & ~n10078;
  assign n10085 = ~n8398 & ~n10084;
  assign n10086 = ~i_StoB_REQ11 & ~n10085;
  assign n10087 = ~n10083 & ~n10086;
  assign n10088 = i_StoB_REQ9 & ~n10087;
  assign n10089 = controllable_BtoS_ACK11 & ~n10078;
  assign n10090 = i_StoB_REQ10 & ~n10073;
  assign n10091 = i_StoB_REQ8 & ~n10066;
  assign n10092 = i_StoB_REQ7 & ~n10055;
  assign n10093 = i_StoB_REQ6 & ~n10050;
  assign n10094 = i_StoB_REQ5 & ~n10043;
  assign n10095 = controllable_BtoS_ACK4 & ~n10032;
  assign n10096 = i_StoB_REQ3 & ~n10027;
  assign n10097 = i_StoB_REQ2 & ~n10020;
  assign n10098 = ~n6671 & ~n8271;
  assign n10099 = n6670 & ~n10098;
  assign n10100 = ~n6670 & n7391;
  assign n10101 = ~n10099 & ~n10100;
  assign n10102 = n6669 & ~n10101;
  assign n10103 = ~n7407 & ~n10102;
  assign n10104 = ~i_StoB_REQ2 & ~n10103;
  assign n10105 = ~n10097 & ~n10104;
  assign n10106 = controllable_BtoS_ACK2 & ~n10105;
  assign n10107 = ~controllable_BtoS_ACK2 & ~n10103;
  assign n10108 = ~n10106 & ~n10107;
  assign n10109 = n6668 & ~n10108;
  assign n10110 = ~n7425 & ~n10109;
  assign n10111 = ~i_StoB_REQ3 & ~n10110;
  assign n10112 = ~n10096 & ~n10111;
  assign n10113 = controllable_BtoS_ACK3 & ~n10112;
  assign n10114 = ~controllable_BtoS_ACK3 & ~n10110;
  assign n10115 = ~n10113 & ~n10114;
  assign n10116 = ~controllable_BtoS_ACK4 & ~n10115;
  assign n10117 = ~n10095 & ~n10116;
  assign n10118 = n6667 & ~n10117;
  assign n10119 = ~n6667 & ~n7473;
  assign n10120 = ~n10118 & ~n10119;
  assign n10121 = i_StoB_REQ4 & ~n10120;
  assign n10122 = n6667 & ~n10115;
  assign n10123 = ~n8294 & ~n10122;
  assign n10124 = ~i_StoB_REQ4 & ~n10123;
  assign n10125 = ~n10121 & ~n10124;
  assign n10126 = n6666 & ~n10125;
  assign n10127 = ~n7477 & ~n10126;
  assign n10128 = ~i_StoB_REQ5 & ~n10127;
  assign n10129 = ~n10094 & ~n10128;
  assign n10130 = controllable_BtoS_ACK5 & ~n10129;
  assign n10131 = ~controllable_BtoS_ACK5 & ~n10127;
  assign n10132 = ~n10130 & ~n10131;
  assign n10133 = n6665 & ~n10132;
  assign n10134 = ~n7497 & ~n10133;
  assign n10135 = ~i_StoB_REQ6 & ~n10134;
  assign n10136 = ~n10093 & ~n10135;
  assign n10137 = controllable_BtoS_ACK6 & ~n10136;
  assign n10138 = ~controllable_BtoS_ACK6 & ~n10134;
  assign n10139 = ~n10137 & ~n10138;
  assign n10140 = ~i_StoB_REQ7 & ~n10139;
  assign n10141 = ~n10092 & ~n10140;
  assign n10142 = n6664 & ~n10141;
  assign n10143 = ~n9443 & ~n10142;
  assign n10144 = controllable_BtoS_ACK7 & ~n10143;
  assign n10145 = n6664 & ~n10139;
  assign n10146 = ~n8327 & ~n10145;
  assign n10147 = ~controllable_BtoS_ACK7 & ~n10146;
  assign n10148 = ~n10144 & ~n10147;
  assign n10149 = n6663 & ~n10148;
  assign n10150 = ~n7546 & ~n10149;
  assign n10151 = ~i_StoB_REQ8 & ~n10150;
  assign n10152 = ~n10091 & ~n10151;
  assign n10153 = controllable_BtoS_ACK8 & ~n10152;
  assign n10154 = ~controllable_BtoS_ACK8 & ~n10150;
  assign n10155 = ~n10153 & ~n10154;
  assign n10156 = n6662 & ~n10155;
  assign n10157 = ~n7568 & ~n10156;
  assign n10158 = ~i_StoB_REQ10 & ~n10157;
  assign n10159 = ~n10090 & ~n10158;
  assign n10160 = controllable_BtoS_ACK10 & ~n10159;
  assign n10161 = ~controllable_BtoS_ACK10 & ~n10157;
  assign n10162 = ~n10160 & ~n10161;
  assign n10163 = ~controllable_BtoS_ACK11 & ~n10162;
  assign n10164 = ~n10089 & ~n10163;
  assign n10165 = n6661 & ~n10164;
  assign n10166 = ~n8227 & ~n10165;
  assign n10167 = i_StoB_REQ11 & ~n10166;
  assign n10168 = ~n8231 & ~n10072;
  assign n10169 = i_StoB_REQ10 & ~n10168;
  assign n10170 = ~n8235 & ~n10065;
  assign n10171 = i_StoB_REQ8 & ~n10170;
  assign n10172 = ~n8239 & ~n10049;
  assign n10173 = i_StoB_REQ6 & ~n10172;
  assign n10174 = ~n8243 & ~n10042;
  assign n10175 = i_StoB_REQ5 & ~n10174;
  assign n10176 = ~n8249 & ~n10118;
  assign n10177 = i_StoB_REQ4 & ~n10176;
  assign n10178 = ~n8253 & ~n10026;
  assign n10179 = i_StoB_REQ3 & ~n10178;
  assign n10180 = ~n8257 & ~n10019;
  assign n10181 = i_StoB_REQ2 & ~n10180;
  assign n10182 = ~n6671 & ~n8265;
  assign n10183 = n6670 & ~n10182;
  assign n10184 = ~n8273 & ~n10183;
  assign n10185 = n6669 & ~n10184;
  assign n10186 = ~n7407 & ~n10185;
  assign n10187 = ~i_StoB_REQ2 & ~n10186;
  assign n10188 = ~n10181 & ~n10187;
  assign n10189 = controllable_BtoS_ACK2 & ~n10188;
  assign n10190 = i_StoB_REQ2 & ~n10103;
  assign n10191 = ~n10187 & ~n10190;
  assign n10192 = ~controllable_BtoS_ACK2 & ~n10191;
  assign n10193 = ~n10189 & ~n10192;
  assign n10194 = n6668 & ~n10193;
  assign n10195 = ~n7425 & ~n10194;
  assign n10196 = ~i_StoB_REQ3 & ~n10195;
  assign n10197 = ~n10179 & ~n10196;
  assign n10198 = controllable_BtoS_ACK3 & ~n10197;
  assign n10199 = i_StoB_REQ3 & ~n10110;
  assign n10200 = ~n10196 & ~n10199;
  assign n10201 = ~controllable_BtoS_ACK3 & ~n10200;
  assign n10202 = ~n10198 & ~n10201;
  assign n10203 = n6667 & ~n10202;
  assign n10204 = ~n8294 & ~n10203;
  assign n10205 = ~i_StoB_REQ4 & ~n10204;
  assign n10206 = ~n10177 & ~n10205;
  assign n10207 = n6666 & ~n10206;
  assign n10208 = ~n7477 & ~n10207;
  assign n10209 = ~i_StoB_REQ5 & ~n10208;
  assign n10210 = ~n10175 & ~n10209;
  assign n10211 = controllable_BtoS_ACK5 & ~n10210;
  assign n10212 = i_StoB_REQ5 & ~n10127;
  assign n10213 = ~n10209 & ~n10212;
  assign n10214 = ~controllable_BtoS_ACK5 & ~n10213;
  assign n10215 = ~n10211 & ~n10214;
  assign n10216 = n6665 & ~n10215;
  assign n10217 = ~n7497 & ~n10216;
  assign n10218 = ~i_StoB_REQ6 & ~n10217;
  assign n10219 = ~n10173 & ~n10218;
  assign n10220 = controllable_BtoS_ACK6 & ~n10219;
  assign n10221 = i_StoB_REQ6 & ~n10134;
  assign n10222 = ~n10218 & ~n10221;
  assign n10223 = ~controllable_BtoS_ACK6 & ~n10222;
  assign n10224 = ~n10220 & ~n10223;
  assign n10225 = ~i_StoB_REQ7 & ~n10224;
  assign n10226 = ~n10092 & ~n10225;
  assign n10227 = n6664 & ~n10226;
  assign n10228 = ~n8321 & ~n10227;
  assign n10229 = controllable_BtoS_ACK7 & ~n10228;
  assign n10230 = i_StoB_REQ7 & ~n10139;
  assign n10231 = ~n10225 & ~n10230;
  assign n10232 = n6664 & ~n10231;
  assign n10233 = ~n8327 & ~n10232;
  assign n10234 = ~controllable_BtoS_ACK7 & ~n10233;
  assign n10235 = ~n10229 & ~n10234;
  assign n10236 = n6663 & ~n10235;
  assign n10237 = ~n7546 & ~n10236;
  assign n10238 = ~i_StoB_REQ8 & ~n10237;
  assign n10239 = ~n10171 & ~n10238;
  assign n10240 = controllable_BtoS_ACK8 & ~n10239;
  assign n10241 = i_StoB_REQ8 & ~n10150;
  assign n10242 = ~n10238 & ~n10241;
  assign n10243 = ~controllable_BtoS_ACK8 & ~n10242;
  assign n10244 = ~n10240 & ~n10243;
  assign n10245 = n6662 & ~n10244;
  assign n10246 = ~n7568 & ~n10245;
  assign n10247 = ~i_StoB_REQ10 & ~n10246;
  assign n10248 = ~n10169 & ~n10247;
  assign n10249 = controllable_BtoS_ACK10 & ~n10248;
  assign n10250 = i_StoB_REQ10 & ~n10157;
  assign n10251 = ~n10247 & ~n10250;
  assign n10252 = ~controllable_BtoS_ACK10 & ~n10251;
  assign n10253 = ~n10249 & ~n10252;
  assign n10254 = n6661 & ~n10253;
  assign n10255 = ~n8350 & ~n10254;
  assign n10256 = ~i_StoB_REQ11 & ~n10255;
  assign n10257 = ~n10167 & ~n10256;
  assign n10258 = ~i_StoB_REQ9 & ~n10257;
  assign n10259 = ~n10088 & ~n10258;
  assign n10260 = controllable_BtoS_ACK9 & ~n10259;
  assign n10261 = ~n6661 & ~n8035;
  assign n10262 = ~n10165 & ~n10261;
  assign n10263 = i_StoB_REQ11 & ~n10262;
  assign n10264 = n6661 & ~n10162;
  assign n10265 = ~n8350 & ~n10264;
  assign n10266 = ~i_StoB_REQ11 & ~n10265;
  assign n10267 = ~n10263 & ~n10266;
  assign n10268 = i_StoB_REQ9 & ~n10267;
  assign n10269 = ~n10258 & ~n10268;
  assign n10270 = ~controllable_BtoS_ACK9 & ~n10269;
  assign n10271 = ~n10260 & ~n10270;
  assign n10272 = ~controllable_DEQ & ~n10271;
  assign n10273 = ~n10015 & ~n10272;
  assign n10274 = i_nEMPTY & ~n10273;
  assign n10275 = ~controllable_ENQ & ~n10005;
  assign n10276 = ~i_StoB_REQ9 & ~n10275;
  assign n10277 = ~i_StoB_REQ9 & ~n10276;
  assign n10278 = controllable_BtoS_ACK9 & ~n10277;
  assign n10279 = ~n9613 & ~n10276;
  assign n10280 = ~controllable_BtoS_ACK9 & ~n10279;
  assign n10281 = ~n10278 & ~n10280;
  assign n10282 = controllable_DEQ & ~n10281;
  assign n10283 = controllable_ENQ & ~n10087;
  assign n10284 = controllable_ENQ & ~n10283;
  assign n10285 = i_StoB_REQ9 & ~n10284;
  assign n10286 = controllable_ENQ & ~n10257;
  assign n10287 = controllable_ENQ & ~n10286;
  assign n10288 = ~i_StoB_REQ9 & ~n10287;
  assign n10289 = ~n10285 & ~n10288;
  assign n10290 = controllable_BtoS_ACK9 & ~n10289;
  assign n10291 = controllable_ENQ & ~n10267;
  assign n10292 = controllable_ENQ & ~n10291;
  assign n10293 = i_StoB_REQ9 & ~n10292;
  assign n10294 = ~n10288 & ~n10293;
  assign n10295 = ~controllable_BtoS_ACK9 & ~n10294;
  assign n10296 = ~n10290 & ~n10295;
  assign n10297 = ~controllable_DEQ & ~n10296;
  assign n10298 = ~n10282 & ~n10297;
  assign n10299 = ~i_nEMPTY & ~n10298;
  assign n10300 = ~n10274 & ~n10299;
  assign n10301 = i_FULL & ~n10300;
  assign n10302 = ~i_StoB_REQ9 & ~n10004;
  assign n10303 = ~i_StoB_REQ9 & ~n10302;
  assign n10304 = controllable_BtoS_ACK9 & ~n10303;
  assign n10305 = ~n8415 & ~n10302;
  assign n10306 = ~controllable_BtoS_ACK9 & ~n10305;
  assign n10307 = ~n10304 & ~n10306;
  assign n10308 = controllable_DEQ & ~n10307;
  assign n10309 = ~n8054 & ~n10286;
  assign n10310 = ~i_StoB_REQ9 & ~n10309;
  assign n10311 = ~n10285 & ~n10310;
  assign n10312 = controllable_BtoS_ACK9 & ~n10311;
  assign n10313 = ~n9771 & ~n10291;
  assign n10314 = i_StoB_REQ9 & ~n10313;
  assign n10315 = ~n10310 & ~n10314;
  assign n10316 = ~controllable_BtoS_ACK9 & ~n10315;
  assign n10317 = ~n10312 & ~n10316;
  assign n10318 = ~controllable_DEQ & ~n10317;
  assign n10319 = ~n10308 & ~n10318;
  assign n10320 = ~i_nEMPTY & ~n10319;
  assign n10321 = ~n10274 & ~n10320;
  assign n10322 = ~i_FULL & ~n10321;
  assign n10323 = ~n10301 & ~n10322;
  assign n10324 = ~i_RtoB_ACK0 & ~n10323;
  assign n10325 = ~n9768 & ~n10324;
  assign n10326 = n6660 & ~n10325;
  assign n10327 = ~n8042 & ~n8408;
  assign n10328 = ~controllable_BtoS_ACK9 & ~n10327;
  assign n10329 = ~n8406 & ~n10328;
  assign n10330 = controllable_DEQ & ~n10329;
  assign n10331 = ~n8420 & ~n10330;
  assign n10332 = i_nEMPTY & ~n10331;
  assign n10333 = ~n8071 & ~n8075;
  assign n10334 = ~controllable_BtoS_ACK9 & ~n10333;
  assign n10335 = ~n8073 & ~n10334;
  assign n10336 = controllable_DEQ & ~n10335;
  assign n10337 = ~n8427 & ~n10336;
  assign n10338 = ~i_nEMPTY & ~n10337;
  assign n10339 = ~n10332 & ~n10338;
  assign n10340 = i_FULL & ~n10339;
  assign n10341 = ~n8010 & ~n8013;
  assign n10342 = ~controllable_BtoS_ACK9 & ~n10341;
  assign n10343 = ~n8012 & ~n10342;
  assign n10344 = controllable_DEQ & ~n10343;
  assign n10345 = ~n8432 & ~n10344;
  assign n10346 = ~i_nEMPTY & ~n10345;
  assign n10347 = ~n10332 & ~n10346;
  assign n10348 = ~i_FULL & ~n10347;
  assign n10349 = ~n10340 & ~n10348;
  assign n10350 = ~i_RtoB_ACK0 & ~n10349;
  assign n10351 = ~n8025 & ~n10350;
  assign n10352 = ~n6660 & ~n10351;
  assign n10353 = ~n10326 & ~n10352;
  assign n10354 = ~n6659 & ~n10353;
  assign n10355 = ~n8149 & ~n10353;
  assign n10356 = ~n8149 & ~n10355;
  assign n10357 = n6659 & ~n10356;
  assign n10358 = ~n10354 & ~n10357;
  assign n10359 = ~n6652 & ~n10358;
  assign n10360 = ~n9833 & ~n10359;
  assign n10361 = n6651 & ~n10360;
  assign n10362 = ~n7987 & ~n7994;
  assign n10363 = ~controllable_BtoS_ACK9 & ~n10362;
  assign n10364 = ~n7989 & ~n10363;
  assign n10365 = controllable_DEQ & ~n10364;
  assign n10366 = ~n9761 & ~n10365;
  assign n10367 = i_nEMPTY & ~n10366;
  assign n10368 = ~n9766 & ~n10367;
  assign n10369 = i_RtoB_ACK0 & ~n10368;
  assign n10370 = ~n8482 & ~n10328;
  assign n10371 = controllable_DEQ & ~n10370;
  assign n10372 = ~i_StoB_REQ9 & ~n10267;
  assign n10373 = ~n10088 & ~n10372;
  assign n10374 = controllable_BtoS_ACK9 & ~n10373;
  assign n10375 = ~controllable_BtoS_ACK9 & ~n10267;
  assign n10376 = ~n10374 & ~n10375;
  assign n10377 = ~controllable_DEQ & ~n10376;
  assign n10378 = ~n10371 & ~n10377;
  assign n10379 = i_nEMPTY & ~n10378;
  assign n10380 = ~i_StoB_REQ9 & ~n10292;
  assign n10381 = ~n10285 & ~n10380;
  assign n10382 = controllable_BtoS_ACK9 & ~n10381;
  assign n10383 = ~controllable_BtoS_ACK9 & ~n10292;
  assign n10384 = ~n10382 & ~n10383;
  assign n10385 = ~controllable_DEQ & ~n10384;
  assign n10386 = ~n10336 & ~n10385;
  assign n10387 = ~i_nEMPTY & ~n10386;
  assign n10388 = ~n10379 & ~n10387;
  assign n10389 = i_FULL & ~n10388;
  assign n10390 = ~n8054 & ~n10291;
  assign n10391 = ~i_StoB_REQ9 & ~n10390;
  assign n10392 = ~n10285 & ~n10391;
  assign n10393 = controllable_BtoS_ACK9 & ~n10392;
  assign n10394 = ~n10314 & ~n10391;
  assign n10395 = ~controllable_BtoS_ACK9 & ~n10394;
  assign n10396 = ~n10393 & ~n10395;
  assign n10397 = ~controllable_DEQ & ~n10396;
  assign n10398 = ~n10344 & ~n10397;
  assign n10399 = ~i_nEMPTY & ~n10398;
  assign n10400 = ~n10379 & ~n10399;
  assign n10401 = ~i_FULL & ~n10400;
  assign n10402 = ~n10389 & ~n10401;
  assign n10403 = ~i_RtoB_ACK0 & ~n10402;
  assign n10404 = ~n10369 & ~n10403;
  assign n10405 = n6660 & ~n10404;
  assign n10406 = ~n8018 & ~n10365;
  assign n10407 = i_nEMPTY & ~n10406;
  assign n10408 = ~n8023 & ~n10407;
  assign n10409 = i_RtoB_ACK0 & ~n10408;
  assign n10410 = ~n8461 & ~n10371;
  assign n10411 = i_nEMPTY & ~n10410;
  assign n10412 = ~n8467 & ~n10336;
  assign n10413 = ~i_nEMPTY & ~n10412;
  assign n10414 = ~n10411 & ~n10413;
  assign n10415 = i_FULL & ~n10414;
  assign n10416 = ~n8491 & ~n10344;
  assign n10417 = ~i_nEMPTY & ~n10416;
  assign n10418 = ~n10411 & ~n10417;
  assign n10419 = ~i_FULL & ~n10418;
  assign n10420 = ~n10415 & ~n10419;
  assign n10421 = ~i_RtoB_ACK0 & ~n10420;
  assign n10422 = ~n10409 & ~n10421;
  assign n10423 = ~n6660 & ~n10422;
  assign n10424 = ~n10405 & ~n10423;
  assign n10425 = ~n6659 & ~n10424;
  assign n10426 = ~n8149 & ~n10424;
  assign n10427 = ~n8149 & ~n10426;
  assign n10428 = n6659 & ~n10427;
  assign n10429 = ~n10425 & ~n10428;
  assign n10430 = ~n6651 & ~n10429;
  assign n10431 = ~n10361 & ~n10430;
  assign n10432 = ~controllable_BtoR_REQ0 & ~n10431;
  assign n10433 = ~controllable_BtoR_REQ0 & ~n10432;
  assign n10434 = i_RtoB_ACK1 & ~n10433;
  assign n10435 = ~n9036 & ~n9058;
  assign n10436 = controllable_BtoS_ACK9 & ~n10435;
  assign n10437 = i_StoB_REQ9 & ~n9176;
  assign n10438 = ~n9058 & ~n10437;
  assign n10439 = ~controllable_BtoS_ACK9 & ~n10438;
  assign n10440 = ~n10436 & ~n10439;
  assign n10441 = controllable_DEQ & ~n10440;
  assign n10442 = ~n9063 & ~n9068;
  assign n10443 = controllable_BtoS_ACK9 & ~n10442;
  assign n10444 = i_StoB_REQ9 & ~n8111;
  assign n10445 = ~n9068 & ~n10444;
  assign n10446 = ~controllable_BtoS_ACK9 & ~n10445;
  assign n10447 = ~n10443 & ~n10446;
  assign n10448 = ~controllable_DEQ & ~n10447;
  assign n10449 = ~n10441 & ~n10448;
  assign n10450 = i_nEMPTY & ~n10449;
  assign n10451 = ~controllable_DEQ & ~n10440;
  assign n10452 = ~controllable_DEQ & ~n10451;
  assign n10453 = ~i_nEMPTY & ~n10452;
  assign n10454 = ~n10450 & ~n10453;
  assign n10455 = i_RtoB_ACK0 & ~n10454;
  assign n10456 = ~n9082 & ~n9090;
  assign n10457 = controllable_BtoS_ACK9 & ~n10456;
  assign n10458 = i_StoB_REQ9 & ~n8123;
  assign n10459 = ~n9090 & ~n10458;
  assign n10460 = ~controllable_BtoS_ACK9 & ~n10459;
  assign n10461 = ~n10457 & ~n10460;
  assign n10462 = controllable_DEQ & ~n10461;
  assign n10463 = ~n9782 & ~n10462;
  assign n10464 = i_nEMPTY & ~n10463;
  assign n10465 = ~n9098 & ~n9106;
  assign n10466 = controllable_BtoS_ACK9 & ~n10465;
  assign n10467 = i_StoB_REQ9 & ~n9308;
  assign n10468 = ~n9106 & ~n10467;
  assign n10469 = ~controllable_BtoS_ACK9 & ~n10468;
  assign n10470 = ~n10466 & ~n10469;
  assign n10471 = controllable_DEQ & ~n10470;
  assign n10472 = ~n9797 & ~n10471;
  assign n10473 = ~i_nEMPTY & ~n10472;
  assign n10474 = ~n10464 & ~n10473;
  assign n10475 = i_FULL & ~n10474;
  assign n10476 = ~n9082 & ~n9116;
  assign n10477 = controllable_BtoS_ACK9 & ~n10476;
  assign n10478 = ~n9116 & ~n10444;
  assign n10479 = ~controllable_BtoS_ACK9 & ~n10478;
  assign n10480 = ~n10477 & ~n10479;
  assign n10481 = controllable_DEQ & ~n10480;
  assign n10482 = ~n9814 & ~n10481;
  assign n10483 = i_nEMPTY & ~n10482;
  assign n10484 = controllable_DEQ & ~n10447;
  assign n10485 = ~controllable_DEQ & ~n10461;
  assign n10486 = ~n10484 & ~n10485;
  assign n10487 = ~i_nEMPTY & ~n10486;
  assign n10488 = ~n10483 & ~n10487;
  assign n10489 = ~i_FULL & ~n10488;
  assign n10490 = ~n10475 & ~n10489;
  assign n10491 = ~i_RtoB_ACK0 & ~n10490;
  assign n10492 = ~n10455 & ~n10491;
  assign n10493 = n6660 & ~n10492;
  assign n10494 = ~n9132 & ~n10493;
  assign n10495 = ~n6659 & ~n10494;
  assign n10496 = ~n8149 & ~n10494;
  assign n10497 = ~n8149 & ~n10496;
  assign n10498 = n6659 & ~n10497;
  assign n10499 = ~n10495 & ~n10498;
  assign n10500 = ~controllable_BtoR_REQ0 & ~n10499;
  assign n10501 = ~controllable_BtoR_REQ0 & ~n10500;
  assign n10502 = ~i_RtoB_ACK1 & ~n10501;
  assign n10503 = ~n10434 & ~n10502;
  assign n10504 = controllable_BtoR_REQ1 & ~n10503;
  assign n10505 = ~i_RtoB_ACK0 & ~n10454;
  assign n10506 = ~n9768 & ~n10505;
  assign n10507 = n6660 & ~n10506;
  assign n10508 = ~n9149 & ~n10507;
  assign n10509 = ~n8149 & ~n10508;
  assign n10510 = ~n8149 & ~n10509;
  assign n10511 = ~n6659 & ~n10510;
  assign n10512 = n6659 & ~n10508;
  assign n10513 = ~n10511 & ~n10512;
  assign n10514 = n6652 & ~n10513;
  assign n10515 = ~n10369 & ~n10505;
  assign n10516 = n6660 & ~n10515;
  assign n10517 = ~n9147 & ~n10409;
  assign n10518 = ~n6660 & ~n10517;
  assign n10519 = ~n10516 & ~n10518;
  assign n10520 = ~n8149 & ~n10519;
  assign n10521 = ~n8149 & ~n10520;
  assign n10522 = ~n6659 & ~n10521;
  assign n10523 = n6659 & ~n10519;
  assign n10524 = ~n10522 & ~n10523;
  assign n10525 = ~n6652 & ~n10524;
  assign n10526 = ~n10514 & ~n10525;
  assign n10527 = controllable_BtoR_REQ0 & ~n10526;
  assign n10528 = ~n8033 & ~n9177;
  assign n10529 = controllable_BtoS_ACK9 & ~n10528;
  assign n10530 = ~controllable_BtoS_ACK9 & ~n9176;
  assign n10531 = ~n10529 & ~n10530;
  assign n10532 = controllable_DEQ & ~n10531;
  assign n10533 = ~n8061 & ~n9182;
  assign n10534 = controllable_BtoS_ACK9 & ~n10533;
  assign n10535 = ~controllable_BtoS_ACK9 & ~n8111;
  assign n10536 = ~n10534 & ~n10535;
  assign n10537 = ~controllable_DEQ & ~n10536;
  assign n10538 = ~n10532 & ~n10537;
  assign n10539 = i_nEMPTY & ~n10538;
  assign n10540 = ~controllable_DEQ & ~n10531;
  assign n10541 = ~controllable_DEQ & ~n10540;
  assign n10542 = ~i_nEMPTY & ~n10541;
  assign n10543 = ~n10539 & ~n10542;
  assign n10544 = n6660 & ~n10543;
  assign n10545 = ~n9193 & ~n10544;
  assign n10546 = n6652 & ~n10545;
  assign n10547 = ~n6659 & ~n10545;
  assign n10548 = i_RtoB_ACK0 & ~n10543;
  assign n10549 = controllable_ENQ & ~n9911;
  assign n10550 = ~i_StoB_REQ9 & ~n10549;
  assign n10551 = ~n8404 & ~n10550;
  assign n10552 = controllable_BtoS_ACK9 & ~n10551;
  assign n10553 = ~n8379 & ~n10550;
  assign n10554 = ~controllable_BtoS_ACK9 & ~n10553;
  assign n10555 = ~n10552 & ~n10554;
  assign n10556 = controllable_DEQ & ~n10555;
  assign n10557 = ~n10272 & ~n10556;
  assign n10558 = i_nEMPTY & ~n10557;
  assign n10559 = ~controllable_DEQ & ~n10297;
  assign n10560 = ~i_nEMPTY & ~n10559;
  assign n10561 = ~n10558 & ~n10560;
  assign n10562 = ~i_RtoB_ACK0 & ~n10561;
  assign n10563 = ~n10548 & ~n10562;
  assign n10564 = n6660 & ~n10563;
  assign n10565 = ~n9216 & ~n10564;
  assign n10566 = n6659 & ~n10565;
  assign n10567 = ~n10547 & ~n10566;
  assign n10568 = ~n6652 & ~n10567;
  assign n10569 = ~n10546 & ~n10568;
  assign n10570 = ~controllable_BtoR_REQ0 & ~n10569;
  assign n10571 = ~n10527 & ~n10570;
  assign n10572 = i_RtoB_ACK1 & ~n10571;
  assign n10573 = i_RtoB_ACK0 & ~n9823;
  assign n10574 = ~n10491 & ~n10573;
  assign n10575 = n6660 & ~n10574;
  assign n10576 = ~n9230 & ~n10575;
  assign n10577 = ~n8149 & ~n10576;
  assign n10578 = ~n8149 & ~n10577;
  assign n10579 = ~n6659 & ~n10578;
  assign n10580 = n6659 & ~n10576;
  assign n10581 = ~n10579 & ~n10580;
  assign n10582 = n6652 & ~n10581;
  assign n10583 = i_RtoB_ACK0 & ~n10402;
  assign n10584 = ~n10491 & ~n10583;
  assign n10585 = n6660 & ~n10584;
  assign n10586 = i_RtoB_ACK0 & ~n10420;
  assign n10587 = ~n9130 & ~n10586;
  assign n10588 = ~n6660 & ~n10587;
  assign n10589 = ~n10585 & ~n10588;
  assign n10590 = ~n8149 & ~n10589;
  assign n10591 = ~n8149 & ~n10590;
  assign n10592 = ~n6659 & ~n10591;
  assign n10593 = n6659 & ~n10589;
  assign n10594 = ~n10592 & ~n10593;
  assign n10595 = ~n6652 & ~n10594;
  assign n10596 = ~n10582 & ~n10595;
  assign n10597 = n6651 & ~n10596;
  assign n10598 = i_RtoB_ACK0 & ~n10323;
  assign n10599 = ~n10491 & ~n10598;
  assign n10600 = n6660 & ~n10599;
  assign n10601 = i_RtoB_ACK0 & ~n10349;
  assign n10602 = ~n9130 & ~n10601;
  assign n10603 = ~n6660 & ~n10602;
  assign n10604 = ~n10600 & ~n10603;
  assign n10605 = ~n8149 & ~n10604;
  assign n10606 = ~n8149 & ~n10605;
  assign n10607 = ~n6659 & ~n10606;
  assign n10608 = n6659 & ~n10604;
  assign n10609 = ~n10607 & ~n10608;
  assign n10610 = n6652 & ~n10609;
  assign n10611 = ~n10595 & ~n10610;
  assign n10612 = ~n6651 & ~n10611;
  assign n10613 = ~n10597 & ~n10612;
  assign n10614 = controllable_BtoR_REQ0 & ~n10613;
  assign n10615 = controllable_DEQ & ~n9813;
  assign n10616 = ~n9782 & ~n10615;
  assign n10617 = i_nEMPTY & ~n10616;
  assign n10618 = ~n9302 & ~n9309;
  assign n10619 = controllable_BtoS_ACK9 & ~n10618;
  assign n10620 = ~controllable_BtoS_ACK9 & ~n9308;
  assign n10621 = ~n10619 & ~n10620;
  assign n10622 = controllable_DEQ & ~n10621;
  assign n10623 = ~n9797 & ~n10622;
  assign n10624 = ~i_nEMPTY & ~n10623;
  assign n10625 = ~n10617 & ~n10624;
  assign n10626 = i_FULL & ~n10625;
  assign n10627 = controllable_DEQ & ~n10536;
  assign n10628 = ~n9814 & ~n10627;
  assign n10629 = i_nEMPTY & ~n10628;
  assign n10630 = ~n10485 & ~n10627;
  assign n10631 = ~i_nEMPTY & ~n10630;
  assign n10632 = ~n10629 & ~n10631;
  assign n10633 = ~i_FULL & ~n10632;
  assign n10634 = ~n10626 & ~n10633;
  assign n10635 = ~i_RtoB_ACK0 & ~n10634;
  assign n10636 = ~n10548 & ~n10635;
  assign n10637 = n6660 & ~n10636;
  assign n10638 = ~n9328 & ~n10637;
  assign n10639 = n6652 & ~n10638;
  assign n10640 = ~n6659 & ~n10638;
  assign n10641 = ~controllable_ENQ & ~n9910;
  assign n10642 = ~n8039 & ~n10641;
  assign n10643 = ~i_StoB_REQ9 & ~n10642;
  assign n10644 = ~n9591 & ~n10643;
  assign n10645 = controllable_BtoS_ACK9 & ~n10644;
  assign n10646 = ~n8368 & ~n10643;
  assign n10647 = ~controllable_BtoS_ACK9 & ~n10646;
  assign n10648 = ~n10645 & ~n10647;
  assign n10649 = controllable_DEQ & ~n10648;
  assign n10650 = ~i_StoB_REQ9 & ~n9601;
  assign n10651 = ~n8061 & ~n10650;
  assign n10652 = controllable_BtoS_ACK9 & ~n10651;
  assign n10653 = ~n9607 & ~n10652;
  assign n10654 = ~controllable_DEQ & ~n10653;
  assign n10655 = ~n10649 & ~n10654;
  assign n10656 = i_nEMPTY & ~n10655;
  assign n10657 = ~controllable_ENQ & ~n10641;
  assign n10658 = ~i_StoB_REQ9 & ~n10657;
  assign n10659 = ~n9613 & ~n10658;
  assign n10660 = controllable_BtoS_ACK9 & ~n10659;
  assign n10661 = ~n9538 & ~n10658;
  assign n10662 = ~controllable_BtoS_ACK9 & ~n10661;
  assign n10663 = ~n10660 & ~n10662;
  assign n10664 = controllable_DEQ & ~n10663;
  assign n10665 = ~i_StoB_REQ9 & ~n9619;
  assign n10666 = ~n8033 & ~n10665;
  assign n10667 = controllable_BtoS_ACK9 & ~n10666;
  assign n10668 = ~n9620 & ~n10667;
  assign n10669 = ~controllable_DEQ & ~n10668;
  assign n10670 = ~n10664 & ~n10669;
  assign n10671 = ~i_nEMPTY & ~n10670;
  assign n10672 = ~n10656 & ~n10671;
  assign n10673 = i_FULL & ~n10672;
  assign n10674 = ~controllable_ENQ & ~n10087;
  assign n10675 = ~n8031 & ~n10674;
  assign n10676 = i_StoB_REQ9 & ~n10675;
  assign n10677 = ~controllable_ENQ & ~n10267;
  assign n10678 = ~n9602 & ~n10677;
  assign n10679 = ~i_StoB_REQ9 & ~n10678;
  assign n10680 = ~n10676 & ~n10679;
  assign n10681 = controllable_BtoS_ACK9 & ~n10680;
  assign n10682 = ~controllable_BtoS_ACK9 & ~n10678;
  assign n10683 = ~n10681 & ~n10682;
  assign n10684 = ~controllable_DEQ & ~n10683;
  assign n10685 = ~n10649 & ~n10684;
  assign n10686 = i_nEMPTY & ~n10685;
  assign n10687 = ~i_StoB_REQ9 & ~n9910;
  assign n10688 = ~n8415 & ~n10687;
  assign n10689 = controllable_BtoS_ACK9 & ~n10688;
  assign n10690 = ~n8368 & ~n10687;
  assign n10691 = ~controllable_BtoS_ACK9 & ~n10690;
  assign n10692 = ~n10689 & ~n10691;
  assign n10693 = controllable_DEQ & ~n10692;
  assign n10694 = ~n6671 & ~n6941;
  assign n10695 = n6670 & ~n10694;
  assign n10696 = ~n9928 & ~n10695;
  assign n10697 = n6669 & ~n10696;
  assign n10698 = ~n6946 & ~n10697;
  assign n10699 = ~i_StoB_REQ2 & ~n10698;
  assign n10700 = ~i_StoB_REQ2 & ~n10699;
  assign n10701 = controllable_BtoS_ACK2 & ~n10700;
  assign n10702 = ~n10097 & ~n10699;
  assign n10703 = ~controllable_BtoS_ACK2 & ~n10702;
  assign n10704 = ~n10701 & ~n10703;
  assign n10705 = n6668 & ~n10704;
  assign n10706 = ~n6968 & ~n10705;
  assign n10707 = ~i_StoB_REQ3 & ~n10706;
  assign n10708 = ~i_StoB_REQ3 & ~n10707;
  assign n10709 = controllable_BtoS_ACK3 & ~n10708;
  assign n10710 = ~n10096 & ~n10707;
  assign n10711 = ~controllable_BtoS_ACK3 & ~n10710;
  assign n10712 = ~n10709 & ~n10711;
  assign n10713 = n6667 & ~n10712;
  assign n10714 = ~n9949 & ~n10713;
  assign n10715 = ~i_StoB_REQ4 & ~n10714;
  assign n10716 = ~n10037 & ~n10715;
  assign n10717 = n6666 & ~n10716;
  assign n10718 = ~n7015 & ~n10717;
  assign n10719 = ~i_StoB_REQ5 & ~n10718;
  assign n10720 = ~i_StoB_REQ5 & ~n10719;
  assign n10721 = controllable_BtoS_ACK5 & ~n10720;
  assign n10722 = ~n10094 & ~n10719;
  assign n10723 = ~controllable_BtoS_ACK5 & ~n10722;
  assign n10724 = ~n10721 & ~n10723;
  assign n10725 = n6665 & ~n10724;
  assign n10726 = ~n7038 & ~n10725;
  assign n10727 = ~i_StoB_REQ6 & ~n10726;
  assign n10728 = ~i_StoB_REQ6 & ~n10727;
  assign n10729 = controllable_BtoS_ACK6 & ~n10728;
  assign n10730 = ~n10093 & ~n10727;
  assign n10731 = ~controllable_BtoS_ACK6 & ~n10730;
  assign n10732 = ~n10729 & ~n10731;
  assign n10733 = ~i_StoB_REQ7 & ~n10732;
  assign n10734 = ~i_StoB_REQ7 & ~n10733;
  assign n10735 = n6664 & ~n10734;
  assign n10736 = ~n7070 & ~n10735;
  assign n10737 = controllable_BtoS_ACK7 & ~n10736;
  assign n10738 = ~n10092 & ~n10733;
  assign n10739 = n6664 & ~n10738;
  assign n10740 = ~n9978 & ~n10739;
  assign n10741 = ~controllable_BtoS_ACK7 & ~n10740;
  assign n10742 = ~n10737 & ~n10741;
  assign n10743 = n6663 & ~n10742;
  assign n10744 = ~n7096 & ~n10743;
  assign n10745 = ~i_StoB_REQ8 & ~n10744;
  assign n10746 = ~i_StoB_REQ8 & ~n10745;
  assign n10747 = controllable_BtoS_ACK8 & ~n10746;
  assign n10748 = ~n10091 & ~n10745;
  assign n10749 = ~controllable_BtoS_ACK8 & ~n10748;
  assign n10750 = ~n10747 & ~n10749;
  assign n10751 = n6662 & ~n10750;
  assign n10752 = ~n7125 & ~n10751;
  assign n10753 = ~i_StoB_REQ10 & ~n10752;
  assign n10754 = ~i_StoB_REQ10 & ~n10753;
  assign n10755 = controllable_BtoS_ACK10 & ~n10754;
  assign n10756 = ~n10090 & ~n10753;
  assign n10757 = ~controllable_BtoS_ACK10 & ~n10756;
  assign n10758 = ~n10755 & ~n10757;
  assign n10759 = n6661 & ~n10758;
  assign n10760 = ~n10001 & ~n10759;
  assign n10761 = ~i_StoB_REQ11 & ~n10760;
  assign n10762 = ~n10083 & ~n10761;
  assign n10763 = ~controllable_ENQ & ~n10762;
  assign n10764 = ~n8031 & ~n10763;
  assign n10765 = i_StoB_REQ9 & ~n10764;
  assign n10766 = controllable_BtoS_ACK11 & ~n10758;
  assign n10767 = ~n10163 & ~n10766;
  assign n10768 = n6661 & ~n10767;
  assign n10769 = ~n6661 & ~n9037;
  assign n10770 = ~n10768 & ~n10769;
  assign n10771 = i_StoB_REQ11 & ~n10770;
  assign n10772 = i_StoB_REQ10 & ~n10752;
  assign n10773 = i_StoB_REQ8 & ~n10744;
  assign n10774 = i_StoB_REQ7 & ~n10732;
  assign n10775 = i_StoB_REQ6 & ~n10726;
  assign n10776 = i_StoB_REQ5 & ~n10718;
  assign n10777 = controllable_BtoS_ACK4 & ~n10712;
  assign n10778 = ~n10116 & ~n10777;
  assign n10779 = n6667 & ~n10778;
  assign n10780 = ~n6667 & ~n8783;
  assign n10781 = ~n10779 & ~n10780;
  assign n10782 = i_StoB_REQ4 & ~n10781;
  assign n10783 = i_StoB_REQ3 & ~n10706;
  assign n10784 = i_StoB_REQ2 & ~n10698;
  assign n10785 = ~n6671 & ~n8714;
  assign n10786 = ~n6671 & ~n10785;
  assign n10787 = n6670 & ~n10786;
  assign n10788 = ~n6670 & ~n8714;
  assign n10789 = ~n10787 & ~n10788;
  assign n10790 = n6669 & ~n10789;
  assign n10791 = ~n8720 & ~n10790;
  assign n10792 = ~i_StoB_REQ2 & ~n10791;
  assign n10793 = ~n10784 & ~n10792;
  assign n10794 = controllable_BtoS_ACK2 & ~n10793;
  assign n10795 = ~n10190 & ~n10792;
  assign n10796 = ~controllable_BtoS_ACK2 & ~n10795;
  assign n10797 = ~n10794 & ~n10796;
  assign n10798 = n6668 & ~n10797;
  assign n10799 = ~n8738 & ~n10798;
  assign n10800 = ~i_StoB_REQ3 & ~n10799;
  assign n10801 = ~n10783 & ~n10800;
  assign n10802 = controllable_BtoS_ACK3 & ~n10801;
  assign n10803 = ~n10199 & ~n10800;
  assign n10804 = ~controllable_BtoS_ACK3 & ~n10803;
  assign n10805 = ~n10802 & ~n10804;
  assign n10806 = n6667 & ~n10805;
  assign n10807 = ~n6667 & ~n8764;
  assign n10808 = ~n10806 & ~n10807;
  assign n10809 = ~i_StoB_REQ4 & ~n10808;
  assign n10810 = ~n10782 & ~n10809;
  assign n10811 = n6666 & ~n10810;
  assign n10812 = ~n8787 & ~n10811;
  assign n10813 = ~i_StoB_REQ5 & ~n10812;
  assign n10814 = ~n10776 & ~n10813;
  assign n10815 = controllable_BtoS_ACK5 & ~n10814;
  assign n10816 = ~n10212 & ~n10813;
  assign n10817 = ~controllable_BtoS_ACK5 & ~n10816;
  assign n10818 = ~n10815 & ~n10817;
  assign n10819 = n6665 & ~n10818;
  assign n10820 = ~n8814 & ~n10819;
  assign n10821 = ~i_StoB_REQ6 & ~n10820;
  assign n10822 = ~n10775 & ~n10821;
  assign n10823 = controllable_BtoS_ACK6 & ~n10822;
  assign n10824 = ~n10221 & ~n10821;
  assign n10825 = ~controllable_BtoS_ACK6 & ~n10824;
  assign n10826 = ~n10823 & ~n10825;
  assign n10827 = ~i_StoB_REQ7 & ~n10826;
  assign n10828 = ~n10774 & ~n10827;
  assign n10829 = n6664 & ~n10828;
  assign n10830 = ~n6664 & ~n8872;
  assign n10831 = ~n10829 & ~n10830;
  assign n10832 = controllable_BtoS_ACK7 & ~n10831;
  assign n10833 = ~n10230 & ~n10827;
  assign n10834 = n6664 & ~n10833;
  assign n10835 = ~n6664 & ~n8874;
  assign n10836 = ~n10834 & ~n10835;
  assign n10837 = ~controllable_BtoS_ACK7 & ~n10836;
  assign n10838 = ~n10832 & ~n10837;
  assign n10839 = n6663 & ~n10838;
  assign n10840 = ~n8877 & ~n10839;
  assign n10841 = ~i_StoB_REQ8 & ~n10840;
  assign n10842 = ~n10773 & ~n10841;
  assign n10843 = controllable_BtoS_ACK8 & ~n10842;
  assign n10844 = ~n10241 & ~n10841;
  assign n10845 = ~controllable_BtoS_ACK8 & ~n10844;
  assign n10846 = ~n10843 & ~n10845;
  assign n10847 = n6662 & ~n10846;
  assign n10848 = ~n8906 & ~n10847;
  assign n10849 = ~i_StoB_REQ10 & ~n10848;
  assign n10850 = ~n10772 & ~n10849;
  assign n10851 = controllable_BtoS_ACK10 & ~n10850;
  assign n10852 = ~n10250 & ~n10849;
  assign n10853 = ~controllable_BtoS_ACK10 & ~n10852;
  assign n10854 = ~n10851 & ~n10853;
  assign n10855 = n6661 & ~n10854;
  assign n10856 = ~n6661 & ~n8934;
  assign n10857 = ~n10855 & ~n10856;
  assign n10858 = ~i_StoB_REQ11 & ~n10857;
  assign n10859 = ~n10771 & ~n10858;
  assign n10860 = ~controllable_ENQ & ~n10859;
  assign n10861 = ~n9602 & ~n10860;
  assign n10862 = ~i_StoB_REQ9 & ~n10861;
  assign n10863 = ~n10765 & ~n10862;
  assign n10864 = controllable_BtoS_ACK9 & ~n10863;
  assign n10865 = i_StoB_REQ9 & ~n10678;
  assign n10866 = ~n10862 & ~n10865;
  assign n10867 = ~controllable_BtoS_ACK9 & ~n10866;
  assign n10868 = ~n10864 & ~n10867;
  assign n10869 = ~controllable_DEQ & ~n10868;
  assign n10870 = ~n10693 & ~n10869;
  assign n10871 = ~i_nEMPTY & ~n10870;
  assign n10872 = ~n10686 & ~n10871;
  assign n10873 = ~i_FULL & ~n10872;
  assign n10874 = ~n10673 & ~n10873;
  assign n10875 = ~i_RtoB_ACK0 & ~n10874;
  assign n10876 = ~n10548 & ~n10875;
  assign n10877 = n6660 & ~n10876;
  assign n10878 = ~n9609 & ~n9628;
  assign n10879 = i_nEMPTY & ~n10878;
  assign n10880 = ~n9624 & ~n10879;
  assign n10881 = i_FULL & ~n10880;
  assign n10882 = ~n9648 & ~n10881;
  assign n10883 = ~i_RtoB_ACK0 & ~n10882;
  assign n10884 = ~n9207 & ~n10883;
  assign n10885 = ~n6660 & ~n10884;
  assign n10886 = ~n10877 & ~n10885;
  assign n10887 = n6659 & ~n10886;
  assign n10888 = ~n10640 & ~n10887;
  assign n10889 = ~n6652 & ~n10888;
  assign n10890 = ~n10639 & ~n10889;
  assign n10891 = n6651 & ~n10890;
  assign n10892 = i_RtoB_ACK0 & ~n10561;
  assign n10893 = ~n10875 & ~n10892;
  assign n10894 = n6660 & ~n10893;
  assign n10895 = ~n9662 & ~n10883;
  assign n10896 = ~n6660 & ~n10895;
  assign n10897 = ~n10894 & ~n10896;
  assign n10898 = ~n6659 & ~n10897;
  assign n10899 = n6659 & ~n10638;
  assign n10900 = ~n10898 & ~n10899;
  assign n10901 = n6652 & ~n10900;
  assign n10902 = ~n10887 & ~n10898;
  assign n10903 = ~n6652 & ~n10902;
  assign n10904 = ~n10901 & ~n10903;
  assign n10905 = ~n6651 & ~n10904;
  assign n10906 = ~n10891 & ~n10905;
  assign n10907 = ~controllable_BtoR_REQ0 & ~n10906;
  assign n10908 = ~n10614 & ~n10907;
  assign n10909 = ~i_RtoB_ACK1 & ~n10908;
  assign n10910 = ~n10572 & ~n10909;
  assign n10911 = ~controllable_BtoR_REQ1 & ~n10910;
  assign n10912 = ~n10504 & ~n10911;
  assign n10913 = n6649 & ~n10912;
  assign n10914 = ~controllable_DEQ & ~n10343;
  assign n10915 = ~n10365 & ~n10914;
  assign n10916 = i_nEMPTY & ~n10915;
  assign n10917 = ~controllable_DEQ & ~n10364;
  assign n10918 = ~controllable_DEQ & ~n10917;
  assign n10919 = ~i_nEMPTY & ~n10918;
  assign n10920 = ~n10916 & ~n10919;
  assign n10921 = i_RtoB_ACK0 & ~n10920;
  assign n10922 = ~controllable_DEQ & ~n10370;
  assign n10923 = ~n10344 & ~n10922;
  assign n10924 = ~i_nEMPTY & ~n10923;
  assign n10925 = ~n10411 & ~n10924;
  assign n10926 = ~i_FULL & ~n10925;
  assign n10927 = ~n10415 & ~n10926;
  assign n10928 = ~i_RtoB_ACK0 & ~n10927;
  assign n10929 = ~n10921 & ~n10928;
  assign n10930 = ~n6659 & ~n10929;
  assign n10931 = ~n8149 & ~n10929;
  assign n10932 = ~n8149 & ~n10931;
  assign n10933 = n6659 & ~n10932;
  assign n10934 = ~n10930 & ~n10933;
  assign n10935 = ~controllable_BtoR_REQ0 & ~n10934;
  assign n10936 = ~controllable_BtoR_REQ0 & ~n10935;
  assign n10937 = i_RtoB_ACK1 & ~n10936;
  assign n10938 = i_StoB_REQ9 & ~n7986;
  assign n10939 = ~n9043 & ~n10938;
  assign n10940 = controllable_BtoS_ACK9 & ~n10939;
  assign n10941 = ~n8379 & ~n9043;
  assign n10942 = ~controllable_BtoS_ACK9 & ~n10941;
  assign n10943 = ~n10940 & ~n10942;
  assign n10944 = controllable_DEQ & ~n10943;
  assign n10945 = i_StoB_REQ9 & ~n7984;
  assign n10946 = ~n9064 & ~n10945;
  assign n10947 = controllable_BtoS_ACK9 & ~n10946;
  assign n10948 = ~n8368 & ~n9064;
  assign n10949 = ~controllable_BtoS_ACK9 & ~n10948;
  assign n10950 = ~n10947 & ~n10949;
  assign n10951 = ~controllable_DEQ & ~n10950;
  assign n10952 = ~n10944 & ~n10951;
  assign n10953 = i_nEMPTY & ~n10952;
  assign n10954 = ~controllable_DEQ & ~n10943;
  assign n10955 = ~controllable_DEQ & ~n10954;
  assign n10956 = ~i_nEMPTY & ~n10955;
  assign n10957 = ~n10953 & ~n10956;
  assign n10958 = i_RtoB_ACK0 & ~n10957;
  assign n10959 = ~n8368 & ~n9085;
  assign n10960 = ~controllable_BtoS_ACK9 & ~n10959;
  assign n10961 = ~n9637 & ~n10960;
  assign n10962 = controllable_DEQ & ~n10961;
  assign n10963 = ~n8461 & ~n10962;
  assign n10964 = i_nEMPTY & ~n10963;
  assign n10965 = i_StoB_REQ9 & ~n8070;
  assign n10966 = ~n9100 & ~n10965;
  assign n10967 = controllable_BtoS_ACK9 & ~n10966;
  assign n10968 = ~n9100 & ~n9538;
  assign n10969 = ~controllable_BtoS_ACK9 & ~n10968;
  assign n10970 = ~n10967 & ~n10969;
  assign n10971 = controllable_DEQ & ~n10970;
  assign n10972 = ~n8467 & ~n10971;
  assign n10973 = ~i_nEMPTY & ~n10972;
  assign n10974 = ~n10964 & ~n10973;
  assign n10975 = i_FULL & ~n10974;
  assign n10976 = controllable_DEQ & ~n10950;
  assign n10977 = ~controllable_DEQ & ~n10961;
  assign n10978 = ~n10976 & ~n10977;
  assign n10979 = ~i_nEMPTY & ~n10978;
  assign n10980 = ~n10964 & ~n10979;
  assign n10981 = ~i_FULL & ~n10980;
  assign n10982 = ~n10975 & ~n10981;
  assign n10983 = ~i_RtoB_ACK0 & ~n10982;
  assign n10984 = ~n10958 & ~n10983;
  assign n10985 = ~n6659 & ~n10984;
  assign n10986 = ~n8149 & ~n10984;
  assign n10987 = ~n8149 & ~n10986;
  assign n10988 = n6659 & ~n10987;
  assign n10989 = ~n10985 & ~n10988;
  assign n10990 = ~controllable_BtoR_REQ0 & ~n10989;
  assign n10991 = ~controllable_BtoR_REQ0 & ~n10990;
  assign n10992 = ~i_RtoB_ACK1 & ~n10991;
  assign n10993 = ~n10937 & ~n10992;
  assign n10994 = controllable_BtoR_REQ1 & ~n10993;
  assign n10995 = ~i_RtoB_ACK0 & ~n10957;
  assign n10996 = ~n10921 & ~n10995;
  assign n10997 = ~n8149 & ~n10996;
  assign n10998 = ~n8149 & ~n10997;
  assign n10999 = ~n6659 & ~n10998;
  assign n11000 = n6659 & ~n10996;
  assign n11001 = ~n10999 & ~n11000;
  assign n11002 = controllable_BtoR_REQ0 & ~n11001;
  assign n11003 = controllable_DEQ & ~n8466;
  assign n11004 = ~n8461 & ~n11003;
  assign n11005 = i_nEMPTY & ~n11004;
  assign n11006 = ~controllable_DEQ & ~n8467;
  assign n11007 = ~i_nEMPTY & ~n11006;
  assign n11008 = ~n11005 & ~n11007;
  assign n11009 = ~controllable_BtoR_REQ0 & ~n11008;
  assign n11010 = ~n11002 & ~n11009;
  assign n11011 = i_RtoB_ACK1 & ~n11010;
  assign n11012 = i_RtoB_ACK0 & ~n10927;
  assign n11013 = ~n10983 & ~n11012;
  assign n11014 = ~n8149 & ~n11013;
  assign n11015 = ~n8149 & ~n11014;
  assign n11016 = ~n6659 & ~n11015;
  assign n11017 = n6659 & ~n11013;
  assign n11018 = ~n11016 & ~n11017;
  assign n11019 = controllable_BtoR_REQ0 & ~n11018;
  assign n11020 = i_RtoB_ACK0 & ~n11008;
  assign n11021 = i_nEMPTY & ~n8460;
  assign n11022 = ~n8075 & ~n9305;
  assign n11023 = controllable_BtoS_ACK9 & ~n11022;
  assign n11024 = ~n9616 & ~n11023;
  assign n11025 = controllable_DEQ & ~n11024;
  assign n11026 = ~n8467 & ~n11025;
  assign n11027 = ~i_nEMPTY & ~n11026;
  assign n11028 = ~n11021 & ~n11027;
  assign n11029 = i_FULL & ~n11028;
  assign n11030 = ~i_FULL & ~n8460;
  assign n11031 = ~n11029 & ~n11030;
  assign n11032 = ~i_RtoB_ACK0 & ~n11031;
  assign n11033 = ~n11020 & ~n11032;
  assign n11034 = ~controllable_BtoR_REQ0 & ~n11033;
  assign n11035 = ~n11019 & ~n11034;
  assign n11036 = ~i_RtoB_ACK1 & ~n11035;
  assign n11037 = ~n11011 & ~n11036;
  assign n11038 = ~controllable_BtoR_REQ1 & ~n11037;
  assign n11039 = ~n10994 & ~n11038;
  assign n11040 = ~n6649 & ~n11039;
  assign n11041 = ~n10913 & ~n11040;
  assign n11042 = ~n6647 & ~n11041;
  assign n11043 = ~n9741 & ~n11042;
  assign n11044 = n6646 & ~n11043;
  assign n11045 = controllable_DEQ & ~n8460;
  assign n11046 = ~n10977 & ~n11045;
  assign n11047 = ~i_nEMPTY & ~n11046;
  assign n11048 = ~n11021 & ~n11047;
  assign n11049 = ~i_FULL & ~n11048;
  assign n11050 = ~n11029 & ~n11049;
  assign n11051 = ~i_RtoB_ACK0 & ~n11050;
  assign n11052 = ~n11020 & ~n11051;
  assign n11053 = ~controllable_BtoR_REQ0 & ~n11052;
  assign n11054 = ~n11019 & ~n11053;
  assign n11055 = ~i_RtoB_ACK1 & ~n11054;
  assign n11056 = ~n11011 & ~n11055;
  assign n11057 = ~controllable_BtoR_REQ1 & ~n11056;
  assign n11058 = ~n10994 & ~n11057;
  assign n11059 = n6649 & ~n11058;
  assign n11060 = ~n11040 & ~n11059;
  assign n11061 = n6647 & ~n11060;
  assign n11062 = n6661 & ~n8226;
  assign n11063 = ~n10261 & ~n11062;
  assign n11064 = i_StoB_REQ11 & ~n11063;
  assign n11065 = n6667 & ~n8248;
  assign n11066 = ~n10119 & ~n11065;
  assign n11067 = i_StoB_REQ4 & ~n11066;
  assign n11068 = ~n8271 & ~n8715;
  assign n11069 = n6670 & ~n11068;
  assign n11070 = ~n10100 & ~n11069;
  assign n11071 = n6669 & ~n11070;
  assign n11072 = ~n7407 & ~n11071;
  assign n11073 = ~i_StoB_REQ2 & ~n11072;
  assign n11074 = ~n9935 & ~n11073;
  assign n11075 = controllable_BtoS_ACK2 & ~n11074;
  assign n11076 = ~n8280 & ~n11073;
  assign n11077 = ~controllable_BtoS_ACK2 & ~n11076;
  assign n11078 = ~n11075 & ~n11077;
  assign n11079 = n6668 & ~n11078;
  assign n11080 = ~n7425 & ~n11079;
  assign n11081 = ~i_StoB_REQ3 & ~n11080;
  assign n11082 = ~n9944 & ~n11081;
  assign n11083 = controllable_BtoS_ACK3 & ~n11082;
  assign n11084 = ~n8289 & ~n11081;
  assign n11085 = ~controllable_BtoS_ACK3 & ~n11084;
  assign n11086 = ~n11083 & ~n11085;
  assign n11087 = n6667 & ~n11086;
  assign n11088 = ~n8294 & ~n11087;
  assign n11089 = ~i_StoB_REQ4 & ~n11088;
  assign n11090 = ~n11067 & ~n11089;
  assign n11091 = n6666 & ~n11090;
  assign n11092 = ~n7477 & ~n11091;
  assign n11093 = ~i_StoB_REQ5 & ~n11092;
  assign n11094 = ~n9958 & ~n11093;
  assign n11095 = controllable_BtoS_ACK5 & ~n11094;
  assign n11096 = ~n8303 & ~n11093;
  assign n11097 = ~controllable_BtoS_ACK5 & ~n11096;
  assign n11098 = ~n11095 & ~n11097;
  assign n11099 = n6665 & ~n11098;
  assign n11100 = ~n7497 & ~n11099;
  assign n11101 = ~i_StoB_REQ6 & ~n11100;
  assign n11102 = ~n9967 & ~n11101;
  assign n11103 = controllable_BtoS_ACK6 & ~n11102;
  assign n11104 = ~n8312 & ~n11101;
  assign n11105 = ~controllable_BtoS_ACK6 & ~n11104;
  assign n11106 = ~n11103 & ~n11105;
  assign n11107 = ~i_StoB_REQ7 & ~n11106;
  assign n11108 = ~n8319 & ~n11107;
  assign n11109 = n6664 & ~n11108;
  assign n11110 = ~n9443 & ~n11109;
  assign n11111 = controllable_BtoS_ACK7 & ~n11110;
  assign n11112 = ~n8324 & ~n11107;
  assign n11113 = n6664 & ~n11112;
  assign n11114 = ~n8327 & ~n11113;
  assign n11115 = ~controllable_BtoS_ACK7 & ~n11114;
  assign n11116 = ~n11111 & ~n11115;
  assign n11117 = n6663 & ~n11116;
  assign n11118 = ~n7546 & ~n11117;
  assign n11119 = ~i_StoB_REQ8 & ~n11118;
  assign n11120 = ~n9987 & ~n11119;
  assign n11121 = controllable_BtoS_ACK8 & ~n11120;
  assign n11122 = ~n8336 & ~n11119;
  assign n11123 = ~controllable_BtoS_ACK8 & ~n11122;
  assign n11124 = ~n11121 & ~n11123;
  assign n11125 = n6662 & ~n11124;
  assign n11126 = ~n7568 & ~n11125;
  assign n11127 = ~i_StoB_REQ10 & ~n11126;
  assign n11128 = ~n9996 & ~n11127;
  assign n11129 = controllable_BtoS_ACK10 & ~n11128;
  assign n11130 = ~n8345 & ~n11127;
  assign n11131 = ~controllable_BtoS_ACK10 & ~n11130;
  assign n11132 = ~n11129 & ~n11131;
  assign n11133 = n6661 & ~n11132;
  assign n11134 = ~n8350 & ~n11133;
  assign n11135 = ~i_StoB_REQ11 & ~n11134;
  assign n11136 = ~n11064 & ~n11135;
  assign n11137 = ~i_StoB_REQ9 & ~n11136;
  assign n11138 = ~n8415 & ~n11137;
  assign n11139 = controllable_BtoS_ACK9 & ~n11138;
  assign n11140 = ~n8368 & ~n11137;
  assign n11141 = ~controllable_BtoS_ACK9 & ~n11140;
  assign n11142 = ~n11139 & ~n11141;
  assign n11143 = ~controllable_DEQ & ~n11142;
  assign n11144 = ~n10371 & ~n11143;
  assign n11145 = i_nEMPTY & ~n11144;
  assign n11146 = controllable_ENQ & ~n11136;
  assign n11147 = controllable_ENQ & ~n11146;
  assign n11148 = ~i_StoB_REQ9 & ~n11147;
  assign n11149 = ~n8404 & ~n11148;
  assign n11150 = controllable_BtoS_ACK9 & ~n11149;
  assign n11151 = ~n8379 & ~n11148;
  assign n11152 = ~controllable_BtoS_ACK9 & ~n11151;
  assign n11153 = ~n11150 & ~n11152;
  assign n11154 = ~controllable_DEQ & ~n11153;
  assign n11155 = ~n10336 & ~n11154;
  assign n11156 = ~i_nEMPTY & ~n11155;
  assign n11157 = ~n11145 & ~n11156;
  assign n11158 = i_FULL & ~n11157;
  assign n11159 = ~n10005 & ~n11146;
  assign n11160 = ~i_StoB_REQ9 & ~n11159;
  assign n11161 = ~n8404 & ~n11160;
  assign n11162 = controllable_BtoS_ACK9 & ~n11161;
  assign n11163 = ~n10011 & ~n11160;
  assign n11164 = ~controllable_BtoS_ACK9 & ~n11163;
  assign n11165 = ~n11162 & ~n11164;
  assign n11166 = ~controllable_DEQ & ~n11165;
  assign n11167 = ~n10344 & ~n11166;
  assign n11168 = ~i_nEMPTY & ~n11167;
  assign n11169 = ~n11145 & ~n11168;
  assign n11170 = ~i_FULL & ~n11169;
  assign n11171 = ~n11158 & ~n11170;
  assign n11172 = ~i_RtoB_ACK0 & ~n11171;
  assign n11173 = ~n10921 & ~n11172;
  assign n11174 = n6660 & ~n11173;
  assign n11175 = ~n6660 & ~n10929;
  assign n11176 = ~n11174 & ~n11175;
  assign n11177 = ~n6659 & ~n11176;
  assign n11178 = ~n8149 & ~n11176;
  assign n11179 = ~n8149 & ~n11178;
  assign n11180 = n6659 & ~n11179;
  assign n11181 = ~n11177 & ~n11180;
  assign n11182 = n6651 & ~n11181;
  assign n11183 = ~n6651 & ~n10934;
  assign n11184 = ~n11182 & ~n11183;
  assign n11185 = ~controllable_BtoR_REQ0 & ~n11184;
  assign n11186 = ~controllable_BtoR_REQ0 & ~n11185;
  assign n11187 = i_RtoB_ACK1 & ~n11186;
  assign n11188 = ~n10377 & ~n10962;
  assign n11189 = i_nEMPTY & ~n11188;
  assign n11190 = ~n10385 & ~n10971;
  assign n11191 = ~i_nEMPTY & ~n11190;
  assign n11192 = ~n11189 & ~n11191;
  assign n11193 = i_FULL & ~n11192;
  assign n11194 = ~n10283 & ~n10763;
  assign n11195 = i_StoB_REQ9 & ~n11194;
  assign n11196 = ~n10291 & ~n10860;
  assign n11197 = ~i_StoB_REQ9 & ~n11196;
  assign n11198 = ~n11195 & ~n11197;
  assign n11199 = controllable_BtoS_ACK9 & ~n11198;
  assign n11200 = ~n10268 & ~n11197;
  assign n11201 = ~controllable_BtoS_ACK9 & ~n11200;
  assign n11202 = ~n11199 & ~n11201;
  assign n11203 = ~controllable_DEQ & ~n11202;
  assign n11204 = ~n10976 & ~n11203;
  assign n11205 = ~i_nEMPTY & ~n11204;
  assign n11206 = ~n11189 & ~n11205;
  assign n11207 = ~i_FULL & ~n11206;
  assign n11208 = ~n11193 & ~n11207;
  assign n11209 = ~i_RtoB_ACK0 & ~n11208;
  assign n11210 = ~n10958 & ~n11209;
  assign n11211 = n6660 & ~n11210;
  assign n11212 = ~n6660 & ~n10984;
  assign n11213 = ~n11211 & ~n11212;
  assign n11214 = ~n6659 & ~n11213;
  assign n11215 = ~n8149 & ~n11213;
  assign n11216 = ~n8149 & ~n11215;
  assign n11217 = n6659 & ~n11216;
  assign n11218 = ~n11214 & ~n11217;
  assign n11219 = n6651 & ~n11218;
  assign n11220 = ~n10962 & ~n11143;
  assign n11221 = i_nEMPTY & ~n11220;
  assign n11222 = ~n10971 & ~n11154;
  assign n11223 = ~i_nEMPTY & ~n11222;
  assign n11224 = ~n11221 & ~n11223;
  assign n11225 = i_FULL & ~n11224;
  assign n11226 = ~n8402 & ~n10005;
  assign n11227 = i_StoB_REQ9 & ~n11226;
  assign n11228 = controllable_BtoS_ACK11 & ~n9999;
  assign n11229 = ~controllable_BtoS_ACK11 & ~n11132;
  assign n11230 = ~n11228 & ~n11229;
  assign n11231 = n6661 & ~n11230;
  assign n11232 = ~n10769 & ~n11231;
  assign n11233 = i_StoB_REQ11 & ~n11232;
  assign n11234 = i_StoB_REQ10 & ~n9992;
  assign n11235 = i_StoB_REQ8 & ~n9983;
  assign n11236 = i_StoB_REQ7 & ~n9970;
  assign n11237 = i_StoB_REQ6 & ~n9963;
  assign n11238 = i_StoB_REQ5 & ~n9954;
  assign n11239 = controllable_BtoS_ACK4 & ~n9947;
  assign n11240 = ~controllable_BtoS_ACK4 & ~n11086;
  assign n11241 = ~n11239 & ~n11240;
  assign n11242 = n6667 & ~n11241;
  assign n11243 = ~n10780 & ~n11242;
  assign n11244 = i_StoB_REQ4 & ~n11243;
  assign n11245 = i_StoB_REQ3 & ~n9940;
  assign n11246 = i_StoB_REQ2 & ~n9931;
  assign n11247 = ~n9925 & ~n10785;
  assign n11248 = n6670 & ~n11247;
  assign n11249 = ~n10788 & ~n11248;
  assign n11250 = n6669 & ~n11249;
  assign n11251 = ~n8720 & ~n11250;
  assign n11252 = ~i_StoB_REQ2 & ~n11251;
  assign n11253 = ~n11246 & ~n11252;
  assign n11254 = controllable_BtoS_ACK2 & ~n11253;
  assign n11255 = i_StoB_REQ2 & ~n11072;
  assign n11256 = ~n11252 & ~n11255;
  assign n11257 = ~controllable_BtoS_ACK2 & ~n11256;
  assign n11258 = ~n11254 & ~n11257;
  assign n11259 = n6668 & ~n11258;
  assign n11260 = ~n8738 & ~n11259;
  assign n11261 = ~i_StoB_REQ3 & ~n11260;
  assign n11262 = ~n11245 & ~n11261;
  assign n11263 = controllable_BtoS_ACK3 & ~n11262;
  assign n11264 = i_StoB_REQ3 & ~n11080;
  assign n11265 = ~n11261 & ~n11264;
  assign n11266 = ~controllable_BtoS_ACK3 & ~n11265;
  assign n11267 = ~n11263 & ~n11266;
  assign n11268 = n6667 & ~n11267;
  assign n11269 = ~n10807 & ~n11268;
  assign n11270 = ~i_StoB_REQ4 & ~n11269;
  assign n11271 = ~n11244 & ~n11270;
  assign n11272 = n6666 & ~n11271;
  assign n11273 = ~n8787 & ~n11272;
  assign n11274 = ~i_StoB_REQ5 & ~n11273;
  assign n11275 = ~n11238 & ~n11274;
  assign n11276 = controllable_BtoS_ACK5 & ~n11275;
  assign n11277 = i_StoB_REQ5 & ~n11092;
  assign n11278 = ~n11274 & ~n11277;
  assign n11279 = ~controllable_BtoS_ACK5 & ~n11278;
  assign n11280 = ~n11276 & ~n11279;
  assign n11281 = n6665 & ~n11280;
  assign n11282 = ~n8814 & ~n11281;
  assign n11283 = ~i_StoB_REQ6 & ~n11282;
  assign n11284 = ~n11237 & ~n11283;
  assign n11285 = controllable_BtoS_ACK6 & ~n11284;
  assign n11286 = i_StoB_REQ6 & ~n11100;
  assign n11287 = ~n11283 & ~n11286;
  assign n11288 = ~controllable_BtoS_ACK6 & ~n11287;
  assign n11289 = ~n11285 & ~n11288;
  assign n11290 = ~i_StoB_REQ7 & ~n11289;
  assign n11291 = ~n11236 & ~n11290;
  assign n11292 = n6664 & ~n11291;
  assign n11293 = ~n10830 & ~n11292;
  assign n11294 = controllable_BtoS_ACK7 & ~n11293;
  assign n11295 = i_StoB_REQ7 & ~n11106;
  assign n11296 = ~n11290 & ~n11295;
  assign n11297 = n6664 & ~n11296;
  assign n11298 = ~n10835 & ~n11297;
  assign n11299 = ~controllable_BtoS_ACK7 & ~n11298;
  assign n11300 = ~n11294 & ~n11299;
  assign n11301 = n6663 & ~n11300;
  assign n11302 = ~n8877 & ~n11301;
  assign n11303 = ~i_StoB_REQ8 & ~n11302;
  assign n11304 = ~n11235 & ~n11303;
  assign n11305 = controllable_BtoS_ACK8 & ~n11304;
  assign n11306 = i_StoB_REQ8 & ~n11118;
  assign n11307 = ~n11303 & ~n11306;
  assign n11308 = ~controllable_BtoS_ACK8 & ~n11307;
  assign n11309 = ~n11305 & ~n11308;
  assign n11310 = n6662 & ~n11309;
  assign n11311 = ~n8906 & ~n11310;
  assign n11312 = ~i_StoB_REQ10 & ~n11311;
  assign n11313 = ~n11234 & ~n11312;
  assign n11314 = controllable_BtoS_ACK10 & ~n11313;
  assign n11315 = i_StoB_REQ10 & ~n11126;
  assign n11316 = ~n11312 & ~n11315;
  assign n11317 = ~controllable_BtoS_ACK10 & ~n11316;
  assign n11318 = ~n11314 & ~n11317;
  assign n11319 = n6661 & ~n11318;
  assign n11320 = ~n10856 & ~n11319;
  assign n11321 = ~i_StoB_REQ11 & ~n11320;
  assign n11322 = ~n11233 & ~n11321;
  assign n11323 = ~controllable_ENQ & ~n11322;
  assign n11324 = ~n11146 & ~n11323;
  assign n11325 = ~i_StoB_REQ9 & ~n11324;
  assign n11326 = ~n11227 & ~n11325;
  assign n11327 = controllable_BtoS_ACK9 & ~n11326;
  assign n11328 = ~controllable_ENQ & ~n11136;
  assign n11329 = ~n8039 & ~n11328;
  assign n11330 = i_StoB_REQ9 & ~n11329;
  assign n11331 = ~n11325 & ~n11330;
  assign n11332 = ~controllable_BtoS_ACK9 & ~n11331;
  assign n11333 = ~n11327 & ~n11332;
  assign n11334 = ~controllable_DEQ & ~n11333;
  assign n11335 = ~n10976 & ~n11334;
  assign n11336 = ~i_nEMPTY & ~n11335;
  assign n11337 = ~n11221 & ~n11336;
  assign n11338 = ~i_FULL & ~n11337;
  assign n11339 = ~n11225 & ~n11338;
  assign n11340 = ~i_RtoB_ACK0 & ~n11339;
  assign n11341 = ~n10958 & ~n11340;
  assign n11342 = n6660 & ~n11341;
  assign n11343 = ~n11212 & ~n11342;
  assign n11344 = ~n6659 & ~n11343;
  assign n11345 = ~n8149 & ~n11343;
  assign n11346 = ~n8149 & ~n11345;
  assign n11347 = n6659 & ~n11346;
  assign n11348 = ~n11344 & ~n11347;
  assign n11349 = ~n6651 & ~n11348;
  assign n11350 = ~n11219 & ~n11349;
  assign n11351 = ~controllable_BtoR_REQ0 & ~n11350;
  assign n11352 = ~controllable_BtoR_REQ0 & ~n11351;
  assign n11353 = ~i_RtoB_ACK1 & ~n11352;
  assign n11354 = ~n11187 & ~n11353;
  assign n11355 = controllable_BtoR_REQ1 & ~n11354;
  assign n11356 = i_RtoB_ACK0 & ~n11171;
  assign n11357 = ~n11209 & ~n11356;
  assign n11358 = n6660 & ~n11357;
  assign n11359 = ~n6660 & ~n11013;
  assign n11360 = ~n11358 & ~n11359;
  assign n11361 = ~n8149 & ~n11360;
  assign n11362 = ~n8149 & ~n11361;
  assign n11363 = ~n6659 & ~n11362;
  assign n11364 = n6659 & ~n11360;
  assign n11365 = ~n11363 & ~n11364;
  assign n11366 = n6652 & ~n11365;
  assign n11367 = ~n11012 & ~n11340;
  assign n11368 = n6660 & ~n11367;
  assign n11369 = ~n11359 & ~n11368;
  assign n11370 = ~n8149 & ~n11369;
  assign n11371 = ~n8149 & ~n11370;
  assign n11372 = ~n6659 & ~n11371;
  assign n11373 = n6659 & ~n11369;
  assign n11374 = ~n11372 & ~n11373;
  assign n11375 = ~n6652 & ~n11374;
  assign n11376 = ~n11366 & ~n11375;
  assign n11377 = controllable_BtoR_REQ0 & ~n11376;
  assign n11378 = ~n10377 & ~n11045;
  assign n11379 = i_nEMPTY & ~n11378;
  assign n11380 = ~n10385 & ~n11025;
  assign n11381 = ~i_nEMPTY & ~n11380;
  assign n11382 = ~n11379 & ~n11381;
  assign n11383 = i_FULL & ~n11382;
  assign n11384 = ~n11045 & ~n11203;
  assign n11385 = ~i_nEMPTY & ~n11384;
  assign n11386 = ~n11379 & ~n11385;
  assign n11387 = ~i_FULL & ~n11386;
  assign n11388 = ~n11383 & ~n11387;
  assign n11389 = ~i_RtoB_ACK0 & ~n11388;
  assign n11390 = ~n11020 & ~n11389;
  assign n11391 = n6660 & ~n11390;
  assign n11392 = ~n6660 & ~n11052;
  assign n11393 = ~n11391 & ~n11392;
  assign n11394 = n6652 & ~n11393;
  assign n11395 = ~n6659 & ~n11393;
  assign n11396 = ~n11045 & ~n11143;
  assign n11397 = i_nEMPTY & ~n11396;
  assign n11398 = ~n11025 & ~n11154;
  assign n11399 = ~i_nEMPTY & ~n11398;
  assign n11400 = ~n11397 & ~n11399;
  assign n11401 = i_FULL & ~n11400;
  assign n11402 = ~n11045 & ~n11334;
  assign n11403 = ~i_nEMPTY & ~n11402;
  assign n11404 = ~n11397 & ~n11403;
  assign n11405 = ~i_FULL & ~n11404;
  assign n11406 = ~n11401 & ~n11405;
  assign n11407 = ~i_RtoB_ACK0 & ~n11406;
  assign n11408 = ~n11020 & ~n11407;
  assign n11409 = n6660 & ~n11408;
  assign n11410 = ~n11392 & ~n11409;
  assign n11411 = n6659 & ~n11410;
  assign n11412 = ~n11395 & ~n11411;
  assign n11413 = ~n6652 & ~n11412;
  assign n11414 = ~n11394 & ~n11413;
  assign n11415 = n6651 & ~n11414;
  assign n11416 = ~n6659 & ~n11410;
  assign n11417 = n6659 & ~n11393;
  assign n11418 = ~n11416 & ~n11417;
  assign n11419 = n6652 & ~n11418;
  assign n11420 = ~n6652 & ~n11410;
  assign n11421 = ~n11419 & ~n11420;
  assign n11422 = ~n6651 & ~n11421;
  assign n11423 = ~n11415 & ~n11422;
  assign n11424 = ~controllable_BtoR_REQ0 & ~n11423;
  assign n11425 = ~n11377 & ~n11424;
  assign n11426 = ~i_RtoB_ACK1 & ~n11425;
  assign n11427 = ~n11011 & ~n11426;
  assign n11428 = ~controllable_BtoR_REQ1 & ~n11427;
  assign n11429 = ~n11355 & ~n11428;
  assign n11430 = n6649 & ~n11429;
  assign n11431 = ~n11040 & ~n11430;
  assign n11432 = ~n6647 & ~n11431;
  assign n11433 = ~n11061 & ~n11432;
  assign n11434 = ~n6646 & ~n11433;
  assign n11435 = ~n11044 & ~n11434;
  assign n11436 = n6642 & ~n11435;
  assign n11437 = controllable_DEQ & ~n9579;
  assign n11438 = ~n9531 & ~n11437;
  assign n11439 = i_nEMPTY & ~n11438;
  assign n11440 = ~n9549 & ~n10971;
  assign n11441 = ~i_nEMPTY & ~n11440;
  assign n11442 = ~n11439 & ~n11441;
  assign n11443 = i_FULL & ~n11442;
  assign n11444 = ~n9567 & ~n10962;
  assign n11445 = i_nEMPTY & ~n11444;
  assign n11446 = ~n9580 & ~n10976;
  assign n11447 = ~i_nEMPTY & ~n11446;
  assign n11448 = ~n11445 & ~n11447;
  assign n11449 = ~i_FULL & ~n11448;
  assign n11450 = ~n11443 & ~n11449;
  assign n11451 = ~i_RtoB_ACK0 & ~n11450;
  assign n11452 = ~n10958 & ~n11451;
  assign n11453 = n6660 & ~n11452;
  assign n11454 = controllable_DEQ & ~n9643;
  assign n11455 = ~n9609 & ~n11454;
  assign n11456 = i_nEMPTY & ~n11455;
  assign n11457 = ~n9622 & ~n10971;
  assign n11458 = ~i_nEMPTY & ~n11457;
  assign n11459 = ~n11456 & ~n11458;
  assign n11460 = i_FULL & ~n11459;
  assign n11461 = ~n9630 & ~n10962;
  assign n11462 = i_nEMPTY & ~n11461;
  assign n11463 = ~n9644 & ~n10976;
  assign n11464 = ~i_nEMPTY & ~n11463;
  assign n11465 = ~n11462 & ~n11464;
  assign n11466 = ~i_FULL & ~n11465;
  assign n11467 = ~n11460 & ~n11466;
  assign n11468 = ~i_RtoB_ACK0 & ~n11467;
  assign n11469 = ~n10958 & ~n11468;
  assign n11470 = ~n6660 & ~n11469;
  assign n11471 = ~n11453 & ~n11470;
  assign n11472 = ~n6659 & ~n11471;
  assign n11473 = ~n8149 & ~n11471;
  assign n11474 = ~n8149 & ~n11473;
  assign n11475 = n6659 & ~n11474;
  assign n11476 = ~n11472 & ~n11475;
  assign n11477 = n6651 & ~n11476;
  assign n11478 = ~n6651 & ~n10989;
  assign n11479 = ~n11477 & ~n11478;
  assign n11480 = ~controllable_BtoR_REQ0 & ~n11479;
  assign n11481 = ~controllable_BtoR_REQ0 & ~n11480;
  assign n11482 = ~i_RtoB_ACK1 & ~n11481;
  assign n11483 = ~n10937 & ~n11482;
  assign n11484 = controllable_BtoR_REQ1 & ~n11483;
  assign n11485 = ~n11012 & ~n11451;
  assign n11486 = n6660 & ~n11485;
  assign n11487 = ~n11012 & ~n11468;
  assign n11488 = ~n6660 & ~n11487;
  assign n11489 = ~n11486 & ~n11488;
  assign n11490 = ~n8149 & ~n11489;
  assign n11491 = ~n8149 & ~n11490;
  assign n11492 = ~n6659 & ~n11491;
  assign n11493 = n6659 & ~n11489;
  assign n11494 = ~n11492 & ~n11493;
  assign n11495 = n6652 & ~n11494;
  assign n11496 = ~n6652 & ~n11018;
  assign n11497 = ~n11495 & ~n11496;
  assign n11498 = controllable_BtoR_REQ0 & ~n11497;
  assign n11499 = controllable_DEQ & ~n9566;
  assign n11500 = ~n9531 & ~n11499;
  assign n11501 = i_nEMPTY & ~n11500;
  assign n11502 = ~n9549 & ~n11025;
  assign n11503 = ~i_nEMPTY & ~n11502;
  assign n11504 = ~n11501 & ~n11503;
  assign n11505 = i_FULL & ~n11504;
  assign n11506 = ~n9567 & ~n11045;
  assign n11507 = i_nEMPTY & ~n11506;
  assign n11508 = ~n9580 & ~n11045;
  assign n11509 = ~i_nEMPTY & ~n11508;
  assign n11510 = ~n11507 & ~n11509;
  assign n11511 = ~i_FULL & ~n11510;
  assign n11512 = ~n11505 & ~n11511;
  assign n11513 = ~i_RtoB_ACK0 & ~n11512;
  assign n11514 = ~n11020 & ~n11513;
  assign n11515 = n6660 & ~n11514;
  assign n11516 = controllable_DEQ & ~n9629;
  assign n11517 = ~n9609 & ~n11516;
  assign n11518 = i_nEMPTY & ~n11517;
  assign n11519 = ~n9622 & ~n11025;
  assign n11520 = ~i_nEMPTY & ~n11519;
  assign n11521 = ~n11518 & ~n11520;
  assign n11522 = i_FULL & ~n11521;
  assign n11523 = ~n9630 & ~n11045;
  assign n11524 = i_nEMPTY & ~n11523;
  assign n11525 = ~n9644 & ~n11045;
  assign n11526 = ~i_nEMPTY & ~n11525;
  assign n11527 = ~n11524 & ~n11526;
  assign n11528 = ~i_FULL & ~n11527;
  assign n11529 = ~n11522 & ~n11528;
  assign n11530 = ~i_RtoB_ACK0 & ~n11529;
  assign n11531 = ~n11020 & ~n11530;
  assign n11532 = ~n6660 & ~n11531;
  assign n11533 = ~n11515 & ~n11532;
  assign n11534 = n6652 & ~n11533;
  assign n11535 = ~n6659 & ~n11533;
  assign n11536 = n6659 & ~n11052;
  assign n11537 = ~n11535 & ~n11536;
  assign n11538 = ~n6652 & ~n11537;
  assign n11539 = ~n11534 & ~n11538;
  assign n11540 = n6651 & ~n11539;
  assign n11541 = ~n6659 & ~n11052;
  assign n11542 = n6659 & ~n11533;
  assign n11543 = ~n11541 & ~n11542;
  assign n11544 = n6652 & ~n11543;
  assign n11545 = ~n6652 & ~n11052;
  assign n11546 = ~n11544 & ~n11545;
  assign n11547 = ~n6651 & ~n11546;
  assign n11548 = ~n11540 & ~n11547;
  assign n11549 = ~controllable_BtoR_REQ0 & ~n11548;
  assign n11550 = ~n11498 & ~n11549;
  assign n11551 = ~i_RtoB_ACK1 & ~n11550;
  assign n11552 = ~n11011 & ~n11551;
  assign n11553 = ~controllable_BtoR_REQ1 & ~n11552;
  assign n11554 = ~n11484 & ~n11553;
  assign n11555 = n6649 & ~n11554;
  assign n11556 = ~i_FULL & ~n11506;
  assign n11557 = ~n11505 & ~n11556;
  assign n11558 = ~i_RtoB_ACK0 & ~n11557;
  assign n11559 = ~n11020 & ~n11558;
  assign n11560 = n6660 & ~n11559;
  assign n11561 = ~i_FULL & ~n11523;
  assign n11562 = ~n11522 & ~n11561;
  assign n11563 = ~i_RtoB_ACK0 & ~n11562;
  assign n11564 = ~n11020 & ~n11563;
  assign n11565 = ~n6660 & ~n11564;
  assign n11566 = ~n11560 & ~n11565;
  assign n11567 = n6652 & ~n11566;
  assign n11568 = ~n6659 & ~n11566;
  assign n11569 = n6659 & ~n11033;
  assign n11570 = ~n11568 & ~n11569;
  assign n11571 = ~n6652 & ~n11570;
  assign n11572 = ~n11567 & ~n11571;
  assign n11573 = n6651 & ~n11572;
  assign n11574 = ~n6659 & ~n11033;
  assign n11575 = n6659 & ~n11566;
  assign n11576 = ~n11574 & ~n11575;
  assign n11577 = n6652 & ~n11576;
  assign n11578 = ~n6652 & ~n11033;
  assign n11579 = ~n11577 & ~n11578;
  assign n11580 = ~n6651 & ~n11579;
  assign n11581 = ~n11573 & ~n11580;
  assign n11582 = ~controllable_BtoR_REQ0 & ~n11581;
  assign n11583 = ~n11498 & ~n11582;
  assign n11584 = ~i_RtoB_ACK1 & ~n11583;
  assign n11585 = ~n11011 & ~n11584;
  assign n11586 = ~controllable_BtoR_REQ1 & ~n11585;
  assign n11587 = ~n11484 & ~n11586;
  assign n11588 = ~n6649 & ~n11587;
  assign n11589 = ~n11555 & ~n11588;
  assign n11590 = n6647 & ~n11589;
  assign n11591 = ~controllable_DEQ & ~n10307;
  assign n11592 = ~n10365 & ~n11591;
  assign n11593 = i_nEMPTY & ~n11592;
  assign n11594 = controllable_ENQ & ~n10004;
  assign n11595 = controllable_ENQ & ~n11594;
  assign n11596 = ~i_StoB_REQ9 & ~n11595;
  assign n11597 = ~i_StoB_REQ9 & ~n11596;
  assign n11598 = controllable_BtoS_ACK9 & ~n11597;
  assign n11599 = ~n8404 & ~n11596;
  assign n11600 = ~controllable_BtoS_ACK9 & ~n11599;
  assign n11601 = ~n11598 & ~n11600;
  assign n11602 = ~controllable_DEQ & ~n11601;
  assign n11603 = ~controllable_DEQ & ~n11602;
  assign n11604 = ~i_nEMPTY & ~n11603;
  assign n11605 = ~n11593 & ~n11604;
  assign n11606 = i_RtoB_ACK0 & ~n11605;
  assign n11607 = ~n10291 & ~n10763;
  assign n11608 = ~i_StoB_REQ9 & ~n11607;
  assign n11609 = ~n10285 & ~n11608;
  assign n11610 = controllable_BtoS_ACK9 & ~n11609;
  assign n11611 = ~n10291 & ~n10674;
  assign n11612 = i_StoB_REQ9 & ~n11611;
  assign n11613 = ~n11608 & ~n11612;
  assign n11614 = ~controllable_BtoS_ACK9 & ~n11613;
  assign n11615 = ~n11610 & ~n11614;
  assign n11616 = ~controllable_DEQ & ~n11615;
  assign n11617 = ~n10344 & ~n11616;
  assign n11618 = ~i_nEMPTY & ~n11617;
  assign n11619 = ~n10379 & ~n11618;
  assign n11620 = ~i_FULL & ~n11619;
  assign n11621 = ~n10389 & ~n11620;
  assign n11622 = ~i_RtoB_ACK0 & ~n11621;
  assign n11623 = ~n11606 & ~n11622;
  assign n11624 = n6660 & ~n11623;
  assign n11625 = ~n11175 & ~n11624;
  assign n11626 = ~n6659 & ~n11625;
  assign n11627 = ~n8149 & ~n11625;
  assign n11628 = ~n8149 & ~n11627;
  assign n11629 = n6659 & ~n11628;
  assign n11630 = ~n11626 & ~n11629;
  assign n11631 = n6652 & ~n11630;
  assign n11632 = ~n11172 & ~n11606;
  assign n11633 = n6660 & ~n11632;
  assign n11634 = ~n11175 & ~n11633;
  assign n11635 = ~n6659 & ~n11634;
  assign n11636 = ~n8149 & ~n11634;
  assign n11637 = ~n8149 & ~n11636;
  assign n11638 = n6659 & ~n11637;
  assign n11639 = ~n11635 & ~n11638;
  assign n11640 = ~n6652 & ~n11639;
  assign n11641 = ~n11631 & ~n11640;
  assign n11642 = n6651 & ~n11641;
  assign n11643 = ~n6651 & ~n11181;
  assign n11644 = ~n11642 & ~n11643;
  assign n11645 = ~controllable_BtoR_REQ0 & ~n11644;
  assign n11646 = ~controllable_BtoR_REQ0 & ~n11645;
  assign n11647 = i_RtoB_ACK1 & ~n11646;
  assign n11648 = i_StoB_REQ9 & ~n10762;
  assign n11649 = ~i_StoB_REQ9 & ~n10859;
  assign n11650 = ~n11648 & ~n11649;
  assign n11651 = controllable_BtoS_ACK9 & ~n11650;
  assign n11652 = ~n10268 & ~n11649;
  assign n11653 = ~controllable_BtoS_ACK9 & ~n11652;
  assign n11654 = ~n11651 & ~n11653;
  assign n11655 = ~controllable_DEQ & ~n11654;
  assign n11656 = ~n10944 & ~n11655;
  assign n11657 = i_nEMPTY & ~n11656;
  assign n11658 = controllable_ENQ & ~n10762;
  assign n11659 = controllable_ENQ & ~n11658;
  assign n11660 = i_StoB_REQ9 & ~n11659;
  assign n11661 = controllable_ENQ & ~n10859;
  assign n11662 = controllable_ENQ & ~n11661;
  assign n11663 = ~i_StoB_REQ9 & ~n11662;
  assign n11664 = ~n11660 & ~n11663;
  assign n11665 = controllable_BtoS_ACK9 & ~n11664;
  assign n11666 = ~n10293 & ~n11663;
  assign n11667 = ~controllable_BtoS_ACK9 & ~n11666;
  assign n11668 = ~n11665 & ~n11667;
  assign n11669 = ~controllable_DEQ & ~n11668;
  assign n11670 = ~controllable_DEQ & ~n11669;
  assign n11671 = ~i_nEMPTY & ~n11670;
  assign n11672 = ~n11657 & ~n11671;
  assign n11673 = i_RtoB_ACK0 & ~n11672;
  assign n11674 = ~n10654 & ~n10962;
  assign n11675 = i_nEMPTY & ~n11674;
  assign n11676 = ~n10669 & ~n10971;
  assign n11677 = ~i_nEMPTY & ~n11676;
  assign n11678 = ~n11675 & ~n11677;
  assign n11679 = i_FULL & ~n11678;
  assign n11680 = ~n10684 & ~n10962;
  assign n11681 = i_nEMPTY & ~n11680;
  assign n11682 = ~n10869 & ~n10976;
  assign n11683 = ~i_nEMPTY & ~n11682;
  assign n11684 = ~n11681 & ~n11683;
  assign n11685 = ~i_FULL & ~n11684;
  assign n11686 = ~n11679 & ~n11685;
  assign n11687 = ~i_RtoB_ACK0 & ~n11686;
  assign n11688 = ~n11673 & ~n11687;
  assign n11689 = n6660 & ~n11688;
  assign n11690 = ~n9609 & ~n10962;
  assign n11691 = i_nEMPTY & ~n11690;
  assign n11692 = ~n11458 & ~n11691;
  assign n11693 = i_FULL & ~n11692;
  assign n11694 = ~n11466 & ~n11693;
  assign n11695 = ~i_RtoB_ACK0 & ~n11694;
  assign n11696 = ~n10958 & ~n11695;
  assign n11697 = ~n6660 & ~n11696;
  assign n11698 = ~n11689 & ~n11697;
  assign n11699 = ~n6659 & ~n11698;
  assign n11700 = ~n8149 & ~n11698;
  assign n11701 = ~n8149 & ~n11700;
  assign n11702 = n6659 & ~n11701;
  assign n11703 = ~n11699 & ~n11702;
  assign n11704 = n6651 & ~n11703;
  assign n11705 = ~n6651 & ~n11218;
  assign n11706 = ~n11704 & ~n11705;
  assign n11707 = ~controllable_BtoR_REQ0 & ~n11706;
  assign n11708 = ~controllable_BtoR_REQ0 & ~n11707;
  assign n11709 = ~i_RtoB_ACK1 & ~n11708;
  assign n11710 = ~n11647 & ~n11709;
  assign n11711 = controllable_BtoR_REQ1 & ~n11710;
  assign n11712 = ~i_RtoB_ACK0 & ~n11672;
  assign n11713 = ~n11606 & ~n11712;
  assign n11714 = n6660 & ~n11713;
  assign n11715 = ~n6660 & ~n10996;
  assign n11716 = ~n11714 & ~n11715;
  assign n11717 = ~n8149 & ~n11716;
  assign n11718 = ~n8149 & ~n11717;
  assign n11719 = ~n6659 & ~n11718;
  assign n11720 = n6659 & ~n11716;
  assign n11721 = ~n11719 & ~n11720;
  assign n11722 = n6652 & ~n11721;
  assign n11723 = ~n6652 & ~n11001;
  assign n11724 = ~n11722 & ~n11723;
  assign n11725 = controllable_BtoR_REQ0 & ~n11724;
  assign n11726 = ~n11003 & ~n11143;
  assign n11727 = i_nEMPTY & ~n11726;
  assign n11728 = ~controllable_DEQ & ~n11154;
  assign n11729 = ~i_nEMPTY & ~n11728;
  assign n11730 = ~n11727 & ~n11729;
  assign n11731 = n6660 & ~n11730;
  assign n11732 = ~n6660 & ~n11008;
  assign n11733 = ~n11731 & ~n11732;
  assign n11734 = ~controllable_BtoR_REQ0 & ~n11733;
  assign n11735 = ~n11725 & ~n11734;
  assign n11736 = i_RtoB_ACK1 & ~n11735;
  assign n11737 = i_RtoB_ACK0 & ~n11621;
  assign n11738 = ~n11687 & ~n11737;
  assign n11739 = n6660 & ~n11738;
  assign n11740 = ~n11012 & ~n11695;
  assign n11741 = ~n6660 & ~n11740;
  assign n11742 = ~n11739 & ~n11741;
  assign n11743 = ~n8149 & ~n11742;
  assign n11744 = ~n8149 & ~n11743;
  assign n11745 = ~n6659 & ~n11744;
  assign n11746 = n6659 & ~n11742;
  assign n11747 = ~n11745 & ~n11746;
  assign n11748 = n6652 & ~n11747;
  assign n11749 = ~n6652 & ~n11365;
  assign n11750 = ~n11748 & ~n11749;
  assign n11751 = n6651 & ~n11750;
  assign n11752 = ~n11356 & ~n11687;
  assign n11753 = n6660 & ~n11752;
  assign n11754 = ~n11741 & ~n11753;
  assign n11755 = ~n8149 & ~n11754;
  assign n11756 = ~n8149 & ~n11755;
  assign n11757 = ~n6659 & ~n11756;
  assign n11758 = n6659 & ~n11754;
  assign n11759 = ~n11757 & ~n11758;
  assign n11760 = n6652 & ~n11759;
  assign n11761 = ~n11749 & ~n11760;
  assign n11762 = ~n6651 & ~n11761;
  assign n11763 = ~n11751 & ~n11762;
  assign n11764 = controllable_BtoR_REQ0 & ~n11763;
  assign n11765 = i_RtoB_ACK0 & ~n11730;
  assign n11766 = ~n10654 & ~n11045;
  assign n11767 = i_nEMPTY & ~n11766;
  assign n11768 = ~n10669 & ~n11025;
  assign n11769 = ~i_nEMPTY & ~n11768;
  assign n11770 = ~n11767 & ~n11769;
  assign n11771 = i_FULL & ~n11770;
  assign n11772 = ~n10684 & ~n11045;
  assign n11773 = i_nEMPTY & ~n11772;
  assign n11774 = ~n10869 & ~n11045;
  assign n11775 = ~i_nEMPTY & ~n11774;
  assign n11776 = ~n11773 & ~n11775;
  assign n11777 = ~i_FULL & ~n11776;
  assign n11778 = ~n11771 & ~n11777;
  assign n11779 = ~i_RtoB_ACK0 & ~n11778;
  assign n11780 = ~n11765 & ~n11779;
  assign n11781 = n6660 & ~n11780;
  assign n11782 = ~n9609 & ~n11045;
  assign n11783 = i_nEMPTY & ~n11782;
  assign n11784 = ~n11520 & ~n11783;
  assign n11785 = i_FULL & ~n11784;
  assign n11786 = ~n11528 & ~n11785;
  assign n11787 = ~i_RtoB_ACK0 & ~n11786;
  assign n11788 = ~n11020 & ~n11787;
  assign n11789 = ~n6660 & ~n11788;
  assign n11790 = ~n11781 & ~n11789;
  assign n11791 = n6652 & ~n11790;
  assign n11792 = ~n6659 & ~n11790;
  assign n11793 = ~n11389 & ~n11765;
  assign n11794 = n6660 & ~n11793;
  assign n11795 = ~n11392 & ~n11794;
  assign n11796 = n6659 & ~n11795;
  assign n11797 = ~n11792 & ~n11796;
  assign n11798 = ~n6652 & ~n11797;
  assign n11799 = ~n11791 & ~n11798;
  assign n11800 = n6651 & ~n11799;
  assign n11801 = ~n6659 & ~n11795;
  assign n11802 = n6659 & ~n11790;
  assign n11803 = ~n11801 & ~n11802;
  assign n11804 = n6652 & ~n11803;
  assign n11805 = ~n6652 & ~n11795;
  assign n11806 = ~n11804 & ~n11805;
  assign n11807 = ~n6651 & ~n11806;
  assign n11808 = ~n11800 & ~n11807;
  assign n11809 = ~controllable_BtoR_REQ0 & ~n11808;
  assign n11810 = ~n11764 & ~n11809;
  assign n11811 = ~i_RtoB_ACK1 & ~n11810;
  assign n11812 = ~n11736 & ~n11811;
  assign n11813 = ~controllable_BtoR_REQ1 & ~n11812;
  assign n11814 = ~n11711 & ~n11813;
  assign n11815 = n6649 & ~n11814;
  assign n11816 = ~n11040 & ~n11815;
  assign n11817 = ~n6647 & ~n11816;
  assign n11818 = ~n11590 & ~n11817;
  assign n11819 = n6646 & ~n11818;
  assign n11820 = n6651 & ~n11348;
  assign n11821 = ~n11478 & ~n11820;
  assign n11822 = ~controllable_BtoR_REQ0 & ~n11821;
  assign n11823 = ~controllable_BtoR_REQ0 & ~n11822;
  assign n11824 = ~i_RtoB_ACK1 & ~n11823;
  assign n11825 = ~n10937 & ~n11824;
  assign n11826 = controllable_BtoR_REQ1 & ~n11825;
  assign n11827 = n6652 & ~n11374;
  assign n11828 = ~n11496 & ~n11827;
  assign n11829 = controllable_BtoR_REQ0 & ~n11828;
  assign n11830 = n6652 & ~n11410;
  assign n11831 = ~n11416 & ~n11536;
  assign n11832 = ~n6652 & ~n11831;
  assign n11833 = ~n11830 & ~n11832;
  assign n11834 = n6651 & ~n11833;
  assign n11835 = ~n11411 & ~n11541;
  assign n11836 = n6652 & ~n11835;
  assign n11837 = ~n11545 & ~n11836;
  assign n11838 = ~n6651 & ~n11837;
  assign n11839 = ~n11834 & ~n11838;
  assign n11840 = ~controllable_BtoR_REQ0 & ~n11839;
  assign n11841 = ~n11829 & ~n11840;
  assign n11842 = ~i_RtoB_ACK1 & ~n11841;
  assign n11843 = ~n11011 & ~n11842;
  assign n11844 = ~controllable_BtoR_REQ1 & ~n11843;
  assign n11845 = ~n11826 & ~n11844;
  assign n11846 = n6649 & ~n11845;
  assign n11847 = ~n11040 & ~n11846;
  assign n11848 = ~n6647 & ~n11847;
  assign n11849 = ~n11061 & ~n11848;
  assign n11850 = ~n6646 & ~n11849;
  assign n11851 = ~n11819 & ~n11850;
  assign n11852 = ~n6642 & ~n11851;
  assign n11853 = ~n11436 & ~n11852;
  assign n11854 = ~n6639 & ~n11853;
  assign n11855 = ~n6639 & ~n11854;
  assign n11856 = n6518 & n11855;
  assign n11857 = n6518 & ~n11856;
  assign inductivity_check  = ~n6399 & n11857;
endmodule


