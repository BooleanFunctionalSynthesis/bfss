// Generated using findDep.cpp 
module rankfunc61_unsigned_64 (v_1, v_2, v_3, v_4, v_5, v_6, v_7, v_8, v_9, v_10, v_11, v_12, v_13, v_14, v_15, v_16, v_17, v_18, v_19, v_20, v_21, v_22, v_23, v_24, v_25, v_26, v_27, v_28, v_29, v_30, v_31, v_32, v_33, v_34, v_35, v_36, v_37, v_38, v_39, v_40, v_41, v_42, v_43, v_44, v_45, v_46, v_47, v_48, v_49, v_50, v_51, v_52, v_53, v_54, v_55, v_56, v_57, v_58, v_59, v_60, v_61, v_62, v_63, v_64, v_65, v_66, v_67, v_68, v_69, v_70, v_71, v_72, v_73, v_74, v_75, v_76, v_77, v_78, v_79, v_80, v_81, v_82, v_83, v_84, v_85, v_86, v_87, v_88, v_89, v_90, v_91, v_92, v_93, v_94, v_95, v_96, v_97, v_98, v_99, v_100, v_101, v_102, v_103, v_104, v_105, v_106, v_107, v_108, v_109, v_110, v_111, v_112, v_113, v_114, v_115, v_116, v_117, v_118, v_119, v_120, v_121, v_122, v_123, v_124, v_125, v_126, v_127, v_128, v_129, v_130, v_131, v_132, v_133, v_134, v_135, v_136, v_137, v_138, v_139, v_140, v_141, v_142, v_143, v_144, v_145, v_146, v_147, v_148, v_149, v_150, v_151, v_152, v_153, v_154, v_155, v_156, v_157, v_158, v_159, v_160, v_161, v_162, v_163, v_164, v_165, v_166, v_167, v_168, v_169, v_170, v_171, v_172, v_173, v_174, v_175, v_176, v_177, v_178, v_179, v_180, v_181, v_182, v_183, v_184, v_185, v_186, v_187, v_188, v_189, v_190, v_191, v_192, v_193, v_194, v_195, v_196, v_197, v_198, v_199, v_200, v_201, v_202, v_203, v_204, v_205, v_206, v_207, v_208, v_209, v_210, v_211, v_212, v_213, v_214, v_215, v_216, v_217, v_218, v_219, v_220, v_221, v_222, v_223, v_224, v_225, v_226, v_227, v_228, v_229, v_230, v_231, v_232, v_233, v_234, v_235, v_236, v_237, v_238, v_239, v_240, v_241, v_242, v_243, v_244, v_245, v_246, v_247, v_248, v_249, v_250, v_251, v_252, v_253, v_254, v_255, v_256, v_257, v_258, v_259, v_260, v_261, v_262, v_263, v_264, v_265, v_266, v_267, v_268, v_269, v_270, v_271, v_272, v_273, v_274, v_275, v_276, v_277, v_278, v_279, v_280, v_281, v_282, v_283, v_284, v_285, v_286, v_287, v_288, v_289, v_290, v_291, v_292, v_293, v_294, v_295, v_296, v_297, v_298, v_299, v_300, v_301, v_302, v_303, v_304, v_305, v_306, v_307, v_308, v_309, v_310, v_311, v_312, v_313, v_314, v_315, v_316, v_317, v_318, v_319, v_320, v_321, v_322, v_323, v_324, v_325, v_326, v_327, v_328, v_329, v_330, v_331, v_332, v_333, v_334, v_335, v_336, v_337, v_338, v_339, v_340, v_341, v_342, v_343, v_344, v_345, v_346, v_347, v_348, v_349, v_350, v_351, v_352, v_353, v_354, v_355, v_356, v_357, v_358, v_359, v_360, v_361, v_362, v_363, v_364, v_365, v_366, v_367, v_368, v_369, v_370, v_371, v_372, v_373, v_374, v_375, v_376, v_377, v_378, v_379, v_380, v_381, v_382, v_383, v_384, v_385, v_386, v_387, v_388, v_389, v_390, v_391, v_392, v_393, v_394, v_395, v_396, v_397, v_398, v_399, v_400, v_401, v_402, v_403, v_404, v_405, v_406, v_407, v_408, v_409, v_410, v_411, v_412, v_413, v_414, v_415, v_416, v_417, v_418, v_419, v_420, v_421, v_422, v_423, v_424, v_425, v_426, v_427, v_428, v_429, v_430, v_431, v_432, v_433, v_434, v_435, v_436, v_437, v_438, v_439, v_440, v_441, v_442, v_443, v_444, v_445, v_446, v_447, v_448, v_450, v_451, v_452, v_453, v_454, v_455, v_456, v_457, v_458, v_459, v_460, v_461, v_462, v_463, v_464, v_465, v_466, v_467, v_468, v_469, v_470, v_471, v_472, v_473, v_474, v_475, v_476, v_477, v_478, v_479, v_480, v_481, v_482, v_483, v_484, v_485, v_486, v_487, v_488, v_489, v_490, v_491, v_492, v_493, v_494, v_495, v_496, v_497, v_498, v_499, v_500, v_501, v_502, v_503, v_504, v_505, v_506, v_507, v_508, v_509, v_510, v_511, v_512, v_513, v_514, v_515, v_516, v_517, v_518, v_519, v_520, v_521, v_522, v_523, v_524, v_525, v_526, v_527, v_528, v_529, v_530, v_531, v_532, v_533, v_534, v_535, v_536, v_537, v_538, v_539, v_540, v_541, v_542, v_543, v_544, v_545, v_546, v_547, v_548, v_549, v_550, v_551, v_552, v_553, v_554, v_555, v_556, v_557, v_558, v_559, v_560, v_561, v_562, v_563, v_564, v_565, v_566, v_567, v_568, v_569, v_570, v_571, v_572, v_573, v_574, v_575, v_576, v_577, v_1087, v_1216, v_1218, v_1219, v_1220, v_1221, v_1222, v_1223, v_1224, v_1225, v_1226, v_1227, v_1228, v_1229, v_1230, v_1231, v_1232, v_1233, v_1234, v_1235, v_1236, v_1237, v_1238, v_1239, v_1240, v_1241, v_1242, v_1243, v_1244, v_1245, v_1246, v_1247, v_1248, v_1249, v_1250, v_1251, v_1252, v_1253, v_1254, v_1255, v_1256, v_1257, v_1258, v_1259, v_1260, v_1261, v_1262, v_1263, v_1264, v_1265, v_1266, v_1267, v_1268, v_1269, v_1270, v_1271, v_1272, v_1273, v_1274, v_1275, v_1276, v_1277, v_1278, v_1279, v_1280, v_1281, v_1347, v_1348, v_1349, v_1350, v_1351, v_1352, v_1353, v_1354, v_1355, v_1356, v_1357, v_1358, v_1359, v_1360, v_1361, v_1362, v_1363, v_1364, v_1365, v_1366, v_1367, v_1368, v_1369, v_1370, v_1371, v_1372, v_1373, v_1374, v_1375, v_1376, v_1377, v_1378, v_1379, v_1380, v_1381, v_1382, v_1383, v_1384, v_1385, v_1386, v_1387, v_1388, v_1389, v_1390, v_1391, v_1392, v_1393, v_1394, v_1395, v_1396, v_1397, v_1398, v_1399, v_1400, v_1401, v_1402, v_1403, v_1404, v_1405, v_1406, v_1407, v_1408, v_1409, v_1410, v_1476, v_1477, v_1478, v_1479, v_1480, v_1481, v_1482, v_1483, v_1484, v_1485, v_1486, v_1487, v_1488, v_1489, v_1490, v_1491, v_1492, v_1493, v_1494, v_1495, v_1496, v_1497, v_1498, v_1499, v_1500, v_1501, v_1502, v_1503, v_1504, v_1505, v_1506, v_1507, v_1508, v_1509, v_1510, v_1511, v_1512, v_1513, v_1514, v_1515, v_1516, v_1517, v_1518, v_1519, v_1520, v_1521, v_1522, v_1523, v_1524, v_1525, v_1526, v_1527, v_1528, v_1529, v_1530, v_1531, v_1532, v_1533, v_1534, v_1535, v_1536, v_1537, v_1538, v_1539, v_2757, v_2758, v_2759, v_2760, v_2761, v_2762, v_2763, v_2764, v_2765, v_2766, v_2767, v_2768, v_2769, v_2770, v_2771, v_2772, v_2773, v_2774, v_2775, v_2776, v_2777, v_2778, v_2779, v_2780, v_2781, v_2782, v_2783, v_2784, v_2785, v_2786, v_2787, v_2788, v_2789, v_2790, v_2791, v_2792, v_2793, v_2794, v_2795, v_2796, v_2797, v_2798, v_2799, v_2800, v_2801, v_2802, v_2803, v_2804, v_2805, v_2806, v_2807, v_2808, v_2809, v_2810, v_2811, v_2812, v_2813, v_2814, v_2815, v_2816, v_2817, v_2818, v_2819, v_2820, v_2821, v_2822, v_2823, v_2824, v_2825, v_2826, v_2827, v_2828, v_2829, v_2830, v_2831, v_2832, v_2833, v_2834, v_2835, v_2836, v_2837, v_2838, v_2839, v_2840, v_2841, v_2842, v_2843, v_2844, v_2845, v_2846, v_2847, v_2848, v_2849, v_2850, v_2851, v_2852, v_2853, v_2854, v_2855, v_2856, v_2857, v_2858, v_2859, v_2860, v_2861, v_2862, v_2863, v_2864, v_2865, v_2866, v_2867, v_2868, v_2869, v_2870, v_2871, v_2872, v_2873, v_2874, v_2875, v_2876, v_2877, v_2878, v_2879, v_2880, v_2881, v_2882, v_2883, v_2884, v_3139, v_3141, v_3142, v_3143, v_3144, v_3145, v_3146, v_3147, v_3148, v_3149, v_3150, v_3151, v_3152, v_3153, v_3154, v_3155, v_3156, v_3157, v_3158, v_3159, v_3160, v_3161, v_3162, v_3163, v_3164, v_3165, v_3166, v_3167, v_3168, v_3169, v_3170, v_3171, v_3172, v_3173, v_3174, v_3175, v_3176, v_3177, v_3178, v_3179, v_3180, v_3181, v_3182, v_3183, v_3184, v_3185, v_3186, v_3187, v_3188, v_3189, v_3190, v_3191, v_3192, v_3193, v_3194, v_3195, v_3196, v_3197, v_3198, v_3199, v_3200, v_3201, v_3202, v_3203, v_3204, v_3205, v_3206, v_3207, v_3208, v_3209, v_3210, v_3211, v_3212, v_3213, v_3214, v_3215, v_3216, v_3217, v_3218, v_3219, v_3220, v_3221, v_3222, v_3223, v_3224, v_3225, v_3226, v_3227, v_3228, v_3229, v_3230, v_3231, v_3232, v_3233, v_3234, v_3235, v_3236, v_3237, v_3238, v_3239, v_3240, v_3241, v_3242, v_3243, v_3244, v_3245, v_3246, v_3247, v_3248, v_3249, v_3250, v_3251, v_3252, v_3253, v_3254, v_3255, v_3256, v_3257, v_3258, v_3259, v_3260, v_3261, v_3262, v_3263, v_3264, v_3265, v_3266, v_3267, v_3268, v_3523, v_3525, v_3526, v_3527, v_3528, v_3529, v_3530, v_3531, v_3532, v_3533, v_3534, v_3535, v_3536, v_3537, v_3538, v_3539, v_3540, v_3541, v_3542, v_3543, v_3544, v_3545, v_3546, v_3547, v_3548, v_3549, v_3550, v_3551, v_3552, v_3553, v_3554, v_3555, v_3556, v_3557, v_3558, v_3559, v_3560, v_3561, v_3562, v_3563, v_3564, v_3565, v_3566, v_3567, v_3568, v_3569, v_3570, v_3571, v_3572, v_3573, v_3574, v_3575, v_3576, v_3577, v_3578, v_3579, v_3580, v_3581, v_3582, v_3583, v_3584, v_3585, v_3586, v_3587, v_3588, v_3589, v_3590, v_3591, v_3592, v_3593, v_3594, v_3595, v_3596, v_3597, v_3598, v_3599, v_3600, v_3601, v_3602, v_3603, v_3604, v_3605, v_3606, v_3607, v_3608, v_3609, v_3610, v_3611, v_3612, v_3613, v_3614, v_3615, v_3616, v_3617, v_3618, v_3619, v_3620, v_3621, v_3622, v_3623, v_3624, v_3625, v_3626, v_3627, v_3628, v_3629, v_3630, v_3631, v_3632, v_3633, v_3634, v_3635, v_3636, v_3637, v_3638, v_3639, v_3640, v_3641, v_3642, v_3643, v_3644, v_3645, v_3646, v_3647, v_3648, v_3649, v_3650, v_3651, v_3652, v_3907, o_1);
input v_1;
input v_2;
input v_3;
input v_4;
input v_5;
input v_6;
input v_7;
input v_8;
input v_9;
input v_10;
input v_11;
input v_12;
input v_13;
input v_14;
input v_15;
input v_16;
input v_17;
input v_18;
input v_19;
input v_20;
input v_21;
input v_22;
input v_23;
input v_24;
input v_25;
input v_26;
input v_27;
input v_28;
input v_29;
input v_30;
input v_31;
input v_32;
input v_33;
input v_34;
input v_35;
input v_36;
input v_37;
input v_38;
input v_39;
input v_40;
input v_41;
input v_42;
input v_43;
input v_44;
input v_45;
input v_46;
input v_47;
input v_48;
input v_49;
input v_50;
input v_51;
input v_52;
input v_53;
input v_54;
input v_55;
input v_56;
input v_57;
input v_58;
input v_59;
input v_60;
input v_61;
input v_62;
input v_63;
input v_64;
input v_65;
input v_66;
input v_67;
input v_68;
input v_69;
input v_70;
input v_71;
input v_72;
input v_73;
input v_74;
input v_75;
input v_76;
input v_77;
input v_78;
input v_79;
input v_80;
input v_81;
input v_82;
input v_83;
input v_84;
input v_85;
input v_86;
input v_87;
input v_88;
input v_89;
input v_90;
input v_91;
input v_92;
input v_93;
input v_94;
input v_95;
input v_96;
input v_97;
input v_98;
input v_99;
input v_100;
input v_101;
input v_102;
input v_103;
input v_104;
input v_105;
input v_106;
input v_107;
input v_108;
input v_109;
input v_110;
input v_111;
input v_112;
input v_113;
input v_114;
input v_115;
input v_116;
input v_117;
input v_118;
input v_119;
input v_120;
input v_121;
input v_122;
input v_123;
input v_124;
input v_125;
input v_126;
input v_127;
input v_128;
input v_129;
input v_130;
input v_131;
input v_132;
input v_133;
input v_134;
input v_135;
input v_136;
input v_137;
input v_138;
input v_139;
input v_140;
input v_141;
input v_142;
input v_143;
input v_144;
input v_145;
input v_146;
input v_147;
input v_148;
input v_149;
input v_150;
input v_151;
input v_152;
input v_153;
input v_154;
input v_155;
input v_156;
input v_157;
input v_158;
input v_159;
input v_160;
input v_161;
input v_162;
input v_163;
input v_164;
input v_165;
input v_166;
input v_167;
input v_168;
input v_169;
input v_170;
input v_171;
input v_172;
input v_173;
input v_174;
input v_175;
input v_176;
input v_177;
input v_178;
input v_179;
input v_180;
input v_181;
input v_182;
input v_183;
input v_184;
input v_185;
input v_186;
input v_187;
input v_188;
input v_189;
input v_190;
input v_191;
input v_192;
input v_193;
input v_194;
input v_195;
input v_196;
input v_197;
input v_198;
input v_199;
input v_200;
input v_201;
input v_202;
input v_203;
input v_204;
input v_205;
input v_206;
input v_207;
input v_208;
input v_209;
input v_210;
input v_211;
input v_212;
input v_213;
input v_214;
input v_215;
input v_216;
input v_217;
input v_218;
input v_219;
input v_220;
input v_221;
input v_222;
input v_223;
input v_224;
input v_225;
input v_226;
input v_227;
input v_228;
input v_229;
input v_230;
input v_231;
input v_232;
input v_233;
input v_234;
input v_235;
input v_236;
input v_237;
input v_238;
input v_239;
input v_240;
input v_241;
input v_242;
input v_243;
input v_244;
input v_245;
input v_246;
input v_247;
input v_248;
input v_249;
input v_250;
input v_251;
input v_252;
input v_253;
input v_254;
input v_255;
input v_256;
input v_257;
input v_258;
input v_259;
input v_260;
input v_261;
input v_262;
input v_263;
input v_264;
input v_265;
input v_266;
input v_267;
input v_268;
input v_269;
input v_270;
input v_271;
input v_272;
input v_273;
input v_274;
input v_275;
input v_276;
input v_277;
input v_278;
input v_279;
input v_280;
input v_281;
input v_282;
input v_283;
input v_284;
input v_285;
input v_286;
input v_287;
input v_288;
input v_289;
input v_290;
input v_291;
input v_292;
input v_293;
input v_294;
input v_295;
input v_296;
input v_297;
input v_298;
input v_299;
input v_300;
input v_301;
input v_302;
input v_303;
input v_304;
input v_305;
input v_306;
input v_307;
input v_308;
input v_309;
input v_310;
input v_311;
input v_312;
input v_313;
input v_314;
input v_315;
input v_316;
input v_317;
input v_318;
input v_319;
input v_320;
input v_321;
input v_322;
input v_323;
input v_324;
input v_325;
input v_326;
input v_327;
input v_328;
input v_329;
input v_330;
input v_331;
input v_332;
input v_333;
input v_334;
input v_335;
input v_336;
input v_337;
input v_338;
input v_339;
input v_340;
input v_341;
input v_342;
input v_343;
input v_344;
input v_345;
input v_346;
input v_347;
input v_348;
input v_349;
input v_350;
input v_351;
input v_352;
input v_353;
input v_354;
input v_355;
input v_356;
input v_357;
input v_358;
input v_359;
input v_360;
input v_361;
input v_362;
input v_363;
input v_364;
input v_365;
input v_366;
input v_367;
input v_368;
input v_369;
input v_370;
input v_371;
input v_372;
input v_373;
input v_374;
input v_375;
input v_376;
input v_377;
input v_378;
input v_379;
input v_380;
input v_381;
input v_382;
input v_383;
input v_384;
input v_385;
input v_386;
input v_387;
input v_388;
input v_389;
input v_390;
input v_391;
input v_392;
input v_393;
input v_394;
input v_395;
input v_396;
input v_397;
input v_398;
input v_399;
input v_400;
input v_401;
input v_402;
input v_403;
input v_404;
input v_405;
input v_406;
input v_407;
input v_408;
input v_409;
input v_410;
input v_411;
input v_412;
input v_413;
input v_414;
input v_415;
input v_416;
input v_417;
input v_418;
input v_419;
input v_420;
input v_421;
input v_422;
input v_423;
input v_424;
input v_425;
input v_426;
input v_427;
input v_428;
input v_429;
input v_430;
input v_431;
input v_432;
input v_433;
input v_434;
input v_435;
input v_436;
input v_437;
input v_438;
input v_439;
input v_440;
input v_441;
input v_442;
input v_443;
input v_444;
input v_445;
input v_446;
input v_447;
input v_448;
input v_450;
input v_451;
input v_452;
input v_453;
input v_454;
input v_455;
input v_456;
input v_457;
input v_458;
input v_459;
input v_460;
input v_461;
input v_462;
input v_463;
input v_464;
input v_465;
input v_466;
input v_467;
input v_468;
input v_469;
input v_470;
input v_471;
input v_472;
input v_473;
input v_474;
input v_475;
input v_476;
input v_477;
input v_478;
input v_479;
input v_480;
input v_481;
input v_482;
input v_483;
input v_484;
input v_485;
input v_486;
input v_487;
input v_488;
input v_489;
input v_490;
input v_491;
input v_492;
input v_493;
input v_494;
input v_495;
input v_496;
input v_497;
input v_498;
input v_499;
input v_500;
input v_501;
input v_502;
input v_503;
input v_504;
input v_505;
input v_506;
input v_507;
input v_508;
input v_509;
input v_510;
input v_511;
input v_512;
input v_513;
input v_514;
input v_515;
input v_516;
input v_517;
input v_518;
input v_519;
input v_520;
input v_521;
input v_522;
input v_523;
input v_524;
input v_525;
input v_526;
input v_527;
input v_528;
input v_529;
input v_530;
input v_531;
input v_532;
input v_533;
input v_534;
input v_535;
input v_536;
input v_537;
input v_538;
input v_539;
input v_540;
input v_541;
input v_542;
input v_543;
input v_544;
input v_545;
input v_546;
input v_547;
input v_548;
input v_549;
input v_550;
input v_551;
input v_552;
input v_553;
input v_554;
input v_555;
input v_556;
input v_557;
input v_558;
input v_559;
input v_560;
input v_561;
input v_562;
input v_563;
input v_564;
input v_565;
input v_566;
input v_567;
input v_568;
input v_569;
input v_570;
input v_571;
input v_572;
input v_573;
input v_574;
input v_575;
input v_576;
input v_577;
input v_1087;
input v_1216;
input v_1218;
input v_1219;
input v_1220;
input v_1221;
input v_1222;
input v_1223;
input v_1224;
input v_1225;
input v_1226;
input v_1227;
input v_1228;
input v_1229;
input v_1230;
input v_1231;
input v_1232;
input v_1233;
input v_1234;
input v_1235;
input v_1236;
input v_1237;
input v_1238;
input v_1239;
input v_1240;
input v_1241;
input v_1242;
input v_1243;
input v_1244;
input v_1245;
input v_1246;
input v_1247;
input v_1248;
input v_1249;
input v_1250;
input v_1251;
input v_1252;
input v_1253;
input v_1254;
input v_1255;
input v_1256;
input v_1257;
input v_1258;
input v_1259;
input v_1260;
input v_1261;
input v_1262;
input v_1263;
input v_1264;
input v_1265;
input v_1266;
input v_1267;
input v_1268;
input v_1269;
input v_1270;
input v_1271;
input v_1272;
input v_1273;
input v_1274;
input v_1275;
input v_1276;
input v_1277;
input v_1278;
input v_1279;
input v_1280;
input v_1281;
input v_1347;
input v_1348;
input v_1349;
input v_1350;
input v_1351;
input v_1352;
input v_1353;
input v_1354;
input v_1355;
input v_1356;
input v_1357;
input v_1358;
input v_1359;
input v_1360;
input v_1361;
input v_1362;
input v_1363;
input v_1364;
input v_1365;
input v_1366;
input v_1367;
input v_1368;
input v_1369;
input v_1370;
input v_1371;
input v_1372;
input v_1373;
input v_1374;
input v_1375;
input v_1376;
input v_1377;
input v_1378;
input v_1379;
input v_1380;
input v_1381;
input v_1382;
input v_1383;
input v_1384;
input v_1385;
input v_1386;
input v_1387;
input v_1388;
input v_1389;
input v_1390;
input v_1391;
input v_1392;
input v_1393;
input v_1394;
input v_1395;
input v_1396;
input v_1397;
input v_1398;
input v_1399;
input v_1400;
input v_1401;
input v_1402;
input v_1403;
input v_1404;
input v_1405;
input v_1406;
input v_1407;
input v_1408;
input v_1409;
input v_1410;
input v_1476;
input v_1477;
input v_1478;
input v_1479;
input v_1480;
input v_1481;
input v_1482;
input v_1483;
input v_1484;
input v_1485;
input v_1486;
input v_1487;
input v_1488;
input v_1489;
input v_1490;
input v_1491;
input v_1492;
input v_1493;
input v_1494;
input v_1495;
input v_1496;
input v_1497;
input v_1498;
input v_1499;
input v_1500;
input v_1501;
input v_1502;
input v_1503;
input v_1504;
input v_1505;
input v_1506;
input v_1507;
input v_1508;
input v_1509;
input v_1510;
input v_1511;
input v_1512;
input v_1513;
input v_1514;
input v_1515;
input v_1516;
input v_1517;
input v_1518;
input v_1519;
input v_1520;
input v_1521;
input v_1522;
input v_1523;
input v_1524;
input v_1525;
input v_1526;
input v_1527;
input v_1528;
input v_1529;
input v_1530;
input v_1531;
input v_1532;
input v_1533;
input v_1534;
input v_1535;
input v_1536;
input v_1537;
input v_1538;
input v_1539;
input v_2757;
input v_2758;
input v_2759;
input v_2760;
input v_2761;
input v_2762;
input v_2763;
input v_2764;
input v_2765;
input v_2766;
input v_2767;
input v_2768;
input v_2769;
input v_2770;
input v_2771;
input v_2772;
input v_2773;
input v_2774;
input v_2775;
input v_2776;
input v_2777;
input v_2778;
input v_2779;
input v_2780;
input v_2781;
input v_2782;
input v_2783;
input v_2784;
input v_2785;
input v_2786;
input v_2787;
input v_2788;
input v_2789;
input v_2790;
input v_2791;
input v_2792;
input v_2793;
input v_2794;
input v_2795;
input v_2796;
input v_2797;
input v_2798;
input v_2799;
input v_2800;
input v_2801;
input v_2802;
input v_2803;
input v_2804;
input v_2805;
input v_2806;
input v_2807;
input v_2808;
input v_2809;
input v_2810;
input v_2811;
input v_2812;
input v_2813;
input v_2814;
input v_2815;
input v_2816;
input v_2817;
input v_2818;
input v_2819;
input v_2820;
input v_2821;
input v_2822;
input v_2823;
input v_2824;
input v_2825;
input v_2826;
input v_2827;
input v_2828;
input v_2829;
input v_2830;
input v_2831;
input v_2832;
input v_2833;
input v_2834;
input v_2835;
input v_2836;
input v_2837;
input v_2838;
input v_2839;
input v_2840;
input v_2841;
input v_2842;
input v_2843;
input v_2844;
input v_2845;
input v_2846;
input v_2847;
input v_2848;
input v_2849;
input v_2850;
input v_2851;
input v_2852;
input v_2853;
input v_2854;
input v_2855;
input v_2856;
input v_2857;
input v_2858;
input v_2859;
input v_2860;
input v_2861;
input v_2862;
input v_2863;
input v_2864;
input v_2865;
input v_2866;
input v_2867;
input v_2868;
input v_2869;
input v_2870;
input v_2871;
input v_2872;
input v_2873;
input v_2874;
input v_2875;
input v_2876;
input v_2877;
input v_2878;
input v_2879;
input v_2880;
input v_2881;
input v_2882;
input v_2883;
input v_2884;
input v_3139;
input v_3141;
input v_3142;
input v_3143;
input v_3144;
input v_3145;
input v_3146;
input v_3147;
input v_3148;
input v_3149;
input v_3150;
input v_3151;
input v_3152;
input v_3153;
input v_3154;
input v_3155;
input v_3156;
input v_3157;
input v_3158;
input v_3159;
input v_3160;
input v_3161;
input v_3162;
input v_3163;
input v_3164;
input v_3165;
input v_3166;
input v_3167;
input v_3168;
input v_3169;
input v_3170;
input v_3171;
input v_3172;
input v_3173;
input v_3174;
input v_3175;
input v_3176;
input v_3177;
input v_3178;
input v_3179;
input v_3180;
input v_3181;
input v_3182;
input v_3183;
input v_3184;
input v_3185;
input v_3186;
input v_3187;
input v_3188;
input v_3189;
input v_3190;
input v_3191;
input v_3192;
input v_3193;
input v_3194;
input v_3195;
input v_3196;
input v_3197;
input v_3198;
input v_3199;
input v_3200;
input v_3201;
input v_3202;
input v_3203;
input v_3204;
input v_3205;
input v_3206;
input v_3207;
input v_3208;
input v_3209;
input v_3210;
input v_3211;
input v_3212;
input v_3213;
input v_3214;
input v_3215;
input v_3216;
input v_3217;
input v_3218;
input v_3219;
input v_3220;
input v_3221;
input v_3222;
input v_3223;
input v_3224;
input v_3225;
input v_3226;
input v_3227;
input v_3228;
input v_3229;
input v_3230;
input v_3231;
input v_3232;
input v_3233;
input v_3234;
input v_3235;
input v_3236;
input v_3237;
input v_3238;
input v_3239;
input v_3240;
input v_3241;
input v_3242;
input v_3243;
input v_3244;
input v_3245;
input v_3246;
input v_3247;
input v_3248;
input v_3249;
input v_3250;
input v_3251;
input v_3252;
input v_3253;
input v_3254;
input v_3255;
input v_3256;
input v_3257;
input v_3258;
input v_3259;
input v_3260;
input v_3261;
input v_3262;
input v_3263;
input v_3264;
input v_3265;
input v_3266;
input v_3267;
input v_3268;
input v_3523;
input v_3525;
input v_3526;
input v_3527;
input v_3528;
input v_3529;
input v_3530;
input v_3531;
input v_3532;
input v_3533;
input v_3534;
input v_3535;
input v_3536;
input v_3537;
input v_3538;
input v_3539;
input v_3540;
input v_3541;
input v_3542;
input v_3543;
input v_3544;
input v_3545;
input v_3546;
input v_3547;
input v_3548;
input v_3549;
input v_3550;
input v_3551;
input v_3552;
input v_3553;
input v_3554;
input v_3555;
input v_3556;
input v_3557;
input v_3558;
input v_3559;
input v_3560;
input v_3561;
input v_3562;
input v_3563;
input v_3564;
input v_3565;
input v_3566;
input v_3567;
input v_3568;
input v_3569;
input v_3570;
input v_3571;
input v_3572;
input v_3573;
input v_3574;
input v_3575;
input v_3576;
input v_3577;
input v_3578;
input v_3579;
input v_3580;
input v_3581;
input v_3582;
input v_3583;
input v_3584;
input v_3585;
input v_3586;
input v_3587;
input v_3588;
input v_3589;
input v_3590;
input v_3591;
input v_3592;
input v_3593;
input v_3594;
input v_3595;
input v_3596;
input v_3597;
input v_3598;
input v_3599;
input v_3600;
input v_3601;
input v_3602;
input v_3603;
input v_3604;
input v_3605;
input v_3606;
input v_3607;
input v_3608;
input v_3609;
input v_3610;
input v_3611;
input v_3612;
input v_3613;
input v_3614;
input v_3615;
input v_3616;
input v_3617;
input v_3618;
input v_3619;
input v_3620;
input v_3621;
input v_3622;
input v_3623;
input v_3624;
input v_3625;
input v_3626;
input v_3627;
input v_3628;
input v_3629;
input v_3630;
input v_3631;
input v_3632;
input v_3633;
input v_3634;
input v_3635;
input v_3636;
input v_3637;
input v_3638;
input v_3639;
input v_3640;
input v_3641;
input v_3642;
input v_3643;
input v_3644;
input v_3645;
input v_3646;
input v_3647;
input v_3648;
input v_3649;
input v_3650;
input v_3651;
input v_3652;
input v_3907;
output o_1;
wire v_578;
wire v_579;
wire v_580;
wire v_581;
wire v_582;
wire v_583;
wire v_584;
wire v_585;
wire v_586;
wire v_587;
wire v_588;
wire v_589;
wire v_590;
wire v_591;
wire v_592;
wire v_593;
wire v_594;
wire v_595;
wire v_596;
wire v_597;
wire v_598;
wire v_599;
wire v_600;
wire v_601;
wire v_602;
wire v_603;
wire v_604;
wire v_605;
wire v_606;
wire v_607;
wire v_608;
wire v_609;
wire v_610;
wire v_611;
wire v_612;
wire v_613;
wire v_614;
wire v_615;
wire v_616;
wire v_617;
wire v_618;
wire v_619;
wire v_620;
wire v_621;
wire v_622;
wire v_623;
wire v_624;
wire v_625;
wire v_626;
wire v_627;
wire v_628;
wire v_629;
wire v_630;
wire v_631;
wire v_632;
wire v_633;
wire v_634;
wire v_635;
wire v_636;
wire v_637;
wire v_638;
wire v_639;
wire v_640;
wire v_641;
wire v_642;
wire v_643;
wire v_644;
wire v_645;
wire v_646;
wire v_647;
wire v_648;
wire v_649;
wire v_650;
wire v_651;
wire v_652;
wire v_653;
wire v_654;
wire v_655;
wire v_656;
wire v_657;
wire v_658;
wire v_659;
wire v_660;
wire v_661;
wire v_662;
wire v_663;
wire v_664;
wire v_665;
wire v_666;
wire v_667;
wire v_668;
wire v_669;
wire v_670;
wire v_671;
wire v_672;
wire v_673;
wire v_674;
wire v_675;
wire v_676;
wire v_677;
wire v_678;
wire v_679;
wire v_680;
wire v_681;
wire v_682;
wire v_683;
wire v_684;
wire v_685;
wire v_686;
wire v_687;
wire v_688;
wire v_689;
wire v_690;
wire v_691;
wire v_692;
wire v_693;
wire v_694;
wire v_695;
wire v_696;
wire v_697;
wire v_698;
wire v_699;
wire v_700;
wire v_701;
wire v_702;
wire v_703;
wire v_704;
wire v_705;
wire v_706;
wire v_707;
wire v_708;
wire v_709;
wire v_710;
wire v_711;
wire v_712;
wire v_713;
wire v_714;
wire v_715;
wire v_716;
wire v_717;
wire v_718;
wire v_719;
wire v_720;
wire v_721;
wire v_722;
wire v_723;
wire v_724;
wire v_725;
wire v_726;
wire v_727;
wire v_728;
wire v_729;
wire v_730;
wire v_731;
wire v_732;
wire v_733;
wire v_734;
wire v_735;
wire v_736;
wire v_737;
wire v_738;
wire v_739;
wire v_740;
wire v_741;
wire v_742;
wire v_743;
wire v_744;
wire v_745;
wire v_746;
wire v_747;
wire v_748;
wire v_749;
wire v_750;
wire v_751;
wire v_752;
wire v_753;
wire v_754;
wire v_755;
wire v_756;
wire v_757;
wire v_758;
wire v_759;
wire v_760;
wire v_761;
wire v_762;
wire v_763;
wire v_764;
wire v_765;
wire v_766;
wire v_767;
wire v_768;
wire v_769;
wire v_770;
wire v_771;
wire v_772;
wire v_773;
wire v_774;
wire v_775;
wire v_776;
wire v_777;
wire v_778;
wire v_779;
wire v_780;
wire v_781;
wire v_782;
wire v_783;
wire v_784;
wire v_785;
wire v_786;
wire v_787;
wire v_788;
wire v_789;
wire v_790;
wire v_791;
wire v_792;
wire v_793;
wire v_794;
wire v_795;
wire v_796;
wire v_797;
wire v_798;
wire v_799;
wire v_800;
wire v_801;
wire v_802;
wire v_803;
wire v_804;
wire v_805;
wire v_806;
wire v_807;
wire v_808;
wire v_809;
wire v_810;
wire v_811;
wire v_812;
wire v_813;
wire v_814;
wire v_815;
wire v_816;
wire v_817;
wire v_818;
wire v_819;
wire v_820;
wire v_821;
wire v_822;
wire v_823;
wire v_824;
wire v_825;
wire v_826;
wire v_827;
wire v_828;
wire v_829;
wire v_830;
wire v_831;
wire v_832;
wire v_833;
wire v_834;
wire v_835;
wire v_836;
wire v_837;
wire v_838;
wire v_839;
wire v_840;
wire v_841;
wire v_842;
wire v_843;
wire v_844;
wire v_845;
wire v_846;
wire v_847;
wire v_848;
wire v_849;
wire v_850;
wire v_851;
wire v_852;
wire v_853;
wire v_854;
wire v_855;
wire v_856;
wire v_857;
wire v_858;
wire v_859;
wire v_860;
wire v_861;
wire v_862;
wire v_863;
wire v_864;
wire v_865;
wire v_866;
wire v_867;
wire v_868;
wire v_869;
wire v_870;
wire v_871;
wire v_872;
wire v_873;
wire v_874;
wire v_875;
wire v_876;
wire v_877;
wire v_878;
wire v_879;
wire v_880;
wire v_881;
wire v_882;
wire v_883;
wire v_884;
wire v_885;
wire v_886;
wire v_887;
wire v_888;
wire v_889;
wire v_890;
wire v_891;
wire v_892;
wire v_893;
wire v_894;
wire v_895;
wire v_896;
wire v_897;
wire v_898;
wire v_899;
wire v_900;
wire v_901;
wire v_902;
wire v_903;
wire v_904;
wire v_905;
wire v_906;
wire v_907;
wire v_908;
wire v_909;
wire v_910;
wire v_911;
wire v_912;
wire v_913;
wire v_914;
wire v_915;
wire v_916;
wire v_917;
wire v_918;
wire v_919;
wire v_920;
wire v_921;
wire v_922;
wire v_923;
wire v_924;
wire v_925;
wire v_926;
wire v_927;
wire v_928;
wire v_929;
wire v_930;
wire v_931;
wire v_932;
wire v_933;
wire v_934;
wire v_935;
wire v_936;
wire v_937;
wire v_938;
wire v_939;
wire v_940;
wire v_941;
wire v_942;
wire v_943;
wire v_944;
wire v_945;
wire v_946;
wire v_947;
wire v_948;
wire v_949;
wire v_950;
wire v_951;
wire v_952;
wire v_953;
wire v_954;
wire v_955;
wire v_956;
wire v_957;
wire v_958;
wire v_959;
wire v_960;
wire v_961;
wire v_962;
wire v_963;
wire v_964;
wire v_965;
wire v_966;
wire v_967;
wire v_968;
wire v_969;
wire v_970;
wire v_971;
wire v_972;
wire v_973;
wire v_974;
wire v_975;
wire v_976;
wire v_977;
wire v_978;
wire v_979;
wire v_980;
wire v_981;
wire v_982;
wire v_983;
wire v_984;
wire v_985;
wire v_986;
wire v_987;
wire v_988;
wire v_989;
wire v_990;
wire v_991;
wire v_992;
wire v_993;
wire v_994;
wire v_995;
wire v_996;
wire v_997;
wire v_998;
wire v_999;
wire v_1000;
wire v_1001;
wire v_1002;
wire v_1003;
wire v_1004;
wire v_1005;
wire v_1006;
wire v_1007;
wire v_1008;
wire v_1009;
wire v_1010;
wire v_1011;
wire v_1012;
wire v_1013;
wire v_1014;
wire v_1015;
wire v_1016;
wire v_1017;
wire v_1018;
wire v_1019;
wire v_1020;
wire v_1021;
wire v_1022;
wire v_1023;
wire v_1024;
wire v_1025;
wire v_1026;
wire v_1027;
wire v_1028;
wire v_1029;
wire v_1030;
wire v_1031;
wire v_1032;
wire v_1033;
wire v_1034;
wire v_1035;
wire v_1036;
wire v_1037;
wire v_1038;
wire v_1039;
wire v_1040;
wire v_1041;
wire v_1042;
wire v_1043;
wire v_1044;
wire v_1045;
wire v_1046;
wire v_1047;
wire v_1048;
wire v_1049;
wire v_1050;
wire v_1051;
wire v_1052;
wire v_1053;
wire v_1054;
wire v_1055;
wire v_1056;
wire v_1057;
wire v_1058;
wire v_1059;
wire v_1060;
wire v_1061;
wire v_1062;
wire v_1063;
wire v_1064;
wire v_1065;
wire v_1066;
wire v_1067;
wire v_1068;
wire v_1069;
wire v_1070;
wire v_1071;
wire v_1072;
wire v_1073;
wire v_1074;
wire v_1075;
wire v_1076;
wire v_1077;
wire v_1078;
wire v_1079;
wire v_1080;
wire v_1081;
wire v_1082;
wire v_1083;
wire v_1084;
wire v_1085;
wire v_1086;
wire v_1088;
wire v_1089;
wire v_1090;
wire v_1091;
wire v_1092;
wire v_1093;
wire v_1094;
wire v_1095;
wire v_1096;
wire v_1097;
wire v_1098;
wire v_1099;
wire v_1100;
wire v_1101;
wire v_1102;
wire v_1103;
wire v_1104;
wire v_1105;
wire v_1106;
wire v_1107;
wire v_1108;
wire v_1109;
wire v_1110;
wire v_1111;
wire v_1112;
wire v_1113;
wire v_1114;
wire v_1115;
wire v_1116;
wire v_1117;
wire v_1118;
wire v_1119;
wire v_1120;
wire v_1121;
wire v_1122;
wire v_1123;
wire v_1124;
wire v_1125;
wire v_1126;
wire v_1127;
wire v_1128;
wire v_1129;
wire v_1130;
wire v_1131;
wire v_1132;
wire v_1133;
wire v_1134;
wire v_1135;
wire v_1136;
wire v_1137;
wire v_1138;
wire v_1139;
wire v_1140;
wire v_1141;
wire v_1142;
wire v_1143;
wire v_1144;
wire v_1145;
wire v_1146;
wire v_1147;
wire v_1148;
wire v_1149;
wire v_1150;
wire v_1151;
wire v_1152;
wire v_1153;
wire v_1154;
wire v_1155;
wire v_1156;
wire v_1157;
wire v_1158;
wire v_1159;
wire v_1160;
wire v_1161;
wire v_1162;
wire v_1163;
wire v_1164;
wire v_1165;
wire v_1166;
wire v_1167;
wire v_1168;
wire v_1169;
wire v_1170;
wire v_1171;
wire v_1172;
wire v_1173;
wire v_1174;
wire v_1175;
wire v_1176;
wire v_1177;
wire v_1178;
wire v_1179;
wire v_1180;
wire v_1181;
wire v_1182;
wire v_1183;
wire v_1184;
wire v_1185;
wire v_1186;
wire v_1187;
wire v_1188;
wire v_1189;
wire v_1190;
wire v_1191;
wire v_1192;
wire v_1193;
wire v_1194;
wire v_1195;
wire v_1196;
wire v_1197;
wire v_1198;
wire v_1199;
wire v_1200;
wire v_1201;
wire v_1202;
wire v_1203;
wire v_1204;
wire v_1205;
wire v_1206;
wire v_1207;
wire v_1208;
wire v_1209;
wire v_1210;
wire v_1211;
wire v_1212;
wire v_1213;
wire v_1214;
wire v_1215;
wire v_1217;
wire v_1282;
wire v_1283;
wire v_1284;
wire v_1285;
wire v_1286;
wire v_1287;
wire v_1288;
wire v_1289;
wire v_1290;
wire v_1291;
wire v_1292;
wire v_1293;
wire v_1294;
wire v_1295;
wire v_1296;
wire v_1297;
wire v_1298;
wire v_1299;
wire v_1300;
wire v_1301;
wire v_1302;
wire v_1303;
wire v_1304;
wire v_1305;
wire v_1306;
wire v_1307;
wire v_1308;
wire v_1309;
wire v_1310;
wire v_1311;
wire v_1312;
wire v_1313;
wire v_1314;
wire v_1315;
wire v_1316;
wire v_1317;
wire v_1318;
wire v_1319;
wire v_1320;
wire v_1321;
wire v_1322;
wire v_1323;
wire v_1324;
wire v_1325;
wire v_1326;
wire v_1327;
wire v_1328;
wire v_1329;
wire v_1330;
wire v_1331;
wire v_1332;
wire v_1333;
wire v_1334;
wire v_1335;
wire v_1336;
wire v_1337;
wire v_1338;
wire v_1339;
wire v_1340;
wire v_1341;
wire v_1342;
wire v_1343;
wire v_1344;
wire v_1345;
wire v_1346;
wire v_1411;
wire v_1412;
wire v_1413;
wire v_1414;
wire v_1415;
wire v_1416;
wire v_1417;
wire v_1418;
wire v_1419;
wire v_1420;
wire v_1421;
wire v_1422;
wire v_1423;
wire v_1424;
wire v_1425;
wire v_1426;
wire v_1427;
wire v_1428;
wire v_1429;
wire v_1430;
wire v_1431;
wire v_1432;
wire v_1433;
wire v_1434;
wire v_1435;
wire v_1436;
wire v_1437;
wire v_1438;
wire v_1439;
wire v_1440;
wire v_1441;
wire v_1442;
wire v_1443;
wire v_1444;
wire v_1445;
wire v_1446;
wire v_1447;
wire v_1448;
wire v_1449;
wire v_1450;
wire v_1451;
wire v_1452;
wire v_1453;
wire v_1454;
wire v_1455;
wire v_1456;
wire v_1457;
wire v_1458;
wire v_1459;
wire v_1460;
wire v_1461;
wire v_1462;
wire v_1463;
wire v_1464;
wire v_1465;
wire v_1466;
wire v_1467;
wire v_1468;
wire v_1469;
wire v_1470;
wire v_1471;
wire v_1472;
wire v_1473;
wire v_1474;
wire v_1475;
wire v_1540;
wire v_1541;
wire v_1542;
wire v_1543;
wire v_1544;
wire v_1545;
wire v_1546;
wire v_1547;
wire v_1548;
wire v_1549;
wire v_1550;
wire v_1551;
wire v_1552;
wire v_1553;
wire v_1554;
wire v_1555;
wire v_1556;
wire v_1557;
wire v_1558;
wire v_1559;
wire v_1560;
wire v_1561;
wire v_1562;
wire v_1563;
wire v_1564;
wire v_1565;
wire v_1566;
wire v_1567;
wire v_1568;
wire v_1569;
wire v_1570;
wire v_1571;
wire v_1572;
wire v_1573;
wire v_1574;
wire v_1575;
wire v_1576;
wire v_1577;
wire v_1578;
wire v_1579;
wire v_1580;
wire v_1581;
wire v_1582;
wire v_1583;
wire v_1584;
wire v_1585;
wire v_1586;
wire v_1587;
wire v_1588;
wire v_1589;
wire v_1590;
wire v_1591;
wire v_1592;
wire v_1593;
wire v_1594;
wire v_1595;
wire v_1596;
wire v_1597;
wire v_1598;
wire v_1599;
wire v_1600;
wire v_1601;
wire v_1602;
wire v_1603;
wire v_1604;
wire v_1605;
wire v_1606;
wire v_1607;
wire v_1608;
wire v_1609;
wire v_1610;
wire v_1611;
wire v_1612;
wire v_1613;
wire v_1614;
wire v_1615;
wire v_1616;
wire v_1617;
wire v_1618;
wire v_1619;
wire v_1620;
wire v_1621;
wire v_1622;
wire v_1623;
wire v_1624;
wire v_1625;
wire v_1626;
wire v_1627;
wire v_1628;
wire v_1629;
wire v_1630;
wire v_1631;
wire v_1632;
wire v_1633;
wire v_1634;
wire v_1635;
wire v_1636;
wire v_1637;
wire v_1638;
wire v_1639;
wire v_1640;
wire v_1641;
wire v_1642;
wire v_1643;
wire v_1644;
wire v_1645;
wire v_1646;
wire v_1647;
wire v_1648;
wire v_1649;
wire v_1650;
wire v_1651;
wire v_1652;
wire v_1653;
wire v_1654;
wire v_1655;
wire v_1656;
wire v_1657;
wire v_1658;
wire v_1659;
wire v_1660;
wire v_1661;
wire v_1662;
wire v_1663;
wire v_1664;
wire v_1665;
wire v_1666;
wire v_1667;
wire v_1668;
wire v_1669;
wire v_1670;
wire v_1671;
wire v_1672;
wire v_1673;
wire v_1674;
wire v_1675;
wire v_1676;
wire v_1677;
wire v_1678;
wire v_1679;
wire v_1680;
wire v_1681;
wire v_1682;
wire v_1683;
wire v_1684;
wire v_1685;
wire v_1686;
wire v_1687;
wire v_1688;
wire v_1689;
wire v_1690;
wire v_1691;
wire v_1692;
wire v_1693;
wire v_1694;
wire v_1695;
wire v_1696;
wire v_1697;
wire v_1698;
wire v_1699;
wire v_1700;
wire v_1701;
wire v_1702;
wire v_1703;
wire v_1704;
wire v_1705;
wire v_1706;
wire v_1707;
wire v_1708;
wire v_1709;
wire v_1710;
wire v_1711;
wire v_1712;
wire v_1713;
wire v_1714;
wire v_1715;
wire v_1716;
wire v_1717;
wire v_1718;
wire v_1719;
wire v_1720;
wire v_1721;
wire v_1722;
wire v_1723;
wire v_1724;
wire v_1725;
wire v_1726;
wire v_1727;
wire v_1728;
wire v_1729;
wire v_1730;
wire v_1731;
wire v_1732;
wire v_1733;
wire v_1734;
wire v_1735;
wire v_1736;
wire v_1737;
wire v_1738;
wire v_1739;
wire v_1740;
wire v_1741;
wire v_1742;
wire v_1743;
wire v_1744;
wire v_1745;
wire v_1746;
wire v_1747;
wire v_1748;
wire v_1749;
wire v_1750;
wire v_1751;
wire v_1752;
wire v_1753;
wire v_1754;
wire v_1755;
wire v_1756;
wire v_1757;
wire v_1758;
wire v_1759;
wire v_1760;
wire v_1761;
wire v_1762;
wire v_1763;
wire v_1764;
wire v_1765;
wire v_1766;
wire v_1767;
wire v_1768;
wire v_1769;
wire v_1770;
wire v_1771;
wire v_1772;
wire v_1773;
wire v_1774;
wire v_1775;
wire v_1776;
wire v_1777;
wire v_1778;
wire v_1779;
wire v_1780;
wire v_1781;
wire v_1782;
wire v_1783;
wire v_1784;
wire v_1785;
wire v_1786;
wire v_1787;
wire v_1788;
wire v_1789;
wire v_1790;
wire v_1791;
wire v_1792;
wire v_1793;
wire v_1794;
wire v_1795;
wire v_1796;
wire v_1797;
wire v_1798;
wire v_1799;
wire v_1800;
wire v_1801;
wire v_1802;
wire v_1803;
wire v_1804;
wire v_1805;
wire v_1806;
wire v_1807;
wire v_1808;
wire v_1809;
wire v_1810;
wire v_1811;
wire v_1812;
wire v_1813;
wire v_1814;
wire v_1815;
wire v_1816;
wire v_1817;
wire v_1818;
wire v_1819;
wire v_1820;
wire v_1821;
wire v_1822;
wire v_1823;
wire v_1824;
wire v_1825;
wire v_1826;
wire v_1827;
wire v_1828;
wire v_1829;
wire v_1830;
wire v_1831;
wire v_1832;
wire v_1833;
wire v_1834;
wire v_1835;
wire v_1836;
wire v_1837;
wire v_1838;
wire v_1839;
wire v_1840;
wire v_1841;
wire v_1842;
wire v_1843;
wire v_1844;
wire v_1845;
wire v_1846;
wire v_1847;
wire v_1848;
wire v_1849;
wire v_1850;
wire v_1851;
wire v_1852;
wire v_1853;
wire v_1854;
wire v_1855;
wire v_1856;
wire v_1857;
wire v_1858;
wire v_1859;
wire v_1860;
wire v_1861;
wire v_1862;
wire v_1863;
wire v_1864;
wire v_1865;
wire v_1866;
wire v_1867;
wire v_1868;
wire v_1869;
wire v_1870;
wire v_1871;
wire v_1872;
wire v_1873;
wire v_1874;
wire v_1875;
wire v_1876;
wire v_1877;
wire v_1878;
wire v_1879;
wire v_1880;
wire v_1881;
wire v_1882;
wire v_1883;
wire v_1884;
wire v_1885;
wire v_1886;
wire v_1887;
wire v_1888;
wire v_1889;
wire v_1890;
wire v_1891;
wire v_1892;
wire v_1893;
wire v_1894;
wire v_1895;
wire v_1896;
wire v_1897;
wire v_1898;
wire v_1899;
wire v_1900;
wire v_1901;
wire v_1902;
wire v_1903;
wire v_1904;
wire v_1905;
wire v_1906;
wire v_1907;
wire v_1908;
wire v_1909;
wire v_1910;
wire v_1911;
wire v_1912;
wire v_1913;
wire v_1914;
wire v_1915;
wire v_1916;
wire v_1917;
wire v_1918;
wire v_1919;
wire v_1920;
wire v_1921;
wire v_1922;
wire v_1923;
wire v_1924;
wire v_1925;
wire v_1926;
wire v_1927;
wire v_1928;
wire v_1929;
wire v_1930;
wire v_1931;
wire v_1932;
wire v_1933;
wire v_1934;
wire v_1935;
wire v_1936;
wire v_1937;
wire v_1938;
wire v_1939;
wire v_1940;
wire v_1941;
wire v_1942;
wire v_1943;
wire v_1944;
wire v_1945;
wire v_1946;
wire v_1947;
wire v_1948;
wire v_1949;
wire v_1950;
wire v_1951;
wire v_1952;
wire v_1953;
wire v_1954;
wire v_1955;
wire v_1956;
wire v_1957;
wire v_1958;
wire v_1959;
wire v_1960;
wire v_1961;
wire v_1962;
wire v_1963;
wire v_1964;
wire v_1965;
wire v_1966;
wire v_1967;
wire v_1968;
wire v_1969;
wire v_1970;
wire v_1971;
wire v_1972;
wire v_1973;
wire v_1974;
wire v_1975;
wire v_1976;
wire v_1977;
wire v_1978;
wire v_1979;
wire v_1980;
wire v_1981;
wire v_1982;
wire v_1983;
wire v_1984;
wire v_1985;
wire v_1986;
wire v_1987;
wire v_1988;
wire v_1989;
wire v_1990;
wire v_1991;
wire v_1992;
wire v_1993;
wire v_1994;
wire v_1995;
wire v_1996;
wire v_1997;
wire v_1998;
wire v_1999;
wire v_2000;
wire v_2001;
wire v_2002;
wire v_2003;
wire v_2004;
wire v_2005;
wire v_2006;
wire v_2007;
wire v_2008;
wire v_2009;
wire v_2010;
wire v_2011;
wire v_2012;
wire v_2013;
wire v_2014;
wire v_2015;
wire v_2016;
wire v_2017;
wire v_2018;
wire v_2019;
wire v_2020;
wire v_2021;
wire v_2022;
wire v_2023;
wire v_2024;
wire v_2025;
wire v_2026;
wire v_2027;
wire v_2028;
wire v_2029;
wire v_2030;
wire v_2031;
wire v_2032;
wire v_2033;
wire v_2034;
wire v_2035;
wire v_2036;
wire v_2037;
wire v_2038;
wire v_2039;
wire v_2040;
wire v_2041;
wire v_2042;
wire v_2043;
wire v_2044;
wire v_2045;
wire v_2046;
wire v_2047;
wire v_2048;
wire v_2049;
wire v_2050;
wire v_2051;
wire v_2052;
wire v_2053;
wire v_2054;
wire v_2055;
wire v_2056;
wire v_2057;
wire v_2058;
wire v_2059;
wire v_2060;
wire v_2061;
wire v_2062;
wire v_2063;
wire v_2064;
wire v_2065;
wire v_2066;
wire v_2067;
wire v_2068;
wire v_2069;
wire v_2070;
wire v_2071;
wire v_2072;
wire v_2073;
wire v_2074;
wire v_2075;
wire v_2076;
wire v_2077;
wire v_2078;
wire v_2079;
wire v_2080;
wire v_2081;
wire v_2082;
wire v_2083;
wire v_2084;
wire v_2085;
wire v_2086;
wire v_2087;
wire v_2088;
wire v_2089;
wire v_2090;
wire v_2091;
wire v_2092;
wire v_2093;
wire v_2094;
wire v_2095;
wire v_2096;
wire v_2097;
wire v_2098;
wire v_2099;
wire v_2100;
wire v_2101;
wire v_2102;
wire v_2103;
wire v_2104;
wire v_2105;
wire v_2106;
wire v_2107;
wire v_2108;
wire v_2109;
wire v_2110;
wire v_2111;
wire v_2112;
wire v_2113;
wire v_2114;
wire v_2115;
wire v_2116;
wire v_2117;
wire v_2118;
wire v_2119;
wire v_2120;
wire v_2121;
wire v_2122;
wire v_2123;
wire v_2124;
wire v_2125;
wire v_2126;
wire v_2127;
wire v_2128;
wire v_2129;
wire v_2130;
wire v_2131;
wire v_2132;
wire v_2133;
wire v_2134;
wire v_2135;
wire v_2136;
wire v_2137;
wire v_2138;
wire v_2139;
wire v_2140;
wire v_2141;
wire v_2142;
wire v_2143;
wire v_2144;
wire v_2145;
wire v_2146;
wire v_2147;
wire v_2148;
wire v_2149;
wire v_2150;
wire v_2151;
wire v_2152;
wire v_2153;
wire v_2154;
wire v_2155;
wire v_2156;
wire v_2157;
wire v_2158;
wire v_2159;
wire v_2160;
wire v_2161;
wire v_2162;
wire v_2163;
wire v_2164;
wire v_2165;
wire v_2166;
wire v_2167;
wire v_2168;
wire v_2169;
wire v_2170;
wire v_2171;
wire v_2172;
wire v_2173;
wire v_2174;
wire v_2175;
wire v_2176;
wire v_2177;
wire v_2178;
wire v_2179;
wire v_2180;
wire v_2181;
wire v_2182;
wire v_2183;
wire v_2184;
wire v_2185;
wire v_2186;
wire v_2187;
wire v_2188;
wire v_2189;
wire v_2190;
wire v_2191;
wire v_2192;
wire v_2193;
wire v_2194;
wire v_2195;
wire v_2196;
wire v_2197;
wire v_2198;
wire v_2199;
wire v_2200;
wire v_2201;
wire v_2202;
wire v_2203;
wire v_2204;
wire v_2205;
wire v_2206;
wire v_2207;
wire v_2208;
wire v_2209;
wire v_2210;
wire v_2211;
wire v_2212;
wire v_2213;
wire v_2214;
wire v_2215;
wire v_2216;
wire v_2217;
wire v_2218;
wire v_2219;
wire v_2220;
wire v_2221;
wire v_2222;
wire v_2223;
wire v_2224;
wire v_2225;
wire v_2226;
wire v_2227;
wire v_2228;
wire v_2229;
wire v_2230;
wire v_2231;
wire v_2232;
wire v_2233;
wire v_2234;
wire v_2235;
wire v_2236;
wire v_2237;
wire v_2238;
wire v_2239;
wire v_2240;
wire v_2241;
wire v_2242;
wire v_2243;
wire v_2244;
wire v_2245;
wire v_2246;
wire v_2247;
wire v_2248;
wire v_2249;
wire v_2250;
wire v_2251;
wire v_2252;
wire v_2253;
wire v_2254;
wire v_2255;
wire v_2256;
wire v_2257;
wire v_2258;
wire v_2259;
wire v_2260;
wire v_2261;
wire v_2262;
wire v_2263;
wire v_2264;
wire v_2265;
wire v_2266;
wire v_2267;
wire v_2268;
wire v_2269;
wire v_2270;
wire v_2271;
wire v_2272;
wire v_2273;
wire v_2274;
wire v_2275;
wire v_2276;
wire v_2277;
wire v_2278;
wire v_2279;
wire v_2280;
wire v_2281;
wire v_2282;
wire v_2283;
wire v_2284;
wire v_2285;
wire v_2286;
wire v_2287;
wire v_2288;
wire v_2289;
wire v_2290;
wire v_2291;
wire v_2292;
wire v_2293;
wire v_2294;
wire v_2295;
wire v_2296;
wire v_2297;
wire v_2298;
wire v_2299;
wire v_2300;
wire v_2301;
wire v_2302;
wire v_2303;
wire v_2304;
wire v_2305;
wire v_2306;
wire v_2307;
wire v_2308;
wire v_2309;
wire v_2310;
wire v_2311;
wire v_2312;
wire v_2313;
wire v_2314;
wire v_2315;
wire v_2316;
wire v_2317;
wire v_2318;
wire v_2319;
wire v_2320;
wire v_2321;
wire v_2322;
wire v_2323;
wire v_2324;
wire v_2325;
wire v_2326;
wire v_2327;
wire v_2328;
wire v_2329;
wire v_2330;
wire v_2331;
wire v_2332;
wire v_2333;
wire v_2334;
wire v_2335;
wire v_2336;
wire v_2337;
wire v_2338;
wire v_2339;
wire v_2340;
wire v_2341;
wire v_2342;
wire v_2343;
wire v_2344;
wire v_2345;
wire v_2346;
wire v_2347;
wire v_2348;
wire v_2349;
wire v_2350;
wire v_2351;
wire v_2352;
wire v_2353;
wire v_2354;
wire v_2355;
wire v_2356;
wire v_2357;
wire v_2358;
wire v_2359;
wire v_2360;
wire v_2361;
wire v_2362;
wire v_2363;
wire v_2364;
wire v_2365;
wire v_2366;
wire v_2367;
wire v_2368;
wire v_2369;
wire v_2370;
wire v_2371;
wire v_2372;
wire v_2373;
wire v_2374;
wire v_2375;
wire v_2376;
wire v_2377;
wire v_2378;
wire v_2379;
wire v_2380;
wire v_2381;
wire v_2382;
wire v_2383;
wire v_2384;
wire v_2385;
wire v_2386;
wire v_2387;
wire v_2388;
wire v_2389;
wire v_2390;
wire v_2391;
wire v_2392;
wire v_2393;
wire v_2394;
wire v_2395;
wire v_2396;
wire v_2397;
wire v_2398;
wire v_2399;
wire v_2400;
wire v_2401;
wire v_2402;
wire v_2403;
wire v_2404;
wire v_2405;
wire v_2406;
wire v_2407;
wire v_2408;
wire v_2409;
wire v_2410;
wire v_2411;
wire v_2412;
wire v_2413;
wire v_2414;
wire v_2415;
wire v_2416;
wire v_2417;
wire v_2418;
wire v_2419;
wire v_2420;
wire v_2421;
wire v_2422;
wire v_2423;
wire v_2424;
wire v_2425;
wire v_2426;
wire v_2427;
wire v_2428;
wire v_2429;
wire v_2430;
wire v_2431;
wire v_2432;
wire v_2433;
wire v_2434;
wire v_2435;
wire v_2436;
wire v_2437;
wire v_2438;
wire v_2439;
wire v_2440;
wire v_2441;
wire v_2442;
wire v_2443;
wire v_2444;
wire v_2445;
wire v_2446;
wire v_2447;
wire v_2448;
wire v_2449;
wire v_2450;
wire v_2451;
wire v_2452;
wire v_2453;
wire v_2454;
wire v_2455;
wire v_2456;
wire v_2457;
wire v_2458;
wire v_2459;
wire v_2460;
wire v_2461;
wire v_2462;
wire v_2463;
wire v_2464;
wire v_2465;
wire v_2466;
wire v_2467;
wire v_2468;
wire v_2469;
wire v_2470;
wire v_2471;
wire v_2472;
wire v_2473;
wire v_2474;
wire v_2475;
wire v_2476;
wire v_2477;
wire v_2478;
wire v_2479;
wire v_2480;
wire v_2481;
wire v_2482;
wire v_2483;
wire v_2484;
wire v_2485;
wire v_2486;
wire v_2487;
wire v_2488;
wire v_2489;
wire v_2490;
wire v_2491;
wire v_2492;
wire v_2493;
wire v_2494;
wire v_2495;
wire v_2496;
wire v_2497;
wire v_2498;
wire v_2499;
wire v_2500;
wire v_2501;
wire v_2502;
wire v_2503;
wire v_2504;
wire v_2505;
wire v_2506;
wire v_2507;
wire v_2508;
wire v_2509;
wire v_2510;
wire v_2511;
wire v_2512;
wire v_2513;
wire v_2514;
wire v_2515;
wire v_2516;
wire v_2517;
wire v_2518;
wire v_2519;
wire v_2520;
wire v_2521;
wire v_2522;
wire v_2523;
wire v_2524;
wire v_2525;
wire v_2526;
wire v_2527;
wire v_2528;
wire v_2529;
wire v_2530;
wire v_2531;
wire v_2532;
wire v_2533;
wire v_2534;
wire v_2535;
wire v_2536;
wire v_2537;
wire v_2538;
wire v_2539;
wire v_2540;
wire v_2541;
wire v_2542;
wire v_2543;
wire v_2544;
wire v_2545;
wire v_2546;
wire v_2547;
wire v_2548;
wire v_2549;
wire v_2550;
wire v_2551;
wire v_2552;
wire v_2553;
wire v_2554;
wire v_2555;
wire v_2556;
wire v_2557;
wire v_2558;
wire v_2559;
wire v_2560;
wire v_2561;
wire v_2562;
wire v_2563;
wire v_2564;
wire v_2565;
wire v_2566;
wire v_2567;
wire v_2568;
wire v_2569;
wire v_2570;
wire v_2571;
wire v_2572;
wire v_2573;
wire v_2574;
wire v_2575;
wire v_2576;
wire v_2577;
wire v_2578;
wire v_2579;
wire v_2580;
wire v_2581;
wire v_2582;
wire v_2583;
wire v_2584;
wire v_2585;
wire v_2586;
wire v_2587;
wire v_2588;
wire v_2589;
wire v_2590;
wire v_2591;
wire v_2592;
wire v_2593;
wire v_2594;
wire v_2595;
wire v_2596;
wire v_2597;
wire v_2598;
wire v_2599;
wire v_2600;
wire v_2601;
wire v_2602;
wire v_2603;
wire v_2604;
wire v_2605;
wire v_2606;
wire v_2607;
wire v_2608;
wire v_2609;
wire v_2610;
wire v_2611;
wire v_2612;
wire v_2613;
wire v_2614;
wire v_2615;
wire v_2616;
wire v_2617;
wire v_2618;
wire v_2619;
wire v_2620;
wire v_2621;
wire v_2622;
wire v_2623;
wire v_2624;
wire v_2625;
wire v_2626;
wire v_2627;
wire v_2628;
wire v_2629;
wire v_2630;
wire v_2631;
wire v_2632;
wire v_2633;
wire v_2634;
wire v_2635;
wire v_2636;
wire v_2637;
wire v_2638;
wire v_2639;
wire v_2640;
wire v_2641;
wire v_2642;
wire v_2643;
wire v_2644;
wire v_2645;
wire v_2646;
wire v_2647;
wire v_2648;
wire v_2649;
wire v_2650;
wire v_2651;
wire v_2652;
wire v_2653;
wire v_2654;
wire v_2655;
wire v_2656;
wire v_2657;
wire v_2658;
wire v_2659;
wire v_2660;
wire v_2661;
wire v_2662;
wire v_2663;
wire v_2664;
wire v_2665;
wire v_2666;
wire v_2667;
wire v_2668;
wire v_2669;
wire v_2670;
wire v_2671;
wire v_2672;
wire v_2673;
wire v_2674;
wire v_2675;
wire v_2676;
wire v_2677;
wire v_2678;
wire v_2679;
wire v_2680;
wire v_2681;
wire v_2682;
wire v_2683;
wire v_2684;
wire v_2685;
wire v_2686;
wire v_2687;
wire v_2688;
wire v_2689;
wire v_2690;
wire v_2691;
wire v_2692;
wire v_2693;
wire v_2694;
wire v_2695;
wire v_2696;
wire v_2697;
wire v_2698;
wire v_2699;
wire v_2700;
wire v_2701;
wire v_2702;
wire v_2703;
wire v_2704;
wire v_2705;
wire v_2706;
wire v_2707;
wire v_2708;
wire v_2709;
wire v_2710;
wire v_2711;
wire v_2712;
wire v_2713;
wire v_2714;
wire v_2715;
wire v_2716;
wire v_2717;
wire v_2718;
wire v_2719;
wire v_2720;
wire v_2721;
wire v_2722;
wire v_2723;
wire v_2724;
wire v_2725;
wire v_2726;
wire v_2727;
wire v_2728;
wire v_2729;
wire v_2730;
wire v_2731;
wire v_2732;
wire v_2733;
wire v_2734;
wire v_2735;
wire v_2736;
wire v_2737;
wire v_2738;
wire v_2739;
wire v_2740;
wire v_2741;
wire v_2742;
wire v_2743;
wire v_2744;
wire v_2745;
wire v_2746;
wire v_2747;
wire v_2748;
wire v_2749;
wire v_2750;
wire v_2751;
wire v_2752;
wire v_2753;
wire v_2754;
wire v_2755;
wire v_2756;
wire v_2885;
wire v_2886;
wire v_2887;
wire v_2888;
wire v_2889;
wire v_2890;
wire v_2891;
wire v_2892;
wire v_2893;
wire v_2894;
wire v_2895;
wire v_2896;
wire v_2897;
wire v_2898;
wire v_2899;
wire v_2900;
wire v_2901;
wire v_2902;
wire v_2903;
wire v_2904;
wire v_2905;
wire v_2906;
wire v_2907;
wire v_2908;
wire v_2909;
wire v_2910;
wire v_2911;
wire v_2912;
wire v_2913;
wire v_2914;
wire v_2915;
wire v_2916;
wire v_2917;
wire v_2918;
wire v_2919;
wire v_2920;
wire v_2921;
wire v_2922;
wire v_2923;
wire v_2924;
wire v_2925;
wire v_2926;
wire v_2927;
wire v_2928;
wire v_2929;
wire v_2930;
wire v_2931;
wire v_2932;
wire v_2933;
wire v_2934;
wire v_2935;
wire v_2936;
wire v_2937;
wire v_2938;
wire v_2939;
wire v_2940;
wire v_2941;
wire v_2942;
wire v_2943;
wire v_2944;
wire v_2945;
wire v_2946;
wire v_2947;
wire v_2948;
wire v_2949;
wire v_2950;
wire v_2951;
wire v_2952;
wire v_2953;
wire v_2954;
wire v_2955;
wire v_2956;
wire v_2957;
wire v_2958;
wire v_2959;
wire v_2960;
wire v_2961;
wire v_2962;
wire v_2963;
wire v_2964;
wire v_2965;
wire v_2966;
wire v_2967;
wire v_2968;
wire v_2969;
wire v_2970;
wire v_2971;
wire v_2972;
wire v_2973;
wire v_2974;
wire v_2975;
wire v_2976;
wire v_2977;
wire v_2978;
wire v_2979;
wire v_2980;
wire v_2981;
wire v_2982;
wire v_2983;
wire v_2984;
wire v_2985;
wire v_2986;
wire v_2987;
wire v_2988;
wire v_2989;
wire v_2990;
wire v_2991;
wire v_2992;
wire v_2993;
wire v_2994;
wire v_2995;
wire v_2996;
wire v_2997;
wire v_2998;
wire v_2999;
wire v_3000;
wire v_3001;
wire v_3002;
wire v_3003;
wire v_3004;
wire v_3005;
wire v_3006;
wire v_3007;
wire v_3008;
wire v_3009;
wire v_3010;
wire v_3011;
wire v_3012;
wire v_3013;
wire v_3014;
wire v_3015;
wire v_3016;
wire v_3017;
wire v_3018;
wire v_3019;
wire v_3020;
wire v_3021;
wire v_3022;
wire v_3023;
wire v_3024;
wire v_3025;
wire v_3026;
wire v_3027;
wire v_3028;
wire v_3029;
wire v_3030;
wire v_3031;
wire v_3032;
wire v_3033;
wire v_3034;
wire v_3035;
wire v_3036;
wire v_3037;
wire v_3038;
wire v_3039;
wire v_3040;
wire v_3041;
wire v_3042;
wire v_3043;
wire v_3044;
wire v_3045;
wire v_3046;
wire v_3047;
wire v_3048;
wire v_3049;
wire v_3050;
wire v_3051;
wire v_3052;
wire v_3053;
wire v_3054;
wire v_3055;
wire v_3056;
wire v_3057;
wire v_3058;
wire v_3059;
wire v_3060;
wire v_3061;
wire v_3062;
wire v_3063;
wire v_3064;
wire v_3065;
wire v_3066;
wire v_3067;
wire v_3068;
wire v_3069;
wire v_3070;
wire v_3071;
wire v_3072;
wire v_3073;
wire v_3074;
wire v_3075;
wire v_3076;
wire v_3077;
wire v_3078;
wire v_3079;
wire v_3080;
wire v_3081;
wire v_3082;
wire v_3083;
wire v_3084;
wire v_3085;
wire v_3086;
wire v_3087;
wire v_3088;
wire v_3089;
wire v_3090;
wire v_3091;
wire v_3092;
wire v_3093;
wire v_3094;
wire v_3095;
wire v_3096;
wire v_3097;
wire v_3098;
wire v_3099;
wire v_3100;
wire v_3101;
wire v_3102;
wire v_3103;
wire v_3104;
wire v_3105;
wire v_3106;
wire v_3107;
wire v_3108;
wire v_3109;
wire v_3110;
wire v_3111;
wire v_3112;
wire v_3113;
wire v_3114;
wire v_3115;
wire v_3116;
wire v_3117;
wire v_3118;
wire v_3119;
wire v_3120;
wire v_3121;
wire v_3122;
wire v_3123;
wire v_3124;
wire v_3125;
wire v_3126;
wire v_3127;
wire v_3128;
wire v_3129;
wire v_3130;
wire v_3131;
wire v_3132;
wire v_3133;
wire v_3134;
wire v_3135;
wire v_3136;
wire v_3137;
wire v_3138;
wire v_3140;
wire v_3269;
wire v_3270;
wire v_3271;
wire v_3272;
wire v_3273;
wire v_3274;
wire v_3275;
wire v_3276;
wire v_3277;
wire v_3278;
wire v_3279;
wire v_3280;
wire v_3281;
wire v_3282;
wire v_3283;
wire v_3284;
wire v_3285;
wire v_3286;
wire v_3287;
wire v_3288;
wire v_3289;
wire v_3290;
wire v_3291;
wire v_3292;
wire v_3293;
wire v_3294;
wire v_3295;
wire v_3296;
wire v_3297;
wire v_3298;
wire v_3299;
wire v_3300;
wire v_3301;
wire v_3302;
wire v_3303;
wire v_3304;
wire v_3305;
wire v_3306;
wire v_3307;
wire v_3308;
wire v_3309;
wire v_3310;
wire v_3311;
wire v_3312;
wire v_3313;
wire v_3314;
wire v_3315;
wire v_3316;
wire v_3317;
wire v_3318;
wire v_3319;
wire v_3320;
wire v_3321;
wire v_3322;
wire v_3323;
wire v_3324;
wire v_3325;
wire v_3326;
wire v_3327;
wire v_3328;
wire v_3329;
wire v_3330;
wire v_3331;
wire v_3332;
wire v_3333;
wire v_3334;
wire v_3335;
wire v_3336;
wire v_3337;
wire v_3338;
wire v_3339;
wire v_3340;
wire v_3341;
wire v_3342;
wire v_3343;
wire v_3344;
wire v_3345;
wire v_3346;
wire v_3347;
wire v_3348;
wire v_3349;
wire v_3350;
wire v_3351;
wire v_3352;
wire v_3353;
wire v_3354;
wire v_3355;
wire v_3356;
wire v_3357;
wire v_3358;
wire v_3359;
wire v_3360;
wire v_3361;
wire v_3362;
wire v_3363;
wire v_3364;
wire v_3365;
wire v_3366;
wire v_3367;
wire v_3368;
wire v_3369;
wire v_3370;
wire v_3371;
wire v_3372;
wire v_3373;
wire v_3374;
wire v_3375;
wire v_3376;
wire v_3377;
wire v_3378;
wire v_3379;
wire v_3380;
wire v_3381;
wire v_3382;
wire v_3383;
wire v_3384;
wire v_3385;
wire v_3386;
wire v_3387;
wire v_3388;
wire v_3389;
wire v_3390;
wire v_3391;
wire v_3392;
wire v_3393;
wire v_3394;
wire v_3395;
wire v_3396;
wire v_3397;
wire v_3398;
wire v_3399;
wire v_3400;
wire v_3401;
wire v_3402;
wire v_3403;
wire v_3404;
wire v_3405;
wire v_3406;
wire v_3407;
wire v_3408;
wire v_3409;
wire v_3410;
wire v_3411;
wire v_3412;
wire v_3413;
wire v_3414;
wire v_3415;
wire v_3416;
wire v_3417;
wire v_3418;
wire v_3419;
wire v_3420;
wire v_3421;
wire v_3422;
wire v_3423;
wire v_3424;
wire v_3425;
wire v_3426;
wire v_3427;
wire v_3428;
wire v_3429;
wire v_3430;
wire v_3431;
wire v_3432;
wire v_3433;
wire v_3434;
wire v_3435;
wire v_3436;
wire v_3437;
wire v_3438;
wire v_3439;
wire v_3440;
wire v_3441;
wire v_3442;
wire v_3443;
wire v_3444;
wire v_3445;
wire v_3446;
wire v_3447;
wire v_3448;
wire v_3449;
wire v_3450;
wire v_3451;
wire v_3452;
wire v_3453;
wire v_3454;
wire v_3455;
wire v_3456;
wire v_3457;
wire v_3458;
wire v_3459;
wire v_3460;
wire v_3461;
wire v_3462;
wire v_3463;
wire v_3464;
wire v_3465;
wire v_3466;
wire v_3467;
wire v_3468;
wire v_3469;
wire v_3470;
wire v_3471;
wire v_3472;
wire v_3473;
wire v_3474;
wire v_3475;
wire v_3476;
wire v_3477;
wire v_3478;
wire v_3479;
wire v_3480;
wire v_3481;
wire v_3482;
wire v_3483;
wire v_3484;
wire v_3485;
wire v_3486;
wire v_3487;
wire v_3488;
wire v_3489;
wire v_3490;
wire v_3491;
wire v_3492;
wire v_3493;
wire v_3494;
wire v_3495;
wire v_3496;
wire v_3497;
wire v_3498;
wire v_3499;
wire v_3500;
wire v_3501;
wire v_3502;
wire v_3503;
wire v_3504;
wire v_3505;
wire v_3506;
wire v_3507;
wire v_3508;
wire v_3509;
wire v_3510;
wire v_3511;
wire v_3512;
wire v_3513;
wire v_3514;
wire v_3515;
wire v_3516;
wire v_3517;
wire v_3518;
wire v_3519;
wire v_3520;
wire v_3521;
wire v_3522;
wire v_3524;
wire v_3653;
wire v_3654;
wire v_3655;
wire v_3656;
wire v_3657;
wire v_3658;
wire v_3659;
wire v_3660;
wire v_3661;
wire v_3662;
wire v_3663;
wire v_3664;
wire v_3665;
wire v_3666;
wire v_3667;
wire v_3668;
wire v_3669;
wire v_3670;
wire v_3671;
wire v_3672;
wire v_3673;
wire v_3674;
wire v_3675;
wire v_3676;
wire v_3677;
wire v_3678;
wire v_3679;
wire v_3680;
wire v_3681;
wire v_3682;
wire v_3683;
wire v_3684;
wire v_3685;
wire v_3686;
wire v_3687;
wire v_3688;
wire v_3689;
wire v_3690;
wire v_3691;
wire v_3692;
wire v_3693;
wire v_3694;
wire v_3695;
wire v_3696;
wire v_3697;
wire v_3698;
wire v_3699;
wire v_3700;
wire v_3701;
wire v_3702;
wire v_3703;
wire v_3704;
wire v_3705;
wire v_3706;
wire v_3707;
wire v_3708;
wire v_3709;
wire v_3710;
wire v_3711;
wire v_3712;
wire v_3713;
wire v_3714;
wire v_3715;
wire v_3716;
wire v_3717;
wire v_3718;
wire v_3719;
wire v_3720;
wire v_3721;
wire v_3722;
wire v_3723;
wire v_3724;
wire v_3725;
wire v_3726;
wire v_3727;
wire v_3728;
wire v_3729;
wire v_3730;
wire v_3731;
wire v_3732;
wire v_3733;
wire v_3734;
wire v_3735;
wire v_3736;
wire v_3737;
wire v_3738;
wire v_3739;
wire v_3740;
wire v_3741;
wire v_3742;
wire v_3743;
wire v_3744;
wire v_3745;
wire v_3746;
wire v_3747;
wire v_3748;
wire v_3749;
wire v_3750;
wire v_3751;
wire v_3752;
wire v_3753;
wire v_3754;
wire v_3755;
wire v_3756;
wire v_3757;
wire v_3758;
wire v_3759;
wire v_3760;
wire v_3761;
wire v_3762;
wire v_3763;
wire v_3764;
wire v_3765;
wire v_3766;
wire v_3767;
wire v_3768;
wire v_3769;
wire v_3770;
wire v_3771;
wire v_3772;
wire v_3773;
wire v_3774;
wire v_3775;
wire v_3776;
wire v_3777;
wire v_3778;
wire v_3779;
wire v_3780;
wire v_3781;
wire v_3782;
wire v_3783;
wire v_3784;
wire v_3785;
wire v_3786;
wire v_3787;
wire v_3788;
wire v_3789;
wire v_3790;
wire v_3791;
wire v_3792;
wire v_3793;
wire v_3794;
wire v_3795;
wire v_3796;
wire v_3797;
wire v_3798;
wire v_3799;
wire v_3800;
wire v_3801;
wire v_3802;
wire v_3803;
wire v_3804;
wire v_3805;
wire v_3806;
wire v_3807;
wire v_3808;
wire v_3809;
wire v_3810;
wire v_3811;
wire v_3812;
wire v_3813;
wire v_3814;
wire v_3815;
wire v_3816;
wire v_3817;
wire v_3818;
wire v_3819;
wire v_3820;
wire v_3821;
wire v_3822;
wire v_3823;
wire v_3824;
wire v_3825;
wire v_3826;
wire v_3827;
wire v_3828;
wire v_3829;
wire v_3830;
wire v_3831;
wire v_3832;
wire v_3833;
wire v_3834;
wire v_3835;
wire v_3836;
wire v_3837;
wire v_3838;
wire v_3839;
wire v_3840;
wire v_3841;
wire v_3842;
wire v_3843;
wire v_3844;
wire v_3845;
wire v_3846;
wire v_3847;
wire v_3848;
wire v_3849;
wire v_3850;
wire v_3851;
wire v_3852;
wire v_3853;
wire v_3854;
wire v_3855;
wire v_3856;
wire v_3857;
wire v_3858;
wire v_3859;
wire v_3860;
wire v_3861;
wire v_3862;
wire v_3863;
wire v_3864;
wire v_3865;
wire v_3866;
wire v_3867;
wire v_3868;
wire v_3869;
wire v_3870;
wire v_3871;
wire v_3872;
wire v_3873;
wire v_3874;
wire v_3875;
wire v_3876;
wire v_3877;
wire v_3878;
wire v_3879;
wire v_3880;
wire v_3881;
wire v_3882;
wire v_3883;
wire v_3884;
wire v_3885;
wire v_3886;
wire v_3887;
wire v_3888;
wire v_3889;
wire v_3890;
wire v_3891;
wire v_3892;
wire v_3893;
wire v_3894;
wire v_3895;
wire v_3896;
wire v_3897;
wire v_3898;
wire v_3899;
wire v_3900;
wire v_3901;
wire v_3902;
wire v_3903;
wire v_3904;
wire v_3905;
wire v_3906;
wire v_3908;
wire v_3909;
wire v_3910;
wire v_3911;
wire v_3912;
wire v_3913;
wire v_3914;
wire v_3915;
wire v_3916;
wire v_3917;
wire v_3918;
wire v_3919;
wire v_3920;
wire v_3921;
wire v_3922;
wire v_3923;
wire v_3924;
wire v_3925;
wire v_3926;
wire v_3927;
wire v_3928;
wire v_3929;
wire v_3930;
wire v_3931;
wire v_3932;
wire v_3933;
wire v_3934;
wire v_3935;
wire v_3936;
wire v_3937;
wire v_3938;
wire v_3939;
wire v_3940;
wire v_3941;
wire v_3942;
wire v_3943;
wire v_3944;
wire v_3945;
wire v_3946;
wire v_3947;
wire v_3948;
wire v_3949;
wire v_3950;
wire v_3951;
wire v_3952;
wire v_3953;
wire v_3954;
wire v_3955;
wire v_3956;
wire v_3957;
wire v_3958;
wire v_3959;
wire v_3960;
wire v_3961;
wire v_3962;
wire v_3963;
wire v_3964;
wire v_3965;
wire v_3966;
wire v_3967;
wire v_3968;
wire v_3969;
wire v_3970;
wire v_3971;
wire v_3972;
wire v_3973;
wire v_3974;
wire v_3975;
wire v_3976;
wire v_3977;
wire v_3978;
wire v_3979;
wire v_3980;
wire v_3981;
wire v_3982;
wire v_3983;
wire v_3984;
wire v_3985;
wire v_3986;
wire v_3987;
wire v_3988;
wire v_3989;
wire v_3990;
wire v_3991;
wire v_3992;
wire v_3993;
wire v_3994;
wire v_3995;
wire v_3996;
wire v_3997;
wire v_3998;
wire v_3999;
wire v_4000;
wire v_4001;
wire v_4002;
wire v_4003;
wire v_4004;
wire v_4005;
wire v_4006;
wire v_4007;
wire v_4008;
wire v_4009;
wire v_4010;
wire v_4011;
wire v_4012;
wire v_4013;
wire v_4014;
wire v_4015;
wire v_4016;
wire v_4017;
wire v_4018;
wire v_4019;
wire v_4020;
wire v_4021;
wire v_4022;
wire v_4023;
wire v_4024;
wire v_4025;
wire v_4026;
wire v_4027;
wire v_4028;
wire v_4029;
wire v_4030;
wire v_4031;
wire v_4032;
wire v_4033;
wire v_4034;
wire v_4035;
wire v_4036;
wire v_4037;
wire v_4038;
wire v_4039;
wire v_4040;
wire v_4041;
wire v_4042;
wire v_4043;
wire v_4044;
wire v_4045;
wire v_4046;
wire v_4047;
wire v_4048;
wire v_4049;
wire v_4050;
wire v_4051;
wire v_4052;
wire v_4053;
wire v_4054;
wire v_4055;
wire v_4056;
wire v_4057;
wire v_4058;
wire v_4059;
wire v_4060;
wire v_4061;
wire v_4062;
wire v_4063;
wire v_4064;
wire v_4065;
wire v_4066;
wire v_4067;
wire v_4068;
wire v_4069;
wire v_4070;
wire v_4071;
wire v_4072;
wire v_4073;
wire v_4074;
wire v_4075;
wire v_4076;
wire v_4077;
wire v_4078;
wire v_4079;
wire v_4080;
wire v_4081;
wire v_4082;
wire v_4083;
wire v_4084;
wire v_4085;
wire v_4086;
wire v_4087;
wire v_4088;
wire v_4089;
wire v_4090;
wire v_4091;
wire v_4092;
wire v_4093;
wire v_4094;
wire v_4095;
wire v_4096;
wire v_4097;
wire v_4098;
wire v_4099;
wire v_4100;
wire v_4101;
wire v_4102;
wire v_4103;
wire v_4104;
wire v_4105;
wire v_4106;
wire v_4107;
wire v_4108;
wire v_4109;
wire v_4110;
wire v_4111;
wire v_4112;
wire v_4113;
wire v_4114;
wire v_4115;
wire v_4116;
wire v_4117;
wire v_4118;
wire v_4119;
wire v_4120;
wire v_4121;
wire v_4122;
wire v_4123;
wire v_4124;
wire v_4125;
wire v_4126;
wire v_4127;
wire v_4128;
wire v_4129;
wire v_4130;
wire v_4131;
wire v_4132;
wire v_4133;
wire v_4134;
wire v_4135;
wire v_4136;
wire v_4137;
wire v_4138;
wire v_4139;
wire v_4140;
wire v_4141;
wire v_4142;
wire v_4143;
wire v_4144;
wire v_4145;
wire v_4146;
wire v_4147;
wire v_4148;
wire v_4149;
wire v_4150;
wire v_4151;
wire v_4152;
wire v_4153;
wire v_4154;
wire v_4155;
wire v_4156;
wire v_4157;
wire v_4158;
wire v_4159;
wire v_4160;
wire v_4161;
wire v_4162;
wire v_4163;
wire v_4164;
wire v_4165;
wire v_4166;
wire v_4167;
wire v_4168;
wire v_4169;
wire v_4170;
wire v_4171;
wire v_4172;
wire v_4173;
wire v_4174;
wire v_4175;
wire v_4176;
wire v_4177;
wire v_4178;
wire v_4179;
wire v_4180;
wire v_4181;
wire v_4182;
wire v_4183;
wire v_4184;
wire v_4185;
wire v_4186;
wire v_4187;
wire v_4188;
wire v_4189;
wire v_4190;
wire v_4191;
wire v_4192;
wire v_4193;
wire v_4194;
wire v_4195;
wire v_4196;
wire v_4197;
wire v_4198;
wire v_4199;
wire v_4200;
wire v_4201;
wire v_4202;
wire v_4203;
wire v_4204;
wire v_4205;
wire v_4206;
wire v_4207;
wire v_4208;
wire v_4209;
wire v_4210;
wire v_4211;
wire v_4212;
wire v_4213;
wire v_4214;
wire v_4215;
wire v_4216;
wire v_4217;
wire v_4218;
wire v_4219;
wire v_4220;
wire v_4221;
wire v_4222;
wire v_4223;
wire v_4224;
wire v_4225;
wire v_4226;
wire v_4227;
wire v_4228;
wire v_4229;
wire v_4230;
wire v_4231;
wire v_4232;
wire v_4233;
wire v_4234;
wire v_4235;
wire v_4236;
wire v_4237;
wire v_4238;
wire v_4239;
wire v_4240;
wire v_4241;
wire v_4242;
wire v_4243;
wire v_4244;
wire v_4245;
wire v_4246;
wire v_4247;
wire v_4248;
wire v_4249;
wire v_4250;
wire v_4251;
wire v_4252;
wire v_4253;
wire v_4254;
wire v_4255;
wire v_4256;
wire v_4257;
wire v_4258;
wire v_4259;
wire v_4260;
wire v_4261;
wire v_4262;
wire v_4263;
wire v_4264;
wire v_4265;
wire v_4266;
wire v_4267;
wire v_4268;
wire v_4269;
wire v_4270;
wire v_4271;
wire v_4272;
wire v_4273;
wire v_4274;
wire v_4275;
wire v_4276;
wire v_4277;
wire v_4278;
wire v_4279;
wire v_4280;
wire v_4281;
wire v_4282;
wire v_4283;
wire v_4284;
wire v_4285;
wire v_4286;
wire v_4287;
wire v_4288;
wire v_4289;
wire v_4290;
wire v_4291;
wire v_4292;
wire v_4293;
wire v_4294;
wire v_4295;
wire v_4296;
wire v_4297;
wire v_4298;
wire v_4299;
wire v_4300;
wire v_4301;
wire v_4302;
wire v_4303;
wire v_4304;
wire v_4305;
wire v_4306;
wire v_4307;
wire v_4308;
wire v_4309;
wire v_4310;
wire v_4311;
wire v_4312;
wire v_4313;
wire v_4314;
wire v_4315;
wire v_4316;
wire v_4317;
wire v_4318;
wire v_4319;
wire v_4320;
wire v_4321;
wire v_4322;
wire v_4323;
wire v_4324;
wire v_4325;
wire v_4326;
wire v_4327;
wire v_4328;
wire v_4329;
wire v_4330;
wire v_4331;
wire v_4332;
wire v_4333;
wire v_4334;
wire v_4335;
wire v_4336;
wire v_4337;
wire v_4338;
wire v_4339;
wire v_4340;
wire v_4341;
wire v_4342;
wire v_4343;
wire v_4344;
wire v_4345;
wire v_4346;
wire v_4347;
wire v_4348;
wire v_4349;
wire v_4350;
wire v_4351;
wire v_4352;
wire v_4353;
wire v_4354;
wire v_4355;
wire v_4356;
wire v_4357;
wire v_4358;
wire v_4359;
wire v_4360;
wire v_4361;
wire v_4362;
wire v_4363;
wire v_4364;
wire v_4365;
wire v_4366;
wire v_4367;
wire v_4368;
wire v_4369;
wire v_4370;
wire v_4371;
wire v_4372;
wire v_4373;
wire v_4374;
wire v_4375;
wire v_4376;
wire v_4377;
wire v_4378;
wire v_4379;
wire v_4380;
wire v_4381;
wire v_4382;
wire v_4383;
wire v_4384;
wire v_4385;
wire v_4386;
wire v_4387;
wire v_4388;
wire v_4389;
wire v_4390;
wire v_4391;
wire v_4392;
wire v_4393;
wire v_4394;
wire v_4395;
wire v_4396;
wire v_4397;
wire v_4398;
wire v_4399;
wire v_4400;
wire v_4401;
wire v_4402;
wire v_4403;
wire v_4404;
wire v_4405;
wire v_4406;
wire v_4407;
wire v_4408;
wire v_4409;
wire v_4410;
wire v_4411;
wire v_4412;
wire v_4413;
wire v_4414;
wire v_4415;
wire v_4416;
wire v_4417;
wire v_4418;
wire v_4419;
wire v_4420;
wire v_4421;
wire v_4422;
wire v_4423;
wire v_4424;
wire v_4425;
wire v_4426;
wire v_4427;
wire v_4428;
wire v_4429;
wire v_4430;
wire v_4431;
wire v_4432;
wire v_4433;
wire v_4434;
wire v_4435;
wire v_4436;
wire v_4437;
wire v_4438;
wire v_4439;
wire v_4440;
wire v_4441;
wire v_4442;
wire v_4443;
wire v_4444;
wire v_4445;
wire v_4446;
wire v_4447;
wire v_4448;
wire v_4449;
wire v_4450;
wire v_4451;
wire v_4452;
wire v_4453;
wire v_4454;
wire v_4455;
wire v_4456;
wire v_4457;
wire v_4458;
wire v_4459;
wire v_4460;
wire v_4461;
wire v_4462;
wire v_4463;
wire v_4464;
wire v_4465;
wire v_4466;
wire v_4467;
wire v_4468;
wire v_4469;
wire v_4470;
wire v_4471;
wire v_4472;
wire v_4473;
wire v_4474;
wire v_4475;
wire v_4476;
wire v_4477;
wire v_4478;
wire v_4479;
wire v_4480;
wire v_4481;
wire v_4482;
wire v_4483;
wire v_4484;
wire v_4485;
wire v_4486;
wire v_4487;
wire v_4488;
wire v_4489;
wire v_4490;
wire v_4491;
wire v_4492;
wire v_4493;
wire v_4494;
wire v_4495;
wire v_4496;
wire v_4497;
wire v_4498;
wire v_4499;
wire v_4500;
wire v_4501;
wire v_4502;
wire v_4503;
wire v_4504;
wire v_4505;
wire v_4506;
wire v_4507;
wire v_4508;
wire v_4509;
wire v_4510;
wire v_4511;
wire v_4512;
wire v_4513;
wire v_4514;
wire v_4515;
wire v_4516;
wire v_4517;
wire v_4518;
wire v_4519;
wire v_4520;
wire v_4521;
wire v_4522;
wire v_4523;
wire v_4524;
wire v_4525;
wire v_4526;
wire v_4527;
wire v_4528;
wire v_4529;
wire v_4530;
wire v_4531;
wire v_4532;
wire v_4533;
wire v_4534;
wire v_4535;
wire v_4536;
wire v_4537;
wire v_4538;
wire v_4539;
wire v_4540;
wire v_4541;
wire v_4542;
wire v_4543;
wire v_4544;
wire v_4545;
wire v_4546;
wire v_4547;
wire v_4548;
wire v_4549;
wire v_4550;
wire v_4551;
wire v_4552;
wire v_4553;
wire v_4554;
wire v_4555;
wire x_1;
wire x_2;
wire x_3;
wire x_4;
wire x_5;
wire x_6;
wire x_7;
wire x_8;
wire x_9;
wire x_10;
wire x_11;
wire x_12;
wire x_13;
wire x_14;
wire x_15;
assign v_1088 = 1;
assign v_1217 = 1;
assign v_3140 = 1;
assign v_3524 = 1;
assign v_3908 = 1;
assign v_578 = ~v_514 & ~v_515;
assign v_580 = ~v_516 & v_578;
assign v_582 = ~v_517 & v_580;
assign v_584 = ~v_518 & v_582;
assign v_586 = ~v_519 & v_584;
assign v_588 = ~v_520 & v_586;
assign v_590 = ~v_521 & v_588;
assign v_592 = ~v_522 & v_590;
assign v_594 = ~v_523 & v_592;
assign v_596 = ~v_524 & v_594;
assign v_598 = ~v_525 & v_596;
assign v_600 = ~v_526 & v_598;
assign v_602 = ~v_527 & v_600;
assign v_604 = ~v_528 & v_602;
assign v_606 = ~v_529 & v_604;
assign v_608 = ~v_530 & v_606;
assign v_610 = ~v_531 & v_608;
assign v_612 = ~v_532 & v_610;
assign v_614 = ~v_533 & v_612;
assign v_616 = ~v_534 & v_614;
assign v_618 = ~v_535 & v_616;
assign v_620 = ~v_536 & v_618;
assign v_622 = ~v_537 & v_620;
assign v_624 = ~v_538 & v_622;
assign v_626 = ~v_539 & v_624;
assign v_628 = ~v_540 & v_626;
assign v_630 = ~v_541 & v_628;
assign v_632 = ~v_542 & v_630;
assign v_634 = ~v_543 & v_632;
assign v_636 = ~v_544 & v_634;
assign v_638 = ~v_545 & v_636;
assign v_640 = ~v_546 & v_638;
assign v_642 = ~v_547 & v_640;
assign v_644 = ~v_548 & v_642;
assign v_646 = ~v_549 & v_644;
assign v_648 = ~v_550 & v_646;
assign v_650 = ~v_551 & v_648;
assign v_652 = ~v_552 & v_650;
assign v_654 = ~v_553 & v_652;
assign v_656 = ~v_554 & v_654;
assign v_658 = ~v_555 & v_656;
assign v_660 = ~v_556 & v_658;
assign v_662 = ~v_557 & v_660;
assign v_664 = ~v_558 & v_662;
assign v_666 = ~v_559 & v_664;
assign v_668 = ~v_560 & v_666;
assign v_670 = ~v_561 & v_668;
assign v_672 = ~v_562 & v_670;
assign v_674 = ~v_563 & v_672;
assign v_676 = ~v_564 & v_674;
assign v_678 = ~v_565 & v_676;
assign v_680 = ~v_566 & v_678;
assign v_682 = ~v_567 & v_680;
assign v_684 = ~v_568 & v_682;
assign v_686 = ~v_569 & v_684;
assign v_688 = ~v_570 & v_686;
assign v_690 = ~v_571 & v_688;
assign v_692 = ~v_572 & v_690;
assign v_694 = ~v_573 & v_692;
assign v_696 = ~v_574 & v_694;
assign v_698 = ~v_575 & v_696;
assign v_700 = ~v_576 & v_698;
assign v_702 = ~v_577 & v_700;
assign v_705 = ~v_514 & v_450;
assign v_709 = ~v_579 & v_451;
assign v_710 = v_451 & v_706;
assign v_711 = ~v_579 & v_706;
assign v_715 = ~v_581 & v_452;
assign v_716 = v_452 & v_712;
assign v_717 = ~v_581 & v_712;
assign v_721 = ~v_583 & v_453;
assign v_722 = v_453 & v_718;
assign v_723 = ~v_583 & v_718;
assign v_727 = ~v_585 & v_454;
assign v_728 = v_454 & v_724;
assign v_729 = ~v_585 & v_724;
assign v_733 = ~v_587 & v_455;
assign v_734 = v_455 & v_730;
assign v_735 = ~v_587 & v_730;
assign v_739 = ~v_589 & v_456;
assign v_740 = v_456 & v_736;
assign v_741 = ~v_589 & v_736;
assign v_745 = ~v_591 & v_457;
assign v_746 = v_457 & v_742;
assign v_747 = ~v_591 & v_742;
assign v_751 = ~v_593 & v_458;
assign v_752 = v_458 & v_748;
assign v_753 = ~v_593 & v_748;
assign v_757 = ~v_595 & v_459;
assign v_758 = v_459 & v_754;
assign v_759 = ~v_595 & v_754;
assign v_763 = ~v_597 & v_460;
assign v_764 = v_460 & v_760;
assign v_765 = ~v_597 & v_760;
assign v_769 = ~v_599 & v_461;
assign v_770 = v_461 & v_766;
assign v_771 = ~v_599 & v_766;
assign v_775 = ~v_601 & v_462;
assign v_776 = v_462 & v_772;
assign v_777 = ~v_601 & v_772;
assign v_781 = ~v_603 & v_463;
assign v_782 = v_463 & v_778;
assign v_783 = ~v_603 & v_778;
assign v_787 = ~v_605 & v_464;
assign v_788 = v_464 & v_784;
assign v_789 = ~v_605 & v_784;
assign v_793 = ~v_607 & v_465;
assign v_794 = v_465 & v_790;
assign v_795 = ~v_607 & v_790;
assign v_799 = ~v_609 & v_466;
assign v_800 = v_466 & v_796;
assign v_801 = ~v_609 & v_796;
assign v_805 = ~v_611 & v_467;
assign v_806 = v_467 & v_802;
assign v_807 = ~v_611 & v_802;
assign v_811 = ~v_613 & v_468;
assign v_812 = v_468 & v_808;
assign v_813 = ~v_613 & v_808;
assign v_817 = ~v_615 & v_469;
assign v_818 = v_469 & v_814;
assign v_819 = ~v_615 & v_814;
assign v_823 = ~v_617 & v_470;
assign v_824 = v_470 & v_820;
assign v_825 = ~v_617 & v_820;
assign v_829 = ~v_619 & v_471;
assign v_830 = v_471 & v_826;
assign v_831 = ~v_619 & v_826;
assign v_835 = ~v_621 & v_472;
assign v_836 = v_472 & v_832;
assign v_837 = ~v_621 & v_832;
assign v_841 = ~v_623 & v_473;
assign v_842 = v_473 & v_838;
assign v_843 = ~v_623 & v_838;
assign v_847 = ~v_625 & v_474;
assign v_848 = v_474 & v_844;
assign v_849 = ~v_625 & v_844;
assign v_853 = ~v_627 & v_475;
assign v_854 = v_475 & v_850;
assign v_855 = ~v_627 & v_850;
assign v_859 = ~v_629 & v_476;
assign v_860 = v_476 & v_856;
assign v_861 = ~v_629 & v_856;
assign v_865 = ~v_631 & v_477;
assign v_866 = v_477 & v_862;
assign v_867 = ~v_631 & v_862;
assign v_871 = ~v_633 & v_478;
assign v_872 = v_478 & v_868;
assign v_873 = ~v_633 & v_868;
assign v_877 = ~v_635 & v_479;
assign v_878 = v_479 & v_874;
assign v_879 = ~v_635 & v_874;
assign v_883 = ~v_637 & v_480;
assign v_884 = v_480 & v_880;
assign v_885 = ~v_637 & v_880;
assign v_889 = ~v_639 & v_481;
assign v_890 = v_481 & v_886;
assign v_891 = ~v_639 & v_886;
assign v_895 = ~v_641 & v_482;
assign v_896 = v_482 & v_892;
assign v_897 = ~v_641 & v_892;
assign v_901 = ~v_643 & v_483;
assign v_902 = v_483 & v_898;
assign v_903 = ~v_643 & v_898;
assign v_907 = ~v_645 & v_484;
assign v_908 = v_484 & v_904;
assign v_909 = ~v_645 & v_904;
assign v_913 = ~v_647 & v_485;
assign v_914 = v_485 & v_910;
assign v_915 = ~v_647 & v_910;
assign v_919 = ~v_649 & v_486;
assign v_920 = v_486 & v_916;
assign v_921 = ~v_649 & v_916;
assign v_925 = ~v_651 & v_487;
assign v_926 = v_487 & v_922;
assign v_927 = ~v_651 & v_922;
assign v_931 = ~v_653 & v_488;
assign v_932 = v_488 & v_928;
assign v_933 = ~v_653 & v_928;
assign v_937 = ~v_655 & v_489;
assign v_938 = v_489 & v_934;
assign v_939 = ~v_655 & v_934;
assign v_943 = ~v_657 & v_490;
assign v_944 = v_490 & v_940;
assign v_945 = ~v_657 & v_940;
assign v_949 = ~v_659 & v_491;
assign v_950 = v_491 & v_946;
assign v_951 = ~v_659 & v_946;
assign v_955 = ~v_661 & v_492;
assign v_956 = v_492 & v_952;
assign v_957 = ~v_661 & v_952;
assign v_961 = ~v_663 & v_493;
assign v_962 = v_493 & v_958;
assign v_963 = ~v_663 & v_958;
assign v_967 = ~v_665 & v_494;
assign v_968 = v_494 & v_964;
assign v_969 = ~v_665 & v_964;
assign v_973 = ~v_667 & v_495;
assign v_974 = v_495 & v_970;
assign v_975 = ~v_667 & v_970;
assign v_979 = ~v_669 & v_496;
assign v_980 = v_496 & v_976;
assign v_981 = ~v_669 & v_976;
assign v_985 = ~v_671 & v_497;
assign v_986 = v_497 & v_982;
assign v_987 = ~v_671 & v_982;
assign v_991 = ~v_673 & v_498;
assign v_992 = v_498 & v_988;
assign v_993 = ~v_673 & v_988;
assign v_997 = ~v_675 & v_499;
assign v_998 = v_499 & v_994;
assign v_999 = ~v_675 & v_994;
assign v_1003 = ~v_677 & v_500;
assign v_1004 = v_500 & v_1000;
assign v_1005 = ~v_677 & v_1000;
assign v_1009 = ~v_679 & v_501;
assign v_1010 = v_501 & v_1006;
assign v_1011 = ~v_679 & v_1006;
assign v_1015 = ~v_681 & v_502;
assign v_1016 = v_502 & v_1012;
assign v_1017 = ~v_681 & v_1012;
assign v_1021 = ~v_683 & v_503;
assign v_1022 = v_503 & v_1018;
assign v_1023 = ~v_683 & v_1018;
assign v_1027 = ~v_685 & v_504;
assign v_1028 = v_504 & v_1024;
assign v_1029 = ~v_685 & v_1024;
assign v_1033 = ~v_687 & v_505;
assign v_1034 = v_505 & v_1030;
assign v_1035 = ~v_687 & v_1030;
assign v_1039 = ~v_689 & v_506;
assign v_1040 = v_506 & v_1036;
assign v_1041 = ~v_689 & v_1036;
assign v_1045 = ~v_691 & v_507;
assign v_1046 = v_507 & v_1042;
assign v_1047 = ~v_691 & v_1042;
assign v_1051 = ~v_693 & v_508;
assign v_1052 = v_508 & v_1048;
assign v_1053 = ~v_693 & v_1048;
assign v_1057 = ~v_695 & v_509;
assign v_1058 = v_509 & v_1054;
assign v_1059 = ~v_695 & v_1054;
assign v_1063 = ~v_697 & v_510;
assign v_1064 = v_510 & v_1060;
assign v_1065 = ~v_697 & v_1060;
assign v_1069 = ~v_699 & v_511;
assign v_1070 = v_511 & v_1066;
assign v_1071 = ~v_699 & v_1066;
assign v_1075 = ~v_701 & v_512;
assign v_1076 = v_512 & v_1072;
assign v_1077 = ~v_701 & v_1072;
assign v_1081 = ~v_703 & v_513;
assign v_1082 = v_513 & v_1078;
assign v_1083 = ~v_703 & v_1078;
assign v_1089 = ~v_514;
assign v_1090 = ~v_515 & v_1089;
assign v_1091 = v_1090;
assign v_1092 = ~v_516 & v_1091;
assign v_1093 = v_1092;
assign v_1094 = ~v_517 & v_1093;
assign v_1095 = v_1094;
assign v_1096 = ~v_518 & v_1095;
assign v_1097 = v_1096;
assign v_1098 = ~v_519 & v_1097;
assign v_1099 = v_1098;
assign v_1100 = ~v_520 & v_1099;
assign v_1101 = v_1100;
assign v_1102 = ~v_521 & v_1101;
assign v_1103 = v_1102;
assign v_1104 = ~v_522 & v_1103;
assign v_1105 = v_1104;
assign v_1106 = ~v_523 & v_1105;
assign v_1107 = v_1106;
assign v_1108 = ~v_524 & v_1107;
assign v_1109 = v_1108;
assign v_1110 = ~v_525 & v_1109;
assign v_1111 = v_1110;
assign v_1112 = ~v_526 & v_1111;
assign v_1113 = v_1112;
assign v_1114 = ~v_527 & v_1113;
assign v_1115 = v_1114;
assign v_1116 = ~v_528 & v_1115;
assign v_1117 = v_1116;
assign v_1118 = ~v_529 & v_1117;
assign v_1119 = v_1118;
assign v_1120 = ~v_530 & v_1119;
assign v_1121 = v_1120;
assign v_1122 = ~v_531 & v_1121;
assign v_1123 = v_1122;
assign v_1124 = ~v_532 & v_1123;
assign v_1125 = v_1124;
assign v_1126 = ~v_533 & v_1125;
assign v_1127 = v_1126;
assign v_1128 = ~v_534 & v_1127;
assign v_1129 = v_1128;
assign v_1130 = ~v_535 & v_1129;
assign v_1131 = v_1130;
assign v_1132 = ~v_536 & v_1131;
assign v_1133 = v_1132;
assign v_1134 = ~v_537 & v_1133;
assign v_1135 = v_1134;
assign v_1136 = ~v_538 & v_1135;
assign v_1137 = v_1136;
assign v_1138 = ~v_539 & v_1137;
assign v_1139 = v_1138;
assign v_1140 = ~v_540 & v_1139;
assign v_1141 = v_1140;
assign v_1142 = ~v_541 & v_1141;
assign v_1143 = v_1142;
assign v_1144 = ~v_542 & v_1143;
assign v_1145 = v_1144;
assign v_1146 = ~v_543 & v_1145;
assign v_1147 = v_1146;
assign v_1148 = ~v_544 & v_1147;
assign v_1149 = v_1148;
assign v_1150 = ~v_545 & v_1149;
assign v_1151 = v_1150;
assign v_1152 = ~v_546 & v_1151;
assign v_1153 = v_1152;
assign v_1154 = ~v_547 & v_1153;
assign v_1155 = v_1154;
assign v_1156 = ~v_548 & v_1155;
assign v_1157 = v_1156;
assign v_1158 = ~v_549 & v_1157;
assign v_1159 = v_1158;
assign v_1160 = ~v_550 & v_1159;
assign v_1161 = v_1160;
assign v_1162 = ~v_551 & v_1161;
assign v_1163 = v_1162;
assign v_1164 = ~v_552 & v_1163;
assign v_1165 = v_1164;
assign v_1166 = ~v_553 & v_1165;
assign v_1167 = v_1166;
assign v_1168 = ~v_554 & v_1167;
assign v_1169 = v_1168;
assign v_1170 = ~v_555 & v_1169;
assign v_1171 = v_1170;
assign v_1172 = ~v_556 & v_1171;
assign v_1173 = v_1172;
assign v_1174 = ~v_557 & v_1173;
assign v_1175 = v_1174;
assign v_1176 = ~v_558 & v_1175;
assign v_1177 = v_1176;
assign v_1178 = ~v_559 & v_1177;
assign v_1179 = v_1178;
assign v_1180 = ~v_560 & v_1179;
assign v_1181 = v_1180;
assign v_1182 = ~v_561 & v_1181;
assign v_1183 = v_1182;
assign v_1184 = ~v_562 & v_1183;
assign v_1185 = v_1184;
assign v_1186 = ~v_563 & v_1185;
assign v_1187 = v_1186;
assign v_1188 = ~v_564 & v_1187;
assign v_1189 = v_1188;
assign v_1190 = ~v_565 & v_1189;
assign v_1191 = v_1190;
assign v_1192 = ~v_566 & v_1191;
assign v_1193 = v_1192;
assign v_1194 = ~v_567 & v_1193;
assign v_1195 = v_1194;
assign v_1196 = ~v_568 & v_1195;
assign v_1197 = v_1196;
assign v_1198 = ~v_569 & v_1197;
assign v_1199 = v_1198;
assign v_1200 = ~v_570 & v_1199;
assign v_1201 = v_1200;
assign v_1202 = ~v_571 & v_1201;
assign v_1203 = v_1202;
assign v_1204 = ~v_572 & v_1203;
assign v_1205 = v_1204;
assign v_1206 = ~v_573 & v_1205;
assign v_1207 = v_1206;
assign v_1208 = ~v_574 & v_1207;
assign v_1209 = v_1208;
assign v_1210 = ~v_575 & v_1209;
assign v_1211 = v_1210;
assign v_1212 = ~v_576 & v_1211;
assign v_1213 = v_1212;
assign v_1214 = ~v_577 & v_1213;
assign v_1215 = v_1214;
assign v_1346 = v_4313 & v_4314 & v_4315;
assign v_1475 = v_4329 & v_4330 & v_4331;
assign v_1604 = v_4345 & v_4346 & v_4347;
assign v_1669 = v_4361 & v_4362 & v_4363;
assign v_1671 = v_450 & v_514;
assign v_1672 = v_1671;
assign v_1675 = v_451 & v_515;
assign v_1676 = v_515 & v_1672;
assign v_1677 = v_451 & v_1672;
assign v_1681 = v_452 & v_516;
assign v_1682 = v_516 & v_1678;
assign v_1683 = v_452 & v_1678;
assign v_1687 = v_453 & v_517;
assign v_1688 = v_517 & v_1684;
assign v_1689 = v_453 & v_1684;
assign v_1693 = v_454 & v_518;
assign v_1694 = v_518 & v_1690;
assign v_1695 = v_454 & v_1690;
assign v_1699 = v_455 & v_519;
assign v_1700 = v_519 & v_1696;
assign v_1701 = v_455 & v_1696;
assign v_1705 = v_456 & v_520;
assign v_1706 = v_520 & v_1702;
assign v_1707 = v_456 & v_1702;
assign v_1711 = v_457 & v_521;
assign v_1712 = v_521 & v_1708;
assign v_1713 = v_457 & v_1708;
assign v_1717 = v_458 & v_522;
assign v_1718 = v_522 & v_1714;
assign v_1719 = v_458 & v_1714;
assign v_1723 = v_459 & v_523;
assign v_1724 = v_523 & v_1720;
assign v_1725 = v_459 & v_1720;
assign v_1729 = v_460 & v_524;
assign v_1730 = v_524 & v_1726;
assign v_1731 = v_460 & v_1726;
assign v_1735 = v_461 & v_525;
assign v_1736 = v_525 & v_1732;
assign v_1737 = v_461 & v_1732;
assign v_1741 = v_462 & v_526;
assign v_1742 = v_526 & v_1738;
assign v_1743 = v_462 & v_1738;
assign v_1747 = v_463 & v_527;
assign v_1748 = v_527 & v_1744;
assign v_1749 = v_463 & v_1744;
assign v_1753 = v_464 & v_528;
assign v_1754 = v_528 & v_1750;
assign v_1755 = v_464 & v_1750;
assign v_1759 = v_465 & v_529;
assign v_1760 = v_529 & v_1756;
assign v_1761 = v_465 & v_1756;
assign v_1765 = v_466 & v_530;
assign v_1766 = v_530 & v_1762;
assign v_1767 = v_466 & v_1762;
assign v_1771 = v_467 & v_531;
assign v_1772 = v_531 & v_1768;
assign v_1773 = v_467 & v_1768;
assign v_1777 = v_468 & v_532;
assign v_1778 = v_532 & v_1774;
assign v_1779 = v_468 & v_1774;
assign v_1783 = v_469 & v_533;
assign v_1784 = v_533 & v_1780;
assign v_1785 = v_469 & v_1780;
assign v_1789 = v_470 & v_534;
assign v_1790 = v_534 & v_1786;
assign v_1791 = v_470 & v_1786;
assign v_1795 = v_471 & v_535;
assign v_1796 = v_535 & v_1792;
assign v_1797 = v_471 & v_1792;
assign v_1801 = v_472 & v_536;
assign v_1802 = v_536 & v_1798;
assign v_1803 = v_472 & v_1798;
assign v_1807 = v_473 & v_537;
assign v_1808 = v_537 & v_1804;
assign v_1809 = v_473 & v_1804;
assign v_1813 = v_474 & v_538;
assign v_1814 = v_538 & v_1810;
assign v_1815 = v_474 & v_1810;
assign v_1819 = v_475 & v_539;
assign v_1820 = v_539 & v_1816;
assign v_1821 = v_475 & v_1816;
assign v_1825 = v_476 & v_540;
assign v_1826 = v_540 & v_1822;
assign v_1827 = v_476 & v_1822;
assign v_1831 = v_477 & v_541;
assign v_1832 = v_541 & v_1828;
assign v_1833 = v_477 & v_1828;
assign v_1837 = v_478 & v_542;
assign v_1838 = v_542 & v_1834;
assign v_1839 = v_478 & v_1834;
assign v_1843 = v_479 & v_543;
assign v_1844 = v_543 & v_1840;
assign v_1845 = v_479 & v_1840;
assign v_1849 = v_480 & v_544;
assign v_1850 = v_544 & v_1846;
assign v_1851 = v_480 & v_1846;
assign v_1855 = v_481 & v_545;
assign v_1856 = v_545 & v_1852;
assign v_1857 = v_481 & v_1852;
assign v_1861 = v_482 & v_546;
assign v_1862 = v_546 & v_1858;
assign v_1863 = v_482 & v_1858;
assign v_1867 = v_483 & v_547;
assign v_1868 = v_547 & v_1864;
assign v_1869 = v_483 & v_1864;
assign v_1873 = v_484 & v_548;
assign v_1874 = v_548 & v_1870;
assign v_1875 = v_484 & v_1870;
assign v_1879 = v_485 & v_549;
assign v_1880 = v_549 & v_1876;
assign v_1881 = v_485 & v_1876;
assign v_1885 = v_486 & v_550;
assign v_1886 = v_550 & v_1882;
assign v_1887 = v_486 & v_1882;
assign v_1891 = v_487 & v_551;
assign v_1892 = v_551 & v_1888;
assign v_1893 = v_487 & v_1888;
assign v_1897 = v_488 & v_552;
assign v_1898 = v_552 & v_1894;
assign v_1899 = v_488 & v_1894;
assign v_1903 = v_489 & v_553;
assign v_1904 = v_553 & v_1900;
assign v_1905 = v_489 & v_1900;
assign v_1909 = v_490 & v_554;
assign v_1910 = v_554 & v_1906;
assign v_1911 = v_490 & v_1906;
assign v_1915 = v_491 & v_555;
assign v_1916 = v_555 & v_1912;
assign v_1917 = v_491 & v_1912;
assign v_1921 = v_492 & v_556;
assign v_1922 = v_556 & v_1918;
assign v_1923 = v_492 & v_1918;
assign v_1927 = v_493 & v_557;
assign v_1928 = v_557 & v_1924;
assign v_1929 = v_493 & v_1924;
assign v_1933 = v_494 & v_558;
assign v_1934 = v_558 & v_1930;
assign v_1935 = v_494 & v_1930;
assign v_1939 = v_495 & v_559;
assign v_1940 = v_559 & v_1936;
assign v_1941 = v_495 & v_1936;
assign v_1945 = v_496 & v_560;
assign v_1946 = v_560 & v_1942;
assign v_1947 = v_496 & v_1942;
assign v_1951 = v_497 & v_561;
assign v_1952 = v_561 & v_1948;
assign v_1953 = v_497 & v_1948;
assign v_1957 = v_498 & v_562;
assign v_1958 = v_562 & v_1954;
assign v_1959 = v_498 & v_1954;
assign v_1963 = v_499 & v_563;
assign v_1964 = v_563 & v_1960;
assign v_1965 = v_499 & v_1960;
assign v_1969 = v_500 & v_564;
assign v_1970 = v_564 & v_1966;
assign v_1971 = v_500 & v_1966;
assign v_1975 = v_501 & v_565;
assign v_1976 = v_565 & v_1972;
assign v_1977 = v_501 & v_1972;
assign v_1981 = v_502 & v_566;
assign v_1982 = v_566 & v_1978;
assign v_1983 = v_502 & v_1978;
assign v_1987 = v_503 & v_567;
assign v_1988 = v_567 & v_1984;
assign v_1989 = v_503 & v_1984;
assign v_1993 = v_504 & v_568;
assign v_1994 = v_568 & v_1990;
assign v_1995 = v_504 & v_1990;
assign v_1999 = v_505 & v_569;
assign v_2000 = v_569 & v_1996;
assign v_2001 = v_505 & v_1996;
assign v_2005 = v_506 & v_570;
assign v_2006 = v_570 & v_2002;
assign v_2007 = v_506 & v_2002;
assign v_2011 = v_507 & v_571;
assign v_2012 = v_571 & v_2008;
assign v_2013 = v_507 & v_2008;
assign v_2017 = v_508 & v_572;
assign v_2018 = v_572 & v_2014;
assign v_2019 = v_508 & v_2014;
assign v_2023 = v_509 & v_573;
assign v_2024 = v_573 & v_2020;
assign v_2025 = v_509 & v_2020;
assign v_2029 = v_510 & v_574;
assign v_2030 = v_574 & v_2026;
assign v_2031 = v_510 & v_2026;
assign v_2035 = v_511 & v_575;
assign v_2036 = v_575 & v_2032;
assign v_2037 = v_511 & v_2032;
assign v_2041 = v_512 & v_576;
assign v_2042 = v_576 & v_2038;
assign v_2043 = v_512 & v_2038;
assign v_2047 = v_513 & v_577;
assign v_2048 = v_577 & v_2044;
assign v_2049 = v_513 & v_2044;
assign v_2115 = v_4377 & v_4378 & v_4379;
assign v_2180 = v_4393 & v_4394 & v_4395;
assign v_2182 = v_385 & v_450;
assign v_2183 = v_2182;
assign v_2186 = v_386 & v_451;
assign v_2187 = v_451 & v_2183;
assign v_2188 = v_386 & v_2183;
assign v_2192 = v_387 & v_452;
assign v_2193 = v_452 & v_2189;
assign v_2194 = v_387 & v_2189;
assign v_2198 = v_388 & v_453;
assign v_2199 = v_453 & v_2195;
assign v_2200 = v_388 & v_2195;
assign v_2204 = v_389 & v_454;
assign v_2205 = v_454 & v_2201;
assign v_2206 = v_389 & v_2201;
assign v_2210 = v_390 & v_455;
assign v_2211 = v_455 & v_2207;
assign v_2212 = v_390 & v_2207;
assign v_2216 = v_391 & v_456;
assign v_2217 = v_456 & v_2213;
assign v_2218 = v_391 & v_2213;
assign v_2222 = v_392 & v_457;
assign v_2223 = v_457 & v_2219;
assign v_2224 = v_392 & v_2219;
assign v_2228 = v_393 & v_458;
assign v_2229 = v_458 & v_2225;
assign v_2230 = v_393 & v_2225;
assign v_2234 = v_394 & v_459;
assign v_2235 = v_459 & v_2231;
assign v_2236 = v_394 & v_2231;
assign v_2240 = v_395 & v_460;
assign v_2241 = v_460 & v_2237;
assign v_2242 = v_395 & v_2237;
assign v_2246 = v_396 & v_461;
assign v_2247 = v_461 & v_2243;
assign v_2248 = v_396 & v_2243;
assign v_2252 = v_397 & v_462;
assign v_2253 = v_462 & v_2249;
assign v_2254 = v_397 & v_2249;
assign v_2258 = v_398 & v_463;
assign v_2259 = v_463 & v_2255;
assign v_2260 = v_398 & v_2255;
assign v_2264 = v_399 & v_464;
assign v_2265 = v_464 & v_2261;
assign v_2266 = v_399 & v_2261;
assign v_2270 = v_400 & v_465;
assign v_2271 = v_465 & v_2267;
assign v_2272 = v_400 & v_2267;
assign v_2276 = v_401 & v_466;
assign v_2277 = v_466 & v_2273;
assign v_2278 = v_401 & v_2273;
assign v_2282 = v_402 & v_467;
assign v_2283 = v_467 & v_2279;
assign v_2284 = v_402 & v_2279;
assign v_2288 = v_403 & v_468;
assign v_2289 = v_468 & v_2285;
assign v_2290 = v_403 & v_2285;
assign v_2294 = v_404 & v_469;
assign v_2295 = v_469 & v_2291;
assign v_2296 = v_404 & v_2291;
assign v_2300 = v_405 & v_470;
assign v_2301 = v_470 & v_2297;
assign v_2302 = v_405 & v_2297;
assign v_2306 = v_406 & v_471;
assign v_2307 = v_471 & v_2303;
assign v_2308 = v_406 & v_2303;
assign v_2312 = v_407 & v_472;
assign v_2313 = v_472 & v_2309;
assign v_2314 = v_407 & v_2309;
assign v_2318 = v_408 & v_473;
assign v_2319 = v_473 & v_2315;
assign v_2320 = v_408 & v_2315;
assign v_2324 = v_409 & v_474;
assign v_2325 = v_474 & v_2321;
assign v_2326 = v_409 & v_2321;
assign v_2330 = v_410 & v_475;
assign v_2331 = v_475 & v_2327;
assign v_2332 = v_410 & v_2327;
assign v_2336 = v_411 & v_476;
assign v_2337 = v_476 & v_2333;
assign v_2338 = v_411 & v_2333;
assign v_2342 = v_412 & v_477;
assign v_2343 = v_477 & v_2339;
assign v_2344 = v_412 & v_2339;
assign v_2348 = v_413 & v_478;
assign v_2349 = v_478 & v_2345;
assign v_2350 = v_413 & v_2345;
assign v_2354 = v_414 & v_479;
assign v_2355 = v_479 & v_2351;
assign v_2356 = v_414 & v_2351;
assign v_2360 = v_415 & v_480;
assign v_2361 = v_480 & v_2357;
assign v_2362 = v_415 & v_2357;
assign v_2366 = v_416 & v_481;
assign v_2367 = v_481 & v_2363;
assign v_2368 = v_416 & v_2363;
assign v_2372 = v_417 & v_482;
assign v_2373 = v_482 & v_2369;
assign v_2374 = v_417 & v_2369;
assign v_2378 = v_418 & v_483;
assign v_2379 = v_483 & v_2375;
assign v_2380 = v_418 & v_2375;
assign v_2384 = v_419 & v_484;
assign v_2385 = v_484 & v_2381;
assign v_2386 = v_419 & v_2381;
assign v_2390 = v_420 & v_485;
assign v_2391 = v_485 & v_2387;
assign v_2392 = v_420 & v_2387;
assign v_2396 = v_421 & v_486;
assign v_2397 = v_486 & v_2393;
assign v_2398 = v_421 & v_2393;
assign v_2402 = v_422 & v_487;
assign v_2403 = v_487 & v_2399;
assign v_2404 = v_422 & v_2399;
assign v_2408 = v_423 & v_488;
assign v_2409 = v_488 & v_2405;
assign v_2410 = v_423 & v_2405;
assign v_2414 = v_424 & v_489;
assign v_2415 = v_489 & v_2411;
assign v_2416 = v_424 & v_2411;
assign v_2420 = v_425 & v_490;
assign v_2421 = v_490 & v_2417;
assign v_2422 = v_425 & v_2417;
assign v_2426 = v_426 & v_491;
assign v_2427 = v_491 & v_2423;
assign v_2428 = v_426 & v_2423;
assign v_2432 = v_427 & v_492;
assign v_2433 = v_492 & v_2429;
assign v_2434 = v_427 & v_2429;
assign v_2438 = v_428 & v_493;
assign v_2439 = v_493 & v_2435;
assign v_2440 = v_428 & v_2435;
assign v_2444 = v_429 & v_494;
assign v_2445 = v_494 & v_2441;
assign v_2446 = v_429 & v_2441;
assign v_2450 = v_430 & v_495;
assign v_2451 = v_495 & v_2447;
assign v_2452 = v_430 & v_2447;
assign v_2456 = v_431 & v_496;
assign v_2457 = v_496 & v_2453;
assign v_2458 = v_431 & v_2453;
assign v_2462 = v_432 & v_497;
assign v_2463 = v_497 & v_2459;
assign v_2464 = v_432 & v_2459;
assign v_2468 = v_433 & v_498;
assign v_2469 = v_498 & v_2465;
assign v_2470 = v_433 & v_2465;
assign v_2474 = v_434 & v_499;
assign v_2475 = v_499 & v_2471;
assign v_2476 = v_434 & v_2471;
assign v_2480 = v_435 & v_500;
assign v_2481 = v_500 & v_2477;
assign v_2482 = v_435 & v_2477;
assign v_2486 = v_436 & v_501;
assign v_2487 = v_501 & v_2483;
assign v_2488 = v_436 & v_2483;
assign v_2492 = v_437 & v_502;
assign v_2493 = v_502 & v_2489;
assign v_2494 = v_437 & v_2489;
assign v_2498 = v_438 & v_503;
assign v_2499 = v_503 & v_2495;
assign v_2500 = v_438 & v_2495;
assign v_2504 = v_439 & v_504;
assign v_2505 = v_504 & v_2501;
assign v_2506 = v_439 & v_2501;
assign v_2510 = v_440 & v_505;
assign v_2511 = v_505 & v_2507;
assign v_2512 = v_440 & v_2507;
assign v_2516 = v_441 & v_506;
assign v_2517 = v_506 & v_2513;
assign v_2518 = v_441 & v_2513;
assign v_2522 = v_442 & v_507;
assign v_2523 = v_507 & v_2519;
assign v_2524 = v_442 & v_2519;
assign v_2528 = v_443 & v_508;
assign v_2529 = v_508 & v_2525;
assign v_2530 = v_443 & v_2525;
assign v_2534 = v_444 & v_509;
assign v_2535 = v_509 & v_2531;
assign v_2536 = v_444 & v_2531;
assign v_2540 = v_445 & v_510;
assign v_2541 = v_510 & v_2537;
assign v_2542 = v_445 & v_2537;
assign v_2546 = v_446 & v_511;
assign v_2547 = v_511 & v_2543;
assign v_2548 = v_446 & v_2543;
assign v_2552 = v_447 & v_512;
assign v_2553 = v_512 & v_2549;
assign v_2554 = v_447 & v_2549;
assign v_2558 = v_448 & v_513;
assign v_2559 = v_513 & v_2555;
assign v_2560 = v_448 & v_2555;
assign v_2626 = v_4409 & v_4410 & v_4411;
assign v_2691 = v_4425 & v_4426 & v_4427;
assign v_2756 = v_4441 & v_4442 & v_4443;
assign v_2885 = ~v_2757 & v_2821;
assign v_2887 = ~v_2758 & v_2822;
assign v_2888 = v_2822 & v_2886;
assign v_2889 = ~v_2758 & v_2886;
assign v_2891 = ~v_2759 & v_2823;
assign v_2892 = v_2823 & v_2890;
assign v_2893 = ~v_2759 & v_2890;
assign v_2895 = ~v_2760 & v_2824;
assign v_2896 = v_2824 & v_2894;
assign v_2897 = ~v_2760 & v_2894;
assign v_2899 = ~v_2761 & v_2825;
assign v_2900 = v_2825 & v_2898;
assign v_2901 = ~v_2761 & v_2898;
assign v_2903 = ~v_2762 & v_2826;
assign v_2904 = v_2826 & v_2902;
assign v_2905 = ~v_2762 & v_2902;
assign v_2907 = ~v_2763 & v_2827;
assign v_2908 = v_2827 & v_2906;
assign v_2909 = ~v_2763 & v_2906;
assign v_2911 = ~v_2764 & v_2828;
assign v_2912 = v_2828 & v_2910;
assign v_2913 = ~v_2764 & v_2910;
assign v_2915 = ~v_2765 & v_2829;
assign v_2916 = v_2829 & v_2914;
assign v_2917 = ~v_2765 & v_2914;
assign v_2919 = ~v_2766 & v_2830;
assign v_2920 = v_2830 & v_2918;
assign v_2921 = ~v_2766 & v_2918;
assign v_2923 = ~v_2767 & v_2831;
assign v_2924 = v_2831 & v_2922;
assign v_2925 = ~v_2767 & v_2922;
assign v_2927 = ~v_2768 & v_2832;
assign v_2928 = v_2832 & v_2926;
assign v_2929 = ~v_2768 & v_2926;
assign v_2931 = ~v_2769 & v_2833;
assign v_2932 = v_2833 & v_2930;
assign v_2933 = ~v_2769 & v_2930;
assign v_2935 = ~v_2770 & v_2834;
assign v_2936 = v_2834 & v_2934;
assign v_2937 = ~v_2770 & v_2934;
assign v_2939 = ~v_2771 & v_2835;
assign v_2940 = v_2835 & v_2938;
assign v_2941 = ~v_2771 & v_2938;
assign v_2943 = ~v_2772 & v_2836;
assign v_2944 = v_2836 & v_2942;
assign v_2945 = ~v_2772 & v_2942;
assign v_2947 = ~v_2773 & v_2837;
assign v_2948 = v_2837 & v_2946;
assign v_2949 = ~v_2773 & v_2946;
assign v_2951 = ~v_2774 & v_2838;
assign v_2952 = v_2838 & v_2950;
assign v_2953 = ~v_2774 & v_2950;
assign v_2955 = ~v_2775 & v_2839;
assign v_2956 = v_2839 & v_2954;
assign v_2957 = ~v_2775 & v_2954;
assign v_2959 = ~v_2776 & v_2840;
assign v_2960 = v_2840 & v_2958;
assign v_2961 = ~v_2776 & v_2958;
assign v_2963 = ~v_2777 & v_2841;
assign v_2964 = v_2841 & v_2962;
assign v_2965 = ~v_2777 & v_2962;
assign v_2967 = ~v_2778 & v_2842;
assign v_2968 = v_2842 & v_2966;
assign v_2969 = ~v_2778 & v_2966;
assign v_2971 = ~v_2779 & v_2843;
assign v_2972 = v_2843 & v_2970;
assign v_2973 = ~v_2779 & v_2970;
assign v_2975 = ~v_2780 & v_2844;
assign v_2976 = v_2844 & v_2974;
assign v_2977 = ~v_2780 & v_2974;
assign v_2979 = ~v_2781 & v_2845;
assign v_2980 = v_2845 & v_2978;
assign v_2981 = ~v_2781 & v_2978;
assign v_2983 = ~v_2782 & v_2846;
assign v_2984 = v_2846 & v_2982;
assign v_2985 = ~v_2782 & v_2982;
assign v_2987 = ~v_2783 & v_2847;
assign v_2988 = v_2847 & v_2986;
assign v_2989 = ~v_2783 & v_2986;
assign v_2991 = ~v_2784 & v_2848;
assign v_2992 = v_2848 & v_2990;
assign v_2993 = ~v_2784 & v_2990;
assign v_2995 = ~v_2785 & v_2849;
assign v_2996 = v_2849 & v_2994;
assign v_2997 = ~v_2785 & v_2994;
assign v_2999 = ~v_2786 & v_2850;
assign v_3000 = v_2850 & v_2998;
assign v_3001 = ~v_2786 & v_2998;
assign v_3003 = ~v_2787 & v_2851;
assign v_3004 = v_2851 & v_3002;
assign v_3005 = ~v_2787 & v_3002;
assign v_3007 = ~v_2788 & v_2852;
assign v_3008 = v_2852 & v_3006;
assign v_3009 = ~v_2788 & v_3006;
assign v_3011 = ~v_2789 & v_2853;
assign v_3012 = v_2853 & v_3010;
assign v_3013 = ~v_2789 & v_3010;
assign v_3015 = ~v_2790 & v_2854;
assign v_3016 = v_2854 & v_3014;
assign v_3017 = ~v_2790 & v_3014;
assign v_3019 = ~v_2791 & v_2855;
assign v_3020 = v_2855 & v_3018;
assign v_3021 = ~v_2791 & v_3018;
assign v_3023 = ~v_2792 & v_2856;
assign v_3024 = v_2856 & v_3022;
assign v_3025 = ~v_2792 & v_3022;
assign v_3027 = ~v_2793 & v_2857;
assign v_3028 = v_2857 & v_3026;
assign v_3029 = ~v_2793 & v_3026;
assign v_3031 = ~v_2794 & v_2858;
assign v_3032 = v_2858 & v_3030;
assign v_3033 = ~v_2794 & v_3030;
assign v_3035 = ~v_2795 & v_2859;
assign v_3036 = v_2859 & v_3034;
assign v_3037 = ~v_2795 & v_3034;
assign v_3039 = ~v_2796 & v_2860;
assign v_3040 = v_2860 & v_3038;
assign v_3041 = ~v_2796 & v_3038;
assign v_3043 = ~v_2797 & v_2861;
assign v_3044 = v_2861 & v_3042;
assign v_3045 = ~v_2797 & v_3042;
assign v_3047 = ~v_2798 & v_2862;
assign v_3048 = v_2862 & v_3046;
assign v_3049 = ~v_2798 & v_3046;
assign v_3051 = ~v_2799 & v_2863;
assign v_3052 = v_2863 & v_3050;
assign v_3053 = ~v_2799 & v_3050;
assign v_3055 = ~v_2800 & v_2864;
assign v_3056 = v_2864 & v_3054;
assign v_3057 = ~v_2800 & v_3054;
assign v_3059 = ~v_2801 & v_2865;
assign v_3060 = v_2865 & v_3058;
assign v_3061 = ~v_2801 & v_3058;
assign v_3063 = ~v_2802 & v_2866;
assign v_3064 = v_2866 & v_3062;
assign v_3065 = ~v_2802 & v_3062;
assign v_3067 = ~v_2803 & v_2867;
assign v_3068 = v_2867 & v_3066;
assign v_3069 = ~v_2803 & v_3066;
assign v_3071 = ~v_2804 & v_2868;
assign v_3072 = v_2868 & v_3070;
assign v_3073 = ~v_2804 & v_3070;
assign v_3075 = ~v_2805 & v_2869;
assign v_3076 = v_2869 & v_3074;
assign v_3077 = ~v_2805 & v_3074;
assign v_3079 = ~v_2806 & v_2870;
assign v_3080 = v_2870 & v_3078;
assign v_3081 = ~v_2806 & v_3078;
assign v_3083 = ~v_2807 & v_2871;
assign v_3084 = v_2871 & v_3082;
assign v_3085 = ~v_2807 & v_3082;
assign v_3087 = ~v_2808 & v_2872;
assign v_3088 = v_2872 & v_3086;
assign v_3089 = ~v_2808 & v_3086;
assign v_3091 = ~v_2809 & v_2873;
assign v_3092 = v_2873 & v_3090;
assign v_3093 = ~v_2809 & v_3090;
assign v_3095 = ~v_2810 & v_2874;
assign v_3096 = v_2874 & v_3094;
assign v_3097 = ~v_2810 & v_3094;
assign v_3099 = ~v_2811 & v_2875;
assign v_3100 = v_2875 & v_3098;
assign v_3101 = ~v_2811 & v_3098;
assign v_3103 = ~v_2812 & v_2876;
assign v_3104 = v_2876 & v_3102;
assign v_3105 = ~v_2812 & v_3102;
assign v_3107 = ~v_2813 & v_2877;
assign v_3108 = v_2877 & v_3106;
assign v_3109 = ~v_2813 & v_3106;
assign v_3111 = ~v_2814 & v_2878;
assign v_3112 = v_2878 & v_3110;
assign v_3113 = ~v_2814 & v_3110;
assign v_3115 = ~v_2815 & v_2879;
assign v_3116 = v_2879 & v_3114;
assign v_3117 = ~v_2815 & v_3114;
assign v_3119 = ~v_2816 & v_2880;
assign v_3120 = v_2880 & v_3118;
assign v_3121 = ~v_2816 & v_3118;
assign v_3123 = ~v_2817 & v_2881;
assign v_3124 = v_2881 & v_3122;
assign v_3125 = ~v_2817 & v_3122;
assign v_3127 = ~v_2818 & v_2882;
assign v_3128 = v_2882 & v_3126;
assign v_3129 = ~v_2818 & v_3126;
assign v_3131 = ~v_2819 & v_2883;
assign v_3132 = v_2883 & v_3130;
assign v_3133 = ~v_2819 & v_3130;
assign v_3135 = ~v_2820 & v_2884;
assign v_3136 = v_2884 & v_3134;
assign v_3137 = ~v_2820 & v_3134;
assign v_3269 = ~v_3141 & v_3205;
assign v_3271 = ~v_3142 & v_3206;
assign v_3272 = v_3206 & v_3270;
assign v_3273 = ~v_3142 & v_3270;
assign v_3275 = ~v_3143 & v_3207;
assign v_3276 = v_3207 & v_3274;
assign v_3277 = ~v_3143 & v_3274;
assign v_3279 = ~v_3144 & v_3208;
assign v_3280 = v_3208 & v_3278;
assign v_3281 = ~v_3144 & v_3278;
assign v_3283 = ~v_3145 & v_3209;
assign v_3284 = v_3209 & v_3282;
assign v_3285 = ~v_3145 & v_3282;
assign v_3287 = ~v_3146 & v_3210;
assign v_3288 = v_3210 & v_3286;
assign v_3289 = ~v_3146 & v_3286;
assign v_3291 = ~v_3147 & v_3211;
assign v_3292 = v_3211 & v_3290;
assign v_3293 = ~v_3147 & v_3290;
assign v_3295 = ~v_3148 & v_3212;
assign v_3296 = v_3212 & v_3294;
assign v_3297 = ~v_3148 & v_3294;
assign v_3299 = ~v_3149 & v_3213;
assign v_3300 = v_3213 & v_3298;
assign v_3301 = ~v_3149 & v_3298;
assign v_3303 = ~v_3150 & v_3214;
assign v_3304 = v_3214 & v_3302;
assign v_3305 = ~v_3150 & v_3302;
assign v_3307 = ~v_3151 & v_3215;
assign v_3308 = v_3215 & v_3306;
assign v_3309 = ~v_3151 & v_3306;
assign v_3311 = ~v_3152 & v_3216;
assign v_3312 = v_3216 & v_3310;
assign v_3313 = ~v_3152 & v_3310;
assign v_3315 = ~v_3153 & v_3217;
assign v_3316 = v_3217 & v_3314;
assign v_3317 = ~v_3153 & v_3314;
assign v_3319 = ~v_3154 & v_3218;
assign v_3320 = v_3218 & v_3318;
assign v_3321 = ~v_3154 & v_3318;
assign v_3323 = ~v_3155 & v_3219;
assign v_3324 = v_3219 & v_3322;
assign v_3325 = ~v_3155 & v_3322;
assign v_3327 = ~v_3156 & v_3220;
assign v_3328 = v_3220 & v_3326;
assign v_3329 = ~v_3156 & v_3326;
assign v_3331 = ~v_3157 & v_3221;
assign v_3332 = v_3221 & v_3330;
assign v_3333 = ~v_3157 & v_3330;
assign v_3335 = ~v_3158 & v_3222;
assign v_3336 = v_3222 & v_3334;
assign v_3337 = ~v_3158 & v_3334;
assign v_3339 = ~v_3159 & v_3223;
assign v_3340 = v_3223 & v_3338;
assign v_3341 = ~v_3159 & v_3338;
assign v_3343 = ~v_3160 & v_3224;
assign v_3344 = v_3224 & v_3342;
assign v_3345 = ~v_3160 & v_3342;
assign v_3347 = ~v_3161 & v_3225;
assign v_3348 = v_3225 & v_3346;
assign v_3349 = ~v_3161 & v_3346;
assign v_3351 = ~v_3162 & v_3226;
assign v_3352 = v_3226 & v_3350;
assign v_3353 = ~v_3162 & v_3350;
assign v_3355 = ~v_3163 & v_3227;
assign v_3356 = v_3227 & v_3354;
assign v_3357 = ~v_3163 & v_3354;
assign v_3359 = ~v_3164 & v_3228;
assign v_3360 = v_3228 & v_3358;
assign v_3361 = ~v_3164 & v_3358;
assign v_3363 = ~v_3165 & v_3229;
assign v_3364 = v_3229 & v_3362;
assign v_3365 = ~v_3165 & v_3362;
assign v_3367 = ~v_3166 & v_3230;
assign v_3368 = v_3230 & v_3366;
assign v_3369 = ~v_3166 & v_3366;
assign v_3371 = ~v_3167 & v_3231;
assign v_3372 = v_3231 & v_3370;
assign v_3373 = ~v_3167 & v_3370;
assign v_3375 = ~v_3168 & v_3232;
assign v_3376 = v_3232 & v_3374;
assign v_3377 = ~v_3168 & v_3374;
assign v_3379 = ~v_3169 & v_3233;
assign v_3380 = v_3233 & v_3378;
assign v_3381 = ~v_3169 & v_3378;
assign v_3383 = ~v_3170 & v_3234;
assign v_3384 = v_3234 & v_3382;
assign v_3385 = ~v_3170 & v_3382;
assign v_3387 = ~v_3171 & v_3235;
assign v_3388 = v_3235 & v_3386;
assign v_3389 = ~v_3171 & v_3386;
assign v_3391 = ~v_3172 & v_3236;
assign v_3392 = v_3236 & v_3390;
assign v_3393 = ~v_3172 & v_3390;
assign v_3395 = ~v_3173 & v_3237;
assign v_3396 = v_3237 & v_3394;
assign v_3397 = ~v_3173 & v_3394;
assign v_3399 = ~v_3174 & v_3238;
assign v_3400 = v_3238 & v_3398;
assign v_3401 = ~v_3174 & v_3398;
assign v_3403 = ~v_3175 & v_3239;
assign v_3404 = v_3239 & v_3402;
assign v_3405 = ~v_3175 & v_3402;
assign v_3407 = ~v_3176 & v_3240;
assign v_3408 = v_3240 & v_3406;
assign v_3409 = ~v_3176 & v_3406;
assign v_3411 = ~v_3177 & v_3241;
assign v_3412 = v_3241 & v_3410;
assign v_3413 = ~v_3177 & v_3410;
assign v_3415 = ~v_3178 & v_3242;
assign v_3416 = v_3242 & v_3414;
assign v_3417 = ~v_3178 & v_3414;
assign v_3419 = ~v_3179 & v_3243;
assign v_3420 = v_3243 & v_3418;
assign v_3421 = ~v_3179 & v_3418;
assign v_3423 = ~v_3180 & v_3244;
assign v_3424 = v_3244 & v_3422;
assign v_3425 = ~v_3180 & v_3422;
assign v_3427 = ~v_3181 & v_3245;
assign v_3428 = v_3245 & v_3426;
assign v_3429 = ~v_3181 & v_3426;
assign v_3431 = ~v_3182 & v_3246;
assign v_3432 = v_3246 & v_3430;
assign v_3433 = ~v_3182 & v_3430;
assign v_3435 = ~v_3183 & v_3247;
assign v_3436 = v_3247 & v_3434;
assign v_3437 = ~v_3183 & v_3434;
assign v_3439 = ~v_3184 & v_3248;
assign v_3440 = v_3248 & v_3438;
assign v_3441 = ~v_3184 & v_3438;
assign v_3443 = ~v_3185 & v_3249;
assign v_3444 = v_3249 & v_3442;
assign v_3445 = ~v_3185 & v_3442;
assign v_3447 = ~v_3186 & v_3250;
assign v_3448 = v_3250 & v_3446;
assign v_3449 = ~v_3186 & v_3446;
assign v_3451 = ~v_3187 & v_3251;
assign v_3452 = v_3251 & v_3450;
assign v_3453 = ~v_3187 & v_3450;
assign v_3455 = ~v_3188 & v_3252;
assign v_3456 = v_3252 & v_3454;
assign v_3457 = ~v_3188 & v_3454;
assign v_3459 = ~v_3189 & v_3253;
assign v_3460 = v_3253 & v_3458;
assign v_3461 = ~v_3189 & v_3458;
assign v_3463 = ~v_3190 & v_3254;
assign v_3464 = v_3254 & v_3462;
assign v_3465 = ~v_3190 & v_3462;
assign v_3467 = ~v_3191 & v_3255;
assign v_3468 = v_3255 & v_3466;
assign v_3469 = ~v_3191 & v_3466;
assign v_3471 = ~v_3192 & v_3256;
assign v_3472 = v_3256 & v_3470;
assign v_3473 = ~v_3192 & v_3470;
assign v_3475 = ~v_3193 & v_3257;
assign v_3476 = v_3257 & v_3474;
assign v_3477 = ~v_3193 & v_3474;
assign v_3479 = ~v_3194 & v_3258;
assign v_3480 = v_3258 & v_3478;
assign v_3481 = ~v_3194 & v_3478;
assign v_3483 = ~v_3195 & v_3259;
assign v_3484 = v_3259 & v_3482;
assign v_3485 = ~v_3195 & v_3482;
assign v_3487 = ~v_3196 & v_3260;
assign v_3488 = v_3260 & v_3486;
assign v_3489 = ~v_3196 & v_3486;
assign v_3491 = ~v_3197 & v_3261;
assign v_3492 = v_3261 & v_3490;
assign v_3493 = ~v_3197 & v_3490;
assign v_3495 = ~v_3198 & v_3262;
assign v_3496 = v_3262 & v_3494;
assign v_3497 = ~v_3198 & v_3494;
assign v_3499 = ~v_3199 & v_3263;
assign v_3500 = v_3263 & v_3498;
assign v_3501 = ~v_3199 & v_3498;
assign v_3503 = ~v_3200 & v_3264;
assign v_3504 = v_3264 & v_3502;
assign v_3505 = ~v_3200 & v_3502;
assign v_3507 = ~v_3201 & v_3265;
assign v_3508 = v_3265 & v_3506;
assign v_3509 = ~v_3201 & v_3506;
assign v_3511 = ~v_3202 & v_3266;
assign v_3512 = v_3266 & v_3510;
assign v_3513 = ~v_3202 & v_3510;
assign v_3515 = ~v_3203 & v_3267;
assign v_3516 = v_3267 & v_3514;
assign v_3517 = ~v_3203 & v_3514;
assign v_3519 = ~v_3204 & v_3268;
assign v_3520 = v_3268 & v_3518;
assign v_3521 = ~v_3204 & v_3518;
assign v_3653 = ~v_3525 & v_3589;
assign v_3655 = ~v_3526 & v_3590;
assign v_3656 = v_3590 & v_3654;
assign v_3657 = ~v_3526 & v_3654;
assign v_3659 = ~v_3527 & v_3591;
assign v_3660 = v_3591 & v_3658;
assign v_3661 = ~v_3527 & v_3658;
assign v_3663 = ~v_3528 & v_3592;
assign v_3664 = v_3592 & v_3662;
assign v_3665 = ~v_3528 & v_3662;
assign v_3667 = ~v_3529 & v_3593;
assign v_3668 = v_3593 & v_3666;
assign v_3669 = ~v_3529 & v_3666;
assign v_3671 = ~v_3530 & v_3594;
assign v_3672 = v_3594 & v_3670;
assign v_3673 = ~v_3530 & v_3670;
assign v_3675 = ~v_3531 & v_3595;
assign v_3676 = v_3595 & v_3674;
assign v_3677 = ~v_3531 & v_3674;
assign v_3679 = ~v_3532 & v_3596;
assign v_3680 = v_3596 & v_3678;
assign v_3681 = ~v_3532 & v_3678;
assign v_3683 = ~v_3533 & v_3597;
assign v_3684 = v_3597 & v_3682;
assign v_3685 = ~v_3533 & v_3682;
assign v_3687 = ~v_3534 & v_3598;
assign v_3688 = v_3598 & v_3686;
assign v_3689 = ~v_3534 & v_3686;
assign v_3691 = ~v_3535 & v_3599;
assign v_3692 = v_3599 & v_3690;
assign v_3693 = ~v_3535 & v_3690;
assign v_3695 = ~v_3536 & v_3600;
assign v_3696 = v_3600 & v_3694;
assign v_3697 = ~v_3536 & v_3694;
assign v_3699 = ~v_3537 & v_3601;
assign v_3700 = v_3601 & v_3698;
assign v_3701 = ~v_3537 & v_3698;
assign v_3703 = ~v_3538 & v_3602;
assign v_3704 = v_3602 & v_3702;
assign v_3705 = ~v_3538 & v_3702;
assign v_3707 = ~v_3539 & v_3603;
assign v_3708 = v_3603 & v_3706;
assign v_3709 = ~v_3539 & v_3706;
assign v_3711 = ~v_3540 & v_3604;
assign v_3712 = v_3604 & v_3710;
assign v_3713 = ~v_3540 & v_3710;
assign v_3715 = ~v_3541 & v_3605;
assign v_3716 = v_3605 & v_3714;
assign v_3717 = ~v_3541 & v_3714;
assign v_3719 = ~v_3542 & v_3606;
assign v_3720 = v_3606 & v_3718;
assign v_3721 = ~v_3542 & v_3718;
assign v_3723 = ~v_3543 & v_3607;
assign v_3724 = v_3607 & v_3722;
assign v_3725 = ~v_3543 & v_3722;
assign v_3727 = ~v_3544 & v_3608;
assign v_3728 = v_3608 & v_3726;
assign v_3729 = ~v_3544 & v_3726;
assign v_3731 = ~v_3545 & v_3609;
assign v_3732 = v_3609 & v_3730;
assign v_3733 = ~v_3545 & v_3730;
assign v_3735 = ~v_3546 & v_3610;
assign v_3736 = v_3610 & v_3734;
assign v_3737 = ~v_3546 & v_3734;
assign v_3739 = ~v_3547 & v_3611;
assign v_3740 = v_3611 & v_3738;
assign v_3741 = ~v_3547 & v_3738;
assign v_3743 = ~v_3548 & v_3612;
assign v_3744 = v_3612 & v_3742;
assign v_3745 = ~v_3548 & v_3742;
assign v_3747 = ~v_3549 & v_3613;
assign v_3748 = v_3613 & v_3746;
assign v_3749 = ~v_3549 & v_3746;
assign v_3751 = ~v_3550 & v_3614;
assign v_3752 = v_3614 & v_3750;
assign v_3753 = ~v_3550 & v_3750;
assign v_3755 = ~v_3551 & v_3615;
assign v_3756 = v_3615 & v_3754;
assign v_3757 = ~v_3551 & v_3754;
assign v_3759 = ~v_3552 & v_3616;
assign v_3760 = v_3616 & v_3758;
assign v_3761 = ~v_3552 & v_3758;
assign v_3763 = ~v_3553 & v_3617;
assign v_3764 = v_3617 & v_3762;
assign v_3765 = ~v_3553 & v_3762;
assign v_3767 = ~v_3554 & v_3618;
assign v_3768 = v_3618 & v_3766;
assign v_3769 = ~v_3554 & v_3766;
assign v_3771 = ~v_3555 & v_3619;
assign v_3772 = v_3619 & v_3770;
assign v_3773 = ~v_3555 & v_3770;
assign v_3775 = ~v_3556 & v_3620;
assign v_3776 = v_3620 & v_3774;
assign v_3777 = ~v_3556 & v_3774;
assign v_3779 = ~v_3557 & v_3621;
assign v_3780 = v_3621 & v_3778;
assign v_3781 = ~v_3557 & v_3778;
assign v_3783 = ~v_3558 & v_3622;
assign v_3784 = v_3622 & v_3782;
assign v_3785 = ~v_3558 & v_3782;
assign v_3787 = ~v_3559 & v_3623;
assign v_3788 = v_3623 & v_3786;
assign v_3789 = ~v_3559 & v_3786;
assign v_3791 = ~v_3560 & v_3624;
assign v_3792 = v_3624 & v_3790;
assign v_3793 = ~v_3560 & v_3790;
assign v_3795 = ~v_3561 & v_3625;
assign v_3796 = v_3625 & v_3794;
assign v_3797 = ~v_3561 & v_3794;
assign v_3799 = ~v_3562 & v_3626;
assign v_3800 = v_3626 & v_3798;
assign v_3801 = ~v_3562 & v_3798;
assign v_3803 = ~v_3563 & v_3627;
assign v_3804 = v_3627 & v_3802;
assign v_3805 = ~v_3563 & v_3802;
assign v_3807 = ~v_3564 & v_3628;
assign v_3808 = v_3628 & v_3806;
assign v_3809 = ~v_3564 & v_3806;
assign v_3811 = ~v_3565 & v_3629;
assign v_3812 = v_3629 & v_3810;
assign v_3813 = ~v_3565 & v_3810;
assign v_3815 = ~v_3566 & v_3630;
assign v_3816 = v_3630 & v_3814;
assign v_3817 = ~v_3566 & v_3814;
assign v_3819 = ~v_3567 & v_3631;
assign v_3820 = v_3631 & v_3818;
assign v_3821 = ~v_3567 & v_3818;
assign v_3823 = ~v_3568 & v_3632;
assign v_3824 = v_3632 & v_3822;
assign v_3825 = ~v_3568 & v_3822;
assign v_3827 = ~v_3569 & v_3633;
assign v_3828 = v_3633 & v_3826;
assign v_3829 = ~v_3569 & v_3826;
assign v_3831 = ~v_3570 & v_3634;
assign v_3832 = v_3634 & v_3830;
assign v_3833 = ~v_3570 & v_3830;
assign v_3835 = ~v_3571 & v_3635;
assign v_3836 = v_3635 & v_3834;
assign v_3837 = ~v_3571 & v_3834;
assign v_3839 = ~v_3572 & v_3636;
assign v_3840 = v_3636 & v_3838;
assign v_3841 = ~v_3572 & v_3838;
assign v_3843 = ~v_3573 & v_3637;
assign v_3844 = v_3637 & v_3842;
assign v_3845 = ~v_3573 & v_3842;
assign v_3847 = ~v_3574 & v_3638;
assign v_3848 = v_3638 & v_3846;
assign v_3849 = ~v_3574 & v_3846;
assign v_3851 = ~v_3575 & v_3639;
assign v_3852 = v_3639 & v_3850;
assign v_3853 = ~v_3575 & v_3850;
assign v_3855 = ~v_3576 & v_3640;
assign v_3856 = v_3640 & v_3854;
assign v_3857 = ~v_3576 & v_3854;
assign v_3859 = ~v_3577 & v_3641;
assign v_3860 = v_3641 & v_3858;
assign v_3861 = ~v_3577 & v_3858;
assign v_3863 = ~v_3578 & v_3642;
assign v_3864 = v_3642 & v_3862;
assign v_3865 = ~v_3578 & v_3862;
assign v_3867 = ~v_3579 & v_3643;
assign v_3868 = v_3643 & v_3866;
assign v_3869 = ~v_3579 & v_3866;
assign v_3871 = ~v_3580 & v_3644;
assign v_3872 = v_3644 & v_3870;
assign v_3873 = ~v_3580 & v_3870;
assign v_3875 = ~v_3581 & v_3645;
assign v_3876 = v_3645 & v_3874;
assign v_3877 = ~v_3581 & v_3874;
assign v_3879 = ~v_3582 & v_3646;
assign v_3880 = v_3646 & v_3878;
assign v_3881 = ~v_3582 & v_3878;
assign v_3883 = ~v_3583 & v_3647;
assign v_3884 = v_3647 & v_3882;
assign v_3885 = ~v_3583 & v_3882;
assign v_3887 = ~v_3584 & v_3648;
assign v_3888 = v_3648 & v_3886;
assign v_3889 = ~v_3584 & v_3886;
assign v_3891 = ~v_3585 & v_3649;
assign v_3892 = v_3649 & v_3890;
assign v_3893 = ~v_3585 & v_3890;
assign v_3895 = ~v_3586 & v_3650;
assign v_3896 = v_3650 & v_3894;
assign v_3897 = ~v_3586 & v_3894;
assign v_3899 = ~v_3587 & v_3651;
assign v_3900 = v_3651 & v_3898;
assign v_3901 = ~v_3587 & v_3898;
assign v_3903 = ~v_3588 & v_3652;
assign v_3904 = v_3652 & v_3902;
assign v_3905 = ~v_3588 & v_3902;
assign v_3909 = ~v_3138 & ~v_3522 & ~v_3906;
assign v_3974 = v_4457 & v_4458 & v_4459;
assign v_4039 = v_4473 & v_4474 & v_4475;
assign v_4104 = v_4489 & v_4490 & v_4491;
assign v_4169 = v_4505 & v_4506 & v_4507;
assign v_4234 = v_4521 & v_4522 & v_4523;
assign v_4299 = v_4537 & v_4538 & v_4539;
assign v_4300 = ~v_1282 & ~v_1283 & ~v_1284 & ~v_1285 & ~v_1286;
assign v_4301 = ~v_1287 & ~v_1288 & ~v_1289 & ~v_1290 & ~v_1291;
assign v_4302 = ~v_1292 & ~v_1293 & ~v_1294 & ~v_1295 & ~v_1296;
assign v_4303 = ~v_1297 & ~v_1298 & ~v_1299 & ~v_1300 & ~v_1301;
assign v_4304 = ~v_1302 & ~v_1303 & ~v_1304 & ~v_1305 & ~v_1306;
assign v_4305 = ~v_1307 & ~v_1308 & ~v_1309 & ~v_1310 & ~v_1311;
assign v_4306 = ~v_1312 & ~v_1313 & ~v_1314 & ~v_1315 & ~v_1316;
assign v_4307 = ~v_1317 & ~v_1318 & ~v_1319 & ~v_1320 & ~v_1321;
assign v_4308 = ~v_1322 & ~v_1323 & ~v_1324 & ~v_1325 & ~v_1326;
assign v_4309 = ~v_1327 & ~v_1328 & ~v_1329 & ~v_1330 & ~v_1331;
assign v_4310 = ~v_1332 & ~v_1333 & ~v_1334 & ~v_1335 & ~v_1336;
assign v_4311 = ~v_1337 & ~v_1338 & ~v_1339 & ~v_1340 & ~v_1341;
assign v_4312 = ~v_1342 & ~v_1343 & ~v_1344 & ~v_1345;
assign v_4313 = v_4300 & v_4301 & v_4302 & v_4303 & v_4304;
assign v_4314 = v_4305 & v_4306 & v_4307 & v_4308 & v_4309;
assign v_4315 = v_4310 & v_4311 & v_4312;
assign v_4316 = ~v_1411 & ~v_1412 & ~v_1413 & ~v_1414 & ~v_1415;
assign v_4317 = ~v_1416 & ~v_1417 & ~v_1418 & ~v_1419 & ~v_1420;
assign v_4318 = ~v_1421 & ~v_1422 & ~v_1423 & ~v_1424 & ~v_1425;
assign v_4319 = ~v_1426 & ~v_1427 & ~v_1428 & ~v_1429 & ~v_1430;
assign v_4320 = ~v_1431 & ~v_1432 & ~v_1433 & ~v_1434 & ~v_1435;
assign v_4321 = ~v_1436 & ~v_1437 & ~v_1438 & ~v_1439 & ~v_1440;
assign v_4322 = ~v_1441 & ~v_1442 & ~v_1443 & ~v_1444 & ~v_1445;
assign v_4323 = ~v_1446 & ~v_1447 & ~v_1448 & ~v_1449 & ~v_1450;
assign v_4324 = ~v_1451 & ~v_1452 & ~v_1453 & ~v_1454 & ~v_1455;
assign v_4325 = ~v_1456 & ~v_1457 & ~v_1458 & ~v_1459 & ~v_1460;
assign v_4326 = ~v_1461 & ~v_1462 & ~v_1463 & ~v_1464 & ~v_1465;
assign v_4327 = ~v_1466 & ~v_1467 & ~v_1468 & ~v_1469 & ~v_1470;
assign v_4328 = ~v_1471 & ~v_1472 & ~v_1473 & ~v_1474;
assign v_4329 = v_4316 & v_4317 & v_4318 & v_4319 & v_4320;
assign v_4330 = v_4321 & v_4322 & v_4323 & v_4324 & v_4325;
assign v_4331 = v_4326 & v_4327 & v_4328;
assign v_4332 = ~v_1540 & ~v_1541 & ~v_1542 & ~v_1543 & ~v_1544;
assign v_4333 = ~v_1545 & ~v_1546 & ~v_1547 & ~v_1548 & ~v_1549;
assign v_4334 = ~v_1550 & ~v_1551 & ~v_1552 & ~v_1553 & ~v_1554;
assign v_4335 = ~v_1555 & ~v_1556 & ~v_1557 & ~v_1558 & ~v_1559;
assign v_4336 = ~v_1560 & ~v_1561 & ~v_1562 & ~v_1563 & ~v_1564;
assign v_4337 = ~v_1565 & ~v_1566 & ~v_1567 & ~v_1568 & ~v_1569;
assign v_4338 = ~v_1570 & ~v_1571 & ~v_1572 & ~v_1573 & ~v_1574;
assign v_4339 = ~v_1575 & ~v_1576 & ~v_1577 & ~v_1578 & ~v_1579;
assign v_4340 = ~v_1580 & ~v_1581 & ~v_1582 & ~v_1583 & ~v_1584;
assign v_4341 = ~v_1585 & ~v_1586 & ~v_1587 & ~v_1588 & ~v_1589;
assign v_4342 = ~v_1590 & ~v_1591 & ~v_1592 & ~v_1593 & ~v_1594;
assign v_4343 = ~v_1595 & ~v_1596 & ~v_1597 & ~v_1598 & ~v_1599;
assign v_4344 = ~v_1600 & ~v_1601 & ~v_1602 & ~v_1603;
assign v_4345 = v_4332 & v_4333 & v_4334 & v_4335 & v_4336;
assign v_4346 = v_4337 & v_4338 & v_4339 & v_4340 & v_4341;
assign v_4347 = v_4342 & v_4343 & v_4344;
assign v_4348 = ~v_1605 & ~v_1606 & ~v_1607 & ~v_1608 & ~v_1609;
assign v_4349 = ~v_1610 & ~v_1611 & ~v_1612 & ~v_1613 & ~v_1614;
assign v_4350 = ~v_1615 & ~v_1616 & ~v_1617 & ~v_1618 & ~v_1619;
assign v_4351 = ~v_1620 & ~v_1621 & ~v_1622 & ~v_1623 & ~v_1624;
assign v_4352 = ~v_1625 & ~v_1626 & ~v_1627 & ~v_1628 & ~v_1629;
assign v_4353 = ~v_1630 & ~v_1631 & ~v_1632 & ~v_1633 & ~v_1634;
assign v_4354 = ~v_1635 & ~v_1636 & ~v_1637 & ~v_1638 & ~v_1639;
assign v_4355 = ~v_1640 & ~v_1641 & ~v_1642 & ~v_1643 & ~v_1644;
assign v_4356 = ~v_1645 & ~v_1646 & ~v_1647 & ~v_1648 & ~v_1649;
assign v_4357 = ~v_1650 & ~v_1651 & ~v_1652 & ~v_1653 & ~v_1654;
assign v_4358 = ~v_1655 & ~v_1656 & ~v_1657 & ~v_1658 & ~v_1659;
assign v_4359 = ~v_1660 & ~v_1661 & ~v_1662 & ~v_1663 & ~v_1664;
assign v_4360 = ~v_1665 & ~v_1666 & ~v_1667 & ~v_1668;
assign v_4361 = v_4348 & v_4349 & v_4350 & v_4351 & v_4352;
assign v_4362 = v_4353 & v_4354 & v_4355 & v_4356 & v_4357;
assign v_4363 = v_4358 & v_4359 & v_4360;
assign v_4364 = ~v_2051 & ~v_2052 & ~v_2053 & ~v_2054 & ~v_2055;
assign v_4365 = ~v_2056 & ~v_2057 & ~v_2058 & ~v_2059 & ~v_2060;
assign v_4366 = ~v_2061 & ~v_2062 & ~v_2063 & ~v_2064 & ~v_2065;
assign v_4367 = ~v_2066 & ~v_2067 & ~v_2068 & ~v_2069 & ~v_2070;
assign v_4368 = ~v_2071 & ~v_2072 & ~v_2073 & ~v_2074 & ~v_2075;
assign v_4369 = ~v_2076 & ~v_2077 & ~v_2078 & ~v_2079 & ~v_2080;
assign v_4370 = ~v_2081 & ~v_2082 & ~v_2083 & ~v_2084 & ~v_2085;
assign v_4371 = ~v_2086 & ~v_2087 & ~v_2088 & ~v_2089 & ~v_2090;
assign v_4372 = ~v_2091 & ~v_2092 & ~v_2093 & ~v_2094 & ~v_2095;
assign v_4373 = ~v_2096 & ~v_2097 & ~v_2098 & ~v_2099 & ~v_2100;
assign v_4374 = ~v_2101 & ~v_2102 & ~v_2103 & ~v_2104 & ~v_2105;
assign v_4375 = ~v_2106 & ~v_2107 & ~v_2108 & ~v_2109 & ~v_2110;
assign v_4376 = ~v_2111 & ~v_2112 & ~v_2113 & ~v_2114;
assign v_4377 = v_4364 & v_4365 & v_4366 & v_4367 & v_4368;
assign v_4378 = v_4369 & v_4370 & v_4371 & v_4372 & v_4373;
assign v_4379 = v_4374 & v_4375 & v_4376;
assign v_4380 = ~v_2116 & ~v_2117 & ~v_2118 & ~v_2119 & ~v_2120;
assign v_4381 = ~v_2121 & ~v_2122 & ~v_2123 & ~v_2124 & ~v_2125;
assign v_4382 = ~v_2126 & ~v_2127 & ~v_2128 & ~v_2129 & ~v_2130;
assign v_4383 = ~v_2131 & ~v_2132 & ~v_2133 & ~v_2134 & ~v_2135;
assign v_4384 = ~v_2136 & ~v_2137 & ~v_2138 & ~v_2139 & ~v_2140;
assign v_4385 = ~v_2141 & ~v_2142 & ~v_2143 & ~v_2144 & ~v_2145;
assign v_4386 = ~v_2146 & ~v_2147 & ~v_2148 & ~v_2149 & ~v_2150;
assign v_4387 = ~v_2151 & ~v_2152 & ~v_2153 & ~v_2154 & ~v_2155;
assign v_4388 = ~v_2156 & ~v_2157 & ~v_2158 & ~v_2159 & ~v_2160;
assign v_4389 = ~v_2161 & ~v_2162 & ~v_2163 & ~v_2164 & ~v_2165;
assign v_4390 = ~v_2166 & ~v_2167 & ~v_2168 & ~v_2169 & ~v_2170;
assign v_4391 = ~v_2171 & ~v_2172 & ~v_2173 & ~v_2174 & ~v_2175;
assign v_4392 = ~v_2176 & ~v_2177 & ~v_2178 & ~v_2179;
assign v_4393 = v_4380 & v_4381 & v_4382 & v_4383 & v_4384;
assign v_4394 = v_4385 & v_4386 & v_4387 & v_4388 & v_4389;
assign v_4395 = v_4390 & v_4391 & v_4392;
assign v_4396 = ~v_2562 & ~v_2563 & ~v_2564 & ~v_2565 & ~v_2566;
assign v_4397 = ~v_2567 & ~v_2568 & ~v_2569 & ~v_2570 & ~v_2571;
assign v_4398 = ~v_2572 & ~v_2573 & ~v_2574 & ~v_2575 & ~v_2576;
assign v_4399 = ~v_2577 & ~v_2578 & ~v_2579 & ~v_2580 & ~v_2581;
assign v_4400 = ~v_2582 & ~v_2583 & ~v_2584 & ~v_2585 & ~v_2586;
assign v_4401 = ~v_2587 & ~v_2588 & ~v_2589 & ~v_2590 & ~v_2591;
assign v_4402 = ~v_2592 & ~v_2593 & ~v_2594 & ~v_2595 & ~v_2596;
assign v_4403 = ~v_2597 & ~v_2598 & ~v_2599 & ~v_2600 & ~v_2601;
assign v_4404 = ~v_2602 & ~v_2603 & ~v_2604 & ~v_2605 & ~v_2606;
assign v_4405 = ~v_2607 & ~v_2608 & ~v_2609 & ~v_2610 & ~v_2611;
assign v_4406 = ~v_2612 & ~v_2613 & ~v_2614 & ~v_2615 & ~v_2616;
assign v_4407 = ~v_2617 & ~v_2618 & ~v_2619 & ~v_2620 & ~v_2621;
assign v_4408 = ~v_2622 & ~v_2623 & ~v_2624 & ~v_2625;
assign v_4409 = v_4396 & v_4397 & v_4398 & v_4399 & v_4400;
assign v_4410 = v_4401 & v_4402 & v_4403 & v_4404 & v_4405;
assign v_4411 = v_4406 & v_4407 & v_4408;
assign v_4412 = ~v_2627 & ~v_2628 & ~v_2629 & ~v_2630 & ~v_2631;
assign v_4413 = ~v_2632 & ~v_2633 & ~v_2634 & ~v_2635 & ~v_2636;
assign v_4414 = ~v_2637 & ~v_2638 & ~v_2639 & ~v_2640 & ~v_2641;
assign v_4415 = ~v_2642 & ~v_2643 & ~v_2644 & ~v_2645 & ~v_2646;
assign v_4416 = ~v_2647 & ~v_2648 & ~v_2649 & ~v_2650 & ~v_2651;
assign v_4417 = ~v_2652 & ~v_2653 & ~v_2654 & ~v_2655 & ~v_2656;
assign v_4418 = ~v_2657 & ~v_2658 & ~v_2659 & ~v_2660 & ~v_2661;
assign v_4419 = ~v_2662 & ~v_2663 & ~v_2664 & ~v_2665 & ~v_2666;
assign v_4420 = ~v_2667 & ~v_2668 & ~v_2669 & ~v_2670 & ~v_2671;
assign v_4421 = ~v_2672 & ~v_2673 & ~v_2674 & ~v_2675 & ~v_2676;
assign v_4422 = ~v_2677 & ~v_2678 & ~v_2679 & ~v_2680 & ~v_2681;
assign v_4423 = ~v_2682 & ~v_2683 & ~v_2684 & ~v_2685 & ~v_2686;
assign v_4424 = ~v_2687 & ~v_2688 & ~v_2689 & ~v_2690;
assign v_4425 = v_4412 & v_4413 & v_4414 & v_4415 & v_4416;
assign v_4426 = v_4417 & v_4418 & v_4419 & v_4420 & v_4421;
assign v_4427 = v_4422 & v_4423 & v_4424;
assign v_4428 = ~v_2692 & ~v_2693 & ~v_2694 & ~v_2695 & ~v_2696;
assign v_4429 = ~v_2697 & ~v_2698 & ~v_2699 & ~v_2700 & ~v_2701;
assign v_4430 = ~v_2702 & ~v_2703 & ~v_2704 & ~v_2705 & ~v_2706;
assign v_4431 = ~v_2707 & ~v_2708 & ~v_2709 & ~v_2710 & ~v_2711;
assign v_4432 = ~v_2712 & ~v_2713 & ~v_2714 & ~v_2715 & ~v_2716;
assign v_4433 = ~v_2717 & ~v_2718 & ~v_2719 & ~v_2720 & ~v_2721;
assign v_4434 = ~v_2722 & ~v_2723 & ~v_2724 & ~v_2725 & ~v_2726;
assign v_4435 = ~v_2727 & ~v_2728 & ~v_2729 & ~v_2730 & ~v_2731;
assign v_4436 = ~v_2732 & ~v_2733 & ~v_2734 & ~v_2735 & ~v_2736;
assign v_4437 = ~v_2737 & ~v_2738 & ~v_2739 & ~v_2740 & ~v_2741;
assign v_4438 = ~v_2742 & ~v_2743 & ~v_2744 & ~v_2745 & ~v_2746;
assign v_4439 = ~v_2747 & ~v_2748 & ~v_2749 & ~v_2750 & ~v_2751;
assign v_4440 = ~v_2752 & ~v_2753 & ~v_2754 & ~v_2755;
assign v_4441 = v_4428 & v_4429 & v_4430 & v_4431 & v_4432;
assign v_4442 = v_4433 & v_4434 & v_4435 & v_4436 & v_4437;
assign v_4443 = v_4438 & v_4439 & v_4440;
assign v_4444 = ~v_3910 & ~v_3911 & ~v_3912 & ~v_3913 & ~v_3914;
assign v_4445 = ~v_3915 & ~v_3916 & ~v_3917 & ~v_3918 & ~v_3919;
assign v_4446 = ~v_3920 & ~v_3921 & ~v_3922 & ~v_3923 & ~v_3924;
assign v_4447 = ~v_3925 & ~v_3926 & ~v_3927 & ~v_3928 & ~v_3929;
assign v_4448 = ~v_3930 & ~v_3931 & ~v_3932 & ~v_3933 & ~v_3934;
assign v_4449 = ~v_3935 & ~v_3936 & ~v_3937 & ~v_3938 & ~v_3939;
assign v_4450 = ~v_3940 & ~v_3941 & ~v_3942 & ~v_3943 & ~v_3944;
assign v_4451 = ~v_3945 & ~v_3946 & ~v_3947 & ~v_3948 & ~v_3949;
assign v_4452 = ~v_3950 & ~v_3951 & ~v_3952 & ~v_3953 & ~v_3954;
assign v_4453 = ~v_3955 & ~v_3956 & ~v_3957 & ~v_3958 & ~v_3959;
assign v_4454 = ~v_3960 & ~v_3961 & ~v_3962 & ~v_3963 & ~v_3964;
assign v_4455 = ~v_3965 & ~v_3966 & ~v_3967 & ~v_3968 & ~v_3969;
assign v_4456 = ~v_3970 & ~v_3971 & ~v_3972 & ~v_3973;
assign v_4457 = v_4444 & v_4445 & v_4446 & v_4447 & v_4448;
assign v_4458 = v_4449 & v_4450 & v_4451 & v_4452 & v_4453;
assign v_4459 = v_4454 & v_4455 & v_4456;
assign v_4460 = ~v_3975 & ~v_3976 & ~v_3977 & ~v_3978 & ~v_3979;
assign v_4461 = ~v_3980 & ~v_3981 & ~v_3982 & ~v_3983 & ~v_3984;
assign v_4462 = ~v_3985 & ~v_3986 & ~v_3987 & ~v_3988 & ~v_3989;
assign v_4463 = ~v_3990 & ~v_3991 & ~v_3992 & ~v_3993 & ~v_3994;
assign v_4464 = ~v_3995 & ~v_3996 & ~v_3997 & ~v_3998 & ~v_3999;
assign v_4465 = ~v_4000 & ~v_4001 & ~v_4002 & ~v_4003 & ~v_4004;
assign v_4466 = ~v_4005 & ~v_4006 & ~v_4007 & ~v_4008 & ~v_4009;
assign v_4467 = ~v_4010 & ~v_4011 & ~v_4012 & ~v_4013 & ~v_4014;
assign v_4468 = ~v_4015 & ~v_4016 & ~v_4017 & ~v_4018 & ~v_4019;
assign v_4469 = ~v_4020 & ~v_4021 & ~v_4022 & ~v_4023 & ~v_4024;
assign v_4470 = ~v_4025 & ~v_4026 & ~v_4027 & ~v_4028 & ~v_4029;
assign v_4471 = ~v_4030 & ~v_4031 & ~v_4032 & ~v_4033 & ~v_4034;
assign v_4472 = ~v_4035 & ~v_4036 & ~v_4037 & ~v_4038;
assign v_4473 = v_4460 & v_4461 & v_4462 & v_4463 & v_4464;
assign v_4474 = v_4465 & v_4466 & v_4467 & v_4468 & v_4469;
assign v_4475 = v_4470 & v_4471 & v_4472;
assign v_4476 = ~v_4040 & ~v_4041 & ~v_4042 & ~v_4043 & ~v_4044;
assign v_4477 = ~v_4045 & ~v_4046 & ~v_4047 & ~v_4048 & ~v_4049;
assign v_4478 = ~v_4050 & ~v_4051 & ~v_4052 & ~v_4053 & ~v_4054;
assign v_4479 = ~v_4055 & ~v_4056 & ~v_4057 & ~v_4058 & ~v_4059;
assign v_4480 = ~v_4060 & ~v_4061 & ~v_4062 & ~v_4063 & ~v_4064;
assign v_4481 = ~v_4065 & ~v_4066 & ~v_4067 & ~v_4068 & ~v_4069;
assign v_4482 = ~v_4070 & ~v_4071 & ~v_4072 & ~v_4073 & ~v_4074;
assign v_4483 = ~v_4075 & ~v_4076 & ~v_4077 & ~v_4078 & ~v_4079;
assign v_4484 = ~v_4080 & ~v_4081 & ~v_4082 & ~v_4083 & ~v_4084;
assign v_4485 = ~v_4085 & ~v_4086 & ~v_4087 & ~v_4088 & ~v_4089;
assign v_4486 = ~v_4090 & ~v_4091 & ~v_4092 & ~v_4093 & ~v_4094;
assign v_4487 = ~v_4095 & ~v_4096 & ~v_4097 & ~v_4098 & ~v_4099;
assign v_4488 = ~v_4100 & ~v_4101 & ~v_4102 & ~v_4103;
assign v_4489 = v_4476 & v_4477 & v_4478 & v_4479 & v_4480;
assign v_4490 = v_4481 & v_4482 & v_4483 & v_4484 & v_4485;
assign v_4491 = v_4486 & v_4487 & v_4488;
assign v_4492 = ~v_4105 & ~v_4106 & ~v_4107 & ~v_4108 & ~v_4109;
assign v_4493 = ~v_4110 & ~v_4111 & ~v_4112 & ~v_4113 & ~v_4114;
assign v_4494 = ~v_4115 & ~v_4116 & ~v_4117 & ~v_4118 & ~v_4119;
assign v_4495 = ~v_4120 & ~v_4121 & ~v_4122 & ~v_4123 & ~v_4124;
assign v_4496 = ~v_4125 & ~v_4126 & ~v_4127 & ~v_4128 & ~v_4129;
assign v_4497 = ~v_4130 & ~v_4131 & ~v_4132 & ~v_4133 & ~v_4134;
assign v_4498 = ~v_4135 & ~v_4136 & ~v_4137 & ~v_4138 & ~v_4139;
assign v_4499 = ~v_4140 & ~v_4141 & ~v_4142 & ~v_4143 & ~v_4144;
assign v_4500 = ~v_4145 & ~v_4146 & ~v_4147 & ~v_4148 & ~v_4149;
assign v_4501 = ~v_4150 & ~v_4151 & ~v_4152 & ~v_4153 & ~v_4154;
assign v_4502 = ~v_4155 & ~v_4156 & ~v_4157 & ~v_4158 & ~v_4159;
assign v_4503 = ~v_4160 & ~v_4161 & ~v_4162 & ~v_4163 & ~v_4164;
assign v_4504 = ~v_4165 & ~v_4166 & ~v_4167 & ~v_4168;
assign v_4505 = v_4492 & v_4493 & v_4494 & v_4495 & v_4496;
assign v_4506 = v_4497 & v_4498 & v_4499 & v_4500 & v_4501;
assign v_4507 = v_4502 & v_4503 & v_4504;
assign v_4508 = ~v_4170 & ~v_4171 & ~v_4172 & ~v_4173 & ~v_4174;
assign v_4509 = ~v_4175 & ~v_4176 & ~v_4177 & ~v_4178 & ~v_4179;
assign v_4510 = ~v_4180 & ~v_4181 & ~v_4182 & ~v_4183 & ~v_4184;
assign v_4511 = ~v_4185 & ~v_4186 & ~v_4187 & ~v_4188 & ~v_4189;
assign v_4512 = ~v_4190 & ~v_4191 & ~v_4192 & ~v_4193 & ~v_4194;
assign v_4513 = ~v_4195 & ~v_4196 & ~v_4197 & ~v_4198 & ~v_4199;
assign v_4514 = ~v_4200 & ~v_4201 & ~v_4202 & ~v_4203 & ~v_4204;
assign v_4515 = ~v_4205 & ~v_4206 & ~v_4207 & ~v_4208 & ~v_4209;
assign v_4516 = ~v_4210 & ~v_4211 & ~v_4212 & ~v_4213 & ~v_4214;
assign v_4517 = ~v_4215 & ~v_4216 & ~v_4217 & ~v_4218 & ~v_4219;
assign v_4518 = ~v_4220 & ~v_4221 & ~v_4222 & ~v_4223 & ~v_4224;
assign v_4519 = ~v_4225 & ~v_4226 & ~v_4227 & ~v_4228 & ~v_4229;
assign v_4520 = ~v_4230 & ~v_4231 & ~v_4232 & ~v_4233;
assign v_4521 = v_4508 & v_4509 & v_4510 & v_4511 & v_4512;
assign v_4522 = v_4513 & v_4514 & v_4515 & v_4516 & v_4517;
assign v_4523 = v_4518 & v_4519 & v_4520;
assign v_4524 = ~v_4235 & ~v_4236 & ~v_4237 & ~v_4238 & ~v_4239;
assign v_4525 = ~v_4240 & ~v_4241 & ~v_4242 & ~v_4243 & ~v_4244;
assign v_4526 = ~v_4245 & ~v_4246 & ~v_4247 & ~v_4248 & ~v_4249;
assign v_4527 = ~v_4250 & ~v_4251 & ~v_4252 & ~v_4253 & ~v_4254;
assign v_4528 = ~v_4255 & ~v_4256 & ~v_4257 & ~v_4258 & ~v_4259;
assign v_4529 = ~v_4260 & ~v_4261 & ~v_4262 & ~v_4263 & ~v_4264;
assign v_4530 = ~v_4265 & ~v_4266 & ~v_4267 & ~v_4268 & ~v_4269;
assign v_4531 = ~v_4270 & ~v_4271 & ~v_4272 & ~v_4273 & ~v_4274;
assign v_4532 = ~v_4275 & ~v_4276 & ~v_4277 & ~v_4278 & ~v_4279;
assign v_4533 = ~v_4280 & ~v_4281 & ~v_4282 & ~v_4283 & ~v_4284;
assign v_4534 = ~v_4285 & ~v_4286 & ~v_4287 & ~v_4288 & ~v_4289;
assign v_4535 = ~v_4290 & ~v_4291 & ~v_4292 & ~v_4293 & ~v_4294;
assign v_4536 = ~v_4295 & ~v_4296 & ~v_4297 & ~v_4298;
assign v_4537 = v_4524 & v_4525 & v_4526 & v_4527 & v_4528;
assign v_4538 = v_4529 & v_4530 & v_4531 & v_4532 & v_4533;
assign v_4539 = v_4534 & v_4535 & v_4536;
assign v_706 = v_450 | v_705 | ~v_514;
assign v_712 = v_709 | v_710 | v_711;
assign v_718 = v_715 | v_716 | v_717;
assign v_724 = v_721 | v_722 | v_723;
assign v_730 = v_727 | v_728 | v_729;
assign v_736 = v_733 | v_734 | v_735;
assign v_742 = v_739 | v_740 | v_741;
assign v_748 = v_745 | v_746 | v_747;
assign v_754 = v_751 | v_752 | v_753;
assign v_760 = v_757 | v_758 | v_759;
assign v_766 = v_763 | v_764 | v_765;
assign v_772 = v_769 | v_770 | v_771;
assign v_778 = v_775 | v_776 | v_777;
assign v_784 = v_781 | v_782 | v_783;
assign v_790 = v_787 | v_788 | v_789;
assign v_796 = v_793 | v_794 | v_795;
assign v_802 = v_799 | v_800 | v_801;
assign v_808 = v_805 | v_806 | v_807;
assign v_814 = v_811 | v_812 | v_813;
assign v_820 = v_817 | v_818 | v_819;
assign v_826 = v_823 | v_824 | v_825;
assign v_832 = v_829 | v_830 | v_831;
assign v_838 = v_835 | v_836 | v_837;
assign v_844 = v_841 | v_842 | v_843;
assign v_850 = v_847 | v_848 | v_849;
assign v_856 = v_853 | v_854 | v_855;
assign v_862 = v_859 | v_860 | v_861;
assign v_868 = v_865 | v_866 | v_867;
assign v_874 = v_871 | v_872 | v_873;
assign v_880 = v_877 | v_878 | v_879;
assign v_886 = v_883 | v_884 | v_885;
assign v_892 = v_889 | v_890 | v_891;
assign v_898 = v_895 | v_896 | v_897;
assign v_904 = v_901 | v_902 | v_903;
assign v_910 = v_907 | v_908 | v_909;
assign v_916 = v_913 | v_914 | v_915;
assign v_922 = v_919 | v_920 | v_921;
assign v_928 = v_925 | v_926 | v_927;
assign v_934 = v_931 | v_932 | v_933;
assign v_940 = v_937 | v_938 | v_939;
assign v_946 = v_943 | v_944 | v_945;
assign v_952 = v_949 | v_950 | v_951;
assign v_958 = v_955 | v_956 | v_957;
assign v_964 = v_961 | v_962 | v_963;
assign v_970 = v_967 | v_968 | v_969;
assign v_976 = v_973 | v_974 | v_975;
assign v_982 = v_979 | v_980 | v_981;
assign v_988 = v_985 | v_986 | v_987;
assign v_994 = v_991 | v_992 | v_993;
assign v_1000 = v_997 | v_998 | v_999;
assign v_1006 = v_1003 | v_1004 | v_1005;
assign v_1012 = v_1009 | v_1010 | v_1011;
assign v_1018 = v_1015 | v_1016 | v_1017;
assign v_1024 = v_1021 | v_1022 | v_1023;
assign v_1030 = v_1027 | v_1028 | v_1029;
assign v_1036 = v_1033 | v_1034 | v_1035;
assign v_1042 = v_1039 | v_1040 | v_1041;
assign v_1048 = v_1045 | v_1046 | v_1047;
assign v_1054 = v_1051 | v_1052 | v_1053;
assign v_1060 = v_1057 | v_1058 | v_1059;
assign v_1066 = v_1063 | v_1064 | v_1065;
assign v_1072 = v_1069 | v_1070 | v_1071;
assign v_1078 = v_1075 | v_1076 | v_1077;
assign v_1084 = v_1081 | v_1082 | v_1083;
assign v_1085 = v_4553 | v_4554 | v_4555;
assign v_1086 = ~v_1084 | ~v_1085;
assign v_1678 = v_1675 | v_1676 | v_1677;
assign v_1684 = v_1681 | v_1682 | v_1683;
assign v_1690 = v_1687 | v_1688 | v_1689;
assign v_1696 = v_1693 | v_1694 | v_1695;
assign v_1702 = v_1699 | v_1700 | v_1701;
assign v_1708 = v_1705 | v_1706 | v_1707;
assign v_1714 = v_1711 | v_1712 | v_1713;
assign v_1720 = v_1717 | v_1718 | v_1719;
assign v_1726 = v_1723 | v_1724 | v_1725;
assign v_1732 = v_1729 | v_1730 | v_1731;
assign v_1738 = v_1735 | v_1736 | v_1737;
assign v_1744 = v_1741 | v_1742 | v_1743;
assign v_1750 = v_1747 | v_1748 | v_1749;
assign v_1756 = v_1753 | v_1754 | v_1755;
assign v_1762 = v_1759 | v_1760 | v_1761;
assign v_1768 = v_1765 | v_1766 | v_1767;
assign v_1774 = v_1771 | v_1772 | v_1773;
assign v_1780 = v_1777 | v_1778 | v_1779;
assign v_1786 = v_1783 | v_1784 | v_1785;
assign v_1792 = v_1789 | v_1790 | v_1791;
assign v_1798 = v_1795 | v_1796 | v_1797;
assign v_1804 = v_1801 | v_1802 | v_1803;
assign v_1810 = v_1807 | v_1808 | v_1809;
assign v_1816 = v_1813 | v_1814 | v_1815;
assign v_1822 = v_1819 | v_1820 | v_1821;
assign v_1828 = v_1825 | v_1826 | v_1827;
assign v_1834 = v_1831 | v_1832 | v_1833;
assign v_1840 = v_1837 | v_1838 | v_1839;
assign v_1846 = v_1843 | v_1844 | v_1845;
assign v_1852 = v_1849 | v_1850 | v_1851;
assign v_1858 = v_1855 | v_1856 | v_1857;
assign v_1864 = v_1861 | v_1862 | v_1863;
assign v_1870 = v_1867 | v_1868 | v_1869;
assign v_1876 = v_1873 | v_1874 | v_1875;
assign v_1882 = v_1879 | v_1880 | v_1881;
assign v_1888 = v_1885 | v_1886 | v_1887;
assign v_1894 = v_1891 | v_1892 | v_1893;
assign v_1900 = v_1897 | v_1898 | v_1899;
assign v_1906 = v_1903 | v_1904 | v_1905;
assign v_1912 = v_1909 | v_1910 | v_1911;
assign v_1918 = v_1915 | v_1916 | v_1917;
assign v_1924 = v_1921 | v_1922 | v_1923;
assign v_1930 = v_1927 | v_1928 | v_1929;
assign v_1936 = v_1933 | v_1934 | v_1935;
assign v_1942 = v_1939 | v_1940 | v_1941;
assign v_1948 = v_1945 | v_1946 | v_1947;
assign v_1954 = v_1951 | v_1952 | v_1953;
assign v_1960 = v_1957 | v_1958 | v_1959;
assign v_1966 = v_1963 | v_1964 | v_1965;
assign v_1972 = v_1969 | v_1970 | v_1971;
assign v_1978 = v_1975 | v_1976 | v_1977;
assign v_1984 = v_1981 | v_1982 | v_1983;
assign v_1990 = v_1987 | v_1988 | v_1989;
assign v_1996 = v_1993 | v_1994 | v_1995;
assign v_2002 = v_1999 | v_2000 | v_2001;
assign v_2008 = v_2005 | v_2006 | v_2007;
assign v_2014 = v_2011 | v_2012 | v_2013;
assign v_2020 = v_2017 | v_2018 | v_2019;
assign v_2026 = v_2023 | v_2024 | v_2025;
assign v_2032 = v_2029 | v_2030 | v_2031;
assign v_2038 = v_2035 | v_2036 | v_2037;
assign v_2044 = v_2041 | v_2042 | v_2043;
assign v_2050 = v_2047 | v_2048 | v_2049;
assign v_2189 = v_2186 | v_2187 | v_2188;
assign v_2195 = v_2192 | v_2193 | v_2194;
assign v_2201 = v_2198 | v_2199 | v_2200;
assign v_2207 = v_2204 | v_2205 | v_2206;
assign v_2213 = v_2210 | v_2211 | v_2212;
assign v_2219 = v_2216 | v_2217 | v_2218;
assign v_2225 = v_2222 | v_2223 | v_2224;
assign v_2231 = v_2228 | v_2229 | v_2230;
assign v_2237 = v_2234 | v_2235 | v_2236;
assign v_2243 = v_2240 | v_2241 | v_2242;
assign v_2249 = v_2246 | v_2247 | v_2248;
assign v_2255 = v_2252 | v_2253 | v_2254;
assign v_2261 = v_2258 | v_2259 | v_2260;
assign v_2267 = v_2264 | v_2265 | v_2266;
assign v_2273 = v_2270 | v_2271 | v_2272;
assign v_2279 = v_2276 | v_2277 | v_2278;
assign v_2285 = v_2282 | v_2283 | v_2284;
assign v_2291 = v_2288 | v_2289 | v_2290;
assign v_2297 = v_2294 | v_2295 | v_2296;
assign v_2303 = v_2300 | v_2301 | v_2302;
assign v_2309 = v_2306 | v_2307 | v_2308;
assign v_2315 = v_2312 | v_2313 | v_2314;
assign v_2321 = v_2318 | v_2319 | v_2320;
assign v_2327 = v_2324 | v_2325 | v_2326;
assign v_2333 = v_2330 | v_2331 | v_2332;
assign v_2339 = v_2336 | v_2337 | v_2338;
assign v_2345 = v_2342 | v_2343 | v_2344;
assign v_2351 = v_2348 | v_2349 | v_2350;
assign v_2357 = v_2354 | v_2355 | v_2356;
assign v_2363 = v_2360 | v_2361 | v_2362;
assign v_2369 = v_2366 | v_2367 | v_2368;
assign v_2375 = v_2372 | v_2373 | v_2374;
assign v_2381 = v_2378 | v_2379 | v_2380;
assign v_2387 = v_2384 | v_2385 | v_2386;
assign v_2393 = v_2390 | v_2391 | v_2392;
assign v_2399 = v_2396 | v_2397 | v_2398;
assign v_2405 = v_2402 | v_2403 | v_2404;
assign v_2411 = v_2408 | v_2409 | v_2410;
assign v_2417 = v_2414 | v_2415 | v_2416;
assign v_2423 = v_2420 | v_2421 | v_2422;
assign v_2429 = v_2426 | v_2427 | v_2428;
assign v_2435 = v_2432 | v_2433 | v_2434;
assign v_2441 = v_2438 | v_2439 | v_2440;
assign v_2447 = v_2444 | v_2445 | v_2446;
assign v_2453 = v_2450 | v_2451 | v_2452;
assign v_2459 = v_2456 | v_2457 | v_2458;
assign v_2465 = v_2462 | v_2463 | v_2464;
assign v_2471 = v_2468 | v_2469 | v_2470;
assign v_2477 = v_2474 | v_2475 | v_2476;
assign v_2483 = v_2480 | v_2481 | v_2482;
assign v_2489 = v_2486 | v_2487 | v_2488;
assign v_2495 = v_2492 | v_2493 | v_2494;
assign v_2501 = v_2498 | v_2499 | v_2500;
assign v_2507 = v_2504 | v_2505 | v_2506;
assign v_2513 = v_2510 | v_2511 | v_2512;
assign v_2519 = v_2516 | v_2517 | v_2518;
assign v_2525 = v_2522 | v_2523 | v_2524;
assign v_2531 = v_2528 | v_2529 | v_2530;
assign v_2537 = v_2534 | v_2535 | v_2536;
assign v_2543 = v_2540 | v_2541 | v_2542;
assign v_2549 = v_2546 | v_2547 | v_2548;
assign v_2555 = v_2552 | v_2553 | v_2554;
assign v_2561 = v_2558 | v_2559 | v_2560;
assign v_2886 = v_2821 | v_2885 | ~v_2757;
assign v_2890 = v_2887 | v_2888 | v_2889;
assign v_2894 = v_2891 | v_2892 | v_2893;
assign v_2898 = v_2895 | v_2896 | v_2897;
assign v_2902 = v_2899 | v_2900 | v_2901;
assign v_2906 = v_2903 | v_2904 | v_2905;
assign v_2910 = v_2907 | v_2908 | v_2909;
assign v_2914 = v_2911 | v_2912 | v_2913;
assign v_2918 = v_2915 | v_2916 | v_2917;
assign v_2922 = v_2919 | v_2920 | v_2921;
assign v_2926 = v_2923 | v_2924 | v_2925;
assign v_2930 = v_2927 | v_2928 | v_2929;
assign v_2934 = v_2931 | v_2932 | v_2933;
assign v_2938 = v_2935 | v_2936 | v_2937;
assign v_2942 = v_2939 | v_2940 | v_2941;
assign v_2946 = v_2943 | v_2944 | v_2945;
assign v_2950 = v_2947 | v_2948 | v_2949;
assign v_2954 = v_2951 | v_2952 | v_2953;
assign v_2958 = v_2955 | v_2956 | v_2957;
assign v_2962 = v_2959 | v_2960 | v_2961;
assign v_2966 = v_2963 | v_2964 | v_2965;
assign v_2970 = v_2967 | v_2968 | v_2969;
assign v_2974 = v_2971 | v_2972 | v_2973;
assign v_2978 = v_2975 | v_2976 | v_2977;
assign v_2982 = v_2979 | v_2980 | v_2981;
assign v_2986 = v_2983 | v_2984 | v_2985;
assign v_2990 = v_2987 | v_2988 | v_2989;
assign v_2994 = v_2991 | v_2992 | v_2993;
assign v_2998 = v_2995 | v_2996 | v_2997;
assign v_3002 = v_2999 | v_3000 | v_3001;
assign v_3006 = v_3003 | v_3004 | v_3005;
assign v_3010 = v_3007 | v_3008 | v_3009;
assign v_3014 = v_3011 | v_3012 | v_3013;
assign v_3018 = v_3015 | v_3016 | v_3017;
assign v_3022 = v_3019 | v_3020 | v_3021;
assign v_3026 = v_3023 | v_3024 | v_3025;
assign v_3030 = v_3027 | v_3028 | v_3029;
assign v_3034 = v_3031 | v_3032 | v_3033;
assign v_3038 = v_3035 | v_3036 | v_3037;
assign v_3042 = v_3039 | v_3040 | v_3041;
assign v_3046 = v_3043 | v_3044 | v_3045;
assign v_3050 = v_3047 | v_3048 | v_3049;
assign v_3054 = v_3051 | v_3052 | v_3053;
assign v_3058 = v_3055 | v_3056 | v_3057;
assign v_3062 = v_3059 | v_3060 | v_3061;
assign v_3066 = v_3063 | v_3064 | v_3065;
assign v_3070 = v_3067 | v_3068 | v_3069;
assign v_3074 = v_3071 | v_3072 | v_3073;
assign v_3078 = v_3075 | v_3076 | v_3077;
assign v_3082 = v_3079 | v_3080 | v_3081;
assign v_3086 = v_3083 | v_3084 | v_3085;
assign v_3090 = v_3087 | v_3088 | v_3089;
assign v_3094 = v_3091 | v_3092 | v_3093;
assign v_3098 = v_3095 | v_3096 | v_3097;
assign v_3102 = v_3099 | v_3100 | v_3101;
assign v_3106 = v_3103 | v_3104 | v_3105;
assign v_3110 = v_3107 | v_3108 | v_3109;
assign v_3114 = v_3111 | v_3112 | v_3113;
assign v_3118 = v_3115 | v_3116 | v_3117;
assign v_3122 = v_3119 | v_3120 | v_3121;
assign v_3126 = v_3123 | v_3124 | v_3125;
assign v_3130 = v_3127 | v_3128 | v_3129;
assign v_3134 = v_3131 | v_3132 | v_3133;
assign v_3138 = v_3135 | v_3136 | v_3137;
assign v_3270 = v_3205 | v_3269 | ~v_3141;
assign v_3274 = v_3271 | v_3272 | v_3273;
assign v_3278 = v_3275 | v_3276 | v_3277;
assign v_3282 = v_3279 | v_3280 | v_3281;
assign v_3286 = v_3283 | v_3284 | v_3285;
assign v_3290 = v_3287 | v_3288 | v_3289;
assign v_3294 = v_3291 | v_3292 | v_3293;
assign v_3298 = v_3295 | v_3296 | v_3297;
assign v_3302 = v_3299 | v_3300 | v_3301;
assign v_3306 = v_3303 | v_3304 | v_3305;
assign v_3310 = v_3307 | v_3308 | v_3309;
assign v_3314 = v_3311 | v_3312 | v_3313;
assign v_3318 = v_3315 | v_3316 | v_3317;
assign v_3322 = v_3319 | v_3320 | v_3321;
assign v_3326 = v_3323 | v_3324 | v_3325;
assign v_3330 = v_3327 | v_3328 | v_3329;
assign v_3334 = v_3331 | v_3332 | v_3333;
assign v_3338 = v_3335 | v_3336 | v_3337;
assign v_3342 = v_3339 | v_3340 | v_3341;
assign v_3346 = v_3343 | v_3344 | v_3345;
assign v_3350 = v_3347 | v_3348 | v_3349;
assign v_3354 = v_3351 | v_3352 | v_3353;
assign v_3358 = v_3355 | v_3356 | v_3357;
assign v_3362 = v_3359 | v_3360 | v_3361;
assign v_3366 = v_3363 | v_3364 | v_3365;
assign v_3370 = v_3367 | v_3368 | v_3369;
assign v_3374 = v_3371 | v_3372 | v_3373;
assign v_3378 = v_3375 | v_3376 | v_3377;
assign v_3382 = v_3379 | v_3380 | v_3381;
assign v_3386 = v_3383 | v_3384 | v_3385;
assign v_3390 = v_3387 | v_3388 | v_3389;
assign v_3394 = v_3391 | v_3392 | v_3393;
assign v_3398 = v_3395 | v_3396 | v_3397;
assign v_3402 = v_3399 | v_3400 | v_3401;
assign v_3406 = v_3403 | v_3404 | v_3405;
assign v_3410 = v_3407 | v_3408 | v_3409;
assign v_3414 = v_3411 | v_3412 | v_3413;
assign v_3418 = v_3415 | v_3416 | v_3417;
assign v_3422 = v_3419 | v_3420 | v_3421;
assign v_3426 = v_3423 | v_3424 | v_3425;
assign v_3430 = v_3427 | v_3428 | v_3429;
assign v_3434 = v_3431 | v_3432 | v_3433;
assign v_3438 = v_3435 | v_3436 | v_3437;
assign v_3442 = v_3439 | v_3440 | v_3441;
assign v_3446 = v_3443 | v_3444 | v_3445;
assign v_3450 = v_3447 | v_3448 | v_3449;
assign v_3454 = v_3451 | v_3452 | v_3453;
assign v_3458 = v_3455 | v_3456 | v_3457;
assign v_3462 = v_3459 | v_3460 | v_3461;
assign v_3466 = v_3463 | v_3464 | v_3465;
assign v_3470 = v_3467 | v_3468 | v_3469;
assign v_3474 = v_3471 | v_3472 | v_3473;
assign v_3478 = v_3475 | v_3476 | v_3477;
assign v_3482 = v_3479 | v_3480 | v_3481;
assign v_3486 = v_3483 | v_3484 | v_3485;
assign v_3490 = v_3487 | v_3488 | v_3489;
assign v_3494 = v_3491 | v_3492 | v_3493;
assign v_3498 = v_3495 | v_3496 | v_3497;
assign v_3502 = v_3499 | v_3500 | v_3501;
assign v_3506 = v_3503 | v_3504 | v_3505;
assign v_3510 = v_3507 | v_3508 | v_3509;
assign v_3514 = v_3511 | v_3512 | v_3513;
assign v_3518 = v_3515 | v_3516 | v_3517;
assign v_3522 = v_3519 | v_3520 | v_3521;
assign v_3654 = v_3589 | v_3653 | ~v_3525;
assign v_3658 = v_3655 | v_3656 | v_3657;
assign v_3662 = v_3659 | v_3660 | v_3661;
assign v_3666 = v_3663 | v_3664 | v_3665;
assign v_3670 = v_3667 | v_3668 | v_3669;
assign v_3674 = v_3671 | v_3672 | v_3673;
assign v_3678 = v_3675 | v_3676 | v_3677;
assign v_3682 = v_3679 | v_3680 | v_3681;
assign v_3686 = v_3683 | v_3684 | v_3685;
assign v_3690 = v_3687 | v_3688 | v_3689;
assign v_3694 = v_3691 | v_3692 | v_3693;
assign v_3698 = v_3695 | v_3696 | v_3697;
assign v_3702 = v_3699 | v_3700 | v_3701;
assign v_3706 = v_3703 | v_3704 | v_3705;
assign v_3710 = v_3707 | v_3708 | v_3709;
assign v_3714 = v_3711 | v_3712 | v_3713;
assign v_3718 = v_3715 | v_3716 | v_3717;
assign v_3722 = v_3719 | v_3720 | v_3721;
assign v_3726 = v_3723 | v_3724 | v_3725;
assign v_3730 = v_3727 | v_3728 | v_3729;
assign v_3734 = v_3731 | v_3732 | v_3733;
assign v_3738 = v_3735 | v_3736 | v_3737;
assign v_3742 = v_3739 | v_3740 | v_3741;
assign v_3746 = v_3743 | v_3744 | v_3745;
assign v_3750 = v_3747 | v_3748 | v_3749;
assign v_3754 = v_3751 | v_3752 | v_3753;
assign v_3758 = v_3755 | v_3756 | v_3757;
assign v_3762 = v_3759 | v_3760 | v_3761;
assign v_3766 = v_3763 | v_3764 | v_3765;
assign v_3770 = v_3767 | v_3768 | v_3769;
assign v_3774 = v_3771 | v_3772 | v_3773;
assign v_3778 = v_3775 | v_3776 | v_3777;
assign v_3782 = v_3779 | v_3780 | v_3781;
assign v_3786 = v_3783 | v_3784 | v_3785;
assign v_3790 = v_3787 | v_3788 | v_3789;
assign v_3794 = v_3791 | v_3792 | v_3793;
assign v_3798 = v_3795 | v_3796 | v_3797;
assign v_3802 = v_3799 | v_3800 | v_3801;
assign v_3806 = v_3803 | v_3804 | v_3805;
assign v_3810 = v_3807 | v_3808 | v_3809;
assign v_3814 = v_3811 | v_3812 | v_3813;
assign v_3818 = v_3815 | v_3816 | v_3817;
assign v_3822 = v_3819 | v_3820 | v_3821;
assign v_3826 = v_3823 | v_3824 | v_3825;
assign v_3830 = v_3827 | v_3828 | v_3829;
assign v_3834 = v_3831 | v_3832 | v_3833;
assign v_3838 = v_3835 | v_3836 | v_3837;
assign v_3842 = v_3839 | v_3840 | v_3841;
assign v_3846 = v_3843 | v_3844 | v_3845;
assign v_3850 = v_3847 | v_3848 | v_3849;
assign v_3854 = v_3851 | v_3852 | v_3853;
assign v_3858 = v_3855 | v_3856 | v_3857;
assign v_3862 = v_3859 | v_3860 | v_3861;
assign v_3866 = v_3863 | v_3864 | v_3865;
assign v_3870 = v_3867 | v_3868 | v_3869;
assign v_3874 = v_3871 | v_3872 | v_3873;
assign v_3878 = v_3875 | v_3876 | v_3877;
assign v_3882 = v_3879 | v_3880 | v_3881;
assign v_3886 = v_3883 | v_3884 | v_3885;
assign v_3890 = v_3887 | v_3888 | v_3889;
assign v_3894 = v_3891 | v_3892 | v_3893;
assign v_3898 = v_3895 | v_3896 | v_3897;
assign v_3902 = v_3899 | v_3900 | v_3901;
assign v_3906 = v_3903 | v_3904 | v_3905;
assign v_4540 = v_708 | v_714 | v_720 | v_726 | v_732;
assign v_4541 = v_738 | v_744 | v_750 | v_756 | v_762;
assign v_4542 = v_768 | v_774 | v_780 | v_786 | v_792;
assign v_4543 = v_798 | v_804 | v_810 | v_816 | v_822;
assign v_4544 = v_828 | v_834 | v_840 | v_846 | v_852;
assign v_4545 = v_858 | v_864 | v_870 | v_876 | v_882;
assign v_4546 = v_888 | v_894 | v_900 | v_906 | v_912;
assign v_4547 = v_918 | v_924 | v_930 | v_936 | v_942;
assign v_4548 = v_948 | v_954 | v_960 | v_966 | v_972;
assign v_4549 = v_978 | v_984 | v_990 | v_996 | v_1002;
assign v_4550 = v_1008 | v_1014 | v_1020 | v_1026 | v_1032;
assign v_4551 = v_1038 | v_1044 | v_1050 | v_1056 | v_1062;
assign v_4552 = v_1068 | v_1074 | v_1080 | ~v_704;
assign v_4553 = v_4540 | v_4541 | v_4542 | v_4543 | v_4544;
assign v_4554 = v_4545 | v_4546 | v_4547 | v_4548 | v_4549;
assign v_4555 = v_4550 | v_4551 | v_4552;
assign v_579 = v_514 ^ v_515;
assign v_581 = ~v_516 ^ v_578;
assign v_583 = ~v_517 ^ v_580;
assign v_585 = ~v_518 ^ v_582;
assign v_587 = ~v_519 ^ v_584;
assign v_589 = ~v_520 ^ v_586;
assign v_591 = ~v_521 ^ v_588;
assign v_593 = ~v_522 ^ v_590;
assign v_595 = ~v_523 ^ v_592;
assign v_597 = ~v_524 ^ v_594;
assign v_599 = ~v_525 ^ v_596;
assign v_601 = ~v_526 ^ v_598;
assign v_603 = ~v_527 ^ v_600;
assign v_605 = ~v_528 ^ v_602;
assign v_607 = ~v_529 ^ v_604;
assign v_609 = ~v_530 ^ v_606;
assign v_611 = ~v_531 ^ v_608;
assign v_613 = ~v_532 ^ v_610;
assign v_615 = ~v_533 ^ v_612;
assign v_617 = ~v_534 ^ v_614;
assign v_619 = ~v_535 ^ v_616;
assign v_621 = ~v_536 ^ v_618;
assign v_623 = ~v_537 ^ v_620;
assign v_625 = ~v_538 ^ v_622;
assign v_627 = ~v_539 ^ v_624;
assign v_629 = ~v_540 ^ v_626;
assign v_631 = ~v_541 ^ v_628;
assign v_633 = ~v_542 ^ v_630;
assign v_635 = ~v_543 ^ v_632;
assign v_637 = ~v_544 ^ v_634;
assign v_639 = ~v_545 ^ v_636;
assign v_641 = ~v_546 ^ v_638;
assign v_643 = ~v_547 ^ v_640;
assign v_645 = ~v_548 ^ v_642;
assign v_647 = ~v_549 ^ v_644;
assign v_649 = ~v_550 ^ v_646;
assign v_651 = ~v_551 ^ v_648;
assign v_653 = ~v_552 ^ v_650;
assign v_655 = ~v_553 ^ v_652;
assign v_657 = ~v_554 ^ v_654;
assign v_659 = ~v_555 ^ v_656;
assign v_661 = ~v_556 ^ v_658;
assign v_663 = ~v_557 ^ v_660;
assign v_665 = ~v_558 ^ v_662;
assign v_667 = ~v_559 ^ v_664;
assign v_669 = ~v_560 ^ v_666;
assign v_671 = ~v_561 ^ v_668;
assign v_673 = ~v_562 ^ v_670;
assign v_675 = ~v_563 ^ v_672;
assign v_677 = ~v_564 ^ v_674;
assign v_679 = ~v_565 ^ v_676;
assign v_681 = ~v_566 ^ v_678;
assign v_683 = ~v_567 ^ v_680;
assign v_685 = ~v_568 ^ v_682;
assign v_687 = ~v_569 ^ v_684;
assign v_689 = ~v_570 ^ v_686;
assign v_691 = ~v_571 ^ v_688;
assign v_693 = ~v_572 ^ v_690;
assign v_695 = ~v_573 ^ v_692;
assign v_697 = ~v_574 ^ v_694;
assign v_699 = ~v_575 ^ v_696;
assign v_701 = ~v_576 ^ v_698;
assign v_703 = ~v_577 ^ v_700;
assign v_704 = v_450 ^ ~v_514;
assign v_707 = v_451 ^ ~v_579;
assign v_708 = v_707 ^ v_706;
assign v_713 = v_452 ^ ~v_581;
assign v_714 = v_713 ^ v_712;
assign v_719 = v_453 ^ ~v_583;
assign v_720 = v_719 ^ v_718;
assign v_725 = v_454 ^ ~v_585;
assign v_726 = v_725 ^ v_724;
assign v_731 = v_455 ^ ~v_587;
assign v_732 = v_731 ^ v_730;
assign v_737 = v_456 ^ ~v_589;
assign v_738 = v_737 ^ v_736;
assign v_743 = v_457 ^ ~v_591;
assign v_744 = v_743 ^ v_742;
assign v_749 = v_458 ^ ~v_593;
assign v_750 = v_749 ^ v_748;
assign v_755 = v_459 ^ ~v_595;
assign v_756 = v_755 ^ v_754;
assign v_761 = v_460 ^ ~v_597;
assign v_762 = v_761 ^ v_760;
assign v_767 = v_461 ^ ~v_599;
assign v_768 = v_767 ^ v_766;
assign v_773 = v_462 ^ ~v_601;
assign v_774 = v_773 ^ v_772;
assign v_779 = v_463 ^ ~v_603;
assign v_780 = v_779 ^ v_778;
assign v_785 = v_464 ^ ~v_605;
assign v_786 = v_785 ^ v_784;
assign v_791 = v_465 ^ ~v_607;
assign v_792 = v_791 ^ v_790;
assign v_797 = v_466 ^ ~v_609;
assign v_798 = v_797 ^ v_796;
assign v_803 = v_467 ^ ~v_611;
assign v_804 = v_803 ^ v_802;
assign v_809 = v_468 ^ ~v_613;
assign v_810 = v_809 ^ v_808;
assign v_815 = v_469 ^ ~v_615;
assign v_816 = v_815 ^ v_814;
assign v_821 = v_470 ^ ~v_617;
assign v_822 = v_821 ^ v_820;
assign v_827 = v_471 ^ ~v_619;
assign v_828 = v_827 ^ v_826;
assign v_833 = v_472 ^ ~v_621;
assign v_834 = v_833 ^ v_832;
assign v_839 = v_473 ^ ~v_623;
assign v_840 = v_839 ^ v_838;
assign v_845 = v_474 ^ ~v_625;
assign v_846 = v_845 ^ v_844;
assign v_851 = v_475 ^ ~v_627;
assign v_852 = v_851 ^ v_850;
assign v_857 = v_476 ^ ~v_629;
assign v_858 = v_857 ^ v_856;
assign v_863 = v_477 ^ ~v_631;
assign v_864 = v_863 ^ v_862;
assign v_869 = v_478 ^ ~v_633;
assign v_870 = v_869 ^ v_868;
assign v_875 = v_479 ^ ~v_635;
assign v_876 = v_875 ^ v_874;
assign v_881 = v_480 ^ ~v_637;
assign v_882 = v_881 ^ v_880;
assign v_887 = v_481 ^ ~v_639;
assign v_888 = v_887 ^ v_886;
assign v_893 = v_482 ^ ~v_641;
assign v_894 = v_893 ^ v_892;
assign v_899 = v_483 ^ ~v_643;
assign v_900 = v_899 ^ v_898;
assign v_905 = v_484 ^ ~v_645;
assign v_906 = v_905 ^ v_904;
assign v_911 = v_485 ^ ~v_647;
assign v_912 = v_911 ^ v_910;
assign v_917 = v_486 ^ ~v_649;
assign v_918 = v_917 ^ v_916;
assign v_923 = v_487 ^ ~v_651;
assign v_924 = v_923 ^ v_922;
assign v_929 = v_488 ^ ~v_653;
assign v_930 = v_929 ^ v_928;
assign v_935 = v_489 ^ ~v_655;
assign v_936 = v_935 ^ v_934;
assign v_941 = v_490 ^ ~v_657;
assign v_942 = v_941 ^ v_940;
assign v_947 = v_491 ^ ~v_659;
assign v_948 = v_947 ^ v_946;
assign v_953 = v_492 ^ ~v_661;
assign v_954 = v_953 ^ v_952;
assign v_959 = v_493 ^ ~v_663;
assign v_960 = v_959 ^ v_958;
assign v_965 = v_494 ^ ~v_665;
assign v_966 = v_965 ^ v_964;
assign v_971 = v_495 ^ ~v_667;
assign v_972 = v_971 ^ v_970;
assign v_977 = v_496 ^ ~v_669;
assign v_978 = v_977 ^ v_976;
assign v_983 = v_497 ^ ~v_671;
assign v_984 = v_983 ^ v_982;
assign v_989 = v_498 ^ ~v_673;
assign v_990 = v_989 ^ v_988;
assign v_995 = v_499 ^ ~v_675;
assign v_996 = v_995 ^ v_994;
assign v_1001 = v_500 ^ ~v_677;
assign v_1002 = v_1001 ^ v_1000;
assign v_1007 = v_501 ^ ~v_679;
assign v_1008 = v_1007 ^ v_1006;
assign v_1013 = v_502 ^ ~v_681;
assign v_1014 = v_1013 ^ v_1012;
assign v_1019 = v_503 ^ ~v_683;
assign v_1020 = v_1019 ^ v_1018;
assign v_1025 = v_504 ^ ~v_685;
assign v_1026 = v_1025 ^ v_1024;
assign v_1031 = v_505 ^ ~v_687;
assign v_1032 = v_1031 ^ v_1030;
assign v_1037 = v_506 ^ ~v_689;
assign v_1038 = v_1037 ^ v_1036;
assign v_1043 = v_507 ^ ~v_691;
assign v_1044 = v_1043 ^ v_1042;
assign v_1049 = v_508 ^ ~v_693;
assign v_1050 = v_1049 ^ v_1048;
assign v_1055 = v_509 ^ ~v_695;
assign v_1056 = v_1055 ^ v_1054;
assign v_1061 = v_510 ^ ~v_697;
assign v_1062 = v_1061 ^ v_1060;
assign v_1067 = v_511 ^ ~v_699;
assign v_1068 = v_1067 ^ v_1066;
assign v_1073 = v_512 ^ ~v_701;
assign v_1074 = v_1073 ^ v_1072;
assign v_1079 = v_513 ^ ~v_703;
assign v_1080 = v_1079 ^ v_1078;
assign v_1282 = v_1218 ^ v_385;
assign v_1283 = v_1219 ^ v_386;
assign v_1284 = v_1220 ^ v_387;
assign v_1285 = v_1221 ^ v_388;
assign v_1286 = v_1222 ^ v_389;
assign v_1287 = v_1223 ^ v_390;
assign v_1288 = v_1224 ^ v_391;
assign v_1289 = v_1225 ^ v_392;
assign v_1290 = v_1226 ^ v_393;
assign v_1291 = v_1227 ^ v_394;
assign v_1292 = v_1228 ^ v_395;
assign v_1293 = v_1229 ^ v_396;
assign v_1294 = v_1230 ^ v_397;
assign v_1295 = v_1231 ^ v_398;
assign v_1296 = v_1232 ^ v_399;
assign v_1297 = v_1233 ^ v_400;
assign v_1298 = v_1234 ^ v_401;
assign v_1299 = v_1235 ^ v_402;
assign v_1300 = v_1236 ^ v_403;
assign v_1301 = v_1237 ^ v_404;
assign v_1302 = v_1238 ^ v_405;
assign v_1303 = v_1239 ^ v_406;
assign v_1304 = v_1240 ^ v_407;
assign v_1305 = v_1241 ^ v_408;
assign v_1306 = v_1242 ^ v_409;
assign v_1307 = v_1243 ^ v_410;
assign v_1308 = v_1244 ^ v_411;
assign v_1309 = v_1245 ^ v_412;
assign v_1310 = v_1246 ^ v_413;
assign v_1311 = v_1247 ^ v_414;
assign v_1312 = v_1248 ^ v_415;
assign v_1313 = v_1249 ^ v_416;
assign v_1314 = v_1250 ^ v_417;
assign v_1315 = v_1251 ^ v_418;
assign v_1316 = v_1252 ^ v_419;
assign v_1317 = v_1253 ^ v_420;
assign v_1318 = v_1254 ^ v_421;
assign v_1319 = v_1255 ^ v_422;
assign v_1320 = v_1256 ^ v_423;
assign v_1321 = v_1257 ^ v_424;
assign v_1322 = v_1258 ^ v_425;
assign v_1323 = v_1259 ^ v_426;
assign v_1324 = v_1260 ^ v_427;
assign v_1325 = v_1261 ^ v_428;
assign v_1326 = v_1262 ^ v_429;
assign v_1327 = v_1263 ^ v_430;
assign v_1328 = v_1264 ^ v_431;
assign v_1329 = v_1265 ^ v_432;
assign v_1330 = v_1266 ^ v_433;
assign v_1331 = v_1267 ^ v_434;
assign v_1332 = v_1268 ^ v_435;
assign v_1333 = v_1269 ^ v_436;
assign v_1334 = v_1270 ^ v_437;
assign v_1335 = v_1271 ^ v_438;
assign v_1336 = v_1272 ^ v_439;
assign v_1337 = v_1273 ^ v_440;
assign v_1338 = v_1274 ^ v_441;
assign v_1339 = v_1275 ^ v_442;
assign v_1340 = v_1276 ^ v_443;
assign v_1341 = v_1277 ^ v_444;
assign v_1342 = v_1278 ^ v_445;
assign v_1343 = v_1279 ^ v_446;
assign v_1344 = v_1280 ^ v_447;
assign v_1345 = v_1281 ^ v_448;
assign v_1411 = v_1347 ^ v_450;
assign v_1412 = v_1348 ^ v_451;
assign v_1413 = v_1349 ^ v_452;
assign v_1414 = v_1350 ^ v_453;
assign v_1415 = v_1351 ^ v_454;
assign v_1416 = v_1352 ^ v_455;
assign v_1417 = v_1353 ^ v_456;
assign v_1418 = v_1354 ^ v_457;
assign v_1419 = v_1355 ^ v_458;
assign v_1420 = v_1356 ^ v_459;
assign v_1421 = v_1357 ^ v_460;
assign v_1422 = v_1358 ^ v_461;
assign v_1423 = v_1359 ^ v_462;
assign v_1424 = v_1360 ^ v_463;
assign v_1425 = v_1361 ^ v_464;
assign v_1426 = v_1362 ^ v_465;
assign v_1427 = v_1363 ^ v_466;
assign v_1428 = v_1364 ^ v_467;
assign v_1429 = v_1365 ^ v_468;
assign v_1430 = v_1366 ^ v_469;
assign v_1431 = v_1367 ^ v_470;
assign v_1432 = v_1368 ^ v_471;
assign v_1433 = v_1369 ^ v_472;
assign v_1434 = v_1370 ^ v_473;
assign v_1435 = v_1371 ^ v_474;
assign v_1436 = v_1372 ^ v_475;
assign v_1437 = v_1373 ^ v_476;
assign v_1438 = v_1374 ^ v_477;
assign v_1439 = v_1375 ^ v_478;
assign v_1440 = v_1376 ^ v_479;
assign v_1441 = v_1377 ^ v_480;
assign v_1442 = v_1378 ^ v_481;
assign v_1443 = v_1379 ^ v_482;
assign v_1444 = v_1380 ^ v_483;
assign v_1445 = v_1381 ^ v_484;
assign v_1446 = v_1382 ^ v_485;
assign v_1447 = v_1383 ^ v_486;
assign v_1448 = v_1384 ^ v_487;
assign v_1449 = v_1385 ^ v_488;
assign v_1450 = v_1386 ^ v_489;
assign v_1451 = v_1387 ^ v_490;
assign v_1452 = v_1388 ^ v_491;
assign v_1453 = v_1389 ^ v_492;
assign v_1454 = v_1390 ^ v_493;
assign v_1455 = v_1391 ^ v_494;
assign v_1456 = v_1392 ^ v_495;
assign v_1457 = v_1393 ^ v_496;
assign v_1458 = v_1394 ^ v_497;
assign v_1459 = v_1395 ^ v_498;
assign v_1460 = v_1396 ^ v_499;
assign v_1461 = v_1397 ^ v_500;
assign v_1462 = v_1398 ^ v_501;
assign v_1463 = v_1399 ^ v_502;
assign v_1464 = v_1400 ^ v_503;
assign v_1465 = v_1401 ^ v_504;
assign v_1466 = v_1402 ^ v_505;
assign v_1467 = v_1403 ^ v_506;
assign v_1468 = v_1404 ^ v_507;
assign v_1469 = v_1405 ^ v_508;
assign v_1470 = v_1406 ^ v_509;
assign v_1471 = v_1407 ^ v_510;
assign v_1472 = v_1408 ^ v_511;
assign v_1473 = v_1409 ^ v_512;
assign v_1474 = v_1410 ^ v_513;
assign v_1540 = v_1476 ^ v_514;
assign v_1541 = v_1477 ^ v_515;
assign v_1542 = v_1478 ^ v_516;
assign v_1543 = v_1479 ^ v_517;
assign v_1544 = v_1480 ^ v_518;
assign v_1545 = v_1481 ^ v_519;
assign v_1546 = v_1482 ^ v_520;
assign v_1547 = v_1483 ^ v_521;
assign v_1548 = v_1484 ^ v_522;
assign v_1549 = v_1485 ^ v_523;
assign v_1550 = v_1486 ^ v_524;
assign v_1551 = v_1487 ^ v_525;
assign v_1552 = v_1488 ^ v_526;
assign v_1553 = v_1489 ^ v_527;
assign v_1554 = v_1490 ^ v_528;
assign v_1555 = v_1491 ^ v_529;
assign v_1556 = v_1492 ^ v_530;
assign v_1557 = v_1493 ^ v_531;
assign v_1558 = v_1494 ^ v_532;
assign v_1559 = v_1495 ^ v_533;
assign v_1560 = v_1496 ^ v_534;
assign v_1561 = v_1497 ^ v_535;
assign v_1562 = v_1498 ^ v_536;
assign v_1563 = v_1499 ^ v_537;
assign v_1564 = v_1500 ^ v_538;
assign v_1565 = v_1501 ^ v_539;
assign v_1566 = v_1502 ^ v_540;
assign v_1567 = v_1503 ^ v_541;
assign v_1568 = v_1504 ^ v_542;
assign v_1569 = v_1505 ^ v_543;
assign v_1570 = v_1506 ^ v_544;
assign v_1571 = v_1507 ^ v_545;
assign v_1572 = v_1508 ^ v_546;
assign v_1573 = v_1509 ^ v_547;
assign v_1574 = v_1510 ^ v_548;
assign v_1575 = v_1511 ^ v_549;
assign v_1576 = v_1512 ^ v_550;
assign v_1577 = v_1513 ^ v_551;
assign v_1578 = v_1514 ^ v_552;
assign v_1579 = v_1515 ^ v_553;
assign v_1580 = v_1516 ^ v_554;
assign v_1581 = v_1517 ^ v_555;
assign v_1582 = v_1518 ^ v_556;
assign v_1583 = v_1519 ^ v_557;
assign v_1584 = v_1520 ^ v_558;
assign v_1585 = v_1521 ^ v_559;
assign v_1586 = v_1522 ^ v_560;
assign v_1587 = v_1523 ^ v_561;
assign v_1588 = v_1524 ^ v_562;
assign v_1589 = v_1525 ^ v_563;
assign v_1590 = v_1526 ^ v_564;
assign v_1591 = v_1527 ^ v_565;
assign v_1592 = v_1528 ^ v_566;
assign v_1593 = v_1529 ^ v_567;
assign v_1594 = v_1530 ^ v_568;
assign v_1595 = v_1531 ^ v_569;
assign v_1596 = v_1532 ^ v_570;
assign v_1597 = v_1533 ^ v_571;
assign v_1598 = v_1534 ^ v_572;
assign v_1599 = v_1535 ^ v_573;
assign v_1600 = v_1536 ^ v_574;
assign v_1601 = v_1537 ^ v_575;
assign v_1602 = v_1538 ^ v_576;
assign v_1603 = v_1539 ^ v_577;
assign v_1605 = v_1 ^ v_1476;
assign v_1606 = v_2 ^ v_1477;
assign v_1607 = v_3 ^ v_1478;
assign v_1608 = v_4 ^ v_1479;
assign v_1609 = v_5 ^ v_1480;
assign v_1610 = v_6 ^ v_1481;
assign v_1611 = v_7 ^ v_1482;
assign v_1612 = v_8 ^ v_1483;
assign v_1613 = v_9 ^ v_1484;
assign v_1614 = v_10 ^ v_1485;
assign v_1615 = v_11 ^ v_1486;
assign v_1616 = v_12 ^ v_1487;
assign v_1617 = v_13 ^ v_1488;
assign v_1618 = v_14 ^ v_1489;
assign v_1619 = v_15 ^ v_1490;
assign v_1620 = v_16 ^ v_1491;
assign v_1621 = v_17 ^ v_1492;
assign v_1622 = v_18 ^ v_1493;
assign v_1623 = v_19 ^ v_1494;
assign v_1624 = v_20 ^ v_1495;
assign v_1625 = v_21 ^ v_1496;
assign v_1626 = v_22 ^ v_1497;
assign v_1627 = v_23 ^ v_1498;
assign v_1628 = v_24 ^ v_1499;
assign v_1629 = v_25 ^ v_1500;
assign v_1630 = v_26 ^ v_1501;
assign v_1631 = v_27 ^ v_1502;
assign v_1632 = v_28 ^ v_1503;
assign v_1633 = v_29 ^ v_1504;
assign v_1634 = v_30 ^ v_1505;
assign v_1635 = v_31 ^ v_1506;
assign v_1636 = v_32 ^ v_1507;
assign v_1637 = v_33 ^ v_1508;
assign v_1638 = v_34 ^ v_1509;
assign v_1639 = v_35 ^ v_1510;
assign v_1640 = v_36 ^ v_1511;
assign v_1641 = v_37 ^ v_1512;
assign v_1642 = v_38 ^ v_1513;
assign v_1643 = v_39 ^ v_1514;
assign v_1644 = v_40 ^ v_1515;
assign v_1645 = v_41 ^ v_1516;
assign v_1646 = v_42 ^ v_1517;
assign v_1647 = v_43 ^ v_1518;
assign v_1648 = v_44 ^ v_1519;
assign v_1649 = v_45 ^ v_1520;
assign v_1650 = v_46 ^ v_1521;
assign v_1651 = v_47 ^ v_1522;
assign v_1652 = v_48 ^ v_1523;
assign v_1653 = v_49 ^ v_1524;
assign v_1654 = v_50 ^ v_1525;
assign v_1655 = v_51 ^ v_1526;
assign v_1656 = v_52 ^ v_1527;
assign v_1657 = v_53 ^ v_1528;
assign v_1658 = v_54 ^ v_1529;
assign v_1659 = v_55 ^ v_1530;
assign v_1660 = v_56 ^ v_1531;
assign v_1661 = v_57 ^ v_1532;
assign v_1662 = v_58 ^ v_1533;
assign v_1663 = v_59 ^ v_1534;
assign v_1664 = v_60 ^ v_1535;
assign v_1665 = v_61 ^ v_1536;
assign v_1666 = v_62 ^ v_1537;
assign v_1667 = v_63 ^ v_1538;
assign v_1668 = v_64 ^ v_1539;
assign v_1670 = v_514 ^ v_450;
assign v_1673 = v_515 ^ v_451;
assign v_1674 = v_1673 ^ v_1672;
assign v_1679 = v_516 ^ v_452;
assign v_1680 = v_1679 ^ v_1678;
assign v_1685 = v_517 ^ v_453;
assign v_1686 = v_1685 ^ v_1684;
assign v_1691 = v_518 ^ v_454;
assign v_1692 = v_1691 ^ v_1690;
assign v_1697 = v_519 ^ v_455;
assign v_1698 = v_1697 ^ v_1696;
assign v_1703 = v_520 ^ v_456;
assign v_1704 = v_1703 ^ v_1702;
assign v_1709 = v_521 ^ v_457;
assign v_1710 = v_1709 ^ v_1708;
assign v_1715 = v_522 ^ v_458;
assign v_1716 = v_1715 ^ v_1714;
assign v_1721 = v_523 ^ v_459;
assign v_1722 = v_1721 ^ v_1720;
assign v_1727 = v_524 ^ v_460;
assign v_1728 = v_1727 ^ v_1726;
assign v_1733 = v_525 ^ v_461;
assign v_1734 = v_1733 ^ v_1732;
assign v_1739 = v_526 ^ v_462;
assign v_1740 = v_1739 ^ v_1738;
assign v_1745 = v_527 ^ v_463;
assign v_1746 = v_1745 ^ v_1744;
assign v_1751 = v_528 ^ v_464;
assign v_1752 = v_1751 ^ v_1750;
assign v_1757 = v_529 ^ v_465;
assign v_1758 = v_1757 ^ v_1756;
assign v_1763 = v_530 ^ v_466;
assign v_1764 = v_1763 ^ v_1762;
assign v_1769 = v_531 ^ v_467;
assign v_1770 = v_1769 ^ v_1768;
assign v_1775 = v_532 ^ v_468;
assign v_1776 = v_1775 ^ v_1774;
assign v_1781 = v_533 ^ v_469;
assign v_1782 = v_1781 ^ v_1780;
assign v_1787 = v_534 ^ v_470;
assign v_1788 = v_1787 ^ v_1786;
assign v_1793 = v_535 ^ v_471;
assign v_1794 = v_1793 ^ v_1792;
assign v_1799 = v_536 ^ v_472;
assign v_1800 = v_1799 ^ v_1798;
assign v_1805 = v_537 ^ v_473;
assign v_1806 = v_1805 ^ v_1804;
assign v_1811 = v_538 ^ v_474;
assign v_1812 = v_1811 ^ v_1810;
assign v_1817 = v_539 ^ v_475;
assign v_1818 = v_1817 ^ v_1816;
assign v_1823 = v_540 ^ v_476;
assign v_1824 = v_1823 ^ v_1822;
assign v_1829 = v_541 ^ v_477;
assign v_1830 = v_1829 ^ v_1828;
assign v_1835 = v_542 ^ v_478;
assign v_1836 = v_1835 ^ v_1834;
assign v_1841 = v_543 ^ v_479;
assign v_1842 = v_1841 ^ v_1840;
assign v_1847 = v_544 ^ v_480;
assign v_1848 = v_1847 ^ v_1846;
assign v_1853 = v_545 ^ v_481;
assign v_1854 = v_1853 ^ v_1852;
assign v_1859 = v_546 ^ v_482;
assign v_1860 = v_1859 ^ v_1858;
assign v_1865 = v_547 ^ v_483;
assign v_1866 = v_1865 ^ v_1864;
assign v_1871 = v_548 ^ v_484;
assign v_1872 = v_1871 ^ v_1870;
assign v_1877 = v_549 ^ v_485;
assign v_1878 = v_1877 ^ v_1876;
assign v_1883 = v_550 ^ v_486;
assign v_1884 = v_1883 ^ v_1882;
assign v_1889 = v_551 ^ v_487;
assign v_1890 = v_1889 ^ v_1888;
assign v_1895 = v_552 ^ v_488;
assign v_1896 = v_1895 ^ v_1894;
assign v_1901 = v_553 ^ v_489;
assign v_1902 = v_1901 ^ v_1900;
assign v_1907 = v_554 ^ v_490;
assign v_1908 = v_1907 ^ v_1906;
assign v_1913 = v_555 ^ v_491;
assign v_1914 = v_1913 ^ v_1912;
assign v_1919 = v_556 ^ v_492;
assign v_1920 = v_1919 ^ v_1918;
assign v_1925 = v_557 ^ v_493;
assign v_1926 = v_1925 ^ v_1924;
assign v_1931 = v_558 ^ v_494;
assign v_1932 = v_1931 ^ v_1930;
assign v_1937 = v_559 ^ v_495;
assign v_1938 = v_1937 ^ v_1936;
assign v_1943 = v_560 ^ v_496;
assign v_1944 = v_1943 ^ v_1942;
assign v_1949 = v_561 ^ v_497;
assign v_1950 = v_1949 ^ v_1948;
assign v_1955 = v_562 ^ v_498;
assign v_1956 = v_1955 ^ v_1954;
assign v_1961 = v_563 ^ v_499;
assign v_1962 = v_1961 ^ v_1960;
assign v_1967 = v_564 ^ v_500;
assign v_1968 = v_1967 ^ v_1966;
assign v_1973 = v_565 ^ v_501;
assign v_1974 = v_1973 ^ v_1972;
assign v_1979 = v_566 ^ v_502;
assign v_1980 = v_1979 ^ v_1978;
assign v_1985 = v_567 ^ v_503;
assign v_1986 = v_1985 ^ v_1984;
assign v_1991 = v_568 ^ v_504;
assign v_1992 = v_1991 ^ v_1990;
assign v_1997 = v_569 ^ v_505;
assign v_1998 = v_1997 ^ v_1996;
assign v_2003 = v_570 ^ v_506;
assign v_2004 = v_2003 ^ v_2002;
assign v_2009 = v_571 ^ v_507;
assign v_2010 = v_2009 ^ v_2008;
assign v_2015 = v_572 ^ v_508;
assign v_2016 = v_2015 ^ v_2014;
assign v_2021 = v_573 ^ v_509;
assign v_2022 = v_2021 ^ v_2020;
assign v_2027 = v_574 ^ v_510;
assign v_2028 = v_2027 ^ v_2026;
assign v_2033 = v_575 ^ v_511;
assign v_2034 = v_2033 ^ v_2032;
assign v_2039 = v_576 ^ v_512;
assign v_2040 = v_2039 ^ v_2038;
assign v_2045 = v_577 ^ v_513;
assign v_2046 = v_2045 ^ v_2044;
assign v_2051 = v_193 ^ v_1670;
assign v_2052 = v_194 ^ v_1674;
assign v_2053 = v_195 ^ v_1680;
assign v_2054 = v_196 ^ v_1686;
assign v_2055 = v_197 ^ v_1692;
assign v_2056 = v_198 ^ v_1698;
assign v_2057 = v_199 ^ v_1704;
assign v_2058 = v_200 ^ v_1710;
assign v_2059 = v_201 ^ v_1716;
assign v_2060 = v_202 ^ v_1722;
assign v_2061 = v_203 ^ v_1728;
assign v_2062 = v_204 ^ v_1734;
assign v_2063 = v_205 ^ v_1740;
assign v_2064 = v_206 ^ v_1746;
assign v_2065 = v_207 ^ v_1752;
assign v_2066 = v_208 ^ v_1758;
assign v_2067 = v_209 ^ v_1764;
assign v_2068 = v_210 ^ v_1770;
assign v_2069 = v_211 ^ v_1776;
assign v_2070 = v_212 ^ v_1782;
assign v_2071 = v_213 ^ v_1788;
assign v_2072 = v_214 ^ v_1794;
assign v_2073 = v_215 ^ v_1800;
assign v_2074 = v_216 ^ v_1806;
assign v_2075 = v_217 ^ v_1812;
assign v_2076 = v_218 ^ v_1818;
assign v_2077 = v_219 ^ v_1824;
assign v_2078 = v_220 ^ v_1830;
assign v_2079 = v_221 ^ v_1836;
assign v_2080 = v_222 ^ v_1842;
assign v_2081 = v_223 ^ v_1848;
assign v_2082 = v_224 ^ v_1854;
assign v_2083 = v_225 ^ v_1860;
assign v_2084 = v_226 ^ v_1866;
assign v_2085 = v_227 ^ v_1872;
assign v_2086 = v_228 ^ v_1878;
assign v_2087 = v_229 ^ v_1884;
assign v_2088 = v_230 ^ v_1890;
assign v_2089 = v_231 ^ v_1896;
assign v_2090 = v_232 ^ v_1902;
assign v_2091 = v_233 ^ v_1908;
assign v_2092 = v_234 ^ v_1914;
assign v_2093 = v_235 ^ v_1920;
assign v_2094 = v_236 ^ v_1926;
assign v_2095 = v_237 ^ v_1932;
assign v_2096 = v_238 ^ v_1938;
assign v_2097 = v_239 ^ v_1944;
assign v_2098 = v_240 ^ v_1950;
assign v_2099 = v_241 ^ v_1956;
assign v_2100 = v_242 ^ v_1962;
assign v_2101 = v_243 ^ v_1968;
assign v_2102 = v_244 ^ v_1974;
assign v_2103 = v_245 ^ v_1980;
assign v_2104 = v_246 ^ v_1986;
assign v_2105 = v_247 ^ v_1992;
assign v_2106 = v_248 ^ v_1998;
assign v_2107 = v_249 ^ v_2004;
assign v_2108 = v_250 ^ v_2010;
assign v_2109 = v_251 ^ v_2016;
assign v_2110 = v_252 ^ v_2022;
assign v_2111 = v_253 ^ v_2028;
assign v_2112 = v_254 ^ v_2034;
assign v_2113 = v_255 ^ v_2040;
assign v_2114 = v_256 ^ v_2046;
assign v_2116 = v_65 ^ v_1347;
assign v_2117 = v_66 ^ v_1348;
assign v_2118 = v_67 ^ v_1349;
assign v_2119 = v_68 ^ v_1350;
assign v_2120 = v_69 ^ v_1351;
assign v_2121 = v_70 ^ v_1352;
assign v_2122 = v_71 ^ v_1353;
assign v_2123 = v_72 ^ v_1354;
assign v_2124 = v_73 ^ v_1355;
assign v_2125 = v_74 ^ v_1356;
assign v_2126 = v_75 ^ v_1357;
assign v_2127 = v_76 ^ v_1358;
assign v_2128 = v_77 ^ v_1359;
assign v_2129 = v_78 ^ v_1360;
assign v_2130 = v_79 ^ v_1361;
assign v_2131 = v_80 ^ v_1362;
assign v_2132 = v_81 ^ v_1363;
assign v_2133 = v_82 ^ v_1364;
assign v_2134 = v_83 ^ v_1365;
assign v_2135 = v_84 ^ v_1366;
assign v_2136 = v_85 ^ v_1367;
assign v_2137 = v_86 ^ v_1368;
assign v_2138 = v_87 ^ v_1369;
assign v_2139 = v_88 ^ v_1370;
assign v_2140 = v_89 ^ v_1371;
assign v_2141 = v_90 ^ v_1372;
assign v_2142 = v_91 ^ v_1373;
assign v_2143 = v_92 ^ v_1374;
assign v_2144 = v_93 ^ v_1375;
assign v_2145 = v_94 ^ v_1376;
assign v_2146 = v_95 ^ v_1377;
assign v_2147 = v_96 ^ v_1378;
assign v_2148 = v_97 ^ v_1379;
assign v_2149 = v_98 ^ v_1380;
assign v_2150 = v_99 ^ v_1381;
assign v_2151 = v_100 ^ v_1382;
assign v_2152 = v_101 ^ v_1383;
assign v_2153 = v_102 ^ v_1384;
assign v_2154 = v_103 ^ v_1385;
assign v_2155 = v_104 ^ v_1386;
assign v_2156 = v_105 ^ v_1387;
assign v_2157 = v_106 ^ v_1388;
assign v_2158 = v_107 ^ v_1389;
assign v_2159 = v_108 ^ v_1390;
assign v_2160 = v_109 ^ v_1391;
assign v_2161 = v_110 ^ v_1392;
assign v_2162 = v_111 ^ v_1393;
assign v_2163 = v_112 ^ v_1394;
assign v_2164 = v_113 ^ v_1395;
assign v_2165 = v_114 ^ v_1396;
assign v_2166 = v_115 ^ v_1397;
assign v_2167 = v_116 ^ v_1398;
assign v_2168 = v_117 ^ v_1399;
assign v_2169 = v_118 ^ v_1400;
assign v_2170 = v_119 ^ v_1401;
assign v_2171 = v_120 ^ v_1402;
assign v_2172 = v_121 ^ v_1403;
assign v_2173 = v_122 ^ v_1404;
assign v_2174 = v_123 ^ v_1405;
assign v_2175 = v_124 ^ v_1406;
assign v_2176 = v_125 ^ v_1407;
assign v_2177 = v_126 ^ v_1408;
assign v_2178 = v_127 ^ v_1409;
assign v_2179 = v_128 ^ v_1410;
assign v_2181 = v_450 ^ v_385;
assign v_2184 = v_451 ^ v_386;
assign v_2185 = v_2184 ^ v_2183;
assign v_2190 = v_452 ^ v_387;
assign v_2191 = v_2190 ^ v_2189;
assign v_2196 = v_453 ^ v_388;
assign v_2197 = v_2196 ^ v_2195;
assign v_2202 = v_454 ^ v_389;
assign v_2203 = v_2202 ^ v_2201;
assign v_2208 = v_455 ^ v_390;
assign v_2209 = v_2208 ^ v_2207;
assign v_2214 = v_456 ^ v_391;
assign v_2215 = v_2214 ^ v_2213;
assign v_2220 = v_457 ^ v_392;
assign v_2221 = v_2220 ^ v_2219;
assign v_2226 = v_458 ^ v_393;
assign v_2227 = v_2226 ^ v_2225;
assign v_2232 = v_459 ^ v_394;
assign v_2233 = v_2232 ^ v_2231;
assign v_2238 = v_460 ^ v_395;
assign v_2239 = v_2238 ^ v_2237;
assign v_2244 = v_461 ^ v_396;
assign v_2245 = v_2244 ^ v_2243;
assign v_2250 = v_462 ^ v_397;
assign v_2251 = v_2250 ^ v_2249;
assign v_2256 = v_463 ^ v_398;
assign v_2257 = v_2256 ^ v_2255;
assign v_2262 = v_464 ^ v_399;
assign v_2263 = v_2262 ^ v_2261;
assign v_2268 = v_465 ^ v_400;
assign v_2269 = v_2268 ^ v_2267;
assign v_2274 = v_466 ^ v_401;
assign v_2275 = v_2274 ^ v_2273;
assign v_2280 = v_467 ^ v_402;
assign v_2281 = v_2280 ^ v_2279;
assign v_2286 = v_468 ^ v_403;
assign v_2287 = v_2286 ^ v_2285;
assign v_2292 = v_469 ^ v_404;
assign v_2293 = v_2292 ^ v_2291;
assign v_2298 = v_470 ^ v_405;
assign v_2299 = v_2298 ^ v_2297;
assign v_2304 = v_471 ^ v_406;
assign v_2305 = v_2304 ^ v_2303;
assign v_2310 = v_472 ^ v_407;
assign v_2311 = v_2310 ^ v_2309;
assign v_2316 = v_473 ^ v_408;
assign v_2317 = v_2316 ^ v_2315;
assign v_2322 = v_474 ^ v_409;
assign v_2323 = v_2322 ^ v_2321;
assign v_2328 = v_475 ^ v_410;
assign v_2329 = v_2328 ^ v_2327;
assign v_2334 = v_476 ^ v_411;
assign v_2335 = v_2334 ^ v_2333;
assign v_2340 = v_477 ^ v_412;
assign v_2341 = v_2340 ^ v_2339;
assign v_2346 = v_478 ^ v_413;
assign v_2347 = v_2346 ^ v_2345;
assign v_2352 = v_479 ^ v_414;
assign v_2353 = v_2352 ^ v_2351;
assign v_2358 = v_480 ^ v_415;
assign v_2359 = v_2358 ^ v_2357;
assign v_2364 = v_481 ^ v_416;
assign v_2365 = v_2364 ^ v_2363;
assign v_2370 = v_482 ^ v_417;
assign v_2371 = v_2370 ^ v_2369;
assign v_2376 = v_483 ^ v_418;
assign v_2377 = v_2376 ^ v_2375;
assign v_2382 = v_484 ^ v_419;
assign v_2383 = v_2382 ^ v_2381;
assign v_2388 = v_485 ^ v_420;
assign v_2389 = v_2388 ^ v_2387;
assign v_2394 = v_486 ^ v_421;
assign v_2395 = v_2394 ^ v_2393;
assign v_2400 = v_487 ^ v_422;
assign v_2401 = v_2400 ^ v_2399;
assign v_2406 = v_488 ^ v_423;
assign v_2407 = v_2406 ^ v_2405;
assign v_2412 = v_489 ^ v_424;
assign v_2413 = v_2412 ^ v_2411;
assign v_2418 = v_490 ^ v_425;
assign v_2419 = v_2418 ^ v_2417;
assign v_2424 = v_491 ^ v_426;
assign v_2425 = v_2424 ^ v_2423;
assign v_2430 = v_492 ^ v_427;
assign v_2431 = v_2430 ^ v_2429;
assign v_2436 = v_493 ^ v_428;
assign v_2437 = v_2436 ^ v_2435;
assign v_2442 = v_494 ^ v_429;
assign v_2443 = v_2442 ^ v_2441;
assign v_2448 = v_495 ^ v_430;
assign v_2449 = v_2448 ^ v_2447;
assign v_2454 = v_496 ^ v_431;
assign v_2455 = v_2454 ^ v_2453;
assign v_2460 = v_497 ^ v_432;
assign v_2461 = v_2460 ^ v_2459;
assign v_2466 = v_498 ^ v_433;
assign v_2467 = v_2466 ^ v_2465;
assign v_2472 = v_499 ^ v_434;
assign v_2473 = v_2472 ^ v_2471;
assign v_2478 = v_500 ^ v_435;
assign v_2479 = v_2478 ^ v_2477;
assign v_2484 = v_501 ^ v_436;
assign v_2485 = v_2484 ^ v_2483;
assign v_2490 = v_502 ^ v_437;
assign v_2491 = v_2490 ^ v_2489;
assign v_2496 = v_503 ^ v_438;
assign v_2497 = v_2496 ^ v_2495;
assign v_2502 = v_504 ^ v_439;
assign v_2503 = v_2502 ^ v_2501;
assign v_2508 = v_505 ^ v_440;
assign v_2509 = v_2508 ^ v_2507;
assign v_2514 = v_506 ^ v_441;
assign v_2515 = v_2514 ^ v_2513;
assign v_2520 = v_507 ^ v_442;
assign v_2521 = v_2520 ^ v_2519;
assign v_2526 = v_508 ^ v_443;
assign v_2527 = v_2526 ^ v_2525;
assign v_2532 = v_509 ^ v_444;
assign v_2533 = v_2532 ^ v_2531;
assign v_2538 = v_510 ^ v_445;
assign v_2539 = v_2538 ^ v_2537;
assign v_2544 = v_511 ^ v_446;
assign v_2545 = v_2544 ^ v_2543;
assign v_2550 = v_512 ^ v_447;
assign v_2551 = v_2550 ^ v_2549;
assign v_2556 = v_513 ^ v_448;
assign v_2557 = v_2556 ^ v_2555;
assign v_2562 = v_257 ^ v_2181;
assign v_2563 = v_258 ^ v_2185;
assign v_2564 = v_259 ^ v_2191;
assign v_2565 = v_260 ^ v_2197;
assign v_2566 = v_261 ^ v_2203;
assign v_2567 = v_262 ^ v_2209;
assign v_2568 = v_263 ^ v_2215;
assign v_2569 = v_264 ^ v_2221;
assign v_2570 = v_265 ^ v_2227;
assign v_2571 = v_266 ^ v_2233;
assign v_2572 = v_267 ^ v_2239;
assign v_2573 = v_268 ^ v_2245;
assign v_2574 = v_269 ^ v_2251;
assign v_2575 = v_270 ^ v_2257;
assign v_2576 = v_271 ^ v_2263;
assign v_2577 = v_272 ^ v_2269;
assign v_2578 = v_273 ^ v_2275;
assign v_2579 = v_274 ^ v_2281;
assign v_2580 = v_275 ^ v_2287;
assign v_2581 = v_276 ^ v_2293;
assign v_2582 = v_277 ^ v_2299;
assign v_2583 = v_278 ^ v_2305;
assign v_2584 = v_279 ^ v_2311;
assign v_2585 = v_280 ^ v_2317;
assign v_2586 = v_281 ^ v_2323;
assign v_2587 = v_282 ^ v_2329;
assign v_2588 = v_283 ^ v_2335;
assign v_2589 = v_284 ^ v_2341;
assign v_2590 = v_285 ^ v_2347;
assign v_2591 = v_286 ^ v_2353;
assign v_2592 = v_287 ^ v_2359;
assign v_2593 = v_288 ^ v_2365;
assign v_2594 = v_289 ^ v_2371;
assign v_2595 = v_290 ^ v_2377;
assign v_2596 = v_291 ^ v_2383;
assign v_2597 = v_292 ^ v_2389;
assign v_2598 = v_293 ^ v_2395;
assign v_2599 = v_294 ^ v_2401;
assign v_2600 = v_295 ^ v_2407;
assign v_2601 = v_296 ^ v_2413;
assign v_2602 = v_297 ^ v_2419;
assign v_2603 = v_298 ^ v_2425;
assign v_2604 = v_299 ^ v_2431;
assign v_2605 = v_300 ^ v_2437;
assign v_2606 = v_301 ^ v_2443;
assign v_2607 = v_302 ^ v_2449;
assign v_2608 = v_303 ^ v_2455;
assign v_2609 = v_304 ^ v_2461;
assign v_2610 = v_305 ^ v_2467;
assign v_2611 = v_306 ^ v_2473;
assign v_2612 = v_307 ^ v_2479;
assign v_2613 = v_308 ^ v_2485;
assign v_2614 = v_309 ^ v_2491;
assign v_2615 = v_310 ^ v_2497;
assign v_2616 = v_311 ^ v_2503;
assign v_2617 = v_312 ^ v_2509;
assign v_2618 = v_313 ^ v_2515;
assign v_2619 = v_314 ^ v_2521;
assign v_2620 = v_315 ^ v_2527;
assign v_2621 = v_316 ^ v_2533;
assign v_2622 = v_317 ^ v_2539;
assign v_2623 = v_318 ^ v_2545;
assign v_2624 = v_319 ^ v_2551;
assign v_2625 = v_320 ^ v_2557;
assign v_2627 = v_129 ^ v_1218;
assign v_2628 = v_130 ^ v_1219;
assign v_2629 = v_131 ^ v_1220;
assign v_2630 = v_132 ^ v_1221;
assign v_2631 = v_133 ^ v_1222;
assign v_2632 = v_134 ^ v_1223;
assign v_2633 = v_135 ^ v_1224;
assign v_2634 = v_136 ^ v_1225;
assign v_2635 = v_137 ^ v_1226;
assign v_2636 = v_138 ^ v_1227;
assign v_2637 = v_139 ^ v_1228;
assign v_2638 = v_140 ^ v_1229;
assign v_2639 = v_141 ^ v_1230;
assign v_2640 = v_142 ^ v_1231;
assign v_2641 = v_143 ^ v_1232;
assign v_2642 = v_144 ^ v_1233;
assign v_2643 = v_145 ^ v_1234;
assign v_2644 = v_146 ^ v_1235;
assign v_2645 = v_147 ^ v_1236;
assign v_2646 = v_148 ^ v_1237;
assign v_2647 = v_149 ^ v_1238;
assign v_2648 = v_150 ^ v_1239;
assign v_2649 = v_151 ^ v_1240;
assign v_2650 = v_152 ^ v_1241;
assign v_2651 = v_153 ^ v_1242;
assign v_2652 = v_154 ^ v_1243;
assign v_2653 = v_155 ^ v_1244;
assign v_2654 = v_156 ^ v_1245;
assign v_2655 = v_157 ^ v_1246;
assign v_2656 = v_158 ^ v_1247;
assign v_2657 = v_159 ^ v_1248;
assign v_2658 = v_160 ^ v_1249;
assign v_2659 = v_161 ^ v_1250;
assign v_2660 = v_162 ^ v_1251;
assign v_2661 = v_163 ^ v_1252;
assign v_2662 = v_164 ^ v_1253;
assign v_2663 = v_165 ^ v_1254;
assign v_2664 = v_166 ^ v_1255;
assign v_2665 = v_167 ^ v_1256;
assign v_2666 = v_168 ^ v_1257;
assign v_2667 = v_169 ^ v_1258;
assign v_2668 = v_170 ^ v_1259;
assign v_2669 = v_171 ^ v_1260;
assign v_2670 = v_172 ^ v_1261;
assign v_2671 = v_173 ^ v_1262;
assign v_2672 = v_174 ^ v_1263;
assign v_2673 = v_175 ^ v_1264;
assign v_2674 = v_176 ^ v_1265;
assign v_2675 = v_177 ^ v_1266;
assign v_2676 = v_178 ^ v_1267;
assign v_2677 = v_179 ^ v_1268;
assign v_2678 = v_180 ^ v_1269;
assign v_2679 = v_181 ^ v_1270;
assign v_2680 = v_182 ^ v_1271;
assign v_2681 = v_183 ^ v_1272;
assign v_2682 = v_184 ^ v_1273;
assign v_2683 = v_185 ^ v_1274;
assign v_2684 = v_186 ^ v_1275;
assign v_2685 = v_187 ^ v_1276;
assign v_2686 = v_188 ^ v_1277;
assign v_2687 = v_189 ^ v_1278;
assign v_2688 = v_190 ^ v_1279;
assign v_2689 = v_191 ^ v_1280;
assign v_2690 = v_192 ^ v_1281;
assign v_2692 = v_321 ^ v_385;
assign v_2693 = v_322 ^ v_386;
assign v_2694 = v_323 ^ v_387;
assign v_2695 = v_324 ^ v_388;
assign v_2696 = v_325 ^ v_389;
assign v_2697 = v_326 ^ v_390;
assign v_2698 = v_327 ^ v_391;
assign v_2699 = v_328 ^ v_392;
assign v_2700 = v_329 ^ v_393;
assign v_2701 = v_330 ^ v_394;
assign v_2702 = v_331 ^ v_395;
assign v_2703 = v_332 ^ v_396;
assign v_2704 = v_333 ^ v_397;
assign v_2705 = v_334 ^ v_398;
assign v_2706 = v_335 ^ v_399;
assign v_2707 = v_336 ^ v_400;
assign v_2708 = v_337 ^ v_401;
assign v_2709 = v_338 ^ v_402;
assign v_2710 = v_339 ^ v_403;
assign v_2711 = v_340 ^ v_404;
assign v_2712 = v_341 ^ v_405;
assign v_2713 = v_342 ^ v_406;
assign v_2714 = v_343 ^ v_407;
assign v_2715 = v_344 ^ v_408;
assign v_2716 = v_345 ^ v_409;
assign v_2717 = v_346 ^ v_410;
assign v_2718 = v_347 ^ v_411;
assign v_2719 = v_348 ^ v_412;
assign v_2720 = v_349 ^ v_413;
assign v_2721 = v_350 ^ v_414;
assign v_2722 = v_351 ^ v_415;
assign v_2723 = v_352 ^ v_416;
assign v_2724 = v_353 ^ v_417;
assign v_2725 = v_354 ^ v_418;
assign v_2726 = v_355 ^ v_419;
assign v_2727 = v_356 ^ v_420;
assign v_2728 = v_357 ^ v_421;
assign v_2729 = v_358 ^ v_422;
assign v_2730 = v_359 ^ v_423;
assign v_2731 = v_360 ^ v_424;
assign v_2732 = v_361 ^ v_425;
assign v_2733 = v_362 ^ v_426;
assign v_2734 = v_363 ^ v_427;
assign v_2735 = v_364 ^ v_428;
assign v_2736 = v_365 ^ v_429;
assign v_2737 = v_366 ^ v_430;
assign v_2738 = v_367 ^ v_431;
assign v_2739 = v_368 ^ v_432;
assign v_2740 = v_369 ^ v_433;
assign v_2741 = v_370 ^ v_434;
assign v_2742 = v_371 ^ v_435;
assign v_2743 = v_372 ^ v_436;
assign v_2744 = v_373 ^ v_437;
assign v_2745 = v_374 ^ v_438;
assign v_2746 = v_375 ^ v_439;
assign v_2747 = v_376 ^ v_440;
assign v_2748 = v_377 ^ v_441;
assign v_2749 = v_378 ^ v_442;
assign v_2750 = v_379 ^ v_443;
assign v_2751 = v_380 ^ v_444;
assign v_2752 = v_381 ^ v_445;
assign v_2753 = v_382 ^ v_446;
assign v_2754 = v_383 ^ v_447;
assign v_2755 = v_384 ^ v_448;
assign v_3910 = v_1 ^ v_193;
assign v_3911 = v_2 ^ v_194;
assign v_3912 = v_3 ^ v_195;
assign v_3913 = v_4 ^ v_196;
assign v_3914 = v_5 ^ v_197;
assign v_3915 = v_6 ^ v_198;
assign v_3916 = v_7 ^ v_199;
assign v_3917 = v_8 ^ v_200;
assign v_3918 = v_9 ^ v_201;
assign v_3919 = v_10 ^ v_202;
assign v_3920 = v_11 ^ v_203;
assign v_3921 = v_12 ^ v_204;
assign v_3922 = v_13 ^ v_205;
assign v_3923 = v_14 ^ v_206;
assign v_3924 = v_15 ^ v_207;
assign v_3925 = v_16 ^ v_208;
assign v_3926 = v_17 ^ v_209;
assign v_3927 = v_18 ^ v_210;
assign v_3928 = v_19 ^ v_211;
assign v_3929 = v_20 ^ v_212;
assign v_3930 = v_21 ^ v_213;
assign v_3931 = v_22 ^ v_214;
assign v_3932 = v_23 ^ v_215;
assign v_3933 = v_24 ^ v_216;
assign v_3934 = v_25 ^ v_217;
assign v_3935 = v_26 ^ v_218;
assign v_3936 = v_27 ^ v_219;
assign v_3937 = v_28 ^ v_220;
assign v_3938 = v_29 ^ v_221;
assign v_3939 = v_30 ^ v_222;
assign v_3940 = v_31 ^ v_223;
assign v_3941 = v_32 ^ v_224;
assign v_3942 = v_33 ^ v_225;
assign v_3943 = v_34 ^ v_226;
assign v_3944 = v_35 ^ v_227;
assign v_3945 = v_36 ^ v_228;
assign v_3946 = v_37 ^ v_229;
assign v_3947 = v_38 ^ v_230;
assign v_3948 = v_39 ^ v_231;
assign v_3949 = v_40 ^ v_232;
assign v_3950 = v_41 ^ v_233;
assign v_3951 = v_42 ^ v_234;
assign v_3952 = v_43 ^ v_235;
assign v_3953 = v_44 ^ v_236;
assign v_3954 = v_45 ^ v_237;
assign v_3955 = v_46 ^ v_238;
assign v_3956 = v_47 ^ v_239;
assign v_3957 = v_48 ^ v_240;
assign v_3958 = v_49 ^ v_241;
assign v_3959 = v_50 ^ v_242;
assign v_3960 = v_51 ^ v_243;
assign v_3961 = v_52 ^ v_244;
assign v_3962 = v_53 ^ v_245;
assign v_3963 = v_54 ^ v_246;
assign v_3964 = v_55 ^ v_247;
assign v_3965 = v_56 ^ v_248;
assign v_3966 = v_57 ^ v_249;
assign v_3967 = v_58 ^ v_250;
assign v_3968 = v_59 ^ v_251;
assign v_3969 = v_60 ^ v_252;
assign v_3970 = v_61 ^ v_253;
assign v_3971 = v_62 ^ v_254;
assign v_3972 = v_63 ^ v_255;
assign v_3973 = v_64 ^ v_256;
assign v_3975 = v_2757 ^ v_2821;
assign v_3976 = v_2758 ^ v_2822;
assign v_3977 = v_2759 ^ v_2823;
assign v_3978 = v_2760 ^ v_2824;
assign v_3979 = v_2761 ^ v_2825;
assign v_3980 = v_2762 ^ v_2826;
assign v_3981 = v_2763 ^ v_2827;
assign v_3982 = v_2764 ^ v_2828;
assign v_3983 = v_2765 ^ v_2829;
assign v_3984 = v_2766 ^ v_2830;
assign v_3985 = v_2767 ^ v_2831;
assign v_3986 = v_2768 ^ v_2832;
assign v_3987 = v_2769 ^ v_2833;
assign v_3988 = v_2770 ^ v_2834;
assign v_3989 = v_2771 ^ v_2835;
assign v_3990 = v_2772 ^ v_2836;
assign v_3991 = v_2773 ^ v_2837;
assign v_3992 = v_2774 ^ v_2838;
assign v_3993 = v_2775 ^ v_2839;
assign v_3994 = v_2776 ^ v_2840;
assign v_3995 = v_2777 ^ v_2841;
assign v_3996 = v_2778 ^ v_2842;
assign v_3997 = v_2779 ^ v_2843;
assign v_3998 = v_2780 ^ v_2844;
assign v_3999 = v_2781 ^ v_2845;
assign v_4000 = v_2782 ^ v_2846;
assign v_4001 = v_2783 ^ v_2847;
assign v_4002 = v_2784 ^ v_2848;
assign v_4003 = v_2785 ^ v_2849;
assign v_4004 = v_2786 ^ v_2850;
assign v_4005 = v_2787 ^ v_2851;
assign v_4006 = v_2788 ^ v_2852;
assign v_4007 = v_2789 ^ v_2853;
assign v_4008 = v_2790 ^ v_2854;
assign v_4009 = v_2791 ^ v_2855;
assign v_4010 = v_2792 ^ v_2856;
assign v_4011 = v_2793 ^ v_2857;
assign v_4012 = v_2794 ^ v_2858;
assign v_4013 = v_2795 ^ v_2859;
assign v_4014 = v_2796 ^ v_2860;
assign v_4015 = v_2797 ^ v_2861;
assign v_4016 = v_2798 ^ v_2862;
assign v_4017 = v_2799 ^ v_2863;
assign v_4018 = v_2800 ^ v_2864;
assign v_4019 = v_2801 ^ v_2865;
assign v_4020 = v_2802 ^ v_2866;
assign v_4021 = v_2803 ^ v_2867;
assign v_4022 = v_2804 ^ v_2868;
assign v_4023 = v_2805 ^ v_2869;
assign v_4024 = v_2806 ^ v_2870;
assign v_4025 = v_2807 ^ v_2871;
assign v_4026 = v_2808 ^ v_2872;
assign v_4027 = v_2809 ^ v_2873;
assign v_4028 = v_2810 ^ v_2874;
assign v_4029 = v_2811 ^ v_2875;
assign v_4030 = v_2812 ^ v_2876;
assign v_4031 = v_2813 ^ v_2877;
assign v_4032 = v_2814 ^ v_2878;
assign v_4033 = v_2815 ^ v_2879;
assign v_4034 = v_2816 ^ v_2880;
assign v_4035 = v_2817 ^ v_2881;
assign v_4036 = v_2818 ^ v_2882;
assign v_4037 = v_2819 ^ v_2883;
assign v_4038 = v_2820 ^ v_2884;
assign v_4040 = v_65 ^ v_257;
assign v_4041 = v_66 ^ v_258;
assign v_4042 = v_67 ^ v_259;
assign v_4043 = v_68 ^ v_260;
assign v_4044 = v_69 ^ v_261;
assign v_4045 = v_70 ^ v_262;
assign v_4046 = v_71 ^ v_263;
assign v_4047 = v_72 ^ v_264;
assign v_4048 = v_73 ^ v_265;
assign v_4049 = v_74 ^ v_266;
assign v_4050 = v_75 ^ v_267;
assign v_4051 = v_76 ^ v_268;
assign v_4052 = v_77 ^ v_269;
assign v_4053 = v_78 ^ v_270;
assign v_4054 = v_79 ^ v_271;
assign v_4055 = v_80 ^ v_272;
assign v_4056 = v_81 ^ v_273;
assign v_4057 = v_82 ^ v_274;
assign v_4058 = v_83 ^ v_275;
assign v_4059 = v_84 ^ v_276;
assign v_4060 = v_85 ^ v_277;
assign v_4061 = v_86 ^ v_278;
assign v_4062 = v_87 ^ v_279;
assign v_4063 = v_88 ^ v_280;
assign v_4064 = v_89 ^ v_281;
assign v_4065 = v_90 ^ v_282;
assign v_4066 = v_91 ^ v_283;
assign v_4067 = v_92 ^ v_284;
assign v_4068 = v_93 ^ v_285;
assign v_4069 = v_94 ^ v_286;
assign v_4070 = v_95 ^ v_287;
assign v_4071 = v_96 ^ v_288;
assign v_4072 = v_97 ^ v_289;
assign v_4073 = v_98 ^ v_290;
assign v_4074 = v_99 ^ v_291;
assign v_4075 = v_100 ^ v_292;
assign v_4076 = v_101 ^ v_293;
assign v_4077 = v_102 ^ v_294;
assign v_4078 = v_103 ^ v_295;
assign v_4079 = v_104 ^ v_296;
assign v_4080 = v_105 ^ v_297;
assign v_4081 = v_106 ^ v_298;
assign v_4082 = v_107 ^ v_299;
assign v_4083 = v_108 ^ v_300;
assign v_4084 = v_109 ^ v_301;
assign v_4085 = v_110 ^ v_302;
assign v_4086 = v_111 ^ v_303;
assign v_4087 = v_112 ^ v_304;
assign v_4088 = v_113 ^ v_305;
assign v_4089 = v_114 ^ v_306;
assign v_4090 = v_115 ^ v_307;
assign v_4091 = v_116 ^ v_308;
assign v_4092 = v_117 ^ v_309;
assign v_4093 = v_118 ^ v_310;
assign v_4094 = v_119 ^ v_311;
assign v_4095 = v_120 ^ v_312;
assign v_4096 = v_121 ^ v_313;
assign v_4097 = v_122 ^ v_314;
assign v_4098 = v_123 ^ v_315;
assign v_4099 = v_124 ^ v_316;
assign v_4100 = v_125 ^ v_317;
assign v_4101 = v_126 ^ v_318;
assign v_4102 = v_127 ^ v_319;
assign v_4103 = v_128 ^ v_320;
assign v_4105 = v_3141 ^ v_3205;
assign v_4106 = v_3142 ^ v_3206;
assign v_4107 = v_3143 ^ v_3207;
assign v_4108 = v_3144 ^ v_3208;
assign v_4109 = v_3145 ^ v_3209;
assign v_4110 = v_3146 ^ v_3210;
assign v_4111 = v_3147 ^ v_3211;
assign v_4112 = v_3148 ^ v_3212;
assign v_4113 = v_3149 ^ v_3213;
assign v_4114 = v_3150 ^ v_3214;
assign v_4115 = v_3151 ^ v_3215;
assign v_4116 = v_3152 ^ v_3216;
assign v_4117 = v_3153 ^ v_3217;
assign v_4118 = v_3154 ^ v_3218;
assign v_4119 = v_3155 ^ v_3219;
assign v_4120 = v_3156 ^ v_3220;
assign v_4121 = v_3157 ^ v_3221;
assign v_4122 = v_3158 ^ v_3222;
assign v_4123 = v_3159 ^ v_3223;
assign v_4124 = v_3160 ^ v_3224;
assign v_4125 = v_3161 ^ v_3225;
assign v_4126 = v_3162 ^ v_3226;
assign v_4127 = v_3163 ^ v_3227;
assign v_4128 = v_3164 ^ v_3228;
assign v_4129 = v_3165 ^ v_3229;
assign v_4130 = v_3166 ^ v_3230;
assign v_4131 = v_3167 ^ v_3231;
assign v_4132 = v_3168 ^ v_3232;
assign v_4133 = v_3169 ^ v_3233;
assign v_4134 = v_3170 ^ v_3234;
assign v_4135 = v_3171 ^ v_3235;
assign v_4136 = v_3172 ^ v_3236;
assign v_4137 = v_3173 ^ v_3237;
assign v_4138 = v_3174 ^ v_3238;
assign v_4139 = v_3175 ^ v_3239;
assign v_4140 = v_3176 ^ v_3240;
assign v_4141 = v_3177 ^ v_3241;
assign v_4142 = v_3178 ^ v_3242;
assign v_4143 = v_3179 ^ v_3243;
assign v_4144 = v_3180 ^ v_3244;
assign v_4145 = v_3181 ^ v_3245;
assign v_4146 = v_3182 ^ v_3246;
assign v_4147 = v_3183 ^ v_3247;
assign v_4148 = v_3184 ^ v_3248;
assign v_4149 = v_3185 ^ v_3249;
assign v_4150 = v_3186 ^ v_3250;
assign v_4151 = v_3187 ^ v_3251;
assign v_4152 = v_3188 ^ v_3252;
assign v_4153 = v_3189 ^ v_3253;
assign v_4154 = v_3190 ^ v_3254;
assign v_4155 = v_3191 ^ v_3255;
assign v_4156 = v_3192 ^ v_3256;
assign v_4157 = v_3193 ^ v_3257;
assign v_4158 = v_3194 ^ v_3258;
assign v_4159 = v_3195 ^ v_3259;
assign v_4160 = v_3196 ^ v_3260;
assign v_4161 = v_3197 ^ v_3261;
assign v_4162 = v_3198 ^ v_3262;
assign v_4163 = v_3199 ^ v_3263;
assign v_4164 = v_3200 ^ v_3264;
assign v_4165 = v_3201 ^ v_3265;
assign v_4166 = v_3202 ^ v_3266;
assign v_4167 = v_3203 ^ v_3267;
assign v_4168 = v_3204 ^ v_3268;
assign v_4170 = v_129 ^ v_321;
assign v_4171 = v_130 ^ v_322;
assign v_4172 = v_131 ^ v_323;
assign v_4173 = v_132 ^ v_324;
assign v_4174 = v_133 ^ v_325;
assign v_4175 = v_134 ^ v_326;
assign v_4176 = v_135 ^ v_327;
assign v_4177 = v_136 ^ v_328;
assign v_4178 = v_137 ^ v_329;
assign v_4179 = v_138 ^ v_330;
assign v_4180 = v_139 ^ v_331;
assign v_4181 = v_140 ^ v_332;
assign v_4182 = v_141 ^ v_333;
assign v_4183 = v_142 ^ v_334;
assign v_4184 = v_143 ^ v_335;
assign v_4185 = v_144 ^ v_336;
assign v_4186 = v_145 ^ v_337;
assign v_4187 = v_146 ^ v_338;
assign v_4188 = v_147 ^ v_339;
assign v_4189 = v_148 ^ v_340;
assign v_4190 = v_149 ^ v_341;
assign v_4191 = v_150 ^ v_342;
assign v_4192 = v_151 ^ v_343;
assign v_4193 = v_152 ^ v_344;
assign v_4194 = v_153 ^ v_345;
assign v_4195 = v_154 ^ v_346;
assign v_4196 = v_155 ^ v_347;
assign v_4197 = v_156 ^ v_348;
assign v_4198 = v_157 ^ v_349;
assign v_4199 = v_158 ^ v_350;
assign v_4200 = v_159 ^ v_351;
assign v_4201 = v_160 ^ v_352;
assign v_4202 = v_161 ^ v_353;
assign v_4203 = v_162 ^ v_354;
assign v_4204 = v_163 ^ v_355;
assign v_4205 = v_164 ^ v_356;
assign v_4206 = v_165 ^ v_357;
assign v_4207 = v_166 ^ v_358;
assign v_4208 = v_167 ^ v_359;
assign v_4209 = v_168 ^ v_360;
assign v_4210 = v_169 ^ v_361;
assign v_4211 = v_170 ^ v_362;
assign v_4212 = v_171 ^ v_363;
assign v_4213 = v_172 ^ v_364;
assign v_4214 = v_173 ^ v_365;
assign v_4215 = v_174 ^ v_366;
assign v_4216 = v_175 ^ v_367;
assign v_4217 = v_176 ^ v_368;
assign v_4218 = v_177 ^ v_369;
assign v_4219 = v_178 ^ v_370;
assign v_4220 = v_179 ^ v_371;
assign v_4221 = v_180 ^ v_372;
assign v_4222 = v_181 ^ v_373;
assign v_4223 = v_182 ^ v_374;
assign v_4224 = v_183 ^ v_375;
assign v_4225 = v_184 ^ v_376;
assign v_4226 = v_185 ^ v_377;
assign v_4227 = v_186 ^ v_378;
assign v_4228 = v_187 ^ v_379;
assign v_4229 = v_188 ^ v_380;
assign v_4230 = v_189 ^ v_381;
assign v_4231 = v_190 ^ v_382;
assign v_4232 = v_191 ^ v_383;
assign v_4233 = v_192 ^ v_384;
assign v_4235 = v_3525 ^ v_3589;
assign v_4236 = v_3526 ^ v_3590;
assign v_4237 = v_3527 ^ v_3591;
assign v_4238 = v_3528 ^ v_3592;
assign v_4239 = v_3529 ^ v_3593;
assign v_4240 = v_3530 ^ v_3594;
assign v_4241 = v_3531 ^ v_3595;
assign v_4242 = v_3532 ^ v_3596;
assign v_4243 = v_3533 ^ v_3597;
assign v_4244 = v_3534 ^ v_3598;
assign v_4245 = v_3535 ^ v_3599;
assign v_4246 = v_3536 ^ v_3600;
assign v_4247 = v_3537 ^ v_3601;
assign v_4248 = v_3538 ^ v_3602;
assign v_4249 = v_3539 ^ v_3603;
assign v_4250 = v_3540 ^ v_3604;
assign v_4251 = v_3541 ^ v_3605;
assign v_4252 = v_3542 ^ v_3606;
assign v_4253 = v_3543 ^ v_3607;
assign v_4254 = v_3544 ^ v_3608;
assign v_4255 = v_3545 ^ v_3609;
assign v_4256 = v_3546 ^ v_3610;
assign v_4257 = v_3547 ^ v_3611;
assign v_4258 = v_3548 ^ v_3612;
assign v_4259 = v_3549 ^ v_3613;
assign v_4260 = v_3550 ^ v_3614;
assign v_4261 = v_3551 ^ v_3615;
assign v_4262 = v_3552 ^ v_3616;
assign v_4263 = v_3553 ^ v_3617;
assign v_4264 = v_3554 ^ v_3618;
assign v_4265 = v_3555 ^ v_3619;
assign v_4266 = v_3556 ^ v_3620;
assign v_4267 = v_3557 ^ v_3621;
assign v_4268 = v_3558 ^ v_3622;
assign v_4269 = v_3559 ^ v_3623;
assign v_4270 = v_3560 ^ v_3624;
assign v_4271 = v_3561 ^ v_3625;
assign v_4272 = v_3562 ^ v_3626;
assign v_4273 = v_3563 ^ v_3627;
assign v_4274 = v_3564 ^ v_3628;
assign v_4275 = v_3565 ^ v_3629;
assign v_4276 = v_3566 ^ v_3630;
assign v_4277 = v_3567 ^ v_3631;
assign v_4278 = v_3568 ^ v_3632;
assign v_4279 = v_3569 ^ v_3633;
assign v_4280 = v_3570 ^ v_3634;
assign v_4281 = v_3571 ^ v_3635;
assign v_4282 = v_3572 ^ v_3636;
assign v_4283 = v_3573 ^ v_3637;
assign v_4284 = v_3574 ^ v_3638;
assign v_4285 = v_3575 ^ v_3639;
assign v_4286 = v_3576 ^ v_3640;
assign v_4287 = v_3577 ^ v_3641;
assign v_4288 = v_3578 ^ v_3642;
assign v_4289 = v_3579 ^ v_3643;
assign v_4290 = v_3580 ^ v_3644;
assign v_4291 = v_3581 ^ v_3645;
assign v_4292 = v_3582 ^ v_3646;
assign v_4293 = v_3583 ^ v_3647;
assign v_4294 = v_3584 ^ v_3648;
assign v_4295 = v_3585 ^ v_3649;
assign v_4296 = v_3586 ^ v_3650;
assign v_4297 = v_3587 ^ v_3651;
assign v_4298 = v_3588 ^ v_3652;
assign x_1 = v_1086 | ~v_1087;
assign x_2 = v_1215 | ~v_1216;
assign x_3 = v_3138 | ~v_3139;
assign x_4 = v_3522 | ~v_3523;
assign x_5 = v_3906 | ~v_3907;
assign x_6 = v_4039 | ~v_3974;
assign x_7 = v_4169 | ~v_4104;
assign x_8 = v_4299 | ~v_4234;
assign x_9 = x_1 & x_2;
assign x_10 = x_3 & x_4;
assign x_11 = x_9 & x_10;
assign x_12 = x_5 & x_6;
assign x_13 = x_7 & x_8;
assign x_14 = x_12 & x_13;
assign x_15 = x_11 & x_14;
assign o_1 = x_15;
endmodule
