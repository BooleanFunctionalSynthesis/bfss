// Generated using findDep.cpp 
module stmt28_89_97 (v_2, v_3, v_4, v_5, v_7, v_8, v_213, v_214, v_219, v_221, v_225, v_227, v_229, v_230, v_232, v_234, v_236, v_237, v_239, v_241, v_243, v_245, v_247, v_249, v_251, v_254, v_255, v_262, v_264, v_268, v_272, v_274, v_279, v_280, v_281, v_283, v_286, v_288, v_292, v_293, v_295, v_297, v_298, v_303, v_308, v_309, v_311, v_312, v_316, v_318, v_322, v_324, v_326, v_333, v_334, v_336, v_338, v_340, v_345, v_346, v_348, v_350, v_352, v_354, v_357, v_359, v_360, v_362, v_364, v_366, v_370, v_372, v_373, v_375, v_377, v_379, v_381, v_385, v_389, v_391, v_392, v_394, v_396, v_398, v_400, v_406, v_410, v_411, v_413, v_415, v_417, v_419, v_422, v_424, v_425, v_427, v_429, v_431, v_435, v_437, v_438, v_440, v_442, v_444, v_446, v_450, v_454, v_456, v_457, v_459, v_461, v_463, v_465, v_471, v_475, v_477, v_481, v_486, v_489, v_491, v_493, v_494, v_496, v_498, v_500, v_501, v_503, v_505, v_507, v_509, v_511, v_513, v_515, v_518, v_519, v_526, v_528, v_532, v_537, v_542, v_543, v_547, v_549, v_551, v_555, v_559, v_561, v_563, v_565, v_569, v_571, v_573, v_574, v_578, v_583, v_584, v_586, v_589, v_591, v_594, v_600, v_601, v_605, v_607, v_609, v_613, v_617, v_619, v_621, v_623, v_627, v_629, v_631, v_632, v_636, v_641, v_643, v_645, v_647, v_649, v_663, v_666, v_669, v_670, v_672, v_674, v_675, v_680, v_682, v_684, v_685, v_687, v_690, v_692, v_695, v_700, v_705, v_706, v_707, v_711, v_713, v_715, v_719, v_723, v_724, v_726, v_727, v_729, v_731, v_733, v_735, v_738, v_739, v_742, v_746, v_747, v_751, v_753, v_755, v_759, v_760, v_764, v_766, v_768, v_772, v_775, v_776, v_780, v_782, v_784, v_788, v_792, v_798, v_799, v_800, v_801, v_805, v_809, v_811, v_815, v_817, v_822, v_823, v_824, v_828, v_832, v_834, v_838, v_840, v_845, v_846, v_847, v_851, v_855, v_857, v_861, v_863, v_868, v_869, v_870, v_872, v_879, v_880, v_881, v_882, v_886, v_890, v_892, v_896, v_898, v_903, v_904, v_905, v_909, v_913, v_915, v_919, v_921, v_926, v_927, v_928, v_932, v_936, v_938, v_942, v_944, v_949, v_950, v_951, v_953, v_960, v_961, v_962, v_963, v_967, v_971, v_973, v_977, v_979, v_984, v_985, v_986, v_990, v_994, v_996, v_1000, v_1002, v_1007, v_1008, v_1009, v_1013, v_1017, v_1019, v_1023, v_1025, v_1030, v_1031, v_1032, v_1034, v_1041, v_1042, v_1043, v_1044, v_1048, v_1052, v_1054, v_1058, v_1060, v_1065, v_1066, v_1067, v_1071, v_1075, v_1077, v_1081, v_1083, v_1088, v_1089, v_1090, v_1094, v_1098, v_1100, v_1104, v_1106, v_1111, v_1112, v_1113, v_1115, v_1122, v_1123, v_1124, v_1125, v_1129, v_1133, v_1135, v_1139, v_1141, v_1146, v_1147, v_1148, v_1152, v_1156, v_1158, v_1162, v_1164, v_1169, v_1170, v_1171, v_1175, v_1179, v_1181, v_1185, v_1187, v_1192, v_1193, v_1194, v_1196, v_1203, v_1204, v_1205, v_1206, v_1210, v_1214, v_1216, v_1220, v_1222, v_1227, v_1228, v_1229, v_1233, v_1237, v_1239, v_1243, v_1245, v_1250, v_1251, v_1252, v_1256, v_1260, v_1262, v_1266, v_1268, v_1273, v_1274, v_1275, v_1277, v_1284, v_1285, v_1286, v_1287, v_1291, v_1295, v_1297, v_1301, v_1303, v_1308, v_1309, v_1310, v_1314, v_1318, v_1320, v_1324, v_1326, v_1331, v_1332, v_1333, v_1337, v_1341, v_1343, v_1347, v_1349, v_1354, v_1355, v_1356, v_1358, v_1365, v_1366, v_1367, v_1368, v_1372, v_1376, v_1378, v_1382, v_1384, v_1389, v_1390, v_1391, v_1395, v_1399, v_1401, v_1405, v_1407, v_1412, v_1413, v_1414, v_1418, v_1422, v_1424, v_1428, v_1430, v_1435, v_1436, v_1437, v_1439, v_1446, v_1447, v_1448, v_1449, v_1453, v_1457, v_1459, v_1463, v_1465, v_1470, v_1471, v_1472, v_1476, v_1480, v_1482, v_1486, v_1488, v_1493, v_1494, v_1495, v_1499, v_1503, v_1505, v_1509, v_1511, v_1516, v_1517, v_1518, v_1520, v_1527, v_1528, v_1529, v_1533, v_1654, v_1655, v_2118, v_2122, v_2218, v_2744, v_2764, v_2815, v_2833, v_3277, v_3297, v_3348, v_3366, v_3688, v_3813, v_3833, v_3884, v_3902, v_4224, v_4349, v_4369, v_4420, v_4438, v_4884, v_4904, v_4955, v_4973, v_5295, v_5420, v_5440, v_5491, v_5509, v_5831, v_5836, v_5931, v_6332, v_6457, v_6477, v_6528, v_6546, v_6868, v_6869, v_6870, v_6871, v_6873, v_6874, v_7079, v_7080, v_7085, v_7087, v_7091, v_7093, v_7095, v_7096, v_7098, v_7100, v_7102, v_7103, v_7105, v_7107, v_7109, v_7111, v_7113, v_7115, v_7117, v_7120, v_7121, v_7128, v_7130, v_7134, v_7138, v_7140, v_7145, v_7146, v_7147, v_7149, v_7152, v_7154, v_7158, v_7159, v_7161, v_7163, v_7164, v_7169, v_7174, v_7175, v_7177, v_7178, v_7182, v_7184, v_7188, v_7190, v_7192, v_7199, v_7200, v_7202, v_7204, v_7206, v_7211, v_7212, v_7214, v_7216, v_7218, v_7220, v_7223, v_7225, v_7226, v_7228, v_7230, v_7232, v_7236, v_7238, v_7239, v_7241, v_7243, v_7245, v_7247, v_7251, v_7255, v_7257, v_7258, v_7260, v_7262, v_7264, v_7266, v_7272, v_7276, v_7277, v_7279, v_7281, v_7283, v_7285, v_7288, v_7290, v_7291, v_7293, v_7295, v_7297, v_7301, v_7303, v_7304, v_7306, v_7308, v_7310, v_7312, v_7316, v_7320, v_7322, v_7323, v_7325, v_7327, v_7329, v_7331, v_7337, v_7341, v_7343, v_7347, v_7352, v_7355, v_7357, v_7359, v_7360, v_7362, v_7364, v_7366, v_7367, v_7369, v_7371, v_7373, v_7375, v_7377, v_7379, v_7381, v_7384, v_7385, v_7392, v_7394, v_7398, v_7403, v_7408, v_7409, v_7413, v_7415, v_7417, v_7421, v_7425, v_7427, v_7429, v_7431, v_7435, v_7437, v_7439, v_7440, v_7444, v_7449, v_7450, v_7452, v_7455, v_7457, v_7460, v_7466, v_7467, v_7471, v_7473, v_7475, v_7479, v_7483, v_7485, v_7487, v_7489, v_7493, v_7495, v_7497, v_7498, v_7502, v_7507, v_7509, v_7511, v_7513, v_7515, v_7529, v_7532, v_7535, v_7536, v_7538, v_7540, v_7541, v_7546, v_7548, v_7550, v_7551, v_7553, v_7556, v_7558, v_7561, v_7566, v_7571, v_7572, v_7573, v_7577, v_7579, v_7581, v_7585, v_7589, v_7590, v_7592, v_7593, v_7595, v_7597, v_7599, v_7601, v_7604, v_7605, v_7608, v_7612, v_7613, v_7617, v_7619, v_7621, v_7625, v_7626, v_7630, v_7632, v_7634, v_7638, v_7641, v_7642, v_7646, v_7648, v_7650, v_7654, v_7658, v_7664, v_7665, v_7666, v_7667, v_7671, v_7675, v_7677, v_7681, v_7683, v_7688, v_7689, v_7690, v_7694, v_7698, v_7700, v_7704, v_7706, v_7711, v_7712, v_7713, v_7717, v_7721, v_7723, v_7727, v_7729, v_7734, v_7735, v_7736, v_7738, v_7745, v_7746, v_7747, v_7748, v_7752, v_7756, v_7758, v_7762, v_7764, v_7769, v_7770, v_7771, v_7775, v_7779, v_7781, v_7785, v_7787, v_7792, v_7793, v_7794, v_7798, v_7802, v_7804, v_7808, v_7810, v_7815, v_7816, v_7817, v_7819, v_7826, v_7827, v_7828, v_7829, v_7833, v_7837, v_7839, v_7843, v_7845, v_7850, v_7851, v_7852, v_7856, v_7860, v_7862, v_7866, v_7868, v_7873, v_7874, v_7875, v_7879, v_7883, v_7885, v_7889, v_7891, v_7896, v_7897, v_7898, v_7900, v_7907, v_7908, v_7909, v_7910, v_7914, v_7918, v_7920, v_7924, v_7926, v_7931, v_7932, v_7933, v_7937, v_7941, v_7943, v_7947, v_7949, v_7954, v_7955, v_7956, v_7960, v_7964, v_7966, v_7970, v_7972, v_7977, v_7978, v_7979, v_7981, v_7988, v_7989, v_7990, v_7991, v_7995, v_7999, v_8001, v_8005, v_8007, v_8012, v_8013, v_8014, v_8018, v_8022, v_8024, v_8028, v_8030, v_8035, v_8036, v_8037, v_8041, v_8045, v_8047, v_8051, v_8053, v_8058, v_8059, v_8060, v_8062, v_8069, v_8070, v_8071, v_8072, v_8076, v_8080, v_8082, v_8086, v_8088, v_8093, v_8094, v_8095, v_8099, v_8103, v_8105, v_8109, v_8111, v_8116, v_8117, v_8118, v_8122, v_8126, v_8128, v_8132, v_8134, v_8139, v_8140, v_8141, v_8143, v_8150, v_8151, v_8152, v_8153, v_8157, v_8161, v_8163, v_8167, v_8169, v_8174, v_8175, v_8176, v_8180, v_8184, v_8186, v_8190, v_8192, v_8197, v_8198, v_8199, v_8203, v_8207, v_8209, v_8213, v_8215, v_8220, v_8221, v_8222, v_8224, v_8231, v_8232, v_8233, v_8237, v_8358, v_8359, v_8744, v_8748, v_8844, v_9300, v_9320, v_9371, v_9389, v_9763, v_9783, v_9834, v_9852, v_10104, v_10229, v_10249, v_10300, v_10318, v_10570, v_10695, v_10715, v_10766, v_10784, v_11160, v_11180, v_11231, v_11249, v_11501, v_11626, v_11646, v_11697, v_11715, v_11967, v_11972, v_12067, v_12398, v_12523, v_12543, v_12594, v_12612, o_1);
input v_2;
input v_3;
input v_4;
input v_5;
input v_7;
input v_8;
input v_213;
input v_214;
input v_219;
input v_221;
input v_225;
input v_227;
input v_229;
input v_230;
input v_232;
input v_234;
input v_236;
input v_237;
input v_239;
input v_241;
input v_243;
input v_245;
input v_247;
input v_249;
input v_251;
input v_254;
input v_255;
input v_262;
input v_264;
input v_268;
input v_272;
input v_274;
input v_279;
input v_280;
input v_281;
input v_283;
input v_286;
input v_288;
input v_292;
input v_293;
input v_295;
input v_297;
input v_298;
input v_303;
input v_308;
input v_309;
input v_311;
input v_312;
input v_316;
input v_318;
input v_322;
input v_324;
input v_326;
input v_333;
input v_334;
input v_336;
input v_338;
input v_340;
input v_345;
input v_346;
input v_348;
input v_350;
input v_352;
input v_354;
input v_357;
input v_359;
input v_360;
input v_362;
input v_364;
input v_366;
input v_370;
input v_372;
input v_373;
input v_375;
input v_377;
input v_379;
input v_381;
input v_385;
input v_389;
input v_391;
input v_392;
input v_394;
input v_396;
input v_398;
input v_400;
input v_406;
input v_410;
input v_411;
input v_413;
input v_415;
input v_417;
input v_419;
input v_422;
input v_424;
input v_425;
input v_427;
input v_429;
input v_431;
input v_435;
input v_437;
input v_438;
input v_440;
input v_442;
input v_444;
input v_446;
input v_450;
input v_454;
input v_456;
input v_457;
input v_459;
input v_461;
input v_463;
input v_465;
input v_471;
input v_475;
input v_477;
input v_481;
input v_486;
input v_489;
input v_491;
input v_493;
input v_494;
input v_496;
input v_498;
input v_500;
input v_501;
input v_503;
input v_505;
input v_507;
input v_509;
input v_511;
input v_513;
input v_515;
input v_518;
input v_519;
input v_526;
input v_528;
input v_532;
input v_537;
input v_542;
input v_543;
input v_547;
input v_549;
input v_551;
input v_555;
input v_559;
input v_561;
input v_563;
input v_565;
input v_569;
input v_571;
input v_573;
input v_574;
input v_578;
input v_583;
input v_584;
input v_586;
input v_589;
input v_591;
input v_594;
input v_600;
input v_601;
input v_605;
input v_607;
input v_609;
input v_613;
input v_617;
input v_619;
input v_621;
input v_623;
input v_627;
input v_629;
input v_631;
input v_632;
input v_636;
input v_641;
input v_643;
input v_645;
input v_647;
input v_649;
input v_663;
input v_666;
input v_669;
input v_670;
input v_672;
input v_674;
input v_675;
input v_680;
input v_682;
input v_684;
input v_685;
input v_687;
input v_690;
input v_692;
input v_695;
input v_700;
input v_705;
input v_706;
input v_707;
input v_711;
input v_713;
input v_715;
input v_719;
input v_723;
input v_724;
input v_726;
input v_727;
input v_729;
input v_731;
input v_733;
input v_735;
input v_738;
input v_739;
input v_742;
input v_746;
input v_747;
input v_751;
input v_753;
input v_755;
input v_759;
input v_760;
input v_764;
input v_766;
input v_768;
input v_772;
input v_775;
input v_776;
input v_780;
input v_782;
input v_784;
input v_788;
input v_792;
input v_798;
input v_799;
input v_800;
input v_801;
input v_805;
input v_809;
input v_811;
input v_815;
input v_817;
input v_822;
input v_823;
input v_824;
input v_828;
input v_832;
input v_834;
input v_838;
input v_840;
input v_845;
input v_846;
input v_847;
input v_851;
input v_855;
input v_857;
input v_861;
input v_863;
input v_868;
input v_869;
input v_870;
input v_872;
input v_879;
input v_880;
input v_881;
input v_882;
input v_886;
input v_890;
input v_892;
input v_896;
input v_898;
input v_903;
input v_904;
input v_905;
input v_909;
input v_913;
input v_915;
input v_919;
input v_921;
input v_926;
input v_927;
input v_928;
input v_932;
input v_936;
input v_938;
input v_942;
input v_944;
input v_949;
input v_950;
input v_951;
input v_953;
input v_960;
input v_961;
input v_962;
input v_963;
input v_967;
input v_971;
input v_973;
input v_977;
input v_979;
input v_984;
input v_985;
input v_986;
input v_990;
input v_994;
input v_996;
input v_1000;
input v_1002;
input v_1007;
input v_1008;
input v_1009;
input v_1013;
input v_1017;
input v_1019;
input v_1023;
input v_1025;
input v_1030;
input v_1031;
input v_1032;
input v_1034;
input v_1041;
input v_1042;
input v_1043;
input v_1044;
input v_1048;
input v_1052;
input v_1054;
input v_1058;
input v_1060;
input v_1065;
input v_1066;
input v_1067;
input v_1071;
input v_1075;
input v_1077;
input v_1081;
input v_1083;
input v_1088;
input v_1089;
input v_1090;
input v_1094;
input v_1098;
input v_1100;
input v_1104;
input v_1106;
input v_1111;
input v_1112;
input v_1113;
input v_1115;
input v_1122;
input v_1123;
input v_1124;
input v_1125;
input v_1129;
input v_1133;
input v_1135;
input v_1139;
input v_1141;
input v_1146;
input v_1147;
input v_1148;
input v_1152;
input v_1156;
input v_1158;
input v_1162;
input v_1164;
input v_1169;
input v_1170;
input v_1171;
input v_1175;
input v_1179;
input v_1181;
input v_1185;
input v_1187;
input v_1192;
input v_1193;
input v_1194;
input v_1196;
input v_1203;
input v_1204;
input v_1205;
input v_1206;
input v_1210;
input v_1214;
input v_1216;
input v_1220;
input v_1222;
input v_1227;
input v_1228;
input v_1229;
input v_1233;
input v_1237;
input v_1239;
input v_1243;
input v_1245;
input v_1250;
input v_1251;
input v_1252;
input v_1256;
input v_1260;
input v_1262;
input v_1266;
input v_1268;
input v_1273;
input v_1274;
input v_1275;
input v_1277;
input v_1284;
input v_1285;
input v_1286;
input v_1287;
input v_1291;
input v_1295;
input v_1297;
input v_1301;
input v_1303;
input v_1308;
input v_1309;
input v_1310;
input v_1314;
input v_1318;
input v_1320;
input v_1324;
input v_1326;
input v_1331;
input v_1332;
input v_1333;
input v_1337;
input v_1341;
input v_1343;
input v_1347;
input v_1349;
input v_1354;
input v_1355;
input v_1356;
input v_1358;
input v_1365;
input v_1366;
input v_1367;
input v_1368;
input v_1372;
input v_1376;
input v_1378;
input v_1382;
input v_1384;
input v_1389;
input v_1390;
input v_1391;
input v_1395;
input v_1399;
input v_1401;
input v_1405;
input v_1407;
input v_1412;
input v_1413;
input v_1414;
input v_1418;
input v_1422;
input v_1424;
input v_1428;
input v_1430;
input v_1435;
input v_1436;
input v_1437;
input v_1439;
input v_1446;
input v_1447;
input v_1448;
input v_1449;
input v_1453;
input v_1457;
input v_1459;
input v_1463;
input v_1465;
input v_1470;
input v_1471;
input v_1472;
input v_1476;
input v_1480;
input v_1482;
input v_1486;
input v_1488;
input v_1493;
input v_1494;
input v_1495;
input v_1499;
input v_1503;
input v_1505;
input v_1509;
input v_1511;
input v_1516;
input v_1517;
input v_1518;
input v_1520;
input v_1527;
input v_1528;
input v_1529;
input v_1533;
input v_1654;
input v_1655;
input v_2118;
input v_2122;
input v_2218;
input v_2744;
input v_2764;
input v_2815;
input v_2833;
input v_3277;
input v_3297;
input v_3348;
input v_3366;
input v_3688;
input v_3813;
input v_3833;
input v_3884;
input v_3902;
input v_4224;
input v_4349;
input v_4369;
input v_4420;
input v_4438;
input v_4884;
input v_4904;
input v_4955;
input v_4973;
input v_5295;
input v_5420;
input v_5440;
input v_5491;
input v_5509;
input v_5831;
input v_5836;
input v_5931;
input v_6332;
input v_6457;
input v_6477;
input v_6528;
input v_6546;
input v_6868;
input v_6869;
input v_6870;
input v_6871;
input v_6873;
input v_6874;
input v_7079;
input v_7080;
input v_7085;
input v_7087;
input v_7091;
input v_7093;
input v_7095;
input v_7096;
input v_7098;
input v_7100;
input v_7102;
input v_7103;
input v_7105;
input v_7107;
input v_7109;
input v_7111;
input v_7113;
input v_7115;
input v_7117;
input v_7120;
input v_7121;
input v_7128;
input v_7130;
input v_7134;
input v_7138;
input v_7140;
input v_7145;
input v_7146;
input v_7147;
input v_7149;
input v_7152;
input v_7154;
input v_7158;
input v_7159;
input v_7161;
input v_7163;
input v_7164;
input v_7169;
input v_7174;
input v_7175;
input v_7177;
input v_7178;
input v_7182;
input v_7184;
input v_7188;
input v_7190;
input v_7192;
input v_7199;
input v_7200;
input v_7202;
input v_7204;
input v_7206;
input v_7211;
input v_7212;
input v_7214;
input v_7216;
input v_7218;
input v_7220;
input v_7223;
input v_7225;
input v_7226;
input v_7228;
input v_7230;
input v_7232;
input v_7236;
input v_7238;
input v_7239;
input v_7241;
input v_7243;
input v_7245;
input v_7247;
input v_7251;
input v_7255;
input v_7257;
input v_7258;
input v_7260;
input v_7262;
input v_7264;
input v_7266;
input v_7272;
input v_7276;
input v_7277;
input v_7279;
input v_7281;
input v_7283;
input v_7285;
input v_7288;
input v_7290;
input v_7291;
input v_7293;
input v_7295;
input v_7297;
input v_7301;
input v_7303;
input v_7304;
input v_7306;
input v_7308;
input v_7310;
input v_7312;
input v_7316;
input v_7320;
input v_7322;
input v_7323;
input v_7325;
input v_7327;
input v_7329;
input v_7331;
input v_7337;
input v_7341;
input v_7343;
input v_7347;
input v_7352;
input v_7355;
input v_7357;
input v_7359;
input v_7360;
input v_7362;
input v_7364;
input v_7366;
input v_7367;
input v_7369;
input v_7371;
input v_7373;
input v_7375;
input v_7377;
input v_7379;
input v_7381;
input v_7384;
input v_7385;
input v_7392;
input v_7394;
input v_7398;
input v_7403;
input v_7408;
input v_7409;
input v_7413;
input v_7415;
input v_7417;
input v_7421;
input v_7425;
input v_7427;
input v_7429;
input v_7431;
input v_7435;
input v_7437;
input v_7439;
input v_7440;
input v_7444;
input v_7449;
input v_7450;
input v_7452;
input v_7455;
input v_7457;
input v_7460;
input v_7466;
input v_7467;
input v_7471;
input v_7473;
input v_7475;
input v_7479;
input v_7483;
input v_7485;
input v_7487;
input v_7489;
input v_7493;
input v_7495;
input v_7497;
input v_7498;
input v_7502;
input v_7507;
input v_7509;
input v_7511;
input v_7513;
input v_7515;
input v_7529;
input v_7532;
input v_7535;
input v_7536;
input v_7538;
input v_7540;
input v_7541;
input v_7546;
input v_7548;
input v_7550;
input v_7551;
input v_7553;
input v_7556;
input v_7558;
input v_7561;
input v_7566;
input v_7571;
input v_7572;
input v_7573;
input v_7577;
input v_7579;
input v_7581;
input v_7585;
input v_7589;
input v_7590;
input v_7592;
input v_7593;
input v_7595;
input v_7597;
input v_7599;
input v_7601;
input v_7604;
input v_7605;
input v_7608;
input v_7612;
input v_7613;
input v_7617;
input v_7619;
input v_7621;
input v_7625;
input v_7626;
input v_7630;
input v_7632;
input v_7634;
input v_7638;
input v_7641;
input v_7642;
input v_7646;
input v_7648;
input v_7650;
input v_7654;
input v_7658;
input v_7664;
input v_7665;
input v_7666;
input v_7667;
input v_7671;
input v_7675;
input v_7677;
input v_7681;
input v_7683;
input v_7688;
input v_7689;
input v_7690;
input v_7694;
input v_7698;
input v_7700;
input v_7704;
input v_7706;
input v_7711;
input v_7712;
input v_7713;
input v_7717;
input v_7721;
input v_7723;
input v_7727;
input v_7729;
input v_7734;
input v_7735;
input v_7736;
input v_7738;
input v_7745;
input v_7746;
input v_7747;
input v_7748;
input v_7752;
input v_7756;
input v_7758;
input v_7762;
input v_7764;
input v_7769;
input v_7770;
input v_7771;
input v_7775;
input v_7779;
input v_7781;
input v_7785;
input v_7787;
input v_7792;
input v_7793;
input v_7794;
input v_7798;
input v_7802;
input v_7804;
input v_7808;
input v_7810;
input v_7815;
input v_7816;
input v_7817;
input v_7819;
input v_7826;
input v_7827;
input v_7828;
input v_7829;
input v_7833;
input v_7837;
input v_7839;
input v_7843;
input v_7845;
input v_7850;
input v_7851;
input v_7852;
input v_7856;
input v_7860;
input v_7862;
input v_7866;
input v_7868;
input v_7873;
input v_7874;
input v_7875;
input v_7879;
input v_7883;
input v_7885;
input v_7889;
input v_7891;
input v_7896;
input v_7897;
input v_7898;
input v_7900;
input v_7907;
input v_7908;
input v_7909;
input v_7910;
input v_7914;
input v_7918;
input v_7920;
input v_7924;
input v_7926;
input v_7931;
input v_7932;
input v_7933;
input v_7937;
input v_7941;
input v_7943;
input v_7947;
input v_7949;
input v_7954;
input v_7955;
input v_7956;
input v_7960;
input v_7964;
input v_7966;
input v_7970;
input v_7972;
input v_7977;
input v_7978;
input v_7979;
input v_7981;
input v_7988;
input v_7989;
input v_7990;
input v_7991;
input v_7995;
input v_7999;
input v_8001;
input v_8005;
input v_8007;
input v_8012;
input v_8013;
input v_8014;
input v_8018;
input v_8022;
input v_8024;
input v_8028;
input v_8030;
input v_8035;
input v_8036;
input v_8037;
input v_8041;
input v_8045;
input v_8047;
input v_8051;
input v_8053;
input v_8058;
input v_8059;
input v_8060;
input v_8062;
input v_8069;
input v_8070;
input v_8071;
input v_8072;
input v_8076;
input v_8080;
input v_8082;
input v_8086;
input v_8088;
input v_8093;
input v_8094;
input v_8095;
input v_8099;
input v_8103;
input v_8105;
input v_8109;
input v_8111;
input v_8116;
input v_8117;
input v_8118;
input v_8122;
input v_8126;
input v_8128;
input v_8132;
input v_8134;
input v_8139;
input v_8140;
input v_8141;
input v_8143;
input v_8150;
input v_8151;
input v_8152;
input v_8153;
input v_8157;
input v_8161;
input v_8163;
input v_8167;
input v_8169;
input v_8174;
input v_8175;
input v_8176;
input v_8180;
input v_8184;
input v_8186;
input v_8190;
input v_8192;
input v_8197;
input v_8198;
input v_8199;
input v_8203;
input v_8207;
input v_8209;
input v_8213;
input v_8215;
input v_8220;
input v_8221;
input v_8222;
input v_8224;
input v_8231;
input v_8232;
input v_8233;
input v_8237;
input v_8358;
input v_8359;
input v_8744;
input v_8748;
input v_8844;
input v_9300;
input v_9320;
input v_9371;
input v_9389;
input v_9763;
input v_9783;
input v_9834;
input v_9852;
input v_10104;
input v_10229;
input v_10249;
input v_10300;
input v_10318;
input v_10570;
input v_10695;
input v_10715;
input v_10766;
input v_10784;
input v_11160;
input v_11180;
input v_11231;
input v_11249;
input v_11501;
input v_11626;
input v_11646;
input v_11697;
input v_11715;
input v_11967;
input v_11972;
input v_12067;
input v_12398;
input v_12523;
input v_12543;
input v_12594;
input v_12612;
output o_1;
wire v_1;
wire v_6;
wire v_9;
wire v_10;
wire v_11;
wire v_12;
wire v_13;
wire v_14;
wire v_15;
wire v_16;
wire v_17;
wire v_18;
wire v_19;
wire v_20;
wire v_21;
wire v_22;
wire v_23;
wire v_24;
wire v_25;
wire v_26;
wire v_27;
wire v_28;
wire v_29;
wire v_30;
wire v_31;
wire v_32;
wire v_33;
wire v_34;
wire v_35;
wire v_36;
wire v_37;
wire v_38;
wire v_39;
wire v_40;
wire v_41;
wire v_42;
wire v_43;
wire v_44;
wire v_45;
wire v_46;
wire v_47;
wire v_48;
wire v_49;
wire v_50;
wire v_51;
wire v_52;
wire v_53;
wire v_54;
wire v_55;
wire v_56;
wire v_57;
wire v_58;
wire v_59;
wire v_60;
wire v_61;
wire v_62;
wire v_63;
wire v_64;
wire v_65;
wire v_66;
wire v_67;
wire v_68;
wire v_69;
wire v_70;
wire v_71;
wire v_72;
wire v_73;
wire v_74;
wire v_75;
wire v_76;
wire v_77;
wire v_78;
wire v_79;
wire v_80;
wire v_81;
wire v_82;
wire v_83;
wire v_84;
wire v_85;
wire v_86;
wire v_87;
wire v_88;
wire v_89;
wire v_90;
wire v_91;
wire v_92;
wire v_93;
wire v_94;
wire v_95;
wire v_96;
wire v_97;
wire v_98;
wire v_99;
wire v_100;
wire v_101;
wire v_102;
wire v_103;
wire v_104;
wire v_105;
wire v_106;
wire v_107;
wire v_108;
wire v_109;
wire v_110;
wire v_111;
wire v_112;
wire v_113;
wire v_114;
wire v_115;
wire v_116;
wire v_117;
wire v_118;
wire v_119;
wire v_120;
wire v_121;
wire v_122;
wire v_123;
wire v_124;
wire v_125;
wire v_126;
wire v_127;
wire v_128;
wire v_129;
wire v_130;
wire v_131;
wire v_132;
wire v_133;
wire v_134;
wire v_135;
wire v_136;
wire v_137;
wire v_138;
wire v_139;
wire v_140;
wire v_141;
wire v_142;
wire v_143;
wire v_144;
wire v_145;
wire v_146;
wire v_147;
wire v_148;
wire v_149;
wire v_150;
wire v_151;
wire v_152;
wire v_153;
wire v_154;
wire v_155;
wire v_156;
wire v_157;
wire v_158;
wire v_159;
wire v_160;
wire v_161;
wire v_162;
wire v_163;
wire v_164;
wire v_165;
wire v_166;
wire v_167;
wire v_168;
wire v_169;
wire v_170;
wire v_171;
wire v_172;
wire v_173;
wire v_174;
wire v_175;
wire v_176;
wire v_177;
wire v_178;
wire v_179;
wire v_180;
wire v_181;
wire v_182;
wire v_183;
wire v_184;
wire v_185;
wire v_186;
wire v_187;
wire v_188;
wire v_189;
wire v_190;
wire v_191;
wire v_192;
wire v_193;
wire v_194;
wire v_195;
wire v_196;
wire v_197;
wire v_198;
wire v_199;
wire v_200;
wire v_201;
wire v_202;
wire v_203;
wire v_204;
wire v_205;
wire v_206;
wire v_207;
wire v_208;
wire v_209;
wire v_210;
wire v_211;
wire v_212;
wire v_215;
wire v_216;
wire v_217;
wire v_218;
wire v_220;
wire v_222;
wire v_223;
wire v_224;
wire v_226;
wire v_228;
wire v_231;
wire v_233;
wire v_235;
wire v_238;
wire v_240;
wire v_242;
wire v_244;
wire v_246;
wire v_248;
wire v_250;
wire v_252;
wire v_253;
wire v_256;
wire v_257;
wire v_258;
wire v_259;
wire v_260;
wire v_261;
wire v_263;
wire v_265;
wire v_266;
wire v_267;
wire v_269;
wire v_270;
wire v_271;
wire v_273;
wire v_275;
wire v_276;
wire v_277;
wire v_278;
wire v_282;
wire v_284;
wire v_285;
wire v_287;
wire v_289;
wire v_290;
wire v_291;
wire v_294;
wire v_296;
wire v_299;
wire v_300;
wire v_301;
wire v_302;
wire v_304;
wire v_305;
wire v_306;
wire v_307;
wire v_310;
wire v_313;
wire v_314;
wire v_315;
wire v_317;
wire v_319;
wire v_320;
wire v_321;
wire v_323;
wire v_325;
wire v_327;
wire v_328;
wire v_329;
wire v_330;
wire v_331;
wire v_332;
wire v_335;
wire v_337;
wire v_339;
wire v_341;
wire v_342;
wire v_343;
wire v_344;
wire v_347;
wire v_349;
wire v_351;
wire v_353;
wire v_355;
wire v_356;
wire v_358;
wire v_361;
wire v_363;
wire v_365;
wire v_367;
wire v_368;
wire v_369;
wire v_371;
wire v_374;
wire v_376;
wire v_378;
wire v_380;
wire v_382;
wire v_383;
wire v_384;
wire v_386;
wire v_387;
wire v_388;
wire v_390;
wire v_393;
wire v_395;
wire v_397;
wire v_399;
wire v_401;
wire v_402;
wire v_403;
wire v_404;
wire v_405;
wire v_407;
wire v_408;
wire v_409;
wire v_412;
wire v_414;
wire v_416;
wire v_418;
wire v_420;
wire v_421;
wire v_423;
wire v_426;
wire v_428;
wire v_430;
wire v_432;
wire v_433;
wire v_434;
wire v_436;
wire v_439;
wire v_441;
wire v_443;
wire v_445;
wire v_447;
wire v_448;
wire v_449;
wire v_451;
wire v_452;
wire v_453;
wire v_455;
wire v_458;
wire v_460;
wire v_462;
wire v_464;
wire v_466;
wire v_467;
wire v_468;
wire v_469;
wire v_470;
wire v_472;
wire v_473;
wire v_474;
wire v_476;
wire v_478;
wire v_479;
wire v_480;
wire v_482;
wire v_483;
wire v_484;
wire v_485;
wire v_487;
wire v_488;
wire v_490;
wire v_492;
wire v_495;
wire v_497;
wire v_499;
wire v_502;
wire v_504;
wire v_506;
wire v_508;
wire v_510;
wire v_512;
wire v_514;
wire v_516;
wire v_517;
wire v_520;
wire v_521;
wire v_522;
wire v_523;
wire v_524;
wire v_525;
wire v_527;
wire v_529;
wire v_530;
wire v_531;
wire v_533;
wire v_534;
wire v_535;
wire v_536;
wire v_538;
wire v_539;
wire v_540;
wire v_541;
wire v_544;
wire v_545;
wire v_546;
wire v_548;
wire v_550;
wire v_552;
wire v_553;
wire v_554;
wire v_556;
wire v_557;
wire v_558;
wire v_560;
wire v_562;
wire v_564;
wire v_566;
wire v_567;
wire v_568;
wire v_570;
wire v_572;
wire v_575;
wire v_576;
wire v_577;
wire v_579;
wire v_580;
wire v_581;
wire v_582;
wire v_585;
wire v_587;
wire v_588;
wire v_590;
wire v_592;
wire v_593;
wire v_595;
wire v_596;
wire v_597;
wire v_598;
wire v_599;
wire v_602;
wire v_603;
wire v_604;
wire v_606;
wire v_608;
wire v_610;
wire v_611;
wire v_612;
wire v_614;
wire v_615;
wire v_616;
wire v_618;
wire v_620;
wire v_622;
wire v_624;
wire v_625;
wire v_626;
wire v_628;
wire v_630;
wire v_633;
wire v_634;
wire v_635;
wire v_637;
wire v_638;
wire v_639;
wire v_640;
wire v_642;
wire v_644;
wire v_646;
wire v_648;
wire v_650;
wire v_651;
wire v_652;
wire v_653;
wire v_654;
wire v_655;
wire v_656;
wire v_657;
wire v_658;
wire v_659;
wire v_660;
wire v_661;
wire v_662;
wire v_664;
wire v_665;
wire v_667;
wire v_668;
wire v_671;
wire v_673;
wire v_676;
wire v_677;
wire v_678;
wire v_679;
wire v_681;
wire v_683;
wire v_686;
wire v_688;
wire v_689;
wire v_691;
wire v_693;
wire v_694;
wire v_696;
wire v_697;
wire v_698;
wire v_699;
wire v_701;
wire v_702;
wire v_703;
wire v_704;
wire v_708;
wire v_709;
wire v_710;
wire v_712;
wire v_714;
wire v_716;
wire v_717;
wire v_718;
wire v_720;
wire v_721;
wire v_722;
wire v_725;
wire v_728;
wire v_730;
wire v_732;
wire v_734;
wire v_736;
wire v_737;
wire v_740;
wire v_741;
wire v_743;
wire v_744;
wire v_745;
wire v_748;
wire v_749;
wire v_750;
wire v_752;
wire v_754;
wire v_756;
wire v_757;
wire v_758;
wire v_761;
wire v_762;
wire v_763;
wire v_765;
wire v_767;
wire v_769;
wire v_770;
wire v_771;
wire v_773;
wire v_774;
wire v_777;
wire v_778;
wire v_779;
wire v_781;
wire v_783;
wire v_785;
wire v_786;
wire v_787;
wire v_789;
wire v_790;
wire v_791;
wire v_793;
wire v_794;
wire v_795;
wire v_796;
wire v_797;
wire v_802;
wire v_803;
wire v_804;
wire v_806;
wire v_807;
wire v_808;
wire v_810;
wire v_812;
wire v_813;
wire v_814;
wire v_816;
wire v_818;
wire v_819;
wire v_820;
wire v_821;
wire v_825;
wire v_826;
wire v_827;
wire v_829;
wire v_830;
wire v_831;
wire v_833;
wire v_835;
wire v_836;
wire v_837;
wire v_839;
wire v_841;
wire v_842;
wire v_843;
wire v_844;
wire v_848;
wire v_849;
wire v_850;
wire v_852;
wire v_853;
wire v_854;
wire v_856;
wire v_858;
wire v_859;
wire v_860;
wire v_862;
wire v_864;
wire v_865;
wire v_866;
wire v_867;
wire v_871;
wire v_873;
wire v_874;
wire v_875;
wire v_876;
wire v_877;
wire v_878;
wire v_883;
wire v_884;
wire v_885;
wire v_887;
wire v_888;
wire v_889;
wire v_891;
wire v_893;
wire v_894;
wire v_895;
wire v_897;
wire v_899;
wire v_900;
wire v_901;
wire v_902;
wire v_906;
wire v_907;
wire v_908;
wire v_910;
wire v_911;
wire v_912;
wire v_914;
wire v_916;
wire v_917;
wire v_918;
wire v_920;
wire v_922;
wire v_923;
wire v_924;
wire v_925;
wire v_929;
wire v_930;
wire v_931;
wire v_933;
wire v_934;
wire v_935;
wire v_937;
wire v_939;
wire v_940;
wire v_941;
wire v_943;
wire v_945;
wire v_946;
wire v_947;
wire v_948;
wire v_952;
wire v_954;
wire v_955;
wire v_956;
wire v_957;
wire v_958;
wire v_959;
wire v_964;
wire v_965;
wire v_966;
wire v_968;
wire v_969;
wire v_970;
wire v_972;
wire v_974;
wire v_975;
wire v_976;
wire v_978;
wire v_980;
wire v_981;
wire v_982;
wire v_983;
wire v_987;
wire v_988;
wire v_989;
wire v_991;
wire v_992;
wire v_993;
wire v_995;
wire v_997;
wire v_998;
wire v_999;
wire v_1001;
wire v_1003;
wire v_1004;
wire v_1005;
wire v_1006;
wire v_1010;
wire v_1011;
wire v_1012;
wire v_1014;
wire v_1015;
wire v_1016;
wire v_1018;
wire v_1020;
wire v_1021;
wire v_1022;
wire v_1024;
wire v_1026;
wire v_1027;
wire v_1028;
wire v_1029;
wire v_1033;
wire v_1035;
wire v_1036;
wire v_1037;
wire v_1038;
wire v_1039;
wire v_1040;
wire v_1045;
wire v_1046;
wire v_1047;
wire v_1049;
wire v_1050;
wire v_1051;
wire v_1053;
wire v_1055;
wire v_1056;
wire v_1057;
wire v_1059;
wire v_1061;
wire v_1062;
wire v_1063;
wire v_1064;
wire v_1068;
wire v_1069;
wire v_1070;
wire v_1072;
wire v_1073;
wire v_1074;
wire v_1076;
wire v_1078;
wire v_1079;
wire v_1080;
wire v_1082;
wire v_1084;
wire v_1085;
wire v_1086;
wire v_1087;
wire v_1091;
wire v_1092;
wire v_1093;
wire v_1095;
wire v_1096;
wire v_1097;
wire v_1099;
wire v_1101;
wire v_1102;
wire v_1103;
wire v_1105;
wire v_1107;
wire v_1108;
wire v_1109;
wire v_1110;
wire v_1114;
wire v_1116;
wire v_1117;
wire v_1118;
wire v_1119;
wire v_1120;
wire v_1121;
wire v_1126;
wire v_1127;
wire v_1128;
wire v_1130;
wire v_1131;
wire v_1132;
wire v_1134;
wire v_1136;
wire v_1137;
wire v_1138;
wire v_1140;
wire v_1142;
wire v_1143;
wire v_1144;
wire v_1145;
wire v_1149;
wire v_1150;
wire v_1151;
wire v_1153;
wire v_1154;
wire v_1155;
wire v_1157;
wire v_1159;
wire v_1160;
wire v_1161;
wire v_1163;
wire v_1165;
wire v_1166;
wire v_1167;
wire v_1168;
wire v_1172;
wire v_1173;
wire v_1174;
wire v_1176;
wire v_1177;
wire v_1178;
wire v_1180;
wire v_1182;
wire v_1183;
wire v_1184;
wire v_1186;
wire v_1188;
wire v_1189;
wire v_1190;
wire v_1191;
wire v_1195;
wire v_1197;
wire v_1198;
wire v_1199;
wire v_1200;
wire v_1201;
wire v_1202;
wire v_1207;
wire v_1208;
wire v_1209;
wire v_1211;
wire v_1212;
wire v_1213;
wire v_1215;
wire v_1217;
wire v_1218;
wire v_1219;
wire v_1221;
wire v_1223;
wire v_1224;
wire v_1225;
wire v_1226;
wire v_1230;
wire v_1231;
wire v_1232;
wire v_1234;
wire v_1235;
wire v_1236;
wire v_1238;
wire v_1240;
wire v_1241;
wire v_1242;
wire v_1244;
wire v_1246;
wire v_1247;
wire v_1248;
wire v_1249;
wire v_1253;
wire v_1254;
wire v_1255;
wire v_1257;
wire v_1258;
wire v_1259;
wire v_1261;
wire v_1263;
wire v_1264;
wire v_1265;
wire v_1267;
wire v_1269;
wire v_1270;
wire v_1271;
wire v_1272;
wire v_1276;
wire v_1278;
wire v_1279;
wire v_1280;
wire v_1281;
wire v_1282;
wire v_1283;
wire v_1288;
wire v_1289;
wire v_1290;
wire v_1292;
wire v_1293;
wire v_1294;
wire v_1296;
wire v_1298;
wire v_1299;
wire v_1300;
wire v_1302;
wire v_1304;
wire v_1305;
wire v_1306;
wire v_1307;
wire v_1311;
wire v_1312;
wire v_1313;
wire v_1315;
wire v_1316;
wire v_1317;
wire v_1319;
wire v_1321;
wire v_1322;
wire v_1323;
wire v_1325;
wire v_1327;
wire v_1328;
wire v_1329;
wire v_1330;
wire v_1334;
wire v_1335;
wire v_1336;
wire v_1338;
wire v_1339;
wire v_1340;
wire v_1342;
wire v_1344;
wire v_1345;
wire v_1346;
wire v_1348;
wire v_1350;
wire v_1351;
wire v_1352;
wire v_1353;
wire v_1357;
wire v_1359;
wire v_1360;
wire v_1361;
wire v_1362;
wire v_1363;
wire v_1364;
wire v_1369;
wire v_1370;
wire v_1371;
wire v_1373;
wire v_1374;
wire v_1375;
wire v_1377;
wire v_1379;
wire v_1380;
wire v_1381;
wire v_1383;
wire v_1385;
wire v_1386;
wire v_1387;
wire v_1388;
wire v_1392;
wire v_1393;
wire v_1394;
wire v_1396;
wire v_1397;
wire v_1398;
wire v_1400;
wire v_1402;
wire v_1403;
wire v_1404;
wire v_1406;
wire v_1408;
wire v_1409;
wire v_1410;
wire v_1411;
wire v_1415;
wire v_1416;
wire v_1417;
wire v_1419;
wire v_1420;
wire v_1421;
wire v_1423;
wire v_1425;
wire v_1426;
wire v_1427;
wire v_1429;
wire v_1431;
wire v_1432;
wire v_1433;
wire v_1434;
wire v_1438;
wire v_1440;
wire v_1441;
wire v_1442;
wire v_1443;
wire v_1444;
wire v_1445;
wire v_1450;
wire v_1451;
wire v_1452;
wire v_1454;
wire v_1455;
wire v_1456;
wire v_1458;
wire v_1460;
wire v_1461;
wire v_1462;
wire v_1464;
wire v_1466;
wire v_1467;
wire v_1468;
wire v_1469;
wire v_1473;
wire v_1474;
wire v_1475;
wire v_1477;
wire v_1478;
wire v_1479;
wire v_1481;
wire v_1483;
wire v_1484;
wire v_1485;
wire v_1487;
wire v_1489;
wire v_1490;
wire v_1491;
wire v_1492;
wire v_1496;
wire v_1497;
wire v_1498;
wire v_1500;
wire v_1501;
wire v_1502;
wire v_1504;
wire v_1506;
wire v_1507;
wire v_1508;
wire v_1510;
wire v_1512;
wire v_1513;
wire v_1514;
wire v_1515;
wire v_1519;
wire v_1521;
wire v_1522;
wire v_1523;
wire v_1524;
wire v_1525;
wire v_1526;
wire v_1530;
wire v_1531;
wire v_1532;
wire v_1534;
wire v_1535;
wire v_1536;
wire v_1537;
wire v_1538;
wire v_1539;
wire v_1540;
wire v_1541;
wire v_1542;
wire v_1543;
wire v_1544;
wire v_1545;
wire v_1546;
wire v_1547;
wire v_1548;
wire v_1549;
wire v_1550;
wire v_1551;
wire v_1552;
wire v_1553;
wire v_1554;
wire v_1555;
wire v_1556;
wire v_1557;
wire v_1558;
wire v_1559;
wire v_1560;
wire v_1561;
wire v_1562;
wire v_1563;
wire v_1564;
wire v_1565;
wire v_1566;
wire v_1567;
wire v_1568;
wire v_1569;
wire v_1570;
wire v_1571;
wire v_1572;
wire v_1573;
wire v_1574;
wire v_1575;
wire v_1576;
wire v_1577;
wire v_1578;
wire v_1579;
wire v_1580;
wire v_1581;
wire v_1582;
wire v_1583;
wire v_1584;
wire v_1585;
wire v_1586;
wire v_1587;
wire v_1588;
wire v_1589;
wire v_1590;
wire v_1591;
wire v_1592;
wire v_1593;
wire v_1594;
wire v_1595;
wire v_1596;
wire v_1597;
wire v_1598;
wire v_1599;
wire v_1600;
wire v_1601;
wire v_1602;
wire v_1603;
wire v_1604;
wire v_1605;
wire v_1606;
wire v_1607;
wire v_1608;
wire v_1609;
wire v_1610;
wire v_1611;
wire v_1612;
wire v_1613;
wire v_1614;
wire v_1615;
wire v_1616;
wire v_1617;
wire v_1618;
wire v_1619;
wire v_1620;
wire v_1621;
wire v_1622;
wire v_1623;
wire v_1624;
wire v_1625;
wire v_1626;
wire v_1627;
wire v_1628;
wire v_1629;
wire v_1630;
wire v_1631;
wire v_1632;
wire v_1633;
wire v_1634;
wire v_1635;
wire v_1636;
wire v_1637;
wire v_1638;
wire v_1639;
wire v_1640;
wire v_1641;
wire v_1642;
wire v_1643;
wire v_1644;
wire v_1645;
wire v_1646;
wire v_1647;
wire v_1648;
wire v_1649;
wire v_1650;
wire v_1651;
wire v_1652;
wire v_1653;
wire v_1656;
wire v_1657;
wire v_1658;
wire v_1659;
wire v_1660;
wire v_1661;
wire v_1662;
wire v_1663;
wire v_1664;
wire v_1665;
wire v_1666;
wire v_1667;
wire v_1668;
wire v_1669;
wire v_1670;
wire v_1671;
wire v_1672;
wire v_1673;
wire v_1674;
wire v_1675;
wire v_1676;
wire v_1677;
wire v_1678;
wire v_1679;
wire v_1680;
wire v_1681;
wire v_1682;
wire v_1683;
wire v_1684;
wire v_1685;
wire v_1686;
wire v_1687;
wire v_1688;
wire v_1689;
wire v_1690;
wire v_1691;
wire v_1692;
wire v_1693;
wire v_1694;
wire v_1695;
wire v_1696;
wire v_1697;
wire v_1698;
wire v_1699;
wire v_1700;
wire v_1701;
wire v_1702;
wire v_1703;
wire v_1704;
wire v_1705;
wire v_1706;
wire v_1707;
wire v_1708;
wire v_1709;
wire v_1710;
wire v_1711;
wire v_1712;
wire v_1713;
wire v_1714;
wire v_1715;
wire v_1716;
wire v_1717;
wire v_1718;
wire v_1719;
wire v_1720;
wire v_1721;
wire v_1722;
wire v_1723;
wire v_1724;
wire v_1725;
wire v_1726;
wire v_1727;
wire v_1728;
wire v_1729;
wire v_1730;
wire v_1731;
wire v_1732;
wire v_1733;
wire v_1734;
wire v_1735;
wire v_1736;
wire v_1737;
wire v_1738;
wire v_1739;
wire v_1740;
wire v_1741;
wire v_1742;
wire v_1743;
wire v_1744;
wire v_1745;
wire v_1746;
wire v_1747;
wire v_1748;
wire v_1749;
wire v_1750;
wire v_1751;
wire v_1752;
wire v_1753;
wire v_1754;
wire v_1755;
wire v_1756;
wire v_1757;
wire v_1758;
wire v_1759;
wire v_1760;
wire v_1761;
wire v_1762;
wire v_1763;
wire v_1764;
wire v_1765;
wire v_1766;
wire v_1767;
wire v_1768;
wire v_1769;
wire v_1770;
wire v_1771;
wire v_1772;
wire v_1773;
wire v_1774;
wire v_1775;
wire v_1776;
wire v_1777;
wire v_1778;
wire v_1779;
wire v_1780;
wire v_1781;
wire v_1782;
wire v_1783;
wire v_1784;
wire v_1785;
wire v_1786;
wire v_1787;
wire v_1788;
wire v_1789;
wire v_1790;
wire v_1791;
wire v_1792;
wire v_1793;
wire v_1794;
wire v_1795;
wire v_1796;
wire v_1797;
wire v_1798;
wire v_1799;
wire v_1800;
wire v_1801;
wire v_1802;
wire v_1803;
wire v_1804;
wire v_1805;
wire v_1806;
wire v_1807;
wire v_1808;
wire v_1809;
wire v_1810;
wire v_1811;
wire v_1812;
wire v_1813;
wire v_1814;
wire v_1815;
wire v_1816;
wire v_1817;
wire v_1818;
wire v_1819;
wire v_1820;
wire v_1821;
wire v_1822;
wire v_1823;
wire v_1824;
wire v_1825;
wire v_1826;
wire v_1827;
wire v_1828;
wire v_1829;
wire v_1830;
wire v_1831;
wire v_1832;
wire v_1833;
wire v_1834;
wire v_1835;
wire v_1836;
wire v_1837;
wire v_1838;
wire v_1839;
wire v_1840;
wire v_1841;
wire v_1842;
wire v_1843;
wire v_1844;
wire v_1845;
wire v_1846;
wire v_1847;
wire v_1848;
wire v_1849;
wire v_1850;
wire v_1851;
wire v_1852;
wire v_1853;
wire v_1854;
wire v_1855;
wire v_1856;
wire v_1857;
wire v_1858;
wire v_1859;
wire v_1860;
wire v_1861;
wire v_1862;
wire v_1863;
wire v_1864;
wire v_1865;
wire v_1866;
wire v_1867;
wire v_1868;
wire v_1869;
wire v_1870;
wire v_1871;
wire v_1872;
wire v_1873;
wire v_1874;
wire v_1875;
wire v_1876;
wire v_1877;
wire v_1878;
wire v_1879;
wire v_1880;
wire v_1881;
wire v_1882;
wire v_1883;
wire v_1884;
wire v_1885;
wire v_1886;
wire v_1887;
wire v_1888;
wire v_1889;
wire v_1890;
wire v_1891;
wire v_1892;
wire v_1893;
wire v_1894;
wire v_1895;
wire v_1896;
wire v_1897;
wire v_1898;
wire v_1899;
wire v_1900;
wire v_1901;
wire v_1902;
wire v_1903;
wire v_1904;
wire v_1905;
wire v_1906;
wire v_1907;
wire v_1908;
wire v_1909;
wire v_1910;
wire v_1911;
wire v_1912;
wire v_1913;
wire v_1914;
wire v_1915;
wire v_1916;
wire v_1917;
wire v_1918;
wire v_1919;
wire v_1920;
wire v_1921;
wire v_1922;
wire v_1923;
wire v_1924;
wire v_1925;
wire v_1926;
wire v_1927;
wire v_1928;
wire v_1929;
wire v_1930;
wire v_1931;
wire v_1932;
wire v_1933;
wire v_1934;
wire v_1935;
wire v_1936;
wire v_1937;
wire v_1938;
wire v_1939;
wire v_1940;
wire v_1941;
wire v_1942;
wire v_1943;
wire v_1944;
wire v_1945;
wire v_1946;
wire v_1947;
wire v_1948;
wire v_1949;
wire v_1950;
wire v_1951;
wire v_1952;
wire v_1953;
wire v_1954;
wire v_1955;
wire v_1956;
wire v_1957;
wire v_1958;
wire v_1959;
wire v_1960;
wire v_1961;
wire v_1962;
wire v_1963;
wire v_1964;
wire v_1965;
wire v_1966;
wire v_1967;
wire v_1968;
wire v_1969;
wire v_1970;
wire v_1971;
wire v_1972;
wire v_1973;
wire v_1974;
wire v_1975;
wire v_1976;
wire v_1977;
wire v_1978;
wire v_1979;
wire v_1980;
wire v_1981;
wire v_1982;
wire v_1983;
wire v_1984;
wire v_1985;
wire v_1986;
wire v_1987;
wire v_1988;
wire v_1989;
wire v_1990;
wire v_1991;
wire v_1992;
wire v_1993;
wire v_1994;
wire v_1995;
wire v_1996;
wire v_1997;
wire v_1998;
wire v_1999;
wire v_2000;
wire v_2001;
wire v_2002;
wire v_2003;
wire v_2004;
wire v_2005;
wire v_2006;
wire v_2007;
wire v_2008;
wire v_2009;
wire v_2010;
wire v_2011;
wire v_2012;
wire v_2013;
wire v_2014;
wire v_2015;
wire v_2016;
wire v_2017;
wire v_2018;
wire v_2019;
wire v_2020;
wire v_2021;
wire v_2022;
wire v_2023;
wire v_2024;
wire v_2025;
wire v_2026;
wire v_2027;
wire v_2028;
wire v_2029;
wire v_2030;
wire v_2031;
wire v_2032;
wire v_2033;
wire v_2034;
wire v_2035;
wire v_2036;
wire v_2037;
wire v_2038;
wire v_2039;
wire v_2040;
wire v_2041;
wire v_2042;
wire v_2043;
wire v_2044;
wire v_2045;
wire v_2046;
wire v_2047;
wire v_2048;
wire v_2049;
wire v_2050;
wire v_2051;
wire v_2052;
wire v_2053;
wire v_2054;
wire v_2055;
wire v_2056;
wire v_2057;
wire v_2058;
wire v_2059;
wire v_2060;
wire v_2061;
wire v_2062;
wire v_2063;
wire v_2064;
wire v_2065;
wire v_2066;
wire v_2067;
wire v_2068;
wire v_2069;
wire v_2070;
wire v_2071;
wire v_2072;
wire v_2073;
wire v_2074;
wire v_2075;
wire v_2076;
wire v_2077;
wire v_2078;
wire v_2079;
wire v_2080;
wire v_2081;
wire v_2082;
wire v_2083;
wire v_2084;
wire v_2085;
wire v_2086;
wire v_2087;
wire v_2088;
wire v_2089;
wire v_2090;
wire v_2091;
wire v_2092;
wire v_2093;
wire v_2094;
wire v_2095;
wire v_2096;
wire v_2097;
wire v_2098;
wire v_2099;
wire v_2100;
wire v_2101;
wire v_2102;
wire v_2103;
wire v_2104;
wire v_2105;
wire v_2106;
wire v_2107;
wire v_2108;
wire v_2109;
wire v_2110;
wire v_2111;
wire v_2112;
wire v_2113;
wire v_2114;
wire v_2115;
wire v_2116;
wire v_2117;
wire v_2119;
wire v_2120;
wire v_2121;
wire v_2123;
wire v_2124;
wire v_2125;
wire v_2126;
wire v_2127;
wire v_2128;
wire v_2129;
wire v_2130;
wire v_2131;
wire v_2132;
wire v_2133;
wire v_2134;
wire v_2135;
wire v_2136;
wire v_2137;
wire v_2138;
wire v_2139;
wire v_2140;
wire v_2141;
wire v_2142;
wire v_2143;
wire v_2144;
wire v_2145;
wire v_2146;
wire v_2147;
wire v_2148;
wire v_2149;
wire v_2150;
wire v_2151;
wire v_2152;
wire v_2153;
wire v_2154;
wire v_2155;
wire v_2156;
wire v_2157;
wire v_2158;
wire v_2159;
wire v_2160;
wire v_2161;
wire v_2162;
wire v_2163;
wire v_2164;
wire v_2165;
wire v_2166;
wire v_2167;
wire v_2168;
wire v_2169;
wire v_2170;
wire v_2171;
wire v_2172;
wire v_2173;
wire v_2174;
wire v_2175;
wire v_2176;
wire v_2177;
wire v_2178;
wire v_2179;
wire v_2180;
wire v_2181;
wire v_2182;
wire v_2183;
wire v_2184;
wire v_2185;
wire v_2186;
wire v_2187;
wire v_2188;
wire v_2189;
wire v_2190;
wire v_2191;
wire v_2192;
wire v_2193;
wire v_2194;
wire v_2195;
wire v_2196;
wire v_2197;
wire v_2198;
wire v_2199;
wire v_2200;
wire v_2201;
wire v_2202;
wire v_2203;
wire v_2204;
wire v_2205;
wire v_2206;
wire v_2207;
wire v_2208;
wire v_2209;
wire v_2210;
wire v_2211;
wire v_2212;
wire v_2213;
wire v_2214;
wire v_2215;
wire v_2216;
wire v_2217;
wire v_2219;
wire v_2220;
wire v_2221;
wire v_2222;
wire v_2223;
wire v_2224;
wire v_2225;
wire v_2226;
wire v_2227;
wire v_2228;
wire v_2229;
wire v_2230;
wire v_2231;
wire v_2232;
wire v_2233;
wire v_2234;
wire v_2235;
wire v_2236;
wire v_2237;
wire v_2238;
wire v_2239;
wire v_2240;
wire v_2241;
wire v_2242;
wire v_2243;
wire v_2244;
wire v_2245;
wire v_2246;
wire v_2247;
wire v_2248;
wire v_2249;
wire v_2250;
wire v_2251;
wire v_2252;
wire v_2253;
wire v_2254;
wire v_2255;
wire v_2256;
wire v_2257;
wire v_2258;
wire v_2259;
wire v_2260;
wire v_2261;
wire v_2262;
wire v_2263;
wire v_2264;
wire v_2265;
wire v_2266;
wire v_2267;
wire v_2268;
wire v_2269;
wire v_2270;
wire v_2271;
wire v_2272;
wire v_2273;
wire v_2274;
wire v_2275;
wire v_2276;
wire v_2277;
wire v_2278;
wire v_2279;
wire v_2280;
wire v_2281;
wire v_2282;
wire v_2283;
wire v_2284;
wire v_2285;
wire v_2286;
wire v_2287;
wire v_2288;
wire v_2289;
wire v_2290;
wire v_2291;
wire v_2292;
wire v_2293;
wire v_2294;
wire v_2295;
wire v_2296;
wire v_2297;
wire v_2298;
wire v_2299;
wire v_2300;
wire v_2301;
wire v_2302;
wire v_2303;
wire v_2304;
wire v_2305;
wire v_2306;
wire v_2307;
wire v_2308;
wire v_2309;
wire v_2310;
wire v_2311;
wire v_2312;
wire v_2313;
wire v_2314;
wire v_2315;
wire v_2316;
wire v_2317;
wire v_2318;
wire v_2319;
wire v_2320;
wire v_2321;
wire v_2322;
wire v_2323;
wire v_2324;
wire v_2325;
wire v_2326;
wire v_2327;
wire v_2328;
wire v_2329;
wire v_2330;
wire v_2331;
wire v_2332;
wire v_2333;
wire v_2334;
wire v_2335;
wire v_2336;
wire v_2337;
wire v_2338;
wire v_2339;
wire v_2340;
wire v_2341;
wire v_2342;
wire v_2343;
wire v_2344;
wire v_2345;
wire v_2346;
wire v_2347;
wire v_2348;
wire v_2349;
wire v_2350;
wire v_2351;
wire v_2352;
wire v_2353;
wire v_2354;
wire v_2355;
wire v_2356;
wire v_2357;
wire v_2358;
wire v_2359;
wire v_2360;
wire v_2361;
wire v_2362;
wire v_2363;
wire v_2364;
wire v_2365;
wire v_2366;
wire v_2367;
wire v_2368;
wire v_2369;
wire v_2370;
wire v_2371;
wire v_2372;
wire v_2373;
wire v_2374;
wire v_2375;
wire v_2376;
wire v_2377;
wire v_2378;
wire v_2379;
wire v_2380;
wire v_2381;
wire v_2382;
wire v_2383;
wire v_2384;
wire v_2385;
wire v_2386;
wire v_2387;
wire v_2388;
wire v_2389;
wire v_2390;
wire v_2391;
wire v_2392;
wire v_2393;
wire v_2394;
wire v_2395;
wire v_2396;
wire v_2397;
wire v_2398;
wire v_2399;
wire v_2400;
wire v_2401;
wire v_2402;
wire v_2403;
wire v_2404;
wire v_2405;
wire v_2406;
wire v_2407;
wire v_2408;
wire v_2409;
wire v_2410;
wire v_2411;
wire v_2412;
wire v_2413;
wire v_2414;
wire v_2415;
wire v_2416;
wire v_2417;
wire v_2418;
wire v_2419;
wire v_2420;
wire v_2421;
wire v_2422;
wire v_2423;
wire v_2424;
wire v_2425;
wire v_2426;
wire v_2427;
wire v_2428;
wire v_2429;
wire v_2430;
wire v_2431;
wire v_2432;
wire v_2433;
wire v_2434;
wire v_2435;
wire v_2436;
wire v_2437;
wire v_2438;
wire v_2439;
wire v_2440;
wire v_2441;
wire v_2442;
wire v_2443;
wire v_2444;
wire v_2445;
wire v_2446;
wire v_2447;
wire v_2448;
wire v_2449;
wire v_2450;
wire v_2451;
wire v_2452;
wire v_2453;
wire v_2454;
wire v_2455;
wire v_2456;
wire v_2457;
wire v_2458;
wire v_2459;
wire v_2460;
wire v_2461;
wire v_2462;
wire v_2463;
wire v_2464;
wire v_2465;
wire v_2466;
wire v_2467;
wire v_2468;
wire v_2469;
wire v_2470;
wire v_2471;
wire v_2472;
wire v_2473;
wire v_2474;
wire v_2475;
wire v_2476;
wire v_2477;
wire v_2478;
wire v_2479;
wire v_2480;
wire v_2481;
wire v_2482;
wire v_2483;
wire v_2484;
wire v_2485;
wire v_2486;
wire v_2487;
wire v_2488;
wire v_2489;
wire v_2490;
wire v_2491;
wire v_2492;
wire v_2493;
wire v_2494;
wire v_2495;
wire v_2496;
wire v_2497;
wire v_2498;
wire v_2499;
wire v_2500;
wire v_2501;
wire v_2502;
wire v_2503;
wire v_2504;
wire v_2505;
wire v_2506;
wire v_2507;
wire v_2508;
wire v_2509;
wire v_2510;
wire v_2511;
wire v_2512;
wire v_2513;
wire v_2514;
wire v_2515;
wire v_2516;
wire v_2517;
wire v_2518;
wire v_2519;
wire v_2520;
wire v_2521;
wire v_2522;
wire v_2523;
wire v_2524;
wire v_2525;
wire v_2526;
wire v_2527;
wire v_2528;
wire v_2529;
wire v_2530;
wire v_2531;
wire v_2532;
wire v_2533;
wire v_2534;
wire v_2535;
wire v_2536;
wire v_2537;
wire v_2538;
wire v_2539;
wire v_2540;
wire v_2541;
wire v_2542;
wire v_2543;
wire v_2544;
wire v_2545;
wire v_2546;
wire v_2547;
wire v_2548;
wire v_2549;
wire v_2550;
wire v_2551;
wire v_2552;
wire v_2553;
wire v_2554;
wire v_2555;
wire v_2556;
wire v_2557;
wire v_2558;
wire v_2559;
wire v_2560;
wire v_2561;
wire v_2562;
wire v_2563;
wire v_2564;
wire v_2565;
wire v_2566;
wire v_2567;
wire v_2568;
wire v_2569;
wire v_2570;
wire v_2571;
wire v_2572;
wire v_2573;
wire v_2574;
wire v_2575;
wire v_2576;
wire v_2577;
wire v_2578;
wire v_2579;
wire v_2580;
wire v_2581;
wire v_2582;
wire v_2583;
wire v_2584;
wire v_2585;
wire v_2586;
wire v_2587;
wire v_2588;
wire v_2589;
wire v_2590;
wire v_2591;
wire v_2592;
wire v_2593;
wire v_2594;
wire v_2595;
wire v_2596;
wire v_2597;
wire v_2598;
wire v_2599;
wire v_2600;
wire v_2601;
wire v_2602;
wire v_2603;
wire v_2604;
wire v_2605;
wire v_2606;
wire v_2607;
wire v_2608;
wire v_2609;
wire v_2610;
wire v_2611;
wire v_2612;
wire v_2613;
wire v_2614;
wire v_2615;
wire v_2616;
wire v_2617;
wire v_2618;
wire v_2619;
wire v_2620;
wire v_2621;
wire v_2622;
wire v_2623;
wire v_2624;
wire v_2625;
wire v_2626;
wire v_2627;
wire v_2628;
wire v_2629;
wire v_2630;
wire v_2631;
wire v_2632;
wire v_2633;
wire v_2634;
wire v_2635;
wire v_2636;
wire v_2637;
wire v_2638;
wire v_2639;
wire v_2640;
wire v_2641;
wire v_2642;
wire v_2643;
wire v_2644;
wire v_2645;
wire v_2646;
wire v_2647;
wire v_2648;
wire v_2649;
wire v_2650;
wire v_2651;
wire v_2652;
wire v_2653;
wire v_2654;
wire v_2655;
wire v_2656;
wire v_2657;
wire v_2658;
wire v_2659;
wire v_2660;
wire v_2661;
wire v_2662;
wire v_2663;
wire v_2664;
wire v_2665;
wire v_2666;
wire v_2667;
wire v_2668;
wire v_2669;
wire v_2670;
wire v_2671;
wire v_2672;
wire v_2673;
wire v_2674;
wire v_2675;
wire v_2676;
wire v_2677;
wire v_2678;
wire v_2679;
wire v_2680;
wire v_2681;
wire v_2682;
wire v_2683;
wire v_2684;
wire v_2685;
wire v_2686;
wire v_2687;
wire v_2688;
wire v_2689;
wire v_2690;
wire v_2691;
wire v_2692;
wire v_2693;
wire v_2694;
wire v_2695;
wire v_2696;
wire v_2697;
wire v_2698;
wire v_2699;
wire v_2700;
wire v_2701;
wire v_2702;
wire v_2703;
wire v_2704;
wire v_2705;
wire v_2706;
wire v_2707;
wire v_2708;
wire v_2709;
wire v_2710;
wire v_2711;
wire v_2712;
wire v_2713;
wire v_2714;
wire v_2715;
wire v_2716;
wire v_2717;
wire v_2718;
wire v_2719;
wire v_2720;
wire v_2721;
wire v_2722;
wire v_2723;
wire v_2724;
wire v_2725;
wire v_2726;
wire v_2727;
wire v_2728;
wire v_2729;
wire v_2730;
wire v_2731;
wire v_2732;
wire v_2733;
wire v_2734;
wire v_2735;
wire v_2736;
wire v_2737;
wire v_2738;
wire v_2739;
wire v_2740;
wire v_2741;
wire v_2742;
wire v_2743;
wire v_2745;
wire v_2746;
wire v_2747;
wire v_2748;
wire v_2749;
wire v_2750;
wire v_2751;
wire v_2752;
wire v_2753;
wire v_2754;
wire v_2755;
wire v_2756;
wire v_2757;
wire v_2758;
wire v_2759;
wire v_2760;
wire v_2761;
wire v_2762;
wire v_2763;
wire v_2765;
wire v_2766;
wire v_2767;
wire v_2768;
wire v_2769;
wire v_2770;
wire v_2771;
wire v_2772;
wire v_2773;
wire v_2774;
wire v_2775;
wire v_2776;
wire v_2777;
wire v_2778;
wire v_2779;
wire v_2780;
wire v_2781;
wire v_2782;
wire v_2783;
wire v_2784;
wire v_2785;
wire v_2786;
wire v_2787;
wire v_2788;
wire v_2789;
wire v_2790;
wire v_2791;
wire v_2792;
wire v_2793;
wire v_2794;
wire v_2795;
wire v_2796;
wire v_2797;
wire v_2798;
wire v_2799;
wire v_2800;
wire v_2801;
wire v_2802;
wire v_2803;
wire v_2804;
wire v_2805;
wire v_2806;
wire v_2807;
wire v_2808;
wire v_2809;
wire v_2810;
wire v_2811;
wire v_2812;
wire v_2813;
wire v_2814;
wire v_2816;
wire v_2817;
wire v_2818;
wire v_2819;
wire v_2820;
wire v_2821;
wire v_2822;
wire v_2823;
wire v_2824;
wire v_2825;
wire v_2826;
wire v_2827;
wire v_2828;
wire v_2829;
wire v_2830;
wire v_2831;
wire v_2832;
wire v_2834;
wire v_2835;
wire v_2836;
wire v_2837;
wire v_2838;
wire v_2839;
wire v_2840;
wire v_2841;
wire v_2842;
wire v_2843;
wire v_2844;
wire v_2845;
wire v_2846;
wire v_2847;
wire v_2848;
wire v_2849;
wire v_2850;
wire v_2851;
wire v_2852;
wire v_2853;
wire v_2854;
wire v_2855;
wire v_2856;
wire v_2857;
wire v_2858;
wire v_2859;
wire v_2860;
wire v_2861;
wire v_2862;
wire v_2863;
wire v_2864;
wire v_2865;
wire v_2866;
wire v_2867;
wire v_2868;
wire v_2869;
wire v_2870;
wire v_2871;
wire v_2872;
wire v_2873;
wire v_2874;
wire v_2875;
wire v_2876;
wire v_2877;
wire v_2878;
wire v_2879;
wire v_2880;
wire v_2881;
wire v_2882;
wire v_2883;
wire v_2884;
wire v_2885;
wire v_2886;
wire v_2887;
wire v_2888;
wire v_2889;
wire v_2890;
wire v_2891;
wire v_2892;
wire v_2893;
wire v_2894;
wire v_2895;
wire v_2896;
wire v_2897;
wire v_2898;
wire v_2899;
wire v_2900;
wire v_2901;
wire v_2902;
wire v_2903;
wire v_2904;
wire v_2905;
wire v_2906;
wire v_2907;
wire v_2908;
wire v_2909;
wire v_2910;
wire v_2911;
wire v_2912;
wire v_2913;
wire v_2914;
wire v_2915;
wire v_2916;
wire v_2917;
wire v_2918;
wire v_2919;
wire v_2920;
wire v_2921;
wire v_2922;
wire v_2923;
wire v_2924;
wire v_2925;
wire v_2926;
wire v_2927;
wire v_2928;
wire v_2929;
wire v_2930;
wire v_2931;
wire v_2932;
wire v_2933;
wire v_2934;
wire v_2935;
wire v_2936;
wire v_2937;
wire v_2938;
wire v_2939;
wire v_2940;
wire v_2941;
wire v_2942;
wire v_2943;
wire v_2944;
wire v_2945;
wire v_2946;
wire v_2947;
wire v_2948;
wire v_2949;
wire v_2950;
wire v_2951;
wire v_2952;
wire v_2953;
wire v_2954;
wire v_2955;
wire v_2956;
wire v_2957;
wire v_2958;
wire v_2959;
wire v_2960;
wire v_2961;
wire v_2962;
wire v_2963;
wire v_2964;
wire v_2965;
wire v_2966;
wire v_2967;
wire v_2968;
wire v_2969;
wire v_2970;
wire v_2971;
wire v_2972;
wire v_2973;
wire v_2974;
wire v_2975;
wire v_2976;
wire v_2977;
wire v_2978;
wire v_2979;
wire v_2980;
wire v_2981;
wire v_2982;
wire v_2983;
wire v_2984;
wire v_2985;
wire v_2986;
wire v_2987;
wire v_2988;
wire v_2989;
wire v_2990;
wire v_2991;
wire v_2992;
wire v_2993;
wire v_2994;
wire v_2995;
wire v_2996;
wire v_2997;
wire v_2998;
wire v_2999;
wire v_3000;
wire v_3001;
wire v_3002;
wire v_3003;
wire v_3004;
wire v_3005;
wire v_3006;
wire v_3007;
wire v_3008;
wire v_3009;
wire v_3010;
wire v_3011;
wire v_3012;
wire v_3013;
wire v_3014;
wire v_3015;
wire v_3016;
wire v_3017;
wire v_3018;
wire v_3019;
wire v_3020;
wire v_3021;
wire v_3022;
wire v_3023;
wire v_3024;
wire v_3025;
wire v_3026;
wire v_3027;
wire v_3028;
wire v_3029;
wire v_3030;
wire v_3031;
wire v_3032;
wire v_3033;
wire v_3034;
wire v_3035;
wire v_3036;
wire v_3037;
wire v_3038;
wire v_3039;
wire v_3040;
wire v_3041;
wire v_3042;
wire v_3043;
wire v_3044;
wire v_3045;
wire v_3046;
wire v_3047;
wire v_3048;
wire v_3049;
wire v_3050;
wire v_3051;
wire v_3052;
wire v_3053;
wire v_3054;
wire v_3055;
wire v_3056;
wire v_3057;
wire v_3058;
wire v_3059;
wire v_3060;
wire v_3061;
wire v_3062;
wire v_3063;
wire v_3064;
wire v_3065;
wire v_3066;
wire v_3067;
wire v_3068;
wire v_3069;
wire v_3070;
wire v_3071;
wire v_3072;
wire v_3073;
wire v_3074;
wire v_3075;
wire v_3076;
wire v_3077;
wire v_3078;
wire v_3079;
wire v_3080;
wire v_3081;
wire v_3082;
wire v_3083;
wire v_3084;
wire v_3085;
wire v_3086;
wire v_3087;
wire v_3088;
wire v_3089;
wire v_3090;
wire v_3091;
wire v_3092;
wire v_3093;
wire v_3094;
wire v_3095;
wire v_3096;
wire v_3097;
wire v_3098;
wire v_3099;
wire v_3100;
wire v_3101;
wire v_3102;
wire v_3103;
wire v_3104;
wire v_3105;
wire v_3106;
wire v_3107;
wire v_3108;
wire v_3109;
wire v_3110;
wire v_3111;
wire v_3112;
wire v_3113;
wire v_3114;
wire v_3115;
wire v_3116;
wire v_3117;
wire v_3118;
wire v_3119;
wire v_3120;
wire v_3121;
wire v_3122;
wire v_3123;
wire v_3124;
wire v_3125;
wire v_3126;
wire v_3127;
wire v_3128;
wire v_3129;
wire v_3130;
wire v_3131;
wire v_3132;
wire v_3133;
wire v_3134;
wire v_3135;
wire v_3136;
wire v_3137;
wire v_3138;
wire v_3139;
wire v_3140;
wire v_3141;
wire v_3142;
wire v_3143;
wire v_3144;
wire v_3145;
wire v_3146;
wire v_3147;
wire v_3148;
wire v_3149;
wire v_3150;
wire v_3151;
wire v_3152;
wire v_3153;
wire v_3154;
wire v_3155;
wire v_3156;
wire v_3157;
wire v_3158;
wire v_3159;
wire v_3160;
wire v_3161;
wire v_3162;
wire v_3163;
wire v_3164;
wire v_3165;
wire v_3166;
wire v_3167;
wire v_3168;
wire v_3169;
wire v_3170;
wire v_3171;
wire v_3172;
wire v_3173;
wire v_3174;
wire v_3175;
wire v_3176;
wire v_3177;
wire v_3178;
wire v_3179;
wire v_3180;
wire v_3181;
wire v_3182;
wire v_3183;
wire v_3184;
wire v_3185;
wire v_3186;
wire v_3187;
wire v_3188;
wire v_3189;
wire v_3190;
wire v_3191;
wire v_3192;
wire v_3193;
wire v_3194;
wire v_3195;
wire v_3196;
wire v_3197;
wire v_3198;
wire v_3199;
wire v_3200;
wire v_3201;
wire v_3202;
wire v_3203;
wire v_3204;
wire v_3205;
wire v_3206;
wire v_3207;
wire v_3208;
wire v_3209;
wire v_3210;
wire v_3211;
wire v_3212;
wire v_3213;
wire v_3214;
wire v_3215;
wire v_3216;
wire v_3217;
wire v_3218;
wire v_3219;
wire v_3220;
wire v_3221;
wire v_3222;
wire v_3223;
wire v_3224;
wire v_3225;
wire v_3226;
wire v_3227;
wire v_3228;
wire v_3229;
wire v_3230;
wire v_3231;
wire v_3232;
wire v_3233;
wire v_3234;
wire v_3235;
wire v_3236;
wire v_3237;
wire v_3238;
wire v_3239;
wire v_3240;
wire v_3241;
wire v_3242;
wire v_3243;
wire v_3244;
wire v_3245;
wire v_3246;
wire v_3247;
wire v_3248;
wire v_3249;
wire v_3250;
wire v_3251;
wire v_3252;
wire v_3253;
wire v_3254;
wire v_3255;
wire v_3256;
wire v_3257;
wire v_3258;
wire v_3259;
wire v_3260;
wire v_3261;
wire v_3262;
wire v_3263;
wire v_3264;
wire v_3265;
wire v_3266;
wire v_3267;
wire v_3268;
wire v_3269;
wire v_3270;
wire v_3271;
wire v_3272;
wire v_3273;
wire v_3274;
wire v_3275;
wire v_3276;
wire v_3278;
wire v_3279;
wire v_3280;
wire v_3281;
wire v_3282;
wire v_3283;
wire v_3284;
wire v_3285;
wire v_3286;
wire v_3287;
wire v_3288;
wire v_3289;
wire v_3290;
wire v_3291;
wire v_3292;
wire v_3293;
wire v_3294;
wire v_3295;
wire v_3296;
wire v_3298;
wire v_3299;
wire v_3300;
wire v_3301;
wire v_3302;
wire v_3303;
wire v_3304;
wire v_3305;
wire v_3306;
wire v_3307;
wire v_3308;
wire v_3309;
wire v_3310;
wire v_3311;
wire v_3312;
wire v_3313;
wire v_3314;
wire v_3315;
wire v_3316;
wire v_3317;
wire v_3318;
wire v_3319;
wire v_3320;
wire v_3321;
wire v_3322;
wire v_3323;
wire v_3324;
wire v_3325;
wire v_3326;
wire v_3327;
wire v_3328;
wire v_3329;
wire v_3330;
wire v_3331;
wire v_3332;
wire v_3333;
wire v_3334;
wire v_3335;
wire v_3336;
wire v_3337;
wire v_3338;
wire v_3339;
wire v_3340;
wire v_3341;
wire v_3342;
wire v_3343;
wire v_3344;
wire v_3345;
wire v_3346;
wire v_3347;
wire v_3349;
wire v_3350;
wire v_3351;
wire v_3352;
wire v_3353;
wire v_3354;
wire v_3355;
wire v_3356;
wire v_3357;
wire v_3358;
wire v_3359;
wire v_3360;
wire v_3361;
wire v_3362;
wire v_3363;
wire v_3364;
wire v_3365;
wire v_3367;
wire v_3368;
wire v_3369;
wire v_3370;
wire v_3371;
wire v_3372;
wire v_3373;
wire v_3374;
wire v_3375;
wire v_3376;
wire v_3377;
wire v_3378;
wire v_3379;
wire v_3380;
wire v_3381;
wire v_3382;
wire v_3383;
wire v_3384;
wire v_3385;
wire v_3386;
wire v_3387;
wire v_3388;
wire v_3389;
wire v_3390;
wire v_3391;
wire v_3392;
wire v_3393;
wire v_3394;
wire v_3395;
wire v_3396;
wire v_3397;
wire v_3398;
wire v_3399;
wire v_3400;
wire v_3401;
wire v_3402;
wire v_3403;
wire v_3404;
wire v_3405;
wire v_3406;
wire v_3407;
wire v_3408;
wire v_3409;
wire v_3410;
wire v_3411;
wire v_3412;
wire v_3413;
wire v_3414;
wire v_3415;
wire v_3416;
wire v_3417;
wire v_3418;
wire v_3419;
wire v_3420;
wire v_3421;
wire v_3422;
wire v_3423;
wire v_3424;
wire v_3425;
wire v_3426;
wire v_3427;
wire v_3428;
wire v_3429;
wire v_3430;
wire v_3431;
wire v_3432;
wire v_3433;
wire v_3434;
wire v_3435;
wire v_3436;
wire v_3437;
wire v_3438;
wire v_3439;
wire v_3440;
wire v_3441;
wire v_3442;
wire v_3443;
wire v_3444;
wire v_3445;
wire v_3446;
wire v_3447;
wire v_3448;
wire v_3449;
wire v_3450;
wire v_3451;
wire v_3452;
wire v_3453;
wire v_3454;
wire v_3455;
wire v_3456;
wire v_3457;
wire v_3458;
wire v_3459;
wire v_3460;
wire v_3461;
wire v_3462;
wire v_3463;
wire v_3464;
wire v_3465;
wire v_3466;
wire v_3467;
wire v_3468;
wire v_3469;
wire v_3470;
wire v_3471;
wire v_3472;
wire v_3473;
wire v_3474;
wire v_3475;
wire v_3476;
wire v_3477;
wire v_3478;
wire v_3479;
wire v_3480;
wire v_3481;
wire v_3482;
wire v_3483;
wire v_3484;
wire v_3485;
wire v_3486;
wire v_3487;
wire v_3488;
wire v_3489;
wire v_3490;
wire v_3491;
wire v_3492;
wire v_3493;
wire v_3494;
wire v_3495;
wire v_3496;
wire v_3497;
wire v_3498;
wire v_3499;
wire v_3500;
wire v_3501;
wire v_3502;
wire v_3503;
wire v_3504;
wire v_3505;
wire v_3506;
wire v_3507;
wire v_3508;
wire v_3509;
wire v_3510;
wire v_3511;
wire v_3512;
wire v_3513;
wire v_3514;
wire v_3515;
wire v_3516;
wire v_3517;
wire v_3518;
wire v_3519;
wire v_3520;
wire v_3521;
wire v_3522;
wire v_3523;
wire v_3524;
wire v_3525;
wire v_3526;
wire v_3527;
wire v_3528;
wire v_3529;
wire v_3530;
wire v_3531;
wire v_3532;
wire v_3533;
wire v_3534;
wire v_3535;
wire v_3536;
wire v_3537;
wire v_3538;
wire v_3539;
wire v_3540;
wire v_3541;
wire v_3542;
wire v_3543;
wire v_3544;
wire v_3545;
wire v_3546;
wire v_3547;
wire v_3548;
wire v_3549;
wire v_3550;
wire v_3551;
wire v_3552;
wire v_3553;
wire v_3554;
wire v_3555;
wire v_3556;
wire v_3557;
wire v_3558;
wire v_3559;
wire v_3560;
wire v_3561;
wire v_3562;
wire v_3563;
wire v_3564;
wire v_3565;
wire v_3566;
wire v_3567;
wire v_3568;
wire v_3569;
wire v_3570;
wire v_3571;
wire v_3572;
wire v_3573;
wire v_3574;
wire v_3575;
wire v_3576;
wire v_3577;
wire v_3578;
wire v_3579;
wire v_3580;
wire v_3581;
wire v_3582;
wire v_3583;
wire v_3584;
wire v_3585;
wire v_3586;
wire v_3587;
wire v_3588;
wire v_3589;
wire v_3590;
wire v_3591;
wire v_3592;
wire v_3593;
wire v_3594;
wire v_3595;
wire v_3596;
wire v_3597;
wire v_3598;
wire v_3599;
wire v_3600;
wire v_3601;
wire v_3602;
wire v_3603;
wire v_3604;
wire v_3605;
wire v_3606;
wire v_3607;
wire v_3608;
wire v_3609;
wire v_3610;
wire v_3611;
wire v_3612;
wire v_3613;
wire v_3614;
wire v_3615;
wire v_3616;
wire v_3617;
wire v_3618;
wire v_3619;
wire v_3620;
wire v_3621;
wire v_3622;
wire v_3623;
wire v_3624;
wire v_3625;
wire v_3626;
wire v_3627;
wire v_3628;
wire v_3629;
wire v_3630;
wire v_3631;
wire v_3632;
wire v_3633;
wire v_3634;
wire v_3635;
wire v_3636;
wire v_3637;
wire v_3638;
wire v_3639;
wire v_3640;
wire v_3641;
wire v_3642;
wire v_3643;
wire v_3644;
wire v_3645;
wire v_3646;
wire v_3647;
wire v_3648;
wire v_3649;
wire v_3650;
wire v_3651;
wire v_3652;
wire v_3653;
wire v_3654;
wire v_3655;
wire v_3656;
wire v_3657;
wire v_3658;
wire v_3659;
wire v_3660;
wire v_3661;
wire v_3662;
wire v_3663;
wire v_3664;
wire v_3665;
wire v_3666;
wire v_3667;
wire v_3668;
wire v_3669;
wire v_3670;
wire v_3671;
wire v_3672;
wire v_3673;
wire v_3674;
wire v_3675;
wire v_3676;
wire v_3677;
wire v_3678;
wire v_3679;
wire v_3680;
wire v_3681;
wire v_3682;
wire v_3683;
wire v_3684;
wire v_3685;
wire v_3686;
wire v_3687;
wire v_3689;
wire v_3690;
wire v_3691;
wire v_3692;
wire v_3693;
wire v_3694;
wire v_3695;
wire v_3696;
wire v_3697;
wire v_3698;
wire v_3699;
wire v_3700;
wire v_3701;
wire v_3702;
wire v_3703;
wire v_3704;
wire v_3705;
wire v_3706;
wire v_3707;
wire v_3708;
wire v_3709;
wire v_3710;
wire v_3711;
wire v_3712;
wire v_3713;
wire v_3714;
wire v_3715;
wire v_3716;
wire v_3717;
wire v_3718;
wire v_3719;
wire v_3720;
wire v_3721;
wire v_3722;
wire v_3723;
wire v_3724;
wire v_3725;
wire v_3726;
wire v_3727;
wire v_3728;
wire v_3729;
wire v_3730;
wire v_3731;
wire v_3732;
wire v_3733;
wire v_3734;
wire v_3735;
wire v_3736;
wire v_3737;
wire v_3738;
wire v_3739;
wire v_3740;
wire v_3741;
wire v_3742;
wire v_3743;
wire v_3744;
wire v_3745;
wire v_3746;
wire v_3747;
wire v_3748;
wire v_3749;
wire v_3750;
wire v_3751;
wire v_3752;
wire v_3753;
wire v_3754;
wire v_3755;
wire v_3756;
wire v_3757;
wire v_3758;
wire v_3759;
wire v_3760;
wire v_3761;
wire v_3762;
wire v_3763;
wire v_3764;
wire v_3765;
wire v_3766;
wire v_3767;
wire v_3768;
wire v_3769;
wire v_3770;
wire v_3771;
wire v_3772;
wire v_3773;
wire v_3774;
wire v_3775;
wire v_3776;
wire v_3777;
wire v_3778;
wire v_3779;
wire v_3780;
wire v_3781;
wire v_3782;
wire v_3783;
wire v_3784;
wire v_3785;
wire v_3786;
wire v_3787;
wire v_3788;
wire v_3789;
wire v_3790;
wire v_3791;
wire v_3792;
wire v_3793;
wire v_3794;
wire v_3795;
wire v_3796;
wire v_3797;
wire v_3798;
wire v_3799;
wire v_3800;
wire v_3801;
wire v_3802;
wire v_3803;
wire v_3804;
wire v_3805;
wire v_3806;
wire v_3807;
wire v_3808;
wire v_3809;
wire v_3810;
wire v_3811;
wire v_3812;
wire v_3814;
wire v_3815;
wire v_3816;
wire v_3817;
wire v_3818;
wire v_3819;
wire v_3820;
wire v_3821;
wire v_3822;
wire v_3823;
wire v_3824;
wire v_3825;
wire v_3826;
wire v_3827;
wire v_3828;
wire v_3829;
wire v_3830;
wire v_3831;
wire v_3832;
wire v_3834;
wire v_3835;
wire v_3836;
wire v_3837;
wire v_3838;
wire v_3839;
wire v_3840;
wire v_3841;
wire v_3842;
wire v_3843;
wire v_3844;
wire v_3845;
wire v_3846;
wire v_3847;
wire v_3848;
wire v_3849;
wire v_3850;
wire v_3851;
wire v_3852;
wire v_3853;
wire v_3854;
wire v_3855;
wire v_3856;
wire v_3857;
wire v_3858;
wire v_3859;
wire v_3860;
wire v_3861;
wire v_3862;
wire v_3863;
wire v_3864;
wire v_3865;
wire v_3866;
wire v_3867;
wire v_3868;
wire v_3869;
wire v_3870;
wire v_3871;
wire v_3872;
wire v_3873;
wire v_3874;
wire v_3875;
wire v_3876;
wire v_3877;
wire v_3878;
wire v_3879;
wire v_3880;
wire v_3881;
wire v_3882;
wire v_3883;
wire v_3885;
wire v_3886;
wire v_3887;
wire v_3888;
wire v_3889;
wire v_3890;
wire v_3891;
wire v_3892;
wire v_3893;
wire v_3894;
wire v_3895;
wire v_3896;
wire v_3897;
wire v_3898;
wire v_3899;
wire v_3900;
wire v_3901;
wire v_3903;
wire v_3904;
wire v_3905;
wire v_3906;
wire v_3907;
wire v_3908;
wire v_3909;
wire v_3910;
wire v_3911;
wire v_3912;
wire v_3913;
wire v_3914;
wire v_3915;
wire v_3916;
wire v_3917;
wire v_3918;
wire v_3919;
wire v_3920;
wire v_3921;
wire v_3922;
wire v_3923;
wire v_3924;
wire v_3925;
wire v_3926;
wire v_3927;
wire v_3928;
wire v_3929;
wire v_3930;
wire v_3931;
wire v_3932;
wire v_3933;
wire v_3934;
wire v_3935;
wire v_3936;
wire v_3937;
wire v_3938;
wire v_3939;
wire v_3940;
wire v_3941;
wire v_3942;
wire v_3943;
wire v_3944;
wire v_3945;
wire v_3946;
wire v_3947;
wire v_3948;
wire v_3949;
wire v_3950;
wire v_3951;
wire v_3952;
wire v_3953;
wire v_3954;
wire v_3955;
wire v_3956;
wire v_3957;
wire v_3958;
wire v_3959;
wire v_3960;
wire v_3961;
wire v_3962;
wire v_3963;
wire v_3964;
wire v_3965;
wire v_3966;
wire v_3967;
wire v_3968;
wire v_3969;
wire v_3970;
wire v_3971;
wire v_3972;
wire v_3973;
wire v_3974;
wire v_3975;
wire v_3976;
wire v_3977;
wire v_3978;
wire v_3979;
wire v_3980;
wire v_3981;
wire v_3982;
wire v_3983;
wire v_3984;
wire v_3985;
wire v_3986;
wire v_3987;
wire v_3988;
wire v_3989;
wire v_3990;
wire v_3991;
wire v_3992;
wire v_3993;
wire v_3994;
wire v_3995;
wire v_3996;
wire v_3997;
wire v_3998;
wire v_3999;
wire v_4000;
wire v_4001;
wire v_4002;
wire v_4003;
wire v_4004;
wire v_4005;
wire v_4006;
wire v_4007;
wire v_4008;
wire v_4009;
wire v_4010;
wire v_4011;
wire v_4012;
wire v_4013;
wire v_4014;
wire v_4015;
wire v_4016;
wire v_4017;
wire v_4018;
wire v_4019;
wire v_4020;
wire v_4021;
wire v_4022;
wire v_4023;
wire v_4024;
wire v_4025;
wire v_4026;
wire v_4027;
wire v_4028;
wire v_4029;
wire v_4030;
wire v_4031;
wire v_4032;
wire v_4033;
wire v_4034;
wire v_4035;
wire v_4036;
wire v_4037;
wire v_4038;
wire v_4039;
wire v_4040;
wire v_4041;
wire v_4042;
wire v_4043;
wire v_4044;
wire v_4045;
wire v_4046;
wire v_4047;
wire v_4048;
wire v_4049;
wire v_4050;
wire v_4051;
wire v_4052;
wire v_4053;
wire v_4054;
wire v_4055;
wire v_4056;
wire v_4057;
wire v_4058;
wire v_4059;
wire v_4060;
wire v_4061;
wire v_4062;
wire v_4063;
wire v_4064;
wire v_4065;
wire v_4066;
wire v_4067;
wire v_4068;
wire v_4069;
wire v_4070;
wire v_4071;
wire v_4072;
wire v_4073;
wire v_4074;
wire v_4075;
wire v_4076;
wire v_4077;
wire v_4078;
wire v_4079;
wire v_4080;
wire v_4081;
wire v_4082;
wire v_4083;
wire v_4084;
wire v_4085;
wire v_4086;
wire v_4087;
wire v_4088;
wire v_4089;
wire v_4090;
wire v_4091;
wire v_4092;
wire v_4093;
wire v_4094;
wire v_4095;
wire v_4096;
wire v_4097;
wire v_4098;
wire v_4099;
wire v_4100;
wire v_4101;
wire v_4102;
wire v_4103;
wire v_4104;
wire v_4105;
wire v_4106;
wire v_4107;
wire v_4108;
wire v_4109;
wire v_4110;
wire v_4111;
wire v_4112;
wire v_4113;
wire v_4114;
wire v_4115;
wire v_4116;
wire v_4117;
wire v_4118;
wire v_4119;
wire v_4120;
wire v_4121;
wire v_4122;
wire v_4123;
wire v_4124;
wire v_4125;
wire v_4126;
wire v_4127;
wire v_4128;
wire v_4129;
wire v_4130;
wire v_4131;
wire v_4132;
wire v_4133;
wire v_4134;
wire v_4135;
wire v_4136;
wire v_4137;
wire v_4138;
wire v_4139;
wire v_4140;
wire v_4141;
wire v_4142;
wire v_4143;
wire v_4144;
wire v_4145;
wire v_4146;
wire v_4147;
wire v_4148;
wire v_4149;
wire v_4150;
wire v_4151;
wire v_4152;
wire v_4153;
wire v_4154;
wire v_4155;
wire v_4156;
wire v_4157;
wire v_4158;
wire v_4159;
wire v_4160;
wire v_4161;
wire v_4162;
wire v_4163;
wire v_4164;
wire v_4165;
wire v_4166;
wire v_4167;
wire v_4168;
wire v_4169;
wire v_4170;
wire v_4171;
wire v_4172;
wire v_4173;
wire v_4174;
wire v_4175;
wire v_4176;
wire v_4177;
wire v_4178;
wire v_4179;
wire v_4180;
wire v_4181;
wire v_4182;
wire v_4183;
wire v_4184;
wire v_4185;
wire v_4186;
wire v_4187;
wire v_4188;
wire v_4189;
wire v_4190;
wire v_4191;
wire v_4192;
wire v_4193;
wire v_4194;
wire v_4195;
wire v_4196;
wire v_4197;
wire v_4198;
wire v_4199;
wire v_4200;
wire v_4201;
wire v_4202;
wire v_4203;
wire v_4204;
wire v_4205;
wire v_4206;
wire v_4207;
wire v_4208;
wire v_4209;
wire v_4210;
wire v_4211;
wire v_4212;
wire v_4213;
wire v_4214;
wire v_4215;
wire v_4216;
wire v_4217;
wire v_4218;
wire v_4219;
wire v_4220;
wire v_4221;
wire v_4222;
wire v_4223;
wire v_4225;
wire v_4226;
wire v_4227;
wire v_4228;
wire v_4229;
wire v_4230;
wire v_4231;
wire v_4232;
wire v_4233;
wire v_4234;
wire v_4235;
wire v_4236;
wire v_4237;
wire v_4238;
wire v_4239;
wire v_4240;
wire v_4241;
wire v_4242;
wire v_4243;
wire v_4244;
wire v_4245;
wire v_4246;
wire v_4247;
wire v_4248;
wire v_4249;
wire v_4250;
wire v_4251;
wire v_4252;
wire v_4253;
wire v_4254;
wire v_4255;
wire v_4256;
wire v_4257;
wire v_4258;
wire v_4259;
wire v_4260;
wire v_4261;
wire v_4262;
wire v_4263;
wire v_4264;
wire v_4265;
wire v_4266;
wire v_4267;
wire v_4268;
wire v_4269;
wire v_4270;
wire v_4271;
wire v_4272;
wire v_4273;
wire v_4274;
wire v_4275;
wire v_4276;
wire v_4277;
wire v_4278;
wire v_4279;
wire v_4280;
wire v_4281;
wire v_4282;
wire v_4283;
wire v_4284;
wire v_4285;
wire v_4286;
wire v_4287;
wire v_4288;
wire v_4289;
wire v_4290;
wire v_4291;
wire v_4292;
wire v_4293;
wire v_4294;
wire v_4295;
wire v_4296;
wire v_4297;
wire v_4298;
wire v_4299;
wire v_4300;
wire v_4301;
wire v_4302;
wire v_4303;
wire v_4304;
wire v_4305;
wire v_4306;
wire v_4307;
wire v_4308;
wire v_4309;
wire v_4310;
wire v_4311;
wire v_4312;
wire v_4313;
wire v_4314;
wire v_4315;
wire v_4316;
wire v_4317;
wire v_4318;
wire v_4319;
wire v_4320;
wire v_4321;
wire v_4322;
wire v_4323;
wire v_4324;
wire v_4325;
wire v_4326;
wire v_4327;
wire v_4328;
wire v_4329;
wire v_4330;
wire v_4331;
wire v_4332;
wire v_4333;
wire v_4334;
wire v_4335;
wire v_4336;
wire v_4337;
wire v_4338;
wire v_4339;
wire v_4340;
wire v_4341;
wire v_4342;
wire v_4343;
wire v_4344;
wire v_4345;
wire v_4346;
wire v_4347;
wire v_4348;
wire v_4350;
wire v_4351;
wire v_4352;
wire v_4353;
wire v_4354;
wire v_4355;
wire v_4356;
wire v_4357;
wire v_4358;
wire v_4359;
wire v_4360;
wire v_4361;
wire v_4362;
wire v_4363;
wire v_4364;
wire v_4365;
wire v_4366;
wire v_4367;
wire v_4368;
wire v_4370;
wire v_4371;
wire v_4372;
wire v_4373;
wire v_4374;
wire v_4375;
wire v_4376;
wire v_4377;
wire v_4378;
wire v_4379;
wire v_4380;
wire v_4381;
wire v_4382;
wire v_4383;
wire v_4384;
wire v_4385;
wire v_4386;
wire v_4387;
wire v_4388;
wire v_4389;
wire v_4390;
wire v_4391;
wire v_4392;
wire v_4393;
wire v_4394;
wire v_4395;
wire v_4396;
wire v_4397;
wire v_4398;
wire v_4399;
wire v_4400;
wire v_4401;
wire v_4402;
wire v_4403;
wire v_4404;
wire v_4405;
wire v_4406;
wire v_4407;
wire v_4408;
wire v_4409;
wire v_4410;
wire v_4411;
wire v_4412;
wire v_4413;
wire v_4414;
wire v_4415;
wire v_4416;
wire v_4417;
wire v_4418;
wire v_4419;
wire v_4421;
wire v_4422;
wire v_4423;
wire v_4424;
wire v_4425;
wire v_4426;
wire v_4427;
wire v_4428;
wire v_4429;
wire v_4430;
wire v_4431;
wire v_4432;
wire v_4433;
wire v_4434;
wire v_4435;
wire v_4436;
wire v_4437;
wire v_4439;
wire v_4440;
wire v_4441;
wire v_4442;
wire v_4443;
wire v_4444;
wire v_4445;
wire v_4446;
wire v_4447;
wire v_4448;
wire v_4449;
wire v_4450;
wire v_4451;
wire v_4452;
wire v_4453;
wire v_4454;
wire v_4455;
wire v_4456;
wire v_4457;
wire v_4458;
wire v_4459;
wire v_4460;
wire v_4461;
wire v_4462;
wire v_4463;
wire v_4464;
wire v_4465;
wire v_4466;
wire v_4467;
wire v_4468;
wire v_4469;
wire v_4470;
wire v_4471;
wire v_4472;
wire v_4473;
wire v_4474;
wire v_4475;
wire v_4476;
wire v_4477;
wire v_4478;
wire v_4479;
wire v_4480;
wire v_4481;
wire v_4482;
wire v_4483;
wire v_4484;
wire v_4485;
wire v_4486;
wire v_4487;
wire v_4488;
wire v_4489;
wire v_4490;
wire v_4491;
wire v_4492;
wire v_4493;
wire v_4494;
wire v_4495;
wire v_4496;
wire v_4497;
wire v_4498;
wire v_4499;
wire v_4500;
wire v_4501;
wire v_4502;
wire v_4503;
wire v_4504;
wire v_4505;
wire v_4506;
wire v_4507;
wire v_4508;
wire v_4509;
wire v_4510;
wire v_4511;
wire v_4512;
wire v_4513;
wire v_4514;
wire v_4515;
wire v_4516;
wire v_4517;
wire v_4518;
wire v_4519;
wire v_4520;
wire v_4521;
wire v_4522;
wire v_4523;
wire v_4524;
wire v_4525;
wire v_4526;
wire v_4527;
wire v_4528;
wire v_4529;
wire v_4530;
wire v_4531;
wire v_4532;
wire v_4533;
wire v_4534;
wire v_4535;
wire v_4536;
wire v_4537;
wire v_4538;
wire v_4539;
wire v_4540;
wire v_4541;
wire v_4542;
wire v_4543;
wire v_4544;
wire v_4545;
wire v_4546;
wire v_4547;
wire v_4548;
wire v_4549;
wire v_4550;
wire v_4551;
wire v_4552;
wire v_4553;
wire v_4554;
wire v_4555;
wire v_4556;
wire v_4557;
wire v_4558;
wire v_4559;
wire v_4560;
wire v_4561;
wire v_4562;
wire v_4563;
wire v_4564;
wire v_4565;
wire v_4566;
wire v_4567;
wire v_4568;
wire v_4569;
wire v_4570;
wire v_4571;
wire v_4572;
wire v_4573;
wire v_4574;
wire v_4575;
wire v_4576;
wire v_4577;
wire v_4578;
wire v_4579;
wire v_4580;
wire v_4581;
wire v_4582;
wire v_4583;
wire v_4584;
wire v_4585;
wire v_4586;
wire v_4587;
wire v_4588;
wire v_4589;
wire v_4590;
wire v_4591;
wire v_4592;
wire v_4593;
wire v_4594;
wire v_4595;
wire v_4596;
wire v_4597;
wire v_4598;
wire v_4599;
wire v_4600;
wire v_4601;
wire v_4602;
wire v_4603;
wire v_4604;
wire v_4605;
wire v_4606;
wire v_4607;
wire v_4608;
wire v_4609;
wire v_4610;
wire v_4611;
wire v_4612;
wire v_4613;
wire v_4614;
wire v_4615;
wire v_4616;
wire v_4617;
wire v_4618;
wire v_4619;
wire v_4620;
wire v_4621;
wire v_4622;
wire v_4623;
wire v_4624;
wire v_4625;
wire v_4626;
wire v_4627;
wire v_4628;
wire v_4629;
wire v_4630;
wire v_4631;
wire v_4632;
wire v_4633;
wire v_4634;
wire v_4635;
wire v_4636;
wire v_4637;
wire v_4638;
wire v_4639;
wire v_4640;
wire v_4641;
wire v_4642;
wire v_4643;
wire v_4644;
wire v_4645;
wire v_4646;
wire v_4647;
wire v_4648;
wire v_4649;
wire v_4650;
wire v_4651;
wire v_4652;
wire v_4653;
wire v_4654;
wire v_4655;
wire v_4656;
wire v_4657;
wire v_4658;
wire v_4659;
wire v_4660;
wire v_4661;
wire v_4662;
wire v_4663;
wire v_4664;
wire v_4665;
wire v_4666;
wire v_4667;
wire v_4668;
wire v_4669;
wire v_4670;
wire v_4671;
wire v_4672;
wire v_4673;
wire v_4674;
wire v_4675;
wire v_4676;
wire v_4677;
wire v_4678;
wire v_4679;
wire v_4680;
wire v_4681;
wire v_4682;
wire v_4683;
wire v_4684;
wire v_4685;
wire v_4686;
wire v_4687;
wire v_4688;
wire v_4689;
wire v_4690;
wire v_4691;
wire v_4692;
wire v_4693;
wire v_4694;
wire v_4695;
wire v_4696;
wire v_4697;
wire v_4698;
wire v_4699;
wire v_4700;
wire v_4701;
wire v_4702;
wire v_4703;
wire v_4704;
wire v_4705;
wire v_4706;
wire v_4707;
wire v_4708;
wire v_4709;
wire v_4710;
wire v_4711;
wire v_4712;
wire v_4713;
wire v_4714;
wire v_4715;
wire v_4716;
wire v_4717;
wire v_4718;
wire v_4719;
wire v_4720;
wire v_4721;
wire v_4722;
wire v_4723;
wire v_4724;
wire v_4725;
wire v_4726;
wire v_4727;
wire v_4728;
wire v_4729;
wire v_4730;
wire v_4731;
wire v_4732;
wire v_4733;
wire v_4734;
wire v_4735;
wire v_4736;
wire v_4737;
wire v_4738;
wire v_4739;
wire v_4740;
wire v_4741;
wire v_4742;
wire v_4743;
wire v_4744;
wire v_4745;
wire v_4746;
wire v_4747;
wire v_4748;
wire v_4749;
wire v_4750;
wire v_4751;
wire v_4752;
wire v_4753;
wire v_4754;
wire v_4755;
wire v_4756;
wire v_4757;
wire v_4758;
wire v_4759;
wire v_4760;
wire v_4761;
wire v_4762;
wire v_4763;
wire v_4764;
wire v_4765;
wire v_4766;
wire v_4767;
wire v_4768;
wire v_4769;
wire v_4770;
wire v_4771;
wire v_4772;
wire v_4773;
wire v_4774;
wire v_4775;
wire v_4776;
wire v_4777;
wire v_4778;
wire v_4779;
wire v_4780;
wire v_4781;
wire v_4782;
wire v_4783;
wire v_4784;
wire v_4785;
wire v_4786;
wire v_4787;
wire v_4788;
wire v_4789;
wire v_4790;
wire v_4791;
wire v_4792;
wire v_4793;
wire v_4794;
wire v_4795;
wire v_4796;
wire v_4797;
wire v_4798;
wire v_4799;
wire v_4800;
wire v_4801;
wire v_4802;
wire v_4803;
wire v_4804;
wire v_4805;
wire v_4806;
wire v_4807;
wire v_4808;
wire v_4809;
wire v_4810;
wire v_4811;
wire v_4812;
wire v_4813;
wire v_4814;
wire v_4815;
wire v_4816;
wire v_4817;
wire v_4818;
wire v_4819;
wire v_4820;
wire v_4821;
wire v_4822;
wire v_4823;
wire v_4824;
wire v_4825;
wire v_4826;
wire v_4827;
wire v_4828;
wire v_4829;
wire v_4830;
wire v_4831;
wire v_4832;
wire v_4833;
wire v_4834;
wire v_4835;
wire v_4836;
wire v_4837;
wire v_4838;
wire v_4839;
wire v_4840;
wire v_4841;
wire v_4842;
wire v_4843;
wire v_4844;
wire v_4845;
wire v_4846;
wire v_4847;
wire v_4848;
wire v_4849;
wire v_4850;
wire v_4851;
wire v_4852;
wire v_4853;
wire v_4854;
wire v_4855;
wire v_4856;
wire v_4857;
wire v_4858;
wire v_4859;
wire v_4860;
wire v_4861;
wire v_4862;
wire v_4863;
wire v_4864;
wire v_4865;
wire v_4866;
wire v_4867;
wire v_4868;
wire v_4869;
wire v_4870;
wire v_4871;
wire v_4872;
wire v_4873;
wire v_4874;
wire v_4875;
wire v_4876;
wire v_4877;
wire v_4878;
wire v_4879;
wire v_4880;
wire v_4881;
wire v_4882;
wire v_4883;
wire v_4885;
wire v_4886;
wire v_4887;
wire v_4888;
wire v_4889;
wire v_4890;
wire v_4891;
wire v_4892;
wire v_4893;
wire v_4894;
wire v_4895;
wire v_4896;
wire v_4897;
wire v_4898;
wire v_4899;
wire v_4900;
wire v_4901;
wire v_4902;
wire v_4903;
wire v_4905;
wire v_4906;
wire v_4907;
wire v_4908;
wire v_4909;
wire v_4910;
wire v_4911;
wire v_4912;
wire v_4913;
wire v_4914;
wire v_4915;
wire v_4916;
wire v_4917;
wire v_4918;
wire v_4919;
wire v_4920;
wire v_4921;
wire v_4922;
wire v_4923;
wire v_4924;
wire v_4925;
wire v_4926;
wire v_4927;
wire v_4928;
wire v_4929;
wire v_4930;
wire v_4931;
wire v_4932;
wire v_4933;
wire v_4934;
wire v_4935;
wire v_4936;
wire v_4937;
wire v_4938;
wire v_4939;
wire v_4940;
wire v_4941;
wire v_4942;
wire v_4943;
wire v_4944;
wire v_4945;
wire v_4946;
wire v_4947;
wire v_4948;
wire v_4949;
wire v_4950;
wire v_4951;
wire v_4952;
wire v_4953;
wire v_4954;
wire v_4956;
wire v_4957;
wire v_4958;
wire v_4959;
wire v_4960;
wire v_4961;
wire v_4962;
wire v_4963;
wire v_4964;
wire v_4965;
wire v_4966;
wire v_4967;
wire v_4968;
wire v_4969;
wire v_4970;
wire v_4971;
wire v_4972;
wire v_4974;
wire v_4975;
wire v_4976;
wire v_4977;
wire v_4978;
wire v_4979;
wire v_4980;
wire v_4981;
wire v_4982;
wire v_4983;
wire v_4984;
wire v_4985;
wire v_4986;
wire v_4987;
wire v_4988;
wire v_4989;
wire v_4990;
wire v_4991;
wire v_4992;
wire v_4993;
wire v_4994;
wire v_4995;
wire v_4996;
wire v_4997;
wire v_4998;
wire v_4999;
wire v_5000;
wire v_5001;
wire v_5002;
wire v_5003;
wire v_5004;
wire v_5005;
wire v_5006;
wire v_5007;
wire v_5008;
wire v_5009;
wire v_5010;
wire v_5011;
wire v_5012;
wire v_5013;
wire v_5014;
wire v_5015;
wire v_5016;
wire v_5017;
wire v_5018;
wire v_5019;
wire v_5020;
wire v_5021;
wire v_5022;
wire v_5023;
wire v_5024;
wire v_5025;
wire v_5026;
wire v_5027;
wire v_5028;
wire v_5029;
wire v_5030;
wire v_5031;
wire v_5032;
wire v_5033;
wire v_5034;
wire v_5035;
wire v_5036;
wire v_5037;
wire v_5038;
wire v_5039;
wire v_5040;
wire v_5041;
wire v_5042;
wire v_5043;
wire v_5044;
wire v_5045;
wire v_5046;
wire v_5047;
wire v_5048;
wire v_5049;
wire v_5050;
wire v_5051;
wire v_5052;
wire v_5053;
wire v_5054;
wire v_5055;
wire v_5056;
wire v_5057;
wire v_5058;
wire v_5059;
wire v_5060;
wire v_5061;
wire v_5062;
wire v_5063;
wire v_5064;
wire v_5065;
wire v_5066;
wire v_5067;
wire v_5068;
wire v_5069;
wire v_5070;
wire v_5071;
wire v_5072;
wire v_5073;
wire v_5074;
wire v_5075;
wire v_5076;
wire v_5077;
wire v_5078;
wire v_5079;
wire v_5080;
wire v_5081;
wire v_5082;
wire v_5083;
wire v_5084;
wire v_5085;
wire v_5086;
wire v_5087;
wire v_5088;
wire v_5089;
wire v_5090;
wire v_5091;
wire v_5092;
wire v_5093;
wire v_5094;
wire v_5095;
wire v_5096;
wire v_5097;
wire v_5098;
wire v_5099;
wire v_5100;
wire v_5101;
wire v_5102;
wire v_5103;
wire v_5104;
wire v_5105;
wire v_5106;
wire v_5107;
wire v_5108;
wire v_5109;
wire v_5110;
wire v_5111;
wire v_5112;
wire v_5113;
wire v_5114;
wire v_5115;
wire v_5116;
wire v_5117;
wire v_5118;
wire v_5119;
wire v_5120;
wire v_5121;
wire v_5122;
wire v_5123;
wire v_5124;
wire v_5125;
wire v_5126;
wire v_5127;
wire v_5128;
wire v_5129;
wire v_5130;
wire v_5131;
wire v_5132;
wire v_5133;
wire v_5134;
wire v_5135;
wire v_5136;
wire v_5137;
wire v_5138;
wire v_5139;
wire v_5140;
wire v_5141;
wire v_5142;
wire v_5143;
wire v_5144;
wire v_5145;
wire v_5146;
wire v_5147;
wire v_5148;
wire v_5149;
wire v_5150;
wire v_5151;
wire v_5152;
wire v_5153;
wire v_5154;
wire v_5155;
wire v_5156;
wire v_5157;
wire v_5158;
wire v_5159;
wire v_5160;
wire v_5161;
wire v_5162;
wire v_5163;
wire v_5164;
wire v_5165;
wire v_5166;
wire v_5167;
wire v_5168;
wire v_5169;
wire v_5170;
wire v_5171;
wire v_5172;
wire v_5173;
wire v_5174;
wire v_5175;
wire v_5176;
wire v_5177;
wire v_5178;
wire v_5179;
wire v_5180;
wire v_5181;
wire v_5182;
wire v_5183;
wire v_5184;
wire v_5185;
wire v_5186;
wire v_5187;
wire v_5188;
wire v_5189;
wire v_5190;
wire v_5191;
wire v_5192;
wire v_5193;
wire v_5194;
wire v_5195;
wire v_5196;
wire v_5197;
wire v_5198;
wire v_5199;
wire v_5200;
wire v_5201;
wire v_5202;
wire v_5203;
wire v_5204;
wire v_5205;
wire v_5206;
wire v_5207;
wire v_5208;
wire v_5209;
wire v_5210;
wire v_5211;
wire v_5212;
wire v_5213;
wire v_5214;
wire v_5215;
wire v_5216;
wire v_5217;
wire v_5218;
wire v_5219;
wire v_5220;
wire v_5221;
wire v_5222;
wire v_5223;
wire v_5224;
wire v_5225;
wire v_5226;
wire v_5227;
wire v_5228;
wire v_5229;
wire v_5230;
wire v_5231;
wire v_5232;
wire v_5233;
wire v_5234;
wire v_5235;
wire v_5236;
wire v_5237;
wire v_5238;
wire v_5239;
wire v_5240;
wire v_5241;
wire v_5242;
wire v_5243;
wire v_5244;
wire v_5245;
wire v_5246;
wire v_5247;
wire v_5248;
wire v_5249;
wire v_5250;
wire v_5251;
wire v_5252;
wire v_5253;
wire v_5254;
wire v_5255;
wire v_5256;
wire v_5257;
wire v_5258;
wire v_5259;
wire v_5260;
wire v_5261;
wire v_5262;
wire v_5263;
wire v_5264;
wire v_5265;
wire v_5266;
wire v_5267;
wire v_5268;
wire v_5269;
wire v_5270;
wire v_5271;
wire v_5272;
wire v_5273;
wire v_5274;
wire v_5275;
wire v_5276;
wire v_5277;
wire v_5278;
wire v_5279;
wire v_5280;
wire v_5281;
wire v_5282;
wire v_5283;
wire v_5284;
wire v_5285;
wire v_5286;
wire v_5287;
wire v_5288;
wire v_5289;
wire v_5290;
wire v_5291;
wire v_5292;
wire v_5293;
wire v_5294;
wire v_5296;
wire v_5297;
wire v_5298;
wire v_5299;
wire v_5300;
wire v_5301;
wire v_5302;
wire v_5303;
wire v_5304;
wire v_5305;
wire v_5306;
wire v_5307;
wire v_5308;
wire v_5309;
wire v_5310;
wire v_5311;
wire v_5312;
wire v_5313;
wire v_5314;
wire v_5315;
wire v_5316;
wire v_5317;
wire v_5318;
wire v_5319;
wire v_5320;
wire v_5321;
wire v_5322;
wire v_5323;
wire v_5324;
wire v_5325;
wire v_5326;
wire v_5327;
wire v_5328;
wire v_5329;
wire v_5330;
wire v_5331;
wire v_5332;
wire v_5333;
wire v_5334;
wire v_5335;
wire v_5336;
wire v_5337;
wire v_5338;
wire v_5339;
wire v_5340;
wire v_5341;
wire v_5342;
wire v_5343;
wire v_5344;
wire v_5345;
wire v_5346;
wire v_5347;
wire v_5348;
wire v_5349;
wire v_5350;
wire v_5351;
wire v_5352;
wire v_5353;
wire v_5354;
wire v_5355;
wire v_5356;
wire v_5357;
wire v_5358;
wire v_5359;
wire v_5360;
wire v_5361;
wire v_5362;
wire v_5363;
wire v_5364;
wire v_5365;
wire v_5366;
wire v_5367;
wire v_5368;
wire v_5369;
wire v_5370;
wire v_5371;
wire v_5372;
wire v_5373;
wire v_5374;
wire v_5375;
wire v_5376;
wire v_5377;
wire v_5378;
wire v_5379;
wire v_5380;
wire v_5381;
wire v_5382;
wire v_5383;
wire v_5384;
wire v_5385;
wire v_5386;
wire v_5387;
wire v_5388;
wire v_5389;
wire v_5390;
wire v_5391;
wire v_5392;
wire v_5393;
wire v_5394;
wire v_5395;
wire v_5396;
wire v_5397;
wire v_5398;
wire v_5399;
wire v_5400;
wire v_5401;
wire v_5402;
wire v_5403;
wire v_5404;
wire v_5405;
wire v_5406;
wire v_5407;
wire v_5408;
wire v_5409;
wire v_5410;
wire v_5411;
wire v_5412;
wire v_5413;
wire v_5414;
wire v_5415;
wire v_5416;
wire v_5417;
wire v_5418;
wire v_5419;
wire v_5421;
wire v_5422;
wire v_5423;
wire v_5424;
wire v_5425;
wire v_5426;
wire v_5427;
wire v_5428;
wire v_5429;
wire v_5430;
wire v_5431;
wire v_5432;
wire v_5433;
wire v_5434;
wire v_5435;
wire v_5436;
wire v_5437;
wire v_5438;
wire v_5439;
wire v_5441;
wire v_5442;
wire v_5443;
wire v_5444;
wire v_5445;
wire v_5446;
wire v_5447;
wire v_5448;
wire v_5449;
wire v_5450;
wire v_5451;
wire v_5452;
wire v_5453;
wire v_5454;
wire v_5455;
wire v_5456;
wire v_5457;
wire v_5458;
wire v_5459;
wire v_5460;
wire v_5461;
wire v_5462;
wire v_5463;
wire v_5464;
wire v_5465;
wire v_5466;
wire v_5467;
wire v_5468;
wire v_5469;
wire v_5470;
wire v_5471;
wire v_5472;
wire v_5473;
wire v_5474;
wire v_5475;
wire v_5476;
wire v_5477;
wire v_5478;
wire v_5479;
wire v_5480;
wire v_5481;
wire v_5482;
wire v_5483;
wire v_5484;
wire v_5485;
wire v_5486;
wire v_5487;
wire v_5488;
wire v_5489;
wire v_5490;
wire v_5492;
wire v_5493;
wire v_5494;
wire v_5495;
wire v_5496;
wire v_5497;
wire v_5498;
wire v_5499;
wire v_5500;
wire v_5501;
wire v_5502;
wire v_5503;
wire v_5504;
wire v_5505;
wire v_5506;
wire v_5507;
wire v_5508;
wire v_5510;
wire v_5511;
wire v_5512;
wire v_5513;
wire v_5514;
wire v_5515;
wire v_5516;
wire v_5517;
wire v_5518;
wire v_5519;
wire v_5520;
wire v_5521;
wire v_5522;
wire v_5523;
wire v_5524;
wire v_5525;
wire v_5526;
wire v_5527;
wire v_5528;
wire v_5529;
wire v_5530;
wire v_5531;
wire v_5532;
wire v_5533;
wire v_5534;
wire v_5535;
wire v_5536;
wire v_5537;
wire v_5538;
wire v_5539;
wire v_5540;
wire v_5541;
wire v_5542;
wire v_5543;
wire v_5544;
wire v_5545;
wire v_5546;
wire v_5547;
wire v_5548;
wire v_5549;
wire v_5550;
wire v_5551;
wire v_5552;
wire v_5553;
wire v_5554;
wire v_5555;
wire v_5556;
wire v_5557;
wire v_5558;
wire v_5559;
wire v_5560;
wire v_5561;
wire v_5562;
wire v_5563;
wire v_5564;
wire v_5565;
wire v_5566;
wire v_5567;
wire v_5568;
wire v_5569;
wire v_5570;
wire v_5571;
wire v_5572;
wire v_5573;
wire v_5574;
wire v_5575;
wire v_5576;
wire v_5577;
wire v_5578;
wire v_5579;
wire v_5580;
wire v_5581;
wire v_5582;
wire v_5583;
wire v_5584;
wire v_5585;
wire v_5586;
wire v_5587;
wire v_5588;
wire v_5589;
wire v_5590;
wire v_5591;
wire v_5592;
wire v_5593;
wire v_5594;
wire v_5595;
wire v_5596;
wire v_5597;
wire v_5598;
wire v_5599;
wire v_5600;
wire v_5601;
wire v_5602;
wire v_5603;
wire v_5604;
wire v_5605;
wire v_5606;
wire v_5607;
wire v_5608;
wire v_5609;
wire v_5610;
wire v_5611;
wire v_5612;
wire v_5613;
wire v_5614;
wire v_5615;
wire v_5616;
wire v_5617;
wire v_5618;
wire v_5619;
wire v_5620;
wire v_5621;
wire v_5622;
wire v_5623;
wire v_5624;
wire v_5625;
wire v_5626;
wire v_5627;
wire v_5628;
wire v_5629;
wire v_5630;
wire v_5631;
wire v_5632;
wire v_5633;
wire v_5634;
wire v_5635;
wire v_5636;
wire v_5637;
wire v_5638;
wire v_5639;
wire v_5640;
wire v_5641;
wire v_5642;
wire v_5643;
wire v_5644;
wire v_5645;
wire v_5646;
wire v_5647;
wire v_5648;
wire v_5649;
wire v_5650;
wire v_5651;
wire v_5652;
wire v_5653;
wire v_5654;
wire v_5655;
wire v_5656;
wire v_5657;
wire v_5658;
wire v_5659;
wire v_5660;
wire v_5661;
wire v_5662;
wire v_5663;
wire v_5664;
wire v_5665;
wire v_5666;
wire v_5667;
wire v_5668;
wire v_5669;
wire v_5670;
wire v_5671;
wire v_5672;
wire v_5673;
wire v_5674;
wire v_5675;
wire v_5676;
wire v_5677;
wire v_5678;
wire v_5679;
wire v_5680;
wire v_5681;
wire v_5682;
wire v_5683;
wire v_5684;
wire v_5685;
wire v_5686;
wire v_5687;
wire v_5688;
wire v_5689;
wire v_5690;
wire v_5691;
wire v_5692;
wire v_5693;
wire v_5694;
wire v_5695;
wire v_5696;
wire v_5697;
wire v_5698;
wire v_5699;
wire v_5700;
wire v_5701;
wire v_5702;
wire v_5703;
wire v_5704;
wire v_5705;
wire v_5706;
wire v_5707;
wire v_5708;
wire v_5709;
wire v_5710;
wire v_5711;
wire v_5712;
wire v_5713;
wire v_5714;
wire v_5715;
wire v_5716;
wire v_5717;
wire v_5718;
wire v_5719;
wire v_5720;
wire v_5721;
wire v_5722;
wire v_5723;
wire v_5724;
wire v_5725;
wire v_5726;
wire v_5727;
wire v_5728;
wire v_5729;
wire v_5730;
wire v_5731;
wire v_5732;
wire v_5733;
wire v_5734;
wire v_5735;
wire v_5736;
wire v_5737;
wire v_5738;
wire v_5739;
wire v_5740;
wire v_5741;
wire v_5742;
wire v_5743;
wire v_5744;
wire v_5745;
wire v_5746;
wire v_5747;
wire v_5748;
wire v_5749;
wire v_5750;
wire v_5751;
wire v_5752;
wire v_5753;
wire v_5754;
wire v_5755;
wire v_5756;
wire v_5757;
wire v_5758;
wire v_5759;
wire v_5760;
wire v_5761;
wire v_5762;
wire v_5763;
wire v_5764;
wire v_5765;
wire v_5766;
wire v_5767;
wire v_5768;
wire v_5769;
wire v_5770;
wire v_5771;
wire v_5772;
wire v_5773;
wire v_5774;
wire v_5775;
wire v_5776;
wire v_5777;
wire v_5778;
wire v_5779;
wire v_5780;
wire v_5781;
wire v_5782;
wire v_5783;
wire v_5784;
wire v_5785;
wire v_5786;
wire v_5787;
wire v_5788;
wire v_5789;
wire v_5790;
wire v_5791;
wire v_5792;
wire v_5793;
wire v_5794;
wire v_5795;
wire v_5796;
wire v_5797;
wire v_5798;
wire v_5799;
wire v_5800;
wire v_5801;
wire v_5802;
wire v_5803;
wire v_5804;
wire v_5805;
wire v_5806;
wire v_5807;
wire v_5808;
wire v_5809;
wire v_5810;
wire v_5811;
wire v_5812;
wire v_5813;
wire v_5814;
wire v_5815;
wire v_5816;
wire v_5817;
wire v_5818;
wire v_5819;
wire v_5820;
wire v_5821;
wire v_5822;
wire v_5823;
wire v_5824;
wire v_5825;
wire v_5826;
wire v_5827;
wire v_5828;
wire v_5829;
wire v_5830;
wire v_5832;
wire v_5833;
wire v_5834;
wire v_5835;
wire v_5837;
wire v_5838;
wire v_5839;
wire v_5840;
wire v_5841;
wire v_5842;
wire v_5843;
wire v_5844;
wire v_5845;
wire v_5846;
wire v_5847;
wire v_5848;
wire v_5849;
wire v_5850;
wire v_5851;
wire v_5852;
wire v_5853;
wire v_5854;
wire v_5855;
wire v_5856;
wire v_5857;
wire v_5858;
wire v_5859;
wire v_5860;
wire v_5861;
wire v_5862;
wire v_5863;
wire v_5864;
wire v_5865;
wire v_5866;
wire v_5867;
wire v_5868;
wire v_5869;
wire v_5870;
wire v_5871;
wire v_5872;
wire v_5873;
wire v_5874;
wire v_5875;
wire v_5876;
wire v_5877;
wire v_5878;
wire v_5879;
wire v_5880;
wire v_5881;
wire v_5882;
wire v_5883;
wire v_5884;
wire v_5885;
wire v_5886;
wire v_5887;
wire v_5888;
wire v_5889;
wire v_5890;
wire v_5891;
wire v_5892;
wire v_5893;
wire v_5894;
wire v_5895;
wire v_5896;
wire v_5897;
wire v_5898;
wire v_5899;
wire v_5900;
wire v_5901;
wire v_5902;
wire v_5903;
wire v_5904;
wire v_5905;
wire v_5906;
wire v_5907;
wire v_5908;
wire v_5909;
wire v_5910;
wire v_5911;
wire v_5912;
wire v_5913;
wire v_5914;
wire v_5915;
wire v_5916;
wire v_5917;
wire v_5918;
wire v_5919;
wire v_5920;
wire v_5921;
wire v_5922;
wire v_5923;
wire v_5924;
wire v_5925;
wire v_5926;
wire v_5927;
wire v_5928;
wire v_5929;
wire v_5930;
wire v_5932;
wire v_5933;
wire v_5934;
wire v_5935;
wire v_5936;
wire v_5937;
wire v_5938;
wire v_5939;
wire v_5940;
wire v_5941;
wire v_5942;
wire v_5943;
wire v_5944;
wire v_5945;
wire v_5946;
wire v_5947;
wire v_5948;
wire v_5949;
wire v_5950;
wire v_5951;
wire v_5952;
wire v_5953;
wire v_5954;
wire v_5955;
wire v_5956;
wire v_5957;
wire v_5958;
wire v_5959;
wire v_5960;
wire v_5961;
wire v_5962;
wire v_5963;
wire v_5964;
wire v_5965;
wire v_5966;
wire v_5967;
wire v_5968;
wire v_5969;
wire v_5970;
wire v_5971;
wire v_5972;
wire v_5973;
wire v_5974;
wire v_5975;
wire v_5976;
wire v_5977;
wire v_5978;
wire v_5979;
wire v_5980;
wire v_5981;
wire v_5982;
wire v_5983;
wire v_5984;
wire v_5985;
wire v_5986;
wire v_5987;
wire v_5988;
wire v_5989;
wire v_5990;
wire v_5991;
wire v_5992;
wire v_5993;
wire v_5994;
wire v_5995;
wire v_5996;
wire v_5997;
wire v_5998;
wire v_5999;
wire v_6000;
wire v_6001;
wire v_6002;
wire v_6003;
wire v_6004;
wire v_6005;
wire v_6006;
wire v_6007;
wire v_6008;
wire v_6009;
wire v_6010;
wire v_6011;
wire v_6012;
wire v_6013;
wire v_6014;
wire v_6015;
wire v_6016;
wire v_6017;
wire v_6018;
wire v_6019;
wire v_6020;
wire v_6021;
wire v_6022;
wire v_6023;
wire v_6024;
wire v_6025;
wire v_6026;
wire v_6027;
wire v_6028;
wire v_6029;
wire v_6030;
wire v_6031;
wire v_6032;
wire v_6033;
wire v_6034;
wire v_6035;
wire v_6036;
wire v_6037;
wire v_6038;
wire v_6039;
wire v_6040;
wire v_6041;
wire v_6042;
wire v_6043;
wire v_6044;
wire v_6045;
wire v_6046;
wire v_6047;
wire v_6048;
wire v_6049;
wire v_6050;
wire v_6051;
wire v_6052;
wire v_6053;
wire v_6054;
wire v_6055;
wire v_6056;
wire v_6057;
wire v_6058;
wire v_6059;
wire v_6060;
wire v_6061;
wire v_6062;
wire v_6063;
wire v_6064;
wire v_6065;
wire v_6066;
wire v_6067;
wire v_6068;
wire v_6069;
wire v_6070;
wire v_6071;
wire v_6072;
wire v_6073;
wire v_6074;
wire v_6075;
wire v_6076;
wire v_6077;
wire v_6078;
wire v_6079;
wire v_6080;
wire v_6081;
wire v_6082;
wire v_6083;
wire v_6084;
wire v_6085;
wire v_6086;
wire v_6087;
wire v_6088;
wire v_6089;
wire v_6090;
wire v_6091;
wire v_6092;
wire v_6093;
wire v_6094;
wire v_6095;
wire v_6096;
wire v_6097;
wire v_6098;
wire v_6099;
wire v_6100;
wire v_6101;
wire v_6102;
wire v_6103;
wire v_6104;
wire v_6105;
wire v_6106;
wire v_6107;
wire v_6108;
wire v_6109;
wire v_6110;
wire v_6111;
wire v_6112;
wire v_6113;
wire v_6114;
wire v_6115;
wire v_6116;
wire v_6117;
wire v_6118;
wire v_6119;
wire v_6120;
wire v_6121;
wire v_6122;
wire v_6123;
wire v_6124;
wire v_6125;
wire v_6126;
wire v_6127;
wire v_6128;
wire v_6129;
wire v_6130;
wire v_6131;
wire v_6132;
wire v_6133;
wire v_6134;
wire v_6135;
wire v_6136;
wire v_6137;
wire v_6138;
wire v_6139;
wire v_6140;
wire v_6141;
wire v_6142;
wire v_6143;
wire v_6144;
wire v_6145;
wire v_6146;
wire v_6147;
wire v_6148;
wire v_6149;
wire v_6150;
wire v_6151;
wire v_6152;
wire v_6153;
wire v_6154;
wire v_6155;
wire v_6156;
wire v_6157;
wire v_6158;
wire v_6159;
wire v_6160;
wire v_6161;
wire v_6162;
wire v_6163;
wire v_6164;
wire v_6165;
wire v_6166;
wire v_6167;
wire v_6168;
wire v_6169;
wire v_6170;
wire v_6171;
wire v_6172;
wire v_6173;
wire v_6174;
wire v_6175;
wire v_6176;
wire v_6177;
wire v_6178;
wire v_6179;
wire v_6180;
wire v_6181;
wire v_6182;
wire v_6183;
wire v_6184;
wire v_6185;
wire v_6186;
wire v_6187;
wire v_6188;
wire v_6189;
wire v_6190;
wire v_6191;
wire v_6192;
wire v_6193;
wire v_6194;
wire v_6195;
wire v_6196;
wire v_6197;
wire v_6198;
wire v_6199;
wire v_6200;
wire v_6201;
wire v_6202;
wire v_6203;
wire v_6204;
wire v_6205;
wire v_6206;
wire v_6207;
wire v_6208;
wire v_6209;
wire v_6210;
wire v_6211;
wire v_6212;
wire v_6213;
wire v_6214;
wire v_6215;
wire v_6216;
wire v_6217;
wire v_6218;
wire v_6219;
wire v_6220;
wire v_6221;
wire v_6222;
wire v_6223;
wire v_6224;
wire v_6225;
wire v_6226;
wire v_6227;
wire v_6228;
wire v_6229;
wire v_6230;
wire v_6231;
wire v_6232;
wire v_6233;
wire v_6234;
wire v_6235;
wire v_6236;
wire v_6237;
wire v_6238;
wire v_6239;
wire v_6240;
wire v_6241;
wire v_6242;
wire v_6243;
wire v_6244;
wire v_6245;
wire v_6246;
wire v_6247;
wire v_6248;
wire v_6249;
wire v_6250;
wire v_6251;
wire v_6252;
wire v_6253;
wire v_6254;
wire v_6255;
wire v_6256;
wire v_6257;
wire v_6258;
wire v_6259;
wire v_6260;
wire v_6261;
wire v_6262;
wire v_6263;
wire v_6264;
wire v_6265;
wire v_6266;
wire v_6267;
wire v_6268;
wire v_6269;
wire v_6270;
wire v_6271;
wire v_6272;
wire v_6273;
wire v_6274;
wire v_6275;
wire v_6276;
wire v_6277;
wire v_6278;
wire v_6279;
wire v_6280;
wire v_6281;
wire v_6282;
wire v_6283;
wire v_6284;
wire v_6285;
wire v_6286;
wire v_6287;
wire v_6288;
wire v_6289;
wire v_6290;
wire v_6291;
wire v_6292;
wire v_6293;
wire v_6294;
wire v_6295;
wire v_6296;
wire v_6297;
wire v_6298;
wire v_6299;
wire v_6300;
wire v_6301;
wire v_6302;
wire v_6303;
wire v_6304;
wire v_6305;
wire v_6306;
wire v_6307;
wire v_6308;
wire v_6309;
wire v_6310;
wire v_6311;
wire v_6312;
wire v_6313;
wire v_6314;
wire v_6315;
wire v_6316;
wire v_6317;
wire v_6318;
wire v_6319;
wire v_6320;
wire v_6321;
wire v_6322;
wire v_6323;
wire v_6324;
wire v_6325;
wire v_6326;
wire v_6327;
wire v_6328;
wire v_6329;
wire v_6330;
wire v_6331;
wire v_6333;
wire v_6334;
wire v_6335;
wire v_6336;
wire v_6337;
wire v_6338;
wire v_6339;
wire v_6340;
wire v_6341;
wire v_6342;
wire v_6343;
wire v_6344;
wire v_6345;
wire v_6346;
wire v_6347;
wire v_6348;
wire v_6349;
wire v_6350;
wire v_6351;
wire v_6352;
wire v_6353;
wire v_6354;
wire v_6355;
wire v_6356;
wire v_6357;
wire v_6358;
wire v_6359;
wire v_6360;
wire v_6361;
wire v_6362;
wire v_6363;
wire v_6364;
wire v_6365;
wire v_6366;
wire v_6367;
wire v_6368;
wire v_6369;
wire v_6370;
wire v_6371;
wire v_6372;
wire v_6373;
wire v_6374;
wire v_6375;
wire v_6376;
wire v_6377;
wire v_6378;
wire v_6379;
wire v_6380;
wire v_6381;
wire v_6382;
wire v_6383;
wire v_6384;
wire v_6385;
wire v_6386;
wire v_6387;
wire v_6388;
wire v_6389;
wire v_6390;
wire v_6391;
wire v_6392;
wire v_6393;
wire v_6394;
wire v_6395;
wire v_6396;
wire v_6397;
wire v_6398;
wire v_6399;
wire v_6400;
wire v_6401;
wire v_6402;
wire v_6403;
wire v_6404;
wire v_6405;
wire v_6406;
wire v_6407;
wire v_6408;
wire v_6409;
wire v_6410;
wire v_6411;
wire v_6412;
wire v_6413;
wire v_6414;
wire v_6415;
wire v_6416;
wire v_6417;
wire v_6418;
wire v_6419;
wire v_6420;
wire v_6421;
wire v_6422;
wire v_6423;
wire v_6424;
wire v_6425;
wire v_6426;
wire v_6427;
wire v_6428;
wire v_6429;
wire v_6430;
wire v_6431;
wire v_6432;
wire v_6433;
wire v_6434;
wire v_6435;
wire v_6436;
wire v_6437;
wire v_6438;
wire v_6439;
wire v_6440;
wire v_6441;
wire v_6442;
wire v_6443;
wire v_6444;
wire v_6445;
wire v_6446;
wire v_6447;
wire v_6448;
wire v_6449;
wire v_6450;
wire v_6451;
wire v_6452;
wire v_6453;
wire v_6454;
wire v_6455;
wire v_6456;
wire v_6458;
wire v_6459;
wire v_6460;
wire v_6461;
wire v_6462;
wire v_6463;
wire v_6464;
wire v_6465;
wire v_6466;
wire v_6467;
wire v_6468;
wire v_6469;
wire v_6470;
wire v_6471;
wire v_6472;
wire v_6473;
wire v_6474;
wire v_6475;
wire v_6476;
wire v_6478;
wire v_6479;
wire v_6480;
wire v_6481;
wire v_6482;
wire v_6483;
wire v_6484;
wire v_6485;
wire v_6486;
wire v_6487;
wire v_6488;
wire v_6489;
wire v_6490;
wire v_6491;
wire v_6492;
wire v_6493;
wire v_6494;
wire v_6495;
wire v_6496;
wire v_6497;
wire v_6498;
wire v_6499;
wire v_6500;
wire v_6501;
wire v_6502;
wire v_6503;
wire v_6504;
wire v_6505;
wire v_6506;
wire v_6507;
wire v_6508;
wire v_6509;
wire v_6510;
wire v_6511;
wire v_6512;
wire v_6513;
wire v_6514;
wire v_6515;
wire v_6516;
wire v_6517;
wire v_6518;
wire v_6519;
wire v_6520;
wire v_6521;
wire v_6522;
wire v_6523;
wire v_6524;
wire v_6525;
wire v_6526;
wire v_6527;
wire v_6529;
wire v_6530;
wire v_6531;
wire v_6532;
wire v_6533;
wire v_6534;
wire v_6535;
wire v_6536;
wire v_6537;
wire v_6538;
wire v_6539;
wire v_6540;
wire v_6541;
wire v_6542;
wire v_6543;
wire v_6544;
wire v_6545;
wire v_6547;
wire v_6548;
wire v_6549;
wire v_6550;
wire v_6551;
wire v_6552;
wire v_6553;
wire v_6554;
wire v_6555;
wire v_6556;
wire v_6557;
wire v_6558;
wire v_6559;
wire v_6560;
wire v_6561;
wire v_6562;
wire v_6563;
wire v_6564;
wire v_6565;
wire v_6566;
wire v_6567;
wire v_6568;
wire v_6569;
wire v_6570;
wire v_6571;
wire v_6572;
wire v_6573;
wire v_6574;
wire v_6575;
wire v_6576;
wire v_6577;
wire v_6578;
wire v_6579;
wire v_6580;
wire v_6581;
wire v_6582;
wire v_6583;
wire v_6584;
wire v_6585;
wire v_6586;
wire v_6587;
wire v_6588;
wire v_6589;
wire v_6590;
wire v_6591;
wire v_6592;
wire v_6593;
wire v_6594;
wire v_6595;
wire v_6596;
wire v_6597;
wire v_6598;
wire v_6599;
wire v_6600;
wire v_6601;
wire v_6602;
wire v_6603;
wire v_6604;
wire v_6605;
wire v_6606;
wire v_6607;
wire v_6608;
wire v_6609;
wire v_6610;
wire v_6611;
wire v_6612;
wire v_6613;
wire v_6614;
wire v_6615;
wire v_6616;
wire v_6617;
wire v_6618;
wire v_6619;
wire v_6620;
wire v_6621;
wire v_6622;
wire v_6623;
wire v_6624;
wire v_6625;
wire v_6626;
wire v_6627;
wire v_6628;
wire v_6629;
wire v_6630;
wire v_6631;
wire v_6632;
wire v_6633;
wire v_6634;
wire v_6635;
wire v_6636;
wire v_6637;
wire v_6638;
wire v_6639;
wire v_6640;
wire v_6641;
wire v_6642;
wire v_6643;
wire v_6644;
wire v_6645;
wire v_6646;
wire v_6647;
wire v_6648;
wire v_6649;
wire v_6650;
wire v_6651;
wire v_6652;
wire v_6653;
wire v_6654;
wire v_6655;
wire v_6656;
wire v_6657;
wire v_6658;
wire v_6659;
wire v_6660;
wire v_6661;
wire v_6662;
wire v_6663;
wire v_6664;
wire v_6665;
wire v_6666;
wire v_6667;
wire v_6668;
wire v_6669;
wire v_6670;
wire v_6671;
wire v_6672;
wire v_6673;
wire v_6674;
wire v_6675;
wire v_6676;
wire v_6677;
wire v_6678;
wire v_6679;
wire v_6680;
wire v_6681;
wire v_6682;
wire v_6683;
wire v_6684;
wire v_6685;
wire v_6686;
wire v_6687;
wire v_6688;
wire v_6689;
wire v_6690;
wire v_6691;
wire v_6692;
wire v_6693;
wire v_6694;
wire v_6695;
wire v_6696;
wire v_6697;
wire v_6698;
wire v_6699;
wire v_6700;
wire v_6701;
wire v_6702;
wire v_6703;
wire v_6704;
wire v_6705;
wire v_6706;
wire v_6707;
wire v_6708;
wire v_6709;
wire v_6710;
wire v_6711;
wire v_6712;
wire v_6713;
wire v_6714;
wire v_6715;
wire v_6716;
wire v_6717;
wire v_6718;
wire v_6719;
wire v_6720;
wire v_6721;
wire v_6722;
wire v_6723;
wire v_6724;
wire v_6725;
wire v_6726;
wire v_6727;
wire v_6728;
wire v_6729;
wire v_6730;
wire v_6731;
wire v_6732;
wire v_6733;
wire v_6734;
wire v_6735;
wire v_6736;
wire v_6737;
wire v_6738;
wire v_6739;
wire v_6740;
wire v_6741;
wire v_6742;
wire v_6743;
wire v_6744;
wire v_6745;
wire v_6746;
wire v_6747;
wire v_6748;
wire v_6749;
wire v_6750;
wire v_6751;
wire v_6752;
wire v_6753;
wire v_6754;
wire v_6755;
wire v_6756;
wire v_6757;
wire v_6758;
wire v_6759;
wire v_6760;
wire v_6761;
wire v_6762;
wire v_6763;
wire v_6764;
wire v_6765;
wire v_6766;
wire v_6767;
wire v_6768;
wire v_6769;
wire v_6770;
wire v_6771;
wire v_6772;
wire v_6773;
wire v_6774;
wire v_6775;
wire v_6776;
wire v_6777;
wire v_6778;
wire v_6779;
wire v_6780;
wire v_6781;
wire v_6782;
wire v_6783;
wire v_6784;
wire v_6785;
wire v_6786;
wire v_6787;
wire v_6788;
wire v_6789;
wire v_6790;
wire v_6791;
wire v_6792;
wire v_6793;
wire v_6794;
wire v_6795;
wire v_6796;
wire v_6797;
wire v_6798;
wire v_6799;
wire v_6800;
wire v_6801;
wire v_6802;
wire v_6803;
wire v_6804;
wire v_6805;
wire v_6806;
wire v_6807;
wire v_6808;
wire v_6809;
wire v_6810;
wire v_6811;
wire v_6812;
wire v_6813;
wire v_6814;
wire v_6815;
wire v_6816;
wire v_6817;
wire v_6818;
wire v_6819;
wire v_6820;
wire v_6821;
wire v_6822;
wire v_6823;
wire v_6824;
wire v_6825;
wire v_6826;
wire v_6827;
wire v_6828;
wire v_6829;
wire v_6830;
wire v_6831;
wire v_6832;
wire v_6833;
wire v_6834;
wire v_6835;
wire v_6836;
wire v_6837;
wire v_6838;
wire v_6839;
wire v_6840;
wire v_6841;
wire v_6842;
wire v_6843;
wire v_6844;
wire v_6845;
wire v_6846;
wire v_6847;
wire v_6848;
wire v_6849;
wire v_6850;
wire v_6851;
wire v_6852;
wire v_6853;
wire v_6854;
wire v_6855;
wire v_6856;
wire v_6857;
wire v_6858;
wire v_6859;
wire v_6860;
wire v_6861;
wire v_6862;
wire v_6863;
wire v_6864;
wire v_6865;
wire v_6866;
wire v_6867;
wire v_6872;
wire v_6875;
wire v_6876;
wire v_6877;
wire v_6878;
wire v_6879;
wire v_6880;
wire v_6881;
wire v_6882;
wire v_6883;
wire v_6884;
wire v_6885;
wire v_6886;
wire v_6887;
wire v_6888;
wire v_6889;
wire v_6890;
wire v_6891;
wire v_6892;
wire v_6893;
wire v_6894;
wire v_6895;
wire v_6896;
wire v_6897;
wire v_6898;
wire v_6899;
wire v_6900;
wire v_6901;
wire v_6902;
wire v_6903;
wire v_6904;
wire v_6905;
wire v_6906;
wire v_6907;
wire v_6908;
wire v_6909;
wire v_6910;
wire v_6911;
wire v_6912;
wire v_6913;
wire v_6914;
wire v_6915;
wire v_6916;
wire v_6917;
wire v_6918;
wire v_6919;
wire v_6920;
wire v_6921;
wire v_6922;
wire v_6923;
wire v_6924;
wire v_6925;
wire v_6926;
wire v_6927;
wire v_6928;
wire v_6929;
wire v_6930;
wire v_6931;
wire v_6932;
wire v_6933;
wire v_6934;
wire v_6935;
wire v_6936;
wire v_6937;
wire v_6938;
wire v_6939;
wire v_6940;
wire v_6941;
wire v_6942;
wire v_6943;
wire v_6944;
wire v_6945;
wire v_6946;
wire v_6947;
wire v_6948;
wire v_6949;
wire v_6950;
wire v_6951;
wire v_6952;
wire v_6953;
wire v_6954;
wire v_6955;
wire v_6956;
wire v_6957;
wire v_6958;
wire v_6959;
wire v_6960;
wire v_6961;
wire v_6962;
wire v_6963;
wire v_6964;
wire v_6965;
wire v_6966;
wire v_6967;
wire v_6968;
wire v_6969;
wire v_6970;
wire v_6971;
wire v_6972;
wire v_6973;
wire v_6974;
wire v_6975;
wire v_6976;
wire v_6977;
wire v_6978;
wire v_6979;
wire v_6980;
wire v_6981;
wire v_6982;
wire v_6983;
wire v_6984;
wire v_6985;
wire v_6986;
wire v_6987;
wire v_6988;
wire v_6989;
wire v_6990;
wire v_6991;
wire v_6992;
wire v_6993;
wire v_6994;
wire v_6995;
wire v_6996;
wire v_6997;
wire v_6998;
wire v_6999;
wire v_7000;
wire v_7001;
wire v_7002;
wire v_7003;
wire v_7004;
wire v_7005;
wire v_7006;
wire v_7007;
wire v_7008;
wire v_7009;
wire v_7010;
wire v_7011;
wire v_7012;
wire v_7013;
wire v_7014;
wire v_7015;
wire v_7016;
wire v_7017;
wire v_7018;
wire v_7019;
wire v_7020;
wire v_7021;
wire v_7022;
wire v_7023;
wire v_7024;
wire v_7025;
wire v_7026;
wire v_7027;
wire v_7028;
wire v_7029;
wire v_7030;
wire v_7031;
wire v_7032;
wire v_7033;
wire v_7034;
wire v_7035;
wire v_7036;
wire v_7037;
wire v_7038;
wire v_7039;
wire v_7040;
wire v_7041;
wire v_7042;
wire v_7043;
wire v_7044;
wire v_7045;
wire v_7046;
wire v_7047;
wire v_7048;
wire v_7049;
wire v_7050;
wire v_7051;
wire v_7052;
wire v_7053;
wire v_7054;
wire v_7055;
wire v_7056;
wire v_7057;
wire v_7058;
wire v_7059;
wire v_7060;
wire v_7061;
wire v_7062;
wire v_7063;
wire v_7064;
wire v_7065;
wire v_7066;
wire v_7067;
wire v_7068;
wire v_7069;
wire v_7070;
wire v_7071;
wire v_7072;
wire v_7073;
wire v_7074;
wire v_7075;
wire v_7076;
wire v_7077;
wire v_7078;
wire v_7081;
wire v_7082;
wire v_7083;
wire v_7084;
wire v_7086;
wire v_7088;
wire v_7089;
wire v_7090;
wire v_7092;
wire v_7094;
wire v_7097;
wire v_7099;
wire v_7101;
wire v_7104;
wire v_7106;
wire v_7108;
wire v_7110;
wire v_7112;
wire v_7114;
wire v_7116;
wire v_7118;
wire v_7119;
wire v_7122;
wire v_7123;
wire v_7124;
wire v_7125;
wire v_7126;
wire v_7127;
wire v_7129;
wire v_7131;
wire v_7132;
wire v_7133;
wire v_7135;
wire v_7136;
wire v_7137;
wire v_7139;
wire v_7141;
wire v_7142;
wire v_7143;
wire v_7144;
wire v_7148;
wire v_7150;
wire v_7151;
wire v_7153;
wire v_7155;
wire v_7156;
wire v_7157;
wire v_7160;
wire v_7162;
wire v_7165;
wire v_7166;
wire v_7167;
wire v_7168;
wire v_7170;
wire v_7171;
wire v_7172;
wire v_7173;
wire v_7176;
wire v_7179;
wire v_7180;
wire v_7181;
wire v_7183;
wire v_7185;
wire v_7186;
wire v_7187;
wire v_7189;
wire v_7191;
wire v_7193;
wire v_7194;
wire v_7195;
wire v_7196;
wire v_7197;
wire v_7198;
wire v_7201;
wire v_7203;
wire v_7205;
wire v_7207;
wire v_7208;
wire v_7209;
wire v_7210;
wire v_7213;
wire v_7215;
wire v_7217;
wire v_7219;
wire v_7221;
wire v_7222;
wire v_7224;
wire v_7227;
wire v_7229;
wire v_7231;
wire v_7233;
wire v_7234;
wire v_7235;
wire v_7237;
wire v_7240;
wire v_7242;
wire v_7244;
wire v_7246;
wire v_7248;
wire v_7249;
wire v_7250;
wire v_7252;
wire v_7253;
wire v_7254;
wire v_7256;
wire v_7259;
wire v_7261;
wire v_7263;
wire v_7265;
wire v_7267;
wire v_7268;
wire v_7269;
wire v_7270;
wire v_7271;
wire v_7273;
wire v_7274;
wire v_7275;
wire v_7278;
wire v_7280;
wire v_7282;
wire v_7284;
wire v_7286;
wire v_7287;
wire v_7289;
wire v_7292;
wire v_7294;
wire v_7296;
wire v_7298;
wire v_7299;
wire v_7300;
wire v_7302;
wire v_7305;
wire v_7307;
wire v_7309;
wire v_7311;
wire v_7313;
wire v_7314;
wire v_7315;
wire v_7317;
wire v_7318;
wire v_7319;
wire v_7321;
wire v_7324;
wire v_7326;
wire v_7328;
wire v_7330;
wire v_7332;
wire v_7333;
wire v_7334;
wire v_7335;
wire v_7336;
wire v_7338;
wire v_7339;
wire v_7340;
wire v_7342;
wire v_7344;
wire v_7345;
wire v_7346;
wire v_7348;
wire v_7349;
wire v_7350;
wire v_7351;
wire v_7353;
wire v_7354;
wire v_7356;
wire v_7358;
wire v_7361;
wire v_7363;
wire v_7365;
wire v_7368;
wire v_7370;
wire v_7372;
wire v_7374;
wire v_7376;
wire v_7378;
wire v_7380;
wire v_7382;
wire v_7383;
wire v_7386;
wire v_7387;
wire v_7388;
wire v_7389;
wire v_7390;
wire v_7391;
wire v_7393;
wire v_7395;
wire v_7396;
wire v_7397;
wire v_7399;
wire v_7400;
wire v_7401;
wire v_7402;
wire v_7404;
wire v_7405;
wire v_7406;
wire v_7407;
wire v_7410;
wire v_7411;
wire v_7412;
wire v_7414;
wire v_7416;
wire v_7418;
wire v_7419;
wire v_7420;
wire v_7422;
wire v_7423;
wire v_7424;
wire v_7426;
wire v_7428;
wire v_7430;
wire v_7432;
wire v_7433;
wire v_7434;
wire v_7436;
wire v_7438;
wire v_7441;
wire v_7442;
wire v_7443;
wire v_7445;
wire v_7446;
wire v_7447;
wire v_7448;
wire v_7451;
wire v_7453;
wire v_7454;
wire v_7456;
wire v_7458;
wire v_7459;
wire v_7461;
wire v_7462;
wire v_7463;
wire v_7464;
wire v_7465;
wire v_7468;
wire v_7469;
wire v_7470;
wire v_7472;
wire v_7474;
wire v_7476;
wire v_7477;
wire v_7478;
wire v_7480;
wire v_7481;
wire v_7482;
wire v_7484;
wire v_7486;
wire v_7488;
wire v_7490;
wire v_7491;
wire v_7492;
wire v_7494;
wire v_7496;
wire v_7499;
wire v_7500;
wire v_7501;
wire v_7503;
wire v_7504;
wire v_7505;
wire v_7506;
wire v_7508;
wire v_7510;
wire v_7512;
wire v_7514;
wire v_7516;
wire v_7517;
wire v_7518;
wire v_7519;
wire v_7520;
wire v_7521;
wire v_7522;
wire v_7523;
wire v_7524;
wire v_7525;
wire v_7526;
wire v_7527;
wire v_7528;
wire v_7530;
wire v_7531;
wire v_7533;
wire v_7534;
wire v_7537;
wire v_7539;
wire v_7542;
wire v_7543;
wire v_7544;
wire v_7545;
wire v_7547;
wire v_7549;
wire v_7552;
wire v_7554;
wire v_7555;
wire v_7557;
wire v_7559;
wire v_7560;
wire v_7562;
wire v_7563;
wire v_7564;
wire v_7565;
wire v_7567;
wire v_7568;
wire v_7569;
wire v_7570;
wire v_7574;
wire v_7575;
wire v_7576;
wire v_7578;
wire v_7580;
wire v_7582;
wire v_7583;
wire v_7584;
wire v_7586;
wire v_7587;
wire v_7588;
wire v_7591;
wire v_7594;
wire v_7596;
wire v_7598;
wire v_7600;
wire v_7602;
wire v_7603;
wire v_7606;
wire v_7607;
wire v_7609;
wire v_7610;
wire v_7611;
wire v_7614;
wire v_7615;
wire v_7616;
wire v_7618;
wire v_7620;
wire v_7622;
wire v_7623;
wire v_7624;
wire v_7627;
wire v_7628;
wire v_7629;
wire v_7631;
wire v_7633;
wire v_7635;
wire v_7636;
wire v_7637;
wire v_7639;
wire v_7640;
wire v_7643;
wire v_7644;
wire v_7645;
wire v_7647;
wire v_7649;
wire v_7651;
wire v_7652;
wire v_7653;
wire v_7655;
wire v_7656;
wire v_7657;
wire v_7659;
wire v_7660;
wire v_7661;
wire v_7662;
wire v_7663;
wire v_7668;
wire v_7669;
wire v_7670;
wire v_7672;
wire v_7673;
wire v_7674;
wire v_7676;
wire v_7678;
wire v_7679;
wire v_7680;
wire v_7682;
wire v_7684;
wire v_7685;
wire v_7686;
wire v_7687;
wire v_7691;
wire v_7692;
wire v_7693;
wire v_7695;
wire v_7696;
wire v_7697;
wire v_7699;
wire v_7701;
wire v_7702;
wire v_7703;
wire v_7705;
wire v_7707;
wire v_7708;
wire v_7709;
wire v_7710;
wire v_7714;
wire v_7715;
wire v_7716;
wire v_7718;
wire v_7719;
wire v_7720;
wire v_7722;
wire v_7724;
wire v_7725;
wire v_7726;
wire v_7728;
wire v_7730;
wire v_7731;
wire v_7732;
wire v_7733;
wire v_7737;
wire v_7739;
wire v_7740;
wire v_7741;
wire v_7742;
wire v_7743;
wire v_7744;
wire v_7749;
wire v_7750;
wire v_7751;
wire v_7753;
wire v_7754;
wire v_7755;
wire v_7757;
wire v_7759;
wire v_7760;
wire v_7761;
wire v_7763;
wire v_7765;
wire v_7766;
wire v_7767;
wire v_7768;
wire v_7772;
wire v_7773;
wire v_7774;
wire v_7776;
wire v_7777;
wire v_7778;
wire v_7780;
wire v_7782;
wire v_7783;
wire v_7784;
wire v_7786;
wire v_7788;
wire v_7789;
wire v_7790;
wire v_7791;
wire v_7795;
wire v_7796;
wire v_7797;
wire v_7799;
wire v_7800;
wire v_7801;
wire v_7803;
wire v_7805;
wire v_7806;
wire v_7807;
wire v_7809;
wire v_7811;
wire v_7812;
wire v_7813;
wire v_7814;
wire v_7818;
wire v_7820;
wire v_7821;
wire v_7822;
wire v_7823;
wire v_7824;
wire v_7825;
wire v_7830;
wire v_7831;
wire v_7832;
wire v_7834;
wire v_7835;
wire v_7836;
wire v_7838;
wire v_7840;
wire v_7841;
wire v_7842;
wire v_7844;
wire v_7846;
wire v_7847;
wire v_7848;
wire v_7849;
wire v_7853;
wire v_7854;
wire v_7855;
wire v_7857;
wire v_7858;
wire v_7859;
wire v_7861;
wire v_7863;
wire v_7864;
wire v_7865;
wire v_7867;
wire v_7869;
wire v_7870;
wire v_7871;
wire v_7872;
wire v_7876;
wire v_7877;
wire v_7878;
wire v_7880;
wire v_7881;
wire v_7882;
wire v_7884;
wire v_7886;
wire v_7887;
wire v_7888;
wire v_7890;
wire v_7892;
wire v_7893;
wire v_7894;
wire v_7895;
wire v_7899;
wire v_7901;
wire v_7902;
wire v_7903;
wire v_7904;
wire v_7905;
wire v_7906;
wire v_7911;
wire v_7912;
wire v_7913;
wire v_7915;
wire v_7916;
wire v_7917;
wire v_7919;
wire v_7921;
wire v_7922;
wire v_7923;
wire v_7925;
wire v_7927;
wire v_7928;
wire v_7929;
wire v_7930;
wire v_7934;
wire v_7935;
wire v_7936;
wire v_7938;
wire v_7939;
wire v_7940;
wire v_7942;
wire v_7944;
wire v_7945;
wire v_7946;
wire v_7948;
wire v_7950;
wire v_7951;
wire v_7952;
wire v_7953;
wire v_7957;
wire v_7958;
wire v_7959;
wire v_7961;
wire v_7962;
wire v_7963;
wire v_7965;
wire v_7967;
wire v_7968;
wire v_7969;
wire v_7971;
wire v_7973;
wire v_7974;
wire v_7975;
wire v_7976;
wire v_7980;
wire v_7982;
wire v_7983;
wire v_7984;
wire v_7985;
wire v_7986;
wire v_7987;
wire v_7992;
wire v_7993;
wire v_7994;
wire v_7996;
wire v_7997;
wire v_7998;
wire v_8000;
wire v_8002;
wire v_8003;
wire v_8004;
wire v_8006;
wire v_8008;
wire v_8009;
wire v_8010;
wire v_8011;
wire v_8015;
wire v_8016;
wire v_8017;
wire v_8019;
wire v_8020;
wire v_8021;
wire v_8023;
wire v_8025;
wire v_8026;
wire v_8027;
wire v_8029;
wire v_8031;
wire v_8032;
wire v_8033;
wire v_8034;
wire v_8038;
wire v_8039;
wire v_8040;
wire v_8042;
wire v_8043;
wire v_8044;
wire v_8046;
wire v_8048;
wire v_8049;
wire v_8050;
wire v_8052;
wire v_8054;
wire v_8055;
wire v_8056;
wire v_8057;
wire v_8061;
wire v_8063;
wire v_8064;
wire v_8065;
wire v_8066;
wire v_8067;
wire v_8068;
wire v_8073;
wire v_8074;
wire v_8075;
wire v_8077;
wire v_8078;
wire v_8079;
wire v_8081;
wire v_8083;
wire v_8084;
wire v_8085;
wire v_8087;
wire v_8089;
wire v_8090;
wire v_8091;
wire v_8092;
wire v_8096;
wire v_8097;
wire v_8098;
wire v_8100;
wire v_8101;
wire v_8102;
wire v_8104;
wire v_8106;
wire v_8107;
wire v_8108;
wire v_8110;
wire v_8112;
wire v_8113;
wire v_8114;
wire v_8115;
wire v_8119;
wire v_8120;
wire v_8121;
wire v_8123;
wire v_8124;
wire v_8125;
wire v_8127;
wire v_8129;
wire v_8130;
wire v_8131;
wire v_8133;
wire v_8135;
wire v_8136;
wire v_8137;
wire v_8138;
wire v_8142;
wire v_8144;
wire v_8145;
wire v_8146;
wire v_8147;
wire v_8148;
wire v_8149;
wire v_8154;
wire v_8155;
wire v_8156;
wire v_8158;
wire v_8159;
wire v_8160;
wire v_8162;
wire v_8164;
wire v_8165;
wire v_8166;
wire v_8168;
wire v_8170;
wire v_8171;
wire v_8172;
wire v_8173;
wire v_8177;
wire v_8178;
wire v_8179;
wire v_8181;
wire v_8182;
wire v_8183;
wire v_8185;
wire v_8187;
wire v_8188;
wire v_8189;
wire v_8191;
wire v_8193;
wire v_8194;
wire v_8195;
wire v_8196;
wire v_8200;
wire v_8201;
wire v_8202;
wire v_8204;
wire v_8205;
wire v_8206;
wire v_8208;
wire v_8210;
wire v_8211;
wire v_8212;
wire v_8214;
wire v_8216;
wire v_8217;
wire v_8218;
wire v_8219;
wire v_8223;
wire v_8225;
wire v_8226;
wire v_8227;
wire v_8228;
wire v_8229;
wire v_8230;
wire v_8234;
wire v_8235;
wire v_8236;
wire v_8238;
wire v_8239;
wire v_8240;
wire v_8241;
wire v_8242;
wire v_8243;
wire v_8244;
wire v_8245;
wire v_8246;
wire v_8247;
wire v_8248;
wire v_8249;
wire v_8250;
wire v_8251;
wire v_8252;
wire v_8253;
wire v_8254;
wire v_8255;
wire v_8256;
wire v_8257;
wire v_8258;
wire v_8259;
wire v_8260;
wire v_8261;
wire v_8262;
wire v_8263;
wire v_8264;
wire v_8265;
wire v_8266;
wire v_8267;
wire v_8268;
wire v_8269;
wire v_8270;
wire v_8271;
wire v_8272;
wire v_8273;
wire v_8274;
wire v_8275;
wire v_8276;
wire v_8277;
wire v_8278;
wire v_8279;
wire v_8280;
wire v_8281;
wire v_8282;
wire v_8283;
wire v_8284;
wire v_8285;
wire v_8286;
wire v_8287;
wire v_8288;
wire v_8289;
wire v_8290;
wire v_8291;
wire v_8292;
wire v_8293;
wire v_8294;
wire v_8295;
wire v_8296;
wire v_8297;
wire v_8298;
wire v_8299;
wire v_8300;
wire v_8301;
wire v_8302;
wire v_8303;
wire v_8304;
wire v_8305;
wire v_8306;
wire v_8307;
wire v_8308;
wire v_8309;
wire v_8310;
wire v_8311;
wire v_8312;
wire v_8313;
wire v_8314;
wire v_8315;
wire v_8316;
wire v_8317;
wire v_8318;
wire v_8319;
wire v_8320;
wire v_8321;
wire v_8322;
wire v_8323;
wire v_8324;
wire v_8325;
wire v_8326;
wire v_8327;
wire v_8328;
wire v_8329;
wire v_8330;
wire v_8331;
wire v_8332;
wire v_8333;
wire v_8334;
wire v_8335;
wire v_8336;
wire v_8337;
wire v_8338;
wire v_8339;
wire v_8340;
wire v_8341;
wire v_8342;
wire v_8343;
wire v_8344;
wire v_8345;
wire v_8346;
wire v_8347;
wire v_8348;
wire v_8349;
wire v_8350;
wire v_8351;
wire v_8352;
wire v_8353;
wire v_8354;
wire v_8355;
wire v_8356;
wire v_8357;
wire v_8360;
wire v_8361;
wire v_8362;
wire v_8363;
wire v_8364;
wire v_8365;
wire v_8366;
wire v_8367;
wire v_8368;
wire v_8369;
wire v_8370;
wire v_8371;
wire v_8372;
wire v_8373;
wire v_8374;
wire v_8375;
wire v_8376;
wire v_8377;
wire v_8378;
wire v_8379;
wire v_8380;
wire v_8381;
wire v_8382;
wire v_8383;
wire v_8384;
wire v_8385;
wire v_8386;
wire v_8387;
wire v_8388;
wire v_8389;
wire v_8390;
wire v_8391;
wire v_8392;
wire v_8393;
wire v_8394;
wire v_8395;
wire v_8396;
wire v_8397;
wire v_8398;
wire v_8399;
wire v_8400;
wire v_8401;
wire v_8402;
wire v_8403;
wire v_8404;
wire v_8405;
wire v_8406;
wire v_8407;
wire v_8408;
wire v_8409;
wire v_8410;
wire v_8411;
wire v_8412;
wire v_8413;
wire v_8414;
wire v_8415;
wire v_8416;
wire v_8417;
wire v_8418;
wire v_8419;
wire v_8420;
wire v_8421;
wire v_8422;
wire v_8423;
wire v_8424;
wire v_8425;
wire v_8426;
wire v_8427;
wire v_8428;
wire v_8429;
wire v_8430;
wire v_8431;
wire v_8432;
wire v_8433;
wire v_8434;
wire v_8435;
wire v_8436;
wire v_8437;
wire v_8438;
wire v_8439;
wire v_8440;
wire v_8441;
wire v_8442;
wire v_8443;
wire v_8444;
wire v_8445;
wire v_8446;
wire v_8447;
wire v_8448;
wire v_8449;
wire v_8450;
wire v_8451;
wire v_8452;
wire v_8453;
wire v_8454;
wire v_8455;
wire v_8456;
wire v_8457;
wire v_8458;
wire v_8459;
wire v_8460;
wire v_8461;
wire v_8462;
wire v_8463;
wire v_8464;
wire v_8465;
wire v_8466;
wire v_8467;
wire v_8468;
wire v_8469;
wire v_8470;
wire v_8471;
wire v_8472;
wire v_8473;
wire v_8474;
wire v_8475;
wire v_8476;
wire v_8477;
wire v_8478;
wire v_8479;
wire v_8480;
wire v_8481;
wire v_8482;
wire v_8483;
wire v_8484;
wire v_8485;
wire v_8486;
wire v_8487;
wire v_8488;
wire v_8489;
wire v_8490;
wire v_8491;
wire v_8492;
wire v_8493;
wire v_8494;
wire v_8495;
wire v_8496;
wire v_8497;
wire v_8498;
wire v_8499;
wire v_8500;
wire v_8501;
wire v_8502;
wire v_8503;
wire v_8504;
wire v_8505;
wire v_8506;
wire v_8507;
wire v_8508;
wire v_8509;
wire v_8510;
wire v_8511;
wire v_8512;
wire v_8513;
wire v_8514;
wire v_8515;
wire v_8516;
wire v_8517;
wire v_8518;
wire v_8519;
wire v_8520;
wire v_8521;
wire v_8522;
wire v_8523;
wire v_8524;
wire v_8525;
wire v_8526;
wire v_8527;
wire v_8528;
wire v_8529;
wire v_8530;
wire v_8531;
wire v_8532;
wire v_8533;
wire v_8534;
wire v_8535;
wire v_8536;
wire v_8537;
wire v_8538;
wire v_8539;
wire v_8540;
wire v_8541;
wire v_8542;
wire v_8543;
wire v_8544;
wire v_8545;
wire v_8546;
wire v_8547;
wire v_8548;
wire v_8549;
wire v_8550;
wire v_8551;
wire v_8552;
wire v_8553;
wire v_8554;
wire v_8555;
wire v_8556;
wire v_8557;
wire v_8558;
wire v_8559;
wire v_8560;
wire v_8561;
wire v_8562;
wire v_8563;
wire v_8564;
wire v_8565;
wire v_8566;
wire v_8567;
wire v_8568;
wire v_8569;
wire v_8570;
wire v_8571;
wire v_8572;
wire v_8573;
wire v_8574;
wire v_8575;
wire v_8576;
wire v_8577;
wire v_8578;
wire v_8579;
wire v_8580;
wire v_8581;
wire v_8582;
wire v_8583;
wire v_8584;
wire v_8585;
wire v_8586;
wire v_8587;
wire v_8588;
wire v_8589;
wire v_8590;
wire v_8591;
wire v_8592;
wire v_8593;
wire v_8594;
wire v_8595;
wire v_8596;
wire v_8597;
wire v_8598;
wire v_8599;
wire v_8600;
wire v_8601;
wire v_8602;
wire v_8603;
wire v_8604;
wire v_8605;
wire v_8606;
wire v_8607;
wire v_8608;
wire v_8609;
wire v_8610;
wire v_8611;
wire v_8612;
wire v_8613;
wire v_8614;
wire v_8615;
wire v_8616;
wire v_8617;
wire v_8618;
wire v_8619;
wire v_8620;
wire v_8621;
wire v_8622;
wire v_8623;
wire v_8624;
wire v_8625;
wire v_8626;
wire v_8627;
wire v_8628;
wire v_8629;
wire v_8630;
wire v_8631;
wire v_8632;
wire v_8633;
wire v_8634;
wire v_8635;
wire v_8636;
wire v_8637;
wire v_8638;
wire v_8639;
wire v_8640;
wire v_8641;
wire v_8642;
wire v_8643;
wire v_8644;
wire v_8645;
wire v_8646;
wire v_8647;
wire v_8648;
wire v_8649;
wire v_8650;
wire v_8651;
wire v_8652;
wire v_8653;
wire v_8654;
wire v_8655;
wire v_8656;
wire v_8657;
wire v_8658;
wire v_8659;
wire v_8660;
wire v_8661;
wire v_8662;
wire v_8663;
wire v_8664;
wire v_8665;
wire v_8666;
wire v_8667;
wire v_8668;
wire v_8669;
wire v_8670;
wire v_8671;
wire v_8672;
wire v_8673;
wire v_8674;
wire v_8675;
wire v_8676;
wire v_8677;
wire v_8678;
wire v_8679;
wire v_8680;
wire v_8681;
wire v_8682;
wire v_8683;
wire v_8684;
wire v_8685;
wire v_8686;
wire v_8687;
wire v_8688;
wire v_8689;
wire v_8690;
wire v_8691;
wire v_8692;
wire v_8693;
wire v_8694;
wire v_8695;
wire v_8696;
wire v_8697;
wire v_8698;
wire v_8699;
wire v_8700;
wire v_8701;
wire v_8702;
wire v_8703;
wire v_8704;
wire v_8705;
wire v_8706;
wire v_8707;
wire v_8708;
wire v_8709;
wire v_8710;
wire v_8711;
wire v_8712;
wire v_8713;
wire v_8714;
wire v_8715;
wire v_8716;
wire v_8717;
wire v_8718;
wire v_8719;
wire v_8720;
wire v_8721;
wire v_8722;
wire v_8723;
wire v_8724;
wire v_8725;
wire v_8726;
wire v_8727;
wire v_8728;
wire v_8729;
wire v_8730;
wire v_8731;
wire v_8732;
wire v_8733;
wire v_8734;
wire v_8735;
wire v_8736;
wire v_8737;
wire v_8738;
wire v_8739;
wire v_8740;
wire v_8741;
wire v_8742;
wire v_8743;
wire v_8745;
wire v_8746;
wire v_8747;
wire v_8749;
wire v_8750;
wire v_8751;
wire v_8752;
wire v_8753;
wire v_8754;
wire v_8755;
wire v_8756;
wire v_8757;
wire v_8758;
wire v_8759;
wire v_8760;
wire v_8761;
wire v_8762;
wire v_8763;
wire v_8764;
wire v_8765;
wire v_8766;
wire v_8767;
wire v_8768;
wire v_8769;
wire v_8770;
wire v_8771;
wire v_8772;
wire v_8773;
wire v_8774;
wire v_8775;
wire v_8776;
wire v_8777;
wire v_8778;
wire v_8779;
wire v_8780;
wire v_8781;
wire v_8782;
wire v_8783;
wire v_8784;
wire v_8785;
wire v_8786;
wire v_8787;
wire v_8788;
wire v_8789;
wire v_8790;
wire v_8791;
wire v_8792;
wire v_8793;
wire v_8794;
wire v_8795;
wire v_8796;
wire v_8797;
wire v_8798;
wire v_8799;
wire v_8800;
wire v_8801;
wire v_8802;
wire v_8803;
wire v_8804;
wire v_8805;
wire v_8806;
wire v_8807;
wire v_8808;
wire v_8809;
wire v_8810;
wire v_8811;
wire v_8812;
wire v_8813;
wire v_8814;
wire v_8815;
wire v_8816;
wire v_8817;
wire v_8818;
wire v_8819;
wire v_8820;
wire v_8821;
wire v_8822;
wire v_8823;
wire v_8824;
wire v_8825;
wire v_8826;
wire v_8827;
wire v_8828;
wire v_8829;
wire v_8830;
wire v_8831;
wire v_8832;
wire v_8833;
wire v_8834;
wire v_8835;
wire v_8836;
wire v_8837;
wire v_8838;
wire v_8839;
wire v_8840;
wire v_8841;
wire v_8842;
wire v_8843;
wire v_8845;
wire v_8846;
wire v_8847;
wire v_8848;
wire v_8849;
wire v_8850;
wire v_8851;
wire v_8852;
wire v_8853;
wire v_8854;
wire v_8855;
wire v_8856;
wire v_8857;
wire v_8858;
wire v_8859;
wire v_8860;
wire v_8861;
wire v_8862;
wire v_8863;
wire v_8864;
wire v_8865;
wire v_8866;
wire v_8867;
wire v_8868;
wire v_8869;
wire v_8870;
wire v_8871;
wire v_8872;
wire v_8873;
wire v_8874;
wire v_8875;
wire v_8876;
wire v_8877;
wire v_8878;
wire v_8879;
wire v_8880;
wire v_8881;
wire v_8882;
wire v_8883;
wire v_8884;
wire v_8885;
wire v_8886;
wire v_8887;
wire v_8888;
wire v_8889;
wire v_8890;
wire v_8891;
wire v_8892;
wire v_8893;
wire v_8894;
wire v_8895;
wire v_8896;
wire v_8897;
wire v_8898;
wire v_8899;
wire v_8900;
wire v_8901;
wire v_8902;
wire v_8903;
wire v_8904;
wire v_8905;
wire v_8906;
wire v_8907;
wire v_8908;
wire v_8909;
wire v_8910;
wire v_8911;
wire v_8912;
wire v_8913;
wire v_8914;
wire v_8915;
wire v_8916;
wire v_8917;
wire v_8918;
wire v_8919;
wire v_8920;
wire v_8921;
wire v_8922;
wire v_8923;
wire v_8924;
wire v_8925;
wire v_8926;
wire v_8927;
wire v_8928;
wire v_8929;
wire v_8930;
wire v_8931;
wire v_8932;
wire v_8933;
wire v_8934;
wire v_8935;
wire v_8936;
wire v_8937;
wire v_8938;
wire v_8939;
wire v_8940;
wire v_8941;
wire v_8942;
wire v_8943;
wire v_8944;
wire v_8945;
wire v_8946;
wire v_8947;
wire v_8948;
wire v_8949;
wire v_8950;
wire v_8951;
wire v_8952;
wire v_8953;
wire v_8954;
wire v_8955;
wire v_8956;
wire v_8957;
wire v_8958;
wire v_8959;
wire v_8960;
wire v_8961;
wire v_8962;
wire v_8963;
wire v_8964;
wire v_8965;
wire v_8966;
wire v_8967;
wire v_8968;
wire v_8969;
wire v_8970;
wire v_8971;
wire v_8972;
wire v_8973;
wire v_8974;
wire v_8975;
wire v_8976;
wire v_8977;
wire v_8978;
wire v_8979;
wire v_8980;
wire v_8981;
wire v_8982;
wire v_8983;
wire v_8984;
wire v_8985;
wire v_8986;
wire v_8987;
wire v_8988;
wire v_8989;
wire v_8990;
wire v_8991;
wire v_8992;
wire v_8993;
wire v_8994;
wire v_8995;
wire v_8996;
wire v_8997;
wire v_8998;
wire v_8999;
wire v_9000;
wire v_9001;
wire v_9002;
wire v_9003;
wire v_9004;
wire v_9005;
wire v_9006;
wire v_9007;
wire v_9008;
wire v_9009;
wire v_9010;
wire v_9011;
wire v_9012;
wire v_9013;
wire v_9014;
wire v_9015;
wire v_9016;
wire v_9017;
wire v_9018;
wire v_9019;
wire v_9020;
wire v_9021;
wire v_9022;
wire v_9023;
wire v_9024;
wire v_9025;
wire v_9026;
wire v_9027;
wire v_9028;
wire v_9029;
wire v_9030;
wire v_9031;
wire v_9032;
wire v_9033;
wire v_9034;
wire v_9035;
wire v_9036;
wire v_9037;
wire v_9038;
wire v_9039;
wire v_9040;
wire v_9041;
wire v_9042;
wire v_9043;
wire v_9044;
wire v_9045;
wire v_9046;
wire v_9047;
wire v_9048;
wire v_9049;
wire v_9050;
wire v_9051;
wire v_9052;
wire v_9053;
wire v_9054;
wire v_9055;
wire v_9056;
wire v_9057;
wire v_9058;
wire v_9059;
wire v_9060;
wire v_9061;
wire v_9062;
wire v_9063;
wire v_9064;
wire v_9065;
wire v_9066;
wire v_9067;
wire v_9068;
wire v_9069;
wire v_9070;
wire v_9071;
wire v_9072;
wire v_9073;
wire v_9074;
wire v_9075;
wire v_9076;
wire v_9077;
wire v_9078;
wire v_9079;
wire v_9080;
wire v_9081;
wire v_9082;
wire v_9083;
wire v_9084;
wire v_9085;
wire v_9086;
wire v_9087;
wire v_9088;
wire v_9089;
wire v_9090;
wire v_9091;
wire v_9092;
wire v_9093;
wire v_9094;
wire v_9095;
wire v_9096;
wire v_9097;
wire v_9098;
wire v_9099;
wire v_9100;
wire v_9101;
wire v_9102;
wire v_9103;
wire v_9104;
wire v_9105;
wire v_9106;
wire v_9107;
wire v_9108;
wire v_9109;
wire v_9110;
wire v_9111;
wire v_9112;
wire v_9113;
wire v_9114;
wire v_9115;
wire v_9116;
wire v_9117;
wire v_9118;
wire v_9119;
wire v_9120;
wire v_9121;
wire v_9122;
wire v_9123;
wire v_9124;
wire v_9125;
wire v_9126;
wire v_9127;
wire v_9128;
wire v_9129;
wire v_9130;
wire v_9131;
wire v_9132;
wire v_9133;
wire v_9134;
wire v_9135;
wire v_9136;
wire v_9137;
wire v_9138;
wire v_9139;
wire v_9140;
wire v_9141;
wire v_9142;
wire v_9143;
wire v_9144;
wire v_9145;
wire v_9146;
wire v_9147;
wire v_9148;
wire v_9149;
wire v_9150;
wire v_9151;
wire v_9152;
wire v_9153;
wire v_9154;
wire v_9155;
wire v_9156;
wire v_9157;
wire v_9158;
wire v_9159;
wire v_9160;
wire v_9161;
wire v_9162;
wire v_9163;
wire v_9164;
wire v_9165;
wire v_9166;
wire v_9167;
wire v_9168;
wire v_9169;
wire v_9170;
wire v_9171;
wire v_9172;
wire v_9173;
wire v_9174;
wire v_9175;
wire v_9176;
wire v_9177;
wire v_9178;
wire v_9179;
wire v_9180;
wire v_9181;
wire v_9182;
wire v_9183;
wire v_9184;
wire v_9185;
wire v_9186;
wire v_9187;
wire v_9188;
wire v_9189;
wire v_9190;
wire v_9191;
wire v_9192;
wire v_9193;
wire v_9194;
wire v_9195;
wire v_9196;
wire v_9197;
wire v_9198;
wire v_9199;
wire v_9200;
wire v_9201;
wire v_9202;
wire v_9203;
wire v_9204;
wire v_9205;
wire v_9206;
wire v_9207;
wire v_9208;
wire v_9209;
wire v_9210;
wire v_9211;
wire v_9212;
wire v_9213;
wire v_9214;
wire v_9215;
wire v_9216;
wire v_9217;
wire v_9218;
wire v_9219;
wire v_9220;
wire v_9221;
wire v_9222;
wire v_9223;
wire v_9224;
wire v_9225;
wire v_9226;
wire v_9227;
wire v_9228;
wire v_9229;
wire v_9230;
wire v_9231;
wire v_9232;
wire v_9233;
wire v_9234;
wire v_9235;
wire v_9236;
wire v_9237;
wire v_9238;
wire v_9239;
wire v_9240;
wire v_9241;
wire v_9242;
wire v_9243;
wire v_9244;
wire v_9245;
wire v_9246;
wire v_9247;
wire v_9248;
wire v_9249;
wire v_9250;
wire v_9251;
wire v_9252;
wire v_9253;
wire v_9254;
wire v_9255;
wire v_9256;
wire v_9257;
wire v_9258;
wire v_9259;
wire v_9260;
wire v_9261;
wire v_9262;
wire v_9263;
wire v_9264;
wire v_9265;
wire v_9266;
wire v_9267;
wire v_9268;
wire v_9269;
wire v_9270;
wire v_9271;
wire v_9272;
wire v_9273;
wire v_9274;
wire v_9275;
wire v_9276;
wire v_9277;
wire v_9278;
wire v_9279;
wire v_9280;
wire v_9281;
wire v_9282;
wire v_9283;
wire v_9284;
wire v_9285;
wire v_9286;
wire v_9287;
wire v_9288;
wire v_9289;
wire v_9290;
wire v_9291;
wire v_9292;
wire v_9293;
wire v_9294;
wire v_9295;
wire v_9296;
wire v_9297;
wire v_9298;
wire v_9299;
wire v_9301;
wire v_9302;
wire v_9303;
wire v_9304;
wire v_9305;
wire v_9306;
wire v_9307;
wire v_9308;
wire v_9309;
wire v_9310;
wire v_9311;
wire v_9312;
wire v_9313;
wire v_9314;
wire v_9315;
wire v_9316;
wire v_9317;
wire v_9318;
wire v_9319;
wire v_9321;
wire v_9322;
wire v_9323;
wire v_9324;
wire v_9325;
wire v_9326;
wire v_9327;
wire v_9328;
wire v_9329;
wire v_9330;
wire v_9331;
wire v_9332;
wire v_9333;
wire v_9334;
wire v_9335;
wire v_9336;
wire v_9337;
wire v_9338;
wire v_9339;
wire v_9340;
wire v_9341;
wire v_9342;
wire v_9343;
wire v_9344;
wire v_9345;
wire v_9346;
wire v_9347;
wire v_9348;
wire v_9349;
wire v_9350;
wire v_9351;
wire v_9352;
wire v_9353;
wire v_9354;
wire v_9355;
wire v_9356;
wire v_9357;
wire v_9358;
wire v_9359;
wire v_9360;
wire v_9361;
wire v_9362;
wire v_9363;
wire v_9364;
wire v_9365;
wire v_9366;
wire v_9367;
wire v_9368;
wire v_9369;
wire v_9370;
wire v_9372;
wire v_9373;
wire v_9374;
wire v_9375;
wire v_9376;
wire v_9377;
wire v_9378;
wire v_9379;
wire v_9380;
wire v_9381;
wire v_9382;
wire v_9383;
wire v_9384;
wire v_9385;
wire v_9386;
wire v_9387;
wire v_9388;
wire v_9390;
wire v_9391;
wire v_9392;
wire v_9393;
wire v_9394;
wire v_9395;
wire v_9396;
wire v_9397;
wire v_9398;
wire v_9399;
wire v_9400;
wire v_9401;
wire v_9402;
wire v_9403;
wire v_9404;
wire v_9405;
wire v_9406;
wire v_9407;
wire v_9408;
wire v_9409;
wire v_9410;
wire v_9411;
wire v_9412;
wire v_9413;
wire v_9414;
wire v_9415;
wire v_9416;
wire v_9417;
wire v_9418;
wire v_9419;
wire v_9420;
wire v_9421;
wire v_9422;
wire v_9423;
wire v_9424;
wire v_9425;
wire v_9426;
wire v_9427;
wire v_9428;
wire v_9429;
wire v_9430;
wire v_9431;
wire v_9432;
wire v_9433;
wire v_9434;
wire v_9435;
wire v_9436;
wire v_9437;
wire v_9438;
wire v_9439;
wire v_9440;
wire v_9441;
wire v_9442;
wire v_9443;
wire v_9444;
wire v_9445;
wire v_9446;
wire v_9447;
wire v_9448;
wire v_9449;
wire v_9450;
wire v_9451;
wire v_9452;
wire v_9453;
wire v_9454;
wire v_9455;
wire v_9456;
wire v_9457;
wire v_9458;
wire v_9459;
wire v_9460;
wire v_9461;
wire v_9462;
wire v_9463;
wire v_9464;
wire v_9465;
wire v_9466;
wire v_9467;
wire v_9468;
wire v_9469;
wire v_9470;
wire v_9471;
wire v_9472;
wire v_9473;
wire v_9474;
wire v_9475;
wire v_9476;
wire v_9477;
wire v_9478;
wire v_9479;
wire v_9480;
wire v_9481;
wire v_9482;
wire v_9483;
wire v_9484;
wire v_9485;
wire v_9486;
wire v_9487;
wire v_9488;
wire v_9489;
wire v_9490;
wire v_9491;
wire v_9492;
wire v_9493;
wire v_9494;
wire v_9495;
wire v_9496;
wire v_9497;
wire v_9498;
wire v_9499;
wire v_9500;
wire v_9501;
wire v_9502;
wire v_9503;
wire v_9504;
wire v_9505;
wire v_9506;
wire v_9507;
wire v_9508;
wire v_9509;
wire v_9510;
wire v_9511;
wire v_9512;
wire v_9513;
wire v_9514;
wire v_9515;
wire v_9516;
wire v_9517;
wire v_9518;
wire v_9519;
wire v_9520;
wire v_9521;
wire v_9522;
wire v_9523;
wire v_9524;
wire v_9525;
wire v_9526;
wire v_9527;
wire v_9528;
wire v_9529;
wire v_9530;
wire v_9531;
wire v_9532;
wire v_9533;
wire v_9534;
wire v_9535;
wire v_9536;
wire v_9537;
wire v_9538;
wire v_9539;
wire v_9540;
wire v_9541;
wire v_9542;
wire v_9543;
wire v_9544;
wire v_9545;
wire v_9546;
wire v_9547;
wire v_9548;
wire v_9549;
wire v_9550;
wire v_9551;
wire v_9552;
wire v_9553;
wire v_9554;
wire v_9555;
wire v_9556;
wire v_9557;
wire v_9558;
wire v_9559;
wire v_9560;
wire v_9561;
wire v_9562;
wire v_9563;
wire v_9564;
wire v_9565;
wire v_9566;
wire v_9567;
wire v_9568;
wire v_9569;
wire v_9570;
wire v_9571;
wire v_9572;
wire v_9573;
wire v_9574;
wire v_9575;
wire v_9576;
wire v_9577;
wire v_9578;
wire v_9579;
wire v_9580;
wire v_9581;
wire v_9582;
wire v_9583;
wire v_9584;
wire v_9585;
wire v_9586;
wire v_9587;
wire v_9588;
wire v_9589;
wire v_9590;
wire v_9591;
wire v_9592;
wire v_9593;
wire v_9594;
wire v_9595;
wire v_9596;
wire v_9597;
wire v_9598;
wire v_9599;
wire v_9600;
wire v_9601;
wire v_9602;
wire v_9603;
wire v_9604;
wire v_9605;
wire v_9606;
wire v_9607;
wire v_9608;
wire v_9609;
wire v_9610;
wire v_9611;
wire v_9612;
wire v_9613;
wire v_9614;
wire v_9615;
wire v_9616;
wire v_9617;
wire v_9618;
wire v_9619;
wire v_9620;
wire v_9621;
wire v_9622;
wire v_9623;
wire v_9624;
wire v_9625;
wire v_9626;
wire v_9627;
wire v_9628;
wire v_9629;
wire v_9630;
wire v_9631;
wire v_9632;
wire v_9633;
wire v_9634;
wire v_9635;
wire v_9636;
wire v_9637;
wire v_9638;
wire v_9639;
wire v_9640;
wire v_9641;
wire v_9642;
wire v_9643;
wire v_9644;
wire v_9645;
wire v_9646;
wire v_9647;
wire v_9648;
wire v_9649;
wire v_9650;
wire v_9651;
wire v_9652;
wire v_9653;
wire v_9654;
wire v_9655;
wire v_9656;
wire v_9657;
wire v_9658;
wire v_9659;
wire v_9660;
wire v_9661;
wire v_9662;
wire v_9663;
wire v_9664;
wire v_9665;
wire v_9666;
wire v_9667;
wire v_9668;
wire v_9669;
wire v_9670;
wire v_9671;
wire v_9672;
wire v_9673;
wire v_9674;
wire v_9675;
wire v_9676;
wire v_9677;
wire v_9678;
wire v_9679;
wire v_9680;
wire v_9681;
wire v_9682;
wire v_9683;
wire v_9684;
wire v_9685;
wire v_9686;
wire v_9687;
wire v_9688;
wire v_9689;
wire v_9690;
wire v_9691;
wire v_9692;
wire v_9693;
wire v_9694;
wire v_9695;
wire v_9696;
wire v_9697;
wire v_9698;
wire v_9699;
wire v_9700;
wire v_9701;
wire v_9702;
wire v_9703;
wire v_9704;
wire v_9705;
wire v_9706;
wire v_9707;
wire v_9708;
wire v_9709;
wire v_9710;
wire v_9711;
wire v_9712;
wire v_9713;
wire v_9714;
wire v_9715;
wire v_9716;
wire v_9717;
wire v_9718;
wire v_9719;
wire v_9720;
wire v_9721;
wire v_9722;
wire v_9723;
wire v_9724;
wire v_9725;
wire v_9726;
wire v_9727;
wire v_9728;
wire v_9729;
wire v_9730;
wire v_9731;
wire v_9732;
wire v_9733;
wire v_9734;
wire v_9735;
wire v_9736;
wire v_9737;
wire v_9738;
wire v_9739;
wire v_9740;
wire v_9741;
wire v_9742;
wire v_9743;
wire v_9744;
wire v_9745;
wire v_9746;
wire v_9747;
wire v_9748;
wire v_9749;
wire v_9750;
wire v_9751;
wire v_9752;
wire v_9753;
wire v_9754;
wire v_9755;
wire v_9756;
wire v_9757;
wire v_9758;
wire v_9759;
wire v_9760;
wire v_9761;
wire v_9762;
wire v_9764;
wire v_9765;
wire v_9766;
wire v_9767;
wire v_9768;
wire v_9769;
wire v_9770;
wire v_9771;
wire v_9772;
wire v_9773;
wire v_9774;
wire v_9775;
wire v_9776;
wire v_9777;
wire v_9778;
wire v_9779;
wire v_9780;
wire v_9781;
wire v_9782;
wire v_9784;
wire v_9785;
wire v_9786;
wire v_9787;
wire v_9788;
wire v_9789;
wire v_9790;
wire v_9791;
wire v_9792;
wire v_9793;
wire v_9794;
wire v_9795;
wire v_9796;
wire v_9797;
wire v_9798;
wire v_9799;
wire v_9800;
wire v_9801;
wire v_9802;
wire v_9803;
wire v_9804;
wire v_9805;
wire v_9806;
wire v_9807;
wire v_9808;
wire v_9809;
wire v_9810;
wire v_9811;
wire v_9812;
wire v_9813;
wire v_9814;
wire v_9815;
wire v_9816;
wire v_9817;
wire v_9818;
wire v_9819;
wire v_9820;
wire v_9821;
wire v_9822;
wire v_9823;
wire v_9824;
wire v_9825;
wire v_9826;
wire v_9827;
wire v_9828;
wire v_9829;
wire v_9830;
wire v_9831;
wire v_9832;
wire v_9833;
wire v_9835;
wire v_9836;
wire v_9837;
wire v_9838;
wire v_9839;
wire v_9840;
wire v_9841;
wire v_9842;
wire v_9843;
wire v_9844;
wire v_9845;
wire v_9846;
wire v_9847;
wire v_9848;
wire v_9849;
wire v_9850;
wire v_9851;
wire v_9853;
wire v_9854;
wire v_9855;
wire v_9856;
wire v_9857;
wire v_9858;
wire v_9859;
wire v_9860;
wire v_9861;
wire v_9862;
wire v_9863;
wire v_9864;
wire v_9865;
wire v_9866;
wire v_9867;
wire v_9868;
wire v_9869;
wire v_9870;
wire v_9871;
wire v_9872;
wire v_9873;
wire v_9874;
wire v_9875;
wire v_9876;
wire v_9877;
wire v_9878;
wire v_9879;
wire v_9880;
wire v_9881;
wire v_9882;
wire v_9883;
wire v_9884;
wire v_9885;
wire v_9886;
wire v_9887;
wire v_9888;
wire v_9889;
wire v_9890;
wire v_9891;
wire v_9892;
wire v_9893;
wire v_9894;
wire v_9895;
wire v_9896;
wire v_9897;
wire v_9898;
wire v_9899;
wire v_9900;
wire v_9901;
wire v_9902;
wire v_9903;
wire v_9904;
wire v_9905;
wire v_9906;
wire v_9907;
wire v_9908;
wire v_9909;
wire v_9910;
wire v_9911;
wire v_9912;
wire v_9913;
wire v_9914;
wire v_9915;
wire v_9916;
wire v_9917;
wire v_9918;
wire v_9919;
wire v_9920;
wire v_9921;
wire v_9922;
wire v_9923;
wire v_9924;
wire v_9925;
wire v_9926;
wire v_9927;
wire v_9928;
wire v_9929;
wire v_9930;
wire v_9931;
wire v_9932;
wire v_9933;
wire v_9934;
wire v_9935;
wire v_9936;
wire v_9937;
wire v_9938;
wire v_9939;
wire v_9940;
wire v_9941;
wire v_9942;
wire v_9943;
wire v_9944;
wire v_9945;
wire v_9946;
wire v_9947;
wire v_9948;
wire v_9949;
wire v_9950;
wire v_9951;
wire v_9952;
wire v_9953;
wire v_9954;
wire v_9955;
wire v_9956;
wire v_9957;
wire v_9958;
wire v_9959;
wire v_9960;
wire v_9961;
wire v_9962;
wire v_9963;
wire v_9964;
wire v_9965;
wire v_9966;
wire v_9967;
wire v_9968;
wire v_9969;
wire v_9970;
wire v_9971;
wire v_9972;
wire v_9973;
wire v_9974;
wire v_9975;
wire v_9976;
wire v_9977;
wire v_9978;
wire v_9979;
wire v_9980;
wire v_9981;
wire v_9982;
wire v_9983;
wire v_9984;
wire v_9985;
wire v_9986;
wire v_9987;
wire v_9988;
wire v_9989;
wire v_9990;
wire v_9991;
wire v_9992;
wire v_9993;
wire v_9994;
wire v_9995;
wire v_9996;
wire v_9997;
wire v_9998;
wire v_9999;
wire v_10000;
wire v_10001;
wire v_10002;
wire v_10003;
wire v_10004;
wire v_10005;
wire v_10006;
wire v_10007;
wire v_10008;
wire v_10009;
wire v_10010;
wire v_10011;
wire v_10012;
wire v_10013;
wire v_10014;
wire v_10015;
wire v_10016;
wire v_10017;
wire v_10018;
wire v_10019;
wire v_10020;
wire v_10021;
wire v_10022;
wire v_10023;
wire v_10024;
wire v_10025;
wire v_10026;
wire v_10027;
wire v_10028;
wire v_10029;
wire v_10030;
wire v_10031;
wire v_10032;
wire v_10033;
wire v_10034;
wire v_10035;
wire v_10036;
wire v_10037;
wire v_10038;
wire v_10039;
wire v_10040;
wire v_10041;
wire v_10042;
wire v_10043;
wire v_10044;
wire v_10045;
wire v_10046;
wire v_10047;
wire v_10048;
wire v_10049;
wire v_10050;
wire v_10051;
wire v_10052;
wire v_10053;
wire v_10054;
wire v_10055;
wire v_10056;
wire v_10057;
wire v_10058;
wire v_10059;
wire v_10060;
wire v_10061;
wire v_10062;
wire v_10063;
wire v_10064;
wire v_10065;
wire v_10066;
wire v_10067;
wire v_10068;
wire v_10069;
wire v_10070;
wire v_10071;
wire v_10072;
wire v_10073;
wire v_10074;
wire v_10075;
wire v_10076;
wire v_10077;
wire v_10078;
wire v_10079;
wire v_10080;
wire v_10081;
wire v_10082;
wire v_10083;
wire v_10084;
wire v_10085;
wire v_10086;
wire v_10087;
wire v_10088;
wire v_10089;
wire v_10090;
wire v_10091;
wire v_10092;
wire v_10093;
wire v_10094;
wire v_10095;
wire v_10096;
wire v_10097;
wire v_10098;
wire v_10099;
wire v_10100;
wire v_10101;
wire v_10102;
wire v_10103;
wire v_10105;
wire v_10106;
wire v_10107;
wire v_10108;
wire v_10109;
wire v_10110;
wire v_10111;
wire v_10112;
wire v_10113;
wire v_10114;
wire v_10115;
wire v_10116;
wire v_10117;
wire v_10118;
wire v_10119;
wire v_10120;
wire v_10121;
wire v_10122;
wire v_10123;
wire v_10124;
wire v_10125;
wire v_10126;
wire v_10127;
wire v_10128;
wire v_10129;
wire v_10130;
wire v_10131;
wire v_10132;
wire v_10133;
wire v_10134;
wire v_10135;
wire v_10136;
wire v_10137;
wire v_10138;
wire v_10139;
wire v_10140;
wire v_10141;
wire v_10142;
wire v_10143;
wire v_10144;
wire v_10145;
wire v_10146;
wire v_10147;
wire v_10148;
wire v_10149;
wire v_10150;
wire v_10151;
wire v_10152;
wire v_10153;
wire v_10154;
wire v_10155;
wire v_10156;
wire v_10157;
wire v_10158;
wire v_10159;
wire v_10160;
wire v_10161;
wire v_10162;
wire v_10163;
wire v_10164;
wire v_10165;
wire v_10166;
wire v_10167;
wire v_10168;
wire v_10169;
wire v_10170;
wire v_10171;
wire v_10172;
wire v_10173;
wire v_10174;
wire v_10175;
wire v_10176;
wire v_10177;
wire v_10178;
wire v_10179;
wire v_10180;
wire v_10181;
wire v_10182;
wire v_10183;
wire v_10184;
wire v_10185;
wire v_10186;
wire v_10187;
wire v_10188;
wire v_10189;
wire v_10190;
wire v_10191;
wire v_10192;
wire v_10193;
wire v_10194;
wire v_10195;
wire v_10196;
wire v_10197;
wire v_10198;
wire v_10199;
wire v_10200;
wire v_10201;
wire v_10202;
wire v_10203;
wire v_10204;
wire v_10205;
wire v_10206;
wire v_10207;
wire v_10208;
wire v_10209;
wire v_10210;
wire v_10211;
wire v_10212;
wire v_10213;
wire v_10214;
wire v_10215;
wire v_10216;
wire v_10217;
wire v_10218;
wire v_10219;
wire v_10220;
wire v_10221;
wire v_10222;
wire v_10223;
wire v_10224;
wire v_10225;
wire v_10226;
wire v_10227;
wire v_10228;
wire v_10230;
wire v_10231;
wire v_10232;
wire v_10233;
wire v_10234;
wire v_10235;
wire v_10236;
wire v_10237;
wire v_10238;
wire v_10239;
wire v_10240;
wire v_10241;
wire v_10242;
wire v_10243;
wire v_10244;
wire v_10245;
wire v_10246;
wire v_10247;
wire v_10248;
wire v_10250;
wire v_10251;
wire v_10252;
wire v_10253;
wire v_10254;
wire v_10255;
wire v_10256;
wire v_10257;
wire v_10258;
wire v_10259;
wire v_10260;
wire v_10261;
wire v_10262;
wire v_10263;
wire v_10264;
wire v_10265;
wire v_10266;
wire v_10267;
wire v_10268;
wire v_10269;
wire v_10270;
wire v_10271;
wire v_10272;
wire v_10273;
wire v_10274;
wire v_10275;
wire v_10276;
wire v_10277;
wire v_10278;
wire v_10279;
wire v_10280;
wire v_10281;
wire v_10282;
wire v_10283;
wire v_10284;
wire v_10285;
wire v_10286;
wire v_10287;
wire v_10288;
wire v_10289;
wire v_10290;
wire v_10291;
wire v_10292;
wire v_10293;
wire v_10294;
wire v_10295;
wire v_10296;
wire v_10297;
wire v_10298;
wire v_10299;
wire v_10301;
wire v_10302;
wire v_10303;
wire v_10304;
wire v_10305;
wire v_10306;
wire v_10307;
wire v_10308;
wire v_10309;
wire v_10310;
wire v_10311;
wire v_10312;
wire v_10313;
wire v_10314;
wire v_10315;
wire v_10316;
wire v_10317;
wire v_10319;
wire v_10320;
wire v_10321;
wire v_10322;
wire v_10323;
wire v_10324;
wire v_10325;
wire v_10326;
wire v_10327;
wire v_10328;
wire v_10329;
wire v_10330;
wire v_10331;
wire v_10332;
wire v_10333;
wire v_10334;
wire v_10335;
wire v_10336;
wire v_10337;
wire v_10338;
wire v_10339;
wire v_10340;
wire v_10341;
wire v_10342;
wire v_10343;
wire v_10344;
wire v_10345;
wire v_10346;
wire v_10347;
wire v_10348;
wire v_10349;
wire v_10350;
wire v_10351;
wire v_10352;
wire v_10353;
wire v_10354;
wire v_10355;
wire v_10356;
wire v_10357;
wire v_10358;
wire v_10359;
wire v_10360;
wire v_10361;
wire v_10362;
wire v_10363;
wire v_10364;
wire v_10365;
wire v_10366;
wire v_10367;
wire v_10368;
wire v_10369;
wire v_10370;
wire v_10371;
wire v_10372;
wire v_10373;
wire v_10374;
wire v_10375;
wire v_10376;
wire v_10377;
wire v_10378;
wire v_10379;
wire v_10380;
wire v_10381;
wire v_10382;
wire v_10383;
wire v_10384;
wire v_10385;
wire v_10386;
wire v_10387;
wire v_10388;
wire v_10389;
wire v_10390;
wire v_10391;
wire v_10392;
wire v_10393;
wire v_10394;
wire v_10395;
wire v_10396;
wire v_10397;
wire v_10398;
wire v_10399;
wire v_10400;
wire v_10401;
wire v_10402;
wire v_10403;
wire v_10404;
wire v_10405;
wire v_10406;
wire v_10407;
wire v_10408;
wire v_10409;
wire v_10410;
wire v_10411;
wire v_10412;
wire v_10413;
wire v_10414;
wire v_10415;
wire v_10416;
wire v_10417;
wire v_10418;
wire v_10419;
wire v_10420;
wire v_10421;
wire v_10422;
wire v_10423;
wire v_10424;
wire v_10425;
wire v_10426;
wire v_10427;
wire v_10428;
wire v_10429;
wire v_10430;
wire v_10431;
wire v_10432;
wire v_10433;
wire v_10434;
wire v_10435;
wire v_10436;
wire v_10437;
wire v_10438;
wire v_10439;
wire v_10440;
wire v_10441;
wire v_10442;
wire v_10443;
wire v_10444;
wire v_10445;
wire v_10446;
wire v_10447;
wire v_10448;
wire v_10449;
wire v_10450;
wire v_10451;
wire v_10452;
wire v_10453;
wire v_10454;
wire v_10455;
wire v_10456;
wire v_10457;
wire v_10458;
wire v_10459;
wire v_10460;
wire v_10461;
wire v_10462;
wire v_10463;
wire v_10464;
wire v_10465;
wire v_10466;
wire v_10467;
wire v_10468;
wire v_10469;
wire v_10470;
wire v_10471;
wire v_10472;
wire v_10473;
wire v_10474;
wire v_10475;
wire v_10476;
wire v_10477;
wire v_10478;
wire v_10479;
wire v_10480;
wire v_10481;
wire v_10482;
wire v_10483;
wire v_10484;
wire v_10485;
wire v_10486;
wire v_10487;
wire v_10488;
wire v_10489;
wire v_10490;
wire v_10491;
wire v_10492;
wire v_10493;
wire v_10494;
wire v_10495;
wire v_10496;
wire v_10497;
wire v_10498;
wire v_10499;
wire v_10500;
wire v_10501;
wire v_10502;
wire v_10503;
wire v_10504;
wire v_10505;
wire v_10506;
wire v_10507;
wire v_10508;
wire v_10509;
wire v_10510;
wire v_10511;
wire v_10512;
wire v_10513;
wire v_10514;
wire v_10515;
wire v_10516;
wire v_10517;
wire v_10518;
wire v_10519;
wire v_10520;
wire v_10521;
wire v_10522;
wire v_10523;
wire v_10524;
wire v_10525;
wire v_10526;
wire v_10527;
wire v_10528;
wire v_10529;
wire v_10530;
wire v_10531;
wire v_10532;
wire v_10533;
wire v_10534;
wire v_10535;
wire v_10536;
wire v_10537;
wire v_10538;
wire v_10539;
wire v_10540;
wire v_10541;
wire v_10542;
wire v_10543;
wire v_10544;
wire v_10545;
wire v_10546;
wire v_10547;
wire v_10548;
wire v_10549;
wire v_10550;
wire v_10551;
wire v_10552;
wire v_10553;
wire v_10554;
wire v_10555;
wire v_10556;
wire v_10557;
wire v_10558;
wire v_10559;
wire v_10560;
wire v_10561;
wire v_10562;
wire v_10563;
wire v_10564;
wire v_10565;
wire v_10566;
wire v_10567;
wire v_10568;
wire v_10569;
wire v_10571;
wire v_10572;
wire v_10573;
wire v_10574;
wire v_10575;
wire v_10576;
wire v_10577;
wire v_10578;
wire v_10579;
wire v_10580;
wire v_10581;
wire v_10582;
wire v_10583;
wire v_10584;
wire v_10585;
wire v_10586;
wire v_10587;
wire v_10588;
wire v_10589;
wire v_10590;
wire v_10591;
wire v_10592;
wire v_10593;
wire v_10594;
wire v_10595;
wire v_10596;
wire v_10597;
wire v_10598;
wire v_10599;
wire v_10600;
wire v_10601;
wire v_10602;
wire v_10603;
wire v_10604;
wire v_10605;
wire v_10606;
wire v_10607;
wire v_10608;
wire v_10609;
wire v_10610;
wire v_10611;
wire v_10612;
wire v_10613;
wire v_10614;
wire v_10615;
wire v_10616;
wire v_10617;
wire v_10618;
wire v_10619;
wire v_10620;
wire v_10621;
wire v_10622;
wire v_10623;
wire v_10624;
wire v_10625;
wire v_10626;
wire v_10627;
wire v_10628;
wire v_10629;
wire v_10630;
wire v_10631;
wire v_10632;
wire v_10633;
wire v_10634;
wire v_10635;
wire v_10636;
wire v_10637;
wire v_10638;
wire v_10639;
wire v_10640;
wire v_10641;
wire v_10642;
wire v_10643;
wire v_10644;
wire v_10645;
wire v_10646;
wire v_10647;
wire v_10648;
wire v_10649;
wire v_10650;
wire v_10651;
wire v_10652;
wire v_10653;
wire v_10654;
wire v_10655;
wire v_10656;
wire v_10657;
wire v_10658;
wire v_10659;
wire v_10660;
wire v_10661;
wire v_10662;
wire v_10663;
wire v_10664;
wire v_10665;
wire v_10666;
wire v_10667;
wire v_10668;
wire v_10669;
wire v_10670;
wire v_10671;
wire v_10672;
wire v_10673;
wire v_10674;
wire v_10675;
wire v_10676;
wire v_10677;
wire v_10678;
wire v_10679;
wire v_10680;
wire v_10681;
wire v_10682;
wire v_10683;
wire v_10684;
wire v_10685;
wire v_10686;
wire v_10687;
wire v_10688;
wire v_10689;
wire v_10690;
wire v_10691;
wire v_10692;
wire v_10693;
wire v_10694;
wire v_10696;
wire v_10697;
wire v_10698;
wire v_10699;
wire v_10700;
wire v_10701;
wire v_10702;
wire v_10703;
wire v_10704;
wire v_10705;
wire v_10706;
wire v_10707;
wire v_10708;
wire v_10709;
wire v_10710;
wire v_10711;
wire v_10712;
wire v_10713;
wire v_10714;
wire v_10716;
wire v_10717;
wire v_10718;
wire v_10719;
wire v_10720;
wire v_10721;
wire v_10722;
wire v_10723;
wire v_10724;
wire v_10725;
wire v_10726;
wire v_10727;
wire v_10728;
wire v_10729;
wire v_10730;
wire v_10731;
wire v_10732;
wire v_10733;
wire v_10734;
wire v_10735;
wire v_10736;
wire v_10737;
wire v_10738;
wire v_10739;
wire v_10740;
wire v_10741;
wire v_10742;
wire v_10743;
wire v_10744;
wire v_10745;
wire v_10746;
wire v_10747;
wire v_10748;
wire v_10749;
wire v_10750;
wire v_10751;
wire v_10752;
wire v_10753;
wire v_10754;
wire v_10755;
wire v_10756;
wire v_10757;
wire v_10758;
wire v_10759;
wire v_10760;
wire v_10761;
wire v_10762;
wire v_10763;
wire v_10764;
wire v_10765;
wire v_10767;
wire v_10768;
wire v_10769;
wire v_10770;
wire v_10771;
wire v_10772;
wire v_10773;
wire v_10774;
wire v_10775;
wire v_10776;
wire v_10777;
wire v_10778;
wire v_10779;
wire v_10780;
wire v_10781;
wire v_10782;
wire v_10783;
wire v_10785;
wire v_10786;
wire v_10787;
wire v_10788;
wire v_10789;
wire v_10790;
wire v_10791;
wire v_10792;
wire v_10793;
wire v_10794;
wire v_10795;
wire v_10796;
wire v_10797;
wire v_10798;
wire v_10799;
wire v_10800;
wire v_10801;
wire v_10802;
wire v_10803;
wire v_10804;
wire v_10805;
wire v_10806;
wire v_10807;
wire v_10808;
wire v_10809;
wire v_10810;
wire v_10811;
wire v_10812;
wire v_10813;
wire v_10814;
wire v_10815;
wire v_10816;
wire v_10817;
wire v_10818;
wire v_10819;
wire v_10820;
wire v_10821;
wire v_10822;
wire v_10823;
wire v_10824;
wire v_10825;
wire v_10826;
wire v_10827;
wire v_10828;
wire v_10829;
wire v_10830;
wire v_10831;
wire v_10832;
wire v_10833;
wire v_10834;
wire v_10835;
wire v_10836;
wire v_10837;
wire v_10838;
wire v_10839;
wire v_10840;
wire v_10841;
wire v_10842;
wire v_10843;
wire v_10844;
wire v_10845;
wire v_10846;
wire v_10847;
wire v_10848;
wire v_10849;
wire v_10850;
wire v_10851;
wire v_10852;
wire v_10853;
wire v_10854;
wire v_10855;
wire v_10856;
wire v_10857;
wire v_10858;
wire v_10859;
wire v_10860;
wire v_10861;
wire v_10862;
wire v_10863;
wire v_10864;
wire v_10865;
wire v_10866;
wire v_10867;
wire v_10868;
wire v_10869;
wire v_10870;
wire v_10871;
wire v_10872;
wire v_10873;
wire v_10874;
wire v_10875;
wire v_10876;
wire v_10877;
wire v_10878;
wire v_10879;
wire v_10880;
wire v_10881;
wire v_10882;
wire v_10883;
wire v_10884;
wire v_10885;
wire v_10886;
wire v_10887;
wire v_10888;
wire v_10889;
wire v_10890;
wire v_10891;
wire v_10892;
wire v_10893;
wire v_10894;
wire v_10895;
wire v_10896;
wire v_10897;
wire v_10898;
wire v_10899;
wire v_10900;
wire v_10901;
wire v_10902;
wire v_10903;
wire v_10904;
wire v_10905;
wire v_10906;
wire v_10907;
wire v_10908;
wire v_10909;
wire v_10910;
wire v_10911;
wire v_10912;
wire v_10913;
wire v_10914;
wire v_10915;
wire v_10916;
wire v_10917;
wire v_10918;
wire v_10919;
wire v_10920;
wire v_10921;
wire v_10922;
wire v_10923;
wire v_10924;
wire v_10925;
wire v_10926;
wire v_10927;
wire v_10928;
wire v_10929;
wire v_10930;
wire v_10931;
wire v_10932;
wire v_10933;
wire v_10934;
wire v_10935;
wire v_10936;
wire v_10937;
wire v_10938;
wire v_10939;
wire v_10940;
wire v_10941;
wire v_10942;
wire v_10943;
wire v_10944;
wire v_10945;
wire v_10946;
wire v_10947;
wire v_10948;
wire v_10949;
wire v_10950;
wire v_10951;
wire v_10952;
wire v_10953;
wire v_10954;
wire v_10955;
wire v_10956;
wire v_10957;
wire v_10958;
wire v_10959;
wire v_10960;
wire v_10961;
wire v_10962;
wire v_10963;
wire v_10964;
wire v_10965;
wire v_10966;
wire v_10967;
wire v_10968;
wire v_10969;
wire v_10970;
wire v_10971;
wire v_10972;
wire v_10973;
wire v_10974;
wire v_10975;
wire v_10976;
wire v_10977;
wire v_10978;
wire v_10979;
wire v_10980;
wire v_10981;
wire v_10982;
wire v_10983;
wire v_10984;
wire v_10985;
wire v_10986;
wire v_10987;
wire v_10988;
wire v_10989;
wire v_10990;
wire v_10991;
wire v_10992;
wire v_10993;
wire v_10994;
wire v_10995;
wire v_10996;
wire v_10997;
wire v_10998;
wire v_10999;
wire v_11000;
wire v_11001;
wire v_11002;
wire v_11003;
wire v_11004;
wire v_11005;
wire v_11006;
wire v_11007;
wire v_11008;
wire v_11009;
wire v_11010;
wire v_11011;
wire v_11012;
wire v_11013;
wire v_11014;
wire v_11015;
wire v_11016;
wire v_11017;
wire v_11018;
wire v_11019;
wire v_11020;
wire v_11021;
wire v_11022;
wire v_11023;
wire v_11024;
wire v_11025;
wire v_11026;
wire v_11027;
wire v_11028;
wire v_11029;
wire v_11030;
wire v_11031;
wire v_11032;
wire v_11033;
wire v_11034;
wire v_11035;
wire v_11036;
wire v_11037;
wire v_11038;
wire v_11039;
wire v_11040;
wire v_11041;
wire v_11042;
wire v_11043;
wire v_11044;
wire v_11045;
wire v_11046;
wire v_11047;
wire v_11048;
wire v_11049;
wire v_11050;
wire v_11051;
wire v_11052;
wire v_11053;
wire v_11054;
wire v_11055;
wire v_11056;
wire v_11057;
wire v_11058;
wire v_11059;
wire v_11060;
wire v_11061;
wire v_11062;
wire v_11063;
wire v_11064;
wire v_11065;
wire v_11066;
wire v_11067;
wire v_11068;
wire v_11069;
wire v_11070;
wire v_11071;
wire v_11072;
wire v_11073;
wire v_11074;
wire v_11075;
wire v_11076;
wire v_11077;
wire v_11078;
wire v_11079;
wire v_11080;
wire v_11081;
wire v_11082;
wire v_11083;
wire v_11084;
wire v_11085;
wire v_11086;
wire v_11087;
wire v_11088;
wire v_11089;
wire v_11090;
wire v_11091;
wire v_11092;
wire v_11093;
wire v_11094;
wire v_11095;
wire v_11096;
wire v_11097;
wire v_11098;
wire v_11099;
wire v_11100;
wire v_11101;
wire v_11102;
wire v_11103;
wire v_11104;
wire v_11105;
wire v_11106;
wire v_11107;
wire v_11108;
wire v_11109;
wire v_11110;
wire v_11111;
wire v_11112;
wire v_11113;
wire v_11114;
wire v_11115;
wire v_11116;
wire v_11117;
wire v_11118;
wire v_11119;
wire v_11120;
wire v_11121;
wire v_11122;
wire v_11123;
wire v_11124;
wire v_11125;
wire v_11126;
wire v_11127;
wire v_11128;
wire v_11129;
wire v_11130;
wire v_11131;
wire v_11132;
wire v_11133;
wire v_11134;
wire v_11135;
wire v_11136;
wire v_11137;
wire v_11138;
wire v_11139;
wire v_11140;
wire v_11141;
wire v_11142;
wire v_11143;
wire v_11144;
wire v_11145;
wire v_11146;
wire v_11147;
wire v_11148;
wire v_11149;
wire v_11150;
wire v_11151;
wire v_11152;
wire v_11153;
wire v_11154;
wire v_11155;
wire v_11156;
wire v_11157;
wire v_11158;
wire v_11159;
wire v_11161;
wire v_11162;
wire v_11163;
wire v_11164;
wire v_11165;
wire v_11166;
wire v_11167;
wire v_11168;
wire v_11169;
wire v_11170;
wire v_11171;
wire v_11172;
wire v_11173;
wire v_11174;
wire v_11175;
wire v_11176;
wire v_11177;
wire v_11178;
wire v_11179;
wire v_11181;
wire v_11182;
wire v_11183;
wire v_11184;
wire v_11185;
wire v_11186;
wire v_11187;
wire v_11188;
wire v_11189;
wire v_11190;
wire v_11191;
wire v_11192;
wire v_11193;
wire v_11194;
wire v_11195;
wire v_11196;
wire v_11197;
wire v_11198;
wire v_11199;
wire v_11200;
wire v_11201;
wire v_11202;
wire v_11203;
wire v_11204;
wire v_11205;
wire v_11206;
wire v_11207;
wire v_11208;
wire v_11209;
wire v_11210;
wire v_11211;
wire v_11212;
wire v_11213;
wire v_11214;
wire v_11215;
wire v_11216;
wire v_11217;
wire v_11218;
wire v_11219;
wire v_11220;
wire v_11221;
wire v_11222;
wire v_11223;
wire v_11224;
wire v_11225;
wire v_11226;
wire v_11227;
wire v_11228;
wire v_11229;
wire v_11230;
wire v_11232;
wire v_11233;
wire v_11234;
wire v_11235;
wire v_11236;
wire v_11237;
wire v_11238;
wire v_11239;
wire v_11240;
wire v_11241;
wire v_11242;
wire v_11243;
wire v_11244;
wire v_11245;
wire v_11246;
wire v_11247;
wire v_11248;
wire v_11250;
wire v_11251;
wire v_11252;
wire v_11253;
wire v_11254;
wire v_11255;
wire v_11256;
wire v_11257;
wire v_11258;
wire v_11259;
wire v_11260;
wire v_11261;
wire v_11262;
wire v_11263;
wire v_11264;
wire v_11265;
wire v_11266;
wire v_11267;
wire v_11268;
wire v_11269;
wire v_11270;
wire v_11271;
wire v_11272;
wire v_11273;
wire v_11274;
wire v_11275;
wire v_11276;
wire v_11277;
wire v_11278;
wire v_11279;
wire v_11280;
wire v_11281;
wire v_11282;
wire v_11283;
wire v_11284;
wire v_11285;
wire v_11286;
wire v_11287;
wire v_11288;
wire v_11289;
wire v_11290;
wire v_11291;
wire v_11292;
wire v_11293;
wire v_11294;
wire v_11295;
wire v_11296;
wire v_11297;
wire v_11298;
wire v_11299;
wire v_11300;
wire v_11301;
wire v_11302;
wire v_11303;
wire v_11304;
wire v_11305;
wire v_11306;
wire v_11307;
wire v_11308;
wire v_11309;
wire v_11310;
wire v_11311;
wire v_11312;
wire v_11313;
wire v_11314;
wire v_11315;
wire v_11316;
wire v_11317;
wire v_11318;
wire v_11319;
wire v_11320;
wire v_11321;
wire v_11322;
wire v_11323;
wire v_11324;
wire v_11325;
wire v_11326;
wire v_11327;
wire v_11328;
wire v_11329;
wire v_11330;
wire v_11331;
wire v_11332;
wire v_11333;
wire v_11334;
wire v_11335;
wire v_11336;
wire v_11337;
wire v_11338;
wire v_11339;
wire v_11340;
wire v_11341;
wire v_11342;
wire v_11343;
wire v_11344;
wire v_11345;
wire v_11346;
wire v_11347;
wire v_11348;
wire v_11349;
wire v_11350;
wire v_11351;
wire v_11352;
wire v_11353;
wire v_11354;
wire v_11355;
wire v_11356;
wire v_11357;
wire v_11358;
wire v_11359;
wire v_11360;
wire v_11361;
wire v_11362;
wire v_11363;
wire v_11364;
wire v_11365;
wire v_11366;
wire v_11367;
wire v_11368;
wire v_11369;
wire v_11370;
wire v_11371;
wire v_11372;
wire v_11373;
wire v_11374;
wire v_11375;
wire v_11376;
wire v_11377;
wire v_11378;
wire v_11379;
wire v_11380;
wire v_11381;
wire v_11382;
wire v_11383;
wire v_11384;
wire v_11385;
wire v_11386;
wire v_11387;
wire v_11388;
wire v_11389;
wire v_11390;
wire v_11391;
wire v_11392;
wire v_11393;
wire v_11394;
wire v_11395;
wire v_11396;
wire v_11397;
wire v_11398;
wire v_11399;
wire v_11400;
wire v_11401;
wire v_11402;
wire v_11403;
wire v_11404;
wire v_11405;
wire v_11406;
wire v_11407;
wire v_11408;
wire v_11409;
wire v_11410;
wire v_11411;
wire v_11412;
wire v_11413;
wire v_11414;
wire v_11415;
wire v_11416;
wire v_11417;
wire v_11418;
wire v_11419;
wire v_11420;
wire v_11421;
wire v_11422;
wire v_11423;
wire v_11424;
wire v_11425;
wire v_11426;
wire v_11427;
wire v_11428;
wire v_11429;
wire v_11430;
wire v_11431;
wire v_11432;
wire v_11433;
wire v_11434;
wire v_11435;
wire v_11436;
wire v_11437;
wire v_11438;
wire v_11439;
wire v_11440;
wire v_11441;
wire v_11442;
wire v_11443;
wire v_11444;
wire v_11445;
wire v_11446;
wire v_11447;
wire v_11448;
wire v_11449;
wire v_11450;
wire v_11451;
wire v_11452;
wire v_11453;
wire v_11454;
wire v_11455;
wire v_11456;
wire v_11457;
wire v_11458;
wire v_11459;
wire v_11460;
wire v_11461;
wire v_11462;
wire v_11463;
wire v_11464;
wire v_11465;
wire v_11466;
wire v_11467;
wire v_11468;
wire v_11469;
wire v_11470;
wire v_11471;
wire v_11472;
wire v_11473;
wire v_11474;
wire v_11475;
wire v_11476;
wire v_11477;
wire v_11478;
wire v_11479;
wire v_11480;
wire v_11481;
wire v_11482;
wire v_11483;
wire v_11484;
wire v_11485;
wire v_11486;
wire v_11487;
wire v_11488;
wire v_11489;
wire v_11490;
wire v_11491;
wire v_11492;
wire v_11493;
wire v_11494;
wire v_11495;
wire v_11496;
wire v_11497;
wire v_11498;
wire v_11499;
wire v_11500;
wire v_11502;
wire v_11503;
wire v_11504;
wire v_11505;
wire v_11506;
wire v_11507;
wire v_11508;
wire v_11509;
wire v_11510;
wire v_11511;
wire v_11512;
wire v_11513;
wire v_11514;
wire v_11515;
wire v_11516;
wire v_11517;
wire v_11518;
wire v_11519;
wire v_11520;
wire v_11521;
wire v_11522;
wire v_11523;
wire v_11524;
wire v_11525;
wire v_11526;
wire v_11527;
wire v_11528;
wire v_11529;
wire v_11530;
wire v_11531;
wire v_11532;
wire v_11533;
wire v_11534;
wire v_11535;
wire v_11536;
wire v_11537;
wire v_11538;
wire v_11539;
wire v_11540;
wire v_11541;
wire v_11542;
wire v_11543;
wire v_11544;
wire v_11545;
wire v_11546;
wire v_11547;
wire v_11548;
wire v_11549;
wire v_11550;
wire v_11551;
wire v_11552;
wire v_11553;
wire v_11554;
wire v_11555;
wire v_11556;
wire v_11557;
wire v_11558;
wire v_11559;
wire v_11560;
wire v_11561;
wire v_11562;
wire v_11563;
wire v_11564;
wire v_11565;
wire v_11566;
wire v_11567;
wire v_11568;
wire v_11569;
wire v_11570;
wire v_11571;
wire v_11572;
wire v_11573;
wire v_11574;
wire v_11575;
wire v_11576;
wire v_11577;
wire v_11578;
wire v_11579;
wire v_11580;
wire v_11581;
wire v_11582;
wire v_11583;
wire v_11584;
wire v_11585;
wire v_11586;
wire v_11587;
wire v_11588;
wire v_11589;
wire v_11590;
wire v_11591;
wire v_11592;
wire v_11593;
wire v_11594;
wire v_11595;
wire v_11596;
wire v_11597;
wire v_11598;
wire v_11599;
wire v_11600;
wire v_11601;
wire v_11602;
wire v_11603;
wire v_11604;
wire v_11605;
wire v_11606;
wire v_11607;
wire v_11608;
wire v_11609;
wire v_11610;
wire v_11611;
wire v_11612;
wire v_11613;
wire v_11614;
wire v_11615;
wire v_11616;
wire v_11617;
wire v_11618;
wire v_11619;
wire v_11620;
wire v_11621;
wire v_11622;
wire v_11623;
wire v_11624;
wire v_11625;
wire v_11627;
wire v_11628;
wire v_11629;
wire v_11630;
wire v_11631;
wire v_11632;
wire v_11633;
wire v_11634;
wire v_11635;
wire v_11636;
wire v_11637;
wire v_11638;
wire v_11639;
wire v_11640;
wire v_11641;
wire v_11642;
wire v_11643;
wire v_11644;
wire v_11645;
wire v_11647;
wire v_11648;
wire v_11649;
wire v_11650;
wire v_11651;
wire v_11652;
wire v_11653;
wire v_11654;
wire v_11655;
wire v_11656;
wire v_11657;
wire v_11658;
wire v_11659;
wire v_11660;
wire v_11661;
wire v_11662;
wire v_11663;
wire v_11664;
wire v_11665;
wire v_11666;
wire v_11667;
wire v_11668;
wire v_11669;
wire v_11670;
wire v_11671;
wire v_11672;
wire v_11673;
wire v_11674;
wire v_11675;
wire v_11676;
wire v_11677;
wire v_11678;
wire v_11679;
wire v_11680;
wire v_11681;
wire v_11682;
wire v_11683;
wire v_11684;
wire v_11685;
wire v_11686;
wire v_11687;
wire v_11688;
wire v_11689;
wire v_11690;
wire v_11691;
wire v_11692;
wire v_11693;
wire v_11694;
wire v_11695;
wire v_11696;
wire v_11698;
wire v_11699;
wire v_11700;
wire v_11701;
wire v_11702;
wire v_11703;
wire v_11704;
wire v_11705;
wire v_11706;
wire v_11707;
wire v_11708;
wire v_11709;
wire v_11710;
wire v_11711;
wire v_11712;
wire v_11713;
wire v_11714;
wire v_11716;
wire v_11717;
wire v_11718;
wire v_11719;
wire v_11720;
wire v_11721;
wire v_11722;
wire v_11723;
wire v_11724;
wire v_11725;
wire v_11726;
wire v_11727;
wire v_11728;
wire v_11729;
wire v_11730;
wire v_11731;
wire v_11732;
wire v_11733;
wire v_11734;
wire v_11735;
wire v_11736;
wire v_11737;
wire v_11738;
wire v_11739;
wire v_11740;
wire v_11741;
wire v_11742;
wire v_11743;
wire v_11744;
wire v_11745;
wire v_11746;
wire v_11747;
wire v_11748;
wire v_11749;
wire v_11750;
wire v_11751;
wire v_11752;
wire v_11753;
wire v_11754;
wire v_11755;
wire v_11756;
wire v_11757;
wire v_11758;
wire v_11759;
wire v_11760;
wire v_11761;
wire v_11762;
wire v_11763;
wire v_11764;
wire v_11765;
wire v_11766;
wire v_11767;
wire v_11768;
wire v_11769;
wire v_11770;
wire v_11771;
wire v_11772;
wire v_11773;
wire v_11774;
wire v_11775;
wire v_11776;
wire v_11777;
wire v_11778;
wire v_11779;
wire v_11780;
wire v_11781;
wire v_11782;
wire v_11783;
wire v_11784;
wire v_11785;
wire v_11786;
wire v_11787;
wire v_11788;
wire v_11789;
wire v_11790;
wire v_11791;
wire v_11792;
wire v_11793;
wire v_11794;
wire v_11795;
wire v_11796;
wire v_11797;
wire v_11798;
wire v_11799;
wire v_11800;
wire v_11801;
wire v_11802;
wire v_11803;
wire v_11804;
wire v_11805;
wire v_11806;
wire v_11807;
wire v_11808;
wire v_11809;
wire v_11810;
wire v_11811;
wire v_11812;
wire v_11813;
wire v_11814;
wire v_11815;
wire v_11816;
wire v_11817;
wire v_11818;
wire v_11819;
wire v_11820;
wire v_11821;
wire v_11822;
wire v_11823;
wire v_11824;
wire v_11825;
wire v_11826;
wire v_11827;
wire v_11828;
wire v_11829;
wire v_11830;
wire v_11831;
wire v_11832;
wire v_11833;
wire v_11834;
wire v_11835;
wire v_11836;
wire v_11837;
wire v_11838;
wire v_11839;
wire v_11840;
wire v_11841;
wire v_11842;
wire v_11843;
wire v_11844;
wire v_11845;
wire v_11846;
wire v_11847;
wire v_11848;
wire v_11849;
wire v_11850;
wire v_11851;
wire v_11852;
wire v_11853;
wire v_11854;
wire v_11855;
wire v_11856;
wire v_11857;
wire v_11858;
wire v_11859;
wire v_11860;
wire v_11861;
wire v_11862;
wire v_11863;
wire v_11864;
wire v_11865;
wire v_11866;
wire v_11867;
wire v_11868;
wire v_11869;
wire v_11870;
wire v_11871;
wire v_11872;
wire v_11873;
wire v_11874;
wire v_11875;
wire v_11876;
wire v_11877;
wire v_11878;
wire v_11879;
wire v_11880;
wire v_11881;
wire v_11882;
wire v_11883;
wire v_11884;
wire v_11885;
wire v_11886;
wire v_11887;
wire v_11888;
wire v_11889;
wire v_11890;
wire v_11891;
wire v_11892;
wire v_11893;
wire v_11894;
wire v_11895;
wire v_11896;
wire v_11897;
wire v_11898;
wire v_11899;
wire v_11900;
wire v_11901;
wire v_11902;
wire v_11903;
wire v_11904;
wire v_11905;
wire v_11906;
wire v_11907;
wire v_11908;
wire v_11909;
wire v_11910;
wire v_11911;
wire v_11912;
wire v_11913;
wire v_11914;
wire v_11915;
wire v_11916;
wire v_11917;
wire v_11918;
wire v_11919;
wire v_11920;
wire v_11921;
wire v_11922;
wire v_11923;
wire v_11924;
wire v_11925;
wire v_11926;
wire v_11927;
wire v_11928;
wire v_11929;
wire v_11930;
wire v_11931;
wire v_11932;
wire v_11933;
wire v_11934;
wire v_11935;
wire v_11936;
wire v_11937;
wire v_11938;
wire v_11939;
wire v_11940;
wire v_11941;
wire v_11942;
wire v_11943;
wire v_11944;
wire v_11945;
wire v_11946;
wire v_11947;
wire v_11948;
wire v_11949;
wire v_11950;
wire v_11951;
wire v_11952;
wire v_11953;
wire v_11954;
wire v_11955;
wire v_11956;
wire v_11957;
wire v_11958;
wire v_11959;
wire v_11960;
wire v_11961;
wire v_11962;
wire v_11963;
wire v_11964;
wire v_11965;
wire v_11966;
wire v_11968;
wire v_11969;
wire v_11970;
wire v_11971;
wire v_11973;
wire v_11974;
wire v_11975;
wire v_11976;
wire v_11977;
wire v_11978;
wire v_11979;
wire v_11980;
wire v_11981;
wire v_11982;
wire v_11983;
wire v_11984;
wire v_11985;
wire v_11986;
wire v_11987;
wire v_11988;
wire v_11989;
wire v_11990;
wire v_11991;
wire v_11992;
wire v_11993;
wire v_11994;
wire v_11995;
wire v_11996;
wire v_11997;
wire v_11998;
wire v_11999;
wire v_12000;
wire v_12001;
wire v_12002;
wire v_12003;
wire v_12004;
wire v_12005;
wire v_12006;
wire v_12007;
wire v_12008;
wire v_12009;
wire v_12010;
wire v_12011;
wire v_12012;
wire v_12013;
wire v_12014;
wire v_12015;
wire v_12016;
wire v_12017;
wire v_12018;
wire v_12019;
wire v_12020;
wire v_12021;
wire v_12022;
wire v_12023;
wire v_12024;
wire v_12025;
wire v_12026;
wire v_12027;
wire v_12028;
wire v_12029;
wire v_12030;
wire v_12031;
wire v_12032;
wire v_12033;
wire v_12034;
wire v_12035;
wire v_12036;
wire v_12037;
wire v_12038;
wire v_12039;
wire v_12040;
wire v_12041;
wire v_12042;
wire v_12043;
wire v_12044;
wire v_12045;
wire v_12046;
wire v_12047;
wire v_12048;
wire v_12049;
wire v_12050;
wire v_12051;
wire v_12052;
wire v_12053;
wire v_12054;
wire v_12055;
wire v_12056;
wire v_12057;
wire v_12058;
wire v_12059;
wire v_12060;
wire v_12061;
wire v_12062;
wire v_12063;
wire v_12064;
wire v_12065;
wire v_12066;
wire v_12068;
wire v_12069;
wire v_12070;
wire v_12071;
wire v_12072;
wire v_12073;
wire v_12074;
wire v_12075;
wire v_12076;
wire v_12077;
wire v_12078;
wire v_12079;
wire v_12080;
wire v_12081;
wire v_12082;
wire v_12083;
wire v_12084;
wire v_12085;
wire v_12086;
wire v_12087;
wire v_12088;
wire v_12089;
wire v_12090;
wire v_12091;
wire v_12092;
wire v_12093;
wire v_12094;
wire v_12095;
wire v_12096;
wire v_12097;
wire v_12098;
wire v_12099;
wire v_12100;
wire v_12101;
wire v_12102;
wire v_12103;
wire v_12104;
wire v_12105;
wire v_12106;
wire v_12107;
wire v_12108;
wire v_12109;
wire v_12110;
wire v_12111;
wire v_12112;
wire v_12113;
wire v_12114;
wire v_12115;
wire v_12116;
wire v_12117;
wire v_12118;
wire v_12119;
wire v_12120;
wire v_12121;
wire v_12122;
wire v_12123;
wire v_12124;
wire v_12125;
wire v_12126;
wire v_12127;
wire v_12128;
wire v_12129;
wire v_12130;
wire v_12131;
wire v_12132;
wire v_12133;
wire v_12134;
wire v_12135;
wire v_12136;
wire v_12137;
wire v_12138;
wire v_12139;
wire v_12140;
wire v_12141;
wire v_12142;
wire v_12143;
wire v_12144;
wire v_12145;
wire v_12146;
wire v_12147;
wire v_12148;
wire v_12149;
wire v_12150;
wire v_12151;
wire v_12152;
wire v_12153;
wire v_12154;
wire v_12155;
wire v_12156;
wire v_12157;
wire v_12158;
wire v_12159;
wire v_12160;
wire v_12161;
wire v_12162;
wire v_12163;
wire v_12164;
wire v_12165;
wire v_12166;
wire v_12167;
wire v_12168;
wire v_12169;
wire v_12170;
wire v_12171;
wire v_12172;
wire v_12173;
wire v_12174;
wire v_12175;
wire v_12176;
wire v_12177;
wire v_12178;
wire v_12179;
wire v_12180;
wire v_12181;
wire v_12182;
wire v_12183;
wire v_12184;
wire v_12185;
wire v_12186;
wire v_12187;
wire v_12188;
wire v_12189;
wire v_12190;
wire v_12191;
wire v_12192;
wire v_12193;
wire v_12194;
wire v_12195;
wire v_12196;
wire v_12197;
wire v_12198;
wire v_12199;
wire v_12200;
wire v_12201;
wire v_12202;
wire v_12203;
wire v_12204;
wire v_12205;
wire v_12206;
wire v_12207;
wire v_12208;
wire v_12209;
wire v_12210;
wire v_12211;
wire v_12212;
wire v_12213;
wire v_12214;
wire v_12215;
wire v_12216;
wire v_12217;
wire v_12218;
wire v_12219;
wire v_12220;
wire v_12221;
wire v_12222;
wire v_12223;
wire v_12224;
wire v_12225;
wire v_12226;
wire v_12227;
wire v_12228;
wire v_12229;
wire v_12230;
wire v_12231;
wire v_12232;
wire v_12233;
wire v_12234;
wire v_12235;
wire v_12236;
wire v_12237;
wire v_12238;
wire v_12239;
wire v_12240;
wire v_12241;
wire v_12242;
wire v_12243;
wire v_12244;
wire v_12245;
wire v_12246;
wire v_12247;
wire v_12248;
wire v_12249;
wire v_12250;
wire v_12251;
wire v_12252;
wire v_12253;
wire v_12254;
wire v_12255;
wire v_12256;
wire v_12257;
wire v_12258;
wire v_12259;
wire v_12260;
wire v_12261;
wire v_12262;
wire v_12263;
wire v_12264;
wire v_12265;
wire v_12266;
wire v_12267;
wire v_12268;
wire v_12269;
wire v_12270;
wire v_12271;
wire v_12272;
wire v_12273;
wire v_12274;
wire v_12275;
wire v_12276;
wire v_12277;
wire v_12278;
wire v_12279;
wire v_12280;
wire v_12281;
wire v_12282;
wire v_12283;
wire v_12284;
wire v_12285;
wire v_12286;
wire v_12287;
wire v_12288;
wire v_12289;
wire v_12290;
wire v_12291;
wire v_12292;
wire v_12293;
wire v_12294;
wire v_12295;
wire v_12296;
wire v_12297;
wire v_12298;
wire v_12299;
wire v_12300;
wire v_12301;
wire v_12302;
wire v_12303;
wire v_12304;
wire v_12305;
wire v_12306;
wire v_12307;
wire v_12308;
wire v_12309;
wire v_12310;
wire v_12311;
wire v_12312;
wire v_12313;
wire v_12314;
wire v_12315;
wire v_12316;
wire v_12317;
wire v_12318;
wire v_12319;
wire v_12320;
wire v_12321;
wire v_12322;
wire v_12323;
wire v_12324;
wire v_12325;
wire v_12326;
wire v_12327;
wire v_12328;
wire v_12329;
wire v_12330;
wire v_12331;
wire v_12332;
wire v_12333;
wire v_12334;
wire v_12335;
wire v_12336;
wire v_12337;
wire v_12338;
wire v_12339;
wire v_12340;
wire v_12341;
wire v_12342;
wire v_12343;
wire v_12344;
wire v_12345;
wire v_12346;
wire v_12347;
wire v_12348;
wire v_12349;
wire v_12350;
wire v_12351;
wire v_12352;
wire v_12353;
wire v_12354;
wire v_12355;
wire v_12356;
wire v_12357;
wire v_12358;
wire v_12359;
wire v_12360;
wire v_12361;
wire v_12362;
wire v_12363;
wire v_12364;
wire v_12365;
wire v_12366;
wire v_12367;
wire v_12368;
wire v_12369;
wire v_12370;
wire v_12371;
wire v_12372;
wire v_12373;
wire v_12374;
wire v_12375;
wire v_12376;
wire v_12377;
wire v_12378;
wire v_12379;
wire v_12380;
wire v_12381;
wire v_12382;
wire v_12383;
wire v_12384;
wire v_12385;
wire v_12386;
wire v_12387;
wire v_12388;
wire v_12389;
wire v_12390;
wire v_12391;
wire v_12392;
wire v_12393;
wire v_12394;
wire v_12395;
wire v_12396;
wire v_12397;
wire v_12399;
wire v_12400;
wire v_12401;
wire v_12402;
wire v_12403;
wire v_12404;
wire v_12405;
wire v_12406;
wire v_12407;
wire v_12408;
wire v_12409;
wire v_12410;
wire v_12411;
wire v_12412;
wire v_12413;
wire v_12414;
wire v_12415;
wire v_12416;
wire v_12417;
wire v_12418;
wire v_12419;
wire v_12420;
wire v_12421;
wire v_12422;
wire v_12423;
wire v_12424;
wire v_12425;
wire v_12426;
wire v_12427;
wire v_12428;
wire v_12429;
wire v_12430;
wire v_12431;
wire v_12432;
wire v_12433;
wire v_12434;
wire v_12435;
wire v_12436;
wire v_12437;
wire v_12438;
wire v_12439;
wire v_12440;
wire v_12441;
wire v_12442;
wire v_12443;
wire v_12444;
wire v_12445;
wire v_12446;
wire v_12447;
wire v_12448;
wire v_12449;
wire v_12450;
wire v_12451;
wire v_12452;
wire v_12453;
wire v_12454;
wire v_12455;
wire v_12456;
wire v_12457;
wire v_12458;
wire v_12459;
wire v_12460;
wire v_12461;
wire v_12462;
wire v_12463;
wire v_12464;
wire v_12465;
wire v_12466;
wire v_12467;
wire v_12468;
wire v_12469;
wire v_12470;
wire v_12471;
wire v_12472;
wire v_12473;
wire v_12474;
wire v_12475;
wire v_12476;
wire v_12477;
wire v_12478;
wire v_12479;
wire v_12480;
wire v_12481;
wire v_12482;
wire v_12483;
wire v_12484;
wire v_12485;
wire v_12486;
wire v_12487;
wire v_12488;
wire v_12489;
wire v_12490;
wire v_12491;
wire v_12492;
wire v_12493;
wire v_12494;
wire v_12495;
wire v_12496;
wire v_12497;
wire v_12498;
wire v_12499;
wire v_12500;
wire v_12501;
wire v_12502;
wire v_12503;
wire v_12504;
wire v_12505;
wire v_12506;
wire v_12507;
wire v_12508;
wire v_12509;
wire v_12510;
wire v_12511;
wire v_12512;
wire v_12513;
wire v_12514;
wire v_12515;
wire v_12516;
wire v_12517;
wire v_12518;
wire v_12519;
wire v_12520;
wire v_12521;
wire v_12522;
wire v_12524;
wire v_12525;
wire v_12526;
wire v_12527;
wire v_12528;
wire v_12529;
wire v_12530;
wire v_12531;
wire v_12532;
wire v_12533;
wire v_12534;
wire v_12535;
wire v_12536;
wire v_12537;
wire v_12538;
wire v_12539;
wire v_12540;
wire v_12541;
wire v_12542;
wire v_12544;
wire v_12545;
wire v_12546;
wire v_12547;
wire v_12548;
wire v_12549;
wire v_12550;
wire v_12551;
wire v_12552;
wire v_12553;
wire v_12554;
wire v_12555;
wire v_12556;
wire v_12557;
wire v_12558;
wire v_12559;
wire v_12560;
wire v_12561;
wire v_12562;
wire v_12563;
wire v_12564;
wire v_12565;
wire v_12566;
wire v_12567;
wire v_12568;
wire v_12569;
wire v_12570;
wire v_12571;
wire v_12572;
wire v_12573;
wire v_12574;
wire v_12575;
wire v_12576;
wire v_12577;
wire v_12578;
wire v_12579;
wire v_12580;
wire v_12581;
wire v_12582;
wire v_12583;
wire v_12584;
wire v_12585;
wire v_12586;
wire v_12587;
wire v_12588;
wire v_12589;
wire v_12590;
wire v_12591;
wire v_12592;
wire v_12593;
wire v_12595;
wire v_12596;
wire v_12597;
wire v_12598;
wire v_12599;
wire v_12600;
wire v_12601;
wire v_12602;
wire v_12603;
wire v_12604;
wire v_12605;
wire v_12606;
wire v_12607;
wire v_12608;
wire v_12609;
wire v_12610;
wire v_12611;
wire v_12613;
wire v_12614;
wire v_12615;
wire v_12616;
wire v_12617;
wire v_12618;
wire v_12619;
wire v_12620;
wire v_12621;
wire v_12622;
wire v_12623;
wire v_12624;
wire v_12625;
wire v_12626;
wire v_12627;
wire v_12628;
wire v_12629;
wire v_12630;
wire v_12631;
wire v_12632;
wire v_12633;
wire v_12634;
wire v_12635;
wire v_12636;
wire v_12637;
wire v_12638;
wire v_12639;
wire v_12640;
wire v_12641;
wire v_12642;
wire v_12643;
wire v_12644;
wire v_12645;
wire v_12646;
wire v_12647;
wire v_12648;
wire v_12649;
wire v_12650;
wire v_12651;
wire v_12652;
wire v_12653;
wire v_12654;
wire v_12655;
wire v_12656;
wire v_12657;
wire v_12658;
wire v_12659;
wire v_12660;
wire v_12661;
wire v_12662;
wire v_12663;
wire v_12664;
wire v_12665;
wire v_12666;
wire v_12667;
wire v_12668;
wire v_12669;
wire v_12670;
wire v_12671;
wire v_12672;
wire v_12673;
wire v_12674;
wire v_12675;
wire v_12676;
wire v_12677;
wire v_12678;
wire v_12679;
wire v_12680;
wire v_12681;
wire v_12682;
wire v_12683;
wire v_12684;
wire v_12685;
wire v_12686;
wire v_12687;
wire v_12688;
wire v_12689;
wire v_12690;
wire v_12691;
wire v_12692;
wire v_12693;
wire v_12694;
wire v_12695;
wire v_12696;
wire v_12697;
wire v_12698;
wire v_12699;
wire v_12700;
wire v_12701;
wire v_12702;
wire v_12703;
wire v_12704;
wire v_12705;
wire v_12706;
wire v_12707;
wire v_12708;
wire v_12709;
wire v_12710;
wire v_12711;
wire v_12712;
wire v_12713;
wire v_12714;
wire v_12715;
wire v_12716;
wire v_12717;
wire v_12718;
wire v_12719;
wire v_12720;
wire v_12721;
wire v_12722;
wire v_12723;
wire v_12724;
wire v_12725;
wire v_12726;
wire v_12727;
wire v_12728;
wire v_12729;
wire v_12730;
wire v_12731;
wire v_12732;
wire v_12733;
wire v_12734;
wire v_12735;
wire v_12736;
wire v_12737;
wire v_12738;
wire v_12739;
wire v_12740;
wire v_12741;
wire v_12742;
wire v_12743;
wire v_12744;
wire v_12745;
wire v_12746;
wire v_12747;
wire v_12748;
wire v_12749;
wire v_12750;
wire v_12751;
wire v_12752;
wire v_12753;
wire v_12754;
wire v_12755;
wire v_12756;
wire v_12757;
wire v_12758;
wire v_12759;
wire v_12760;
wire v_12761;
wire v_12762;
wire v_12763;
wire v_12764;
wire v_12765;
wire v_12766;
wire v_12767;
wire v_12768;
wire v_12769;
wire v_12770;
wire v_12771;
wire v_12772;
wire v_12773;
wire v_12774;
wire v_12775;
wire v_12776;
wire v_12777;
wire v_12778;
wire v_12779;
wire v_12780;
wire v_12781;
wire v_12782;
wire v_12783;
wire v_12784;
wire v_12785;
wire v_12786;
wire v_12787;
wire v_12788;
wire v_12789;
wire v_12790;
wire v_12791;
wire v_12792;
wire v_12793;
wire v_12794;
wire v_12795;
wire v_12796;
wire v_12797;
wire v_12798;
wire v_12799;
wire v_12800;
wire v_12801;
wire v_12802;
wire v_12803;
wire v_12804;
wire v_12805;
wire v_12806;
wire v_12807;
wire v_12808;
wire v_12809;
wire v_12810;
wire v_12811;
wire v_12812;
wire v_12813;
wire v_12814;
wire v_12815;
wire v_12816;
wire v_12817;
wire v_12818;
wire v_12819;
wire v_12820;
wire v_12821;
wire v_12822;
wire v_12823;
wire v_12824;
wire v_12825;
wire v_12826;
wire v_12827;
wire v_12828;
wire v_12829;
wire v_12830;
wire v_12831;
wire v_12832;
wire v_12833;
wire v_12834;
wire v_12835;
wire v_12836;
wire v_12837;
wire v_12838;
wire v_12839;
wire v_12840;
wire v_12841;
wire v_12842;
wire v_12843;
wire v_12844;
wire v_12845;
wire v_12846;
wire v_12847;
wire v_12848;
wire v_12849;
wire v_12850;
wire v_12851;
wire v_12852;
wire v_12853;
wire v_12854;
wire v_12855;
wire v_12856;
wire v_12857;
wire v_12858;
wire v_12859;
wire v_12860;
wire v_12861;
wire v_12862;
wire v_12863;
wire v_12864;
wire v_12865;
wire v_12866;
wire v_12867;
wire v_12868;
wire v_12869;
wire v_12870;
wire v_12871;
wire v_12872;
wire v_12873;
wire v_12874;
wire v_12875;
wire v_12876;
wire v_12877;
wire v_12878;
wire v_12879;
wire v_12880;
wire v_12881;
wire v_12882;
wire v_12883;
wire v_12884;
wire v_12885;
wire v_12886;
wire v_12887;
wire v_12888;
wire v_12889;
wire v_12890;
wire v_12891;
wire v_12892;
wire v_12893;
wire v_12894;
wire v_12895;
wire v_12896;
wire v_12897;
wire v_12898;
wire v_12899;
wire v_12900;
wire v_12901;
wire v_12902;
wire v_12903;
wire v_12904;
wire v_12905;
wire v_12906;
wire v_12907;
wire v_12908;
wire v_12909;
wire v_12910;
wire v_12911;
wire v_12912;
wire v_12913;
wire v_12914;
wire v_12915;
wire v_12916;
wire v_12917;
wire v_12918;
wire v_12919;
wire v_12920;
wire v_12921;
wire v_12922;
wire v_12923;
wire v_12924;
wire v_12925;
wire v_12926;
wire v_12927;
wire v_12928;
wire v_12929;
wire v_12930;
wire v_12931;
wire v_12932;
wire v_12933;
wire v_12934;
wire v_12935;
wire v_12936;
wire v_12937;
wire v_12938;
wire v_12939;
wire v_12940;
wire v_12941;
wire v_12942;
wire v_12943;
wire v_12944;
wire v_12945;
wire v_12946;
wire v_12947;
wire v_12948;
wire v_12949;
wire v_12950;
wire v_12951;
wire v_12952;
wire v_12953;
wire v_12954;
wire v_12955;
wire v_12956;
wire v_12957;
wire v_12958;
wire v_12959;
wire v_12960;
wire v_12961;
wire v_12962;
wire v_12963;
wire v_12964;
wire v_12965;
wire v_12966;
wire v_12967;
wire v_12968;
wire v_12969;
wire v_12970;
wire v_12971;
wire v_12972;
wire v_12973;
wire v_12974;
wire v_12975;
wire v_12976;
wire v_12977;
wire v_12978;
wire v_12979;
wire v_12980;
wire v_12981;
wire v_12982;
wire v_12983;
wire v_12984;
wire v_12985;
wire v_12986;
wire v_12987;
wire v_12988;
wire v_12989;
wire v_12990;
wire v_12991;
wire v_12992;
wire v_12993;
wire v_12994;
wire v_12995;
wire v_12996;
wire v_12997;
wire v_12998;
wire v_12999;
wire v_13000;
wire v_13001;
wire v_13002;
wire v_13003;
wire v_13004;
wire v_13005;
wire v_13006;
wire v_13007;
wire v_13008;
wire v_13009;
wire v_13010;
wire v_13011;
wire v_13012;
wire v_13013;
wire v_13014;
wire v_13015;
wire v_13016;
wire v_13017;
wire v_13018;
wire v_13019;
wire v_13020;
wire v_13021;
wire v_13022;
wire v_13023;
wire v_13024;
wire v_13025;
wire v_13026;
wire v_13027;
wire v_13028;
wire v_13029;
wire v_13030;
wire v_13031;
wire v_13032;
wire v_13033;
wire v_13034;
wire v_13035;
wire v_13036;
wire v_13037;
wire v_13038;
wire v_13039;
wire v_13040;
wire v_13041;
wire v_13042;
wire v_13043;
wire v_13044;
wire v_13045;
wire v_13046;
wire v_13047;
wire v_13048;
wire v_13049;
wire v_13050;
wire v_13051;
wire v_13052;
wire v_13053;
wire v_13054;
wire v_13055;
wire v_13056;
wire v_13057;
wire v_13058;
wire v_13059;
wire v_13060;
wire v_13061;
wire v_13062;
wire v_13063;
wire v_13064;
wire v_13065;
wire v_13066;
wire v_13067;
wire v_13068;
wire v_13069;
wire v_13070;
wire v_13071;
wire v_13072;
wire v_13073;
wire v_13074;
wire v_13075;
wire v_13076;
wire v_13077;
wire v_13078;
wire v_13079;
wire v_13080;
wire v_13081;
wire v_13082;
wire v_13083;
wire v_13084;
wire v_13085;
wire v_13086;
wire v_13087;
wire v_13088;
wire v_13089;
wire v_13090;
wire v_13091;
wire v_13092;
wire v_13093;
wire v_13094;
wire v_13095;
wire v_13096;
wire v_13097;
wire v_13098;
wire v_13099;
wire v_13100;
wire v_13101;
wire v_13102;
wire v_13103;
wire v_13104;
wire v_13105;
wire v_13106;
wire v_13107;
wire v_13108;
wire v_13109;
wire v_13110;
wire v_13111;
wire v_13112;
wire v_13113;
wire v_13114;
wire v_13115;
wire v_13116;
wire v_13117;
wire v_13118;
wire v_13119;
wire v_13120;
wire v_13121;
wire v_13122;
wire v_13123;
wire v_13124;
wire v_13125;
wire v_13126;
wire v_13127;
wire v_13128;
wire v_13129;
wire v_13130;
wire v_13131;
wire v_13132;
wire v_13133;
wire v_13134;
wire v_13135;
wire v_13136;
wire v_13137;
wire v_13138;
wire v_13139;
wire v_13140;
wire v_13141;
wire v_13142;
wire v_13143;
wire v_13144;
wire v_13145;
wire v_13146;
wire v_13147;
wire v_13148;
wire v_13149;
wire v_13150;
wire v_13151;
wire v_13152;
wire v_13153;
wire v_13154;
wire v_13155;
wire v_13156;
wire v_13157;
wire v_13158;
wire v_13159;
wire v_13160;
wire v_13161;
wire v_13162;
wire v_13163;
wire v_13164;
wire v_13165;
wire v_13166;
wire v_13167;
wire v_13168;
wire v_13169;
wire v_13170;
wire v_13171;
wire v_13172;
wire v_13173;
wire v_13174;
wire v_13175;
wire v_13176;
wire v_13177;
wire v_13178;
wire v_13179;
wire v_13180;
wire v_13181;
wire v_13182;
wire v_13183;
wire v_13184;
wire v_13185;
wire v_13186;
wire v_13187;
wire v_13188;
wire v_13189;
wire v_13190;
wire v_13191;
wire v_13192;
wire v_13193;
wire v_13194;
wire v_13195;
wire v_13196;
wire v_13197;
wire v_13198;
wire v_13199;
wire v_13200;
wire v_13201;
wire v_13202;
wire v_13203;
wire v_13204;
wire v_13205;
wire v_13206;
wire v_13207;
wire v_13208;
wire v_13209;
wire v_13210;
wire v_13211;
wire v_13212;
wire v_13213;
wire v_13214;
wire v_13215;
wire v_13216;
wire v_13217;
wire v_13218;
wire v_13219;
wire v_13220;
wire v_13221;
wire v_13222;
wire v_13223;
wire v_13224;
wire v_13225;
wire v_13226;
wire v_13227;
wire v_13228;
wire v_13229;
wire v_13230;
wire v_13231;
wire v_13232;
wire v_13233;
wire v_13234;
wire v_13235;
wire v_13236;
wire v_13237;
wire v_13238;
wire v_13239;
wire v_13240;
wire v_13241;
wire v_13242;
wire v_13243;
wire v_13244;
wire v_13245;
wire v_13246;
wire v_13247;
wire v_13248;
wire v_13249;
wire v_13250;
wire v_13251;
wire v_13252;
wire v_13253;
wire v_13254;
wire v_13255;
wire v_13256;
wire v_13257;
wire v_13258;
wire v_13259;
wire v_13260;
wire v_13261;
wire v_13262;
wire v_13263;
wire v_13264;
wire v_13265;
wire v_13266;
wire v_13267;
wire v_13268;
wire v_13269;
wire v_13270;
wire v_13271;
wire v_13272;
wire v_13273;
wire v_13274;
wire v_13275;
wire v_13276;
wire v_13277;
wire v_13278;
wire v_13279;
wire v_13280;
wire v_13281;
wire v_13282;
wire v_13283;
wire v_13284;
wire v_13285;
wire v_13286;
wire v_13287;
wire v_13288;
wire v_13289;
wire v_13290;
wire v_13291;
wire v_13292;
wire v_13293;
wire v_13294;
wire v_13295;
wire v_13296;
wire v_13297;
wire v_13298;
wire v_13299;
wire v_13300;
wire v_13301;
wire v_13302;
wire v_13303;
wire v_13304;
wire v_13305;
wire v_13306;
wire v_13307;
wire v_13308;
wire v_13309;
wire v_13310;
wire v_13311;
wire v_13312;
wire v_13313;
wire v_13314;
wire v_13315;
wire v_13316;
wire v_13317;
wire v_13318;
wire v_13319;
wire v_13320;
wire v_13321;
wire v_13322;
wire v_13323;
wire v_13324;
wire v_13325;
wire v_13326;
wire v_13327;
wire v_13328;
wire v_13329;
wire v_13330;
wire v_13331;
wire v_13332;
wire v_13333;
wire v_13334;
wire v_13335;
wire v_13336;
wire v_13337;
wire v_13338;
wire v_13339;
wire v_13340;
wire v_13341;
wire v_13342;
wire v_13343;
wire v_13344;
wire v_13345;
wire v_13346;
wire v_13347;
wire v_13348;
wire v_13349;
wire v_13350;
wire v_13351;
wire v_13352;
wire v_13353;
wire v_13354;
wire v_13355;
wire v_13356;
wire v_13357;
wire v_13358;
wire v_13359;
wire v_13360;
wire v_13361;
wire v_13362;
wire v_13363;
wire v_13364;
wire v_13365;
wire v_13366;
wire v_13367;
wire v_13368;
wire v_13369;
wire v_13370;
wire v_13371;
wire v_13372;
wire v_13373;
wire v_13374;
wire v_13375;
wire v_13376;
wire v_13377;
wire v_13378;
wire v_13379;
wire v_13380;
wire v_13381;
wire v_13382;
wire v_13383;
wire v_13384;
wire v_13385;
wire v_13386;
wire v_13387;
wire v_13388;
wire v_13389;
wire v_13390;
wire v_13391;
wire v_13392;
wire v_13393;
wire v_13394;
wire v_13395;
wire v_13396;
wire v_13397;
wire v_13398;
wire v_13399;
wire v_13400;
wire v_13401;
wire v_13402;
wire v_13403;
wire v_13404;
wire v_13405;
wire v_13406;
wire v_13407;
wire v_13408;
wire v_13409;
wire v_13410;
wire v_13411;
wire v_13412;
wire v_13413;
wire v_13414;
wire v_13415;
wire v_13416;
wire v_13417;
wire v_13418;
wire v_13419;
wire v_13420;
wire v_13421;
wire v_13422;
wire v_13423;
wire v_13424;
wire v_13425;
wire v_13426;
wire v_13427;
wire v_13428;
wire v_13429;
wire v_13430;
wire v_13431;
wire v_13432;
wire v_13433;
wire v_13434;
wire v_13435;
wire v_13436;
wire v_13437;
wire v_13438;
wire v_13439;
wire v_13440;
wire v_13441;
wire v_13442;
wire v_13443;
wire v_13444;
wire v_13445;
wire v_13446;
wire v_13447;
wire v_13448;
wire v_13449;
wire v_13450;
wire v_13451;
wire v_13452;
wire v_13453;
wire v_13454;
wire v_13455;
wire v_13456;
wire v_13457;
wire v_13458;
wire v_13459;
wire v_13460;
wire v_13461;
wire v_13462;
wire v_13463;
wire v_13464;
wire v_13465;
wire v_13466;
wire v_13467;
wire v_13468;
wire v_13469;
wire v_13470;
wire v_13471;
wire v_13472;
wire v_13473;
wire v_13474;
wire v_13475;
wire v_13476;
wire v_13477;
wire v_13478;
wire v_13479;
wire v_13480;
wire v_13481;
wire v_13482;
wire v_13483;
wire v_13484;
wire v_13485;
wire v_13486;
wire v_13487;
wire v_13488;
wire v_13489;
wire v_13490;
wire v_13491;
wire v_13492;
wire v_13493;
wire v_13494;
wire v_13495;
wire v_13496;
wire v_13497;
wire v_13498;
wire v_13499;
wire v_13500;
wire v_13501;
wire v_13502;
wire v_13503;
wire v_13504;
wire v_13505;
wire v_13506;
wire v_13507;
wire v_13508;
wire v_13509;
wire v_13510;
wire v_13511;
wire v_13512;
wire v_13513;
wire v_13514;
wire v_13515;
wire v_13516;
wire v_13517;
wire v_13518;
wire v_13519;
wire v_13520;
wire v_13521;
wire v_13522;
wire v_13523;
wire v_13524;
wire v_13525;
wire v_13526;
wire v_13527;
wire v_13528;
wire v_13529;
wire v_13530;
wire v_13531;
wire v_13532;
wire v_13533;
wire v_13534;
wire v_13535;
wire v_13536;
wire v_13537;
wire v_13538;
wire v_13539;
wire v_13540;
wire v_13541;
wire v_13542;
wire v_13543;
wire v_13544;
wire v_13545;
wire v_13546;
wire v_13547;
wire v_13548;
wire v_13549;
wire v_13550;
wire v_13551;
wire v_13552;
wire v_13553;
wire v_13554;
wire v_13555;
wire v_13556;
wire v_13557;
wire v_13558;
wire v_13559;
wire v_13560;
wire v_13561;
wire v_13562;
wire v_13563;
wire v_13564;
wire v_13565;
wire v_13566;
wire v_13567;
wire v_13568;
wire v_13569;
wire v_13570;
wire v_13571;
wire v_13572;
wire v_13573;
wire v_13574;
wire v_13575;
wire v_13576;
wire v_13577;
wire v_13578;
wire v_13579;
wire v_13580;
wire v_13581;
wire v_13582;
wire v_13583;
wire v_13584;
wire v_13585;
wire v_13586;
wire v_13587;
wire v_13588;
wire v_13589;
wire v_13590;
wire v_13591;
wire v_13592;
wire v_13593;
wire v_13594;
wire v_13595;
wire v_13596;
wire v_13597;
wire v_13598;
wire v_13599;
wire v_13600;
wire v_13601;
wire v_13602;
wire v_13603;
wire v_13604;
wire v_13605;
wire v_13606;
wire v_13607;
wire v_13608;
wire v_13609;
wire v_13610;
wire v_13611;
wire v_13612;
wire v_13613;
wire v_13614;
wire v_13615;
wire v_13616;
wire v_13617;
wire v_13618;
wire v_13619;
wire v_13620;
wire v_13621;
wire v_13622;
wire v_13623;
wire v_13624;
wire v_13625;
wire v_13626;
wire v_13627;
wire v_13628;
wire v_13629;
wire v_13630;
wire v_13631;
wire v_13632;
wire v_13633;
wire v_13634;
wire v_13635;
wire v_13636;
wire v_13637;
wire v_13638;
wire v_13639;
wire v_13640;
wire v_13641;
wire v_13642;
wire v_13643;
wire v_13644;
wire v_13645;
wire v_13646;
wire v_13647;
wire v_13648;
wire v_13649;
wire v_13650;
wire v_13651;
wire v_13652;
wire v_13653;
wire v_13654;
wire v_13655;
wire v_13656;
wire v_13657;
wire v_13658;
wire v_13659;
wire v_13660;
wire v_13661;
wire v_13662;
wire v_13663;
wire v_13664;
wire v_13665;
wire v_13666;
wire v_13667;
wire v_13668;
wire v_13669;
wire v_13670;
wire v_13671;
wire v_13672;
wire v_13673;
wire v_13674;
wire v_13675;
wire v_13676;
wire v_13677;
wire v_13678;
wire v_13679;
wire v_13680;
wire v_13681;
wire v_13682;
wire v_13683;
wire v_13684;
wire v_13685;
wire v_13686;
wire v_13687;
wire v_13688;
wire v_13689;
wire v_13690;
wire v_13691;
wire v_13692;
wire v_13693;
wire v_13694;
wire v_13695;
wire v_13696;
wire v_13697;
wire v_13698;
wire v_13699;
wire v_13700;
wire v_13701;
wire v_13702;
wire v_13703;
wire v_13704;
wire v_13705;
wire v_13706;
wire v_13707;
wire v_13708;
wire v_13709;
wire v_13710;
wire v_13711;
wire v_13712;
wire v_13713;
wire v_13714;
wire v_13715;
wire v_13716;
wire v_13717;
wire v_13718;
wire v_13719;
wire v_13720;
wire v_13721;
wire v_13722;
wire v_13723;
wire v_13724;
wire v_13725;
wire v_13726;
wire v_13727;
wire v_13728;
wire v_13729;
wire v_13730;
wire v_13731;
wire v_13732;
wire v_13733;
wire v_13734;
wire v_13735;
wire v_13736;
wire v_13737;
wire v_13738;
wire v_13739;
wire v_13740;
wire v_13741;
wire v_13742;
wire v_13743;
wire v_13744;
wire v_13745;
wire v_13746;
wire v_13747;
wire v_13748;
wire v_13749;
wire v_13750;
wire v_13751;
wire v_13752;
wire v_13753;
wire v_13754;
wire v_13755;
wire v_13756;
wire v_13757;
wire v_13758;
wire v_13759;
wire v_13760;
wire v_13761;
wire v_13762;
wire v_13763;
wire v_13764;
wire v_13765;
wire v_13766;
wire v_13767;
wire v_13768;
wire v_13769;
wire v_13770;
wire v_13771;
wire v_13772;
wire v_13773;
wire v_13774;
wire v_13775;
wire v_13776;
wire v_13777;
wire v_13778;
wire v_13779;
wire v_13780;
wire v_13781;
wire v_13782;
wire v_13783;
wire v_13784;
wire v_13785;
wire v_13786;
wire v_13787;
wire v_13788;
wire v_13789;
wire v_13790;
wire v_13791;
wire v_13792;
wire v_13793;
wire v_13794;
wire v_13795;
wire v_13796;
wire v_13797;
wire v_13798;
wire v_13799;
wire v_13800;
wire v_13801;
wire v_13802;
wire v_13803;
wire v_13804;
wire v_13805;
wire v_13806;
wire v_13807;
wire v_13808;
wire v_13809;
wire v_13810;
wire v_13811;
wire v_13812;
wire v_13813;
wire v_13814;
wire v_13815;
wire v_13816;
wire v_13817;
wire v_13818;
wire v_13819;
wire v_13820;
wire v_13821;
wire v_13822;
wire v_13823;
wire v_13824;
wire v_13825;
wire v_13826;
wire v_13827;
wire v_13828;
wire v_13829;
wire v_13830;
wire v_13831;
wire v_13832;
wire v_13833;
wire v_13834;
wire v_13835;
wire v_13836;
wire v_13837;
wire v_13838;
wire v_13839;
wire v_13840;
wire v_13841;
wire v_13842;
wire v_13843;
wire v_13844;
wire v_13845;
wire v_13846;
wire v_13847;
wire v_13848;
wire v_13849;
wire v_13850;
wire v_13851;
wire v_13852;
wire v_13853;
wire v_13854;
wire v_13855;
wire v_13856;
wire v_13857;
wire v_13858;
wire v_13859;
wire v_13860;
wire v_13861;
wire v_13862;
wire v_13863;
wire v_13864;
wire v_13865;
wire v_13866;
wire v_13867;
wire v_13868;
wire v_13869;
wire v_13870;
wire v_13871;
wire v_13872;
wire v_13873;
wire v_13874;
wire v_13875;
wire v_13876;
wire v_13877;
wire v_13878;
wire v_13879;
wire v_13880;
wire v_13881;
wire v_13882;
wire v_13883;
wire v_13884;
wire v_13885;
wire v_13886;
wire v_13887;
wire v_13888;
wire v_13889;
wire v_13890;
wire v_13891;
wire v_13892;
wire v_13893;
wire v_13894;
wire v_13895;
wire v_13896;
wire v_13897;
wire v_13898;
wire v_13899;
wire v_13900;
wire v_13901;
wire v_13902;
wire v_13903;
wire v_13904;
wire v_13905;
wire v_13906;
wire v_13907;
wire v_13908;
wire v_13909;
wire v_13910;
wire v_13911;
wire v_13912;
wire v_13913;
wire v_13914;
wire v_13915;
wire v_13916;
wire v_13917;
wire v_13918;
wire v_13919;
wire v_13920;
wire v_13921;
wire x_1;
assign v_1 = 1;
assign v_220 = 1;
assign v_226 = 1;
assign v_231 = 1;
assign v_250 = 1;
assign v_273 = 1;
assign v_339 = 1;
assign v_487 = 1;
assign v_490 = 1;
assign v_495 = 1;
assign v_514 = 1;
assign v_538 = 1;
assign v_550 = 1;
assign v_556 = 1;
assign v_564 = 1;
assign v_608 = 1;
assign v_614 = 1;
assign v_622 = 1;
assign v_664 = 1;
assign v_667 = 1;
assign v_714 = 1;
assign v_720 = 1;
assign v_728 = 1;
assign v_754 = 1;
assign v_756 = 1;
assign v_767 = 1;
assign v_769 = 1;
assign v_773 = 1;
assign v_783 = 1;
assign v_789 = 1;
assign v_1537 = 1;
assign v_3159 = 1;
assign v_7086 = 1;
assign v_7092 = 1;
assign v_7097 = 1;
assign v_7116 = 1;
assign v_7139 = 1;
assign v_7205 = 1;
assign v_7353 = 1;
assign v_7356 = 1;
assign v_7361 = 1;
assign v_7380 = 1;
assign v_7404 = 1;
assign v_7416 = 1;
assign v_7422 = 1;
assign v_7430 = 1;
assign v_7474 = 1;
assign v_7480 = 1;
assign v_7488 = 1;
assign v_7530 = 1;
assign v_7533 = 1;
assign v_7580 = 1;
assign v_7586 = 1;
assign v_7594 = 1;
assign v_7620 = 1;
assign v_7622 = 1;
assign v_7633 = 1;
assign v_7635 = 1;
assign v_7639 = 1;
assign v_7649 = 1;
assign v_7655 = 1;
assign v_8241 = 1;
assign v_9645 = 1;
assign v_6 = ~v_4 & ~v_5;
assign v_9 = ~v_7 & v_8;
assign v_10 = ~v_6 & ~v_9;
assign v_11 = ~v_4 & ~v_5;
assign v_12 = ~v_7 & v_8;
assign v_13 = ~v_11 & ~v_12;
assign v_14 = v_10 & v_13;
assign v_15 = ~v_4 & ~v_5;
assign v_16 = ~v_7 & v_8;
assign v_17 = ~v_15 & ~v_16;
assign v_18 = v_14 & v_17;
assign v_19 = ~v_4 & ~v_5;
assign v_20 = ~v_7 & v_8;
assign v_21 = ~v_19 & ~v_20;
assign v_22 = v_18 & v_21;
assign v_23 = ~v_4 & ~v_5;
assign v_24 = ~v_7 & v_8;
assign v_25 = ~v_23 & ~v_24;
assign v_26 = v_22 & v_25;
assign v_27 = ~v_4 & ~v_5;
assign v_28 = ~v_7 & v_8;
assign v_29 = ~v_27 & ~v_28;
assign v_30 = v_26 & v_29;
assign v_31 = ~v_4 & ~v_5;
assign v_32 = ~v_7 & v_8;
assign v_33 = ~v_31 & ~v_32;
assign v_34 = v_30 & v_33;
assign v_35 = ~v_4 & ~v_5;
assign v_36 = ~v_7 & v_8;
assign v_37 = ~v_35 & ~v_36;
assign v_38 = v_34 & v_37;
assign v_39 = ~v_4 & ~v_5;
assign v_40 = ~v_7 & v_8;
assign v_41 = ~v_39 & ~v_40;
assign v_42 = v_38 & v_41;
assign v_43 = ~v_4 & ~v_5;
assign v_44 = ~v_7 & v_8;
assign v_45 = ~v_43 & ~v_44;
assign v_46 = v_42 & v_45;
assign v_47 = ~v_4 & ~v_5;
assign v_48 = ~v_7 & v_8;
assign v_49 = ~v_47 & ~v_48;
assign v_50 = v_46 & v_49;
assign v_51 = ~v_4 & ~v_5;
assign v_52 = ~v_7 & v_8;
assign v_53 = ~v_51 & ~v_52;
assign v_54 = v_50 & v_53;
assign v_55 = ~v_4 & ~v_5;
assign v_56 = ~v_7 & v_8;
assign v_57 = ~v_55 & ~v_56;
assign v_58 = v_54 & v_57;
assign v_59 = ~v_4 & ~v_5;
assign v_60 = ~v_7 & v_8;
assign v_61 = ~v_59 & ~v_60;
assign v_62 = v_58 & v_61;
assign v_63 = ~v_4 & ~v_5;
assign v_64 = ~v_7 & v_8;
assign v_65 = ~v_63 & ~v_64;
assign v_66 = v_62 & v_65;
assign v_67 = ~v_4 & ~v_5;
assign v_68 = ~v_7 & v_8;
assign v_69 = ~v_67 & ~v_68;
assign v_70 = v_66 & v_69;
assign v_71 = ~v_4 & ~v_5;
assign v_72 = ~v_7 & v_8;
assign v_73 = ~v_71 & ~v_72;
assign v_74 = v_70 & v_73;
assign v_75 = ~v_4 & ~v_5;
assign v_76 = ~v_7 & v_8;
assign v_77 = ~v_75 & ~v_76;
assign v_78 = v_74 & v_77;
assign v_79 = ~v_4 & ~v_5;
assign v_80 = ~v_7 & v_8;
assign v_81 = ~v_79 & ~v_80;
assign v_82 = v_78 & v_81;
assign v_83 = ~v_4 & ~v_5;
assign v_84 = ~v_7 & v_8;
assign v_85 = ~v_83 & ~v_84;
assign v_86 = v_82 & v_85;
assign v_87 = ~v_4 & ~v_5;
assign v_88 = ~v_7 & v_8;
assign v_89 = ~v_87 & ~v_88;
assign v_90 = v_86 & v_89;
assign v_91 = ~v_4 & ~v_5;
assign v_92 = ~v_7 & v_8;
assign v_93 = ~v_91 & ~v_92;
assign v_94 = v_90 & v_93;
assign v_95 = ~v_4 & ~v_5;
assign v_96 = ~v_7 & v_8;
assign v_97 = ~v_95 & ~v_96;
assign v_98 = v_94 & v_97;
assign v_99 = ~v_4 & ~v_5;
assign v_100 = ~v_7 & v_8;
assign v_101 = ~v_99 & ~v_100;
assign v_102 = v_98 & v_101;
assign v_103 = ~v_4 & ~v_5;
assign v_104 = ~v_7 & v_8;
assign v_105 = ~v_103 & ~v_104;
assign v_106 = v_102 & v_105;
assign v_107 = ~v_4 & ~v_5;
assign v_108 = ~v_7 & v_8;
assign v_109 = ~v_107 & ~v_108;
assign v_110 = v_106 & v_109;
assign v_111 = ~v_4 & ~v_5;
assign v_112 = ~v_7 & v_8;
assign v_113 = ~v_111 & ~v_112;
assign v_114 = v_110 & v_113;
assign v_115 = ~v_4 & ~v_5;
assign v_116 = ~v_7 & v_8;
assign v_117 = ~v_115 & ~v_116;
assign v_118 = v_114 & v_117;
assign v_119 = ~v_4 & ~v_5;
assign v_120 = ~v_7 & v_8;
assign v_121 = ~v_119 & ~v_120;
assign v_122 = v_118 & v_121;
assign v_123 = ~v_4 & ~v_5;
assign v_124 = ~v_7 & v_8;
assign v_125 = ~v_123 & ~v_124;
assign v_126 = v_122 & v_125;
assign v_127 = ~v_4 & ~v_5;
assign v_128 = ~v_7 & v_8;
assign v_129 = ~v_127 & ~v_128;
assign v_130 = v_126 & v_129;
assign v_131 = ~v_4 & ~v_5;
assign v_132 = ~v_7 & v_8;
assign v_133 = ~v_131 & ~v_132;
assign v_134 = v_130 & v_133;
assign v_135 = ~v_4 & ~v_5;
assign v_136 = ~v_7 & v_8;
assign v_137 = ~v_135 & ~v_136;
assign v_138 = v_134 & v_137;
assign v_139 = ~v_4 & ~v_5;
assign v_140 = ~v_7 & v_8;
assign v_141 = ~v_139 & ~v_140;
assign v_142 = v_138 & v_141;
assign v_143 = ~v_4 & ~v_5;
assign v_144 = ~v_7 & v_8;
assign v_145 = ~v_143 & ~v_144;
assign v_146 = v_142 & v_145;
assign v_147 = ~v_4 & ~v_5;
assign v_148 = ~v_7 & v_8;
assign v_149 = ~v_147 & ~v_148;
assign v_150 = v_146 & v_149;
assign v_151 = ~v_4 & ~v_5;
assign v_152 = ~v_7 & v_8;
assign v_153 = ~v_151 & ~v_152;
assign v_154 = v_150 & v_153;
assign v_155 = ~v_4 & ~v_5;
assign v_156 = ~v_7 & v_8;
assign v_157 = ~v_155 & ~v_156;
assign v_158 = v_154 & v_157;
assign v_159 = ~v_4 & ~v_5;
assign v_160 = ~v_7 & v_8;
assign v_161 = ~v_159 & ~v_160;
assign v_162 = v_158 & v_161;
assign v_163 = ~v_4 & ~v_5;
assign v_164 = ~v_7 & v_8;
assign v_165 = ~v_163 & ~v_164;
assign v_166 = v_162 & v_165;
assign v_167 = ~v_4 & ~v_5;
assign v_168 = ~v_7 & v_8;
assign v_169 = ~v_167 & ~v_168;
assign v_170 = v_166 & v_169;
assign v_171 = ~v_4 & ~v_5;
assign v_172 = ~v_7 & v_8;
assign v_173 = ~v_171 & ~v_172;
assign v_174 = v_170 & v_173;
assign v_175 = ~v_4 & ~v_5;
assign v_176 = ~v_7 & v_8;
assign v_177 = ~v_175 & ~v_176;
assign v_178 = v_174 & v_177;
assign v_179 = ~v_4 & ~v_5;
assign v_180 = ~v_7 & v_8;
assign v_181 = ~v_179 & ~v_180;
assign v_182 = v_178 & v_181;
assign v_183 = ~v_4 & ~v_5;
assign v_184 = ~v_7 & v_8;
assign v_185 = ~v_183 & ~v_184;
assign v_186 = v_182 & v_185;
assign v_187 = ~v_4 & ~v_5;
assign v_188 = ~v_7 & v_8;
assign v_189 = ~v_187 & ~v_188;
assign v_190 = v_186 & v_189;
assign v_191 = ~v_4 & ~v_5;
assign v_192 = ~v_7 & v_8;
assign v_193 = ~v_191 & ~v_192;
assign v_194 = v_190 & v_193;
assign v_195 = ~v_4 & ~v_5;
assign v_196 = ~v_7 & v_8;
assign v_197 = ~v_195 & ~v_196;
assign v_198 = v_194 & v_197;
assign v_199 = ~v_4 & ~v_5;
assign v_200 = ~v_7 & v_8;
assign v_201 = ~v_199 & ~v_200;
assign v_202 = v_198 & v_201;
assign v_203 = ~v_7 & v_8;
assign v_204 = v_202 & ~v_203;
assign v_205 = ~v_7 & v_8;
assign v_206 = v_204 & ~v_205;
assign v_207 = ~v_7 & v_8;
assign v_208 = v_206 & ~v_207;
assign v_209 = ~v_7 & v_8;
assign v_210 = v_208 & ~v_209;
assign v_211 = ~v_7 & v_8;
assign v_212 = v_210 & ~v_211;
assign v_215 = v_213 & v_214;
assign v_216 = v_213 & ~v_214;
assign v_218 = v_212 & v_217;
assign v_222 = v_221;
assign v_223 = ~v_221;
assign v_228 = v_227;
assign v_233 = ~v_232;
assign v_235 = v_232 & v_234;
assign v_238 = v_232 & ~v_234 & v_236 & v_237;
assign v_240 = v_232 & ~v_234 & v_236 & ~v_237 & ~v_239;
assign v_242 = v_232 & ~v_234 & ~v_236 & ~v_241;
assign v_244 = v_232 & ~v_234 & ~v_236 & v_241 & v_243;
assign v_246 = v_12875 & v_12876;
assign v_248 = v_12877 & v_12878;
assign v_252 = v_12879 & v_12880;
assign v_253 = v_12881 & v_12882;
assign v_256 = v_254 & v_255;
assign v_257 = v_254 & ~v_255;
assign v_259 = v_12883 & v_12884;
assign v_261 = ~v_227 & ~v_229 & v_260;
assign v_263 = ~v_227 & v_229 & ~v_262;
assign v_265 = ~v_227 & v_229 & v_262 & ~v_264;
assign v_266 = ~v_227 & v_229 & v_262 & v_264;
assign v_269 = v_267 & v_268;
assign v_270 = v_267 & ~v_268;
assign v_275 = v_224 & v_271 & v_274;
assign v_276 = v_224 & v_271 & ~v_274;
assign v_278 = v_218 & v_277;
assign v_282 = v_280 & v_281;
assign v_284 = v_280 & ~v_281 & v_283;
assign v_287 = v_285 & ~v_286;
assign v_289 = v_285 & v_286 & v_288;
assign v_290 = v_285 & v_286 & ~v_288;
assign v_294 = v_279 & v_291 & v_292 & v_293;
assign v_296 = v_279 & v_291 & v_292 & ~v_293 & v_295;
assign v_299 = ~v_297 & v_298;
assign v_301 = v_279 & v_291 & ~v_292 & v_300;
assign v_304 = v_302 & v_303;
assign v_305 = v_302 & ~v_303;
assign v_307 = v_278 & v_306;
assign v_310 = ~v_308 & ~v_309;
assign v_313 = v_311 & v_312;
assign v_314 = v_311 & ~v_312;
assign v_317 = v_315 & ~v_316;
assign v_319 = v_315 & v_316 & v_318;
assign v_320 = v_315 & v_316 & ~v_318;
assign v_323 = v_321 & v_322;
assign v_325 = v_321 & ~v_322 & v_324;
assign v_327 = v_321 & ~v_322 & ~v_324 & v_326;
assign v_328 = v_321 & ~v_322 & ~v_324 & ~v_326;
assign v_330 = ~v_308 & v_309 & v_329;
assign v_332 = v_307 & v_331;
assign v_335 = v_333 & ~v_334;
assign v_337 = v_333 & v_334 & ~v_336;
assign v_341 = v_333 & v_334 & v_336 & v_340;
assign v_342 = v_333 & v_334 & v_336 & ~v_340;
assign v_344 = v_332 & v_343;
assign v_347 = v_345 & v_346;
assign v_349 = v_345 & ~v_346 & v_348;
assign v_351 = v_345 & ~v_346 & ~v_348 & v_350;
assign v_353 = v_345 & ~v_346 & ~v_348 & ~v_350 & v_352;
assign v_355 = v_12885 & v_12886;
assign v_358 = v_356 & v_357;
assign v_361 = v_359 & v_360;
assign v_363 = v_359 & ~v_360 & v_362;
assign v_365 = v_359 & ~v_360 & ~v_362 & v_364;
assign v_367 = v_359 & ~v_360 & ~v_362 & ~v_364 & v_366;
assign v_368 = v_359 & ~v_360 & ~v_362 & ~v_364 & ~v_366;
assign v_371 = v_356 & ~v_357 & v_369 & v_370;
assign v_374 = v_372 & v_373;
assign v_376 = v_372 & ~v_373 & v_375;
assign v_378 = v_372 & ~v_373 & ~v_375 & v_377;
assign v_380 = v_372 & ~v_373 & ~v_375 & ~v_377 & v_379;
assign v_382 = v_12887 & v_12888;
assign v_383 = v_12889 & v_12890;
assign v_386 = v_384 & v_385;
assign v_387 = v_384 & ~v_385;
assign v_390 = v_12891 & v_12892;
assign v_393 = v_391 & v_392;
assign v_395 = v_391 & ~v_392 & v_394;
assign v_397 = v_391 & ~v_392 & ~v_394 & v_396;
assign v_399 = v_391 & ~v_392 & ~v_394 & ~v_396 & ~v_398;
assign v_401 = v_12893 & v_12894;
assign v_402 = v_12895 & v_12896;
assign v_404 = v_12897 & v_12898;
assign v_407 = v_405 & v_406;
assign v_408 = v_405 & ~v_406;
assign v_412 = v_410 & v_411;
assign v_414 = v_410 & ~v_411 & v_413;
assign v_416 = v_410 & ~v_411 & ~v_413 & v_415;
assign v_418 = v_410 & ~v_411 & ~v_413 & ~v_415 & v_417;
assign v_420 = v_12899 & v_12900;
assign v_423 = v_421 & v_422;
assign v_426 = v_424 & v_425;
assign v_428 = v_424 & ~v_425 & v_427;
assign v_430 = v_424 & ~v_425 & ~v_427 & v_429;
assign v_432 = v_424 & ~v_425 & ~v_427 & ~v_429 & v_431;
assign v_433 = v_424 & ~v_425 & ~v_427 & ~v_429 & ~v_431;
assign v_436 = v_421 & ~v_422 & v_434 & v_435;
assign v_439 = v_437 & v_438;
assign v_441 = v_437 & ~v_438 & v_440;
assign v_443 = v_437 & ~v_438 & ~v_440 & v_442;
assign v_445 = v_437 & ~v_438 & ~v_440 & ~v_442 & v_444;
assign v_447 = v_12901 & v_12902;
assign v_448 = v_12903 & v_12904;
assign v_451 = v_449 & v_450;
assign v_452 = v_449 & ~v_450;
assign v_455 = v_12905 & v_12906;
assign v_458 = v_456 & v_457;
assign v_460 = v_456 & ~v_457 & v_459;
assign v_462 = v_456 & ~v_457 & ~v_459 & v_461;
assign v_464 = v_456 & ~v_457 & ~v_459 & ~v_461 & ~v_463;
assign v_466 = v_12907 & v_12908;
assign v_467 = v_12909 & v_12910;
assign v_469 = v_12911 & v_12912;
assign v_472 = v_470 & v_471;
assign v_473 = v_470 & ~v_471;
assign v_476 = v_409 & v_474 & v_475;
assign v_478 = v_409 & v_474 & ~v_475 & v_477;
assign v_479 = v_409 & v_474 & ~v_475 & ~v_477;
assign v_482 = v_480 & v_481;
assign v_483 = v_480 & ~v_481;
assign v_485 = v_344 & v_484;
assign v_488 = v_485;
assign v_492 = v_491;
assign v_497 = ~v_496;
assign v_499 = v_496 & v_498;
assign v_502 = v_496 & ~v_498 & v_500 & v_501;
assign v_504 = v_496 & ~v_498 & v_500 & ~v_501 & ~v_503;
assign v_506 = v_496 & ~v_498 & ~v_500 & ~v_505;
assign v_508 = v_496 & ~v_498 & ~v_500 & v_505 & v_507;
assign v_510 = v_12913 & v_12914;
assign v_512 = v_12915 & v_12916;
assign v_516 = v_12917 & v_12918;
assign v_517 = v_12919 & v_12920;
assign v_520 = v_518 & v_519;
assign v_521 = v_518 & ~v_519;
assign v_523 = v_12921 & v_12922;
assign v_525 = ~v_491 & ~v_493 & v_524;
assign v_527 = ~v_491 & v_493 & ~v_526;
assign v_529 = ~v_491 & v_493 & v_526 & ~v_528;
assign v_530 = ~v_491 & v_493 & v_526 & v_528;
assign v_533 = v_531 & v_532;
assign v_534 = v_531 & ~v_532;
assign v_536 = v_488 & v_535;
assign v_539 = v_3 & v_536;
assign v_540 = ~v_3 & v_488 & v_535;
assign v_544 = v_542 & v_543;
assign v_545 = v_542 & ~v_543;
assign v_548 = v_546 & v_547;
assign v_552 = v_546 & ~v_547 & ~v_551;
assign v_553 = v_546 & ~v_547 & v_551;
assign v_557 = v_554;
assign v_560 = v_558 & v_559;
assign v_562 = v_558 & ~v_559 & v_561;
assign v_566 = v_558 & ~v_559 & ~v_561 & v_565;
assign v_567 = v_558 & ~v_559 & ~v_561 & ~v_565;
assign v_570 = v_568 & v_569;
assign v_572 = v_568 & ~v_569 & v_571;
assign v_575 = v_573 & v_574;
assign v_576 = v_573 & ~v_574;
assign v_579 = v_568 & ~v_569 & ~v_571 & v_577 & v_578;
assign v_580 = v_568 & ~v_569 & ~v_571 & v_577 & ~v_578;
assign v_582 = v_541 & v_581;
assign v_585 = ~v_583 & v_584;
assign v_587 = ~v_583 & ~v_584 & v_586;
assign v_590 = v_588 & v_589;
assign v_592 = v_588 & ~v_589 & v_591;
assign v_595 = v_593 & ~v_594;
assign v_596 = v_588 & ~v_589 & ~v_591;
assign v_597 = v_593 & v_594;
assign v_599 = v_582 & v_598;
assign v_602 = v_600 & v_601;
assign v_603 = v_600 & ~v_601;
assign v_606 = v_604 & v_605;
assign v_610 = v_604 & ~v_605 & ~v_609;
assign v_611 = v_604 & ~v_605 & v_609;
assign v_615 = v_612;
assign v_618 = v_616 & v_617;
assign v_620 = v_616 & ~v_617 & v_619;
assign v_624 = v_616 & ~v_617 & ~v_619 & v_623;
assign v_625 = v_616 & ~v_617 & ~v_619 & ~v_623;
assign v_628 = v_626 & v_627;
assign v_630 = v_626 & ~v_627 & v_629;
assign v_633 = v_631 & v_632;
assign v_634 = v_631 & ~v_632;
assign v_637 = v_626 & ~v_627 & ~v_629 & v_635 & v_636;
assign v_638 = v_626 & ~v_627 & ~v_629 & v_635 & ~v_636;
assign v_640 = v_2 & v_599 & v_639;
assign v_642 = v_641 & v_541 & v_581;
assign v_644 = v_643 & v_536;
assign v_646 = v_645 & v_536;
assign v_648 = v_647 & v_488 & v_535;
assign v_650 = v_649 & v_488 & v_535;
assign v_651 = ~v_649 & v_485;
assign v_653 = ~v_647 & v_652;
assign v_655 = ~v_645 & v_654;
assign v_657 = ~v_643 & v_656;
assign v_659 = ~v_641 & v_658;
assign v_661 = ~v_2 & v_660;
assign v_665 = v_662;
assign v_668 = v_665;
assign v_671 = v_669 & ~v_670;
assign v_673 = v_669 & v_670 & ~v_672;
assign v_676 = v_669 & v_670 & v_672 & ~v_674 & ~v_675;
assign v_677 = v_669 & v_670 & v_672 & v_674;
assign v_678 = v_669 & v_670 & v_672 & ~v_674 & v_675;
assign v_681 = v_679 & v_680;
assign v_683 = v_679 & ~v_680 & v_682;
assign v_686 = ~v_684 & v_685;
assign v_688 = ~v_684 & ~v_685 & v_687;
assign v_691 = v_689 & v_690;
assign v_693 = v_689 & ~v_690 & v_692;
assign v_696 = v_694 & ~v_695;
assign v_697 = v_689 & ~v_690 & ~v_692;
assign v_698 = v_694 & v_695;
assign v_701 = v_679 & ~v_680 & ~v_682 & v_699 & v_700;
assign v_702 = v_679 & ~v_680 & ~v_682 & v_699 & ~v_700;
assign v_704 = v_668 & v_703;
assign v_708 = v_706 & v_707;
assign v_709 = v_706 & ~v_707;
assign v_712 = v_710 & v_711;
assign v_716 = v_710 & ~v_711 & ~v_715;
assign v_717 = v_710 & ~v_711 & v_715;
assign v_721 = v_718;
assign v_725 = v_705 & v_722 & v_723 & ~v_724;
assign v_730 = v_12923 & v_12924;
assign v_732 = v_12925 & v_12926;
assign v_734 = v_12927 & v_12928;
assign v_736 = v_12929 & v_12930;
assign v_740 = v_737 & ~v_738 & v_739;
assign v_741 = v_737 & ~v_738 & ~v_739;
assign v_743 = v_737 & v_738 & v_742;
assign v_744 = v_737 & v_738 & ~v_742;
assign v_748 = v_746 & v_747;
assign v_749 = v_746 & ~v_747;
assign v_752 = v_750 & v_751;
assign v_757 = v_750 & ~v_751;
assign v_761 = v_759 & v_760;
assign v_762 = v_759 & ~v_760;
assign v_765 = v_763 & v_764;
assign v_770 = v_763 & ~v_764;
assign v_774 = v_745 & v_758 & v_771;
assign v_777 = v_775 & v_776;
assign v_778 = v_775 & ~v_776;
assign v_781 = v_779 & v_780;
assign v_785 = v_779 & ~v_780 & ~v_784;
assign v_786 = v_779 & ~v_780 & v_784;
assign v_790 = v_787;
assign v_793 = v_705 & v_722 & ~v_723 & v_791 & v_792;
assign v_794 = v_705 & v_722 & ~v_723 & v_791 & ~v_792;
assign v_795 = v_705 & v_722 & v_723 & v_724 & v_726;
assign v_797 = v_704 & v_796;
assign v_802 = v_800 & v_801;
assign v_803 = v_800 & ~v_801;
assign v_806 = v_804 & v_805;
assign v_807 = v_804 & ~v_805;
assign v_810 = v_808 & ~v_809;
assign v_812 = v_808 & v_809 & v_811;
assign v_813 = v_808 & v_809 & ~v_811;
assign v_816 = v_798 & v_799 & v_814 & v_815;
assign v_818 = v_798 & ~v_799 & v_817;
assign v_819 = v_798 & v_799 & v_814 & ~v_815;
assign v_820 = v_798 & ~v_799 & ~v_817;
assign v_825 = v_823 & v_824;
assign v_826 = v_823 & ~v_824;
assign v_829 = v_827 & v_828;
assign v_830 = v_827 & ~v_828;
assign v_833 = v_831 & ~v_832;
assign v_835 = v_831 & v_832 & v_834;
assign v_836 = v_831 & v_832 & ~v_834;
assign v_839 = v_821 & v_822 & v_837 & v_838;
assign v_841 = v_821 & ~v_822 & v_840;
assign v_842 = v_821 & v_822 & v_837 & ~v_838;
assign v_843 = v_821 & ~v_822 & ~v_840;
assign v_848 = v_846 & v_847;
assign v_849 = v_846 & ~v_847;
assign v_852 = v_850 & v_851;
assign v_853 = v_850 & ~v_851;
assign v_856 = v_854 & ~v_855;
assign v_858 = v_854 & v_855 & v_857;
assign v_859 = v_854 & v_855 & ~v_857;
assign v_862 = v_844 & v_845 & v_860 & v_861;
assign v_864 = v_844 & ~v_845 & v_863;
assign v_865 = v_844 & v_845 & v_860 & ~v_861;
assign v_866 = v_844 & ~v_845 & ~v_863;
assign v_871 = v_867 & v_868 & ~v_869 & v_870;
assign v_873 = v_867 & ~v_868 & v_872;
assign v_874 = v_867 & ~v_868 & ~v_872;
assign v_875 = v_867 & v_868 & ~v_869 & ~v_870;
assign v_876 = v_867 & v_868 & v_869;
assign v_878 = v_797 & v_877;
assign v_883 = v_881 & v_882;
assign v_884 = v_881 & ~v_882;
assign v_887 = v_885 & v_886;
assign v_888 = v_885 & ~v_886;
assign v_891 = v_889 & ~v_890;
assign v_893 = v_889 & v_890 & v_892;
assign v_894 = v_889 & v_890 & ~v_892;
assign v_897 = v_879 & v_880 & v_895 & v_896;
assign v_899 = v_879 & ~v_880 & v_898;
assign v_900 = v_879 & v_880 & v_895 & ~v_896;
assign v_901 = v_879 & ~v_880 & ~v_898;
assign v_906 = v_904 & v_905;
assign v_907 = v_904 & ~v_905;
assign v_910 = v_908 & v_909;
assign v_911 = v_908 & ~v_909;
assign v_914 = v_912 & ~v_913;
assign v_916 = v_912 & v_913 & v_915;
assign v_917 = v_912 & v_913 & ~v_915;
assign v_920 = v_902 & v_903 & v_918 & v_919;
assign v_922 = v_902 & ~v_903 & v_921;
assign v_923 = v_902 & v_903 & v_918 & ~v_919;
assign v_924 = v_902 & ~v_903 & ~v_921;
assign v_929 = v_927 & v_928;
assign v_930 = v_927 & ~v_928;
assign v_933 = v_931 & v_932;
assign v_934 = v_931 & ~v_932;
assign v_937 = v_935 & ~v_936;
assign v_939 = v_935 & v_936 & v_938;
assign v_940 = v_935 & v_936 & ~v_938;
assign v_943 = v_925 & v_926 & v_941 & v_942;
assign v_945 = v_925 & ~v_926 & v_944;
assign v_946 = v_925 & v_926 & v_941 & ~v_942;
assign v_947 = v_925 & ~v_926 & ~v_944;
assign v_952 = v_948 & v_949 & ~v_950 & v_951;
assign v_954 = v_948 & ~v_949 & v_953;
assign v_955 = v_948 & ~v_949 & ~v_953;
assign v_956 = v_948 & v_949 & ~v_950 & ~v_951;
assign v_957 = v_948 & v_949 & v_950;
assign v_959 = v_878 & v_958;
assign v_964 = v_962 & v_963;
assign v_965 = v_962 & ~v_963;
assign v_968 = v_966 & v_967;
assign v_969 = v_966 & ~v_967;
assign v_972 = v_970 & ~v_971;
assign v_974 = v_970 & v_971 & v_973;
assign v_975 = v_970 & v_971 & ~v_973;
assign v_978 = v_960 & v_961 & v_976 & v_977;
assign v_980 = v_960 & ~v_961 & v_979;
assign v_981 = v_960 & v_961 & v_976 & ~v_977;
assign v_982 = v_960 & ~v_961 & ~v_979;
assign v_987 = v_985 & v_986;
assign v_988 = v_985 & ~v_986;
assign v_991 = v_989 & v_990;
assign v_992 = v_989 & ~v_990;
assign v_995 = v_993 & ~v_994;
assign v_997 = v_993 & v_994 & v_996;
assign v_998 = v_993 & v_994 & ~v_996;
assign v_1001 = v_983 & v_984 & v_999 & v_1000;
assign v_1003 = v_983 & ~v_984 & v_1002;
assign v_1004 = v_983 & v_984 & v_999 & ~v_1000;
assign v_1005 = v_983 & ~v_984 & ~v_1002;
assign v_1010 = v_1008 & v_1009;
assign v_1011 = v_1008 & ~v_1009;
assign v_1014 = v_1012 & v_1013;
assign v_1015 = v_1012 & ~v_1013;
assign v_1018 = v_1016 & ~v_1017;
assign v_1020 = v_1016 & v_1017 & v_1019;
assign v_1021 = v_1016 & v_1017 & ~v_1019;
assign v_1024 = v_1006 & v_1007 & v_1022 & v_1023;
assign v_1026 = v_1006 & ~v_1007 & v_1025;
assign v_1027 = v_1006 & v_1007 & v_1022 & ~v_1023;
assign v_1028 = v_1006 & ~v_1007 & ~v_1025;
assign v_1033 = v_1029 & v_1030 & ~v_1031 & v_1032;
assign v_1035 = v_1029 & ~v_1030 & v_1034;
assign v_1036 = v_1029 & ~v_1030 & ~v_1034;
assign v_1037 = v_1029 & v_1030 & ~v_1031 & ~v_1032;
assign v_1038 = v_1029 & v_1030 & v_1031;
assign v_1040 = v_959 & v_1039;
assign v_1045 = v_1043 & v_1044;
assign v_1046 = v_1043 & ~v_1044;
assign v_1049 = v_1047 & v_1048;
assign v_1050 = v_1047 & ~v_1048;
assign v_1053 = v_1051 & ~v_1052;
assign v_1055 = v_1051 & v_1052 & v_1054;
assign v_1056 = v_1051 & v_1052 & ~v_1054;
assign v_1059 = v_1041 & v_1042 & v_1057 & v_1058;
assign v_1061 = v_1041 & ~v_1042 & v_1060;
assign v_1062 = v_1041 & v_1042 & v_1057 & ~v_1058;
assign v_1063 = v_1041 & ~v_1042 & ~v_1060;
assign v_1068 = v_1066 & v_1067;
assign v_1069 = v_1066 & ~v_1067;
assign v_1072 = v_1070 & v_1071;
assign v_1073 = v_1070 & ~v_1071;
assign v_1076 = v_1074 & ~v_1075;
assign v_1078 = v_1074 & v_1075 & v_1077;
assign v_1079 = v_1074 & v_1075 & ~v_1077;
assign v_1082 = v_1064 & v_1065 & v_1080 & v_1081;
assign v_1084 = v_1064 & ~v_1065 & v_1083;
assign v_1085 = v_1064 & v_1065 & v_1080 & ~v_1081;
assign v_1086 = v_1064 & ~v_1065 & ~v_1083;
assign v_1091 = v_1089 & v_1090;
assign v_1092 = v_1089 & ~v_1090;
assign v_1095 = v_1093 & v_1094;
assign v_1096 = v_1093 & ~v_1094;
assign v_1099 = v_1097 & ~v_1098;
assign v_1101 = v_1097 & v_1098 & v_1100;
assign v_1102 = v_1097 & v_1098 & ~v_1100;
assign v_1105 = v_1087 & v_1088 & v_1103 & v_1104;
assign v_1107 = v_1087 & ~v_1088 & v_1106;
assign v_1108 = v_1087 & v_1088 & v_1103 & ~v_1104;
assign v_1109 = v_1087 & ~v_1088 & ~v_1106;
assign v_1114 = v_1110 & v_1111 & ~v_1112 & v_1113;
assign v_1116 = v_1110 & ~v_1111 & v_1115;
assign v_1117 = v_1110 & ~v_1111 & ~v_1115;
assign v_1118 = v_1110 & v_1111 & ~v_1112 & ~v_1113;
assign v_1119 = v_1110 & v_1111 & v_1112;
assign v_1121 = v_1040 & v_1120;
assign v_1126 = v_1124 & v_1125;
assign v_1127 = v_1124 & ~v_1125;
assign v_1130 = v_1128 & v_1129;
assign v_1131 = v_1128 & ~v_1129;
assign v_1134 = v_1132 & ~v_1133;
assign v_1136 = v_1132 & v_1133 & v_1135;
assign v_1137 = v_1132 & v_1133 & ~v_1135;
assign v_1140 = v_1122 & v_1123 & v_1138 & v_1139;
assign v_1142 = v_1122 & ~v_1123 & v_1141;
assign v_1143 = v_1122 & v_1123 & v_1138 & ~v_1139;
assign v_1144 = v_1122 & ~v_1123 & ~v_1141;
assign v_1149 = v_1147 & v_1148;
assign v_1150 = v_1147 & ~v_1148;
assign v_1153 = v_1151 & v_1152;
assign v_1154 = v_1151 & ~v_1152;
assign v_1157 = v_1155 & ~v_1156;
assign v_1159 = v_1155 & v_1156 & v_1158;
assign v_1160 = v_1155 & v_1156 & ~v_1158;
assign v_1163 = v_1145 & v_1146 & v_1161 & v_1162;
assign v_1165 = v_1145 & ~v_1146 & v_1164;
assign v_1166 = v_1145 & v_1146 & v_1161 & ~v_1162;
assign v_1167 = v_1145 & ~v_1146 & ~v_1164;
assign v_1172 = v_1170 & v_1171;
assign v_1173 = v_1170 & ~v_1171;
assign v_1176 = v_1174 & v_1175;
assign v_1177 = v_1174 & ~v_1175;
assign v_1180 = v_1178 & ~v_1179;
assign v_1182 = v_1178 & v_1179 & v_1181;
assign v_1183 = v_1178 & v_1179 & ~v_1181;
assign v_1186 = v_1168 & v_1169 & v_1184 & v_1185;
assign v_1188 = v_1168 & ~v_1169 & v_1187;
assign v_1189 = v_1168 & v_1169 & v_1184 & ~v_1185;
assign v_1190 = v_1168 & ~v_1169 & ~v_1187;
assign v_1195 = v_1191 & v_1192 & ~v_1193 & v_1194;
assign v_1197 = v_1191 & ~v_1192 & v_1196;
assign v_1198 = v_1191 & ~v_1192 & ~v_1196;
assign v_1199 = v_1191 & v_1192 & ~v_1193 & ~v_1194;
assign v_1200 = v_1191 & v_1192 & v_1193;
assign v_1202 = v_1121 & v_1201;
assign v_1207 = v_1205 & v_1206;
assign v_1208 = v_1205 & ~v_1206;
assign v_1211 = v_1209 & v_1210;
assign v_1212 = v_1209 & ~v_1210;
assign v_1215 = v_1213 & ~v_1214;
assign v_1217 = v_1213 & v_1214 & v_1216;
assign v_1218 = v_1213 & v_1214 & ~v_1216;
assign v_1221 = v_1203 & v_1204 & v_1219 & v_1220;
assign v_1223 = v_1203 & ~v_1204 & v_1222;
assign v_1224 = v_1203 & v_1204 & v_1219 & ~v_1220;
assign v_1225 = v_1203 & ~v_1204 & ~v_1222;
assign v_1230 = v_1228 & v_1229;
assign v_1231 = v_1228 & ~v_1229;
assign v_1234 = v_1232 & v_1233;
assign v_1235 = v_1232 & ~v_1233;
assign v_1238 = v_1236 & ~v_1237;
assign v_1240 = v_1236 & v_1237 & v_1239;
assign v_1241 = v_1236 & v_1237 & ~v_1239;
assign v_1244 = v_1226 & v_1227 & v_1242 & v_1243;
assign v_1246 = v_1226 & ~v_1227 & v_1245;
assign v_1247 = v_1226 & v_1227 & v_1242 & ~v_1243;
assign v_1248 = v_1226 & ~v_1227 & ~v_1245;
assign v_1253 = v_1251 & v_1252;
assign v_1254 = v_1251 & ~v_1252;
assign v_1257 = v_1255 & v_1256;
assign v_1258 = v_1255 & ~v_1256;
assign v_1261 = v_1259 & ~v_1260;
assign v_1263 = v_1259 & v_1260 & v_1262;
assign v_1264 = v_1259 & v_1260 & ~v_1262;
assign v_1267 = v_1249 & v_1250 & v_1265 & v_1266;
assign v_1269 = v_1249 & ~v_1250 & v_1268;
assign v_1270 = v_1249 & v_1250 & v_1265 & ~v_1266;
assign v_1271 = v_1249 & ~v_1250 & ~v_1268;
assign v_1276 = v_1272 & v_1273 & ~v_1274 & v_1275;
assign v_1278 = v_1272 & ~v_1273 & v_1277;
assign v_1279 = v_1272 & ~v_1273 & ~v_1277;
assign v_1280 = v_1272 & v_1273 & ~v_1274 & ~v_1275;
assign v_1281 = v_1272 & v_1273 & v_1274;
assign v_1283 = v_1202 & v_1282;
assign v_1288 = v_1286 & v_1287;
assign v_1289 = v_1286 & ~v_1287;
assign v_1292 = v_1290 & v_1291;
assign v_1293 = v_1290 & ~v_1291;
assign v_1296 = v_1294 & ~v_1295;
assign v_1298 = v_1294 & v_1295 & v_1297;
assign v_1299 = v_1294 & v_1295 & ~v_1297;
assign v_1302 = v_1284 & v_1285 & v_1300 & v_1301;
assign v_1304 = v_1284 & ~v_1285 & v_1303;
assign v_1305 = v_1284 & v_1285 & v_1300 & ~v_1301;
assign v_1306 = v_1284 & ~v_1285 & ~v_1303;
assign v_1311 = v_1309 & v_1310;
assign v_1312 = v_1309 & ~v_1310;
assign v_1315 = v_1313 & v_1314;
assign v_1316 = v_1313 & ~v_1314;
assign v_1319 = v_1317 & ~v_1318;
assign v_1321 = v_1317 & v_1318 & v_1320;
assign v_1322 = v_1317 & v_1318 & ~v_1320;
assign v_1325 = v_1307 & v_1308 & v_1323 & v_1324;
assign v_1327 = v_1307 & ~v_1308 & v_1326;
assign v_1328 = v_1307 & v_1308 & v_1323 & ~v_1324;
assign v_1329 = v_1307 & ~v_1308 & ~v_1326;
assign v_1334 = v_1332 & v_1333;
assign v_1335 = v_1332 & ~v_1333;
assign v_1338 = v_1336 & v_1337;
assign v_1339 = v_1336 & ~v_1337;
assign v_1342 = v_1340 & ~v_1341;
assign v_1344 = v_1340 & v_1341 & v_1343;
assign v_1345 = v_1340 & v_1341 & ~v_1343;
assign v_1348 = v_1330 & v_1331 & v_1346 & v_1347;
assign v_1350 = v_1330 & ~v_1331 & v_1349;
assign v_1351 = v_1330 & v_1331 & v_1346 & ~v_1347;
assign v_1352 = v_1330 & ~v_1331 & ~v_1349;
assign v_1357 = v_1353 & v_1354 & ~v_1355 & v_1356;
assign v_1359 = v_1353 & ~v_1354 & v_1358;
assign v_1360 = v_1353 & ~v_1354 & ~v_1358;
assign v_1361 = v_1353 & v_1354 & ~v_1355 & ~v_1356;
assign v_1362 = v_1353 & v_1354 & v_1355;
assign v_1364 = v_1283 & v_1363;
assign v_1369 = v_1367 & v_1368;
assign v_1370 = v_1367 & ~v_1368;
assign v_1373 = v_1371 & v_1372;
assign v_1374 = v_1371 & ~v_1372;
assign v_1377 = v_1375 & ~v_1376;
assign v_1379 = v_1375 & v_1376 & v_1378;
assign v_1380 = v_1375 & v_1376 & ~v_1378;
assign v_1383 = v_1365 & v_1366 & v_1381 & v_1382;
assign v_1385 = v_1365 & ~v_1366 & v_1384;
assign v_1386 = v_1365 & v_1366 & v_1381 & ~v_1382;
assign v_1387 = v_1365 & ~v_1366 & ~v_1384;
assign v_1392 = v_1390 & v_1391;
assign v_1393 = v_1390 & ~v_1391;
assign v_1396 = v_1394 & v_1395;
assign v_1397 = v_1394 & ~v_1395;
assign v_1400 = v_1398 & ~v_1399;
assign v_1402 = v_1398 & v_1399 & v_1401;
assign v_1403 = v_1398 & v_1399 & ~v_1401;
assign v_1406 = v_1388 & v_1389 & v_1404 & v_1405;
assign v_1408 = v_1388 & ~v_1389 & v_1407;
assign v_1409 = v_1388 & v_1389 & v_1404 & ~v_1405;
assign v_1410 = v_1388 & ~v_1389 & ~v_1407;
assign v_1415 = v_1413 & v_1414;
assign v_1416 = v_1413 & ~v_1414;
assign v_1419 = v_1417 & v_1418;
assign v_1420 = v_1417 & ~v_1418;
assign v_1423 = v_1421 & ~v_1422;
assign v_1425 = v_1421 & v_1422 & v_1424;
assign v_1426 = v_1421 & v_1422 & ~v_1424;
assign v_1429 = v_1411 & v_1412 & v_1427 & v_1428;
assign v_1431 = v_1411 & ~v_1412 & v_1430;
assign v_1432 = v_1411 & v_1412 & v_1427 & ~v_1428;
assign v_1433 = v_1411 & ~v_1412 & ~v_1430;
assign v_1438 = v_1434 & v_1435 & ~v_1436 & v_1437;
assign v_1440 = v_1434 & ~v_1435 & v_1439;
assign v_1441 = v_1434 & ~v_1435 & ~v_1439;
assign v_1442 = v_1434 & v_1435 & ~v_1436 & ~v_1437;
assign v_1443 = v_1434 & v_1435 & v_1436;
assign v_1445 = v_1364 & v_1444;
assign v_1450 = v_1448 & v_1449;
assign v_1451 = v_1448 & ~v_1449;
assign v_1454 = v_1452 & v_1453;
assign v_1455 = v_1452 & ~v_1453;
assign v_1458 = v_1456 & ~v_1457;
assign v_1460 = v_1456 & v_1457 & v_1459;
assign v_1461 = v_1456 & v_1457 & ~v_1459;
assign v_1464 = v_1446 & v_1447 & v_1462 & v_1463;
assign v_1466 = v_1446 & ~v_1447 & v_1465;
assign v_1467 = v_1446 & v_1447 & v_1462 & ~v_1463;
assign v_1468 = v_1446 & ~v_1447 & ~v_1465;
assign v_1473 = v_1471 & v_1472;
assign v_1474 = v_1471 & ~v_1472;
assign v_1477 = v_1475 & v_1476;
assign v_1478 = v_1475 & ~v_1476;
assign v_1481 = v_1479 & ~v_1480;
assign v_1483 = v_1479 & v_1480 & v_1482;
assign v_1484 = v_1479 & v_1480 & ~v_1482;
assign v_1487 = v_1469 & v_1470 & v_1485 & v_1486;
assign v_1489 = v_1469 & ~v_1470 & v_1488;
assign v_1490 = v_1469 & v_1470 & v_1485 & ~v_1486;
assign v_1491 = v_1469 & ~v_1470 & ~v_1488;
assign v_1496 = v_1494 & v_1495;
assign v_1497 = v_1494 & ~v_1495;
assign v_1500 = v_1498 & v_1499;
assign v_1501 = v_1498 & ~v_1499;
assign v_1504 = v_1502 & ~v_1503;
assign v_1506 = v_1502 & v_1503 & v_1505;
assign v_1507 = v_1502 & v_1503 & ~v_1505;
assign v_1510 = v_1492 & v_1493 & v_1508 & v_1509;
assign v_1512 = v_1492 & ~v_1493 & v_1511;
assign v_1513 = v_1492 & v_1493 & v_1508 & ~v_1509;
assign v_1514 = v_1492 & ~v_1493 & ~v_1511;
assign v_1519 = v_1515 & v_1516 & ~v_1517 & v_1518;
assign v_1521 = v_1515 & ~v_1516 & v_1520;
assign v_1522 = v_1515 & ~v_1516 & ~v_1520;
assign v_1523 = v_1515 & v_1516 & ~v_1517 & ~v_1518;
assign v_1524 = v_1515 & v_1516 & v_1517;
assign v_1526 = v_1445 & v_1525;
assign v_1530 = v_1528 & ~v_1529;
assign v_1532 = v_1527 & v_1531;
assign v_1534 = ~v_227 & v_229 & v_262 & ~v_264;
assign v_1535 = ~v_227 & v_229 & v_262 & v_264;
assign v_1536 = ~v_227 & v_229 & ~v_262;
assign v_1539 = v_1538;
assign v_1541 = v_1540;
assign v_1542 = v_12931 & v_12932;
assign v_1544 = v_1543 & ~v_227 & ~v_229 & v_260;
assign v_1546 = v_1533 & ~v_1545;
assign v_1548 = v_1547 & v_267 & v_268;
assign v_1549 = v_1547 & v_267 & ~v_268;
assign v_1551 = v_1550 & ~v_279;
assign v_1553 = v_1550 & v_1552;
assign v_1554 = v_1550 & v_279 & v_291 & ~v_292 & v_300;
assign v_1557 = v_1555 & v_1556;
assign v_1558 = v_1555 & v_321 & v_322;
assign v_1559 = v_1555 & v_321 & ~v_322 & v_324;
assign v_1560 = v_1555 & v_321 & ~v_322 & ~v_324 & v_326;
assign v_1561 = v_1555 & v_321 & ~v_322 & ~v_324 & ~v_326;
assign v_1564 = v_1562 & v_1563;
assign v_1566 = v_1565 & ~v_308 & v_309 & v_329;
assign v_1569 = v_1567 & v_1568;
assign v_1571 = v_1567 & v_1570;
assign v_1573 = ~v_1527 & v_1572;
assign v_1575 = v_1574 & v_345 & v_346;
assign v_1576 = v_1574 & v_345 & ~v_346 & v_348;
assign v_1577 = v_1574 & v_345 & ~v_346 & ~v_348 & v_350;
assign v_1578 = v_1574 & v_356 & v_357;
assign v_1579 = v_1574 & v_359 & v_360;
assign v_1580 = v_1574 & v_359 & ~v_360 & v_362;
assign v_1581 = v_1574 & v_359 & ~v_360 & ~v_362 & v_364;
assign v_1583 = v_1574 & v_1582;
assign v_1586 = v_1584 & v_1585;
assign v_1588 = v_1587 & v_356 & ~v_357 & v_369 & v_370;
assign v_1589 = v_1587 & v_372 & v_373;
assign v_1590 = v_1587 & v_372 & ~v_373 & v_375;
assign v_1591 = v_1587 & v_372 & ~v_373 & ~v_375 & v_377;
assign v_1593 = v_1587 & v_1592;
assign v_1594 = v_12933 & v_12934;
assign v_1596 = v_1595 & v_384 & v_385;
assign v_1597 = v_1595 & v_384 & ~v_385;
assign v_1600 = v_1598 & v_1599;
assign v_1602 = v_12935 & v_12936;
assign v_1603 = v_1601 & v_391 & v_392;
assign v_1604 = v_1601 & v_391 & ~v_392 & v_394;
assign v_1605 = v_1601 & v_391 & ~v_392 & ~v_394 & v_396;
assign v_1607 = v_1601 & v_1606;
assign v_1609 = v_12937 & v_12938;
assign v_1612 = v_1610 & v_1611;
assign v_1614 = v_1613 & v_410 & v_411;
assign v_1615 = v_1613 & v_410 & ~v_411 & v_413;
assign v_1616 = v_1613 & v_410 & ~v_411 & ~v_413 & v_415;
assign v_1617 = v_1613 & v_421 & v_422;
assign v_1618 = v_1613 & v_424 & v_425;
assign v_1619 = v_1613 & v_424 & ~v_425 & v_427;
assign v_1620 = v_1613 & v_424 & ~v_425 & ~v_427 & v_429;
assign v_1622 = v_1613 & v_1621;
assign v_1625 = v_1623 & v_1624;
assign v_1627 = v_1626 & v_421 & ~v_422 & v_434 & v_435;
assign v_1628 = v_1626 & v_437 & v_438;
assign v_1629 = v_1626 & v_437 & ~v_438 & v_440;
assign v_1630 = v_1626 & v_437 & ~v_438 & ~v_440 & v_442;
assign v_1632 = v_1626 & v_1631;
assign v_1633 = v_12939 & v_12940;
assign v_1635 = v_1634 & v_449 & v_450;
assign v_1636 = v_1634 & v_449 & ~v_450;
assign v_1639 = v_1637 & v_1638;
assign v_1641 = v_12941 & v_12942;
assign v_1642 = v_1640 & v_456 & v_457;
assign v_1643 = v_1640 & v_456 & ~v_457 & v_459;
assign v_1644 = v_1640 & v_456 & ~v_457 & ~v_459 & v_461;
assign v_1646 = v_1640 & v_1645;
assign v_1648 = v_12943 & v_12944;
assign v_1651 = v_1649 & v_1650;
assign v_1653 = v_1652 & v_491;
assign v_1656 = v_1655 & ~v_1652;
assign v_1658 = v_1657 & ~v_491 & v_493 & v_526 & ~v_528;
assign v_1659 = v_1657 & ~v_491 & v_493 & v_526 & v_528;
assign v_1660 = v_1657 & ~v_491 & v_493 & ~v_526;
assign v_1661 = v_1657 & v_494;
assign v_1662 = v_1657 & ~v_494;
assign v_1665 = v_1663 & v_1664;
assign v_1667 = v_1663 & v_1666;
assign v_1668 = v_12945 & v_12946;
assign v_1670 = v_1669 & ~v_491 & ~v_493 & v_524;
assign v_1672 = v_1654 & ~v_1671;
assign v_1674 = v_1673 & v_531 & v_532;
assign v_1675 = v_1673 & v_531 & ~v_532;
assign v_1677 = v_1676 & v_546 & v_547;
assign v_1678 = v_1676 & v_554;
assign v_1680 = v_1679 & v_558 & v_559;
assign v_1681 = v_1679 & v_558 & ~v_559 & v_561;
assign v_1683 = v_1679 & v_1682;
assign v_1686 = v_1684 & v_1685;
assign v_1688 = v_1684 & v_1687;
assign v_1690 = v_1689 & v_588 & ~v_589 & ~v_591;
assign v_1691 = v_1689 & v_593 & ~v_594;
assign v_1692 = v_1689 & v_593 & v_594;
assign v_1693 = v_1689 & v_583;
assign v_1695 = v_1694 & v_604 & v_605;
assign v_1696 = v_1694 & v_612;
assign v_1698 = v_1697 & v_616 & v_617;
assign v_1699 = v_1697 & v_616 & ~v_617 & v_619;
assign v_1701 = v_1697 & v_1700;
assign v_1704 = v_1702 & v_1703;
assign v_1706 = v_1702 & v_1705;
assign v_1708 = v_2 & v_1707;
assign v_1709 = v_641 & v_1689;
assign v_1710 = v_643 & v_1676;
assign v_1711 = v_645 & v_1676;
assign v_1712 = v_647 & v_1676;
assign v_1713 = v_649 & v_1676;
assign v_1714 = ~v_649 & v_1652;
assign v_1716 = ~v_647 & v_1715;
assign v_1718 = ~v_645 & v_1717;
assign v_1720 = ~v_643 & v_1719;
assign v_1722 = ~v_641 & v_1721;
assign v_1724 = ~v_2 & v_1723;
assign v_1726 = v_1725 & ~v_669;
assign v_1727 = v_12947 & v_12948;
assign v_1728 = v_1725 & v_669 & v_670 & v_672 & v_674;
assign v_1729 = v_12949 & v_12950;
assign v_1731 = v_1730 & v_679 & ~v_680 & v_682;
assign v_1732 = v_1730 & v_689 & ~v_690 & ~v_692;
assign v_1733 = v_1730 & v_694 & ~v_695;
assign v_1734 = v_1730 & v_694 & v_695;
assign v_1735 = v_1730 & v_684;
assign v_1738 = v_1736 & v_1737;
assign v_1741 = v_1739 & v_1740;
assign v_1742 = v_1730 & v_679 & v_680;
assign v_1744 = v_1725 & v_1743;
assign v_1746 = v_1745 & ~v_705;
assign v_1747 = v_1745 & v_710 & v_711;
assign v_1748 = v_1745 & v_718;
assign v_1750 = v_1749 & v_705 & v_722 & v_723 & ~v_724;
assign v_1752 = v_1749 & v_1751;
assign v_1753 = v_1749 & v_750 & v_751;
assign v_1754 = v_1749 & v_750 & ~v_751;
assign v_1756 = v_1755 & v_763 & v_764;
assign v_1757 = v_1755 & v_763 & ~v_764;
assign v_1759 = v_1758 & v_745 & v_758 & v_771;
assign v_1760 = v_12951 & v_12952;
assign v_1761 = v_1749 & v_779 & v_780;
assign v_1762 = v_1749 & v_787;
assign v_1765 = v_1763 & v_1764;
assign v_1767 = v_1766 & v_798 & ~v_799 & v_817;
assign v_1768 = v_1766 & v_798 & ~v_799 & ~v_817;
assign v_1769 = v_1766 & ~v_800;
assign v_1770 = v_1766 & v_808 & ~v_809;
assign v_1772 = v_1766 & v_1771;
assign v_1774 = v_1773 & v_798 & v_799 & v_814 & ~v_815;
assign v_1776 = v_1775 & v_821 & ~v_822 & v_840;
assign v_1777 = v_1775 & v_821 & ~v_822 & ~v_840;
assign v_1778 = v_1775 & ~v_823;
assign v_1779 = v_1775 & v_831 & ~v_832;
assign v_1781 = v_1775 & v_1780;
assign v_1783 = v_1782 & v_821 & v_822 & v_837 & ~v_838;
assign v_1785 = v_1784 & v_844 & ~v_845 & v_863;
assign v_1786 = v_1784 & ~v_846;
assign v_1787 = v_1784 & v_854 & ~v_855;
assign v_1789 = v_1784 & v_1788;
assign v_1791 = v_1790 & v_844 & v_845 & v_860 & v_861;
assign v_1792 = v_1784 & v_844 & ~v_845 & ~v_863;
assign v_1793 = v_1790 & v_844 & v_845 & v_860 & ~v_861;
assign v_1796 = v_1794 & v_1795;
assign v_1797 = v_1794 & v_867 & v_868 & ~v_869 & ~v_870;
assign v_1798 = v_1794 & v_867 & v_868 & v_869;
assign v_1799 = v_1794 & v_867 & ~v_868 & ~v_872;
assign v_1802 = v_1800 & v_1801;
assign v_1803 = v_1782 & v_821 & v_822 & v_837 & v_838;
assign v_1804 = v_1773 & v_798 & v_799 & v_814 & v_815;
assign v_1806 = v_1805 & v_879 & ~v_880 & v_898;
assign v_1807 = v_1805 & v_879 & ~v_880 & ~v_898;
assign v_1808 = v_1805 & ~v_881;
assign v_1809 = v_1805 & v_889 & ~v_890;
assign v_1811 = v_1805 & v_1810;
assign v_1813 = v_1812 & v_879 & v_880 & v_895 & ~v_896;
assign v_1815 = v_1814 & v_902 & ~v_903 & v_921;
assign v_1816 = v_1814 & v_902 & ~v_903 & ~v_921;
assign v_1817 = v_1814 & ~v_904;
assign v_1818 = v_1814 & v_912 & ~v_913;
assign v_1820 = v_1814 & v_1819;
assign v_1822 = v_1821 & v_902 & v_903 & v_918 & ~v_919;
assign v_1824 = v_1823 & v_925 & ~v_926 & v_944;
assign v_1825 = v_1823 & ~v_927;
assign v_1826 = v_1823 & v_935 & ~v_936;
assign v_1828 = v_1823 & v_1827;
assign v_1830 = v_1829 & v_925 & v_926 & v_941 & v_942;
assign v_1831 = v_1823 & v_925 & ~v_926 & ~v_944;
assign v_1832 = v_1829 & v_925 & v_926 & v_941 & ~v_942;
assign v_1835 = v_1833 & v_1834;
assign v_1836 = v_1833 & v_948 & v_949 & ~v_950 & ~v_951;
assign v_1837 = v_1833 & v_948 & v_949 & v_950;
assign v_1838 = v_1833 & v_948 & ~v_949 & ~v_953;
assign v_1841 = v_1839 & v_1840;
assign v_1842 = v_1821 & v_902 & v_903 & v_918 & v_919;
assign v_1843 = v_1812 & v_879 & v_880 & v_895 & v_896;
assign v_1845 = v_1844 & v_960 & ~v_961 & v_979;
assign v_1846 = v_1844 & v_960 & ~v_961 & ~v_979;
assign v_1847 = v_1844 & ~v_962;
assign v_1848 = v_1844 & v_970 & ~v_971;
assign v_1850 = v_1844 & v_1849;
assign v_1852 = v_1851 & v_960 & v_961 & v_976 & ~v_977;
assign v_1854 = v_1853 & v_983 & ~v_984 & v_1002;
assign v_1855 = v_1853 & v_983 & ~v_984 & ~v_1002;
assign v_1856 = v_1853 & ~v_985;
assign v_1857 = v_1853 & v_993 & ~v_994;
assign v_1859 = v_1853 & v_1858;
assign v_1861 = v_1860 & v_983 & v_984 & v_999 & ~v_1000;
assign v_1863 = v_1862 & v_1006 & ~v_1007 & v_1025;
assign v_1864 = v_1862 & ~v_1008;
assign v_1865 = v_1862 & v_1016 & ~v_1017;
assign v_1867 = v_1862 & v_1866;
assign v_1869 = v_1868 & v_1006 & v_1007 & v_1022 & v_1023;
assign v_1870 = v_1862 & v_1006 & ~v_1007 & ~v_1025;
assign v_1871 = v_1868 & v_1006 & v_1007 & v_1022 & ~v_1023;
assign v_1874 = v_1872 & v_1873;
assign v_1875 = v_1872 & v_1029 & v_1030 & ~v_1031 & ~v_1032;
assign v_1876 = v_1872 & v_1029 & v_1030 & v_1031;
assign v_1877 = v_1872 & v_1029 & ~v_1030 & ~v_1034;
assign v_1880 = v_1878 & v_1879;
assign v_1881 = v_1860 & v_983 & v_984 & v_999 & v_1000;
assign v_1882 = v_1851 & v_960 & v_961 & v_976 & v_977;
assign v_1884 = v_1883 & v_1041 & ~v_1042 & v_1060;
assign v_1885 = v_1883 & v_1041 & ~v_1042 & ~v_1060;
assign v_1886 = v_1883 & ~v_1043;
assign v_1887 = v_1883 & v_1051 & ~v_1052;
assign v_1889 = v_1883 & v_1888;
assign v_1891 = v_1890 & v_1041 & v_1042 & v_1057 & ~v_1058;
assign v_1893 = v_1892 & v_1064 & ~v_1065 & v_1083;
assign v_1894 = v_1892 & v_1064 & ~v_1065 & ~v_1083;
assign v_1895 = v_1892 & ~v_1066;
assign v_1896 = v_1892 & v_1074 & ~v_1075;
assign v_1898 = v_1892 & v_1897;
assign v_1900 = v_1899 & v_1064 & v_1065 & v_1080 & ~v_1081;
assign v_1902 = v_1901 & v_1087 & ~v_1088 & v_1106;
assign v_1903 = v_1901 & ~v_1089;
assign v_1904 = v_1901 & v_1097 & ~v_1098;
assign v_1906 = v_1901 & v_1905;
assign v_1908 = v_1907 & v_1087 & v_1088 & v_1103 & v_1104;
assign v_1909 = v_1901 & v_1087 & ~v_1088 & ~v_1106;
assign v_1910 = v_1907 & v_1087 & v_1088 & v_1103 & ~v_1104;
assign v_1913 = v_1911 & v_1912;
assign v_1914 = v_1911 & v_1110 & v_1111 & ~v_1112 & ~v_1113;
assign v_1915 = v_1911 & v_1110 & v_1111 & v_1112;
assign v_1916 = v_1911 & v_1110 & ~v_1111 & ~v_1115;
assign v_1919 = v_1917 & v_1918;
assign v_1920 = v_1899 & v_1064 & v_1065 & v_1080 & v_1081;
assign v_1921 = v_1890 & v_1041 & v_1042 & v_1057 & v_1058;
assign v_1923 = v_1922 & v_1122 & ~v_1123 & v_1141;
assign v_1924 = v_1922 & v_1122 & ~v_1123 & ~v_1141;
assign v_1925 = v_1922 & ~v_1124;
assign v_1926 = v_1922 & v_1132 & ~v_1133;
assign v_1928 = v_1922 & v_1927;
assign v_1930 = v_1929 & v_1122 & v_1123 & v_1138 & ~v_1139;
assign v_1932 = v_1931 & v_1145 & ~v_1146 & v_1164;
assign v_1933 = v_1931 & v_1145 & ~v_1146 & ~v_1164;
assign v_1934 = v_1931 & ~v_1147;
assign v_1935 = v_1931 & v_1155 & ~v_1156;
assign v_1937 = v_1931 & v_1936;
assign v_1939 = v_1938 & v_1145 & v_1146 & v_1161 & ~v_1162;
assign v_1941 = v_1940 & v_1168 & ~v_1169 & v_1187;
assign v_1942 = v_1940 & ~v_1170;
assign v_1943 = v_1940 & v_1178 & ~v_1179;
assign v_1945 = v_1940 & v_1944;
assign v_1947 = v_1946 & v_1168 & v_1169 & v_1184 & v_1185;
assign v_1948 = v_1940 & v_1168 & ~v_1169 & ~v_1187;
assign v_1949 = v_1946 & v_1168 & v_1169 & v_1184 & ~v_1185;
assign v_1952 = v_1950 & v_1951;
assign v_1953 = v_1950 & v_1191 & v_1192 & ~v_1193 & ~v_1194;
assign v_1954 = v_1950 & v_1191 & v_1192 & v_1193;
assign v_1955 = v_1950 & v_1191 & ~v_1192 & ~v_1196;
assign v_1958 = v_1956 & v_1957;
assign v_1959 = v_1938 & v_1145 & v_1146 & v_1161 & v_1162;
assign v_1960 = v_1929 & v_1122 & v_1123 & v_1138 & v_1139;
assign v_1962 = v_1961 & v_1203 & ~v_1204 & v_1222;
assign v_1963 = v_1961 & v_1203 & ~v_1204 & ~v_1222;
assign v_1964 = v_1961 & ~v_1205;
assign v_1965 = v_1961 & v_1213 & ~v_1214;
assign v_1967 = v_1961 & v_1966;
assign v_1969 = v_1968 & v_1203 & v_1204 & v_1219 & ~v_1220;
assign v_1971 = v_1970 & v_1226 & ~v_1227 & v_1245;
assign v_1972 = v_1970 & v_1226 & ~v_1227 & ~v_1245;
assign v_1973 = v_1970 & ~v_1228;
assign v_1974 = v_1970 & v_1236 & ~v_1237;
assign v_1976 = v_1970 & v_1975;
assign v_1978 = v_1977 & v_1226 & v_1227 & v_1242 & ~v_1243;
assign v_1980 = v_1979 & v_1249 & ~v_1250 & v_1268;
assign v_1981 = v_1979 & ~v_1251;
assign v_1982 = v_1979 & v_1259 & ~v_1260;
assign v_1984 = v_1979 & v_1983;
assign v_1986 = v_1985 & v_1249 & v_1250 & v_1265 & v_1266;
assign v_1987 = v_1979 & v_1249 & ~v_1250 & ~v_1268;
assign v_1988 = v_1985 & v_1249 & v_1250 & v_1265 & ~v_1266;
assign v_1991 = v_1989 & v_1990;
assign v_1992 = v_1989 & v_1272 & v_1273 & ~v_1274 & ~v_1275;
assign v_1993 = v_1989 & v_1272 & v_1273 & v_1274;
assign v_1994 = v_1989 & v_1272 & ~v_1273 & ~v_1277;
assign v_1997 = v_1995 & v_1996;
assign v_1998 = v_1977 & v_1226 & v_1227 & v_1242 & v_1243;
assign v_1999 = v_1968 & v_1203 & v_1204 & v_1219 & v_1220;
assign v_2001 = v_2000 & v_1284 & ~v_1285 & v_1303;
assign v_2002 = v_2000 & v_1284 & ~v_1285 & ~v_1303;
assign v_2003 = v_2000 & ~v_1286;
assign v_2004 = v_2000 & v_1294 & ~v_1295;
assign v_2006 = v_2000 & v_2005;
assign v_2008 = v_2007 & v_1284 & v_1285 & v_1300 & ~v_1301;
assign v_2010 = v_2009 & v_1307 & ~v_1308 & v_1326;
assign v_2011 = v_2009 & v_1307 & ~v_1308 & ~v_1326;
assign v_2012 = v_2009 & ~v_1309;
assign v_2013 = v_2009 & v_1317 & ~v_1318;
assign v_2015 = v_2009 & v_2014;
assign v_2017 = v_2016 & v_1307 & v_1308 & v_1323 & ~v_1324;
assign v_2019 = v_2018 & v_1330 & ~v_1331 & v_1349;
assign v_2020 = v_2018 & ~v_1332;
assign v_2021 = v_2018 & v_1340 & ~v_1341;
assign v_2023 = v_2018 & v_2022;
assign v_2025 = v_2024 & v_1330 & v_1331 & v_1346 & v_1347;
assign v_2026 = v_2018 & v_1330 & ~v_1331 & ~v_1349;
assign v_2027 = v_2024 & v_1330 & v_1331 & v_1346 & ~v_1347;
assign v_2030 = v_2028 & v_2029;
assign v_2031 = v_2028 & v_1353 & v_1354 & ~v_1355 & ~v_1356;
assign v_2032 = v_2028 & v_1353 & v_1354 & v_1355;
assign v_2033 = v_2028 & v_1353 & ~v_1354 & ~v_1358;
assign v_2036 = v_2034 & v_2035;
assign v_2037 = v_2016 & v_1307 & v_1308 & v_1323 & v_1324;
assign v_2038 = v_2007 & v_1284 & v_1285 & v_1300 & v_1301;
assign v_2040 = v_2039 & v_1365 & ~v_1366 & v_1384;
assign v_2041 = v_2039 & v_1365 & ~v_1366 & ~v_1384;
assign v_2042 = v_2039 & ~v_1367;
assign v_2043 = v_2039 & v_1375 & ~v_1376;
assign v_2045 = v_2039 & v_2044;
assign v_2047 = v_2046 & v_1365 & v_1366 & v_1381 & ~v_1382;
assign v_2049 = v_2048 & v_1388 & ~v_1389 & v_1407;
assign v_2050 = v_2048 & v_1388 & ~v_1389 & ~v_1407;
assign v_2051 = v_2048 & ~v_1390;
assign v_2052 = v_2048 & v_1398 & ~v_1399;
assign v_2054 = v_2048 & v_2053;
assign v_2056 = v_2055 & v_1388 & v_1389 & v_1404 & ~v_1405;
assign v_2058 = v_2057 & v_1411 & ~v_1412 & v_1430;
assign v_2059 = v_2057 & ~v_1413;
assign v_2060 = v_2057 & v_1421 & ~v_1422;
assign v_2062 = v_2057 & v_2061;
assign v_2064 = v_2063 & v_1411 & v_1412 & v_1427 & v_1428;
assign v_2065 = v_2057 & v_1411 & ~v_1412 & ~v_1430;
assign v_2066 = v_2063 & v_1411 & v_1412 & v_1427 & ~v_1428;
assign v_2069 = v_2067 & v_2068;
assign v_2070 = v_2067 & v_1434 & v_1435 & ~v_1436 & ~v_1437;
assign v_2071 = v_2067 & v_1434 & v_1435 & v_1436;
assign v_2072 = v_2067 & v_1434 & ~v_1435 & ~v_1439;
assign v_2075 = v_2073 & v_2074;
assign v_2076 = v_2055 & v_1388 & v_1389 & v_1404 & v_1405;
assign v_2077 = v_2046 & v_1365 & v_1366 & v_1381 & v_1382;
assign v_2079 = v_2078 & v_1446 & ~v_1447 & v_1465;
assign v_2080 = v_2078 & v_1446 & ~v_1447 & ~v_1465;
assign v_2081 = v_2078 & ~v_1448;
assign v_2082 = v_2078 & v_1456 & ~v_1457;
assign v_2084 = v_2078 & v_2083;
assign v_2086 = v_2085 & v_1446 & v_1447 & v_1462 & ~v_1463;
assign v_2088 = v_2087 & v_1469 & ~v_1470 & v_1488;
assign v_2089 = v_2087 & v_1469 & ~v_1470 & ~v_1488;
assign v_2090 = v_2087 & ~v_1471;
assign v_2091 = v_2087 & v_1479 & ~v_1480;
assign v_2093 = v_2087 & v_2092;
assign v_2095 = v_2094 & v_1469 & v_1470 & v_1485 & ~v_1486;
assign v_2097 = v_2096 & v_1492 & ~v_1493 & v_1511;
assign v_2098 = v_2096 & ~v_1494;
assign v_2099 = v_2096 & v_1502 & ~v_1503;
assign v_2101 = v_2096 & v_2100;
assign v_2103 = v_2102 & v_1492 & v_1493 & v_1508 & v_1509;
assign v_2104 = v_2096 & v_1492 & ~v_1493 & ~v_1511;
assign v_2105 = v_2102 & v_1492 & v_1493 & v_1508 & ~v_1509;
assign v_2108 = v_2106 & v_2107;
assign v_2109 = v_2106 & v_1515 & v_1516 & ~v_1517 & ~v_1518;
assign v_2110 = v_2106 & v_1515 & v_1516 & v_1517;
assign v_2111 = v_2106 & v_1515 & ~v_1516 & ~v_1520;
assign v_2114 = v_2112 & v_2113;
assign v_2115 = v_2094 & v_1469 & v_1470 & v_1485 & v_1486;
assign v_2116 = v_2085 & v_1446 & v_1447 & v_1462 & v_1463;
assign v_2120 = v_1527 & v_2119;
assign v_2121 = v_227;
assign v_2124 = v_2123 & v_267 & v_268;
assign v_2125 = v_2123 & v_267 & ~v_268;
assign v_2127 = v_2126 & ~v_279;
assign v_2129 = v_2126 & v_2128;
assign v_2130 = v_2126 & v_279 & v_291 & ~v_292 & v_300;
assign v_2133 = v_2131 & v_2132;
assign v_2134 = v_2131 & v_321 & v_322;
assign v_2135 = v_2131 & v_321 & ~v_322 & v_324;
assign v_2136 = v_2131 & v_321 & ~v_322 & ~v_324 & v_326;
assign v_2137 = v_2131 & v_321 & ~v_322 & ~v_324 & ~v_326;
assign v_2139 = v_2138 & v_1563;
assign v_2141 = v_2140 & ~v_308 & v_309 & v_329;
assign v_2144 = v_2142 & v_2143;
assign v_2145 = v_2142 & v_1570;
assign v_2147 = ~v_1527 & v_2146;
assign v_2149 = v_2148 & v_345 & v_346;
assign v_2150 = v_2148 & v_345 & ~v_346 & v_348;
assign v_2151 = v_2148 & v_345 & ~v_346 & ~v_348 & v_350;
assign v_2152 = v_2148 & v_356 & v_357;
assign v_2153 = v_2148 & v_359 & v_360;
assign v_2154 = v_2148 & v_359 & ~v_360 & v_362;
assign v_2155 = v_2148 & v_359 & ~v_360 & ~v_362 & v_364;
assign v_2156 = v_2148 & v_1582;
assign v_2158 = v_2157 & v_1585;
assign v_2160 = v_2159 & v_356 & ~v_357 & v_369 & v_370;
assign v_2161 = v_2159 & v_372 & v_373;
assign v_2162 = v_2159 & v_372 & ~v_373 & v_375;
assign v_2163 = v_2159 & v_372 & ~v_373 & ~v_375 & v_377;
assign v_2165 = v_2159 & v_2164;
assign v_2166 = v_12953 & v_12954;
assign v_2168 = v_2167 & v_384 & v_385;
assign v_2169 = v_2167 & v_384 & ~v_385;
assign v_2171 = v_2170 & v_1599;
assign v_2173 = v_12955 & v_12956;
assign v_2174 = v_2172 & v_391 & v_392;
assign v_2175 = v_2172 & v_391 & ~v_392 & v_394;
assign v_2176 = v_2172 & v_391 & ~v_392 & ~v_394 & v_396;
assign v_2177 = v_2172 & v_1606;
assign v_2179 = v_12957 & v_12958;
assign v_2181 = v_2180 & v_1611;
assign v_2183 = v_2182 & v_410 & v_411;
assign v_2184 = v_2182 & v_410 & ~v_411 & v_413;
assign v_2185 = v_2182 & v_410 & ~v_411 & ~v_413 & v_415;
assign v_2186 = v_2182 & v_421 & v_422;
assign v_2187 = v_2182 & v_424 & v_425;
assign v_2188 = v_2182 & v_424 & ~v_425 & v_427;
assign v_2189 = v_2182 & v_424 & ~v_425 & ~v_427 & v_429;
assign v_2190 = v_2182 & v_1621;
assign v_2192 = v_2191 & v_1624;
assign v_2194 = v_2193 & v_421 & ~v_422 & v_434 & v_435;
assign v_2195 = v_2193 & v_437 & v_438;
assign v_2196 = v_2193 & v_437 & ~v_438 & v_440;
assign v_2197 = v_2193 & v_437 & ~v_438 & ~v_440 & v_442;
assign v_2199 = v_2193 & v_2198;
assign v_2200 = v_12959 & v_12960;
assign v_2202 = v_2201 & v_449 & v_450;
assign v_2203 = v_2201 & v_449 & ~v_450;
assign v_2205 = v_2204 & v_1638;
assign v_2207 = v_12961 & v_12962;
assign v_2208 = v_2206 & v_456 & v_457;
assign v_2209 = v_2206 & v_456 & ~v_457 & v_459;
assign v_2210 = v_2206 & v_456 & ~v_457 & ~v_459 & v_461;
assign v_2211 = v_2206 & v_1645;
assign v_2213 = v_12963 & v_12964;
assign v_2215 = v_2214 & v_1650;
assign v_2217 = v_2216 & v_491;
assign v_2220 = v_2219 & v_531 & v_532;
assign v_2221 = v_2219 & v_531 & ~v_532;
assign v_2223 = v_2222 & v_546 & v_547;
assign v_2224 = v_2222 & v_554;
assign v_2226 = v_2225 & v_558 & v_559;
assign v_2227 = v_2225 & v_558 & ~v_559 & v_561;
assign v_2228 = v_2225 & v_1682;
assign v_2231 = v_2229 & v_2230;
assign v_2232 = v_2229 & v_1687;
assign v_2234 = v_2233 & v_588 & ~v_589 & ~v_591;
assign v_2235 = v_2233 & v_593 & ~v_594;
assign v_2236 = v_2233 & v_593 & v_594;
assign v_2237 = v_2233 & v_583;
assign v_2239 = v_2238 & v_604 & v_605;
assign v_2240 = v_2238 & v_612;
assign v_2242 = v_2241 & v_616 & v_617;
assign v_2243 = v_2241 & v_616 & ~v_617 & v_619;
assign v_2244 = v_2241 & v_1700;
assign v_2247 = v_2245 & v_2246;
assign v_2248 = v_2245 & v_1705;
assign v_2250 = v_2 & v_2249;
assign v_2251 = v_641 & v_2233;
assign v_2252 = v_643 & v_2222;
assign v_2253 = v_645 & v_2222;
assign v_2254 = v_647 & v_2222;
assign v_2255 = v_649 & v_2222;
assign v_2256 = ~v_649 & v_2216;
assign v_2258 = ~v_647 & v_2257;
assign v_2260 = ~v_645 & v_2259;
assign v_2262 = ~v_643 & v_2261;
assign v_2264 = ~v_641 & v_2263;
assign v_2266 = ~v_2 & v_2265;
assign v_2268 = v_2267 & ~v_669;
assign v_2269 = v_12965 & v_12966;
assign v_2270 = v_2267 & v_669 & v_670 & v_672 & v_674;
assign v_2271 = v_12967 & v_12968;
assign v_2273 = v_2272 & v_679 & ~v_680 & v_682;
assign v_2274 = v_2272 & v_689 & ~v_690 & ~v_692;
assign v_2275 = v_2272 & v_694 & ~v_695;
assign v_2276 = v_2272 & v_694 & v_695;
assign v_2277 = v_2272 & v_684;
assign v_2279 = v_2278 & v_1737;
assign v_2281 = v_2280 & v_1740;
assign v_2282 = v_2272 & v_679 & v_680;
assign v_2283 = v_2267 & v_1743;
assign v_2285 = v_2284 & ~v_705;
assign v_2286 = v_2284 & v_710 & v_711;
assign v_2287 = v_2284 & v_718;
assign v_2289 = v_2288 & v_705 & v_722 & v_723 & ~v_724;
assign v_2291 = v_2288 & v_2290;
assign v_2292 = v_2288 & v_750 & v_751;
assign v_2293 = v_2288 & v_750 & ~v_751;
assign v_2295 = v_2294 & v_763 & v_764;
assign v_2296 = v_2294 & v_763 & ~v_764;
assign v_2298 = v_2297 & v_745 & v_758 & v_771;
assign v_2299 = v_12969 & v_12970;
assign v_2300 = v_2288 & v_779 & v_780;
assign v_2301 = v_2288 & v_787;
assign v_2303 = v_2302 & v_1764;
assign v_2305 = v_2304 & v_798 & ~v_799 & v_817;
assign v_2306 = v_2304 & v_798 & ~v_799 & ~v_817;
assign v_2307 = v_2304 & ~v_800;
assign v_2308 = v_2304 & v_808 & ~v_809;
assign v_2309 = v_2304 & v_1771;
assign v_2311 = v_2310 & v_798 & v_799 & v_814 & ~v_815;
assign v_2313 = v_2312 & v_821 & ~v_822 & v_840;
assign v_2314 = v_2312 & v_821 & ~v_822 & ~v_840;
assign v_2315 = v_2312 & ~v_823;
assign v_2316 = v_2312 & v_831 & ~v_832;
assign v_2317 = v_2312 & v_1780;
assign v_2319 = v_2318 & v_821 & v_822 & v_837 & ~v_838;
assign v_2321 = v_2320 & v_844 & ~v_845 & v_863;
assign v_2322 = v_2320 & ~v_846;
assign v_2323 = v_2320 & v_854 & ~v_855;
assign v_2324 = v_2320 & v_1788;
assign v_2326 = v_2325 & v_844 & v_845 & v_860 & v_861;
assign v_2327 = v_2320 & v_844 & ~v_845 & ~v_863;
assign v_2328 = v_2325 & v_844 & v_845 & v_860 & ~v_861;
assign v_2331 = v_2329 & v_2330;
assign v_2332 = v_2329 & v_867 & v_868 & ~v_869 & ~v_870;
assign v_2333 = v_2329 & v_867 & v_868 & v_869;
assign v_2334 = v_2329 & v_867 & ~v_868 & ~v_872;
assign v_2336 = v_2335 & v_1801;
assign v_2337 = v_2318 & v_821 & v_822 & v_837 & v_838;
assign v_2338 = v_2310 & v_798 & v_799 & v_814 & v_815;
assign v_2340 = v_2339 & v_879 & ~v_880 & v_898;
assign v_2341 = v_2339 & v_879 & ~v_880 & ~v_898;
assign v_2342 = v_2339 & ~v_881;
assign v_2343 = v_2339 & v_889 & ~v_890;
assign v_2344 = v_2339 & v_1810;
assign v_2346 = v_2345 & v_879 & v_880 & v_895 & ~v_896;
assign v_2348 = v_2347 & v_902 & ~v_903 & v_921;
assign v_2349 = v_2347 & v_902 & ~v_903 & ~v_921;
assign v_2350 = v_2347 & ~v_904;
assign v_2351 = v_2347 & v_912 & ~v_913;
assign v_2352 = v_2347 & v_1819;
assign v_2354 = v_2353 & v_902 & v_903 & v_918 & ~v_919;
assign v_2356 = v_2355 & v_925 & ~v_926 & v_944;
assign v_2357 = v_2355 & ~v_927;
assign v_2358 = v_2355 & v_935 & ~v_936;
assign v_2359 = v_2355 & v_1827;
assign v_2361 = v_2360 & v_925 & v_926 & v_941 & v_942;
assign v_2362 = v_2355 & v_925 & ~v_926 & ~v_944;
assign v_2363 = v_2360 & v_925 & v_926 & v_941 & ~v_942;
assign v_2366 = v_2364 & v_2365;
assign v_2367 = v_2364 & v_948 & v_949 & ~v_950 & ~v_951;
assign v_2368 = v_2364 & v_948 & v_949 & v_950;
assign v_2369 = v_2364 & v_948 & ~v_949 & ~v_953;
assign v_2371 = v_2370 & v_1840;
assign v_2372 = v_2353 & v_902 & v_903 & v_918 & v_919;
assign v_2373 = v_2345 & v_879 & v_880 & v_895 & v_896;
assign v_2375 = v_2374 & v_960 & ~v_961 & v_979;
assign v_2376 = v_2374 & v_960 & ~v_961 & ~v_979;
assign v_2377 = v_2374 & ~v_962;
assign v_2378 = v_2374 & v_970 & ~v_971;
assign v_2379 = v_2374 & v_1849;
assign v_2381 = v_2380 & v_960 & v_961 & v_976 & ~v_977;
assign v_2383 = v_2382 & v_983 & ~v_984 & v_1002;
assign v_2384 = v_2382 & v_983 & ~v_984 & ~v_1002;
assign v_2385 = v_2382 & ~v_985;
assign v_2386 = v_2382 & v_993 & ~v_994;
assign v_2387 = v_2382 & v_1858;
assign v_2389 = v_2388 & v_983 & v_984 & v_999 & ~v_1000;
assign v_2391 = v_2390 & v_1006 & ~v_1007 & v_1025;
assign v_2392 = v_2390 & ~v_1008;
assign v_2393 = v_2390 & v_1016 & ~v_1017;
assign v_2394 = v_2390 & v_1866;
assign v_2396 = v_2395 & v_1006 & v_1007 & v_1022 & v_1023;
assign v_2397 = v_2390 & v_1006 & ~v_1007 & ~v_1025;
assign v_2398 = v_2395 & v_1006 & v_1007 & v_1022 & ~v_1023;
assign v_2401 = v_2399 & v_2400;
assign v_2402 = v_2399 & v_1029 & v_1030 & ~v_1031 & ~v_1032;
assign v_2403 = v_2399 & v_1029 & v_1030 & v_1031;
assign v_2404 = v_2399 & v_1029 & ~v_1030 & ~v_1034;
assign v_2406 = v_2405 & v_1879;
assign v_2407 = v_2388 & v_983 & v_984 & v_999 & v_1000;
assign v_2408 = v_2380 & v_960 & v_961 & v_976 & v_977;
assign v_2410 = v_2409 & v_1041 & ~v_1042 & v_1060;
assign v_2411 = v_2409 & v_1041 & ~v_1042 & ~v_1060;
assign v_2412 = v_2409 & ~v_1043;
assign v_2413 = v_2409 & v_1051 & ~v_1052;
assign v_2414 = v_2409 & v_1888;
assign v_2416 = v_2415 & v_1041 & v_1042 & v_1057 & ~v_1058;
assign v_2418 = v_2417 & v_1064 & ~v_1065 & v_1083;
assign v_2419 = v_2417 & v_1064 & ~v_1065 & ~v_1083;
assign v_2420 = v_2417 & ~v_1066;
assign v_2421 = v_2417 & v_1074 & ~v_1075;
assign v_2422 = v_2417 & v_1897;
assign v_2424 = v_2423 & v_1064 & v_1065 & v_1080 & ~v_1081;
assign v_2426 = v_2425 & v_1087 & ~v_1088 & v_1106;
assign v_2427 = v_2425 & ~v_1089;
assign v_2428 = v_2425 & v_1097 & ~v_1098;
assign v_2429 = v_2425 & v_1905;
assign v_2431 = v_2430 & v_1087 & v_1088 & v_1103 & v_1104;
assign v_2432 = v_2425 & v_1087 & ~v_1088 & ~v_1106;
assign v_2433 = v_2430 & v_1087 & v_1088 & v_1103 & ~v_1104;
assign v_2436 = v_2434 & v_2435;
assign v_2437 = v_2434 & v_1110 & v_1111 & ~v_1112 & ~v_1113;
assign v_2438 = v_2434 & v_1110 & v_1111 & v_1112;
assign v_2439 = v_2434 & v_1110 & ~v_1111 & ~v_1115;
assign v_2441 = v_2440 & v_1918;
assign v_2442 = v_2423 & v_1064 & v_1065 & v_1080 & v_1081;
assign v_2443 = v_2415 & v_1041 & v_1042 & v_1057 & v_1058;
assign v_2445 = v_2444 & v_1122 & ~v_1123 & v_1141;
assign v_2446 = v_2444 & v_1122 & ~v_1123 & ~v_1141;
assign v_2447 = v_2444 & ~v_1124;
assign v_2448 = v_2444 & v_1132 & ~v_1133;
assign v_2449 = v_2444 & v_1927;
assign v_2451 = v_2450 & v_1122 & v_1123 & v_1138 & ~v_1139;
assign v_2453 = v_2452 & v_1145 & ~v_1146 & v_1164;
assign v_2454 = v_2452 & v_1145 & ~v_1146 & ~v_1164;
assign v_2455 = v_2452 & ~v_1147;
assign v_2456 = v_2452 & v_1155 & ~v_1156;
assign v_2457 = v_2452 & v_1936;
assign v_2459 = v_2458 & v_1145 & v_1146 & v_1161 & ~v_1162;
assign v_2461 = v_2460 & v_1168 & ~v_1169 & v_1187;
assign v_2462 = v_2460 & ~v_1170;
assign v_2463 = v_2460 & v_1178 & ~v_1179;
assign v_2464 = v_2460 & v_1944;
assign v_2466 = v_2465 & v_1168 & v_1169 & v_1184 & v_1185;
assign v_2467 = v_2460 & v_1168 & ~v_1169 & ~v_1187;
assign v_2468 = v_2465 & v_1168 & v_1169 & v_1184 & ~v_1185;
assign v_2471 = v_2469 & v_2470;
assign v_2472 = v_2469 & v_1191 & v_1192 & ~v_1193 & ~v_1194;
assign v_2473 = v_2469 & v_1191 & v_1192 & v_1193;
assign v_2474 = v_2469 & v_1191 & ~v_1192 & ~v_1196;
assign v_2476 = v_2475 & v_1957;
assign v_2477 = v_2458 & v_1145 & v_1146 & v_1161 & v_1162;
assign v_2478 = v_2450 & v_1122 & v_1123 & v_1138 & v_1139;
assign v_2480 = v_2479 & v_1203 & ~v_1204 & v_1222;
assign v_2481 = v_2479 & v_1203 & ~v_1204 & ~v_1222;
assign v_2482 = v_2479 & ~v_1205;
assign v_2483 = v_2479 & v_1213 & ~v_1214;
assign v_2484 = v_2479 & v_1966;
assign v_2486 = v_2485 & v_1203 & v_1204 & v_1219 & ~v_1220;
assign v_2488 = v_2487 & v_1226 & ~v_1227 & v_1245;
assign v_2489 = v_2487 & v_1226 & ~v_1227 & ~v_1245;
assign v_2490 = v_2487 & ~v_1228;
assign v_2491 = v_2487 & v_1236 & ~v_1237;
assign v_2492 = v_2487 & v_1975;
assign v_2494 = v_2493 & v_1226 & v_1227 & v_1242 & ~v_1243;
assign v_2496 = v_2495 & v_1249 & ~v_1250 & v_1268;
assign v_2497 = v_2495 & ~v_1251;
assign v_2498 = v_2495 & v_1259 & ~v_1260;
assign v_2499 = v_2495 & v_1983;
assign v_2501 = v_2500 & v_1249 & v_1250 & v_1265 & v_1266;
assign v_2502 = v_2495 & v_1249 & ~v_1250 & ~v_1268;
assign v_2503 = v_2500 & v_1249 & v_1250 & v_1265 & ~v_1266;
assign v_2506 = v_2504 & v_2505;
assign v_2507 = v_2504 & v_1272 & v_1273 & ~v_1274 & ~v_1275;
assign v_2508 = v_2504 & v_1272 & v_1273 & v_1274;
assign v_2509 = v_2504 & v_1272 & ~v_1273 & ~v_1277;
assign v_2511 = v_2510 & v_1996;
assign v_2512 = v_2493 & v_1226 & v_1227 & v_1242 & v_1243;
assign v_2513 = v_2485 & v_1203 & v_1204 & v_1219 & v_1220;
assign v_2515 = v_2514 & v_1284 & ~v_1285 & v_1303;
assign v_2516 = v_2514 & v_1284 & ~v_1285 & ~v_1303;
assign v_2517 = v_2514 & ~v_1286;
assign v_2518 = v_2514 & v_1294 & ~v_1295;
assign v_2519 = v_2514 & v_2005;
assign v_2521 = v_2520 & v_1284 & v_1285 & v_1300 & ~v_1301;
assign v_2523 = v_2522 & v_1307 & ~v_1308 & v_1326;
assign v_2524 = v_2522 & v_1307 & ~v_1308 & ~v_1326;
assign v_2525 = v_2522 & ~v_1309;
assign v_2526 = v_2522 & v_1317 & ~v_1318;
assign v_2527 = v_2522 & v_2014;
assign v_2529 = v_2528 & v_1307 & v_1308 & v_1323 & ~v_1324;
assign v_2531 = v_2530 & v_1330 & ~v_1331 & v_1349;
assign v_2532 = v_2530 & ~v_1332;
assign v_2533 = v_2530 & v_1340 & ~v_1341;
assign v_2534 = v_2530 & v_2022;
assign v_2536 = v_2535 & v_1330 & v_1331 & v_1346 & v_1347;
assign v_2537 = v_2530 & v_1330 & ~v_1331 & ~v_1349;
assign v_2538 = v_2535 & v_1330 & v_1331 & v_1346 & ~v_1347;
assign v_2541 = v_2539 & v_2540;
assign v_2542 = v_2539 & v_1353 & v_1354 & ~v_1355 & ~v_1356;
assign v_2543 = v_2539 & v_1353 & v_1354 & v_1355;
assign v_2544 = v_2539 & v_1353 & ~v_1354 & ~v_1358;
assign v_2546 = v_2545 & v_2035;
assign v_2547 = v_2528 & v_1307 & v_1308 & v_1323 & v_1324;
assign v_2548 = v_2520 & v_1284 & v_1285 & v_1300 & v_1301;
assign v_2550 = v_2549 & v_1365 & ~v_1366 & v_1384;
assign v_2551 = v_2549 & v_1365 & ~v_1366 & ~v_1384;
assign v_2552 = v_2549 & ~v_1367;
assign v_2553 = v_2549 & v_1375 & ~v_1376;
assign v_2554 = v_2549 & v_2044;
assign v_2556 = v_2555 & v_1365 & v_1366 & v_1381 & ~v_1382;
assign v_2558 = v_2557 & v_1388 & ~v_1389 & v_1407;
assign v_2559 = v_2557 & v_1388 & ~v_1389 & ~v_1407;
assign v_2560 = v_2557 & ~v_1390;
assign v_2561 = v_2557 & v_1398 & ~v_1399;
assign v_2562 = v_2557 & v_2053;
assign v_2564 = v_2563 & v_1388 & v_1389 & v_1404 & ~v_1405;
assign v_2566 = v_2565 & v_1411 & ~v_1412 & v_1430;
assign v_2567 = v_2565 & ~v_1413;
assign v_2568 = v_2565 & v_1421 & ~v_1422;
assign v_2569 = v_2565 & v_2061;
assign v_2571 = v_2570 & v_1411 & v_1412 & v_1427 & v_1428;
assign v_2572 = v_2565 & v_1411 & ~v_1412 & ~v_1430;
assign v_2573 = v_2570 & v_1411 & v_1412 & v_1427 & ~v_1428;
assign v_2576 = v_2574 & v_2575;
assign v_2577 = v_2574 & v_1434 & v_1435 & ~v_1436 & ~v_1437;
assign v_2578 = v_2574 & v_1434 & v_1435 & v_1436;
assign v_2579 = v_2574 & v_1434 & ~v_1435 & ~v_1439;
assign v_2581 = v_2580 & v_2074;
assign v_2582 = v_2563 & v_1388 & v_1389 & v_1404 & v_1405;
assign v_2583 = v_2555 & v_1365 & v_1366 & v_1381 & v_1382;
assign v_2585 = v_2584 & v_1446 & ~v_1447 & v_1465;
assign v_2586 = v_2584 & v_1446 & ~v_1447 & ~v_1465;
assign v_2587 = v_2584 & ~v_1448;
assign v_2588 = v_2584 & v_1456 & ~v_1457;
assign v_2589 = v_2584 & v_2083;
assign v_2591 = v_2590 & v_1446 & v_1447 & v_1462 & ~v_1463;
assign v_2593 = v_2592 & v_1469 & ~v_1470 & v_1488;
assign v_2594 = v_2592 & v_1469 & ~v_1470 & ~v_1488;
assign v_2595 = v_2592 & ~v_1471;
assign v_2596 = v_2592 & v_1479 & ~v_1480;
assign v_2597 = v_2592 & v_2092;
assign v_2599 = v_2598 & v_1469 & v_1470 & v_1485 & ~v_1486;
assign v_2601 = v_2600 & v_1492 & ~v_1493 & v_1511;
assign v_2602 = v_2600 & ~v_1494;
assign v_2603 = v_2600 & v_1502 & ~v_1503;
assign v_2604 = v_2600 & v_2100;
assign v_2606 = v_2605 & v_1492 & v_1493 & v_1508 & v_1509;
assign v_2607 = v_2600 & v_1492 & ~v_1493 & ~v_1511;
assign v_2608 = v_2605 & v_1492 & v_1493 & v_1508 & ~v_1509;
assign v_2611 = v_2609 & v_2610;
assign v_2612 = v_2609 & v_1515 & v_1516 & ~v_1517 & ~v_1518;
assign v_2613 = v_2609 & v_1515 & v_1516 & v_1517;
assign v_2614 = v_2609 & v_1515 & ~v_1516 & ~v_1520;
assign v_2616 = v_2615 & v_2113;
assign v_2617 = v_2598 & v_1469 & v_1470 & v_1485 & v_1486;
assign v_2618 = v_2590 & v_1446 & v_1447 & v_1462 & v_1463;
assign v_2620 = v_8 & v_227;
assign v_2621 = v_8 & ~v_227 & v_229 & v_262 & ~v_264;
assign v_2622 = v_8 & ~v_227 & v_229 & v_262 & v_264;
assign v_2623 = v_8 & ~v_227 & v_229 & ~v_262;
assign v_2624 = v_8 & v_230;
assign v_2625 = v_8 & ~v_230;
assign v_2628 = v_2626 & v_2627;
assign v_2629 = v_2626 & v_1540;
assign v_2630 = v_12971 & v_12972;
assign v_2632 = v_2631 & ~v_227 & ~v_229 & v_260;
assign v_2634 = v_2633 & v_267 & v_268;
assign v_2635 = v_2633 & v_267 & ~v_268;
assign v_2637 = v_2636 & ~v_279;
assign v_2639 = v_2636 & v_2638;
assign v_2640 = v_2636 & v_279 & v_291 & ~v_292 & v_300;
assign v_2643 = v_2641 & v_2642;
assign v_2644 = v_2641 & v_321 & v_322;
assign v_2645 = v_2641 & v_321 & ~v_322 & v_324;
assign v_2646 = v_2641 & v_321 & ~v_322 & ~v_324 & v_326;
assign v_2647 = v_2641 & v_321 & ~v_322 & ~v_324 & ~v_326;
assign v_2649 = v_2648 & v_1563;
assign v_2651 = v_2650 & ~v_308 & v_309 & v_329;
assign v_2654 = v_2652 & v_2653;
assign v_2655 = v_2652 & v_1570;
assign v_2657 = v_2656 & v_345 & v_346;
assign v_2658 = v_2656 & v_345 & ~v_346 & v_348;
assign v_2659 = v_2656 & v_345 & ~v_346 & ~v_348 & v_350;
assign v_2660 = v_2656 & v_356 & v_357;
assign v_2661 = v_2656 & v_359 & v_360;
assign v_2662 = v_2656 & v_359 & ~v_360 & v_362;
assign v_2663 = v_2656 & v_359 & ~v_360 & ~v_362 & v_364;
assign v_2664 = v_2656 & v_1582;
assign v_2666 = v_2665 & v_1585;
assign v_2668 = v_2667 & v_356 & ~v_357 & v_369 & v_370;
assign v_2669 = v_2667 & v_372 & v_373;
assign v_2670 = v_2667 & v_372 & ~v_373 & v_375;
assign v_2671 = v_2667 & v_372 & ~v_373 & ~v_375 & v_377;
assign v_2673 = v_2667 & v_2672;
assign v_2674 = v_12973 & v_12974;
assign v_2676 = v_2675 & v_384 & v_385;
assign v_2677 = v_2675 & v_384 & ~v_385;
assign v_2679 = v_2678 & v_1599;
assign v_2681 = v_12975 & v_12976;
assign v_2682 = v_2680 & v_391 & v_392;
assign v_2683 = v_2680 & v_391 & ~v_392 & v_394;
assign v_2684 = v_2680 & v_391 & ~v_392 & ~v_394 & v_396;
assign v_2685 = v_2680 & v_1606;
assign v_2687 = v_12977 & v_12978;
assign v_2689 = v_2688 & v_1611;
assign v_2691 = v_2690 & v_410 & v_411;
assign v_2692 = v_2690 & v_410 & ~v_411 & v_413;
assign v_2693 = v_2690 & v_410 & ~v_411 & ~v_413 & v_415;
assign v_2694 = v_2690 & v_421 & v_422;
assign v_2695 = v_2690 & v_424 & v_425;
assign v_2696 = v_2690 & v_424 & ~v_425 & v_427;
assign v_2697 = v_2690 & v_424 & ~v_425 & ~v_427 & v_429;
assign v_2698 = v_2690 & v_1621;
assign v_2700 = v_2699 & v_1624;
assign v_2702 = v_2701 & v_421 & ~v_422 & v_434 & v_435;
assign v_2703 = v_2701 & v_437 & v_438;
assign v_2704 = v_2701 & v_437 & ~v_438 & v_440;
assign v_2705 = v_2701 & v_437 & ~v_438 & ~v_440 & v_442;
assign v_2707 = v_2701 & v_2706;
assign v_2708 = v_12979 & v_12980;
assign v_2710 = v_2709 & v_449 & v_450;
assign v_2711 = v_2709 & v_449 & ~v_450;
assign v_2713 = v_2712 & v_1638;
assign v_2715 = v_12981 & v_12982;
assign v_2716 = v_2714 & v_456 & v_457;
assign v_2717 = v_2714 & v_456 & ~v_457 & v_459;
assign v_2718 = v_2714 & v_456 & ~v_457 & ~v_459 & v_461;
assign v_2719 = v_2714 & v_1645;
assign v_2721 = v_12983 & v_12984;
assign v_2723 = v_2722 & v_1650;
assign v_2725 = v_2724 & v_491;
assign v_2726 = v_2724 & ~v_491 & v_493 & v_526 & ~v_528;
assign v_2727 = v_2724 & ~v_491 & v_493 & v_526 & v_528;
assign v_2728 = v_2724 & ~v_491 & v_493 & ~v_526;
assign v_2729 = v_2724 & v_494;
assign v_2730 = v_2724 & ~v_494;
assign v_2733 = v_2731 & v_2732;
assign v_2734 = v_2731 & v_1666;
assign v_2735 = v_12985 & v_12986;
assign v_2737 = v_2736 & ~v_491 & ~v_493 & v_524;
assign v_2739 = v_2738 & v_531 & v_532;
assign v_2740 = v_2738 & v_531 & ~v_532;
assign v_2742 = v_2741 & v_546 & v_547;
assign v_2743 = v_2741 & v_546 & ~v_547 & ~v_551;
assign v_2745 = v_2744 & v_546 & ~v_547 & v_551;
assign v_2747 = v_2746 & v_554;
assign v_2749 = v_2748 & v_558 & v_559;
assign v_2750 = v_2748 & v_558 & ~v_559 & v_561;
assign v_2751 = v_2748 & v_1682;
assign v_2754 = v_2752 & v_2753;
assign v_2755 = v_2752 & v_1687;
assign v_2757 = v_2756 & v_588 & ~v_589 & ~v_591;
assign v_2758 = v_2756 & v_593 & ~v_594;
assign v_2759 = v_2756 & v_593 & v_594;
assign v_2760 = v_2756 & v_583;
assign v_2762 = v_2761 & v_604 & v_605;
assign v_2763 = v_2761 & v_604 & ~v_605 & ~v_609;
assign v_2765 = v_2764 & v_604 & ~v_605 & v_609;
assign v_2767 = v_2766 & v_612;
assign v_2769 = v_2768 & v_616 & v_617;
assign v_2770 = v_2768 & v_616 & ~v_617 & v_619;
assign v_2771 = v_2768 & v_1700;
assign v_2774 = v_2772 & v_2773;
assign v_2775 = v_2772 & v_1705;
assign v_2777 = v_2 & v_2776;
assign v_2778 = v_641 & v_2756;
assign v_2779 = v_643 & v_2741;
assign v_2780 = v_645 & v_2741;
assign v_2781 = v_647 & v_2741;
assign v_2782 = v_649 & v_2741;
assign v_2783 = ~v_649 & v_2724;
assign v_2785 = ~v_647 & v_2784;
assign v_2787 = ~v_645 & v_2786;
assign v_2789 = ~v_643 & v_2788;
assign v_2791 = ~v_641 & v_2790;
assign v_2793 = ~v_2 & v_2792;
assign v_2795 = v_2794 & ~v_669;
assign v_2796 = v_12987 & v_12988;
assign v_2797 = v_2794 & v_669 & v_670 & v_672 & v_674;
assign v_2798 = v_12989 & v_12990;
assign v_2800 = v_2799 & v_679 & ~v_680 & v_682;
assign v_2801 = v_2799 & v_689 & ~v_690 & ~v_692;
assign v_2802 = v_2799 & v_694 & ~v_695;
assign v_2803 = v_2799 & v_694 & v_695;
assign v_2804 = v_2799 & v_684;
assign v_2806 = v_2805 & v_1737;
assign v_2808 = v_2807 & v_1740;
assign v_2809 = v_2799 & v_679 & v_680;
assign v_2810 = v_2794 & v_1743;
assign v_2812 = v_2811 & ~v_705;
assign v_2813 = v_2811 & v_710 & v_711;
assign v_2814 = v_2811 & v_710 & ~v_711 & ~v_715;
assign v_2816 = v_2815 & v_710 & ~v_711 & v_715;
assign v_2818 = v_2817 & v_718;
assign v_2820 = v_2819 & v_705 & v_722 & v_723 & ~v_724;
assign v_2822 = v_2819 & v_2821;
assign v_2823 = v_2819 & v_750 & v_751;
assign v_2824 = v_2819 & v_750 & ~v_751;
assign v_2826 = v_2825 & v_763 & v_764;
assign v_2827 = v_2825 & v_763 & ~v_764;
assign v_2829 = v_2828 & v_745 & v_758 & v_771;
assign v_2830 = v_12991 & v_12992;
assign v_2831 = v_2819 & v_779 & v_780;
assign v_2832 = v_2819 & v_779 & ~v_780 & ~v_784;
assign v_2834 = v_2833 & v_779 & ~v_780 & v_784;
assign v_2836 = v_2835 & v_787;
assign v_2838 = v_2837 & v_1764;
assign v_2840 = v_2839 & v_798 & ~v_799 & v_817;
assign v_2841 = v_2839 & v_798 & ~v_799 & ~v_817;
assign v_2842 = v_2839 & ~v_800;
assign v_2843 = v_2839 & v_808 & ~v_809;
assign v_2844 = v_2839 & v_1771;
assign v_2846 = v_2845 & v_798 & v_799 & v_814 & ~v_815;
assign v_2848 = v_2847 & v_821 & ~v_822 & v_840;
assign v_2849 = v_2847 & v_821 & ~v_822 & ~v_840;
assign v_2850 = v_2847 & ~v_823;
assign v_2851 = v_2847 & v_831 & ~v_832;
assign v_2852 = v_2847 & v_1780;
assign v_2854 = v_2853 & v_821 & v_822 & v_837 & ~v_838;
assign v_2856 = v_2855 & v_844 & ~v_845 & v_863;
assign v_2857 = v_2855 & ~v_846;
assign v_2858 = v_2855 & v_854 & ~v_855;
assign v_2859 = v_2855 & v_1788;
assign v_2861 = v_2860 & v_844 & v_845 & v_860 & v_861;
assign v_2862 = v_2855 & v_844 & ~v_845 & ~v_863;
assign v_2863 = v_2860 & v_844 & v_845 & v_860 & ~v_861;
assign v_2866 = v_2864 & v_2865;
assign v_2867 = v_2864 & v_867 & v_868 & ~v_869 & ~v_870;
assign v_2868 = v_2864 & v_867 & v_868 & v_869;
assign v_2869 = v_2864 & v_867 & ~v_868 & ~v_872;
assign v_2871 = v_2870 & v_1801;
assign v_2872 = v_2853 & v_821 & v_822 & v_837 & v_838;
assign v_2873 = v_2845 & v_798 & v_799 & v_814 & v_815;
assign v_2875 = v_2874 & v_879 & ~v_880 & v_898;
assign v_2876 = v_2874 & v_879 & ~v_880 & ~v_898;
assign v_2877 = v_2874 & ~v_881;
assign v_2878 = v_2874 & v_889 & ~v_890;
assign v_2879 = v_2874 & v_1810;
assign v_2881 = v_2880 & v_879 & v_880 & v_895 & ~v_896;
assign v_2883 = v_2882 & v_902 & ~v_903 & v_921;
assign v_2884 = v_2882 & v_902 & ~v_903 & ~v_921;
assign v_2885 = v_2882 & ~v_904;
assign v_2886 = v_2882 & v_912 & ~v_913;
assign v_2887 = v_2882 & v_1819;
assign v_2889 = v_2888 & v_902 & v_903 & v_918 & ~v_919;
assign v_2891 = v_2890 & v_925 & ~v_926 & v_944;
assign v_2892 = v_2890 & ~v_927;
assign v_2893 = v_2890 & v_935 & ~v_936;
assign v_2894 = v_2890 & v_1827;
assign v_2896 = v_2895 & v_925 & v_926 & v_941 & v_942;
assign v_2897 = v_2890 & v_925 & ~v_926 & ~v_944;
assign v_2898 = v_2895 & v_925 & v_926 & v_941 & ~v_942;
assign v_2901 = v_2899 & v_2900;
assign v_2902 = v_2899 & v_948 & v_949 & ~v_950 & ~v_951;
assign v_2903 = v_2899 & v_948 & v_949 & v_950;
assign v_2904 = v_2899 & v_948 & ~v_949 & ~v_953;
assign v_2906 = v_2905 & v_1840;
assign v_2907 = v_2888 & v_902 & v_903 & v_918 & v_919;
assign v_2908 = v_2880 & v_879 & v_880 & v_895 & v_896;
assign v_2910 = v_2909 & v_960 & ~v_961 & v_979;
assign v_2911 = v_2909 & v_960 & ~v_961 & ~v_979;
assign v_2912 = v_2909 & ~v_962;
assign v_2913 = v_2909 & v_970 & ~v_971;
assign v_2914 = v_2909 & v_1849;
assign v_2916 = v_2915 & v_960 & v_961 & v_976 & ~v_977;
assign v_2918 = v_2917 & v_983 & ~v_984 & v_1002;
assign v_2919 = v_2917 & v_983 & ~v_984 & ~v_1002;
assign v_2920 = v_2917 & ~v_985;
assign v_2921 = v_2917 & v_993 & ~v_994;
assign v_2922 = v_2917 & v_1858;
assign v_2924 = v_2923 & v_983 & v_984 & v_999 & ~v_1000;
assign v_2926 = v_2925 & v_1006 & ~v_1007 & v_1025;
assign v_2927 = v_2925 & ~v_1008;
assign v_2928 = v_2925 & v_1016 & ~v_1017;
assign v_2929 = v_2925 & v_1866;
assign v_2931 = v_2930 & v_1006 & v_1007 & v_1022 & v_1023;
assign v_2932 = v_2925 & v_1006 & ~v_1007 & ~v_1025;
assign v_2933 = v_2930 & v_1006 & v_1007 & v_1022 & ~v_1023;
assign v_2936 = v_2934 & v_2935;
assign v_2937 = v_2934 & v_1029 & v_1030 & ~v_1031 & ~v_1032;
assign v_2938 = v_2934 & v_1029 & v_1030 & v_1031;
assign v_2939 = v_2934 & v_1029 & ~v_1030 & ~v_1034;
assign v_2941 = v_2940 & v_1879;
assign v_2942 = v_2923 & v_983 & v_984 & v_999 & v_1000;
assign v_2943 = v_2915 & v_960 & v_961 & v_976 & v_977;
assign v_2945 = v_2944 & v_1041 & ~v_1042 & v_1060;
assign v_2946 = v_2944 & v_1041 & ~v_1042 & ~v_1060;
assign v_2947 = v_2944 & ~v_1043;
assign v_2948 = v_2944 & v_1051 & ~v_1052;
assign v_2949 = v_2944 & v_1888;
assign v_2951 = v_2950 & v_1041 & v_1042 & v_1057 & ~v_1058;
assign v_2953 = v_2952 & v_1064 & ~v_1065 & v_1083;
assign v_2954 = v_2952 & v_1064 & ~v_1065 & ~v_1083;
assign v_2955 = v_2952 & ~v_1066;
assign v_2956 = v_2952 & v_1074 & ~v_1075;
assign v_2957 = v_2952 & v_1897;
assign v_2959 = v_2958 & v_1064 & v_1065 & v_1080 & ~v_1081;
assign v_2961 = v_2960 & v_1087 & ~v_1088 & v_1106;
assign v_2962 = v_2960 & ~v_1089;
assign v_2963 = v_2960 & v_1097 & ~v_1098;
assign v_2964 = v_2960 & v_1905;
assign v_2966 = v_2965 & v_1087 & v_1088 & v_1103 & v_1104;
assign v_2967 = v_2960 & v_1087 & ~v_1088 & ~v_1106;
assign v_2968 = v_2965 & v_1087 & v_1088 & v_1103 & ~v_1104;
assign v_2971 = v_2969 & v_2970;
assign v_2972 = v_2969 & v_1110 & v_1111 & ~v_1112 & ~v_1113;
assign v_2973 = v_2969 & v_1110 & v_1111 & v_1112;
assign v_2974 = v_2969 & v_1110 & ~v_1111 & ~v_1115;
assign v_2976 = v_2975 & v_1918;
assign v_2977 = v_2958 & v_1064 & v_1065 & v_1080 & v_1081;
assign v_2978 = v_2950 & v_1041 & v_1042 & v_1057 & v_1058;
assign v_2980 = v_2979 & v_1122 & ~v_1123 & v_1141;
assign v_2981 = v_2979 & v_1122 & ~v_1123 & ~v_1141;
assign v_2982 = v_2979 & ~v_1124;
assign v_2983 = v_2979 & v_1132 & ~v_1133;
assign v_2984 = v_2979 & v_1927;
assign v_2986 = v_2985 & v_1122 & v_1123 & v_1138 & ~v_1139;
assign v_2988 = v_2987 & v_1145 & ~v_1146 & v_1164;
assign v_2989 = v_2987 & v_1145 & ~v_1146 & ~v_1164;
assign v_2990 = v_2987 & ~v_1147;
assign v_2991 = v_2987 & v_1155 & ~v_1156;
assign v_2992 = v_2987 & v_1936;
assign v_2994 = v_2993 & v_1145 & v_1146 & v_1161 & ~v_1162;
assign v_2996 = v_2995 & v_1168 & ~v_1169 & v_1187;
assign v_2997 = v_2995 & ~v_1170;
assign v_2998 = v_2995 & v_1178 & ~v_1179;
assign v_2999 = v_2995 & v_1944;
assign v_3001 = v_3000 & v_1168 & v_1169 & v_1184 & v_1185;
assign v_3002 = v_2995 & v_1168 & ~v_1169 & ~v_1187;
assign v_3003 = v_3000 & v_1168 & v_1169 & v_1184 & ~v_1185;
assign v_3006 = v_3004 & v_3005;
assign v_3007 = v_3004 & v_1191 & v_1192 & ~v_1193 & ~v_1194;
assign v_3008 = v_3004 & v_1191 & v_1192 & v_1193;
assign v_3009 = v_3004 & v_1191 & ~v_1192 & ~v_1196;
assign v_3011 = v_3010 & v_1957;
assign v_3012 = v_2993 & v_1145 & v_1146 & v_1161 & v_1162;
assign v_3013 = v_2985 & v_1122 & v_1123 & v_1138 & v_1139;
assign v_3015 = v_3014 & v_1203 & ~v_1204 & v_1222;
assign v_3016 = v_3014 & v_1203 & ~v_1204 & ~v_1222;
assign v_3017 = v_3014 & ~v_1205;
assign v_3018 = v_3014 & v_1213 & ~v_1214;
assign v_3019 = v_3014 & v_1966;
assign v_3021 = v_3020 & v_1203 & v_1204 & v_1219 & ~v_1220;
assign v_3023 = v_3022 & v_1226 & ~v_1227 & v_1245;
assign v_3024 = v_3022 & v_1226 & ~v_1227 & ~v_1245;
assign v_3025 = v_3022 & ~v_1228;
assign v_3026 = v_3022 & v_1236 & ~v_1237;
assign v_3027 = v_3022 & v_1975;
assign v_3029 = v_3028 & v_1226 & v_1227 & v_1242 & ~v_1243;
assign v_3031 = v_3030 & v_1249 & ~v_1250 & v_1268;
assign v_3032 = v_3030 & ~v_1251;
assign v_3033 = v_3030 & v_1259 & ~v_1260;
assign v_3034 = v_3030 & v_1983;
assign v_3036 = v_3035 & v_1249 & v_1250 & v_1265 & v_1266;
assign v_3037 = v_3030 & v_1249 & ~v_1250 & ~v_1268;
assign v_3038 = v_3035 & v_1249 & v_1250 & v_1265 & ~v_1266;
assign v_3041 = v_3039 & v_3040;
assign v_3042 = v_3039 & v_1272 & v_1273 & ~v_1274 & ~v_1275;
assign v_3043 = v_3039 & v_1272 & v_1273 & v_1274;
assign v_3044 = v_3039 & v_1272 & ~v_1273 & ~v_1277;
assign v_3046 = v_3045 & v_1996;
assign v_3047 = v_3028 & v_1226 & v_1227 & v_1242 & v_1243;
assign v_3048 = v_3020 & v_1203 & v_1204 & v_1219 & v_1220;
assign v_3050 = v_3049 & v_1284 & ~v_1285 & v_1303;
assign v_3051 = v_3049 & v_1284 & ~v_1285 & ~v_1303;
assign v_3052 = v_3049 & ~v_1286;
assign v_3053 = v_3049 & v_1294 & ~v_1295;
assign v_3054 = v_3049 & v_2005;
assign v_3056 = v_3055 & v_1284 & v_1285 & v_1300 & ~v_1301;
assign v_3058 = v_3057 & v_1307 & ~v_1308 & v_1326;
assign v_3059 = v_3057 & v_1307 & ~v_1308 & ~v_1326;
assign v_3060 = v_3057 & ~v_1309;
assign v_3061 = v_3057 & v_1317 & ~v_1318;
assign v_3062 = v_3057 & v_2014;
assign v_3064 = v_3063 & v_1307 & v_1308 & v_1323 & ~v_1324;
assign v_3066 = v_3065 & v_1330 & ~v_1331 & v_1349;
assign v_3067 = v_3065 & ~v_1332;
assign v_3068 = v_3065 & v_1340 & ~v_1341;
assign v_3069 = v_3065 & v_2022;
assign v_3071 = v_3070 & v_1330 & v_1331 & v_1346 & v_1347;
assign v_3072 = v_3065 & v_1330 & ~v_1331 & ~v_1349;
assign v_3073 = v_3070 & v_1330 & v_1331 & v_1346 & ~v_1347;
assign v_3076 = v_3074 & v_3075;
assign v_3077 = v_3074 & v_1353 & v_1354 & ~v_1355 & ~v_1356;
assign v_3078 = v_3074 & v_1353 & v_1354 & v_1355;
assign v_3079 = v_3074 & v_1353 & ~v_1354 & ~v_1358;
assign v_3081 = v_3080 & v_2035;
assign v_3082 = v_3063 & v_1307 & v_1308 & v_1323 & v_1324;
assign v_3083 = v_3055 & v_1284 & v_1285 & v_1300 & v_1301;
assign v_3085 = v_3084 & v_1365 & ~v_1366 & v_1384;
assign v_3086 = v_3084 & v_1365 & ~v_1366 & ~v_1384;
assign v_3087 = v_3084 & ~v_1367;
assign v_3088 = v_3084 & v_1375 & ~v_1376;
assign v_3089 = v_3084 & v_2044;
assign v_3091 = v_3090 & v_1365 & v_1366 & v_1381 & ~v_1382;
assign v_3093 = v_3092 & v_1388 & ~v_1389 & v_1407;
assign v_3094 = v_3092 & v_1388 & ~v_1389 & ~v_1407;
assign v_3095 = v_3092 & ~v_1390;
assign v_3096 = v_3092 & v_1398 & ~v_1399;
assign v_3097 = v_3092 & v_2053;
assign v_3099 = v_3098 & v_1388 & v_1389 & v_1404 & ~v_1405;
assign v_3101 = v_3100 & v_1411 & ~v_1412 & v_1430;
assign v_3102 = v_3100 & ~v_1413;
assign v_3103 = v_3100 & v_1421 & ~v_1422;
assign v_3104 = v_3100 & v_2061;
assign v_3106 = v_3105 & v_1411 & v_1412 & v_1427 & v_1428;
assign v_3107 = v_3100 & v_1411 & ~v_1412 & ~v_1430;
assign v_3108 = v_3105 & v_1411 & v_1412 & v_1427 & ~v_1428;
assign v_3111 = v_3109 & v_3110;
assign v_3112 = v_3109 & v_1434 & v_1435 & ~v_1436 & ~v_1437;
assign v_3113 = v_3109 & v_1434 & v_1435 & v_1436;
assign v_3114 = v_3109 & v_1434 & ~v_1435 & ~v_1439;
assign v_3116 = v_3115 & v_2074;
assign v_3117 = v_3098 & v_1388 & v_1389 & v_1404 & v_1405;
assign v_3118 = v_3090 & v_1365 & v_1366 & v_1381 & v_1382;
assign v_3120 = v_3119 & v_1446 & ~v_1447 & v_1465;
assign v_3121 = v_3119 & v_1446 & ~v_1447 & ~v_1465;
assign v_3122 = v_3119 & ~v_1448;
assign v_3123 = v_3119 & v_1456 & ~v_1457;
assign v_3124 = v_3119 & v_2083;
assign v_3126 = v_3125 & v_1446 & v_1447 & v_1462 & ~v_1463;
assign v_3128 = v_3127 & v_1469 & ~v_1470 & v_1488;
assign v_3129 = v_3127 & v_1469 & ~v_1470 & ~v_1488;
assign v_3130 = v_3127 & ~v_1471;
assign v_3131 = v_3127 & v_1479 & ~v_1480;
assign v_3132 = v_3127 & v_2092;
assign v_3134 = v_3133 & v_1469 & v_1470 & v_1485 & ~v_1486;
assign v_3136 = v_3135 & v_1492 & ~v_1493 & v_1511;
assign v_3137 = v_3135 & ~v_1494;
assign v_3138 = v_3135 & v_1502 & ~v_1503;
assign v_3139 = v_3135 & v_2100;
assign v_3141 = v_3140 & v_1492 & v_1493 & v_1508 & v_1509;
assign v_3142 = v_3135 & v_1492 & ~v_1493 & ~v_1511;
assign v_3143 = v_3140 & v_1492 & v_1493 & v_1508 & ~v_1509;
assign v_3146 = v_3144 & v_3145;
assign v_3147 = v_3144 & v_1515 & v_1516 & ~v_1517 & ~v_1518;
assign v_3148 = v_3144 & v_1515 & v_1516 & v_1517;
assign v_3149 = v_3144 & v_1515 & ~v_1516 & ~v_1520;
assign v_3151 = v_3150 & v_2113;
assign v_3152 = v_3133 & v_1469 & v_1470 & v_1485 & v_1486;
assign v_3153 = v_3125 & v_1446 & v_1447 & v_1462 & v_1463;
assign v_3155 = v_227;
assign v_3156 = ~v_227 & v_229 & v_262 & ~v_264;
assign v_3157 = ~v_227 & v_229 & v_262 & v_264;
assign v_3158 = ~v_227 & v_229 & ~v_262;
assign v_3161 = v_3160;
assign v_3162 = v_1540;
assign v_3163 = v_12993 & v_12994;
assign v_3165 = v_3164 & ~v_227 & ~v_229 & v_260;
assign v_3167 = v_3166 & v_267 & v_268;
assign v_3168 = v_3166 & v_267 & ~v_268;
assign v_3170 = v_3169 & ~v_279;
assign v_3172 = v_3169 & v_3171;
assign v_3173 = v_3169 & v_279 & v_291 & ~v_292 & v_300;
assign v_3176 = v_3174 & v_3175;
assign v_3177 = v_3174 & v_321 & v_322;
assign v_3178 = v_3174 & v_321 & ~v_322 & v_324;
assign v_3179 = v_3174 & v_321 & ~v_322 & ~v_324 & v_326;
assign v_3180 = v_3174 & v_321 & ~v_322 & ~v_324 & ~v_326;
assign v_3182 = v_3181 & v_1563;
assign v_3184 = v_3183 & ~v_308 & v_309 & v_329;
assign v_3187 = v_3185 & v_3186;
assign v_3188 = v_3185 & v_1570;
assign v_3190 = v_3189 & v_345 & v_346;
assign v_3191 = v_3189 & v_345 & ~v_346 & v_348;
assign v_3192 = v_3189 & v_345 & ~v_346 & ~v_348 & v_350;
assign v_3193 = v_3189 & v_356 & v_357;
assign v_3194 = v_3189 & v_359 & v_360;
assign v_3195 = v_3189 & v_359 & ~v_360 & v_362;
assign v_3196 = v_3189 & v_359 & ~v_360 & ~v_362 & v_364;
assign v_3197 = v_3189 & v_1582;
assign v_3199 = v_3198 & v_1585;
assign v_3201 = v_3200 & v_356 & ~v_357 & v_369 & v_370;
assign v_3202 = v_3200 & v_372 & v_373;
assign v_3203 = v_3200 & v_372 & ~v_373 & v_375;
assign v_3204 = v_3200 & v_372 & ~v_373 & ~v_375 & v_377;
assign v_3206 = v_3200 & v_3205;
assign v_3207 = v_12995 & v_12996;
assign v_3209 = v_3208 & v_384 & v_385;
assign v_3210 = v_3208 & v_384 & ~v_385;
assign v_3212 = v_3211 & v_1599;
assign v_3214 = v_12997 & v_12998;
assign v_3215 = v_3213 & v_391 & v_392;
assign v_3216 = v_3213 & v_391 & ~v_392 & v_394;
assign v_3217 = v_3213 & v_391 & ~v_392 & ~v_394 & v_396;
assign v_3218 = v_3213 & v_1606;
assign v_3220 = v_12999 & v_13000;
assign v_3222 = v_3221 & v_1611;
assign v_3224 = v_3223 & v_410 & v_411;
assign v_3225 = v_3223 & v_410 & ~v_411 & v_413;
assign v_3226 = v_3223 & v_410 & ~v_411 & ~v_413 & v_415;
assign v_3227 = v_3223 & v_421 & v_422;
assign v_3228 = v_3223 & v_424 & v_425;
assign v_3229 = v_3223 & v_424 & ~v_425 & v_427;
assign v_3230 = v_3223 & v_424 & ~v_425 & ~v_427 & v_429;
assign v_3231 = v_3223 & v_1621;
assign v_3233 = v_3232 & v_1624;
assign v_3235 = v_3234 & v_421 & ~v_422 & v_434 & v_435;
assign v_3236 = v_3234 & v_437 & v_438;
assign v_3237 = v_3234 & v_437 & ~v_438 & v_440;
assign v_3238 = v_3234 & v_437 & ~v_438 & ~v_440 & v_442;
assign v_3240 = v_3234 & v_3239;
assign v_3241 = v_13001 & v_13002;
assign v_3243 = v_3242 & v_449 & v_450;
assign v_3244 = v_3242 & v_449 & ~v_450;
assign v_3246 = v_3245 & v_1638;
assign v_3248 = v_13003 & v_13004;
assign v_3249 = v_3247 & v_456 & v_457;
assign v_3250 = v_3247 & v_456 & ~v_457 & v_459;
assign v_3251 = v_3247 & v_456 & ~v_457 & ~v_459 & v_461;
assign v_3252 = v_3247 & v_1645;
assign v_3254 = v_13005 & v_13006;
assign v_3256 = v_3255 & v_1650;
assign v_3258 = v_3257 & v_491;
assign v_3259 = v_3257 & ~v_491 & v_493 & v_526 & ~v_528;
assign v_3260 = v_3257 & ~v_491 & v_493 & v_526 & v_528;
assign v_3261 = v_3257 & ~v_491 & v_493 & ~v_526;
assign v_3262 = v_3257 & v_494;
assign v_3263 = v_3257 & ~v_494;
assign v_3266 = v_3264 & v_3265;
assign v_3267 = v_3264 & v_1666;
assign v_3268 = v_13007 & v_13008;
assign v_3270 = v_3269 & ~v_491 & ~v_493 & v_524;
assign v_3272 = v_3271 & v_531 & v_532;
assign v_3273 = v_3271 & v_531 & ~v_532;
assign v_3275 = v_3274 & v_546 & v_547;
assign v_3276 = v_3274 & v_546 & ~v_547 & ~v_551;
assign v_3278 = v_3277 & v_546 & ~v_547 & v_551;
assign v_3280 = v_3279 & v_554;
assign v_3282 = v_3281 & v_558 & v_559;
assign v_3283 = v_3281 & v_558 & ~v_559 & v_561;
assign v_3284 = v_3281 & v_1682;
assign v_3287 = v_3285 & v_3286;
assign v_3288 = v_3285 & v_1687;
assign v_3290 = v_3289 & v_588 & ~v_589 & ~v_591;
assign v_3291 = v_3289 & v_593 & ~v_594;
assign v_3292 = v_3289 & v_593 & v_594;
assign v_3293 = v_3289 & v_583;
assign v_3295 = v_3294 & v_604 & v_605;
assign v_3296 = v_3294 & v_604 & ~v_605 & ~v_609;
assign v_3298 = v_3297 & v_604 & ~v_605 & v_609;
assign v_3300 = v_3299 & v_612;
assign v_3302 = v_3301 & v_616 & v_617;
assign v_3303 = v_3301 & v_616 & ~v_617 & v_619;
assign v_3304 = v_3301 & v_1700;
assign v_3307 = v_3305 & v_3306;
assign v_3308 = v_3305 & v_1705;
assign v_3310 = v_2 & v_3309;
assign v_3311 = v_641 & v_3289;
assign v_3312 = v_643 & v_3274;
assign v_3313 = v_645 & v_3274;
assign v_3314 = v_647 & v_3274;
assign v_3315 = v_649 & v_3274;
assign v_3316 = ~v_649 & v_3257;
assign v_3318 = ~v_647 & v_3317;
assign v_3320 = ~v_645 & v_3319;
assign v_3322 = ~v_643 & v_3321;
assign v_3324 = ~v_641 & v_3323;
assign v_3326 = ~v_2 & v_3325;
assign v_3328 = v_3327 & ~v_669;
assign v_3329 = v_13009 & v_13010;
assign v_3330 = v_3327 & v_669 & v_670 & v_672 & v_674;
assign v_3331 = v_13011 & v_13012;
assign v_3333 = v_3332 & v_679 & ~v_680 & v_682;
assign v_3334 = v_3332 & v_689 & ~v_690 & ~v_692;
assign v_3335 = v_3332 & v_694 & ~v_695;
assign v_3336 = v_3332 & v_694 & v_695;
assign v_3337 = v_3332 & v_684;
assign v_3339 = v_3338 & v_1737;
assign v_3341 = v_3340 & v_1740;
assign v_3342 = v_3332 & v_679 & v_680;
assign v_3343 = v_3327 & v_1743;
assign v_3345 = v_3344 & ~v_705;
assign v_3346 = v_3344 & v_710 & v_711;
assign v_3347 = v_3344 & v_710 & ~v_711 & ~v_715;
assign v_3349 = v_3348 & v_710 & ~v_711 & v_715;
assign v_3351 = v_3350 & v_718;
assign v_3353 = v_3352 & v_705 & v_722 & v_723 & ~v_724;
assign v_3355 = v_3352 & v_3354;
assign v_3356 = v_3352 & v_750 & v_751;
assign v_3357 = v_3352 & v_750 & ~v_751;
assign v_3359 = v_3358 & v_763 & v_764;
assign v_3360 = v_3358 & v_763 & ~v_764;
assign v_3362 = v_3361 & v_745 & v_758 & v_771;
assign v_3363 = v_13013 & v_13014;
assign v_3364 = v_3352 & v_779 & v_780;
assign v_3365 = v_3352 & v_779 & ~v_780 & ~v_784;
assign v_3367 = v_3366 & v_779 & ~v_780 & v_784;
assign v_3369 = v_3368 & v_787;
assign v_3371 = v_3370 & v_1764;
assign v_3373 = v_3372 & v_798 & ~v_799 & v_817;
assign v_3374 = v_3372 & v_798 & ~v_799 & ~v_817;
assign v_3375 = v_3372 & ~v_800;
assign v_3376 = v_3372 & v_808 & ~v_809;
assign v_3377 = v_3372 & v_1771;
assign v_3379 = v_3378 & v_798 & v_799 & v_814 & ~v_815;
assign v_3381 = v_3380 & v_821 & ~v_822 & v_840;
assign v_3382 = v_3380 & v_821 & ~v_822 & ~v_840;
assign v_3383 = v_3380 & ~v_823;
assign v_3384 = v_3380 & v_831 & ~v_832;
assign v_3385 = v_3380 & v_1780;
assign v_3387 = v_3386 & v_821 & v_822 & v_837 & ~v_838;
assign v_3389 = v_3388 & v_844 & ~v_845 & v_863;
assign v_3390 = v_3388 & ~v_846;
assign v_3391 = v_3388 & v_854 & ~v_855;
assign v_3392 = v_3388 & v_1788;
assign v_3394 = v_3393 & v_844 & v_845 & v_860 & v_861;
assign v_3395 = v_3388 & v_844 & ~v_845 & ~v_863;
assign v_3396 = v_3393 & v_844 & v_845 & v_860 & ~v_861;
assign v_3399 = v_3397 & v_3398;
assign v_3400 = v_3397 & v_867 & v_868 & ~v_869 & ~v_870;
assign v_3401 = v_3397 & v_867 & v_868 & v_869;
assign v_3402 = v_3397 & v_867 & ~v_868 & ~v_872;
assign v_3404 = v_3403 & v_1801;
assign v_3405 = v_3386 & v_821 & v_822 & v_837 & v_838;
assign v_3406 = v_3378 & v_798 & v_799 & v_814 & v_815;
assign v_3408 = v_3407 & v_879 & ~v_880 & v_898;
assign v_3409 = v_3407 & v_879 & ~v_880 & ~v_898;
assign v_3410 = v_3407 & ~v_881;
assign v_3411 = v_3407 & v_889 & ~v_890;
assign v_3412 = v_3407 & v_1810;
assign v_3414 = v_3413 & v_879 & v_880 & v_895 & ~v_896;
assign v_3416 = v_3415 & v_902 & ~v_903 & v_921;
assign v_3417 = v_3415 & v_902 & ~v_903 & ~v_921;
assign v_3418 = v_3415 & ~v_904;
assign v_3419 = v_3415 & v_912 & ~v_913;
assign v_3420 = v_3415 & v_1819;
assign v_3422 = v_3421 & v_902 & v_903 & v_918 & ~v_919;
assign v_3424 = v_3423 & v_925 & ~v_926 & v_944;
assign v_3425 = v_3423 & ~v_927;
assign v_3426 = v_3423 & v_935 & ~v_936;
assign v_3427 = v_3423 & v_1827;
assign v_3429 = v_3428 & v_925 & v_926 & v_941 & v_942;
assign v_3430 = v_3423 & v_925 & ~v_926 & ~v_944;
assign v_3431 = v_3428 & v_925 & v_926 & v_941 & ~v_942;
assign v_3434 = v_3432 & v_3433;
assign v_3435 = v_3432 & v_948 & v_949 & ~v_950 & ~v_951;
assign v_3436 = v_3432 & v_948 & v_949 & v_950;
assign v_3437 = v_3432 & v_948 & ~v_949 & ~v_953;
assign v_3439 = v_3438 & v_1840;
assign v_3440 = v_3421 & v_902 & v_903 & v_918 & v_919;
assign v_3441 = v_3413 & v_879 & v_880 & v_895 & v_896;
assign v_3443 = v_3442 & v_960 & ~v_961 & v_979;
assign v_3444 = v_3442 & v_960 & ~v_961 & ~v_979;
assign v_3445 = v_3442 & ~v_962;
assign v_3446 = v_3442 & v_970 & ~v_971;
assign v_3447 = v_3442 & v_1849;
assign v_3449 = v_3448 & v_960 & v_961 & v_976 & ~v_977;
assign v_3451 = v_3450 & v_983 & ~v_984 & v_1002;
assign v_3452 = v_3450 & v_983 & ~v_984 & ~v_1002;
assign v_3453 = v_3450 & ~v_985;
assign v_3454 = v_3450 & v_993 & ~v_994;
assign v_3455 = v_3450 & v_1858;
assign v_3457 = v_3456 & v_983 & v_984 & v_999 & ~v_1000;
assign v_3459 = v_3458 & v_1006 & ~v_1007 & v_1025;
assign v_3460 = v_3458 & ~v_1008;
assign v_3461 = v_3458 & v_1016 & ~v_1017;
assign v_3462 = v_3458 & v_1866;
assign v_3464 = v_3463 & v_1006 & v_1007 & v_1022 & v_1023;
assign v_3465 = v_3458 & v_1006 & ~v_1007 & ~v_1025;
assign v_3466 = v_3463 & v_1006 & v_1007 & v_1022 & ~v_1023;
assign v_3469 = v_3467 & v_3468;
assign v_3470 = v_3467 & v_1029 & v_1030 & ~v_1031 & ~v_1032;
assign v_3471 = v_3467 & v_1029 & v_1030 & v_1031;
assign v_3472 = v_3467 & v_1029 & ~v_1030 & ~v_1034;
assign v_3474 = v_3473 & v_1879;
assign v_3475 = v_3456 & v_983 & v_984 & v_999 & v_1000;
assign v_3476 = v_3448 & v_960 & v_961 & v_976 & v_977;
assign v_3478 = v_3477 & v_1041 & ~v_1042 & v_1060;
assign v_3479 = v_3477 & v_1041 & ~v_1042 & ~v_1060;
assign v_3480 = v_3477 & ~v_1043;
assign v_3481 = v_3477 & v_1051 & ~v_1052;
assign v_3482 = v_3477 & v_1888;
assign v_3484 = v_3483 & v_1041 & v_1042 & v_1057 & ~v_1058;
assign v_3486 = v_3485 & v_1064 & ~v_1065 & v_1083;
assign v_3487 = v_3485 & v_1064 & ~v_1065 & ~v_1083;
assign v_3488 = v_3485 & ~v_1066;
assign v_3489 = v_3485 & v_1074 & ~v_1075;
assign v_3490 = v_3485 & v_1897;
assign v_3492 = v_3491 & v_1064 & v_1065 & v_1080 & ~v_1081;
assign v_3494 = v_3493 & v_1087 & ~v_1088 & v_1106;
assign v_3495 = v_3493 & ~v_1089;
assign v_3496 = v_3493 & v_1097 & ~v_1098;
assign v_3497 = v_3493 & v_1905;
assign v_3499 = v_3498 & v_1087 & v_1088 & v_1103 & v_1104;
assign v_3500 = v_3493 & v_1087 & ~v_1088 & ~v_1106;
assign v_3501 = v_3498 & v_1087 & v_1088 & v_1103 & ~v_1104;
assign v_3504 = v_3502 & v_3503;
assign v_3505 = v_3502 & v_1110 & v_1111 & ~v_1112 & ~v_1113;
assign v_3506 = v_3502 & v_1110 & v_1111 & v_1112;
assign v_3507 = v_3502 & v_1110 & ~v_1111 & ~v_1115;
assign v_3509 = v_3508 & v_1918;
assign v_3510 = v_3491 & v_1064 & v_1065 & v_1080 & v_1081;
assign v_3511 = v_3483 & v_1041 & v_1042 & v_1057 & v_1058;
assign v_3513 = v_3512 & v_1122 & ~v_1123 & v_1141;
assign v_3514 = v_3512 & v_1122 & ~v_1123 & ~v_1141;
assign v_3515 = v_3512 & ~v_1124;
assign v_3516 = v_3512 & v_1132 & ~v_1133;
assign v_3517 = v_3512 & v_1927;
assign v_3519 = v_3518 & v_1122 & v_1123 & v_1138 & ~v_1139;
assign v_3521 = v_3520 & v_1145 & ~v_1146 & v_1164;
assign v_3522 = v_3520 & v_1145 & ~v_1146 & ~v_1164;
assign v_3523 = v_3520 & ~v_1147;
assign v_3524 = v_3520 & v_1155 & ~v_1156;
assign v_3525 = v_3520 & v_1936;
assign v_3527 = v_3526 & v_1145 & v_1146 & v_1161 & ~v_1162;
assign v_3529 = v_3528 & v_1168 & ~v_1169 & v_1187;
assign v_3530 = v_3528 & ~v_1170;
assign v_3531 = v_3528 & v_1178 & ~v_1179;
assign v_3532 = v_3528 & v_1944;
assign v_3534 = v_3533 & v_1168 & v_1169 & v_1184 & v_1185;
assign v_3535 = v_3528 & v_1168 & ~v_1169 & ~v_1187;
assign v_3536 = v_3533 & v_1168 & v_1169 & v_1184 & ~v_1185;
assign v_3539 = v_3537 & v_3538;
assign v_3540 = v_3537 & v_1191 & v_1192 & ~v_1193 & ~v_1194;
assign v_3541 = v_3537 & v_1191 & v_1192 & v_1193;
assign v_3542 = v_3537 & v_1191 & ~v_1192 & ~v_1196;
assign v_3544 = v_3543 & v_1957;
assign v_3545 = v_3526 & v_1145 & v_1146 & v_1161 & v_1162;
assign v_3546 = v_3518 & v_1122 & v_1123 & v_1138 & v_1139;
assign v_3548 = v_3547 & v_1203 & ~v_1204 & v_1222;
assign v_3549 = v_3547 & v_1203 & ~v_1204 & ~v_1222;
assign v_3550 = v_3547 & ~v_1205;
assign v_3551 = v_3547 & v_1213 & ~v_1214;
assign v_3552 = v_3547 & v_1966;
assign v_3554 = v_3553 & v_1203 & v_1204 & v_1219 & ~v_1220;
assign v_3556 = v_3555 & v_1226 & ~v_1227 & v_1245;
assign v_3557 = v_3555 & v_1226 & ~v_1227 & ~v_1245;
assign v_3558 = v_3555 & ~v_1228;
assign v_3559 = v_3555 & v_1236 & ~v_1237;
assign v_3560 = v_3555 & v_1975;
assign v_3562 = v_3561 & v_1226 & v_1227 & v_1242 & ~v_1243;
assign v_3564 = v_3563 & v_1249 & ~v_1250 & v_1268;
assign v_3565 = v_3563 & ~v_1251;
assign v_3566 = v_3563 & v_1259 & ~v_1260;
assign v_3567 = v_3563 & v_1983;
assign v_3569 = v_3568 & v_1249 & v_1250 & v_1265 & v_1266;
assign v_3570 = v_3563 & v_1249 & ~v_1250 & ~v_1268;
assign v_3571 = v_3568 & v_1249 & v_1250 & v_1265 & ~v_1266;
assign v_3574 = v_3572 & v_3573;
assign v_3575 = v_3572 & v_1272 & v_1273 & ~v_1274 & ~v_1275;
assign v_3576 = v_3572 & v_1272 & v_1273 & v_1274;
assign v_3577 = v_3572 & v_1272 & ~v_1273 & ~v_1277;
assign v_3579 = v_3578 & v_1996;
assign v_3580 = v_3561 & v_1226 & v_1227 & v_1242 & v_1243;
assign v_3581 = v_3553 & v_1203 & v_1204 & v_1219 & v_1220;
assign v_3583 = v_3582 & v_1284 & ~v_1285 & v_1303;
assign v_3584 = v_3582 & v_1284 & ~v_1285 & ~v_1303;
assign v_3585 = v_3582 & ~v_1286;
assign v_3586 = v_3582 & v_1294 & ~v_1295;
assign v_3587 = v_3582 & v_2005;
assign v_3589 = v_3588 & v_1284 & v_1285 & v_1300 & ~v_1301;
assign v_3591 = v_3590 & v_1307 & ~v_1308 & v_1326;
assign v_3592 = v_3590 & v_1307 & ~v_1308 & ~v_1326;
assign v_3593 = v_3590 & ~v_1309;
assign v_3594 = v_3590 & v_1317 & ~v_1318;
assign v_3595 = v_3590 & v_2014;
assign v_3597 = v_3596 & v_1307 & v_1308 & v_1323 & ~v_1324;
assign v_3599 = v_3598 & v_1330 & ~v_1331 & v_1349;
assign v_3600 = v_3598 & ~v_1332;
assign v_3601 = v_3598 & v_1340 & ~v_1341;
assign v_3602 = v_3598 & v_2022;
assign v_3604 = v_3603 & v_1330 & v_1331 & v_1346 & v_1347;
assign v_3605 = v_3598 & v_1330 & ~v_1331 & ~v_1349;
assign v_3606 = v_3603 & v_1330 & v_1331 & v_1346 & ~v_1347;
assign v_3609 = v_3607 & v_3608;
assign v_3610 = v_3607 & v_1353 & v_1354 & ~v_1355 & ~v_1356;
assign v_3611 = v_3607 & v_1353 & v_1354 & v_1355;
assign v_3612 = v_3607 & v_1353 & ~v_1354 & ~v_1358;
assign v_3614 = v_3613 & v_2035;
assign v_3615 = v_3596 & v_1307 & v_1308 & v_1323 & v_1324;
assign v_3616 = v_3588 & v_1284 & v_1285 & v_1300 & v_1301;
assign v_3618 = v_3617 & v_1365 & ~v_1366 & v_1384;
assign v_3619 = v_3617 & v_1365 & ~v_1366 & ~v_1384;
assign v_3620 = v_3617 & ~v_1367;
assign v_3621 = v_3617 & v_1375 & ~v_1376;
assign v_3622 = v_3617 & v_2044;
assign v_3624 = v_3623 & v_1365 & v_1366 & v_1381 & ~v_1382;
assign v_3626 = v_3625 & v_1388 & ~v_1389 & v_1407;
assign v_3627 = v_3625 & v_1388 & ~v_1389 & ~v_1407;
assign v_3628 = v_3625 & ~v_1390;
assign v_3629 = v_3625 & v_1398 & ~v_1399;
assign v_3630 = v_3625 & v_2053;
assign v_3632 = v_3631 & v_1388 & v_1389 & v_1404 & ~v_1405;
assign v_3634 = v_3633 & v_1411 & ~v_1412 & v_1430;
assign v_3635 = v_3633 & ~v_1413;
assign v_3636 = v_3633 & v_1421 & ~v_1422;
assign v_3637 = v_3633 & v_2061;
assign v_3639 = v_3638 & v_1411 & v_1412 & v_1427 & v_1428;
assign v_3640 = v_3633 & v_1411 & ~v_1412 & ~v_1430;
assign v_3641 = v_3638 & v_1411 & v_1412 & v_1427 & ~v_1428;
assign v_3644 = v_3642 & v_3643;
assign v_3645 = v_3642 & v_1434 & v_1435 & ~v_1436 & ~v_1437;
assign v_3646 = v_3642 & v_1434 & v_1435 & v_1436;
assign v_3647 = v_3642 & v_1434 & ~v_1435 & ~v_1439;
assign v_3649 = v_3648 & v_2074;
assign v_3650 = v_3631 & v_1388 & v_1389 & v_1404 & v_1405;
assign v_3651 = v_3623 & v_1365 & v_1366 & v_1381 & v_1382;
assign v_3653 = v_3652 & v_1446 & ~v_1447 & v_1465;
assign v_3654 = v_3652 & v_1446 & ~v_1447 & ~v_1465;
assign v_3655 = v_3652 & ~v_1448;
assign v_3656 = v_3652 & v_1456 & ~v_1457;
assign v_3657 = v_3652 & v_2083;
assign v_3659 = v_3658 & v_1446 & v_1447 & v_1462 & ~v_1463;
assign v_3661 = v_3660 & v_1469 & ~v_1470 & v_1488;
assign v_3662 = v_3660 & v_1469 & ~v_1470 & ~v_1488;
assign v_3663 = v_3660 & ~v_1471;
assign v_3664 = v_3660 & v_1479 & ~v_1480;
assign v_3665 = v_3660 & v_2092;
assign v_3667 = v_3666 & v_1469 & v_1470 & v_1485 & ~v_1486;
assign v_3669 = v_3668 & v_1492 & ~v_1493 & v_1511;
assign v_3670 = v_3668 & ~v_1494;
assign v_3671 = v_3668 & v_1502 & ~v_1503;
assign v_3672 = v_3668 & v_2100;
assign v_3674 = v_3673 & v_1492 & v_1493 & v_1508 & v_1509;
assign v_3675 = v_3668 & v_1492 & ~v_1493 & ~v_1511;
assign v_3676 = v_3673 & v_1492 & v_1493 & v_1508 & ~v_1509;
assign v_3679 = v_3677 & v_3678;
assign v_3680 = v_3677 & v_1515 & v_1516 & ~v_1517 & ~v_1518;
assign v_3681 = v_3677 & v_1515 & v_1516 & v_1517;
assign v_3682 = v_3677 & v_1515 & ~v_1516 & ~v_1520;
assign v_3684 = v_3683 & v_2113;
assign v_3685 = v_3666 & v_1469 & v_1470 & v_1485 & v_1486;
assign v_3686 = v_3658 & v_1446 & v_1447 & v_1462 & v_1463;
assign v_3689 = v_3688 & v_227;
assign v_3690 = v_3688 & ~v_227 & v_229 & v_262 & ~v_264;
assign v_3691 = v_3688 & ~v_227 & v_229 & v_262 & v_264;
assign v_3692 = v_3688 & ~v_227 & v_229 & ~v_262;
assign v_3693 = v_3688 & v_230;
assign v_3694 = v_3688 & ~v_230;
assign v_3697 = v_3695 & v_3696;
assign v_3698 = v_3695 & v_1540;
assign v_3699 = v_13015 & v_13016;
assign v_3701 = v_3700 & ~v_227 & ~v_229 & v_260;
assign v_3703 = v_3702 & v_267 & v_268;
assign v_3704 = v_3702 & v_267 & ~v_268;
assign v_3706 = v_3705 & ~v_279;
assign v_3708 = v_3705 & v_3707;
assign v_3709 = v_3705 & v_279 & v_291 & ~v_292 & v_300;
assign v_3712 = v_3710 & v_3711;
assign v_3713 = v_3710 & v_321 & v_322;
assign v_3714 = v_3710 & v_321 & ~v_322 & v_324;
assign v_3715 = v_3710 & v_321 & ~v_322 & ~v_324 & v_326;
assign v_3716 = v_3710 & v_321 & ~v_322 & ~v_324 & ~v_326;
assign v_3718 = v_3717 & v_1563;
assign v_3720 = v_3719 & ~v_308 & v_309 & v_329;
assign v_3723 = v_3721 & v_3722;
assign v_3724 = v_3721 & v_1570;
assign v_3726 = v_3725 & v_345 & v_346;
assign v_3727 = v_3725 & v_345 & ~v_346 & v_348;
assign v_3728 = v_3725 & v_345 & ~v_346 & ~v_348 & v_350;
assign v_3729 = v_3725 & v_356 & v_357;
assign v_3730 = v_3725 & v_359 & v_360;
assign v_3731 = v_3725 & v_359 & ~v_360 & v_362;
assign v_3732 = v_3725 & v_359 & ~v_360 & ~v_362 & v_364;
assign v_3733 = v_3725 & v_1582;
assign v_3735 = v_3734 & v_1585;
assign v_3737 = v_3736 & v_356 & ~v_357 & v_369 & v_370;
assign v_3738 = v_3736 & v_372 & v_373;
assign v_3739 = v_3736 & v_372 & ~v_373 & v_375;
assign v_3740 = v_3736 & v_372 & ~v_373 & ~v_375 & v_377;
assign v_3742 = v_3736 & v_3741;
assign v_3743 = v_13017 & v_13018;
assign v_3745 = v_3744 & v_384 & v_385;
assign v_3746 = v_3744 & v_384 & ~v_385;
assign v_3748 = v_3747 & v_1599;
assign v_3750 = v_13019 & v_13020;
assign v_3751 = v_3749 & v_391 & v_392;
assign v_3752 = v_3749 & v_391 & ~v_392 & v_394;
assign v_3753 = v_3749 & v_391 & ~v_392 & ~v_394 & v_396;
assign v_3754 = v_3749 & v_1606;
assign v_3756 = v_13021 & v_13022;
assign v_3758 = v_3757 & v_1611;
assign v_3760 = v_3759 & v_410 & v_411;
assign v_3761 = v_3759 & v_410 & ~v_411 & v_413;
assign v_3762 = v_3759 & v_410 & ~v_411 & ~v_413 & v_415;
assign v_3763 = v_3759 & v_421 & v_422;
assign v_3764 = v_3759 & v_424 & v_425;
assign v_3765 = v_3759 & v_424 & ~v_425 & v_427;
assign v_3766 = v_3759 & v_424 & ~v_425 & ~v_427 & v_429;
assign v_3767 = v_3759 & v_1621;
assign v_3769 = v_3768 & v_1624;
assign v_3771 = v_3770 & v_421 & ~v_422 & v_434 & v_435;
assign v_3772 = v_3770 & v_437 & v_438;
assign v_3773 = v_3770 & v_437 & ~v_438 & v_440;
assign v_3774 = v_3770 & v_437 & ~v_438 & ~v_440 & v_442;
assign v_3776 = v_3770 & v_3775;
assign v_3777 = v_13023 & v_13024;
assign v_3779 = v_3778 & v_449 & v_450;
assign v_3780 = v_3778 & v_449 & ~v_450;
assign v_3782 = v_3781 & v_1638;
assign v_3784 = v_13025 & v_13026;
assign v_3785 = v_3783 & v_456 & v_457;
assign v_3786 = v_3783 & v_456 & ~v_457 & v_459;
assign v_3787 = v_3783 & v_456 & ~v_457 & ~v_459 & v_461;
assign v_3788 = v_3783 & v_1645;
assign v_3790 = v_13027 & v_13028;
assign v_3792 = v_3791 & v_1650;
assign v_3794 = v_3793 & v_491;
assign v_3795 = v_3793 & ~v_491 & v_493 & v_526 & ~v_528;
assign v_3796 = v_3793 & ~v_491 & v_493 & v_526 & v_528;
assign v_3797 = v_3793 & ~v_491 & v_493 & ~v_526;
assign v_3798 = v_3793 & v_494;
assign v_3799 = v_3793 & ~v_494;
assign v_3802 = v_3800 & v_3801;
assign v_3803 = v_3800 & v_1666;
assign v_3804 = v_13029 & v_13030;
assign v_3806 = v_3805 & ~v_491 & ~v_493 & v_524;
assign v_3808 = v_3807 & v_531 & v_532;
assign v_3809 = v_3807 & v_531 & ~v_532;
assign v_3811 = v_3810 & v_546 & v_547;
assign v_3812 = v_3810 & v_546 & ~v_547 & ~v_551;
assign v_3814 = v_3813 & v_546 & ~v_547 & v_551;
assign v_3816 = v_3815 & v_554;
assign v_3818 = v_3817 & v_558 & v_559;
assign v_3819 = v_3817 & v_558 & ~v_559 & v_561;
assign v_3820 = v_3817 & v_1682;
assign v_3823 = v_3821 & v_3822;
assign v_3824 = v_3821 & v_1687;
assign v_3826 = v_3825 & v_588 & ~v_589 & ~v_591;
assign v_3827 = v_3825 & v_593 & ~v_594;
assign v_3828 = v_3825 & v_593 & v_594;
assign v_3829 = v_3825 & v_583;
assign v_3831 = v_3830 & v_604 & v_605;
assign v_3832 = v_3830 & v_604 & ~v_605 & ~v_609;
assign v_3834 = v_3833 & v_604 & ~v_605 & v_609;
assign v_3836 = v_3835 & v_612;
assign v_3838 = v_3837 & v_616 & v_617;
assign v_3839 = v_3837 & v_616 & ~v_617 & v_619;
assign v_3840 = v_3837 & v_1700;
assign v_3843 = v_3841 & v_3842;
assign v_3844 = v_3841 & v_1705;
assign v_3846 = v_2 & v_3845;
assign v_3847 = v_641 & v_3825;
assign v_3848 = v_643 & v_3810;
assign v_3849 = v_645 & v_3810;
assign v_3850 = v_647 & v_3810;
assign v_3851 = v_649 & v_3810;
assign v_3852 = ~v_649 & v_3793;
assign v_3854 = ~v_647 & v_3853;
assign v_3856 = ~v_645 & v_3855;
assign v_3858 = ~v_643 & v_3857;
assign v_3860 = ~v_641 & v_3859;
assign v_3862 = ~v_2 & v_3861;
assign v_3864 = v_3863 & ~v_669;
assign v_3865 = v_13031 & v_13032;
assign v_3866 = v_3863 & v_669 & v_670 & v_672 & v_674;
assign v_3867 = v_13033 & v_13034;
assign v_3869 = v_3868 & v_679 & ~v_680 & v_682;
assign v_3870 = v_3868 & v_689 & ~v_690 & ~v_692;
assign v_3871 = v_3868 & v_694 & ~v_695;
assign v_3872 = v_3868 & v_694 & v_695;
assign v_3873 = v_3868 & v_684;
assign v_3875 = v_3874 & v_1737;
assign v_3877 = v_3876 & v_1740;
assign v_3878 = v_3868 & v_679 & v_680;
assign v_3879 = v_3863 & v_1743;
assign v_3881 = v_3880 & ~v_705;
assign v_3882 = v_3880 & v_710 & v_711;
assign v_3883 = v_3880 & v_710 & ~v_711 & ~v_715;
assign v_3885 = v_3884 & v_710 & ~v_711 & v_715;
assign v_3887 = v_3886 & v_718;
assign v_3889 = v_3888 & v_705 & v_722 & v_723 & ~v_724;
assign v_3891 = v_3888 & v_3890;
assign v_3892 = v_3888 & v_750 & v_751;
assign v_3893 = v_3888 & v_750 & ~v_751;
assign v_3895 = v_3894 & v_763 & v_764;
assign v_3896 = v_3894 & v_763 & ~v_764;
assign v_3898 = v_3897 & v_745 & v_758 & v_771;
assign v_3899 = v_13035 & v_13036;
assign v_3900 = v_3888 & v_779 & v_780;
assign v_3901 = v_3888 & v_779 & ~v_780 & ~v_784;
assign v_3903 = v_3902 & v_779 & ~v_780 & v_784;
assign v_3905 = v_3904 & v_787;
assign v_3907 = v_3906 & v_1764;
assign v_3909 = v_3908 & v_798 & ~v_799 & v_817;
assign v_3910 = v_3908 & v_798 & ~v_799 & ~v_817;
assign v_3911 = v_3908 & ~v_800;
assign v_3912 = v_3908 & v_808 & ~v_809;
assign v_3913 = v_3908 & v_1771;
assign v_3915 = v_3914 & v_798 & v_799 & v_814 & ~v_815;
assign v_3917 = v_3916 & v_821 & ~v_822 & v_840;
assign v_3918 = v_3916 & v_821 & ~v_822 & ~v_840;
assign v_3919 = v_3916 & ~v_823;
assign v_3920 = v_3916 & v_831 & ~v_832;
assign v_3921 = v_3916 & v_1780;
assign v_3923 = v_3922 & v_821 & v_822 & v_837 & ~v_838;
assign v_3925 = v_3924 & v_844 & ~v_845 & v_863;
assign v_3926 = v_3924 & ~v_846;
assign v_3927 = v_3924 & v_854 & ~v_855;
assign v_3928 = v_3924 & v_1788;
assign v_3930 = v_3929 & v_844 & v_845 & v_860 & v_861;
assign v_3931 = v_3924 & v_844 & ~v_845 & ~v_863;
assign v_3932 = v_3929 & v_844 & v_845 & v_860 & ~v_861;
assign v_3935 = v_3933 & v_3934;
assign v_3936 = v_3933 & v_867 & v_868 & ~v_869 & ~v_870;
assign v_3937 = v_3933 & v_867 & v_868 & v_869;
assign v_3938 = v_3933 & v_867 & ~v_868 & ~v_872;
assign v_3940 = v_3939 & v_1801;
assign v_3941 = v_3922 & v_821 & v_822 & v_837 & v_838;
assign v_3942 = v_3914 & v_798 & v_799 & v_814 & v_815;
assign v_3944 = v_3943 & v_879 & ~v_880 & v_898;
assign v_3945 = v_3943 & v_879 & ~v_880 & ~v_898;
assign v_3946 = v_3943 & ~v_881;
assign v_3947 = v_3943 & v_889 & ~v_890;
assign v_3948 = v_3943 & v_1810;
assign v_3950 = v_3949 & v_879 & v_880 & v_895 & ~v_896;
assign v_3952 = v_3951 & v_902 & ~v_903 & v_921;
assign v_3953 = v_3951 & v_902 & ~v_903 & ~v_921;
assign v_3954 = v_3951 & ~v_904;
assign v_3955 = v_3951 & v_912 & ~v_913;
assign v_3956 = v_3951 & v_1819;
assign v_3958 = v_3957 & v_902 & v_903 & v_918 & ~v_919;
assign v_3960 = v_3959 & v_925 & ~v_926 & v_944;
assign v_3961 = v_3959 & ~v_927;
assign v_3962 = v_3959 & v_935 & ~v_936;
assign v_3963 = v_3959 & v_1827;
assign v_3965 = v_3964 & v_925 & v_926 & v_941 & v_942;
assign v_3966 = v_3959 & v_925 & ~v_926 & ~v_944;
assign v_3967 = v_3964 & v_925 & v_926 & v_941 & ~v_942;
assign v_3970 = v_3968 & v_3969;
assign v_3971 = v_3968 & v_948 & v_949 & ~v_950 & ~v_951;
assign v_3972 = v_3968 & v_948 & v_949 & v_950;
assign v_3973 = v_3968 & v_948 & ~v_949 & ~v_953;
assign v_3975 = v_3974 & v_1840;
assign v_3976 = v_3957 & v_902 & v_903 & v_918 & v_919;
assign v_3977 = v_3949 & v_879 & v_880 & v_895 & v_896;
assign v_3979 = v_3978 & v_960 & ~v_961 & v_979;
assign v_3980 = v_3978 & v_960 & ~v_961 & ~v_979;
assign v_3981 = v_3978 & ~v_962;
assign v_3982 = v_3978 & v_970 & ~v_971;
assign v_3983 = v_3978 & v_1849;
assign v_3985 = v_3984 & v_960 & v_961 & v_976 & ~v_977;
assign v_3987 = v_3986 & v_983 & ~v_984 & v_1002;
assign v_3988 = v_3986 & v_983 & ~v_984 & ~v_1002;
assign v_3989 = v_3986 & ~v_985;
assign v_3990 = v_3986 & v_993 & ~v_994;
assign v_3991 = v_3986 & v_1858;
assign v_3993 = v_3992 & v_983 & v_984 & v_999 & ~v_1000;
assign v_3995 = v_3994 & v_1006 & ~v_1007 & v_1025;
assign v_3996 = v_3994 & ~v_1008;
assign v_3997 = v_3994 & v_1016 & ~v_1017;
assign v_3998 = v_3994 & v_1866;
assign v_4000 = v_3999 & v_1006 & v_1007 & v_1022 & v_1023;
assign v_4001 = v_3994 & v_1006 & ~v_1007 & ~v_1025;
assign v_4002 = v_3999 & v_1006 & v_1007 & v_1022 & ~v_1023;
assign v_4005 = v_4003 & v_4004;
assign v_4006 = v_4003 & v_1029 & v_1030 & ~v_1031 & ~v_1032;
assign v_4007 = v_4003 & v_1029 & v_1030 & v_1031;
assign v_4008 = v_4003 & v_1029 & ~v_1030 & ~v_1034;
assign v_4010 = v_4009 & v_1879;
assign v_4011 = v_3992 & v_983 & v_984 & v_999 & v_1000;
assign v_4012 = v_3984 & v_960 & v_961 & v_976 & v_977;
assign v_4014 = v_4013 & v_1041 & ~v_1042 & v_1060;
assign v_4015 = v_4013 & v_1041 & ~v_1042 & ~v_1060;
assign v_4016 = v_4013 & ~v_1043;
assign v_4017 = v_4013 & v_1051 & ~v_1052;
assign v_4018 = v_4013 & v_1888;
assign v_4020 = v_4019 & v_1041 & v_1042 & v_1057 & ~v_1058;
assign v_4022 = v_4021 & v_1064 & ~v_1065 & v_1083;
assign v_4023 = v_4021 & v_1064 & ~v_1065 & ~v_1083;
assign v_4024 = v_4021 & ~v_1066;
assign v_4025 = v_4021 & v_1074 & ~v_1075;
assign v_4026 = v_4021 & v_1897;
assign v_4028 = v_4027 & v_1064 & v_1065 & v_1080 & ~v_1081;
assign v_4030 = v_4029 & v_1087 & ~v_1088 & v_1106;
assign v_4031 = v_4029 & ~v_1089;
assign v_4032 = v_4029 & v_1097 & ~v_1098;
assign v_4033 = v_4029 & v_1905;
assign v_4035 = v_4034 & v_1087 & v_1088 & v_1103 & v_1104;
assign v_4036 = v_4029 & v_1087 & ~v_1088 & ~v_1106;
assign v_4037 = v_4034 & v_1087 & v_1088 & v_1103 & ~v_1104;
assign v_4040 = v_4038 & v_4039;
assign v_4041 = v_4038 & v_1110 & v_1111 & ~v_1112 & ~v_1113;
assign v_4042 = v_4038 & v_1110 & v_1111 & v_1112;
assign v_4043 = v_4038 & v_1110 & ~v_1111 & ~v_1115;
assign v_4045 = v_4044 & v_1918;
assign v_4046 = v_4027 & v_1064 & v_1065 & v_1080 & v_1081;
assign v_4047 = v_4019 & v_1041 & v_1042 & v_1057 & v_1058;
assign v_4049 = v_4048 & v_1122 & ~v_1123 & v_1141;
assign v_4050 = v_4048 & v_1122 & ~v_1123 & ~v_1141;
assign v_4051 = v_4048 & ~v_1124;
assign v_4052 = v_4048 & v_1132 & ~v_1133;
assign v_4053 = v_4048 & v_1927;
assign v_4055 = v_4054 & v_1122 & v_1123 & v_1138 & ~v_1139;
assign v_4057 = v_4056 & v_1145 & ~v_1146 & v_1164;
assign v_4058 = v_4056 & v_1145 & ~v_1146 & ~v_1164;
assign v_4059 = v_4056 & ~v_1147;
assign v_4060 = v_4056 & v_1155 & ~v_1156;
assign v_4061 = v_4056 & v_1936;
assign v_4063 = v_4062 & v_1145 & v_1146 & v_1161 & ~v_1162;
assign v_4065 = v_4064 & v_1168 & ~v_1169 & v_1187;
assign v_4066 = v_4064 & ~v_1170;
assign v_4067 = v_4064 & v_1178 & ~v_1179;
assign v_4068 = v_4064 & v_1944;
assign v_4070 = v_4069 & v_1168 & v_1169 & v_1184 & v_1185;
assign v_4071 = v_4064 & v_1168 & ~v_1169 & ~v_1187;
assign v_4072 = v_4069 & v_1168 & v_1169 & v_1184 & ~v_1185;
assign v_4075 = v_4073 & v_4074;
assign v_4076 = v_4073 & v_1191 & v_1192 & ~v_1193 & ~v_1194;
assign v_4077 = v_4073 & v_1191 & v_1192 & v_1193;
assign v_4078 = v_4073 & v_1191 & ~v_1192 & ~v_1196;
assign v_4080 = v_4079 & v_1957;
assign v_4081 = v_4062 & v_1145 & v_1146 & v_1161 & v_1162;
assign v_4082 = v_4054 & v_1122 & v_1123 & v_1138 & v_1139;
assign v_4084 = v_4083 & v_1203 & ~v_1204 & v_1222;
assign v_4085 = v_4083 & v_1203 & ~v_1204 & ~v_1222;
assign v_4086 = v_4083 & ~v_1205;
assign v_4087 = v_4083 & v_1213 & ~v_1214;
assign v_4088 = v_4083 & v_1966;
assign v_4090 = v_4089 & v_1203 & v_1204 & v_1219 & ~v_1220;
assign v_4092 = v_4091 & v_1226 & ~v_1227 & v_1245;
assign v_4093 = v_4091 & v_1226 & ~v_1227 & ~v_1245;
assign v_4094 = v_4091 & ~v_1228;
assign v_4095 = v_4091 & v_1236 & ~v_1237;
assign v_4096 = v_4091 & v_1975;
assign v_4098 = v_4097 & v_1226 & v_1227 & v_1242 & ~v_1243;
assign v_4100 = v_4099 & v_1249 & ~v_1250 & v_1268;
assign v_4101 = v_4099 & ~v_1251;
assign v_4102 = v_4099 & v_1259 & ~v_1260;
assign v_4103 = v_4099 & v_1983;
assign v_4105 = v_4104 & v_1249 & v_1250 & v_1265 & v_1266;
assign v_4106 = v_4099 & v_1249 & ~v_1250 & ~v_1268;
assign v_4107 = v_4104 & v_1249 & v_1250 & v_1265 & ~v_1266;
assign v_4110 = v_4108 & v_4109;
assign v_4111 = v_4108 & v_1272 & v_1273 & ~v_1274 & ~v_1275;
assign v_4112 = v_4108 & v_1272 & v_1273 & v_1274;
assign v_4113 = v_4108 & v_1272 & ~v_1273 & ~v_1277;
assign v_4115 = v_4114 & v_1996;
assign v_4116 = v_4097 & v_1226 & v_1227 & v_1242 & v_1243;
assign v_4117 = v_4089 & v_1203 & v_1204 & v_1219 & v_1220;
assign v_4119 = v_4118 & v_1284 & ~v_1285 & v_1303;
assign v_4120 = v_4118 & v_1284 & ~v_1285 & ~v_1303;
assign v_4121 = v_4118 & ~v_1286;
assign v_4122 = v_4118 & v_1294 & ~v_1295;
assign v_4123 = v_4118 & v_2005;
assign v_4125 = v_4124 & v_1284 & v_1285 & v_1300 & ~v_1301;
assign v_4127 = v_4126 & v_1307 & ~v_1308 & v_1326;
assign v_4128 = v_4126 & v_1307 & ~v_1308 & ~v_1326;
assign v_4129 = v_4126 & ~v_1309;
assign v_4130 = v_4126 & v_1317 & ~v_1318;
assign v_4131 = v_4126 & v_2014;
assign v_4133 = v_4132 & v_1307 & v_1308 & v_1323 & ~v_1324;
assign v_4135 = v_4134 & v_1330 & ~v_1331 & v_1349;
assign v_4136 = v_4134 & ~v_1332;
assign v_4137 = v_4134 & v_1340 & ~v_1341;
assign v_4138 = v_4134 & v_2022;
assign v_4140 = v_4139 & v_1330 & v_1331 & v_1346 & v_1347;
assign v_4141 = v_4134 & v_1330 & ~v_1331 & ~v_1349;
assign v_4142 = v_4139 & v_1330 & v_1331 & v_1346 & ~v_1347;
assign v_4145 = v_4143 & v_4144;
assign v_4146 = v_4143 & v_1353 & v_1354 & ~v_1355 & ~v_1356;
assign v_4147 = v_4143 & v_1353 & v_1354 & v_1355;
assign v_4148 = v_4143 & v_1353 & ~v_1354 & ~v_1358;
assign v_4150 = v_4149 & v_2035;
assign v_4151 = v_4132 & v_1307 & v_1308 & v_1323 & v_1324;
assign v_4152 = v_4124 & v_1284 & v_1285 & v_1300 & v_1301;
assign v_4154 = v_4153 & v_1365 & ~v_1366 & v_1384;
assign v_4155 = v_4153 & v_1365 & ~v_1366 & ~v_1384;
assign v_4156 = v_4153 & ~v_1367;
assign v_4157 = v_4153 & v_1375 & ~v_1376;
assign v_4158 = v_4153 & v_2044;
assign v_4160 = v_4159 & v_1365 & v_1366 & v_1381 & ~v_1382;
assign v_4162 = v_4161 & v_1388 & ~v_1389 & v_1407;
assign v_4163 = v_4161 & v_1388 & ~v_1389 & ~v_1407;
assign v_4164 = v_4161 & ~v_1390;
assign v_4165 = v_4161 & v_1398 & ~v_1399;
assign v_4166 = v_4161 & v_2053;
assign v_4168 = v_4167 & v_1388 & v_1389 & v_1404 & ~v_1405;
assign v_4170 = v_4169 & v_1411 & ~v_1412 & v_1430;
assign v_4171 = v_4169 & ~v_1413;
assign v_4172 = v_4169 & v_1421 & ~v_1422;
assign v_4173 = v_4169 & v_2061;
assign v_4175 = v_4174 & v_1411 & v_1412 & v_1427 & v_1428;
assign v_4176 = v_4169 & v_1411 & ~v_1412 & ~v_1430;
assign v_4177 = v_4174 & v_1411 & v_1412 & v_1427 & ~v_1428;
assign v_4180 = v_4178 & v_4179;
assign v_4181 = v_4178 & v_1434 & v_1435 & ~v_1436 & ~v_1437;
assign v_4182 = v_4178 & v_1434 & v_1435 & v_1436;
assign v_4183 = v_4178 & v_1434 & ~v_1435 & ~v_1439;
assign v_4185 = v_4184 & v_2074;
assign v_4186 = v_4167 & v_1388 & v_1389 & v_1404 & v_1405;
assign v_4187 = v_4159 & v_1365 & v_1366 & v_1381 & v_1382;
assign v_4189 = v_4188 & v_1446 & ~v_1447 & v_1465;
assign v_4190 = v_4188 & v_1446 & ~v_1447 & ~v_1465;
assign v_4191 = v_4188 & ~v_1448;
assign v_4192 = v_4188 & v_1456 & ~v_1457;
assign v_4193 = v_4188 & v_2083;
assign v_4195 = v_4194 & v_1446 & v_1447 & v_1462 & ~v_1463;
assign v_4197 = v_4196 & v_1469 & ~v_1470 & v_1488;
assign v_4198 = v_4196 & v_1469 & ~v_1470 & ~v_1488;
assign v_4199 = v_4196 & ~v_1471;
assign v_4200 = v_4196 & v_1479 & ~v_1480;
assign v_4201 = v_4196 & v_2092;
assign v_4203 = v_4202 & v_1469 & v_1470 & v_1485 & ~v_1486;
assign v_4205 = v_4204 & v_1492 & ~v_1493 & v_1511;
assign v_4206 = v_4204 & ~v_1494;
assign v_4207 = v_4204 & v_1502 & ~v_1503;
assign v_4208 = v_4204 & v_2100;
assign v_4210 = v_4209 & v_1492 & v_1493 & v_1508 & v_1509;
assign v_4211 = v_4204 & v_1492 & ~v_1493 & ~v_1511;
assign v_4212 = v_4209 & v_1492 & v_1493 & v_1508 & ~v_1509;
assign v_4215 = v_4213 & v_4214;
assign v_4216 = v_4213 & v_1515 & v_1516 & ~v_1517 & ~v_1518;
assign v_4217 = v_4213 & v_1515 & v_1516 & v_1517;
assign v_4218 = v_4213 & v_1515 & ~v_1516 & ~v_1520;
assign v_4220 = v_4219 & v_2113;
assign v_4221 = v_4202 & v_1469 & v_1470 & v_1485 & v_1486;
assign v_4222 = v_4194 & v_1446 & v_1447 & v_1462 & v_1463;
assign v_4225 = v_4224 & v_227;
assign v_4226 = v_4224 & ~v_227 & v_229 & v_262 & ~v_264;
assign v_4227 = v_4224 & ~v_227 & v_229 & v_262 & v_264;
assign v_4228 = v_4224 & ~v_227 & v_229 & ~v_262;
assign v_4229 = v_4224 & v_230;
assign v_4230 = v_4224 & ~v_230;
assign v_4233 = v_4231 & v_4232;
assign v_4234 = v_4231 & v_1540;
assign v_4235 = v_13037 & v_13038;
assign v_4237 = v_4236 & ~v_227 & ~v_229 & v_260;
assign v_4239 = v_4238 & v_267 & v_268;
assign v_4240 = v_4238 & v_267 & ~v_268;
assign v_4242 = v_4241 & ~v_279;
assign v_4244 = v_4241 & v_4243;
assign v_4245 = v_4241 & v_279 & v_291 & ~v_292 & v_300;
assign v_4248 = v_4246 & v_4247;
assign v_4249 = v_4246 & v_321 & v_322;
assign v_4250 = v_4246 & v_321 & ~v_322 & v_324;
assign v_4251 = v_4246 & v_321 & ~v_322 & ~v_324 & v_326;
assign v_4252 = v_4246 & v_321 & ~v_322 & ~v_324 & ~v_326;
assign v_4254 = v_4253 & v_1563;
assign v_4256 = v_4255 & ~v_308 & v_309 & v_329;
assign v_4259 = v_4257 & v_4258;
assign v_4260 = v_4257 & v_1570;
assign v_4262 = v_4261 & v_345 & v_346;
assign v_4263 = v_4261 & v_345 & ~v_346 & v_348;
assign v_4264 = v_4261 & v_345 & ~v_346 & ~v_348 & v_350;
assign v_4265 = v_4261 & v_356 & v_357;
assign v_4266 = v_4261 & v_359 & v_360;
assign v_4267 = v_4261 & v_359 & ~v_360 & v_362;
assign v_4268 = v_4261 & v_359 & ~v_360 & ~v_362 & v_364;
assign v_4269 = v_4261 & v_1582;
assign v_4271 = v_4270 & v_1585;
assign v_4273 = v_4272 & v_356 & ~v_357 & v_369 & v_370;
assign v_4274 = v_4272 & v_372 & v_373;
assign v_4275 = v_4272 & v_372 & ~v_373 & v_375;
assign v_4276 = v_4272 & v_372 & ~v_373 & ~v_375 & v_377;
assign v_4278 = v_4272 & v_4277;
assign v_4279 = v_13039 & v_13040;
assign v_4281 = v_4280 & v_384 & v_385;
assign v_4282 = v_4280 & v_384 & ~v_385;
assign v_4284 = v_4283 & v_1599;
assign v_4286 = v_13041 & v_13042;
assign v_4287 = v_4285 & v_391 & v_392;
assign v_4288 = v_4285 & v_391 & ~v_392 & v_394;
assign v_4289 = v_4285 & v_391 & ~v_392 & ~v_394 & v_396;
assign v_4290 = v_4285 & v_1606;
assign v_4292 = v_13043 & v_13044;
assign v_4294 = v_4293 & v_1611;
assign v_4296 = v_4295 & v_410 & v_411;
assign v_4297 = v_4295 & v_410 & ~v_411 & v_413;
assign v_4298 = v_4295 & v_410 & ~v_411 & ~v_413 & v_415;
assign v_4299 = v_4295 & v_421 & v_422;
assign v_4300 = v_4295 & v_424 & v_425;
assign v_4301 = v_4295 & v_424 & ~v_425 & v_427;
assign v_4302 = v_4295 & v_424 & ~v_425 & ~v_427 & v_429;
assign v_4303 = v_4295 & v_1621;
assign v_4305 = v_4304 & v_1624;
assign v_4307 = v_4306 & v_421 & ~v_422 & v_434 & v_435;
assign v_4308 = v_4306 & v_437 & v_438;
assign v_4309 = v_4306 & v_437 & ~v_438 & v_440;
assign v_4310 = v_4306 & v_437 & ~v_438 & ~v_440 & v_442;
assign v_4312 = v_4306 & v_4311;
assign v_4313 = v_13045 & v_13046;
assign v_4315 = v_4314 & v_449 & v_450;
assign v_4316 = v_4314 & v_449 & ~v_450;
assign v_4318 = v_4317 & v_1638;
assign v_4320 = v_13047 & v_13048;
assign v_4321 = v_4319 & v_456 & v_457;
assign v_4322 = v_4319 & v_456 & ~v_457 & v_459;
assign v_4323 = v_4319 & v_456 & ~v_457 & ~v_459 & v_461;
assign v_4324 = v_4319 & v_1645;
assign v_4326 = v_13049 & v_13050;
assign v_4328 = v_4327 & v_1650;
assign v_4330 = v_4329 & v_491;
assign v_4331 = v_4329 & ~v_491 & v_493 & v_526 & ~v_528;
assign v_4332 = v_4329 & ~v_491 & v_493 & v_526 & v_528;
assign v_4333 = v_4329 & ~v_491 & v_493 & ~v_526;
assign v_4334 = v_4329 & v_494;
assign v_4335 = v_4329 & ~v_494;
assign v_4338 = v_4336 & v_4337;
assign v_4339 = v_4336 & v_1666;
assign v_4340 = v_13051 & v_13052;
assign v_4342 = v_4341 & ~v_491 & ~v_493 & v_524;
assign v_4344 = v_4343 & v_531 & v_532;
assign v_4345 = v_4343 & v_531 & ~v_532;
assign v_4347 = v_4346 & v_546 & v_547;
assign v_4348 = v_4346 & v_546 & ~v_547 & ~v_551;
assign v_4350 = v_4349 & v_546 & ~v_547 & v_551;
assign v_4352 = v_4351 & v_554;
assign v_4354 = v_4353 & v_558 & v_559;
assign v_4355 = v_4353 & v_558 & ~v_559 & v_561;
assign v_4356 = v_4353 & v_1682;
assign v_4359 = v_4357 & v_4358;
assign v_4360 = v_4357 & v_1687;
assign v_4362 = v_4361 & v_588 & ~v_589 & ~v_591;
assign v_4363 = v_4361 & v_593 & ~v_594;
assign v_4364 = v_4361 & v_593 & v_594;
assign v_4365 = v_4361 & v_583;
assign v_4367 = v_4366 & v_604 & v_605;
assign v_4368 = v_4366 & v_604 & ~v_605 & ~v_609;
assign v_4370 = v_4369 & v_604 & ~v_605 & v_609;
assign v_4372 = v_4371 & v_612;
assign v_4374 = v_4373 & v_616 & v_617;
assign v_4375 = v_4373 & v_616 & ~v_617 & v_619;
assign v_4376 = v_4373 & v_1700;
assign v_4379 = v_4377 & v_4378;
assign v_4380 = v_4377 & v_1705;
assign v_4382 = v_2 & v_4381;
assign v_4383 = v_641 & v_4361;
assign v_4384 = v_643 & v_4346;
assign v_4385 = v_645 & v_4346;
assign v_4386 = v_647 & v_4346;
assign v_4387 = v_649 & v_4346;
assign v_4388 = ~v_649 & v_4329;
assign v_4390 = ~v_647 & v_4389;
assign v_4392 = ~v_645 & v_4391;
assign v_4394 = ~v_643 & v_4393;
assign v_4396 = ~v_641 & v_4395;
assign v_4398 = ~v_2 & v_4397;
assign v_4400 = v_4399 & ~v_669;
assign v_4401 = v_13053 & v_13054;
assign v_4402 = v_4399 & v_669 & v_670 & v_672 & v_674;
assign v_4403 = v_13055 & v_13056;
assign v_4405 = v_4404 & v_679 & ~v_680 & v_682;
assign v_4406 = v_4404 & v_689 & ~v_690 & ~v_692;
assign v_4407 = v_4404 & v_694 & ~v_695;
assign v_4408 = v_4404 & v_694 & v_695;
assign v_4409 = v_4404 & v_684;
assign v_4411 = v_4410 & v_1737;
assign v_4413 = v_4412 & v_1740;
assign v_4414 = v_4404 & v_679 & v_680;
assign v_4415 = v_4399 & v_1743;
assign v_4417 = v_4416 & ~v_705;
assign v_4418 = v_4416 & v_710 & v_711;
assign v_4419 = v_4416 & v_710 & ~v_711 & ~v_715;
assign v_4421 = v_4420 & v_710 & ~v_711 & v_715;
assign v_4423 = v_4422 & v_718;
assign v_4425 = v_4424 & v_705 & v_722 & v_723 & ~v_724;
assign v_4427 = v_4424 & v_4426;
assign v_4428 = v_4424 & v_750 & v_751;
assign v_4429 = v_4424 & v_750 & ~v_751;
assign v_4431 = v_4430 & v_763 & v_764;
assign v_4432 = v_4430 & v_763 & ~v_764;
assign v_4434 = v_4433 & v_745 & v_758 & v_771;
assign v_4435 = v_13057 & v_13058;
assign v_4436 = v_4424 & v_779 & v_780;
assign v_4437 = v_4424 & v_779 & ~v_780 & ~v_784;
assign v_4439 = v_4438 & v_779 & ~v_780 & v_784;
assign v_4441 = v_4440 & v_787;
assign v_4443 = v_4442 & v_1764;
assign v_4445 = v_4444 & v_798 & ~v_799 & v_817;
assign v_4446 = v_4444 & v_798 & ~v_799 & ~v_817;
assign v_4447 = v_4444 & ~v_800;
assign v_4448 = v_4444 & v_808 & ~v_809;
assign v_4449 = v_4444 & v_1771;
assign v_4451 = v_4450 & v_798 & v_799 & v_814 & ~v_815;
assign v_4453 = v_4452 & v_821 & ~v_822 & v_840;
assign v_4454 = v_4452 & v_821 & ~v_822 & ~v_840;
assign v_4455 = v_4452 & ~v_823;
assign v_4456 = v_4452 & v_831 & ~v_832;
assign v_4457 = v_4452 & v_1780;
assign v_4459 = v_4458 & v_821 & v_822 & v_837 & ~v_838;
assign v_4461 = v_4460 & v_844 & ~v_845 & v_863;
assign v_4462 = v_4460 & ~v_846;
assign v_4463 = v_4460 & v_854 & ~v_855;
assign v_4464 = v_4460 & v_1788;
assign v_4466 = v_4465 & v_844 & v_845 & v_860 & v_861;
assign v_4467 = v_4460 & v_844 & ~v_845 & ~v_863;
assign v_4468 = v_4465 & v_844 & v_845 & v_860 & ~v_861;
assign v_4471 = v_4469 & v_4470;
assign v_4472 = v_4469 & v_867 & v_868 & ~v_869 & ~v_870;
assign v_4473 = v_4469 & v_867 & v_868 & v_869;
assign v_4474 = v_4469 & v_867 & ~v_868 & ~v_872;
assign v_4476 = v_4475 & v_1801;
assign v_4477 = v_4458 & v_821 & v_822 & v_837 & v_838;
assign v_4478 = v_4450 & v_798 & v_799 & v_814 & v_815;
assign v_4480 = v_4479 & v_879 & ~v_880 & v_898;
assign v_4481 = v_4479 & v_879 & ~v_880 & ~v_898;
assign v_4482 = v_4479 & ~v_881;
assign v_4483 = v_4479 & v_889 & ~v_890;
assign v_4484 = v_4479 & v_1810;
assign v_4486 = v_4485 & v_879 & v_880 & v_895 & ~v_896;
assign v_4488 = v_4487 & v_902 & ~v_903 & v_921;
assign v_4489 = v_4487 & v_902 & ~v_903 & ~v_921;
assign v_4490 = v_4487 & ~v_904;
assign v_4491 = v_4487 & v_912 & ~v_913;
assign v_4492 = v_4487 & v_1819;
assign v_4494 = v_4493 & v_902 & v_903 & v_918 & ~v_919;
assign v_4496 = v_4495 & v_925 & ~v_926 & v_944;
assign v_4497 = v_4495 & ~v_927;
assign v_4498 = v_4495 & v_935 & ~v_936;
assign v_4499 = v_4495 & v_1827;
assign v_4501 = v_4500 & v_925 & v_926 & v_941 & v_942;
assign v_4502 = v_4495 & v_925 & ~v_926 & ~v_944;
assign v_4503 = v_4500 & v_925 & v_926 & v_941 & ~v_942;
assign v_4506 = v_4504 & v_4505;
assign v_4507 = v_4504 & v_948 & v_949 & ~v_950 & ~v_951;
assign v_4508 = v_4504 & v_948 & v_949 & v_950;
assign v_4509 = v_4504 & v_948 & ~v_949 & ~v_953;
assign v_4511 = v_4510 & v_1840;
assign v_4512 = v_4493 & v_902 & v_903 & v_918 & v_919;
assign v_4513 = v_4485 & v_879 & v_880 & v_895 & v_896;
assign v_4515 = v_4514 & v_960 & ~v_961 & v_979;
assign v_4516 = v_4514 & v_960 & ~v_961 & ~v_979;
assign v_4517 = v_4514 & ~v_962;
assign v_4518 = v_4514 & v_970 & ~v_971;
assign v_4519 = v_4514 & v_1849;
assign v_4521 = v_4520 & v_960 & v_961 & v_976 & ~v_977;
assign v_4523 = v_4522 & v_983 & ~v_984 & v_1002;
assign v_4524 = v_4522 & v_983 & ~v_984 & ~v_1002;
assign v_4525 = v_4522 & ~v_985;
assign v_4526 = v_4522 & v_993 & ~v_994;
assign v_4527 = v_4522 & v_1858;
assign v_4529 = v_4528 & v_983 & v_984 & v_999 & ~v_1000;
assign v_4531 = v_4530 & v_1006 & ~v_1007 & v_1025;
assign v_4532 = v_4530 & ~v_1008;
assign v_4533 = v_4530 & v_1016 & ~v_1017;
assign v_4534 = v_4530 & v_1866;
assign v_4536 = v_4535 & v_1006 & v_1007 & v_1022 & v_1023;
assign v_4537 = v_4530 & v_1006 & ~v_1007 & ~v_1025;
assign v_4538 = v_4535 & v_1006 & v_1007 & v_1022 & ~v_1023;
assign v_4541 = v_4539 & v_4540;
assign v_4542 = v_4539 & v_1029 & v_1030 & ~v_1031 & ~v_1032;
assign v_4543 = v_4539 & v_1029 & v_1030 & v_1031;
assign v_4544 = v_4539 & v_1029 & ~v_1030 & ~v_1034;
assign v_4546 = v_4545 & v_1879;
assign v_4547 = v_4528 & v_983 & v_984 & v_999 & v_1000;
assign v_4548 = v_4520 & v_960 & v_961 & v_976 & v_977;
assign v_4550 = v_4549 & v_1041 & ~v_1042 & v_1060;
assign v_4551 = v_4549 & v_1041 & ~v_1042 & ~v_1060;
assign v_4552 = v_4549 & ~v_1043;
assign v_4553 = v_4549 & v_1051 & ~v_1052;
assign v_4554 = v_4549 & v_1888;
assign v_4556 = v_4555 & v_1041 & v_1042 & v_1057 & ~v_1058;
assign v_4558 = v_4557 & v_1064 & ~v_1065 & v_1083;
assign v_4559 = v_4557 & v_1064 & ~v_1065 & ~v_1083;
assign v_4560 = v_4557 & ~v_1066;
assign v_4561 = v_4557 & v_1074 & ~v_1075;
assign v_4562 = v_4557 & v_1897;
assign v_4564 = v_4563 & v_1064 & v_1065 & v_1080 & ~v_1081;
assign v_4566 = v_4565 & v_1087 & ~v_1088 & v_1106;
assign v_4567 = v_4565 & ~v_1089;
assign v_4568 = v_4565 & v_1097 & ~v_1098;
assign v_4569 = v_4565 & v_1905;
assign v_4571 = v_4570 & v_1087 & v_1088 & v_1103 & v_1104;
assign v_4572 = v_4565 & v_1087 & ~v_1088 & ~v_1106;
assign v_4573 = v_4570 & v_1087 & v_1088 & v_1103 & ~v_1104;
assign v_4576 = v_4574 & v_4575;
assign v_4577 = v_4574 & v_1110 & v_1111 & ~v_1112 & ~v_1113;
assign v_4578 = v_4574 & v_1110 & v_1111 & v_1112;
assign v_4579 = v_4574 & v_1110 & ~v_1111 & ~v_1115;
assign v_4581 = v_4580 & v_1918;
assign v_4582 = v_4563 & v_1064 & v_1065 & v_1080 & v_1081;
assign v_4583 = v_4555 & v_1041 & v_1042 & v_1057 & v_1058;
assign v_4585 = v_4584 & v_1122 & ~v_1123 & v_1141;
assign v_4586 = v_4584 & v_1122 & ~v_1123 & ~v_1141;
assign v_4587 = v_4584 & ~v_1124;
assign v_4588 = v_4584 & v_1132 & ~v_1133;
assign v_4589 = v_4584 & v_1927;
assign v_4591 = v_4590 & v_1122 & v_1123 & v_1138 & ~v_1139;
assign v_4593 = v_4592 & v_1145 & ~v_1146 & v_1164;
assign v_4594 = v_4592 & v_1145 & ~v_1146 & ~v_1164;
assign v_4595 = v_4592 & ~v_1147;
assign v_4596 = v_4592 & v_1155 & ~v_1156;
assign v_4597 = v_4592 & v_1936;
assign v_4599 = v_4598 & v_1145 & v_1146 & v_1161 & ~v_1162;
assign v_4601 = v_4600 & v_1168 & ~v_1169 & v_1187;
assign v_4602 = v_4600 & ~v_1170;
assign v_4603 = v_4600 & v_1178 & ~v_1179;
assign v_4604 = v_4600 & v_1944;
assign v_4606 = v_4605 & v_1168 & v_1169 & v_1184 & v_1185;
assign v_4607 = v_4600 & v_1168 & ~v_1169 & ~v_1187;
assign v_4608 = v_4605 & v_1168 & v_1169 & v_1184 & ~v_1185;
assign v_4611 = v_4609 & v_4610;
assign v_4612 = v_4609 & v_1191 & v_1192 & ~v_1193 & ~v_1194;
assign v_4613 = v_4609 & v_1191 & v_1192 & v_1193;
assign v_4614 = v_4609 & v_1191 & ~v_1192 & ~v_1196;
assign v_4616 = v_4615 & v_1957;
assign v_4617 = v_4598 & v_1145 & v_1146 & v_1161 & v_1162;
assign v_4618 = v_4590 & v_1122 & v_1123 & v_1138 & v_1139;
assign v_4620 = v_4619 & v_1203 & ~v_1204 & v_1222;
assign v_4621 = v_4619 & v_1203 & ~v_1204 & ~v_1222;
assign v_4622 = v_4619 & ~v_1205;
assign v_4623 = v_4619 & v_1213 & ~v_1214;
assign v_4624 = v_4619 & v_1966;
assign v_4626 = v_4625 & v_1203 & v_1204 & v_1219 & ~v_1220;
assign v_4628 = v_4627 & v_1226 & ~v_1227 & v_1245;
assign v_4629 = v_4627 & v_1226 & ~v_1227 & ~v_1245;
assign v_4630 = v_4627 & ~v_1228;
assign v_4631 = v_4627 & v_1236 & ~v_1237;
assign v_4632 = v_4627 & v_1975;
assign v_4634 = v_4633 & v_1226 & v_1227 & v_1242 & ~v_1243;
assign v_4636 = v_4635 & v_1249 & ~v_1250 & v_1268;
assign v_4637 = v_4635 & ~v_1251;
assign v_4638 = v_4635 & v_1259 & ~v_1260;
assign v_4639 = v_4635 & v_1983;
assign v_4641 = v_4640 & v_1249 & v_1250 & v_1265 & v_1266;
assign v_4642 = v_4635 & v_1249 & ~v_1250 & ~v_1268;
assign v_4643 = v_4640 & v_1249 & v_1250 & v_1265 & ~v_1266;
assign v_4646 = v_4644 & v_4645;
assign v_4647 = v_4644 & v_1272 & v_1273 & ~v_1274 & ~v_1275;
assign v_4648 = v_4644 & v_1272 & v_1273 & v_1274;
assign v_4649 = v_4644 & v_1272 & ~v_1273 & ~v_1277;
assign v_4651 = v_4650 & v_1996;
assign v_4652 = v_4633 & v_1226 & v_1227 & v_1242 & v_1243;
assign v_4653 = v_4625 & v_1203 & v_1204 & v_1219 & v_1220;
assign v_4655 = v_4654 & v_1284 & ~v_1285 & v_1303;
assign v_4656 = v_4654 & v_1284 & ~v_1285 & ~v_1303;
assign v_4657 = v_4654 & ~v_1286;
assign v_4658 = v_4654 & v_1294 & ~v_1295;
assign v_4659 = v_4654 & v_2005;
assign v_4661 = v_4660 & v_1284 & v_1285 & v_1300 & ~v_1301;
assign v_4663 = v_4662 & v_1307 & ~v_1308 & v_1326;
assign v_4664 = v_4662 & v_1307 & ~v_1308 & ~v_1326;
assign v_4665 = v_4662 & ~v_1309;
assign v_4666 = v_4662 & v_1317 & ~v_1318;
assign v_4667 = v_4662 & v_2014;
assign v_4669 = v_4668 & v_1307 & v_1308 & v_1323 & ~v_1324;
assign v_4671 = v_4670 & v_1330 & ~v_1331 & v_1349;
assign v_4672 = v_4670 & ~v_1332;
assign v_4673 = v_4670 & v_1340 & ~v_1341;
assign v_4674 = v_4670 & v_2022;
assign v_4676 = v_4675 & v_1330 & v_1331 & v_1346 & v_1347;
assign v_4677 = v_4670 & v_1330 & ~v_1331 & ~v_1349;
assign v_4678 = v_4675 & v_1330 & v_1331 & v_1346 & ~v_1347;
assign v_4681 = v_4679 & v_4680;
assign v_4682 = v_4679 & v_1353 & v_1354 & ~v_1355 & ~v_1356;
assign v_4683 = v_4679 & v_1353 & v_1354 & v_1355;
assign v_4684 = v_4679 & v_1353 & ~v_1354 & ~v_1358;
assign v_4686 = v_4685 & v_2035;
assign v_4687 = v_4668 & v_1307 & v_1308 & v_1323 & v_1324;
assign v_4688 = v_4660 & v_1284 & v_1285 & v_1300 & v_1301;
assign v_4690 = v_4689 & v_1365 & ~v_1366 & v_1384;
assign v_4691 = v_4689 & v_1365 & ~v_1366 & ~v_1384;
assign v_4692 = v_4689 & ~v_1367;
assign v_4693 = v_4689 & v_1375 & ~v_1376;
assign v_4694 = v_4689 & v_2044;
assign v_4696 = v_4695 & v_1365 & v_1366 & v_1381 & ~v_1382;
assign v_4698 = v_4697 & v_1388 & ~v_1389 & v_1407;
assign v_4699 = v_4697 & v_1388 & ~v_1389 & ~v_1407;
assign v_4700 = v_4697 & ~v_1390;
assign v_4701 = v_4697 & v_1398 & ~v_1399;
assign v_4702 = v_4697 & v_2053;
assign v_4704 = v_4703 & v_1388 & v_1389 & v_1404 & ~v_1405;
assign v_4706 = v_4705 & v_1411 & ~v_1412 & v_1430;
assign v_4707 = v_4705 & ~v_1413;
assign v_4708 = v_4705 & v_1421 & ~v_1422;
assign v_4709 = v_4705 & v_2061;
assign v_4711 = v_4710 & v_1411 & v_1412 & v_1427 & v_1428;
assign v_4712 = v_4705 & v_1411 & ~v_1412 & ~v_1430;
assign v_4713 = v_4710 & v_1411 & v_1412 & v_1427 & ~v_1428;
assign v_4716 = v_4714 & v_4715;
assign v_4717 = v_4714 & v_1434 & v_1435 & ~v_1436 & ~v_1437;
assign v_4718 = v_4714 & v_1434 & v_1435 & v_1436;
assign v_4719 = v_4714 & v_1434 & ~v_1435 & ~v_1439;
assign v_4721 = v_4720 & v_2074;
assign v_4722 = v_4703 & v_1388 & v_1389 & v_1404 & v_1405;
assign v_4723 = v_4695 & v_1365 & v_1366 & v_1381 & v_1382;
assign v_4725 = v_4724 & v_1446 & ~v_1447 & v_1465;
assign v_4726 = v_4724 & v_1446 & ~v_1447 & ~v_1465;
assign v_4727 = v_4724 & ~v_1448;
assign v_4728 = v_4724 & v_1456 & ~v_1457;
assign v_4729 = v_4724 & v_2083;
assign v_4731 = v_4730 & v_1446 & v_1447 & v_1462 & ~v_1463;
assign v_4733 = v_4732 & v_1469 & ~v_1470 & v_1488;
assign v_4734 = v_4732 & v_1469 & ~v_1470 & ~v_1488;
assign v_4735 = v_4732 & ~v_1471;
assign v_4736 = v_4732 & v_1479 & ~v_1480;
assign v_4737 = v_4732 & v_2092;
assign v_4739 = v_4738 & v_1469 & v_1470 & v_1485 & ~v_1486;
assign v_4741 = v_4740 & v_1492 & ~v_1493 & v_1511;
assign v_4742 = v_4740 & ~v_1494;
assign v_4743 = v_4740 & v_1502 & ~v_1503;
assign v_4744 = v_4740 & v_2100;
assign v_4746 = v_4745 & v_1492 & v_1493 & v_1508 & v_1509;
assign v_4747 = v_4740 & v_1492 & ~v_1493 & ~v_1511;
assign v_4748 = v_4745 & v_1492 & v_1493 & v_1508 & ~v_1509;
assign v_4751 = v_4749 & v_4750;
assign v_4752 = v_4749 & v_1515 & v_1516 & ~v_1517 & ~v_1518;
assign v_4753 = v_4749 & v_1515 & v_1516 & v_1517;
assign v_4754 = v_4749 & v_1515 & ~v_1516 & ~v_1520;
assign v_4756 = v_4755 & v_2113;
assign v_4757 = v_4738 & v_1469 & v_1470 & v_1485 & v_1486;
assign v_4758 = v_4730 & v_1446 & v_1447 & v_1462 & v_1463;
assign v_4760 = v_7 & v_227;
assign v_4761 = v_7 & ~v_227 & v_229 & v_262 & ~v_264;
assign v_4762 = v_7 & ~v_227 & v_229 & v_262 & v_264;
assign v_4763 = v_7 & ~v_227 & v_229 & ~v_262;
assign v_4764 = v_7 & v_230;
assign v_4765 = v_7 & ~v_230;
assign v_4768 = v_4766 & v_4767;
assign v_4769 = v_4766 & v_1540;
assign v_4770 = v_13059 & v_13060;
assign v_4772 = v_4771 & ~v_227 & ~v_229 & v_260;
assign v_4774 = v_4773 & v_267 & v_268;
assign v_4775 = v_4773 & v_267 & ~v_268;
assign v_4777 = v_4776 & ~v_279;
assign v_4779 = v_4776 & v_4778;
assign v_4780 = v_4776 & v_279 & v_291 & ~v_292 & v_300;
assign v_4783 = v_4781 & v_4782;
assign v_4784 = v_4781 & v_321 & v_322;
assign v_4785 = v_4781 & v_321 & ~v_322 & v_324;
assign v_4786 = v_4781 & v_321 & ~v_322 & ~v_324 & v_326;
assign v_4787 = v_4781 & v_321 & ~v_322 & ~v_324 & ~v_326;
assign v_4789 = v_4788 & v_1563;
assign v_4791 = v_4790 & ~v_308 & v_309 & v_329;
assign v_4794 = v_4792 & v_4793;
assign v_4795 = v_4792 & v_1570;
assign v_4797 = v_4796 & v_345 & v_346;
assign v_4798 = v_4796 & v_345 & ~v_346 & v_348;
assign v_4799 = v_4796 & v_345 & ~v_346 & ~v_348 & v_350;
assign v_4800 = v_4796 & v_356 & v_357;
assign v_4801 = v_4796 & v_359 & v_360;
assign v_4802 = v_4796 & v_359 & ~v_360 & v_362;
assign v_4803 = v_4796 & v_359 & ~v_360 & ~v_362 & v_364;
assign v_4804 = v_4796 & v_1582;
assign v_4806 = v_4805 & v_1585;
assign v_4808 = v_4807 & v_356 & ~v_357 & v_369 & v_370;
assign v_4809 = v_4807 & v_372 & v_373;
assign v_4810 = v_4807 & v_372 & ~v_373 & v_375;
assign v_4811 = v_4807 & v_372 & ~v_373 & ~v_375 & v_377;
assign v_4813 = v_4807 & v_4812;
assign v_4814 = v_13061 & v_13062;
assign v_4816 = v_4815 & v_384 & v_385;
assign v_4817 = v_4815 & v_384 & ~v_385;
assign v_4819 = v_4818 & v_1599;
assign v_4821 = v_13063 & v_13064;
assign v_4822 = v_4820 & v_391 & v_392;
assign v_4823 = v_4820 & v_391 & ~v_392 & v_394;
assign v_4824 = v_4820 & v_391 & ~v_392 & ~v_394 & v_396;
assign v_4825 = v_4820 & v_1606;
assign v_4827 = v_13065 & v_13066;
assign v_4829 = v_4828 & v_1611;
assign v_4831 = v_4830 & v_410 & v_411;
assign v_4832 = v_4830 & v_410 & ~v_411 & v_413;
assign v_4833 = v_4830 & v_410 & ~v_411 & ~v_413 & v_415;
assign v_4834 = v_4830 & v_421 & v_422;
assign v_4835 = v_4830 & v_424 & v_425;
assign v_4836 = v_4830 & v_424 & ~v_425 & v_427;
assign v_4837 = v_4830 & v_424 & ~v_425 & ~v_427 & v_429;
assign v_4838 = v_4830 & v_1621;
assign v_4840 = v_4839 & v_1624;
assign v_4842 = v_4841 & v_421 & ~v_422 & v_434 & v_435;
assign v_4843 = v_4841 & v_437 & v_438;
assign v_4844 = v_4841 & v_437 & ~v_438 & v_440;
assign v_4845 = v_4841 & v_437 & ~v_438 & ~v_440 & v_442;
assign v_4847 = v_4841 & v_4846;
assign v_4848 = v_13067 & v_13068;
assign v_4850 = v_4849 & v_449 & v_450;
assign v_4851 = v_4849 & v_449 & ~v_450;
assign v_4853 = v_4852 & v_1638;
assign v_4855 = v_13069 & v_13070;
assign v_4856 = v_4854 & v_456 & v_457;
assign v_4857 = v_4854 & v_456 & ~v_457 & v_459;
assign v_4858 = v_4854 & v_456 & ~v_457 & ~v_459 & v_461;
assign v_4859 = v_4854 & v_1645;
assign v_4861 = v_13071 & v_13072;
assign v_4863 = v_4862 & v_1650;
assign v_4865 = v_4864 & v_491;
assign v_4866 = v_4864 & ~v_491 & v_493 & v_526 & ~v_528;
assign v_4867 = v_4864 & ~v_491 & v_493 & v_526 & v_528;
assign v_4868 = v_4864 & ~v_491 & v_493 & ~v_526;
assign v_4869 = v_4864 & v_494;
assign v_4870 = v_4864 & ~v_494;
assign v_4873 = v_4871 & v_4872;
assign v_4874 = v_4871 & v_1666;
assign v_4875 = v_13073 & v_13074;
assign v_4877 = v_4876 & ~v_491 & ~v_493 & v_524;
assign v_4879 = v_4878 & v_531 & v_532;
assign v_4880 = v_4878 & v_531 & ~v_532;
assign v_4882 = v_4881 & v_546 & v_547;
assign v_4883 = v_4881 & v_546 & ~v_547 & ~v_551;
assign v_4885 = v_4884 & v_546 & ~v_547 & v_551;
assign v_4887 = v_4886 & v_554;
assign v_4889 = v_4888 & v_558 & v_559;
assign v_4890 = v_4888 & v_558 & ~v_559 & v_561;
assign v_4891 = v_4888 & v_1682;
assign v_4894 = v_4892 & v_4893;
assign v_4895 = v_4892 & v_1687;
assign v_4897 = v_4896 & v_588 & ~v_589 & ~v_591;
assign v_4898 = v_4896 & v_593 & ~v_594;
assign v_4899 = v_4896 & v_593 & v_594;
assign v_4900 = v_4896 & v_583;
assign v_4902 = v_4901 & v_604 & v_605;
assign v_4903 = v_4901 & v_604 & ~v_605 & ~v_609;
assign v_4905 = v_4904 & v_604 & ~v_605 & v_609;
assign v_4907 = v_4906 & v_612;
assign v_4909 = v_4908 & v_616 & v_617;
assign v_4910 = v_4908 & v_616 & ~v_617 & v_619;
assign v_4911 = v_4908 & v_1700;
assign v_4914 = v_4912 & v_4913;
assign v_4915 = v_4912 & v_1705;
assign v_4917 = v_2 & v_4916;
assign v_4918 = v_641 & v_4896;
assign v_4919 = v_643 & v_4881;
assign v_4920 = v_645 & v_4881;
assign v_4921 = v_647 & v_4881;
assign v_4922 = v_649 & v_4881;
assign v_4923 = ~v_649 & v_4864;
assign v_4925 = ~v_647 & v_4924;
assign v_4927 = ~v_645 & v_4926;
assign v_4929 = ~v_643 & v_4928;
assign v_4931 = ~v_641 & v_4930;
assign v_4933 = ~v_2 & v_4932;
assign v_4935 = v_4934 & ~v_669;
assign v_4936 = v_13075 & v_13076;
assign v_4937 = v_4934 & v_669 & v_670 & v_672 & v_674;
assign v_4938 = v_13077 & v_13078;
assign v_4940 = v_4939 & v_679 & ~v_680 & v_682;
assign v_4941 = v_4939 & v_689 & ~v_690 & ~v_692;
assign v_4942 = v_4939 & v_694 & ~v_695;
assign v_4943 = v_4939 & v_694 & v_695;
assign v_4944 = v_4939 & v_684;
assign v_4946 = v_4945 & v_1737;
assign v_4948 = v_4947 & v_1740;
assign v_4949 = v_4939 & v_679 & v_680;
assign v_4950 = v_4934 & v_1743;
assign v_4952 = v_4951 & ~v_705;
assign v_4953 = v_4951 & v_710 & v_711;
assign v_4954 = v_4951 & v_710 & ~v_711 & ~v_715;
assign v_4956 = v_4955 & v_710 & ~v_711 & v_715;
assign v_4958 = v_4957 & v_718;
assign v_4960 = v_4959 & v_705 & v_722 & v_723 & ~v_724;
assign v_4962 = v_4959 & v_4961;
assign v_4963 = v_4959 & v_750 & v_751;
assign v_4964 = v_4959 & v_750 & ~v_751;
assign v_4966 = v_4965 & v_763 & v_764;
assign v_4967 = v_4965 & v_763 & ~v_764;
assign v_4969 = v_4968 & v_745 & v_758 & v_771;
assign v_4970 = v_13079 & v_13080;
assign v_4971 = v_4959 & v_779 & v_780;
assign v_4972 = v_4959 & v_779 & ~v_780 & ~v_784;
assign v_4974 = v_4973 & v_779 & ~v_780 & v_784;
assign v_4976 = v_4975 & v_787;
assign v_4978 = v_4977 & v_1764;
assign v_4980 = v_4979 & v_798 & ~v_799 & v_817;
assign v_4981 = v_4979 & v_798 & ~v_799 & ~v_817;
assign v_4982 = v_4979 & ~v_800;
assign v_4983 = v_4979 & v_808 & ~v_809;
assign v_4984 = v_4979 & v_1771;
assign v_4986 = v_4985 & v_798 & v_799 & v_814 & ~v_815;
assign v_4988 = v_4987 & v_821 & ~v_822 & v_840;
assign v_4989 = v_4987 & v_821 & ~v_822 & ~v_840;
assign v_4990 = v_4987 & ~v_823;
assign v_4991 = v_4987 & v_831 & ~v_832;
assign v_4992 = v_4987 & v_1780;
assign v_4994 = v_4993 & v_821 & v_822 & v_837 & ~v_838;
assign v_4996 = v_4995 & v_844 & ~v_845 & v_863;
assign v_4997 = v_4995 & ~v_846;
assign v_4998 = v_4995 & v_854 & ~v_855;
assign v_4999 = v_4995 & v_1788;
assign v_5001 = v_5000 & v_844 & v_845 & v_860 & v_861;
assign v_5002 = v_4995 & v_844 & ~v_845 & ~v_863;
assign v_5003 = v_5000 & v_844 & v_845 & v_860 & ~v_861;
assign v_5006 = v_5004 & v_5005;
assign v_5007 = v_5004 & v_867 & v_868 & ~v_869 & ~v_870;
assign v_5008 = v_5004 & v_867 & v_868 & v_869;
assign v_5009 = v_5004 & v_867 & ~v_868 & ~v_872;
assign v_5011 = v_5010 & v_1801;
assign v_5012 = v_4993 & v_821 & v_822 & v_837 & v_838;
assign v_5013 = v_4985 & v_798 & v_799 & v_814 & v_815;
assign v_5015 = v_5014 & v_879 & ~v_880 & v_898;
assign v_5016 = v_5014 & v_879 & ~v_880 & ~v_898;
assign v_5017 = v_5014 & ~v_881;
assign v_5018 = v_5014 & v_889 & ~v_890;
assign v_5019 = v_5014 & v_1810;
assign v_5021 = v_5020 & v_879 & v_880 & v_895 & ~v_896;
assign v_5023 = v_5022 & v_902 & ~v_903 & v_921;
assign v_5024 = v_5022 & v_902 & ~v_903 & ~v_921;
assign v_5025 = v_5022 & ~v_904;
assign v_5026 = v_5022 & v_912 & ~v_913;
assign v_5027 = v_5022 & v_1819;
assign v_5029 = v_5028 & v_902 & v_903 & v_918 & ~v_919;
assign v_5031 = v_5030 & v_925 & ~v_926 & v_944;
assign v_5032 = v_5030 & ~v_927;
assign v_5033 = v_5030 & v_935 & ~v_936;
assign v_5034 = v_5030 & v_1827;
assign v_5036 = v_5035 & v_925 & v_926 & v_941 & v_942;
assign v_5037 = v_5030 & v_925 & ~v_926 & ~v_944;
assign v_5038 = v_5035 & v_925 & v_926 & v_941 & ~v_942;
assign v_5041 = v_5039 & v_5040;
assign v_5042 = v_5039 & v_948 & v_949 & ~v_950 & ~v_951;
assign v_5043 = v_5039 & v_948 & v_949 & v_950;
assign v_5044 = v_5039 & v_948 & ~v_949 & ~v_953;
assign v_5046 = v_5045 & v_1840;
assign v_5047 = v_5028 & v_902 & v_903 & v_918 & v_919;
assign v_5048 = v_5020 & v_879 & v_880 & v_895 & v_896;
assign v_5050 = v_5049 & v_960 & ~v_961 & v_979;
assign v_5051 = v_5049 & v_960 & ~v_961 & ~v_979;
assign v_5052 = v_5049 & ~v_962;
assign v_5053 = v_5049 & v_970 & ~v_971;
assign v_5054 = v_5049 & v_1849;
assign v_5056 = v_5055 & v_960 & v_961 & v_976 & ~v_977;
assign v_5058 = v_5057 & v_983 & ~v_984 & v_1002;
assign v_5059 = v_5057 & v_983 & ~v_984 & ~v_1002;
assign v_5060 = v_5057 & ~v_985;
assign v_5061 = v_5057 & v_993 & ~v_994;
assign v_5062 = v_5057 & v_1858;
assign v_5064 = v_5063 & v_983 & v_984 & v_999 & ~v_1000;
assign v_5066 = v_5065 & v_1006 & ~v_1007 & v_1025;
assign v_5067 = v_5065 & ~v_1008;
assign v_5068 = v_5065 & v_1016 & ~v_1017;
assign v_5069 = v_5065 & v_1866;
assign v_5071 = v_5070 & v_1006 & v_1007 & v_1022 & v_1023;
assign v_5072 = v_5065 & v_1006 & ~v_1007 & ~v_1025;
assign v_5073 = v_5070 & v_1006 & v_1007 & v_1022 & ~v_1023;
assign v_5076 = v_5074 & v_5075;
assign v_5077 = v_5074 & v_1029 & v_1030 & ~v_1031 & ~v_1032;
assign v_5078 = v_5074 & v_1029 & v_1030 & v_1031;
assign v_5079 = v_5074 & v_1029 & ~v_1030 & ~v_1034;
assign v_5081 = v_5080 & v_1879;
assign v_5082 = v_5063 & v_983 & v_984 & v_999 & v_1000;
assign v_5083 = v_5055 & v_960 & v_961 & v_976 & v_977;
assign v_5085 = v_5084 & v_1041 & ~v_1042 & v_1060;
assign v_5086 = v_5084 & v_1041 & ~v_1042 & ~v_1060;
assign v_5087 = v_5084 & ~v_1043;
assign v_5088 = v_5084 & v_1051 & ~v_1052;
assign v_5089 = v_5084 & v_1888;
assign v_5091 = v_5090 & v_1041 & v_1042 & v_1057 & ~v_1058;
assign v_5093 = v_5092 & v_1064 & ~v_1065 & v_1083;
assign v_5094 = v_5092 & v_1064 & ~v_1065 & ~v_1083;
assign v_5095 = v_5092 & ~v_1066;
assign v_5096 = v_5092 & v_1074 & ~v_1075;
assign v_5097 = v_5092 & v_1897;
assign v_5099 = v_5098 & v_1064 & v_1065 & v_1080 & ~v_1081;
assign v_5101 = v_5100 & v_1087 & ~v_1088 & v_1106;
assign v_5102 = v_5100 & ~v_1089;
assign v_5103 = v_5100 & v_1097 & ~v_1098;
assign v_5104 = v_5100 & v_1905;
assign v_5106 = v_5105 & v_1087 & v_1088 & v_1103 & v_1104;
assign v_5107 = v_5100 & v_1087 & ~v_1088 & ~v_1106;
assign v_5108 = v_5105 & v_1087 & v_1088 & v_1103 & ~v_1104;
assign v_5111 = v_5109 & v_5110;
assign v_5112 = v_5109 & v_1110 & v_1111 & ~v_1112 & ~v_1113;
assign v_5113 = v_5109 & v_1110 & v_1111 & v_1112;
assign v_5114 = v_5109 & v_1110 & ~v_1111 & ~v_1115;
assign v_5116 = v_5115 & v_1918;
assign v_5117 = v_5098 & v_1064 & v_1065 & v_1080 & v_1081;
assign v_5118 = v_5090 & v_1041 & v_1042 & v_1057 & v_1058;
assign v_5120 = v_5119 & v_1122 & ~v_1123 & v_1141;
assign v_5121 = v_5119 & v_1122 & ~v_1123 & ~v_1141;
assign v_5122 = v_5119 & ~v_1124;
assign v_5123 = v_5119 & v_1132 & ~v_1133;
assign v_5124 = v_5119 & v_1927;
assign v_5126 = v_5125 & v_1122 & v_1123 & v_1138 & ~v_1139;
assign v_5128 = v_5127 & v_1145 & ~v_1146 & v_1164;
assign v_5129 = v_5127 & v_1145 & ~v_1146 & ~v_1164;
assign v_5130 = v_5127 & ~v_1147;
assign v_5131 = v_5127 & v_1155 & ~v_1156;
assign v_5132 = v_5127 & v_1936;
assign v_5134 = v_5133 & v_1145 & v_1146 & v_1161 & ~v_1162;
assign v_5136 = v_5135 & v_1168 & ~v_1169 & v_1187;
assign v_5137 = v_5135 & ~v_1170;
assign v_5138 = v_5135 & v_1178 & ~v_1179;
assign v_5139 = v_5135 & v_1944;
assign v_5141 = v_5140 & v_1168 & v_1169 & v_1184 & v_1185;
assign v_5142 = v_5135 & v_1168 & ~v_1169 & ~v_1187;
assign v_5143 = v_5140 & v_1168 & v_1169 & v_1184 & ~v_1185;
assign v_5146 = v_5144 & v_5145;
assign v_5147 = v_5144 & v_1191 & v_1192 & ~v_1193 & ~v_1194;
assign v_5148 = v_5144 & v_1191 & v_1192 & v_1193;
assign v_5149 = v_5144 & v_1191 & ~v_1192 & ~v_1196;
assign v_5151 = v_5150 & v_1957;
assign v_5152 = v_5133 & v_1145 & v_1146 & v_1161 & v_1162;
assign v_5153 = v_5125 & v_1122 & v_1123 & v_1138 & v_1139;
assign v_5155 = v_5154 & v_1203 & ~v_1204 & v_1222;
assign v_5156 = v_5154 & v_1203 & ~v_1204 & ~v_1222;
assign v_5157 = v_5154 & ~v_1205;
assign v_5158 = v_5154 & v_1213 & ~v_1214;
assign v_5159 = v_5154 & v_1966;
assign v_5161 = v_5160 & v_1203 & v_1204 & v_1219 & ~v_1220;
assign v_5163 = v_5162 & v_1226 & ~v_1227 & v_1245;
assign v_5164 = v_5162 & v_1226 & ~v_1227 & ~v_1245;
assign v_5165 = v_5162 & ~v_1228;
assign v_5166 = v_5162 & v_1236 & ~v_1237;
assign v_5167 = v_5162 & v_1975;
assign v_5169 = v_5168 & v_1226 & v_1227 & v_1242 & ~v_1243;
assign v_5171 = v_5170 & v_1249 & ~v_1250 & v_1268;
assign v_5172 = v_5170 & ~v_1251;
assign v_5173 = v_5170 & v_1259 & ~v_1260;
assign v_5174 = v_5170 & v_1983;
assign v_5176 = v_5175 & v_1249 & v_1250 & v_1265 & v_1266;
assign v_5177 = v_5170 & v_1249 & ~v_1250 & ~v_1268;
assign v_5178 = v_5175 & v_1249 & v_1250 & v_1265 & ~v_1266;
assign v_5181 = v_5179 & v_5180;
assign v_5182 = v_5179 & v_1272 & v_1273 & ~v_1274 & ~v_1275;
assign v_5183 = v_5179 & v_1272 & v_1273 & v_1274;
assign v_5184 = v_5179 & v_1272 & ~v_1273 & ~v_1277;
assign v_5186 = v_5185 & v_1996;
assign v_5187 = v_5168 & v_1226 & v_1227 & v_1242 & v_1243;
assign v_5188 = v_5160 & v_1203 & v_1204 & v_1219 & v_1220;
assign v_5190 = v_5189 & v_1284 & ~v_1285 & v_1303;
assign v_5191 = v_5189 & v_1284 & ~v_1285 & ~v_1303;
assign v_5192 = v_5189 & ~v_1286;
assign v_5193 = v_5189 & v_1294 & ~v_1295;
assign v_5194 = v_5189 & v_2005;
assign v_5196 = v_5195 & v_1284 & v_1285 & v_1300 & ~v_1301;
assign v_5198 = v_5197 & v_1307 & ~v_1308 & v_1326;
assign v_5199 = v_5197 & v_1307 & ~v_1308 & ~v_1326;
assign v_5200 = v_5197 & ~v_1309;
assign v_5201 = v_5197 & v_1317 & ~v_1318;
assign v_5202 = v_5197 & v_2014;
assign v_5204 = v_5203 & v_1307 & v_1308 & v_1323 & ~v_1324;
assign v_5206 = v_5205 & v_1330 & ~v_1331 & v_1349;
assign v_5207 = v_5205 & ~v_1332;
assign v_5208 = v_5205 & v_1340 & ~v_1341;
assign v_5209 = v_5205 & v_2022;
assign v_5211 = v_5210 & v_1330 & v_1331 & v_1346 & v_1347;
assign v_5212 = v_5205 & v_1330 & ~v_1331 & ~v_1349;
assign v_5213 = v_5210 & v_1330 & v_1331 & v_1346 & ~v_1347;
assign v_5216 = v_5214 & v_5215;
assign v_5217 = v_5214 & v_1353 & v_1354 & ~v_1355 & ~v_1356;
assign v_5218 = v_5214 & v_1353 & v_1354 & v_1355;
assign v_5219 = v_5214 & v_1353 & ~v_1354 & ~v_1358;
assign v_5221 = v_5220 & v_2035;
assign v_5222 = v_5203 & v_1307 & v_1308 & v_1323 & v_1324;
assign v_5223 = v_5195 & v_1284 & v_1285 & v_1300 & v_1301;
assign v_5225 = v_5224 & v_1365 & ~v_1366 & v_1384;
assign v_5226 = v_5224 & v_1365 & ~v_1366 & ~v_1384;
assign v_5227 = v_5224 & ~v_1367;
assign v_5228 = v_5224 & v_1375 & ~v_1376;
assign v_5229 = v_5224 & v_2044;
assign v_5231 = v_5230 & v_1365 & v_1366 & v_1381 & ~v_1382;
assign v_5233 = v_5232 & v_1388 & ~v_1389 & v_1407;
assign v_5234 = v_5232 & v_1388 & ~v_1389 & ~v_1407;
assign v_5235 = v_5232 & ~v_1390;
assign v_5236 = v_5232 & v_1398 & ~v_1399;
assign v_5237 = v_5232 & v_2053;
assign v_5239 = v_5238 & v_1388 & v_1389 & v_1404 & ~v_1405;
assign v_5241 = v_5240 & v_1411 & ~v_1412 & v_1430;
assign v_5242 = v_5240 & ~v_1413;
assign v_5243 = v_5240 & v_1421 & ~v_1422;
assign v_5244 = v_5240 & v_2061;
assign v_5246 = v_5245 & v_1411 & v_1412 & v_1427 & v_1428;
assign v_5247 = v_5240 & v_1411 & ~v_1412 & ~v_1430;
assign v_5248 = v_5245 & v_1411 & v_1412 & v_1427 & ~v_1428;
assign v_5251 = v_5249 & v_5250;
assign v_5252 = v_5249 & v_1434 & v_1435 & ~v_1436 & ~v_1437;
assign v_5253 = v_5249 & v_1434 & v_1435 & v_1436;
assign v_5254 = v_5249 & v_1434 & ~v_1435 & ~v_1439;
assign v_5256 = v_5255 & v_2074;
assign v_5257 = v_5238 & v_1388 & v_1389 & v_1404 & v_1405;
assign v_5258 = v_5230 & v_1365 & v_1366 & v_1381 & v_1382;
assign v_5260 = v_5259 & v_1446 & ~v_1447 & v_1465;
assign v_5261 = v_5259 & v_1446 & ~v_1447 & ~v_1465;
assign v_5262 = v_5259 & ~v_1448;
assign v_5263 = v_5259 & v_1456 & ~v_1457;
assign v_5264 = v_5259 & v_2083;
assign v_5266 = v_5265 & v_1446 & v_1447 & v_1462 & ~v_1463;
assign v_5268 = v_5267 & v_1469 & ~v_1470 & v_1488;
assign v_5269 = v_5267 & v_1469 & ~v_1470 & ~v_1488;
assign v_5270 = v_5267 & ~v_1471;
assign v_5271 = v_5267 & v_1479 & ~v_1480;
assign v_5272 = v_5267 & v_2092;
assign v_5274 = v_5273 & v_1469 & v_1470 & v_1485 & ~v_1486;
assign v_5276 = v_5275 & v_1492 & ~v_1493 & v_1511;
assign v_5277 = v_5275 & ~v_1494;
assign v_5278 = v_5275 & v_1502 & ~v_1503;
assign v_5279 = v_5275 & v_2100;
assign v_5281 = v_5280 & v_1492 & v_1493 & v_1508 & v_1509;
assign v_5282 = v_5275 & v_1492 & ~v_1493 & ~v_1511;
assign v_5283 = v_5280 & v_1492 & v_1493 & v_1508 & ~v_1509;
assign v_5286 = v_5284 & v_5285;
assign v_5287 = v_5284 & v_1515 & v_1516 & ~v_1517 & ~v_1518;
assign v_5288 = v_5284 & v_1515 & v_1516 & v_1517;
assign v_5289 = v_5284 & v_1515 & ~v_1516 & ~v_1520;
assign v_5291 = v_5290 & v_2113;
assign v_5292 = v_5273 & v_1469 & v_1470 & v_1485 & v_1486;
assign v_5293 = v_5265 & v_1446 & v_1447 & v_1462 & v_1463;
assign v_5296 = v_5295 & v_227;
assign v_5297 = v_5295 & ~v_227 & v_229 & v_262 & ~v_264;
assign v_5298 = v_5295 & ~v_227 & v_229 & v_262 & v_264;
assign v_5299 = v_5295 & ~v_227 & v_229 & ~v_262;
assign v_5300 = v_5295 & v_230;
assign v_5301 = v_5295 & ~v_230;
assign v_5304 = v_5302 & v_5303;
assign v_5305 = v_5302 & v_1540;
assign v_5306 = v_13081 & v_13082;
assign v_5308 = v_5307 & ~v_227 & ~v_229 & v_260;
assign v_5310 = v_5309 & v_267 & v_268;
assign v_5311 = v_5309 & v_267 & ~v_268;
assign v_5313 = v_5312 & ~v_279;
assign v_5315 = v_5312 & v_5314;
assign v_5316 = v_5312 & v_279 & v_291 & ~v_292 & v_300;
assign v_5319 = v_5317 & v_5318;
assign v_5320 = v_5317 & v_321 & v_322;
assign v_5321 = v_5317 & v_321 & ~v_322 & v_324;
assign v_5322 = v_5317 & v_321 & ~v_322 & ~v_324 & v_326;
assign v_5323 = v_5317 & v_321 & ~v_322 & ~v_324 & ~v_326;
assign v_5325 = v_5324 & v_1563;
assign v_5327 = v_5326 & ~v_308 & v_309 & v_329;
assign v_5330 = v_5328 & v_5329;
assign v_5331 = v_5328 & v_1570;
assign v_5333 = v_5332 & v_345 & v_346;
assign v_5334 = v_5332 & v_345 & ~v_346 & v_348;
assign v_5335 = v_5332 & v_345 & ~v_346 & ~v_348 & v_350;
assign v_5336 = v_5332 & v_356 & v_357;
assign v_5337 = v_5332 & v_359 & v_360;
assign v_5338 = v_5332 & v_359 & ~v_360 & v_362;
assign v_5339 = v_5332 & v_359 & ~v_360 & ~v_362 & v_364;
assign v_5340 = v_5332 & v_1582;
assign v_5342 = v_5341 & v_1585;
assign v_5344 = v_5343 & v_356 & ~v_357 & v_369 & v_370;
assign v_5345 = v_5343 & v_372 & v_373;
assign v_5346 = v_5343 & v_372 & ~v_373 & v_375;
assign v_5347 = v_5343 & v_372 & ~v_373 & ~v_375 & v_377;
assign v_5349 = v_5343 & v_5348;
assign v_5350 = v_13083 & v_13084;
assign v_5352 = v_5351 & v_384 & v_385;
assign v_5353 = v_5351 & v_384 & ~v_385;
assign v_5355 = v_5354 & v_1599;
assign v_5357 = v_13085 & v_13086;
assign v_5358 = v_5356 & v_391 & v_392;
assign v_5359 = v_5356 & v_391 & ~v_392 & v_394;
assign v_5360 = v_5356 & v_391 & ~v_392 & ~v_394 & v_396;
assign v_5361 = v_5356 & v_1606;
assign v_5363 = v_13087 & v_13088;
assign v_5365 = v_5364 & v_1611;
assign v_5367 = v_5366 & v_410 & v_411;
assign v_5368 = v_5366 & v_410 & ~v_411 & v_413;
assign v_5369 = v_5366 & v_410 & ~v_411 & ~v_413 & v_415;
assign v_5370 = v_5366 & v_421 & v_422;
assign v_5371 = v_5366 & v_424 & v_425;
assign v_5372 = v_5366 & v_424 & ~v_425 & v_427;
assign v_5373 = v_5366 & v_424 & ~v_425 & ~v_427 & v_429;
assign v_5374 = v_5366 & v_1621;
assign v_5376 = v_5375 & v_1624;
assign v_5378 = v_5377 & v_421 & ~v_422 & v_434 & v_435;
assign v_5379 = v_5377 & v_437 & v_438;
assign v_5380 = v_5377 & v_437 & ~v_438 & v_440;
assign v_5381 = v_5377 & v_437 & ~v_438 & ~v_440 & v_442;
assign v_5383 = v_5377 & v_5382;
assign v_5384 = v_13089 & v_13090;
assign v_5386 = v_5385 & v_449 & v_450;
assign v_5387 = v_5385 & v_449 & ~v_450;
assign v_5389 = v_5388 & v_1638;
assign v_5391 = v_13091 & v_13092;
assign v_5392 = v_5390 & v_456 & v_457;
assign v_5393 = v_5390 & v_456 & ~v_457 & v_459;
assign v_5394 = v_5390 & v_456 & ~v_457 & ~v_459 & v_461;
assign v_5395 = v_5390 & v_1645;
assign v_5397 = v_13093 & v_13094;
assign v_5399 = v_5398 & v_1650;
assign v_5401 = v_5400 & v_491;
assign v_5402 = v_5400 & ~v_491 & v_493 & v_526 & ~v_528;
assign v_5403 = v_5400 & ~v_491 & v_493 & v_526 & v_528;
assign v_5404 = v_5400 & ~v_491 & v_493 & ~v_526;
assign v_5405 = v_5400 & v_494;
assign v_5406 = v_5400 & ~v_494;
assign v_5409 = v_5407 & v_5408;
assign v_5410 = v_5407 & v_1666;
assign v_5411 = v_13095 & v_13096;
assign v_5413 = v_5412 & ~v_491 & ~v_493 & v_524;
assign v_5415 = v_5414 & v_531 & v_532;
assign v_5416 = v_5414 & v_531 & ~v_532;
assign v_5418 = v_5417 & v_546 & v_547;
assign v_5419 = v_5417 & v_546 & ~v_547 & ~v_551;
assign v_5421 = v_5420 & v_546 & ~v_547 & v_551;
assign v_5423 = v_5422 & v_554;
assign v_5425 = v_5424 & v_558 & v_559;
assign v_5426 = v_5424 & v_558 & ~v_559 & v_561;
assign v_5427 = v_5424 & v_1682;
assign v_5430 = v_5428 & v_5429;
assign v_5431 = v_5428 & v_1687;
assign v_5433 = v_5432 & v_588 & ~v_589 & ~v_591;
assign v_5434 = v_5432 & v_593 & ~v_594;
assign v_5435 = v_5432 & v_593 & v_594;
assign v_5436 = v_5432 & v_583;
assign v_5438 = v_5437 & v_604 & v_605;
assign v_5439 = v_5437 & v_604 & ~v_605 & ~v_609;
assign v_5441 = v_5440 & v_604 & ~v_605 & v_609;
assign v_5443 = v_5442 & v_612;
assign v_5445 = v_5444 & v_616 & v_617;
assign v_5446 = v_5444 & v_616 & ~v_617 & v_619;
assign v_5447 = v_5444 & v_1700;
assign v_5450 = v_5448 & v_5449;
assign v_5451 = v_5448 & v_1705;
assign v_5453 = v_2 & v_5452;
assign v_5454 = v_641 & v_5432;
assign v_5455 = v_643 & v_5417;
assign v_5456 = v_645 & v_5417;
assign v_5457 = v_647 & v_5417;
assign v_5458 = v_649 & v_5417;
assign v_5459 = ~v_649 & v_5400;
assign v_5461 = ~v_647 & v_5460;
assign v_5463 = ~v_645 & v_5462;
assign v_5465 = ~v_643 & v_5464;
assign v_5467 = ~v_641 & v_5466;
assign v_5469 = ~v_2 & v_5468;
assign v_5471 = v_5470 & ~v_669;
assign v_5472 = v_13097 & v_13098;
assign v_5473 = v_5470 & v_669 & v_670 & v_672 & v_674;
assign v_5474 = v_13099 & v_13100;
assign v_5476 = v_5475 & v_679 & ~v_680 & v_682;
assign v_5477 = v_5475 & v_689 & ~v_690 & ~v_692;
assign v_5478 = v_5475 & v_694 & ~v_695;
assign v_5479 = v_5475 & v_694 & v_695;
assign v_5480 = v_5475 & v_684;
assign v_5482 = v_5481 & v_1737;
assign v_5484 = v_5483 & v_1740;
assign v_5485 = v_5475 & v_679 & v_680;
assign v_5486 = v_5470 & v_1743;
assign v_5488 = v_5487 & ~v_705;
assign v_5489 = v_5487 & v_710 & v_711;
assign v_5490 = v_5487 & v_710 & ~v_711 & ~v_715;
assign v_5492 = v_5491 & v_710 & ~v_711 & v_715;
assign v_5494 = v_5493 & v_718;
assign v_5496 = v_5495 & v_705 & v_722 & v_723 & ~v_724;
assign v_5498 = v_5495 & v_5497;
assign v_5499 = v_5495 & v_750 & v_751;
assign v_5500 = v_5495 & v_750 & ~v_751;
assign v_5502 = v_5501 & v_763 & v_764;
assign v_5503 = v_5501 & v_763 & ~v_764;
assign v_5505 = v_5504 & v_745 & v_758 & v_771;
assign v_5506 = v_13101 & v_13102;
assign v_5507 = v_5495 & v_779 & v_780;
assign v_5508 = v_5495 & v_779 & ~v_780 & ~v_784;
assign v_5510 = v_5509 & v_779 & ~v_780 & v_784;
assign v_5512 = v_5511 & v_787;
assign v_5514 = v_5513 & v_1764;
assign v_5516 = v_5515 & v_798 & ~v_799 & v_817;
assign v_5517 = v_5515 & v_798 & ~v_799 & ~v_817;
assign v_5518 = v_5515 & ~v_800;
assign v_5519 = v_5515 & v_808 & ~v_809;
assign v_5520 = v_5515 & v_1771;
assign v_5522 = v_5521 & v_798 & v_799 & v_814 & ~v_815;
assign v_5524 = v_5523 & v_821 & ~v_822 & v_840;
assign v_5525 = v_5523 & v_821 & ~v_822 & ~v_840;
assign v_5526 = v_5523 & ~v_823;
assign v_5527 = v_5523 & v_831 & ~v_832;
assign v_5528 = v_5523 & v_1780;
assign v_5530 = v_5529 & v_821 & v_822 & v_837 & ~v_838;
assign v_5532 = v_5531 & v_844 & ~v_845 & v_863;
assign v_5533 = v_5531 & ~v_846;
assign v_5534 = v_5531 & v_854 & ~v_855;
assign v_5535 = v_5531 & v_1788;
assign v_5537 = v_5536 & v_844 & v_845 & v_860 & v_861;
assign v_5538 = v_5531 & v_844 & ~v_845 & ~v_863;
assign v_5539 = v_5536 & v_844 & v_845 & v_860 & ~v_861;
assign v_5542 = v_5540 & v_5541;
assign v_5543 = v_5540 & v_867 & v_868 & ~v_869 & ~v_870;
assign v_5544 = v_5540 & v_867 & v_868 & v_869;
assign v_5545 = v_5540 & v_867 & ~v_868 & ~v_872;
assign v_5547 = v_5546 & v_1801;
assign v_5548 = v_5529 & v_821 & v_822 & v_837 & v_838;
assign v_5549 = v_5521 & v_798 & v_799 & v_814 & v_815;
assign v_5551 = v_5550 & v_879 & ~v_880 & v_898;
assign v_5552 = v_5550 & v_879 & ~v_880 & ~v_898;
assign v_5553 = v_5550 & ~v_881;
assign v_5554 = v_5550 & v_889 & ~v_890;
assign v_5555 = v_5550 & v_1810;
assign v_5557 = v_5556 & v_879 & v_880 & v_895 & ~v_896;
assign v_5559 = v_5558 & v_902 & ~v_903 & v_921;
assign v_5560 = v_5558 & v_902 & ~v_903 & ~v_921;
assign v_5561 = v_5558 & ~v_904;
assign v_5562 = v_5558 & v_912 & ~v_913;
assign v_5563 = v_5558 & v_1819;
assign v_5565 = v_5564 & v_902 & v_903 & v_918 & ~v_919;
assign v_5567 = v_5566 & v_925 & ~v_926 & v_944;
assign v_5568 = v_5566 & ~v_927;
assign v_5569 = v_5566 & v_935 & ~v_936;
assign v_5570 = v_5566 & v_1827;
assign v_5572 = v_5571 & v_925 & v_926 & v_941 & v_942;
assign v_5573 = v_5566 & v_925 & ~v_926 & ~v_944;
assign v_5574 = v_5571 & v_925 & v_926 & v_941 & ~v_942;
assign v_5577 = v_5575 & v_5576;
assign v_5578 = v_5575 & v_948 & v_949 & ~v_950 & ~v_951;
assign v_5579 = v_5575 & v_948 & v_949 & v_950;
assign v_5580 = v_5575 & v_948 & ~v_949 & ~v_953;
assign v_5582 = v_5581 & v_1840;
assign v_5583 = v_5564 & v_902 & v_903 & v_918 & v_919;
assign v_5584 = v_5556 & v_879 & v_880 & v_895 & v_896;
assign v_5586 = v_5585 & v_960 & ~v_961 & v_979;
assign v_5587 = v_5585 & v_960 & ~v_961 & ~v_979;
assign v_5588 = v_5585 & ~v_962;
assign v_5589 = v_5585 & v_970 & ~v_971;
assign v_5590 = v_5585 & v_1849;
assign v_5592 = v_5591 & v_960 & v_961 & v_976 & ~v_977;
assign v_5594 = v_5593 & v_983 & ~v_984 & v_1002;
assign v_5595 = v_5593 & v_983 & ~v_984 & ~v_1002;
assign v_5596 = v_5593 & ~v_985;
assign v_5597 = v_5593 & v_993 & ~v_994;
assign v_5598 = v_5593 & v_1858;
assign v_5600 = v_5599 & v_983 & v_984 & v_999 & ~v_1000;
assign v_5602 = v_5601 & v_1006 & ~v_1007 & v_1025;
assign v_5603 = v_5601 & ~v_1008;
assign v_5604 = v_5601 & v_1016 & ~v_1017;
assign v_5605 = v_5601 & v_1866;
assign v_5607 = v_5606 & v_1006 & v_1007 & v_1022 & v_1023;
assign v_5608 = v_5601 & v_1006 & ~v_1007 & ~v_1025;
assign v_5609 = v_5606 & v_1006 & v_1007 & v_1022 & ~v_1023;
assign v_5612 = v_5610 & v_5611;
assign v_5613 = v_5610 & v_1029 & v_1030 & ~v_1031 & ~v_1032;
assign v_5614 = v_5610 & v_1029 & v_1030 & v_1031;
assign v_5615 = v_5610 & v_1029 & ~v_1030 & ~v_1034;
assign v_5617 = v_5616 & v_1879;
assign v_5618 = v_5599 & v_983 & v_984 & v_999 & v_1000;
assign v_5619 = v_5591 & v_960 & v_961 & v_976 & v_977;
assign v_5621 = v_5620 & v_1041 & ~v_1042 & v_1060;
assign v_5622 = v_5620 & v_1041 & ~v_1042 & ~v_1060;
assign v_5623 = v_5620 & ~v_1043;
assign v_5624 = v_5620 & v_1051 & ~v_1052;
assign v_5625 = v_5620 & v_1888;
assign v_5627 = v_5626 & v_1041 & v_1042 & v_1057 & ~v_1058;
assign v_5629 = v_5628 & v_1064 & ~v_1065 & v_1083;
assign v_5630 = v_5628 & v_1064 & ~v_1065 & ~v_1083;
assign v_5631 = v_5628 & ~v_1066;
assign v_5632 = v_5628 & v_1074 & ~v_1075;
assign v_5633 = v_5628 & v_1897;
assign v_5635 = v_5634 & v_1064 & v_1065 & v_1080 & ~v_1081;
assign v_5637 = v_5636 & v_1087 & ~v_1088 & v_1106;
assign v_5638 = v_5636 & ~v_1089;
assign v_5639 = v_5636 & v_1097 & ~v_1098;
assign v_5640 = v_5636 & v_1905;
assign v_5642 = v_5641 & v_1087 & v_1088 & v_1103 & v_1104;
assign v_5643 = v_5636 & v_1087 & ~v_1088 & ~v_1106;
assign v_5644 = v_5641 & v_1087 & v_1088 & v_1103 & ~v_1104;
assign v_5647 = v_5645 & v_5646;
assign v_5648 = v_5645 & v_1110 & v_1111 & ~v_1112 & ~v_1113;
assign v_5649 = v_5645 & v_1110 & v_1111 & v_1112;
assign v_5650 = v_5645 & v_1110 & ~v_1111 & ~v_1115;
assign v_5652 = v_5651 & v_1918;
assign v_5653 = v_5634 & v_1064 & v_1065 & v_1080 & v_1081;
assign v_5654 = v_5626 & v_1041 & v_1042 & v_1057 & v_1058;
assign v_5656 = v_5655 & v_1122 & ~v_1123 & v_1141;
assign v_5657 = v_5655 & v_1122 & ~v_1123 & ~v_1141;
assign v_5658 = v_5655 & ~v_1124;
assign v_5659 = v_5655 & v_1132 & ~v_1133;
assign v_5660 = v_5655 & v_1927;
assign v_5662 = v_5661 & v_1122 & v_1123 & v_1138 & ~v_1139;
assign v_5664 = v_5663 & v_1145 & ~v_1146 & v_1164;
assign v_5665 = v_5663 & v_1145 & ~v_1146 & ~v_1164;
assign v_5666 = v_5663 & ~v_1147;
assign v_5667 = v_5663 & v_1155 & ~v_1156;
assign v_5668 = v_5663 & v_1936;
assign v_5670 = v_5669 & v_1145 & v_1146 & v_1161 & ~v_1162;
assign v_5672 = v_5671 & v_1168 & ~v_1169 & v_1187;
assign v_5673 = v_5671 & ~v_1170;
assign v_5674 = v_5671 & v_1178 & ~v_1179;
assign v_5675 = v_5671 & v_1944;
assign v_5677 = v_5676 & v_1168 & v_1169 & v_1184 & v_1185;
assign v_5678 = v_5671 & v_1168 & ~v_1169 & ~v_1187;
assign v_5679 = v_5676 & v_1168 & v_1169 & v_1184 & ~v_1185;
assign v_5682 = v_5680 & v_5681;
assign v_5683 = v_5680 & v_1191 & v_1192 & ~v_1193 & ~v_1194;
assign v_5684 = v_5680 & v_1191 & v_1192 & v_1193;
assign v_5685 = v_5680 & v_1191 & ~v_1192 & ~v_1196;
assign v_5687 = v_5686 & v_1957;
assign v_5688 = v_5669 & v_1145 & v_1146 & v_1161 & v_1162;
assign v_5689 = v_5661 & v_1122 & v_1123 & v_1138 & v_1139;
assign v_5691 = v_5690 & v_1203 & ~v_1204 & v_1222;
assign v_5692 = v_5690 & v_1203 & ~v_1204 & ~v_1222;
assign v_5693 = v_5690 & ~v_1205;
assign v_5694 = v_5690 & v_1213 & ~v_1214;
assign v_5695 = v_5690 & v_1966;
assign v_5697 = v_5696 & v_1203 & v_1204 & v_1219 & ~v_1220;
assign v_5699 = v_5698 & v_1226 & ~v_1227 & v_1245;
assign v_5700 = v_5698 & v_1226 & ~v_1227 & ~v_1245;
assign v_5701 = v_5698 & ~v_1228;
assign v_5702 = v_5698 & v_1236 & ~v_1237;
assign v_5703 = v_5698 & v_1975;
assign v_5705 = v_5704 & v_1226 & v_1227 & v_1242 & ~v_1243;
assign v_5707 = v_5706 & v_1249 & ~v_1250 & v_1268;
assign v_5708 = v_5706 & ~v_1251;
assign v_5709 = v_5706 & v_1259 & ~v_1260;
assign v_5710 = v_5706 & v_1983;
assign v_5712 = v_5711 & v_1249 & v_1250 & v_1265 & v_1266;
assign v_5713 = v_5706 & v_1249 & ~v_1250 & ~v_1268;
assign v_5714 = v_5711 & v_1249 & v_1250 & v_1265 & ~v_1266;
assign v_5717 = v_5715 & v_5716;
assign v_5718 = v_5715 & v_1272 & v_1273 & ~v_1274 & ~v_1275;
assign v_5719 = v_5715 & v_1272 & v_1273 & v_1274;
assign v_5720 = v_5715 & v_1272 & ~v_1273 & ~v_1277;
assign v_5722 = v_5721 & v_1996;
assign v_5723 = v_5704 & v_1226 & v_1227 & v_1242 & v_1243;
assign v_5724 = v_5696 & v_1203 & v_1204 & v_1219 & v_1220;
assign v_5726 = v_5725 & v_1284 & ~v_1285 & v_1303;
assign v_5727 = v_5725 & v_1284 & ~v_1285 & ~v_1303;
assign v_5728 = v_5725 & ~v_1286;
assign v_5729 = v_5725 & v_1294 & ~v_1295;
assign v_5730 = v_5725 & v_2005;
assign v_5732 = v_5731 & v_1284 & v_1285 & v_1300 & ~v_1301;
assign v_5734 = v_5733 & v_1307 & ~v_1308 & v_1326;
assign v_5735 = v_5733 & v_1307 & ~v_1308 & ~v_1326;
assign v_5736 = v_5733 & ~v_1309;
assign v_5737 = v_5733 & v_1317 & ~v_1318;
assign v_5738 = v_5733 & v_2014;
assign v_5740 = v_5739 & v_1307 & v_1308 & v_1323 & ~v_1324;
assign v_5742 = v_5741 & v_1330 & ~v_1331 & v_1349;
assign v_5743 = v_5741 & ~v_1332;
assign v_5744 = v_5741 & v_1340 & ~v_1341;
assign v_5745 = v_5741 & v_2022;
assign v_5747 = v_5746 & v_1330 & v_1331 & v_1346 & v_1347;
assign v_5748 = v_5741 & v_1330 & ~v_1331 & ~v_1349;
assign v_5749 = v_5746 & v_1330 & v_1331 & v_1346 & ~v_1347;
assign v_5752 = v_5750 & v_5751;
assign v_5753 = v_5750 & v_1353 & v_1354 & ~v_1355 & ~v_1356;
assign v_5754 = v_5750 & v_1353 & v_1354 & v_1355;
assign v_5755 = v_5750 & v_1353 & ~v_1354 & ~v_1358;
assign v_5757 = v_5756 & v_2035;
assign v_5758 = v_5739 & v_1307 & v_1308 & v_1323 & v_1324;
assign v_5759 = v_5731 & v_1284 & v_1285 & v_1300 & v_1301;
assign v_5761 = v_5760 & v_1365 & ~v_1366 & v_1384;
assign v_5762 = v_5760 & v_1365 & ~v_1366 & ~v_1384;
assign v_5763 = v_5760 & ~v_1367;
assign v_5764 = v_5760 & v_1375 & ~v_1376;
assign v_5765 = v_5760 & v_2044;
assign v_5767 = v_5766 & v_1365 & v_1366 & v_1381 & ~v_1382;
assign v_5769 = v_5768 & v_1388 & ~v_1389 & v_1407;
assign v_5770 = v_5768 & v_1388 & ~v_1389 & ~v_1407;
assign v_5771 = v_5768 & ~v_1390;
assign v_5772 = v_5768 & v_1398 & ~v_1399;
assign v_5773 = v_5768 & v_2053;
assign v_5775 = v_5774 & v_1388 & v_1389 & v_1404 & ~v_1405;
assign v_5777 = v_5776 & v_1411 & ~v_1412 & v_1430;
assign v_5778 = v_5776 & ~v_1413;
assign v_5779 = v_5776 & v_1421 & ~v_1422;
assign v_5780 = v_5776 & v_2061;
assign v_5782 = v_5781 & v_1411 & v_1412 & v_1427 & v_1428;
assign v_5783 = v_5776 & v_1411 & ~v_1412 & ~v_1430;
assign v_5784 = v_5781 & v_1411 & v_1412 & v_1427 & ~v_1428;
assign v_5787 = v_5785 & v_5786;
assign v_5788 = v_5785 & v_1434 & v_1435 & ~v_1436 & ~v_1437;
assign v_5789 = v_5785 & v_1434 & v_1435 & v_1436;
assign v_5790 = v_5785 & v_1434 & ~v_1435 & ~v_1439;
assign v_5792 = v_5791 & v_2074;
assign v_5793 = v_5774 & v_1388 & v_1389 & v_1404 & v_1405;
assign v_5794 = v_5766 & v_1365 & v_1366 & v_1381 & v_1382;
assign v_5796 = v_5795 & v_1446 & ~v_1447 & v_1465;
assign v_5797 = v_5795 & v_1446 & ~v_1447 & ~v_1465;
assign v_5798 = v_5795 & ~v_1448;
assign v_5799 = v_5795 & v_1456 & ~v_1457;
assign v_5800 = v_5795 & v_2083;
assign v_5802 = v_5801 & v_1446 & v_1447 & v_1462 & ~v_1463;
assign v_5804 = v_5803 & v_1469 & ~v_1470 & v_1488;
assign v_5805 = v_5803 & v_1469 & ~v_1470 & ~v_1488;
assign v_5806 = v_5803 & ~v_1471;
assign v_5807 = v_5803 & v_1479 & ~v_1480;
assign v_5808 = v_5803 & v_2092;
assign v_5810 = v_5809 & v_1469 & v_1470 & v_1485 & ~v_1486;
assign v_5812 = v_5811 & v_1492 & ~v_1493 & v_1511;
assign v_5813 = v_5811 & ~v_1494;
assign v_5814 = v_5811 & v_1502 & ~v_1503;
assign v_5815 = v_5811 & v_2100;
assign v_5817 = v_5816 & v_1492 & v_1493 & v_1508 & v_1509;
assign v_5818 = v_5811 & v_1492 & ~v_1493 & ~v_1511;
assign v_5819 = v_5816 & v_1492 & v_1493 & v_1508 & ~v_1509;
assign v_5822 = v_5820 & v_5821;
assign v_5823 = v_5820 & v_1515 & v_1516 & ~v_1517 & ~v_1518;
assign v_5824 = v_5820 & v_1515 & v_1516 & v_1517;
assign v_5825 = v_5820 & v_1515 & ~v_1516 & ~v_1520;
assign v_5827 = v_5826 & v_2113;
assign v_5828 = v_5809 & v_1469 & v_1470 & v_1485 & v_1486;
assign v_5829 = v_5801 & v_1446 & v_1447 & v_1462 & v_1463;
assign v_5832 = v_5831 & ~v_1572;
assign v_5834 = v_1527 & v_5833;
assign v_5835 = v_227;
assign v_5837 = v_5836 & v_267 & v_268;
assign v_5838 = v_5836 & v_267 & ~v_268;
assign v_5840 = v_5839 & ~v_279;
assign v_5842 = v_5839 & v_5841;
assign v_5843 = v_5839 & v_279 & v_291 & ~v_292 & v_300;
assign v_5846 = v_5844 & v_5845;
assign v_5847 = v_5844 & v_321 & v_322;
assign v_5848 = v_5844 & v_321 & ~v_322 & v_324;
assign v_5849 = v_5844 & v_321 & ~v_322 & ~v_324 & v_326;
assign v_5850 = v_5844 & v_321 & ~v_322 & ~v_324 & ~v_326;
assign v_5852 = v_5851 & v_1563;
assign v_5854 = v_5853 & ~v_308 & v_309 & v_329;
assign v_5857 = v_5855 & v_5856;
assign v_5858 = v_5855 & v_1570;
assign v_5860 = ~v_1527 & v_5859;
assign v_5862 = v_5861 & v_345 & v_346;
assign v_5863 = v_5861 & v_345 & ~v_346 & v_348;
assign v_5864 = v_5861 & v_345 & ~v_346 & ~v_348 & v_350;
assign v_5865 = v_5861 & v_356 & v_357;
assign v_5866 = v_5861 & v_359 & v_360;
assign v_5867 = v_5861 & v_359 & ~v_360 & v_362;
assign v_5868 = v_5861 & v_359 & ~v_360 & ~v_362 & v_364;
assign v_5869 = v_5861 & v_1582;
assign v_5871 = v_5870 & v_1585;
assign v_5873 = v_5872 & v_356 & ~v_357 & v_369 & v_370;
assign v_5874 = v_5872 & v_372 & v_373;
assign v_5875 = v_5872 & v_372 & ~v_373 & v_375;
assign v_5876 = v_5872 & v_372 & ~v_373 & ~v_375 & v_377;
assign v_5878 = v_5872 & v_5877;
assign v_5879 = v_13103 & v_13104;
assign v_5881 = v_5880 & v_384 & v_385;
assign v_5882 = v_5880 & v_384 & ~v_385;
assign v_5884 = v_5883 & v_1599;
assign v_5886 = v_13105 & v_13106;
assign v_5887 = v_5885 & v_391 & v_392;
assign v_5888 = v_5885 & v_391 & ~v_392 & v_394;
assign v_5889 = v_5885 & v_391 & ~v_392 & ~v_394 & v_396;
assign v_5890 = v_5885 & v_1606;
assign v_5892 = v_13107 & v_13108;
assign v_5894 = v_5893 & v_1611;
assign v_5896 = v_5895 & v_410 & v_411;
assign v_5897 = v_5895 & v_410 & ~v_411 & v_413;
assign v_5898 = v_5895 & v_410 & ~v_411 & ~v_413 & v_415;
assign v_5899 = v_5895 & v_421 & v_422;
assign v_5900 = v_5895 & v_424 & v_425;
assign v_5901 = v_5895 & v_424 & ~v_425 & v_427;
assign v_5902 = v_5895 & v_424 & ~v_425 & ~v_427 & v_429;
assign v_5903 = v_5895 & v_1621;
assign v_5905 = v_5904 & v_1624;
assign v_5907 = v_5906 & v_421 & ~v_422 & v_434 & v_435;
assign v_5908 = v_5906 & v_437 & v_438;
assign v_5909 = v_5906 & v_437 & ~v_438 & v_440;
assign v_5910 = v_5906 & v_437 & ~v_438 & ~v_440 & v_442;
assign v_5912 = v_5906 & v_5911;
assign v_5913 = v_13109 & v_13110;
assign v_5915 = v_5914 & v_449 & v_450;
assign v_5916 = v_5914 & v_449 & ~v_450;
assign v_5918 = v_5917 & v_1638;
assign v_5920 = v_13111 & v_13112;
assign v_5921 = v_5919 & v_456 & v_457;
assign v_5922 = v_5919 & v_456 & ~v_457 & v_459;
assign v_5923 = v_5919 & v_456 & ~v_457 & ~v_459 & v_461;
assign v_5924 = v_5919 & v_1645;
assign v_5926 = v_13113 & v_13114;
assign v_5928 = v_5927 & v_1650;
assign v_5930 = v_5929 & v_491;
assign v_5932 = v_5931 & v_531 & v_532;
assign v_5933 = v_5931 & v_531 & ~v_532;
assign v_5935 = v_5934 & v_546 & v_547;
assign v_5936 = v_5934 & v_554;
assign v_5938 = v_5937 & v_558 & v_559;
assign v_5939 = v_5937 & v_558 & ~v_559 & v_561;
assign v_5940 = v_5937 & v_1682;
assign v_5943 = v_5941 & v_5942;
assign v_5944 = v_5941 & v_1687;
assign v_5946 = v_5945 & v_588 & ~v_589 & ~v_591;
assign v_5947 = v_5945 & v_593 & ~v_594;
assign v_5948 = v_5945 & v_593 & v_594;
assign v_5949 = v_5945 & v_583;
assign v_5951 = v_5950 & v_604 & v_605;
assign v_5952 = v_5950 & v_612;
assign v_5954 = v_5953 & v_616 & v_617;
assign v_5955 = v_5953 & v_616 & ~v_617 & v_619;
assign v_5956 = v_5953 & v_1700;
assign v_5959 = v_5957 & v_5958;
assign v_5960 = v_5957 & v_1705;
assign v_5962 = v_2 & v_5961;
assign v_5963 = v_641 & v_5945;
assign v_5964 = v_643 & v_5934;
assign v_5965 = v_645 & v_5934;
assign v_5966 = v_647 & v_5934;
assign v_5967 = v_649 & v_5934;
assign v_5968 = ~v_649 & v_5929;
assign v_5970 = ~v_647 & v_5969;
assign v_5972 = ~v_645 & v_5971;
assign v_5974 = ~v_643 & v_5973;
assign v_5976 = ~v_641 & v_5975;
assign v_5978 = ~v_2 & v_5977;
assign v_5980 = v_5979 & ~v_669;
assign v_5981 = v_13115 & v_13116;
assign v_5982 = v_5979 & v_669 & v_670 & v_672 & v_674;
assign v_5983 = v_13117 & v_13118;
assign v_5985 = v_5984 & v_679 & ~v_680 & v_682;
assign v_5986 = v_5984 & v_689 & ~v_690 & ~v_692;
assign v_5987 = v_5984 & v_694 & ~v_695;
assign v_5988 = v_5984 & v_694 & v_695;
assign v_5989 = v_5984 & v_684;
assign v_5991 = v_5990 & v_1737;
assign v_5993 = v_5992 & v_1740;
assign v_5994 = v_5984 & v_679 & v_680;
assign v_5995 = v_5979 & v_1743;
assign v_5997 = v_5996 & ~v_705;
assign v_5998 = v_5996 & v_710 & v_711;
assign v_5999 = v_5996 & v_718;
assign v_6001 = v_6000 & v_705 & v_722 & v_723 & ~v_724;
assign v_6003 = v_6000 & v_6002;
assign v_6004 = v_6000 & v_750 & v_751;
assign v_6005 = v_6000 & v_750 & ~v_751;
assign v_6007 = v_6006 & v_763 & v_764;
assign v_6008 = v_6006 & v_763 & ~v_764;
assign v_6010 = v_6009 & v_745 & v_758 & v_771;
assign v_6011 = v_13119 & v_13120;
assign v_6012 = v_6000 & v_779 & v_780;
assign v_6013 = v_6000 & v_787;
assign v_6015 = v_6014 & v_1764;
assign v_6017 = v_6016 & v_798 & ~v_799 & v_817;
assign v_6018 = v_6016 & v_798 & ~v_799 & ~v_817;
assign v_6019 = v_6016 & ~v_800;
assign v_6020 = v_6016 & v_808 & ~v_809;
assign v_6021 = v_6016 & v_1771;
assign v_6023 = v_6022 & v_798 & v_799 & v_814 & ~v_815;
assign v_6025 = v_6024 & v_821 & ~v_822 & v_840;
assign v_6026 = v_6024 & v_821 & ~v_822 & ~v_840;
assign v_6027 = v_6024 & ~v_823;
assign v_6028 = v_6024 & v_831 & ~v_832;
assign v_6029 = v_6024 & v_1780;
assign v_6031 = v_6030 & v_821 & v_822 & v_837 & ~v_838;
assign v_6033 = v_6032 & v_844 & ~v_845 & v_863;
assign v_6034 = v_6032 & ~v_846;
assign v_6035 = v_6032 & v_854 & ~v_855;
assign v_6036 = v_6032 & v_1788;
assign v_6038 = v_6037 & v_844 & v_845 & v_860 & v_861;
assign v_6039 = v_6032 & v_844 & ~v_845 & ~v_863;
assign v_6040 = v_6037 & v_844 & v_845 & v_860 & ~v_861;
assign v_6043 = v_6041 & v_6042;
assign v_6044 = v_6041 & v_867 & v_868 & ~v_869 & ~v_870;
assign v_6045 = v_6041 & v_867 & v_868 & v_869;
assign v_6046 = v_6041 & v_867 & ~v_868 & ~v_872;
assign v_6048 = v_6047 & v_1801;
assign v_6049 = v_6030 & v_821 & v_822 & v_837 & v_838;
assign v_6050 = v_6022 & v_798 & v_799 & v_814 & v_815;
assign v_6052 = v_6051 & v_879 & ~v_880 & v_898;
assign v_6053 = v_6051 & v_879 & ~v_880 & ~v_898;
assign v_6054 = v_6051 & ~v_881;
assign v_6055 = v_6051 & v_889 & ~v_890;
assign v_6056 = v_6051 & v_1810;
assign v_6058 = v_6057 & v_879 & v_880 & v_895 & ~v_896;
assign v_6060 = v_6059 & v_902 & ~v_903 & v_921;
assign v_6061 = v_6059 & v_902 & ~v_903 & ~v_921;
assign v_6062 = v_6059 & ~v_904;
assign v_6063 = v_6059 & v_912 & ~v_913;
assign v_6064 = v_6059 & v_1819;
assign v_6066 = v_6065 & v_902 & v_903 & v_918 & ~v_919;
assign v_6068 = v_6067 & v_925 & ~v_926 & v_944;
assign v_6069 = v_6067 & ~v_927;
assign v_6070 = v_6067 & v_935 & ~v_936;
assign v_6071 = v_6067 & v_1827;
assign v_6073 = v_6072 & v_925 & v_926 & v_941 & v_942;
assign v_6074 = v_6067 & v_925 & ~v_926 & ~v_944;
assign v_6075 = v_6072 & v_925 & v_926 & v_941 & ~v_942;
assign v_6078 = v_6076 & v_6077;
assign v_6079 = v_6076 & v_948 & v_949 & ~v_950 & ~v_951;
assign v_6080 = v_6076 & v_948 & v_949 & v_950;
assign v_6081 = v_6076 & v_948 & ~v_949 & ~v_953;
assign v_6083 = v_6082 & v_1840;
assign v_6084 = v_6065 & v_902 & v_903 & v_918 & v_919;
assign v_6085 = v_6057 & v_879 & v_880 & v_895 & v_896;
assign v_6087 = v_6086 & v_960 & ~v_961 & v_979;
assign v_6088 = v_6086 & v_960 & ~v_961 & ~v_979;
assign v_6089 = v_6086 & ~v_962;
assign v_6090 = v_6086 & v_970 & ~v_971;
assign v_6091 = v_6086 & v_1849;
assign v_6093 = v_6092 & v_960 & v_961 & v_976 & ~v_977;
assign v_6095 = v_6094 & v_983 & ~v_984 & v_1002;
assign v_6096 = v_6094 & v_983 & ~v_984 & ~v_1002;
assign v_6097 = v_6094 & ~v_985;
assign v_6098 = v_6094 & v_993 & ~v_994;
assign v_6099 = v_6094 & v_1858;
assign v_6101 = v_6100 & v_983 & v_984 & v_999 & ~v_1000;
assign v_6103 = v_6102 & v_1006 & ~v_1007 & v_1025;
assign v_6104 = v_6102 & ~v_1008;
assign v_6105 = v_6102 & v_1016 & ~v_1017;
assign v_6106 = v_6102 & v_1866;
assign v_6108 = v_6107 & v_1006 & v_1007 & v_1022 & v_1023;
assign v_6109 = v_6102 & v_1006 & ~v_1007 & ~v_1025;
assign v_6110 = v_6107 & v_1006 & v_1007 & v_1022 & ~v_1023;
assign v_6113 = v_6111 & v_6112;
assign v_6114 = v_6111 & v_1029 & v_1030 & ~v_1031 & ~v_1032;
assign v_6115 = v_6111 & v_1029 & v_1030 & v_1031;
assign v_6116 = v_6111 & v_1029 & ~v_1030 & ~v_1034;
assign v_6118 = v_6117 & v_1879;
assign v_6119 = v_6100 & v_983 & v_984 & v_999 & v_1000;
assign v_6120 = v_6092 & v_960 & v_961 & v_976 & v_977;
assign v_6122 = v_6121 & v_1041 & ~v_1042 & v_1060;
assign v_6123 = v_6121 & v_1041 & ~v_1042 & ~v_1060;
assign v_6124 = v_6121 & ~v_1043;
assign v_6125 = v_6121 & v_1051 & ~v_1052;
assign v_6126 = v_6121 & v_1888;
assign v_6128 = v_6127 & v_1041 & v_1042 & v_1057 & ~v_1058;
assign v_6130 = v_6129 & v_1064 & ~v_1065 & v_1083;
assign v_6131 = v_6129 & v_1064 & ~v_1065 & ~v_1083;
assign v_6132 = v_6129 & ~v_1066;
assign v_6133 = v_6129 & v_1074 & ~v_1075;
assign v_6134 = v_6129 & v_1897;
assign v_6136 = v_6135 & v_1064 & v_1065 & v_1080 & ~v_1081;
assign v_6138 = v_6137 & v_1087 & ~v_1088 & v_1106;
assign v_6139 = v_6137 & ~v_1089;
assign v_6140 = v_6137 & v_1097 & ~v_1098;
assign v_6141 = v_6137 & v_1905;
assign v_6143 = v_6142 & v_1087 & v_1088 & v_1103 & v_1104;
assign v_6144 = v_6137 & v_1087 & ~v_1088 & ~v_1106;
assign v_6145 = v_6142 & v_1087 & v_1088 & v_1103 & ~v_1104;
assign v_6148 = v_6146 & v_6147;
assign v_6149 = v_6146 & v_1110 & v_1111 & ~v_1112 & ~v_1113;
assign v_6150 = v_6146 & v_1110 & v_1111 & v_1112;
assign v_6151 = v_6146 & v_1110 & ~v_1111 & ~v_1115;
assign v_6153 = v_6152 & v_1918;
assign v_6154 = v_6135 & v_1064 & v_1065 & v_1080 & v_1081;
assign v_6155 = v_6127 & v_1041 & v_1042 & v_1057 & v_1058;
assign v_6157 = v_6156 & v_1122 & ~v_1123 & v_1141;
assign v_6158 = v_6156 & v_1122 & ~v_1123 & ~v_1141;
assign v_6159 = v_6156 & ~v_1124;
assign v_6160 = v_6156 & v_1132 & ~v_1133;
assign v_6161 = v_6156 & v_1927;
assign v_6163 = v_6162 & v_1122 & v_1123 & v_1138 & ~v_1139;
assign v_6165 = v_6164 & v_1145 & ~v_1146 & v_1164;
assign v_6166 = v_6164 & v_1145 & ~v_1146 & ~v_1164;
assign v_6167 = v_6164 & ~v_1147;
assign v_6168 = v_6164 & v_1155 & ~v_1156;
assign v_6169 = v_6164 & v_1936;
assign v_6171 = v_6170 & v_1145 & v_1146 & v_1161 & ~v_1162;
assign v_6173 = v_6172 & v_1168 & ~v_1169 & v_1187;
assign v_6174 = v_6172 & ~v_1170;
assign v_6175 = v_6172 & v_1178 & ~v_1179;
assign v_6176 = v_6172 & v_1944;
assign v_6178 = v_6177 & v_1168 & v_1169 & v_1184 & v_1185;
assign v_6179 = v_6172 & v_1168 & ~v_1169 & ~v_1187;
assign v_6180 = v_6177 & v_1168 & v_1169 & v_1184 & ~v_1185;
assign v_6183 = v_6181 & v_6182;
assign v_6184 = v_6181 & v_1191 & v_1192 & ~v_1193 & ~v_1194;
assign v_6185 = v_6181 & v_1191 & v_1192 & v_1193;
assign v_6186 = v_6181 & v_1191 & ~v_1192 & ~v_1196;
assign v_6188 = v_6187 & v_1957;
assign v_6189 = v_6170 & v_1145 & v_1146 & v_1161 & v_1162;
assign v_6190 = v_6162 & v_1122 & v_1123 & v_1138 & v_1139;
assign v_6192 = v_6191 & v_1203 & ~v_1204 & v_1222;
assign v_6193 = v_6191 & v_1203 & ~v_1204 & ~v_1222;
assign v_6194 = v_6191 & ~v_1205;
assign v_6195 = v_6191 & v_1213 & ~v_1214;
assign v_6196 = v_6191 & v_1966;
assign v_6198 = v_6197 & v_1203 & v_1204 & v_1219 & ~v_1220;
assign v_6200 = v_6199 & v_1226 & ~v_1227 & v_1245;
assign v_6201 = v_6199 & v_1226 & ~v_1227 & ~v_1245;
assign v_6202 = v_6199 & ~v_1228;
assign v_6203 = v_6199 & v_1236 & ~v_1237;
assign v_6204 = v_6199 & v_1975;
assign v_6206 = v_6205 & v_1226 & v_1227 & v_1242 & ~v_1243;
assign v_6208 = v_6207 & v_1249 & ~v_1250 & v_1268;
assign v_6209 = v_6207 & ~v_1251;
assign v_6210 = v_6207 & v_1259 & ~v_1260;
assign v_6211 = v_6207 & v_1983;
assign v_6213 = v_6212 & v_1249 & v_1250 & v_1265 & v_1266;
assign v_6214 = v_6207 & v_1249 & ~v_1250 & ~v_1268;
assign v_6215 = v_6212 & v_1249 & v_1250 & v_1265 & ~v_1266;
assign v_6218 = v_6216 & v_6217;
assign v_6219 = v_6216 & v_1272 & v_1273 & ~v_1274 & ~v_1275;
assign v_6220 = v_6216 & v_1272 & v_1273 & v_1274;
assign v_6221 = v_6216 & v_1272 & ~v_1273 & ~v_1277;
assign v_6223 = v_6222 & v_1996;
assign v_6224 = v_6205 & v_1226 & v_1227 & v_1242 & v_1243;
assign v_6225 = v_6197 & v_1203 & v_1204 & v_1219 & v_1220;
assign v_6227 = v_6226 & v_1284 & ~v_1285 & v_1303;
assign v_6228 = v_6226 & v_1284 & ~v_1285 & ~v_1303;
assign v_6229 = v_6226 & ~v_1286;
assign v_6230 = v_6226 & v_1294 & ~v_1295;
assign v_6231 = v_6226 & v_2005;
assign v_6233 = v_6232 & v_1284 & v_1285 & v_1300 & ~v_1301;
assign v_6235 = v_6234 & v_1307 & ~v_1308 & v_1326;
assign v_6236 = v_6234 & v_1307 & ~v_1308 & ~v_1326;
assign v_6237 = v_6234 & ~v_1309;
assign v_6238 = v_6234 & v_1317 & ~v_1318;
assign v_6239 = v_6234 & v_2014;
assign v_6241 = v_6240 & v_1307 & v_1308 & v_1323 & ~v_1324;
assign v_6243 = v_6242 & v_1330 & ~v_1331 & v_1349;
assign v_6244 = v_6242 & ~v_1332;
assign v_6245 = v_6242 & v_1340 & ~v_1341;
assign v_6246 = v_6242 & v_2022;
assign v_6248 = v_6247 & v_1330 & v_1331 & v_1346 & v_1347;
assign v_6249 = v_6242 & v_1330 & ~v_1331 & ~v_1349;
assign v_6250 = v_6247 & v_1330 & v_1331 & v_1346 & ~v_1347;
assign v_6253 = v_6251 & v_6252;
assign v_6254 = v_6251 & v_1353 & v_1354 & ~v_1355 & ~v_1356;
assign v_6255 = v_6251 & v_1353 & v_1354 & v_1355;
assign v_6256 = v_6251 & v_1353 & ~v_1354 & ~v_1358;
assign v_6258 = v_6257 & v_2035;
assign v_6259 = v_6240 & v_1307 & v_1308 & v_1323 & v_1324;
assign v_6260 = v_6232 & v_1284 & v_1285 & v_1300 & v_1301;
assign v_6262 = v_6261 & v_1365 & ~v_1366 & v_1384;
assign v_6263 = v_6261 & v_1365 & ~v_1366 & ~v_1384;
assign v_6264 = v_6261 & ~v_1367;
assign v_6265 = v_6261 & v_1375 & ~v_1376;
assign v_6266 = v_6261 & v_2044;
assign v_6268 = v_6267 & v_1365 & v_1366 & v_1381 & ~v_1382;
assign v_6270 = v_6269 & v_1388 & ~v_1389 & v_1407;
assign v_6271 = v_6269 & v_1388 & ~v_1389 & ~v_1407;
assign v_6272 = v_6269 & ~v_1390;
assign v_6273 = v_6269 & v_1398 & ~v_1399;
assign v_6274 = v_6269 & v_2053;
assign v_6276 = v_6275 & v_1388 & v_1389 & v_1404 & ~v_1405;
assign v_6278 = v_6277 & v_1411 & ~v_1412 & v_1430;
assign v_6279 = v_6277 & ~v_1413;
assign v_6280 = v_6277 & v_1421 & ~v_1422;
assign v_6281 = v_6277 & v_2061;
assign v_6283 = v_6282 & v_1411 & v_1412 & v_1427 & v_1428;
assign v_6284 = v_6277 & v_1411 & ~v_1412 & ~v_1430;
assign v_6285 = v_6282 & v_1411 & v_1412 & v_1427 & ~v_1428;
assign v_6288 = v_6286 & v_6287;
assign v_6289 = v_6286 & v_1434 & v_1435 & ~v_1436 & ~v_1437;
assign v_6290 = v_6286 & v_1434 & v_1435 & v_1436;
assign v_6291 = v_6286 & v_1434 & ~v_1435 & ~v_1439;
assign v_6293 = v_6292 & v_2074;
assign v_6294 = v_6275 & v_1388 & v_1389 & v_1404 & v_1405;
assign v_6295 = v_6267 & v_1365 & v_1366 & v_1381 & v_1382;
assign v_6297 = v_6296 & v_1446 & ~v_1447 & v_1465;
assign v_6298 = v_6296 & v_1446 & ~v_1447 & ~v_1465;
assign v_6299 = v_6296 & ~v_1448;
assign v_6300 = v_6296 & v_1456 & ~v_1457;
assign v_6301 = v_6296 & v_2083;
assign v_6303 = v_6302 & v_1446 & v_1447 & v_1462 & ~v_1463;
assign v_6305 = v_6304 & v_1469 & ~v_1470 & v_1488;
assign v_6306 = v_6304 & v_1469 & ~v_1470 & ~v_1488;
assign v_6307 = v_6304 & ~v_1471;
assign v_6308 = v_6304 & v_1479 & ~v_1480;
assign v_6309 = v_6304 & v_2092;
assign v_6311 = v_6310 & v_1469 & v_1470 & v_1485 & ~v_1486;
assign v_6313 = v_6312 & v_1492 & ~v_1493 & v_1511;
assign v_6314 = v_6312 & ~v_1494;
assign v_6315 = v_6312 & v_1502 & ~v_1503;
assign v_6316 = v_6312 & v_2100;
assign v_6318 = v_6317 & v_1492 & v_1493 & v_1508 & v_1509;
assign v_6319 = v_6312 & v_1492 & ~v_1493 & ~v_1511;
assign v_6320 = v_6317 & v_1492 & v_1493 & v_1508 & ~v_1509;
assign v_6323 = v_6321 & v_6322;
assign v_6324 = v_6321 & v_1515 & v_1516 & ~v_1517 & ~v_1518;
assign v_6325 = v_6321 & v_1515 & v_1516 & v_1517;
assign v_6326 = v_6321 & v_1515 & ~v_1516 & ~v_1520;
assign v_6328 = v_6327 & v_2113;
assign v_6329 = v_6310 & v_1469 & v_1470 & v_1485 & v_1486;
assign v_6330 = v_6302 & v_1446 & v_1447 & v_1462 & v_1463;
assign v_6333 = v_6332 & v_227;
assign v_6334 = v_6332 & ~v_227 & v_229 & v_262 & ~v_264;
assign v_6335 = v_6332 & ~v_227 & v_229 & v_262 & v_264;
assign v_6336 = v_6332 & ~v_227 & v_229 & ~v_262;
assign v_6337 = v_6332 & v_230;
assign v_6338 = v_6332 & ~v_230;
assign v_6341 = v_6339 & v_6340;
assign v_6342 = v_6339 & v_1540;
assign v_6343 = v_13121 & v_13122;
assign v_6345 = v_6344 & ~v_227 & ~v_229 & v_260;
assign v_6347 = v_6346 & v_267 & v_268;
assign v_6348 = v_6346 & v_267 & ~v_268;
assign v_6350 = v_6349 & ~v_279;
assign v_6352 = v_6349 & v_6351;
assign v_6353 = v_6349 & v_279 & v_291 & ~v_292 & v_300;
assign v_6356 = v_6354 & v_6355;
assign v_6357 = v_6354 & v_321 & v_322;
assign v_6358 = v_6354 & v_321 & ~v_322 & v_324;
assign v_6359 = v_6354 & v_321 & ~v_322 & ~v_324 & v_326;
assign v_6360 = v_6354 & v_321 & ~v_322 & ~v_324 & ~v_326;
assign v_6362 = v_6361 & v_1563;
assign v_6364 = v_6363 & ~v_308 & v_309 & v_329;
assign v_6367 = v_6365 & v_6366;
assign v_6368 = v_6365 & v_1570;
assign v_6370 = v_6369 & v_345 & v_346;
assign v_6371 = v_6369 & v_345 & ~v_346 & v_348;
assign v_6372 = v_6369 & v_345 & ~v_346 & ~v_348 & v_350;
assign v_6373 = v_6369 & v_356 & v_357;
assign v_6374 = v_6369 & v_359 & v_360;
assign v_6375 = v_6369 & v_359 & ~v_360 & v_362;
assign v_6376 = v_6369 & v_359 & ~v_360 & ~v_362 & v_364;
assign v_6377 = v_6369 & v_1582;
assign v_6379 = v_6378 & v_1585;
assign v_6381 = v_6380 & v_356 & ~v_357 & v_369 & v_370;
assign v_6382 = v_6380 & v_372 & v_373;
assign v_6383 = v_6380 & v_372 & ~v_373 & v_375;
assign v_6384 = v_6380 & v_372 & ~v_373 & ~v_375 & v_377;
assign v_6386 = v_6380 & v_6385;
assign v_6387 = v_13123 & v_13124;
assign v_6389 = v_6388 & v_384 & v_385;
assign v_6390 = v_6388 & v_384 & ~v_385;
assign v_6392 = v_6391 & v_1599;
assign v_6394 = v_13125 & v_13126;
assign v_6395 = v_6393 & v_391 & v_392;
assign v_6396 = v_6393 & v_391 & ~v_392 & v_394;
assign v_6397 = v_6393 & v_391 & ~v_392 & ~v_394 & v_396;
assign v_6398 = v_6393 & v_1606;
assign v_6400 = v_13127 & v_13128;
assign v_6402 = v_6401 & v_1611;
assign v_6404 = v_6403 & v_410 & v_411;
assign v_6405 = v_6403 & v_410 & ~v_411 & v_413;
assign v_6406 = v_6403 & v_410 & ~v_411 & ~v_413 & v_415;
assign v_6407 = v_6403 & v_421 & v_422;
assign v_6408 = v_6403 & v_424 & v_425;
assign v_6409 = v_6403 & v_424 & ~v_425 & v_427;
assign v_6410 = v_6403 & v_424 & ~v_425 & ~v_427 & v_429;
assign v_6411 = v_6403 & v_1621;
assign v_6413 = v_6412 & v_1624;
assign v_6415 = v_6414 & v_421 & ~v_422 & v_434 & v_435;
assign v_6416 = v_6414 & v_437 & v_438;
assign v_6417 = v_6414 & v_437 & ~v_438 & v_440;
assign v_6418 = v_6414 & v_437 & ~v_438 & ~v_440 & v_442;
assign v_6420 = v_6414 & v_6419;
assign v_6421 = v_13129 & v_13130;
assign v_6423 = v_6422 & v_449 & v_450;
assign v_6424 = v_6422 & v_449 & ~v_450;
assign v_6426 = v_6425 & v_1638;
assign v_6428 = v_13131 & v_13132;
assign v_6429 = v_6427 & v_456 & v_457;
assign v_6430 = v_6427 & v_456 & ~v_457 & v_459;
assign v_6431 = v_6427 & v_456 & ~v_457 & ~v_459 & v_461;
assign v_6432 = v_6427 & v_1645;
assign v_6434 = v_13133 & v_13134;
assign v_6436 = v_6435 & v_1650;
assign v_6438 = v_6437 & v_491;
assign v_6439 = v_6437 & ~v_491 & v_493 & v_526 & ~v_528;
assign v_6440 = v_6437 & ~v_491 & v_493 & v_526 & v_528;
assign v_6441 = v_6437 & ~v_491 & v_493 & ~v_526;
assign v_6442 = v_6437 & v_494;
assign v_6443 = v_6437 & ~v_494;
assign v_6446 = v_6444 & v_6445;
assign v_6447 = v_6444 & v_1666;
assign v_6448 = v_13135 & v_13136;
assign v_6450 = v_6449 & ~v_491 & ~v_493 & v_524;
assign v_6452 = v_6451 & v_531 & v_532;
assign v_6453 = v_6451 & v_531 & ~v_532;
assign v_6455 = v_6454 & v_546 & v_547;
assign v_6456 = v_6454 & v_546 & ~v_547 & ~v_551;
assign v_6458 = v_6457 & v_546 & ~v_547 & v_551;
assign v_6460 = v_6459 & v_554;
assign v_6462 = v_6461 & v_558 & v_559;
assign v_6463 = v_6461 & v_558 & ~v_559 & v_561;
assign v_6464 = v_6461 & v_1682;
assign v_6467 = v_6465 & v_6466;
assign v_6468 = v_6465 & v_1687;
assign v_6470 = v_6469 & v_588 & ~v_589 & ~v_591;
assign v_6471 = v_6469 & v_593 & ~v_594;
assign v_6472 = v_6469 & v_593 & v_594;
assign v_6473 = v_6469 & v_583;
assign v_6475 = v_6474 & v_604 & v_605;
assign v_6476 = v_6474 & v_604 & ~v_605 & ~v_609;
assign v_6478 = v_6477 & v_604 & ~v_605 & v_609;
assign v_6480 = v_6479 & v_612;
assign v_6482 = v_6481 & v_616 & v_617;
assign v_6483 = v_6481 & v_616 & ~v_617 & v_619;
assign v_6484 = v_6481 & v_1700;
assign v_6487 = v_6485 & v_6486;
assign v_6488 = v_6485 & v_1705;
assign v_6490 = v_2 & v_6489;
assign v_6491 = v_641 & v_6469;
assign v_6492 = v_643 & v_6454;
assign v_6493 = v_645 & v_6454;
assign v_6494 = v_647 & v_6454;
assign v_6495 = v_649 & v_6454;
assign v_6496 = ~v_649 & v_6437;
assign v_6498 = ~v_647 & v_6497;
assign v_6500 = ~v_645 & v_6499;
assign v_6502 = ~v_643 & v_6501;
assign v_6504 = ~v_641 & v_6503;
assign v_6506 = ~v_2 & v_6505;
assign v_6508 = v_6507 & ~v_669;
assign v_6509 = v_13137 & v_13138;
assign v_6510 = v_6507 & v_669 & v_670 & v_672 & v_674;
assign v_6511 = v_13139 & v_13140;
assign v_6513 = v_6512 & v_679 & ~v_680 & v_682;
assign v_6514 = v_6512 & v_689 & ~v_690 & ~v_692;
assign v_6515 = v_6512 & v_694 & ~v_695;
assign v_6516 = v_6512 & v_694 & v_695;
assign v_6517 = v_6512 & v_684;
assign v_6519 = v_6518 & v_1737;
assign v_6521 = v_6520 & v_1740;
assign v_6522 = v_6512 & v_679 & v_680;
assign v_6523 = v_6507 & v_1743;
assign v_6525 = v_6524 & ~v_705;
assign v_6526 = v_6524 & v_710 & v_711;
assign v_6527 = v_6524 & v_710 & ~v_711 & ~v_715;
assign v_6529 = v_6528 & v_710 & ~v_711 & v_715;
assign v_6531 = v_6530 & v_718;
assign v_6533 = v_6532 & v_705 & v_722 & v_723 & ~v_724;
assign v_6535 = v_6532 & v_6534;
assign v_6536 = v_6532 & v_750 & v_751;
assign v_6537 = v_6532 & v_750 & ~v_751;
assign v_6539 = v_6538 & v_763 & v_764;
assign v_6540 = v_6538 & v_763 & ~v_764;
assign v_6542 = v_6541 & v_745 & v_758 & v_771;
assign v_6543 = v_13141 & v_13142;
assign v_6544 = v_6532 & v_779 & v_780;
assign v_6545 = v_6532 & v_779 & ~v_780 & ~v_784;
assign v_6547 = v_6546 & v_779 & ~v_780 & v_784;
assign v_6549 = v_6548 & v_787;
assign v_6551 = v_6550 & v_1764;
assign v_6553 = v_6552 & v_798 & ~v_799 & v_817;
assign v_6554 = v_6552 & v_798 & ~v_799 & ~v_817;
assign v_6555 = v_6552 & ~v_800;
assign v_6556 = v_6552 & v_808 & ~v_809;
assign v_6557 = v_6552 & v_1771;
assign v_6559 = v_6558 & v_798 & v_799 & v_814 & ~v_815;
assign v_6561 = v_6560 & v_821 & ~v_822 & v_840;
assign v_6562 = v_6560 & v_821 & ~v_822 & ~v_840;
assign v_6563 = v_6560 & ~v_823;
assign v_6564 = v_6560 & v_831 & ~v_832;
assign v_6565 = v_6560 & v_1780;
assign v_6567 = v_6566 & v_821 & v_822 & v_837 & ~v_838;
assign v_6569 = v_6568 & v_844 & ~v_845 & v_863;
assign v_6570 = v_6568 & ~v_846;
assign v_6571 = v_6568 & v_854 & ~v_855;
assign v_6572 = v_6568 & v_1788;
assign v_6574 = v_6573 & v_844 & v_845 & v_860 & v_861;
assign v_6575 = v_6568 & v_844 & ~v_845 & ~v_863;
assign v_6576 = v_6573 & v_844 & v_845 & v_860 & ~v_861;
assign v_6579 = v_6577 & v_6578;
assign v_6580 = v_6577 & v_867 & v_868 & ~v_869 & ~v_870;
assign v_6581 = v_6577 & v_867 & v_868 & v_869;
assign v_6582 = v_6577 & v_867 & ~v_868 & ~v_872;
assign v_6584 = v_6583 & v_1801;
assign v_6585 = v_6566 & v_821 & v_822 & v_837 & v_838;
assign v_6586 = v_6558 & v_798 & v_799 & v_814 & v_815;
assign v_6588 = v_6587 & v_879 & ~v_880 & v_898;
assign v_6589 = v_6587 & v_879 & ~v_880 & ~v_898;
assign v_6590 = v_6587 & ~v_881;
assign v_6591 = v_6587 & v_889 & ~v_890;
assign v_6592 = v_6587 & v_1810;
assign v_6594 = v_6593 & v_879 & v_880 & v_895 & ~v_896;
assign v_6596 = v_6595 & v_902 & ~v_903 & v_921;
assign v_6597 = v_6595 & v_902 & ~v_903 & ~v_921;
assign v_6598 = v_6595 & ~v_904;
assign v_6599 = v_6595 & v_912 & ~v_913;
assign v_6600 = v_6595 & v_1819;
assign v_6602 = v_6601 & v_902 & v_903 & v_918 & ~v_919;
assign v_6604 = v_6603 & v_925 & ~v_926 & v_944;
assign v_6605 = v_6603 & ~v_927;
assign v_6606 = v_6603 & v_935 & ~v_936;
assign v_6607 = v_6603 & v_1827;
assign v_6609 = v_6608 & v_925 & v_926 & v_941 & v_942;
assign v_6610 = v_6603 & v_925 & ~v_926 & ~v_944;
assign v_6611 = v_6608 & v_925 & v_926 & v_941 & ~v_942;
assign v_6614 = v_6612 & v_6613;
assign v_6615 = v_6612 & v_948 & v_949 & ~v_950 & ~v_951;
assign v_6616 = v_6612 & v_948 & v_949 & v_950;
assign v_6617 = v_6612 & v_948 & ~v_949 & ~v_953;
assign v_6619 = v_6618 & v_1840;
assign v_6620 = v_6601 & v_902 & v_903 & v_918 & v_919;
assign v_6621 = v_6593 & v_879 & v_880 & v_895 & v_896;
assign v_6623 = v_6622 & v_960 & ~v_961 & v_979;
assign v_6624 = v_6622 & v_960 & ~v_961 & ~v_979;
assign v_6625 = v_6622 & ~v_962;
assign v_6626 = v_6622 & v_970 & ~v_971;
assign v_6627 = v_6622 & v_1849;
assign v_6629 = v_6628 & v_960 & v_961 & v_976 & ~v_977;
assign v_6631 = v_6630 & v_983 & ~v_984 & v_1002;
assign v_6632 = v_6630 & v_983 & ~v_984 & ~v_1002;
assign v_6633 = v_6630 & ~v_985;
assign v_6634 = v_6630 & v_993 & ~v_994;
assign v_6635 = v_6630 & v_1858;
assign v_6637 = v_6636 & v_983 & v_984 & v_999 & ~v_1000;
assign v_6639 = v_6638 & v_1006 & ~v_1007 & v_1025;
assign v_6640 = v_6638 & ~v_1008;
assign v_6641 = v_6638 & v_1016 & ~v_1017;
assign v_6642 = v_6638 & v_1866;
assign v_6644 = v_6643 & v_1006 & v_1007 & v_1022 & v_1023;
assign v_6645 = v_6638 & v_1006 & ~v_1007 & ~v_1025;
assign v_6646 = v_6643 & v_1006 & v_1007 & v_1022 & ~v_1023;
assign v_6649 = v_6647 & v_6648;
assign v_6650 = v_6647 & v_1029 & v_1030 & ~v_1031 & ~v_1032;
assign v_6651 = v_6647 & v_1029 & v_1030 & v_1031;
assign v_6652 = v_6647 & v_1029 & ~v_1030 & ~v_1034;
assign v_6654 = v_6653 & v_1879;
assign v_6655 = v_6636 & v_983 & v_984 & v_999 & v_1000;
assign v_6656 = v_6628 & v_960 & v_961 & v_976 & v_977;
assign v_6658 = v_6657 & v_1041 & ~v_1042 & v_1060;
assign v_6659 = v_6657 & v_1041 & ~v_1042 & ~v_1060;
assign v_6660 = v_6657 & ~v_1043;
assign v_6661 = v_6657 & v_1051 & ~v_1052;
assign v_6662 = v_6657 & v_1888;
assign v_6664 = v_6663 & v_1041 & v_1042 & v_1057 & ~v_1058;
assign v_6666 = v_6665 & v_1064 & ~v_1065 & v_1083;
assign v_6667 = v_6665 & v_1064 & ~v_1065 & ~v_1083;
assign v_6668 = v_6665 & ~v_1066;
assign v_6669 = v_6665 & v_1074 & ~v_1075;
assign v_6670 = v_6665 & v_1897;
assign v_6672 = v_6671 & v_1064 & v_1065 & v_1080 & ~v_1081;
assign v_6674 = v_6673 & v_1087 & ~v_1088 & v_1106;
assign v_6675 = v_6673 & ~v_1089;
assign v_6676 = v_6673 & v_1097 & ~v_1098;
assign v_6677 = v_6673 & v_1905;
assign v_6679 = v_6678 & v_1087 & v_1088 & v_1103 & v_1104;
assign v_6680 = v_6673 & v_1087 & ~v_1088 & ~v_1106;
assign v_6681 = v_6678 & v_1087 & v_1088 & v_1103 & ~v_1104;
assign v_6684 = v_6682 & v_6683;
assign v_6685 = v_6682 & v_1110 & v_1111 & ~v_1112 & ~v_1113;
assign v_6686 = v_6682 & v_1110 & v_1111 & v_1112;
assign v_6687 = v_6682 & v_1110 & ~v_1111 & ~v_1115;
assign v_6689 = v_6688 & v_1918;
assign v_6690 = v_6671 & v_1064 & v_1065 & v_1080 & v_1081;
assign v_6691 = v_6663 & v_1041 & v_1042 & v_1057 & v_1058;
assign v_6693 = v_6692 & v_1122 & ~v_1123 & v_1141;
assign v_6694 = v_6692 & v_1122 & ~v_1123 & ~v_1141;
assign v_6695 = v_6692 & ~v_1124;
assign v_6696 = v_6692 & v_1132 & ~v_1133;
assign v_6697 = v_6692 & v_1927;
assign v_6699 = v_6698 & v_1122 & v_1123 & v_1138 & ~v_1139;
assign v_6701 = v_6700 & v_1145 & ~v_1146 & v_1164;
assign v_6702 = v_6700 & v_1145 & ~v_1146 & ~v_1164;
assign v_6703 = v_6700 & ~v_1147;
assign v_6704 = v_6700 & v_1155 & ~v_1156;
assign v_6705 = v_6700 & v_1936;
assign v_6707 = v_6706 & v_1145 & v_1146 & v_1161 & ~v_1162;
assign v_6709 = v_6708 & v_1168 & ~v_1169 & v_1187;
assign v_6710 = v_6708 & ~v_1170;
assign v_6711 = v_6708 & v_1178 & ~v_1179;
assign v_6712 = v_6708 & v_1944;
assign v_6714 = v_6713 & v_1168 & v_1169 & v_1184 & v_1185;
assign v_6715 = v_6708 & v_1168 & ~v_1169 & ~v_1187;
assign v_6716 = v_6713 & v_1168 & v_1169 & v_1184 & ~v_1185;
assign v_6719 = v_6717 & v_6718;
assign v_6720 = v_6717 & v_1191 & v_1192 & ~v_1193 & ~v_1194;
assign v_6721 = v_6717 & v_1191 & v_1192 & v_1193;
assign v_6722 = v_6717 & v_1191 & ~v_1192 & ~v_1196;
assign v_6724 = v_6723 & v_1957;
assign v_6725 = v_6706 & v_1145 & v_1146 & v_1161 & v_1162;
assign v_6726 = v_6698 & v_1122 & v_1123 & v_1138 & v_1139;
assign v_6728 = v_6727 & v_1203 & ~v_1204 & v_1222;
assign v_6729 = v_6727 & v_1203 & ~v_1204 & ~v_1222;
assign v_6730 = v_6727 & ~v_1205;
assign v_6731 = v_6727 & v_1213 & ~v_1214;
assign v_6732 = v_6727 & v_1966;
assign v_6734 = v_6733 & v_1203 & v_1204 & v_1219 & ~v_1220;
assign v_6736 = v_6735 & v_1226 & ~v_1227 & v_1245;
assign v_6737 = v_6735 & v_1226 & ~v_1227 & ~v_1245;
assign v_6738 = v_6735 & ~v_1228;
assign v_6739 = v_6735 & v_1236 & ~v_1237;
assign v_6740 = v_6735 & v_1975;
assign v_6742 = v_6741 & v_1226 & v_1227 & v_1242 & ~v_1243;
assign v_6744 = v_6743 & v_1249 & ~v_1250 & v_1268;
assign v_6745 = v_6743 & ~v_1251;
assign v_6746 = v_6743 & v_1259 & ~v_1260;
assign v_6747 = v_6743 & v_1983;
assign v_6749 = v_6748 & v_1249 & v_1250 & v_1265 & v_1266;
assign v_6750 = v_6743 & v_1249 & ~v_1250 & ~v_1268;
assign v_6751 = v_6748 & v_1249 & v_1250 & v_1265 & ~v_1266;
assign v_6754 = v_6752 & v_6753;
assign v_6755 = v_6752 & v_1272 & v_1273 & ~v_1274 & ~v_1275;
assign v_6756 = v_6752 & v_1272 & v_1273 & v_1274;
assign v_6757 = v_6752 & v_1272 & ~v_1273 & ~v_1277;
assign v_6759 = v_6758 & v_1996;
assign v_6760 = v_6741 & v_1226 & v_1227 & v_1242 & v_1243;
assign v_6761 = v_6733 & v_1203 & v_1204 & v_1219 & v_1220;
assign v_6763 = v_6762 & v_1284 & ~v_1285 & v_1303;
assign v_6764 = v_6762 & v_1284 & ~v_1285 & ~v_1303;
assign v_6765 = v_6762 & ~v_1286;
assign v_6766 = v_6762 & v_1294 & ~v_1295;
assign v_6767 = v_6762 & v_2005;
assign v_6769 = v_6768 & v_1284 & v_1285 & v_1300 & ~v_1301;
assign v_6771 = v_6770 & v_1307 & ~v_1308 & v_1326;
assign v_6772 = v_6770 & v_1307 & ~v_1308 & ~v_1326;
assign v_6773 = v_6770 & ~v_1309;
assign v_6774 = v_6770 & v_1317 & ~v_1318;
assign v_6775 = v_6770 & v_2014;
assign v_6777 = v_6776 & v_1307 & v_1308 & v_1323 & ~v_1324;
assign v_6779 = v_6778 & v_1330 & ~v_1331 & v_1349;
assign v_6780 = v_6778 & ~v_1332;
assign v_6781 = v_6778 & v_1340 & ~v_1341;
assign v_6782 = v_6778 & v_2022;
assign v_6784 = v_6783 & v_1330 & v_1331 & v_1346 & v_1347;
assign v_6785 = v_6778 & v_1330 & ~v_1331 & ~v_1349;
assign v_6786 = v_6783 & v_1330 & v_1331 & v_1346 & ~v_1347;
assign v_6789 = v_6787 & v_6788;
assign v_6790 = v_6787 & v_1353 & v_1354 & ~v_1355 & ~v_1356;
assign v_6791 = v_6787 & v_1353 & v_1354 & v_1355;
assign v_6792 = v_6787 & v_1353 & ~v_1354 & ~v_1358;
assign v_6794 = v_6793 & v_2035;
assign v_6795 = v_6776 & v_1307 & v_1308 & v_1323 & v_1324;
assign v_6796 = v_6768 & v_1284 & v_1285 & v_1300 & v_1301;
assign v_6798 = v_6797 & v_1365 & ~v_1366 & v_1384;
assign v_6799 = v_6797 & v_1365 & ~v_1366 & ~v_1384;
assign v_6800 = v_6797 & ~v_1367;
assign v_6801 = v_6797 & v_1375 & ~v_1376;
assign v_6802 = v_6797 & v_2044;
assign v_6804 = v_6803 & v_1365 & v_1366 & v_1381 & ~v_1382;
assign v_6806 = v_6805 & v_1388 & ~v_1389 & v_1407;
assign v_6807 = v_6805 & v_1388 & ~v_1389 & ~v_1407;
assign v_6808 = v_6805 & ~v_1390;
assign v_6809 = v_6805 & v_1398 & ~v_1399;
assign v_6810 = v_6805 & v_2053;
assign v_6812 = v_6811 & v_1388 & v_1389 & v_1404 & ~v_1405;
assign v_6814 = v_6813 & v_1411 & ~v_1412 & v_1430;
assign v_6815 = v_6813 & ~v_1413;
assign v_6816 = v_6813 & v_1421 & ~v_1422;
assign v_6817 = v_6813 & v_2061;
assign v_6819 = v_6818 & v_1411 & v_1412 & v_1427 & v_1428;
assign v_6820 = v_6813 & v_1411 & ~v_1412 & ~v_1430;
assign v_6821 = v_6818 & v_1411 & v_1412 & v_1427 & ~v_1428;
assign v_6824 = v_6822 & v_6823;
assign v_6825 = v_6822 & v_1434 & v_1435 & ~v_1436 & ~v_1437;
assign v_6826 = v_6822 & v_1434 & v_1435 & v_1436;
assign v_6827 = v_6822 & v_1434 & ~v_1435 & ~v_1439;
assign v_6829 = v_6828 & v_2074;
assign v_6830 = v_6811 & v_1388 & v_1389 & v_1404 & v_1405;
assign v_6831 = v_6803 & v_1365 & v_1366 & v_1381 & v_1382;
assign v_6833 = v_6832 & v_1446 & ~v_1447 & v_1465;
assign v_6834 = v_6832 & v_1446 & ~v_1447 & ~v_1465;
assign v_6835 = v_6832 & ~v_1448;
assign v_6836 = v_6832 & v_1456 & ~v_1457;
assign v_6837 = v_6832 & v_2083;
assign v_6839 = v_6838 & v_1446 & v_1447 & v_1462 & ~v_1463;
assign v_6841 = v_6840 & v_1469 & ~v_1470 & v_1488;
assign v_6842 = v_6840 & v_1469 & ~v_1470 & ~v_1488;
assign v_6843 = v_6840 & ~v_1471;
assign v_6844 = v_6840 & v_1479 & ~v_1480;
assign v_6845 = v_6840 & v_2092;
assign v_6847 = v_6846 & v_1469 & v_1470 & v_1485 & ~v_1486;
assign v_6849 = v_6848 & v_1492 & ~v_1493 & v_1511;
assign v_6850 = v_6848 & ~v_1494;
assign v_6851 = v_6848 & v_1502 & ~v_1503;
assign v_6852 = v_6848 & v_2100;
assign v_6854 = v_6853 & v_1492 & v_1493 & v_1508 & v_1509;
assign v_6855 = v_6848 & v_1492 & ~v_1493 & ~v_1511;
assign v_6856 = v_6853 & v_1492 & v_1493 & v_1508 & ~v_1509;
assign v_6859 = v_6857 & v_6858;
assign v_6860 = v_6857 & v_1515 & v_1516 & ~v_1517 & ~v_1518;
assign v_6861 = v_6857 & v_1515 & v_1516 & v_1517;
assign v_6862 = v_6857 & v_1515 & ~v_1516 & ~v_1520;
assign v_6864 = v_6863 & v_2113;
assign v_6865 = v_6846 & v_1469 & v_1470 & v_1485 & v_1486;
assign v_6866 = v_6838 & v_1446 & v_1447 & v_1462 & v_1463;
assign v_6872 = ~v_6870 & ~v_6871;
assign v_6875 = ~v_6873 & v_6874;
assign v_6876 = ~v_6872 & ~v_6875;
assign v_6877 = ~v_6870 & ~v_6871;
assign v_6878 = ~v_6873 & v_6874;
assign v_6879 = ~v_6877 & ~v_6878;
assign v_6880 = v_6876 & v_6879;
assign v_6881 = ~v_6870 & ~v_6871;
assign v_6882 = ~v_6873 & v_6874;
assign v_6883 = ~v_6881 & ~v_6882;
assign v_6884 = v_6880 & v_6883;
assign v_6885 = ~v_6870 & ~v_6871;
assign v_6886 = ~v_6873 & v_6874;
assign v_6887 = ~v_6885 & ~v_6886;
assign v_6888 = v_6884 & v_6887;
assign v_6889 = ~v_6870 & ~v_6871;
assign v_6890 = ~v_6873 & v_6874;
assign v_6891 = ~v_6889 & ~v_6890;
assign v_6892 = v_6888 & v_6891;
assign v_6893 = ~v_6870 & ~v_6871;
assign v_6894 = ~v_6873 & v_6874;
assign v_6895 = ~v_6893 & ~v_6894;
assign v_6896 = v_6892 & v_6895;
assign v_6897 = ~v_6870 & ~v_6871;
assign v_6898 = ~v_6873 & v_6874;
assign v_6899 = ~v_6897 & ~v_6898;
assign v_6900 = v_6896 & v_6899;
assign v_6901 = ~v_6870 & ~v_6871;
assign v_6902 = ~v_6873 & v_6874;
assign v_6903 = ~v_6901 & ~v_6902;
assign v_6904 = v_6900 & v_6903;
assign v_6905 = ~v_6870 & ~v_6871;
assign v_6906 = ~v_6873 & v_6874;
assign v_6907 = ~v_6905 & ~v_6906;
assign v_6908 = v_6904 & v_6907;
assign v_6909 = ~v_6870 & ~v_6871;
assign v_6910 = ~v_6873 & v_6874;
assign v_6911 = ~v_6909 & ~v_6910;
assign v_6912 = v_6908 & v_6911;
assign v_6913 = ~v_6870 & ~v_6871;
assign v_6914 = ~v_6873 & v_6874;
assign v_6915 = ~v_6913 & ~v_6914;
assign v_6916 = v_6912 & v_6915;
assign v_6917 = ~v_6870 & ~v_6871;
assign v_6918 = ~v_6873 & v_6874;
assign v_6919 = ~v_6917 & ~v_6918;
assign v_6920 = v_6916 & v_6919;
assign v_6921 = ~v_6870 & ~v_6871;
assign v_6922 = ~v_6873 & v_6874;
assign v_6923 = ~v_6921 & ~v_6922;
assign v_6924 = v_6920 & v_6923;
assign v_6925 = ~v_6870 & ~v_6871;
assign v_6926 = ~v_6873 & v_6874;
assign v_6927 = ~v_6925 & ~v_6926;
assign v_6928 = v_6924 & v_6927;
assign v_6929 = ~v_6870 & ~v_6871;
assign v_6930 = ~v_6873 & v_6874;
assign v_6931 = ~v_6929 & ~v_6930;
assign v_6932 = v_6928 & v_6931;
assign v_6933 = ~v_6870 & ~v_6871;
assign v_6934 = ~v_6873 & v_6874;
assign v_6935 = ~v_6933 & ~v_6934;
assign v_6936 = v_6932 & v_6935;
assign v_6937 = ~v_6870 & ~v_6871;
assign v_6938 = ~v_6873 & v_6874;
assign v_6939 = ~v_6937 & ~v_6938;
assign v_6940 = v_6936 & v_6939;
assign v_6941 = ~v_6870 & ~v_6871;
assign v_6942 = ~v_6873 & v_6874;
assign v_6943 = ~v_6941 & ~v_6942;
assign v_6944 = v_6940 & v_6943;
assign v_6945 = ~v_6870 & ~v_6871;
assign v_6946 = ~v_6873 & v_6874;
assign v_6947 = ~v_6945 & ~v_6946;
assign v_6948 = v_6944 & v_6947;
assign v_6949 = ~v_6870 & ~v_6871;
assign v_6950 = ~v_6873 & v_6874;
assign v_6951 = ~v_6949 & ~v_6950;
assign v_6952 = v_6948 & v_6951;
assign v_6953 = ~v_6870 & ~v_6871;
assign v_6954 = ~v_6873 & v_6874;
assign v_6955 = ~v_6953 & ~v_6954;
assign v_6956 = v_6952 & v_6955;
assign v_6957 = ~v_6870 & ~v_6871;
assign v_6958 = ~v_6873 & v_6874;
assign v_6959 = ~v_6957 & ~v_6958;
assign v_6960 = v_6956 & v_6959;
assign v_6961 = ~v_6870 & ~v_6871;
assign v_6962 = ~v_6873 & v_6874;
assign v_6963 = ~v_6961 & ~v_6962;
assign v_6964 = v_6960 & v_6963;
assign v_6965 = ~v_6870 & ~v_6871;
assign v_6966 = ~v_6873 & v_6874;
assign v_6967 = ~v_6965 & ~v_6966;
assign v_6968 = v_6964 & v_6967;
assign v_6969 = ~v_6870 & ~v_6871;
assign v_6970 = ~v_6873 & v_6874;
assign v_6971 = ~v_6969 & ~v_6970;
assign v_6972 = v_6968 & v_6971;
assign v_6973 = ~v_6870 & ~v_6871;
assign v_6974 = ~v_6873 & v_6874;
assign v_6975 = ~v_6973 & ~v_6974;
assign v_6976 = v_6972 & v_6975;
assign v_6977 = ~v_6870 & ~v_6871;
assign v_6978 = ~v_6873 & v_6874;
assign v_6979 = ~v_6977 & ~v_6978;
assign v_6980 = v_6976 & v_6979;
assign v_6981 = ~v_6870 & ~v_6871;
assign v_6982 = ~v_6873 & v_6874;
assign v_6983 = ~v_6981 & ~v_6982;
assign v_6984 = v_6980 & v_6983;
assign v_6985 = ~v_6870 & ~v_6871;
assign v_6986 = ~v_6873 & v_6874;
assign v_6987 = ~v_6985 & ~v_6986;
assign v_6988 = v_6984 & v_6987;
assign v_6989 = ~v_6870 & ~v_6871;
assign v_6990 = ~v_6873 & v_6874;
assign v_6991 = ~v_6989 & ~v_6990;
assign v_6992 = v_6988 & v_6991;
assign v_6993 = ~v_6870 & ~v_6871;
assign v_6994 = ~v_6873 & v_6874;
assign v_6995 = ~v_6993 & ~v_6994;
assign v_6996 = v_6992 & v_6995;
assign v_6997 = ~v_6870 & ~v_6871;
assign v_6998 = ~v_6873 & v_6874;
assign v_6999 = ~v_6997 & ~v_6998;
assign v_7000 = v_6996 & v_6999;
assign v_7001 = ~v_6870 & ~v_6871;
assign v_7002 = ~v_6873 & v_6874;
assign v_7003 = ~v_7001 & ~v_7002;
assign v_7004 = v_7000 & v_7003;
assign v_7005 = ~v_6870 & ~v_6871;
assign v_7006 = ~v_6873 & v_6874;
assign v_7007 = ~v_7005 & ~v_7006;
assign v_7008 = v_7004 & v_7007;
assign v_7009 = ~v_6870 & ~v_6871;
assign v_7010 = ~v_6873 & v_6874;
assign v_7011 = ~v_7009 & ~v_7010;
assign v_7012 = v_7008 & v_7011;
assign v_7013 = ~v_6870 & ~v_6871;
assign v_7014 = ~v_6873 & v_6874;
assign v_7015 = ~v_7013 & ~v_7014;
assign v_7016 = v_7012 & v_7015;
assign v_7017 = ~v_6870 & ~v_6871;
assign v_7018 = ~v_6873 & v_6874;
assign v_7019 = ~v_7017 & ~v_7018;
assign v_7020 = v_7016 & v_7019;
assign v_7021 = ~v_6870 & ~v_6871;
assign v_7022 = ~v_6873 & v_6874;
assign v_7023 = ~v_7021 & ~v_7022;
assign v_7024 = v_7020 & v_7023;
assign v_7025 = ~v_6870 & ~v_6871;
assign v_7026 = ~v_6873 & v_6874;
assign v_7027 = ~v_7025 & ~v_7026;
assign v_7028 = v_7024 & v_7027;
assign v_7029 = ~v_6870 & ~v_6871;
assign v_7030 = ~v_6873 & v_6874;
assign v_7031 = ~v_7029 & ~v_7030;
assign v_7032 = v_7028 & v_7031;
assign v_7033 = ~v_6870 & ~v_6871;
assign v_7034 = ~v_6873 & v_6874;
assign v_7035 = ~v_7033 & ~v_7034;
assign v_7036 = v_7032 & v_7035;
assign v_7037 = ~v_6870 & ~v_6871;
assign v_7038 = ~v_6873 & v_6874;
assign v_7039 = ~v_7037 & ~v_7038;
assign v_7040 = v_7036 & v_7039;
assign v_7041 = ~v_6870 & ~v_6871;
assign v_7042 = ~v_6873 & v_6874;
assign v_7043 = ~v_7041 & ~v_7042;
assign v_7044 = v_7040 & v_7043;
assign v_7045 = ~v_6870 & ~v_6871;
assign v_7046 = ~v_6873 & v_6874;
assign v_7047 = ~v_7045 & ~v_7046;
assign v_7048 = v_7044 & v_7047;
assign v_7049 = ~v_6870 & ~v_6871;
assign v_7050 = ~v_6873 & v_6874;
assign v_7051 = ~v_7049 & ~v_7050;
assign v_7052 = v_7048 & v_7051;
assign v_7053 = ~v_6870 & ~v_6871;
assign v_7054 = ~v_6873 & v_6874;
assign v_7055 = ~v_7053 & ~v_7054;
assign v_7056 = v_7052 & v_7055;
assign v_7057 = ~v_6870 & ~v_6871;
assign v_7058 = ~v_6873 & v_6874;
assign v_7059 = ~v_7057 & ~v_7058;
assign v_7060 = v_7056 & v_7059;
assign v_7061 = ~v_6870 & ~v_6871;
assign v_7062 = ~v_6873 & v_6874;
assign v_7063 = ~v_7061 & ~v_7062;
assign v_7064 = v_7060 & v_7063;
assign v_7065 = ~v_6870 & ~v_6871;
assign v_7066 = ~v_6873 & v_6874;
assign v_7067 = ~v_7065 & ~v_7066;
assign v_7068 = v_7064 & v_7067;
assign v_7069 = ~v_6873 & v_6874;
assign v_7070 = v_7068 & ~v_7069;
assign v_7071 = ~v_6873 & v_6874;
assign v_7072 = v_7070 & ~v_7071;
assign v_7073 = ~v_6873 & v_6874;
assign v_7074 = v_7072 & ~v_7073;
assign v_7075 = ~v_6873 & v_6874;
assign v_7076 = v_7074 & ~v_7075;
assign v_7077 = ~v_6873 & v_6874;
assign v_7078 = v_7076 & ~v_7077;
assign v_7081 = v_7079 & v_7080;
assign v_7082 = v_7079 & ~v_7080;
assign v_7084 = v_7078 & v_7083;
assign v_7088 = v_7087;
assign v_7089 = ~v_7087;
assign v_7094 = v_7093;
assign v_7099 = ~v_7098;
assign v_7101 = v_7098 & v_7100;
assign v_7104 = v_7098 & ~v_7100 & v_7102 & v_7103;
assign v_7106 = v_7098 & ~v_7100 & v_7102 & ~v_7103 & ~v_7105;
assign v_7108 = v_7098 & ~v_7100 & ~v_7102 & ~v_7107;
assign v_7110 = v_7098 & ~v_7100 & ~v_7102 & v_7107 & v_7109;
assign v_7112 = v_13143 & v_13144;
assign v_7114 = v_13145 & v_13146;
assign v_7118 = v_13147 & v_13148;
assign v_7119 = v_13149 & v_13150;
assign v_7122 = v_7120 & v_7121;
assign v_7123 = v_7120 & ~v_7121;
assign v_7125 = v_13151 & v_13152;
assign v_7127 = ~v_7093 & ~v_7095 & v_7126;
assign v_7129 = ~v_7093 & v_7095 & ~v_7128;
assign v_7131 = ~v_7093 & v_7095 & v_7128 & ~v_7130;
assign v_7132 = ~v_7093 & v_7095 & v_7128 & v_7130;
assign v_7135 = v_7133 & v_7134;
assign v_7136 = v_7133 & ~v_7134;
assign v_7141 = v_7090 & v_7137 & v_7140;
assign v_7142 = v_7090 & v_7137 & ~v_7140;
assign v_7144 = v_7084 & v_7143;
assign v_7148 = v_7146 & v_7147;
assign v_7150 = v_7146 & ~v_7147 & v_7149;
assign v_7153 = v_7151 & ~v_7152;
assign v_7155 = v_7151 & v_7152 & v_7154;
assign v_7156 = v_7151 & v_7152 & ~v_7154;
assign v_7160 = v_7145 & v_7157 & v_7158 & v_7159;
assign v_7162 = v_7145 & v_7157 & v_7158 & ~v_7159 & v_7161;
assign v_7165 = ~v_7163 & v_7164;
assign v_7167 = v_7145 & v_7157 & ~v_7158 & v_7166;
assign v_7170 = v_7168 & v_7169;
assign v_7171 = v_7168 & ~v_7169;
assign v_7173 = v_7144 & v_7172;
assign v_7176 = ~v_7174 & ~v_7175;
assign v_7179 = v_7177 & v_7178;
assign v_7180 = v_7177 & ~v_7178;
assign v_7183 = v_7181 & ~v_7182;
assign v_7185 = v_7181 & v_7182 & v_7184;
assign v_7186 = v_7181 & v_7182 & ~v_7184;
assign v_7189 = v_7187 & v_7188;
assign v_7191 = v_7187 & ~v_7188 & v_7190;
assign v_7193 = v_7187 & ~v_7188 & ~v_7190 & v_7192;
assign v_7194 = v_7187 & ~v_7188 & ~v_7190 & ~v_7192;
assign v_7196 = ~v_7174 & v_7175 & v_7195;
assign v_7198 = v_7173 & v_7197;
assign v_7201 = v_7199 & ~v_7200;
assign v_7203 = v_7199 & v_7200 & ~v_7202;
assign v_7207 = v_7199 & v_7200 & v_7202 & v_7206;
assign v_7208 = v_7199 & v_7200 & v_7202 & ~v_7206;
assign v_7210 = v_7198 & v_7209;
assign v_7213 = v_7211 & v_7212;
assign v_7215 = v_7211 & ~v_7212 & v_7214;
assign v_7217 = v_7211 & ~v_7212 & ~v_7214 & v_7216;
assign v_7219 = v_7211 & ~v_7212 & ~v_7214 & ~v_7216 & v_7218;
assign v_7221 = v_13153 & v_13154;
assign v_7224 = v_7222 & v_7223;
assign v_7227 = v_7225 & v_7226;
assign v_7229 = v_7225 & ~v_7226 & v_7228;
assign v_7231 = v_7225 & ~v_7226 & ~v_7228 & v_7230;
assign v_7233 = v_7225 & ~v_7226 & ~v_7228 & ~v_7230 & v_7232;
assign v_7234 = v_7225 & ~v_7226 & ~v_7228 & ~v_7230 & ~v_7232;
assign v_7237 = v_7222 & ~v_7223 & v_7235 & v_7236;
assign v_7240 = v_7238 & v_7239;
assign v_7242 = v_7238 & ~v_7239 & v_7241;
assign v_7244 = v_7238 & ~v_7239 & ~v_7241 & v_7243;
assign v_7246 = v_7238 & ~v_7239 & ~v_7241 & ~v_7243 & v_7245;
assign v_7248 = v_13155 & v_13156;
assign v_7249 = v_13157 & v_13158;
assign v_7252 = v_7250 & v_7251;
assign v_7253 = v_7250 & ~v_7251;
assign v_7256 = v_13159 & v_13160;
assign v_7259 = v_7257 & v_7258;
assign v_7261 = v_7257 & ~v_7258 & v_7260;
assign v_7263 = v_7257 & ~v_7258 & ~v_7260 & v_7262;
assign v_7265 = v_7257 & ~v_7258 & ~v_7260 & ~v_7262 & ~v_7264;
assign v_7267 = v_13161 & v_13162;
assign v_7268 = v_13163 & v_13164;
assign v_7270 = v_13165 & v_13166;
assign v_7273 = v_7271 & v_7272;
assign v_7274 = v_7271 & ~v_7272;
assign v_7278 = v_7276 & v_7277;
assign v_7280 = v_7276 & ~v_7277 & v_7279;
assign v_7282 = v_7276 & ~v_7277 & ~v_7279 & v_7281;
assign v_7284 = v_7276 & ~v_7277 & ~v_7279 & ~v_7281 & v_7283;
assign v_7286 = v_13167 & v_13168;
assign v_7289 = v_7287 & v_7288;
assign v_7292 = v_7290 & v_7291;
assign v_7294 = v_7290 & ~v_7291 & v_7293;
assign v_7296 = v_7290 & ~v_7291 & ~v_7293 & v_7295;
assign v_7298 = v_7290 & ~v_7291 & ~v_7293 & ~v_7295 & v_7297;
assign v_7299 = v_7290 & ~v_7291 & ~v_7293 & ~v_7295 & ~v_7297;
assign v_7302 = v_7287 & ~v_7288 & v_7300 & v_7301;
assign v_7305 = v_7303 & v_7304;
assign v_7307 = v_7303 & ~v_7304 & v_7306;
assign v_7309 = v_7303 & ~v_7304 & ~v_7306 & v_7308;
assign v_7311 = v_7303 & ~v_7304 & ~v_7306 & ~v_7308 & v_7310;
assign v_7313 = v_13169 & v_13170;
assign v_7314 = v_13171 & v_13172;
assign v_7317 = v_7315 & v_7316;
assign v_7318 = v_7315 & ~v_7316;
assign v_7321 = v_13173 & v_13174;
assign v_7324 = v_7322 & v_7323;
assign v_7326 = v_7322 & ~v_7323 & v_7325;
assign v_7328 = v_7322 & ~v_7323 & ~v_7325 & v_7327;
assign v_7330 = v_7322 & ~v_7323 & ~v_7325 & ~v_7327 & ~v_7329;
assign v_7332 = v_13175 & v_13176;
assign v_7333 = v_13177 & v_13178;
assign v_7335 = v_13179 & v_13180;
assign v_7338 = v_7336 & v_7337;
assign v_7339 = v_7336 & ~v_7337;
assign v_7342 = v_7275 & v_7340 & v_7341;
assign v_7344 = v_7275 & v_7340 & ~v_7341 & v_7343;
assign v_7345 = v_7275 & v_7340 & ~v_7341 & ~v_7343;
assign v_7348 = v_7346 & v_7347;
assign v_7349 = v_7346 & ~v_7347;
assign v_7351 = v_7210 & v_7350;
assign v_7354 = v_7351;
assign v_7358 = v_7357;
assign v_7363 = ~v_7362;
assign v_7365 = v_7362 & v_7364;
assign v_7368 = v_7362 & ~v_7364 & v_7366 & v_7367;
assign v_7370 = v_7362 & ~v_7364 & v_7366 & ~v_7367 & ~v_7369;
assign v_7372 = v_7362 & ~v_7364 & ~v_7366 & ~v_7371;
assign v_7374 = v_7362 & ~v_7364 & ~v_7366 & v_7371 & v_7373;
assign v_7376 = v_13181 & v_13182;
assign v_7378 = v_13183 & v_13184;
assign v_7382 = v_13185 & v_13186;
assign v_7383 = v_13187 & v_13188;
assign v_7386 = v_7384 & v_7385;
assign v_7387 = v_7384 & ~v_7385;
assign v_7389 = v_13189 & v_13190;
assign v_7391 = ~v_7357 & ~v_7359 & v_7390;
assign v_7393 = ~v_7357 & v_7359 & ~v_7392;
assign v_7395 = ~v_7357 & v_7359 & v_7392 & ~v_7394;
assign v_7396 = ~v_7357 & v_7359 & v_7392 & v_7394;
assign v_7399 = v_7397 & v_7398;
assign v_7400 = v_7397 & ~v_7398;
assign v_7402 = v_7354 & v_7401;
assign v_7405 = v_6869 & v_7402;
assign v_7406 = ~v_6869 & v_7354 & v_7401;
assign v_7410 = v_7408 & v_7409;
assign v_7411 = v_7408 & ~v_7409;
assign v_7414 = v_7412 & v_7413;
assign v_7418 = v_7412 & ~v_7413 & ~v_7417;
assign v_7419 = v_7412 & ~v_7413 & v_7417;
assign v_7423 = v_7420;
assign v_7426 = v_7424 & v_7425;
assign v_7428 = v_7424 & ~v_7425 & v_7427;
assign v_7432 = v_7424 & ~v_7425 & ~v_7427 & v_7431;
assign v_7433 = v_7424 & ~v_7425 & ~v_7427 & ~v_7431;
assign v_7436 = v_7434 & v_7435;
assign v_7438 = v_7434 & ~v_7435 & v_7437;
assign v_7441 = v_7439 & v_7440;
assign v_7442 = v_7439 & ~v_7440;
assign v_7445 = v_7434 & ~v_7435 & ~v_7437 & v_7443 & v_7444;
assign v_7446 = v_7434 & ~v_7435 & ~v_7437 & v_7443 & ~v_7444;
assign v_7448 = v_7407 & v_7447;
assign v_7451 = ~v_7449 & v_7450;
assign v_7453 = ~v_7449 & ~v_7450 & v_7452;
assign v_7456 = v_7454 & v_7455;
assign v_7458 = v_7454 & ~v_7455 & v_7457;
assign v_7461 = v_7459 & ~v_7460;
assign v_7462 = v_7454 & ~v_7455 & ~v_7457;
assign v_7463 = v_7459 & v_7460;
assign v_7465 = v_7448 & v_7464;
assign v_7468 = v_7466 & v_7467;
assign v_7469 = v_7466 & ~v_7467;
assign v_7472 = v_7470 & v_7471;
assign v_7476 = v_7470 & ~v_7471 & ~v_7475;
assign v_7477 = v_7470 & ~v_7471 & v_7475;
assign v_7481 = v_7478;
assign v_7484 = v_7482 & v_7483;
assign v_7486 = v_7482 & ~v_7483 & v_7485;
assign v_7490 = v_7482 & ~v_7483 & ~v_7485 & v_7489;
assign v_7491 = v_7482 & ~v_7483 & ~v_7485 & ~v_7489;
assign v_7494 = v_7492 & v_7493;
assign v_7496 = v_7492 & ~v_7493 & v_7495;
assign v_7499 = v_7497 & v_7498;
assign v_7500 = v_7497 & ~v_7498;
assign v_7503 = v_7492 & ~v_7493 & ~v_7495 & v_7501 & v_7502;
assign v_7504 = v_7492 & ~v_7493 & ~v_7495 & v_7501 & ~v_7502;
assign v_7506 = v_6868 & v_7465 & v_7505;
assign v_7508 = v_7507 & v_7407 & v_7447;
assign v_7510 = v_7509 & v_7402;
assign v_7512 = v_7511 & v_7402;
assign v_7514 = v_7513 & v_7354 & v_7401;
assign v_7516 = v_7515 & v_7354 & v_7401;
assign v_7517 = ~v_7515 & v_7351;
assign v_7519 = ~v_7513 & v_7518;
assign v_7521 = ~v_7511 & v_7520;
assign v_7523 = ~v_7509 & v_7522;
assign v_7525 = ~v_7507 & v_7524;
assign v_7527 = ~v_6868 & v_7526;
assign v_7531 = v_7528;
assign v_7534 = v_7531;
assign v_7537 = v_7535 & ~v_7536;
assign v_7539 = v_7535 & v_7536 & ~v_7538;
assign v_7542 = v_7535 & v_7536 & v_7538 & ~v_7540 & ~v_7541;
assign v_7543 = v_7535 & v_7536 & v_7538 & v_7540;
assign v_7544 = v_7535 & v_7536 & v_7538 & ~v_7540 & v_7541;
assign v_7547 = v_7545 & v_7546;
assign v_7549 = v_7545 & ~v_7546 & v_7548;
assign v_7552 = ~v_7550 & v_7551;
assign v_7554 = ~v_7550 & ~v_7551 & v_7553;
assign v_7557 = v_7555 & v_7556;
assign v_7559 = v_7555 & ~v_7556 & v_7558;
assign v_7562 = v_7560 & ~v_7561;
assign v_7563 = v_7555 & ~v_7556 & ~v_7558;
assign v_7564 = v_7560 & v_7561;
assign v_7567 = v_7545 & ~v_7546 & ~v_7548 & v_7565 & v_7566;
assign v_7568 = v_7545 & ~v_7546 & ~v_7548 & v_7565 & ~v_7566;
assign v_7570 = v_7534 & v_7569;
assign v_7574 = v_7572 & v_7573;
assign v_7575 = v_7572 & ~v_7573;
assign v_7578 = v_7576 & v_7577;
assign v_7582 = v_7576 & ~v_7577 & ~v_7581;
assign v_7583 = v_7576 & ~v_7577 & v_7581;
assign v_7587 = v_7584;
assign v_7591 = v_7571 & v_7588 & v_7589 & ~v_7590;
assign v_7596 = v_13191 & v_13192;
assign v_7598 = v_13193 & v_13194;
assign v_7600 = v_13195 & v_13196;
assign v_7602 = v_13197 & v_13198;
assign v_7606 = v_7603 & ~v_7604 & v_7605;
assign v_7607 = v_7603 & ~v_7604 & ~v_7605;
assign v_7609 = v_7603 & v_7604 & v_7608;
assign v_7610 = v_7603 & v_7604 & ~v_7608;
assign v_7614 = v_7612 & v_7613;
assign v_7615 = v_7612 & ~v_7613;
assign v_7618 = v_7616 & v_7617;
assign v_7623 = v_7616 & ~v_7617;
assign v_7627 = v_7625 & v_7626;
assign v_7628 = v_7625 & ~v_7626;
assign v_7631 = v_7629 & v_7630;
assign v_7636 = v_7629 & ~v_7630;
assign v_7640 = v_7611 & v_7624 & v_7637;
assign v_7643 = v_7641 & v_7642;
assign v_7644 = v_7641 & ~v_7642;
assign v_7647 = v_7645 & v_7646;
assign v_7651 = v_7645 & ~v_7646 & ~v_7650;
assign v_7652 = v_7645 & ~v_7646 & v_7650;
assign v_7656 = v_7653;
assign v_7659 = v_7571 & v_7588 & ~v_7589 & v_7657 & v_7658;
assign v_7660 = v_7571 & v_7588 & ~v_7589 & v_7657 & ~v_7658;
assign v_7661 = v_7571 & v_7588 & v_7589 & v_7590 & v_7592;
assign v_7663 = v_7570 & v_7662;
assign v_7668 = v_7666 & v_7667;
assign v_7669 = v_7666 & ~v_7667;
assign v_7672 = v_7670 & v_7671;
assign v_7673 = v_7670 & ~v_7671;
assign v_7676 = v_7674 & ~v_7675;
assign v_7678 = v_7674 & v_7675 & v_7677;
assign v_7679 = v_7674 & v_7675 & ~v_7677;
assign v_7682 = v_7664 & v_7665 & v_7680 & v_7681;
assign v_7684 = v_7664 & ~v_7665 & v_7683;
assign v_7685 = v_7664 & v_7665 & v_7680 & ~v_7681;
assign v_7686 = v_7664 & ~v_7665 & ~v_7683;
assign v_7691 = v_7689 & v_7690;
assign v_7692 = v_7689 & ~v_7690;
assign v_7695 = v_7693 & v_7694;
assign v_7696 = v_7693 & ~v_7694;
assign v_7699 = v_7697 & ~v_7698;
assign v_7701 = v_7697 & v_7698 & v_7700;
assign v_7702 = v_7697 & v_7698 & ~v_7700;
assign v_7705 = v_7687 & v_7688 & v_7703 & v_7704;
assign v_7707 = v_7687 & ~v_7688 & v_7706;
assign v_7708 = v_7687 & v_7688 & v_7703 & ~v_7704;
assign v_7709 = v_7687 & ~v_7688 & ~v_7706;
assign v_7714 = v_7712 & v_7713;
assign v_7715 = v_7712 & ~v_7713;
assign v_7718 = v_7716 & v_7717;
assign v_7719 = v_7716 & ~v_7717;
assign v_7722 = v_7720 & ~v_7721;
assign v_7724 = v_7720 & v_7721 & v_7723;
assign v_7725 = v_7720 & v_7721 & ~v_7723;
assign v_7728 = v_7710 & v_7711 & v_7726 & v_7727;
assign v_7730 = v_7710 & ~v_7711 & v_7729;
assign v_7731 = v_7710 & v_7711 & v_7726 & ~v_7727;
assign v_7732 = v_7710 & ~v_7711 & ~v_7729;
assign v_7737 = v_7733 & v_7734 & ~v_7735 & v_7736;
assign v_7739 = v_7733 & ~v_7734 & v_7738;
assign v_7740 = v_7733 & ~v_7734 & ~v_7738;
assign v_7741 = v_7733 & v_7734 & ~v_7735 & ~v_7736;
assign v_7742 = v_7733 & v_7734 & v_7735;
assign v_7744 = v_7663 & v_7743;
assign v_7749 = v_7747 & v_7748;
assign v_7750 = v_7747 & ~v_7748;
assign v_7753 = v_7751 & v_7752;
assign v_7754 = v_7751 & ~v_7752;
assign v_7757 = v_7755 & ~v_7756;
assign v_7759 = v_7755 & v_7756 & v_7758;
assign v_7760 = v_7755 & v_7756 & ~v_7758;
assign v_7763 = v_7745 & v_7746 & v_7761 & v_7762;
assign v_7765 = v_7745 & ~v_7746 & v_7764;
assign v_7766 = v_7745 & v_7746 & v_7761 & ~v_7762;
assign v_7767 = v_7745 & ~v_7746 & ~v_7764;
assign v_7772 = v_7770 & v_7771;
assign v_7773 = v_7770 & ~v_7771;
assign v_7776 = v_7774 & v_7775;
assign v_7777 = v_7774 & ~v_7775;
assign v_7780 = v_7778 & ~v_7779;
assign v_7782 = v_7778 & v_7779 & v_7781;
assign v_7783 = v_7778 & v_7779 & ~v_7781;
assign v_7786 = v_7768 & v_7769 & v_7784 & v_7785;
assign v_7788 = v_7768 & ~v_7769 & v_7787;
assign v_7789 = v_7768 & v_7769 & v_7784 & ~v_7785;
assign v_7790 = v_7768 & ~v_7769 & ~v_7787;
assign v_7795 = v_7793 & v_7794;
assign v_7796 = v_7793 & ~v_7794;
assign v_7799 = v_7797 & v_7798;
assign v_7800 = v_7797 & ~v_7798;
assign v_7803 = v_7801 & ~v_7802;
assign v_7805 = v_7801 & v_7802 & v_7804;
assign v_7806 = v_7801 & v_7802 & ~v_7804;
assign v_7809 = v_7791 & v_7792 & v_7807 & v_7808;
assign v_7811 = v_7791 & ~v_7792 & v_7810;
assign v_7812 = v_7791 & v_7792 & v_7807 & ~v_7808;
assign v_7813 = v_7791 & ~v_7792 & ~v_7810;
assign v_7818 = v_7814 & v_7815 & ~v_7816 & v_7817;
assign v_7820 = v_7814 & ~v_7815 & v_7819;
assign v_7821 = v_7814 & ~v_7815 & ~v_7819;
assign v_7822 = v_7814 & v_7815 & ~v_7816 & ~v_7817;
assign v_7823 = v_7814 & v_7815 & v_7816;
assign v_7825 = v_7744 & v_7824;
assign v_7830 = v_7828 & v_7829;
assign v_7831 = v_7828 & ~v_7829;
assign v_7834 = v_7832 & v_7833;
assign v_7835 = v_7832 & ~v_7833;
assign v_7838 = v_7836 & ~v_7837;
assign v_7840 = v_7836 & v_7837 & v_7839;
assign v_7841 = v_7836 & v_7837 & ~v_7839;
assign v_7844 = v_7826 & v_7827 & v_7842 & v_7843;
assign v_7846 = v_7826 & ~v_7827 & v_7845;
assign v_7847 = v_7826 & v_7827 & v_7842 & ~v_7843;
assign v_7848 = v_7826 & ~v_7827 & ~v_7845;
assign v_7853 = v_7851 & v_7852;
assign v_7854 = v_7851 & ~v_7852;
assign v_7857 = v_7855 & v_7856;
assign v_7858 = v_7855 & ~v_7856;
assign v_7861 = v_7859 & ~v_7860;
assign v_7863 = v_7859 & v_7860 & v_7862;
assign v_7864 = v_7859 & v_7860 & ~v_7862;
assign v_7867 = v_7849 & v_7850 & v_7865 & v_7866;
assign v_7869 = v_7849 & ~v_7850 & v_7868;
assign v_7870 = v_7849 & v_7850 & v_7865 & ~v_7866;
assign v_7871 = v_7849 & ~v_7850 & ~v_7868;
assign v_7876 = v_7874 & v_7875;
assign v_7877 = v_7874 & ~v_7875;
assign v_7880 = v_7878 & v_7879;
assign v_7881 = v_7878 & ~v_7879;
assign v_7884 = v_7882 & ~v_7883;
assign v_7886 = v_7882 & v_7883 & v_7885;
assign v_7887 = v_7882 & v_7883 & ~v_7885;
assign v_7890 = v_7872 & v_7873 & v_7888 & v_7889;
assign v_7892 = v_7872 & ~v_7873 & v_7891;
assign v_7893 = v_7872 & v_7873 & v_7888 & ~v_7889;
assign v_7894 = v_7872 & ~v_7873 & ~v_7891;
assign v_7899 = v_7895 & v_7896 & ~v_7897 & v_7898;
assign v_7901 = v_7895 & ~v_7896 & v_7900;
assign v_7902 = v_7895 & ~v_7896 & ~v_7900;
assign v_7903 = v_7895 & v_7896 & ~v_7897 & ~v_7898;
assign v_7904 = v_7895 & v_7896 & v_7897;
assign v_7906 = v_7825 & v_7905;
assign v_7911 = v_7909 & v_7910;
assign v_7912 = v_7909 & ~v_7910;
assign v_7915 = v_7913 & v_7914;
assign v_7916 = v_7913 & ~v_7914;
assign v_7919 = v_7917 & ~v_7918;
assign v_7921 = v_7917 & v_7918 & v_7920;
assign v_7922 = v_7917 & v_7918 & ~v_7920;
assign v_7925 = v_7907 & v_7908 & v_7923 & v_7924;
assign v_7927 = v_7907 & ~v_7908 & v_7926;
assign v_7928 = v_7907 & v_7908 & v_7923 & ~v_7924;
assign v_7929 = v_7907 & ~v_7908 & ~v_7926;
assign v_7934 = v_7932 & v_7933;
assign v_7935 = v_7932 & ~v_7933;
assign v_7938 = v_7936 & v_7937;
assign v_7939 = v_7936 & ~v_7937;
assign v_7942 = v_7940 & ~v_7941;
assign v_7944 = v_7940 & v_7941 & v_7943;
assign v_7945 = v_7940 & v_7941 & ~v_7943;
assign v_7948 = v_7930 & v_7931 & v_7946 & v_7947;
assign v_7950 = v_7930 & ~v_7931 & v_7949;
assign v_7951 = v_7930 & v_7931 & v_7946 & ~v_7947;
assign v_7952 = v_7930 & ~v_7931 & ~v_7949;
assign v_7957 = v_7955 & v_7956;
assign v_7958 = v_7955 & ~v_7956;
assign v_7961 = v_7959 & v_7960;
assign v_7962 = v_7959 & ~v_7960;
assign v_7965 = v_7963 & ~v_7964;
assign v_7967 = v_7963 & v_7964 & v_7966;
assign v_7968 = v_7963 & v_7964 & ~v_7966;
assign v_7971 = v_7953 & v_7954 & v_7969 & v_7970;
assign v_7973 = v_7953 & ~v_7954 & v_7972;
assign v_7974 = v_7953 & v_7954 & v_7969 & ~v_7970;
assign v_7975 = v_7953 & ~v_7954 & ~v_7972;
assign v_7980 = v_7976 & v_7977 & ~v_7978 & v_7979;
assign v_7982 = v_7976 & ~v_7977 & v_7981;
assign v_7983 = v_7976 & ~v_7977 & ~v_7981;
assign v_7984 = v_7976 & v_7977 & ~v_7978 & ~v_7979;
assign v_7985 = v_7976 & v_7977 & v_7978;
assign v_7987 = v_7906 & v_7986;
assign v_7992 = v_7990 & v_7991;
assign v_7993 = v_7990 & ~v_7991;
assign v_7996 = v_7994 & v_7995;
assign v_7997 = v_7994 & ~v_7995;
assign v_8000 = v_7998 & ~v_7999;
assign v_8002 = v_7998 & v_7999 & v_8001;
assign v_8003 = v_7998 & v_7999 & ~v_8001;
assign v_8006 = v_7988 & v_7989 & v_8004 & v_8005;
assign v_8008 = v_7988 & ~v_7989 & v_8007;
assign v_8009 = v_7988 & v_7989 & v_8004 & ~v_8005;
assign v_8010 = v_7988 & ~v_7989 & ~v_8007;
assign v_8015 = v_8013 & v_8014;
assign v_8016 = v_8013 & ~v_8014;
assign v_8019 = v_8017 & v_8018;
assign v_8020 = v_8017 & ~v_8018;
assign v_8023 = v_8021 & ~v_8022;
assign v_8025 = v_8021 & v_8022 & v_8024;
assign v_8026 = v_8021 & v_8022 & ~v_8024;
assign v_8029 = v_8011 & v_8012 & v_8027 & v_8028;
assign v_8031 = v_8011 & ~v_8012 & v_8030;
assign v_8032 = v_8011 & v_8012 & v_8027 & ~v_8028;
assign v_8033 = v_8011 & ~v_8012 & ~v_8030;
assign v_8038 = v_8036 & v_8037;
assign v_8039 = v_8036 & ~v_8037;
assign v_8042 = v_8040 & v_8041;
assign v_8043 = v_8040 & ~v_8041;
assign v_8046 = v_8044 & ~v_8045;
assign v_8048 = v_8044 & v_8045 & v_8047;
assign v_8049 = v_8044 & v_8045 & ~v_8047;
assign v_8052 = v_8034 & v_8035 & v_8050 & v_8051;
assign v_8054 = v_8034 & ~v_8035 & v_8053;
assign v_8055 = v_8034 & v_8035 & v_8050 & ~v_8051;
assign v_8056 = v_8034 & ~v_8035 & ~v_8053;
assign v_8061 = v_8057 & v_8058 & ~v_8059 & v_8060;
assign v_8063 = v_8057 & ~v_8058 & v_8062;
assign v_8064 = v_8057 & ~v_8058 & ~v_8062;
assign v_8065 = v_8057 & v_8058 & ~v_8059 & ~v_8060;
assign v_8066 = v_8057 & v_8058 & v_8059;
assign v_8068 = v_7987 & v_8067;
assign v_8073 = v_8071 & v_8072;
assign v_8074 = v_8071 & ~v_8072;
assign v_8077 = v_8075 & v_8076;
assign v_8078 = v_8075 & ~v_8076;
assign v_8081 = v_8079 & ~v_8080;
assign v_8083 = v_8079 & v_8080 & v_8082;
assign v_8084 = v_8079 & v_8080 & ~v_8082;
assign v_8087 = v_8069 & v_8070 & v_8085 & v_8086;
assign v_8089 = v_8069 & ~v_8070 & v_8088;
assign v_8090 = v_8069 & v_8070 & v_8085 & ~v_8086;
assign v_8091 = v_8069 & ~v_8070 & ~v_8088;
assign v_8096 = v_8094 & v_8095;
assign v_8097 = v_8094 & ~v_8095;
assign v_8100 = v_8098 & v_8099;
assign v_8101 = v_8098 & ~v_8099;
assign v_8104 = v_8102 & ~v_8103;
assign v_8106 = v_8102 & v_8103 & v_8105;
assign v_8107 = v_8102 & v_8103 & ~v_8105;
assign v_8110 = v_8092 & v_8093 & v_8108 & v_8109;
assign v_8112 = v_8092 & ~v_8093 & v_8111;
assign v_8113 = v_8092 & v_8093 & v_8108 & ~v_8109;
assign v_8114 = v_8092 & ~v_8093 & ~v_8111;
assign v_8119 = v_8117 & v_8118;
assign v_8120 = v_8117 & ~v_8118;
assign v_8123 = v_8121 & v_8122;
assign v_8124 = v_8121 & ~v_8122;
assign v_8127 = v_8125 & ~v_8126;
assign v_8129 = v_8125 & v_8126 & v_8128;
assign v_8130 = v_8125 & v_8126 & ~v_8128;
assign v_8133 = v_8115 & v_8116 & v_8131 & v_8132;
assign v_8135 = v_8115 & ~v_8116 & v_8134;
assign v_8136 = v_8115 & v_8116 & v_8131 & ~v_8132;
assign v_8137 = v_8115 & ~v_8116 & ~v_8134;
assign v_8142 = v_8138 & v_8139 & ~v_8140 & v_8141;
assign v_8144 = v_8138 & ~v_8139 & v_8143;
assign v_8145 = v_8138 & ~v_8139 & ~v_8143;
assign v_8146 = v_8138 & v_8139 & ~v_8140 & ~v_8141;
assign v_8147 = v_8138 & v_8139 & v_8140;
assign v_8149 = v_8068 & v_8148;
assign v_8154 = v_8152 & v_8153;
assign v_8155 = v_8152 & ~v_8153;
assign v_8158 = v_8156 & v_8157;
assign v_8159 = v_8156 & ~v_8157;
assign v_8162 = v_8160 & ~v_8161;
assign v_8164 = v_8160 & v_8161 & v_8163;
assign v_8165 = v_8160 & v_8161 & ~v_8163;
assign v_8168 = v_8150 & v_8151 & v_8166 & v_8167;
assign v_8170 = v_8150 & ~v_8151 & v_8169;
assign v_8171 = v_8150 & v_8151 & v_8166 & ~v_8167;
assign v_8172 = v_8150 & ~v_8151 & ~v_8169;
assign v_8177 = v_8175 & v_8176;
assign v_8178 = v_8175 & ~v_8176;
assign v_8181 = v_8179 & v_8180;
assign v_8182 = v_8179 & ~v_8180;
assign v_8185 = v_8183 & ~v_8184;
assign v_8187 = v_8183 & v_8184 & v_8186;
assign v_8188 = v_8183 & v_8184 & ~v_8186;
assign v_8191 = v_8173 & v_8174 & v_8189 & v_8190;
assign v_8193 = v_8173 & ~v_8174 & v_8192;
assign v_8194 = v_8173 & v_8174 & v_8189 & ~v_8190;
assign v_8195 = v_8173 & ~v_8174 & ~v_8192;
assign v_8200 = v_8198 & v_8199;
assign v_8201 = v_8198 & ~v_8199;
assign v_8204 = v_8202 & v_8203;
assign v_8205 = v_8202 & ~v_8203;
assign v_8208 = v_8206 & ~v_8207;
assign v_8210 = v_8206 & v_8207 & v_8209;
assign v_8211 = v_8206 & v_8207 & ~v_8209;
assign v_8214 = v_8196 & v_8197 & v_8212 & v_8213;
assign v_8216 = v_8196 & ~v_8197 & v_8215;
assign v_8217 = v_8196 & v_8197 & v_8212 & ~v_8213;
assign v_8218 = v_8196 & ~v_8197 & ~v_8215;
assign v_8223 = v_8219 & v_8220 & ~v_8221 & v_8222;
assign v_8225 = v_8219 & ~v_8220 & v_8224;
assign v_8226 = v_8219 & ~v_8220 & ~v_8224;
assign v_8227 = v_8219 & v_8220 & ~v_8221 & ~v_8222;
assign v_8228 = v_8219 & v_8220 & v_8221;
assign v_8230 = v_8149 & v_8229;
assign v_8234 = v_8232 & ~v_8233;
assign v_8236 = v_8231 & v_8235;
assign v_8238 = ~v_7093 & v_7095 & v_7128 & ~v_7130;
assign v_8239 = ~v_7093 & v_7095 & v_7128 & v_7130;
assign v_8240 = ~v_7093 & v_7095 & ~v_7128;
assign v_8243 = v_8242;
assign v_8245 = v_8244;
assign v_8246 = v_13199 & v_13200;
assign v_8248 = v_8247 & ~v_7093 & ~v_7095 & v_7126;
assign v_8250 = v_8237 & ~v_8249;
assign v_8252 = v_8251 & v_7133 & v_7134;
assign v_8253 = v_8251 & v_7133 & ~v_7134;
assign v_8255 = v_8254 & ~v_7145;
assign v_8257 = v_8254 & v_8256;
assign v_8258 = v_8254 & v_7145 & v_7157 & ~v_7158 & v_7166;
assign v_8261 = v_8259 & v_8260;
assign v_8262 = v_8259 & v_7187 & v_7188;
assign v_8263 = v_8259 & v_7187 & ~v_7188 & v_7190;
assign v_8264 = v_8259 & v_7187 & ~v_7188 & ~v_7190 & v_7192;
assign v_8265 = v_8259 & v_7187 & ~v_7188 & ~v_7190 & ~v_7192;
assign v_8268 = v_8266 & v_8267;
assign v_8270 = v_8269 & ~v_7174 & v_7175 & v_7195;
assign v_8273 = v_8271 & v_8272;
assign v_8275 = v_8271 & v_8274;
assign v_8277 = ~v_8231 & v_8276;
assign v_8279 = v_8278 & v_7211 & v_7212;
assign v_8280 = v_8278 & v_7211 & ~v_7212 & v_7214;
assign v_8281 = v_8278 & v_7211 & ~v_7212 & ~v_7214 & v_7216;
assign v_8282 = v_8278 & v_7222 & v_7223;
assign v_8283 = v_8278 & v_7225 & v_7226;
assign v_8284 = v_8278 & v_7225 & ~v_7226 & v_7228;
assign v_8285 = v_8278 & v_7225 & ~v_7226 & ~v_7228 & v_7230;
assign v_8287 = v_8278 & v_8286;
assign v_8290 = v_8288 & v_8289;
assign v_8292 = v_8291 & v_7222 & ~v_7223 & v_7235 & v_7236;
assign v_8293 = v_8291 & v_7238 & v_7239;
assign v_8294 = v_8291 & v_7238 & ~v_7239 & v_7241;
assign v_8295 = v_8291 & v_7238 & ~v_7239 & ~v_7241 & v_7243;
assign v_8297 = v_8291 & v_8296;
assign v_8298 = v_13201 & v_13202;
assign v_8300 = v_8299 & v_7250 & v_7251;
assign v_8301 = v_8299 & v_7250 & ~v_7251;
assign v_8304 = v_8302 & v_8303;
assign v_8306 = v_13203 & v_13204;
assign v_8307 = v_8305 & v_7257 & v_7258;
assign v_8308 = v_8305 & v_7257 & ~v_7258 & v_7260;
assign v_8309 = v_8305 & v_7257 & ~v_7258 & ~v_7260 & v_7262;
assign v_8311 = v_8305 & v_8310;
assign v_8313 = v_13205 & v_13206;
assign v_8316 = v_8314 & v_8315;
assign v_8318 = v_8317 & v_7276 & v_7277;
assign v_8319 = v_8317 & v_7276 & ~v_7277 & v_7279;
assign v_8320 = v_8317 & v_7276 & ~v_7277 & ~v_7279 & v_7281;
assign v_8321 = v_8317 & v_7287 & v_7288;
assign v_8322 = v_8317 & v_7290 & v_7291;
assign v_8323 = v_8317 & v_7290 & ~v_7291 & v_7293;
assign v_8324 = v_8317 & v_7290 & ~v_7291 & ~v_7293 & v_7295;
assign v_8326 = v_8317 & v_8325;
assign v_8329 = v_8327 & v_8328;
assign v_8331 = v_8330 & v_7287 & ~v_7288 & v_7300 & v_7301;
assign v_8332 = v_8330 & v_7303 & v_7304;
assign v_8333 = v_8330 & v_7303 & ~v_7304 & v_7306;
assign v_8334 = v_8330 & v_7303 & ~v_7304 & ~v_7306 & v_7308;
assign v_8336 = v_8330 & v_8335;
assign v_8337 = v_13207 & v_13208;
assign v_8339 = v_8338 & v_7315 & v_7316;
assign v_8340 = v_8338 & v_7315 & ~v_7316;
assign v_8343 = v_8341 & v_8342;
assign v_8345 = v_13209 & v_13210;
assign v_8346 = v_8344 & v_7322 & v_7323;
assign v_8347 = v_8344 & v_7322 & ~v_7323 & v_7325;
assign v_8348 = v_8344 & v_7322 & ~v_7323 & ~v_7325 & v_7327;
assign v_8350 = v_8344 & v_8349;
assign v_8352 = v_13211 & v_13212;
assign v_8355 = v_8353 & v_8354;
assign v_8357 = v_8356 & v_7357;
assign v_8360 = v_8359 & ~v_8356;
assign v_8362 = v_8361 & ~v_7357 & v_7359 & v_7392 & ~v_7394;
assign v_8363 = v_8361 & ~v_7357 & v_7359 & v_7392 & v_7394;
assign v_8364 = v_8361 & ~v_7357 & v_7359 & ~v_7392;
assign v_8365 = v_8361 & v_7360;
assign v_8366 = v_8361 & ~v_7360;
assign v_8369 = v_8367 & v_8368;
assign v_8371 = v_8367 & v_8370;
assign v_8372 = v_13213 & v_13214;
assign v_8374 = v_8373 & ~v_7357 & ~v_7359 & v_7390;
assign v_8376 = v_8358 & ~v_8375;
assign v_8378 = v_8377 & v_7397 & v_7398;
assign v_8379 = v_8377 & v_7397 & ~v_7398;
assign v_8381 = v_8380 & v_7412 & v_7413;
assign v_8382 = v_8380 & v_7420;
assign v_8384 = v_8383 & v_7424 & v_7425;
assign v_8385 = v_8383 & v_7424 & ~v_7425 & v_7427;
assign v_8387 = v_8383 & v_8386;
assign v_8390 = v_8388 & v_8389;
assign v_8392 = v_8388 & v_8391;
assign v_8394 = v_8393 & v_7454 & ~v_7455 & ~v_7457;
assign v_8395 = v_8393 & v_7459 & ~v_7460;
assign v_8396 = v_8393 & v_7459 & v_7460;
assign v_8397 = v_8393 & v_7449;
assign v_8399 = v_8398 & v_7470 & v_7471;
assign v_8400 = v_8398 & v_7478;
assign v_8402 = v_8401 & v_7482 & v_7483;
assign v_8403 = v_8401 & v_7482 & ~v_7483 & v_7485;
assign v_8405 = v_8401 & v_8404;
assign v_8408 = v_8406 & v_8407;
assign v_8410 = v_8406 & v_8409;
assign v_8412 = v_6868 & v_8411;
assign v_8413 = v_7507 & v_8393;
assign v_8414 = v_7509 & v_8380;
assign v_8415 = v_7511 & v_8380;
assign v_8416 = v_7513 & v_8380;
assign v_8417 = v_7515 & v_8380;
assign v_8418 = ~v_7515 & v_8356;
assign v_8420 = ~v_7513 & v_8419;
assign v_8422 = ~v_7511 & v_8421;
assign v_8424 = ~v_7509 & v_8423;
assign v_8426 = ~v_7507 & v_8425;
assign v_8428 = ~v_6868 & v_8427;
assign v_8430 = v_8429 & ~v_7535;
assign v_8431 = v_13215 & v_13216;
assign v_8432 = v_8429 & v_7535 & v_7536 & v_7538 & v_7540;
assign v_8433 = v_13217 & v_13218;
assign v_8435 = v_8434 & v_7545 & ~v_7546 & v_7548;
assign v_8436 = v_8434 & v_7555 & ~v_7556 & ~v_7558;
assign v_8437 = v_8434 & v_7560 & ~v_7561;
assign v_8438 = v_8434 & v_7560 & v_7561;
assign v_8439 = v_8434 & v_7550;
assign v_8442 = v_8440 & v_8441;
assign v_8445 = v_8443 & v_8444;
assign v_8446 = v_8434 & v_7545 & v_7546;
assign v_8448 = v_8429 & v_8447;
assign v_8450 = v_8449 & ~v_7571;
assign v_8451 = v_8449 & v_7576 & v_7577;
assign v_8452 = v_8449 & v_7584;
assign v_8454 = v_8453 & v_7571 & v_7588 & v_7589 & ~v_7590;
assign v_8456 = v_8453 & v_8455;
assign v_8457 = v_8453 & v_7616 & v_7617;
assign v_8458 = v_8453 & v_7616 & ~v_7617;
assign v_8460 = v_8459 & v_7629 & v_7630;
assign v_8461 = v_8459 & v_7629 & ~v_7630;
assign v_8463 = v_8462 & v_7611 & v_7624 & v_7637;
assign v_8464 = v_13219 & v_13220;
assign v_8465 = v_8453 & v_7645 & v_7646;
assign v_8466 = v_8453 & v_7653;
assign v_8469 = v_8467 & v_8468;
assign v_8471 = v_8470 & v_7664 & ~v_7665 & v_7683;
assign v_8472 = v_8470 & v_7664 & ~v_7665 & ~v_7683;
assign v_8473 = v_8470 & ~v_7666;
assign v_8474 = v_8470 & v_7674 & ~v_7675;
assign v_8476 = v_8470 & v_8475;
assign v_8478 = v_8477 & v_7664 & v_7665 & v_7680 & ~v_7681;
assign v_8480 = v_8479 & v_7687 & ~v_7688 & v_7706;
assign v_8481 = v_8479 & v_7687 & ~v_7688 & ~v_7706;
assign v_8482 = v_8479 & ~v_7689;
assign v_8483 = v_8479 & v_7697 & ~v_7698;
assign v_8485 = v_8479 & v_8484;
assign v_8487 = v_8486 & v_7687 & v_7688 & v_7703 & ~v_7704;
assign v_8489 = v_8488 & v_7710 & ~v_7711 & v_7729;
assign v_8490 = v_8488 & ~v_7712;
assign v_8491 = v_8488 & v_7720 & ~v_7721;
assign v_8493 = v_8488 & v_8492;
assign v_8495 = v_8494 & v_7710 & v_7711 & v_7726 & v_7727;
assign v_8496 = v_8488 & v_7710 & ~v_7711 & ~v_7729;
assign v_8497 = v_8494 & v_7710 & v_7711 & v_7726 & ~v_7727;
assign v_8500 = v_8498 & v_8499;
assign v_8501 = v_8498 & v_7733 & v_7734 & ~v_7735 & ~v_7736;
assign v_8502 = v_8498 & v_7733 & v_7734 & v_7735;
assign v_8503 = v_8498 & v_7733 & ~v_7734 & ~v_7738;
assign v_8506 = v_8504 & v_8505;
assign v_8507 = v_8486 & v_7687 & v_7688 & v_7703 & v_7704;
assign v_8508 = v_8477 & v_7664 & v_7665 & v_7680 & v_7681;
assign v_8510 = v_8509 & v_7745 & ~v_7746 & v_7764;
assign v_8511 = v_8509 & v_7745 & ~v_7746 & ~v_7764;
assign v_8512 = v_8509 & ~v_7747;
assign v_8513 = v_8509 & v_7755 & ~v_7756;
assign v_8515 = v_8509 & v_8514;
assign v_8517 = v_8516 & v_7745 & v_7746 & v_7761 & ~v_7762;
assign v_8519 = v_8518 & v_7768 & ~v_7769 & v_7787;
assign v_8520 = v_8518 & v_7768 & ~v_7769 & ~v_7787;
assign v_8521 = v_8518 & ~v_7770;
assign v_8522 = v_8518 & v_7778 & ~v_7779;
assign v_8524 = v_8518 & v_8523;
assign v_8526 = v_8525 & v_7768 & v_7769 & v_7784 & ~v_7785;
assign v_8528 = v_8527 & v_7791 & ~v_7792 & v_7810;
assign v_8529 = v_8527 & ~v_7793;
assign v_8530 = v_8527 & v_7801 & ~v_7802;
assign v_8532 = v_8527 & v_8531;
assign v_8534 = v_8533 & v_7791 & v_7792 & v_7807 & v_7808;
assign v_8535 = v_8527 & v_7791 & ~v_7792 & ~v_7810;
assign v_8536 = v_8533 & v_7791 & v_7792 & v_7807 & ~v_7808;
assign v_8539 = v_8537 & v_8538;
assign v_8540 = v_8537 & v_7814 & v_7815 & ~v_7816 & ~v_7817;
assign v_8541 = v_8537 & v_7814 & v_7815 & v_7816;
assign v_8542 = v_8537 & v_7814 & ~v_7815 & ~v_7819;
assign v_8545 = v_8543 & v_8544;
assign v_8546 = v_8525 & v_7768 & v_7769 & v_7784 & v_7785;
assign v_8547 = v_8516 & v_7745 & v_7746 & v_7761 & v_7762;
assign v_8549 = v_8548 & v_7826 & ~v_7827 & v_7845;
assign v_8550 = v_8548 & v_7826 & ~v_7827 & ~v_7845;
assign v_8551 = v_8548 & ~v_7828;
assign v_8552 = v_8548 & v_7836 & ~v_7837;
assign v_8554 = v_8548 & v_8553;
assign v_8556 = v_8555 & v_7826 & v_7827 & v_7842 & ~v_7843;
assign v_8558 = v_8557 & v_7849 & ~v_7850 & v_7868;
assign v_8559 = v_8557 & v_7849 & ~v_7850 & ~v_7868;
assign v_8560 = v_8557 & ~v_7851;
assign v_8561 = v_8557 & v_7859 & ~v_7860;
assign v_8563 = v_8557 & v_8562;
assign v_8565 = v_8564 & v_7849 & v_7850 & v_7865 & ~v_7866;
assign v_8567 = v_8566 & v_7872 & ~v_7873 & v_7891;
assign v_8568 = v_8566 & ~v_7874;
assign v_8569 = v_8566 & v_7882 & ~v_7883;
assign v_8571 = v_8566 & v_8570;
assign v_8573 = v_8572 & v_7872 & v_7873 & v_7888 & v_7889;
assign v_8574 = v_8566 & v_7872 & ~v_7873 & ~v_7891;
assign v_8575 = v_8572 & v_7872 & v_7873 & v_7888 & ~v_7889;
assign v_8578 = v_8576 & v_8577;
assign v_8579 = v_8576 & v_7895 & v_7896 & ~v_7897 & ~v_7898;
assign v_8580 = v_8576 & v_7895 & v_7896 & v_7897;
assign v_8581 = v_8576 & v_7895 & ~v_7896 & ~v_7900;
assign v_8584 = v_8582 & v_8583;
assign v_8585 = v_8564 & v_7849 & v_7850 & v_7865 & v_7866;
assign v_8586 = v_8555 & v_7826 & v_7827 & v_7842 & v_7843;
assign v_8588 = v_8587 & v_7907 & ~v_7908 & v_7926;
assign v_8589 = v_8587 & v_7907 & ~v_7908 & ~v_7926;
assign v_8590 = v_8587 & ~v_7909;
assign v_8591 = v_8587 & v_7917 & ~v_7918;
assign v_8593 = v_8587 & v_8592;
assign v_8595 = v_8594 & v_7907 & v_7908 & v_7923 & ~v_7924;
assign v_8597 = v_8596 & v_7930 & ~v_7931 & v_7949;
assign v_8598 = v_8596 & v_7930 & ~v_7931 & ~v_7949;
assign v_8599 = v_8596 & ~v_7932;
assign v_8600 = v_8596 & v_7940 & ~v_7941;
assign v_8602 = v_8596 & v_8601;
assign v_8604 = v_8603 & v_7930 & v_7931 & v_7946 & ~v_7947;
assign v_8606 = v_8605 & v_7953 & ~v_7954 & v_7972;
assign v_8607 = v_8605 & ~v_7955;
assign v_8608 = v_8605 & v_7963 & ~v_7964;
assign v_8610 = v_8605 & v_8609;
assign v_8612 = v_8611 & v_7953 & v_7954 & v_7969 & v_7970;
assign v_8613 = v_8605 & v_7953 & ~v_7954 & ~v_7972;
assign v_8614 = v_8611 & v_7953 & v_7954 & v_7969 & ~v_7970;
assign v_8617 = v_8615 & v_8616;
assign v_8618 = v_8615 & v_7976 & v_7977 & ~v_7978 & ~v_7979;
assign v_8619 = v_8615 & v_7976 & v_7977 & v_7978;
assign v_8620 = v_8615 & v_7976 & ~v_7977 & ~v_7981;
assign v_8623 = v_8621 & v_8622;
assign v_8624 = v_8603 & v_7930 & v_7931 & v_7946 & v_7947;
assign v_8625 = v_8594 & v_7907 & v_7908 & v_7923 & v_7924;
assign v_8627 = v_8626 & v_7988 & ~v_7989 & v_8007;
assign v_8628 = v_8626 & v_7988 & ~v_7989 & ~v_8007;
assign v_8629 = v_8626 & ~v_7990;
assign v_8630 = v_8626 & v_7998 & ~v_7999;
assign v_8632 = v_8626 & v_8631;
assign v_8634 = v_8633 & v_7988 & v_7989 & v_8004 & ~v_8005;
assign v_8636 = v_8635 & v_8011 & ~v_8012 & v_8030;
assign v_8637 = v_8635 & v_8011 & ~v_8012 & ~v_8030;
assign v_8638 = v_8635 & ~v_8013;
assign v_8639 = v_8635 & v_8021 & ~v_8022;
assign v_8641 = v_8635 & v_8640;
assign v_8643 = v_8642 & v_8011 & v_8012 & v_8027 & ~v_8028;
assign v_8645 = v_8644 & v_8034 & ~v_8035 & v_8053;
assign v_8646 = v_8644 & ~v_8036;
assign v_8647 = v_8644 & v_8044 & ~v_8045;
assign v_8649 = v_8644 & v_8648;
assign v_8651 = v_8650 & v_8034 & v_8035 & v_8050 & v_8051;
assign v_8652 = v_8644 & v_8034 & ~v_8035 & ~v_8053;
assign v_8653 = v_8650 & v_8034 & v_8035 & v_8050 & ~v_8051;
assign v_8656 = v_8654 & v_8655;
assign v_8657 = v_8654 & v_8057 & v_8058 & ~v_8059 & ~v_8060;
assign v_8658 = v_8654 & v_8057 & v_8058 & v_8059;
assign v_8659 = v_8654 & v_8057 & ~v_8058 & ~v_8062;
assign v_8662 = v_8660 & v_8661;
assign v_8663 = v_8642 & v_8011 & v_8012 & v_8027 & v_8028;
assign v_8664 = v_8633 & v_7988 & v_7989 & v_8004 & v_8005;
assign v_8666 = v_8665 & v_8069 & ~v_8070 & v_8088;
assign v_8667 = v_8665 & v_8069 & ~v_8070 & ~v_8088;
assign v_8668 = v_8665 & ~v_8071;
assign v_8669 = v_8665 & v_8079 & ~v_8080;
assign v_8671 = v_8665 & v_8670;
assign v_8673 = v_8672 & v_8069 & v_8070 & v_8085 & ~v_8086;
assign v_8675 = v_8674 & v_8092 & ~v_8093 & v_8111;
assign v_8676 = v_8674 & v_8092 & ~v_8093 & ~v_8111;
assign v_8677 = v_8674 & ~v_8094;
assign v_8678 = v_8674 & v_8102 & ~v_8103;
assign v_8680 = v_8674 & v_8679;
assign v_8682 = v_8681 & v_8092 & v_8093 & v_8108 & ~v_8109;
assign v_8684 = v_8683 & v_8115 & ~v_8116 & v_8134;
assign v_8685 = v_8683 & ~v_8117;
assign v_8686 = v_8683 & v_8125 & ~v_8126;
assign v_8688 = v_8683 & v_8687;
assign v_8690 = v_8689 & v_8115 & v_8116 & v_8131 & v_8132;
assign v_8691 = v_8683 & v_8115 & ~v_8116 & ~v_8134;
assign v_8692 = v_8689 & v_8115 & v_8116 & v_8131 & ~v_8132;
assign v_8695 = v_8693 & v_8694;
assign v_8696 = v_8693 & v_8138 & v_8139 & ~v_8140 & ~v_8141;
assign v_8697 = v_8693 & v_8138 & v_8139 & v_8140;
assign v_8698 = v_8693 & v_8138 & ~v_8139 & ~v_8143;
assign v_8701 = v_8699 & v_8700;
assign v_8702 = v_8681 & v_8092 & v_8093 & v_8108 & v_8109;
assign v_8703 = v_8672 & v_8069 & v_8070 & v_8085 & v_8086;
assign v_8705 = v_8704 & v_8150 & ~v_8151 & v_8169;
assign v_8706 = v_8704 & v_8150 & ~v_8151 & ~v_8169;
assign v_8707 = v_8704 & ~v_8152;
assign v_8708 = v_8704 & v_8160 & ~v_8161;
assign v_8710 = v_8704 & v_8709;
assign v_8712 = v_8711 & v_8150 & v_8151 & v_8166 & ~v_8167;
assign v_8714 = v_8713 & v_8173 & ~v_8174 & v_8192;
assign v_8715 = v_8713 & v_8173 & ~v_8174 & ~v_8192;
assign v_8716 = v_8713 & ~v_8175;
assign v_8717 = v_8713 & v_8183 & ~v_8184;
assign v_8719 = v_8713 & v_8718;
assign v_8721 = v_8720 & v_8173 & v_8174 & v_8189 & ~v_8190;
assign v_8723 = v_8722 & v_8196 & ~v_8197 & v_8215;
assign v_8724 = v_8722 & ~v_8198;
assign v_8725 = v_8722 & v_8206 & ~v_8207;
assign v_8727 = v_8722 & v_8726;
assign v_8729 = v_8728 & v_8196 & v_8197 & v_8212 & v_8213;
assign v_8730 = v_8722 & v_8196 & ~v_8197 & ~v_8215;
assign v_8731 = v_8728 & v_8196 & v_8197 & v_8212 & ~v_8213;
assign v_8734 = v_8732 & v_8733;
assign v_8735 = v_8732 & v_8219 & v_8220 & ~v_8221 & ~v_8222;
assign v_8736 = v_8732 & v_8219 & v_8220 & v_8221;
assign v_8737 = v_8732 & v_8219 & ~v_8220 & ~v_8224;
assign v_8740 = v_8738 & v_8739;
assign v_8741 = v_8720 & v_8173 & v_8174 & v_8189 & v_8190;
assign v_8742 = v_8711 & v_8150 & v_8151 & v_8166 & v_8167;
assign v_8746 = v_8231 & v_8745;
assign v_8747 = v_7093;
assign v_8750 = v_8749 & v_7133 & v_7134;
assign v_8751 = v_8749 & v_7133 & ~v_7134;
assign v_8753 = v_8752 & ~v_7145;
assign v_8755 = v_8752 & v_8754;
assign v_8756 = v_8752 & v_7145 & v_7157 & ~v_7158 & v_7166;
assign v_8759 = v_8757 & v_8758;
assign v_8760 = v_8757 & v_7187 & v_7188;
assign v_8761 = v_8757 & v_7187 & ~v_7188 & v_7190;
assign v_8762 = v_8757 & v_7187 & ~v_7188 & ~v_7190 & v_7192;
assign v_8763 = v_8757 & v_7187 & ~v_7188 & ~v_7190 & ~v_7192;
assign v_8765 = v_8764 & v_8267;
assign v_8767 = v_8766 & ~v_7174 & v_7175 & v_7195;
assign v_8770 = v_8768 & v_8769;
assign v_8771 = v_8768 & v_8274;
assign v_8773 = ~v_8231 & v_8772;
assign v_8775 = v_8774 & v_7211 & v_7212;
assign v_8776 = v_8774 & v_7211 & ~v_7212 & v_7214;
assign v_8777 = v_8774 & v_7211 & ~v_7212 & ~v_7214 & v_7216;
assign v_8778 = v_8774 & v_7222 & v_7223;
assign v_8779 = v_8774 & v_7225 & v_7226;
assign v_8780 = v_8774 & v_7225 & ~v_7226 & v_7228;
assign v_8781 = v_8774 & v_7225 & ~v_7226 & ~v_7228 & v_7230;
assign v_8782 = v_8774 & v_8286;
assign v_8784 = v_8783 & v_8289;
assign v_8786 = v_8785 & v_7222 & ~v_7223 & v_7235 & v_7236;
assign v_8787 = v_8785 & v_7238 & v_7239;
assign v_8788 = v_8785 & v_7238 & ~v_7239 & v_7241;
assign v_8789 = v_8785 & v_7238 & ~v_7239 & ~v_7241 & v_7243;
assign v_8791 = v_8785 & v_8790;
assign v_8792 = v_13221 & v_13222;
assign v_8794 = v_8793 & v_7250 & v_7251;
assign v_8795 = v_8793 & v_7250 & ~v_7251;
assign v_8797 = v_8796 & v_8303;
assign v_8799 = v_13223 & v_13224;
assign v_8800 = v_8798 & v_7257 & v_7258;
assign v_8801 = v_8798 & v_7257 & ~v_7258 & v_7260;
assign v_8802 = v_8798 & v_7257 & ~v_7258 & ~v_7260 & v_7262;
assign v_8803 = v_8798 & v_8310;
assign v_8805 = v_13225 & v_13226;
assign v_8807 = v_8806 & v_8315;
assign v_8809 = v_8808 & v_7276 & v_7277;
assign v_8810 = v_8808 & v_7276 & ~v_7277 & v_7279;
assign v_8811 = v_8808 & v_7276 & ~v_7277 & ~v_7279 & v_7281;
assign v_8812 = v_8808 & v_7287 & v_7288;
assign v_8813 = v_8808 & v_7290 & v_7291;
assign v_8814 = v_8808 & v_7290 & ~v_7291 & v_7293;
assign v_8815 = v_8808 & v_7290 & ~v_7291 & ~v_7293 & v_7295;
assign v_8816 = v_8808 & v_8325;
assign v_8818 = v_8817 & v_8328;
assign v_8820 = v_8819 & v_7287 & ~v_7288 & v_7300 & v_7301;
assign v_8821 = v_8819 & v_7303 & v_7304;
assign v_8822 = v_8819 & v_7303 & ~v_7304 & v_7306;
assign v_8823 = v_8819 & v_7303 & ~v_7304 & ~v_7306 & v_7308;
assign v_8825 = v_8819 & v_8824;
assign v_8826 = v_13227 & v_13228;
assign v_8828 = v_8827 & v_7315 & v_7316;
assign v_8829 = v_8827 & v_7315 & ~v_7316;
assign v_8831 = v_8830 & v_8342;
assign v_8833 = v_13229 & v_13230;
assign v_8834 = v_8832 & v_7322 & v_7323;
assign v_8835 = v_8832 & v_7322 & ~v_7323 & v_7325;
assign v_8836 = v_8832 & v_7322 & ~v_7323 & ~v_7325 & v_7327;
assign v_8837 = v_8832 & v_8349;
assign v_8839 = v_13231 & v_13232;
assign v_8841 = v_8840 & v_8354;
assign v_8843 = v_8842 & v_7357;
assign v_8846 = v_8845 & v_7397 & v_7398;
assign v_8847 = v_8845 & v_7397 & ~v_7398;
assign v_8849 = v_8848 & v_7412 & v_7413;
assign v_8850 = v_8848 & v_7420;
assign v_8852 = v_8851 & v_7424 & v_7425;
assign v_8853 = v_8851 & v_7424 & ~v_7425 & v_7427;
assign v_8854 = v_8851 & v_8386;
assign v_8857 = v_8855 & v_8856;
assign v_8858 = v_8855 & v_8391;
assign v_8860 = v_8859 & v_7454 & ~v_7455 & ~v_7457;
assign v_8861 = v_8859 & v_7459 & ~v_7460;
assign v_8862 = v_8859 & v_7459 & v_7460;
assign v_8863 = v_8859 & v_7449;
assign v_8865 = v_8864 & v_7470 & v_7471;
assign v_8866 = v_8864 & v_7478;
assign v_8868 = v_8867 & v_7482 & v_7483;
assign v_8869 = v_8867 & v_7482 & ~v_7483 & v_7485;
assign v_8870 = v_8867 & v_8404;
assign v_8873 = v_8871 & v_8872;
assign v_8874 = v_8871 & v_8409;
assign v_8876 = v_6868 & v_8875;
assign v_8877 = v_7507 & v_8859;
assign v_8878 = v_7509 & v_8848;
assign v_8879 = v_7511 & v_8848;
assign v_8880 = v_7513 & v_8848;
assign v_8881 = v_7515 & v_8848;
assign v_8882 = ~v_7515 & v_8842;
assign v_8884 = ~v_7513 & v_8883;
assign v_8886 = ~v_7511 & v_8885;
assign v_8888 = ~v_7509 & v_8887;
assign v_8890 = ~v_7507 & v_8889;
assign v_8892 = ~v_6868 & v_8891;
assign v_8894 = v_8893 & ~v_7535;
assign v_8895 = v_13233 & v_13234;
assign v_8896 = v_8893 & v_7535 & v_7536 & v_7538 & v_7540;
assign v_8897 = v_13235 & v_13236;
assign v_8899 = v_8898 & v_7545 & ~v_7546 & v_7548;
assign v_8900 = v_8898 & v_7555 & ~v_7556 & ~v_7558;
assign v_8901 = v_8898 & v_7560 & ~v_7561;
assign v_8902 = v_8898 & v_7560 & v_7561;
assign v_8903 = v_8898 & v_7550;
assign v_8905 = v_8904 & v_8441;
assign v_8907 = v_8906 & v_8444;
assign v_8908 = v_8898 & v_7545 & v_7546;
assign v_8909 = v_8893 & v_8447;
assign v_8911 = v_8910 & ~v_7571;
assign v_8912 = v_8910 & v_7576 & v_7577;
assign v_8913 = v_8910 & v_7584;
assign v_8915 = v_8914 & v_7571 & v_7588 & v_7589 & ~v_7590;
assign v_8917 = v_8914 & v_8916;
assign v_8918 = v_8914 & v_7616 & v_7617;
assign v_8919 = v_8914 & v_7616 & ~v_7617;
assign v_8921 = v_8920 & v_7629 & v_7630;
assign v_8922 = v_8920 & v_7629 & ~v_7630;
assign v_8924 = v_8923 & v_7611 & v_7624 & v_7637;
assign v_8925 = v_13237 & v_13238;
assign v_8926 = v_8914 & v_7645 & v_7646;
assign v_8927 = v_8914 & v_7653;
assign v_8929 = v_8928 & v_8468;
assign v_8931 = v_8930 & v_7664 & ~v_7665 & v_7683;
assign v_8932 = v_8930 & v_7664 & ~v_7665 & ~v_7683;
assign v_8933 = v_8930 & ~v_7666;
assign v_8934 = v_8930 & v_7674 & ~v_7675;
assign v_8935 = v_8930 & v_8475;
assign v_8937 = v_8936 & v_7664 & v_7665 & v_7680 & ~v_7681;
assign v_8939 = v_8938 & v_7687 & ~v_7688 & v_7706;
assign v_8940 = v_8938 & v_7687 & ~v_7688 & ~v_7706;
assign v_8941 = v_8938 & ~v_7689;
assign v_8942 = v_8938 & v_7697 & ~v_7698;
assign v_8943 = v_8938 & v_8484;
assign v_8945 = v_8944 & v_7687 & v_7688 & v_7703 & ~v_7704;
assign v_8947 = v_8946 & v_7710 & ~v_7711 & v_7729;
assign v_8948 = v_8946 & ~v_7712;
assign v_8949 = v_8946 & v_7720 & ~v_7721;
assign v_8950 = v_8946 & v_8492;
assign v_8952 = v_8951 & v_7710 & v_7711 & v_7726 & v_7727;
assign v_8953 = v_8946 & v_7710 & ~v_7711 & ~v_7729;
assign v_8954 = v_8951 & v_7710 & v_7711 & v_7726 & ~v_7727;
assign v_8957 = v_8955 & v_8956;
assign v_8958 = v_8955 & v_7733 & v_7734 & ~v_7735 & ~v_7736;
assign v_8959 = v_8955 & v_7733 & v_7734 & v_7735;
assign v_8960 = v_8955 & v_7733 & ~v_7734 & ~v_7738;
assign v_8962 = v_8961 & v_8505;
assign v_8963 = v_8944 & v_7687 & v_7688 & v_7703 & v_7704;
assign v_8964 = v_8936 & v_7664 & v_7665 & v_7680 & v_7681;
assign v_8966 = v_8965 & v_7745 & ~v_7746 & v_7764;
assign v_8967 = v_8965 & v_7745 & ~v_7746 & ~v_7764;
assign v_8968 = v_8965 & ~v_7747;
assign v_8969 = v_8965 & v_7755 & ~v_7756;
assign v_8970 = v_8965 & v_8514;
assign v_8972 = v_8971 & v_7745 & v_7746 & v_7761 & ~v_7762;
assign v_8974 = v_8973 & v_7768 & ~v_7769 & v_7787;
assign v_8975 = v_8973 & v_7768 & ~v_7769 & ~v_7787;
assign v_8976 = v_8973 & ~v_7770;
assign v_8977 = v_8973 & v_7778 & ~v_7779;
assign v_8978 = v_8973 & v_8523;
assign v_8980 = v_8979 & v_7768 & v_7769 & v_7784 & ~v_7785;
assign v_8982 = v_8981 & v_7791 & ~v_7792 & v_7810;
assign v_8983 = v_8981 & ~v_7793;
assign v_8984 = v_8981 & v_7801 & ~v_7802;
assign v_8985 = v_8981 & v_8531;
assign v_8987 = v_8986 & v_7791 & v_7792 & v_7807 & v_7808;
assign v_8988 = v_8981 & v_7791 & ~v_7792 & ~v_7810;
assign v_8989 = v_8986 & v_7791 & v_7792 & v_7807 & ~v_7808;
assign v_8992 = v_8990 & v_8991;
assign v_8993 = v_8990 & v_7814 & v_7815 & ~v_7816 & ~v_7817;
assign v_8994 = v_8990 & v_7814 & v_7815 & v_7816;
assign v_8995 = v_8990 & v_7814 & ~v_7815 & ~v_7819;
assign v_8997 = v_8996 & v_8544;
assign v_8998 = v_8979 & v_7768 & v_7769 & v_7784 & v_7785;
assign v_8999 = v_8971 & v_7745 & v_7746 & v_7761 & v_7762;
assign v_9001 = v_9000 & v_7826 & ~v_7827 & v_7845;
assign v_9002 = v_9000 & v_7826 & ~v_7827 & ~v_7845;
assign v_9003 = v_9000 & ~v_7828;
assign v_9004 = v_9000 & v_7836 & ~v_7837;
assign v_9005 = v_9000 & v_8553;
assign v_9007 = v_9006 & v_7826 & v_7827 & v_7842 & ~v_7843;
assign v_9009 = v_9008 & v_7849 & ~v_7850 & v_7868;
assign v_9010 = v_9008 & v_7849 & ~v_7850 & ~v_7868;
assign v_9011 = v_9008 & ~v_7851;
assign v_9012 = v_9008 & v_7859 & ~v_7860;
assign v_9013 = v_9008 & v_8562;
assign v_9015 = v_9014 & v_7849 & v_7850 & v_7865 & ~v_7866;
assign v_9017 = v_9016 & v_7872 & ~v_7873 & v_7891;
assign v_9018 = v_9016 & ~v_7874;
assign v_9019 = v_9016 & v_7882 & ~v_7883;
assign v_9020 = v_9016 & v_8570;
assign v_9022 = v_9021 & v_7872 & v_7873 & v_7888 & v_7889;
assign v_9023 = v_9016 & v_7872 & ~v_7873 & ~v_7891;
assign v_9024 = v_9021 & v_7872 & v_7873 & v_7888 & ~v_7889;
assign v_9027 = v_9025 & v_9026;
assign v_9028 = v_9025 & v_7895 & v_7896 & ~v_7897 & ~v_7898;
assign v_9029 = v_9025 & v_7895 & v_7896 & v_7897;
assign v_9030 = v_9025 & v_7895 & ~v_7896 & ~v_7900;
assign v_9032 = v_9031 & v_8583;
assign v_9033 = v_9014 & v_7849 & v_7850 & v_7865 & v_7866;
assign v_9034 = v_9006 & v_7826 & v_7827 & v_7842 & v_7843;
assign v_9036 = v_9035 & v_7907 & ~v_7908 & v_7926;
assign v_9037 = v_9035 & v_7907 & ~v_7908 & ~v_7926;
assign v_9038 = v_9035 & ~v_7909;
assign v_9039 = v_9035 & v_7917 & ~v_7918;
assign v_9040 = v_9035 & v_8592;
assign v_9042 = v_9041 & v_7907 & v_7908 & v_7923 & ~v_7924;
assign v_9044 = v_9043 & v_7930 & ~v_7931 & v_7949;
assign v_9045 = v_9043 & v_7930 & ~v_7931 & ~v_7949;
assign v_9046 = v_9043 & ~v_7932;
assign v_9047 = v_9043 & v_7940 & ~v_7941;
assign v_9048 = v_9043 & v_8601;
assign v_9050 = v_9049 & v_7930 & v_7931 & v_7946 & ~v_7947;
assign v_9052 = v_9051 & v_7953 & ~v_7954 & v_7972;
assign v_9053 = v_9051 & ~v_7955;
assign v_9054 = v_9051 & v_7963 & ~v_7964;
assign v_9055 = v_9051 & v_8609;
assign v_9057 = v_9056 & v_7953 & v_7954 & v_7969 & v_7970;
assign v_9058 = v_9051 & v_7953 & ~v_7954 & ~v_7972;
assign v_9059 = v_9056 & v_7953 & v_7954 & v_7969 & ~v_7970;
assign v_9062 = v_9060 & v_9061;
assign v_9063 = v_9060 & v_7976 & v_7977 & ~v_7978 & ~v_7979;
assign v_9064 = v_9060 & v_7976 & v_7977 & v_7978;
assign v_9065 = v_9060 & v_7976 & ~v_7977 & ~v_7981;
assign v_9067 = v_9066 & v_8622;
assign v_9068 = v_9049 & v_7930 & v_7931 & v_7946 & v_7947;
assign v_9069 = v_9041 & v_7907 & v_7908 & v_7923 & v_7924;
assign v_9071 = v_9070 & v_7988 & ~v_7989 & v_8007;
assign v_9072 = v_9070 & v_7988 & ~v_7989 & ~v_8007;
assign v_9073 = v_9070 & ~v_7990;
assign v_9074 = v_9070 & v_7998 & ~v_7999;
assign v_9075 = v_9070 & v_8631;
assign v_9077 = v_9076 & v_7988 & v_7989 & v_8004 & ~v_8005;
assign v_9079 = v_9078 & v_8011 & ~v_8012 & v_8030;
assign v_9080 = v_9078 & v_8011 & ~v_8012 & ~v_8030;
assign v_9081 = v_9078 & ~v_8013;
assign v_9082 = v_9078 & v_8021 & ~v_8022;
assign v_9083 = v_9078 & v_8640;
assign v_9085 = v_9084 & v_8011 & v_8012 & v_8027 & ~v_8028;
assign v_9087 = v_9086 & v_8034 & ~v_8035 & v_8053;
assign v_9088 = v_9086 & ~v_8036;
assign v_9089 = v_9086 & v_8044 & ~v_8045;
assign v_9090 = v_9086 & v_8648;
assign v_9092 = v_9091 & v_8034 & v_8035 & v_8050 & v_8051;
assign v_9093 = v_9086 & v_8034 & ~v_8035 & ~v_8053;
assign v_9094 = v_9091 & v_8034 & v_8035 & v_8050 & ~v_8051;
assign v_9097 = v_9095 & v_9096;
assign v_9098 = v_9095 & v_8057 & v_8058 & ~v_8059 & ~v_8060;
assign v_9099 = v_9095 & v_8057 & v_8058 & v_8059;
assign v_9100 = v_9095 & v_8057 & ~v_8058 & ~v_8062;
assign v_9102 = v_9101 & v_8661;
assign v_9103 = v_9084 & v_8011 & v_8012 & v_8027 & v_8028;
assign v_9104 = v_9076 & v_7988 & v_7989 & v_8004 & v_8005;
assign v_9106 = v_9105 & v_8069 & ~v_8070 & v_8088;
assign v_9107 = v_9105 & v_8069 & ~v_8070 & ~v_8088;
assign v_9108 = v_9105 & ~v_8071;
assign v_9109 = v_9105 & v_8079 & ~v_8080;
assign v_9110 = v_9105 & v_8670;
assign v_9112 = v_9111 & v_8069 & v_8070 & v_8085 & ~v_8086;
assign v_9114 = v_9113 & v_8092 & ~v_8093 & v_8111;
assign v_9115 = v_9113 & v_8092 & ~v_8093 & ~v_8111;
assign v_9116 = v_9113 & ~v_8094;
assign v_9117 = v_9113 & v_8102 & ~v_8103;
assign v_9118 = v_9113 & v_8679;
assign v_9120 = v_9119 & v_8092 & v_8093 & v_8108 & ~v_8109;
assign v_9122 = v_9121 & v_8115 & ~v_8116 & v_8134;
assign v_9123 = v_9121 & ~v_8117;
assign v_9124 = v_9121 & v_8125 & ~v_8126;
assign v_9125 = v_9121 & v_8687;
assign v_9127 = v_9126 & v_8115 & v_8116 & v_8131 & v_8132;
assign v_9128 = v_9121 & v_8115 & ~v_8116 & ~v_8134;
assign v_9129 = v_9126 & v_8115 & v_8116 & v_8131 & ~v_8132;
assign v_9132 = v_9130 & v_9131;
assign v_9133 = v_9130 & v_8138 & v_8139 & ~v_8140 & ~v_8141;
assign v_9134 = v_9130 & v_8138 & v_8139 & v_8140;
assign v_9135 = v_9130 & v_8138 & ~v_8139 & ~v_8143;
assign v_9137 = v_9136 & v_8700;
assign v_9138 = v_9119 & v_8092 & v_8093 & v_8108 & v_8109;
assign v_9139 = v_9111 & v_8069 & v_8070 & v_8085 & v_8086;
assign v_9141 = v_9140 & v_8150 & ~v_8151 & v_8169;
assign v_9142 = v_9140 & v_8150 & ~v_8151 & ~v_8169;
assign v_9143 = v_9140 & ~v_8152;
assign v_9144 = v_9140 & v_8160 & ~v_8161;
assign v_9145 = v_9140 & v_8709;
assign v_9147 = v_9146 & v_8150 & v_8151 & v_8166 & ~v_8167;
assign v_9149 = v_9148 & v_8173 & ~v_8174 & v_8192;
assign v_9150 = v_9148 & v_8173 & ~v_8174 & ~v_8192;
assign v_9151 = v_9148 & ~v_8175;
assign v_9152 = v_9148 & v_8183 & ~v_8184;
assign v_9153 = v_9148 & v_8718;
assign v_9155 = v_9154 & v_8173 & v_8174 & v_8189 & ~v_8190;
assign v_9157 = v_9156 & v_8196 & ~v_8197 & v_8215;
assign v_9158 = v_9156 & ~v_8198;
assign v_9159 = v_9156 & v_8206 & ~v_8207;
assign v_9160 = v_9156 & v_8726;
assign v_9162 = v_9161 & v_8196 & v_8197 & v_8212 & v_8213;
assign v_9163 = v_9156 & v_8196 & ~v_8197 & ~v_8215;
assign v_9164 = v_9161 & v_8196 & v_8197 & v_8212 & ~v_8213;
assign v_9167 = v_9165 & v_9166;
assign v_9168 = v_9165 & v_8219 & v_8220 & ~v_8221 & ~v_8222;
assign v_9169 = v_9165 & v_8219 & v_8220 & v_8221;
assign v_9170 = v_9165 & v_8219 & ~v_8220 & ~v_8224;
assign v_9172 = v_9171 & v_8739;
assign v_9173 = v_9154 & v_8173 & v_8174 & v_8189 & v_8190;
assign v_9174 = v_9146 & v_8150 & v_8151 & v_8166 & v_8167;
assign v_9176 = v_6874 & v_7093;
assign v_9177 = v_6874 & ~v_7093 & v_7095 & v_7128 & ~v_7130;
assign v_9178 = v_6874 & ~v_7093 & v_7095 & v_7128 & v_7130;
assign v_9179 = v_6874 & ~v_7093 & v_7095 & ~v_7128;
assign v_9180 = v_6874 & v_7096;
assign v_9181 = v_6874 & ~v_7096;
assign v_9184 = v_9182 & v_9183;
assign v_9185 = v_9182 & v_8244;
assign v_9186 = v_13239 & v_13240;
assign v_9188 = v_9187 & ~v_7093 & ~v_7095 & v_7126;
assign v_9190 = v_9189 & v_7133 & v_7134;
assign v_9191 = v_9189 & v_7133 & ~v_7134;
assign v_9193 = v_9192 & ~v_7145;
assign v_9195 = v_9192 & v_9194;
assign v_9196 = v_9192 & v_7145 & v_7157 & ~v_7158 & v_7166;
assign v_9199 = v_9197 & v_9198;
assign v_9200 = v_9197 & v_7187 & v_7188;
assign v_9201 = v_9197 & v_7187 & ~v_7188 & v_7190;
assign v_9202 = v_9197 & v_7187 & ~v_7188 & ~v_7190 & v_7192;
assign v_9203 = v_9197 & v_7187 & ~v_7188 & ~v_7190 & ~v_7192;
assign v_9205 = v_9204 & v_8267;
assign v_9207 = v_9206 & ~v_7174 & v_7175 & v_7195;
assign v_9210 = v_9208 & v_9209;
assign v_9211 = v_9208 & v_8274;
assign v_9213 = v_9212 & v_7211 & v_7212;
assign v_9214 = v_9212 & v_7211 & ~v_7212 & v_7214;
assign v_9215 = v_9212 & v_7211 & ~v_7212 & ~v_7214 & v_7216;
assign v_9216 = v_9212 & v_7222 & v_7223;
assign v_9217 = v_9212 & v_7225 & v_7226;
assign v_9218 = v_9212 & v_7225 & ~v_7226 & v_7228;
assign v_9219 = v_9212 & v_7225 & ~v_7226 & ~v_7228 & v_7230;
assign v_9220 = v_9212 & v_8286;
assign v_9222 = v_9221 & v_8289;
assign v_9224 = v_9223 & v_7222 & ~v_7223 & v_7235 & v_7236;
assign v_9225 = v_9223 & v_7238 & v_7239;
assign v_9226 = v_9223 & v_7238 & ~v_7239 & v_7241;
assign v_9227 = v_9223 & v_7238 & ~v_7239 & ~v_7241 & v_7243;
assign v_9229 = v_9223 & v_9228;
assign v_9230 = v_13241 & v_13242;
assign v_9232 = v_9231 & v_7250 & v_7251;
assign v_9233 = v_9231 & v_7250 & ~v_7251;
assign v_9235 = v_9234 & v_8303;
assign v_9237 = v_13243 & v_13244;
assign v_9238 = v_9236 & v_7257 & v_7258;
assign v_9239 = v_9236 & v_7257 & ~v_7258 & v_7260;
assign v_9240 = v_9236 & v_7257 & ~v_7258 & ~v_7260 & v_7262;
assign v_9241 = v_9236 & v_8310;
assign v_9243 = v_13245 & v_13246;
assign v_9245 = v_9244 & v_8315;
assign v_9247 = v_9246 & v_7276 & v_7277;
assign v_9248 = v_9246 & v_7276 & ~v_7277 & v_7279;
assign v_9249 = v_9246 & v_7276 & ~v_7277 & ~v_7279 & v_7281;
assign v_9250 = v_9246 & v_7287 & v_7288;
assign v_9251 = v_9246 & v_7290 & v_7291;
assign v_9252 = v_9246 & v_7290 & ~v_7291 & v_7293;
assign v_9253 = v_9246 & v_7290 & ~v_7291 & ~v_7293 & v_7295;
assign v_9254 = v_9246 & v_8325;
assign v_9256 = v_9255 & v_8328;
assign v_9258 = v_9257 & v_7287 & ~v_7288 & v_7300 & v_7301;
assign v_9259 = v_9257 & v_7303 & v_7304;
assign v_9260 = v_9257 & v_7303 & ~v_7304 & v_7306;
assign v_9261 = v_9257 & v_7303 & ~v_7304 & ~v_7306 & v_7308;
assign v_9263 = v_9257 & v_9262;
assign v_9264 = v_13247 & v_13248;
assign v_9266 = v_9265 & v_7315 & v_7316;
assign v_9267 = v_9265 & v_7315 & ~v_7316;
assign v_9269 = v_9268 & v_8342;
assign v_9271 = v_13249 & v_13250;
assign v_9272 = v_9270 & v_7322 & v_7323;
assign v_9273 = v_9270 & v_7322 & ~v_7323 & v_7325;
assign v_9274 = v_9270 & v_7322 & ~v_7323 & ~v_7325 & v_7327;
assign v_9275 = v_9270 & v_8349;
assign v_9277 = v_13251 & v_13252;
assign v_9279 = v_9278 & v_8354;
assign v_9281 = v_9280 & v_7357;
assign v_9282 = v_9280 & ~v_7357 & v_7359 & v_7392 & ~v_7394;
assign v_9283 = v_9280 & ~v_7357 & v_7359 & v_7392 & v_7394;
assign v_9284 = v_9280 & ~v_7357 & v_7359 & ~v_7392;
assign v_9285 = v_9280 & v_7360;
assign v_9286 = v_9280 & ~v_7360;
assign v_9289 = v_9287 & v_9288;
assign v_9290 = v_9287 & v_8370;
assign v_9291 = v_13253 & v_13254;
assign v_9293 = v_9292 & ~v_7357 & ~v_7359 & v_7390;
assign v_9295 = v_9294 & v_7397 & v_7398;
assign v_9296 = v_9294 & v_7397 & ~v_7398;
assign v_9298 = v_9297 & v_7412 & v_7413;
assign v_9299 = v_9297 & v_7412 & ~v_7413 & ~v_7417;
assign v_9301 = v_9300 & v_7412 & ~v_7413 & v_7417;
assign v_9303 = v_9302 & v_7420;
assign v_9305 = v_9304 & v_7424 & v_7425;
assign v_9306 = v_9304 & v_7424 & ~v_7425 & v_7427;
assign v_9307 = v_9304 & v_8386;
assign v_9310 = v_9308 & v_9309;
assign v_9311 = v_9308 & v_8391;
assign v_9313 = v_9312 & v_7454 & ~v_7455 & ~v_7457;
assign v_9314 = v_9312 & v_7459 & ~v_7460;
assign v_9315 = v_9312 & v_7459 & v_7460;
assign v_9316 = v_9312 & v_7449;
assign v_9318 = v_9317 & v_7470 & v_7471;
assign v_9319 = v_9317 & v_7470 & ~v_7471 & ~v_7475;
assign v_9321 = v_9320 & v_7470 & ~v_7471 & v_7475;
assign v_9323 = v_9322 & v_7478;
assign v_9325 = v_9324 & v_7482 & v_7483;
assign v_9326 = v_9324 & v_7482 & ~v_7483 & v_7485;
assign v_9327 = v_9324 & v_8404;
assign v_9330 = v_9328 & v_9329;
assign v_9331 = v_9328 & v_8409;
assign v_9333 = v_6868 & v_9332;
assign v_9334 = v_7507 & v_9312;
assign v_9335 = v_7509 & v_9297;
assign v_9336 = v_7511 & v_9297;
assign v_9337 = v_7513 & v_9297;
assign v_9338 = v_7515 & v_9297;
assign v_9339 = ~v_7515 & v_9280;
assign v_9341 = ~v_7513 & v_9340;
assign v_9343 = ~v_7511 & v_9342;
assign v_9345 = ~v_7509 & v_9344;
assign v_9347 = ~v_7507 & v_9346;
assign v_9349 = ~v_6868 & v_9348;
assign v_9351 = v_9350 & ~v_7535;
assign v_9352 = v_13255 & v_13256;
assign v_9353 = v_9350 & v_7535 & v_7536 & v_7538 & v_7540;
assign v_9354 = v_13257 & v_13258;
assign v_9356 = v_9355 & v_7545 & ~v_7546 & v_7548;
assign v_9357 = v_9355 & v_7555 & ~v_7556 & ~v_7558;
assign v_9358 = v_9355 & v_7560 & ~v_7561;
assign v_9359 = v_9355 & v_7560 & v_7561;
assign v_9360 = v_9355 & v_7550;
assign v_9362 = v_9361 & v_8441;
assign v_9364 = v_9363 & v_8444;
assign v_9365 = v_9355 & v_7545 & v_7546;
assign v_9366 = v_9350 & v_8447;
assign v_9368 = v_9367 & ~v_7571;
assign v_9369 = v_9367 & v_7576 & v_7577;
assign v_9370 = v_9367 & v_7576 & ~v_7577 & ~v_7581;
assign v_9372 = v_9371 & v_7576 & ~v_7577 & v_7581;
assign v_9374 = v_9373 & v_7584;
assign v_9376 = v_9375 & v_7571 & v_7588 & v_7589 & ~v_7590;
assign v_9378 = v_9375 & v_9377;
assign v_9379 = v_9375 & v_7616 & v_7617;
assign v_9380 = v_9375 & v_7616 & ~v_7617;
assign v_9382 = v_9381 & v_7629 & v_7630;
assign v_9383 = v_9381 & v_7629 & ~v_7630;
assign v_9385 = v_9384 & v_7611 & v_7624 & v_7637;
assign v_9386 = v_13259 & v_13260;
assign v_9387 = v_9375 & v_7645 & v_7646;
assign v_9388 = v_9375 & v_7645 & ~v_7646 & ~v_7650;
assign v_9390 = v_9389 & v_7645 & ~v_7646 & v_7650;
assign v_9392 = v_9391 & v_7653;
assign v_9394 = v_9393 & v_8468;
assign v_9396 = v_9395 & v_7664 & ~v_7665 & v_7683;
assign v_9397 = v_9395 & v_7664 & ~v_7665 & ~v_7683;
assign v_9398 = v_9395 & ~v_7666;
assign v_9399 = v_9395 & v_7674 & ~v_7675;
assign v_9400 = v_9395 & v_8475;
assign v_9402 = v_9401 & v_7664 & v_7665 & v_7680 & ~v_7681;
assign v_9404 = v_9403 & v_7687 & ~v_7688 & v_7706;
assign v_9405 = v_9403 & v_7687 & ~v_7688 & ~v_7706;
assign v_9406 = v_9403 & ~v_7689;
assign v_9407 = v_9403 & v_7697 & ~v_7698;
assign v_9408 = v_9403 & v_8484;
assign v_9410 = v_9409 & v_7687 & v_7688 & v_7703 & ~v_7704;
assign v_9412 = v_9411 & v_7710 & ~v_7711 & v_7729;
assign v_9413 = v_9411 & ~v_7712;
assign v_9414 = v_9411 & v_7720 & ~v_7721;
assign v_9415 = v_9411 & v_8492;
assign v_9417 = v_9416 & v_7710 & v_7711 & v_7726 & v_7727;
assign v_9418 = v_9411 & v_7710 & ~v_7711 & ~v_7729;
assign v_9419 = v_9416 & v_7710 & v_7711 & v_7726 & ~v_7727;
assign v_9422 = v_9420 & v_9421;
assign v_9423 = v_9420 & v_7733 & v_7734 & ~v_7735 & ~v_7736;
assign v_9424 = v_9420 & v_7733 & v_7734 & v_7735;
assign v_9425 = v_9420 & v_7733 & ~v_7734 & ~v_7738;
assign v_9427 = v_9426 & v_8505;
assign v_9428 = v_9409 & v_7687 & v_7688 & v_7703 & v_7704;
assign v_9429 = v_9401 & v_7664 & v_7665 & v_7680 & v_7681;
assign v_9431 = v_9430 & v_7745 & ~v_7746 & v_7764;
assign v_9432 = v_9430 & v_7745 & ~v_7746 & ~v_7764;
assign v_9433 = v_9430 & ~v_7747;
assign v_9434 = v_9430 & v_7755 & ~v_7756;
assign v_9435 = v_9430 & v_8514;
assign v_9437 = v_9436 & v_7745 & v_7746 & v_7761 & ~v_7762;
assign v_9439 = v_9438 & v_7768 & ~v_7769 & v_7787;
assign v_9440 = v_9438 & v_7768 & ~v_7769 & ~v_7787;
assign v_9441 = v_9438 & ~v_7770;
assign v_9442 = v_9438 & v_7778 & ~v_7779;
assign v_9443 = v_9438 & v_8523;
assign v_9445 = v_9444 & v_7768 & v_7769 & v_7784 & ~v_7785;
assign v_9447 = v_9446 & v_7791 & ~v_7792 & v_7810;
assign v_9448 = v_9446 & ~v_7793;
assign v_9449 = v_9446 & v_7801 & ~v_7802;
assign v_9450 = v_9446 & v_8531;
assign v_9452 = v_9451 & v_7791 & v_7792 & v_7807 & v_7808;
assign v_9453 = v_9446 & v_7791 & ~v_7792 & ~v_7810;
assign v_9454 = v_9451 & v_7791 & v_7792 & v_7807 & ~v_7808;
assign v_9457 = v_9455 & v_9456;
assign v_9458 = v_9455 & v_7814 & v_7815 & ~v_7816 & ~v_7817;
assign v_9459 = v_9455 & v_7814 & v_7815 & v_7816;
assign v_9460 = v_9455 & v_7814 & ~v_7815 & ~v_7819;
assign v_9462 = v_9461 & v_8544;
assign v_9463 = v_9444 & v_7768 & v_7769 & v_7784 & v_7785;
assign v_9464 = v_9436 & v_7745 & v_7746 & v_7761 & v_7762;
assign v_9466 = v_9465 & v_7826 & ~v_7827 & v_7845;
assign v_9467 = v_9465 & v_7826 & ~v_7827 & ~v_7845;
assign v_9468 = v_9465 & ~v_7828;
assign v_9469 = v_9465 & v_7836 & ~v_7837;
assign v_9470 = v_9465 & v_8553;
assign v_9472 = v_9471 & v_7826 & v_7827 & v_7842 & ~v_7843;
assign v_9474 = v_9473 & v_7849 & ~v_7850 & v_7868;
assign v_9475 = v_9473 & v_7849 & ~v_7850 & ~v_7868;
assign v_9476 = v_9473 & ~v_7851;
assign v_9477 = v_9473 & v_7859 & ~v_7860;
assign v_9478 = v_9473 & v_8562;
assign v_9480 = v_9479 & v_7849 & v_7850 & v_7865 & ~v_7866;
assign v_9482 = v_9481 & v_7872 & ~v_7873 & v_7891;
assign v_9483 = v_9481 & ~v_7874;
assign v_9484 = v_9481 & v_7882 & ~v_7883;
assign v_9485 = v_9481 & v_8570;
assign v_9487 = v_9486 & v_7872 & v_7873 & v_7888 & v_7889;
assign v_9488 = v_9481 & v_7872 & ~v_7873 & ~v_7891;
assign v_9489 = v_9486 & v_7872 & v_7873 & v_7888 & ~v_7889;
assign v_9492 = v_9490 & v_9491;
assign v_9493 = v_9490 & v_7895 & v_7896 & ~v_7897 & ~v_7898;
assign v_9494 = v_9490 & v_7895 & v_7896 & v_7897;
assign v_9495 = v_9490 & v_7895 & ~v_7896 & ~v_7900;
assign v_9497 = v_9496 & v_8583;
assign v_9498 = v_9479 & v_7849 & v_7850 & v_7865 & v_7866;
assign v_9499 = v_9471 & v_7826 & v_7827 & v_7842 & v_7843;
assign v_9501 = v_9500 & v_7907 & ~v_7908 & v_7926;
assign v_9502 = v_9500 & v_7907 & ~v_7908 & ~v_7926;
assign v_9503 = v_9500 & ~v_7909;
assign v_9504 = v_9500 & v_7917 & ~v_7918;
assign v_9505 = v_9500 & v_8592;
assign v_9507 = v_9506 & v_7907 & v_7908 & v_7923 & ~v_7924;
assign v_9509 = v_9508 & v_7930 & ~v_7931 & v_7949;
assign v_9510 = v_9508 & v_7930 & ~v_7931 & ~v_7949;
assign v_9511 = v_9508 & ~v_7932;
assign v_9512 = v_9508 & v_7940 & ~v_7941;
assign v_9513 = v_9508 & v_8601;
assign v_9515 = v_9514 & v_7930 & v_7931 & v_7946 & ~v_7947;
assign v_9517 = v_9516 & v_7953 & ~v_7954 & v_7972;
assign v_9518 = v_9516 & ~v_7955;
assign v_9519 = v_9516 & v_7963 & ~v_7964;
assign v_9520 = v_9516 & v_8609;
assign v_9522 = v_9521 & v_7953 & v_7954 & v_7969 & v_7970;
assign v_9523 = v_9516 & v_7953 & ~v_7954 & ~v_7972;
assign v_9524 = v_9521 & v_7953 & v_7954 & v_7969 & ~v_7970;
assign v_9527 = v_9525 & v_9526;
assign v_9528 = v_9525 & v_7976 & v_7977 & ~v_7978 & ~v_7979;
assign v_9529 = v_9525 & v_7976 & v_7977 & v_7978;
assign v_9530 = v_9525 & v_7976 & ~v_7977 & ~v_7981;
assign v_9532 = v_9531 & v_8622;
assign v_9533 = v_9514 & v_7930 & v_7931 & v_7946 & v_7947;
assign v_9534 = v_9506 & v_7907 & v_7908 & v_7923 & v_7924;
assign v_9536 = v_9535 & v_7988 & ~v_7989 & v_8007;
assign v_9537 = v_9535 & v_7988 & ~v_7989 & ~v_8007;
assign v_9538 = v_9535 & ~v_7990;
assign v_9539 = v_9535 & v_7998 & ~v_7999;
assign v_9540 = v_9535 & v_8631;
assign v_9542 = v_9541 & v_7988 & v_7989 & v_8004 & ~v_8005;
assign v_9544 = v_9543 & v_8011 & ~v_8012 & v_8030;
assign v_9545 = v_9543 & v_8011 & ~v_8012 & ~v_8030;
assign v_9546 = v_9543 & ~v_8013;
assign v_9547 = v_9543 & v_8021 & ~v_8022;
assign v_9548 = v_9543 & v_8640;
assign v_9550 = v_9549 & v_8011 & v_8012 & v_8027 & ~v_8028;
assign v_9552 = v_9551 & v_8034 & ~v_8035 & v_8053;
assign v_9553 = v_9551 & ~v_8036;
assign v_9554 = v_9551 & v_8044 & ~v_8045;
assign v_9555 = v_9551 & v_8648;
assign v_9557 = v_9556 & v_8034 & v_8035 & v_8050 & v_8051;
assign v_9558 = v_9551 & v_8034 & ~v_8035 & ~v_8053;
assign v_9559 = v_9556 & v_8034 & v_8035 & v_8050 & ~v_8051;
assign v_9562 = v_9560 & v_9561;
assign v_9563 = v_9560 & v_8057 & v_8058 & ~v_8059 & ~v_8060;
assign v_9564 = v_9560 & v_8057 & v_8058 & v_8059;
assign v_9565 = v_9560 & v_8057 & ~v_8058 & ~v_8062;
assign v_9567 = v_9566 & v_8661;
assign v_9568 = v_9549 & v_8011 & v_8012 & v_8027 & v_8028;
assign v_9569 = v_9541 & v_7988 & v_7989 & v_8004 & v_8005;
assign v_9571 = v_9570 & v_8069 & ~v_8070 & v_8088;
assign v_9572 = v_9570 & v_8069 & ~v_8070 & ~v_8088;
assign v_9573 = v_9570 & ~v_8071;
assign v_9574 = v_9570 & v_8079 & ~v_8080;
assign v_9575 = v_9570 & v_8670;
assign v_9577 = v_9576 & v_8069 & v_8070 & v_8085 & ~v_8086;
assign v_9579 = v_9578 & v_8092 & ~v_8093 & v_8111;
assign v_9580 = v_9578 & v_8092 & ~v_8093 & ~v_8111;
assign v_9581 = v_9578 & ~v_8094;
assign v_9582 = v_9578 & v_8102 & ~v_8103;
assign v_9583 = v_9578 & v_8679;
assign v_9585 = v_9584 & v_8092 & v_8093 & v_8108 & ~v_8109;
assign v_9587 = v_9586 & v_8115 & ~v_8116 & v_8134;
assign v_9588 = v_9586 & ~v_8117;
assign v_9589 = v_9586 & v_8125 & ~v_8126;
assign v_9590 = v_9586 & v_8687;
assign v_9592 = v_9591 & v_8115 & v_8116 & v_8131 & v_8132;
assign v_9593 = v_9586 & v_8115 & ~v_8116 & ~v_8134;
assign v_9594 = v_9591 & v_8115 & v_8116 & v_8131 & ~v_8132;
assign v_9597 = v_9595 & v_9596;
assign v_9598 = v_9595 & v_8138 & v_8139 & ~v_8140 & ~v_8141;
assign v_9599 = v_9595 & v_8138 & v_8139 & v_8140;
assign v_9600 = v_9595 & v_8138 & ~v_8139 & ~v_8143;
assign v_9602 = v_9601 & v_8700;
assign v_9603 = v_9584 & v_8092 & v_8093 & v_8108 & v_8109;
assign v_9604 = v_9576 & v_8069 & v_8070 & v_8085 & v_8086;
assign v_9606 = v_9605 & v_8150 & ~v_8151 & v_8169;
assign v_9607 = v_9605 & v_8150 & ~v_8151 & ~v_8169;
assign v_9608 = v_9605 & ~v_8152;
assign v_9609 = v_9605 & v_8160 & ~v_8161;
assign v_9610 = v_9605 & v_8709;
assign v_9612 = v_9611 & v_8150 & v_8151 & v_8166 & ~v_8167;
assign v_9614 = v_9613 & v_8173 & ~v_8174 & v_8192;
assign v_9615 = v_9613 & v_8173 & ~v_8174 & ~v_8192;
assign v_9616 = v_9613 & ~v_8175;
assign v_9617 = v_9613 & v_8183 & ~v_8184;
assign v_9618 = v_9613 & v_8718;
assign v_9620 = v_9619 & v_8173 & v_8174 & v_8189 & ~v_8190;
assign v_9622 = v_9621 & v_8196 & ~v_8197 & v_8215;
assign v_9623 = v_9621 & ~v_8198;
assign v_9624 = v_9621 & v_8206 & ~v_8207;
assign v_9625 = v_9621 & v_8726;
assign v_9627 = v_9626 & v_8196 & v_8197 & v_8212 & v_8213;
assign v_9628 = v_9621 & v_8196 & ~v_8197 & ~v_8215;
assign v_9629 = v_9626 & v_8196 & v_8197 & v_8212 & ~v_8213;
assign v_9632 = v_9630 & v_9631;
assign v_9633 = v_9630 & v_8219 & v_8220 & ~v_8221 & ~v_8222;
assign v_9634 = v_9630 & v_8219 & v_8220 & v_8221;
assign v_9635 = v_9630 & v_8219 & ~v_8220 & ~v_8224;
assign v_9637 = v_9636 & v_8739;
assign v_9638 = v_9619 & v_8173 & v_8174 & v_8189 & v_8190;
assign v_9639 = v_9611 & v_8150 & v_8151 & v_8166 & v_8167;
assign v_9641 = v_7093;
assign v_9642 = ~v_7093 & v_7095 & v_7128 & ~v_7130;
assign v_9643 = ~v_7093 & v_7095 & v_7128 & v_7130;
assign v_9644 = ~v_7093 & v_7095 & ~v_7128;
assign v_9647 = v_9646;
assign v_9648 = v_8244;
assign v_9649 = v_13261 & v_13262;
assign v_9651 = v_9650 & ~v_7093 & ~v_7095 & v_7126;
assign v_9653 = v_9652 & v_7133 & v_7134;
assign v_9654 = v_9652 & v_7133 & ~v_7134;
assign v_9656 = v_9655 & ~v_7145;
assign v_9658 = v_9655 & v_9657;
assign v_9659 = v_9655 & v_7145 & v_7157 & ~v_7158 & v_7166;
assign v_9662 = v_9660 & v_9661;
assign v_9663 = v_9660 & v_7187 & v_7188;
assign v_9664 = v_9660 & v_7187 & ~v_7188 & v_7190;
assign v_9665 = v_9660 & v_7187 & ~v_7188 & ~v_7190 & v_7192;
assign v_9666 = v_9660 & v_7187 & ~v_7188 & ~v_7190 & ~v_7192;
assign v_9668 = v_9667 & v_8267;
assign v_9670 = v_9669 & ~v_7174 & v_7175 & v_7195;
assign v_9673 = v_9671 & v_9672;
assign v_9674 = v_9671 & v_8274;
assign v_9676 = v_9675 & v_7211 & v_7212;
assign v_9677 = v_9675 & v_7211 & ~v_7212 & v_7214;
assign v_9678 = v_9675 & v_7211 & ~v_7212 & ~v_7214 & v_7216;
assign v_9679 = v_9675 & v_7222 & v_7223;
assign v_9680 = v_9675 & v_7225 & v_7226;
assign v_9681 = v_9675 & v_7225 & ~v_7226 & v_7228;
assign v_9682 = v_9675 & v_7225 & ~v_7226 & ~v_7228 & v_7230;
assign v_9683 = v_9675 & v_8286;
assign v_9685 = v_9684 & v_8289;
assign v_9687 = v_9686 & v_7222 & ~v_7223 & v_7235 & v_7236;
assign v_9688 = v_9686 & v_7238 & v_7239;
assign v_9689 = v_9686 & v_7238 & ~v_7239 & v_7241;
assign v_9690 = v_9686 & v_7238 & ~v_7239 & ~v_7241 & v_7243;
assign v_9692 = v_9686 & v_9691;
assign v_9693 = v_13263 & v_13264;
assign v_9695 = v_9694 & v_7250 & v_7251;
assign v_9696 = v_9694 & v_7250 & ~v_7251;
assign v_9698 = v_9697 & v_8303;
assign v_9700 = v_13265 & v_13266;
assign v_9701 = v_9699 & v_7257 & v_7258;
assign v_9702 = v_9699 & v_7257 & ~v_7258 & v_7260;
assign v_9703 = v_9699 & v_7257 & ~v_7258 & ~v_7260 & v_7262;
assign v_9704 = v_9699 & v_8310;
assign v_9706 = v_13267 & v_13268;
assign v_9708 = v_9707 & v_8315;
assign v_9710 = v_9709 & v_7276 & v_7277;
assign v_9711 = v_9709 & v_7276 & ~v_7277 & v_7279;
assign v_9712 = v_9709 & v_7276 & ~v_7277 & ~v_7279 & v_7281;
assign v_9713 = v_9709 & v_7287 & v_7288;
assign v_9714 = v_9709 & v_7290 & v_7291;
assign v_9715 = v_9709 & v_7290 & ~v_7291 & v_7293;
assign v_9716 = v_9709 & v_7290 & ~v_7291 & ~v_7293 & v_7295;
assign v_9717 = v_9709 & v_8325;
assign v_9719 = v_9718 & v_8328;
assign v_9721 = v_9720 & v_7287 & ~v_7288 & v_7300 & v_7301;
assign v_9722 = v_9720 & v_7303 & v_7304;
assign v_9723 = v_9720 & v_7303 & ~v_7304 & v_7306;
assign v_9724 = v_9720 & v_7303 & ~v_7304 & ~v_7306 & v_7308;
assign v_9726 = v_9720 & v_9725;
assign v_9727 = v_13269 & v_13270;
assign v_9729 = v_9728 & v_7315 & v_7316;
assign v_9730 = v_9728 & v_7315 & ~v_7316;
assign v_9732 = v_9731 & v_8342;
assign v_9734 = v_13271 & v_13272;
assign v_9735 = v_9733 & v_7322 & v_7323;
assign v_9736 = v_9733 & v_7322 & ~v_7323 & v_7325;
assign v_9737 = v_9733 & v_7322 & ~v_7323 & ~v_7325 & v_7327;
assign v_9738 = v_9733 & v_8349;
assign v_9740 = v_13273 & v_13274;
assign v_9742 = v_9741 & v_8354;
assign v_9744 = v_9743 & v_7357;
assign v_9745 = v_9743 & ~v_7357 & v_7359 & v_7392 & ~v_7394;
assign v_9746 = v_9743 & ~v_7357 & v_7359 & v_7392 & v_7394;
assign v_9747 = v_9743 & ~v_7357 & v_7359 & ~v_7392;
assign v_9748 = v_9743 & v_7360;
assign v_9749 = v_9743 & ~v_7360;
assign v_9752 = v_9750 & v_9751;
assign v_9753 = v_9750 & v_8370;
assign v_9754 = v_13275 & v_13276;
assign v_9756 = v_9755 & ~v_7357 & ~v_7359 & v_7390;
assign v_9758 = v_9757 & v_7397 & v_7398;
assign v_9759 = v_9757 & v_7397 & ~v_7398;
assign v_9761 = v_9760 & v_7412 & v_7413;
assign v_9762 = v_9760 & v_7412 & ~v_7413 & ~v_7417;
assign v_9764 = v_9763 & v_7412 & ~v_7413 & v_7417;
assign v_9766 = v_9765 & v_7420;
assign v_9768 = v_9767 & v_7424 & v_7425;
assign v_9769 = v_9767 & v_7424 & ~v_7425 & v_7427;
assign v_9770 = v_9767 & v_8386;
assign v_9773 = v_9771 & v_9772;
assign v_9774 = v_9771 & v_8391;
assign v_9776 = v_9775 & v_7454 & ~v_7455 & ~v_7457;
assign v_9777 = v_9775 & v_7459 & ~v_7460;
assign v_9778 = v_9775 & v_7459 & v_7460;
assign v_9779 = v_9775 & v_7449;
assign v_9781 = v_9780 & v_7470 & v_7471;
assign v_9782 = v_9780 & v_7470 & ~v_7471 & ~v_7475;
assign v_9784 = v_9783 & v_7470 & ~v_7471 & v_7475;
assign v_9786 = v_9785 & v_7478;
assign v_9788 = v_9787 & v_7482 & v_7483;
assign v_9789 = v_9787 & v_7482 & ~v_7483 & v_7485;
assign v_9790 = v_9787 & v_8404;
assign v_9793 = v_9791 & v_9792;
assign v_9794 = v_9791 & v_8409;
assign v_9796 = v_6868 & v_9795;
assign v_9797 = v_7507 & v_9775;
assign v_9798 = v_7509 & v_9760;
assign v_9799 = v_7511 & v_9760;
assign v_9800 = v_7513 & v_9760;
assign v_9801 = v_7515 & v_9760;
assign v_9802 = ~v_7515 & v_9743;
assign v_9804 = ~v_7513 & v_9803;
assign v_9806 = ~v_7511 & v_9805;
assign v_9808 = ~v_7509 & v_9807;
assign v_9810 = ~v_7507 & v_9809;
assign v_9812 = ~v_6868 & v_9811;
assign v_9814 = v_9813 & ~v_7535;
assign v_9815 = v_13277 & v_13278;
assign v_9816 = v_9813 & v_7535 & v_7536 & v_7538 & v_7540;
assign v_9817 = v_13279 & v_13280;
assign v_9819 = v_9818 & v_7545 & ~v_7546 & v_7548;
assign v_9820 = v_9818 & v_7555 & ~v_7556 & ~v_7558;
assign v_9821 = v_9818 & v_7560 & ~v_7561;
assign v_9822 = v_9818 & v_7560 & v_7561;
assign v_9823 = v_9818 & v_7550;
assign v_9825 = v_9824 & v_8441;
assign v_9827 = v_9826 & v_8444;
assign v_9828 = v_9818 & v_7545 & v_7546;
assign v_9829 = v_9813 & v_8447;
assign v_9831 = v_9830 & ~v_7571;
assign v_9832 = v_9830 & v_7576 & v_7577;
assign v_9833 = v_9830 & v_7576 & ~v_7577 & ~v_7581;
assign v_9835 = v_9834 & v_7576 & ~v_7577 & v_7581;
assign v_9837 = v_9836 & v_7584;
assign v_9839 = v_9838 & v_7571 & v_7588 & v_7589 & ~v_7590;
assign v_9841 = v_9838 & v_9840;
assign v_9842 = v_9838 & v_7616 & v_7617;
assign v_9843 = v_9838 & v_7616 & ~v_7617;
assign v_9845 = v_9844 & v_7629 & v_7630;
assign v_9846 = v_9844 & v_7629 & ~v_7630;
assign v_9848 = v_9847 & v_7611 & v_7624 & v_7637;
assign v_9849 = v_13281 & v_13282;
assign v_9850 = v_9838 & v_7645 & v_7646;
assign v_9851 = v_9838 & v_7645 & ~v_7646 & ~v_7650;
assign v_9853 = v_9852 & v_7645 & ~v_7646 & v_7650;
assign v_9855 = v_9854 & v_7653;
assign v_9857 = v_9856 & v_8468;
assign v_9859 = v_9858 & v_7664 & ~v_7665 & v_7683;
assign v_9860 = v_9858 & v_7664 & ~v_7665 & ~v_7683;
assign v_9861 = v_9858 & ~v_7666;
assign v_9862 = v_9858 & v_7674 & ~v_7675;
assign v_9863 = v_9858 & v_8475;
assign v_9865 = v_9864 & v_7664 & v_7665 & v_7680 & ~v_7681;
assign v_9867 = v_9866 & v_7687 & ~v_7688 & v_7706;
assign v_9868 = v_9866 & v_7687 & ~v_7688 & ~v_7706;
assign v_9869 = v_9866 & ~v_7689;
assign v_9870 = v_9866 & v_7697 & ~v_7698;
assign v_9871 = v_9866 & v_8484;
assign v_9873 = v_9872 & v_7687 & v_7688 & v_7703 & ~v_7704;
assign v_9875 = v_9874 & v_7710 & ~v_7711 & v_7729;
assign v_9876 = v_9874 & ~v_7712;
assign v_9877 = v_9874 & v_7720 & ~v_7721;
assign v_9878 = v_9874 & v_8492;
assign v_9880 = v_9879 & v_7710 & v_7711 & v_7726 & v_7727;
assign v_9881 = v_9874 & v_7710 & ~v_7711 & ~v_7729;
assign v_9882 = v_9879 & v_7710 & v_7711 & v_7726 & ~v_7727;
assign v_9885 = v_9883 & v_9884;
assign v_9886 = v_9883 & v_7733 & v_7734 & ~v_7735 & ~v_7736;
assign v_9887 = v_9883 & v_7733 & v_7734 & v_7735;
assign v_9888 = v_9883 & v_7733 & ~v_7734 & ~v_7738;
assign v_9890 = v_9889 & v_8505;
assign v_9891 = v_9872 & v_7687 & v_7688 & v_7703 & v_7704;
assign v_9892 = v_9864 & v_7664 & v_7665 & v_7680 & v_7681;
assign v_9894 = v_9893 & v_7745 & ~v_7746 & v_7764;
assign v_9895 = v_9893 & v_7745 & ~v_7746 & ~v_7764;
assign v_9896 = v_9893 & ~v_7747;
assign v_9897 = v_9893 & v_7755 & ~v_7756;
assign v_9898 = v_9893 & v_8514;
assign v_9900 = v_9899 & v_7745 & v_7746 & v_7761 & ~v_7762;
assign v_9902 = v_9901 & v_7768 & ~v_7769 & v_7787;
assign v_9903 = v_9901 & v_7768 & ~v_7769 & ~v_7787;
assign v_9904 = v_9901 & ~v_7770;
assign v_9905 = v_9901 & v_7778 & ~v_7779;
assign v_9906 = v_9901 & v_8523;
assign v_9908 = v_9907 & v_7768 & v_7769 & v_7784 & ~v_7785;
assign v_9910 = v_9909 & v_7791 & ~v_7792 & v_7810;
assign v_9911 = v_9909 & ~v_7793;
assign v_9912 = v_9909 & v_7801 & ~v_7802;
assign v_9913 = v_9909 & v_8531;
assign v_9915 = v_9914 & v_7791 & v_7792 & v_7807 & v_7808;
assign v_9916 = v_9909 & v_7791 & ~v_7792 & ~v_7810;
assign v_9917 = v_9914 & v_7791 & v_7792 & v_7807 & ~v_7808;
assign v_9920 = v_9918 & v_9919;
assign v_9921 = v_9918 & v_7814 & v_7815 & ~v_7816 & ~v_7817;
assign v_9922 = v_9918 & v_7814 & v_7815 & v_7816;
assign v_9923 = v_9918 & v_7814 & ~v_7815 & ~v_7819;
assign v_9925 = v_9924 & v_8544;
assign v_9926 = v_9907 & v_7768 & v_7769 & v_7784 & v_7785;
assign v_9927 = v_9899 & v_7745 & v_7746 & v_7761 & v_7762;
assign v_9929 = v_9928 & v_7826 & ~v_7827 & v_7845;
assign v_9930 = v_9928 & v_7826 & ~v_7827 & ~v_7845;
assign v_9931 = v_9928 & ~v_7828;
assign v_9932 = v_9928 & v_7836 & ~v_7837;
assign v_9933 = v_9928 & v_8553;
assign v_9935 = v_9934 & v_7826 & v_7827 & v_7842 & ~v_7843;
assign v_9937 = v_9936 & v_7849 & ~v_7850 & v_7868;
assign v_9938 = v_9936 & v_7849 & ~v_7850 & ~v_7868;
assign v_9939 = v_9936 & ~v_7851;
assign v_9940 = v_9936 & v_7859 & ~v_7860;
assign v_9941 = v_9936 & v_8562;
assign v_9943 = v_9942 & v_7849 & v_7850 & v_7865 & ~v_7866;
assign v_9945 = v_9944 & v_7872 & ~v_7873 & v_7891;
assign v_9946 = v_9944 & ~v_7874;
assign v_9947 = v_9944 & v_7882 & ~v_7883;
assign v_9948 = v_9944 & v_8570;
assign v_9950 = v_9949 & v_7872 & v_7873 & v_7888 & v_7889;
assign v_9951 = v_9944 & v_7872 & ~v_7873 & ~v_7891;
assign v_9952 = v_9949 & v_7872 & v_7873 & v_7888 & ~v_7889;
assign v_9955 = v_9953 & v_9954;
assign v_9956 = v_9953 & v_7895 & v_7896 & ~v_7897 & ~v_7898;
assign v_9957 = v_9953 & v_7895 & v_7896 & v_7897;
assign v_9958 = v_9953 & v_7895 & ~v_7896 & ~v_7900;
assign v_9960 = v_9959 & v_8583;
assign v_9961 = v_9942 & v_7849 & v_7850 & v_7865 & v_7866;
assign v_9962 = v_9934 & v_7826 & v_7827 & v_7842 & v_7843;
assign v_9964 = v_9963 & v_7907 & ~v_7908 & v_7926;
assign v_9965 = v_9963 & v_7907 & ~v_7908 & ~v_7926;
assign v_9966 = v_9963 & ~v_7909;
assign v_9967 = v_9963 & v_7917 & ~v_7918;
assign v_9968 = v_9963 & v_8592;
assign v_9970 = v_9969 & v_7907 & v_7908 & v_7923 & ~v_7924;
assign v_9972 = v_9971 & v_7930 & ~v_7931 & v_7949;
assign v_9973 = v_9971 & v_7930 & ~v_7931 & ~v_7949;
assign v_9974 = v_9971 & ~v_7932;
assign v_9975 = v_9971 & v_7940 & ~v_7941;
assign v_9976 = v_9971 & v_8601;
assign v_9978 = v_9977 & v_7930 & v_7931 & v_7946 & ~v_7947;
assign v_9980 = v_9979 & v_7953 & ~v_7954 & v_7972;
assign v_9981 = v_9979 & ~v_7955;
assign v_9982 = v_9979 & v_7963 & ~v_7964;
assign v_9983 = v_9979 & v_8609;
assign v_9985 = v_9984 & v_7953 & v_7954 & v_7969 & v_7970;
assign v_9986 = v_9979 & v_7953 & ~v_7954 & ~v_7972;
assign v_9987 = v_9984 & v_7953 & v_7954 & v_7969 & ~v_7970;
assign v_9990 = v_9988 & v_9989;
assign v_9991 = v_9988 & v_7976 & v_7977 & ~v_7978 & ~v_7979;
assign v_9992 = v_9988 & v_7976 & v_7977 & v_7978;
assign v_9993 = v_9988 & v_7976 & ~v_7977 & ~v_7981;
assign v_9995 = v_9994 & v_8622;
assign v_9996 = v_9977 & v_7930 & v_7931 & v_7946 & v_7947;
assign v_9997 = v_9969 & v_7907 & v_7908 & v_7923 & v_7924;
assign v_9999 = v_9998 & v_7988 & ~v_7989 & v_8007;
assign v_10000 = v_9998 & v_7988 & ~v_7989 & ~v_8007;
assign v_10001 = v_9998 & ~v_7990;
assign v_10002 = v_9998 & v_7998 & ~v_7999;
assign v_10003 = v_9998 & v_8631;
assign v_10005 = v_10004 & v_7988 & v_7989 & v_8004 & ~v_8005;
assign v_10007 = v_10006 & v_8011 & ~v_8012 & v_8030;
assign v_10008 = v_10006 & v_8011 & ~v_8012 & ~v_8030;
assign v_10009 = v_10006 & ~v_8013;
assign v_10010 = v_10006 & v_8021 & ~v_8022;
assign v_10011 = v_10006 & v_8640;
assign v_10013 = v_10012 & v_8011 & v_8012 & v_8027 & ~v_8028;
assign v_10015 = v_10014 & v_8034 & ~v_8035 & v_8053;
assign v_10016 = v_10014 & ~v_8036;
assign v_10017 = v_10014 & v_8044 & ~v_8045;
assign v_10018 = v_10014 & v_8648;
assign v_10020 = v_10019 & v_8034 & v_8035 & v_8050 & v_8051;
assign v_10021 = v_10014 & v_8034 & ~v_8035 & ~v_8053;
assign v_10022 = v_10019 & v_8034 & v_8035 & v_8050 & ~v_8051;
assign v_10025 = v_10023 & v_10024;
assign v_10026 = v_10023 & v_8057 & v_8058 & ~v_8059 & ~v_8060;
assign v_10027 = v_10023 & v_8057 & v_8058 & v_8059;
assign v_10028 = v_10023 & v_8057 & ~v_8058 & ~v_8062;
assign v_10030 = v_10029 & v_8661;
assign v_10031 = v_10012 & v_8011 & v_8012 & v_8027 & v_8028;
assign v_10032 = v_10004 & v_7988 & v_7989 & v_8004 & v_8005;
assign v_10034 = v_10033 & v_8069 & ~v_8070 & v_8088;
assign v_10035 = v_10033 & v_8069 & ~v_8070 & ~v_8088;
assign v_10036 = v_10033 & ~v_8071;
assign v_10037 = v_10033 & v_8079 & ~v_8080;
assign v_10038 = v_10033 & v_8670;
assign v_10040 = v_10039 & v_8069 & v_8070 & v_8085 & ~v_8086;
assign v_10042 = v_10041 & v_8092 & ~v_8093 & v_8111;
assign v_10043 = v_10041 & v_8092 & ~v_8093 & ~v_8111;
assign v_10044 = v_10041 & ~v_8094;
assign v_10045 = v_10041 & v_8102 & ~v_8103;
assign v_10046 = v_10041 & v_8679;
assign v_10048 = v_10047 & v_8092 & v_8093 & v_8108 & ~v_8109;
assign v_10050 = v_10049 & v_8115 & ~v_8116 & v_8134;
assign v_10051 = v_10049 & ~v_8117;
assign v_10052 = v_10049 & v_8125 & ~v_8126;
assign v_10053 = v_10049 & v_8687;
assign v_10055 = v_10054 & v_8115 & v_8116 & v_8131 & v_8132;
assign v_10056 = v_10049 & v_8115 & ~v_8116 & ~v_8134;
assign v_10057 = v_10054 & v_8115 & v_8116 & v_8131 & ~v_8132;
assign v_10060 = v_10058 & v_10059;
assign v_10061 = v_10058 & v_8138 & v_8139 & ~v_8140 & ~v_8141;
assign v_10062 = v_10058 & v_8138 & v_8139 & v_8140;
assign v_10063 = v_10058 & v_8138 & ~v_8139 & ~v_8143;
assign v_10065 = v_10064 & v_8700;
assign v_10066 = v_10047 & v_8092 & v_8093 & v_8108 & v_8109;
assign v_10067 = v_10039 & v_8069 & v_8070 & v_8085 & v_8086;
assign v_10069 = v_10068 & v_8150 & ~v_8151 & v_8169;
assign v_10070 = v_10068 & v_8150 & ~v_8151 & ~v_8169;
assign v_10071 = v_10068 & ~v_8152;
assign v_10072 = v_10068 & v_8160 & ~v_8161;
assign v_10073 = v_10068 & v_8709;
assign v_10075 = v_10074 & v_8150 & v_8151 & v_8166 & ~v_8167;
assign v_10077 = v_10076 & v_8173 & ~v_8174 & v_8192;
assign v_10078 = v_10076 & v_8173 & ~v_8174 & ~v_8192;
assign v_10079 = v_10076 & ~v_8175;
assign v_10080 = v_10076 & v_8183 & ~v_8184;
assign v_10081 = v_10076 & v_8718;
assign v_10083 = v_10082 & v_8173 & v_8174 & v_8189 & ~v_8190;
assign v_10085 = v_10084 & v_8196 & ~v_8197 & v_8215;
assign v_10086 = v_10084 & ~v_8198;
assign v_10087 = v_10084 & v_8206 & ~v_8207;
assign v_10088 = v_10084 & v_8726;
assign v_10090 = v_10089 & v_8196 & v_8197 & v_8212 & v_8213;
assign v_10091 = v_10084 & v_8196 & ~v_8197 & ~v_8215;
assign v_10092 = v_10089 & v_8196 & v_8197 & v_8212 & ~v_8213;
assign v_10095 = v_10093 & v_10094;
assign v_10096 = v_10093 & v_8219 & v_8220 & ~v_8221 & ~v_8222;
assign v_10097 = v_10093 & v_8219 & v_8220 & v_8221;
assign v_10098 = v_10093 & v_8219 & ~v_8220 & ~v_8224;
assign v_10100 = v_10099 & v_8739;
assign v_10101 = v_10082 & v_8173 & v_8174 & v_8189 & v_8190;
assign v_10102 = v_10074 & v_8150 & v_8151 & v_8166 & v_8167;
assign v_10105 = v_10104 & v_7093;
assign v_10106 = v_10104 & ~v_7093 & v_7095 & v_7128 & ~v_7130;
assign v_10107 = v_10104 & ~v_7093 & v_7095 & v_7128 & v_7130;
assign v_10108 = v_10104 & ~v_7093 & v_7095 & ~v_7128;
assign v_10109 = v_10104 & v_7096;
assign v_10110 = v_10104 & ~v_7096;
assign v_10113 = v_10111 & v_10112;
assign v_10114 = v_10111 & v_8244;
assign v_10115 = v_13283 & v_13284;
assign v_10117 = v_10116 & ~v_7093 & ~v_7095 & v_7126;
assign v_10119 = v_10118 & v_7133 & v_7134;
assign v_10120 = v_10118 & v_7133 & ~v_7134;
assign v_10122 = v_10121 & ~v_7145;
assign v_10124 = v_10121 & v_10123;
assign v_10125 = v_10121 & v_7145 & v_7157 & ~v_7158 & v_7166;
assign v_10128 = v_10126 & v_10127;
assign v_10129 = v_10126 & v_7187 & v_7188;
assign v_10130 = v_10126 & v_7187 & ~v_7188 & v_7190;
assign v_10131 = v_10126 & v_7187 & ~v_7188 & ~v_7190 & v_7192;
assign v_10132 = v_10126 & v_7187 & ~v_7188 & ~v_7190 & ~v_7192;
assign v_10134 = v_10133 & v_8267;
assign v_10136 = v_10135 & ~v_7174 & v_7175 & v_7195;
assign v_10139 = v_10137 & v_10138;
assign v_10140 = v_10137 & v_8274;
assign v_10142 = v_10141 & v_7211 & v_7212;
assign v_10143 = v_10141 & v_7211 & ~v_7212 & v_7214;
assign v_10144 = v_10141 & v_7211 & ~v_7212 & ~v_7214 & v_7216;
assign v_10145 = v_10141 & v_7222 & v_7223;
assign v_10146 = v_10141 & v_7225 & v_7226;
assign v_10147 = v_10141 & v_7225 & ~v_7226 & v_7228;
assign v_10148 = v_10141 & v_7225 & ~v_7226 & ~v_7228 & v_7230;
assign v_10149 = v_10141 & v_8286;
assign v_10151 = v_10150 & v_8289;
assign v_10153 = v_10152 & v_7222 & ~v_7223 & v_7235 & v_7236;
assign v_10154 = v_10152 & v_7238 & v_7239;
assign v_10155 = v_10152 & v_7238 & ~v_7239 & v_7241;
assign v_10156 = v_10152 & v_7238 & ~v_7239 & ~v_7241 & v_7243;
assign v_10158 = v_10152 & v_10157;
assign v_10159 = v_13285 & v_13286;
assign v_10161 = v_10160 & v_7250 & v_7251;
assign v_10162 = v_10160 & v_7250 & ~v_7251;
assign v_10164 = v_10163 & v_8303;
assign v_10166 = v_13287 & v_13288;
assign v_10167 = v_10165 & v_7257 & v_7258;
assign v_10168 = v_10165 & v_7257 & ~v_7258 & v_7260;
assign v_10169 = v_10165 & v_7257 & ~v_7258 & ~v_7260 & v_7262;
assign v_10170 = v_10165 & v_8310;
assign v_10172 = v_13289 & v_13290;
assign v_10174 = v_10173 & v_8315;
assign v_10176 = v_10175 & v_7276 & v_7277;
assign v_10177 = v_10175 & v_7276 & ~v_7277 & v_7279;
assign v_10178 = v_10175 & v_7276 & ~v_7277 & ~v_7279 & v_7281;
assign v_10179 = v_10175 & v_7287 & v_7288;
assign v_10180 = v_10175 & v_7290 & v_7291;
assign v_10181 = v_10175 & v_7290 & ~v_7291 & v_7293;
assign v_10182 = v_10175 & v_7290 & ~v_7291 & ~v_7293 & v_7295;
assign v_10183 = v_10175 & v_8325;
assign v_10185 = v_10184 & v_8328;
assign v_10187 = v_10186 & v_7287 & ~v_7288 & v_7300 & v_7301;
assign v_10188 = v_10186 & v_7303 & v_7304;
assign v_10189 = v_10186 & v_7303 & ~v_7304 & v_7306;
assign v_10190 = v_10186 & v_7303 & ~v_7304 & ~v_7306 & v_7308;
assign v_10192 = v_10186 & v_10191;
assign v_10193 = v_13291 & v_13292;
assign v_10195 = v_10194 & v_7315 & v_7316;
assign v_10196 = v_10194 & v_7315 & ~v_7316;
assign v_10198 = v_10197 & v_8342;
assign v_10200 = v_13293 & v_13294;
assign v_10201 = v_10199 & v_7322 & v_7323;
assign v_10202 = v_10199 & v_7322 & ~v_7323 & v_7325;
assign v_10203 = v_10199 & v_7322 & ~v_7323 & ~v_7325 & v_7327;
assign v_10204 = v_10199 & v_8349;
assign v_10206 = v_13295 & v_13296;
assign v_10208 = v_10207 & v_8354;
assign v_10210 = v_10209 & v_7357;
assign v_10211 = v_10209 & ~v_7357 & v_7359 & v_7392 & ~v_7394;
assign v_10212 = v_10209 & ~v_7357 & v_7359 & v_7392 & v_7394;
assign v_10213 = v_10209 & ~v_7357 & v_7359 & ~v_7392;
assign v_10214 = v_10209 & v_7360;
assign v_10215 = v_10209 & ~v_7360;
assign v_10218 = v_10216 & v_10217;
assign v_10219 = v_10216 & v_8370;
assign v_10220 = v_13297 & v_13298;
assign v_10222 = v_10221 & ~v_7357 & ~v_7359 & v_7390;
assign v_10224 = v_10223 & v_7397 & v_7398;
assign v_10225 = v_10223 & v_7397 & ~v_7398;
assign v_10227 = v_10226 & v_7412 & v_7413;
assign v_10228 = v_10226 & v_7412 & ~v_7413 & ~v_7417;
assign v_10230 = v_10229 & v_7412 & ~v_7413 & v_7417;
assign v_10232 = v_10231 & v_7420;
assign v_10234 = v_10233 & v_7424 & v_7425;
assign v_10235 = v_10233 & v_7424 & ~v_7425 & v_7427;
assign v_10236 = v_10233 & v_8386;
assign v_10239 = v_10237 & v_10238;
assign v_10240 = v_10237 & v_8391;
assign v_10242 = v_10241 & v_7454 & ~v_7455 & ~v_7457;
assign v_10243 = v_10241 & v_7459 & ~v_7460;
assign v_10244 = v_10241 & v_7459 & v_7460;
assign v_10245 = v_10241 & v_7449;
assign v_10247 = v_10246 & v_7470 & v_7471;
assign v_10248 = v_10246 & v_7470 & ~v_7471 & ~v_7475;
assign v_10250 = v_10249 & v_7470 & ~v_7471 & v_7475;
assign v_10252 = v_10251 & v_7478;
assign v_10254 = v_10253 & v_7482 & v_7483;
assign v_10255 = v_10253 & v_7482 & ~v_7483 & v_7485;
assign v_10256 = v_10253 & v_8404;
assign v_10259 = v_10257 & v_10258;
assign v_10260 = v_10257 & v_8409;
assign v_10262 = v_6868 & v_10261;
assign v_10263 = v_7507 & v_10241;
assign v_10264 = v_7509 & v_10226;
assign v_10265 = v_7511 & v_10226;
assign v_10266 = v_7513 & v_10226;
assign v_10267 = v_7515 & v_10226;
assign v_10268 = ~v_7515 & v_10209;
assign v_10270 = ~v_7513 & v_10269;
assign v_10272 = ~v_7511 & v_10271;
assign v_10274 = ~v_7509 & v_10273;
assign v_10276 = ~v_7507 & v_10275;
assign v_10278 = ~v_6868 & v_10277;
assign v_10280 = v_10279 & ~v_7535;
assign v_10281 = v_13299 & v_13300;
assign v_10282 = v_10279 & v_7535 & v_7536 & v_7538 & v_7540;
assign v_10283 = v_13301 & v_13302;
assign v_10285 = v_10284 & v_7545 & ~v_7546 & v_7548;
assign v_10286 = v_10284 & v_7555 & ~v_7556 & ~v_7558;
assign v_10287 = v_10284 & v_7560 & ~v_7561;
assign v_10288 = v_10284 & v_7560 & v_7561;
assign v_10289 = v_10284 & v_7550;
assign v_10291 = v_10290 & v_8441;
assign v_10293 = v_10292 & v_8444;
assign v_10294 = v_10284 & v_7545 & v_7546;
assign v_10295 = v_10279 & v_8447;
assign v_10297 = v_10296 & ~v_7571;
assign v_10298 = v_10296 & v_7576 & v_7577;
assign v_10299 = v_10296 & v_7576 & ~v_7577 & ~v_7581;
assign v_10301 = v_10300 & v_7576 & ~v_7577 & v_7581;
assign v_10303 = v_10302 & v_7584;
assign v_10305 = v_10304 & v_7571 & v_7588 & v_7589 & ~v_7590;
assign v_10307 = v_10304 & v_10306;
assign v_10308 = v_10304 & v_7616 & v_7617;
assign v_10309 = v_10304 & v_7616 & ~v_7617;
assign v_10311 = v_10310 & v_7629 & v_7630;
assign v_10312 = v_10310 & v_7629 & ~v_7630;
assign v_10314 = v_10313 & v_7611 & v_7624 & v_7637;
assign v_10315 = v_13303 & v_13304;
assign v_10316 = v_10304 & v_7645 & v_7646;
assign v_10317 = v_10304 & v_7645 & ~v_7646 & ~v_7650;
assign v_10319 = v_10318 & v_7645 & ~v_7646 & v_7650;
assign v_10321 = v_10320 & v_7653;
assign v_10323 = v_10322 & v_8468;
assign v_10325 = v_10324 & v_7664 & ~v_7665 & v_7683;
assign v_10326 = v_10324 & v_7664 & ~v_7665 & ~v_7683;
assign v_10327 = v_10324 & ~v_7666;
assign v_10328 = v_10324 & v_7674 & ~v_7675;
assign v_10329 = v_10324 & v_8475;
assign v_10331 = v_10330 & v_7664 & v_7665 & v_7680 & ~v_7681;
assign v_10333 = v_10332 & v_7687 & ~v_7688 & v_7706;
assign v_10334 = v_10332 & v_7687 & ~v_7688 & ~v_7706;
assign v_10335 = v_10332 & ~v_7689;
assign v_10336 = v_10332 & v_7697 & ~v_7698;
assign v_10337 = v_10332 & v_8484;
assign v_10339 = v_10338 & v_7687 & v_7688 & v_7703 & ~v_7704;
assign v_10341 = v_10340 & v_7710 & ~v_7711 & v_7729;
assign v_10342 = v_10340 & ~v_7712;
assign v_10343 = v_10340 & v_7720 & ~v_7721;
assign v_10344 = v_10340 & v_8492;
assign v_10346 = v_10345 & v_7710 & v_7711 & v_7726 & v_7727;
assign v_10347 = v_10340 & v_7710 & ~v_7711 & ~v_7729;
assign v_10348 = v_10345 & v_7710 & v_7711 & v_7726 & ~v_7727;
assign v_10351 = v_10349 & v_10350;
assign v_10352 = v_10349 & v_7733 & v_7734 & ~v_7735 & ~v_7736;
assign v_10353 = v_10349 & v_7733 & v_7734 & v_7735;
assign v_10354 = v_10349 & v_7733 & ~v_7734 & ~v_7738;
assign v_10356 = v_10355 & v_8505;
assign v_10357 = v_10338 & v_7687 & v_7688 & v_7703 & v_7704;
assign v_10358 = v_10330 & v_7664 & v_7665 & v_7680 & v_7681;
assign v_10360 = v_10359 & v_7745 & ~v_7746 & v_7764;
assign v_10361 = v_10359 & v_7745 & ~v_7746 & ~v_7764;
assign v_10362 = v_10359 & ~v_7747;
assign v_10363 = v_10359 & v_7755 & ~v_7756;
assign v_10364 = v_10359 & v_8514;
assign v_10366 = v_10365 & v_7745 & v_7746 & v_7761 & ~v_7762;
assign v_10368 = v_10367 & v_7768 & ~v_7769 & v_7787;
assign v_10369 = v_10367 & v_7768 & ~v_7769 & ~v_7787;
assign v_10370 = v_10367 & ~v_7770;
assign v_10371 = v_10367 & v_7778 & ~v_7779;
assign v_10372 = v_10367 & v_8523;
assign v_10374 = v_10373 & v_7768 & v_7769 & v_7784 & ~v_7785;
assign v_10376 = v_10375 & v_7791 & ~v_7792 & v_7810;
assign v_10377 = v_10375 & ~v_7793;
assign v_10378 = v_10375 & v_7801 & ~v_7802;
assign v_10379 = v_10375 & v_8531;
assign v_10381 = v_10380 & v_7791 & v_7792 & v_7807 & v_7808;
assign v_10382 = v_10375 & v_7791 & ~v_7792 & ~v_7810;
assign v_10383 = v_10380 & v_7791 & v_7792 & v_7807 & ~v_7808;
assign v_10386 = v_10384 & v_10385;
assign v_10387 = v_10384 & v_7814 & v_7815 & ~v_7816 & ~v_7817;
assign v_10388 = v_10384 & v_7814 & v_7815 & v_7816;
assign v_10389 = v_10384 & v_7814 & ~v_7815 & ~v_7819;
assign v_10391 = v_10390 & v_8544;
assign v_10392 = v_10373 & v_7768 & v_7769 & v_7784 & v_7785;
assign v_10393 = v_10365 & v_7745 & v_7746 & v_7761 & v_7762;
assign v_10395 = v_10394 & v_7826 & ~v_7827 & v_7845;
assign v_10396 = v_10394 & v_7826 & ~v_7827 & ~v_7845;
assign v_10397 = v_10394 & ~v_7828;
assign v_10398 = v_10394 & v_7836 & ~v_7837;
assign v_10399 = v_10394 & v_8553;
assign v_10401 = v_10400 & v_7826 & v_7827 & v_7842 & ~v_7843;
assign v_10403 = v_10402 & v_7849 & ~v_7850 & v_7868;
assign v_10404 = v_10402 & v_7849 & ~v_7850 & ~v_7868;
assign v_10405 = v_10402 & ~v_7851;
assign v_10406 = v_10402 & v_7859 & ~v_7860;
assign v_10407 = v_10402 & v_8562;
assign v_10409 = v_10408 & v_7849 & v_7850 & v_7865 & ~v_7866;
assign v_10411 = v_10410 & v_7872 & ~v_7873 & v_7891;
assign v_10412 = v_10410 & ~v_7874;
assign v_10413 = v_10410 & v_7882 & ~v_7883;
assign v_10414 = v_10410 & v_8570;
assign v_10416 = v_10415 & v_7872 & v_7873 & v_7888 & v_7889;
assign v_10417 = v_10410 & v_7872 & ~v_7873 & ~v_7891;
assign v_10418 = v_10415 & v_7872 & v_7873 & v_7888 & ~v_7889;
assign v_10421 = v_10419 & v_10420;
assign v_10422 = v_10419 & v_7895 & v_7896 & ~v_7897 & ~v_7898;
assign v_10423 = v_10419 & v_7895 & v_7896 & v_7897;
assign v_10424 = v_10419 & v_7895 & ~v_7896 & ~v_7900;
assign v_10426 = v_10425 & v_8583;
assign v_10427 = v_10408 & v_7849 & v_7850 & v_7865 & v_7866;
assign v_10428 = v_10400 & v_7826 & v_7827 & v_7842 & v_7843;
assign v_10430 = v_10429 & v_7907 & ~v_7908 & v_7926;
assign v_10431 = v_10429 & v_7907 & ~v_7908 & ~v_7926;
assign v_10432 = v_10429 & ~v_7909;
assign v_10433 = v_10429 & v_7917 & ~v_7918;
assign v_10434 = v_10429 & v_8592;
assign v_10436 = v_10435 & v_7907 & v_7908 & v_7923 & ~v_7924;
assign v_10438 = v_10437 & v_7930 & ~v_7931 & v_7949;
assign v_10439 = v_10437 & v_7930 & ~v_7931 & ~v_7949;
assign v_10440 = v_10437 & ~v_7932;
assign v_10441 = v_10437 & v_7940 & ~v_7941;
assign v_10442 = v_10437 & v_8601;
assign v_10444 = v_10443 & v_7930 & v_7931 & v_7946 & ~v_7947;
assign v_10446 = v_10445 & v_7953 & ~v_7954 & v_7972;
assign v_10447 = v_10445 & ~v_7955;
assign v_10448 = v_10445 & v_7963 & ~v_7964;
assign v_10449 = v_10445 & v_8609;
assign v_10451 = v_10450 & v_7953 & v_7954 & v_7969 & v_7970;
assign v_10452 = v_10445 & v_7953 & ~v_7954 & ~v_7972;
assign v_10453 = v_10450 & v_7953 & v_7954 & v_7969 & ~v_7970;
assign v_10456 = v_10454 & v_10455;
assign v_10457 = v_10454 & v_7976 & v_7977 & ~v_7978 & ~v_7979;
assign v_10458 = v_10454 & v_7976 & v_7977 & v_7978;
assign v_10459 = v_10454 & v_7976 & ~v_7977 & ~v_7981;
assign v_10461 = v_10460 & v_8622;
assign v_10462 = v_10443 & v_7930 & v_7931 & v_7946 & v_7947;
assign v_10463 = v_10435 & v_7907 & v_7908 & v_7923 & v_7924;
assign v_10465 = v_10464 & v_7988 & ~v_7989 & v_8007;
assign v_10466 = v_10464 & v_7988 & ~v_7989 & ~v_8007;
assign v_10467 = v_10464 & ~v_7990;
assign v_10468 = v_10464 & v_7998 & ~v_7999;
assign v_10469 = v_10464 & v_8631;
assign v_10471 = v_10470 & v_7988 & v_7989 & v_8004 & ~v_8005;
assign v_10473 = v_10472 & v_8011 & ~v_8012 & v_8030;
assign v_10474 = v_10472 & v_8011 & ~v_8012 & ~v_8030;
assign v_10475 = v_10472 & ~v_8013;
assign v_10476 = v_10472 & v_8021 & ~v_8022;
assign v_10477 = v_10472 & v_8640;
assign v_10479 = v_10478 & v_8011 & v_8012 & v_8027 & ~v_8028;
assign v_10481 = v_10480 & v_8034 & ~v_8035 & v_8053;
assign v_10482 = v_10480 & ~v_8036;
assign v_10483 = v_10480 & v_8044 & ~v_8045;
assign v_10484 = v_10480 & v_8648;
assign v_10486 = v_10485 & v_8034 & v_8035 & v_8050 & v_8051;
assign v_10487 = v_10480 & v_8034 & ~v_8035 & ~v_8053;
assign v_10488 = v_10485 & v_8034 & v_8035 & v_8050 & ~v_8051;
assign v_10491 = v_10489 & v_10490;
assign v_10492 = v_10489 & v_8057 & v_8058 & ~v_8059 & ~v_8060;
assign v_10493 = v_10489 & v_8057 & v_8058 & v_8059;
assign v_10494 = v_10489 & v_8057 & ~v_8058 & ~v_8062;
assign v_10496 = v_10495 & v_8661;
assign v_10497 = v_10478 & v_8011 & v_8012 & v_8027 & v_8028;
assign v_10498 = v_10470 & v_7988 & v_7989 & v_8004 & v_8005;
assign v_10500 = v_10499 & v_8069 & ~v_8070 & v_8088;
assign v_10501 = v_10499 & v_8069 & ~v_8070 & ~v_8088;
assign v_10502 = v_10499 & ~v_8071;
assign v_10503 = v_10499 & v_8079 & ~v_8080;
assign v_10504 = v_10499 & v_8670;
assign v_10506 = v_10505 & v_8069 & v_8070 & v_8085 & ~v_8086;
assign v_10508 = v_10507 & v_8092 & ~v_8093 & v_8111;
assign v_10509 = v_10507 & v_8092 & ~v_8093 & ~v_8111;
assign v_10510 = v_10507 & ~v_8094;
assign v_10511 = v_10507 & v_8102 & ~v_8103;
assign v_10512 = v_10507 & v_8679;
assign v_10514 = v_10513 & v_8092 & v_8093 & v_8108 & ~v_8109;
assign v_10516 = v_10515 & v_8115 & ~v_8116 & v_8134;
assign v_10517 = v_10515 & ~v_8117;
assign v_10518 = v_10515 & v_8125 & ~v_8126;
assign v_10519 = v_10515 & v_8687;
assign v_10521 = v_10520 & v_8115 & v_8116 & v_8131 & v_8132;
assign v_10522 = v_10515 & v_8115 & ~v_8116 & ~v_8134;
assign v_10523 = v_10520 & v_8115 & v_8116 & v_8131 & ~v_8132;
assign v_10526 = v_10524 & v_10525;
assign v_10527 = v_10524 & v_8138 & v_8139 & ~v_8140 & ~v_8141;
assign v_10528 = v_10524 & v_8138 & v_8139 & v_8140;
assign v_10529 = v_10524 & v_8138 & ~v_8139 & ~v_8143;
assign v_10531 = v_10530 & v_8700;
assign v_10532 = v_10513 & v_8092 & v_8093 & v_8108 & v_8109;
assign v_10533 = v_10505 & v_8069 & v_8070 & v_8085 & v_8086;
assign v_10535 = v_10534 & v_8150 & ~v_8151 & v_8169;
assign v_10536 = v_10534 & v_8150 & ~v_8151 & ~v_8169;
assign v_10537 = v_10534 & ~v_8152;
assign v_10538 = v_10534 & v_8160 & ~v_8161;
assign v_10539 = v_10534 & v_8709;
assign v_10541 = v_10540 & v_8150 & v_8151 & v_8166 & ~v_8167;
assign v_10543 = v_10542 & v_8173 & ~v_8174 & v_8192;
assign v_10544 = v_10542 & v_8173 & ~v_8174 & ~v_8192;
assign v_10545 = v_10542 & ~v_8175;
assign v_10546 = v_10542 & v_8183 & ~v_8184;
assign v_10547 = v_10542 & v_8718;
assign v_10549 = v_10548 & v_8173 & v_8174 & v_8189 & ~v_8190;
assign v_10551 = v_10550 & v_8196 & ~v_8197 & v_8215;
assign v_10552 = v_10550 & ~v_8198;
assign v_10553 = v_10550 & v_8206 & ~v_8207;
assign v_10554 = v_10550 & v_8726;
assign v_10556 = v_10555 & v_8196 & v_8197 & v_8212 & v_8213;
assign v_10557 = v_10550 & v_8196 & ~v_8197 & ~v_8215;
assign v_10558 = v_10555 & v_8196 & v_8197 & v_8212 & ~v_8213;
assign v_10561 = v_10559 & v_10560;
assign v_10562 = v_10559 & v_8219 & v_8220 & ~v_8221 & ~v_8222;
assign v_10563 = v_10559 & v_8219 & v_8220 & v_8221;
assign v_10564 = v_10559 & v_8219 & ~v_8220 & ~v_8224;
assign v_10566 = v_10565 & v_8739;
assign v_10567 = v_10548 & v_8173 & v_8174 & v_8189 & v_8190;
assign v_10568 = v_10540 & v_8150 & v_8151 & v_8166 & v_8167;
assign v_10571 = v_10570 & v_7093;
assign v_10572 = v_10570 & ~v_7093 & v_7095 & v_7128 & ~v_7130;
assign v_10573 = v_10570 & ~v_7093 & v_7095 & v_7128 & v_7130;
assign v_10574 = v_10570 & ~v_7093 & v_7095 & ~v_7128;
assign v_10575 = v_10570 & v_7096;
assign v_10576 = v_10570 & ~v_7096;
assign v_10579 = v_10577 & v_10578;
assign v_10580 = v_10577 & v_8244;
assign v_10581 = v_13305 & v_13306;
assign v_10583 = v_10582 & ~v_7093 & ~v_7095 & v_7126;
assign v_10585 = v_10584 & v_7133 & v_7134;
assign v_10586 = v_10584 & v_7133 & ~v_7134;
assign v_10588 = v_10587 & ~v_7145;
assign v_10590 = v_10587 & v_10589;
assign v_10591 = v_10587 & v_7145 & v_7157 & ~v_7158 & v_7166;
assign v_10594 = v_10592 & v_10593;
assign v_10595 = v_10592 & v_7187 & v_7188;
assign v_10596 = v_10592 & v_7187 & ~v_7188 & v_7190;
assign v_10597 = v_10592 & v_7187 & ~v_7188 & ~v_7190 & v_7192;
assign v_10598 = v_10592 & v_7187 & ~v_7188 & ~v_7190 & ~v_7192;
assign v_10600 = v_10599 & v_8267;
assign v_10602 = v_10601 & ~v_7174 & v_7175 & v_7195;
assign v_10605 = v_10603 & v_10604;
assign v_10606 = v_10603 & v_8274;
assign v_10608 = v_10607 & v_7211 & v_7212;
assign v_10609 = v_10607 & v_7211 & ~v_7212 & v_7214;
assign v_10610 = v_10607 & v_7211 & ~v_7212 & ~v_7214 & v_7216;
assign v_10611 = v_10607 & v_7222 & v_7223;
assign v_10612 = v_10607 & v_7225 & v_7226;
assign v_10613 = v_10607 & v_7225 & ~v_7226 & v_7228;
assign v_10614 = v_10607 & v_7225 & ~v_7226 & ~v_7228 & v_7230;
assign v_10615 = v_10607 & v_8286;
assign v_10617 = v_10616 & v_8289;
assign v_10619 = v_10618 & v_7222 & ~v_7223 & v_7235 & v_7236;
assign v_10620 = v_10618 & v_7238 & v_7239;
assign v_10621 = v_10618 & v_7238 & ~v_7239 & v_7241;
assign v_10622 = v_10618 & v_7238 & ~v_7239 & ~v_7241 & v_7243;
assign v_10624 = v_10618 & v_10623;
assign v_10625 = v_13307 & v_13308;
assign v_10627 = v_10626 & v_7250 & v_7251;
assign v_10628 = v_10626 & v_7250 & ~v_7251;
assign v_10630 = v_10629 & v_8303;
assign v_10632 = v_13309 & v_13310;
assign v_10633 = v_10631 & v_7257 & v_7258;
assign v_10634 = v_10631 & v_7257 & ~v_7258 & v_7260;
assign v_10635 = v_10631 & v_7257 & ~v_7258 & ~v_7260 & v_7262;
assign v_10636 = v_10631 & v_8310;
assign v_10638 = v_13311 & v_13312;
assign v_10640 = v_10639 & v_8315;
assign v_10642 = v_10641 & v_7276 & v_7277;
assign v_10643 = v_10641 & v_7276 & ~v_7277 & v_7279;
assign v_10644 = v_10641 & v_7276 & ~v_7277 & ~v_7279 & v_7281;
assign v_10645 = v_10641 & v_7287 & v_7288;
assign v_10646 = v_10641 & v_7290 & v_7291;
assign v_10647 = v_10641 & v_7290 & ~v_7291 & v_7293;
assign v_10648 = v_10641 & v_7290 & ~v_7291 & ~v_7293 & v_7295;
assign v_10649 = v_10641 & v_8325;
assign v_10651 = v_10650 & v_8328;
assign v_10653 = v_10652 & v_7287 & ~v_7288 & v_7300 & v_7301;
assign v_10654 = v_10652 & v_7303 & v_7304;
assign v_10655 = v_10652 & v_7303 & ~v_7304 & v_7306;
assign v_10656 = v_10652 & v_7303 & ~v_7304 & ~v_7306 & v_7308;
assign v_10658 = v_10652 & v_10657;
assign v_10659 = v_13313 & v_13314;
assign v_10661 = v_10660 & v_7315 & v_7316;
assign v_10662 = v_10660 & v_7315 & ~v_7316;
assign v_10664 = v_10663 & v_8342;
assign v_10666 = v_13315 & v_13316;
assign v_10667 = v_10665 & v_7322 & v_7323;
assign v_10668 = v_10665 & v_7322 & ~v_7323 & v_7325;
assign v_10669 = v_10665 & v_7322 & ~v_7323 & ~v_7325 & v_7327;
assign v_10670 = v_10665 & v_8349;
assign v_10672 = v_13317 & v_13318;
assign v_10674 = v_10673 & v_8354;
assign v_10676 = v_10675 & v_7357;
assign v_10677 = v_10675 & ~v_7357 & v_7359 & v_7392 & ~v_7394;
assign v_10678 = v_10675 & ~v_7357 & v_7359 & v_7392 & v_7394;
assign v_10679 = v_10675 & ~v_7357 & v_7359 & ~v_7392;
assign v_10680 = v_10675 & v_7360;
assign v_10681 = v_10675 & ~v_7360;
assign v_10684 = v_10682 & v_10683;
assign v_10685 = v_10682 & v_8370;
assign v_10686 = v_13319 & v_13320;
assign v_10688 = v_10687 & ~v_7357 & ~v_7359 & v_7390;
assign v_10690 = v_10689 & v_7397 & v_7398;
assign v_10691 = v_10689 & v_7397 & ~v_7398;
assign v_10693 = v_10692 & v_7412 & v_7413;
assign v_10694 = v_10692 & v_7412 & ~v_7413 & ~v_7417;
assign v_10696 = v_10695 & v_7412 & ~v_7413 & v_7417;
assign v_10698 = v_10697 & v_7420;
assign v_10700 = v_10699 & v_7424 & v_7425;
assign v_10701 = v_10699 & v_7424 & ~v_7425 & v_7427;
assign v_10702 = v_10699 & v_8386;
assign v_10705 = v_10703 & v_10704;
assign v_10706 = v_10703 & v_8391;
assign v_10708 = v_10707 & v_7454 & ~v_7455 & ~v_7457;
assign v_10709 = v_10707 & v_7459 & ~v_7460;
assign v_10710 = v_10707 & v_7459 & v_7460;
assign v_10711 = v_10707 & v_7449;
assign v_10713 = v_10712 & v_7470 & v_7471;
assign v_10714 = v_10712 & v_7470 & ~v_7471 & ~v_7475;
assign v_10716 = v_10715 & v_7470 & ~v_7471 & v_7475;
assign v_10718 = v_10717 & v_7478;
assign v_10720 = v_10719 & v_7482 & v_7483;
assign v_10721 = v_10719 & v_7482 & ~v_7483 & v_7485;
assign v_10722 = v_10719 & v_8404;
assign v_10725 = v_10723 & v_10724;
assign v_10726 = v_10723 & v_8409;
assign v_10728 = v_6868 & v_10727;
assign v_10729 = v_7507 & v_10707;
assign v_10730 = v_7509 & v_10692;
assign v_10731 = v_7511 & v_10692;
assign v_10732 = v_7513 & v_10692;
assign v_10733 = v_7515 & v_10692;
assign v_10734 = ~v_7515 & v_10675;
assign v_10736 = ~v_7513 & v_10735;
assign v_10738 = ~v_7511 & v_10737;
assign v_10740 = ~v_7509 & v_10739;
assign v_10742 = ~v_7507 & v_10741;
assign v_10744 = ~v_6868 & v_10743;
assign v_10746 = v_10745 & ~v_7535;
assign v_10747 = v_13321 & v_13322;
assign v_10748 = v_10745 & v_7535 & v_7536 & v_7538 & v_7540;
assign v_10749 = v_13323 & v_13324;
assign v_10751 = v_10750 & v_7545 & ~v_7546 & v_7548;
assign v_10752 = v_10750 & v_7555 & ~v_7556 & ~v_7558;
assign v_10753 = v_10750 & v_7560 & ~v_7561;
assign v_10754 = v_10750 & v_7560 & v_7561;
assign v_10755 = v_10750 & v_7550;
assign v_10757 = v_10756 & v_8441;
assign v_10759 = v_10758 & v_8444;
assign v_10760 = v_10750 & v_7545 & v_7546;
assign v_10761 = v_10745 & v_8447;
assign v_10763 = v_10762 & ~v_7571;
assign v_10764 = v_10762 & v_7576 & v_7577;
assign v_10765 = v_10762 & v_7576 & ~v_7577 & ~v_7581;
assign v_10767 = v_10766 & v_7576 & ~v_7577 & v_7581;
assign v_10769 = v_10768 & v_7584;
assign v_10771 = v_10770 & v_7571 & v_7588 & v_7589 & ~v_7590;
assign v_10773 = v_10770 & v_10772;
assign v_10774 = v_10770 & v_7616 & v_7617;
assign v_10775 = v_10770 & v_7616 & ~v_7617;
assign v_10777 = v_10776 & v_7629 & v_7630;
assign v_10778 = v_10776 & v_7629 & ~v_7630;
assign v_10780 = v_10779 & v_7611 & v_7624 & v_7637;
assign v_10781 = v_13325 & v_13326;
assign v_10782 = v_10770 & v_7645 & v_7646;
assign v_10783 = v_10770 & v_7645 & ~v_7646 & ~v_7650;
assign v_10785 = v_10784 & v_7645 & ~v_7646 & v_7650;
assign v_10787 = v_10786 & v_7653;
assign v_10789 = v_10788 & v_8468;
assign v_10791 = v_10790 & v_7664 & ~v_7665 & v_7683;
assign v_10792 = v_10790 & v_7664 & ~v_7665 & ~v_7683;
assign v_10793 = v_10790 & ~v_7666;
assign v_10794 = v_10790 & v_7674 & ~v_7675;
assign v_10795 = v_10790 & v_8475;
assign v_10797 = v_10796 & v_7664 & v_7665 & v_7680 & ~v_7681;
assign v_10799 = v_10798 & v_7687 & ~v_7688 & v_7706;
assign v_10800 = v_10798 & v_7687 & ~v_7688 & ~v_7706;
assign v_10801 = v_10798 & ~v_7689;
assign v_10802 = v_10798 & v_7697 & ~v_7698;
assign v_10803 = v_10798 & v_8484;
assign v_10805 = v_10804 & v_7687 & v_7688 & v_7703 & ~v_7704;
assign v_10807 = v_10806 & v_7710 & ~v_7711 & v_7729;
assign v_10808 = v_10806 & ~v_7712;
assign v_10809 = v_10806 & v_7720 & ~v_7721;
assign v_10810 = v_10806 & v_8492;
assign v_10812 = v_10811 & v_7710 & v_7711 & v_7726 & v_7727;
assign v_10813 = v_10806 & v_7710 & ~v_7711 & ~v_7729;
assign v_10814 = v_10811 & v_7710 & v_7711 & v_7726 & ~v_7727;
assign v_10817 = v_10815 & v_10816;
assign v_10818 = v_10815 & v_7733 & v_7734 & ~v_7735 & ~v_7736;
assign v_10819 = v_10815 & v_7733 & v_7734 & v_7735;
assign v_10820 = v_10815 & v_7733 & ~v_7734 & ~v_7738;
assign v_10822 = v_10821 & v_8505;
assign v_10823 = v_10804 & v_7687 & v_7688 & v_7703 & v_7704;
assign v_10824 = v_10796 & v_7664 & v_7665 & v_7680 & v_7681;
assign v_10826 = v_10825 & v_7745 & ~v_7746 & v_7764;
assign v_10827 = v_10825 & v_7745 & ~v_7746 & ~v_7764;
assign v_10828 = v_10825 & ~v_7747;
assign v_10829 = v_10825 & v_7755 & ~v_7756;
assign v_10830 = v_10825 & v_8514;
assign v_10832 = v_10831 & v_7745 & v_7746 & v_7761 & ~v_7762;
assign v_10834 = v_10833 & v_7768 & ~v_7769 & v_7787;
assign v_10835 = v_10833 & v_7768 & ~v_7769 & ~v_7787;
assign v_10836 = v_10833 & ~v_7770;
assign v_10837 = v_10833 & v_7778 & ~v_7779;
assign v_10838 = v_10833 & v_8523;
assign v_10840 = v_10839 & v_7768 & v_7769 & v_7784 & ~v_7785;
assign v_10842 = v_10841 & v_7791 & ~v_7792 & v_7810;
assign v_10843 = v_10841 & ~v_7793;
assign v_10844 = v_10841 & v_7801 & ~v_7802;
assign v_10845 = v_10841 & v_8531;
assign v_10847 = v_10846 & v_7791 & v_7792 & v_7807 & v_7808;
assign v_10848 = v_10841 & v_7791 & ~v_7792 & ~v_7810;
assign v_10849 = v_10846 & v_7791 & v_7792 & v_7807 & ~v_7808;
assign v_10852 = v_10850 & v_10851;
assign v_10853 = v_10850 & v_7814 & v_7815 & ~v_7816 & ~v_7817;
assign v_10854 = v_10850 & v_7814 & v_7815 & v_7816;
assign v_10855 = v_10850 & v_7814 & ~v_7815 & ~v_7819;
assign v_10857 = v_10856 & v_8544;
assign v_10858 = v_10839 & v_7768 & v_7769 & v_7784 & v_7785;
assign v_10859 = v_10831 & v_7745 & v_7746 & v_7761 & v_7762;
assign v_10861 = v_10860 & v_7826 & ~v_7827 & v_7845;
assign v_10862 = v_10860 & v_7826 & ~v_7827 & ~v_7845;
assign v_10863 = v_10860 & ~v_7828;
assign v_10864 = v_10860 & v_7836 & ~v_7837;
assign v_10865 = v_10860 & v_8553;
assign v_10867 = v_10866 & v_7826 & v_7827 & v_7842 & ~v_7843;
assign v_10869 = v_10868 & v_7849 & ~v_7850 & v_7868;
assign v_10870 = v_10868 & v_7849 & ~v_7850 & ~v_7868;
assign v_10871 = v_10868 & ~v_7851;
assign v_10872 = v_10868 & v_7859 & ~v_7860;
assign v_10873 = v_10868 & v_8562;
assign v_10875 = v_10874 & v_7849 & v_7850 & v_7865 & ~v_7866;
assign v_10877 = v_10876 & v_7872 & ~v_7873 & v_7891;
assign v_10878 = v_10876 & ~v_7874;
assign v_10879 = v_10876 & v_7882 & ~v_7883;
assign v_10880 = v_10876 & v_8570;
assign v_10882 = v_10881 & v_7872 & v_7873 & v_7888 & v_7889;
assign v_10883 = v_10876 & v_7872 & ~v_7873 & ~v_7891;
assign v_10884 = v_10881 & v_7872 & v_7873 & v_7888 & ~v_7889;
assign v_10887 = v_10885 & v_10886;
assign v_10888 = v_10885 & v_7895 & v_7896 & ~v_7897 & ~v_7898;
assign v_10889 = v_10885 & v_7895 & v_7896 & v_7897;
assign v_10890 = v_10885 & v_7895 & ~v_7896 & ~v_7900;
assign v_10892 = v_10891 & v_8583;
assign v_10893 = v_10874 & v_7849 & v_7850 & v_7865 & v_7866;
assign v_10894 = v_10866 & v_7826 & v_7827 & v_7842 & v_7843;
assign v_10896 = v_10895 & v_7907 & ~v_7908 & v_7926;
assign v_10897 = v_10895 & v_7907 & ~v_7908 & ~v_7926;
assign v_10898 = v_10895 & ~v_7909;
assign v_10899 = v_10895 & v_7917 & ~v_7918;
assign v_10900 = v_10895 & v_8592;
assign v_10902 = v_10901 & v_7907 & v_7908 & v_7923 & ~v_7924;
assign v_10904 = v_10903 & v_7930 & ~v_7931 & v_7949;
assign v_10905 = v_10903 & v_7930 & ~v_7931 & ~v_7949;
assign v_10906 = v_10903 & ~v_7932;
assign v_10907 = v_10903 & v_7940 & ~v_7941;
assign v_10908 = v_10903 & v_8601;
assign v_10910 = v_10909 & v_7930 & v_7931 & v_7946 & ~v_7947;
assign v_10912 = v_10911 & v_7953 & ~v_7954 & v_7972;
assign v_10913 = v_10911 & ~v_7955;
assign v_10914 = v_10911 & v_7963 & ~v_7964;
assign v_10915 = v_10911 & v_8609;
assign v_10917 = v_10916 & v_7953 & v_7954 & v_7969 & v_7970;
assign v_10918 = v_10911 & v_7953 & ~v_7954 & ~v_7972;
assign v_10919 = v_10916 & v_7953 & v_7954 & v_7969 & ~v_7970;
assign v_10922 = v_10920 & v_10921;
assign v_10923 = v_10920 & v_7976 & v_7977 & ~v_7978 & ~v_7979;
assign v_10924 = v_10920 & v_7976 & v_7977 & v_7978;
assign v_10925 = v_10920 & v_7976 & ~v_7977 & ~v_7981;
assign v_10927 = v_10926 & v_8622;
assign v_10928 = v_10909 & v_7930 & v_7931 & v_7946 & v_7947;
assign v_10929 = v_10901 & v_7907 & v_7908 & v_7923 & v_7924;
assign v_10931 = v_10930 & v_7988 & ~v_7989 & v_8007;
assign v_10932 = v_10930 & v_7988 & ~v_7989 & ~v_8007;
assign v_10933 = v_10930 & ~v_7990;
assign v_10934 = v_10930 & v_7998 & ~v_7999;
assign v_10935 = v_10930 & v_8631;
assign v_10937 = v_10936 & v_7988 & v_7989 & v_8004 & ~v_8005;
assign v_10939 = v_10938 & v_8011 & ~v_8012 & v_8030;
assign v_10940 = v_10938 & v_8011 & ~v_8012 & ~v_8030;
assign v_10941 = v_10938 & ~v_8013;
assign v_10942 = v_10938 & v_8021 & ~v_8022;
assign v_10943 = v_10938 & v_8640;
assign v_10945 = v_10944 & v_8011 & v_8012 & v_8027 & ~v_8028;
assign v_10947 = v_10946 & v_8034 & ~v_8035 & v_8053;
assign v_10948 = v_10946 & ~v_8036;
assign v_10949 = v_10946 & v_8044 & ~v_8045;
assign v_10950 = v_10946 & v_8648;
assign v_10952 = v_10951 & v_8034 & v_8035 & v_8050 & v_8051;
assign v_10953 = v_10946 & v_8034 & ~v_8035 & ~v_8053;
assign v_10954 = v_10951 & v_8034 & v_8035 & v_8050 & ~v_8051;
assign v_10957 = v_10955 & v_10956;
assign v_10958 = v_10955 & v_8057 & v_8058 & ~v_8059 & ~v_8060;
assign v_10959 = v_10955 & v_8057 & v_8058 & v_8059;
assign v_10960 = v_10955 & v_8057 & ~v_8058 & ~v_8062;
assign v_10962 = v_10961 & v_8661;
assign v_10963 = v_10944 & v_8011 & v_8012 & v_8027 & v_8028;
assign v_10964 = v_10936 & v_7988 & v_7989 & v_8004 & v_8005;
assign v_10966 = v_10965 & v_8069 & ~v_8070 & v_8088;
assign v_10967 = v_10965 & v_8069 & ~v_8070 & ~v_8088;
assign v_10968 = v_10965 & ~v_8071;
assign v_10969 = v_10965 & v_8079 & ~v_8080;
assign v_10970 = v_10965 & v_8670;
assign v_10972 = v_10971 & v_8069 & v_8070 & v_8085 & ~v_8086;
assign v_10974 = v_10973 & v_8092 & ~v_8093 & v_8111;
assign v_10975 = v_10973 & v_8092 & ~v_8093 & ~v_8111;
assign v_10976 = v_10973 & ~v_8094;
assign v_10977 = v_10973 & v_8102 & ~v_8103;
assign v_10978 = v_10973 & v_8679;
assign v_10980 = v_10979 & v_8092 & v_8093 & v_8108 & ~v_8109;
assign v_10982 = v_10981 & v_8115 & ~v_8116 & v_8134;
assign v_10983 = v_10981 & ~v_8117;
assign v_10984 = v_10981 & v_8125 & ~v_8126;
assign v_10985 = v_10981 & v_8687;
assign v_10987 = v_10986 & v_8115 & v_8116 & v_8131 & v_8132;
assign v_10988 = v_10981 & v_8115 & ~v_8116 & ~v_8134;
assign v_10989 = v_10986 & v_8115 & v_8116 & v_8131 & ~v_8132;
assign v_10992 = v_10990 & v_10991;
assign v_10993 = v_10990 & v_8138 & v_8139 & ~v_8140 & ~v_8141;
assign v_10994 = v_10990 & v_8138 & v_8139 & v_8140;
assign v_10995 = v_10990 & v_8138 & ~v_8139 & ~v_8143;
assign v_10997 = v_10996 & v_8700;
assign v_10998 = v_10979 & v_8092 & v_8093 & v_8108 & v_8109;
assign v_10999 = v_10971 & v_8069 & v_8070 & v_8085 & v_8086;
assign v_11001 = v_11000 & v_8150 & ~v_8151 & v_8169;
assign v_11002 = v_11000 & v_8150 & ~v_8151 & ~v_8169;
assign v_11003 = v_11000 & ~v_8152;
assign v_11004 = v_11000 & v_8160 & ~v_8161;
assign v_11005 = v_11000 & v_8709;
assign v_11007 = v_11006 & v_8150 & v_8151 & v_8166 & ~v_8167;
assign v_11009 = v_11008 & v_8173 & ~v_8174 & v_8192;
assign v_11010 = v_11008 & v_8173 & ~v_8174 & ~v_8192;
assign v_11011 = v_11008 & ~v_8175;
assign v_11012 = v_11008 & v_8183 & ~v_8184;
assign v_11013 = v_11008 & v_8718;
assign v_11015 = v_11014 & v_8173 & v_8174 & v_8189 & ~v_8190;
assign v_11017 = v_11016 & v_8196 & ~v_8197 & v_8215;
assign v_11018 = v_11016 & ~v_8198;
assign v_11019 = v_11016 & v_8206 & ~v_8207;
assign v_11020 = v_11016 & v_8726;
assign v_11022 = v_11021 & v_8196 & v_8197 & v_8212 & v_8213;
assign v_11023 = v_11016 & v_8196 & ~v_8197 & ~v_8215;
assign v_11024 = v_11021 & v_8196 & v_8197 & v_8212 & ~v_8213;
assign v_11027 = v_11025 & v_11026;
assign v_11028 = v_11025 & v_8219 & v_8220 & ~v_8221 & ~v_8222;
assign v_11029 = v_11025 & v_8219 & v_8220 & v_8221;
assign v_11030 = v_11025 & v_8219 & ~v_8220 & ~v_8224;
assign v_11032 = v_11031 & v_8739;
assign v_11033 = v_11014 & v_8173 & v_8174 & v_8189 & v_8190;
assign v_11034 = v_11006 & v_8150 & v_8151 & v_8166 & v_8167;
assign v_11036 = v_6873 & v_7093;
assign v_11037 = v_6873 & ~v_7093 & v_7095 & v_7128 & ~v_7130;
assign v_11038 = v_6873 & ~v_7093 & v_7095 & v_7128 & v_7130;
assign v_11039 = v_6873 & ~v_7093 & v_7095 & ~v_7128;
assign v_11040 = v_6873 & v_7096;
assign v_11041 = v_6873 & ~v_7096;
assign v_11044 = v_11042 & v_11043;
assign v_11045 = v_11042 & v_8244;
assign v_11046 = v_13327 & v_13328;
assign v_11048 = v_11047 & ~v_7093 & ~v_7095 & v_7126;
assign v_11050 = v_11049 & v_7133 & v_7134;
assign v_11051 = v_11049 & v_7133 & ~v_7134;
assign v_11053 = v_11052 & ~v_7145;
assign v_11055 = v_11052 & v_11054;
assign v_11056 = v_11052 & v_7145 & v_7157 & ~v_7158 & v_7166;
assign v_11059 = v_11057 & v_11058;
assign v_11060 = v_11057 & v_7187 & v_7188;
assign v_11061 = v_11057 & v_7187 & ~v_7188 & v_7190;
assign v_11062 = v_11057 & v_7187 & ~v_7188 & ~v_7190 & v_7192;
assign v_11063 = v_11057 & v_7187 & ~v_7188 & ~v_7190 & ~v_7192;
assign v_11065 = v_11064 & v_8267;
assign v_11067 = v_11066 & ~v_7174 & v_7175 & v_7195;
assign v_11070 = v_11068 & v_11069;
assign v_11071 = v_11068 & v_8274;
assign v_11073 = v_11072 & v_7211 & v_7212;
assign v_11074 = v_11072 & v_7211 & ~v_7212 & v_7214;
assign v_11075 = v_11072 & v_7211 & ~v_7212 & ~v_7214 & v_7216;
assign v_11076 = v_11072 & v_7222 & v_7223;
assign v_11077 = v_11072 & v_7225 & v_7226;
assign v_11078 = v_11072 & v_7225 & ~v_7226 & v_7228;
assign v_11079 = v_11072 & v_7225 & ~v_7226 & ~v_7228 & v_7230;
assign v_11080 = v_11072 & v_8286;
assign v_11082 = v_11081 & v_8289;
assign v_11084 = v_11083 & v_7222 & ~v_7223 & v_7235 & v_7236;
assign v_11085 = v_11083 & v_7238 & v_7239;
assign v_11086 = v_11083 & v_7238 & ~v_7239 & v_7241;
assign v_11087 = v_11083 & v_7238 & ~v_7239 & ~v_7241 & v_7243;
assign v_11089 = v_11083 & v_11088;
assign v_11090 = v_13329 & v_13330;
assign v_11092 = v_11091 & v_7250 & v_7251;
assign v_11093 = v_11091 & v_7250 & ~v_7251;
assign v_11095 = v_11094 & v_8303;
assign v_11097 = v_13331 & v_13332;
assign v_11098 = v_11096 & v_7257 & v_7258;
assign v_11099 = v_11096 & v_7257 & ~v_7258 & v_7260;
assign v_11100 = v_11096 & v_7257 & ~v_7258 & ~v_7260 & v_7262;
assign v_11101 = v_11096 & v_8310;
assign v_11103 = v_13333 & v_13334;
assign v_11105 = v_11104 & v_8315;
assign v_11107 = v_11106 & v_7276 & v_7277;
assign v_11108 = v_11106 & v_7276 & ~v_7277 & v_7279;
assign v_11109 = v_11106 & v_7276 & ~v_7277 & ~v_7279 & v_7281;
assign v_11110 = v_11106 & v_7287 & v_7288;
assign v_11111 = v_11106 & v_7290 & v_7291;
assign v_11112 = v_11106 & v_7290 & ~v_7291 & v_7293;
assign v_11113 = v_11106 & v_7290 & ~v_7291 & ~v_7293 & v_7295;
assign v_11114 = v_11106 & v_8325;
assign v_11116 = v_11115 & v_8328;
assign v_11118 = v_11117 & v_7287 & ~v_7288 & v_7300 & v_7301;
assign v_11119 = v_11117 & v_7303 & v_7304;
assign v_11120 = v_11117 & v_7303 & ~v_7304 & v_7306;
assign v_11121 = v_11117 & v_7303 & ~v_7304 & ~v_7306 & v_7308;
assign v_11123 = v_11117 & v_11122;
assign v_11124 = v_13335 & v_13336;
assign v_11126 = v_11125 & v_7315 & v_7316;
assign v_11127 = v_11125 & v_7315 & ~v_7316;
assign v_11129 = v_11128 & v_8342;
assign v_11131 = v_13337 & v_13338;
assign v_11132 = v_11130 & v_7322 & v_7323;
assign v_11133 = v_11130 & v_7322 & ~v_7323 & v_7325;
assign v_11134 = v_11130 & v_7322 & ~v_7323 & ~v_7325 & v_7327;
assign v_11135 = v_11130 & v_8349;
assign v_11137 = v_13339 & v_13340;
assign v_11139 = v_11138 & v_8354;
assign v_11141 = v_11140 & v_7357;
assign v_11142 = v_11140 & ~v_7357 & v_7359 & v_7392 & ~v_7394;
assign v_11143 = v_11140 & ~v_7357 & v_7359 & v_7392 & v_7394;
assign v_11144 = v_11140 & ~v_7357 & v_7359 & ~v_7392;
assign v_11145 = v_11140 & v_7360;
assign v_11146 = v_11140 & ~v_7360;
assign v_11149 = v_11147 & v_11148;
assign v_11150 = v_11147 & v_8370;
assign v_11151 = v_13341 & v_13342;
assign v_11153 = v_11152 & ~v_7357 & ~v_7359 & v_7390;
assign v_11155 = v_11154 & v_7397 & v_7398;
assign v_11156 = v_11154 & v_7397 & ~v_7398;
assign v_11158 = v_11157 & v_7412 & v_7413;
assign v_11159 = v_11157 & v_7412 & ~v_7413 & ~v_7417;
assign v_11161 = v_11160 & v_7412 & ~v_7413 & v_7417;
assign v_11163 = v_11162 & v_7420;
assign v_11165 = v_11164 & v_7424 & v_7425;
assign v_11166 = v_11164 & v_7424 & ~v_7425 & v_7427;
assign v_11167 = v_11164 & v_8386;
assign v_11170 = v_11168 & v_11169;
assign v_11171 = v_11168 & v_8391;
assign v_11173 = v_11172 & v_7454 & ~v_7455 & ~v_7457;
assign v_11174 = v_11172 & v_7459 & ~v_7460;
assign v_11175 = v_11172 & v_7459 & v_7460;
assign v_11176 = v_11172 & v_7449;
assign v_11178 = v_11177 & v_7470 & v_7471;
assign v_11179 = v_11177 & v_7470 & ~v_7471 & ~v_7475;
assign v_11181 = v_11180 & v_7470 & ~v_7471 & v_7475;
assign v_11183 = v_11182 & v_7478;
assign v_11185 = v_11184 & v_7482 & v_7483;
assign v_11186 = v_11184 & v_7482 & ~v_7483 & v_7485;
assign v_11187 = v_11184 & v_8404;
assign v_11190 = v_11188 & v_11189;
assign v_11191 = v_11188 & v_8409;
assign v_11193 = v_6868 & v_11192;
assign v_11194 = v_7507 & v_11172;
assign v_11195 = v_7509 & v_11157;
assign v_11196 = v_7511 & v_11157;
assign v_11197 = v_7513 & v_11157;
assign v_11198 = v_7515 & v_11157;
assign v_11199 = ~v_7515 & v_11140;
assign v_11201 = ~v_7513 & v_11200;
assign v_11203 = ~v_7511 & v_11202;
assign v_11205 = ~v_7509 & v_11204;
assign v_11207 = ~v_7507 & v_11206;
assign v_11209 = ~v_6868 & v_11208;
assign v_11211 = v_11210 & ~v_7535;
assign v_11212 = v_13343 & v_13344;
assign v_11213 = v_11210 & v_7535 & v_7536 & v_7538 & v_7540;
assign v_11214 = v_13345 & v_13346;
assign v_11216 = v_11215 & v_7545 & ~v_7546 & v_7548;
assign v_11217 = v_11215 & v_7555 & ~v_7556 & ~v_7558;
assign v_11218 = v_11215 & v_7560 & ~v_7561;
assign v_11219 = v_11215 & v_7560 & v_7561;
assign v_11220 = v_11215 & v_7550;
assign v_11222 = v_11221 & v_8441;
assign v_11224 = v_11223 & v_8444;
assign v_11225 = v_11215 & v_7545 & v_7546;
assign v_11226 = v_11210 & v_8447;
assign v_11228 = v_11227 & ~v_7571;
assign v_11229 = v_11227 & v_7576 & v_7577;
assign v_11230 = v_11227 & v_7576 & ~v_7577 & ~v_7581;
assign v_11232 = v_11231 & v_7576 & ~v_7577 & v_7581;
assign v_11234 = v_11233 & v_7584;
assign v_11236 = v_11235 & v_7571 & v_7588 & v_7589 & ~v_7590;
assign v_11238 = v_11235 & v_11237;
assign v_11239 = v_11235 & v_7616 & v_7617;
assign v_11240 = v_11235 & v_7616 & ~v_7617;
assign v_11242 = v_11241 & v_7629 & v_7630;
assign v_11243 = v_11241 & v_7629 & ~v_7630;
assign v_11245 = v_11244 & v_7611 & v_7624 & v_7637;
assign v_11246 = v_13347 & v_13348;
assign v_11247 = v_11235 & v_7645 & v_7646;
assign v_11248 = v_11235 & v_7645 & ~v_7646 & ~v_7650;
assign v_11250 = v_11249 & v_7645 & ~v_7646 & v_7650;
assign v_11252 = v_11251 & v_7653;
assign v_11254 = v_11253 & v_8468;
assign v_11256 = v_11255 & v_7664 & ~v_7665 & v_7683;
assign v_11257 = v_11255 & v_7664 & ~v_7665 & ~v_7683;
assign v_11258 = v_11255 & ~v_7666;
assign v_11259 = v_11255 & v_7674 & ~v_7675;
assign v_11260 = v_11255 & v_8475;
assign v_11262 = v_11261 & v_7664 & v_7665 & v_7680 & ~v_7681;
assign v_11264 = v_11263 & v_7687 & ~v_7688 & v_7706;
assign v_11265 = v_11263 & v_7687 & ~v_7688 & ~v_7706;
assign v_11266 = v_11263 & ~v_7689;
assign v_11267 = v_11263 & v_7697 & ~v_7698;
assign v_11268 = v_11263 & v_8484;
assign v_11270 = v_11269 & v_7687 & v_7688 & v_7703 & ~v_7704;
assign v_11272 = v_11271 & v_7710 & ~v_7711 & v_7729;
assign v_11273 = v_11271 & ~v_7712;
assign v_11274 = v_11271 & v_7720 & ~v_7721;
assign v_11275 = v_11271 & v_8492;
assign v_11277 = v_11276 & v_7710 & v_7711 & v_7726 & v_7727;
assign v_11278 = v_11271 & v_7710 & ~v_7711 & ~v_7729;
assign v_11279 = v_11276 & v_7710 & v_7711 & v_7726 & ~v_7727;
assign v_11282 = v_11280 & v_11281;
assign v_11283 = v_11280 & v_7733 & v_7734 & ~v_7735 & ~v_7736;
assign v_11284 = v_11280 & v_7733 & v_7734 & v_7735;
assign v_11285 = v_11280 & v_7733 & ~v_7734 & ~v_7738;
assign v_11287 = v_11286 & v_8505;
assign v_11288 = v_11269 & v_7687 & v_7688 & v_7703 & v_7704;
assign v_11289 = v_11261 & v_7664 & v_7665 & v_7680 & v_7681;
assign v_11291 = v_11290 & v_7745 & ~v_7746 & v_7764;
assign v_11292 = v_11290 & v_7745 & ~v_7746 & ~v_7764;
assign v_11293 = v_11290 & ~v_7747;
assign v_11294 = v_11290 & v_7755 & ~v_7756;
assign v_11295 = v_11290 & v_8514;
assign v_11297 = v_11296 & v_7745 & v_7746 & v_7761 & ~v_7762;
assign v_11299 = v_11298 & v_7768 & ~v_7769 & v_7787;
assign v_11300 = v_11298 & v_7768 & ~v_7769 & ~v_7787;
assign v_11301 = v_11298 & ~v_7770;
assign v_11302 = v_11298 & v_7778 & ~v_7779;
assign v_11303 = v_11298 & v_8523;
assign v_11305 = v_11304 & v_7768 & v_7769 & v_7784 & ~v_7785;
assign v_11307 = v_11306 & v_7791 & ~v_7792 & v_7810;
assign v_11308 = v_11306 & ~v_7793;
assign v_11309 = v_11306 & v_7801 & ~v_7802;
assign v_11310 = v_11306 & v_8531;
assign v_11312 = v_11311 & v_7791 & v_7792 & v_7807 & v_7808;
assign v_11313 = v_11306 & v_7791 & ~v_7792 & ~v_7810;
assign v_11314 = v_11311 & v_7791 & v_7792 & v_7807 & ~v_7808;
assign v_11317 = v_11315 & v_11316;
assign v_11318 = v_11315 & v_7814 & v_7815 & ~v_7816 & ~v_7817;
assign v_11319 = v_11315 & v_7814 & v_7815 & v_7816;
assign v_11320 = v_11315 & v_7814 & ~v_7815 & ~v_7819;
assign v_11322 = v_11321 & v_8544;
assign v_11323 = v_11304 & v_7768 & v_7769 & v_7784 & v_7785;
assign v_11324 = v_11296 & v_7745 & v_7746 & v_7761 & v_7762;
assign v_11326 = v_11325 & v_7826 & ~v_7827 & v_7845;
assign v_11327 = v_11325 & v_7826 & ~v_7827 & ~v_7845;
assign v_11328 = v_11325 & ~v_7828;
assign v_11329 = v_11325 & v_7836 & ~v_7837;
assign v_11330 = v_11325 & v_8553;
assign v_11332 = v_11331 & v_7826 & v_7827 & v_7842 & ~v_7843;
assign v_11334 = v_11333 & v_7849 & ~v_7850 & v_7868;
assign v_11335 = v_11333 & v_7849 & ~v_7850 & ~v_7868;
assign v_11336 = v_11333 & ~v_7851;
assign v_11337 = v_11333 & v_7859 & ~v_7860;
assign v_11338 = v_11333 & v_8562;
assign v_11340 = v_11339 & v_7849 & v_7850 & v_7865 & ~v_7866;
assign v_11342 = v_11341 & v_7872 & ~v_7873 & v_7891;
assign v_11343 = v_11341 & ~v_7874;
assign v_11344 = v_11341 & v_7882 & ~v_7883;
assign v_11345 = v_11341 & v_8570;
assign v_11347 = v_11346 & v_7872 & v_7873 & v_7888 & v_7889;
assign v_11348 = v_11341 & v_7872 & ~v_7873 & ~v_7891;
assign v_11349 = v_11346 & v_7872 & v_7873 & v_7888 & ~v_7889;
assign v_11352 = v_11350 & v_11351;
assign v_11353 = v_11350 & v_7895 & v_7896 & ~v_7897 & ~v_7898;
assign v_11354 = v_11350 & v_7895 & v_7896 & v_7897;
assign v_11355 = v_11350 & v_7895 & ~v_7896 & ~v_7900;
assign v_11357 = v_11356 & v_8583;
assign v_11358 = v_11339 & v_7849 & v_7850 & v_7865 & v_7866;
assign v_11359 = v_11331 & v_7826 & v_7827 & v_7842 & v_7843;
assign v_11361 = v_11360 & v_7907 & ~v_7908 & v_7926;
assign v_11362 = v_11360 & v_7907 & ~v_7908 & ~v_7926;
assign v_11363 = v_11360 & ~v_7909;
assign v_11364 = v_11360 & v_7917 & ~v_7918;
assign v_11365 = v_11360 & v_8592;
assign v_11367 = v_11366 & v_7907 & v_7908 & v_7923 & ~v_7924;
assign v_11369 = v_11368 & v_7930 & ~v_7931 & v_7949;
assign v_11370 = v_11368 & v_7930 & ~v_7931 & ~v_7949;
assign v_11371 = v_11368 & ~v_7932;
assign v_11372 = v_11368 & v_7940 & ~v_7941;
assign v_11373 = v_11368 & v_8601;
assign v_11375 = v_11374 & v_7930 & v_7931 & v_7946 & ~v_7947;
assign v_11377 = v_11376 & v_7953 & ~v_7954 & v_7972;
assign v_11378 = v_11376 & ~v_7955;
assign v_11379 = v_11376 & v_7963 & ~v_7964;
assign v_11380 = v_11376 & v_8609;
assign v_11382 = v_11381 & v_7953 & v_7954 & v_7969 & v_7970;
assign v_11383 = v_11376 & v_7953 & ~v_7954 & ~v_7972;
assign v_11384 = v_11381 & v_7953 & v_7954 & v_7969 & ~v_7970;
assign v_11387 = v_11385 & v_11386;
assign v_11388 = v_11385 & v_7976 & v_7977 & ~v_7978 & ~v_7979;
assign v_11389 = v_11385 & v_7976 & v_7977 & v_7978;
assign v_11390 = v_11385 & v_7976 & ~v_7977 & ~v_7981;
assign v_11392 = v_11391 & v_8622;
assign v_11393 = v_11374 & v_7930 & v_7931 & v_7946 & v_7947;
assign v_11394 = v_11366 & v_7907 & v_7908 & v_7923 & v_7924;
assign v_11396 = v_11395 & v_7988 & ~v_7989 & v_8007;
assign v_11397 = v_11395 & v_7988 & ~v_7989 & ~v_8007;
assign v_11398 = v_11395 & ~v_7990;
assign v_11399 = v_11395 & v_7998 & ~v_7999;
assign v_11400 = v_11395 & v_8631;
assign v_11402 = v_11401 & v_7988 & v_7989 & v_8004 & ~v_8005;
assign v_11404 = v_11403 & v_8011 & ~v_8012 & v_8030;
assign v_11405 = v_11403 & v_8011 & ~v_8012 & ~v_8030;
assign v_11406 = v_11403 & ~v_8013;
assign v_11407 = v_11403 & v_8021 & ~v_8022;
assign v_11408 = v_11403 & v_8640;
assign v_11410 = v_11409 & v_8011 & v_8012 & v_8027 & ~v_8028;
assign v_11412 = v_11411 & v_8034 & ~v_8035 & v_8053;
assign v_11413 = v_11411 & ~v_8036;
assign v_11414 = v_11411 & v_8044 & ~v_8045;
assign v_11415 = v_11411 & v_8648;
assign v_11417 = v_11416 & v_8034 & v_8035 & v_8050 & v_8051;
assign v_11418 = v_11411 & v_8034 & ~v_8035 & ~v_8053;
assign v_11419 = v_11416 & v_8034 & v_8035 & v_8050 & ~v_8051;
assign v_11422 = v_11420 & v_11421;
assign v_11423 = v_11420 & v_8057 & v_8058 & ~v_8059 & ~v_8060;
assign v_11424 = v_11420 & v_8057 & v_8058 & v_8059;
assign v_11425 = v_11420 & v_8057 & ~v_8058 & ~v_8062;
assign v_11427 = v_11426 & v_8661;
assign v_11428 = v_11409 & v_8011 & v_8012 & v_8027 & v_8028;
assign v_11429 = v_11401 & v_7988 & v_7989 & v_8004 & v_8005;
assign v_11431 = v_11430 & v_8069 & ~v_8070 & v_8088;
assign v_11432 = v_11430 & v_8069 & ~v_8070 & ~v_8088;
assign v_11433 = v_11430 & ~v_8071;
assign v_11434 = v_11430 & v_8079 & ~v_8080;
assign v_11435 = v_11430 & v_8670;
assign v_11437 = v_11436 & v_8069 & v_8070 & v_8085 & ~v_8086;
assign v_11439 = v_11438 & v_8092 & ~v_8093 & v_8111;
assign v_11440 = v_11438 & v_8092 & ~v_8093 & ~v_8111;
assign v_11441 = v_11438 & ~v_8094;
assign v_11442 = v_11438 & v_8102 & ~v_8103;
assign v_11443 = v_11438 & v_8679;
assign v_11445 = v_11444 & v_8092 & v_8093 & v_8108 & ~v_8109;
assign v_11447 = v_11446 & v_8115 & ~v_8116 & v_8134;
assign v_11448 = v_11446 & ~v_8117;
assign v_11449 = v_11446 & v_8125 & ~v_8126;
assign v_11450 = v_11446 & v_8687;
assign v_11452 = v_11451 & v_8115 & v_8116 & v_8131 & v_8132;
assign v_11453 = v_11446 & v_8115 & ~v_8116 & ~v_8134;
assign v_11454 = v_11451 & v_8115 & v_8116 & v_8131 & ~v_8132;
assign v_11457 = v_11455 & v_11456;
assign v_11458 = v_11455 & v_8138 & v_8139 & ~v_8140 & ~v_8141;
assign v_11459 = v_11455 & v_8138 & v_8139 & v_8140;
assign v_11460 = v_11455 & v_8138 & ~v_8139 & ~v_8143;
assign v_11462 = v_11461 & v_8700;
assign v_11463 = v_11444 & v_8092 & v_8093 & v_8108 & v_8109;
assign v_11464 = v_11436 & v_8069 & v_8070 & v_8085 & v_8086;
assign v_11466 = v_11465 & v_8150 & ~v_8151 & v_8169;
assign v_11467 = v_11465 & v_8150 & ~v_8151 & ~v_8169;
assign v_11468 = v_11465 & ~v_8152;
assign v_11469 = v_11465 & v_8160 & ~v_8161;
assign v_11470 = v_11465 & v_8709;
assign v_11472 = v_11471 & v_8150 & v_8151 & v_8166 & ~v_8167;
assign v_11474 = v_11473 & v_8173 & ~v_8174 & v_8192;
assign v_11475 = v_11473 & v_8173 & ~v_8174 & ~v_8192;
assign v_11476 = v_11473 & ~v_8175;
assign v_11477 = v_11473 & v_8183 & ~v_8184;
assign v_11478 = v_11473 & v_8718;
assign v_11480 = v_11479 & v_8173 & v_8174 & v_8189 & ~v_8190;
assign v_11482 = v_11481 & v_8196 & ~v_8197 & v_8215;
assign v_11483 = v_11481 & ~v_8198;
assign v_11484 = v_11481 & v_8206 & ~v_8207;
assign v_11485 = v_11481 & v_8726;
assign v_11487 = v_11486 & v_8196 & v_8197 & v_8212 & v_8213;
assign v_11488 = v_11481 & v_8196 & ~v_8197 & ~v_8215;
assign v_11489 = v_11486 & v_8196 & v_8197 & v_8212 & ~v_8213;
assign v_11492 = v_11490 & v_11491;
assign v_11493 = v_11490 & v_8219 & v_8220 & ~v_8221 & ~v_8222;
assign v_11494 = v_11490 & v_8219 & v_8220 & v_8221;
assign v_11495 = v_11490 & v_8219 & ~v_8220 & ~v_8224;
assign v_11497 = v_11496 & v_8739;
assign v_11498 = v_11479 & v_8173 & v_8174 & v_8189 & v_8190;
assign v_11499 = v_11471 & v_8150 & v_8151 & v_8166 & v_8167;
assign v_11502 = v_11501 & v_7093;
assign v_11503 = v_11501 & ~v_7093 & v_7095 & v_7128 & ~v_7130;
assign v_11504 = v_11501 & ~v_7093 & v_7095 & v_7128 & v_7130;
assign v_11505 = v_11501 & ~v_7093 & v_7095 & ~v_7128;
assign v_11506 = v_11501 & v_7096;
assign v_11507 = v_11501 & ~v_7096;
assign v_11510 = v_11508 & v_11509;
assign v_11511 = v_11508 & v_8244;
assign v_11512 = v_13349 & v_13350;
assign v_11514 = v_11513 & ~v_7093 & ~v_7095 & v_7126;
assign v_11516 = v_11515 & v_7133 & v_7134;
assign v_11517 = v_11515 & v_7133 & ~v_7134;
assign v_11519 = v_11518 & ~v_7145;
assign v_11521 = v_11518 & v_11520;
assign v_11522 = v_11518 & v_7145 & v_7157 & ~v_7158 & v_7166;
assign v_11525 = v_11523 & v_11524;
assign v_11526 = v_11523 & v_7187 & v_7188;
assign v_11527 = v_11523 & v_7187 & ~v_7188 & v_7190;
assign v_11528 = v_11523 & v_7187 & ~v_7188 & ~v_7190 & v_7192;
assign v_11529 = v_11523 & v_7187 & ~v_7188 & ~v_7190 & ~v_7192;
assign v_11531 = v_11530 & v_8267;
assign v_11533 = v_11532 & ~v_7174 & v_7175 & v_7195;
assign v_11536 = v_11534 & v_11535;
assign v_11537 = v_11534 & v_8274;
assign v_11539 = v_11538 & v_7211 & v_7212;
assign v_11540 = v_11538 & v_7211 & ~v_7212 & v_7214;
assign v_11541 = v_11538 & v_7211 & ~v_7212 & ~v_7214 & v_7216;
assign v_11542 = v_11538 & v_7222 & v_7223;
assign v_11543 = v_11538 & v_7225 & v_7226;
assign v_11544 = v_11538 & v_7225 & ~v_7226 & v_7228;
assign v_11545 = v_11538 & v_7225 & ~v_7226 & ~v_7228 & v_7230;
assign v_11546 = v_11538 & v_8286;
assign v_11548 = v_11547 & v_8289;
assign v_11550 = v_11549 & v_7222 & ~v_7223 & v_7235 & v_7236;
assign v_11551 = v_11549 & v_7238 & v_7239;
assign v_11552 = v_11549 & v_7238 & ~v_7239 & v_7241;
assign v_11553 = v_11549 & v_7238 & ~v_7239 & ~v_7241 & v_7243;
assign v_11555 = v_11549 & v_11554;
assign v_11556 = v_13351 & v_13352;
assign v_11558 = v_11557 & v_7250 & v_7251;
assign v_11559 = v_11557 & v_7250 & ~v_7251;
assign v_11561 = v_11560 & v_8303;
assign v_11563 = v_13353 & v_13354;
assign v_11564 = v_11562 & v_7257 & v_7258;
assign v_11565 = v_11562 & v_7257 & ~v_7258 & v_7260;
assign v_11566 = v_11562 & v_7257 & ~v_7258 & ~v_7260 & v_7262;
assign v_11567 = v_11562 & v_8310;
assign v_11569 = v_13355 & v_13356;
assign v_11571 = v_11570 & v_8315;
assign v_11573 = v_11572 & v_7276 & v_7277;
assign v_11574 = v_11572 & v_7276 & ~v_7277 & v_7279;
assign v_11575 = v_11572 & v_7276 & ~v_7277 & ~v_7279 & v_7281;
assign v_11576 = v_11572 & v_7287 & v_7288;
assign v_11577 = v_11572 & v_7290 & v_7291;
assign v_11578 = v_11572 & v_7290 & ~v_7291 & v_7293;
assign v_11579 = v_11572 & v_7290 & ~v_7291 & ~v_7293 & v_7295;
assign v_11580 = v_11572 & v_8325;
assign v_11582 = v_11581 & v_8328;
assign v_11584 = v_11583 & v_7287 & ~v_7288 & v_7300 & v_7301;
assign v_11585 = v_11583 & v_7303 & v_7304;
assign v_11586 = v_11583 & v_7303 & ~v_7304 & v_7306;
assign v_11587 = v_11583 & v_7303 & ~v_7304 & ~v_7306 & v_7308;
assign v_11589 = v_11583 & v_11588;
assign v_11590 = v_13357 & v_13358;
assign v_11592 = v_11591 & v_7315 & v_7316;
assign v_11593 = v_11591 & v_7315 & ~v_7316;
assign v_11595 = v_11594 & v_8342;
assign v_11597 = v_13359 & v_13360;
assign v_11598 = v_11596 & v_7322 & v_7323;
assign v_11599 = v_11596 & v_7322 & ~v_7323 & v_7325;
assign v_11600 = v_11596 & v_7322 & ~v_7323 & ~v_7325 & v_7327;
assign v_11601 = v_11596 & v_8349;
assign v_11603 = v_13361 & v_13362;
assign v_11605 = v_11604 & v_8354;
assign v_11607 = v_11606 & v_7357;
assign v_11608 = v_11606 & ~v_7357 & v_7359 & v_7392 & ~v_7394;
assign v_11609 = v_11606 & ~v_7357 & v_7359 & v_7392 & v_7394;
assign v_11610 = v_11606 & ~v_7357 & v_7359 & ~v_7392;
assign v_11611 = v_11606 & v_7360;
assign v_11612 = v_11606 & ~v_7360;
assign v_11615 = v_11613 & v_11614;
assign v_11616 = v_11613 & v_8370;
assign v_11617 = v_13363 & v_13364;
assign v_11619 = v_11618 & ~v_7357 & ~v_7359 & v_7390;
assign v_11621 = v_11620 & v_7397 & v_7398;
assign v_11622 = v_11620 & v_7397 & ~v_7398;
assign v_11624 = v_11623 & v_7412 & v_7413;
assign v_11625 = v_11623 & v_7412 & ~v_7413 & ~v_7417;
assign v_11627 = v_11626 & v_7412 & ~v_7413 & v_7417;
assign v_11629 = v_11628 & v_7420;
assign v_11631 = v_11630 & v_7424 & v_7425;
assign v_11632 = v_11630 & v_7424 & ~v_7425 & v_7427;
assign v_11633 = v_11630 & v_8386;
assign v_11636 = v_11634 & v_11635;
assign v_11637 = v_11634 & v_8391;
assign v_11639 = v_11638 & v_7454 & ~v_7455 & ~v_7457;
assign v_11640 = v_11638 & v_7459 & ~v_7460;
assign v_11641 = v_11638 & v_7459 & v_7460;
assign v_11642 = v_11638 & v_7449;
assign v_11644 = v_11643 & v_7470 & v_7471;
assign v_11645 = v_11643 & v_7470 & ~v_7471 & ~v_7475;
assign v_11647 = v_11646 & v_7470 & ~v_7471 & v_7475;
assign v_11649 = v_11648 & v_7478;
assign v_11651 = v_11650 & v_7482 & v_7483;
assign v_11652 = v_11650 & v_7482 & ~v_7483 & v_7485;
assign v_11653 = v_11650 & v_8404;
assign v_11656 = v_11654 & v_11655;
assign v_11657 = v_11654 & v_8409;
assign v_11659 = v_6868 & v_11658;
assign v_11660 = v_7507 & v_11638;
assign v_11661 = v_7509 & v_11623;
assign v_11662 = v_7511 & v_11623;
assign v_11663 = v_7513 & v_11623;
assign v_11664 = v_7515 & v_11623;
assign v_11665 = ~v_7515 & v_11606;
assign v_11667 = ~v_7513 & v_11666;
assign v_11669 = ~v_7511 & v_11668;
assign v_11671 = ~v_7509 & v_11670;
assign v_11673 = ~v_7507 & v_11672;
assign v_11675 = ~v_6868 & v_11674;
assign v_11677 = v_11676 & ~v_7535;
assign v_11678 = v_13365 & v_13366;
assign v_11679 = v_11676 & v_7535 & v_7536 & v_7538 & v_7540;
assign v_11680 = v_13367 & v_13368;
assign v_11682 = v_11681 & v_7545 & ~v_7546 & v_7548;
assign v_11683 = v_11681 & v_7555 & ~v_7556 & ~v_7558;
assign v_11684 = v_11681 & v_7560 & ~v_7561;
assign v_11685 = v_11681 & v_7560 & v_7561;
assign v_11686 = v_11681 & v_7550;
assign v_11688 = v_11687 & v_8441;
assign v_11690 = v_11689 & v_8444;
assign v_11691 = v_11681 & v_7545 & v_7546;
assign v_11692 = v_11676 & v_8447;
assign v_11694 = v_11693 & ~v_7571;
assign v_11695 = v_11693 & v_7576 & v_7577;
assign v_11696 = v_11693 & v_7576 & ~v_7577 & ~v_7581;
assign v_11698 = v_11697 & v_7576 & ~v_7577 & v_7581;
assign v_11700 = v_11699 & v_7584;
assign v_11702 = v_11701 & v_7571 & v_7588 & v_7589 & ~v_7590;
assign v_11704 = v_11701 & v_11703;
assign v_11705 = v_11701 & v_7616 & v_7617;
assign v_11706 = v_11701 & v_7616 & ~v_7617;
assign v_11708 = v_11707 & v_7629 & v_7630;
assign v_11709 = v_11707 & v_7629 & ~v_7630;
assign v_11711 = v_11710 & v_7611 & v_7624 & v_7637;
assign v_11712 = v_13369 & v_13370;
assign v_11713 = v_11701 & v_7645 & v_7646;
assign v_11714 = v_11701 & v_7645 & ~v_7646 & ~v_7650;
assign v_11716 = v_11715 & v_7645 & ~v_7646 & v_7650;
assign v_11718 = v_11717 & v_7653;
assign v_11720 = v_11719 & v_8468;
assign v_11722 = v_11721 & v_7664 & ~v_7665 & v_7683;
assign v_11723 = v_11721 & v_7664 & ~v_7665 & ~v_7683;
assign v_11724 = v_11721 & ~v_7666;
assign v_11725 = v_11721 & v_7674 & ~v_7675;
assign v_11726 = v_11721 & v_8475;
assign v_11728 = v_11727 & v_7664 & v_7665 & v_7680 & ~v_7681;
assign v_11730 = v_11729 & v_7687 & ~v_7688 & v_7706;
assign v_11731 = v_11729 & v_7687 & ~v_7688 & ~v_7706;
assign v_11732 = v_11729 & ~v_7689;
assign v_11733 = v_11729 & v_7697 & ~v_7698;
assign v_11734 = v_11729 & v_8484;
assign v_11736 = v_11735 & v_7687 & v_7688 & v_7703 & ~v_7704;
assign v_11738 = v_11737 & v_7710 & ~v_7711 & v_7729;
assign v_11739 = v_11737 & ~v_7712;
assign v_11740 = v_11737 & v_7720 & ~v_7721;
assign v_11741 = v_11737 & v_8492;
assign v_11743 = v_11742 & v_7710 & v_7711 & v_7726 & v_7727;
assign v_11744 = v_11737 & v_7710 & ~v_7711 & ~v_7729;
assign v_11745 = v_11742 & v_7710 & v_7711 & v_7726 & ~v_7727;
assign v_11748 = v_11746 & v_11747;
assign v_11749 = v_11746 & v_7733 & v_7734 & ~v_7735 & ~v_7736;
assign v_11750 = v_11746 & v_7733 & v_7734 & v_7735;
assign v_11751 = v_11746 & v_7733 & ~v_7734 & ~v_7738;
assign v_11753 = v_11752 & v_8505;
assign v_11754 = v_11735 & v_7687 & v_7688 & v_7703 & v_7704;
assign v_11755 = v_11727 & v_7664 & v_7665 & v_7680 & v_7681;
assign v_11757 = v_11756 & v_7745 & ~v_7746 & v_7764;
assign v_11758 = v_11756 & v_7745 & ~v_7746 & ~v_7764;
assign v_11759 = v_11756 & ~v_7747;
assign v_11760 = v_11756 & v_7755 & ~v_7756;
assign v_11761 = v_11756 & v_8514;
assign v_11763 = v_11762 & v_7745 & v_7746 & v_7761 & ~v_7762;
assign v_11765 = v_11764 & v_7768 & ~v_7769 & v_7787;
assign v_11766 = v_11764 & v_7768 & ~v_7769 & ~v_7787;
assign v_11767 = v_11764 & ~v_7770;
assign v_11768 = v_11764 & v_7778 & ~v_7779;
assign v_11769 = v_11764 & v_8523;
assign v_11771 = v_11770 & v_7768 & v_7769 & v_7784 & ~v_7785;
assign v_11773 = v_11772 & v_7791 & ~v_7792 & v_7810;
assign v_11774 = v_11772 & ~v_7793;
assign v_11775 = v_11772 & v_7801 & ~v_7802;
assign v_11776 = v_11772 & v_8531;
assign v_11778 = v_11777 & v_7791 & v_7792 & v_7807 & v_7808;
assign v_11779 = v_11772 & v_7791 & ~v_7792 & ~v_7810;
assign v_11780 = v_11777 & v_7791 & v_7792 & v_7807 & ~v_7808;
assign v_11783 = v_11781 & v_11782;
assign v_11784 = v_11781 & v_7814 & v_7815 & ~v_7816 & ~v_7817;
assign v_11785 = v_11781 & v_7814 & v_7815 & v_7816;
assign v_11786 = v_11781 & v_7814 & ~v_7815 & ~v_7819;
assign v_11788 = v_11787 & v_8544;
assign v_11789 = v_11770 & v_7768 & v_7769 & v_7784 & v_7785;
assign v_11790 = v_11762 & v_7745 & v_7746 & v_7761 & v_7762;
assign v_11792 = v_11791 & v_7826 & ~v_7827 & v_7845;
assign v_11793 = v_11791 & v_7826 & ~v_7827 & ~v_7845;
assign v_11794 = v_11791 & ~v_7828;
assign v_11795 = v_11791 & v_7836 & ~v_7837;
assign v_11796 = v_11791 & v_8553;
assign v_11798 = v_11797 & v_7826 & v_7827 & v_7842 & ~v_7843;
assign v_11800 = v_11799 & v_7849 & ~v_7850 & v_7868;
assign v_11801 = v_11799 & v_7849 & ~v_7850 & ~v_7868;
assign v_11802 = v_11799 & ~v_7851;
assign v_11803 = v_11799 & v_7859 & ~v_7860;
assign v_11804 = v_11799 & v_8562;
assign v_11806 = v_11805 & v_7849 & v_7850 & v_7865 & ~v_7866;
assign v_11808 = v_11807 & v_7872 & ~v_7873 & v_7891;
assign v_11809 = v_11807 & ~v_7874;
assign v_11810 = v_11807 & v_7882 & ~v_7883;
assign v_11811 = v_11807 & v_8570;
assign v_11813 = v_11812 & v_7872 & v_7873 & v_7888 & v_7889;
assign v_11814 = v_11807 & v_7872 & ~v_7873 & ~v_7891;
assign v_11815 = v_11812 & v_7872 & v_7873 & v_7888 & ~v_7889;
assign v_11818 = v_11816 & v_11817;
assign v_11819 = v_11816 & v_7895 & v_7896 & ~v_7897 & ~v_7898;
assign v_11820 = v_11816 & v_7895 & v_7896 & v_7897;
assign v_11821 = v_11816 & v_7895 & ~v_7896 & ~v_7900;
assign v_11823 = v_11822 & v_8583;
assign v_11824 = v_11805 & v_7849 & v_7850 & v_7865 & v_7866;
assign v_11825 = v_11797 & v_7826 & v_7827 & v_7842 & v_7843;
assign v_11827 = v_11826 & v_7907 & ~v_7908 & v_7926;
assign v_11828 = v_11826 & v_7907 & ~v_7908 & ~v_7926;
assign v_11829 = v_11826 & ~v_7909;
assign v_11830 = v_11826 & v_7917 & ~v_7918;
assign v_11831 = v_11826 & v_8592;
assign v_11833 = v_11832 & v_7907 & v_7908 & v_7923 & ~v_7924;
assign v_11835 = v_11834 & v_7930 & ~v_7931 & v_7949;
assign v_11836 = v_11834 & v_7930 & ~v_7931 & ~v_7949;
assign v_11837 = v_11834 & ~v_7932;
assign v_11838 = v_11834 & v_7940 & ~v_7941;
assign v_11839 = v_11834 & v_8601;
assign v_11841 = v_11840 & v_7930 & v_7931 & v_7946 & ~v_7947;
assign v_11843 = v_11842 & v_7953 & ~v_7954 & v_7972;
assign v_11844 = v_11842 & ~v_7955;
assign v_11845 = v_11842 & v_7963 & ~v_7964;
assign v_11846 = v_11842 & v_8609;
assign v_11848 = v_11847 & v_7953 & v_7954 & v_7969 & v_7970;
assign v_11849 = v_11842 & v_7953 & ~v_7954 & ~v_7972;
assign v_11850 = v_11847 & v_7953 & v_7954 & v_7969 & ~v_7970;
assign v_11853 = v_11851 & v_11852;
assign v_11854 = v_11851 & v_7976 & v_7977 & ~v_7978 & ~v_7979;
assign v_11855 = v_11851 & v_7976 & v_7977 & v_7978;
assign v_11856 = v_11851 & v_7976 & ~v_7977 & ~v_7981;
assign v_11858 = v_11857 & v_8622;
assign v_11859 = v_11840 & v_7930 & v_7931 & v_7946 & v_7947;
assign v_11860 = v_11832 & v_7907 & v_7908 & v_7923 & v_7924;
assign v_11862 = v_11861 & v_7988 & ~v_7989 & v_8007;
assign v_11863 = v_11861 & v_7988 & ~v_7989 & ~v_8007;
assign v_11864 = v_11861 & ~v_7990;
assign v_11865 = v_11861 & v_7998 & ~v_7999;
assign v_11866 = v_11861 & v_8631;
assign v_11868 = v_11867 & v_7988 & v_7989 & v_8004 & ~v_8005;
assign v_11870 = v_11869 & v_8011 & ~v_8012 & v_8030;
assign v_11871 = v_11869 & v_8011 & ~v_8012 & ~v_8030;
assign v_11872 = v_11869 & ~v_8013;
assign v_11873 = v_11869 & v_8021 & ~v_8022;
assign v_11874 = v_11869 & v_8640;
assign v_11876 = v_11875 & v_8011 & v_8012 & v_8027 & ~v_8028;
assign v_11878 = v_11877 & v_8034 & ~v_8035 & v_8053;
assign v_11879 = v_11877 & ~v_8036;
assign v_11880 = v_11877 & v_8044 & ~v_8045;
assign v_11881 = v_11877 & v_8648;
assign v_11883 = v_11882 & v_8034 & v_8035 & v_8050 & v_8051;
assign v_11884 = v_11877 & v_8034 & ~v_8035 & ~v_8053;
assign v_11885 = v_11882 & v_8034 & v_8035 & v_8050 & ~v_8051;
assign v_11888 = v_11886 & v_11887;
assign v_11889 = v_11886 & v_8057 & v_8058 & ~v_8059 & ~v_8060;
assign v_11890 = v_11886 & v_8057 & v_8058 & v_8059;
assign v_11891 = v_11886 & v_8057 & ~v_8058 & ~v_8062;
assign v_11893 = v_11892 & v_8661;
assign v_11894 = v_11875 & v_8011 & v_8012 & v_8027 & v_8028;
assign v_11895 = v_11867 & v_7988 & v_7989 & v_8004 & v_8005;
assign v_11897 = v_11896 & v_8069 & ~v_8070 & v_8088;
assign v_11898 = v_11896 & v_8069 & ~v_8070 & ~v_8088;
assign v_11899 = v_11896 & ~v_8071;
assign v_11900 = v_11896 & v_8079 & ~v_8080;
assign v_11901 = v_11896 & v_8670;
assign v_11903 = v_11902 & v_8069 & v_8070 & v_8085 & ~v_8086;
assign v_11905 = v_11904 & v_8092 & ~v_8093 & v_8111;
assign v_11906 = v_11904 & v_8092 & ~v_8093 & ~v_8111;
assign v_11907 = v_11904 & ~v_8094;
assign v_11908 = v_11904 & v_8102 & ~v_8103;
assign v_11909 = v_11904 & v_8679;
assign v_11911 = v_11910 & v_8092 & v_8093 & v_8108 & ~v_8109;
assign v_11913 = v_11912 & v_8115 & ~v_8116 & v_8134;
assign v_11914 = v_11912 & ~v_8117;
assign v_11915 = v_11912 & v_8125 & ~v_8126;
assign v_11916 = v_11912 & v_8687;
assign v_11918 = v_11917 & v_8115 & v_8116 & v_8131 & v_8132;
assign v_11919 = v_11912 & v_8115 & ~v_8116 & ~v_8134;
assign v_11920 = v_11917 & v_8115 & v_8116 & v_8131 & ~v_8132;
assign v_11923 = v_11921 & v_11922;
assign v_11924 = v_11921 & v_8138 & v_8139 & ~v_8140 & ~v_8141;
assign v_11925 = v_11921 & v_8138 & v_8139 & v_8140;
assign v_11926 = v_11921 & v_8138 & ~v_8139 & ~v_8143;
assign v_11928 = v_11927 & v_8700;
assign v_11929 = v_11910 & v_8092 & v_8093 & v_8108 & v_8109;
assign v_11930 = v_11902 & v_8069 & v_8070 & v_8085 & v_8086;
assign v_11932 = v_11931 & v_8150 & ~v_8151 & v_8169;
assign v_11933 = v_11931 & v_8150 & ~v_8151 & ~v_8169;
assign v_11934 = v_11931 & ~v_8152;
assign v_11935 = v_11931 & v_8160 & ~v_8161;
assign v_11936 = v_11931 & v_8709;
assign v_11938 = v_11937 & v_8150 & v_8151 & v_8166 & ~v_8167;
assign v_11940 = v_11939 & v_8173 & ~v_8174 & v_8192;
assign v_11941 = v_11939 & v_8173 & ~v_8174 & ~v_8192;
assign v_11942 = v_11939 & ~v_8175;
assign v_11943 = v_11939 & v_8183 & ~v_8184;
assign v_11944 = v_11939 & v_8718;
assign v_11946 = v_11945 & v_8173 & v_8174 & v_8189 & ~v_8190;
assign v_11948 = v_11947 & v_8196 & ~v_8197 & v_8215;
assign v_11949 = v_11947 & ~v_8198;
assign v_11950 = v_11947 & v_8206 & ~v_8207;
assign v_11951 = v_11947 & v_8726;
assign v_11953 = v_11952 & v_8196 & v_8197 & v_8212 & v_8213;
assign v_11954 = v_11947 & v_8196 & ~v_8197 & ~v_8215;
assign v_11955 = v_11952 & v_8196 & v_8197 & v_8212 & ~v_8213;
assign v_11958 = v_11956 & v_11957;
assign v_11959 = v_11956 & v_8219 & v_8220 & ~v_8221 & ~v_8222;
assign v_11960 = v_11956 & v_8219 & v_8220 & v_8221;
assign v_11961 = v_11956 & v_8219 & ~v_8220 & ~v_8224;
assign v_11963 = v_11962 & v_8739;
assign v_11964 = v_11945 & v_8173 & v_8174 & v_8189 & v_8190;
assign v_11965 = v_11937 & v_8150 & v_8151 & v_8166 & v_8167;
assign v_11968 = v_11967 & ~v_8276;
assign v_11970 = v_8231 & v_11969;
assign v_11971 = v_7093;
assign v_11973 = v_11972 & v_7133 & v_7134;
assign v_11974 = v_11972 & v_7133 & ~v_7134;
assign v_11976 = v_11975 & ~v_7145;
assign v_11978 = v_11975 & v_11977;
assign v_11979 = v_11975 & v_7145 & v_7157 & ~v_7158 & v_7166;
assign v_11982 = v_11980 & v_11981;
assign v_11983 = v_11980 & v_7187 & v_7188;
assign v_11984 = v_11980 & v_7187 & ~v_7188 & v_7190;
assign v_11985 = v_11980 & v_7187 & ~v_7188 & ~v_7190 & v_7192;
assign v_11986 = v_11980 & v_7187 & ~v_7188 & ~v_7190 & ~v_7192;
assign v_11988 = v_11987 & v_8267;
assign v_11990 = v_11989 & ~v_7174 & v_7175 & v_7195;
assign v_11993 = v_11991 & v_11992;
assign v_11994 = v_11991 & v_8274;
assign v_11996 = ~v_8231 & v_11995;
assign v_11998 = v_11997 & v_7211 & v_7212;
assign v_11999 = v_11997 & v_7211 & ~v_7212 & v_7214;
assign v_12000 = v_11997 & v_7211 & ~v_7212 & ~v_7214 & v_7216;
assign v_12001 = v_11997 & v_7222 & v_7223;
assign v_12002 = v_11997 & v_7225 & v_7226;
assign v_12003 = v_11997 & v_7225 & ~v_7226 & v_7228;
assign v_12004 = v_11997 & v_7225 & ~v_7226 & ~v_7228 & v_7230;
assign v_12005 = v_11997 & v_8286;
assign v_12007 = v_12006 & v_8289;
assign v_12009 = v_12008 & v_7222 & ~v_7223 & v_7235 & v_7236;
assign v_12010 = v_12008 & v_7238 & v_7239;
assign v_12011 = v_12008 & v_7238 & ~v_7239 & v_7241;
assign v_12012 = v_12008 & v_7238 & ~v_7239 & ~v_7241 & v_7243;
assign v_12014 = v_12008 & v_12013;
assign v_12015 = v_13371 & v_13372;
assign v_12017 = v_12016 & v_7250 & v_7251;
assign v_12018 = v_12016 & v_7250 & ~v_7251;
assign v_12020 = v_12019 & v_8303;
assign v_12022 = v_13373 & v_13374;
assign v_12023 = v_12021 & v_7257 & v_7258;
assign v_12024 = v_12021 & v_7257 & ~v_7258 & v_7260;
assign v_12025 = v_12021 & v_7257 & ~v_7258 & ~v_7260 & v_7262;
assign v_12026 = v_12021 & v_8310;
assign v_12028 = v_13375 & v_13376;
assign v_12030 = v_12029 & v_8315;
assign v_12032 = v_12031 & v_7276 & v_7277;
assign v_12033 = v_12031 & v_7276 & ~v_7277 & v_7279;
assign v_12034 = v_12031 & v_7276 & ~v_7277 & ~v_7279 & v_7281;
assign v_12035 = v_12031 & v_7287 & v_7288;
assign v_12036 = v_12031 & v_7290 & v_7291;
assign v_12037 = v_12031 & v_7290 & ~v_7291 & v_7293;
assign v_12038 = v_12031 & v_7290 & ~v_7291 & ~v_7293 & v_7295;
assign v_12039 = v_12031 & v_8325;
assign v_12041 = v_12040 & v_8328;
assign v_12043 = v_12042 & v_7287 & ~v_7288 & v_7300 & v_7301;
assign v_12044 = v_12042 & v_7303 & v_7304;
assign v_12045 = v_12042 & v_7303 & ~v_7304 & v_7306;
assign v_12046 = v_12042 & v_7303 & ~v_7304 & ~v_7306 & v_7308;
assign v_12048 = v_12042 & v_12047;
assign v_12049 = v_13377 & v_13378;
assign v_12051 = v_12050 & v_7315 & v_7316;
assign v_12052 = v_12050 & v_7315 & ~v_7316;
assign v_12054 = v_12053 & v_8342;
assign v_12056 = v_13379 & v_13380;
assign v_12057 = v_12055 & v_7322 & v_7323;
assign v_12058 = v_12055 & v_7322 & ~v_7323 & v_7325;
assign v_12059 = v_12055 & v_7322 & ~v_7323 & ~v_7325 & v_7327;
assign v_12060 = v_12055 & v_8349;
assign v_12062 = v_13381 & v_13382;
assign v_12064 = v_12063 & v_8354;
assign v_12066 = v_12065 & v_7357;
assign v_12068 = v_12067 & v_7397 & v_7398;
assign v_12069 = v_12067 & v_7397 & ~v_7398;
assign v_12071 = v_12070 & v_7412 & v_7413;
assign v_12072 = v_12070 & v_7420;
assign v_12074 = v_12073 & v_7424 & v_7425;
assign v_12075 = v_12073 & v_7424 & ~v_7425 & v_7427;
assign v_12076 = v_12073 & v_8386;
assign v_12079 = v_12077 & v_12078;
assign v_12080 = v_12077 & v_8391;
assign v_12082 = v_12081 & v_7454 & ~v_7455 & ~v_7457;
assign v_12083 = v_12081 & v_7459 & ~v_7460;
assign v_12084 = v_12081 & v_7459 & v_7460;
assign v_12085 = v_12081 & v_7449;
assign v_12087 = v_12086 & v_7470 & v_7471;
assign v_12088 = v_12086 & v_7478;
assign v_12090 = v_12089 & v_7482 & v_7483;
assign v_12091 = v_12089 & v_7482 & ~v_7483 & v_7485;
assign v_12092 = v_12089 & v_8404;
assign v_12095 = v_12093 & v_12094;
assign v_12096 = v_12093 & v_8409;
assign v_12098 = v_6868 & v_12097;
assign v_12099 = v_7507 & v_12081;
assign v_12100 = v_7509 & v_12070;
assign v_12101 = v_7511 & v_12070;
assign v_12102 = v_7513 & v_12070;
assign v_12103 = v_7515 & v_12070;
assign v_12104 = ~v_7515 & v_12065;
assign v_12106 = ~v_7513 & v_12105;
assign v_12108 = ~v_7511 & v_12107;
assign v_12110 = ~v_7509 & v_12109;
assign v_12112 = ~v_7507 & v_12111;
assign v_12114 = ~v_6868 & v_12113;
assign v_12116 = v_12115 & ~v_7535;
assign v_12117 = v_13383 & v_13384;
assign v_12118 = v_12115 & v_7535 & v_7536 & v_7538 & v_7540;
assign v_12119 = v_13385 & v_13386;
assign v_12121 = v_12120 & v_7545 & ~v_7546 & v_7548;
assign v_12122 = v_12120 & v_7555 & ~v_7556 & ~v_7558;
assign v_12123 = v_12120 & v_7560 & ~v_7561;
assign v_12124 = v_12120 & v_7560 & v_7561;
assign v_12125 = v_12120 & v_7550;
assign v_12127 = v_12126 & v_8441;
assign v_12129 = v_12128 & v_8444;
assign v_12130 = v_12120 & v_7545 & v_7546;
assign v_12131 = v_12115 & v_8447;
assign v_12133 = v_12132 & ~v_7571;
assign v_12134 = v_12132 & v_7576 & v_7577;
assign v_12135 = v_12132 & v_7584;
assign v_12137 = v_12136 & v_7571 & v_7588 & v_7589 & ~v_7590;
assign v_12139 = v_12136 & v_12138;
assign v_12140 = v_12136 & v_7616 & v_7617;
assign v_12141 = v_12136 & v_7616 & ~v_7617;
assign v_12143 = v_12142 & v_7629 & v_7630;
assign v_12144 = v_12142 & v_7629 & ~v_7630;
assign v_12146 = v_12145 & v_7611 & v_7624 & v_7637;
assign v_12147 = v_13387 & v_13388;
assign v_12148 = v_12136 & v_7645 & v_7646;
assign v_12149 = v_12136 & v_7653;
assign v_12151 = v_12150 & v_8468;
assign v_12153 = v_12152 & v_7664 & ~v_7665 & v_7683;
assign v_12154 = v_12152 & v_7664 & ~v_7665 & ~v_7683;
assign v_12155 = v_12152 & ~v_7666;
assign v_12156 = v_12152 & v_7674 & ~v_7675;
assign v_12157 = v_12152 & v_8475;
assign v_12159 = v_12158 & v_7664 & v_7665 & v_7680 & ~v_7681;
assign v_12161 = v_12160 & v_7687 & ~v_7688 & v_7706;
assign v_12162 = v_12160 & v_7687 & ~v_7688 & ~v_7706;
assign v_12163 = v_12160 & ~v_7689;
assign v_12164 = v_12160 & v_7697 & ~v_7698;
assign v_12165 = v_12160 & v_8484;
assign v_12167 = v_12166 & v_7687 & v_7688 & v_7703 & ~v_7704;
assign v_12169 = v_12168 & v_7710 & ~v_7711 & v_7729;
assign v_12170 = v_12168 & ~v_7712;
assign v_12171 = v_12168 & v_7720 & ~v_7721;
assign v_12172 = v_12168 & v_8492;
assign v_12174 = v_12173 & v_7710 & v_7711 & v_7726 & v_7727;
assign v_12175 = v_12168 & v_7710 & ~v_7711 & ~v_7729;
assign v_12176 = v_12173 & v_7710 & v_7711 & v_7726 & ~v_7727;
assign v_12179 = v_12177 & v_12178;
assign v_12180 = v_12177 & v_7733 & v_7734 & ~v_7735 & ~v_7736;
assign v_12181 = v_12177 & v_7733 & v_7734 & v_7735;
assign v_12182 = v_12177 & v_7733 & ~v_7734 & ~v_7738;
assign v_12184 = v_12183 & v_8505;
assign v_12185 = v_12166 & v_7687 & v_7688 & v_7703 & v_7704;
assign v_12186 = v_12158 & v_7664 & v_7665 & v_7680 & v_7681;
assign v_12188 = v_12187 & v_7745 & ~v_7746 & v_7764;
assign v_12189 = v_12187 & v_7745 & ~v_7746 & ~v_7764;
assign v_12190 = v_12187 & ~v_7747;
assign v_12191 = v_12187 & v_7755 & ~v_7756;
assign v_12192 = v_12187 & v_8514;
assign v_12194 = v_12193 & v_7745 & v_7746 & v_7761 & ~v_7762;
assign v_12196 = v_12195 & v_7768 & ~v_7769 & v_7787;
assign v_12197 = v_12195 & v_7768 & ~v_7769 & ~v_7787;
assign v_12198 = v_12195 & ~v_7770;
assign v_12199 = v_12195 & v_7778 & ~v_7779;
assign v_12200 = v_12195 & v_8523;
assign v_12202 = v_12201 & v_7768 & v_7769 & v_7784 & ~v_7785;
assign v_12204 = v_12203 & v_7791 & ~v_7792 & v_7810;
assign v_12205 = v_12203 & ~v_7793;
assign v_12206 = v_12203 & v_7801 & ~v_7802;
assign v_12207 = v_12203 & v_8531;
assign v_12209 = v_12208 & v_7791 & v_7792 & v_7807 & v_7808;
assign v_12210 = v_12203 & v_7791 & ~v_7792 & ~v_7810;
assign v_12211 = v_12208 & v_7791 & v_7792 & v_7807 & ~v_7808;
assign v_12214 = v_12212 & v_12213;
assign v_12215 = v_12212 & v_7814 & v_7815 & ~v_7816 & ~v_7817;
assign v_12216 = v_12212 & v_7814 & v_7815 & v_7816;
assign v_12217 = v_12212 & v_7814 & ~v_7815 & ~v_7819;
assign v_12219 = v_12218 & v_8544;
assign v_12220 = v_12201 & v_7768 & v_7769 & v_7784 & v_7785;
assign v_12221 = v_12193 & v_7745 & v_7746 & v_7761 & v_7762;
assign v_12223 = v_12222 & v_7826 & ~v_7827 & v_7845;
assign v_12224 = v_12222 & v_7826 & ~v_7827 & ~v_7845;
assign v_12225 = v_12222 & ~v_7828;
assign v_12226 = v_12222 & v_7836 & ~v_7837;
assign v_12227 = v_12222 & v_8553;
assign v_12229 = v_12228 & v_7826 & v_7827 & v_7842 & ~v_7843;
assign v_12231 = v_12230 & v_7849 & ~v_7850 & v_7868;
assign v_12232 = v_12230 & v_7849 & ~v_7850 & ~v_7868;
assign v_12233 = v_12230 & ~v_7851;
assign v_12234 = v_12230 & v_7859 & ~v_7860;
assign v_12235 = v_12230 & v_8562;
assign v_12237 = v_12236 & v_7849 & v_7850 & v_7865 & ~v_7866;
assign v_12239 = v_12238 & v_7872 & ~v_7873 & v_7891;
assign v_12240 = v_12238 & ~v_7874;
assign v_12241 = v_12238 & v_7882 & ~v_7883;
assign v_12242 = v_12238 & v_8570;
assign v_12244 = v_12243 & v_7872 & v_7873 & v_7888 & v_7889;
assign v_12245 = v_12238 & v_7872 & ~v_7873 & ~v_7891;
assign v_12246 = v_12243 & v_7872 & v_7873 & v_7888 & ~v_7889;
assign v_12249 = v_12247 & v_12248;
assign v_12250 = v_12247 & v_7895 & v_7896 & ~v_7897 & ~v_7898;
assign v_12251 = v_12247 & v_7895 & v_7896 & v_7897;
assign v_12252 = v_12247 & v_7895 & ~v_7896 & ~v_7900;
assign v_12254 = v_12253 & v_8583;
assign v_12255 = v_12236 & v_7849 & v_7850 & v_7865 & v_7866;
assign v_12256 = v_12228 & v_7826 & v_7827 & v_7842 & v_7843;
assign v_12258 = v_12257 & v_7907 & ~v_7908 & v_7926;
assign v_12259 = v_12257 & v_7907 & ~v_7908 & ~v_7926;
assign v_12260 = v_12257 & ~v_7909;
assign v_12261 = v_12257 & v_7917 & ~v_7918;
assign v_12262 = v_12257 & v_8592;
assign v_12264 = v_12263 & v_7907 & v_7908 & v_7923 & ~v_7924;
assign v_12266 = v_12265 & v_7930 & ~v_7931 & v_7949;
assign v_12267 = v_12265 & v_7930 & ~v_7931 & ~v_7949;
assign v_12268 = v_12265 & ~v_7932;
assign v_12269 = v_12265 & v_7940 & ~v_7941;
assign v_12270 = v_12265 & v_8601;
assign v_12272 = v_12271 & v_7930 & v_7931 & v_7946 & ~v_7947;
assign v_12274 = v_12273 & v_7953 & ~v_7954 & v_7972;
assign v_12275 = v_12273 & ~v_7955;
assign v_12276 = v_12273 & v_7963 & ~v_7964;
assign v_12277 = v_12273 & v_8609;
assign v_12279 = v_12278 & v_7953 & v_7954 & v_7969 & v_7970;
assign v_12280 = v_12273 & v_7953 & ~v_7954 & ~v_7972;
assign v_12281 = v_12278 & v_7953 & v_7954 & v_7969 & ~v_7970;
assign v_12284 = v_12282 & v_12283;
assign v_12285 = v_12282 & v_7976 & v_7977 & ~v_7978 & ~v_7979;
assign v_12286 = v_12282 & v_7976 & v_7977 & v_7978;
assign v_12287 = v_12282 & v_7976 & ~v_7977 & ~v_7981;
assign v_12289 = v_12288 & v_8622;
assign v_12290 = v_12271 & v_7930 & v_7931 & v_7946 & v_7947;
assign v_12291 = v_12263 & v_7907 & v_7908 & v_7923 & v_7924;
assign v_12293 = v_12292 & v_7988 & ~v_7989 & v_8007;
assign v_12294 = v_12292 & v_7988 & ~v_7989 & ~v_8007;
assign v_12295 = v_12292 & ~v_7990;
assign v_12296 = v_12292 & v_7998 & ~v_7999;
assign v_12297 = v_12292 & v_8631;
assign v_12299 = v_12298 & v_7988 & v_7989 & v_8004 & ~v_8005;
assign v_12301 = v_12300 & v_8011 & ~v_8012 & v_8030;
assign v_12302 = v_12300 & v_8011 & ~v_8012 & ~v_8030;
assign v_12303 = v_12300 & ~v_8013;
assign v_12304 = v_12300 & v_8021 & ~v_8022;
assign v_12305 = v_12300 & v_8640;
assign v_12307 = v_12306 & v_8011 & v_8012 & v_8027 & ~v_8028;
assign v_12309 = v_12308 & v_8034 & ~v_8035 & v_8053;
assign v_12310 = v_12308 & ~v_8036;
assign v_12311 = v_12308 & v_8044 & ~v_8045;
assign v_12312 = v_12308 & v_8648;
assign v_12314 = v_12313 & v_8034 & v_8035 & v_8050 & v_8051;
assign v_12315 = v_12308 & v_8034 & ~v_8035 & ~v_8053;
assign v_12316 = v_12313 & v_8034 & v_8035 & v_8050 & ~v_8051;
assign v_12319 = v_12317 & v_12318;
assign v_12320 = v_12317 & v_8057 & v_8058 & ~v_8059 & ~v_8060;
assign v_12321 = v_12317 & v_8057 & v_8058 & v_8059;
assign v_12322 = v_12317 & v_8057 & ~v_8058 & ~v_8062;
assign v_12324 = v_12323 & v_8661;
assign v_12325 = v_12306 & v_8011 & v_8012 & v_8027 & v_8028;
assign v_12326 = v_12298 & v_7988 & v_7989 & v_8004 & v_8005;
assign v_12328 = v_12327 & v_8069 & ~v_8070 & v_8088;
assign v_12329 = v_12327 & v_8069 & ~v_8070 & ~v_8088;
assign v_12330 = v_12327 & ~v_8071;
assign v_12331 = v_12327 & v_8079 & ~v_8080;
assign v_12332 = v_12327 & v_8670;
assign v_12334 = v_12333 & v_8069 & v_8070 & v_8085 & ~v_8086;
assign v_12336 = v_12335 & v_8092 & ~v_8093 & v_8111;
assign v_12337 = v_12335 & v_8092 & ~v_8093 & ~v_8111;
assign v_12338 = v_12335 & ~v_8094;
assign v_12339 = v_12335 & v_8102 & ~v_8103;
assign v_12340 = v_12335 & v_8679;
assign v_12342 = v_12341 & v_8092 & v_8093 & v_8108 & ~v_8109;
assign v_12344 = v_12343 & v_8115 & ~v_8116 & v_8134;
assign v_12345 = v_12343 & ~v_8117;
assign v_12346 = v_12343 & v_8125 & ~v_8126;
assign v_12347 = v_12343 & v_8687;
assign v_12349 = v_12348 & v_8115 & v_8116 & v_8131 & v_8132;
assign v_12350 = v_12343 & v_8115 & ~v_8116 & ~v_8134;
assign v_12351 = v_12348 & v_8115 & v_8116 & v_8131 & ~v_8132;
assign v_12354 = v_12352 & v_12353;
assign v_12355 = v_12352 & v_8138 & v_8139 & ~v_8140 & ~v_8141;
assign v_12356 = v_12352 & v_8138 & v_8139 & v_8140;
assign v_12357 = v_12352 & v_8138 & ~v_8139 & ~v_8143;
assign v_12359 = v_12358 & v_8700;
assign v_12360 = v_12341 & v_8092 & v_8093 & v_8108 & v_8109;
assign v_12361 = v_12333 & v_8069 & v_8070 & v_8085 & v_8086;
assign v_12363 = v_12362 & v_8150 & ~v_8151 & v_8169;
assign v_12364 = v_12362 & v_8150 & ~v_8151 & ~v_8169;
assign v_12365 = v_12362 & ~v_8152;
assign v_12366 = v_12362 & v_8160 & ~v_8161;
assign v_12367 = v_12362 & v_8709;
assign v_12369 = v_12368 & v_8150 & v_8151 & v_8166 & ~v_8167;
assign v_12371 = v_12370 & v_8173 & ~v_8174 & v_8192;
assign v_12372 = v_12370 & v_8173 & ~v_8174 & ~v_8192;
assign v_12373 = v_12370 & ~v_8175;
assign v_12374 = v_12370 & v_8183 & ~v_8184;
assign v_12375 = v_12370 & v_8718;
assign v_12377 = v_12376 & v_8173 & v_8174 & v_8189 & ~v_8190;
assign v_12379 = v_12378 & v_8196 & ~v_8197 & v_8215;
assign v_12380 = v_12378 & ~v_8198;
assign v_12381 = v_12378 & v_8206 & ~v_8207;
assign v_12382 = v_12378 & v_8726;
assign v_12384 = v_12383 & v_8196 & v_8197 & v_8212 & v_8213;
assign v_12385 = v_12378 & v_8196 & ~v_8197 & ~v_8215;
assign v_12386 = v_12383 & v_8196 & v_8197 & v_8212 & ~v_8213;
assign v_12389 = v_12387 & v_12388;
assign v_12390 = v_12387 & v_8219 & v_8220 & ~v_8221 & ~v_8222;
assign v_12391 = v_12387 & v_8219 & v_8220 & v_8221;
assign v_12392 = v_12387 & v_8219 & ~v_8220 & ~v_8224;
assign v_12394 = v_12393 & v_8739;
assign v_12395 = v_12376 & v_8173 & v_8174 & v_8189 & v_8190;
assign v_12396 = v_12368 & v_8150 & v_8151 & v_8166 & v_8167;
assign v_12399 = v_12398 & v_7093;
assign v_12400 = v_12398 & ~v_7093 & v_7095 & v_7128 & ~v_7130;
assign v_12401 = v_12398 & ~v_7093 & v_7095 & v_7128 & v_7130;
assign v_12402 = v_12398 & ~v_7093 & v_7095 & ~v_7128;
assign v_12403 = v_12398 & v_7096;
assign v_12404 = v_12398 & ~v_7096;
assign v_12407 = v_12405 & v_12406;
assign v_12408 = v_12405 & v_8244;
assign v_12409 = v_13389 & v_13390;
assign v_12411 = v_12410 & ~v_7093 & ~v_7095 & v_7126;
assign v_12413 = v_12412 & v_7133 & v_7134;
assign v_12414 = v_12412 & v_7133 & ~v_7134;
assign v_12416 = v_12415 & ~v_7145;
assign v_12418 = v_12415 & v_12417;
assign v_12419 = v_12415 & v_7145 & v_7157 & ~v_7158 & v_7166;
assign v_12422 = v_12420 & v_12421;
assign v_12423 = v_12420 & v_7187 & v_7188;
assign v_12424 = v_12420 & v_7187 & ~v_7188 & v_7190;
assign v_12425 = v_12420 & v_7187 & ~v_7188 & ~v_7190 & v_7192;
assign v_12426 = v_12420 & v_7187 & ~v_7188 & ~v_7190 & ~v_7192;
assign v_12428 = v_12427 & v_8267;
assign v_12430 = v_12429 & ~v_7174 & v_7175 & v_7195;
assign v_12433 = v_12431 & v_12432;
assign v_12434 = v_12431 & v_8274;
assign v_12436 = v_12435 & v_7211 & v_7212;
assign v_12437 = v_12435 & v_7211 & ~v_7212 & v_7214;
assign v_12438 = v_12435 & v_7211 & ~v_7212 & ~v_7214 & v_7216;
assign v_12439 = v_12435 & v_7222 & v_7223;
assign v_12440 = v_12435 & v_7225 & v_7226;
assign v_12441 = v_12435 & v_7225 & ~v_7226 & v_7228;
assign v_12442 = v_12435 & v_7225 & ~v_7226 & ~v_7228 & v_7230;
assign v_12443 = v_12435 & v_8286;
assign v_12445 = v_12444 & v_8289;
assign v_12447 = v_12446 & v_7222 & ~v_7223 & v_7235 & v_7236;
assign v_12448 = v_12446 & v_7238 & v_7239;
assign v_12449 = v_12446 & v_7238 & ~v_7239 & v_7241;
assign v_12450 = v_12446 & v_7238 & ~v_7239 & ~v_7241 & v_7243;
assign v_12452 = v_12446 & v_12451;
assign v_12453 = v_13391 & v_13392;
assign v_12455 = v_12454 & v_7250 & v_7251;
assign v_12456 = v_12454 & v_7250 & ~v_7251;
assign v_12458 = v_12457 & v_8303;
assign v_12460 = v_13393 & v_13394;
assign v_12461 = v_12459 & v_7257 & v_7258;
assign v_12462 = v_12459 & v_7257 & ~v_7258 & v_7260;
assign v_12463 = v_12459 & v_7257 & ~v_7258 & ~v_7260 & v_7262;
assign v_12464 = v_12459 & v_8310;
assign v_12466 = v_13395 & v_13396;
assign v_12468 = v_12467 & v_8315;
assign v_12470 = v_12469 & v_7276 & v_7277;
assign v_12471 = v_12469 & v_7276 & ~v_7277 & v_7279;
assign v_12472 = v_12469 & v_7276 & ~v_7277 & ~v_7279 & v_7281;
assign v_12473 = v_12469 & v_7287 & v_7288;
assign v_12474 = v_12469 & v_7290 & v_7291;
assign v_12475 = v_12469 & v_7290 & ~v_7291 & v_7293;
assign v_12476 = v_12469 & v_7290 & ~v_7291 & ~v_7293 & v_7295;
assign v_12477 = v_12469 & v_8325;
assign v_12479 = v_12478 & v_8328;
assign v_12481 = v_12480 & v_7287 & ~v_7288 & v_7300 & v_7301;
assign v_12482 = v_12480 & v_7303 & v_7304;
assign v_12483 = v_12480 & v_7303 & ~v_7304 & v_7306;
assign v_12484 = v_12480 & v_7303 & ~v_7304 & ~v_7306 & v_7308;
assign v_12486 = v_12480 & v_12485;
assign v_12487 = v_13397 & v_13398;
assign v_12489 = v_12488 & v_7315 & v_7316;
assign v_12490 = v_12488 & v_7315 & ~v_7316;
assign v_12492 = v_12491 & v_8342;
assign v_12494 = v_13399 & v_13400;
assign v_12495 = v_12493 & v_7322 & v_7323;
assign v_12496 = v_12493 & v_7322 & ~v_7323 & v_7325;
assign v_12497 = v_12493 & v_7322 & ~v_7323 & ~v_7325 & v_7327;
assign v_12498 = v_12493 & v_8349;
assign v_12500 = v_13401 & v_13402;
assign v_12502 = v_12501 & v_8354;
assign v_12504 = v_12503 & v_7357;
assign v_12505 = v_12503 & ~v_7357 & v_7359 & v_7392 & ~v_7394;
assign v_12506 = v_12503 & ~v_7357 & v_7359 & v_7392 & v_7394;
assign v_12507 = v_12503 & ~v_7357 & v_7359 & ~v_7392;
assign v_12508 = v_12503 & v_7360;
assign v_12509 = v_12503 & ~v_7360;
assign v_12512 = v_12510 & v_12511;
assign v_12513 = v_12510 & v_8370;
assign v_12514 = v_13403 & v_13404;
assign v_12516 = v_12515 & ~v_7357 & ~v_7359 & v_7390;
assign v_12518 = v_12517 & v_7397 & v_7398;
assign v_12519 = v_12517 & v_7397 & ~v_7398;
assign v_12521 = v_12520 & v_7412 & v_7413;
assign v_12522 = v_12520 & v_7412 & ~v_7413 & ~v_7417;
assign v_12524 = v_12523 & v_7412 & ~v_7413 & v_7417;
assign v_12526 = v_12525 & v_7420;
assign v_12528 = v_12527 & v_7424 & v_7425;
assign v_12529 = v_12527 & v_7424 & ~v_7425 & v_7427;
assign v_12530 = v_12527 & v_8386;
assign v_12533 = v_12531 & v_12532;
assign v_12534 = v_12531 & v_8391;
assign v_12536 = v_12535 & v_7454 & ~v_7455 & ~v_7457;
assign v_12537 = v_12535 & v_7459 & ~v_7460;
assign v_12538 = v_12535 & v_7459 & v_7460;
assign v_12539 = v_12535 & v_7449;
assign v_12541 = v_12540 & v_7470 & v_7471;
assign v_12542 = v_12540 & v_7470 & ~v_7471 & ~v_7475;
assign v_12544 = v_12543 & v_7470 & ~v_7471 & v_7475;
assign v_12546 = v_12545 & v_7478;
assign v_12548 = v_12547 & v_7482 & v_7483;
assign v_12549 = v_12547 & v_7482 & ~v_7483 & v_7485;
assign v_12550 = v_12547 & v_8404;
assign v_12553 = v_12551 & v_12552;
assign v_12554 = v_12551 & v_8409;
assign v_12556 = v_6868 & v_12555;
assign v_12557 = v_7507 & v_12535;
assign v_12558 = v_7509 & v_12520;
assign v_12559 = v_7511 & v_12520;
assign v_12560 = v_7513 & v_12520;
assign v_12561 = v_7515 & v_12520;
assign v_12562 = ~v_7515 & v_12503;
assign v_12564 = ~v_7513 & v_12563;
assign v_12566 = ~v_7511 & v_12565;
assign v_12568 = ~v_7509 & v_12567;
assign v_12570 = ~v_7507 & v_12569;
assign v_12572 = ~v_6868 & v_12571;
assign v_12574 = v_12573 & ~v_7535;
assign v_12575 = v_13405 & v_13406;
assign v_12576 = v_12573 & v_7535 & v_7536 & v_7538 & v_7540;
assign v_12577 = v_13407 & v_13408;
assign v_12579 = v_12578 & v_7545 & ~v_7546 & v_7548;
assign v_12580 = v_12578 & v_7555 & ~v_7556 & ~v_7558;
assign v_12581 = v_12578 & v_7560 & ~v_7561;
assign v_12582 = v_12578 & v_7560 & v_7561;
assign v_12583 = v_12578 & v_7550;
assign v_12585 = v_12584 & v_8441;
assign v_12587 = v_12586 & v_8444;
assign v_12588 = v_12578 & v_7545 & v_7546;
assign v_12589 = v_12573 & v_8447;
assign v_12591 = v_12590 & ~v_7571;
assign v_12592 = v_12590 & v_7576 & v_7577;
assign v_12593 = v_12590 & v_7576 & ~v_7577 & ~v_7581;
assign v_12595 = v_12594 & v_7576 & ~v_7577 & v_7581;
assign v_12597 = v_12596 & v_7584;
assign v_12599 = v_12598 & v_7571 & v_7588 & v_7589 & ~v_7590;
assign v_12601 = v_12598 & v_12600;
assign v_12602 = v_12598 & v_7616 & v_7617;
assign v_12603 = v_12598 & v_7616 & ~v_7617;
assign v_12605 = v_12604 & v_7629 & v_7630;
assign v_12606 = v_12604 & v_7629 & ~v_7630;
assign v_12608 = v_12607 & v_7611 & v_7624 & v_7637;
assign v_12609 = v_13409 & v_13410;
assign v_12610 = v_12598 & v_7645 & v_7646;
assign v_12611 = v_12598 & v_7645 & ~v_7646 & ~v_7650;
assign v_12613 = v_12612 & v_7645 & ~v_7646 & v_7650;
assign v_12615 = v_12614 & v_7653;
assign v_12617 = v_12616 & v_8468;
assign v_12619 = v_12618 & v_7664 & ~v_7665 & v_7683;
assign v_12620 = v_12618 & v_7664 & ~v_7665 & ~v_7683;
assign v_12621 = v_12618 & ~v_7666;
assign v_12622 = v_12618 & v_7674 & ~v_7675;
assign v_12623 = v_12618 & v_8475;
assign v_12625 = v_12624 & v_7664 & v_7665 & v_7680 & ~v_7681;
assign v_12627 = v_12626 & v_7687 & ~v_7688 & v_7706;
assign v_12628 = v_12626 & v_7687 & ~v_7688 & ~v_7706;
assign v_12629 = v_12626 & ~v_7689;
assign v_12630 = v_12626 & v_7697 & ~v_7698;
assign v_12631 = v_12626 & v_8484;
assign v_12633 = v_12632 & v_7687 & v_7688 & v_7703 & ~v_7704;
assign v_12635 = v_12634 & v_7710 & ~v_7711 & v_7729;
assign v_12636 = v_12634 & ~v_7712;
assign v_12637 = v_12634 & v_7720 & ~v_7721;
assign v_12638 = v_12634 & v_8492;
assign v_12640 = v_12639 & v_7710 & v_7711 & v_7726 & v_7727;
assign v_12641 = v_12634 & v_7710 & ~v_7711 & ~v_7729;
assign v_12642 = v_12639 & v_7710 & v_7711 & v_7726 & ~v_7727;
assign v_12645 = v_12643 & v_12644;
assign v_12646 = v_12643 & v_7733 & v_7734 & ~v_7735 & ~v_7736;
assign v_12647 = v_12643 & v_7733 & v_7734 & v_7735;
assign v_12648 = v_12643 & v_7733 & ~v_7734 & ~v_7738;
assign v_12650 = v_12649 & v_8505;
assign v_12651 = v_12632 & v_7687 & v_7688 & v_7703 & v_7704;
assign v_12652 = v_12624 & v_7664 & v_7665 & v_7680 & v_7681;
assign v_12654 = v_12653 & v_7745 & ~v_7746 & v_7764;
assign v_12655 = v_12653 & v_7745 & ~v_7746 & ~v_7764;
assign v_12656 = v_12653 & ~v_7747;
assign v_12657 = v_12653 & v_7755 & ~v_7756;
assign v_12658 = v_12653 & v_8514;
assign v_12660 = v_12659 & v_7745 & v_7746 & v_7761 & ~v_7762;
assign v_12662 = v_12661 & v_7768 & ~v_7769 & v_7787;
assign v_12663 = v_12661 & v_7768 & ~v_7769 & ~v_7787;
assign v_12664 = v_12661 & ~v_7770;
assign v_12665 = v_12661 & v_7778 & ~v_7779;
assign v_12666 = v_12661 & v_8523;
assign v_12668 = v_12667 & v_7768 & v_7769 & v_7784 & ~v_7785;
assign v_12670 = v_12669 & v_7791 & ~v_7792 & v_7810;
assign v_12671 = v_12669 & ~v_7793;
assign v_12672 = v_12669 & v_7801 & ~v_7802;
assign v_12673 = v_12669 & v_8531;
assign v_12675 = v_12674 & v_7791 & v_7792 & v_7807 & v_7808;
assign v_12676 = v_12669 & v_7791 & ~v_7792 & ~v_7810;
assign v_12677 = v_12674 & v_7791 & v_7792 & v_7807 & ~v_7808;
assign v_12680 = v_12678 & v_12679;
assign v_12681 = v_12678 & v_7814 & v_7815 & ~v_7816 & ~v_7817;
assign v_12682 = v_12678 & v_7814 & v_7815 & v_7816;
assign v_12683 = v_12678 & v_7814 & ~v_7815 & ~v_7819;
assign v_12685 = v_12684 & v_8544;
assign v_12686 = v_12667 & v_7768 & v_7769 & v_7784 & v_7785;
assign v_12687 = v_12659 & v_7745 & v_7746 & v_7761 & v_7762;
assign v_12689 = v_12688 & v_7826 & ~v_7827 & v_7845;
assign v_12690 = v_12688 & v_7826 & ~v_7827 & ~v_7845;
assign v_12691 = v_12688 & ~v_7828;
assign v_12692 = v_12688 & v_7836 & ~v_7837;
assign v_12693 = v_12688 & v_8553;
assign v_12695 = v_12694 & v_7826 & v_7827 & v_7842 & ~v_7843;
assign v_12697 = v_12696 & v_7849 & ~v_7850 & v_7868;
assign v_12698 = v_12696 & v_7849 & ~v_7850 & ~v_7868;
assign v_12699 = v_12696 & ~v_7851;
assign v_12700 = v_12696 & v_7859 & ~v_7860;
assign v_12701 = v_12696 & v_8562;
assign v_12703 = v_12702 & v_7849 & v_7850 & v_7865 & ~v_7866;
assign v_12705 = v_12704 & v_7872 & ~v_7873 & v_7891;
assign v_12706 = v_12704 & ~v_7874;
assign v_12707 = v_12704 & v_7882 & ~v_7883;
assign v_12708 = v_12704 & v_8570;
assign v_12710 = v_12709 & v_7872 & v_7873 & v_7888 & v_7889;
assign v_12711 = v_12704 & v_7872 & ~v_7873 & ~v_7891;
assign v_12712 = v_12709 & v_7872 & v_7873 & v_7888 & ~v_7889;
assign v_12715 = v_12713 & v_12714;
assign v_12716 = v_12713 & v_7895 & v_7896 & ~v_7897 & ~v_7898;
assign v_12717 = v_12713 & v_7895 & v_7896 & v_7897;
assign v_12718 = v_12713 & v_7895 & ~v_7896 & ~v_7900;
assign v_12720 = v_12719 & v_8583;
assign v_12721 = v_12702 & v_7849 & v_7850 & v_7865 & v_7866;
assign v_12722 = v_12694 & v_7826 & v_7827 & v_7842 & v_7843;
assign v_12724 = v_12723 & v_7907 & ~v_7908 & v_7926;
assign v_12725 = v_12723 & v_7907 & ~v_7908 & ~v_7926;
assign v_12726 = v_12723 & ~v_7909;
assign v_12727 = v_12723 & v_7917 & ~v_7918;
assign v_12728 = v_12723 & v_8592;
assign v_12730 = v_12729 & v_7907 & v_7908 & v_7923 & ~v_7924;
assign v_12732 = v_12731 & v_7930 & ~v_7931 & v_7949;
assign v_12733 = v_12731 & v_7930 & ~v_7931 & ~v_7949;
assign v_12734 = v_12731 & ~v_7932;
assign v_12735 = v_12731 & v_7940 & ~v_7941;
assign v_12736 = v_12731 & v_8601;
assign v_12738 = v_12737 & v_7930 & v_7931 & v_7946 & ~v_7947;
assign v_12740 = v_12739 & v_7953 & ~v_7954 & v_7972;
assign v_12741 = v_12739 & ~v_7955;
assign v_12742 = v_12739 & v_7963 & ~v_7964;
assign v_12743 = v_12739 & v_8609;
assign v_12745 = v_12744 & v_7953 & v_7954 & v_7969 & v_7970;
assign v_12746 = v_12739 & v_7953 & ~v_7954 & ~v_7972;
assign v_12747 = v_12744 & v_7953 & v_7954 & v_7969 & ~v_7970;
assign v_12750 = v_12748 & v_12749;
assign v_12751 = v_12748 & v_7976 & v_7977 & ~v_7978 & ~v_7979;
assign v_12752 = v_12748 & v_7976 & v_7977 & v_7978;
assign v_12753 = v_12748 & v_7976 & ~v_7977 & ~v_7981;
assign v_12755 = v_12754 & v_8622;
assign v_12756 = v_12737 & v_7930 & v_7931 & v_7946 & v_7947;
assign v_12757 = v_12729 & v_7907 & v_7908 & v_7923 & v_7924;
assign v_12759 = v_12758 & v_7988 & ~v_7989 & v_8007;
assign v_12760 = v_12758 & v_7988 & ~v_7989 & ~v_8007;
assign v_12761 = v_12758 & ~v_7990;
assign v_12762 = v_12758 & v_7998 & ~v_7999;
assign v_12763 = v_12758 & v_8631;
assign v_12765 = v_12764 & v_7988 & v_7989 & v_8004 & ~v_8005;
assign v_12767 = v_12766 & v_8011 & ~v_8012 & v_8030;
assign v_12768 = v_12766 & v_8011 & ~v_8012 & ~v_8030;
assign v_12769 = v_12766 & ~v_8013;
assign v_12770 = v_12766 & v_8021 & ~v_8022;
assign v_12771 = v_12766 & v_8640;
assign v_12773 = v_12772 & v_8011 & v_8012 & v_8027 & ~v_8028;
assign v_12775 = v_12774 & v_8034 & ~v_8035 & v_8053;
assign v_12776 = v_12774 & ~v_8036;
assign v_12777 = v_12774 & v_8044 & ~v_8045;
assign v_12778 = v_12774 & v_8648;
assign v_12780 = v_12779 & v_8034 & v_8035 & v_8050 & v_8051;
assign v_12781 = v_12774 & v_8034 & ~v_8035 & ~v_8053;
assign v_12782 = v_12779 & v_8034 & v_8035 & v_8050 & ~v_8051;
assign v_12785 = v_12783 & v_12784;
assign v_12786 = v_12783 & v_8057 & v_8058 & ~v_8059 & ~v_8060;
assign v_12787 = v_12783 & v_8057 & v_8058 & v_8059;
assign v_12788 = v_12783 & v_8057 & ~v_8058 & ~v_8062;
assign v_12790 = v_12789 & v_8661;
assign v_12791 = v_12772 & v_8011 & v_8012 & v_8027 & v_8028;
assign v_12792 = v_12764 & v_7988 & v_7989 & v_8004 & v_8005;
assign v_12794 = v_12793 & v_8069 & ~v_8070 & v_8088;
assign v_12795 = v_12793 & v_8069 & ~v_8070 & ~v_8088;
assign v_12796 = v_12793 & ~v_8071;
assign v_12797 = v_12793 & v_8079 & ~v_8080;
assign v_12798 = v_12793 & v_8670;
assign v_12800 = v_12799 & v_8069 & v_8070 & v_8085 & ~v_8086;
assign v_12802 = v_12801 & v_8092 & ~v_8093 & v_8111;
assign v_12803 = v_12801 & v_8092 & ~v_8093 & ~v_8111;
assign v_12804 = v_12801 & ~v_8094;
assign v_12805 = v_12801 & v_8102 & ~v_8103;
assign v_12806 = v_12801 & v_8679;
assign v_12808 = v_12807 & v_8092 & v_8093 & v_8108 & ~v_8109;
assign v_12810 = v_12809 & v_8115 & ~v_8116 & v_8134;
assign v_12811 = v_12809 & ~v_8117;
assign v_12812 = v_12809 & v_8125 & ~v_8126;
assign v_12813 = v_12809 & v_8687;
assign v_12815 = v_12814 & v_8115 & v_8116 & v_8131 & v_8132;
assign v_12816 = v_12809 & v_8115 & ~v_8116 & ~v_8134;
assign v_12817 = v_12814 & v_8115 & v_8116 & v_8131 & ~v_8132;
assign v_12820 = v_12818 & v_12819;
assign v_12821 = v_12818 & v_8138 & v_8139 & ~v_8140 & ~v_8141;
assign v_12822 = v_12818 & v_8138 & v_8139 & v_8140;
assign v_12823 = v_12818 & v_8138 & ~v_8139 & ~v_8143;
assign v_12825 = v_12824 & v_8700;
assign v_12826 = v_12807 & v_8092 & v_8093 & v_8108 & v_8109;
assign v_12827 = v_12799 & v_8069 & v_8070 & v_8085 & v_8086;
assign v_12829 = v_12828 & v_8150 & ~v_8151 & v_8169;
assign v_12830 = v_12828 & v_8150 & ~v_8151 & ~v_8169;
assign v_12831 = v_12828 & ~v_8152;
assign v_12832 = v_12828 & v_8160 & ~v_8161;
assign v_12833 = v_12828 & v_8709;
assign v_12835 = v_12834 & v_8150 & v_8151 & v_8166 & ~v_8167;
assign v_12837 = v_12836 & v_8173 & ~v_8174 & v_8192;
assign v_12838 = v_12836 & v_8173 & ~v_8174 & ~v_8192;
assign v_12839 = v_12836 & ~v_8175;
assign v_12840 = v_12836 & v_8183 & ~v_8184;
assign v_12841 = v_12836 & v_8718;
assign v_12843 = v_12842 & v_8173 & v_8174 & v_8189 & ~v_8190;
assign v_12845 = v_12844 & v_8196 & ~v_8197 & v_8215;
assign v_12846 = v_12844 & ~v_8198;
assign v_12847 = v_12844 & v_8206 & ~v_8207;
assign v_12848 = v_12844 & v_8726;
assign v_12850 = v_12849 & v_8196 & v_8197 & v_8212 & v_8213;
assign v_12851 = v_12844 & v_8196 & ~v_8197 & ~v_8215;
assign v_12852 = v_12849 & v_8196 & v_8197 & v_8212 & ~v_8213;
assign v_12855 = v_12853 & v_12854;
assign v_12856 = v_12853 & v_8219 & v_8220 & ~v_8221 & ~v_8222;
assign v_12857 = v_12853 & v_8219 & v_8220 & v_8221;
assign v_12858 = v_12853 & v_8219 & ~v_8220 & ~v_8224;
assign v_12860 = v_12859 & v_8739;
assign v_12861 = v_12842 & v_8173 & v_8174 & v_8189 & v_8190;
assign v_12862 = v_12834 & v_8150 & v_8151 & v_8166 & v_8167;
assign v_12874 = v_13411 & v_13412 & v_13413;
assign v_12875 = v_232 & ~v_234 & v_236 & ~v_237 & v_239;
assign v_12876 = v_245;
assign v_12877 = v_232 & ~v_234 & v_236 & ~v_237 & v_239;
assign v_12878 = ~v_245 & v_247;
assign v_12879 = v_232 & ~v_234 & ~v_236 & v_241 & ~v_243;
assign v_12880 = v_251;
assign v_12881 = v_232 & ~v_234 & ~v_236 & v_241 & ~v_243;
assign v_12882 = ~v_251;
assign v_12883 = v_232 & ~v_234 & v_236 & ~v_237 & v_239;
assign v_12884 = ~v_245 & ~v_247 & v_258;
assign v_12885 = v_345 & ~v_346 & ~v_348 & ~v_350 & ~v_352;
assign v_12886 = ~v_354;
assign v_12887 = v_372 & ~v_373 & ~v_375 & ~v_377 & ~v_379;
assign v_12888 = v_381;
assign v_12889 = v_372 & ~v_373 & ~v_375 & ~v_377 & ~v_379;
assign v_12890 = ~v_381;
assign v_12891 = v_356 & ~v_357 & v_369 & ~v_370 & v_388;
assign v_12892 = v_389;
assign v_12893 = v_391 & ~v_392 & ~v_394 & ~v_396 & v_398;
assign v_12894 = v_400;
assign v_12895 = v_391 & ~v_392 & ~v_394 & ~v_396 & v_398;
assign v_12896 = ~v_400;
assign v_12897 = v_356 & ~v_357 & v_369 & ~v_370 & v_388;
assign v_12898 = ~v_389 & v_403;
assign v_12899 = v_410 & ~v_411 & ~v_413 & ~v_415 & ~v_417;
assign v_12900 = ~v_419;
assign v_12901 = v_437 & ~v_438 & ~v_440 & ~v_442 & ~v_444;
assign v_12902 = v_446;
assign v_12903 = v_437 & ~v_438 & ~v_440 & ~v_442 & ~v_444;
assign v_12904 = ~v_446;
assign v_12905 = v_421 & ~v_422 & v_434 & ~v_435 & v_453;
assign v_12906 = v_454;
assign v_12907 = v_456 & ~v_457 & ~v_459 & ~v_461 & v_463;
assign v_12908 = v_465;
assign v_12909 = v_456 & ~v_457 & ~v_459 & ~v_461 & v_463;
assign v_12910 = ~v_465;
assign v_12911 = v_421 & ~v_422 & v_434 & ~v_435 & v_453;
assign v_12912 = ~v_454 & v_468;
assign v_12913 = v_496 & ~v_498 & v_500 & ~v_501 & v_503;
assign v_12914 = v_509;
assign v_12915 = v_496 & ~v_498 & v_500 & ~v_501 & v_503;
assign v_12916 = ~v_509 & v_511;
assign v_12917 = v_496 & ~v_498 & ~v_500 & v_505 & ~v_507;
assign v_12918 = v_515;
assign v_12919 = v_496 & ~v_498 & ~v_500 & v_505 & ~v_507;
assign v_12920 = ~v_515;
assign v_12921 = v_496 & ~v_498 & v_500 & ~v_501 & v_503;
assign v_12922 = ~v_509 & ~v_511 & v_522;
assign v_12923 = v_705 & v_722 & v_723 & v_724 & ~v_726;
assign v_12924 = v_729;
assign v_12925 = v_705 & v_722 & v_723 & v_724 & ~v_726;
assign v_12926 = ~v_729 & ~v_731;
assign v_12927 = v_705 & v_722 & v_723 & v_724 & ~v_726;
assign v_12928 = ~v_729 & v_731 & ~v_733;
assign v_12929 = v_705 & v_722 & v_723 & v_724 & ~v_726;
assign v_12930 = ~v_729 & v_731 & v_733 & v_735;
assign v_12931 = v_258 & v_232 & ~v_234 & v_236 & ~v_237;
assign v_12932 = v_239 & ~v_245 & ~v_247;
assign v_12933 = v_1587 & v_372 & ~v_373 & ~v_375 & ~v_377;
assign v_12934 = ~v_379 & ~v_381;
assign v_12935 = v_1601 & v_356 & ~v_357 & v_369 & ~v_370;
assign v_12936 = v_388 & v_389;
assign v_12937 = v_1608 & v_356 & ~v_357 & v_369 & ~v_370;
assign v_12938 = v_388 & ~v_389 & v_403;
assign v_12939 = v_1626 & v_437 & ~v_438 & ~v_440 & ~v_442;
assign v_12940 = ~v_444 & ~v_446;
assign v_12941 = v_1640 & v_421 & ~v_422 & v_434 & ~v_435;
assign v_12942 = v_453 & v_454;
assign v_12943 = v_1647 & v_421 & ~v_422 & v_434 & ~v_435;
assign v_12944 = v_453 & ~v_454 & v_468;
assign v_12945 = v_1663 & v_496 & ~v_498 & v_500 & ~v_501;
assign v_12946 = v_503 & ~v_509 & ~v_511 & v_522;
assign v_12947 = v_1725 & v_669 & v_670 & v_672 & ~v_674;
assign v_12948 = ~v_675;
assign v_12949 = v_1725 & v_669 & v_670 & v_672 & ~v_674;
assign v_12950 = v_675;
assign v_12951 = v_1749 & v_705 & v_722 & v_723 & v_724;
assign v_12952 = v_726;
assign v_12953 = v_2159 & v_372 & ~v_373 & ~v_375 & ~v_377;
assign v_12954 = ~v_379 & ~v_381;
assign v_12955 = v_2172 & v_356 & ~v_357 & v_369 & ~v_370;
assign v_12956 = v_388 & v_389;
assign v_12957 = v_2178 & v_356 & ~v_357 & v_369 & ~v_370;
assign v_12958 = v_388 & ~v_389 & v_403;
assign v_12959 = v_2193 & v_437 & ~v_438 & ~v_440 & ~v_442;
assign v_12960 = ~v_444 & ~v_446;
assign v_12961 = v_2206 & v_421 & ~v_422 & v_434 & ~v_435;
assign v_12962 = v_453 & v_454;
assign v_12963 = v_2212 & v_421 & ~v_422 & v_434 & ~v_435;
assign v_12964 = v_453 & ~v_454 & v_468;
assign v_12965 = v_2267 & v_669 & v_670 & v_672 & ~v_674;
assign v_12966 = ~v_675;
assign v_12967 = v_2267 & v_669 & v_670 & v_672 & ~v_674;
assign v_12968 = v_675;
assign v_12969 = v_2288 & v_705 & v_722 & v_723 & v_724;
assign v_12970 = v_726;
assign v_12971 = v_2626 & v_232 & ~v_234 & v_236 & ~v_237;
assign v_12972 = v_239 & ~v_245 & ~v_247 & v_258;
assign v_12973 = v_2667 & v_372 & ~v_373 & ~v_375 & ~v_377;
assign v_12974 = ~v_379 & ~v_381;
assign v_12975 = v_2680 & v_356 & ~v_357 & v_369 & ~v_370;
assign v_12976 = v_388 & v_389;
assign v_12977 = v_2686 & v_356 & ~v_357 & v_369 & ~v_370;
assign v_12978 = v_388 & ~v_389 & v_403;
assign v_12979 = v_2701 & v_437 & ~v_438 & ~v_440 & ~v_442;
assign v_12980 = ~v_444 & ~v_446;
assign v_12981 = v_2714 & v_421 & ~v_422 & v_434 & ~v_435;
assign v_12982 = v_453 & v_454;
assign v_12983 = v_2720 & v_421 & ~v_422 & v_434 & ~v_435;
assign v_12984 = v_453 & ~v_454 & v_468;
assign v_12985 = v_2731 & v_496 & ~v_498 & v_500 & ~v_501;
assign v_12986 = v_503 & ~v_509 & ~v_511 & v_522;
assign v_12987 = v_2794 & v_669 & v_670 & v_672 & ~v_674;
assign v_12988 = ~v_675;
assign v_12989 = v_2794 & v_669 & v_670 & v_672 & ~v_674;
assign v_12990 = v_675;
assign v_12991 = v_2819 & v_705 & v_722 & v_723 & v_724;
assign v_12992 = v_726;
assign v_12993 = v_258 & v_232 & ~v_234 & v_236 & ~v_237;
assign v_12994 = v_239 & ~v_245 & ~v_247;
assign v_12995 = v_3200 & v_372 & ~v_373 & ~v_375 & ~v_377;
assign v_12996 = ~v_379 & ~v_381;
assign v_12997 = v_3213 & v_356 & ~v_357 & v_369 & ~v_370;
assign v_12998 = v_388 & v_389;
assign v_12999 = v_3219 & v_356 & ~v_357 & v_369 & ~v_370;
assign v_13000 = v_388 & ~v_389 & v_403;
assign v_13001 = v_3234 & v_437 & ~v_438 & ~v_440 & ~v_442;
assign v_13002 = ~v_444 & ~v_446;
assign v_13003 = v_3247 & v_421 & ~v_422 & v_434 & ~v_435;
assign v_13004 = v_453 & v_454;
assign v_13005 = v_3253 & v_421 & ~v_422 & v_434 & ~v_435;
assign v_13006 = v_453 & ~v_454 & v_468;
assign v_13007 = v_3264 & v_496 & ~v_498 & v_500 & ~v_501;
assign v_13008 = v_503 & ~v_509 & ~v_511 & v_522;
assign v_13009 = v_3327 & v_669 & v_670 & v_672 & ~v_674;
assign v_13010 = ~v_675;
assign v_13011 = v_3327 & v_669 & v_670 & v_672 & ~v_674;
assign v_13012 = v_675;
assign v_13013 = v_3352 & v_705 & v_722 & v_723 & v_724;
assign v_13014 = v_726;
assign v_13015 = v_3695 & v_232 & ~v_234 & v_236 & ~v_237;
assign v_13016 = v_239 & ~v_245 & ~v_247 & v_258;
assign v_13017 = v_3736 & v_372 & ~v_373 & ~v_375 & ~v_377;
assign v_13018 = ~v_379 & ~v_381;
assign v_13019 = v_3749 & v_356 & ~v_357 & v_369 & ~v_370;
assign v_13020 = v_388 & v_389;
assign v_13021 = v_3755 & v_356 & ~v_357 & v_369 & ~v_370;
assign v_13022 = v_388 & ~v_389 & v_403;
assign v_13023 = v_3770 & v_437 & ~v_438 & ~v_440 & ~v_442;
assign v_13024 = ~v_444 & ~v_446;
assign v_13025 = v_3783 & v_421 & ~v_422 & v_434 & ~v_435;
assign v_13026 = v_453 & v_454;
assign v_13027 = v_3789 & v_421 & ~v_422 & v_434 & ~v_435;
assign v_13028 = v_453 & ~v_454 & v_468;
assign v_13029 = v_3800 & v_496 & ~v_498 & v_500 & ~v_501;
assign v_13030 = v_503 & ~v_509 & ~v_511 & v_522;
assign v_13031 = v_3863 & v_669 & v_670 & v_672 & ~v_674;
assign v_13032 = ~v_675;
assign v_13033 = v_3863 & v_669 & v_670 & v_672 & ~v_674;
assign v_13034 = v_675;
assign v_13035 = v_3888 & v_705 & v_722 & v_723 & v_724;
assign v_13036 = v_726;
assign v_13037 = v_4231 & v_232 & ~v_234 & v_236 & ~v_237;
assign v_13038 = v_239 & ~v_245 & ~v_247 & v_258;
assign v_13039 = v_4272 & v_372 & ~v_373 & ~v_375 & ~v_377;
assign v_13040 = ~v_379 & ~v_381;
assign v_13041 = v_4285 & v_356 & ~v_357 & v_369 & ~v_370;
assign v_13042 = v_388 & v_389;
assign v_13043 = v_4291 & v_356 & ~v_357 & v_369 & ~v_370;
assign v_13044 = v_388 & ~v_389 & v_403;
assign v_13045 = v_4306 & v_437 & ~v_438 & ~v_440 & ~v_442;
assign v_13046 = ~v_444 & ~v_446;
assign v_13047 = v_4319 & v_421 & ~v_422 & v_434 & ~v_435;
assign v_13048 = v_453 & v_454;
assign v_13049 = v_4325 & v_421 & ~v_422 & v_434 & ~v_435;
assign v_13050 = v_453 & ~v_454 & v_468;
assign v_13051 = v_4336 & v_496 & ~v_498 & v_500 & ~v_501;
assign v_13052 = v_503 & ~v_509 & ~v_511 & v_522;
assign v_13053 = v_4399 & v_669 & v_670 & v_672 & ~v_674;
assign v_13054 = ~v_675;
assign v_13055 = v_4399 & v_669 & v_670 & v_672 & ~v_674;
assign v_13056 = v_675;
assign v_13057 = v_4424 & v_705 & v_722 & v_723 & v_724;
assign v_13058 = v_726;
assign v_13059 = v_4766 & v_232 & ~v_234 & v_236 & ~v_237;
assign v_13060 = v_239 & ~v_245 & ~v_247 & v_258;
assign v_13061 = v_4807 & v_372 & ~v_373 & ~v_375 & ~v_377;
assign v_13062 = ~v_379 & ~v_381;
assign v_13063 = v_4820 & v_356 & ~v_357 & v_369 & ~v_370;
assign v_13064 = v_388 & v_389;
assign v_13065 = v_4826 & v_356 & ~v_357 & v_369 & ~v_370;
assign v_13066 = v_388 & ~v_389 & v_403;
assign v_13067 = v_4841 & v_437 & ~v_438 & ~v_440 & ~v_442;
assign v_13068 = ~v_444 & ~v_446;
assign v_13069 = v_4854 & v_421 & ~v_422 & v_434 & ~v_435;
assign v_13070 = v_453 & v_454;
assign v_13071 = v_4860 & v_421 & ~v_422 & v_434 & ~v_435;
assign v_13072 = v_453 & ~v_454 & v_468;
assign v_13073 = v_4871 & v_496 & ~v_498 & v_500 & ~v_501;
assign v_13074 = v_503 & ~v_509 & ~v_511 & v_522;
assign v_13075 = v_4934 & v_669 & v_670 & v_672 & ~v_674;
assign v_13076 = ~v_675;
assign v_13077 = v_4934 & v_669 & v_670 & v_672 & ~v_674;
assign v_13078 = v_675;
assign v_13079 = v_4959 & v_705 & v_722 & v_723 & v_724;
assign v_13080 = v_726;
assign v_13081 = v_5302 & v_232 & ~v_234 & v_236 & ~v_237;
assign v_13082 = v_239 & ~v_245 & ~v_247 & v_258;
assign v_13083 = v_5343 & v_372 & ~v_373 & ~v_375 & ~v_377;
assign v_13084 = ~v_379 & ~v_381;
assign v_13085 = v_5356 & v_356 & ~v_357 & v_369 & ~v_370;
assign v_13086 = v_388 & v_389;
assign v_13087 = v_5362 & v_356 & ~v_357 & v_369 & ~v_370;
assign v_13088 = v_388 & ~v_389 & v_403;
assign v_13089 = v_5377 & v_437 & ~v_438 & ~v_440 & ~v_442;
assign v_13090 = ~v_444 & ~v_446;
assign v_13091 = v_5390 & v_421 & ~v_422 & v_434 & ~v_435;
assign v_13092 = v_453 & v_454;
assign v_13093 = v_5396 & v_421 & ~v_422 & v_434 & ~v_435;
assign v_13094 = v_453 & ~v_454 & v_468;
assign v_13095 = v_5407 & v_496 & ~v_498 & v_500 & ~v_501;
assign v_13096 = v_503 & ~v_509 & ~v_511 & v_522;
assign v_13097 = v_5470 & v_669 & v_670 & v_672 & ~v_674;
assign v_13098 = ~v_675;
assign v_13099 = v_5470 & v_669 & v_670 & v_672 & ~v_674;
assign v_13100 = v_675;
assign v_13101 = v_5495 & v_705 & v_722 & v_723 & v_724;
assign v_13102 = v_726;
assign v_13103 = v_5872 & v_372 & ~v_373 & ~v_375 & ~v_377;
assign v_13104 = ~v_379 & ~v_381;
assign v_13105 = v_5885 & v_356 & ~v_357 & v_369 & ~v_370;
assign v_13106 = v_388 & v_389;
assign v_13107 = v_5891 & v_356 & ~v_357 & v_369 & ~v_370;
assign v_13108 = v_388 & ~v_389 & v_403;
assign v_13109 = v_5906 & v_437 & ~v_438 & ~v_440 & ~v_442;
assign v_13110 = ~v_444 & ~v_446;
assign v_13111 = v_5919 & v_421 & ~v_422 & v_434 & ~v_435;
assign v_13112 = v_453 & v_454;
assign v_13113 = v_5925 & v_421 & ~v_422 & v_434 & ~v_435;
assign v_13114 = v_453 & ~v_454 & v_468;
assign v_13115 = v_5979 & v_669 & v_670 & v_672 & ~v_674;
assign v_13116 = ~v_675;
assign v_13117 = v_5979 & v_669 & v_670 & v_672 & ~v_674;
assign v_13118 = v_675;
assign v_13119 = v_6000 & v_705 & v_722 & v_723 & v_724;
assign v_13120 = v_726;
assign v_13121 = v_6339 & v_232 & ~v_234 & v_236 & ~v_237;
assign v_13122 = v_239 & ~v_245 & ~v_247 & v_258;
assign v_13123 = v_6380 & v_372 & ~v_373 & ~v_375 & ~v_377;
assign v_13124 = ~v_379 & ~v_381;
assign v_13125 = v_6393 & v_356 & ~v_357 & v_369 & ~v_370;
assign v_13126 = v_388 & v_389;
assign v_13127 = v_6399 & v_356 & ~v_357 & v_369 & ~v_370;
assign v_13128 = v_388 & ~v_389 & v_403;
assign v_13129 = v_6414 & v_437 & ~v_438 & ~v_440 & ~v_442;
assign v_13130 = ~v_444 & ~v_446;
assign v_13131 = v_6427 & v_421 & ~v_422 & v_434 & ~v_435;
assign v_13132 = v_453 & v_454;
assign v_13133 = v_6433 & v_421 & ~v_422 & v_434 & ~v_435;
assign v_13134 = v_453 & ~v_454 & v_468;
assign v_13135 = v_6444 & v_496 & ~v_498 & v_500 & ~v_501;
assign v_13136 = v_503 & ~v_509 & ~v_511 & v_522;
assign v_13137 = v_6507 & v_669 & v_670 & v_672 & ~v_674;
assign v_13138 = ~v_675;
assign v_13139 = v_6507 & v_669 & v_670 & v_672 & ~v_674;
assign v_13140 = v_675;
assign v_13141 = v_6532 & v_705 & v_722 & v_723 & v_724;
assign v_13142 = v_726;
assign v_13143 = v_7098 & ~v_7100 & v_7102 & ~v_7103 & v_7105;
assign v_13144 = v_7111;
assign v_13145 = v_7098 & ~v_7100 & v_7102 & ~v_7103 & v_7105;
assign v_13146 = ~v_7111 & v_7113;
assign v_13147 = v_7098 & ~v_7100 & ~v_7102 & v_7107 & ~v_7109;
assign v_13148 = v_7117;
assign v_13149 = v_7098 & ~v_7100 & ~v_7102 & v_7107 & ~v_7109;
assign v_13150 = ~v_7117;
assign v_13151 = v_7098 & ~v_7100 & v_7102 & ~v_7103 & v_7105;
assign v_13152 = ~v_7111 & ~v_7113 & v_7124;
assign v_13153 = v_7211 & ~v_7212 & ~v_7214 & ~v_7216 & ~v_7218;
assign v_13154 = ~v_7220;
assign v_13155 = v_7238 & ~v_7239 & ~v_7241 & ~v_7243 & ~v_7245;
assign v_13156 = v_7247;
assign v_13157 = v_7238 & ~v_7239 & ~v_7241 & ~v_7243 & ~v_7245;
assign v_13158 = ~v_7247;
assign v_13159 = v_7222 & ~v_7223 & v_7235 & ~v_7236 & v_7254;
assign v_13160 = v_7255;
assign v_13161 = v_7257 & ~v_7258 & ~v_7260 & ~v_7262 & v_7264;
assign v_13162 = v_7266;
assign v_13163 = v_7257 & ~v_7258 & ~v_7260 & ~v_7262 & v_7264;
assign v_13164 = ~v_7266;
assign v_13165 = v_7222 & ~v_7223 & v_7235 & ~v_7236 & v_7254;
assign v_13166 = ~v_7255 & v_7269;
assign v_13167 = v_7276 & ~v_7277 & ~v_7279 & ~v_7281 & ~v_7283;
assign v_13168 = ~v_7285;
assign v_13169 = v_7303 & ~v_7304 & ~v_7306 & ~v_7308 & ~v_7310;
assign v_13170 = v_7312;
assign v_13171 = v_7303 & ~v_7304 & ~v_7306 & ~v_7308 & ~v_7310;
assign v_13172 = ~v_7312;
assign v_13173 = v_7287 & ~v_7288 & v_7300 & ~v_7301 & v_7319;
assign v_13174 = v_7320;
assign v_13175 = v_7322 & ~v_7323 & ~v_7325 & ~v_7327 & v_7329;
assign v_13176 = v_7331;
assign v_13177 = v_7322 & ~v_7323 & ~v_7325 & ~v_7327 & v_7329;
assign v_13178 = ~v_7331;
assign v_13179 = v_7287 & ~v_7288 & v_7300 & ~v_7301 & v_7319;
assign v_13180 = ~v_7320 & v_7334;
assign v_13181 = v_7362 & ~v_7364 & v_7366 & ~v_7367 & v_7369;
assign v_13182 = v_7375;
assign v_13183 = v_7362 & ~v_7364 & v_7366 & ~v_7367 & v_7369;
assign v_13184 = ~v_7375 & v_7377;
assign v_13185 = v_7362 & ~v_7364 & ~v_7366 & v_7371 & ~v_7373;
assign v_13186 = v_7381;
assign v_13187 = v_7362 & ~v_7364 & ~v_7366 & v_7371 & ~v_7373;
assign v_13188 = ~v_7381;
assign v_13189 = v_7362 & ~v_7364 & v_7366 & ~v_7367 & v_7369;
assign v_13190 = ~v_7375 & ~v_7377 & v_7388;
assign v_13191 = v_7571 & v_7588 & v_7589 & v_7590 & ~v_7592;
assign v_13192 = v_7595;
assign v_13193 = v_7571 & v_7588 & v_7589 & v_7590 & ~v_7592;
assign v_13194 = ~v_7595 & ~v_7597;
assign v_13195 = v_7571 & v_7588 & v_7589 & v_7590 & ~v_7592;
assign v_13196 = ~v_7595 & v_7597 & ~v_7599;
assign v_13197 = v_7571 & v_7588 & v_7589 & v_7590 & ~v_7592;
assign v_13198 = ~v_7595 & v_7597 & v_7599 & v_7601;
assign v_13199 = v_7124 & v_7098 & ~v_7100 & v_7102 & ~v_7103;
assign v_13200 = v_7105 & ~v_7111 & ~v_7113;
assign v_13201 = v_8291 & v_7238 & ~v_7239 & ~v_7241 & ~v_7243;
assign v_13202 = ~v_7245 & ~v_7247;
assign v_13203 = v_8305 & v_7222 & ~v_7223 & v_7235 & ~v_7236;
assign v_13204 = v_7254 & v_7255;
assign v_13205 = v_8312 & v_7222 & ~v_7223 & v_7235 & ~v_7236;
assign v_13206 = v_7254 & ~v_7255 & v_7269;
assign v_13207 = v_8330 & v_7303 & ~v_7304 & ~v_7306 & ~v_7308;
assign v_13208 = ~v_7310 & ~v_7312;
assign v_13209 = v_8344 & v_7287 & ~v_7288 & v_7300 & ~v_7301;
assign v_13210 = v_7319 & v_7320;
assign v_13211 = v_8351 & v_7287 & ~v_7288 & v_7300 & ~v_7301;
assign v_13212 = v_7319 & ~v_7320 & v_7334;
assign v_13213 = v_8367 & v_7362 & ~v_7364 & v_7366 & ~v_7367;
assign v_13214 = v_7369 & ~v_7375 & ~v_7377 & v_7388;
assign v_13215 = v_8429 & v_7535 & v_7536 & v_7538 & ~v_7540;
assign v_13216 = ~v_7541;
assign v_13217 = v_8429 & v_7535 & v_7536 & v_7538 & ~v_7540;
assign v_13218 = v_7541;
assign v_13219 = v_8453 & v_7571 & v_7588 & v_7589 & v_7590;
assign v_13220 = v_7592;
assign v_13221 = v_8785 & v_7238 & ~v_7239 & ~v_7241 & ~v_7243;
assign v_13222 = ~v_7245 & ~v_7247;
assign v_13223 = v_8798 & v_7222 & ~v_7223 & v_7235 & ~v_7236;
assign v_13224 = v_7254 & v_7255;
assign v_13225 = v_8804 & v_7222 & ~v_7223 & v_7235 & ~v_7236;
assign v_13226 = v_7254 & ~v_7255 & v_7269;
assign v_13227 = v_8819 & v_7303 & ~v_7304 & ~v_7306 & ~v_7308;
assign v_13228 = ~v_7310 & ~v_7312;
assign v_13229 = v_8832 & v_7287 & ~v_7288 & v_7300 & ~v_7301;
assign v_13230 = v_7319 & v_7320;
assign v_13231 = v_8838 & v_7287 & ~v_7288 & v_7300 & ~v_7301;
assign v_13232 = v_7319 & ~v_7320 & v_7334;
assign v_13233 = v_8893 & v_7535 & v_7536 & v_7538 & ~v_7540;
assign v_13234 = ~v_7541;
assign v_13235 = v_8893 & v_7535 & v_7536 & v_7538 & ~v_7540;
assign v_13236 = v_7541;
assign v_13237 = v_8914 & v_7571 & v_7588 & v_7589 & v_7590;
assign v_13238 = v_7592;
assign v_13239 = v_9182 & v_7098 & ~v_7100 & v_7102 & ~v_7103;
assign v_13240 = v_7105 & ~v_7111 & ~v_7113 & v_7124;
assign v_13241 = v_9223 & v_7238 & ~v_7239 & ~v_7241 & ~v_7243;
assign v_13242 = ~v_7245 & ~v_7247;
assign v_13243 = v_9236 & v_7222 & ~v_7223 & v_7235 & ~v_7236;
assign v_13244 = v_7254 & v_7255;
assign v_13245 = v_9242 & v_7222 & ~v_7223 & v_7235 & ~v_7236;
assign v_13246 = v_7254 & ~v_7255 & v_7269;
assign v_13247 = v_9257 & v_7303 & ~v_7304 & ~v_7306 & ~v_7308;
assign v_13248 = ~v_7310 & ~v_7312;
assign v_13249 = v_9270 & v_7287 & ~v_7288 & v_7300 & ~v_7301;
assign v_13250 = v_7319 & v_7320;
assign v_13251 = v_9276 & v_7287 & ~v_7288 & v_7300 & ~v_7301;
assign v_13252 = v_7319 & ~v_7320 & v_7334;
assign v_13253 = v_9287 & v_7362 & ~v_7364 & v_7366 & ~v_7367;
assign v_13254 = v_7369 & ~v_7375 & ~v_7377 & v_7388;
assign v_13255 = v_9350 & v_7535 & v_7536 & v_7538 & ~v_7540;
assign v_13256 = ~v_7541;
assign v_13257 = v_9350 & v_7535 & v_7536 & v_7538 & ~v_7540;
assign v_13258 = v_7541;
assign v_13259 = v_9375 & v_7571 & v_7588 & v_7589 & v_7590;
assign v_13260 = v_7592;
assign v_13261 = v_7124 & v_7098 & ~v_7100 & v_7102 & ~v_7103;
assign v_13262 = v_7105 & ~v_7111 & ~v_7113;
assign v_13263 = v_9686 & v_7238 & ~v_7239 & ~v_7241 & ~v_7243;
assign v_13264 = ~v_7245 & ~v_7247;
assign v_13265 = v_9699 & v_7222 & ~v_7223 & v_7235 & ~v_7236;
assign v_13266 = v_7254 & v_7255;
assign v_13267 = v_9705 & v_7222 & ~v_7223 & v_7235 & ~v_7236;
assign v_13268 = v_7254 & ~v_7255 & v_7269;
assign v_13269 = v_9720 & v_7303 & ~v_7304 & ~v_7306 & ~v_7308;
assign v_13270 = ~v_7310 & ~v_7312;
assign v_13271 = v_9733 & v_7287 & ~v_7288 & v_7300 & ~v_7301;
assign v_13272 = v_7319 & v_7320;
assign v_13273 = v_9739 & v_7287 & ~v_7288 & v_7300 & ~v_7301;
assign v_13274 = v_7319 & ~v_7320 & v_7334;
assign v_13275 = v_9750 & v_7362 & ~v_7364 & v_7366 & ~v_7367;
assign v_13276 = v_7369 & ~v_7375 & ~v_7377 & v_7388;
assign v_13277 = v_9813 & v_7535 & v_7536 & v_7538 & ~v_7540;
assign v_13278 = ~v_7541;
assign v_13279 = v_9813 & v_7535 & v_7536 & v_7538 & ~v_7540;
assign v_13280 = v_7541;
assign v_13281 = v_9838 & v_7571 & v_7588 & v_7589 & v_7590;
assign v_13282 = v_7592;
assign v_13283 = v_10111 & v_7098 & ~v_7100 & v_7102 & ~v_7103;
assign v_13284 = v_7105 & ~v_7111 & ~v_7113 & v_7124;
assign v_13285 = v_10152 & v_7238 & ~v_7239 & ~v_7241 & ~v_7243;
assign v_13286 = ~v_7245 & ~v_7247;
assign v_13287 = v_10165 & v_7222 & ~v_7223 & v_7235 & ~v_7236;
assign v_13288 = v_7254 & v_7255;
assign v_13289 = v_10171 & v_7222 & ~v_7223 & v_7235 & ~v_7236;
assign v_13290 = v_7254 & ~v_7255 & v_7269;
assign v_13291 = v_10186 & v_7303 & ~v_7304 & ~v_7306 & ~v_7308;
assign v_13292 = ~v_7310 & ~v_7312;
assign v_13293 = v_10199 & v_7287 & ~v_7288 & v_7300 & ~v_7301;
assign v_13294 = v_7319 & v_7320;
assign v_13295 = v_10205 & v_7287 & ~v_7288 & v_7300 & ~v_7301;
assign v_13296 = v_7319 & ~v_7320 & v_7334;
assign v_13297 = v_10216 & v_7362 & ~v_7364 & v_7366 & ~v_7367;
assign v_13298 = v_7369 & ~v_7375 & ~v_7377 & v_7388;
assign v_13299 = v_10279 & v_7535 & v_7536 & v_7538 & ~v_7540;
assign v_13300 = ~v_7541;
assign v_13301 = v_10279 & v_7535 & v_7536 & v_7538 & ~v_7540;
assign v_13302 = v_7541;
assign v_13303 = v_10304 & v_7571 & v_7588 & v_7589 & v_7590;
assign v_13304 = v_7592;
assign v_13305 = v_10577 & v_7098 & ~v_7100 & v_7102 & ~v_7103;
assign v_13306 = v_7105 & ~v_7111 & ~v_7113 & v_7124;
assign v_13307 = v_10618 & v_7238 & ~v_7239 & ~v_7241 & ~v_7243;
assign v_13308 = ~v_7245 & ~v_7247;
assign v_13309 = v_10631 & v_7222 & ~v_7223 & v_7235 & ~v_7236;
assign v_13310 = v_7254 & v_7255;
assign v_13311 = v_10637 & v_7222 & ~v_7223 & v_7235 & ~v_7236;
assign v_13312 = v_7254 & ~v_7255 & v_7269;
assign v_13313 = v_10652 & v_7303 & ~v_7304 & ~v_7306 & ~v_7308;
assign v_13314 = ~v_7310 & ~v_7312;
assign v_13315 = v_10665 & v_7287 & ~v_7288 & v_7300 & ~v_7301;
assign v_13316 = v_7319 & v_7320;
assign v_13317 = v_10671 & v_7287 & ~v_7288 & v_7300 & ~v_7301;
assign v_13318 = v_7319 & ~v_7320 & v_7334;
assign v_13319 = v_10682 & v_7362 & ~v_7364 & v_7366 & ~v_7367;
assign v_13320 = v_7369 & ~v_7375 & ~v_7377 & v_7388;
assign v_13321 = v_10745 & v_7535 & v_7536 & v_7538 & ~v_7540;
assign v_13322 = ~v_7541;
assign v_13323 = v_10745 & v_7535 & v_7536 & v_7538 & ~v_7540;
assign v_13324 = v_7541;
assign v_13325 = v_10770 & v_7571 & v_7588 & v_7589 & v_7590;
assign v_13326 = v_7592;
assign v_13327 = v_11042 & v_7098 & ~v_7100 & v_7102 & ~v_7103;
assign v_13328 = v_7105 & ~v_7111 & ~v_7113 & v_7124;
assign v_13329 = v_11083 & v_7238 & ~v_7239 & ~v_7241 & ~v_7243;
assign v_13330 = ~v_7245 & ~v_7247;
assign v_13331 = v_11096 & v_7222 & ~v_7223 & v_7235 & ~v_7236;
assign v_13332 = v_7254 & v_7255;
assign v_13333 = v_11102 & v_7222 & ~v_7223 & v_7235 & ~v_7236;
assign v_13334 = v_7254 & ~v_7255 & v_7269;
assign v_13335 = v_11117 & v_7303 & ~v_7304 & ~v_7306 & ~v_7308;
assign v_13336 = ~v_7310 & ~v_7312;
assign v_13337 = v_11130 & v_7287 & ~v_7288 & v_7300 & ~v_7301;
assign v_13338 = v_7319 & v_7320;
assign v_13339 = v_11136 & v_7287 & ~v_7288 & v_7300 & ~v_7301;
assign v_13340 = v_7319 & ~v_7320 & v_7334;
assign v_13341 = v_11147 & v_7362 & ~v_7364 & v_7366 & ~v_7367;
assign v_13342 = v_7369 & ~v_7375 & ~v_7377 & v_7388;
assign v_13343 = v_11210 & v_7535 & v_7536 & v_7538 & ~v_7540;
assign v_13344 = ~v_7541;
assign v_13345 = v_11210 & v_7535 & v_7536 & v_7538 & ~v_7540;
assign v_13346 = v_7541;
assign v_13347 = v_11235 & v_7571 & v_7588 & v_7589 & v_7590;
assign v_13348 = v_7592;
assign v_13349 = v_11508 & v_7098 & ~v_7100 & v_7102 & ~v_7103;
assign v_13350 = v_7105 & ~v_7111 & ~v_7113 & v_7124;
assign v_13351 = v_11549 & v_7238 & ~v_7239 & ~v_7241 & ~v_7243;
assign v_13352 = ~v_7245 & ~v_7247;
assign v_13353 = v_11562 & v_7222 & ~v_7223 & v_7235 & ~v_7236;
assign v_13354 = v_7254 & v_7255;
assign v_13355 = v_11568 & v_7222 & ~v_7223 & v_7235 & ~v_7236;
assign v_13356 = v_7254 & ~v_7255 & v_7269;
assign v_13357 = v_11583 & v_7303 & ~v_7304 & ~v_7306 & ~v_7308;
assign v_13358 = ~v_7310 & ~v_7312;
assign v_13359 = v_11596 & v_7287 & ~v_7288 & v_7300 & ~v_7301;
assign v_13360 = v_7319 & v_7320;
assign v_13361 = v_11602 & v_7287 & ~v_7288 & v_7300 & ~v_7301;
assign v_13362 = v_7319 & ~v_7320 & v_7334;
assign v_13363 = v_11613 & v_7362 & ~v_7364 & v_7366 & ~v_7367;
assign v_13364 = v_7369 & ~v_7375 & ~v_7377 & v_7388;
assign v_13365 = v_11676 & v_7535 & v_7536 & v_7538 & ~v_7540;
assign v_13366 = ~v_7541;
assign v_13367 = v_11676 & v_7535 & v_7536 & v_7538 & ~v_7540;
assign v_13368 = v_7541;
assign v_13369 = v_11701 & v_7571 & v_7588 & v_7589 & v_7590;
assign v_13370 = v_7592;
assign v_13371 = v_12008 & v_7238 & ~v_7239 & ~v_7241 & ~v_7243;
assign v_13372 = ~v_7245 & ~v_7247;
assign v_13373 = v_12021 & v_7222 & ~v_7223 & v_7235 & ~v_7236;
assign v_13374 = v_7254 & v_7255;
assign v_13375 = v_12027 & v_7222 & ~v_7223 & v_7235 & ~v_7236;
assign v_13376 = v_7254 & ~v_7255 & v_7269;
assign v_13377 = v_12042 & v_7303 & ~v_7304 & ~v_7306 & ~v_7308;
assign v_13378 = ~v_7310 & ~v_7312;
assign v_13379 = v_12055 & v_7287 & ~v_7288 & v_7300 & ~v_7301;
assign v_13380 = v_7319 & v_7320;
assign v_13381 = v_12061 & v_7287 & ~v_7288 & v_7300 & ~v_7301;
assign v_13382 = v_7319 & ~v_7320 & v_7334;
assign v_13383 = v_12115 & v_7535 & v_7536 & v_7538 & ~v_7540;
assign v_13384 = ~v_7541;
assign v_13385 = v_12115 & v_7535 & v_7536 & v_7538 & ~v_7540;
assign v_13386 = v_7541;
assign v_13387 = v_12136 & v_7571 & v_7588 & v_7589 & v_7590;
assign v_13388 = v_7592;
assign v_13389 = v_12405 & v_7098 & ~v_7100 & v_7102 & ~v_7103;
assign v_13390 = v_7105 & ~v_7111 & ~v_7113 & v_7124;
assign v_13391 = v_12446 & v_7238 & ~v_7239 & ~v_7241 & ~v_7243;
assign v_13392 = ~v_7245 & ~v_7247;
assign v_13393 = v_12459 & v_7222 & ~v_7223 & v_7235 & ~v_7236;
assign v_13394 = v_7254 & v_7255;
assign v_13395 = v_12465 & v_7222 & ~v_7223 & v_7235 & ~v_7236;
assign v_13396 = v_7254 & ~v_7255 & v_7269;
assign v_13397 = v_12480 & v_7303 & ~v_7304 & ~v_7306 & ~v_7308;
assign v_13398 = ~v_7310 & ~v_7312;
assign v_13399 = v_12493 & v_7287 & ~v_7288 & v_7300 & ~v_7301;
assign v_13400 = v_7319 & v_7320;
assign v_13401 = v_12499 & v_7287 & ~v_7288 & v_7300 & ~v_7301;
assign v_13402 = v_7319 & ~v_7320 & v_7334;
assign v_13403 = v_12510 & v_7362 & ~v_7364 & v_7366 & ~v_7367;
assign v_13404 = v_7369 & ~v_7375 & ~v_7377 & v_7388;
assign v_13405 = v_12573 & v_7535 & v_7536 & v_7538 & ~v_7540;
assign v_13406 = ~v_7541;
assign v_13407 = v_12573 & v_7535 & v_7536 & v_7538 & ~v_7540;
assign v_13408 = v_7541;
assign v_13409 = v_12598 & v_7571 & v_7588 & v_7589 & v_7590;
assign v_13410 = v_7592;
assign v_13411 = ~v_12864 & ~v_12865 & ~v_12866 & ~v_12867 & ~v_12868;
assign v_13412 = ~v_12869 & ~v_12870 & ~v_12871 & ~v_12872 & ~v_12873;
assign v_13413 = v_8230;
assign v_217 = ~v_213 | v_215 | v_216;
assign v_224 = v_222 | v_223;
assign v_258 = ~v_254 | v_256 | v_257;
assign v_260 = v_13414 | v_13415 | v_13416;
assign v_267 = v_261 | v_263 | v_265 | v_266;
assign v_271 = v_228 | v_269 | v_270;
assign v_277 = v_275 | v_276;
assign v_285 = v_282 | v_284;
assign v_291 = ~v_280 | v_287 | v_289 | v_290;
assign v_300 = v_297 | v_299;
assign v_302 = ~v_279 | v_294 | v_296 | v_301;
assign v_306 = v_304 | v_305;
assign v_315 = ~v_311 | v_313 | v_314;
assign v_321 = v_317 | v_319 | v_320;
assign v_329 = v_323 | v_325 | v_327 | v_328;
assign v_331 = v_308 | v_310 | v_330;
assign v_343 = ~v_333 | v_335 | v_337 | v_341 | v_342;
assign v_356 = v_353 | v_355;
assign v_369 = v_361 | v_363 | v_365 | v_367 | v_368;
assign v_384 = v_380 | v_382 | v_383;
assign v_388 = v_374 | v_376 | v_378 | v_386 | v_387;
assign v_403 = v_13417 | v_13418;
assign v_405 = v_371 | v_390 | v_404;
assign v_409 = v_13419 | v_13420;
assign v_421 = v_418 | v_420;
assign v_434 = v_426 | v_428 | v_430 | v_432 | v_433;
assign v_449 = v_445 | v_447 | v_448;
assign v_453 = v_439 | v_441 | v_443 | v_451 | v_452;
assign v_468 = v_13421 | v_13422;
assign v_470 = v_436 | v_455 | v_469;
assign v_474 = v_13423 | v_13424;
assign v_480 = v_476 | v_478 | v_479;
assign v_484 = v_482 | v_483;
assign v_522 = ~v_518 | v_520 | v_521;
assign v_524 = v_13425 | v_13426 | v_13427;
assign v_531 = v_525 | v_527 | v_529 | v_530;
assign v_535 = v_492 | v_533 | v_534;
assign v_541 = v_539 | v_540;
assign v_546 = ~v_542 | v_544 | v_545;
assign v_554 = v_552 | v_553;
assign v_558 = v_548 | v_557;
assign v_568 = v_562 | v_566 | v_567;
assign v_577 = ~v_573 | v_575 | v_576;
assign v_581 = v_560 | v_570 | v_572 | v_579 | v_580;
assign v_588 = v_585 | v_587;
assign v_593 = v_590 | v_592;
assign v_598 = v_595 | v_583 | v_596 | v_597;
assign v_604 = ~v_600 | v_602 | v_603;
assign v_612 = v_610 | v_611;
assign v_616 = v_606 | v_615;
assign v_626 = v_620 | v_624 | v_625;
assign v_635 = ~v_631 | v_633 | v_634;
assign v_639 = v_618 | v_628 | v_630 | v_637 | v_638;
assign v_652 = v_650 | v_651;
assign v_654 = v_648 | v_653;
assign v_656 = v_646 | v_655;
assign v_658 = v_644 | v_657;
assign v_660 = v_642 | v_659;
assign v_662 = v_640 | v_661;
assign v_679 = v_677 | v_678;
assign v_689 = v_686 | v_688;
assign v_694 = v_691 | v_693;
assign v_699 = v_696 | v_684 | v_697 | v_698;
assign v_703 = v_13428 | v_13429;
assign v_710 = ~v_706 | v_708 | v_709;
assign v_718 = v_716 | v_717;
assign v_722 = v_712 | v_721;
assign v_737 = v_734 | v_736;
assign v_745 = v_740 | v_741 | v_743 | v_744;
assign v_750 = ~v_746 | v_748 | v_749;
assign v_758 = v_752 | v_757;
assign v_763 = ~v_759 | v_761 | v_762;
assign v_771 = v_765 | v_770;
assign v_779 = ~v_775 | v_777 | v_778;
assign v_787 = v_785 | v_786;
assign v_791 = v_781 | v_790;
assign v_796 = v_13430 | v_13431;
assign v_804 = v_802 | v_803;
assign v_808 = v_806 | v_807;
assign v_814 = ~v_800 | v_810 | v_812 | v_813;
assign v_821 = v_819 | v_820;
assign v_827 = v_825 | v_826;
assign v_831 = v_829 | v_830;
assign v_837 = ~v_823 | v_833 | v_835 | v_836;
assign v_844 = v_842 | v_843;
assign v_850 = v_848 | v_849;
assign v_854 = v_852 | v_853;
assign v_860 = ~v_846 | v_856 | v_858 | v_859;
assign v_867 = v_865 | v_866;
assign v_877 = v_13432 | v_13433 | v_13434;
assign v_885 = v_883 | v_884;
assign v_889 = v_887 | v_888;
assign v_895 = ~v_881 | v_891 | v_893 | v_894;
assign v_902 = v_900 | v_901;
assign v_908 = v_906 | v_907;
assign v_912 = v_910 | v_911;
assign v_918 = ~v_904 | v_914 | v_916 | v_917;
assign v_925 = v_923 | v_924;
assign v_931 = v_929 | v_930;
assign v_935 = v_933 | v_934;
assign v_941 = ~v_927 | v_937 | v_939 | v_940;
assign v_948 = v_946 | v_947;
assign v_958 = v_13435 | v_13436 | v_13437;
assign v_966 = v_964 | v_965;
assign v_970 = v_968 | v_969;
assign v_976 = ~v_962 | v_972 | v_974 | v_975;
assign v_983 = v_981 | v_982;
assign v_989 = v_987 | v_988;
assign v_993 = v_991 | v_992;
assign v_999 = ~v_985 | v_995 | v_997 | v_998;
assign v_1006 = v_1004 | v_1005;
assign v_1012 = v_1010 | v_1011;
assign v_1016 = v_1014 | v_1015;
assign v_1022 = ~v_1008 | v_1018 | v_1020 | v_1021;
assign v_1029 = v_1027 | v_1028;
assign v_1039 = v_13438 | v_13439 | v_13440;
assign v_1047 = v_1045 | v_1046;
assign v_1051 = v_1049 | v_1050;
assign v_1057 = ~v_1043 | v_1053 | v_1055 | v_1056;
assign v_1064 = v_1062 | v_1063;
assign v_1070 = v_1068 | v_1069;
assign v_1074 = v_1072 | v_1073;
assign v_1080 = ~v_1066 | v_1076 | v_1078 | v_1079;
assign v_1087 = v_1085 | v_1086;
assign v_1093 = v_1091 | v_1092;
assign v_1097 = v_1095 | v_1096;
assign v_1103 = ~v_1089 | v_1099 | v_1101 | v_1102;
assign v_1110 = v_1108 | v_1109;
assign v_1120 = v_13441 | v_13442 | v_13443;
assign v_1128 = v_1126 | v_1127;
assign v_1132 = v_1130 | v_1131;
assign v_1138 = ~v_1124 | v_1134 | v_1136 | v_1137;
assign v_1145 = v_1143 | v_1144;
assign v_1151 = v_1149 | v_1150;
assign v_1155 = v_1153 | v_1154;
assign v_1161 = ~v_1147 | v_1157 | v_1159 | v_1160;
assign v_1168 = v_1166 | v_1167;
assign v_1174 = v_1172 | v_1173;
assign v_1178 = v_1176 | v_1177;
assign v_1184 = ~v_1170 | v_1180 | v_1182 | v_1183;
assign v_1191 = v_1189 | v_1190;
assign v_1201 = v_13444 | v_13445 | v_13446;
assign v_1209 = v_1207 | v_1208;
assign v_1213 = v_1211 | v_1212;
assign v_1219 = ~v_1205 | v_1215 | v_1217 | v_1218;
assign v_1226 = v_1224 | v_1225;
assign v_1232 = v_1230 | v_1231;
assign v_1236 = v_1234 | v_1235;
assign v_1242 = ~v_1228 | v_1238 | v_1240 | v_1241;
assign v_1249 = v_1247 | v_1248;
assign v_1255 = v_1253 | v_1254;
assign v_1259 = v_1257 | v_1258;
assign v_1265 = ~v_1251 | v_1261 | v_1263 | v_1264;
assign v_1272 = v_1270 | v_1271;
assign v_1282 = v_13447 | v_13448 | v_13449;
assign v_1290 = v_1288 | v_1289;
assign v_1294 = v_1292 | v_1293;
assign v_1300 = ~v_1286 | v_1296 | v_1298 | v_1299;
assign v_1307 = v_1305 | v_1306;
assign v_1313 = v_1311 | v_1312;
assign v_1317 = v_1315 | v_1316;
assign v_1323 = ~v_1309 | v_1319 | v_1321 | v_1322;
assign v_1330 = v_1328 | v_1329;
assign v_1336 = v_1334 | v_1335;
assign v_1340 = v_1338 | v_1339;
assign v_1346 = ~v_1332 | v_1342 | v_1344 | v_1345;
assign v_1353 = v_1351 | v_1352;
assign v_1363 = v_13450 | v_13451 | v_13452;
assign v_1371 = v_1369 | v_1370;
assign v_1375 = v_1373 | v_1374;
assign v_1381 = ~v_1367 | v_1377 | v_1379 | v_1380;
assign v_1388 = v_1386 | v_1387;
assign v_1394 = v_1392 | v_1393;
assign v_1398 = v_1396 | v_1397;
assign v_1404 = ~v_1390 | v_1400 | v_1402 | v_1403;
assign v_1411 = v_1409 | v_1410;
assign v_1417 = v_1415 | v_1416;
assign v_1421 = v_1419 | v_1420;
assign v_1427 = ~v_1413 | v_1423 | v_1425 | v_1426;
assign v_1434 = v_1432 | v_1433;
assign v_1444 = v_13453 | v_13454 | v_13455;
assign v_1452 = v_1450 | v_1451;
assign v_1456 = v_1454 | v_1455;
assign v_1462 = ~v_1448 | v_1458 | v_1460 | v_1461;
assign v_1469 = v_1467 | v_1468;
assign v_1475 = v_1473 | v_1474;
assign v_1479 = v_1477 | v_1478;
assign v_1485 = ~v_1471 | v_1481 | v_1483 | v_1484;
assign v_1492 = v_1490 | v_1491;
assign v_1498 = v_1496 | v_1497;
assign v_1502 = v_1500 | v_1501;
assign v_1508 = ~v_1494 | v_1504 | v_1506 | v_1507;
assign v_1515 = v_1513 | v_1514;
assign v_1525 = v_13456 | v_13457 | v_13458;
assign v_1531 = v_1530 | ~v_1529;
assign v_1538 = v_13459 | v_13460;
assign v_1540 = v_252 | v_253;
assign v_1543 = v_1539 | v_1541 | v_1542;
assign v_1545 = v_1534 | v_1535 | v_1536 | v_1544;
assign v_1547 = v_1546 | ~v_1545;
assign v_1550 = v_1548 | v_1549;
assign v_1552 = v_294 | v_296;
assign v_1555 = v_1551 | v_1553 | v_1554;
assign v_1556 = v_308 | v_310;
assign v_1562 = v_1559 | v_1560 | v_1561;
assign v_1563 = v_325 | v_327 | v_328;
assign v_1565 = v_1558 | v_1564;
assign v_1567 = v_1557 | v_1566;
assign v_1568 = ~v_333 | v_335 | v_337;
assign v_1570 = v_341 | v_342;
assign v_1572 = v_1569 | v_1571;
assign v_1574 = v_1532 | v_1573;
assign v_1582 = v_367 | v_368;
assign v_1584 = v_1581 | v_1583;
assign v_1585 = v_365 | v_367 | v_368;
assign v_1587 = v_1579 | v_1580 | v_1586;
assign v_1592 = v_380 | v_382;
assign v_1595 = v_1593 | v_1594;
assign v_1598 = v_1596 | v_1597;
assign v_1599 = v_386 | v_387;
assign v_1601 = v_1589 | v_1590 | v_1591 | v_1600;
assign v_1606 = v_399 | v_401 | v_402;
assign v_1608 = v_1603 | v_1604 | v_1605 | v_1607;
assign v_1610 = v_1588 | v_1602 | v_1609;
assign v_1611 = v_407 | v_408;
assign v_1613 = v_1575 | v_1576 | v_1577 | v_1578 | v_1612;
assign v_1621 = v_432 | v_433;
assign v_1623 = v_1620 | v_1622;
assign v_1624 = v_430 | v_432 | v_433;
assign v_1626 = v_1618 | v_1619 | v_1625;
assign v_1631 = v_445 | v_447;
assign v_1634 = v_1632 | v_1633;
assign v_1637 = v_1635 | v_1636;
assign v_1638 = v_451 | v_452;
assign v_1640 = v_1628 | v_1629 | v_1630 | v_1639;
assign v_1645 = v_464 | v_466 | v_467;
assign v_1647 = v_1642 | v_1643 | v_1644 | v_1646;
assign v_1649 = v_1627 | v_1641 | v_1648;
assign v_1650 = v_472 | v_473;
assign v_1652 = v_1614 | v_1615 | v_1616 | v_1617 | v_1651;
assign v_1657 = v_1656 | ~v_1652;
assign v_1663 = v_1661 | v_1662;
assign v_1664 = v_13461 | v_13462;
assign v_1666 = v_516 | v_517;
assign v_1669 = v_1665 | v_1667 | v_1668;
assign v_1671 = v_1658 | v_1659 | v_1660 | v_1670;
assign v_1673 = v_1672 | ~v_1671;
assign v_1676 = v_1653 | v_1674 | v_1675;
assign v_1679 = v_1677 | v_1678;
assign v_1682 = v_566 | v_567;
assign v_1684 = v_1681 | v_1683;
assign v_1685 = v_570 | v_572;
assign v_1687 = v_579 | v_580;
assign v_1689 = v_1680 | v_1686 | v_1688;
assign v_1694 = v_1690 | v_1691 | v_1692 | v_1693;
assign v_1697 = v_1695 | v_1696;
assign v_1700 = v_624 | v_625;
assign v_1702 = v_1699 | v_1701;
assign v_1703 = v_628 | v_630;
assign v_1705 = v_637 | v_638;
assign v_1707 = v_1698 | v_1704 | v_1706;
assign v_1715 = v_1713 | v_1714;
assign v_1717 = v_1712 | v_1716;
assign v_1719 = v_1711 | v_1718;
assign v_1721 = v_1710 | v_1720;
assign v_1723 = v_1709 | v_1722;
assign v_1725 = v_1708 | v_1724;
assign v_1730 = v_1728 | v_1729;
assign v_1736 = v_1732 | v_1733 | v_1734 | v_1735;
assign v_1737 = v_701 | v_702;
assign v_1739 = v_1731 | v_1738;
assign v_1740 = v_683 | v_701 | v_702;
assign v_1743 = v_671 | v_673;
assign v_1745 = v_1726 | v_1727 | v_1741 | v_1742 | v_1744;
assign v_1749 = v_1747 | v_1748;
assign v_1751 = v_730 | v_732;
assign v_1755 = v_1753 | v_1754;
assign v_1758 = v_1756 | v_1757;
assign v_1763 = v_1761 | v_1762;
assign v_1764 = v_793 | v_794;
assign v_1766 = v_13463 | v_13464;
assign v_1771 = v_812 | v_813;
assign v_1773 = v_1769 | v_1770 | v_1772;
assign v_1775 = v_1768 | v_1774;
assign v_1780 = v_835 | v_836;
assign v_1782 = v_1778 | v_1779 | v_1781;
assign v_1784 = v_1777 | v_1783;
assign v_1788 = v_858 | v_859;
assign v_1790 = v_1786 | v_1787 | v_1789;
assign v_1794 = v_1792 | v_1793;
assign v_1795 = v_873 | v_871;
assign v_1800 = v_1796 | v_1797 | v_1798 | v_1799;
assign v_1801 = v_871 | v_873 | v_874 | v_875 | v_876;
assign v_1805 = v_13465 | v_13466;
assign v_1810 = v_893 | v_894;
assign v_1812 = v_1808 | v_1809 | v_1811;
assign v_1814 = v_1807 | v_1813;
assign v_1819 = v_916 | v_917;
assign v_1821 = v_1817 | v_1818 | v_1820;
assign v_1823 = v_1816 | v_1822;
assign v_1827 = v_939 | v_940;
assign v_1829 = v_1825 | v_1826 | v_1828;
assign v_1833 = v_1831 | v_1832;
assign v_1834 = v_954 | v_952;
assign v_1839 = v_1835 | v_1836 | v_1837 | v_1838;
assign v_1840 = v_952 | v_954 | v_955 | v_956 | v_957;
assign v_1844 = v_13467 | v_13468;
assign v_1849 = v_974 | v_975;
assign v_1851 = v_1847 | v_1848 | v_1850;
assign v_1853 = v_1846 | v_1852;
assign v_1858 = v_997 | v_998;
assign v_1860 = v_1856 | v_1857 | v_1859;
assign v_1862 = v_1855 | v_1861;
assign v_1866 = v_1020 | v_1021;
assign v_1868 = v_1864 | v_1865 | v_1867;
assign v_1872 = v_1870 | v_1871;
assign v_1873 = v_1035 | v_1033;
assign v_1878 = v_1874 | v_1875 | v_1876 | v_1877;
assign v_1879 = v_1033 | v_1035 | v_1036 | v_1037 | v_1038;
assign v_1883 = v_13469 | v_13470;
assign v_1888 = v_1055 | v_1056;
assign v_1890 = v_1886 | v_1887 | v_1889;
assign v_1892 = v_1885 | v_1891;
assign v_1897 = v_1078 | v_1079;
assign v_1899 = v_1895 | v_1896 | v_1898;
assign v_1901 = v_1894 | v_1900;
assign v_1905 = v_1101 | v_1102;
assign v_1907 = v_1903 | v_1904 | v_1906;
assign v_1911 = v_1909 | v_1910;
assign v_1912 = v_1116 | v_1114;
assign v_1917 = v_1913 | v_1914 | v_1915 | v_1916;
assign v_1918 = v_1114 | v_1116 | v_1117 | v_1118 | v_1119;
assign v_1922 = v_13471 | v_13472;
assign v_1927 = v_1136 | v_1137;
assign v_1929 = v_1925 | v_1926 | v_1928;
assign v_1931 = v_1924 | v_1930;
assign v_1936 = v_1159 | v_1160;
assign v_1938 = v_1934 | v_1935 | v_1937;
assign v_1940 = v_1933 | v_1939;
assign v_1944 = v_1182 | v_1183;
assign v_1946 = v_1942 | v_1943 | v_1945;
assign v_1950 = v_1948 | v_1949;
assign v_1951 = v_1197 | v_1195;
assign v_1956 = v_1952 | v_1953 | v_1954 | v_1955;
assign v_1957 = v_1195 | v_1197 | v_1198 | v_1199 | v_1200;
assign v_1961 = v_13473 | v_13474;
assign v_1966 = v_1217 | v_1218;
assign v_1968 = v_1964 | v_1965 | v_1967;
assign v_1970 = v_1963 | v_1969;
assign v_1975 = v_1240 | v_1241;
assign v_1977 = v_1973 | v_1974 | v_1976;
assign v_1979 = v_1972 | v_1978;
assign v_1983 = v_1263 | v_1264;
assign v_1985 = v_1981 | v_1982 | v_1984;
assign v_1989 = v_1987 | v_1988;
assign v_1990 = v_1278 | v_1276;
assign v_1995 = v_1991 | v_1992 | v_1993 | v_1994;
assign v_1996 = v_1276 | v_1278 | v_1279 | v_1280 | v_1281;
assign v_2000 = v_13475 | v_13476;
assign v_2005 = v_1298 | v_1299;
assign v_2007 = v_2003 | v_2004 | v_2006;
assign v_2009 = v_2002 | v_2008;
assign v_2014 = v_1321 | v_1322;
assign v_2016 = v_2012 | v_2013 | v_2015;
assign v_2018 = v_2011 | v_2017;
assign v_2022 = v_1344 | v_1345;
assign v_2024 = v_2020 | v_2021 | v_2023;
assign v_2028 = v_2026 | v_2027;
assign v_2029 = v_1359 | v_1357;
assign v_2034 = v_2030 | v_2031 | v_2032 | v_2033;
assign v_2035 = v_1357 | v_1359 | v_1360 | v_1361 | v_1362;
assign v_2039 = v_13477 | v_13478;
assign v_2044 = v_1379 | v_1380;
assign v_2046 = v_2042 | v_2043 | v_2045;
assign v_2048 = v_2041 | v_2047;
assign v_2053 = v_1402 | v_1403;
assign v_2055 = v_2051 | v_2052 | v_2054;
assign v_2057 = v_2050 | v_2056;
assign v_2061 = v_1425 | v_1426;
assign v_2063 = v_2059 | v_2060 | v_2062;
assign v_2067 = v_2065 | v_2066;
assign v_2068 = v_1440 | v_1438;
assign v_2073 = v_2069 | v_2070 | v_2071 | v_2072;
assign v_2074 = v_1438 | v_1440 | v_1441 | v_1442 | v_1443;
assign v_2078 = v_13479 | v_13480;
assign v_2083 = v_1460 | v_1461;
assign v_2085 = v_2081 | v_2082 | v_2084;
assign v_2087 = v_2080 | v_2086;
assign v_2092 = v_1483 | v_1484;
assign v_2094 = v_2090 | v_2091 | v_2093;
assign v_2096 = v_2089 | v_2095;
assign v_2100 = v_1506 | v_1507;
assign v_2102 = v_2098 | v_2099 | v_2101;
assign v_2106 = v_2104 | v_2105;
assign v_2107 = v_1521 | v_1519;
assign v_2112 = v_2108 | v_2109 | v_2110 | v_2111;
assign v_2113 = v_1519 | v_1521 | v_1522 | v_1523 | v_1524;
assign v_2117 = v_13481 | v_13482;
assign v_2119 = v_2118 | v_1529;
assign v_2123 = v_2122 | v_1545;
assign v_2126 = v_2121 | v_2124 | v_2125;
assign v_2128 = v_294 | v_296;
assign v_2131 = v_2127 | v_2129 | v_2130;
assign v_2132 = v_308 | v_310;
assign v_2138 = v_2135 | v_2136 | v_2137;
assign v_2140 = v_2134 | v_2139;
assign v_2142 = v_2133 | v_2141;
assign v_2143 = ~v_333 | v_335 | v_337;
assign v_2146 = v_2144 | v_2145;
assign v_2148 = v_2120 | v_2147;
assign v_2157 = v_2155 | v_2156;
assign v_2159 = v_2153 | v_2154 | v_2158;
assign v_2164 = v_380 | v_382;
assign v_2167 = v_2165 | v_2166;
assign v_2170 = v_2168 | v_2169;
assign v_2172 = v_2161 | v_2162 | v_2163 | v_2171;
assign v_2178 = v_2174 | v_2175 | v_2176 | v_2177;
assign v_2180 = v_2160 | v_2173 | v_2179;
assign v_2182 = v_2149 | v_2150 | v_2151 | v_2152 | v_2181;
assign v_2191 = v_2189 | v_2190;
assign v_2193 = v_2187 | v_2188 | v_2192;
assign v_2198 = v_445 | v_447;
assign v_2201 = v_2199 | v_2200;
assign v_2204 = v_2202 | v_2203;
assign v_2206 = v_2195 | v_2196 | v_2197 | v_2205;
assign v_2212 = v_2208 | v_2209 | v_2210 | v_2211;
assign v_2214 = v_2194 | v_2207 | v_2213;
assign v_2216 = v_2183 | v_2184 | v_2185 | v_2186 | v_2215;
assign v_2219 = v_2218 | v_1671;
assign v_2222 = v_2217 | v_2220 | v_2221;
assign v_2225 = v_2223 | v_2224;
assign v_2229 = v_2227 | v_2228;
assign v_2230 = v_570 | v_572;
assign v_2233 = v_2226 | v_2231 | v_2232;
assign v_2238 = v_2234 | v_2235 | v_2236 | v_2237;
assign v_2241 = v_2239 | v_2240;
assign v_2245 = v_2243 | v_2244;
assign v_2246 = v_628 | v_630;
assign v_2249 = v_2242 | v_2247 | v_2248;
assign v_2257 = v_2255 | v_2256;
assign v_2259 = v_2254 | v_2258;
assign v_2261 = v_2253 | v_2260;
assign v_2263 = v_2252 | v_2262;
assign v_2265 = v_2251 | v_2264;
assign v_2267 = v_2250 | v_2266;
assign v_2272 = v_2270 | v_2271;
assign v_2278 = v_2274 | v_2275 | v_2276 | v_2277;
assign v_2280 = v_2273 | v_2279;
assign v_2284 = v_2268 | v_2269 | v_2281 | v_2282 | v_2283;
assign v_2288 = v_2286 | v_2287;
assign v_2290 = v_730 | v_732;
assign v_2294 = v_2292 | v_2293;
assign v_2297 = v_2295 | v_2296;
assign v_2302 = v_2300 | v_2301;
assign v_2304 = v_13483 | v_13484;
assign v_2310 = v_2307 | v_2308 | v_2309;
assign v_2312 = v_2306 | v_2311;
assign v_2318 = v_2315 | v_2316 | v_2317;
assign v_2320 = v_2314 | v_2319;
assign v_2325 = v_2322 | v_2323 | v_2324;
assign v_2329 = v_2327 | v_2328;
assign v_2330 = v_873 | v_871;
assign v_2335 = v_2331 | v_2332 | v_2333 | v_2334;
assign v_2339 = v_13485 | v_13486;
assign v_2345 = v_2342 | v_2343 | v_2344;
assign v_2347 = v_2341 | v_2346;
assign v_2353 = v_2350 | v_2351 | v_2352;
assign v_2355 = v_2349 | v_2354;
assign v_2360 = v_2357 | v_2358 | v_2359;
assign v_2364 = v_2362 | v_2363;
assign v_2365 = v_954 | v_952;
assign v_2370 = v_2366 | v_2367 | v_2368 | v_2369;
assign v_2374 = v_13487 | v_13488;
assign v_2380 = v_2377 | v_2378 | v_2379;
assign v_2382 = v_2376 | v_2381;
assign v_2388 = v_2385 | v_2386 | v_2387;
assign v_2390 = v_2384 | v_2389;
assign v_2395 = v_2392 | v_2393 | v_2394;
assign v_2399 = v_2397 | v_2398;
assign v_2400 = v_1035 | v_1033;
assign v_2405 = v_2401 | v_2402 | v_2403 | v_2404;
assign v_2409 = v_13489 | v_13490;
assign v_2415 = v_2412 | v_2413 | v_2414;
assign v_2417 = v_2411 | v_2416;
assign v_2423 = v_2420 | v_2421 | v_2422;
assign v_2425 = v_2419 | v_2424;
assign v_2430 = v_2427 | v_2428 | v_2429;
assign v_2434 = v_2432 | v_2433;
assign v_2435 = v_1116 | v_1114;
assign v_2440 = v_2436 | v_2437 | v_2438 | v_2439;
assign v_2444 = v_13491 | v_13492;
assign v_2450 = v_2447 | v_2448 | v_2449;
assign v_2452 = v_2446 | v_2451;
assign v_2458 = v_2455 | v_2456 | v_2457;
assign v_2460 = v_2454 | v_2459;
assign v_2465 = v_2462 | v_2463 | v_2464;
assign v_2469 = v_2467 | v_2468;
assign v_2470 = v_1197 | v_1195;
assign v_2475 = v_2471 | v_2472 | v_2473 | v_2474;
assign v_2479 = v_13493 | v_13494;
assign v_2485 = v_2482 | v_2483 | v_2484;
assign v_2487 = v_2481 | v_2486;
assign v_2493 = v_2490 | v_2491 | v_2492;
assign v_2495 = v_2489 | v_2494;
assign v_2500 = v_2497 | v_2498 | v_2499;
assign v_2504 = v_2502 | v_2503;
assign v_2505 = v_1278 | v_1276;
assign v_2510 = v_2506 | v_2507 | v_2508 | v_2509;
assign v_2514 = v_13495 | v_13496;
assign v_2520 = v_2517 | v_2518 | v_2519;
assign v_2522 = v_2516 | v_2521;
assign v_2528 = v_2525 | v_2526 | v_2527;
assign v_2530 = v_2524 | v_2529;
assign v_2535 = v_2532 | v_2533 | v_2534;
assign v_2539 = v_2537 | v_2538;
assign v_2540 = v_1359 | v_1357;
assign v_2545 = v_2541 | v_2542 | v_2543 | v_2544;
assign v_2549 = v_13497 | v_13498;
assign v_2555 = v_2552 | v_2553 | v_2554;
assign v_2557 = v_2551 | v_2556;
assign v_2563 = v_2560 | v_2561 | v_2562;
assign v_2565 = v_2559 | v_2564;
assign v_2570 = v_2567 | v_2568 | v_2569;
assign v_2574 = v_2572 | v_2573;
assign v_2575 = v_1440 | v_1438;
assign v_2580 = v_2576 | v_2577 | v_2578 | v_2579;
assign v_2584 = v_13499 | v_13500;
assign v_2590 = v_2587 | v_2588 | v_2589;
assign v_2592 = v_2586 | v_2591;
assign v_2598 = v_2595 | v_2596 | v_2597;
assign v_2600 = v_2594 | v_2599;
assign v_2605 = v_2602 | v_2603 | v_2604;
assign v_2609 = v_2607 | v_2608;
assign v_2610 = v_1521 | v_1519;
assign v_2615 = v_2611 | v_2612 | v_2613 | v_2614;
assign v_2619 = v_13501 | v_13502;
assign v_2626 = v_2624 | v_2625;
assign v_2627 = v_13503 | v_13504;
assign v_2631 = v_2628 | v_2629 | v_2630;
assign v_2633 = v_2621 | v_2622 | v_2623 | v_2632;
assign v_2636 = v_2620 | v_2634 | v_2635;
assign v_2638 = v_294 | v_296;
assign v_2641 = v_2637 | v_2639 | v_2640;
assign v_2642 = v_308 | v_310;
assign v_2648 = v_2645 | v_2646 | v_2647;
assign v_2650 = v_2644 | v_2649;
assign v_2652 = v_2643 | v_2651;
assign v_2653 = ~v_333 | v_335 | v_337;
assign v_2656 = v_2654 | v_2655;
assign v_2665 = v_2663 | v_2664;
assign v_2667 = v_2661 | v_2662 | v_2666;
assign v_2672 = v_380 | v_382;
assign v_2675 = v_2673 | v_2674;
assign v_2678 = v_2676 | v_2677;
assign v_2680 = v_2669 | v_2670 | v_2671 | v_2679;
assign v_2686 = v_2682 | v_2683 | v_2684 | v_2685;
assign v_2688 = v_2668 | v_2681 | v_2687;
assign v_2690 = v_2657 | v_2658 | v_2659 | v_2660 | v_2689;
assign v_2699 = v_2697 | v_2698;
assign v_2701 = v_2695 | v_2696 | v_2700;
assign v_2706 = v_445 | v_447;
assign v_2709 = v_2707 | v_2708;
assign v_2712 = v_2710 | v_2711;
assign v_2714 = v_2703 | v_2704 | v_2705 | v_2713;
assign v_2720 = v_2716 | v_2717 | v_2718 | v_2719;
assign v_2722 = v_2702 | v_2715 | v_2721;
assign v_2724 = v_2691 | v_2692 | v_2693 | v_2694 | v_2723;
assign v_2731 = v_2729 | v_2730;
assign v_2732 = v_13505 | v_13506;
assign v_2736 = v_2733 | v_2734 | v_2735;
assign v_2738 = v_2726 | v_2727 | v_2728 | v_2737;
assign v_2741 = v_2725 | v_2739 | v_2740;
assign v_2746 = v_2743 | v_2745;
assign v_2748 = v_2742 | v_2747;
assign v_2752 = v_2750 | v_2751;
assign v_2753 = v_570 | v_572;
assign v_2756 = v_2749 | v_2754 | v_2755;
assign v_2761 = v_2757 | v_2758 | v_2759 | v_2760;
assign v_2766 = v_2763 | v_2765;
assign v_2768 = v_2762 | v_2767;
assign v_2772 = v_2770 | v_2771;
assign v_2773 = v_628 | v_630;
assign v_2776 = v_2769 | v_2774 | v_2775;
assign v_2784 = v_2782 | v_2783;
assign v_2786 = v_2781 | v_2785;
assign v_2788 = v_2780 | v_2787;
assign v_2790 = v_2779 | v_2789;
assign v_2792 = v_2778 | v_2791;
assign v_2794 = v_2777 | v_2793;
assign v_2799 = v_2797 | v_2798;
assign v_2805 = v_2801 | v_2802 | v_2803 | v_2804;
assign v_2807 = v_2800 | v_2806;
assign v_2811 = v_2795 | v_2796 | v_2808 | v_2809 | v_2810;
assign v_2817 = v_2814 | v_2816;
assign v_2819 = v_2813 | v_2818;
assign v_2821 = v_730 | v_732;
assign v_2825 = v_2823 | v_2824;
assign v_2828 = v_2826 | v_2827;
assign v_2835 = v_2832 | v_2834;
assign v_2837 = v_2831 | v_2836;
assign v_2839 = v_13507 | v_13508;
assign v_2845 = v_2842 | v_2843 | v_2844;
assign v_2847 = v_2841 | v_2846;
assign v_2853 = v_2850 | v_2851 | v_2852;
assign v_2855 = v_2849 | v_2854;
assign v_2860 = v_2857 | v_2858 | v_2859;
assign v_2864 = v_2862 | v_2863;
assign v_2865 = v_873 | v_871;
assign v_2870 = v_2866 | v_2867 | v_2868 | v_2869;
assign v_2874 = v_13509 | v_13510;
assign v_2880 = v_2877 | v_2878 | v_2879;
assign v_2882 = v_2876 | v_2881;
assign v_2888 = v_2885 | v_2886 | v_2887;
assign v_2890 = v_2884 | v_2889;
assign v_2895 = v_2892 | v_2893 | v_2894;
assign v_2899 = v_2897 | v_2898;
assign v_2900 = v_954 | v_952;
assign v_2905 = v_2901 | v_2902 | v_2903 | v_2904;
assign v_2909 = v_13511 | v_13512;
assign v_2915 = v_2912 | v_2913 | v_2914;
assign v_2917 = v_2911 | v_2916;
assign v_2923 = v_2920 | v_2921 | v_2922;
assign v_2925 = v_2919 | v_2924;
assign v_2930 = v_2927 | v_2928 | v_2929;
assign v_2934 = v_2932 | v_2933;
assign v_2935 = v_1035 | v_1033;
assign v_2940 = v_2936 | v_2937 | v_2938 | v_2939;
assign v_2944 = v_13513 | v_13514;
assign v_2950 = v_2947 | v_2948 | v_2949;
assign v_2952 = v_2946 | v_2951;
assign v_2958 = v_2955 | v_2956 | v_2957;
assign v_2960 = v_2954 | v_2959;
assign v_2965 = v_2962 | v_2963 | v_2964;
assign v_2969 = v_2967 | v_2968;
assign v_2970 = v_1116 | v_1114;
assign v_2975 = v_2971 | v_2972 | v_2973 | v_2974;
assign v_2979 = v_13515 | v_13516;
assign v_2985 = v_2982 | v_2983 | v_2984;
assign v_2987 = v_2981 | v_2986;
assign v_2993 = v_2990 | v_2991 | v_2992;
assign v_2995 = v_2989 | v_2994;
assign v_3000 = v_2997 | v_2998 | v_2999;
assign v_3004 = v_3002 | v_3003;
assign v_3005 = v_1197 | v_1195;
assign v_3010 = v_3006 | v_3007 | v_3008 | v_3009;
assign v_3014 = v_13517 | v_13518;
assign v_3020 = v_3017 | v_3018 | v_3019;
assign v_3022 = v_3016 | v_3021;
assign v_3028 = v_3025 | v_3026 | v_3027;
assign v_3030 = v_3024 | v_3029;
assign v_3035 = v_3032 | v_3033 | v_3034;
assign v_3039 = v_3037 | v_3038;
assign v_3040 = v_1278 | v_1276;
assign v_3045 = v_3041 | v_3042 | v_3043 | v_3044;
assign v_3049 = v_13519 | v_13520;
assign v_3055 = v_3052 | v_3053 | v_3054;
assign v_3057 = v_3051 | v_3056;
assign v_3063 = v_3060 | v_3061 | v_3062;
assign v_3065 = v_3059 | v_3064;
assign v_3070 = v_3067 | v_3068 | v_3069;
assign v_3074 = v_3072 | v_3073;
assign v_3075 = v_1359 | v_1357;
assign v_3080 = v_3076 | v_3077 | v_3078 | v_3079;
assign v_3084 = v_13521 | v_13522;
assign v_3090 = v_3087 | v_3088 | v_3089;
assign v_3092 = v_3086 | v_3091;
assign v_3098 = v_3095 | v_3096 | v_3097;
assign v_3100 = v_3094 | v_3099;
assign v_3105 = v_3102 | v_3103 | v_3104;
assign v_3109 = v_3107 | v_3108;
assign v_3110 = v_1440 | v_1438;
assign v_3115 = v_3111 | v_3112 | v_3113 | v_3114;
assign v_3119 = v_13523 | v_13524;
assign v_3125 = v_3122 | v_3123 | v_3124;
assign v_3127 = v_3121 | v_3126;
assign v_3133 = v_3130 | v_3131 | v_3132;
assign v_3135 = v_3129 | v_3134;
assign v_3140 = v_3137 | v_3138 | v_3139;
assign v_3144 = v_3142 | v_3143;
assign v_3145 = v_1521 | v_1519;
assign v_3150 = v_3146 | v_3147 | v_3148 | v_3149;
assign v_3154 = v_13525 | v_13526;
assign v_3160 = v_13527 | v_13528;
assign v_3164 = v_3161 | v_3162 | v_3163;
assign v_3166 = v_3156 | v_3157 | v_3158 | v_3165;
assign v_3169 = v_3155 | v_3167 | v_3168;
assign v_3171 = v_294 | v_296;
assign v_3174 = v_3170 | v_3172 | v_3173;
assign v_3175 = v_308 | v_310;
assign v_3181 = v_3178 | v_3179 | v_3180;
assign v_3183 = v_3177 | v_3182;
assign v_3185 = v_3176 | v_3184;
assign v_3186 = ~v_333 | v_335 | v_337;
assign v_3189 = v_3187 | v_3188;
assign v_3198 = v_3196 | v_3197;
assign v_3200 = v_3194 | v_3195 | v_3199;
assign v_3205 = v_380 | v_382;
assign v_3208 = v_3206 | v_3207;
assign v_3211 = v_3209 | v_3210;
assign v_3213 = v_3202 | v_3203 | v_3204 | v_3212;
assign v_3219 = v_3215 | v_3216 | v_3217 | v_3218;
assign v_3221 = v_3201 | v_3214 | v_3220;
assign v_3223 = v_3190 | v_3191 | v_3192 | v_3193 | v_3222;
assign v_3232 = v_3230 | v_3231;
assign v_3234 = v_3228 | v_3229 | v_3233;
assign v_3239 = v_445 | v_447;
assign v_3242 = v_3240 | v_3241;
assign v_3245 = v_3243 | v_3244;
assign v_3247 = v_3236 | v_3237 | v_3238 | v_3246;
assign v_3253 = v_3249 | v_3250 | v_3251 | v_3252;
assign v_3255 = v_3235 | v_3248 | v_3254;
assign v_3257 = v_3224 | v_3225 | v_3226 | v_3227 | v_3256;
assign v_3264 = v_3262 | v_3263;
assign v_3265 = v_13529 | v_13530;
assign v_3269 = v_3266 | v_3267 | v_3268;
assign v_3271 = v_3259 | v_3260 | v_3261 | v_3270;
assign v_3274 = v_3258 | v_3272 | v_3273;
assign v_3279 = v_3276 | v_3278;
assign v_3281 = v_3275 | v_3280;
assign v_3285 = v_3283 | v_3284;
assign v_3286 = v_570 | v_572;
assign v_3289 = v_3282 | v_3287 | v_3288;
assign v_3294 = v_3290 | v_3291 | v_3292 | v_3293;
assign v_3299 = v_3296 | v_3298;
assign v_3301 = v_3295 | v_3300;
assign v_3305 = v_3303 | v_3304;
assign v_3306 = v_628 | v_630;
assign v_3309 = v_3302 | v_3307 | v_3308;
assign v_3317 = v_3315 | v_3316;
assign v_3319 = v_3314 | v_3318;
assign v_3321 = v_3313 | v_3320;
assign v_3323 = v_3312 | v_3322;
assign v_3325 = v_3311 | v_3324;
assign v_3327 = v_3310 | v_3326;
assign v_3332 = v_3330 | v_3331;
assign v_3338 = v_3334 | v_3335 | v_3336 | v_3337;
assign v_3340 = v_3333 | v_3339;
assign v_3344 = v_3328 | v_3329 | v_3341 | v_3342 | v_3343;
assign v_3350 = v_3347 | v_3349;
assign v_3352 = v_3346 | v_3351;
assign v_3354 = v_730 | v_732;
assign v_3358 = v_3356 | v_3357;
assign v_3361 = v_3359 | v_3360;
assign v_3368 = v_3365 | v_3367;
assign v_3370 = v_3364 | v_3369;
assign v_3372 = v_13531 | v_13532;
assign v_3378 = v_3375 | v_3376 | v_3377;
assign v_3380 = v_3374 | v_3379;
assign v_3386 = v_3383 | v_3384 | v_3385;
assign v_3388 = v_3382 | v_3387;
assign v_3393 = v_3390 | v_3391 | v_3392;
assign v_3397 = v_3395 | v_3396;
assign v_3398 = v_873 | v_871;
assign v_3403 = v_3399 | v_3400 | v_3401 | v_3402;
assign v_3407 = v_13533 | v_13534;
assign v_3413 = v_3410 | v_3411 | v_3412;
assign v_3415 = v_3409 | v_3414;
assign v_3421 = v_3418 | v_3419 | v_3420;
assign v_3423 = v_3417 | v_3422;
assign v_3428 = v_3425 | v_3426 | v_3427;
assign v_3432 = v_3430 | v_3431;
assign v_3433 = v_954 | v_952;
assign v_3438 = v_3434 | v_3435 | v_3436 | v_3437;
assign v_3442 = v_13535 | v_13536;
assign v_3448 = v_3445 | v_3446 | v_3447;
assign v_3450 = v_3444 | v_3449;
assign v_3456 = v_3453 | v_3454 | v_3455;
assign v_3458 = v_3452 | v_3457;
assign v_3463 = v_3460 | v_3461 | v_3462;
assign v_3467 = v_3465 | v_3466;
assign v_3468 = v_1035 | v_1033;
assign v_3473 = v_3469 | v_3470 | v_3471 | v_3472;
assign v_3477 = v_13537 | v_13538;
assign v_3483 = v_3480 | v_3481 | v_3482;
assign v_3485 = v_3479 | v_3484;
assign v_3491 = v_3488 | v_3489 | v_3490;
assign v_3493 = v_3487 | v_3492;
assign v_3498 = v_3495 | v_3496 | v_3497;
assign v_3502 = v_3500 | v_3501;
assign v_3503 = v_1116 | v_1114;
assign v_3508 = v_3504 | v_3505 | v_3506 | v_3507;
assign v_3512 = v_13539 | v_13540;
assign v_3518 = v_3515 | v_3516 | v_3517;
assign v_3520 = v_3514 | v_3519;
assign v_3526 = v_3523 | v_3524 | v_3525;
assign v_3528 = v_3522 | v_3527;
assign v_3533 = v_3530 | v_3531 | v_3532;
assign v_3537 = v_3535 | v_3536;
assign v_3538 = v_1197 | v_1195;
assign v_3543 = v_3539 | v_3540 | v_3541 | v_3542;
assign v_3547 = v_13541 | v_13542;
assign v_3553 = v_3550 | v_3551 | v_3552;
assign v_3555 = v_3549 | v_3554;
assign v_3561 = v_3558 | v_3559 | v_3560;
assign v_3563 = v_3557 | v_3562;
assign v_3568 = v_3565 | v_3566 | v_3567;
assign v_3572 = v_3570 | v_3571;
assign v_3573 = v_1278 | v_1276;
assign v_3578 = v_3574 | v_3575 | v_3576 | v_3577;
assign v_3582 = v_13543 | v_13544;
assign v_3588 = v_3585 | v_3586 | v_3587;
assign v_3590 = v_3584 | v_3589;
assign v_3596 = v_3593 | v_3594 | v_3595;
assign v_3598 = v_3592 | v_3597;
assign v_3603 = v_3600 | v_3601 | v_3602;
assign v_3607 = v_3605 | v_3606;
assign v_3608 = v_1359 | v_1357;
assign v_3613 = v_3609 | v_3610 | v_3611 | v_3612;
assign v_3617 = v_13545 | v_13546;
assign v_3623 = v_3620 | v_3621 | v_3622;
assign v_3625 = v_3619 | v_3624;
assign v_3631 = v_3628 | v_3629 | v_3630;
assign v_3633 = v_3627 | v_3632;
assign v_3638 = v_3635 | v_3636 | v_3637;
assign v_3642 = v_3640 | v_3641;
assign v_3643 = v_1440 | v_1438;
assign v_3648 = v_3644 | v_3645 | v_3646 | v_3647;
assign v_3652 = v_13547 | v_13548;
assign v_3658 = v_3655 | v_3656 | v_3657;
assign v_3660 = v_3654 | v_3659;
assign v_3666 = v_3663 | v_3664 | v_3665;
assign v_3668 = v_3662 | v_3667;
assign v_3673 = v_3670 | v_3671 | v_3672;
assign v_3677 = v_3675 | v_3676;
assign v_3678 = v_1521 | v_1519;
assign v_3683 = v_3679 | v_3680 | v_3681 | v_3682;
assign v_3687 = v_13549 | v_13550;
assign v_3695 = v_3693 | v_3694;
assign v_3696 = v_13551 | v_13552;
assign v_3700 = v_3697 | v_3698 | v_3699;
assign v_3702 = v_3690 | v_3691 | v_3692 | v_3701;
assign v_3705 = v_3689 | v_3703 | v_3704;
assign v_3707 = v_294 | v_296;
assign v_3710 = v_3706 | v_3708 | v_3709;
assign v_3711 = v_308 | v_310;
assign v_3717 = v_3714 | v_3715 | v_3716;
assign v_3719 = v_3713 | v_3718;
assign v_3721 = v_3712 | v_3720;
assign v_3722 = ~v_333 | v_335 | v_337;
assign v_3725 = v_3723 | v_3724;
assign v_3734 = v_3732 | v_3733;
assign v_3736 = v_3730 | v_3731 | v_3735;
assign v_3741 = v_380 | v_382;
assign v_3744 = v_3742 | v_3743;
assign v_3747 = v_3745 | v_3746;
assign v_3749 = v_3738 | v_3739 | v_3740 | v_3748;
assign v_3755 = v_3751 | v_3752 | v_3753 | v_3754;
assign v_3757 = v_3737 | v_3750 | v_3756;
assign v_3759 = v_3726 | v_3727 | v_3728 | v_3729 | v_3758;
assign v_3768 = v_3766 | v_3767;
assign v_3770 = v_3764 | v_3765 | v_3769;
assign v_3775 = v_445 | v_447;
assign v_3778 = v_3776 | v_3777;
assign v_3781 = v_3779 | v_3780;
assign v_3783 = v_3772 | v_3773 | v_3774 | v_3782;
assign v_3789 = v_3785 | v_3786 | v_3787 | v_3788;
assign v_3791 = v_3771 | v_3784 | v_3790;
assign v_3793 = v_3760 | v_3761 | v_3762 | v_3763 | v_3792;
assign v_3800 = v_3798 | v_3799;
assign v_3801 = v_13553 | v_13554;
assign v_3805 = v_3802 | v_3803 | v_3804;
assign v_3807 = v_3795 | v_3796 | v_3797 | v_3806;
assign v_3810 = v_3794 | v_3808 | v_3809;
assign v_3815 = v_3812 | v_3814;
assign v_3817 = v_3811 | v_3816;
assign v_3821 = v_3819 | v_3820;
assign v_3822 = v_570 | v_572;
assign v_3825 = v_3818 | v_3823 | v_3824;
assign v_3830 = v_3826 | v_3827 | v_3828 | v_3829;
assign v_3835 = v_3832 | v_3834;
assign v_3837 = v_3831 | v_3836;
assign v_3841 = v_3839 | v_3840;
assign v_3842 = v_628 | v_630;
assign v_3845 = v_3838 | v_3843 | v_3844;
assign v_3853 = v_3851 | v_3852;
assign v_3855 = v_3850 | v_3854;
assign v_3857 = v_3849 | v_3856;
assign v_3859 = v_3848 | v_3858;
assign v_3861 = v_3847 | v_3860;
assign v_3863 = v_3846 | v_3862;
assign v_3868 = v_3866 | v_3867;
assign v_3874 = v_3870 | v_3871 | v_3872 | v_3873;
assign v_3876 = v_3869 | v_3875;
assign v_3880 = v_3864 | v_3865 | v_3877 | v_3878 | v_3879;
assign v_3886 = v_3883 | v_3885;
assign v_3888 = v_3882 | v_3887;
assign v_3890 = v_730 | v_732;
assign v_3894 = v_3892 | v_3893;
assign v_3897 = v_3895 | v_3896;
assign v_3904 = v_3901 | v_3903;
assign v_3906 = v_3900 | v_3905;
assign v_3908 = v_13555 | v_13556;
assign v_3914 = v_3911 | v_3912 | v_3913;
assign v_3916 = v_3910 | v_3915;
assign v_3922 = v_3919 | v_3920 | v_3921;
assign v_3924 = v_3918 | v_3923;
assign v_3929 = v_3926 | v_3927 | v_3928;
assign v_3933 = v_3931 | v_3932;
assign v_3934 = v_873 | v_871;
assign v_3939 = v_3935 | v_3936 | v_3937 | v_3938;
assign v_3943 = v_13557 | v_13558;
assign v_3949 = v_3946 | v_3947 | v_3948;
assign v_3951 = v_3945 | v_3950;
assign v_3957 = v_3954 | v_3955 | v_3956;
assign v_3959 = v_3953 | v_3958;
assign v_3964 = v_3961 | v_3962 | v_3963;
assign v_3968 = v_3966 | v_3967;
assign v_3969 = v_954 | v_952;
assign v_3974 = v_3970 | v_3971 | v_3972 | v_3973;
assign v_3978 = v_13559 | v_13560;
assign v_3984 = v_3981 | v_3982 | v_3983;
assign v_3986 = v_3980 | v_3985;
assign v_3992 = v_3989 | v_3990 | v_3991;
assign v_3994 = v_3988 | v_3993;
assign v_3999 = v_3996 | v_3997 | v_3998;
assign v_4003 = v_4001 | v_4002;
assign v_4004 = v_1035 | v_1033;
assign v_4009 = v_4005 | v_4006 | v_4007 | v_4008;
assign v_4013 = v_13561 | v_13562;
assign v_4019 = v_4016 | v_4017 | v_4018;
assign v_4021 = v_4015 | v_4020;
assign v_4027 = v_4024 | v_4025 | v_4026;
assign v_4029 = v_4023 | v_4028;
assign v_4034 = v_4031 | v_4032 | v_4033;
assign v_4038 = v_4036 | v_4037;
assign v_4039 = v_1116 | v_1114;
assign v_4044 = v_4040 | v_4041 | v_4042 | v_4043;
assign v_4048 = v_13563 | v_13564;
assign v_4054 = v_4051 | v_4052 | v_4053;
assign v_4056 = v_4050 | v_4055;
assign v_4062 = v_4059 | v_4060 | v_4061;
assign v_4064 = v_4058 | v_4063;
assign v_4069 = v_4066 | v_4067 | v_4068;
assign v_4073 = v_4071 | v_4072;
assign v_4074 = v_1197 | v_1195;
assign v_4079 = v_4075 | v_4076 | v_4077 | v_4078;
assign v_4083 = v_13565 | v_13566;
assign v_4089 = v_4086 | v_4087 | v_4088;
assign v_4091 = v_4085 | v_4090;
assign v_4097 = v_4094 | v_4095 | v_4096;
assign v_4099 = v_4093 | v_4098;
assign v_4104 = v_4101 | v_4102 | v_4103;
assign v_4108 = v_4106 | v_4107;
assign v_4109 = v_1278 | v_1276;
assign v_4114 = v_4110 | v_4111 | v_4112 | v_4113;
assign v_4118 = v_13567 | v_13568;
assign v_4124 = v_4121 | v_4122 | v_4123;
assign v_4126 = v_4120 | v_4125;
assign v_4132 = v_4129 | v_4130 | v_4131;
assign v_4134 = v_4128 | v_4133;
assign v_4139 = v_4136 | v_4137 | v_4138;
assign v_4143 = v_4141 | v_4142;
assign v_4144 = v_1359 | v_1357;
assign v_4149 = v_4145 | v_4146 | v_4147 | v_4148;
assign v_4153 = v_13569 | v_13570;
assign v_4159 = v_4156 | v_4157 | v_4158;
assign v_4161 = v_4155 | v_4160;
assign v_4167 = v_4164 | v_4165 | v_4166;
assign v_4169 = v_4163 | v_4168;
assign v_4174 = v_4171 | v_4172 | v_4173;
assign v_4178 = v_4176 | v_4177;
assign v_4179 = v_1440 | v_1438;
assign v_4184 = v_4180 | v_4181 | v_4182 | v_4183;
assign v_4188 = v_13571 | v_13572;
assign v_4194 = v_4191 | v_4192 | v_4193;
assign v_4196 = v_4190 | v_4195;
assign v_4202 = v_4199 | v_4200 | v_4201;
assign v_4204 = v_4198 | v_4203;
assign v_4209 = v_4206 | v_4207 | v_4208;
assign v_4213 = v_4211 | v_4212;
assign v_4214 = v_1521 | v_1519;
assign v_4219 = v_4215 | v_4216 | v_4217 | v_4218;
assign v_4223 = v_13573 | v_13574;
assign v_4231 = v_4229 | v_4230;
assign v_4232 = v_13575 | v_13576;
assign v_4236 = v_4233 | v_4234 | v_4235;
assign v_4238 = v_4226 | v_4227 | v_4228 | v_4237;
assign v_4241 = v_4225 | v_4239 | v_4240;
assign v_4243 = v_294 | v_296;
assign v_4246 = v_4242 | v_4244 | v_4245;
assign v_4247 = v_308 | v_310;
assign v_4253 = v_4250 | v_4251 | v_4252;
assign v_4255 = v_4249 | v_4254;
assign v_4257 = v_4248 | v_4256;
assign v_4258 = ~v_333 | v_335 | v_337;
assign v_4261 = v_4259 | v_4260;
assign v_4270 = v_4268 | v_4269;
assign v_4272 = v_4266 | v_4267 | v_4271;
assign v_4277 = v_380 | v_382;
assign v_4280 = v_4278 | v_4279;
assign v_4283 = v_4281 | v_4282;
assign v_4285 = v_4274 | v_4275 | v_4276 | v_4284;
assign v_4291 = v_4287 | v_4288 | v_4289 | v_4290;
assign v_4293 = v_4273 | v_4286 | v_4292;
assign v_4295 = v_4262 | v_4263 | v_4264 | v_4265 | v_4294;
assign v_4304 = v_4302 | v_4303;
assign v_4306 = v_4300 | v_4301 | v_4305;
assign v_4311 = v_445 | v_447;
assign v_4314 = v_4312 | v_4313;
assign v_4317 = v_4315 | v_4316;
assign v_4319 = v_4308 | v_4309 | v_4310 | v_4318;
assign v_4325 = v_4321 | v_4322 | v_4323 | v_4324;
assign v_4327 = v_4307 | v_4320 | v_4326;
assign v_4329 = v_4296 | v_4297 | v_4298 | v_4299 | v_4328;
assign v_4336 = v_4334 | v_4335;
assign v_4337 = v_13577 | v_13578;
assign v_4341 = v_4338 | v_4339 | v_4340;
assign v_4343 = v_4331 | v_4332 | v_4333 | v_4342;
assign v_4346 = v_4330 | v_4344 | v_4345;
assign v_4351 = v_4348 | v_4350;
assign v_4353 = v_4347 | v_4352;
assign v_4357 = v_4355 | v_4356;
assign v_4358 = v_570 | v_572;
assign v_4361 = v_4354 | v_4359 | v_4360;
assign v_4366 = v_4362 | v_4363 | v_4364 | v_4365;
assign v_4371 = v_4368 | v_4370;
assign v_4373 = v_4367 | v_4372;
assign v_4377 = v_4375 | v_4376;
assign v_4378 = v_628 | v_630;
assign v_4381 = v_4374 | v_4379 | v_4380;
assign v_4389 = v_4387 | v_4388;
assign v_4391 = v_4386 | v_4390;
assign v_4393 = v_4385 | v_4392;
assign v_4395 = v_4384 | v_4394;
assign v_4397 = v_4383 | v_4396;
assign v_4399 = v_4382 | v_4398;
assign v_4404 = v_4402 | v_4403;
assign v_4410 = v_4406 | v_4407 | v_4408 | v_4409;
assign v_4412 = v_4405 | v_4411;
assign v_4416 = v_4400 | v_4401 | v_4413 | v_4414 | v_4415;
assign v_4422 = v_4419 | v_4421;
assign v_4424 = v_4418 | v_4423;
assign v_4426 = v_730 | v_732;
assign v_4430 = v_4428 | v_4429;
assign v_4433 = v_4431 | v_4432;
assign v_4440 = v_4437 | v_4439;
assign v_4442 = v_4436 | v_4441;
assign v_4444 = v_13579 | v_13580;
assign v_4450 = v_4447 | v_4448 | v_4449;
assign v_4452 = v_4446 | v_4451;
assign v_4458 = v_4455 | v_4456 | v_4457;
assign v_4460 = v_4454 | v_4459;
assign v_4465 = v_4462 | v_4463 | v_4464;
assign v_4469 = v_4467 | v_4468;
assign v_4470 = v_873 | v_871;
assign v_4475 = v_4471 | v_4472 | v_4473 | v_4474;
assign v_4479 = v_13581 | v_13582;
assign v_4485 = v_4482 | v_4483 | v_4484;
assign v_4487 = v_4481 | v_4486;
assign v_4493 = v_4490 | v_4491 | v_4492;
assign v_4495 = v_4489 | v_4494;
assign v_4500 = v_4497 | v_4498 | v_4499;
assign v_4504 = v_4502 | v_4503;
assign v_4505 = v_954 | v_952;
assign v_4510 = v_4506 | v_4507 | v_4508 | v_4509;
assign v_4514 = v_13583 | v_13584;
assign v_4520 = v_4517 | v_4518 | v_4519;
assign v_4522 = v_4516 | v_4521;
assign v_4528 = v_4525 | v_4526 | v_4527;
assign v_4530 = v_4524 | v_4529;
assign v_4535 = v_4532 | v_4533 | v_4534;
assign v_4539 = v_4537 | v_4538;
assign v_4540 = v_1035 | v_1033;
assign v_4545 = v_4541 | v_4542 | v_4543 | v_4544;
assign v_4549 = v_13585 | v_13586;
assign v_4555 = v_4552 | v_4553 | v_4554;
assign v_4557 = v_4551 | v_4556;
assign v_4563 = v_4560 | v_4561 | v_4562;
assign v_4565 = v_4559 | v_4564;
assign v_4570 = v_4567 | v_4568 | v_4569;
assign v_4574 = v_4572 | v_4573;
assign v_4575 = v_1116 | v_1114;
assign v_4580 = v_4576 | v_4577 | v_4578 | v_4579;
assign v_4584 = v_13587 | v_13588;
assign v_4590 = v_4587 | v_4588 | v_4589;
assign v_4592 = v_4586 | v_4591;
assign v_4598 = v_4595 | v_4596 | v_4597;
assign v_4600 = v_4594 | v_4599;
assign v_4605 = v_4602 | v_4603 | v_4604;
assign v_4609 = v_4607 | v_4608;
assign v_4610 = v_1197 | v_1195;
assign v_4615 = v_4611 | v_4612 | v_4613 | v_4614;
assign v_4619 = v_13589 | v_13590;
assign v_4625 = v_4622 | v_4623 | v_4624;
assign v_4627 = v_4621 | v_4626;
assign v_4633 = v_4630 | v_4631 | v_4632;
assign v_4635 = v_4629 | v_4634;
assign v_4640 = v_4637 | v_4638 | v_4639;
assign v_4644 = v_4642 | v_4643;
assign v_4645 = v_1278 | v_1276;
assign v_4650 = v_4646 | v_4647 | v_4648 | v_4649;
assign v_4654 = v_13591 | v_13592;
assign v_4660 = v_4657 | v_4658 | v_4659;
assign v_4662 = v_4656 | v_4661;
assign v_4668 = v_4665 | v_4666 | v_4667;
assign v_4670 = v_4664 | v_4669;
assign v_4675 = v_4672 | v_4673 | v_4674;
assign v_4679 = v_4677 | v_4678;
assign v_4680 = v_1359 | v_1357;
assign v_4685 = v_4681 | v_4682 | v_4683 | v_4684;
assign v_4689 = v_13593 | v_13594;
assign v_4695 = v_4692 | v_4693 | v_4694;
assign v_4697 = v_4691 | v_4696;
assign v_4703 = v_4700 | v_4701 | v_4702;
assign v_4705 = v_4699 | v_4704;
assign v_4710 = v_4707 | v_4708 | v_4709;
assign v_4714 = v_4712 | v_4713;
assign v_4715 = v_1440 | v_1438;
assign v_4720 = v_4716 | v_4717 | v_4718 | v_4719;
assign v_4724 = v_13595 | v_13596;
assign v_4730 = v_4727 | v_4728 | v_4729;
assign v_4732 = v_4726 | v_4731;
assign v_4738 = v_4735 | v_4736 | v_4737;
assign v_4740 = v_4734 | v_4739;
assign v_4745 = v_4742 | v_4743 | v_4744;
assign v_4749 = v_4747 | v_4748;
assign v_4750 = v_1521 | v_1519;
assign v_4755 = v_4751 | v_4752 | v_4753 | v_4754;
assign v_4759 = v_13597 | v_13598;
assign v_4766 = v_4764 | v_4765;
assign v_4767 = v_13599 | v_13600;
assign v_4771 = v_4768 | v_4769 | v_4770;
assign v_4773 = v_4761 | v_4762 | v_4763 | v_4772;
assign v_4776 = v_4760 | v_4774 | v_4775;
assign v_4778 = v_294 | v_296;
assign v_4781 = v_4777 | v_4779 | v_4780;
assign v_4782 = v_308 | v_310;
assign v_4788 = v_4785 | v_4786 | v_4787;
assign v_4790 = v_4784 | v_4789;
assign v_4792 = v_4783 | v_4791;
assign v_4793 = ~v_333 | v_335 | v_337;
assign v_4796 = v_4794 | v_4795;
assign v_4805 = v_4803 | v_4804;
assign v_4807 = v_4801 | v_4802 | v_4806;
assign v_4812 = v_380 | v_382;
assign v_4815 = v_4813 | v_4814;
assign v_4818 = v_4816 | v_4817;
assign v_4820 = v_4809 | v_4810 | v_4811 | v_4819;
assign v_4826 = v_4822 | v_4823 | v_4824 | v_4825;
assign v_4828 = v_4808 | v_4821 | v_4827;
assign v_4830 = v_4797 | v_4798 | v_4799 | v_4800 | v_4829;
assign v_4839 = v_4837 | v_4838;
assign v_4841 = v_4835 | v_4836 | v_4840;
assign v_4846 = v_445 | v_447;
assign v_4849 = v_4847 | v_4848;
assign v_4852 = v_4850 | v_4851;
assign v_4854 = v_4843 | v_4844 | v_4845 | v_4853;
assign v_4860 = v_4856 | v_4857 | v_4858 | v_4859;
assign v_4862 = v_4842 | v_4855 | v_4861;
assign v_4864 = v_4831 | v_4832 | v_4833 | v_4834 | v_4863;
assign v_4871 = v_4869 | v_4870;
assign v_4872 = v_13601 | v_13602;
assign v_4876 = v_4873 | v_4874 | v_4875;
assign v_4878 = v_4866 | v_4867 | v_4868 | v_4877;
assign v_4881 = v_4865 | v_4879 | v_4880;
assign v_4886 = v_4883 | v_4885;
assign v_4888 = v_4882 | v_4887;
assign v_4892 = v_4890 | v_4891;
assign v_4893 = v_570 | v_572;
assign v_4896 = v_4889 | v_4894 | v_4895;
assign v_4901 = v_4897 | v_4898 | v_4899 | v_4900;
assign v_4906 = v_4903 | v_4905;
assign v_4908 = v_4902 | v_4907;
assign v_4912 = v_4910 | v_4911;
assign v_4913 = v_628 | v_630;
assign v_4916 = v_4909 | v_4914 | v_4915;
assign v_4924 = v_4922 | v_4923;
assign v_4926 = v_4921 | v_4925;
assign v_4928 = v_4920 | v_4927;
assign v_4930 = v_4919 | v_4929;
assign v_4932 = v_4918 | v_4931;
assign v_4934 = v_4917 | v_4933;
assign v_4939 = v_4937 | v_4938;
assign v_4945 = v_4941 | v_4942 | v_4943 | v_4944;
assign v_4947 = v_4940 | v_4946;
assign v_4951 = v_4935 | v_4936 | v_4948 | v_4949 | v_4950;
assign v_4957 = v_4954 | v_4956;
assign v_4959 = v_4953 | v_4958;
assign v_4961 = v_730 | v_732;
assign v_4965 = v_4963 | v_4964;
assign v_4968 = v_4966 | v_4967;
assign v_4975 = v_4972 | v_4974;
assign v_4977 = v_4971 | v_4976;
assign v_4979 = v_13603 | v_13604;
assign v_4985 = v_4982 | v_4983 | v_4984;
assign v_4987 = v_4981 | v_4986;
assign v_4993 = v_4990 | v_4991 | v_4992;
assign v_4995 = v_4989 | v_4994;
assign v_5000 = v_4997 | v_4998 | v_4999;
assign v_5004 = v_5002 | v_5003;
assign v_5005 = v_873 | v_871;
assign v_5010 = v_5006 | v_5007 | v_5008 | v_5009;
assign v_5014 = v_13605 | v_13606;
assign v_5020 = v_5017 | v_5018 | v_5019;
assign v_5022 = v_5016 | v_5021;
assign v_5028 = v_5025 | v_5026 | v_5027;
assign v_5030 = v_5024 | v_5029;
assign v_5035 = v_5032 | v_5033 | v_5034;
assign v_5039 = v_5037 | v_5038;
assign v_5040 = v_954 | v_952;
assign v_5045 = v_5041 | v_5042 | v_5043 | v_5044;
assign v_5049 = v_13607 | v_13608;
assign v_5055 = v_5052 | v_5053 | v_5054;
assign v_5057 = v_5051 | v_5056;
assign v_5063 = v_5060 | v_5061 | v_5062;
assign v_5065 = v_5059 | v_5064;
assign v_5070 = v_5067 | v_5068 | v_5069;
assign v_5074 = v_5072 | v_5073;
assign v_5075 = v_1035 | v_1033;
assign v_5080 = v_5076 | v_5077 | v_5078 | v_5079;
assign v_5084 = v_13609 | v_13610;
assign v_5090 = v_5087 | v_5088 | v_5089;
assign v_5092 = v_5086 | v_5091;
assign v_5098 = v_5095 | v_5096 | v_5097;
assign v_5100 = v_5094 | v_5099;
assign v_5105 = v_5102 | v_5103 | v_5104;
assign v_5109 = v_5107 | v_5108;
assign v_5110 = v_1116 | v_1114;
assign v_5115 = v_5111 | v_5112 | v_5113 | v_5114;
assign v_5119 = v_13611 | v_13612;
assign v_5125 = v_5122 | v_5123 | v_5124;
assign v_5127 = v_5121 | v_5126;
assign v_5133 = v_5130 | v_5131 | v_5132;
assign v_5135 = v_5129 | v_5134;
assign v_5140 = v_5137 | v_5138 | v_5139;
assign v_5144 = v_5142 | v_5143;
assign v_5145 = v_1197 | v_1195;
assign v_5150 = v_5146 | v_5147 | v_5148 | v_5149;
assign v_5154 = v_13613 | v_13614;
assign v_5160 = v_5157 | v_5158 | v_5159;
assign v_5162 = v_5156 | v_5161;
assign v_5168 = v_5165 | v_5166 | v_5167;
assign v_5170 = v_5164 | v_5169;
assign v_5175 = v_5172 | v_5173 | v_5174;
assign v_5179 = v_5177 | v_5178;
assign v_5180 = v_1278 | v_1276;
assign v_5185 = v_5181 | v_5182 | v_5183 | v_5184;
assign v_5189 = v_13615 | v_13616;
assign v_5195 = v_5192 | v_5193 | v_5194;
assign v_5197 = v_5191 | v_5196;
assign v_5203 = v_5200 | v_5201 | v_5202;
assign v_5205 = v_5199 | v_5204;
assign v_5210 = v_5207 | v_5208 | v_5209;
assign v_5214 = v_5212 | v_5213;
assign v_5215 = v_1359 | v_1357;
assign v_5220 = v_5216 | v_5217 | v_5218 | v_5219;
assign v_5224 = v_13617 | v_13618;
assign v_5230 = v_5227 | v_5228 | v_5229;
assign v_5232 = v_5226 | v_5231;
assign v_5238 = v_5235 | v_5236 | v_5237;
assign v_5240 = v_5234 | v_5239;
assign v_5245 = v_5242 | v_5243 | v_5244;
assign v_5249 = v_5247 | v_5248;
assign v_5250 = v_1440 | v_1438;
assign v_5255 = v_5251 | v_5252 | v_5253 | v_5254;
assign v_5259 = v_13619 | v_13620;
assign v_5265 = v_5262 | v_5263 | v_5264;
assign v_5267 = v_5261 | v_5266;
assign v_5273 = v_5270 | v_5271 | v_5272;
assign v_5275 = v_5269 | v_5274;
assign v_5280 = v_5277 | v_5278 | v_5279;
assign v_5284 = v_5282 | v_5283;
assign v_5285 = v_1521 | v_1519;
assign v_5290 = v_5286 | v_5287 | v_5288 | v_5289;
assign v_5294 = v_13621 | v_13622;
assign v_5302 = v_5300 | v_5301;
assign v_5303 = v_13623 | v_13624;
assign v_5307 = v_5304 | v_5305 | v_5306;
assign v_5309 = v_5297 | v_5298 | v_5299 | v_5308;
assign v_5312 = v_5296 | v_5310 | v_5311;
assign v_5314 = v_294 | v_296;
assign v_5317 = v_5313 | v_5315 | v_5316;
assign v_5318 = v_308 | v_310;
assign v_5324 = v_5321 | v_5322 | v_5323;
assign v_5326 = v_5320 | v_5325;
assign v_5328 = v_5319 | v_5327;
assign v_5329 = ~v_333 | v_335 | v_337;
assign v_5332 = v_5330 | v_5331;
assign v_5341 = v_5339 | v_5340;
assign v_5343 = v_5337 | v_5338 | v_5342;
assign v_5348 = v_380 | v_382;
assign v_5351 = v_5349 | v_5350;
assign v_5354 = v_5352 | v_5353;
assign v_5356 = v_5345 | v_5346 | v_5347 | v_5355;
assign v_5362 = v_5358 | v_5359 | v_5360 | v_5361;
assign v_5364 = v_5344 | v_5357 | v_5363;
assign v_5366 = v_5333 | v_5334 | v_5335 | v_5336 | v_5365;
assign v_5375 = v_5373 | v_5374;
assign v_5377 = v_5371 | v_5372 | v_5376;
assign v_5382 = v_445 | v_447;
assign v_5385 = v_5383 | v_5384;
assign v_5388 = v_5386 | v_5387;
assign v_5390 = v_5379 | v_5380 | v_5381 | v_5389;
assign v_5396 = v_5392 | v_5393 | v_5394 | v_5395;
assign v_5398 = v_5378 | v_5391 | v_5397;
assign v_5400 = v_5367 | v_5368 | v_5369 | v_5370 | v_5399;
assign v_5407 = v_5405 | v_5406;
assign v_5408 = v_13625 | v_13626;
assign v_5412 = v_5409 | v_5410 | v_5411;
assign v_5414 = v_5402 | v_5403 | v_5404 | v_5413;
assign v_5417 = v_5401 | v_5415 | v_5416;
assign v_5422 = v_5419 | v_5421;
assign v_5424 = v_5418 | v_5423;
assign v_5428 = v_5426 | v_5427;
assign v_5429 = v_570 | v_572;
assign v_5432 = v_5425 | v_5430 | v_5431;
assign v_5437 = v_5433 | v_5434 | v_5435 | v_5436;
assign v_5442 = v_5439 | v_5441;
assign v_5444 = v_5438 | v_5443;
assign v_5448 = v_5446 | v_5447;
assign v_5449 = v_628 | v_630;
assign v_5452 = v_5445 | v_5450 | v_5451;
assign v_5460 = v_5458 | v_5459;
assign v_5462 = v_5457 | v_5461;
assign v_5464 = v_5456 | v_5463;
assign v_5466 = v_5455 | v_5465;
assign v_5468 = v_5454 | v_5467;
assign v_5470 = v_5453 | v_5469;
assign v_5475 = v_5473 | v_5474;
assign v_5481 = v_5477 | v_5478 | v_5479 | v_5480;
assign v_5483 = v_5476 | v_5482;
assign v_5487 = v_5471 | v_5472 | v_5484 | v_5485 | v_5486;
assign v_5493 = v_5490 | v_5492;
assign v_5495 = v_5489 | v_5494;
assign v_5497 = v_730 | v_732;
assign v_5501 = v_5499 | v_5500;
assign v_5504 = v_5502 | v_5503;
assign v_5511 = v_5508 | v_5510;
assign v_5513 = v_5507 | v_5512;
assign v_5515 = v_13627 | v_13628;
assign v_5521 = v_5518 | v_5519 | v_5520;
assign v_5523 = v_5517 | v_5522;
assign v_5529 = v_5526 | v_5527 | v_5528;
assign v_5531 = v_5525 | v_5530;
assign v_5536 = v_5533 | v_5534 | v_5535;
assign v_5540 = v_5538 | v_5539;
assign v_5541 = v_873 | v_871;
assign v_5546 = v_5542 | v_5543 | v_5544 | v_5545;
assign v_5550 = v_13629 | v_13630;
assign v_5556 = v_5553 | v_5554 | v_5555;
assign v_5558 = v_5552 | v_5557;
assign v_5564 = v_5561 | v_5562 | v_5563;
assign v_5566 = v_5560 | v_5565;
assign v_5571 = v_5568 | v_5569 | v_5570;
assign v_5575 = v_5573 | v_5574;
assign v_5576 = v_954 | v_952;
assign v_5581 = v_5577 | v_5578 | v_5579 | v_5580;
assign v_5585 = v_13631 | v_13632;
assign v_5591 = v_5588 | v_5589 | v_5590;
assign v_5593 = v_5587 | v_5592;
assign v_5599 = v_5596 | v_5597 | v_5598;
assign v_5601 = v_5595 | v_5600;
assign v_5606 = v_5603 | v_5604 | v_5605;
assign v_5610 = v_5608 | v_5609;
assign v_5611 = v_1035 | v_1033;
assign v_5616 = v_5612 | v_5613 | v_5614 | v_5615;
assign v_5620 = v_13633 | v_13634;
assign v_5626 = v_5623 | v_5624 | v_5625;
assign v_5628 = v_5622 | v_5627;
assign v_5634 = v_5631 | v_5632 | v_5633;
assign v_5636 = v_5630 | v_5635;
assign v_5641 = v_5638 | v_5639 | v_5640;
assign v_5645 = v_5643 | v_5644;
assign v_5646 = v_1116 | v_1114;
assign v_5651 = v_5647 | v_5648 | v_5649 | v_5650;
assign v_5655 = v_13635 | v_13636;
assign v_5661 = v_5658 | v_5659 | v_5660;
assign v_5663 = v_5657 | v_5662;
assign v_5669 = v_5666 | v_5667 | v_5668;
assign v_5671 = v_5665 | v_5670;
assign v_5676 = v_5673 | v_5674 | v_5675;
assign v_5680 = v_5678 | v_5679;
assign v_5681 = v_1197 | v_1195;
assign v_5686 = v_5682 | v_5683 | v_5684 | v_5685;
assign v_5690 = v_13637 | v_13638;
assign v_5696 = v_5693 | v_5694 | v_5695;
assign v_5698 = v_5692 | v_5697;
assign v_5704 = v_5701 | v_5702 | v_5703;
assign v_5706 = v_5700 | v_5705;
assign v_5711 = v_5708 | v_5709 | v_5710;
assign v_5715 = v_5713 | v_5714;
assign v_5716 = v_1278 | v_1276;
assign v_5721 = v_5717 | v_5718 | v_5719 | v_5720;
assign v_5725 = v_13639 | v_13640;
assign v_5731 = v_5728 | v_5729 | v_5730;
assign v_5733 = v_5727 | v_5732;
assign v_5739 = v_5736 | v_5737 | v_5738;
assign v_5741 = v_5735 | v_5740;
assign v_5746 = v_5743 | v_5744 | v_5745;
assign v_5750 = v_5748 | v_5749;
assign v_5751 = v_1359 | v_1357;
assign v_5756 = v_5752 | v_5753 | v_5754 | v_5755;
assign v_5760 = v_13641 | v_13642;
assign v_5766 = v_5763 | v_5764 | v_5765;
assign v_5768 = v_5762 | v_5767;
assign v_5774 = v_5771 | v_5772 | v_5773;
assign v_5776 = v_5770 | v_5775;
assign v_5781 = v_5778 | v_5779 | v_5780;
assign v_5785 = v_5783 | v_5784;
assign v_5786 = v_1440 | v_1438;
assign v_5791 = v_5787 | v_5788 | v_5789 | v_5790;
assign v_5795 = v_13643 | v_13644;
assign v_5801 = v_5798 | v_5799 | v_5800;
assign v_5803 = v_5797 | v_5802;
assign v_5809 = v_5806 | v_5807 | v_5808;
assign v_5811 = v_5805 | v_5810;
assign v_5816 = v_5813 | v_5814 | v_5815;
assign v_5820 = v_5818 | v_5819;
assign v_5821 = v_1521 | v_1519;
assign v_5826 = v_5822 | v_5823 | v_5824 | v_5825;
assign v_5830 = v_13645 | v_13646;
assign v_5833 = v_5832 | ~v_1572;
assign v_5839 = v_5835 | v_5837 | v_5838;
assign v_5841 = v_294 | v_296;
assign v_5844 = v_5840 | v_5842 | v_5843;
assign v_5845 = v_308 | v_310;
assign v_5851 = v_5848 | v_5849 | v_5850;
assign v_5853 = v_5847 | v_5852;
assign v_5855 = v_5846 | v_5854;
assign v_5856 = ~v_333 | v_335 | v_337;
assign v_5859 = v_5857 | v_5858;
assign v_5861 = v_5834 | v_5860;
assign v_5870 = v_5868 | v_5869;
assign v_5872 = v_5866 | v_5867 | v_5871;
assign v_5877 = v_380 | v_382;
assign v_5880 = v_5878 | v_5879;
assign v_5883 = v_5881 | v_5882;
assign v_5885 = v_5874 | v_5875 | v_5876 | v_5884;
assign v_5891 = v_5887 | v_5888 | v_5889 | v_5890;
assign v_5893 = v_5873 | v_5886 | v_5892;
assign v_5895 = v_5862 | v_5863 | v_5864 | v_5865 | v_5894;
assign v_5904 = v_5902 | v_5903;
assign v_5906 = v_5900 | v_5901 | v_5905;
assign v_5911 = v_445 | v_447;
assign v_5914 = v_5912 | v_5913;
assign v_5917 = v_5915 | v_5916;
assign v_5919 = v_5908 | v_5909 | v_5910 | v_5918;
assign v_5925 = v_5921 | v_5922 | v_5923 | v_5924;
assign v_5927 = v_5907 | v_5920 | v_5926;
assign v_5929 = v_5896 | v_5897 | v_5898 | v_5899 | v_5928;
assign v_5934 = v_5930 | v_5932 | v_5933;
assign v_5937 = v_5935 | v_5936;
assign v_5941 = v_5939 | v_5940;
assign v_5942 = v_570 | v_572;
assign v_5945 = v_5938 | v_5943 | v_5944;
assign v_5950 = v_5946 | v_5947 | v_5948 | v_5949;
assign v_5953 = v_5951 | v_5952;
assign v_5957 = v_5955 | v_5956;
assign v_5958 = v_628 | v_630;
assign v_5961 = v_5954 | v_5959 | v_5960;
assign v_5969 = v_5967 | v_5968;
assign v_5971 = v_5966 | v_5970;
assign v_5973 = v_5965 | v_5972;
assign v_5975 = v_5964 | v_5974;
assign v_5977 = v_5963 | v_5976;
assign v_5979 = v_5962 | v_5978;
assign v_5984 = v_5982 | v_5983;
assign v_5990 = v_5986 | v_5987 | v_5988 | v_5989;
assign v_5992 = v_5985 | v_5991;
assign v_5996 = v_5980 | v_5981 | v_5993 | v_5994 | v_5995;
assign v_6000 = v_5998 | v_5999;
assign v_6002 = v_730 | v_732;
assign v_6006 = v_6004 | v_6005;
assign v_6009 = v_6007 | v_6008;
assign v_6014 = v_6012 | v_6013;
assign v_6016 = v_13647 | v_13648;
assign v_6022 = v_6019 | v_6020 | v_6021;
assign v_6024 = v_6018 | v_6023;
assign v_6030 = v_6027 | v_6028 | v_6029;
assign v_6032 = v_6026 | v_6031;
assign v_6037 = v_6034 | v_6035 | v_6036;
assign v_6041 = v_6039 | v_6040;
assign v_6042 = v_873 | v_871;
assign v_6047 = v_6043 | v_6044 | v_6045 | v_6046;
assign v_6051 = v_13649 | v_13650;
assign v_6057 = v_6054 | v_6055 | v_6056;
assign v_6059 = v_6053 | v_6058;
assign v_6065 = v_6062 | v_6063 | v_6064;
assign v_6067 = v_6061 | v_6066;
assign v_6072 = v_6069 | v_6070 | v_6071;
assign v_6076 = v_6074 | v_6075;
assign v_6077 = v_954 | v_952;
assign v_6082 = v_6078 | v_6079 | v_6080 | v_6081;
assign v_6086 = v_13651 | v_13652;
assign v_6092 = v_6089 | v_6090 | v_6091;
assign v_6094 = v_6088 | v_6093;
assign v_6100 = v_6097 | v_6098 | v_6099;
assign v_6102 = v_6096 | v_6101;
assign v_6107 = v_6104 | v_6105 | v_6106;
assign v_6111 = v_6109 | v_6110;
assign v_6112 = v_1035 | v_1033;
assign v_6117 = v_6113 | v_6114 | v_6115 | v_6116;
assign v_6121 = v_13653 | v_13654;
assign v_6127 = v_6124 | v_6125 | v_6126;
assign v_6129 = v_6123 | v_6128;
assign v_6135 = v_6132 | v_6133 | v_6134;
assign v_6137 = v_6131 | v_6136;
assign v_6142 = v_6139 | v_6140 | v_6141;
assign v_6146 = v_6144 | v_6145;
assign v_6147 = v_1116 | v_1114;
assign v_6152 = v_6148 | v_6149 | v_6150 | v_6151;
assign v_6156 = v_13655 | v_13656;
assign v_6162 = v_6159 | v_6160 | v_6161;
assign v_6164 = v_6158 | v_6163;
assign v_6170 = v_6167 | v_6168 | v_6169;
assign v_6172 = v_6166 | v_6171;
assign v_6177 = v_6174 | v_6175 | v_6176;
assign v_6181 = v_6179 | v_6180;
assign v_6182 = v_1197 | v_1195;
assign v_6187 = v_6183 | v_6184 | v_6185 | v_6186;
assign v_6191 = v_13657 | v_13658;
assign v_6197 = v_6194 | v_6195 | v_6196;
assign v_6199 = v_6193 | v_6198;
assign v_6205 = v_6202 | v_6203 | v_6204;
assign v_6207 = v_6201 | v_6206;
assign v_6212 = v_6209 | v_6210 | v_6211;
assign v_6216 = v_6214 | v_6215;
assign v_6217 = v_1278 | v_1276;
assign v_6222 = v_6218 | v_6219 | v_6220 | v_6221;
assign v_6226 = v_13659 | v_13660;
assign v_6232 = v_6229 | v_6230 | v_6231;
assign v_6234 = v_6228 | v_6233;
assign v_6240 = v_6237 | v_6238 | v_6239;
assign v_6242 = v_6236 | v_6241;
assign v_6247 = v_6244 | v_6245 | v_6246;
assign v_6251 = v_6249 | v_6250;
assign v_6252 = v_1359 | v_1357;
assign v_6257 = v_6253 | v_6254 | v_6255 | v_6256;
assign v_6261 = v_13661 | v_13662;
assign v_6267 = v_6264 | v_6265 | v_6266;
assign v_6269 = v_6263 | v_6268;
assign v_6275 = v_6272 | v_6273 | v_6274;
assign v_6277 = v_6271 | v_6276;
assign v_6282 = v_6279 | v_6280 | v_6281;
assign v_6286 = v_6284 | v_6285;
assign v_6287 = v_1440 | v_1438;
assign v_6292 = v_6288 | v_6289 | v_6290 | v_6291;
assign v_6296 = v_13663 | v_13664;
assign v_6302 = v_6299 | v_6300 | v_6301;
assign v_6304 = v_6298 | v_6303;
assign v_6310 = v_6307 | v_6308 | v_6309;
assign v_6312 = v_6306 | v_6311;
assign v_6317 = v_6314 | v_6315 | v_6316;
assign v_6321 = v_6319 | v_6320;
assign v_6322 = v_1521 | v_1519;
assign v_6327 = v_6323 | v_6324 | v_6325 | v_6326;
assign v_6331 = v_13665 | v_13666;
assign v_6339 = v_6337 | v_6338;
assign v_6340 = v_13667 | v_13668;
assign v_6344 = v_6341 | v_6342 | v_6343;
assign v_6346 = v_6334 | v_6335 | v_6336 | v_6345;
assign v_6349 = v_6333 | v_6347 | v_6348;
assign v_6351 = v_294 | v_296;
assign v_6354 = v_6350 | v_6352 | v_6353;
assign v_6355 = v_308 | v_310;
assign v_6361 = v_6358 | v_6359 | v_6360;
assign v_6363 = v_6357 | v_6362;
assign v_6365 = v_6356 | v_6364;
assign v_6366 = ~v_333 | v_335 | v_337;
assign v_6369 = v_6367 | v_6368;
assign v_6378 = v_6376 | v_6377;
assign v_6380 = v_6374 | v_6375 | v_6379;
assign v_6385 = v_380 | v_382;
assign v_6388 = v_6386 | v_6387;
assign v_6391 = v_6389 | v_6390;
assign v_6393 = v_6382 | v_6383 | v_6384 | v_6392;
assign v_6399 = v_6395 | v_6396 | v_6397 | v_6398;
assign v_6401 = v_6381 | v_6394 | v_6400;
assign v_6403 = v_6370 | v_6371 | v_6372 | v_6373 | v_6402;
assign v_6412 = v_6410 | v_6411;
assign v_6414 = v_6408 | v_6409 | v_6413;
assign v_6419 = v_445 | v_447;
assign v_6422 = v_6420 | v_6421;
assign v_6425 = v_6423 | v_6424;
assign v_6427 = v_6416 | v_6417 | v_6418 | v_6426;
assign v_6433 = v_6429 | v_6430 | v_6431 | v_6432;
assign v_6435 = v_6415 | v_6428 | v_6434;
assign v_6437 = v_6404 | v_6405 | v_6406 | v_6407 | v_6436;
assign v_6444 = v_6442 | v_6443;
assign v_6445 = v_13669 | v_13670;
assign v_6449 = v_6446 | v_6447 | v_6448;
assign v_6451 = v_6439 | v_6440 | v_6441 | v_6450;
assign v_6454 = v_6438 | v_6452 | v_6453;
assign v_6459 = v_6456 | v_6458;
assign v_6461 = v_6455 | v_6460;
assign v_6465 = v_6463 | v_6464;
assign v_6466 = v_570 | v_572;
assign v_6469 = v_6462 | v_6467 | v_6468;
assign v_6474 = v_6470 | v_6471 | v_6472 | v_6473;
assign v_6479 = v_6476 | v_6478;
assign v_6481 = v_6475 | v_6480;
assign v_6485 = v_6483 | v_6484;
assign v_6486 = v_628 | v_630;
assign v_6489 = v_6482 | v_6487 | v_6488;
assign v_6497 = v_6495 | v_6496;
assign v_6499 = v_6494 | v_6498;
assign v_6501 = v_6493 | v_6500;
assign v_6503 = v_6492 | v_6502;
assign v_6505 = v_6491 | v_6504;
assign v_6507 = v_6490 | v_6506;
assign v_6512 = v_6510 | v_6511;
assign v_6518 = v_6514 | v_6515 | v_6516 | v_6517;
assign v_6520 = v_6513 | v_6519;
assign v_6524 = v_6508 | v_6509 | v_6521 | v_6522 | v_6523;
assign v_6530 = v_6527 | v_6529;
assign v_6532 = v_6526 | v_6531;
assign v_6534 = v_730 | v_732;
assign v_6538 = v_6536 | v_6537;
assign v_6541 = v_6539 | v_6540;
assign v_6548 = v_6545 | v_6547;
assign v_6550 = v_6544 | v_6549;
assign v_6552 = v_13671 | v_13672;
assign v_6558 = v_6555 | v_6556 | v_6557;
assign v_6560 = v_6554 | v_6559;
assign v_6566 = v_6563 | v_6564 | v_6565;
assign v_6568 = v_6562 | v_6567;
assign v_6573 = v_6570 | v_6571 | v_6572;
assign v_6577 = v_6575 | v_6576;
assign v_6578 = v_873 | v_871;
assign v_6583 = v_6579 | v_6580 | v_6581 | v_6582;
assign v_6587 = v_13673 | v_13674;
assign v_6593 = v_6590 | v_6591 | v_6592;
assign v_6595 = v_6589 | v_6594;
assign v_6601 = v_6598 | v_6599 | v_6600;
assign v_6603 = v_6597 | v_6602;
assign v_6608 = v_6605 | v_6606 | v_6607;
assign v_6612 = v_6610 | v_6611;
assign v_6613 = v_954 | v_952;
assign v_6618 = v_6614 | v_6615 | v_6616 | v_6617;
assign v_6622 = v_13675 | v_13676;
assign v_6628 = v_6625 | v_6626 | v_6627;
assign v_6630 = v_6624 | v_6629;
assign v_6636 = v_6633 | v_6634 | v_6635;
assign v_6638 = v_6632 | v_6637;
assign v_6643 = v_6640 | v_6641 | v_6642;
assign v_6647 = v_6645 | v_6646;
assign v_6648 = v_1035 | v_1033;
assign v_6653 = v_6649 | v_6650 | v_6651 | v_6652;
assign v_6657 = v_13677 | v_13678;
assign v_6663 = v_6660 | v_6661 | v_6662;
assign v_6665 = v_6659 | v_6664;
assign v_6671 = v_6668 | v_6669 | v_6670;
assign v_6673 = v_6667 | v_6672;
assign v_6678 = v_6675 | v_6676 | v_6677;
assign v_6682 = v_6680 | v_6681;
assign v_6683 = v_1116 | v_1114;
assign v_6688 = v_6684 | v_6685 | v_6686 | v_6687;
assign v_6692 = v_13679 | v_13680;
assign v_6698 = v_6695 | v_6696 | v_6697;
assign v_6700 = v_6694 | v_6699;
assign v_6706 = v_6703 | v_6704 | v_6705;
assign v_6708 = v_6702 | v_6707;
assign v_6713 = v_6710 | v_6711 | v_6712;
assign v_6717 = v_6715 | v_6716;
assign v_6718 = v_1197 | v_1195;
assign v_6723 = v_6719 | v_6720 | v_6721 | v_6722;
assign v_6727 = v_13681 | v_13682;
assign v_6733 = v_6730 | v_6731 | v_6732;
assign v_6735 = v_6729 | v_6734;
assign v_6741 = v_6738 | v_6739 | v_6740;
assign v_6743 = v_6737 | v_6742;
assign v_6748 = v_6745 | v_6746 | v_6747;
assign v_6752 = v_6750 | v_6751;
assign v_6753 = v_1278 | v_1276;
assign v_6758 = v_6754 | v_6755 | v_6756 | v_6757;
assign v_6762 = v_13683 | v_13684;
assign v_6768 = v_6765 | v_6766 | v_6767;
assign v_6770 = v_6764 | v_6769;
assign v_6776 = v_6773 | v_6774 | v_6775;
assign v_6778 = v_6772 | v_6777;
assign v_6783 = v_6780 | v_6781 | v_6782;
assign v_6787 = v_6785 | v_6786;
assign v_6788 = v_1359 | v_1357;
assign v_6793 = v_6789 | v_6790 | v_6791 | v_6792;
assign v_6797 = v_13685 | v_13686;
assign v_6803 = v_6800 | v_6801 | v_6802;
assign v_6805 = v_6799 | v_6804;
assign v_6811 = v_6808 | v_6809 | v_6810;
assign v_6813 = v_6807 | v_6812;
assign v_6818 = v_6815 | v_6816 | v_6817;
assign v_6822 = v_6820 | v_6821;
assign v_6823 = v_1440 | v_1438;
assign v_6828 = v_6824 | v_6825 | v_6826 | v_6827;
assign v_6832 = v_13687 | v_13688;
assign v_6838 = v_6835 | v_6836 | v_6837;
assign v_6840 = v_6834 | v_6839;
assign v_6846 = v_6843 | v_6844 | v_6845;
assign v_6848 = v_6842 | v_6847;
assign v_6853 = v_6850 | v_6851 | v_6852;
assign v_6857 = v_6855 | v_6856;
assign v_6858 = v_1521 | v_1519;
assign v_6863 = v_6859 | v_6860 | v_6861 | v_6862;
assign v_6867 = v_13689 | v_13690;
assign v_7083 = ~v_7079 | v_7081 | v_7082;
assign v_7090 = v_7088 | v_7089;
assign v_7124 = ~v_7120 | v_7122 | v_7123;
assign v_7126 = v_13691 | v_13692 | v_13693;
assign v_7133 = v_7127 | v_7129 | v_7131 | v_7132;
assign v_7137 = v_7094 | v_7135 | v_7136;
assign v_7143 = v_7141 | v_7142;
assign v_7151 = v_7148 | v_7150;
assign v_7157 = ~v_7146 | v_7153 | v_7155 | v_7156;
assign v_7166 = v_7163 | v_7165;
assign v_7168 = ~v_7145 | v_7160 | v_7162 | v_7167;
assign v_7172 = v_7170 | v_7171;
assign v_7181 = ~v_7177 | v_7179 | v_7180;
assign v_7187 = v_7183 | v_7185 | v_7186;
assign v_7195 = v_7189 | v_7191 | v_7193 | v_7194;
assign v_7197 = v_7174 | v_7176 | v_7196;
assign v_7209 = ~v_7199 | v_7201 | v_7203 | v_7207 | v_7208;
assign v_7222 = v_7219 | v_7221;
assign v_7235 = v_7227 | v_7229 | v_7231 | v_7233 | v_7234;
assign v_7250 = v_7246 | v_7248 | v_7249;
assign v_7254 = v_7240 | v_7242 | v_7244 | v_7252 | v_7253;
assign v_7269 = v_13694 | v_13695;
assign v_7271 = v_7237 | v_7256 | v_7270;
assign v_7275 = v_13696 | v_13697;
assign v_7287 = v_7284 | v_7286;
assign v_7300 = v_7292 | v_7294 | v_7296 | v_7298 | v_7299;
assign v_7315 = v_7311 | v_7313 | v_7314;
assign v_7319 = v_7305 | v_7307 | v_7309 | v_7317 | v_7318;
assign v_7334 = v_13698 | v_13699;
assign v_7336 = v_7302 | v_7321 | v_7335;
assign v_7340 = v_13700 | v_13701;
assign v_7346 = v_7342 | v_7344 | v_7345;
assign v_7350 = v_7348 | v_7349;
assign v_7388 = ~v_7384 | v_7386 | v_7387;
assign v_7390 = v_13702 | v_13703 | v_13704;
assign v_7397 = v_7391 | v_7393 | v_7395 | v_7396;
assign v_7401 = v_7358 | v_7399 | v_7400;
assign v_7407 = v_7405 | v_7406;
assign v_7412 = ~v_7408 | v_7410 | v_7411;
assign v_7420 = v_7418 | v_7419;
assign v_7424 = v_7414 | v_7423;
assign v_7434 = v_7428 | v_7432 | v_7433;
assign v_7443 = ~v_7439 | v_7441 | v_7442;
assign v_7447 = v_7426 | v_7436 | v_7438 | v_7445 | v_7446;
assign v_7454 = v_7451 | v_7453;
assign v_7459 = v_7456 | v_7458;
assign v_7464 = v_7461 | v_7449 | v_7462 | v_7463;
assign v_7470 = ~v_7466 | v_7468 | v_7469;
assign v_7478 = v_7476 | v_7477;
assign v_7482 = v_7472 | v_7481;
assign v_7492 = v_7486 | v_7490 | v_7491;
assign v_7501 = ~v_7497 | v_7499 | v_7500;
assign v_7505 = v_7484 | v_7494 | v_7496 | v_7503 | v_7504;
assign v_7518 = v_7516 | v_7517;
assign v_7520 = v_7514 | v_7519;
assign v_7522 = v_7512 | v_7521;
assign v_7524 = v_7510 | v_7523;
assign v_7526 = v_7508 | v_7525;
assign v_7528 = v_7506 | v_7527;
assign v_7545 = v_7543 | v_7544;
assign v_7555 = v_7552 | v_7554;
assign v_7560 = v_7557 | v_7559;
assign v_7565 = v_7562 | v_7550 | v_7563 | v_7564;
assign v_7569 = v_13705 | v_13706;
assign v_7576 = ~v_7572 | v_7574 | v_7575;
assign v_7584 = v_7582 | v_7583;
assign v_7588 = v_7578 | v_7587;
assign v_7603 = v_7600 | v_7602;
assign v_7611 = v_7606 | v_7607 | v_7609 | v_7610;
assign v_7616 = ~v_7612 | v_7614 | v_7615;
assign v_7624 = v_7618 | v_7623;
assign v_7629 = ~v_7625 | v_7627 | v_7628;
assign v_7637 = v_7631 | v_7636;
assign v_7645 = ~v_7641 | v_7643 | v_7644;
assign v_7653 = v_7651 | v_7652;
assign v_7657 = v_7647 | v_7656;
assign v_7662 = v_13707 | v_13708;
assign v_7670 = v_7668 | v_7669;
assign v_7674 = v_7672 | v_7673;
assign v_7680 = ~v_7666 | v_7676 | v_7678 | v_7679;
assign v_7687 = v_7685 | v_7686;
assign v_7693 = v_7691 | v_7692;
assign v_7697 = v_7695 | v_7696;
assign v_7703 = ~v_7689 | v_7699 | v_7701 | v_7702;
assign v_7710 = v_7708 | v_7709;
assign v_7716 = v_7714 | v_7715;
assign v_7720 = v_7718 | v_7719;
assign v_7726 = ~v_7712 | v_7722 | v_7724 | v_7725;
assign v_7733 = v_7731 | v_7732;
assign v_7743 = v_13709 | v_13710 | v_13711;
assign v_7751 = v_7749 | v_7750;
assign v_7755 = v_7753 | v_7754;
assign v_7761 = ~v_7747 | v_7757 | v_7759 | v_7760;
assign v_7768 = v_7766 | v_7767;
assign v_7774 = v_7772 | v_7773;
assign v_7778 = v_7776 | v_7777;
assign v_7784 = ~v_7770 | v_7780 | v_7782 | v_7783;
assign v_7791 = v_7789 | v_7790;
assign v_7797 = v_7795 | v_7796;
assign v_7801 = v_7799 | v_7800;
assign v_7807 = ~v_7793 | v_7803 | v_7805 | v_7806;
assign v_7814 = v_7812 | v_7813;
assign v_7824 = v_13712 | v_13713 | v_13714;
assign v_7832 = v_7830 | v_7831;
assign v_7836 = v_7834 | v_7835;
assign v_7842 = ~v_7828 | v_7838 | v_7840 | v_7841;
assign v_7849 = v_7847 | v_7848;
assign v_7855 = v_7853 | v_7854;
assign v_7859 = v_7857 | v_7858;
assign v_7865 = ~v_7851 | v_7861 | v_7863 | v_7864;
assign v_7872 = v_7870 | v_7871;
assign v_7878 = v_7876 | v_7877;
assign v_7882 = v_7880 | v_7881;
assign v_7888 = ~v_7874 | v_7884 | v_7886 | v_7887;
assign v_7895 = v_7893 | v_7894;
assign v_7905 = v_13715 | v_13716 | v_13717;
assign v_7913 = v_7911 | v_7912;
assign v_7917 = v_7915 | v_7916;
assign v_7923 = ~v_7909 | v_7919 | v_7921 | v_7922;
assign v_7930 = v_7928 | v_7929;
assign v_7936 = v_7934 | v_7935;
assign v_7940 = v_7938 | v_7939;
assign v_7946 = ~v_7932 | v_7942 | v_7944 | v_7945;
assign v_7953 = v_7951 | v_7952;
assign v_7959 = v_7957 | v_7958;
assign v_7963 = v_7961 | v_7962;
assign v_7969 = ~v_7955 | v_7965 | v_7967 | v_7968;
assign v_7976 = v_7974 | v_7975;
assign v_7986 = v_13718 | v_13719 | v_13720;
assign v_7994 = v_7992 | v_7993;
assign v_7998 = v_7996 | v_7997;
assign v_8004 = ~v_7990 | v_8000 | v_8002 | v_8003;
assign v_8011 = v_8009 | v_8010;
assign v_8017 = v_8015 | v_8016;
assign v_8021 = v_8019 | v_8020;
assign v_8027 = ~v_8013 | v_8023 | v_8025 | v_8026;
assign v_8034 = v_8032 | v_8033;
assign v_8040 = v_8038 | v_8039;
assign v_8044 = v_8042 | v_8043;
assign v_8050 = ~v_8036 | v_8046 | v_8048 | v_8049;
assign v_8057 = v_8055 | v_8056;
assign v_8067 = v_13721 | v_13722 | v_13723;
assign v_8075 = v_8073 | v_8074;
assign v_8079 = v_8077 | v_8078;
assign v_8085 = ~v_8071 | v_8081 | v_8083 | v_8084;
assign v_8092 = v_8090 | v_8091;
assign v_8098 = v_8096 | v_8097;
assign v_8102 = v_8100 | v_8101;
assign v_8108 = ~v_8094 | v_8104 | v_8106 | v_8107;
assign v_8115 = v_8113 | v_8114;
assign v_8121 = v_8119 | v_8120;
assign v_8125 = v_8123 | v_8124;
assign v_8131 = ~v_8117 | v_8127 | v_8129 | v_8130;
assign v_8138 = v_8136 | v_8137;
assign v_8148 = v_13724 | v_13725 | v_13726;
assign v_8156 = v_8154 | v_8155;
assign v_8160 = v_8158 | v_8159;
assign v_8166 = ~v_8152 | v_8162 | v_8164 | v_8165;
assign v_8173 = v_8171 | v_8172;
assign v_8179 = v_8177 | v_8178;
assign v_8183 = v_8181 | v_8182;
assign v_8189 = ~v_8175 | v_8185 | v_8187 | v_8188;
assign v_8196 = v_8194 | v_8195;
assign v_8202 = v_8200 | v_8201;
assign v_8206 = v_8204 | v_8205;
assign v_8212 = ~v_8198 | v_8208 | v_8210 | v_8211;
assign v_8219 = v_8217 | v_8218;
assign v_8229 = v_13727 | v_13728 | v_13729;
assign v_8235 = v_8234 | ~v_8233;
assign v_8242 = v_13730 | v_13731;
assign v_8244 = v_7118 | v_7119;
assign v_8247 = v_8243 | v_8245 | v_8246;
assign v_8249 = v_8238 | v_8239 | v_8240 | v_8248;
assign v_8251 = v_8250 | ~v_8249;
assign v_8254 = v_8252 | v_8253;
assign v_8256 = v_7160 | v_7162;
assign v_8259 = v_8255 | v_8257 | v_8258;
assign v_8260 = v_7174 | v_7176;
assign v_8266 = v_8263 | v_8264 | v_8265;
assign v_8267 = v_7191 | v_7193 | v_7194;
assign v_8269 = v_8262 | v_8268;
assign v_8271 = v_8261 | v_8270;
assign v_8272 = ~v_7199 | v_7201 | v_7203;
assign v_8274 = v_7207 | v_7208;
assign v_8276 = v_8273 | v_8275;
assign v_8278 = v_8236 | v_8277;
assign v_8286 = v_7233 | v_7234;
assign v_8288 = v_8285 | v_8287;
assign v_8289 = v_7231 | v_7233 | v_7234;
assign v_8291 = v_8283 | v_8284 | v_8290;
assign v_8296 = v_7246 | v_7248;
assign v_8299 = v_8297 | v_8298;
assign v_8302 = v_8300 | v_8301;
assign v_8303 = v_7252 | v_7253;
assign v_8305 = v_8293 | v_8294 | v_8295 | v_8304;
assign v_8310 = v_7265 | v_7267 | v_7268;
assign v_8312 = v_8307 | v_8308 | v_8309 | v_8311;
assign v_8314 = v_8292 | v_8306 | v_8313;
assign v_8315 = v_7273 | v_7274;
assign v_8317 = v_8279 | v_8280 | v_8281 | v_8282 | v_8316;
assign v_8325 = v_7298 | v_7299;
assign v_8327 = v_8324 | v_8326;
assign v_8328 = v_7296 | v_7298 | v_7299;
assign v_8330 = v_8322 | v_8323 | v_8329;
assign v_8335 = v_7311 | v_7313;
assign v_8338 = v_8336 | v_8337;
assign v_8341 = v_8339 | v_8340;
assign v_8342 = v_7317 | v_7318;
assign v_8344 = v_8332 | v_8333 | v_8334 | v_8343;
assign v_8349 = v_7330 | v_7332 | v_7333;
assign v_8351 = v_8346 | v_8347 | v_8348 | v_8350;
assign v_8353 = v_8331 | v_8345 | v_8352;
assign v_8354 = v_7338 | v_7339;
assign v_8356 = v_8318 | v_8319 | v_8320 | v_8321 | v_8355;
assign v_8361 = v_8360 | ~v_8356;
assign v_8367 = v_8365 | v_8366;
assign v_8368 = v_13732 | v_13733;
assign v_8370 = v_7382 | v_7383;
assign v_8373 = v_8369 | v_8371 | v_8372;
assign v_8375 = v_8362 | v_8363 | v_8364 | v_8374;
assign v_8377 = v_8376 | ~v_8375;
assign v_8380 = v_8357 | v_8378 | v_8379;
assign v_8383 = v_8381 | v_8382;
assign v_8386 = v_7432 | v_7433;
assign v_8388 = v_8385 | v_8387;
assign v_8389 = v_7436 | v_7438;
assign v_8391 = v_7445 | v_7446;
assign v_8393 = v_8384 | v_8390 | v_8392;
assign v_8398 = v_8394 | v_8395 | v_8396 | v_8397;
assign v_8401 = v_8399 | v_8400;
assign v_8404 = v_7490 | v_7491;
assign v_8406 = v_8403 | v_8405;
assign v_8407 = v_7494 | v_7496;
assign v_8409 = v_7503 | v_7504;
assign v_8411 = v_8402 | v_8408 | v_8410;
assign v_8419 = v_8417 | v_8418;
assign v_8421 = v_8416 | v_8420;
assign v_8423 = v_8415 | v_8422;
assign v_8425 = v_8414 | v_8424;
assign v_8427 = v_8413 | v_8426;
assign v_8429 = v_8412 | v_8428;
assign v_8434 = v_8432 | v_8433;
assign v_8440 = v_8436 | v_8437 | v_8438 | v_8439;
assign v_8441 = v_7567 | v_7568;
assign v_8443 = v_8435 | v_8442;
assign v_8444 = v_7549 | v_7567 | v_7568;
assign v_8447 = v_7537 | v_7539;
assign v_8449 = v_8430 | v_8431 | v_8445 | v_8446 | v_8448;
assign v_8453 = v_8451 | v_8452;
assign v_8455 = v_7596 | v_7598;
assign v_8459 = v_8457 | v_8458;
assign v_8462 = v_8460 | v_8461;
assign v_8467 = v_8465 | v_8466;
assign v_8468 = v_7659 | v_7660;
assign v_8470 = v_13734 | v_13735;
assign v_8475 = v_7678 | v_7679;
assign v_8477 = v_8473 | v_8474 | v_8476;
assign v_8479 = v_8472 | v_8478;
assign v_8484 = v_7701 | v_7702;
assign v_8486 = v_8482 | v_8483 | v_8485;
assign v_8488 = v_8481 | v_8487;
assign v_8492 = v_7724 | v_7725;
assign v_8494 = v_8490 | v_8491 | v_8493;
assign v_8498 = v_8496 | v_8497;
assign v_8499 = v_7739 | v_7737;
assign v_8504 = v_8500 | v_8501 | v_8502 | v_8503;
assign v_8505 = v_7737 | v_7739 | v_7740 | v_7741 | v_7742;
assign v_8509 = v_13736 | v_13737;
assign v_8514 = v_7759 | v_7760;
assign v_8516 = v_8512 | v_8513 | v_8515;
assign v_8518 = v_8511 | v_8517;
assign v_8523 = v_7782 | v_7783;
assign v_8525 = v_8521 | v_8522 | v_8524;
assign v_8527 = v_8520 | v_8526;
assign v_8531 = v_7805 | v_7806;
assign v_8533 = v_8529 | v_8530 | v_8532;
assign v_8537 = v_8535 | v_8536;
assign v_8538 = v_7820 | v_7818;
assign v_8543 = v_8539 | v_8540 | v_8541 | v_8542;
assign v_8544 = v_7818 | v_7820 | v_7821 | v_7822 | v_7823;
assign v_8548 = v_13738 | v_13739;
assign v_8553 = v_7840 | v_7841;
assign v_8555 = v_8551 | v_8552 | v_8554;
assign v_8557 = v_8550 | v_8556;
assign v_8562 = v_7863 | v_7864;
assign v_8564 = v_8560 | v_8561 | v_8563;
assign v_8566 = v_8559 | v_8565;
assign v_8570 = v_7886 | v_7887;
assign v_8572 = v_8568 | v_8569 | v_8571;
assign v_8576 = v_8574 | v_8575;
assign v_8577 = v_7901 | v_7899;
assign v_8582 = v_8578 | v_8579 | v_8580 | v_8581;
assign v_8583 = v_7899 | v_7901 | v_7902 | v_7903 | v_7904;
assign v_8587 = v_13740 | v_13741;
assign v_8592 = v_7921 | v_7922;
assign v_8594 = v_8590 | v_8591 | v_8593;
assign v_8596 = v_8589 | v_8595;
assign v_8601 = v_7944 | v_7945;
assign v_8603 = v_8599 | v_8600 | v_8602;
assign v_8605 = v_8598 | v_8604;
assign v_8609 = v_7967 | v_7968;
assign v_8611 = v_8607 | v_8608 | v_8610;
assign v_8615 = v_8613 | v_8614;
assign v_8616 = v_7982 | v_7980;
assign v_8621 = v_8617 | v_8618 | v_8619 | v_8620;
assign v_8622 = v_7980 | v_7982 | v_7983 | v_7984 | v_7985;
assign v_8626 = v_13742 | v_13743;
assign v_8631 = v_8002 | v_8003;
assign v_8633 = v_8629 | v_8630 | v_8632;
assign v_8635 = v_8628 | v_8634;
assign v_8640 = v_8025 | v_8026;
assign v_8642 = v_8638 | v_8639 | v_8641;
assign v_8644 = v_8637 | v_8643;
assign v_8648 = v_8048 | v_8049;
assign v_8650 = v_8646 | v_8647 | v_8649;
assign v_8654 = v_8652 | v_8653;
assign v_8655 = v_8063 | v_8061;
assign v_8660 = v_8656 | v_8657 | v_8658 | v_8659;
assign v_8661 = v_8061 | v_8063 | v_8064 | v_8065 | v_8066;
assign v_8665 = v_13744 | v_13745;
assign v_8670 = v_8083 | v_8084;
assign v_8672 = v_8668 | v_8669 | v_8671;
assign v_8674 = v_8667 | v_8673;
assign v_8679 = v_8106 | v_8107;
assign v_8681 = v_8677 | v_8678 | v_8680;
assign v_8683 = v_8676 | v_8682;
assign v_8687 = v_8129 | v_8130;
assign v_8689 = v_8685 | v_8686 | v_8688;
assign v_8693 = v_8691 | v_8692;
assign v_8694 = v_8144 | v_8142;
assign v_8699 = v_8695 | v_8696 | v_8697 | v_8698;
assign v_8700 = v_8142 | v_8144 | v_8145 | v_8146 | v_8147;
assign v_8704 = v_13746 | v_13747;
assign v_8709 = v_8164 | v_8165;
assign v_8711 = v_8707 | v_8708 | v_8710;
assign v_8713 = v_8706 | v_8712;
assign v_8718 = v_8187 | v_8188;
assign v_8720 = v_8716 | v_8717 | v_8719;
assign v_8722 = v_8715 | v_8721;
assign v_8726 = v_8210 | v_8211;
assign v_8728 = v_8724 | v_8725 | v_8727;
assign v_8732 = v_8730 | v_8731;
assign v_8733 = v_8225 | v_8223;
assign v_8738 = v_8734 | v_8735 | v_8736 | v_8737;
assign v_8739 = v_8223 | v_8225 | v_8226 | v_8227 | v_8228;
assign v_8743 = v_13748 | v_13749;
assign v_8745 = v_8744 | v_8233;
assign v_8749 = v_8748 | v_8249;
assign v_8752 = v_8747 | v_8750 | v_8751;
assign v_8754 = v_7160 | v_7162;
assign v_8757 = v_8753 | v_8755 | v_8756;
assign v_8758 = v_7174 | v_7176;
assign v_8764 = v_8761 | v_8762 | v_8763;
assign v_8766 = v_8760 | v_8765;
assign v_8768 = v_8759 | v_8767;
assign v_8769 = ~v_7199 | v_7201 | v_7203;
assign v_8772 = v_8770 | v_8771;
assign v_8774 = v_8746 | v_8773;
assign v_8783 = v_8781 | v_8782;
assign v_8785 = v_8779 | v_8780 | v_8784;
assign v_8790 = v_7246 | v_7248;
assign v_8793 = v_8791 | v_8792;
assign v_8796 = v_8794 | v_8795;
assign v_8798 = v_8787 | v_8788 | v_8789 | v_8797;
assign v_8804 = v_8800 | v_8801 | v_8802 | v_8803;
assign v_8806 = v_8786 | v_8799 | v_8805;
assign v_8808 = v_8775 | v_8776 | v_8777 | v_8778 | v_8807;
assign v_8817 = v_8815 | v_8816;
assign v_8819 = v_8813 | v_8814 | v_8818;
assign v_8824 = v_7311 | v_7313;
assign v_8827 = v_8825 | v_8826;
assign v_8830 = v_8828 | v_8829;
assign v_8832 = v_8821 | v_8822 | v_8823 | v_8831;
assign v_8838 = v_8834 | v_8835 | v_8836 | v_8837;
assign v_8840 = v_8820 | v_8833 | v_8839;
assign v_8842 = v_8809 | v_8810 | v_8811 | v_8812 | v_8841;
assign v_8845 = v_8844 | v_8375;
assign v_8848 = v_8843 | v_8846 | v_8847;
assign v_8851 = v_8849 | v_8850;
assign v_8855 = v_8853 | v_8854;
assign v_8856 = v_7436 | v_7438;
assign v_8859 = v_8852 | v_8857 | v_8858;
assign v_8864 = v_8860 | v_8861 | v_8862 | v_8863;
assign v_8867 = v_8865 | v_8866;
assign v_8871 = v_8869 | v_8870;
assign v_8872 = v_7494 | v_7496;
assign v_8875 = v_8868 | v_8873 | v_8874;
assign v_8883 = v_8881 | v_8882;
assign v_8885 = v_8880 | v_8884;
assign v_8887 = v_8879 | v_8886;
assign v_8889 = v_8878 | v_8888;
assign v_8891 = v_8877 | v_8890;
assign v_8893 = v_8876 | v_8892;
assign v_8898 = v_8896 | v_8897;
assign v_8904 = v_8900 | v_8901 | v_8902 | v_8903;
assign v_8906 = v_8899 | v_8905;
assign v_8910 = v_8894 | v_8895 | v_8907 | v_8908 | v_8909;
assign v_8914 = v_8912 | v_8913;
assign v_8916 = v_7596 | v_7598;
assign v_8920 = v_8918 | v_8919;
assign v_8923 = v_8921 | v_8922;
assign v_8928 = v_8926 | v_8927;
assign v_8930 = v_13750 | v_13751;
assign v_8936 = v_8933 | v_8934 | v_8935;
assign v_8938 = v_8932 | v_8937;
assign v_8944 = v_8941 | v_8942 | v_8943;
assign v_8946 = v_8940 | v_8945;
assign v_8951 = v_8948 | v_8949 | v_8950;
assign v_8955 = v_8953 | v_8954;
assign v_8956 = v_7739 | v_7737;
assign v_8961 = v_8957 | v_8958 | v_8959 | v_8960;
assign v_8965 = v_13752 | v_13753;
assign v_8971 = v_8968 | v_8969 | v_8970;
assign v_8973 = v_8967 | v_8972;
assign v_8979 = v_8976 | v_8977 | v_8978;
assign v_8981 = v_8975 | v_8980;
assign v_8986 = v_8983 | v_8984 | v_8985;
assign v_8990 = v_8988 | v_8989;
assign v_8991 = v_7820 | v_7818;
assign v_8996 = v_8992 | v_8993 | v_8994 | v_8995;
assign v_9000 = v_13754 | v_13755;
assign v_9006 = v_9003 | v_9004 | v_9005;
assign v_9008 = v_9002 | v_9007;
assign v_9014 = v_9011 | v_9012 | v_9013;
assign v_9016 = v_9010 | v_9015;
assign v_9021 = v_9018 | v_9019 | v_9020;
assign v_9025 = v_9023 | v_9024;
assign v_9026 = v_7901 | v_7899;
assign v_9031 = v_9027 | v_9028 | v_9029 | v_9030;
assign v_9035 = v_13756 | v_13757;
assign v_9041 = v_9038 | v_9039 | v_9040;
assign v_9043 = v_9037 | v_9042;
assign v_9049 = v_9046 | v_9047 | v_9048;
assign v_9051 = v_9045 | v_9050;
assign v_9056 = v_9053 | v_9054 | v_9055;
assign v_9060 = v_9058 | v_9059;
assign v_9061 = v_7982 | v_7980;
assign v_9066 = v_9062 | v_9063 | v_9064 | v_9065;
assign v_9070 = v_13758 | v_13759;
assign v_9076 = v_9073 | v_9074 | v_9075;
assign v_9078 = v_9072 | v_9077;
assign v_9084 = v_9081 | v_9082 | v_9083;
assign v_9086 = v_9080 | v_9085;
assign v_9091 = v_9088 | v_9089 | v_9090;
assign v_9095 = v_9093 | v_9094;
assign v_9096 = v_8063 | v_8061;
assign v_9101 = v_9097 | v_9098 | v_9099 | v_9100;
assign v_9105 = v_13760 | v_13761;
assign v_9111 = v_9108 | v_9109 | v_9110;
assign v_9113 = v_9107 | v_9112;
assign v_9119 = v_9116 | v_9117 | v_9118;
assign v_9121 = v_9115 | v_9120;
assign v_9126 = v_9123 | v_9124 | v_9125;
assign v_9130 = v_9128 | v_9129;
assign v_9131 = v_8144 | v_8142;
assign v_9136 = v_9132 | v_9133 | v_9134 | v_9135;
assign v_9140 = v_13762 | v_13763;
assign v_9146 = v_9143 | v_9144 | v_9145;
assign v_9148 = v_9142 | v_9147;
assign v_9154 = v_9151 | v_9152 | v_9153;
assign v_9156 = v_9150 | v_9155;
assign v_9161 = v_9158 | v_9159 | v_9160;
assign v_9165 = v_9163 | v_9164;
assign v_9166 = v_8225 | v_8223;
assign v_9171 = v_9167 | v_9168 | v_9169 | v_9170;
assign v_9175 = v_13764 | v_13765;
assign v_9182 = v_9180 | v_9181;
assign v_9183 = v_13766 | v_13767;
assign v_9187 = v_9184 | v_9185 | v_9186;
assign v_9189 = v_9177 | v_9178 | v_9179 | v_9188;
assign v_9192 = v_9176 | v_9190 | v_9191;
assign v_9194 = v_7160 | v_7162;
assign v_9197 = v_9193 | v_9195 | v_9196;
assign v_9198 = v_7174 | v_7176;
assign v_9204 = v_9201 | v_9202 | v_9203;
assign v_9206 = v_9200 | v_9205;
assign v_9208 = v_9199 | v_9207;
assign v_9209 = ~v_7199 | v_7201 | v_7203;
assign v_9212 = v_9210 | v_9211;
assign v_9221 = v_9219 | v_9220;
assign v_9223 = v_9217 | v_9218 | v_9222;
assign v_9228 = v_7246 | v_7248;
assign v_9231 = v_9229 | v_9230;
assign v_9234 = v_9232 | v_9233;
assign v_9236 = v_9225 | v_9226 | v_9227 | v_9235;
assign v_9242 = v_9238 | v_9239 | v_9240 | v_9241;
assign v_9244 = v_9224 | v_9237 | v_9243;
assign v_9246 = v_9213 | v_9214 | v_9215 | v_9216 | v_9245;
assign v_9255 = v_9253 | v_9254;
assign v_9257 = v_9251 | v_9252 | v_9256;
assign v_9262 = v_7311 | v_7313;
assign v_9265 = v_9263 | v_9264;
assign v_9268 = v_9266 | v_9267;
assign v_9270 = v_9259 | v_9260 | v_9261 | v_9269;
assign v_9276 = v_9272 | v_9273 | v_9274 | v_9275;
assign v_9278 = v_9258 | v_9271 | v_9277;
assign v_9280 = v_9247 | v_9248 | v_9249 | v_9250 | v_9279;
assign v_9287 = v_9285 | v_9286;
assign v_9288 = v_13768 | v_13769;
assign v_9292 = v_9289 | v_9290 | v_9291;
assign v_9294 = v_9282 | v_9283 | v_9284 | v_9293;
assign v_9297 = v_9281 | v_9295 | v_9296;
assign v_9302 = v_9299 | v_9301;
assign v_9304 = v_9298 | v_9303;
assign v_9308 = v_9306 | v_9307;
assign v_9309 = v_7436 | v_7438;
assign v_9312 = v_9305 | v_9310 | v_9311;
assign v_9317 = v_9313 | v_9314 | v_9315 | v_9316;
assign v_9322 = v_9319 | v_9321;
assign v_9324 = v_9318 | v_9323;
assign v_9328 = v_9326 | v_9327;
assign v_9329 = v_7494 | v_7496;
assign v_9332 = v_9325 | v_9330 | v_9331;
assign v_9340 = v_9338 | v_9339;
assign v_9342 = v_9337 | v_9341;
assign v_9344 = v_9336 | v_9343;
assign v_9346 = v_9335 | v_9345;
assign v_9348 = v_9334 | v_9347;
assign v_9350 = v_9333 | v_9349;
assign v_9355 = v_9353 | v_9354;
assign v_9361 = v_9357 | v_9358 | v_9359 | v_9360;
assign v_9363 = v_9356 | v_9362;
assign v_9367 = v_9351 | v_9352 | v_9364 | v_9365 | v_9366;
assign v_9373 = v_9370 | v_9372;
assign v_9375 = v_9369 | v_9374;
assign v_9377 = v_7596 | v_7598;
assign v_9381 = v_9379 | v_9380;
assign v_9384 = v_9382 | v_9383;
assign v_9391 = v_9388 | v_9390;
assign v_9393 = v_9387 | v_9392;
assign v_9395 = v_13770 | v_13771;
assign v_9401 = v_9398 | v_9399 | v_9400;
assign v_9403 = v_9397 | v_9402;
assign v_9409 = v_9406 | v_9407 | v_9408;
assign v_9411 = v_9405 | v_9410;
assign v_9416 = v_9413 | v_9414 | v_9415;
assign v_9420 = v_9418 | v_9419;
assign v_9421 = v_7739 | v_7737;
assign v_9426 = v_9422 | v_9423 | v_9424 | v_9425;
assign v_9430 = v_13772 | v_13773;
assign v_9436 = v_9433 | v_9434 | v_9435;
assign v_9438 = v_9432 | v_9437;
assign v_9444 = v_9441 | v_9442 | v_9443;
assign v_9446 = v_9440 | v_9445;
assign v_9451 = v_9448 | v_9449 | v_9450;
assign v_9455 = v_9453 | v_9454;
assign v_9456 = v_7820 | v_7818;
assign v_9461 = v_9457 | v_9458 | v_9459 | v_9460;
assign v_9465 = v_13774 | v_13775;
assign v_9471 = v_9468 | v_9469 | v_9470;
assign v_9473 = v_9467 | v_9472;
assign v_9479 = v_9476 | v_9477 | v_9478;
assign v_9481 = v_9475 | v_9480;
assign v_9486 = v_9483 | v_9484 | v_9485;
assign v_9490 = v_9488 | v_9489;
assign v_9491 = v_7901 | v_7899;
assign v_9496 = v_9492 | v_9493 | v_9494 | v_9495;
assign v_9500 = v_13776 | v_13777;
assign v_9506 = v_9503 | v_9504 | v_9505;
assign v_9508 = v_9502 | v_9507;
assign v_9514 = v_9511 | v_9512 | v_9513;
assign v_9516 = v_9510 | v_9515;
assign v_9521 = v_9518 | v_9519 | v_9520;
assign v_9525 = v_9523 | v_9524;
assign v_9526 = v_7982 | v_7980;
assign v_9531 = v_9527 | v_9528 | v_9529 | v_9530;
assign v_9535 = v_13778 | v_13779;
assign v_9541 = v_9538 | v_9539 | v_9540;
assign v_9543 = v_9537 | v_9542;
assign v_9549 = v_9546 | v_9547 | v_9548;
assign v_9551 = v_9545 | v_9550;
assign v_9556 = v_9553 | v_9554 | v_9555;
assign v_9560 = v_9558 | v_9559;
assign v_9561 = v_8063 | v_8061;
assign v_9566 = v_9562 | v_9563 | v_9564 | v_9565;
assign v_9570 = v_13780 | v_13781;
assign v_9576 = v_9573 | v_9574 | v_9575;
assign v_9578 = v_9572 | v_9577;
assign v_9584 = v_9581 | v_9582 | v_9583;
assign v_9586 = v_9580 | v_9585;
assign v_9591 = v_9588 | v_9589 | v_9590;
assign v_9595 = v_9593 | v_9594;
assign v_9596 = v_8144 | v_8142;
assign v_9601 = v_9597 | v_9598 | v_9599 | v_9600;
assign v_9605 = v_13782 | v_13783;
assign v_9611 = v_9608 | v_9609 | v_9610;
assign v_9613 = v_9607 | v_9612;
assign v_9619 = v_9616 | v_9617 | v_9618;
assign v_9621 = v_9615 | v_9620;
assign v_9626 = v_9623 | v_9624 | v_9625;
assign v_9630 = v_9628 | v_9629;
assign v_9631 = v_8225 | v_8223;
assign v_9636 = v_9632 | v_9633 | v_9634 | v_9635;
assign v_9640 = v_13784 | v_13785;
assign v_9646 = v_13786 | v_13787;
assign v_9650 = v_9647 | v_9648 | v_9649;
assign v_9652 = v_9642 | v_9643 | v_9644 | v_9651;
assign v_9655 = v_9641 | v_9653 | v_9654;
assign v_9657 = v_7160 | v_7162;
assign v_9660 = v_9656 | v_9658 | v_9659;
assign v_9661 = v_7174 | v_7176;
assign v_9667 = v_9664 | v_9665 | v_9666;
assign v_9669 = v_9663 | v_9668;
assign v_9671 = v_9662 | v_9670;
assign v_9672 = ~v_7199 | v_7201 | v_7203;
assign v_9675 = v_9673 | v_9674;
assign v_9684 = v_9682 | v_9683;
assign v_9686 = v_9680 | v_9681 | v_9685;
assign v_9691 = v_7246 | v_7248;
assign v_9694 = v_9692 | v_9693;
assign v_9697 = v_9695 | v_9696;
assign v_9699 = v_9688 | v_9689 | v_9690 | v_9698;
assign v_9705 = v_9701 | v_9702 | v_9703 | v_9704;
assign v_9707 = v_9687 | v_9700 | v_9706;
assign v_9709 = v_9676 | v_9677 | v_9678 | v_9679 | v_9708;
assign v_9718 = v_9716 | v_9717;
assign v_9720 = v_9714 | v_9715 | v_9719;
assign v_9725 = v_7311 | v_7313;
assign v_9728 = v_9726 | v_9727;
assign v_9731 = v_9729 | v_9730;
assign v_9733 = v_9722 | v_9723 | v_9724 | v_9732;
assign v_9739 = v_9735 | v_9736 | v_9737 | v_9738;
assign v_9741 = v_9721 | v_9734 | v_9740;
assign v_9743 = v_9710 | v_9711 | v_9712 | v_9713 | v_9742;
assign v_9750 = v_9748 | v_9749;
assign v_9751 = v_13788 | v_13789;
assign v_9755 = v_9752 | v_9753 | v_9754;
assign v_9757 = v_9745 | v_9746 | v_9747 | v_9756;
assign v_9760 = v_9744 | v_9758 | v_9759;
assign v_9765 = v_9762 | v_9764;
assign v_9767 = v_9761 | v_9766;
assign v_9771 = v_9769 | v_9770;
assign v_9772 = v_7436 | v_7438;
assign v_9775 = v_9768 | v_9773 | v_9774;
assign v_9780 = v_9776 | v_9777 | v_9778 | v_9779;
assign v_9785 = v_9782 | v_9784;
assign v_9787 = v_9781 | v_9786;
assign v_9791 = v_9789 | v_9790;
assign v_9792 = v_7494 | v_7496;
assign v_9795 = v_9788 | v_9793 | v_9794;
assign v_9803 = v_9801 | v_9802;
assign v_9805 = v_9800 | v_9804;
assign v_9807 = v_9799 | v_9806;
assign v_9809 = v_9798 | v_9808;
assign v_9811 = v_9797 | v_9810;
assign v_9813 = v_9796 | v_9812;
assign v_9818 = v_9816 | v_9817;
assign v_9824 = v_9820 | v_9821 | v_9822 | v_9823;
assign v_9826 = v_9819 | v_9825;
assign v_9830 = v_9814 | v_9815 | v_9827 | v_9828 | v_9829;
assign v_9836 = v_9833 | v_9835;
assign v_9838 = v_9832 | v_9837;
assign v_9840 = v_7596 | v_7598;
assign v_9844 = v_9842 | v_9843;
assign v_9847 = v_9845 | v_9846;
assign v_9854 = v_9851 | v_9853;
assign v_9856 = v_9850 | v_9855;
assign v_9858 = v_13790 | v_13791;
assign v_9864 = v_9861 | v_9862 | v_9863;
assign v_9866 = v_9860 | v_9865;
assign v_9872 = v_9869 | v_9870 | v_9871;
assign v_9874 = v_9868 | v_9873;
assign v_9879 = v_9876 | v_9877 | v_9878;
assign v_9883 = v_9881 | v_9882;
assign v_9884 = v_7739 | v_7737;
assign v_9889 = v_9885 | v_9886 | v_9887 | v_9888;
assign v_9893 = v_13792 | v_13793;
assign v_9899 = v_9896 | v_9897 | v_9898;
assign v_9901 = v_9895 | v_9900;
assign v_9907 = v_9904 | v_9905 | v_9906;
assign v_9909 = v_9903 | v_9908;
assign v_9914 = v_9911 | v_9912 | v_9913;
assign v_9918 = v_9916 | v_9917;
assign v_9919 = v_7820 | v_7818;
assign v_9924 = v_9920 | v_9921 | v_9922 | v_9923;
assign v_9928 = v_13794 | v_13795;
assign v_9934 = v_9931 | v_9932 | v_9933;
assign v_9936 = v_9930 | v_9935;
assign v_9942 = v_9939 | v_9940 | v_9941;
assign v_9944 = v_9938 | v_9943;
assign v_9949 = v_9946 | v_9947 | v_9948;
assign v_9953 = v_9951 | v_9952;
assign v_9954 = v_7901 | v_7899;
assign v_9959 = v_9955 | v_9956 | v_9957 | v_9958;
assign v_9963 = v_13796 | v_13797;
assign v_9969 = v_9966 | v_9967 | v_9968;
assign v_9971 = v_9965 | v_9970;
assign v_9977 = v_9974 | v_9975 | v_9976;
assign v_9979 = v_9973 | v_9978;
assign v_9984 = v_9981 | v_9982 | v_9983;
assign v_9988 = v_9986 | v_9987;
assign v_9989 = v_7982 | v_7980;
assign v_9994 = v_9990 | v_9991 | v_9992 | v_9993;
assign v_9998 = v_13798 | v_13799;
assign v_10004 = v_10001 | v_10002 | v_10003;
assign v_10006 = v_10000 | v_10005;
assign v_10012 = v_10009 | v_10010 | v_10011;
assign v_10014 = v_10008 | v_10013;
assign v_10019 = v_10016 | v_10017 | v_10018;
assign v_10023 = v_10021 | v_10022;
assign v_10024 = v_8063 | v_8061;
assign v_10029 = v_10025 | v_10026 | v_10027 | v_10028;
assign v_10033 = v_13800 | v_13801;
assign v_10039 = v_10036 | v_10037 | v_10038;
assign v_10041 = v_10035 | v_10040;
assign v_10047 = v_10044 | v_10045 | v_10046;
assign v_10049 = v_10043 | v_10048;
assign v_10054 = v_10051 | v_10052 | v_10053;
assign v_10058 = v_10056 | v_10057;
assign v_10059 = v_8144 | v_8142;
assign v_10064 = v_10060 | v_10061 | v_10062 | v_10063;
assign v_10068 = v_13802 | v_13803;
assign v_10074 = v_10071 | v_10072 | v_10073;
assign v_10076 = v_10070 | v_10075;
assign v_10082 = v_10079 | v_10080 | v_10081;
assign v_10084 = v_10078 | v_10083;
assign v_10089 = v_10086 | v_10087 | v_10088;
assign v_10093 = v_10091 | v_10092;
assign v_10094 = v_8225 | v_8223;
assign v_10099 = v_10095 | v_10096 | v_10097 | v_10098;
assign v_10103 = v_13804 | v_13805;
assign v_10111 = v_10109 | v_10110;
assign v_10112 = v_13806 | v_13807;
assign v_10116 = v_10113 | v_10114 | v_10115;
assign v_10118 = v_10106 | v_10107 | v_10108 | v_10117;
assign v_10121 = v_10105 | v_10119 | v_10120;
assign v_10123 = v_7160 | v_7162;
assign v_10126 = v_10122 | v_10124 | v_10125;
assign v_10127 = v_7174 | v_7176;
assign v_10133 = v_10130 | v_10131 | v_10132;
assign v_10135 = v_10129 | v_10134;
assign v_10137 = v_10128 | v_10136;
assign v_10138 = ~v_7199 | v_7201 | v_7203;
assign v_10141 = v_10139 | v_10140;
assign v_10150 = v_10148 | v_10149;
assign v_10152 = v_10146 | v_10147 | v_10151;
assign v_10157 = v_7246 | v_7248;
assign v_10160 = v_10158 | v_10159;
assign v_10163 = v_10161 | v_10162;
assign v_10165 = v_10154 | v_10155 | v_10156 | v_10164;
assign v_10171 = v_10167 | v_10168 | v_10169 | v_10170;
assign v_10173 = v_10153 | v_10166 | v_10172;
assign v_10175 = v_10142 | v_10143 | v_10144 | v_10145 | v_10174;
assign v_10184 = v_10182 | v_10183;
assign v_10186 = v_10180 | v_10181 | v_10185;
assign v_10191 = v_7311 | v_7313;
assign v_10194 = v_10192 | v_10193;
assign v_10197 = v_10195 | v_10196;
assign v_10199 = v_10188 | v_10189 | v_10190 | v_10198;
assign v_10205 = v_10201 | v_10202 | v_10203 | v_10204;
assign v_10207 = v_10187 | v_10200 | v_10206;
assign v_10209 = v_10176 | v_10177 | v_10178 | v_10179 | v_10208;
assign v_10216 = v_10214 | v_10215;
assign v_10217 = v_13808 | v_13809;
assign v_10221 = v_10218 | v_10219 | v_10220;
assign v_10223 = v_10211 | v_10212 | v_10213 | v_10222;
assign v_10226 = v_10210 | v_10224 | v_10225;
assign v_10231 = v_10228 | v_10230;
assign v_10233 = v_10227 | v_10232;
assign v_10237 = v_10235 | v_10236;
assign v_10238 = v_7436 | v_7438;
assign v_10241 = v_10234 | v_10239 | v_10240;
assign v_10246 = v_10242 | v_10243 | v_10244 | v_10245;
assign v_10251 = v_10248 | v_10250;
assign v_10253 = v_10247 | v_10252;
assign v_10257 = v_10255 | v_10256;
assign v_10258 = v_7494 | v_7496;
assign v_10261 = v_10254 | v_10259 | v_10260;
assign v_10269 = v_10267 | v_10268;
assign v_10271 = v_10266 | v_10270;
assign v_10273 = v_10265 | v_10272;
assign v_10275 = v_10264 | v_10274;
assign v_10277 = v_10263 | v_10276;
assign v_10279 = v_10262 | v_10278;
assign v_10284 = v_10282 | v_10283;
assign v_10290 = v_10286 | v_10287 | v_10288 | v_10289;
assign v_10292 = v_10285 | v_10291;
assign v_10296 = v_10280 | v_10281 | v_10293 | v_10294 | v_10295;
assign v_10302 = v_10299 | v_10301;
assign v_10304 = v_10298 | v_10303;
assign v_10306 = v_7596 | v_7598;
assign v_10310 = v_10308 | v_10309;
assign v_10313 = v_10311 | v_10312;
assign v_10320 = v_10317 | v_10319;
assign v_10322 = v_10316 | v_10321;
assign v_10324 = v_13810 | v_13811;
assign v_10330 = v_10327 | v_10328 | v_10329;
assign v_10332 = v_10326 | v_10331;
assign v_10338 = v_10335 | v_10336 | v_10337;
assign v_10340 = v_10334 | v_10339;
assign v_10345 = v_10342 | v_10343 | v_10344;
assign v_10349 = v_10347 | v_10348;
assign v_10350 = v_7739 | v_7737;
assign v_10355 = v_10351 | v_10352 | v_10353 | v_10354;
assign v_10359 = v_13812 | v_13813;
assign v_10365 = v_10362 | v_10363 | v_10364;
assign v_10367 = v_10361 | v_10366;
assign v_10373 = v_10370 | v_10371 | v_10372;
assign v_10375 = v_10369 | v_10374;
assign v_10380 = v_10377 | v_10378 | v_10379;
assign v_10384 = v_10382 | v_10383;
assign v_10385 = v_7820 | v_7818;
assign v_10390 = v_10386 | v_10387 | v_10388 | v_10389;
assign v_10394 = v_13814 | v_13815;
assign v_10400 = v_10397 | v_10398 | v_10399;
assign v_10402 = v_10396 | v_10401;
assign v_10408 = v_10405 | v_10406 | v_10407;
assign v_10410 = v_10404 | v_10409;
assign v_10415 = v_10412 | v_10413 | v_10414;
assign v_10419 = v_10417 | v_10418;
assign v_10420 = v_7901 | v_7899;
assign v_10425 = v_10421 | v_10422 | v_10423 | v_10424;
assign v_10429 = v_13816 | v_13817;
assign v_10435 = v_10432 | v_10433 | v_10434;
assign v_10437 = v_10431 | v_10436;
assign v_10443 = v_10440 | v_10441 | v_10442;
assign v_10445 = v_10439 | v_10444;
assign v_10450 = v_10447 | v_10448 | v_10449;
assign v_10454 = v_10452 | v_10453;
assign v_10455 = v_7982 | v_7980;
assign v_10460 = v_10456 | v_10457 | v_10458 | v_10459;
assign v_10464 = v_13818 | v_13819;
assign v_10470 = v_10467 | v_10468 | v_10469;
assign v_10472 = v_10466 | v_10471;
assign v_10478 = v_10475 | v_10476 | v_10477;
assign v_10480 = v_10474 | v_10479;
assign v_10485 = v_10482 | v_10483 | v_10484;
assign v_10489 = v_10487 | v_10488;
assign v_10490 = v_8063 | v_8061;
assign v_10495 = v_10491 | v_10492 | v_10493 | v_10494;
assign v_10499 = v_13820 | v_13821;
assign v_10505 = v_10502 | v_10503 | v_10504;
assign v_10507 = v_10501 | v_10506;
assign v_10513 = v_10510 | v_10511 | v_10512;
assign v_10515 = v_10509 | v_10514;
assign v_10520 = v_10517 | v_10518 | v_10519;
assign v_10524 = v_10522 | v_10523;
assign v_10525 = v_8144 | v_8142;
assign v_10530 = v_10526 | v_10527 | v_10528 | v_10529;
assign v_10534 = v_13822 | v_13823;
assign v_10540 = v_10537 | v_10538 | v_10539;
assign v_10542 = v_10536 | v_10541;
assign v_10548 = v_10545 | v_10546 | v_10547;
assign v_10550 = v_10544 | v_10549;
assign v_10555 = v_10552 | v_10553 | v_10554;
assign v_10559 = v_10557 | v_10558;
assign v_10560 = v_8225 | v_8223;
assign v_10565 = v_10561 | v_10562 | v_10563 | v_10564;
assign v_10569 = v_13824 | v_13825;
assign v_10577 = v_10575 | v_10576;
assign v_10578 = v_13826 | v_13827;
assign v_10582 = v_10579 | v_10580 | v_10581;
assign v_10584 = v_10572 | v_10573 | v_10574 | v_10583;
assign v_10587 = v_10571 | v_10585 | v_10586;
assign v_10589 = v_7160 | v_7162;
assign v_10592 = v_10588 | v_10590 | v_10591;
assign v_10593 = v_7174 | v_7176;
assign v_10599 = v_10596 | v_10597 | v_10598;
assign v_10601 = v_10595 | v_10600;
assign v_10603 = v_10594 | v_10602;
assign v_10604 = ~v_7199 | v_7201 | v_7203;
assign v_10607 = v_10605 | v_10606;
assign v_10616 = v_10614 | v_10615;
assign v_10618 = v_10612 | v_10613 | v_10617;
assign v_10623 = v_7246 | v_7248;
assign v_10626 = v_10624 | v_10625;
assign v_10629 = v_10627 | v_10628;
assign v_10631 = v_10620 | v_10621 | v_10622 | v_10630;
assign v_10637 = v_10633 | v_10634 | v_10635 | v_10636;
assign v_10639 = v_10619 | v_10632 | v_10638;
assign v_10641 = v_10608 | v_10609 | v_10610 | v_10611 | v_10640;
assign v_10650 = v_10648 | v_10649;
assign v_10652 = v_10646 | v_10647 | v_10651;
assign v_10657 = v_7311 | v_7313;
assign v_10660 = v_10658 | v_10659;
assign v_10663 = v_10661 | v_10662;
assign v_10665 = v_10654 | v_10655 | v_10656 | v_10664;
assign v_10671 = v_10667 | v_10668 | v_10669 | v_10670;
assign v_10673 = v_10653 | v_10666 | v_10672;
assign v_10675 = v_10642 | v_10643 | v_10644 | v_10645 | v_10674;
assign v_10682 = v_10680 | v_10681;
assign v_10683 = v_13828 | v_13829;
assign v_10687 = v_10684 | v_10685 | v_10686;
assign v_10689 = v_10677 | v_10678 | v_10679 | v_10688;
assign v_10692 = v_10676 | v_10690 | v_10691;
assign v_10697 = v_10694 | v_10696;
assign v_10699 = v_10693 | v_10698;
assign v_10703 = v_10701 | v_10702;
assign v_10704 = v_7436 | v_7438;
assign v_10707 = v_10700 | v_10705 | v_10706;
assign v_10712 = v_10708 | v_10709 | v_10710 | v_10711;
assign v_10717 = v_10714 | v_10716;
assign v_10719 = v_10713 | v_10718;
assign v_10723 = v_10721 | v_10722;
assign v_10724 = v_7494 | v_7496;
assign v_10727 = v_10720 | v_10725 | v_10726;
assign v_10735 = v_10733 | v_10734;
assign v_10737 = v_10732 | v_10736;
assign v_10739 = v_10731 | v_10738;
assign v_10741 = v_10730 | v_10740;
assign v_10743 = v_10729 | v_10742;
assign v_10745 = v_10728 | v_10744;
assign v_10750 = v_10748 | v_10749;
assign v_10756 = v_10752 | v_10753 | v_10754 | v_10755;
assign v_10758 = v_10751 | v_10757;
assign v_10762 = v_10746 | v_10747 | v_10759 | v_10760 | v_10761;
assign v_10768 = v_10765 | v_10767;
assign v_10770 = v_10764 | v_10769;
assign v_10772 = v_7596 | v_7598;
assign v_10776 = v_10774 | v_10775;
assign v_10779 = v_10777 | v_10778;
assign v_10786 = v_10783 | v_10785;
assign v_10788 = v_10782 | v_10787;
assign v_10790 = v_13830 | v_13831;
assign v_10796 = v_10793 | v_10794 | v_10795;
assign v_10798 = v_10792 | v_10797;
assign v_10804 = v_10801 | v_10802 | v_10803;
assign v_10806 = v_10800 | v_10805;
assign v_10811 = v_10808 | v_10809 | v_10810;
assign v_10815 = v_10813 | v_10814;
assign v_10816 = v_7739 | v_7737;
assign v_10821 = v_10817 | v_10818 | v_10819 | v_10820;
assign v_10825 = v_13832 | v_13833;
assign v_10831 = v_10828 | v_10829 | v_10830;
assign v_10833 = v_10827 | v_10832;
assign v_10839 = v_10836 | v_10837 | v_10838;
assign v_10841 = v_10835 | v_10840;
assign v_10846 = v_10843 | v_10844 | v_10845;
assign v_10850 = v_10848 | v_10849;
assign v_10851 = v_7820 | v_7818;
assign v_10856 = v_10852 | v_10853 | v_10854 | v_10855;
assign v_10860 = v_13834 | v_13835;
assign v_10866 = v_10863 | v_10864 | v_10865;
assign v_10868 = v_10862 | v_10867;
assign v_10874 = v_10871 | v_10872 | v_10873;
assign v_10876 = v_10870 | v_10875;
assign v_10881 = v_10878 | v_10879 | v_10880;
assign v_10885 = v_10883 | v_10884;
assign v_10886 = v_7901 | v_7899;
assign v_10891 = v_10887 | v_10888 | v_10889 | v_10890;
assign v_10895 = v_13836 | v_13837;
assign v_10901 = v_10898 | v_10899 | v_10900;
assign v_10903 = v_10897 | v_10902;
assign v_10909 = v_10906 | v_10907 | v_10908;
assign v_10911 = v_10905 | v_10910;
assign v_10916 = v_10913 | v_10914 | v_10915;
assign v_10920 = v_10918 | v_10919;
assign v_10921 = v_7982 | v_7980;
assign v_10926 = v_10922 | v_10923 | v_10924 | v_10925;
assign v_10930 = v_13838 | v_13839;
assign v_10936 = v_10933 | v_10934 | v_10935;
assign v_10938 = v_10932 | v_10937;
assign v_10944 = v_10941 | v_10942 | v_10943;
assign v_10946 = v_10940 | v_10945;
assign v_10951 = v_10948 | v_10949 | v_10950;
assign v_10955 = v_10953 | v_10954;
assign v_10956 = v_8063 | v_8061;
assign v_10961 = v_10957 | v_10958 | v_10959 | v_10960;
assign v_10965 = v_13840 | v_13841;
assign v_10971 = v_10968 | v_10969 | v_10970;
assign v_10973 = v_10967 | v_10972;
assign v_10979 = v_10976 | v_10977 | v_10978;
assign v_10981 = v_10975 | v_10980;
assign v_10986 = v_10983 | v_10984 | v_10985;
assign v_10990 = v_10988 | v_10989;
assign v_10991 = v_8144 | v_8142;
assign v_10996 = v_10992 | v_10993 | v_10994 | v_10995;
assign v_11000 = v_13842 | v_13843;
assign v_11006 = v_11003 | v_11004 | v_11005;
assign v_11008 = v_11002 | v_11007;
assign v_11014 = v_11011 | v_11012 | v_11013;
assign v_11016 = v_11010 | v_11015;
assign v_11021 = v_11018 | v_11019 | v_11020;
assign v_11025 = v_11023 | v_11024;
assign v_11026 = v_8225 | v_8223;
assign v_11031 = v_11027 | v_11028 | v_11029 | v_11030;
assign v_11035 = v_13844 | v_13845;
assign v_11042 = v_11040 | v_11041;
assign v_11043 = v_13846 | v_13847;
assign v_11047 = v_11044 | v_11045 | v_11046;
assign v_11049 = v_11037 | v_11038 | v_11039 | v_11048;
assign v_11052 = v_11036 | v_11050 | v_11051;
assign v_11054 = v_7160 | v_7162;
assign v_11057 = v_11053 | v_11055 | v_11056;
assign v_11058 = v_7174 | v_7176;
assign v_11064 = v_11061 | v_11062 | v_11063;
assign v_11066 = v_11060 | v_11065;
assign v_11068 = v_11059 | v_11067;
assign v_11069 = ~v_7199 | v_7201 | v_7203;
assign v_11072 = v_11070 | v_11071;
assign v_11081 = v_11079 | v_11080;
assign v_11083 = v_11077 | v_11078 | v_11082;
assign v_11088 = v_7246 | v_7248;
assign v_11091 = v_11089 | v_11090;
assign v_11094 = v_11092 | v_11093;
assign v_11096 = v_11085 | v_11086 | v_11087 | v_11095;
assign v_11102 = v_11098 | v_11099 | v_11100 | v_11101;
assign v_11104 = v_11084 | v_11097 | v_11103;
assign v_11106 = v_11073 | v_11074 | v_11075 | v_11076 | v_11105;
assign v_11115 = v_11113 | v_11114;
assign v_11117 = v_11111 | v_11112 | v_11116;
assign v_11122 = v_7311 | v_7313;
assign v_11125 = v_11123 | v_11124;
assign v_11128 = v_11126 | v_11127;
assign v_11130 = v_11119 | v_11120 | v_11121 | v_11129;
assign v_11136 = v_11132 | v_11133 | v_11134 | v_11135;
assign v_11138 = v_11118 | v_11131 | v_11137;
assign v_11140 = v_11107 | v_11108 | v_11109 | v_11110 | v_11139;
assign v_11147 = v_11145 | v_11146;
assign v_11148 = v_13848 | v_13849;
assign v_11152 = v_11149 | v_11150 | v_11151;
assign v_11154 = v_11142 | v_11143 | v_11144 | v_11153;
assign v_11157 = v_11141 | v_11155 | v_11156;
assign v_11162 = v_11159 | v_11161;
assign v_11164 = v_11158 | v_11163;
assign v_11168 = v_11166 | v_11167;
assign v_11169 = v_7436 | v_7438;
assign v_11172 = v_11165 | v_11170 | v_11171;
assign v_11177 = v_11173 | v_11174 | v_11175 | v_11176;
assign v_11182 = v_11179 | v_11181;
assign v_11184 = v_11178 | v_11183;
assign v_11188 = v_11186 | v_11187;
assign v_11189 = v_7494 | v_7496;
assign v_11192 = v_11185 | v_11190 | v_11191;
assign v_11200 = v_11198 | v_11199;
assign v_11202 = v_11197 | v_11201;
assign v_11204 = v_11196 | v_11203;
assign v_11206 = v_11195 | v_11205;
assign v_11208 = v_11194 | v_11207;
assign v_11210 = v_11193 | v_11209;
assign v_11215 = v_11213 | v_11214;
assign v_11221 = v_11217 | v_11218 | v_11219 | v_11220;
assign v_11223 = v_11216 | v_11222;
assign v_11227 = v_11211 | v_11212 | v_11224 | v_11225 | v_11226;
assign v_11233 = v_11230 | v_11232;
assign v_11235 = v_11229 | v_11234;
assign v_11237 = v_7596 | v_7598;
assign v_11241 = v_11239 | v_11240;
assign v_11244 = v_11242 | v_11243;
assign v_11251 = v_11248 | v_11250;
assign v_11253 = v_11247 | v_11252;
assign v_11255 = v_13850 | v_13851;
assign v_11261 = v_11258 | v_11259 | v_11260;
assign v_11263 = v_11257 | v_11262;
assign v_11269 = v_11266 | v_11267 | v_11268;
assign v_11271 = v_11265 | v_11270;
assign v_11276 = v_11273 | v_11274 | v_11275;
assign v_11280 = v_11278 | v_11279;
assign v_11281 = v_7739 | v_7737;
assign v_11286 = v_11282 | v_11283 | v_11284 | v_11285;
assign v_11290 = v_13852 | v_13853;
assign v_11296 = v_11293 | v_11294 | v_11295;
assign v_11298 = v_11292 | v_11297;
assign v_11304 = v_11301 | v_11302 | v_11303;
assign v_11306 = v_11300 | v_11305;
assign v_11311 = v_11308 | v_11309 | v_11310;
assign v_11315 = v_11313 | v_11314;
assign v_11316 = v_7820 | v_7818;
assign v_11321 = v_11317 | v_11318 | v_11319 | v_11320;
assign v_11325 = v_13854 | v_13855;
assign v_11331 = v_11328 | v_11329 | v_11330;
assign v_11333 = v_11327 | v_11332;
assign v_11339 = v_11336 | v_11337 | v_11338;
assign v_11341 = v_11335 | v_11340;
assign v_11346 = v_11343 | v_11344 | v_11345;
assign v_11350 = v_11348 | v_11349;
assign v_11351 = v_7901 | v_7899;
assign v_11356 = v_11352 | v_11353 | v_11354 | v_11355;
assign v_11360 = v_13856 | v_13857;
assign v_11366 = v_11363 | v_11364 | v_11365;
assign v_11368 = v_11362 | v_11367;
assign v_11374 = v_11371 | v_11372 | v_11373;
assign v_11376 = v_11370 | v_11375;
assign v_11381 = v_11378 | v_11379 | v_11380;
assign v_11385 = v_11383 | v_11384;
assign v_11386 = v_7982 | v_7980;
assign v_11391 = v_11387 | v_11388 | v_11389 | v_11390;
assign v_11395 = v_13858 | v_13859;
assign v_11401 = v_11398 | v_11399 | v_11400;
assign v_11403 = v_11397 | v_11402;
assign v_11409 = v_11406 | v_11407 | v_11408;
assign v_11411 = v_11405 | v_11410;
assign v_11416 = v_11413 | v_11414 | v_11415;
assign v_11420 = v_11418 | v_11419;
assign v_11421 = v_8063 | v_8061;
assign v_11426 = v_11422 | v_11423 | v_11424 | v_11425;
assign v_11430 = v_13860 | v_13861;
assign v_11436 = v_11433 | v_11434 | v_11435;
assign v_11438 = v_11432 | v_11437;
assign v_11444 = v_11441 | v_11442 | v_11443;
assign v_11446 = v_11440 | v_11445;
assign v_11451 = v_11448 | v_11449 | v_11450;
assign v_11455 = v_11453 | v_11454;
assign v_11456 = v_8144 | v_8142;
assign v_11461 = v_11457 | v_11458 | v_11459 | v_11460;
assign v_11465 = v_13862 | v_13863;
assign v_11471 = v_11468 | v_11469 | v_11470;
assign v_11473 = v_11467 | v_11472;
assign v_11479 = v_11476 | v_11477 | v_11478;
assign v_11481 = v_11475 | v_11480;
assign v_11486 = v_11483 | v_11484 | v_11485;
assign v_11490 = v_11488 | v_11489;
assign v_11491 = v_8225 | v_8223;
assign v_11496 = v_11492 | v_11493 | v_11494 | v_11495;
assign v_11500 = v_13864 | v_13865;
assign v_11508 = v_11506 | v_11507;
assign v_11509 = v_13866 | v_13867;
assign v_11513 = v_11510 | v_11511 | v_11512;
assign v_11515 = v_11503 | v_11504 | v_11505 | v_11514;
assign v_11518 = v_11502 | v_11516 | v_11517;
assign v_11520 = v_7160 | v_7162;
assign v_11523 = v_11519 | v_11521 | v_11522;
assign v_11524 = v_7174 | v_7176;
assign v_11530 = v_11527 | v_11528 | v_11529;
assign v_11532 = v_11526 | v_11531;
assign v_11534 = v_11525 | v_11533;
assign v_11535 = ~v_7199 | v_7201 | v_7203;
assign v_11538 = v_11536 | v_11537;
assign v_11547 = v_11545 | v_11546;
assign v_11549 = v_11543 | v_11544 | v_11548;
assign v_11554 = v_7246 | v_7248;
assign v_11557 = v_11555 | v_11556;
assign v_11560 = v_11558 | v_11559;
assign v_11562 = v_11551 | v_11552 | v_11553 | v_11561;
assign v_11568 = v_11564 | v_11565 | v_11566 | v_11567;
assign v_11570 = v_11550 | v_11563 | v_11569;
assign v_11572 = v_11539 | v_11540 | v_11541 | v_11542 | v_11571;
assign v_11581 = v_11579 | v_11580;
assign v_11583 = v_11577 | v_11578 | v_11582;
assign v_11588 = v_7311 | v_7313;
assign v_11591 = v_11589 | v_11590;
assign v_11594 = v_11592 | v_11593;
assign v_11596 = v_11585 | v_11586 | v_11587 | v_11595;
assign v_11602 = v_11598 | v_11599 | v_11600 | v_11601;
assign v_11604 = v_11584 | v_11597 | v_11603;
assign v_11606 = v_11573 | v_11574 | v_11575 | v_11576 | v_11605;
assign v_11613 = v_11611 | v_11612;
assign v_11614 = v_13868 | v_13869;
assign v_11618 = v_11615 | v_11616 | v_11617;
assign v_11620 = v_11608 | v_11609 | v_11610 | v_11619;
assign v_11623 = v_11607 | v_11621 | v_11622;
assign v_11628 = v_11625 | v_11627;
assign v_11630 = v_11624 | v_11629;
assign v_11634 = v_11632 | v_11633;
assign v_11635 = v_7436 | v_7438;
assign v_11638 = v_11631 | v_11636 | v_11637;
assign v_11643 = v_11639 | v_11640 | v_11641 | v_11642;
assign v_11648 = v_11645 | v_11647;
assign v_11650 = v_11644 | v_11649;
assign v_11654 = v_11652 | v_11653;
assign v_11655 = v_7494 | v_7496;
assign v_11658 = v_11651 | v_11656 | v_11657;
assign v_11666 = v_11664 | v_11665;
assign v_11668 = v_11663 | v_11667;
assign v_11670 = v_11662 | v_11669;
assign v_11672 = v_11661 | v_11671;
assign v_11674 = v_11660 | v_11673;
assign v_11676 = v_11659 | v_11675;
assign v_11681 = v_11679 | v_11680;
assign v_11687 = v_11683 | v_11684 | v_11685 | v_11686;
assign v_11689 = v_11682 | v_11688;
assign v_11693 = v_11677 | v_11678 | v_11690 | v_11691 | v_11692;
assign v_11699 = v_11696 | v_11698;
assign v_11701 = v_11695 | v_11700;
assign v_11703 = v_7596 | v_7598;
assign v_11707 = v_11705 | v_11706;
assign v_11710 = v_11708 | v_11709;
assign v_11717 = v_11714 | v_11716;
assign v_11719 = v_11713 | v_11718;
assign v_11721 = v_13870 | v_13871;
assign v_11727 = v_11724 | v_11725 | v_11726;
assign v_11729 = v_11723 | v_11728;
assign v_11735 = v_11732 | v_11733 | v_11734;
assign v_11737 = v_11731 | v_11736;
assign v_11742 = v_11739 | v_11740 | v_11741;
assign v_11746 = v_11744 | v_11745;
assign v_11747 = v_7739 | v_7737;
assign v_11752 = v_11748 | v_11749 | v_11750 | v_11751;
assign v_11756 = v_13872 | v_13873;
assign v_11762 = v_11759 | v_11760 | v_11761;
assign v_11764 = v_11758 | v_11763;
assign v_11770 = v_11767 | v_11768 | v_11769;
assign v_11772 = v_11766 | v_11771;
assign v_11777 = v_11774 | v_11775 | v_11776;
assign v_11781 = v_11779 | v_11780;
assign v_11782 = v_7820 | v_7818;
assign v_11787 = v_11783 | v_11784 | v_11785 | v_11786;
assign v_11791 = v_13874 | v_13875;
assign v_11797 = v_11794 | v_11795 | v_11796;
assign v_11799 = v_11793 | v_11798;
assign v_11805 = v_11802 | v_11803 | v_11804;
assign v_11807 = v_11801 | v_11806;
assign v_11812 = v_11809 | v_11810 | v_11811;
assign v_11816 = v_11814 | v_11815;
assign v_11817 = v_7901 | v_7899;
assign v_11822 = v_11818 | v_11819 | v_11820 | v_11821;
assign v_11826 = v_13876 | v_13877;
assign v_11832 = v_11829 | v_11830 | v_11831;
assign v_11834 = v_11828 | v_11833;
assign v_11840 = v_11837 | v_11838 | v_11839;
assign v_11842 = v_11836 | v_11841;
assign v_11847 = v_11844 | v_11845 | v_11846;
assign v_11851 = v_11849 | v_11850;
assign v_11852 = v_7982 | v_7980;
assign v_11857 = v_11853 | v_11854 | v_11855 | v_11856;
assign v_11861 = v_13878 | v_13879;
assign v_11867 = v_11864 | v_11865 | v_11866;
assign v_11869 = v_11863 | v_11868;
assign v_11875 = v_11872 | v_11873 | v_11874;
assign v_11877 = v_11871 | v_11876;
assign v_11882 = v_11879 | v_11880 | v_11881;
assign v_11886 = v_11884 | v_11885;
assign v_11887 = v_8063 | v_8061;
assign v_11892 = v_11888 | v_11889 | v_11890 | v_11891;
assign v_11896 = v_13880 | v_13881;
assign v_11902 = v_11899 | v_11900 | v_11901;
assign v_11904 = v_11898 | v_11903;
assign v_11910 = v_11907 | v_11908 | v_11909;
assign v_11912 = v_11906 | v_11911;
assign v_11917 = v_11914 | v_11915 | v_11916;
assign v_11921 = v_11919 | v_11920;
assign v_11922 = v_8144 | v_8142;
assign v_11927 = v_11923 | v_11924 | v_11925 | v_11926;
assign v_11931 = v_13882 | v_13883;
assign v_11937 = v_11934 | v_11935 | v_11936;
assign v_11939 = v_11933 | v_11938;
assign v_11945 = v_11942 | v_11943 | v_11944;
assign v_11947 = v_11941 | v_11946;
assign v_11952 = v_11949 | v_11950 | v_11951;
assign v_11956 = v_11954 | v_11955;
assign v_11957 = v_8225 | v_8223;
assign v_11962 = v_11958 | v_11959 | v_11960 | v_11961;
assign v_11966 = v_13884 | v_13885;
assign v_11969 = v_11968 | ~v_8276;
assign v_11975 = v_11971 | v_11973 | v_11974;
assign v_11977 = v_7160 | v_7162;
assign v_11980 = v_11976 | v_11978 | v_11979;
assign v_11981 = v_7174 | v_7176;
assign v_11987 = v_11984 | v_11985 | v_11986;
assign v_11989 = v_11983 | v_11988;
assign v_11991 = v_11982 | v_11990;
assign v_11992 = ~v_7199 | v_7201 | v_7203;
assign v_11995 = v_11993 | v_11994;
assign v_11997 = v_11970 | v_11996;
assign v_12006 = v_12004 | v_12005;
assign v_12008 = v_12002 | v_12003 | v_12007;
assign v_12013 = v_7246 | v_7248;
assign v_12016 = v_12014 | v_12015;
assign v_12019 = v_12017 | v_12018;
assign v_12021 = v_12010 | v_12011 | v_12012 | v_12020;
assign v_12027 = v_12023 | v_12024 | v_12025 | v_12026;
assign v_12029 = v_12009 | v_12022 | v_12028;
assign v_12031 = v_11998 | v_11999 | v_12000 | v_12001 | v_12030;
assign v_12040 = v_12038 | v_12039;
assign v_12042 = v_12036 | v_12037 | v_12041;
assign v_12047 = v_7311 | v_7313;
assign v_12050 = v_12048 | v_12049;
assign v_12053 = v_12051 | v_12052;
assign v_12055 = v_12044 | v_12045 | v_12046 | v_12054;
assign v_12061 = v_12057 | v_12058 | v_12059 | v_12060;
assign v_12063 = v_12043 | v_12056 | v_12062;
assign v_12065 = v_12032 | v_12033 | v_12034 | v_12035 | v_12064;
assign v_12070 = v_12066 | v_12068 | v_12069;
assign v_12073 = v_12071 | v_12072;
assign v_12077 = v_12075 | v_12076;
assign v_12078 = v_7436 | v_7438;
assign v_12081 = v_12074 | v_12079 | v_12080;
assign v_12086 = v_12082 | v_12083 | v_12084 | v_12085;
assign v_12089 = v_12087 | v_12088;
assign v_12093 = v_12091 | v_12092;
assign v_12094 = v_7494 | v_7496;
assign v_12097 = v_12090 | v_12095 | v_12096;
assign v_12105 = v_12103 | v_12104;
assign v_12107 = v_12102 | v_12106;
assign v_12109 = v_12101 | v_12108;
assign v_12111 = v_12100 | v_12110;
assign v_12113 = v_12099 | v_12112;
assign v_12115 = v_12098 | v_12114;
assign v_12120 = v_12118 | v_12119;
assign v_12126 = v_12122 | v_12123 | v_12124 | v_12125;
assign v_12128 = v_12121 | v_12127;
assign v_12132 = v_12116 | v_12117 | v_12129 | v_12130 | v_12131;
assign v_12136 = v_12134 | v_12135;
assign v_12138 = v_7596 | v_7598;
assign v_12142 = v_12140 | v_12141;
assign v_12145 = v_12143 | v_12144;
assign v_12150 = v_12148 | v_12149;
assign v_12152 = v_13886 | v_13887;
assign v_12158 = v_12155 | v_12156 | v_12157;
assign v_12160 = v_12154 | v_12159;
assign v_12166 = v_12163 | v_12164 | v_12165;
assign v_12168 = v_12162 | v_12167;
assign v_12173 = v_12170 | v_12171 | v_12172;
assign v_12177 = v_12175 | v_12176;
assign v_12178 = v_7739 | v_7737;
assign v_12183 = v_12179 | v_12180 | v_12181 | v_12182;
assign v_12187 = v_13888 | v_13889;
assign v_12193 = v_12190 | v_12191 | v_12192;
assign v_12195 = v_12189 | v_12194;
assign v_12201 = v_12198 | v_12199 | v_12200;
assign v_12203 = v_12197 | v_12202;
assign v_12208 = v_12205 | v_12206 | v_12207;
assign v_12212 = v_12210 | v_12211;
assign v_12213 = v_7820 | v_7818;
assign v_12218 = v_12214 | v_12215 | v_12216 | v_12217;
assign v_12222 = v_13890 | v_13891;
assign v_12228 = v_12225 | v_12226 | v_12227;
assign v_12230 = v_12224 | v_12229;
assign v_12236 = v_12233 | v_12234 | v_12235;
assign v_12238 = v_12232 | v_12237;
assign v_12243 = v_12240 | v_12241 | v_12242;
assign v_12247 = v_12245 | v_12246;
assign v_12248 = v_7901 | v_7899;
assign v_12253 = v_12249 | v_12250 | v_12251 | v_12252;
assign v_12257 = v_13892 | v_13893;
assign v_12263 = v_12260 | v_12261 | v_12262;
assign v_12265 = v_12259 | v_12264;
assign v_12271 = v_12268 | v_12269 | v_12270;
assign v_12273 = v_12267 | v_12272;
assign v_12278 = v_12275 | v_12276 | v_12277;
assign v_12282 = v_12280 | v_12281;
assign v_12283 = v_7982 | v_7980;
assign v_12288 = v_12284 | v_12285 | v_12286 | v_12287;
assign v_12292 = v_13894 | v_13895;
assign v_12298 = v_12295 | v_12296 | v_12297;
assign v_12300 = v_12294 | v_12299;
assign v_12306 = v_12303 | v_12304 | v_12305;
assign v_12308 = v_12302 | v_12307;
assign v_12313 = v_12310 | v_12311 | v_12312;
assign v_12317 = v_12315 | v_12316;
assign v_12318 = v_8063 | v_8061;
assign v_12323 = v_12319 | v_12320 | v_12321 | v_12322;
assign v_12327 = v_13896 | v_13897;
assign v_12333 = v_12330 | v_12331 | v_12332;
assign v_12335 = v_12329 | v_12334;
assign v_12341 = v_12338 | v_12339 | v_12340;
assign v_12343 = v_12337 | v_12342;
assign v_12348 = v_12345 | v_12346 | v_12347;
assign v_12352 = v_12350 | v_12351;
assign v_12353 = v_8144 | v_8142;
assign v_12358 = v_12354 | v_12355 | v_12356 | v_12357;
assign v_12362 = v_13898 | v_13899;
assign v_12368 = v_12365 | v_12366 | v_12367;
assign v_12370 = v_12364 | v_12369;
assign v_12376 = v_12373 | v_12374 | v_12375;
assign v_12378 = v_12372 | v_12377;
assign v_12383 = v_12380 | v_12381 | v_12382;
assign v_12387 = v_12385 | v_12386;
assign v_12388 = v_8225 | v_8223;
assign v_12393 = v_12389 | v_12390 | v_12391 | v_12392;
assign v_12397 = v_13900 | v_13901;
assign v_12405 = v_12403 | v_12404;
assign v_12406 = v_13902 | v_13903;
assign v_12410 = v_12407 | v_12408 | v_12409;
assign v_12412 = v_12400 | v_12401 | v_12402 | v_12411;
assign v_12415 = v_12399 | v_12413 | v_12414;
assign v_12417 = v_7160 | v_7162;
assign v_12420 = v_12416 | v_12418 | v_12419;
assign v_12421 = v_7174 | v_7176;
assign v_12427 = v_12424 | v_12425 | v_12426;
assign v_12429 = v_12423 | v_12428;
assign v_12431 = v_12422 | v_12430;
assign v_12432 = ~v_7199 | v_7201 | v_7203;
assign v_12435 = v_12433 | v_12434;
assign v_12444 = v_12442 | v_12443;
assign v_12446 = v_12440 | v_12441 | v_12445;
assign v_12451 = v_7246 | v_7248;
assign v_12454 = v_12452 | v_12453;
assign v_12457 = v_12455 | v_12456;
assign v_12459 = v_12448 | v_12449 | v_12450 | v_12458;
assign v_12465 = v_12461 | v_12462 | v_12463 | v_12464;
assign v_12467 = v_12447 | v_12460 | v_12466;
assign v_12469 = v_12436 | v_12437 | v_12438 | v_12439 | v_12468;
assign v_12478 = v_12476 | v_12477;
assign v_12480 = v_12474 | v_12475 | v_12479;
assign v_12485 = v_7311 | v_7313;
assign v_12488 = v_12486 | v_12487;
assign v_12491 = v_12489 | v_12490;
assign v_12493 = v_12482 | v_12483 | v_12484 | v_12492;
assign v_12499 = v_12495 | v_12496 | v_12497 | v_12498;
assign v_12501 = v_12481 | v_12494 | v_12500;
assign v_12503 = v_12470 | v_12471 | v_12472 | v_12473 | v_12502;
assign v_12510 = v_12508 | v_12509;
assign v_12511 = v_13904 | v_13905;
assign v_12515 = v_12512 | v_12513 | v_12514;
assign v_12517 = v_12505 | v_12506 | v_12507 | v_12516;
assign v_12520 = v_12504 | v_12518 | v_12519;
assign v_12525 = v_12522 | v_12524;
assign v_12527 = v_12521 | v_12526;
assign v_12531 = v_12529 | v_12530;
assign v_12532 = v_7436 | v_7438;
assign v_12535 = v_12528 | v_12533 | v_12534;
assign v_12540 = v_12536 | v_12537 | v_12538 | v_12539;
assign v_12545 = v_12542 | v_12544;
assign v_12547 = v_12541 | v_12546;
assign v_12551 = v_12549 | v_12550;
assign v_12552 = v_7494 | v_7496;
assign v_12555 = v_12548 | v_12553 | v_12554;
assign v_12563 = v_12561 | v_12562;
assign v_12565 = v_12560 | v_12564;
assign v_12567 = v_12559 | v_12566;
assign v_12569 = v_12558 | v_12568;
assign v_12571 = v_12557 | v_12570;
assign v_12573 = v_12556 | v_12572;
assign v_12578 = v_12576 | v_12577;
assign v_12584 = v_12580 | v_12581 | v_12582 | v_12583;
assign v_12586 = v_12579 | v_12585;
assign v_12590 = v_12574 | v_12575 | v_12587 | v_12588 | v_12589;
assign v_12596 = v_12593 | v_12595;
assign v_12598 = v_12592 | v_12597;
assign v_12600 = v_7596 | v_7598;
assign v_12604 = v_12602 | v_12603;
assign v_12607 = v_12605 | v_12606;
assign v_12614 = v_12611 | v_12613;
assign v_12616 = v_12610 | v_12615;
assign v_12618 = v_13906 | v_13907;
assign v_12624 = v_12621 | v_12622 | v_12623;
assign v_12626 = v_12620 | v_12625;
assign v_12632 = v_12629 | v_12630 | v_12631;
assign v_12634 = v_12628 | v_12633;
assign v_12639 = v_12636 | v_12637 | v_12638;
assign v_12643 = v_12641 | v_12642;
assign v_12644 = v_7739 | v_7737;
assign v_12649 = v_12645 | v_12646 | v_12647 | v_12648;
assign v_12653 = v_13908 | v_13909;
assign v_12659 = v_12656 | v_12657 | v_12658;
assign v_12661 = v_12655 | v_12660;
assign v_12667 = v_12664 | v_12665 | v_12666;
assign v_12669 = v_12663 | v_12668;
assign v_12674 = v_12671 | v_12672 | v_12673;
assign v_12678 = v_12676 | v_12677;
assign v_12679 = v_7820 | v_7818;
assign v_12684 = v_12680 | v_12681 | v_12682 | v_12683;
assign v_12688 = v_13910 | v_13911;
assign v_12694 = v_12691 | v_12692 | v_12693;
assign v_12696 = v_12690 | v_12695;
assign v_12702 = v_12699 | v_12700 | v_12701;
assign v_12704 = v_12698 | v_12703;
assign v_12709 = v_12706 | v_12707 | v_12708;
assign v_12713 = v_12711 | v_12712;
assign v_12714 = v_7901 | v_7899;
assign v_12719 = v_12715 | v_12716 | v_12717 | v_12718;
assign v_12723 = v_13912 | v_13913;
assign v_12729 = v_12726 | v_12727 | v_12728;
assign v_12731 = v_12725 | v_12730;
assign v_12737 = v_12734 | v_12735 | v_12736;
assign v_12739 = v_12733 | v_12738;
assign v_12744 = v_12741 | v_12742 | v_12743;
assign v_12748 = v_12746 | v_12747;
assign v_12749 = v_7982 | v_7980;
assign v_12754 = v_12750 | v_12751 | v_12752 | v_12753;
assign v_12758 = v_13914 | v_13915;
assign v_12764 = v_12761 | v_12762 | v_12763;
assign v_12766 = v_12760 | v_12765;
assign v_12772 = v_12769 | v_12770 | v_12771;
assign v_12774 = v_12768 | v_12773;
assign v_12779 = v_12776 | v_12777 | v_12778;
assign v_12783 = v_12781 | v_12782;
assign v_12784 = v_8063 | v_8061;
assign v_12789 = v_12785 | v_12786 | v_12787 | v_12788;
assign v_12793 = v_13916 | v_13917;
assign v_12799 = v_12796 | v_12797 | v_12798;
assign v_12801 = v_12795 | v_12800;
assign v_12807 = v_12804 | v_12805 | v_12806;
assign v_12809 = v_12803 | v_12808;
assign v_12814 = v_12811 | v_12812 | v_12813;
assign v_12818 = v_12816 | v_12817;
assign v_12819 = v_8144 | v_8142;
assign v_12824 = v_12820 | v_12821 | v_12822 | v_12823;
assign v_12828 = v_13918 | v_13919;
assign v_12834 = v_12831 | v_12832 | v_12833;
assign v_12836 = v_12830 | v_12835;
assign v_12842 = v_12839 | v_12840 | v_12841;
assign v_12844 = v_12838 | v_12843;
assign v_12849 = v_12846 | v_12847 | v_12848;
assign v_12853 = v_12851 | v_12852;
assign v_12854 = v_8225 | v_8223;
assign v_12859 = v_12855 | v_12856 | v_12857 | v_12858;
assign v_12863 = v_13920 | v_13921;
assign v_13414 = v_233 | v_235 | v_238 | v_240 | v_242;
assign v_13415 = v_244 | v_246 | v_248 | v_252 | v_253;
assign v_13416 = v_259;
assign v_13417 = v_393 | v_395 | v_397 | v_399 | v_401;
assign v_13418 = v_402;
assign v_13419 = v_347 | v_349 | v_351 | v_358 | v_407;
assign v_13420 = v_408;
assign v_13421 = v_458 | v_460 | v_462 | v_464 | v_466;
assign v_13422 = v_467;
assign v_13423 = v_412 | v_414 | v_416 | v_423 | v_472;
assign v_13424 = v_473;
assign v_13425 = v_497 | v_499 | v_502 | v_504 | v_506;
assign v_13426 = v_508 | v_510 | v_512 | v_516 | v_517;
assign v_13427 = v_523;
assign v_13428 = ~v_669 | v_671 | v_673 | v_676 | v_681;
assign v_13429 = v_683 | v_701 | v_702;
assign v_13430 = ~v_705 | v_725 | v_730 | v_732 | v_774;
assign v_13431 = v_793 | v_794 | v_795;
assign v_13432 = v_816 | v_818 | v_839 | v_841 | v_862;
assign v_13433 = v_864 | v_871 | v_873 | v_874 | v_875;
assign v_13434 = v_876;
assign v_13435 = v_897 | v_899 | v_920 | v_922 | v_943;
assign v_13436 = v_945 | v_952 | v_954 | v_955 | v_956;
assign v_13437 = v_957;
assign v_13438 = v_978 | v_980 | v_1001 | v_1003 | v_1024;
assign v_13439 = v_1026 | v_1033 | v_1035 | v_1036 | v_1037;
assign v_13440 = v_1038;
assign v_13441 = v_1059 | v_1061 | v_1082 | v_1084 | v_1105;
assign v_13442 = v_1107 | v_1114 | v_1116 | v_1117 | v_1118;
assign v_13443 = v_1119;
assign v_13444 = v_1140 | v_1142 | v_1163 | v_1165 | v_1186;
assign v_13445 = v_1188 | v_1195 | v_1197 | v_1198 | v_1199;
assign v_13446 = v_1200;
assign v_13447 = v_1221 | v_1223 | v_1244 | v_1246 | v_1267;
assign v_13448 = v_1269 | v_1276 | v_1278 | v_1279 | v_1280;
assign v_13449 = v_1281;
assign v_13450 = v_1302 | v_1304 | v_1325 | v_1327 | v_1348;
assign v_13451 = v_1350 | v_1357 | v_1359 | v_1360 | v_1361;
assign v_13452 = v_1362;
assign v_13453 = v_1383 | v_1385 | v_1406 | v_1408 | v_1429;
assign v_13454 = v_1431 | v_1438 | v_1440 | v_1441 | v_1442;
assign v_13455 = v_1443;
assign v_13456 = v_1464 | v_1466 | v_1487 | v_1489 | v_1510;
assign v_13457 = v_1512 | v_1519 | v_1521 | v_1522 | v_1523;
assign v_13458 = v_1524;
assign v_13459 = v_233 | v_235 | v_238 | v_240 | v_242;
assign v_13460 = v_244 | v_246 | v_248;
assign v_13461 = v_497 | v_499 | v_502 | v_504 | v_506;
assign v_13462 = v_508 | v_510 | v_512;
assign v_13463 = v_1746 | v_1750 | v_1752 | v_1759 | v_1760;
assign v_13464 = v_1765;
assign v_13465 = v_1767 | v_1776 | v_1785 | v_1791 | v_1802;
assign v_13466 = v_1803 | v_1804;
assign v_13467 = v_1806 | v_1815 | v_1824 | v_1830 | v_1841;
assign v_13468 = v_1842 | v_1843;
assign v_13469 = v_1845 | v_1854 | v_1863 | v_1869 | v_1880;
assign v_13470 = v_1881 | v_1882;
assign v_13471 = v_1884 | v_1893 | v_1902 | v_1908 | v_1919;
assign v_13472 = v_1920 | v_1921;
assign v_13473 = v_1923 | v_1932 | v_1941 | v_1947 | v_1958;
assign v_13474 = v_1959 | v_1960;
assign v_13475 = v_1962 | v_1971 | v_1980 | v_1986 | v_1997;
assign v_13476 = v_1998 | v_1999;
assign v_13477 = v_2001 | v_2010 | v_2019 | v_2025 | v_2036;
assign v_13478 = v_2037 | v_2038;
assign v_13479 = v_2040 | v_2049 | v_2058 | v_2064 | v_2075;
assign v_13480 = v_2076 | v_2077;
assign v_13481 = v_2079 | v_2088 | v_2097 | v_2103 | v_2114;
assign v_13482 = v_2115 | v_2116;
assign v_13483 = v_2285 | v_2289 | v_2291 | v_2298 | v_2299;
assign v_13484 = v_2303;
assign v_13485 = v_2305 | v_2313 | v_2321 | v_2326 | v_2336;
assign v_13486 = v_2337 | v_2338;
assign v_13487 = v_2340 | v_2348 | v_2356 | v_2361 | v_2371;
assign v_13488 = v_2372 | v_2373;
assign v_13489 = v_2375 | v_2383 | v_2391 | v_2396 | v_2406;
assign v_13490 = v_2407 | v_2408;
assign v_13491 = v_2410 | v_2418 | v_2426 | v_2431 | v_2441;
assign v_13492 = v_2442 | v_2443;
assign v_13493 = v_2445 | v_2453 | v_2461 | v_2466 | v_2476;
assign v_13494 = v_2477 | v_2478;
assign v_13495 = v_2480 | v_2488 | v_2496 | v_2501 | v_2511;
assign v_13496 = v_2512 | v_2513;
assign v_13497 = v_2515 | v_2523 | v_2531 | v_2536 | v_2546;
assign v_13498 = v_2547 | v_2548;
assign v_13499 = v_2550 | v_2558 | v_2566 | v_2571 | v_2581;
assign v_13500 = v_2582 | v_2583;
assign v_13501 = v_2585 | v_2593 | v_2601 | v_2606 | v_2616;
assign v_13502 = v_2617 | v_2618;
assign v_13503 = v_233 | v_235 | v_238 | v_240 | v_242;
assign v_13504 = v_244 | v_246 | v_248;
assign v_13505 = v_497 | v_499 | v_502 | v_504 | v_506;
assign v_13506 = v_508 | v_510 | v_512;
assign v_13507 = v_2812 | v_2820 | v_2822 | v_2829 | v_2830;
assign v_13508 = v_2838;
assign v_13509 = v_2840 | v_2848 | v_2856 | v_2861 | v_2871;
assign v_13510 = v_2872 | v_2873;
assign v_13511 = v_2875 | v_2883 | v_2891 | v_2896 | v_2906;
assign v_13512 = v_2907 | v_2908;
assign v_13513 = v_2910 | v_2918 | v_2926 | v_2931 | v_2941;
assign v_13514 = v_2942 | v_2943;
assign v_13515 = v_2945 | v_2953 | v_2961 | v_2966 | v_2976;
assign v_13516 = v_2977 | v_2978;
assign v_13517 = v_2980 | v_2988 | v_2996 | v_3001 | v_3011;
assign v_13518 = v_3012 | v_3013;
assign v_13519 = v_3015 | v_3023 | v_3031 | v_3036 | v_3046;
assign v_13520 = v_3047 | v_3048;
assign v_13521 = v_3050 | v_3058 | v_3066 | v_3071 | v_3081;
assign v_13522 = v_3082 | v_3083;
assign v_13523 = v_3085 | v_3093 | v_3101 | v_3106 | v_3116;
assign v_13524 = v_3117 | v_3118;
assign v_13525 = v_3120 | v_3128 | v_3136 | v_3141 | v_3151;
assign v_13526 = v_3152 | v_3153;
assign v_13527 = v_233 | v_235 | v_238 | v_240 | v_242;
assign v_13528 = v_244 | v_246 | v_248;
assign v_13529 = v_497 | v_499 | v_502 | v_504 | v_506;
assign v_13530 = v_508 | v_510 | v_512;
assign v_13531 = v_3345 | v_3353 | v_3355 | v_3362 | v_3363;
assign v_13532 = v_3371;
assign v_13533 = v_3373 | v_3381 | v_3389 | v_3394 | v_3404;
assign v_13534 = v_3405 | v_3406;
assign v_13535 = v_3408 | v_3416 | v_3424 | v_3429 | v_3439;
assign v_13536 = v_3440 | v_3441;
assign v_13537 = v_3443 | v_3451 | v_3459 | v_3464 | v_3474;
assign v_13538 = v_3475 | v_3476;
assign v_13539 = v_3478 | v_3486 | v_3494 | v_3499 | v_3509;
assign v_13540 = v_3510 | v_3511;
assign v_13541 = v_3513 | v_3521 | v_3529 | v_3534 | v_3544;
assign v_13542 = v_3545 | v_3546;
assign v_13543 = v_3548 | v_3556 | v_3564 | v_3569 | v_3579;
assign v_13544 = v_3580 | v_3581;
assign v_13545 = v_3583 | v_3591 | v_3599 | v_3604 | v_3614;
assign v_13546 = v_3615 | v_3616;
assign v_13547 = v_3618 | v_3626 | v_3634 | v_3639 | v_3649;
assign v_13548 = v_3650 | v_3651;
assign v_13549 = v_3653 | v_3661 | v_3669 | v_3674 | v_3684;
assign v_13550 = v_3685 | v_3686;
assign v_13551 = v_233 | v_235 | v_238 | v_240 | v_242;
assign v_13552 = v_244 | v_246 | v_248;
assign v_13553 = v_497 | v_499 | v_502 | v_504 | v_506;
assign v_13554 = v_508 | v_510 | v_512;
assign v_13555 = v_3881 | v_3889 | v_3891 | v_3898 | v_3899;
assign v_13556 = v_3907;
assign v_13557 = v_3909 | v_3917 | v_3925 | v_3930 | v_3940;
assign v_13558 = v_3941 | v_3942;
assign v_13559 = v_3944 | v_3952 | v_3960 | v_3965 | v_3975;
assign v_13560 = v_3976 | v_3977;
assign v_13561 = v_3979 | v_3987 | v_3995 | v_4000 | v_4010;
assign v_13562 = v_4011 | v_4012;
assign v_13563 = v_4014 | v_4022 | v_4030 | v_4035 | v_4045;
assign v_13564 = v_4046 | v_4047;
assign v_13565 = v_4049 | v_4057 | v_4065 | v_4070 | v_4080;
assign v_13566 = v_4081 | v_4082;
assign v_13567 = v_4084 | v_4092 | v_4100 | v_4105 | v_4115;
assign v_13568 = v_4116 | v_4117;
assign v_13569 = v_4119 | v_4127 | v_4135 | v_4140 | v_4150;
assign v_13570 = v_4151 | v_4152;
assign v_13571 = v_4154 | v_4162 | v_4170 | v_4175 | v_4185;
assign v_13572 = v_4186 | v_4187;
assign v_13573 = v_4189 | v_4197 | v_4205 | v_4210 | v_4220;
assign v_13574 = v_4221 | v_4222;
assign v_13575 = v_233 | v_235 | v_238 | v_240 | v_242;
assign v_13576 = v_244 | v_246 | v_248;
assign v_13577 = v_497 | v_499 | v_502 | v_504 | v_506;
assign v_13578 = v_508 | v_510 | v_512;
assign v_13579 = v_4417 | v_4425 | v_4427 | v_4434 | v_4435;
assign v_13580 = v_4443;
assign v_13581 = v_4445 | v_4453 | v_4461 | v_4466 | v_4476;
assign v_13582 = v_4477 | v_4478;
assign v_13583 = v_4480 | v_4488 | v_4496 | v_4501 | v_4511;
assign v_13584 = v_4512 | v_4513;
assign v_13585 = v_4515 | v_4523 | v_4531 | v_4536 | v_4546;
assign v_13586 = v_4547 | v_4548;
assign v_13587 = v_4550 | v_4558 | v_4566 | v_4571 | v_4581;
assign v_13588 = v_4582 | v_4583;
assign v_13589 = v_4585 | v_4593 | v_4601 | v_4606 | v_4616;
assign v_13590 = v_4617 | v_4618;
assign v_13591 = v_4620 | v_4628 | v_4636 | v_4641 | v_4651;
assign v_13592 = v_4652 | v_4653;
assign v_13593 = v_4655 | v_4663 | v_4671 | v_4676 | v_4686;
assign v_13594 = v_4687 | v_4688;
assign v_13595 = v_4690 | v_4698 | v_4706 | v_4711 | v_4721;
assign v_13596 = v_4722 | v_4723;
assign v_13597 = v_4725 | v_4733 | v_4741 | v_4746 | v_4756;
assign v_13598 = v_4757 | v_4758;
assign v_13599 = v_233 | v_235 | v_238 | v_240 | v_242;
assign v_13600 = v_244 | v_246 | v_248;
assign v_13601 = v_497 | v_499 | v_502 | v_504 | v_506;
assign v_13602 = v_508 | v_510 | v_512;
assign v_13603 = v_4952 | v_4960 | v_4962 | v_4969 | v_4970;
assign v_13604 = v_4978;
assign v_13605 = v_4980 | v_4988 | v_4996 | v_5001 | v_5011;
assign v_13606 = v_5012 | v_5013;
assign v_13607 = v_5015 | v_5023 | v_5031 | v_5036 | v_5046;
assign v_13608 = v_5047 | v_5048;
assign v_13609 = v_5050 | v_5058 | v_5066 | v_5071 | v_5081;
assign v_13610 = v_5082 | v_5083;
assign v_13611 = v_5085 | v_5093 | v_5101 | v_5106 | v_5116;
assign v_13612 = v_5117 | v_5118;
assign v_13613 = v_5120 | v_5128 | v_5136 | v_5141 | v_5151;
assign v_13614 = v_5152 | v_5153;
assign v_13615 = v_5155 | v_5163 | v_5171 | v_5176 | v_5186;
assign v_13616 = v_5187 | v_5188;
assign v_13617 = v_5190 | v_5198 | v_5206 | v_5211 | v_5221;
assign v_13618 = v_5222 | v_5223;
assign v_13619 = v_5225 | v_5233 | v_5241 | v_5246 | v_5256;
assign v_13620 = v_5257 | v_5258;
assign v_13621 = v_5260 | v_5268 | v_5276 | v_5281 | v_5291;
assign v_13622 = v_5292 | v_5293;
assign v_13623 = v_233 | v_235 | v_238 | v_240 | v_242;
assign v_13624 = v_244 | v_246 | v_248;
assign v_13625 = v_497 | v_499 | v_502 | v_504 | v_506;
assign v_13626 = v_508 | v_510 | v_512;
assign v_13627 = v_5488 | v_5496 | v_5498 | v_5505 | v_5506;
assign v_13628 = v_5514;
assign v_13629 = v_5516 | v_5524 | v_5532 | v_5537 | v_5547;
assign v_13630 = v_5548 | v_5549;
assign v_13631 = v_5551 | v_5559 | v_5567 | v_5572 | v_5582;
assign v_13632 = v_5583 | v_5584;
assign v_13633 = v_5586 | v_5594 | v_5602 | v_5607 | v_5617;
assign v_13634 = v_5618 | v_5619;
assign v_13635 = v_5621 | v_5629 | v_5637 | v_5642 | v_5652;
assign v_13636 = v_5653 | v_5654;
assign v_13637 = v_5656 | v_5664 | v_5672 | v_5677 | v_5687;
assign v_13638 = v_5688 | v_5689;
assign v_13639 = v_5691 | v_5699 | v_5707 | v_5712 | v_5722;
assign v_13640 = v_5723 | v_5724;
assign v_13641 = v_5726 | v_5734 | v_5742 | v_5747 | v_5757;
assign v_13642 = v_5758 | v_5759;
assign v_13643 = v_5761 | v_5769 | v_5777 | v_5782 | v_5792;
assign v_13644 = v_5793 | v_5794;
assign v_13645 = v_5796 | v_5804 | v_5812 | v_5817 | v_5827;
assign v_13646 = v_5828 | v_5829;
assign v_13647 = v_5997 | v_6001 | v_6003 | v_6010 | v_6011;
assign v_13648 = v_6015;
assign v_13649 = v_6017 | v_6025 | v_6033 | v_6038 | v_6048;
assign v_13650 = v_6049 | v_6050;
assign v_13651 = v_6052 | v_6060 | v_6068 | v_6073 | v_6083;
assign v_13652 = v_6084 | v_6085;
assign v_13653 = v_6087 | v_6095 | v_6103 | v_6108 | v_6118;
assign v_13654 = v_6119 | v_6120;
assign v_13655 = v_6122 | v_6130 | v_6138 | v_6143 | v_6153;
assign v_13656 = v_6154 | v_6155;
assign v_13657 = v_6157 | v_6165 | v_6173 | v_6178 | v_6188;
assign v_13658 = v_6189 | v_6190;
assign v_13659 = v_6192 | v_6200 | v_6208 | v_6213 | v_6223;
assign v_13660 = v_6224 | v_6225;
assign v_13661 = v_6227 | v_6235 | v_6243 | v_6248 | v_6258;
assign v_13662 = v_6259 | v_6260;
assign v_13663 = v_6262 | v_6270 | v_6278 | v_6283 | v_6293;
assign v_13664 = v_6294 | v_6295;
assign v_13665 = v_6297 | v_6305 | v_6313 | v_6318 | v_6328;
assign v_13666 = v_6329 | v_6330;
assign v_13667 = v_233 | v_235 | v_238 | v_240 | v_242;
assign v_13668 = v_244 | v_246 | v_248;
assign v_13669 = v_497 | v_499 | v_502 | v_504 | v_506;
assign v_13670 = v_508 | v_510 | v_512;
assign v_13671 = v_6525 | v_6533 | v_6535 | v_6542 | v_6543;
assign v_13672 = v_6551;
assign v_13673 = v_6553 | v_6561 | v_6569 | v_6574 | v_6584;
assign v_13674 = v_6585 | v_6586;
assign v_13675 = v_6588 | v_6596 | v_6604 | v_6609 | v_6619;
assign v_13676 = v_6620 | v_6621;
assign v_13677 = v_6623 | v_6631 | v_6639 | v_6644 | v_6654;
assign v_13678 = v_6655 | v_6656;
assign v_13679 = v_6658 | v_6666 | v_6674 | v_6679 | v_6689;
assign v_13680 = v_6690 | v_6691;
assign v_13681 = v_6693 | v_6701 | v_6709 | v_6714 | v_6724;
assign v_13682 = v_6725 | v_6726;
assign v_13683 = v_6728 | v_6736 | v_6744 | v_6749 | v_6759;
assign v_13684 = v_6760 | v_6761;
assign v_13685 = v_6763 | v_6771 | v_6779 | v_6784 | v_6794;
assign v_13686 = v_6795 | v_6796;
assign v_13687 = v_6798 | v_6806 | v_6814 | v_6819 | v_6829;
assign v_13688 = v_6830 | v_6831;
assign v_13689 = v_6833 | v_6841 | v_6849 | v_6854 | v_6864;
assign v_13690 = v_6865 | v_6866;
assign v_13691 = v_7099 | v_7101 | v_7104 | v_7106 | v_7108;
assign v_13692 = v_7110 | v_7112 | v_7114 | v_7118 | v_7119;
assign v_13693 = v_7125;
assign v_13694 = v_7259 | v_7261 | v_7263 | v_7265 | v_7267;
assign v_13695 = v_7268;
assign v_13696 = v_7213 | v_7215 | v_7217 | v_7224 | v_7273;
assign v_13697 = v_7274;
assign v_13698 = v_7324 | v_7326 | v_7328 | v_7330 | v_7332;
assign v_13699 = v_7333;
assign v_13700 = v_7278 | v_7280 | v_7282 | v_7289 | v_7338;
assign v_13701 = v_7339;
assign v_13702 = v_7363 | v_7365 | v_7368 | v_7370 | v_7372;
assign v_13703 = v_7374 | v_7376 | v_7378 | v_7382 | v_7383;
assign v_13704 = v_7389;
assign v_13705 = ~v_7535 | v_7537 | v_7539 | v_7542 | v_7547;
assign v_13706 = v_7549 | v_7567 | v_7568;
assign v_13707 = ~v_7571 | v_7591 | v_7596 | v_7598 | v_7640;
assign v_13708 = v_7659 | v_7660 | v_7661;
assign v_13709 = v_7682 | v_7684 | v_7705 | v_7707 | v_7728;
assign v_13710 = v_7730 | v_7737 | v_7739 | v_7740 | v_7741;
assign v_13711 = v_7742;
assign v_13712 = v_7763 | v_7765 | v_7786 | v_7788 | v_7809;
assign v_13713 = v_7811 | v_7818 | v_7820 | v_7821 | v_7822;
assign v_13714 = v_7823;
assign v_13715 = v_7844 | v_7846 | v_7867 | v_7869 | v_7890;
assign v_13716 = v_7892 | v_7899 | v_7901 | v_7902 | v_7903;
assign v_13717 = v_7904;
assign v_13718 = v_7925 | v_7927 | v_7948 | v_7950 | v_7971;
assign v_13719 = v_7973 | v_7980 | v_7982 | v_7983 | v_7984;
assign v_13720 = v_7985;
assign v_13721 = v_8006 | v_8008 | v_8029 | v_8031 | v_8052;
assign v_13722 = v_8054 | v_8061 | v_8063 | v_8064 | v_8065;
assign v_13723 = v_8066;
assign v_13724 = v_8087 | v_8089 | v_8110 | v_8112 | v_8133;
assign v_13725 = v_8135 | v_8142 | v_8144 | v_8145 | v_8146;
assign v_13726 = v_8147;
assign v_13727 = v_8168 | v_8170 | v_8191 | v_8193 | v_8214;
assign v_13728 = v_8216 | v_8223 | v_8225 | v_8226 | v_8227;
assign v_13729 = v_8228;
assign v_13730 = v_7099 | v_7101 | v_7104 | v_7106 | v_7108;
assign v_13731 = v_7110 | v_7112 | v_7114;
assign v_13732 = v_7363 | v_7365 | v_7368 | v_7370 | v_7372;
assign v_13733 = v_7374 | v_7376 | v_7378;
assign v_13734 = v_8450 | v_8454 | v_8456 | v_8463 | v_8464;
assign v_13735 = v_8469;
assign v_13736 = v_8471 | v_8480 | v_8489 | v_8495 | v_8506;
assign v_13737 = v_8507 | v_8508;
assign v_13738 = v_8510 | v_8519 | v_8528 | v_8534 | v_8545;
assign v_13739 = v_8546 | v_8547;
assign v_13740 = v_8549 | v_8558 | v_8567 | v_8573 | v_8584;
assign v_13741 = v_8585 | v_8586;
assign v_13742 = v_8588 | v_8597 | v_8606 | v_8612 | v_8623;
assign v_13743 = v_8624 | v_8625;
assign v_13744 = v_8627 | v_8636 | v_8645 | v_8651 | v_8662;
assign v_13745 = v_8663 | v_8664;
assign v_13746 = v_8666 | v_8675 | v_8684 | v_8690 | v_8701;
assign v_13747 = v_8702 | v_8703;
assign v_13748 = v_8705 | v_8714 | v_8723 | v_8729 | v_8740;
assign v_13749 = v_8741 | v_8742;
assign v_13750 = v_8911 | v_8915 | v_8917 | v_8924 | v_8925;
assign v_13751 = v_8929;
assign v_13752 = v_8931 | v_8939 | v_8947 | v_8952 | v_8962;
assign v_13753 = v_8963 | v_8964;
assign v_13754 = v_8966 | v_8974 | v_8982 | v_8987 | v_8997;
assign v_13755 = v_8998 | v_8999;
assign v_13756 = v_9001 | v_9009 | v_9017 | v_9022 | v_9032;
assign v_13757 = v_9033 | v_9034;
assign v_13758 = v_9036 | v_9044 | v_9052 | v_9057 | v_9067;
assign v_13759 = v_9068 | v_9069;
assign v_13760 = v_9071 | v_9079 | v_9087 | v_9092 | v_9102;
assign v_13761 = v_9103 | v_9104;
assign v_13762 = v_9106 | v_9114 | v_9122 | v_9127 | v_9137;
assign v_13763 = v_9138 | v_9139;
assign v_13764 = v_9141 | v_9149 | v_9157 | v_9162 | v_9172;
assign v_13765 = v_9173 | v_9174;
assign v_13766 = v_7099 | v_7101 | v_7104 | v_7106 | v_7108;
assign v_13767 = v_7110 | v_7112 | v_7114;
assign v_13768 = v_7363 | v_7365 | v_7368 | v_7370 | v_7372;
assign v_13769 = v_7374 | v_7376 | v_7378;
assign v_13770 = v_9368 | v_9376 | v_9378 | v_9385 | v_9386;
assign v_13771 = v_9394;
assign v_13772 = v_9396 | v_9404 | v_9412 | v_9417 | v_9427;
assign v_13773 = v_9428 | v_9429;
assign v_13774 = v_9431 | v_9439 | v_9447 | v_9452 | v_9462;
assign v_13775 = v_9463 | v_9464;
assign v_13776 = v_9466 | v_9474 | v_9482 | v_9487 | v_9497;
assign v_13777 = v_9498 | v_9499;
assign v_13778 = v_9501 | v_9509 | v_9517 | v_9522 | v_9532;
assign v_13779 = v_9533 | v_9534;
assign v_13780 = v_9536 | v_9544 | v_9552 | v_9557 | v_9567;
assign v_13781 = v_9568 | v_9569;
assign v_13782 = v_9571 | v_9579 | v_9587 | v_9592 | v_9602;
assign v_13783 = v_9603 | v_9604;
assign v_13784 = v_9606 | v_9614 | v_9622 | v_9627 | v_9637;
assign v_13785 = v_9638 | v_9639;
assign v_13786 = v_7099 | v_7101 | v_7104 | v_7106 | v_7108;
assign v_13787 = v_7110 | v_7112 | v_7114;
assign v_13788 = v_7363 | v_7365 | v_7368 | v_7370 | v_7372;
assign v_13789 = v_7374 | v_7376 | v_7378;
assign v_13790 = v_9831 | v_9839 | v_9841 | v_9848 | v_9849;
assign v_13791 = v_9857;
assign v_13792 = v_9859 | v_9867 | v_9875 | v_9880 | v_9890;
assign v_13793 = v_9891 | v_9892;
assign v_13794 = v_9894 | v_9902 | v_9910 | v_9915 | v_9925;
assign v_13795 = v_9926 | v_9927;
assign v_13796 = v_9929 | v_9937 | v_9945 | v_9950 | v_9960;
assign v_13797 = v_9961 | v_9962;
assign v_13798 = v_9964 | v_9972 | v_9980 | v_9985 | v_9995;
assign v_13799 = v_9996 | v_9997;
assign v_13800 = v_9999 | v_10007 | v_10015 | v_10020 | v_10030;
assign v_13801 = v_10031 | v_10032;
assign v_13802 = v_10034 | v_10042 | v_10050 | v_10055 | v_10065;
assign v_13803 = v_10066 | v_10067;
assign v_13804 = v_10069 | v_10077 | v_10085 | v_10090 | v_10100;
assign v_13805 = v_10101 | v_10102;
assign v_13806 = v_7099 | v_7101 | v_7104 | v_7106 | v_7108;
assign v_13807 = v_7110 | v_7112 | v_7114;
assign v_13808 = v_7363 | v_7365 | v_7368 | v_7370 | v_7372;
assign v_13809 = v_7374 | v_7376 | v_7378;
assign v_13810 = v_10297 | v_10305 | v_10307 | v_10314 | v_10315;
assign v_13811 = v_10323;
assign v_13812 = v_10325 | v_10333 | v_10341 | v_10346 | v_10356;
assign v_13813 = v_10357 | v_10358;
assign v_13814 = v_10360 | v_10368 | v_10376 | v_10381 | v_10391;
assign v_13815 = v_10392 | v_10393;
assign v_13816 = v_10395 | v_10403 | v_10411 | v_10416 | v_10426;
assign v_13817 = v_10427 | v_10428;
assign v_13818 = v_10430 | v_10438 | v_10446 | v_10451 | v_10461;
assign v_13819 = v_10462 | v_10463;
assign v_13820 = v_10465 | v_10473 | v_10481 | v_10486 | v_10496;
assign v_13821 = v_10497 | v_10498;
assign v_13822 = v_10500 | v_10508 | v_10516 | v_10521 | v_10531;
assign v_13823 = v_10532 | v_10533;
assign v_13824 = v_10535 | v_10543 | v_10551 | v_10556 | v_10566;
assign v_13825 = v_10567 | v_10568;
assign v_13826 = v_7099 | v_7101 | v_7104 | v_7106 | v_7108;
assign v_13827 = v_7110 | v_7112 | v_7114;
assign v_13828 = v_7363 | v_7365 | v_7368 | v_7370 | v_7372;
assign v_13829 = v_7374 | v_7376 | v_7378;
assign v_13830 = v_10763 | v_10771 | v_10773 | v_10780 | v_10781;
assign v_13831 = v_10789;
assign v_13832 = v_10791 | v_10799 | v_10807 | v_10812 | v_10822;
assign v_13833 = v_10823 | v_10824;
assign v_13834 = v_10826 | v_10834 | v_10842 | v_10847 | v_10857;
assign v_13835 = v_10858 | v_10859;
assign v_13836 = v_10861 | v_10869 | v_10877 | v_10882 | v_10892;
assign v_13837 = v_10893 | v_10894;
assign v_13838 = v_10896 | v_10904 | v_10912 | v_10917 | v_10927;
assign v_13839 = v_10928 | v_10929;
assign v_13840 = v_10931 | v_10939 | v_10947 | v_10952 | v_10962;
assign v_13841 = v_10963 | v_10964;
assign v_13842 = v_10966 | v_10974 | v_10982 | v_10987 | v_10997;
assign v_13843 = v_10998 | v_10999;
assign v_13844 = v_11001 | v_11009 | v_11017 | v_11022 | v_11032;
assign v_13845 = v_11033 | v_11034;
assign v_13846 = v_7099 | v_7101 | v_7104 | v_7106 | v_7108;
assign v_13847 = v_7110 | v_7112 | v_7114;
assign v_13848 = v_7363 | v_7365 | v_7368 | v_7370 | v_7372;
assign v_13849 = v_7374 | v_7376 | v_7378;
assign v_13850 = v_11228 | v_11236 | v_11238 | v_11245 | v_11246;
assign v_13851 = v_11254;
assign v_13852 = v_11256 | v_11264 | v_11272 | v_11277 | v_11287;
assign v_13853 = v_11288 | v_11289;
assign v_13854 = v_11291 | v_11299 | v_11307 | v_11312 | v_11322;
assign v_13855 = v_11323 | v_11324;
assign v_13856 = v_11326 | v_11334 | v_11342 | v_11347 | v_11357;
assign v_13857 = v_11358 | v_11359;
assign v_13858 = v_11361 | v_11369 | v_11377 | v_11382 | v_11392;
assign v_13859 = v_11393 | v_11394;
assign v_13860 = v_11396 | v_11404 | v_11412 | v_11417 | v_11427;
assign v_13861 = v_11428 | v_11429;
assign v_13862 = v_11431 | v_11439 | v_11447 | v_11452 | v_11462;
assign v_13863 = v_11463 | v_11464;
assign v_13864 = v_11466 | v_11474 | v_11482 | v_11487 | v_11497;
assign v_13865 = v_11498 | v_11499;
assign v_13866 = v_7099 | v_7101 | v_7104 | v_7106 | v_7108;
assign v_13867 = v_7110 | v_7112 | v_7114;
assign v_13868 = v_7363 | v_7365 | v_7368 | v_7370 | v_7372;
assign v_13869 = v_7374 | v_7376 | v_7378;
assign v_13870 = v_11694 | v_11702 | v_11704 | v_11711 | v_11712;
assign v_13871 = v_11720;
assign v_13872 = v_11722 | v_11730 | v_11738 | v_11743 | v_11753;
assign v_13873 = v_11754 | v_11755;
assign v_13874 = v_11757 | v_11765 | v_11773 | v_11778 | v_11788;
assign v_13875 = v_11789 | v_11790;
assign v_13876 = v_11792 | v_11800 | v_11808 | v_11813 | v_11823;
assign v_13877 = v_11824 | v_11825;
assign v_13878 = v_11827 | v_11835 | v_11843 | v_11848 | v_11858;
assign v_13879 = v_11859 | v_11860;
assign v_13880 = v_11862 | v_11870 | v_11878 | v_11883 | v_11893;
assign v_13881 = v_11894 | v_11895;
assign v_13882 = v_11897 | v_11905 | v_11913 | v_11918 | v_11928;
assign v_13883 = v_11929 | v_11930;
assign v_13884 = v_11932 | v_11940 | v_11948 | v_11953 | v_11963;
assign v_13885 = v_11964 | v_11965;
assign v_13886 = v_12133 | v_12137 | v_12139 | v_12146 | v_12147;
assign v_13887 = v_12151;
assign v_13888 = v_12153 | v_12161 | v_12169 | v_12174 | v_12184;
assign v_13889 = v_12185 | v_12186;
assign v_13890 = v_12188 | v_12196 | v_12204 | v_12209 | v_12219;
assign v_13891 = v_12220 | v_12221;
assign v_13892 = v_12223 | v_12231 | v_12239 | v_12244 | v_12254;
assign v_13893 = v_12255 | v_12256;
assign v_13894 = v_12258 | v_12266 | v_12274 | v_12279 | v_12289;
assign v_13895 = v_12290 | v_12291;
assign v_13896 = v_12293 | v_12301 | v_12309 | v_12314 | v_12324;
assign v_13897 = v_12325 | v_12326;
assign v_13898 = v_12328 | v_12336 | v_12344 | v_12349 | v_12359;
assign v_13899 = v_12360 | v_12361;
assign v_13900 = v_12363 | v_12371 | v_12379 | v_12384 | v_12394;
assign v_13901 = v_12395 | v_12396;
assign v_13902 = v_7099 | v_7101 | v_7104 | v_7106 | v_7108;
assign v_13903 = v_7110 | v_7112 | v_7114;
assign v_13904 = v_7363 | v_7365 | v_7368 | v_7370 | v_7372;
assign v_13905 = v_7374 | v_7376 | v_7378;
assign v_13906 = v_12591 | v_12599 | v_12601 | v_12608 | v_12609;
assign v_13907 = v_12617;
assign v_13908 = v_12619 | v_12627 | v_12635 | v_12640 | v_12650;
assign v_13909 = v_12651 | v_12652;
assign v_13910 = v_12654 | v_12662 | v_12670 | v_12675 | v_12685;
assign v_13911 = v_12686 | v_12687;
assign v_13912 = v_12689 | v_12697 | v_12705 | v_12710 | v_12720;
assign v_13913 = v_12721 | v_12722;
assign v_13914 = v_12724 | v_12732 | v_12740 | v_12745 | v_12755;
assign v_13915 = v_12756 | v_12757;
assign v_13916 = v_12759 | v_12767 | v_12775 | v_12780 | v_12790;
assign v_13917 = v_12791 | v_12792;
assign v_13918 = v_12794 | v_12802 | v_12810 | v_12815 | v_12825;
assign v_13919 = v_12826 | v_12827;
assign v_13920 = v_12829 | v_12837 | v_12845 | v_12850 | v_12860;
assign v_13921 = v_12861 | v_12862;
assign v_12864 = ~v_8743 ^ ~v_2117;
assign v_12865 = ~v_9175 ^ ~v_2619;
assign v_12866 = ~v_9640 ^ ~v_3154;
assign v_12867 = ~v_10103 ^ ~v_3687;
assign v_12868 = ~v_10569 ^ ~v_4223;
assign v_12869 = ~v_11035 ^ ~v_4759;
assign v_12870 = ~v_11500 ^ ~v_5294;
assign v_12871 = ~v_11966 ^ ~v_5830;
assign v_12872 = ~v_12397 ^ ~v_6331;
assign v_12873 = ~v_12863 ^ ~v_6867;
assign x_1 = ~v_1526 | v_12874;
assign o_1 = x_1;
endmodule
