// Verilog file written by procedure writeCombinationalCircuitInVerilog
//Skolem functions to be generated for i_ variables
module neclaftp2002_all_bit_differing_from_cycle ( i_1, i_2, i_3, i_4, i_5, i_6, i_7, i_8, i_9, i_10, i_11, i_12, i_13, i_14, i_15, i_16, i_17, i_18, i_19, i_20, i_21, i_22, i_23, i_24, i_25, i_26, i_27, i_28, i_29, i_30, i_31, i_32, x_33, x_34, x_35, x_36, x_37, x_38, x_39, x_40, x_41, x_42, x_43, x_44, x_45, x_46, x_47, x_48, x_49, x_50, x_51, x_52, x_53, x_54, x_55, x_56, x_57, x_58, x_59, x_60, x_61, x_62, x_63, x_64, x_65, x_66, x_67, x_68, x_69, x_70, x_71, x_72, x_73, x_74, x_75, x_76, x_77, x_78, x_79, x_80, x_81, x_82, x_83, x_84, x_85, x_86, x_87, x_88, x_89, x_90, x_91, x_92, x_93, x_94, x_95, x_96, x_97, x_98, x_99, x_100, x_101, x_102, x_103, x_104, x_105, x_106, x_107, x_108, x_109, x_110, x_111, x_112, x_113, x_114, x_115, x_116, x_117, x_118, x_119, x_120, x_121, x_122, x_123, x_124, x_125, x_126, x_127, x_128, x_129, x_130, x_131, x_132, x_133, x_134, x_135, x_136, x_137, x_138, x_139, x_140, x_141, x_142, x_143, x_144, x_145, x_146, x_147, x_148, x_149, x_150, x_151, x_152, x_153, x_154, x_155, x_156, x_157, x_158, x_159, x_160, x_161, x_162, x_163, x_164, x_165, x_166, x_167, x_168, x_169, x_170, x_171, x_172, x_173, x_174, x_175, x_176, x_177, x_178, x_179, x_180, x_181, x_182, x_183, x_184, x_185, x_186, x_187, x_188, x_189, x_190, x_191, x_192, x_193, x_194, x_195, x_196, x_197, x_198, x_199, x_200, x_201, x_202, x_203, x_204, x_205, x_206, x_207, x_208, x_209, x_210, x_211, x_212, x_213, x_214, x_215, x_216, x_217, x_218, x_219, x_220, x_221, x_222, x_223, x_224, x_225, x_226, x_227, x_228, x_229, x_230, x_231, x_232, x_233, x_234, x_235, x_236, x_237, x_238, x_239, x_240, x_241, x_242, x_243, x_244, x_245, x_246, x_247, x_248, x_249, x_250, x_251, x_252, x_253, x_254, x_255, x_256, x_257, x_258, x_259, x_260, x_261, x_262, x_263, x_264, x_265, x_266, x_267, x_268, x_269, x_270, x_271, x_272, x_273, x_274, x_275, x_276, x_277, x_278, x_279, x_280, x_281, x_282, x_283, x_284, x_285, x_286, x_287, x_288, x_289, x_290, x_291, x_292, x_293, x_294, x_295, x_296, x_297, x_298, x_299, x_300, x_301, x_302, x_303, x_304, x_305, x_306, x_307, x_308, x_309, x_310, x_311, x_312, x_313, x_314, x_315, x_316, x_317, x_318, x_319, x_320, x_321, x_322, x_323, x_324, x_325, x_326, x_327, x_328, x_329, x_330, x_331, x_332, x_333, x_334, x_335, x_336, x_337, x_338, x_339, x_340, x_341, x_342, x_343, x_344, x_345, x_346, x_347, x_348, x_349, x_350, x_351, x_352, x_353, x_354, x_355, x_356, x_357, x_358, x_359, x_360, x_361, x_362, x_363, x_364, x_365, x_366, x_367, x_368, x_369, x_370, x_371, x_372, x_373, x_374, x_375, x_376, x_377, x_378, x_379, x_380, x_381, x_382, x_383, x_384, x_385, x_386, x_387, x_388, x_389, x_390, x_391, x_392, x_393, x_394, x_395, x_396, x_397, x_398, x_399, x_400, x_401, x_402, x_403, x_404, x_405, x_406, x_407, x_408, x_409, x_410, x_411, x_412, x_413, x_414, x_415, x_416, x_417, x_418, x_419, x_420, x_421, x_422, x_423, x_424, x_425, x_426, x_427, x_428, x_429, x_430, x_431, x_432, x_433, x_434, x_435, x_436, x_437, x_438, x_439, x_440, x_441, x_442, x_443, x_444, x_445, x_446, x_447, x_448, x_449, x_450, x_451, x_452, x_453, x_454, x_455, x_456, x_457, x_458, x_459, x_460, x_461, x_462, x_463, x_464, x_465, x_466, x_467, x_468, x_469, x_470, x_471, x_472, x_473, x_474, x_475, x_476, x_477, x_478, x_479, x_480, x_481, x_482, x_483, x_484, x_485, x_486, x_487, x_488, x_489, x_490, x_491, x_492, x_493, x_494, x_495, x_496, x_497, x_498, x_499, x_500, x_501, x_502, x_503, x_504, x_505, x_506, x_507, x_508, x_509, x_510, x_511, x_512, x_513, x_514, x_515, x_516, x_517, x_518, x_519, x_520, x_521, x_522, x_523, x_524, x_525, x_526, x_527, x_528, x_529, x_530, x_531, x_532, x_533, x_534, x_535, x_536, x_537, x_538, x_539, x_540, x_541, x_542, x_543, x_544, x_545, x_546, x_547, x_548, x_549, x_550, x_551, x_552, x_553, x_554, x_555, x_556, x_557, x_558, x_559, x_560, x_561, x_562, x_563, x_564, x_565, x_566, x_567, x_568, x_569, x_570, x_571, x_572, x_573, x_574, x_575, x_576, x_577, x_578, x_579, x_580, x_581, x_582, x_583, x_584, x_585, x_586, x_587, x_588, x_589, x_590, x_591, x_592, x_593, x_594, x_595, x_596, x_597, x_598, x_599, x_600, x_601, x_602, x_603, x_604, x_605, x_606, x_607, x_608, x_609, x_610, x_611, x_612, x_613, x_614, x_615, x_616, x_617, x_618, x_619, x_620, x_621, x_622, x_623, x_624, x_625, x_626, x_627, x_628, x_629, x_630, x_631, x_632, x_633, x_634, x_635, x_636, x_637, x_638, x_639, x_640, x_641, x_642, x_643, x_644, x_645, x_646, x_647, x_648, x_649, x_650, x_651, x_652, x_653, x_654, x_655, x_656, x_657, x_658, x_659, x_660, x_661, x_662, x_663, x_664, x_665, x_666, x_667, x_668, x_669, x_670, x_671, x_672, x_673, x_674, x_675, x_676, x_677, x_678, x_679, x_680, x_681, x_682, x_683, x_684, x_685, x_686, x_687, x_688, x_689, x_690, x_691, x_692, x_693, x_694, x_695, x_696, x_697, x_698, x_699, x_700, x_701, x_702, x_703, x_704, x_705, x_706, x_707, x_708, x_709, x_710, x_711, x_712, x_713, x_714, x_715, x_716, x_717, x_718, x_719, x_720, x_721, x_722, x_723, x_724, x_725, x_726, x_727, x_728, x_729, x_730, x_731, x_732, x_733, x_734, x_735, x_736, x_737, x_738, x_739, x_740, x_741, x_742, x_743, x_744, x_745, x_746, x_747, x_748, x_749, x_750, x_751, x_752, x_753, x_754, x_755, x_756, x_757, x_758, x_759, x_760, x_761, x_762, x_763, x_764, x_765, x_766, x_767, x_768, x_769, x_770, x_771, x_772, x_773, x_774, x_775, x_776, x_777, x_778, x_779, x_780, x_781, x_782, x_783, x_784, x_785, x_786, x_787, x_788, x_789, x_790, x_791, x_792, x_793, x_794, x_795, x_796, x_797, x_798, x_799, x_800, x_801, x_802, x_803, x_804, x_805, x_806, x_807, x_808, x_809, x_810, x_811, x_812, x_813, x_814, x_815, x_816, x_817, x_818, x_819, x_820, x_821, x_822, x_823, x_824, x_825, x_826, x_827, x_828, x_829, x_830, x_831, x_832, x_833, x_834, x_835, x_836, x_837, x_838, x_839, x_840, x_841, x_842, x_843, x_844, x_845, x_846, x_847, x_848, x_849, x_850, x_851, x_852, x_853, x_854, x_855, x_856, x_857, x_858, x_859, x_860, x_861, x_862, x_863, x_864, x_865, x_866, x_867, x_868, x_869, x_870, x_871, x_872, x_873, x_874, x_875, x_876, x_877, x_878, x_879, x_880, x_881, x_882, x_883, x_884, x_885, x_886, x_887, x_888, x_889, x_890, x_891, x_892, x_893, x_894, x_895, x_896, x_897, x_898, x_899, x_900, x_901, x_902, x_903, x_904, x_905, x_906, x_907, x_908, x_909, x_910, x_911, x_912, x_913, x_914, x_915, x_916, x_917, x_918, x_919, x_920, x_921, x_922, x_923, x_924, x_925, x_926, x_927, x_928, x_929, x_930, x_931, x_932, x_933, x_934, x_935, x_936, x_937, x_938, x_939, x_940, x_941, x_942, x_943, x_944, x_945, x_946, x_947, x_948, x_949, x_950, x_951, x_952, x_953, x_954, x_955, x_956, x_957, x_958, x_959, x_960, x_961, x_962, x_963, x_964, x_965, x_966, x_967, x_968, x_969, x_970, x_971, x_972, x_973, x_974, x_975, x_976, x_977, x_978, x_979, x_980, x_981, x_982, x_983, x_984, x_985, x_986, x_987, x_988, x_989, x_990, x_991, x_992, x_993, x_994, x_995, x_996, x_997, x_998, x_999, x_1000, x_1001, x_1002, x_1003, x_1004, x_1005, x_1006, x_1007, x_1008, x_1009, x_1010, x_1011, x_1012, x_1013, x_1014, x_1015, x_1016, x_1017, x_1018, x_1019, x_1020, x_1021, x_1022, x_1023, x_1024, x_1025, x_1026, x_1027, x_1028, x_1029, x_1030, x_1031, x_1032, x_1033, x_1034, x_1035, x_1036, x_1037, x_1038, x_1039, x_1040, x_1041, x_1042, x_1043, x_1044, x_1045, x_1046, x_1047, x_1048, x_1049, x_1050, x_1051, x_1052, x_1053, x_1054, x_1055, x_1056, x_1057, x_1058, x_1059, x_1060, x_1061, x_1062, x_1063, x_1064, x_1065, x_1066, x_1067, x_1068, x_1069, x_1070, x_1071, x_1072, x_1073, x_1074, x_1075, x_1076, x_1077, x_1078, x_1079, x_1080, x_1081, x_1082, x_1083, x_1084, x_1085, x_1086, x_1087, x_1088, x_1089, x_1090, x_1091, x_1092, x_1093, x_1094, x_1095, x_1096, x_1097, x_1098, x_1099, x_1100, x_1101, x_1102, x_1103, x_1104, x_1105, x_1106, x_1107, x_1108, x_1109, x_1110, x_1111, x_1112, x_1113, x_1114, x_1115, x_1116, x_1117, x_1118, x_1119, x_1120, x_1121, x_1122, x_1123, x_1124, x_1125, x_1126, x_1127, x_1128, x_1129, x_1130, x_1131, x_1132, x_1133, x_1134, x_1135, x_1136, x_1137, x_1138, x_1139, x_1140, x_1141, x_1142, x_1143, x_1144, x_1145, x_1146, x_1147, x_1148, x_1149, x_1150, x_1151, x_1152, x_1153, x_1154, x_1155, x_1156, x_1157, x_1158, x_1159, x_1160, x_1161, x_1162, x_1163, x_1164, x_1165, x_1166, x_1167, x_1168, x_1169, x_1170, x_1171, x_1172, x_1173, x_1174, x_1175, x_1176, x_1177, x_1178, x_1179, x_1180, x_1181, x_1182, x_1183, x_1184, x_1185, x_1186, x_1187, x_1188, x_1189, x_1190, x_1191, x_1192, x_1193, x_1194, x_1195, x_1196, x_1197, x_1198, x_1199, x_1200, x_1201, x_1202, x_1203, x_1204, x_1205, x_1206, x_1207, x_1208, x_1209, x_1210, x_1211, x_1212, x_1213, x_1214, x_1215, x_1216, x_1217, x_1218, x_1219, x_1220, x_1221, x_1222, x_1223, x_1224, x_1225, x_1226, x_1227, x_1228, x_1229, x_1230, x_1231, x_1232, x_1233, x_1234, x_1235, x_1236, x_1237, x_1238, x_1239, x_1240, x_1241, x_1242, x_1243, x_1244, x_1245, x_1246, x_1247, x_1248, x_1249, x_1250, x_1251, x_1252, x_1253, x_1254, x_1255, x_1256, x_1257, x_1258, x_1259, x_1260, x_1261, x_1262, x_1263, x_1264, x_1265, x_1266, x_1267, x_1268, x_1269, x_1270, x_1271, x_1272, x_1273, x_1274, x_1275, x_1276, x_1277, x_1278, x_1279, x_1280, x_1281, x_1282, x_1283, x_1284, x_1285, x_1286, x_1287, x_1288, x_1289, x_1290, x_1291, x_1292, x_1293, x_1294, x_1295, x_1296, x_1297, x_1298, x_1299, x_1300, x_1301, x_1302, x_1303, x_1304, x_1305, x_1306, x_1307, x_1308, x_1309, x_1310, x_1311, x_1312, x_1313, x_1314, x_1315, x_1316, x_1317, x_1318, x_1319, x_1320, x_1321, x_1322, x_1323, x_1324, x_1325, x_1326, x_1327, x_1328, x_1329, x_1330, x_1331, x_1332, x_1333, x_1334, x_1335, x_1336, x_1337, x_1338, x_1339, x_1340, x_1341, x_1342, x_1343, x_1344, x_1345, x_1346, x_1347, x_1348, x_1349, x_1350, x_1351, x_1352, x_1353, x_1354, x_1355, x_1356, x_1357, x_1358, x_1359, x_1360, x_1361, x_1362, x_1363, x_1364, x_1365, x_1366, x_1367, x_1368, x_1369, x_1370, x_1371, x_1372, x_1373, x_1374, x_1375, x_1376, x_1377, x_1378, x_1379, x_1380, x_1381, x_1382, x_1383, x_1384, x_1385, x_1386, x_1387, x_1388, x_1389, x_1390, x_1391, x_1392, x_1393, x_1394, x_1395, x_1396, x_1397, x_1398, x_1399, x_1400, x_1401, x_1402, x_1403, x_1404, x_1405, x_1406, x_1407, x_1408, x_1409, x_1410, x_1411, x_1412, x_1413, x_1414, x_1415, x_1416, x_1417, x_1418, x_1419, x_1420, x_1421, x_1422, x_1423, x_1424, x_1425, x_1426, x_1427, x_1428, x_1429, x_1430, x_1431, x_1432, x_1433, x_1434, x_1435, x_1436, x_1437, x_1438, x_1439, x_1440, x_1441, x_1442, x_1443, x_1444, x_1445, x_1446, x_1447, x_1448, x_1449, x_1450, x_1451, x_1452, x_1453, x_1454, x_1455, x_1456, x_1457, x_1458, x_1459, x_1460, x_1461, x_1462, x_1463, x_1464, x_1465, x_1466, x_1467, x_1468, x_1469, x_1470, x_1471, x_1472, x_1473, x_1474, x_1475, x_1476, x_1477, x_1478, x_1479, x_1480, x_1481, x_1482, x_1483, x_1484, x_1485, x_1486, x_1487, x_1488, x_1489, x_1490, x_1491, x_1492, x_1493, x_1494, x_1495, x_1496, x_1497, x_1498, x_1499, x_1500, x_1501, x_1502, x_1503, x_1504, x_1505, x_1506, x_1507, x_1508, x_1509, x_1510, x_1511, x_1512, x_1513, x_1514, x_1515, x_1516, x_1517, x_1518, x_1519, x_1520, x_1521, x_1522, x_1523, x_1524, x_1525, x_1526, x_1527, x_1528, x_1529, x_1530, x_1531, x_1532, x_1533, x_1534, x_1535, x_1536, x_1537, x_1538, x_1539, x_1540, x_1541, x_1542, x_1543, x_1544, x_1545, x_1546, x_1547, x_1548, x_1549, x_1550, x_1551, x_1552, x_1553, x_1554, x_1555, x_1556, x_1557, x_1558, x_1559, x_1560, x_1561, x_1562, x_1563, x_1564, x_1565, x_1566, x_1567, x_1568, x_1569, x_1570, x_1571, x_1572, x_1573, x_1574, x_1575, x_1576, x_1577, x_1578, x_1579, x_1580, x_1581, x_1582, x_1583, x_1584, x_1585, x_1586, x_1587, x_1588, x_1589, x_1590, x_1591, x_1592, x_1593, x_1594, x_1595, x_1596, x_1597, x_1598, x_1599, x_1600, x_1601, x_1602, x_1603, x_1604, x_1605, x_1606, x_1607, x_1608, x_1609, x_1610, x_1611, x_1612, x_1613, x_1614, x_1615, x_1616, x_1617, x_1618, x_1619, x_1620, x_1621, x_1622, x_1623, x_1624, x_1625, x_1626, x_1627, x_1628, x_1629, x_1630, x_1631, x_1632, x_1633, x_1634, x_1635, x_1636, x_1637, x_1638, x_1639, x_1640, x_1641, x_1642, x_1643, x_1644, x_1645, x_1646, x_1647, x_1648, x_1649, x_1650, x_1651, x_1652, x_1653, x_1654, x_1655, x_1656, x_1657, x_1658, x_1659, x_1660, x_1661, x_1662, x_1663, x_1664, x_1665, x_1666, x_1667, x_1668, x_1669, x_1670, x_1671, x_1672, x_1673, x_1674, x_1675, x_1676, x_1677, x_1678, x_1679, x_1680, x_1681, x_1682, x_1683, x_1684, x_1685, x_1686, x_1687, x_1688, x_1689, x_1690, x_1691, x_1692, x_1693, x_1694, x_1695, x_1696, x_1697, x_1698, x_1699, x_1700, x_1701, x_1702, x_1703, x_1704, x_1705, x_1706, x_1707, x_1708, x_1709, x_1710, x_1711, x_1712, x_1713, x_1714, x_1715, x_1716, x_1717, x_1718, x_1719, x_1720, x_1721, x_1722, x_1723, x_1724, x_1725, x_1726, x_1727, x_1728, x_1729, x_1730, x_1731, x_1732, x_1733, x_1734, x_1735, x_1736, x_1737, x_1738, x_1739, x_1740, x_1741, x_1742, x_1743, x_1744, x_1745, x_1746, x_1747, x_1748, x_1749, x_1750, x_1751, x_1752, x_1753, x_1754, x_1755, x_1756, x_1757, x_1758, x_1759, x_1760, x_1761, x_1762, x_1763, x_1764, x_1765, x_1766, x_1767, x_1768, x_1769, x_1770, x_1771, x_1772, x_1773, x_1774, x_1775, x_1776, x_1777, x_1778, x_1779, x_1780, x_1781, x_1782, x_1783, x_1784, x_1785, x_1786, x_1787, x_1788, x_1789, x_1790, x_1791, x_1792, x_1793, x_1794, x_1795, x_1796, x_1797, x_1798, x_1799, x_1800, x_1801, x_1802, x_1803, x_1804, x_1805, x_1806, x_1807, x_1808, x_1809, x_1810, x_1811, x_1812, x_1813, x_1814, x_1815, x_1816, x_1817, x_1818, x_1819, x_1820, x_1821, x_1822, x_1823, x_1824, x_1825, x_1826, x_1827, x_1828, x_1829, x_1830, x_1831, x_1832, x_1833, x_1834, x_1835, x_1836, x_1837, x_1838, x_1839, x_1840, x_1841, x_1842, x_1843, x_1844, x_1845, x_1846, x_1847, x_1848, x_1849, x_1850, x_1851, x_1852, x_1853, x_1854, x_1855, x_1856, x_1857, x_1858, x_1859, x_1860, x_1861, x_1862, x_1863, x_1864, x_1865, x_1866, x_1867, x_1868, x_1869, x_1870, x_1871, x_1872, x_1873, x_1874, x_1875, x_1876, x_1877, x_1878, x_1879, x_1880, x_1881, x_1882, x_1883, x_1884, x_1885, x_1886, x_1887, x_1888, x_1889, x_1890, x_1891, x_1892, x_1893, x_1894, x_1895, x_1896, x_1897, x_1898, x_1899, x_1900, x_1901, x_1902, x_1903, x_1904, x_1905, x_1906, x_1907, x_1908, x_1909, x_1910, x_1911, x_1912, x_1913, x_1914, x_1915, x_1916, x_1917, x_1918, x_1919, x_1920, x_1921, x_1922, x_1923, x_1924, x_1925, x_1926, x_1927, x_1928, x_1929, x_1930, x_1931, x_1932, x_1933, x_1934, x_1935, x_1936, x_1937, x_1938, x_1939, x_1940, x_1941, x_1942, x_1943, x_1944, x_1945, x_1946, x_1947, x_1948, x_1949, x_1950, x_1951, x_1952, x_1953, x_1954, x_1955, x_1956, x_1957, x_1958, x_1959, x_1960, x_1961, x_1962, x_1963, x_1964, x_1965, x_1966, x_1967, x_1968, x_1969, x_1970, x_1971, x_1972, x_1973, x_1974, x_1975, x_1976, x_1977, x_1978, x_1979, x_1980, x_1981, x_1982, x_1983, x_1984, x_1985, x_1986, x_1987, x_1988, x_1989, x_1990, x_1991, x_1992, x_1993, x_1994, x_1995, x_1996, x_1997, x_1998, x_1999, x_2000, x_2001, x_2002, x_2003, x_2004, x_2005, x_2006, x_2007, x_2008, x_2009, x_2010, x_2011, x_2012, x_2013, x_2014, x_2015, x_2016, x_2017, x_2018, x_2019, x_2020, x_2021, x_2022, x_2023, x_2024, x_2025, x_2026, x_2027, x_2028, x_2029, x_2030, x_2031, x_2032, x_2033, x_2034, x_2035, x_2036, x_2037, x_2038, x_2039, x_2040, x_2041, x_2042, x_2043, x_2044, x_2045, x_2046, x_2047, x_2048, x_2049, x_2050, x_2051, x_2052, x_2053, x_2054, x_2055, x_2056, x_2057, x_2058, x_2059, x_2060, x_2061, x_2062, x_2063, x_2064, x_2065, x_2066, x_2067, x_2068, x_2069, x_2070, x_2071, x_2072, x_2073, x_2074, x_2075, x_2076, x_2077, x_2078, x_2079, x_2080, x_2081, x_2082, x_2083, x_2084, x_2085, x_2086, x_2087, x_2088, x_2089, x_2090, x_2091, x_2092, x_2093, x_2094, x_2095, x_2096, x_2097, x_2098, x_2099, x_2100, x_2101, x_2102, x_2103, x_2104, x_2105, x_2106, x_2107, x_2108, x_2109, x_2110, x_2111, x_2112, x_2113, x_2114, x_2115, x_2116, x_2117, x_2118, x_2119, x_2120, x_2121, x_2122, x_2123, x_2124, x_2125, x_2126, x_2127, x_2128, x_2129, x_2130, x_2131, x_2132, x_2133, x_2134, x_2135, x_2136, x_2137, x_2138, x_2139, x_2140, x_2141, x_2142, x_2143, x_2144, x_2145, x_2146, x_2147, x_2148, x_2149, x_2150, x_2151, x_2152, x_2153, x_2154, x_2155, x_2156, x_2157, x_2158, x_2159, x_2160, x_2161, x_2162, x_2163, x_2164, x_2165, x_2166, x_2167, x_2168, x_2169, x_2170, x_2171, x_2172, x_2173, x_2174, x_2175, x_2176, x_2177, x_2178, x_2179, x_2180, x_2181, x_2182, x_2183, x_2184, x_2185, x_2186, x_2187, x_2188, x_2189, x_2190, x_2191, x_2192, x_2193, x_2194, x_2195, x_2196, x_2197, x_2198, x_2199, x_2200, x_2201, x_2202, x_2203, x_2204, x_2205, x_2206, x_2207, x_2208, x_2209, x_2210, x_2211, x_2212, x_2213, x_2214, x_2215, x_2216, x_2217, x_2218, x_2219, x_2220, x_2221, x_2222, x_2223, x_2224, x_2225, x_2226, x_2227, x_2228, x_2229, x_2230, x_2231, x_2232, x_2233, x_2234, x_2235, x_2236, x_2237, x_2238, x_2239, x_2240, x_2241, x_2242, x_2243, x_2244, x_2245, x_2246, x_2247, x_2248, x_2249, x_2250, x_2251, x_2252, x_2253, x_2254, x_2255, x_2256, x_2257, x_2258, x_2259, x_2260, x_2261, x_2262, x_2263, x_2264, x_2265, x_2266, x_2267, x_2268, x_2269, x_2270, x_2271, x_2272, x_2273, x_2274, x_2275, x_2276, x_2277, x_2278, x_2279, x_2280, x_2281, x_2282, x_2283, x_2284, x_2285, x_2286, x_2287, x_2288, x_2289, x_2290, x_2291, x_2292, x_2293, x_2294, x_2295, x_2296, x_2297, x_2298, x_2299, x_2300, x_2301, x_2302, x_2303, x_2304, x_2305, x_2306, x_2307, x_2308, x_2309, x_2310, x_2311, x_2312, x_2313, x_2314, x_2315, x_2316, x_2317, x_2318, x_2319, x_2320, x_2321, x_2322, x_2323, x_2324, x_2325, x_2326, x_2327, x_2328, x_2329, x_2330, x_2331, x_2332, x_2333, x_2334, x_2335, x_2336, x_2337, x_2338, x_2339, x_2340, x_2341, x_2342, x_2343, x_2344, x_2345, x_2346, x_2347, x_2348, x_2349, x_2350, x_2351, x_2352, x_2353, x_2354, x_2355, x_2356, x_2357, x_2358, x_2359, x_2360, x_2361, x_2362, x_2363, x_2364, x_2365, x_2366, x_2367, x_2368, x_2369, x_2370, x_2371, x_2372, x_2373, x_2374, x_2375, x_2376, x_2377, x_2378, x_2379, x_2380, x_2381, x_2382, x_2383, x_2384, x_2385, x_2386, x_2387, x_2388, x_2389, x_2390, x_2391, x_2392, x_2393, x_2394, x_2395, x_2396, x_2397, x_2398, x_2399, x_2400, x_2401, x_2402, x_2403, x_2404, x_2405, x_2406, x_2407, x_2408, x_2409, x_2410, x_2411, x_2412, x_2413, x_2414, x_2415, x_2416, x_2417, x_2418, x_2419, x_2420, x_2421, x_2422, x_2423, x_2424, x_2425, x_2426, x_2427, x_2428, x_2429, x_2430, x_2431, x_2432, x_2433, x_2434, x_2435, x_2436, x_2437, x_2438, x_2439, x_2440, x_2441, x_2442, x_2443, x_2444, x_2445, x_2446, x_2447, x_2448, x_2449, x_2450, x_2451, x_2452, x_2453, x_2454, x_2455, x_2456, x_2457, x_2458, x_2459, x_2460, x_2461, x_2462, x_2463, x_2464, x_2465, x_2466, x_2467, x_2468, x_2469, x_2470, x_2471, x_2472, x_2473, x_2474, x_2475, x_2476, x_2477, x_2478, x_2479, x_2480, x_2481, x_2482, x_2483, x_2484, x_2485, x_2486, x_2487, x_2488, x_2489, x_2490, x_2491, x_2492, x_2493, x_2494, x_2495, x_2496, x_2497, x_2498, x_2499, x_2500, x_2501, x_2502, x_2503, x_2504, x_2505, x_2506, x_2507, x_2508, x_2509, x_2510, x_2511, x_2512, x_2513, x_2514, x_2515, x_2516, x_2517, x_2518, x_2519, x_2520, x_2521, x_2522, x_2523, x_2524, x_2525, x_2526, x_2527, x_2528, x_2529, x_2530, x_2531, x_2532, x_2533, x_2534, x_2535, x_2536, x_2537, x_2538, x_2539, x_2540, x_2541, x_2542, x_2543, x_2544, x_2545, x_2546, x_2547, x_2548, x_2549, x_2550, x_2551, x_2552, x_2553, x_2554, x_2555, x_2556, x_2557, x_2558, x_2559, x_2560, x_2561, x_2562, x_2563, x_2564, x_2565, x_2566, x_2567, x_2568, x_2569, x_2570, x_2571, x_2572, x_2573, x_2574, x_2575, x_2576, x_2577, x_2578, x_2579, x_2580, x_2581, x_2582, x_2583, x_2584, x_2585, x_2586, x_2587, x_2588, x_2589, x_2590, x_2591, x_2592, x_2593, x_2594, x_2595, x_2596, x_2597, x_2598, x_2599, x_2600, x_2601, x_2602, x_2603, x_2604, x_2605, x_2606, x_2607, x_2608, x_2609, x_2610, x_2611, x_2612, x_2613, x_2614, x_2615, x_2616, x_2617, x_2618, x_2619, x_2620, x_2621, x_2622, x_2623, x_2624, x_2625, x_2626, x_2627, x_2628, x_2629, x_2630, x_2631, x_2632, x_2633, x_2634, x_2635, x_2636, x_2637, x_2638, x_2639, x_2640, x_2641, x_2642, x_2643, x_2644, x_2645, x_2646, x_2647, x_2648, x_2649, x_2650, x_2651, x_2652, x_2653, x_2654, x_2655, x_2656, x_2657, x_2658, x_2659, x_2660, x_2661, x_2662, x_2663, x_2664, x_2665, x_2666, x_2667, x_2668, x_2669, x_2670, x_2671, x_2672, x_2673, x_2674, x_2675, x_2676, x_2677, x_2678, x_2679, x_2680, x_2681, x_2682, x_2683, x_2684, x_2685, x_2686, x_2687, x_2688, x_2689, x_2690, x_2691, x_2692, x_2693, x_2694, x_2695, x_2696, x_2697, x_2698, x_2699, x_2700, x_2701, x_2702, x_2703, x_2704, x_2705, x_2706, x_2707, x_2708, x_2709, x_2710, x_2711, x_2712, x_2713, x_2714, x_2715, x_2716, x_2717, x_2718, x_2719, x_2720, x_2721, x_2722, x_2723, x_2724, x_2725, x_2726, x_2727, x_2728, x_2729, x_2730, x_2731, x_2732, x_2733, x_2734, x_2735, x_2736, x_2737, x_2738, x_2739, x_2740, x_2741, x_2742, x_2743, x_2744, x_2745, x_2746, x_2747, x_2748, x_2749, x_2750, x_2751, x_2752, x_2753, x_2754, x_2755, x_2756, x_2757, x_2758, x_2759, x_2760, x_2761, x_2762, x_2763, x_2764, x_2765, x_2766, x_2767, x_2768, x_2769, x_2770, x_2771, x_2772, x_2773, x_2774, x_2775, x_2776, x_2777, x_2778, x_2779, x_2780, x_2781, x_2782, x_2783, x_2784, x_2785, x_2786, x_2787, x_2788, x_2789, x_2790, x_2791, x_2792, x_2793, x_2794, x_2795, x_2796, x_2797, x_2798, x_2799, x_2800, x_2801, x_2802, x_2803, x_2804, x_2805, x_2806, x_2807, x_2808, x_2809, x_2810, x_2811, x_2812, x_2813, x_2814, x_2815, x_2816, x_2817, x_2818, x_2819, x_2820, x_2821, x_2822, x_2823, x_2824, x_2825, x_2826, x_2827, x_2828, x_2829, x_2830, x_2831, x_2832, x_2833, x_2834, x_2835, x_2836, x_2837, x_2838, x_2839, x_2840, x_2841, x_2842, x_2843, x_2844, x_2845, x_2846, x_2847, x_2848, x_2849, x_2850, x_2851, x_2852, x_2853, x_2854, x_2855, x_2856, x_2857, x_2858, x_2859, x_2860, x_2861, x_2862, x_2863, x_2864, x_2865, x_2866, x_2867, x_2868, x_2869, x_2870, x_2871, x_2872, x_2873, x_2874, x_2875, x_2876, x_2877, x_2878, x_2879, x_2880, x_2881, x_2882, x_2883, x_2884, x_2885, x_2886, x_2887, x_2888, x_2889, x_2890, x_2891, x_2892, x_2893, x_2894, x_2895, x_2896, x_2897, x_2898, x_2899, x_2900, x_2901, x_2902, x_2903, x_2904, x_2905, x_2906, x_2907, x_2908, x_2909, x_2910, x_2911, x_2912, x_2913, x_2914, x_2915, x_2916, x_2917, x_2918, x_2919, x_2920, x_2921, x_2922, x_2923, x_2924, x_2925, x_2926, x_2927, x_2928, x_2929, x_2930, x_2931, x_2932, x_2933, x_2934, x_2935, x_2936, x_2937, x_2938, x_2939, x_2940, x_2941, x_2942, x_2943, x_2944, x_2945, x_2946, x_2947, x_2948, x_2949, x_2950, x_2951, x_2952, x_2953, x_2954, x_2955, x_2956, x_2957, x_2958, x_2959, x_2960, x_2961, x_2962, x_2963, x_2964, x_2965, x_2966, x_2967, x_2968, x_2969, x_2970, x_2971, x_2972, x_2973, x_2974, x_2975, x_2976, x_2977, x_2978, x_2979, x_2980, x_2981, x_2982, x_2983, x_2984, x_2985, x_2986, x_2987, x_2988, x_2989, x_2990, x_2991, x_2992, x_2993, x_2994, x_2995, x_2996, x_2997, x_2998, x_2999, x_3000, x_3001, x_3002, x_3003, x_3004, x_3005, x_3006, x_3007, x_3008, x_3009, x_3010, x_3011, x_3012, x_3013, x_3014, x_3015, x_3016, x_3017, x_3018, x_3019, x_3020, x_3021, x_3022, x_3023, x_3024, x_3025, x_3026, x_3027, x_3028, x_3029, x_3030, x_3031, x_3032, x_3033, x_3034, x_3035, x_3036, x_3037, x_3038, x_3039, x_3040, x_3041, x_3042, x_3043, x_3044, x_3045, x_3046, x_3047, x_3048, x_3049, x_3050, x_3051, x_3052, x_3053, x_3054, x_3055, x_3056, x_3057, x_3058, x_3059, x_3060, x_3061, x_3062, x_3063, x_3064, x_3065, x_3066, x_3067, x_3068, x_3069, x_3070, x_3071, x_3072, x_3073, x_3074, x_3075, x_3076, x_3077, x_3078, x_3079, x_3080, x_3081, x_3082, x_3083, x_3084, x_3085, x_3086, x_3087, x_3088, x_3089, x_3090, x_3091, x_3092, x_3093, x_3094, x_3095, x_3096, x_3097, x_3098, x_3099, x_3100, x_3101, x_3102, x_3103, x_3104, x_3105, x_3106, x_3107, x_3108, x_3109, x_3110, x_3111, x_3112, x_3113, x_3114, x_3115, x_3116, x_3117, x_3118, x_3119, x_3120, x_3121, x_3122, x_3123, x_3124, x_3125, x_3126, x_3127, x_3128, x_3129, x_3130, x_3131, x_3132, x_3133, x_3134, x_3135, x_3136, x_3137, x_3138, x_3139, x_3140, x_3141, x_3142, x_3143, x_3144, x_3145, x_3146, x_3147, x_3148, x_3149, x_3150, x_3151, x_3152, x_3153, x_3154, x_3155, x_3156, x_3157, x_3158, x_3159, x_3160, x_3161, x_3162, x_3163, x_3164, x_3165, x_3166, x_3167, x_3168, x_3169, x_3170, x_3171, x_3172, x_3173, x_3174, x_3175, x_3176, x_3177, x_3178, x_3179, x_3180, x_3181, x_3182, x_3183, x_3184, x_3185, x_3186, x_3187, x_3188, x_3189, x_3190, x_3191, x_3192, x_3193, x_3194, x_3195, x_3196, x_3197, x_3198, x_3199, x_3200, x_3201, x_3202, x_3203, x_3204, x_3205, x_3206, x_3207, x_3208, x_3209, x_3210, x_3211, x_3212, x_3213, x_3214, x_3215, x_3216, x_3217, x_3218, x_3219, x_3220, x_3221, x_3222, x_3223, x_3224, x_3225, x_3226, x_3227, x_3228, x_3229, x_3230, x_3231, x_3232, x_3233, x_3234, x_3235, x_3236, x_3237, x_3238, x_3239, x_3240, x_3241, x_3242, x_3243, x_3244, x_3245, x_3246, x_3247, x_3248, x_3249, x_3250, x_3251, x_3252, x_3253, x_3254, x_3255, x_3256, x_3257, x_3258, x_3259, x_3260, x_3261, x_3262, x_3263, x_3264, x_3265, x_3266, x_3267, x_3268, x_3269, x_3270, x_3271, x_3272, x_3273, x_3274, x_3275, x_3276, x_3277, x_3278, x_3279, x_3280, x_3281, x_3282, x_3283, x_3284, x_3285, x_3286, x_3287, x_3288, x_3289, x_3290, x_3291, x_3292, x_3293, x_3294, x_3295, x_3296, x_3297, x_3298, x_3299, x_3300, x_3301, x_3302, x_3303, x_3304, x_3305, x_3306, x_3307, x_3308, x_3309, x_3310, x_3311, x_3312, x_3313, x_3314, x_3315, x_3316, x_3317, x_3318, x_3319, x_3320, x_3321, x_3322, x_3323, x_3324, x_3325, x_3326, x_3327, x_3328, x_3329, x_3330, x_3331, x_3332, x_3333, x_3334, x_3335, x_3336, x_3337, x_3338, x_3339, x_3340, x_3341, x_3342, x_3343, x_3344, x_3345, x_3346, x_3347, x_3348, x_3349, x_3350, x_3351, x_3352, x_3353, x_3354, x_3355, x_3356, x_3357, x_3358, x_3359, x_3360, x_3361, x_3362, x_3363, x_3364, x_3365, x_3366, x_3367, x_3368, x_3369, x_3370, x_3371, x_3372, x_3373, x_3374, x_3375, x_3376, x_3377, x_3378, x_3379, x_3380, x_3381, x_3382, x_3383, x_3384, x_3385, x_3386, x_3387, x_3388, x_3389, x_3390, x_3391, x_3392, x_3393, x_3394, x_3395, x_3396, x_3397, x_3398, x_3399, x_3400, x_3401, x_3402, x_3403, x_3404, x_3405, x_3406, x_3407, x_3408, x_3409, x_3410, x_3411, x_3412, x_3413, x_3414, x_3415, x_3416, x_3417, x_3418, x_3419, x_3420, x_3421, x_3422, x_3423, x_3424, x_3425, x_3426, x_3427, x_3428, x_3429, x_3430, x_3431, x_3432, x_3433, x_3434, x_3435, x_3436, x_3437, x_3438, x_3439, x_3440, x_3441, x_3442, x_3443, x_3444, x_3445, x_3446, x_3447, x_3448, x_3449, x_3450, x_3451, x_3452, x_3453, x_3454, x_3455, x_3456, x_3457, x_3458, x_3459, x_3460, x_3461, x_3462, x_3463, x_3464, x_3465, x_3466, x_3467, x_3468, x_3469, x_3470, x_3471, x_3472, x_3473, x_3474, x_3475, x_3476, x_3477, x_3478, x_3479, x_3480, x_3481, x_3482, x_3483, x_3484, x_3485, x_3486, x_3487, x_3488, x_3489, x_3490, x_3491, x_3492, x_3493, x_3494, x_3495, x_3496, x_3497, x_3498, x_3499, x_3500, x_3501, x_3502, x_3503, x_3504, x_3505, x_3506, x_3507, x_3508, x_3509, x_3510, x_3511, x_3512, x_3513, x_3514, x_3515, x_3516, x_3517, x_3518, x_3519, x_3520, x_3521, x_3522, x_3523, x_3524, x_3525, x_3526, x_3527, x_3528, x_3529, x_3530, x_3531, x_3532, x_3533, x_3534, x_3535, x_3536, x_3537, x_3538, x_3539, x_3540, x_3541, x_3542, x_3543, x_3544, x_3545, x_3546, x_3547, x_3548, x_3549, x_3550, x_3551, x_3552, x_3553, x_3554, x_3555, x_3556, x_3557, x_3558, x_3559, x_3560, x_3561, x_3562, x_3563, x_3564, x_3565, x_3566, x_3567, x_3568, x_3569, x_3570, x_3571, x_3572, x_3573, x_3574, x_3575, x_3576, x_3577, x_3578, x_3579, x_3580, x_3581, x_3582, x_3583, x_3584, x_3585, x_3586, x_3587, x_3588, x_3589, x_3590, x_3591, x_3592, x_3593, x_3594, x_3595, x_3596, x_3597, x_3598, x_3599, x_3600, x_3601, x_3602, x_3603, x_3604, x_3605, x_3606, x_3607, x_3608, x_3609, x_3610, x_3611, x_3612, x_3613, x_3614, x_3615, x_3616, x_3617, x_3618, x_3619, x_3620, x_3621, x_3622, x_3623, x_3624, x_3625, x_3626, x_3627, x_3628, x_3629, x_3630, x_3631, x_3632, x_3633, x_3634, x_3635, x_3636, x_3637, x_3638, x_3639, x_3640, x_3641, x_3642, x_3643, x_3644, x_3645, x_3646, x_3647, x_3648, x_3649, x_3650, x_3651, x_3652, x_3653, x_3654, x_3655, x_3656, x_3657, x_3658, x_3659, x_3660, x_3661, x_3662, x_3663, x_3664, x_3665, x_3666, x_3667, x_3668, x_3669, x_3670, x_3671, x_3672, x_3673, x_3674, x_3675, x_3676, x_3677, x_3678, x_3679, x_3680, x_3681, x_3682, x_3683, x_3684, x_3685, x_3686, x_3687, x_3688, x_3689, x_3690, x_3691, x_3692, x_3693, x_3694, x_3695, x_3696, x_3697, x_3698, x_3699, x_3700, x_3701, x_3702, x_3703, x_3704, x_3705, x_3706, x_3707, x_3708, x_3709, x_3710, x_3711, x_3712, x_3713, x_3714, x_3715, x_3716, x_3717, x_3718, x_3719, x_3720, x_3721, x_3722, x_3723, x_3724, x_3725, x_3726, x_3727, x_3728, x_3729, x_3730, x_3731, x_3732, x_3733, x_3734, x_3735, x_3736, x_3737, x_3738, x_3739, x_3740, x_3741, x_3742, x_3743, x_3744, x_3745, x_3746, x_3747, x_3748, x_3749, x_3750, x_3751, x_3752, x_3753, x_3754, x_3755, x_3756, x_3757, x_3758, x_3759, x_3760, x_3761, x_3762, x_3763, x_3764, x_3765, x_3766, x_3767, x_3768, x_3769, x_3770, x_3771, x_3772, x_3773, x_3774, x_3775, x_3776, x_3777, x_3778, x_3779, x_3780, x_3781, x_3782, x_3783, x_3784, x_3785, x_3786, x_3787, x_3788, x_3789, x_3790, x_3791, x_3792, x_3793, x_3794, x_3795, x_3796, x_3797, x_3798, x_3799, x_3800, x_3801, x_3802, x_3803, x_3804, x_3805, x_3806, x_3807, x_3808, x_3809, x_3810, x_3811, x_3812, x_3813, x_3814, x_3815, x_3816, x_3817, x_3818, x_3819, x_3820, x_3821, x_3822, x_3823, x_3824, x_3825, x_3826, x_3827, x_3828, x_3829, x_3830, x_3831, x_3832, x_3833, x_3834, x_3835, x_3836, x_3837, x_3838, x_3839, x_3840, x_3841, x_3842, x_3843, x_3844, x_3845, x_3846, x_3847, x_3848, x_3849, x_3850, x_3851, x_3852, x_3853, x_3854, x_3855, x_3856, x_3857, x_3858, x_3859, x_3860, x_3861, x_3862, x_3863, x_3864, x_3865, x_3866, x_3867, x_3868, x_3869, x_3870, x_3871, x_3872, x_3873, x_3874, x_3875, x_3876, x_3877, x_3878, x_3879, x_3880, x_3881, x_3882, x_3883, x_3884, x_3885, x_3886, x_3887, x_3888, x_3889, x_3890, x_3891, x_3892, x_3893, x_3894, x_3895, x_3896, x_3897, x_3898, x_3899, x_3900, x_3901, x_3902, x_3903, x_3904, x_3905, x_3906, x_3907, x_3908, x_3909, x_3910, x_3911, x_3912, x_3913, x_3914, x_3915, x_3916, x_3917, x_3918, x_3919, x_3920, x_3921, x_3922, x_3923, x_3924, x_3925, x_3926, x_3927, x_3928, x_3929, x_3930, x_3931, x_3932, x_3933, x_3934, x_3935, x_3936, x_3937, x_3938, x_3939, x_3940, x_3941, x_3942, x_3943, x_3944, x_3945, x_3946, x_3947, x_3948, x_3949, x_3950, x_3951, x_3952, x_3953, x_3954, x_3955, x_3956, x_3957, x_3958, x_3959, x_3960, x_3961, x_3962, x_3963, x_3964, x_3965, x_3966, x_3967, x_3968, x_3969, x_3970, x_3971, x_3972, x_3973, x_3974, x_3975, x_3976, x_3977, x_3978, x_3979, x_3980, x_3981, x_3982, x_3983, x_3984, x_3985, x_3986, x_3987, x_3988, x_3989, x_3990, x_3991, x_3992, x_3993, x_3994, x_3995, x_3996, x_3997, x_3998, x_3999, x_4000, x_4001, x_4002, x_4003, x_4004, x_4005, x_4006, x_4007, x_4008, x_4009, x_4010, x_4011, x_4012, x_4013, x_4014, x_4015, x_4016, x_4017, x_4018, x_4019, x_4020, x_4021, x_4022, x_4023, x_4024, x_4025, x_4026, x_4027, x_4028, x_4029, x_4030, x_4031, x_4032, x_4033, x_4034, x_4035, x_4036, x_4037, x_4038, x_4039, x_4040, x_4041, x_4042, x_4043, x_4044, x_4045, x_4046, x_4047, x_4048, x_4049, x_4050, x_4051, x_4052, x_4053, x_4054, x_4055, x_4056, x_4057, x_4058, x_4059, x_4060, x_4061, x_4062, x_4063, x_4064, x_4065, x_4066, x_4067, x_4068, x_4069, x_4070, x_4071, x_4072, x_4073, x_4074, x_4075, x_4076, x_4077, x_4078, x_4079, x_4080, x_4081, x_4082, x_4083, x_4084, x_4085, x_4086, x_4087, x_4088, x_4089, x_4090, x_4091, x_4092, x_4093, x_4094, x_4095, x_4096, x_4097, x_4098, x_4099, x_4100, x_4101, x_4102, x_4103, x_4104, x_4105, x_4106, x_4107, x_4108, x_4109, x_4110, x_4111, x_4112, x_4113, x_4114, x_4115, x_4116, x_4117, x_4118, x_4119, x_4120, x_4121, x_4122, x_4123, x_4124, x_4125, x_4126, x_4127, x_4128, x_4129, x_4130, x_4131, x_4132, x_4133, x_4134, x_4135, x_4136, x_4137, x_4138, x_4139, x_4140, x_4141, x_4142, x_4143, x_4144, x_4145, x_4146, x_4147, x_4148, x_4149, x_4150, x_4151, x_4152, x_4153, x_4154, x_4155, x_4156, x_4157, x_4158, x_4159, x_4160, x_4161, x_4162, x_4163, x_4164, x_4165, x_4166, x_4167, x_4168, x_4169, x_4170, x_4171, x_4172, x_4173, x_4174, x_4175, x_4176, x_4177, x_4178, x_4179, x_4180, x_4181, x_4182, x_4183, x_4184, x_4185, x_4186, x_4187, x_4188, x_4189, x_4190, x_4191, x_4192, x_4193, x_4194, x_4195, x_4196, x_4197, x_4198, x_4199, x_4200, x_4201, x_4202, x_4203, x_4204, x_4205, x_4206, x_4207, x_4208, x_4209, x_4210, x_4211, x_4212, x_4213, x_4214, x_4215, x_4216, x_4217, x_4218, x_4219, x_4220, x_4221, x_4222, x_4223, x_4224, x_4225, x_4226, x_4227, x_4228, x_4229, x_4230, x_4231, x_4232, x_4233, x_4234, x_4235, x_4236, x_4237, x_4238, x_4239, x_4240, x_4241, x_4242, x_4243, x_4244, x_4245, x_4246, x_4247, x_4248, x_4249, x_4250, x_4251, x_4252, x_4253, x_4254, x_4255, x_4256, x_4257, x_4258, x_4259, x_4260, x_4261, x_4262, x_4263, x_4264, x_4265, x_4266, x_4267, x_4268, x_4269, x_4270, x_4271, x_4272, x_4273, x_4274, x_4275, x_4276, x_4277, x_4278, x_4279, x_4280, x_4281, x_4282, x_4283, x_4284, x_4285, x_4286, x_4287, x_4288, x_4289, x_4290, x_4291, x_4292, x_4293, x_4294, x_4295, x_4296, x_4297, x_4298, x_4299, x_4300, x_4301, x_4302, x_4303, x_4304, x_4305, x_4306, x_4307, x_4308, x_4309, x_4310, x_4311, x_4312, x_4313, x_4314, x_4315, x_4316, x_4317, x_4318, x_4319, x_4320, x_4321, x_4322, x_4323, x_4324, x_4325, x_4326, x_4327, x_4328, x_4329, x_4330, x_4331, x_4332, x_4333, x_4334, x_4335, x_4336, x_4337, x_4338, x_4339, x_4340, x_4341, x_4342, x_4343, x_4344, x_4345, x_4346, x_4347, x_4348, x_4349, x_4350, x_4351, x_4352, x_4353, x_4354, x_4355, x_4356, x_4357, x_4358, x_4359, x_4360, x_4361, x_4362, x_4363, x_4364, x_4365, x_4366, x_4367, x_4368, x_4369, x_4370, x_4371, x_4372, x_4373, x_4374, x_4375, x_4376, x_4377, x_4378, x_4379, x_4380, x_4381, x_4382, x_4383, x_4384, x_4385, x_4386, x_4387, x_4388, x_4389, x_4390, x_4391, x_4392, x_4393, x_4394, x_4395, x_4396, x_4397, x_4398, x_4399, x_4400, x_4401, x_4402, x_4403, x_4404, x_4405, x_4406, x_4407, x_4408, x_4409, x_4410, x_4411, x_4412, x_4413, x_4414, x_4415, x_4416, x_4417, x_4418, x_4419, x_4420, x_4421, x_4422, x_4423, x_4424, x_4425, x_4426, x_4427, x_4428, x_4429, x_4430, x_4431, x_4432, x_4433, x_4434, x_4435, x_4436, x_4437, x_4438, x_4439, x_4440, x_4441, x_4442, x_4443, x_4444, x_4445, x_4446, x_4447, x_4448, x_4449, x_4450, x_4451, x_4452, x_4453, x_4454, x_4455, x_4456, x_4457, x_4458, x_4459, x_4460, x_4461, x_4462, x_4463, x_4464, x_4465, x_4466, x_4467, x_4468, x_4469, x_4470, x_4471, x_4472, x_4473, x_4474, x_4475, x_4476, x_4477, x_4478, x_4479, x_4480, x_4481, x_4482, x_4483, x_4484, x_4485, x_4486, x_4487, x_4488, x_4489, x_4490, x_4491, x_4492, x_4493, x_4494, x_4495, x_4496, x_4497, x_4498, x_4499, x_4500, x_4501, x_4502, x_4503, x_4504, x_4505, x_4506, x_4507, x_4508, x_4509, x_4510, x_4511, x_4512, x_4513, x_4514, x_4515, x_4516, x_4517, x_4518, x_4519, x_4520, x_4521, x_4522, x_4523, x_4524, x_4525, x_4526, x_4527, x_4528, x_4529, x_4530, x_4531, x_4532, x_4533, x_4534, x_4535, x_4536, x_4537, x_4538, x_4539, x_4540, x_4541, x_4542, x_4543, x_4544, x_4545, x_4546, x_4547, x_4548, x_4549, x_4550, x_4551, x_4552, x_4553, x_4554, x_4555, x_4556, x_4557, x_4558, x_4559, x_4560, x_4561, x_4562, x_4563, x_4564, x_4565, x_4566, x_4567, x_4568, x_4569, x_4570, x_4571, x_4572, x_4573, x_4574, x_4575, x_4576, x_4577, x_4578, x_4579, x_4580, x_4581, x_4582, x_4583, x_4584, x_4585, x_4586, x_4587, x_4588, x_4589, x_4590, x_4591, x_4592, x_4593, x_4594, x_4595, x_4596, x_4597, x_4598, x_4599, x_4600, x_4601, x_4602, x_4603, x_4604, x_4605, x_4606, x_4607, x_4608, x_4609, x_4610, x_4611, x_4612, x_4613, x_4614, x_4615, x_4616, x_4617, x_4618, x_4619, x_4620, x_4621, x_4622, x_4623, x_4624, x_4625, x_4626, x_4627, x_4628, x_4629, x_4630, x_4631, x_4632, x_4633, x_4634, x_4635, x_4636, x_4637, x_4638, x_4639, x_4640, x_4641, x_4642, x_4643, x_4644, x_4645, x_4646, x_4647, x_4648, x_4649, x_4650, x_4651, x_4652, x_4653, x_4654, x_4655, x_4656, x_4657, x_4658, x_4659, x_4660, x_4661, x_4662, x_4663, x_4664, x_4665, x_4666, x_4667, x_4668, x_4669, x_4670, x_4671, x_4672, x_4673, x_4674, x_4675, x_4676, x_4677, x_4678, x_4679, x_4680, x_4681, x_4682, x_4683, x_4684, x_4685, x_4686, x_4687, x_4688, x_4689, x_4690, x_4691, x_4692, x_4693, x_4694, x_4695, x_4696, x_4697, x_4698, x_4699, x_4700, x_4701, x_4702, x_4703, x_4704, x_4705, x_4706, x_4707, x_4708, x_4709, x_4710, x_4711, x_4712, x_4713, x_4714, x_4715, x_4716, x_4717, x_4718, x_4719, x_4720, x_4721, x_4722, x_4723, x_4724, x_4725, x_4726, x_4727, x_4728, x_4729, x_4730, x_4731, x_4732, x_4733, x_4734, x_4735, x_4736, x_4737, x_4738, x_4739, x_4740, x_4741, x_4742, x_4743, x_4744, x_4745, x_4746, x_4747, x_4748, x_4749, x_4750, x_4751, x_4752, x_4753, x_4754, x_4755, x_4756, x_4757, x_4758, x_4759, x_4760, x_4761, x_4762, x_4763, x_4764, x_4765, x_4766, x_4767, x_4768, x_4769, x_4770, x_4771, x_4772, x_4773, x_4774, x_4775, x_4776, x_4777, x_4778, x_4779, x_4780, x_4781, x_4782, x_4783, x_4784, x_4785, x_4786, x_4787, x_4788, x_4789, x_4790, x_4791, x_4792, x_4793, x_4794, x_4795, x_4796, x_4797, x_4798, x_4799, x_4800, x_4801, x_4802, x_4803, x_4804, x_4805, x_4806, x_4807, x_4808, x_4809, x_4810, x_4811, x_4812, x_4813, x_4814, x_4815, x_4816, x_4817, x_4818, x_4819, x_4820, x_4821, x_4822, x_4823, x_4824, x_4825, x_4826, x_4827, x_4828, x_4829, x_4830, x_4831, x_4832, x_4833, x_4834, x_4835, x_4836, x_4837, x_4838, x_4839, x_4840, x_4841, x_4842, x_4843, x_4844, x_4845, x_4846, x_4847, x_4848, x_4849, x_4850, x_4851, x_4852, x_4853, x_4854, x_4855, x_4856, x_4857, x_4858, x_4859, x_4860, x_4861, x_4862, x_4863, x_4864, x_4865, x_4866, x_4867, x_4868, x_4869, x_4870, x_4871, x_4872, x_4873, x_4874, x_4875, x_4876, x_4877, x_4878, x_4879, x_4880, x_4881, x_4882, x_4883, x_4884, x_4885, x_4886, x_4887, x_4888, x_4889, x_4890, x_4891, x_4892, x_4893, x_4894, x_4895, x_4896, x_4897, x_4898, x_4899, x_4900, x_4901, x_4902, x_4903, x_4904, x_4905, x_4906, x_4907, x_4908, x_4909, x_4910, x_4911, x_4912, x_4913, x_4914, x_4915, x_4916, x_4917, x_4918, x_4919, x_4920, x_4921, x_4922, x_4923, x_4924, x_4925, x_4926, x_4927, x_4928, x_4929, x_4930, x_4931, x_4932, x_4933, x_4934, x_4935, x_4936, x_4937, x_4938, x_4939, x_4940, x_4941, x_4942, x_4943, x_4944, x_4945, x_4946, x_4947, x_4948, x_4949, x_4950, x_4951, x_4952, x_4953, x_4954, x_4955, x_4956, x_4957, x_4958, x_4959, x_4960, x_4961, x_4962, x_4963, x_4964, x_4965, x_4966, x_4967, x_4968, x_4969, x_4970, x_4971, x_4972, x_4973, x_4974, x_4975, x_4976, x_4977, x_4978, x_4979, x_4980, x_4981, x_4982, x_4983, x_4984, x_4985, x_4986, x_4987, x_4988, x_4989, x_4990, x_4991, x_4992, x_4993, x_4994, x_4995, x_4996, x_4997, x_4998, x_4999, x_5000, x_5001, x_5002, x_5003, x_5004, x_5005, x_5006, x_5007, x_5008, x_5009, x_5010, x_5011, x_5012, x_5013, x_5014, x_5015, x_5016, x_5017, x_5018, x_5019, x_5020, x_5021, x_5022, x_5023, x_5024, x_5025, x_5026, x_5027, x_5028, x_5029, x_5030, x_5031, x_5032, x_5033, x_5034, x_5035, x_5036, x_5037, x_5038, x_5039, x_5040, x_5041, x_5042, x_5043, x_5044, x_5045, x_5046, x_5047, x_5048, x_5049, x_5050, x_5051, x_5052, x_5053, x_5054, x_5055, x_5056, x_5057, x_5058, x_5059, x_5060, x_5061, x_5062, x_5063, x_5064, x_5065, x_5066, x_5067, x_5068, x_5069, x_5070, x_5071, x_5072, x_5073, x_5074, x_5075, x_5076, x_5077, x_5078, x_5079, x_5080, x_5081, x_5082, x_5083, x_5084, x_5085, x_5086, x_5087, x_5088, x_5089, x_5090, x_5091, x_5092, x_5093, x_5094, x_5095, x_5096, x_5097, x_5098, x_5099, x_5100, x_5101, x_5102, x_5103, x_5104, x_5105, x_5106, x_5107, x_5108, x_5109, x_5110, x_5111, x_5112, x_5113, x_5114, x_5115, x_5116, x_5117, x_5118, x_5119, x_5120, x_5121, x_5122, x_5123, x_5124, x_5125, x_5126, x_5127, x_5128, x_5129, x_5130, x_5131, x_5132, x_5133, x_5134, x_5135, x_5136, x_5137, x_5138, x_5139, x_5140, x_5141, x_5142, x_5143, x_5144, x_5145, x_5146, x_5147, x_5148, x_5149, x_5150, x_5151, x_5152, x_5153, x_5154, x_5155, x_5156, x_5157, x_5158, x_5159, x_5160, x_5161, x_5162, x_5163, x_5164, x_5165, x_5166, x_5167, x_5168, x_5169, x_5170, x_5171, x_5172, x_5173, x_5174, x_5175, x_5176, x_5177, x_5178, x_5179, x_5180, x_5181, x_5182, x_5183, x_5184, x_5185, x_5186, x_5187, x_5188, x_5189, x_5190, x_5191, x_5192, x_5193, x_5194, x_5195, x_5196, x_5197, x_5198, x_5199, x_5200, x_5201, x_5202, x_5203, x_5204, x_5205, x_5206, x_5207, x_5208, x_5209, x_5210, x_5211, x_5212, x_5213, x_5214, x_5215, x_5216, x_5217, x_5218, x_5219, x_5220, x_5221, x_5222, x_5223, x_5224, x_5225, x_5226, x_5227, x_5228, x_5229, x_5230, x_5231, x_5232, x_5233, x_5234, x_5235, x_5236, x_5237, x_5238, x_5239, x_5240, x_5241, x_5242, x_5243, x_5244, x_5245, x_5246, x_5247, x_5248, x_5249, x_5250, x_5251, x_5252, x_5253, x_5254, x_5255, x_5256, x_5257, x_5258, x_5259, x_5260, x_5261, x_5262, x_5263, x_5264, x_5265, x_5266, x_5267, x_5268, x_5269, x_5270, x_5271, x_5272, x_5273, x_5274, x_5275, x_5276, x_5277, x_5278, x_5279, x_5280, x_5281, x_5282, x_5283, x_5284, x_5285, x_5286, x_5287, x_5288, x_5289, x_5290, x_5291, x_5292, x_5293, x_5294, x_5295, x_5296, x_5297, x_5298, x_5299, x_5300, x_5301, x_5302, x_5303, x_5304, x_5305, x_5306, x_5307, x_5308, x_5309, x_5310, x_5311, x_5312, x_5313, x_5314, x_5315, x_5316, x_5317, x_5318, x_5319, x_5320, x_5321, x_5322, x_5323, x_5324, x_5325, x_5326, x_5327, x_5328, x_5329, x_5330, x_5331, x_5332, x_5333, x_5334, x_5335, x_5336, x_5337, x_5338, x_5339, x_5340, x_5341, x_5342, x_5343, x_5344, x_5345, x_5346, x_5347, x_5348, x_5349, x_5350, x_5351, x_5352, x_5353, x_5354, x_5355, x_5356, x_5357, x_5358, x_5359, x_5360, x_5361, x_5362, x_5363, x_5364, x_5365, x_5366, x_5367, x_5368, x_5369, x_5370, x_5371, x_5372, x_5373, x_5374, x_5375, x_5376, x_5377, x_5378, x_5379, x_5380, x_5381, x_5382, x_5383, x_5384, x_5385, x_5386, x_5387, x_5388, x_5389, x_5390, x_5391, x_5392, x_5393, x_5394, x_5395, x_5396, x_5397, x_5398, x_5399, x_5400, x_5401, x_5402, x_5403, x_5404, x_5405, x_5406, x_5407, x_5408, x_5409, x_5410, x_5411, x_5412, x_5413, x_5414, x_5415, x_5416, x_5417, x_5418, x_5419, x_5420, x_5421, x_5422, x_5423, x_5424, x_5425, x_5426, x_5427, x_5428, x_5429, x_5430, x_5431, x_5432, x_5433, x_5434, x_5435, x_5436, x_5437, x_5438, x_5439, x_5440, x_5441, x_5442, x_5443, x_5444, x_5445, x_5446, x_5447, x_5448, x_5449, x_5450, x_5451, x_5452, x_5453, x_5454, x_5455, x_5456, x_5457, x_5458, x_5459, x_5460, x_5461, x_5462, x_5463, x_5464, x_5465, x_5466, x_5467, x_5468, x_5469, x_5470, x_5471, x_5472, x_5473, x_5474, x_5475, x_5476, x_5477, x_5478, x_5479, x_5480, x_5481, x_5482, x_5483, x_5484, x_5485, x_5486, x_5487, x_5488, x_5489, x_5490, x_5491, x_5492, x_5493, x_5494, x_5495, x_5496, x_5497, x_5498, x_5499, x_5500, x_5501, x_5502, x_5503, x_5504, x_5505, x_5506, x_5507, x_5508, x_5509, x_5510, x_5511, x_5512, x_5513, x_5514, x_5515, x_5516, x_5517, x_5518, x_5519, x_5520, x_5521, x_5522, x_5523, x_5524, x_5525, x_5526, x_5527, x_5528, x_5529, x_5530, x_5531, x_5532, x_5533, x_5534, x_5535, x_5536, x_5537, x_5538, x_5539, x_5540, x_5541, x_5542, x_5543, x_5544, x_5545, x_5546, x_5547, x_5548, x_5549, x_5550, x_5551, x_5552, x_5553, x_5554, x_5555, x_5556, x_5557, x_5558, x_5559, x_5560, x_5561, x_5562, x_5563, x_5564, x_5565, x_5566, x_5567, x_5568, x_5569, x_5570, x_5571, x_5572, x_5573, x_5574, x_5575, x_5576, x_5577, x_5578, x_5579, x_5580, x_5581, x_5582, x_5583, x_5584, x_5585, x_5586, x_5587, x_5588, x_5589, x_5590, x_5591, x_5592, x_5593, x_5594, x_5595, x_5596, x_5597, x_5598, x_5599, x_5600, x_5601, x_5602, x_5603, x_5604, x_5605, x_5606, x_5607, x_5608, x_5609, x_5610, x_5611, x_5612, x_5613, x_5614, x_5615, x_5616, x_5617, x_5618, x_5619, x_5620, x_5621, x_5622, x_5623, x_5624, x_5625, x_5626, x_5627, x_5628, x_5629, x_5630, x_5631, x_5632, x_5633, x_5634, x_5635, x_5636, x_5637, x_5638, x_5639, x_5640, x_5641, x_5642, x_5643, x_5644, x_5645, x_5646, x_5647, x_5648, x_5649, x_5650, x_5651, x_5652, x_5653, x_5654, x_5655, x_5656, x_5657, x_5658, x_5659, x_5660, x_5661, x_5662, x_5663, x_5664, x_5665, x_5666, x_5667, x_5668, x_5669, x_5670, x_5671, x_5672, x_5673, x_5674, x_5675, x_5676, x_5677, x_5678, x_5679, x_5680, x_5681, x_5682, x_5683, x_5684, x_5685, x_5686, x_5687, x_5688, x_5689, x_5690, x_5691, x_5692, x_5693, x_5694, x_5695, x_5696, x_5697, x_5698, x_5699, x_5700, x_5701, x_5702, x_5703, x_5704, x_5705, x_5706, x_5707, x_5708, x_5709, x_5710, x_5711, x_5712, x_5713, x_5714, x_5715, x_5716, x_5717, x_5718, x_5719, x_5720, x_5721, x_5722, x_5723, x_5724, x_5725, x_5726, x_5727, x_5728, x_5729, x_5730, x_5731, x_5732, x_5733, x_5734, x_5735, x_5736, x_5737, x_5738, x_5739, x_5740, x_5741, x_5742, x_5743, x_5744, x_5745, x_5746, x_5747, x_5748, x_5749, x_5750, x_5751, x_5752, x_5753, x_5754, x_5755, x_5756, x_5757, x_5758, x_5759, x_5760, x_5761, x_5762, x_5763, x_5764, x_5765, x_5766, x_5767, x_5768, x_5769, x_5770, x_5771, x_5772, x_5773, x_5774, x_5775, x_5776, x_5777, x_5778, x_5779, x_5780, x_5781, x_5782, x_5783, x_5784, x_5785, x_5786, x_5787, x_5788, x_5789, x_5790, x_5791, x_5792, x_5793, x_5794, x_5795, x_5796, x_5797, x_5798, x_5799, x_5800, x_5801, x_5802, x_5803, x_5804, x_5805, x_5806, x_5807, x_5808, x_5809, x_5810, x_5811, x_5812, x_5813, x_5814, x_5815, x_5816, x_5817, x_5818, x_5819, x_5820, x_5821, x_5822, x_5823, x_5824, x_5825, x_5826, x_5827, x_5828, x_5829, x_5830, x_5831, x_5832, x_5833, x_5834, x_5835, x_5836, x_5837, x_5838, x_5839, x_5840, x_5841, x_5842, x_5843, x_5844, x_5845, x_5846, x_5847, x_5848, x_5849, x_5850, x_5851, x_5852, x_5853, x_5854, x_5855, x_5856, x_5857, x_5858, x_5859, x_5860, x_5861, x_5862, x_5863, x_5864, x_5865, x_5866, x_5867, x_5868, x_5869, x_5870, x_5871, x_5872, x_5873, x_5874, x_5875, x_5876, x_5877, x_5878, x_5879, x_5880, x_5881, x_5882, x_5883, x_5884, x_5885, x_5886, x_5887, x_5888, x_5889, x_5890, x_5891, x_5892, x_5893, x_5894, x_5895, x_5896, x_5897, x_5898, x_5899, x_5900, x_5901, x_5902, x_5903, x_5904, x_5905, x_5906, x_5907, x_5908, x_5909, x_5910, x_5911, x_5912, x_5913, x_5914, x_5915, x_5916, x_5917, x_5918, x_5919, x_5920, x_5921, x_5922, x_5923, x_5924, x_5925, x_5926, x_5927, x_5928, x_5929, x_5930, x_5931, x_5932, x_5933, x_5934, x_5935, x_5936, x_5937, x_5938, x_5939, x_5940, x_5941, x_5942, x_5943, x_5944, x_5945, x_5946, x_5947, x_5948, x_5949, x_5950, x_5951, x_5952, x_5953, x_5954, x_5955, x_5956, x_5957, x_5958, x_5959, x_5960, x_5961, x_5962, x_5963, x_5964, x_5965, x_5966, x_5967, x_5968, x_5969, x_5970, x_5971, x_5972, x_5973, x_5974, x_5975, x_5976, x_5977, x_5978, x_5979, x_5980, x_5981, x_5982, x_5983, x_5984, x_5985, x_5986, x_5987, x_5988, x_5989, x_5990, x_5991, x_5992, x_5993, x_5994, x_5995, x_5996, x_5997, x_5998, x_5999, x_6000, x_6001, x_6002, x_6003, x_6004, x_6005, x_6006, x_6007, x_6008, x_6009, x_6010, x_6011, x_6012, x_6013, x_6014, x_6015, x_6016, x_6017, x_6018, x_6019, x_6020, x_6021, x_6022, x_6023, x_6024, x_6025, x_6026, x_6027, x_6028, x_6029, x_6030, x_6031, x_6032, x_6033, x_6034, x_6035, x_6036, x_6037, x_6038, x_6039, x_6040, x_6041, x_6042, x_6043, x_6044, x_6045, x_6046, x_6047, x_6048, x_6049, x_6050, x_6051, x_6052, x_6053, x_6054, x_6055, x_6056, x_6057, x_6058, x_6059, x_6060, x_6061, x_6062, x_6063, x_6064, x_6065, x_6066, x_6067, x_6068, x_6069, x_6070, x_6071, x_6072, x_6073, x_6074, x_6075, x_6076, x_6077, x_6078, x_6079, x_6080, x_6081, x_6082, x_6083, x_6084, x_6085, x_6086, x_6087, x_6088, x_6089, x_6090, x_6091, x_6092, x_6093, x_6094, x_6095, x_6096, x_6097, x_6098, x_6099, x_6100, x_6101, x_6102, x_6103, x_6104, x_6105, x_6106, x_6107, x_6108, x_6109, x_6110, x_6111, x_6112, x_6113, x_6114, x_6115, x_6116, x_6117, x_6118, x_6119, x_6120, x_6121, x_6122, x_6123, x_6124, x_6125, x_6126, x_6127, x_6128, x_6129, x_6130, x_6131, x_6132, x_6133, x_6134, x_6135, x_6136, x_6137, x_6138, x_6139, x_6140, x_6141, x_6142, x_6143, x_6144, x_6145, x_6146, x_6147, x_6148, x_6149, x_6150, x_6151, x_6152, x_6153, x_6154, x_6155, x_6156, x_6157, x_6158, x_6159, x_6160, x_6161, x_6162, x_6163, x_6164, x_6165, x_6166, x_6167, x_6168, x_6169, x_6170, x_6171, x_6172, x_6173, x_6174, x_6175, x_6176, x_6177, x_6178, x_6179, x_6180, x_6181, x_6182, x_6183, x_6184, x_6185, x_6186, x_6187, x_6188, x_6189, x_6190, x_6191, x_6192, x_6193, x_6194, x_6195, x_6196, x_6197, x_6198, x_6199, x_6200, x_6201, x_6202, x_6203, x_6204, x_6205, x_6206, x_6207, x_6208, x_6209, x_6210, x_6211, x_6212, x_6213, x_6214, x_6215, x_6216, x_6217, x_6218, x_6219, x_6220, x_6221, x_6222, x_6223, x_6224, x_6225, x_6226, x_6227, x_6228, x_6229, x_6230, x_6231, x_6232, x_6233, x_6234, x_6235, x_6236, x_6237, x_6238, x_6239, x_6240, x_6241, x_6242, x_6243, x_6244, x_6245, x_6246, x_6247, x_6248, x_6249, x_6250, x_6251, x_6252, x_6253, x_6254, x_6255, x_6256, x_6257, x_6258, x_6259, x_6260, x_6261, x_6262, x_6263, x_6264, x_6265, x_6266, x_6267, x_6268, x_6269, x_6270, x_6271, x_6272, x_6273, x_6274, x_6275, x_6276, x_6277, x_6278, x_6279, x_6280, x_6281, x_6282, x_6283, x_6284, x_6285, x_6286, x_6287, x_6288, x_6289, x_6290, x_6291, x_6292, x_6293, x_6294, x_6295, x_6296, x_6297, x_6298, x_6299, x_6300, x_6301, x_6302, x_6303, x_6304, x_6305, x_6306, x_6307, x_6308, x_6309, x_6310, x_6311, x_6312, x_6313, x_6314, x_6315, x_6316, x_6317, x_6318, x_6319, x_6320, x_6321, x_6322, x_6323, x_6324, x_6325, x_6326, x_6327, x_6328, x_6329, x_6330, x_6331, x_6332, x_6333, x_6334, x_6335, x_6336, x_6337, x_6338, x_6339, x_6340, x_6341, x_6342, x_6343, x_6344, x_6345, x_6346, x_6347, x_6348, x_6349, x_6350, x_6351, x_6352, x_6353, x_6354, x_6355, x_6356, x_6357, x_6358, x_6359, x_6360, x_6361, x_6362, x_6363, x_6364, x_6365, x_6366, x_6367, x_6368, x_6369, x_6370, x_6371, x_6372, x_6373, x_6374, x_6375, x_6376, x_6377, x_6378, x_6379, x_6380, x_6381, x_6382, x_6383, x_6384, x_6385, x_6386, x_6387, x_6388, x_6389, x_6390, x_6391, x_6392, x_6393, x_6394, x_6395, x_6396, x_6397, x_6398, x_6399, x_6400, x_6401, x_6402, x_6403, x_6404, x_6405, x_6406, x_6407, x_6408, x_6409, x_6410, x_6411, x_6412, x_6413, x_6414, x_6415, x_6416, x_6417, x_6418, x_6419, x_6420, x_6421, x_6422, x_6423, x_6424, x_6425, x_6426, x_6427, x_6428, x_6429, x_6430, x_6431, x_6432, x_6433, x_6434, x_6435, x_6436, x_6437, x_6438, x_6439, x_6440, x_6441, x_6442, x_6443, x_6444, x_6445, x_6446, x_6447, x_6448, x_6449, x_6450, x_6451, x_6452, x_6453, x_6454, x_6455, x_6456, x_6457, x_6458, x_6459, x_6460, x_6461, x_6462, x_6463, x_6464, x_6465, x_6466, x_6467, x_6468, x_6469, x_6470, x_6471, x_6472, x_6473, x_6474, x_6475, x_6476, x_6477, x_6478, x_6479, x_6480, x_6481, x_6482, x_6483, x_6484, x_6485, x_6486, x_6487, x_6488, x_6489, x_6490, x_6491, x_6492, x_6493, x_6494, x_6495, x_6496, x_6497, x_6498, x_6499, x_6500, x_6501, x_6502, x_6503, x_6504, x_6505, x_6506, x_6507, x_6508, x_6509, x_6510, x_6511, x_6512, x_6513, x_6514, x_6515, x_6516, x_6517, x_6518, x_6519, x_6520, x_6521, x_6522, x_6523, x_6524, x_6525, x_6526, x_6527, x_6528, x_6529, x_6530, x_6531, x_6532, x_6533, x_6534, x_6535, x_6536, x_6537, x_6538, x_6539, x_6540, x_6541, x_6542, x_6543, x_6544, x_6545, x_6546, x_6547, x_6548, x_6549, x_6550, x_6551, x_6552, x_6553, x_6554, x_6555, x_6556, x_6557, x_6558, x_6559, x_6560, x_6561, x_6562, x_6563, x_6564, x_6565, x_6566, x_6567, x_6568, x_6569, x_6570, x_6571, x_6572, x_6573, x_6574, x_6575, x_6576, x_6577, x_6578, x_6579, x_6580, x_6581, x_6582, x_6583, x_6584, x_6585, x_6586, x_6587, x_6588, x_6589, x_6590, x_6591, x_6592, x_6593, x_6594, x_6595, x_6596, x_6597, x_6598, x_6599, x_6600, x_6601, x_6602, x_6603, x_6604, x_6605, x_6606, x_6607, x_6608, x_6609, x_6610, x_6611, x_6612, x_6613, x_6614, x_6615, x_6616, x_6617, x_6618, x_6619, x_6620, x_6621, x_6622, x_6623, x_6624, x_6625, x_6626, x_6627, x_6628, x_6629, x_6630, x_6631, x_6632, x_6633, x_6634, x_6635, x_6636, x_6637, x_6638, x_6639, x_6640, x_6641, x_6642, x_6643, x_6644, x_6645, x_6646, x_6647, x_6648, x_6649, x_6650, x_6651, x_6652, x_6653, x_6654, x_6655, x_6656, x_6657, x_6658, x_6659, x_6660, x_6661, x_6662, x_6663, x_6664, x_6665, x_6666, x_6667, x_6668, x_6669, x_6670, x_6671, x_6672, x_6673, x_6674, x_6675, x_6676, x_6677, x_6678, x_6679, x_6680, x_6681, x_6682, x_6683, x_6684, x_6685, x_6686, x_6687, x_6688, x_6689, x_6690, x_6691, x_6692, x_6693, x_6694, x_6695, x_6696, x_6697, x_6698, x_6699, x_6700, x_6701, x_6702, x_6703, x_6704, x_6705, x_6706, x_6707, x_6708, x_6709, x_6710, x_6711, x_6712, x_6713, x_6714, x_6715, x_6716, x_6717, x_6718, x_6719, x_6720, x_6721, x_6722, x_6723, x_6724, x_6725, x_6726, x_6727, x_6728, x_6729, x_6730, x_6731, x_6732, x_6733, x_6734, x_6735, x_6736, x_6737, x_6738, x_6739, x_6740, x_6741, x_6742, x_6743, x_6744, x_6745, x_6746, x_6747, x_6748, x_6749, x_6750, x_6751, x_6752, x_6753, x_6754, x_6755, x_6756, x_6757, x_6758, x_6759, x_6760, x_6761, x_6762, x_6763, x_6764, x_6765, x_6766, x_6767, x_6768, x_6769, x_6770, x_6771, x_6772, x_6773, x_6774, x_6775, x_6776, x_6777, x_6778, x_6779, x_6780, x_6781, x_6782, x_6783, x_6784, x_6785, x_6786, x_6787, x_6788, x_6789, x_6790, x_6791, x_6792, x_6793, x_6794, x_6795, x_6796, x_6797, x_6798, x_6799, x_6800, x_6801, x_6802, x_6803, x_6804, x_6805, x_6806, x_6807, x_6808, x_6809, x_6810, x_6811, x_6812, x_6813, x_6814, x_6815, x_6816, x_6817, x_6818, x_6819, x_6820, x_6821, x_6822, x_6823, x_6824, x_6825, x_6826, x_6827, x_6828, x_6829, x_6830, x_6831, x_6832, x_6833, x_6834, x_6835, x_6836, x_6837, x_6838, x_6839, x_6840, x_6841, x_6842, x_6843, x_6844, x_6845, x_6846, x_6847, x_6848, x_6849, x_6850, x_6851, x_6852, x_6853, x_6854, x_6855, x_6856, x_6857, x_6858, x_6859, x_6860, x_6861, x_6862, x_6863, x_6864, x_6865, x_6866, x_6867, x_6868, x_6869, x_6870, x_6871, x_6872, x_6873, x_6874, x_6875, x_6876, x_6877, x_6878, x_6879, x_6880, x_6881, x_6882, x_6883, x_6884, x_6885, x_6886, x_6887, x_6888, x_6889, x_6890, x_6891, x_6892, x_6893, x_6894, x_6895, x_6896, x_6897, x_6898, x_6899, x_6900, x_6901, x_6902, x_6903, x_6904, x_6905, x_6906, x_6907, x_6908, x_6909, x_6910, x_6911, x_6912, x_6913, x_6914, x_6915, x_6916, x_6917, x_6918, x_6919, x_6920, x_6921, x_6922, x_6923, x_6924, x_6925, x_6926, x_6927, x_6928, x_6929, x_6930, x_6931, x_6932, x_6933, x_6934, x_6935, x_6936, x_6937, x_6938, x_6939, x_6940, x_6941, x_6942, x_6943, x_6944, x_6945, x_6946, x_6947, x_6948, x_6949, x_6950, x_6951, x_6952, x_6953, x_6954, x_6955, x_6956, x_6957, x_6958, x_6959, x_6960, x_6961, x_6962, x_6963, x_6964, x_6965, x_6966, x_6967, x_6968, x_6969, x_6970, x_6971, x_6972, x_6973, x_6974, x_6975, x_6976, x_6977, x_6978, x_6979, x_6980, x_6981, x_6982, x_6983, x_6984, x_6985, x_6986, x_6987, x_6988, x_6989, x_6990, x_6991, x_6992, x_6993, x_6994, x_6995, x_6996, x_6997, x_6998, x_6999, x_7000, x_7001, x_7002, x_7003, x_7004, x_7005, x_7006, x_7007, x_7008, x_7009, x_7010, x_7011, x_7012, x_7013, x_7014, x_7015, x_7016, x_7017, x_7018, x_7019, x_7020, x_7021, x_7022, x_7023, x_7024, x_7025, x_7026, x_7027, x_7028, x_7029, x_7030, x_7031, x_7032, x_7033, x_7034, x_7035, x_7036, x_7037, x_7038, x_7039, x_7040, x_7041, x_7042, x_7043, x_7044, x_7045, x_7046, x_7047, x_7048, x_7049, x_7050, x_7051, x_7052, x_7053, x_7054, x_7055, x_7056, x_7057, x_7058, x_7059, x_7060, x_7061, x_7062, x_7063, x_7064, x_7065, x_7066, x_7067, x_7068, x_7069, x_7070, x_7071, x_7072, x_7073, x_7074, x_7075, x_7076, x_7077, x_7078, x_7079, x_7080, x_7081, x_7082, x_7083, x_7084, x_7085, x_7086, x_7087, x_7088, x_7089, x_7090, x_7091, x_7092, x_7093, x_7094, x_7095, x_7096, x_7097, x_7098, x_7099, x_7100, x_7101, x_7102, x_7103, x_7104, x_7105, x_7106, x_7107, x_7108, x_7109, x_7110, x_7111, x_7112, x_7113, x_7114, x_7115, x_7116, x_7117, x_7118, x_7119, x_7120, x_7121, x_7122, x_7123, x_7124, x_7125, x_7126, x_7127, x_7128, x_7129, x_7130, x_7131, x_7132, x_7133, x_7134, x_7135, x_7136, x_7137, x_7138, x_7139, x_7140, x_7141, x_7142, x_7143, x_7144, x_7145, x_7146, x_7147, x_7148, x_7149, x_7150, x_7151, x_7152, x_7153, x_7154, x_7155, x_7156, x_7157, x_7158, x_7159, x_7160, x_7161, x_7162, x_7163, x_7164, x_7165, x_7166, x_7167, x_7168, x_7169, x_7170, x_7171, x_7172, x_7173, x_7174, x_7175, x_7176, x_7177, x_7178, x_7179, x_7180, x_7181, x_7182, x_7183, x_7184, x_7185, x_7186, x_7187, x_7188, x_7189, x_7190, x_7191, x_7192, x_7193, x_7194, x_7195, x_7196, x_7197, x_7198, x_7199, x_7200, x_7201, x_7202, x_7203, x_7204, x_7205, x_7206, x_7207, x_7208, x_7209, x_7210, x_7211, x_7212, x_7213, x_7214, x_7215, x_7216, x_7217, x_7218, x_7219, x_7220, x_7221, x_7222, x_7223, x_7224, x_7225, x_7226, x_7227, x_7228, x_7229, x_7230, x_7231, x_7232, x_7233, x_7234, x_7235, x_7236, x_7237, x_7238, x_7239, x_7240, x_7241, x_7242, x_7243, x_7244, x_7245, x_7246, x_7247, x_7248, x_7249, x_7250, x_7251, x_7252, x_7253, x_7254, x_7255, x_7256, x_7257, x_7258, x_7259, x_7260, x_7261, x_7262, x_7263, x_7264, x_7265, x_7266, x_7267, x_7268, x_7269, x_7270, x_7271, x_7272, x_7273, x_7274, x_7275, x_7276, x_7277, x_7278, x_7279, x_7280, x_7281, x_7282, x_7283, x_7284, x_7285, x_7286, x_7287, x_7288, x_7289, x_7290, x_7291, x_7292, x_7293, x_7294, x_7295, x_7296, x_7297, x_7298, x_7299, x_7300, x_7301, x_7302, x_7303, x_7304, x_7305, x_7306, x_7307, x_7308, x_7309, x_7310, x_7311, x_7312, x_7313, x_7314, x_7315, x_7316, x_7317, x_7318, x_7319, x_7320, x_7321, x_7322, x_7323, x_7324, x_7325, x_7326, x_7327, x_7328, x_7329, x_7330, x_7331, x_7332, x_7333, x_7334, x_7335, x_7336, x_7337, x_7338, x_7339, x_7340, x_7341, x_7342, x_7343, x_7344, x_7345, x_7346, x_7347, x_7348, x_7349, x_7350, x_7351, x_7352, x_7353, x_7354, x_7355, x_7356, x_7357, x_7358, x_7359, x_7360, x_7361, x_7362, x_7363, x_7364, x_7365, x_7366, x_7367, x_7368, x_7369, x_7370, x_7371, x_7372, x_7373, x_7374, x_7375, x_7376, x_7377, x_7378, x_7379, x_7380, x_7381, x_7382, x_7383, x_7384, x_7385, x_7386, x_7387, x_7388, x_7389, x_7390, x_7391, x_7392, x_7393, x_7394, x_7395, x_7396, x_7397, x_7398, x_7399, x_7400, x_7401, x_7402, x_7403, x_7404, x_7405, x_7406, x_7407, x_7408, x_7409, x_7410, x_7411, x_7412, x_7413, x_7414, x_7415, x_7416, x_7417, x_7418, x_7419, x_7420, x_7421, x_7422, x_7423, x_7424, x_7425, x_7426, x_7427, x_7428, x_7429, x_7430, x_7431, x_7432, x_7433, x_7434, x_7435, x_7436, x_7437, x_7438, x_7439, x_7440, x_7441, x_7442, x_7443, x_7444, x_7445, x_7446, x_7447, x_7448, x_7449, x_7450, x_7451, x_7452, x_7453, x_7454, x_7455, x_7456, x_7457, x_7458, x_7459, x_7460, x_7461, x_7462, x_7463, x_7464, x_7465, x_7466, x_7467, x_7468, x_7469, x_7470, x_7471, x_7472, x_7473, x_7474, x_7475, x_7476, x_7477, x_7478, x_7479, x_7480, x_7481, x_7482, x_7483, x_7484, x_7485, x_7486, x_7487, x_7488, x_7489, x_7490, x_7491, x_7492, x_7493, x_7494, x_7495, x_7496, x_7497, x_7498, x_7499, x_7500, x_7501, x_7502, x_7503, x_7504, x_7505, x_7506, x_7507, x_7508, x_7509, x_7510, x_7511, x_7512, x_7513, x_7514, x_7515, x_7516, x_7517, x_7518, x_7519, x_7520, x_7521, x_7522, x_7523, x_7524, x_7525, x_7526, x_7527, x_7528, x_7529, x_7530, x_7531, x_7532, x_7533, x_7534, x_7535, x_7536, x_7537, x_7538, x_7539, x_7540, x_7541, x_7542, x_7543, x_7544, x_7545, x_7546, x_7547, x_7548, x_7549, x_7550, x_7551, x_7552, x_7553, x_7554, x_7555, x_7556, x_7557, x_7558, x_7559, x_7560, x_7561, x_7562, x_7563, x_7564, x_7565, x_7566, x_7567, x_7568, x_7569, x_7570, x_7571, x_7572, x_7573, x_7574, x_7575, x_7576, x_7577, x_7578, x_7579, x_7580, x_7581, x_7582, x_7583, x_7584, x_7585, x_7586, x_7587, x_7588, x_7589, x_7590, x_7591, x_7592, x_7593, x_7594, x_7595, x_7596, x_7597, x_7598, x_7599, x_7600, x_7601, x_7602, x_7603, x_7604, x_7605, x_7606, x_7607, x_7608, x_7609, x_7610, x_7611, x_7612, x_7613, x_7614, x_7615, x_7616, x_7617, x_7618, x_7619, x_7620, x_7621, x_7622, x_7623, x_7624, x_7625, x_7626, x_7627, x_7628, x_7629, x_7630, x_7631, x_7632, x_7633, x_7634, x_7635, x_7636, x_7637, x_7638, x_7639, x_7640, x_7641, x_7642, x_7643, x_7644, x_7645, x_7646, x_7647, x_7648, x_7649, x_7650, x_7651, x_7652, x_7653, x_7654, x_7655, x_7656, x_7657, x_7658, x_7659, x_7660, x_7661, x_7662, x_7663, x_7664, x_7665, x_7666, x_7667, x_7668, x_7669, x_7670, x_7671, x_7672, x_7673, x_7674, x_7675, x_7676, x_7677, x_7678, x_7679, x_7680, x_7681, x_7682, x_7683, x_7684, x_7685, x_7686, x_7687, x_7688, x_7689, x_7690, x_7691, x_7692, x_7693, x_7694, x_7695, x_7696, x_7697, x_7698, x_7699, x_7700, x_7701, x_7702, x_7703, x_7704, x_7705, x_7706, x_7707, x_7708, x_7709, x_7710, x_7711, x_7712, x_7713, x_7714, x_7715, x_7716, x_7717, x_7718, x_7719, x_7720, x_7721, x_7722, x_7723, x_7724, x_7725, x_7726, x_7727, x_7728, x_7729, x_7730, x_7731, x_7732, x_7733, x_7734, x_7735, x_7736, x_7737, x_7738, x_7739, x_7740, x_7741, x_7742, x_7743, x_7744, x_7745, x_7746, x_7747, x_7748, x_7749, x_7750, x_7751, x_7752, x_7753, x_7754, x_7755, x_7756, x_7757, x_7758, x_7759, x_7760, x_7761, x_7762, x_7763, x_7764, x_7765, x_7766, x_7767, x_7768, x_7769, x_7770, x_7771, x_7772, x_7773, x_7774, x_7775, x_7776, x_7777, x_7778, x_7779, x_7780, x_7781, x_7782, x_7783, x_7784, x_7785, x_7786, x_7787, x_7788, x_7789, x_7790, x_7791, x_7792, x_7793, x_7794, x_7795, x_7796, x_7797, x_7798, x_7799, x_7800, x_7801, x_7802, x_7803, x_7804, x_7805, x_7806, x_7807, x_7808, x_7809, x_7810, x_7811, x_7812, x_7813, x_7814, x_7815, x_7816, x_7817, x_7818, x_7819, x_7820, x_7821, x_7822, x_7823, x_7824, x_7825, x_7826, x_7827, x_7828, x_7829, x_7830, x_7831, x_7832, x_7833, x_7834, x_7835, x_7836, x_7837, x_7838, x_7839, x_7840, x_7841, x_7842, x_7843, x_7844, x_7845, x_7846, x_7847, x_7848, x_7849, x_7850, x_7851, x_7852, x_7853, x_7854, x_7855, x_7856, x_7857, x_7858, x_7859, x_7860, x_7861, x_7862, x_7863, x_7864, x_7865, x_7866, x_7867, x_7868, x_7869, x_7870, x_7871, x_7872, x_7873, x_7874, x_7875, x_7876, x_7877, x_7878, x_7879, x_7880, x_7881, x_7882, x_7883, x_7884, x_7885, x_7886, x_7887, x_7888, x_7889, x_7890, x_7891, x_7892, x_7893, x_7894, x_7895, x_7896, x_7897, x_7898, x_7899, x_7900, x_7901, x_7902, x_7903, x_7904, x_7905, x_7906, x_7907, x_7908, x_7909, x_7910, x_7911, x_7912, x_7913, x_7914, x_7915, x_7916, x_7917, x_7918, x_7919, x_7920, x_7921, x_7922, x_7923, x_7924, x_7925, x_7926, x_7927, x_7928, x_7929, x_7930, x_7931, x_7932, x_7933, x_7934, x_7935, x_7936, x_7937, x_7938, x_7939, x_7940, x_7941, x_7942, x_7943, x_7944, x_7945, x_7946, x_7947, x_7948, x_7949, x_7950, x_7951, x_7952, x_7953, x_7954, x_7955, x_7956, x_7957, x_7958, x_7959, x_7960, x_7961, x_7962, x_7963, x_7964, x_7965, x_7966, x_7967, x_7968, x_7969, x_7970, x_7971, x_7972, x_7973, x_7974, x_7975, x_7976, x_7977, x_7978, x_7979, x_7980, x_7981, x_7982, x_7983, x_7984, x_7985, x_7986, x_7987, x_7988, x_7989, x_7990, x_7991, x_7992, x_7993, x_7994, x_7995, x_7996, x_7997, x_7998, x_7999, x_8000, x_8001, x_8002, x_8003, x_8004, x_8005, x_8006, x_8007, x_8008, x_8009, x_8010, x_8011, x_8012, x_8013, x_8014, x_8015, x_8016, x_8017, x_8018, x_8019, x_8020, x_8021, x_8022, x_8023, x_8024, x_8025, x_8026, x_8027, x_8028, x_8029, x_8030, x_8031, x_8032, x_8033, x_8034, x_8035, x_8036, x_8037, x_8038, x_8039, x_8040, x_8041, x_8042, x_8043, x_8044, x_8045, x_8046, x_8047, x_8048, x_8049, x_8050, x_8051, x_8052, x_8053, x_8054, x_8055, x_8056, x_8057, x_8058, x_8059, x_8060, x_8061, x_8062, x_8063, x_8064, x_8065, x_8066, x_8067, x_8068, x_8069, x_8070, x_8071, x_8072, x_8073, x_8074, x_8075, x_8076, x_8077, x_8078, x_8079, x_8080, x_8081, x_8082, x_8083, x_8084, x_8085, x_8086, x_8087, x_8088, x_8089, x_8090, x_8091, x_8092, x_8093, x_8094, x_8095, x_8096, x_8097, x_8098, x_8099, x_8100, x_8101, x_8102, x_8103, x_8104, x_8105, x_8106, x_8107, x_8108, x_8109, x_8110, x_8111, x_8112, x_8113, x_8114, x_8115, x_8116, x_8117, x_8118, x_8119, x_8120, x_8121, x_8122, x_8123, x_8124, x_8125, x_8126, x_8127, x_8128, x_8129, x_8130, x_8131, x_8132, x_8133, x_8134, x_8135, x_8136, x_8137, x_8138, x_8139, x_8140, x_8141, x_8142, x_8143, x_8144, x_8145, x_8146, x_8147, x_8148, x_8149, x_8150, x_8151, x_8152, x_8153, x_8154, x_8155, x_8156, x_8157, x_8158, x_8159, x_8160, x_8161, x_8162, x_8163, x_8164, x_8165, x_8166, x_8167, x_8168, x_8169, x_8170, x_8171, x_8172, x_8173, x_8174, x_8175, x_8176, x_8177, x_8178, x_8179, x_8180, x_8181, x_8182, x_8183, x_8184, x_8185, x_8186, x_8187, x_8188, x_8189, x_8190, x_8191, x_8192, x_8193, x_8194, x_8195, x_8196, x_8197, x_8198, x_8199, x_8200, x_8201, x_8202, x_8203, x_8204, x_8205, x_8206, x_8207, x_8208, x_8209, x_8210, x_8211, x_8212, x_8213, x_8214, x_8215, x_8216, x_8217, x_8218, x_8219, x_8220, x_8221, x_8222, x_8223, x_8224, x_8225, x_8226, x_8227, x_8228, x_8229, x_8230, x_8231, x_8232, x_8233, x_8234, x_8235, x_8236, x_8237, x_8238, x_8239, x_8240, x_8241, x_8242, x_8243, x_8244, x_8245, x_8246, x_8247, x_8248, x_8249, x_8250, x_8251, x_8252, x_8253, x_8254, x_8255, x_8256, x_8257, x_8258, x_8259, x_8260, x_8261, x_8262, x_8263, x_8264, x_8265, x_8266, x_8267, x_8268, x_8269, x_8270, x_8271, x_8272, x_8273, x_8274, x_8275, x_8276, x_8277, x_8278, x_8279, x_8280, x_8281, x_8282, x_8283, x_8284, x_8285, x_8286, x_8287, x_8288, x_8289, x_8290, x_8291, x_8292, x_8293, x_8294, x_8295, x_8296, x_8297, x_8298, x_8299, x_8300, x_8301, x_8302, x_8303, x_8304, x_8305, x_8306, x_8307, x_8308, x_8309, x_8310, x_8311, x_8312, x_8313, x_8314, x_8315, x_8316, x_8317, x_8318, x_8319, x_8320, x_8321, x_8322, x_8323, x_8324, x_8325, x_8326, x_8327, x_8328, x_8329, x_8330, x_8331, x_8332, x_8333, x_8334, x_8335, x_8336, x_8337, x_8338, x_8339, x_8340, x_8341, x_8342, x_8343, x_8344, x_8345, x_8346, x_8347, x_8348, x_8349, x_8350, x_8351, x_8352, x_8353, x_8354, x_8355, x_8356, x_8357, x_8358, x_8359, x_8360, x_8361, x_8362, x_8363, x_8364, x_8365, x_8366, x_8367, x_8368, x_8369, x_8370, x_8371, x_8372, x_8373, x_8374, x_8375, x_8376, x_8377, x_8378, x_8379, x_8380, x_8381, x_8382, x_8383, x_8384, x_8385, x_8386, x_8387, x_8388, x_8389, x_8390, x_8391, x_8392, x_8393, x_8394, x_8395, x_8396, x_8397, x_8398, x_8399, x_8400, x_8401, x_8402, x_8403, x_8404, x_8405, x_8406, x_8407, x_8408, x_8409, x_8410, x_8411, x_8412, x_8413, x_8414, x_8415, x_8416, x_8417, x_8418, x_8419, x_8420, x_8421, x_8422, x_8423, x_8424, x_8425, x_8426, x_8427, x_8428, x_8429, x_8430, x_8431, x_8432, x_8433, x_8434, x_8435, x_8436, x_8437, x_8438, x_8439, x_8440, x_8441, x_8442, x_8443, x_8444, x_8445, x_8446, x_8447, x_8448, x_8449, x_8450, x_8451, x_8452, x_8453, x_8454, x_8455, x_8456, x_8457, x_8458, x_8459, x_8460, x_8461, x_8462, x_8463, x_8464, x_8465, x_8466, x_8467, x_8468, x_8469, x_8470, x_8471, x_8472, x_8473, x_8474, x_8475, x_8476, x_8477, x_8478, x_8479, x_8480, x_8481, x_8482, x_8483, x_8484, x_8485, x_8486, x_8487, x_8488, x_8489, x_8490, x_8491, x_8492, x_8493, x_8494, x_8495, x_8496, x_8497, x_8498, x_8499, x_8500, x_8501, x_8502, x_8503, x_8504, x_8505, x_8506, x_8507, x_8508, x_8509, x_8510, x_8511, x_8512, x_8513, x_8514, x_8515, x_8516, x_8517, x_8518, x_8519, x_8520, x_8521, x_8522, x_8523, x_8524, x_8525, x_8526, x_8527, x_8528, x_8529, x_8530, x_8531, x_8532, x_8533, x_8534, x_8535, x_8536, x_8537, x_8538, x_8539, x_8540, x_8541, x_8542, x_8543, x_8544, x_8545, x_8546, x_8547, x_8548, x_8549, x_8550, x_8551, x_8552, x_8553, x_8554, x_8555, x_8556, x_8557, x_8558, x_8559, x_8560, x_8561, x_8562, x_8563, x_8564, x_8565, x_8566, x_8567, x_8568, x_8569, x_8570, x_8571, x_8572, x_8573, x_8574, x_8575, x_8576, x_8577, x_8578, x_8579, x_8580, x_8581, x_8582, x_8583, x_8584, x_8585, x_8586, x_8587, x_8588, x_8589, x_8590, x_8591, x_8592, x_8593, x_8594, x_8595, x_8596, x_8597, x_8598, x_8599, x_8600, x_8601, x_8602, x_8603, x_8604, x_8605, x_8606, x_8607, x_8608, x_8609, x_8610, x_8611, x_8612, x_8613, x_8614, x_8615, x_8616, x_8617, x_8618, x_8619, x_8620, x_8621, x_8622, x_8623, x_8624, x_8625, x_8626, x_8627, x_8628, x_8629, x_8630, x_8631, x_8632, x_8633, x_8634, x_8635, x_8636, x_8637, x_8638, x_8639, x_8640, x_8641, x_8642, x_8643, x_8644, x_8645, x_8646, x_8647, x_8648, x_8649, x_8650, x_8651, x_8652, x_8653, x_8654, x_8655, x_8656, x_8657, x_8658, x_8659, x_8660, x_8661, x_8662, x_8663, x_8664, x_8665, x_8666, x_8667, x_8668, x_8669, x_8670, x_8671, x_8672, x_8673, x_8674, x_8675, x_8676, x_8677, x_8678, x_8679, x_8680, x_8681, x_8682, x_8683, x_8684, x_8685, x_8686, x_8687, x_8688, x_8689, x_8690, x_8691, x_8692, x_8693, x_8694, x_8695, x_8696, x_8697, x_8698, x_8699, x_8700, x_8701, x_8702, x_8703, x_8704, x_8705, x_8706, x_8707, x_8708, x_8709, x_8710, x_8711, x_8712, x_8713, x_8714, x_8715, x_8716, x_8717, x_8718, x_8719, x_8720, x_8721, x_8722, x_8723, x_8724, x_8725, x_8726, x_8727, x_8728, x_8729, x_8730, x_8731, x_8732, x_8733, x_8734, x_8735, x_8736, x_8737, x_8738, x_8739, x_8740, x_8741, x_8742, x_8743, x_8744, x_8745, x_8746, x_8747, x_8748, x_8749, x_8750, x_8751, x_8752, x_8753, x_8754, x_8755, x_8756, x_8757, x_8758, x_8759, x_8760, x_8761, x_8762, x_8763, x_8764, x_8765, x_8766, x_8767, x_8768, x_8769, x_8770, x_8771, x_8772, x_8773, x_8774, x_8775, x_8776, x_8777, x_8778, x_8779, x_8780, x_8781, x_8782, x_8783, x_8784, x_8785, x_8786, x_8787, x_8788, x_8789, x_8790, x_8791, x_8792, x_8793, x_8794, x_8795, x_8796, x_8797, x_8798, x_8799, x_8800, x_8801, x_8802, x_8803, x_8804, x_8805, x_8806, x_8807, x_8808, x_8809, x_8810, x_8811, x_8812, x_8813, x_8814, x_8815, x_8816, x_8817, x_8818, x_8819, x_8820, x_8821, x_8822, x_8823, x_8824, x_8825, x_8826, x_8827, x_8828, x_8829, x_8830, x_8831, x_8832, x_8833, x_8834, x_8835, x_8836, x_8837, x_8838, x_8839, x_8840, x_8841, x_8842, x_8843, x_8844, x_8845, x_8846, x_8847, x_8848, x_8849, x_8850, x_8851, x_8852, x_8853, x_8854, x_8855, x_8856, x_8857, x_8858, x_8859, x_8860, x_8861, x_8862, x_8863, x_8864, x_8865, x_8866, x_8867, x_8868, x_8869, x_8870, x_8871, x_8872, x_8873, x_8874, x_8875, x_8876, x_8877, x_8878, x_8879, x_8880, x_8881, x_8882, x_8883, x_8884, x_8885, x_8886, x_8887, x_8888, x_8889, x_8890, x_8891, x_8892, x_8893, x_8894, x_8895, x_8896, x_8897, x_8898, x_8899, x_8900, x_8901, x_8902, x_8903, x_8904, x_8905, x_8906, x_8907, x_8908, x_8909, x_8910, x_8911, x_8912, x_8913, x_8914, x_8915, x_8916, x_8917, x_8918, x_8919, x_8920, x_8921, x_8922, x_8923, x_8924, x_8925, x_8926, x_8927, x_8928, x_8929, x_8930, x_8931, x_8932, x_8933, x_8934, x_8935, x_8936, x_8937, x_8938, x_8939, x_8940, x_8941, x_8942, x_8943, x_8944, x_8945, x_8946, x_8947, x_8948, x_8949, x_8950, x_8951, x_8952, x_8953, x_8954, x_8955, x_8956, x_8957, x_8958, x_8959, x_8960, x_8961, x_8962, x_8963, x_8964, x_8965, x_8966, x_8967, x_8968, x_8969, x_8970, x_8971, x_8972, x_8973, x_8974, x_8975, x_8976, x_8977, x_8978, x_8979, x_8980, x_8981, x_8982, x_8983, x_8984, x_8985, x_8986, x_8987, x_8988, x_8989, x_8990, x_8991, x_8992, x_8993, x_8994, x_8995, x_8996, x_8997, x_8998, x_8999, x_9000, x_9001, x_9002, x_9003, x_9004, x_9005, x_9006, x_9007, x_9008, x_9009, x_9010, x_9011, x_9012, x_9013, x_9014, x_9015, x_9016, x_9017, x_9018, x_9019, x_9020, x_9021, x_9022, x_9023, x_9024, x_9025, x_9026, x_9027, x_9028, x_9029, x_9030, x_9031, x_9032, x_9033, x_9034, x_9035, x_9036, x_9037, x_9038, x_9039, x_9040, x_9041, x_9042, x_9043, x_9044, x_9045, x_9046, x_9047, x_9048, x_9049, x_9050, x_9051, x_9052, x_9053, x_9054, x_9055, x_9056, x_9057, x_9058, x_9059, x_9060, x_9061, x_9062, x_9063, x_9064, x_9065, x_9066, x_9067, x_9068, x_9069, x_9070, x_9071, x_9072, x_9073, x_9074, x_9075, x_9076, x_9077, x_9078, x_9079, x_9080, x_9081, x_9082, x_9083, x_9084, x_9085, x_9086, x_9087, x_9088, x_9089, x_9090, x_9091, x_9092, x_9093, x_9094, x_9095, x_9096, x_9097, x_9098, x_9099, x_9100, x_9101, x_9102, x_9103, x_9104, x_9105, x_9106, x_9107, x_9108, x_9109, x_9110, x_9111, x_9112, x_9113, x_9114, x_9115, x_9116, x_9117, x_9118, x_9119, x_9120, x_9121, x_9122, x_9123, x_9124, x_9125, x_9126, x_9127, x_9128, x_9129, x_9130, x_9131, x_9132, x_9133, x_9134, x_9135, x_9136, x_9137, x_9138, x_9139, x_9140, x_9141, x_9142, x_9143, x_9144, x_9145, x_9146, x_9147, x_9148, x_9149, x_9150, x_9151, x_9152, x_9153, x_9154, x_9155, x_9156, x_9157, x_9158, x_9159, x_9160, x_9161, x_9162, x_9163, x_9164, x_9165, x_9166, x_9167, x_9168, x_9169, x_9170, x_9171, x_9172, x_9173, x_9174, x_9175, x_9176, x_9177, x_9178, x_9179, x_9180, x_9181, x_9182, x_9183, x_9184, x_9185, x_9186, x_9187, x_9188, x_9189, x_9190, x_9191, x_9192, x_9193, x_9194, x_9195, x_9196, x_9197, x_9198, x_9199, x_9200, x_9201, x_9202, x_9203, x_9204, x_9205, x_9206, x_9207, x_9208, x_9209, x_9210, x_9211, x_9212, x_9213, x_9214, x_9215, x_9216, x_9217, x_9218, x_9219, x_9220, x_9221, x_9222, x_9223, x_9224, x_9225, x_9226, x_9227, x_9228, x_9229, x_9230, x_9231, x_9232, x_9233, x_9234, x_9235, x_9236, x_9237, x_9238, x_9239, x_9240, x_9241, x_9242, x_9243, x_9244, x_9245, x_9246, x_9247, x_9248, x_9249, x_9250, x_9251, x_9252, x_9253, x_9254, x_9255, x_9256, x_9257, x_9258, x_9259, x_9260, x_9261, x_9262, x_9263, x_9264, x_9265, x_9266, x_9267, x_9268, x_9269, x_9270, x_9271, x_9272, x_9273, x_9274, x_9275, x_9276, x_9277, x_9278, x_9279, x_9280, x_9281, x_9282, x_9283, x_9284, x_9285, x_9286, x_9287, x_9288, x_9289, x_9290, x_9291, x_9292, x_9293, x_9294, x_9295, x_9296, x_9297, x_9298, x_9299, x_9300, x_9301, x_9302, x_9303, x_9304, x_9305, x_9306, x_9307, x_9308, x_9309, x_9310, x_9311, x_9312, x_9313, x_9314, x_9315, x_9316, x_9317, x_9318, x_9319, x_9320, x_9321, x_9322, x_9323, x_9324, x_9325, x_9326, x_9327, x_9328, x_9329, x_9330, x_9331, x_9332, x_9333, x_9334, x_9335, x_9336, x_9337, x_9338, x_9339, x_9340, x_9341, x_9342, x_9343, x_9344, x_9345, x_9346, x_9347, x_9348, x_9349, x_9350, x_9351, x_9352, x_9353, x_9354, x_9355, x_9356, x_9357, x_9358, x_9359, x_9360, x_9361, x_9362, x_9363, x_9364, x_9365, x_9366, x_9367, x_9368, x_9369, x_9370, x_9371, x_9372, x_9373, x_9374, x_9375, x_9376, x_9377, x_9378, x_9379, x_9380, x_9381, x_9382, x_9383, x_9384, x_9385, x_9386, x_9387, x_9388, x_9389, x_9390, x_9391, x_9392, x_9393, x_9394, x_9395, x_9396, x_9397, x_9398, x_9399, x_9400, x_9401, x_9402, x_9403, x_9404, x_9405, x_9406, x_9407, x_9408, x_9409, x_9410, x_9411, x_9412, x_9413, x_9414, x_9415, x_9416, x_9417, x_9418, x_9419, x_9420, x_9421, x_9422, x_9423, x_9424, x_9425, x_9426, x_9427, x_9428, x_9429, x_9430, x_9431, x_9432, x_9433, x_9434, x_9435, x_9436, x_9437, x_9438, x_9439, x_9440, x_9441, x_9442, x_9443, x_9444, x_9445, x_9446, x_9447, x_9448, x_9449, x_9450, x_9451, x_9452, x_9453, x_9454, x_9455, x_9456, x_9457, x_9458, x_9459, x_9460, x_9461, x_9462, x_9463, x_9464, x_9465, x_9466, x_9467, x_9468, x_9469, x_9470, x_9471, x_9472, x_9473, x_9474, x_9475, x_9476, x_9477, x_9478, x_9479, x_9480, x_9481, x_9482, x_9483, x_9484, x_9485, x_9486, x_9487, x_9488, x_9489, x_9490, x_9491, x_9492, x_9493, x_9494, x_9495, x_9496, x_9497, x_9498, x_9499, x_9500, x_9501, x_9502, x_9503, x_9504, x_9505, x_9506, x_9507, x_9508, x_9509, x_9510, x_9511, x_9512, x_9513, x_9514, x_9515, x_9516, x_9517, x_9518, x_9519, x_9520, x_9521, x_9522, x_9523, x_9524, x_9525, x_9526, x_9527, x_9528, x_9529, x_9530, x_9531, x_9532, x_9533, x_9534, x_9535, x_9536, x_9537, x_9538, x_9539, x_9540, x_9541, x_9542, x_9543, x_9544, x_9545, x_9546, x_9547, x_9548, x_9549, x_9550, x_9551, x_9552, x_9553, x_9554, x_9555, x_9556, x_9557, x_9558, x_9559, x_9560, x_9561, x_9562, x_9563, x_9564, x_9565, x_9566, x_9567, x_9568, x_9569, x_9570, x_9571, x_9572, x_9573, x_9574, x_9575, x_9576, x_9577, x_9578, x_9579, x_9580, x_9581, x_9582, x_9583, x_9584, x_9585, x_9586, x_9587, x_9588, x_9589, x_9590, x_9591, x_9592, x_9593, x_9594, x_9595, x_9596, x_9597, x_9598, x_9599, x_9600, x_9601, x_9602, x_9603, x_9604, x_9605, x_9606, x_9607, x_9608, x_9609, x_9610, x_9611, x_9612, x_9613, x_9614, x_9615, x_9616, x_9617, x_9618, x_9619, x_9620, x_9621, x_9622, x_9623, x_9624, x_9625, x_9626, x_9627, x_9628, x_9629, x_9630, x_9631, x_9632, x_9633, x_9634, x_9635, x_9636, x_9637, x_9638, x_9639, x_9640, x_9641, x_9642, x_9643, x_9644, x_9645, x_9646, x_9647, x_9648, x_9649, x_9650, x_9651, x_9652, x_9653, x_9654, x_9655, x_9656, x_9657, x_9658, x_9659, x_9660, x_9661, x_9662, x_9663, x_9664, x_9665, x_9666, x_9667, x_9668, x_9669, x_9670, x_9671, x_9672, x_9673, x_9674, x_9675, x_9676, x_9677, x_9678, x_9679, x_9680, x_9681, x_9682, x_9683, x_9684, x_9685, x_9686, x_9687, x_9688, x_9689, x_9690, x_9691, x_9692, x_9693, x_9694, x_9695, x_9696, x_9697, x_9698, x_9699, x_9700, x_9701, x_9702, x_9703, x_9704, x_9705, x_9706, x_9707, x_9708, x_9709, x_9710, x_9711, x_9712, x_9713, x_9714, x_9715, x_9716, x_9717, x_9718, x_9719, x_9720, x_9721, x_9722, x_9723, x_9724, x_9725, x_9726, x_9727, x_9728, x_9729, x_9730, x_9731, x_9732, x_9733, x_9734, x_9735, x_9736, x_9737, x_9738, x_9739, x_9740, x_9741, x_9742, x_9743, x_9744, x_9745, x_9746, x_9747, x_9748, x_9749, x_9750, x_9751, x_9752, x_9753, x_9754, x_9755, x_9756, x_9757, x_9758, x_9759, x_9760, x_9761, x_9762, x_9763, x_9764, x_9765, x_9766, x_9767, x_9768, x_9769, x_9770, x_9771, x_9772, x_9773, x_9774, x_9775, x_9776, x_9777, x_9778, x_9779, x_9780, x_9781, x_9782, x_9783, x_9784, x_9785, x_9786, x_9787, x_9788, x_9789, x_9790, x_9791, x_9792, x_9793, x_9794, x_9795, x_9796, x_9797, x_9798, x_9799, x_9800, x_9801, x_9802, x_9803, x_9804, x_9805, x_9806, x_9807, x_9808, x_9809, x_9810, x_9811, x_9812, x_9813, x_9814, x_9815, x_9816, x_9817, x_9818, x_9819, x_9820, x_9821, x_9822, x_9823, x_9824, x_9825, x_9826, x_9827, x_9828, x_9829, x_9830, x_9831, x_9832, x_9833, x_9834, x_9835, x_9836, x_9837, x_9838, x_9839, x_9840, x_9841, x_9842, x_9843, x_9844, x_9845, x_9846, x_9847, x_9848, x_9849, x_9850, x_9851, x_9852, x_9853, x_9854, x_9855, x_9856, x_9857, x_9858, x_9859, x_9860, x_9861, x_9862, x_9863, x_9864, x_9865, x_9866, x_9867, x_9868, x_9869, x_9870, x_9871, x_9872, x_9873, x_9874, x_9875, x_9876, x_9877, x_9878, x_9879, x_9880, x_9881, x_9882, x_9883, x_9884, x_9885, x_9886, x_9887, x_9888, x_9889, x_9890, x_9891, x_9892, x_9893, x_9894, x_9895, x_9896, x_9897, x_9898, x_9899, x_9900, x_9901, x_9902, x_9903, x_9904, x_9905, x_9906, x_9907, x_9908, x_9909, x_9910, x_9911, x_9912, x_9913, x_9914, x_9915, x_9916, x_9917, x_9918, x_9919, x_9920, x_9921, x_9922, x_9923, x_9924, x_9925, x_9926, x_9927, x_9928, x_9929, x_9930, x_9931, x_9932, x_9933, x_9934, x_9935, x_9936, x_9937, x_9938, x_9939, x_9940, x_9941, x_9942, x_9943, x_9944, x_9945, x_9946, x_9947, x_9948, x_9949, x_9950, x_9951, x_9952, x_9953, x_9954, x_9955, x_9956, x_9957, x_9958, x_9959, x_9960, x_9961, x_9962, x_9963, x_9964, x_9965, x_9966, x_9967, x_9968, x_9969, x_9970, x_9971, x_9972, x_9973, x_9974, x_9975, x_9976, x_9977, x_9978, x_9979, x_9980, x_9981, x_9982, x_9983, x_9984, x_9985, x_9986, x_9987, x_9988, x_9989, x_9990, x_9991, x_9992, x_9993, x_9994, x_9995, x_9996, x_9997, x_9998, x_9999, x_10000, x_10001, x_10002, x_10003, x_10004, x_10005, x_10006, x_10007, x_10008, x_10009, x_10010, x_10011, x_10012, x_10013, x_10014, x_10015, x_10016, x_10017, x_10018, x_10019, x_10020, x_10021, x_10022, x_10023, x_10024, x_10025, x_10026, x_10027, x_10028, x_10029, x_10030, x_10031, x_10032, x_10033, x_10034, x_10035, x_10036, x_10037, x_10038, x_10039, x_10040, x_10041, x_10042, x_10043, x_10044, x_10045, x_10046, x_10047, x_10048, x_10049, x_10050, x_10051, x_10052, x_10053, x_10054, x_10055, x_10056, x_10057, x_10058, x_10059, x_10060, x_10061, x_10062, x_10063, x_10064, x_10065, x_10066, x_10067, x_10068, x_10069, x_10070, x_10071, x_10072, x_10073, x_10074, x_10075, x_10076, x_10077, x_10078, x_10079, x_10080, x_10081, x_10082, x_10083, x_10084, x_10085, x_10086, x_10087, x_10088, x_10089, x_10090, x_10091, x_10092, x_10093, x_10094, o_1 );
input i_1;
input i_2;
input i_3;
input i_4;
input i_5;
input i_6;
input i_7;
input i_8;
input i_9;
input i_10;
input i_11;
input i_12;
input i_13;
input i_14;
input i_15;
input i_16;
input i_17;
input i_18;
input i_19;
input i_20;
input i_21;
input i_22;
input i_23;
input i_24;
input i_25;
input i_26;
input i_27;
input i_28;
input i_29;
input i_30;
input i_31;
input i_32;
input x_33;
input x_34;
input x_35;
input x_36;
input x_37;
input x_38;
input x_39;
input x_40;
input x_41;
input x_42;
input x_43;
input x_44;
input x_45;
input x_46;
input x_47;
input x_48;
input x_49;
input x_50;
input x_51;
input x_52;
input x_53;
input x_54;
input x_55;
input x_56;
input x_57;
input x_58;
input x_59;
input x_60;
input x_61;
input x_62;
input x_63;
input x_64;
input x_65;
input x_66;
input x_67;
input x_68;
input x_69;
input x_70;
input x_71;
input x_72;
input x_73;
input x_74;
input x_75;
input x_76;
input x_77;
input x_78;
input x_79;
input x_80;
input x_81;
input x_82;
input x_83;
input x_84;
input x_85;
input x_86;
input x_87;
input x_88;
input x_89;
input x_90;
input x_91;
input x_92;
input x_93;
input x_94;
input x_95;
input x_96;
input x_97;
input x_98;
input x_99;
input x_100;
input x_101;
input x_102;
input x_103;
input x_104;
input x_105;
input x_106;
input x_107;
input x_108;
input x_109;
input x_110;
input x_111;
input x_112;
input x_113;
input x_114;
input x_115;
input x_116;
input x_117;
input x_118;
input x_119;
input x_120;
input x_121;
input x_122;
input x_123;
input x_124;
input x_125;
input x_126;
input x_127;
input x_128;
input x_129;
input x_130;
input x_131;
input x_132;
input x_133;
input x_134;
input x_135;
input x_136;
input x_137;
input x_138;
input x_139;
input x_140;
input x_141;
input x_142;
input x_143;
input x_144;
input x_145;
input x_146;
input x_147;
input x_148;
input x_149;
input x_150;
input x_151;
input x_152;
input x_153;
input x_154;
input x_155;
input x_156;
input x_157;
input x_158;
input x_159;
input x_160;
input x_161;
input x_162;
input x_163;
input x_164;
input x_165;
input x_166;
input x_167;
input x_168;
input x_169;
input x_170;
input x_171;
input x_172;
input x_173;
input x_174;
input x_175;
input x_176;
input x_177;
input x_178;
input x_179;
input x_180;
input x_181;
input x_182;
input x_183;
input x_184;
input x_185;
input x_186;
input x_187;
input x_188;
input x_189;
input x_190;
input x_191;
input x_192;
input x_193;
input x_194;
input x_195;
input x_196;
input x_197;
input x_198;
input x_199;
input x_200;
input x_201;
input x_202;
input x_203;
input x_204;
input x_205;
input x_206;
input x_207;
input x_208;
input x_209;
input x_210;
input x_211;
input x_212;
input x_213;
input x_214;
input x_215;
input x_216;
input x_217;
input x_218;
input x_219;
input x_220;
input x_221;
input x_222;
input x_223;
input x_224;
input x_225;
input x_226;
input x_227;
input x_228;
input x_229;
input x_230;
input x_231;
input x_232;
input x_233;
input x_234;
input x_235;
input x_236;
input x_237;
input x_238;
input x_239;
input x_240;
input x_241;
input x_242;
input x_243;
input x_244;
input x_245;
input x_246;
input x_247;
input x_248;
input x_249;
input x_250;
input x_251;
input x_252;
input x_253;
input x_254;
input x_255;
input x_256;
input x_257;
input x_258;
input x_259;
input x_260;
input x_261;
input x_262;
input x_263;
input x_264;
input x_265;
input x_266;
input x_267;
input x_268;
input x_269;
input x_270;
input x_271;
input x_272;
input x_273;
input x_274;
input x_275;
input x_276;
input x_277;
input x_278;
input x_279;
input x_280;
input x_281;
input x_282;
input x_283;
input x_284;
input x_285;
input x_286;
input x_287;
input x_288;
input x_289;
input x_290;
input x_291;
input x_292;
input x_293;
input x_294;
input x_295;
input x_296;
input x_297;
input x_298;
input x_299;
input x_300;
input x_301;
input x_302;
input x_303;
input x_304;
input x_305;
input x_306;
input x_307;
input x_308;
input x_309;
input x_310;
input x_311;
input x_312;
input x_313;
input x_314;
input x_315;
input x_316;
input x_317;
input x_318;
input x_319;
input x_320;
input x_321;
input x_322;
input x_323;
input x_324;
input x_325;
input x_326;
input x_327;
input x_328;
input x_329;
input x_330;
input x_331;
input x_332;
input x_333;
input x_334;
input x_335;
input x_336;
input x_337;
input x_338;
input x_339;
input x_340;
input x_341;
input x_342;
input x_343;
input x_344;
input x_345;
input x_346;
input x_347;
input x_348;
input x_349;
input x_350;
input x_351;
input x_352;
input x_353;
input x_354;
input x_355;
input x_356;
input x_357;
input x_358;
input x_359;
input x_360;
input x_361;
input x_362;
input x_363;
input x_364;
input x_365;
input x_366;
input x_367;
input x_368;
input x_369;
input x_370;
input x_371;
input x_372;
input x_373;
input x_374;
input x_375;
input x_376;
input x_377;
input x_378;
input x_379;
input x_380;
input x_381;
input x_382;
input x_383;
input x_384;
input x_385;
input x_386;
input x_387;
input x_388;
input x_389;
input x_390;
input x_391;
input x_392;
input x_393;
input x_394;
input x_395;
input x_396;
input x_397;
input x_398;
input x_399;
input x_400;
input x_401;
input x_402;
input x_403;
input x_404;
input x_405;
input x_406;
input x_407;
input x_408;
input x_409;
input x_410;
input x_411;
input x_412;
input x_413;
input x_414;
input x_415;
input x_416;
input x_417;
input x_418;
input x_419;
input x_420;
input x_421;
input x_422;
input x_423;
input x_424;
input x_425;
input x_426;
input x_427;
input x_428;
input x_429;
input x_430;
input x_431;
input x_432;
input x_433;
input x_434;
input x_435;
input x_436;
input x_437;
input x_438;
input x_439;
input x_440;
input x_441;
input x_442;
input x_443;
input x_444;
input x_445;
input x_446;
input x_447;
input x_448;
input x_449;
input x_450;
input x_451;
input x_452;
input x_453;
input x_454;
input x_455;
input x_456;
input x_457;
input x_458;
input x_459;
input x_460;
input x_461;
input x_462;
input x_463;
input x_464;
input x_465;
input x_466;
input x_467;
input x_468;
input x_469;
input x_470;
input x_471;
input x_472;
input x_473;
input x_474;
input x_475;
input x_476;
input x_477;
input x_478;
input x_479;
input x_480;
input x_481;
input x_482;
input x_483;
input x_484;
input x_485;
input x_486;
input x_487;
input x_488;
input x_489;
input x_490;
input x_491;
input x_492;
input x_493;
input x_494;
input x_495;
input x_496;
input x_497;
input x_498;
input x_499;
input x_500;
input x_501;
input x_502;
input x_503;
input x_504;
input x_505;
input x_506;
input x_507;
input x_508;
input x_509;
input x_510;
input x_511;
input x_512;
input x_513;
input x_514;
input x_515;
input x_516;
input x_517;
input x_518;
input x_519;
input x_520;
input x_521;
input x_522;
input x_523;
input x_524;
input x_525;
input x_526;
input x_527;
input x_528;
input x_529;
input x_530;
input x_531;
input x_532;
input x_533;
input x_534;
input x_535;
input x_536;
input x_537;
input x_538;
input x_539;
input x_540;
input x_541;
input x_542;
input x_543;
input x_544;
input x_545;
input x_546;
input x_547;
input x_548;
input x_549;
input x_550;
input x_551;
input x_552;
input x_553;
input x_554;
input x_555;
input x_556;
input x_557;
input x_558;
input x_559;
input x_560;
input x_561;
input x_562;
input x_563;
input x_564;
input x_565;
input x_566;
input x_567;
input x_568;
input x_569;
input x_570;
input x_571;
input x_572;
input x_573;
input x_574;
input x_575;
input x_576;
input x_577;
input x_578;
input x_579;
input x_580;
input x_581;
input x_582;
input x_583;
input x_584;
input x_585;
input x_586;
input x_587;
input x_588;
input x_589;
input x_590;
input x_591;
input x_592;
input x_593;
input x_594;
input x_595;
input x_596;
input x_597;
input x_598;
input x_599;
input x_600;
input x_601;
input x_602;
input x_603;
input x_604;
input x_605;
input x_606;
input x_607;
input x_608;
input x_609;
input x_610;
input x_611;
input x_612;
input x_613;
input x_614;
input x_615;
input x_616;
input x_617;
input x_618;
input x_619;
input x_620;
input x_621;
input x_622;
input x_623;
input x_624;
input x_625;
input x_626;
input x_627;
input x_628;
input x_629;
input x_630;
input x_631;
input x_632;
input x_633;
input x_634;
input x_635;
input x_636;
input x_637;
input x_638;
input x_639;
input x_640;
input x_641;
input x_642;
input x_643;
input x_644;
input x_645;
input x_646;
input x_647;
input x_648;
input x_649;
input x_650;
input x_651;
input x_652;
input x_653;
input x_654;
input x_655;
input x_656;
input x_657;
input x_658;
input x_659;
input x_660;
input x_661;
input x_662;
input x_663;
input x_664;
input x_665;
input x_666;
input x_667;
input x_668;
input x_669;
input x_670;
input x_671;
input x_672;
input x_673;
input x_674;
input x_675;
input x_676;
input x_677;
input x_678;
input x_679;
input x_680;
input x_681;
input x_682;
input x_683;
input x_684;
input x_685;
input x_686;
input x_687;
input x_688;
input x_689;
input x_690;
input x_691;
input x_692;
input x_693;
input x_694;
input x_695;
input x_696;
input x_697;
input x_698;
input x_699;
input x_700;
input x_701;
input x_702;
input x_703;
input x_704;
input x_705;
input x_706;
input x_707;
input x_708;
input x_709;
input x_710;
input x_711;
input x_712;
input x_713;
input x_714;
input x_715;
input x_716;
input x_717;
input x_718;
input x_719;
input x_720;
input x_721;
input x_722;
input x_723;
input x_724;
input x_725;
input x_726;
input x_727;
input x_728;
input x_729;
input x_730;
input x_731;
input x_732;
input x_733;
input x_734;
input x_735;
input x_736;
input x_737;
input x_738;
input x_739;
input x_740;
input x_741;
input x_742;
input x_743;
input x_744;
input x_745;
input x_746;
input x_747;
input x_748;
input x_749;
input x_750;
input x_751;
input x_752;
input x_753;
input x_754;
input x_755;
input x_756;
input x_757;
input x_758;
input x_759;
input x_760;
input x_761;
input x_762;
input x_763;
input x_764;
input x_765;
input x_766;
input x_767;
input x_768;
input x_769;
input x_770;
input x_771;
input x_772;
input x_773;
input x_774;
input x_775;
input x_776;
input x_777;
input x_778;
input x_779;
input x_780;
input x_781;
input x_782;
input x_783;
input x_784;
input x_785;
input x_786;
input x_787;
input x_788;
input x_789;
input x_790;
input x_791;
input x_792;
input x_793;
input x_794;
input x_795;
input x_796;
input x_797;
input x_798;
input x_799;
input x_800;
input x_801;
input x_802;
input x_803;
input x_804;
input x_805;
input x_806;
input x_807;
input x_808;
input x_809;
input x_810;
input x_811;
input x_812;
input x_813;
input x_814;
input x_815;
input x_816;
input x_817;
input x_818;
input x_819;
input x_820;
input x_821;
input x_822;
input x_823;
input x_824;
input x_825;
input x_826;
input x_827;
input x_828;
input x_829;
input x_830;
input x_831;
input x_832;
input x_833;
input x_834;
input x_835;
input x_836;
input x_837;
input x_838;
input x_839;
input x_840;
input x_841;
input x_842;
input x_843;
input x_844;
input x_845;
input x_846;
input x_847;
input x_848;
input x_849;
input x_850;
input x_851;
input x_852;
input x_853;
input x_854;
input x_855;
input x_856;
input x_857;
input x_858;
input x_859;
input x_860;
input x_861;
input x_862;
input x_863;
input x_864;
input x_865;
input x_866;
input x_867;
input x_868;
input x_869;
input x_870;
input x_871;
input x_872;
input x_873;
input x_874;
input x_875;
input x_876;
input x_877;
input x_878;
input x_879;
input x_880;
input x_881;
input x_882;
input x_883;
input x_884;
input x_885;
input x_886;
input x_887;
input x_888;
input x_889;
input x_890;
input x_891;
input x_892;
input x_893;
input x_894;
input x_895;
input x_896;
input x_897;
input x_898;
input x_899;
input x_900;
input x_901;
input x_902;
input x_903;
input x_904;
input x_905;
input x_906;
input x_907;
input x_908;
input x_909;
input x_910;
input x_911;
input x_912;
input x_913;
input x_914;
input x_915;
input x_916;
input x_917;
input x_918;
input x_919;
input x_920;
input x_921;
input x_922;
input x_923;
input x_924;
input x_925;
input x_926;
input x_927;
input x_928;
input x_929;
input x_930;
input x_931;
input x_932;
input x_933;
input x_934;
input x_935;
input x_936;
input x_937;
input x_938;
input x_939;
input x_940;
input x_941;
input x_942;
input x_943;
input x_944;
input x_945;
input x_946;
input x_947;
input x_948;
input x_949;
input x_950;
input x_951;
input x_952;
input x_953;
input x_954;
input x_955;
input x_956;
input x_957;
input x_958;
input x_959;
input x_960;
input x_961;
input x_962;
input x_963;
input x_964;
input x_965;
input x_966;
input x_967;
input x_968;
input x_969;
input x_970;
input x_971;
input x_972;
input x_973;
input x_974;
input x_975;
input x_976;
input x_977;
input x_978;
input x_979;
input x_980;
input x_981;
input x_982;
input x_983;
input x_984;
input x_985;
input x_986;
input x_987;
input x_988;
input x_989;
input x_990;
input x_991;
input x_992;
input x_993;
input x_994;
input x_995;
input x_996;
input x_997;
input x_998;
input x_999;
input x_1000;
input x_1001;
input x_1002;
input x_1003;
input x_1004;
input x_1005;
input x_1006;
input x_1007;
input x_1008;
input x_1009;
input x_1010;
input x_1011;
input x_1012;
input x_1013;
input x_1014;
input x_1015;
input x_1016;
input x_1017;
input x_1018;
input x_1019;
input x_1020;
input x_1021;
input x_1022;
input x_1023;
input x_1024;
input x_1025;
input x_1026;
input x_1027;
input x_1028;
input x_1029;
input x_1030;
input x_1031;
input x_1032;
input x_1033;
input x_1034;
input x_1035;
input x_1036;
input x_1037;
input x_1038;
input x_1039;
input x_1040;
input x_1041;
input x_1042;
input x_1043;
input x_1044;
input x_1045;
input x_1046;
input x_1047;
input x_1048;
input x_1049;
input x_1050;
input x_1051;
input x_1052;
input x_1053;
input x_1054;
input x_1055;
input x_1056;
input x_1057;
input x_1058;
input x_1059;
input x_1060;
input x_1061;
input x_1062;
input x_1063;
input x_1064;
input x_1065;
input x_1066;
input x_1067;
input x_1068;
input x_1069;
input x_1070;
input x_1071;
input x_1072;
input x_1073;
input x_1074;
input x_1075;
input x_1076;
input x_1077;
input x_1078;
input x_1079;
input x_1080;
input x_1081;
input x_1082;
input x_1083;
input x_1084;
input x_1085;
input x_1086;
input x_1087;
input x_1088;
input x_1089;
input x_1090;
input x_1091;
input x_1092;
input x_1093;
input x_1094;
input x_1095;
input x_1096;
input x_1097;
input x_1098;
input x_1099;
input x_1100;
input x_1101;
input x_1102;
input x_1103;
input x_1104;
input x_1105;
input x_1106;
input x_1107;
input x_1108;
input x_1109;
input x_1110;
input x_1111;
input x_1112;
input x_1113;
input x_1114;
input x_1115;
input x_1116;
input x_1117;
input x_1118;
input x_1119;
input x_1120;
input x_1121;
input x_1122;
input x_1123;
input x_1124;
input x_1125;
input x_1126;
input x_1127;
input x_1128;
input x_1129;
input x_1130;
input x_1131;
input x_1132;
input x_1133;
input x_1134;
input x_1135;
input x_1136;
input x_1137;
input x_1138;
input x_1139;
input x_1140;
input x_1141;
input x_1142;
input x_1143;
input x_1144;
input x_1145;
input x_1146;
input x_1147;
input x_1148;
input x_1149;
input x_1150;
input x_1151;
input x_1152;
input x_1153;
input x_1154;
input x_1155;
input x_1156;
input x_1157;
input x_1158;
input x_1159;
input x_1160;
input x_1161;
input x_1162;
input x_1163;
input x_1164;
input x_1165;
input x_1166;
input x_1167;
input x_1168;
input x_1169;
input x_1170;
input x_1171;
input x_1172;
input x_1173;
input x_1174;
input x_1175;
input x_1176;
input x_1177;
input x_1178;
input x_1179;
input x_1180;
input x_1181;
input x_1182;
input x_1183;
input x_1184;
input x_1185;
input x_1186;
input x_1187;
input x_1188;
input x_1189;
input x_1190;
input x_1191;
input x_1192;
input x_1193;
input x_1194;
input x_1195;
input x_1196;
input x_1197;
input x_1198;
input x_1199;
input x_1200;
input x_1201;
input x_1202;
input x_1203;
input x_1204;
input x_1205;
input x_1206;
input x_1207;
input x_1208;
input x_1209;
input x_1210;
input x_1211;
input x_1212;
input x_1213;
input x_1214;
input x_1215;
input x_1216;
input x_1217;
input x_1218;
input x_1219;
input x_1220;
input x_1221;
input x_1222;
input x_1223;
input x_1224;
input x_1225;
input x_1226;
input x_1227;
input x_1228;
input x_1229;
input x_1230;
input x_1231;
input x_1232;
input x_1233;
input x_1234;
input x_1235;
input x_1236;
input x_1237;
input x_1238;
input x_1239;
input x_1240;
input x_1241;
input x_1242;
input x_1243;
input x_1244;
input x_1245;
input x_1246;
input x_1247;
input x_1248;
input x_1249;
input x_1250;
input x_1251;
input x_1252;
input x_1253;
input x_1254;
input x_1255;
input x_1256;
input x_1257;
input x_1258;
input x_1259;
input x_1260;
input x_1261;
input x_1262;
input x_1263;
input x_1264;
input x_1265;
input x_1266;
input x_1267;
input x_1268;
input x_1269;
input x_1270;
input x_1271;
input x_1272;
input x_1273;
input x_1274;
input x_1275;
input x_1276;
input x_1277;
input x_1278;
input x_1279;
input x_1280;
input x_1281;
input x_1282;
input x_1283;
input x_1284;
input x_1285;
input x_1286;
input x_1287;
input x_1288;
input x_1289;
input x_1290;
input x_1291;
input x_1292;
input x_1293;
input x_1294;
input x_1295;
input x_1296;
input x_1297;
input x_1298;
input x_1299;
input x_1300;
input x_1301;
input x_1302;
input x_1303;
input x_1304;
input x_1305;
input x_1306;
input x_1307;
input x_1308;
input x_1309;
input x_1310;
input x_1311;
input x_1312;
input x_1313;
input x_1314;
input x_1315;
input x_1316;
input x_1317;
input x_1318;
input x_1319;
input x_1320;
input x_1321;
input x_1322;
input x_1323;
input x_1324;
input x_1325;
input x_1326;
input x_1327;
input x_1328;
input x_1329;
input x_1330;
input x_1331;
input x_1332;
input x_1333;
input x_1334;
input x_1335;
input x_1336;
input x_1337;
input x_1338;
input x_1339;
input x_1340;
input x_1341;
input x_1342;
input x_1343;
input x_1344;
input x_1345;
input x_1346;
input x_1347;
input x_1348;
input x_1349;
input x_1350;
input x_1351;
input x_1352;
input x_1353;
input x_1354;
input x_1355;
input x_1356;
input x_1357;
input x_1358;
input x_1359;
input x_1360;
input x_1361;
input x_1362;
input x_1363;
input x_1364;
input x_1365;
input x_1366;
input x_1367;
input x_1368;
input x_1369;
input x_1370;
input x_1371;
input x_1372;
input x_1373;
input x_1374;
input x_1375;
input x_1376;
input x_1377;
input x_1378;
input x_1379;
input x_1380;
input x_1381;
input x_1382;
input x_1383;
input x_1384;
input x_1385;
input x_1386;
input x_1387;
input x_1388;
input x_1389;
input x_1390;
input x_1391;
input x_1392;
input x_1393;
input x_1394;
input x_1395;
input x_1396;
input x_1397;
input x_1398;
input x_1399;
input x_1400;
input x_1401;
input x_1402;
input x_1403;
input x_1404;
input x_1405;
input x_1406;
input x_1407;
input x_1408;
input x_1409;
input x_1410;
input x_1411;
input x_1412;
input x_1413;
input x_1414;
input x_1415;
input x_1416;
input x_1417;
input x_1418;
input x_1419;
input x_1420;
input x_1421;
input x_1422;
input x_1423;
input x_1424;
input x_1425;
input x_1426;
input x_1427;
input x_1428;
input x_1429;
input x_1430;
input x_1431;
input x_1432;
input x_1433;
input x_1434;
input x_1435;
input x_1436;
input x_1437;
input x_1438;
input x_1439;
input x_1440;
input x_1441;
input x_1442;
input x_1443;
input x_1444;
input x_1445;
input x_1446;
input x_1447;
input x_1448;
input x_1449;
input x_1450;
input x_1451;
input x_1452;
input x_1453;
input x_1454;
input x_1455;
input x_1456;
input x_1457;
input x_1458;
input x_1459;
input x_1460;
input x_1461;
input x_1462;
input x_1463;
input x_1464;
input x_1465;
input x_1466;
input x_1467;
input x_1468;
input x_1469;
input x_1470;
input x_1471;
input x_1472;
input x_1473;
input x_1474;
input x_1475;
input x_1476;
input x_1477;
input x_1478;
input x_1479;
input x_1480;
input x_1481;
input x_1482;
input x_1483;
input x_1484;
input x_1485;
input x_1486;
input x_1487;
input x_1488;
input x_1489;
input x_1490;
input x_1491;
input x_1492;
input x_1493;
input x_1494;
input x_1495;
input x_1496;
input x_1497;
input x_1498;
input x_1499;
input x_1500;
input x_1501;
input x_1502;
input x_1503;
input x_1504;
input x_1505;
input x_1506;
input x_1507;
input x_1508;
input x_1509;
input x_1510;
input x_1511;
input x_1512;
input x_1513;
input x_1514;
input x_1515;
input x_1516;
input x_1517;
input x_1518;
input x_1519;
input x_1520;
input x_1521;
input x_1522;
input x_1523;
input x_1524;
input x_1525;
input x_1526;
input x_1527;
input x_1528;
input x_1529;
input x_1530;
input x_1531;
input x_1532;
input x_1533;
input x_1534;
input x_1535;
input x_1536;
input x_1537;
input x_1538;
input x_1539;
input x_1540;
input x_1541;
input x_1542;
input x_1543;
input x_1544;
input x_1545;
input x_1546;
input x_1547;
input x_1548;
input x_1549;
input x_1550;
input x_1551;
input x_1552;
input x_1553;
input x_1554;
input x_1555;
input x_1556;
input x_1557;
input x_1558;
input x_1559;
input x_1560;
input x_1561;
input x_1562;
input x_1563;
input x_1564;
input x_1565;
input x_1566;
input x_1567;
input x_1568;
input x_1569;
input x_1570;
input x_1571;
input x_1572;
input x_1573;
input x_1574;
input x_1575;
input x_1576;
input x_1577;
input x_1578;
input x_1579;
input x_1580;
input x_1581;
input x_1582;
input x_1583;
input x_1584;
input x_1585;
input x_1586;
input x_1587;
input x_1588;
input x_1589;
input x_1590;
input x_1591;
input x_1592;
input x_1593;
input x_1594;
input x_1595;
input x_1596;
input x_1597;
input x_1598;
input x_1599;
input x_1600;
input x_1601;
input x_1602;
input x_1603;
input x_1604;
input x_1605;
input x_1606;
input x_1607;
input x_1608;
input x_1609;
input x_1610;
input x_1611;
input x_1612;
input x_1613;
input x_1614;
input x_1615;
input x_1616;
input x_1617;
input x_1618;
input x_1619;
input x_1620;
input x_1621;
input x_1622;
input x_1623;
input x_1624;
input x_1625;
input x_1626;
input x_1627;
input x_1628;
input x_1629;
input x_1630;
input x_1631;
input x_1632;
input x_1633;
input x_1634;
input x_1635;
input x_1636;
input x_1637;
input x_1638;
input x_1639;
input x_1640;
input x_1641;
input x_1642;
input x_1643;
input x_1644;
input x_1645;
input x_1646;
input x_1647;
input x_1648;
input x_1649;
input x_1650;
input x_1651;
input x_1652;
input x_1653;
input x_1654;
input x_1655;
input x_1656;
input x_1657;
input x_1658;
input x_1659;
input x_1660;
input x_1661;
input x_1662;
input x_1663;
input x_1664;
input x_1665;
input x_1666;
input x_1667;
input x_1668;
input x_1669;
input x_1670;
input x_1671;
input x_1672;
input x_1673;
input x_1674;
input x_1675;
input x_1676;
input x_1677;
input x_1678;
input x_1679;
input x_1680;
input x_1681;
input x_1682;
input x_1683;
input x_1684;
input x_1685;
input x_1686;
input x_1687;
input x_1688;
input x_1689;
input x_1690;
input x_1691;
input x_1692;
input x_1693;
input x_1694;
input x_1695;
input x_1696;
input x_1697;
input x_1698;
input x_1699;
input x_1700;
input x_1701;
input x_1702;
input x_1703;
input x_1704;
input x_1705;
input x_1706;
input x_1707;
input x_1708;
input x_1709;
input x_1710;
input x_1711;
input x_1712;
input x_1713;
input x_1714;
input x_1715;
input x_1716;
input x_1717;
input x_1718;
input x_1719;
input x_1720;
input x_1721;
input x_1722;
input x_1723;
input x_1724;
input x_1725;
input x_1726;
input x_1727;
input x_1728;
input x_1729;
input x_1730;
input x_1731;
input x_1732;
input x_1733;
input x_1734;
input x_1735;
input x_1736;
input x_1737;
input x_1738;
input x_1739;
input x_1740;
input x_1741;
input x_1742;
input x_1743;
input x_1744;
input x_1745;
input x_1746;
input x_1747;
input x_1748;
input x_1749;
input x_1750;
input x_1751;
input x_1752;
input x_1753;
input x_1754;
input x_1755;
input x_1756;
input x_1757;
input x_1758;
input x_1759;
input x_1760;
input x_1761;
input x_1762;
input x_1763;
input x_1764;
input x_1765;
input x_1766;
input x_1767;
input x_1768;
input x_1769;
input x_1770;
input x_1771;
input x_1772;
input x_1773;
input x_1774;
input x_1775;
input x_1776;
input x_1777;
input x_1778;
input x_1779;
input x_1780;
input x_1781;
input x_1782;
input x_1783;
input x_1784;
input x_1785;
input x_1786;
input x_1787;
input x_1788;
input x_1789;
input x_1790;
input x_1791;
input x_1792;
input x_1793;
input x_1794;
input x_1795;
input x_1796;
input x_1797;
input x_1798;
input x_1799;
input x_1800;
input x_1801;
input x_1802;
input x_1803;
input x_1804;
input x_1805;
input x_1806;
input x_1807;
input x_1808;
input x_1809;
input x_1810;
input x_1811;
input x_1812;
input x_1813;
input x_1814;
input x_1815;
input x_1816;
input x_1817;
input x_1818;
input x_1819;
input x_1820;
input x_1821;
input x_1822;
input x_1823;
input x_1824;
input x_1825;
input x_1826;
input x_1827;
input x_1828;
input x_1829;
input x_1830;
input x_1831;
input x_1832;
input x_1833;
input x_1834;
input x_1835;
input x_1836;
input x_1837;
input x_1838;
input x_1839;
input x_1840;
input x_1841;
input x_1842;
input x_1843;
input x_1844;
input x_1845;
input x_1846;
input x_1847;
input x_1848;
input x_1849;
input x_1850;
input x_1851;
input x_1852;
input x_1853;
input x_1854;
input x_1855;
input x_1856;
input x_1857;
input x_1858;
input x_1859;
input x_1860;
input x_1861;
input x_1862;
input x_1863;
input x_1864;
input x_1865;
input x_1866;
input x_1867;
input x_1868;
input x_1869;
input x_1870;
input x_1871;
input x_1872;
input x_1873;
input x_1874;
input x_1875;
input x_1876;
input x_1877;
input x_1878;
input x_1879;
input x_1880;
input x_1881;
input x_1882;
input x_1883;
input x_1884;
input x_1885;
input x_1886;
input x_1887;
input x_1888;
input x_1889;
input x_1890;
input x_1891;
input x_1892;
input x_1893;
input x_1894;
input x_1895;
input x_1896;
input x_1897;
input x_1898;
input x_1899;
input x_1900;
input x_1901;
input x_1902;
input x_1903;
input x_1904;
input x_1905;
input x_1906;
input x_1907;
input x_1908;
input x_1909;
input x_1910;
input x_1911;
input x_1912;
input x_1913;
input x_1914;
input x_1915;
input x_1916;
input x_1917;
input x_1918;
input x_1919;
input x_1920;
input x_1921;
input x_1922;
input x_1923;
input x_1924;
input x_1925;
input x_1926;
input x_1927;
input x_1928;
input x_1929;
input x_1930;
input x_1931;
input x_1932;
input x_1933;
input x_1934;
input x_1935;
input x_1936;
input x_1937;
input x_1938;
input x_1939;
input x_1940;
input x_1941;
input x_1942;
input x_1943;
input x_1944;
input x_1945;
input x_1946;
input x_1947;
input x_1948;
input x_1949;
input x_1950;
input x_1951;
input x_1952;
input x_1953;
input x_1954;
input x_1955;
input x_1956;
input x_1957;
input x_1958;
input x_1959;
input x_1960;
input x_1961;
input x_1962;
input x_1963;
input x_1964;
input x_1965;
input x_1966;
input x_1967;
input x_1968;
input x_1969;
input x_1970;
input x_1971;
input x_1972;
input x_1973;
input x_1974;
input x_1975;
input x_1976;
input x_1977;
input x_1978;
input x_1979;
input x_1980;
input x_1981;
input x_1982;
input x_1983;
input x_1984;
input x_1985;
input x_1986;
input x_1987;
input x_1988;
input x_1989;
input x_1990;
input x_1991;
input x_1992;
input x_1993;
input x_1994;
input x_1995;
input x_1996;
input x_1997;
input x_1998;
input x_1999;
input x_2000;
input x_2001;
input x_2002;
input x_2003;
input x_2004;
input x_2005;
input x_2006;
input x_2007;
input x_2008;
input x_2009;
input x_2010;
input x_2011;
input x_2012;
input x_2013;
input x_2014;
input x_2015;
input x_2016;
input x_2017;
input x_2018;
input x_2019;
input x_2020;
input x_2021;
input x_2022;
input x_2023;
input x_2024;
input x_2025;
input x_2026;
input x_2027;
input x_2028;
input x_2029;
input x_2030;
input x_2031;
input x_2032;
input x_2033;
input x_2034;
input x_2035;
input x_2036;
input x_2037;
input x_2038;
input x_2039;
input x_2040;
input x_2041;
input x_2042;
input x_2043;
input x_2044;
input x_2045;
input x_2046;
input x_2047;
input x_2048;
input x_2049;
input x_2050;
input x_2051;
input x_2052;
input x_2053;
input x_2054;
input x_2055;
input x_2056;
input x_2057;
input x_2058;
input x_2059;
input x_2060;
input x_2061;
input x_2062;
input x_2063;
input x_2064;
input x_2065;
input x_2066;
input x_2067;
input x_2068;
input x_2069;
input x_2070;
input x_2071;
input x_2072;
input x_2073;
input x_2074;
input x_2075;
input x_2076;
input x_2077;
input x_2078;
input x_2079;
input x_2080;
input x_2081;
input x_2082;
input x_2083;
input x_2084;
input x_2085;
input x_2086;
input x_2087;
input x_2088;
input x_2089;
input x_2090;
input x_2091;
input x_2092;
input x_2093;
input x_2094;
input x_2095;
input x_2096;
input x_2097;
input x_2098;
input x_2099;
input x_2100;
input x_2101;
input x_2102;
input x_2103;
input x_2104;
input x_2105;
input x_2106;
input x_2107;
input x_2108;
input x_2109;
input x_2110;
input x_2111;
input x_2112;
input x_2113;
input x_2114;
input x_2115;
input x_2116;
input x_2117;
input x_2118;
input x_2119;
input x_2120;
input x_2121;
input x_2122;
input x_2123;
input x_2124;
input x_2125;
input x_2126;
input x_2127;
input x_2128;
input x_2129;
input x_2130;
input x_2131;
input x_2132;
input x_2133;
input x_2134;
input x_2135;
input x_2136;
input x_2137;
input x_2138;
input x_2139;
input x_2140;
input x_2141;
input x_2142;
input x_2143;
input x_2144;
input x_2145;
input x_2146;
input x_2147;
input x_2148;
input x_2149;
input x_2150;
input x_2151;
input x_2152;
input x_2153;
input x_2154;
input x_2155;
input x_2156;
input x_2157;
input x_2158;
input x_2159;
input x_2160;
input x_2161;
input x_2162;
input x_2163;
input x_2164;
input x_2165;
input x_2166;
input x_2167;
input x_2168;
input x_2169;
input x_2170;
input x_2171;
input x_2172;
input x_2173;
input x_2174;
input x_2175;
input x_2176;
input x_2177;
input x_2178;
input x_2179;
input x_2180;
input x_2181;
input x_2182;
input x_2183;
input x_2184;
input x_2185;
input x_2186;
input x_2187;
input x_2188;
input x_2189;
input x_2190;
input x_2191;
input x_2192;
input x_2193;
input x_2194;
input x_2195;
input x_2196;
input x_2197;
input x_2198;
input x_2199;
input x_2200;
input x_2201;
input x_2202;
input x_2203;
input x_2204;
input x_2205;
input x_2206;
input x_2207;
input x_2208;
input x_2209;
input x_2210;
input x_2211;
input x_2212;
input x_2213;
input x_2214;
input x_2215;
input x_2216;
input x_2217;
input x_2218;
input x_2219;
input x_2220;
input x_2221;
input x_2222;
input x_2223;
input x_2224;
input x_2225;
input x_2226;
input x_2227;
input x_2228;
input x_2229;
input x_2230;
input x_2231;
input x_2232;
input x_2233;
input x_2234;
input x_2235;
input x_2236;
input x_2237;
input x_2238;
input x_2239;
input x_2240;
input x_2241;
input x_2242;
input x_2243;
input x_2244;
input x_2245;
input x_2246;
input x_2247;
input x_2248;
input x_2249;
input x_2250;
input x_2251;
input x_2252;
input x_2253;
input x_2254;
input x_2255;
input x_2256;
input x_2257;
input x_2258;
input x_2259;
input x_2260;
input x_2261;
input x_2262;
input x_2263;
input x_2264;
input x_2265;
input x_2266;
input x_2267;
input x_2268;
input x_2269;
input x_2270;
input x_2271;
input x_2272;
input x_2273;
input x_2274;
input x_2275;
input x_2276;
input x_2277;
input x_2278;
input x_2279;
input x_2280;
input x_2281;
input x_2282;
input x_2283;
input x_2284;
input x_2285;
input x_2286;
input x_2287;
input x_2288;
input x_2289;
input x_2290;
input x_2291;
input x_2292;
input x_2293;
input x_2294;
input x_2295;
input x_2296;
input x_2297;
input x_2298;
input x_2299;
input x_2300;
input x_2301;
input x_2302;
input x_2303;
input x_2304;
input x_2305;
input x_2306;
input x_2307;
input x_2308;
input x_2309;
input x_2310;
input x_2311;
input x_2312;
input x_2313;
input x_2314;
input x_2315;
input x_2316;
input x_2317;
input x_2318;
input x_2319;
input x_2320;
input x_2321;
input x_2322;
input x_2323;
input x_2324;
input x_2325;
input x_2326;
input x_2327;
input x_2328;
input x_2329;
input x_2330;
input x_2331;
input x_2332;
input x_2333;
input x_2334;
input x_2335;
input x_2336;
input x_2337;
input x_2338;
input x_2339;
input x_2340;
input x_2341;
input x_2342;
input x_2343;
input x_2344;
input x_2345;
input x_2346;
input x_2347;
input x_2348;
input x_2349;
input x_2350;
input x_2351;
input x_2352;
input x_2353;
input x_2354;
input x_2355;
input x_2356;
input x_2357;
input x_2358;
input x_2359;
input x_2360;
input x_2361;
input x_2362;
input x_2363;
input x_2364;
input x_2365;
input x_2366;
input x_2367;
input x_2368;
input x_2369;
input x_2370;
input x_2371;
input x_2372;
input x_2373;
input x_2374;
input x_2375;
input x_2376;
input x_2377;
input x_2378;
input x_2379;
input x_2380;
input x_2381;
input x_2382;
input x_2383;
input x_2384;
input x_2385;
input x_2386;
input x_2387;
input x_2388;
input x_2389;
input x_2390;
input x_2391;
input x_2392;
input x_2393;
input x_2394;
input x_2395;
input x_2396;
input x_2397;
input x_2398;
input x_2399;
input x_2400;
input x_2401;
input x_2402;
input x_2403;
input x_2404;
input x_2405;
input x_2406;
input x_2407;
input x_2408;
input x_2409;
input x_2410;
input x_2411;
input x_2412;
input x_2413;
input x_2414;
input x_2415;
input x_2416;
input x_2417;
input x_2418;
input x_2419;
input x_2420;
input x_2421;
input x_2422;
input x_2423;
input x_2424;
input x_2425;
input x_2426;
input x_2427;
input x_2428;
input x_2429;
input x_2430;
input x_2431;
input x_2432;
input x_2433;
input x_2434;
input x_2435;
input x_2436;
input x_2437;
input x_2438;
input x_2439;
input x_2440;
input x_2441;
input x_2442;
input x_2443;
input x_2444;
input x_2445;
input x_2446;
input x_2447;
input x_2448;
input x_2449;
input x_2450;
input x_2451;
input x_2452;
input x_2453;
input x_2454;
input x_2455;
input x_2456;
input x_2457;
input x_2458;
input x_2459;
input x_2460;
input x_2461;
input x_2462;
input x_2463;
input x_2464;
input x_2465;
input x_2466;
input x_2467;
input x_2468;
input x_2469;
input x_2470;
input x_2471;
input x_2472;
input x_2473;
input x_2474;
input x_2475;
input x_2476;
input x_2477;
input x_2478;
input x_2479;
input x_2480;
input x_2481;
input x_2482;
input x_2483;
input x_2484;
input x_2485;
input x_2486;
input x_2487;
input x_2488;
input x_2489;
input x_2490;
input x_2491;
input x_2492;
input x_2493;
input x_2494;
input x_2495;
input x_2496;
input x_2497;
input x_2498;
input x_2499;
input x_2500;
input x_2501;
input x_2502;
input x_2503;
input x_2504;
input x_2505;
input x_2506;
input x_2507;
input x_2508;
input x_2509;
input x_2510;
input x_2511;
input x_2512;
input x_2513;
input x_2514;
input x_2515;
input x_2516;
input x_2517;
input x_2518;
input x_2519;
input x_2520;
input x_2521;
input x_2522;
input x_2523;
input x_2524;
input x_2525;
input x_2526;
input x_2527;
input x_2528;
input x_2529;
input x_2530;
input x_2531;
input x_2532;
input x_2533;
input x_2534;
input x_2535;
input x_2536;
input x_2537;
input x_2538;
input x_2539;
input x_2540;
input x_2541;
input x_2542;
input x_2543;
input x_2544;
input x_2545;
input x_2546;
input x_2547;
input x_2548;
input x_2549;
input x_2550;
input x_2551;
input x_2552;
input x_2553;
input x_2554;
input x_2555;
input x_2556;
input x_2557;
input x_2558;
input x_2559;
input x_2560;
input x_2561;
input x_2562;
input x_2563;
input x_2564;
input x_2565;
input x_2566;
input x_2567;
input x_2568;
input x_2569;
input x_2570;
input x_2571;
input x_2572;
input x_2573;
input x_2574;
input x_2575;
input x_2576;
input x_2577;
input x_2578;
input x_2579;
input x_2580;
input x_2581;
input x_2582;
input x_2583;
input x_2584;
input x_2585;
input x_2586;
input x_2587;
input x_2588;
input x_2589;
input x_2590;
input x_2591;
input x_2592;
input x_2593;
input x_2594;
input x_2595;
input x_2596;
input x_2597;
input x_2598;
input x_2599;
input x_2600;
input x_2601;
input x_2602;
input x_2603;
input x_2604;
input x_2605;
input x_2606;
input x_2607;
input x_2608;
input x_2609;
input x_2610;
input x_2611;
input x_2612;
input x_2613;
input x_2614;
input x_2615;
input x_2616;
input x_2617;
input x_2618;
input x_2619;
input x_2620;
input x_2621;
input x_2622;
input x_2623;
input x_2624;
input x_2625;
input x_2626;
input x_2627;
input x_2628;
input x_2629;
input x_2630;
input x_2631;
input x_2632;
input x_2633;
input x_2634;
input x_2635;
input x_2636;
input x_2637;
input x_2638;
input x_2639;
input x_2640;
input x_2641;
input x_2642;
input x_2643;
input x_2644;
input x_2645;
input x_2646;
input x_2647;
input x_2648;
input x_2649;
input x_2650;
input x_2651;
input x_2652;
input x_2653;
input x_2654;
input x_2655;
input x_2656;
input x_2657;
input x_2658;
input x_2659;
input x_2660;
input x_2661;
input x_2662;
input x_2663;
input x_2664;
input x_2665;
input x_2666;
input x_2667;
input x_2668;
input x_2669;
input x_2670;
input x_2671;
input x_2672;
input x_2673;
input x_2674;
input x_2675;
input x_2676;
input x_2677;
input x_2678;
input x_2679;
input x_2680;
input x_2681;
input x_2682;
input x_2683;
input x_2684;
input x_2685;
input x_2686;
input x_2687;
input x_2688;
input x_2689;
input x_2690;
input x_2691;
input x_2692;
input x_2693;
input x_2694;
input x_2695;
input x_2696;
input x_2697;
input x_2698;
input x_2699;
input x_2700;
input x_2701;
input x_2702;
input x_2703;
input x_2704;
input x_2705;
input x_2706;
input x_2707;
input x_2708;
input x_2709;
input x_2710;
input x_2711;
input x_2712;
input x_2713;
input x_2714;
input x_2715;
input x_2716;
input x_2717;
input x_2718;
input x_2719;
input x_2720;
input x_2721;
input x_2722;
input x_2723;
input x_2724;
input x_2725;
input x_2726;
input x_2727;
input x_2728;
input x_2729;
input x_2730;
input x_2731;
input x_2732;
input x_2733;
input x_2734;
input x_2735;
input x_2736;
input x_2737;
input x_2738;
input x_2739;
input x_2740;
input x_2741;
input x_2742;
input x_2743;
input x_2744;
input x_2745;
input x_2746;
input x_2747;
input x_2748;
input x_2749;
input x_2750;
input x_2751;
input x_2752;
input x_2753;
input x_2754;
input x_2755;
input x_2756;
input x_2757;
input x_2758;
input x_2759;
input x_2760;
input x_2761;
input x_2762;
input x_2763;
input x_2764;
input x_2765;
input x_2766;
input x_2767;
input x_2768;
input x_2769;
input x_2770;
input x_2771;
input x_2772;
input x_2773;
input x_2774;
input x_2775;
input x_2776;
input x_2777;
input x_2778;
input x_2779;
input x_2780;
input x_2781;
input x_2782;
input x_2783;
input x_2784;
input x_2785;
input x_2786;
input x_2787;
input x_2788;
input x_2789;
input x_2790;
input x_2791;
input x_2792;
input x_2793;
input x_2794;
input x_2795;
input x_2796;
input x_2797;
input x_2798;
input x_2799;
input x_2800;
input x_2801;
input x_2802;
input x_2803;
input x_2804;
input x_2805;
input x_2806;
input x_2807;
input x_2808;
input x_2809;
input x_2810;
input x_2811;
input x_2812;
input x_2813;
input x_2814;
input x_2815;
input x_2816;
input x_2817;
input x_2818;
input x_2819;
input x_2820;
input x_2821;
input x_2822;
input x_2823;
input x_2824;
input x_2825;
input x_2826;
input x_2827;
input x_2828;
input x_2829;
input x_2830;
input x_2831;
input x_2832;
input x_2833;
input x_2834;
input x_2835;
input x_2836;
input x_2837;
input x_2838;
input x_2839;
input x_2840;
input x_2841;
input x_2842;
input x_2843;
input x_2844;
input x_2845;
input x_2846;
input x_2847;
input x_2848;
input x_2849;
input x_2850;
input x_2851;
input x_2852;
input x_2853;
input x_2854;
input x_2855;
input x_2856;
input x_2857;
input x_2858;
input x_2859;
input x_2860;
input x_2861;
input x_2862;
input x_2863;
input x_2864;
input x_2865;
input x_2866;
input x_2867;
input x_2868;
input x_2869;
input x_2870;
input x_2871;
input x_2872;
input x_2873;
input x_2874;
input x_2875;
input x_2876;
input x_2877;
input x_2878;
input x_2879;
input x_2880;
input x_2881;
input x_2882;
input x_2883;
input x_2884;
input x_2885;
input x_2886;
input x_2887;
input x_2888;
input x_2889;
input x_2890;
input x_2891;
input x_2892;
input x_2893;
input x_2894;
input x_2895;
input x_2896;
input x_2897;
input x_2898;
input x_2899;
input x_2900;
input x_2901;
input x_2902;
input x_2903;
input x_2904;
input x_2905;
input x_2906;
input x_2907;
input x_2908;
input x_2909;
input x_2910;
input x_2911;
input x_2912;
input x_2913;
input x_2914;
input x_2915;
input x_2916;
input x_2917;
input x_2918;
input x_2919;
input x_2920;
input x_2921;
input x_2922;
input x_2923;
input x_2924;
input x_2925;
input x_2926;
input x_2927;
input x_2928;
input x_2929;
input x_2930;
input x_2931;
input x_2932;
input x_2933;
input x_2934;
input x_2935;
input x_2936;
input x_2937;
input x_2938;
input x_2939;
input x_2940;
input x_2941;
input x_2942;
input x_2943;
input x_2944;
input x_2945;
input x_2946;
input x_2947;
input x_2948;
input x_2949;
input x_2950;
input x_2951;
input x_2952;
input x_2953;
input x_2954;
input x_2955;
input x_2956;
input x_2957;
input x_2958;
input x_2959;
input x_2960;
input x_2961;
input x_2962;
input x_2963;
input x_2964;
input x_2965;
input x_2966;
input x_2967;
input x_2968;
input x_2969;
input x_2970;
input x_2971;
input x_2972;
input x_2973;
input x_2974;
input x_2975;
input x_2976;
input x_2977;
input x_2978;
input x_2979;
input x_2980;
input x_2981;
input x_2982;
input x_2983;
input x_2984;
input x_2985;
input x_2986;
input x_2987;
input x_2988;
input x_2989;
input x_2990;
input x_2991;
input x_2992;
input x_2993;
input x_2994;
input x_2995;
input x_2996;
input x_2997;
input x_2998;
input x_2999;
input x_3000;
input x_3001;
input x_3002;
input x_3003;
input x_3004;
input x_3005;
input x_3006;
input x_3007;
input x_3008;
input x_3009;
input x_3010;
input x_3011;
input x_3012;
input x_3013;
input x_3014;
input x_3015;
input x_3016;
input x_3017;
input x_3018;
input x_3019;
input x_3020;
input x_3021;
input x_3022;
input x_3023;
input x_3024;
input x_3025;
input x_3026;
input x_3027;
input x_3028;
input x_3029;
input x_3030;
input x_3031;
input x_3032;
input x_3033;
input x_3034;
input x_3035;
input x_3036;
input x_3037;
input x_3038;
input x_3039;
input x_3040;
input x_3041;
input x_3042;
input x_3043;
input x_3044;
input x_3045;
input x_3046;
input x_3047;
input x_3048;
input x_3049;
input x_3050;
input x_3051;
input x_3052;
input x_3053;
input x_3054;
input x_3055;
input x_3056;
input x_3057;
input x_3058;
input x_3059;
input x_3060;
input x_3061;
input x_3062;
input x_3063;
input x_3064;
input x_3065;
input x_3066;
input x_3067;
input x_3068;
input x_3069;
input x_3070;
input x_3071;
input x_3072;
input x_3073;
input x_3074;
input x_3075;
input x_3076;
input x_3077;
input x_3078;
input x_3079;
input x_3080;
input x_3081;
input x_3082;
input x_3083;
input x_3084;
input x_3085;
input x_3086;
input x_3087;
input x_3088;
input x_3089;
input x_3090;
input x_3091;
input x_3092;
input x_3093;
input x_3094;
input x_3095;
input x_3096;
input x_3097;
input x_3098;
input x_3099;
input x_3100;
input x_3101;
input x_3102;
input x_3103;
input x_3104;
input x_3105;
input x_3106;
input x_3107;
input x_3108;
input x_3109;
input x_3110;
input x_3111;
input x_3112;
input x_3113;
input x_3114;
input x_3115;
input x_3116;
input x_3117;
input x_3118;
input x_3119;
input x_3120;
input x_3121;
input x_3122;
input x_3123;
input x_3124;
input x_3125;
input x_3126;
input x_3127;
input x_3128;
input x_3129;
input x_3130;
input x_3131;
input x_3132;
input x_3133;
input x_3134;
input x_3135;
input x_3136;
input x_3137;
input x_3138;
input x_3139;
input x_3140;
input x_3141;
input x_3142;
input x_3143;
input x_3144;
input x_3145;
input x_3146;
input x_3147;
input x_3148;
input x_3149;
input x_3150;
input x_3151;
input x_3152;
input x_3153;
input x_3154;
input x_3155;
input x_3156;
input x_3157;
input x_3158;
input x_3159;
input x_3160;
input x_3161;
input x_3162;
input x_3163;
input x_3164;
input x_3165;
input x_3166;
input x_3167;
input x_3168;
input x_3169;
input x_3170;
input x_3171;
input x_3172;
input x_3173;
input x_3174;
input x_3175;
input x_3176;
input x_3177;
input x_3178;
input x_3179;
input x_3180;
input x_3181;
input x_3182;
input x_3183;
input x_3184;
input x_3185;
input x_3186;
input x_3187;
input x_3188;
input x_3189;
input x_3190;
input x_3191;
input x_3192;
input x_3193;
input x_3194;
input x_3195;
input x_3196;
input x_3197;
input x_3198;
input x_3199;
input x_3200;
input x_3201;
input x_3202;
input x_3203;
input x_3204;
input x_3205;
input x_3206;
input x_3207;
input x_3208;
input x_3209;
input x_3210;
input x_3211;
input x_3212;
input x_3213;
input x_3214;
input x_3215;
input x_3216;
input x_3217;
input x_3218;
input x_3219;
input x_3220;
input x_3221;
input x_3222;
input x_3223;
input x_3224;
input x_3225;
input x_3226;
input x_3227;
input x_3228;
input x_3229;
input x_3230;
input x_3231;
input x_3232;
input x_3233;
input x_3234;
input x_3235;
input x_3236;
input x_3237;
input x_3238;
input x_3239;
input x_3240;
input x_3241;
input x_3242;
input x_3243;
input x_3244;
input x_3245;
input x_3246;
input x_3247;
input x_3248;
input x_3249;
input x_3250;
input x_3251;
input x_3252;
input x_3253;
input x_3254;
input x_3255;
input x_3256;
input x_3257;
input x_3258;
input x_3259;
input x_3260;
input x_3261;
input x_3262;
input x_3263;
input x_3264;
input x_3265;
input x_3266;
input x_3267;
input x_3268;
input x_3269;
input x_3270;
input x_3271;
input x_3272;
input x_3273;
input x_3274;
input x_3275;
input x_3276;
input x_3277;
input x_3278;
input x_3279;
input x_3280;
input x_3281;
input x_3282;
input x_3283;
input x_3284;
input x_3285;
input x_3286;
input x_3287;
input x_3288;
input x_3289;
input x_3290;
input x_3291;
input x_3292;
input x_3293;
input x_3294;
input x_3295;
input x_3296;
input x_3297;
input x_3298;
input x_3299;
input x_3300;
input x_3301;
input x_3302;
input x_3303;
input x_3304;
input x_3305;
input x_3306;
input x_3307;
input x_3308;
input x_3309;
input x_3310;
input x_3311;
input x_3312;
input x_3313;
input x_3314;
input x_3315;
input x_3316;
input x_3317;
input x_3318;
input x_3319;
input x_3320;
input x_3321;
input x_3322;
input x_3323;
input x_3324;
input x_3325;
input x_3326;
input x_3327;
input x_3328;
input x_3329;
input x_3330;
input x_3331;
input x_3332;
input x_3333;
input x_3334;
input x_3335;
input x_3336;
input x_3337;
input x_3338;
input x_3339;
input x_3340;
input x_3341;
input x_3342;
input x_3343;
input x_3344;
input x_3345;
input x_3346;
input x_3347;
input x_3348;
input x_3349;
input x_3350;
input x_3351;
input x_3352;
input x_3353;
input x_3354;
input x_3355;
input x_3356;
input x_3357;
input x_3358;
input x_3359;
input x_3360;
input x_3361;
input x_3362;
input x_3363;
input x_3364;
input x_3365;
input x_3366;
input x_3367;
input x_3368;
input x_3369;
input x_3370;
input x_3371;
input x_3372;
input x_3373;
input x_3374;
input x_3375;
input x_3376;
input x_3377;
input x_3378;
input x_3379;
input x_3380;
input x_3381;
input x_3382;
input x_3383;
input x_3384;
input x_3385;
input x_3386;
input x_3387;
input x_3388;
input x_3389;
input x_3390;
input x_3391;
input x_3392;
input x_3393;
input x_3394;
input x_3395;
input x_3396;
input x_3397;
input x_3398;
input x_3399;
input x_3400;
input x_3401;
input x_3402;
input x_3403;
input x_3404;
input x_3405;
input x_3406;
input x_3407;
input x_3408;
input x_3409;
input x_3410;
input x_3411;
input x_3412;
input x_3413;
input x_3414;
input x_3415;
input x_3416;
input x_3417;
input x_3418;
input x_3419;
input x_3420;
input x_3421;
input x_3422;
input x_3423;
input x_3424;
input x_3425;
input x_3426;
input x_3427;
input x_3428;
input x_3429;
input x_3430;
input x_3431;
input x_3432;
input x_3433;
input x_3434;
input x_3435;
input x_3436;
input x_3437;
input x_3438;
input x_3439;
input x_3440;
input x_3441;
input x_3442;
input x_3443;
input x_3444;
input x_3445;
input x_3446;
input x_3447;
input x_3448;
input x_3449;
input x_3450;
input x_3451;
input x_3452;
input x_3453;
input x_3454;
input x_3455;
input x_3456;
input x_3457;
input x_3458;
input x_3459;
input x_3460;
input x_3461;
input x_3462;
input x_3463;
input x_3464;
input x_3465;
input x_3466;
input x_3467;
input x_3468;
input x_3469;
input x_3470;
input x_3471;
input x_3472;
input x_3473;
input x_3474;
input x_3475;
input x_3476;
input x_3477;
input x_3478;
input x_3479;
input x_3480;
input x_3481;
input x_3482;
input x_3483;
input x_3484;
input x_3485;
input x_3486;
input x_3487;
input x_3488;
input x_3489;
input x_3490;
input x_3491;
input x_3492;
input x_3493;
input x_3494;
input x_3495;
input x_3496;
input x_3497;
input x_3498;
input x_3499;
input x_3500;
input x_3501;
input x_3502;
input x_3503;
input x_3504;
input x_3505;
input x_3506;
input x_3507;
input x_3508;
input x_3509;
input x_3510;
input x_3511;
input x_3512;
input x_3513;
input x_3514;
input x_3515;
input x_3516;
input x_3517;
input x_3518;
input x_3519;
input x_3520;
input x_3521;
input x_3522;
input x_3523;
input x_3524;
input x_3525;
input x_3526;
input x_3527;
input x_3528;
input x_3529;
input x_3530;
input x_3531;
input x_3532;
input x_3533;
input x_3534;
input x_3535;
input x_3536;
input x_3537;
input x_3538;
input x_3539;
input x_3540;
input x_3541;
input x_3542;
input x_3543;
input x_3544;
input x_3545;
input x_3546;
input x_3547;
input x_3548;
input x_3549;
input x_3550;
input x_3551;
input x_3552;
input x_3553;
input x_3554;
input x_3555;
input x_3556;
input x_3557;
input x_3558;
input x_3559;
input x_3560;
input x_3561;
input x_3562;
input x_3563;
input x_3564;
input x_3565;
input x_3566;
input x_3567;
input x_3568;
input x_3569;
input x_3570;
input x_3571;
input x_3572;
input x_3573;
input x_3574;
input x_3575;
input x_3576;
input x_3577;
input x_3578;
input x_3579;
input x_3580;
input x_3581;
input x_3582;
input x_3583;
input x_3584;
input x_3585;
input x_3586;
input x_3587;
input x_3588;
input x_3589;
input x_3590;
input x_3591;
input x_3592;
input x_3593;
input x_3594;
input x_3595;
input x_3596;
input x_3597;
input x_3598;
input x_3599;
input x_3600;
input x_3601;
input x_3602;
input x_3603;
input x_3604;
input x_3605;
input x_3606;
input x_3607;
input x_3608;
input x_3609;
input x_3610;
input x_3611;
input x_3612;
input x_3613;
input x_3614;
input x_3615;
input x_3616;
input x_3617;
input x_3618;
input x_3619;
input x_3620;
input x_3621;
input x_3622;
input x_3623;
input x_3624;
input x_3625;
input x_3626;
input x_3627;
input x_3628;
input x_3629;
input x_3630;
input x_3631;
input x_3632;
input x_3633;
input x_3634;
input x_3635;
input x_3636;
input x_3637;
input x_3638;
input x_3639;
input x_3640;
input x_3641;
input x_3642;
input x_3643;
input x_3644;
input x_3645;
input x_3646;
input x_3647;
input x_3648;
input x_3649;
input x_3650;
input x_3651;
input x_3652;
input x_3653;
input x_3654;
input x_3655;
input x_3656;
input x_3657;
input x_3658;
input x_3659;
input x_3660;
input x_3661;
input x_3662;
input x_3663;
input x_3664;
input x_3665;
input x_3666;
input x_3667;
input x_3668;
input x_3669;
input x_3670;
input x_3671;
input x_3672;
input x_3673;
input x_3674;
input x_3675;
input x_3676;
input x_3677;
input x_3678;
input x_3679;
input x_3680;
input x_3681;
input x_3682;
input x_3683;
input x_3684;
input x_3685;
input x_3686;
input x_3687;
input x_3688;
input x_3689;
input x_3690;
input x_3691;
input x_3692;
input x_3693;
input x_3694;
input x_3695;
input x_3696;
input x_3697;
input x_3698;
input x_3699;
input x_3700;
input x_3701;
input x_3702;
input x_3703;
input x_3704;
input x_3705;
input x_3706;
input x_3707;
input x_3708;
input x_3709;
input x_3710;
input x_3711;
input x_3712;
input x_3713;
input x_3714;
input x_3715;
input x_3716;
input x_3717;
input x_3718;
input x_3719;
input x_3720;
input x_3721;
input x_3722;
input x_3723;
input x_3724;
input x_3725;
input x_3726;
input x_3727;
input x_3728;
input x_3729;
input x_3730;
input x_3731;
input x_3732;
input x_3733;
input x_3734;
input x_3735;
input x_3736;
input x_3737;
input x_3738;
input x_3739;
input x_3740;
input x_3741;
input x_3742;
input x_3743;
input x_3744;
input x_3745;
input x_3746;
input x_3747;
input x_3748;
input x_3749;
input x_3750;
input x_3751;
input x_3752;
input x_3753;
input x_3754;
input x_3755;
input x_3756;
input x_3757;
input x_3758;
input x_3759;
input x_3760;
input x_3761;
input x_3762;
input x_3763;
input x_3764;
input x_3765;
input x_3766;
input x_3767;
input x_3768;
input x_3769;
input x_3770;
input x_3771;
input x_3772;
input x_3773;
input x_3774;
input x_3775;
input x_3776;
input x_3777;
input x_3778;
input x_3779;
input x_3780;
input x_3781;
input x_3782;
input x_3783;
input x_3784;
input x_3785;
input x_3786;
input x_3787;
input x_3788;
input x_3789;
input x_3790;
input x_3791;
input x_3792;
input x_3793;
input x_3794;
input x_3795;
input x_3796;
input x_3797;
input x_3798;
input x_3799;
input x_3800;
input x_3801;
input x_3802;
input x_3803;
input x_3804;
input x_3805;
input x_3806;
input x_3807;
input x_3808;
input x_3809;
input x_3810;
input x_3811;
input x_3812;
input x_3813;
input x_3814;
input x_3815;
input x_3816;
input x_3817;
input x_3818;
input x_3819;
input x_3820;
input x_3821;
input x_3822;
input x_3823;
input x_3824;
input x_3825;
input x_3826;
input x_3827;
input x_3828;
input x_3829;
input x_3830;
input x_3831;
input x_3832;
input x_3833;
input x_3834;
input x_3835;
input x_3836;
input x_3837;
input x_3838;
input x_3839;
input x_3840;
input x_3841;
input x_3842;
input x_3843;
input x_3844;
input x_3845;
input x_3846;
input x_3847;
input x_3848;
input x_3849;
input x_3850;
input x_3851;
input x_3852;
input x_3853;
input x_3854;
input x_3855;
input x_3856;
input x_3857;
input x_3858;
input x_3859;
input x_3860;
input x_3861;
input x_3862;
input x_3863;
input x_3864;
input x_3865;
input x_3866;
input x_3867;
input x_3868;
input x_3869;
input x_3870;
input x_3871;
input x_3872;
input x_3873;
input x_3874;
input x_3875;
input x_3876;
input x_3877;
input x_3878;
input x_3879;
input x_3880;
input x_3881;
input x_3882;
input x_3883;
input x_3884;
input x_3885;
input x_3886;
input x_3887;
input x_3888;
input x_3889;
input x_3890;
input x_3891;
input x_3892;
input x_3893;
input x_3894;
input x_3895;
input x_3896;
input x_3897;
input x_3898;
input x_3899;
input x_3900;
input x_3901;
input x_3902;
input x_3903;
input x_3904;
input x_3905;
input x_3906;
input x_3907;
input x_3908;
input x_3909;
input x_3910;
input x_3911;
input x_3912;
input x_3913;
input x_3914;
input x_3915;
input x_3916;
input x_3917;
input x_3918;
input x_3919;
input x_3920;
input x_3921;
input x_3922;
input x_3923;
input x_3924;
input x_3925;
input x_3926;
input x_3927;
input x_3928;
input x_3929;
input x_3930;
input x_3931;
input x_3932;
input x_3933;
input x_3934;
input x_3935;
input x_3936;
input x_3937;
input x_3938;
input x_3939;
input x_3940;
input x_3941;
input x_3942;
input x_3943;
input x_3944;
input x_3945;
input x_3946;
input x_3947;
input x_3948;
input x_3949;
input x_3950;
input x_3951;
input x_3952;
input x_3953;
input x_3954;
input x_3955;
input x_3956;
input x_3957;
input x_3958;
input x_3959;
input x_3960;
input x_3961;
input x_3962;
input x_3963;
input x_3964;
input x_3965;
input x_3966;
input x_3967;
input x_3968;
input x_3969;
input x_3970;
input x_3971;
input x_3972;
input x_3973;
input x_3974;
input x_3975;
input x_3976;
input x_3977;
input x_3978;
input x_3979;
input x_3980;
input x_3981;
input x_3982;
input x_3983;
input x_3984;
input x_3985;
input x_3986;
input x_3987;
input x_3988;
input x_3989;
input x_3990;
input x_3991;
input x_3992;
input x_3993;
input x_3994;
input x_3995;
input x_3996;
input x_3997;
input x_3998;
input x_3999;
input x_4000;
input x_4001;
input x_4002;
input x_4003;
input x_4004;
input x_4005;
input x_4006;
input x_4007;
input x_4008;
input x_4009;
input x_4010;
input x_4011;
input x_4012;
input x_4013;
input x_4014;
input x_4015;
input x_4016;
input x_4017;
input x_4018;
input x_4019;
input x_4020;
input x_4021;
input x_4022;
input x_4023;
input x_4024;
input x_4025;
input x_4026;
input x_4027;
input x_4028;
input x_4029;
input x_4030;
input x_4031;
input x_4032;
input x_4033;
input x_4034;
input x_4035;
input x_4036;
input x_4037;
input x_4038;
input x_4039;
input x_4040;
input x_4041;
input x_4042;
input x_4043;
input x_4044;
input x_4045;
input x_4046;
input x_4047;
input x_4048;
input x_4049;
input x_4050;
input x_4051;
input x_4052;
input x_4053;
input x_4054;
input x_4055;
input x_4056;
input x_4057;
input x_4058;
input x_4059;
input x_4060;
input x_4061;
input x_4062;
input x_4063;
input x_4064;
input x_4065;
input x_4066;
input x_4067;
input x_4068;
input x_4069;
input x_4070;
input x_4071;
input x_4072;
input x_4073;
input x_4074;
input x_4075;
input x_4076;
input x_4077;
input x_4078;
input x_4079;
input x_4080;
input x_4081;
input x_4082;
input x_4083;
input x_4084;
input x_4085;
input x_4086;
input x_4087;
input x_4088;
input x_4089;
input x_4090;
input x_4091;
input x_4092;
input x_4093;
input x_4094;
input x_4095;
input x_4096;
input x_4097;
input x_4098;
input x_4099;
input x_4100;
input x_4101;
input x_4102;
input x_4103;
input x_4104;
input x_4105;
input x_4106;
input x_4107;
input x_4108;
input x_4109;
input x_4110;
input x_4111;
input x_4112;
input x_4113;
input x_4114;
input x_4115;
input x_4116;
input x_4117;
input x_4118;
input x_4119;
input x_4120;
input x_4121;
input x_4122;
input x_4123;
input x_4124;
input x_4125;
input x_4126;
input x_4127;
input x_4128;
input x_4129;
input x_4130;
input x_4131;
input x_4132;
input x_4133;
input x_4134;
input x_4135;
input x_4136;
input x_4137;
input x_4138;
input x_4139;
input x_4140;
input x_4141;
input x_4142;
input x_4143;
input x_4144;
input x_4145;
input x_4146;
input x_4147;
input x_4148;
input x_4149;
input x_4150;
input x_4151;
input x_4152;
input x_4153;
input x_4154;
input x_4155;
input x_4156;
input x_4157;
input x_4158;
input x_4159;
input x_4160;
input x_4161;
input x_4162;
input x_4163;
input x_4164;
input x_4165;
input x_4166;
input x_4167;
input x_4168;
input x_4169;
input x_4170;
input x_4171;
input x_4172;
input x_4173;
input x_4174;
input x_4175;
input x_4176;
input x_4177;
input x_4178;
input x_4179;
input x_4180;
input x_4181;
input x_4182;
input x_4183;
input x_4184;
input x_4185;
input x_4186;
input x_4187;
input x_4188;
input x_4189;
input x_4190;
input x_4191;
input x_4192;
input x_4193;
input x_4194;
input x_4195;
input x_4196;
input x_4197;
input x_4198;
input x_4199;
input x_4200;
input x_4201;
input x_4202;
input x_4203;
input x_4204;
input x_4205;
input x_4206;
input x_4207;
input x_4208;
input x_4209;
input x_4210;
input x_4211;
input x_4212;
input x_4213;
input x_4214;
input x_4215;
input x_4216;
input x_4217;
input x_4218;
input x_4219;
input x_4220;
input x_4221;
input x_4222;
input x_4223;
input x_4224;
input x_4225;
input x_4226;
input x_4227;
input x_4228;
input x_4229;
input x_4230;
input x_4231;
input x_4232;
input x_4233;
input x_4234;
input x_4235;
input x_4236;
input x_4237;
input x_4238;
input x_4239;
input x_4240;
input x_4241;
input x_4242;
input x_4243;
input x_4244;
input x_4245;
input x_4246;
input x_4247;
input x_4248;
input x_4249;
input x_4250;
input x_4251;
input x_4252;
input x_4253;
input x_4254;
input x_4255;
input x_4256;
input x_4257;
input x_4258;
input x_4259;
input x_4260;
input x_4261;
input x_4262;
input x_4263;
input x_4264;
input x_4265;
input x_4266;
input x_4267;
input x_4268;
input x_4269;
input x_4270;
input x_4271;
input x_4272;
input x_4273;
input x_4274;
input x_4275;
input x_4276;
input x_4277;
input x_4278;
input x_4279;
input x_4280;
input x_4281;
input x_4282;
input x_4283;
input x_4284;
input x_4285;
input x_4286;
input x_4287;
input x_4288;
input x_4289;
input x_4290;
input x_4291;
input x_4292;
input x_4293;
input x_4294;
input x_4295;
input x_4296;
input x_4297;
input x_4298;
input x_4299;
input x_4300;
input x_4301;
input x_4302;
input x_4303;
input x_4304;
input x_4305;
input x_4306;
input x_4307;
input x_4308;
input x_4309;
input x_4310;
input x_4311;
input x_4312;
input x_4313;
input x_4314;
input x_4315;
input x_4316;
input x_4317;
input x_4318;
input x_4319;
input x_4320;
input x_4321;
input x_4322;
input x_4323;
input x_4324;
input x_4325;
input x_4326;
input x_4327;
input x_4328;
input x_4329;
input x_4330;
input x_4331;
input x_4332;
input x_4333;
input x_4334;
input x_4335;
input x_4336;
input x_4337;
input x_4338;
input x_4339;
input x_4340;
input x_4341;
input x_4342;
input x_4343;
input x_4344;
input x_4345;
input x_4346;
input x_4347;
input x_4348;
input x_4349;
input x_4350;
input x_4351;
input x_4352;
input x_4353;
input x_4354;
input x_4355;
input x_4356;
input x_4357;
input x_4358;
input x_4359;
input x_4360;
input x_4361;
input x_4362;
input x_4363;
input x_4364;
input x_4365;
input x_4366;
input x_4367;
input x_4368;
input x_4369;
input x_4370;
input x_4371;
input x_4372;
input x_4373;
input x_4374;
input x_4375;
input x_4376;
input x_4377;
input x_4378;
input x_4379;
input x_4380;
input x_4381;
input x_4382;
input x_4383;
input x_4384;
input x_4385;
input x_4386;
input x_4387;
input x_4388;
input x_4389;
input x_4390;
input x_4391;
input x_4392;
input x_4393;
input x_4394;
input x_4395;
input x_4396;
input x_4397;
input x_4398;
input x_4399;
input x_4400;
input x_4401;
input x_4402;
input x_4403;
input x_4404;
input x_4405;
input x_4406;
input x_4407;
input x_4408;
input x_4409;
input x_4410;
input x_4411;
input x_4412;
input x_4413;
input x_4414;
input x_4415;
input x_4416;
input x_4417;
input x_4418;
input x_4419;
input x_4420;
input x_4421;
input x_4422;
input x_4423;
input x_4424;
input x_4425;
input x_4426;
input x_4427;
input x_4428;
input x_4429;
input x_4430;
input x_4431;
input x_4432;
input x_4433;
input x_4434;
input x_4435;
input x_4436;
input x_4437;
input x_4438;
input x_4439;
input x_4440;
input x_4441;
input x_4442;
input x_4443;
input x_4444;
input x_4445;
input x_4446;
input x_4447;
input x_4448;
input x_4449;
input x_4450;
input x_4451;
input x_4452;
input x_4453;
input x_4454;
input x_4455;
input x_4456;
input x_4457;
input x_4458;
input x_4459;
input x_4460;
input x_4461;
input x_4462;
input x_4463;
input x_4464;
input x_4465;
input x_4466;
input x_4467;
input x_4468;
input x_4469;
input x_4470;
input x_4471;
input x_4472;
input x_4473;
input x_4474;
input x_4475;
input x_4476;
input x_4477;
input x_4478;
input x_4479;
input x_4480;
input x_4481;
input x_4482;
input x_4483;
input x_4484;
input x_4485;
input x_4486;
input x_4487;
input x_4488;
input x_4489;
input x_4490;
input x_4491;
input x_4492;
input x_4493;
input x_4494;
input x_4495;
input x_4496;
input x_4497;
input x_4498;
input x_4499;
input x_4500;
input x_4501;
input x_4502;
input x_4503;
input x_4504;
input x_4505;
input x_4506;
input x_4507;
input x_4508;
input x_4509;
input x_4510;
input x_4511;
input x_4512;
input x_4513;
input x_4514;
input x_4515;
input x_4516;
input x_4517;
input x_4518;
input x_4519;
input x_4520;
input x_4521;
input x_4522;
input x_4523;
input x_4524;
input x_4525;
input x_4526;
input x_4527;
input x_4528;
input x_4529;
input x_4530;
input x_4531;
input x_4532;
input x_4533;
input x_4534;
input x_4535;
input x_4536;
input x_4537;
input x_4538;
input x_4539;
input x_4540;
input x_4541;
input x_4542;
input x_4543;
input x_4544;
input x_4545;
input x_4546;
input x_4547;
input x_4548;
input x_4549;
input x_4550;
input x_4551;
input x_4552;
input x_4553;
input x_4554;
input x_4555;
input x_4556;
input x_4557;
input x_4558;
input x_4559;
input x_4560;
input x_4561;
input x_4562;
input x_4563;
input x_4564;
input x_4565;
input x_4566;
input x_4567;
input x_4568;
input x_4569;
input x_4570;
input x_4571;
input x_4572;
input x_4573;
input x_4574;
input x_4575;
input x_4576;
input x_4577;
input x_4578;
input x_4579;
input x_4580;
input x_4581;
input x_4582;
input x_4583;
input x_4584;
input x_4585;
input x_4586;
input x_4587;
input x_4588;
input x_4589;
input x_4590;
input x_4591;
input x_4592;
input x_4593;
input x_4594;
input x_4595;
input x_4596;
input x_4597;
input x_4598;
input x_4599;
input x_4600;
input x_4601;
input x_4602;
input x_4603;
input x_4604;
input x_4605;
input x_4606;
input x_4607;
input x_4608;
input x_4609;
input x_4610;
input x_4611;
input x_4612;
input x_4613;
input x_4614;
input x_4615;
input x_4616;
input x_4617;
input x_4618;
input x_4619;
input x_4620;
input x_4621;
input x_4622;
input x_4623;
input x_4624;
input x_4625;
input x_4626;
input x_4627;
input x_4628;
input x_4629;
input x_4630;
input x_4631;
input x_4632;
input x_4633;
input x_4634;
input x_4635;
input x_4636;
input x_4637;
input x_4638;
input x_4639;
input x_4640;
input x_4641;
input x_4642;
input x_4643;
input x_4644;
input x_4645;
input x_4646;
input x_4647;
input x_4648;
input x_4649;
input x_4650;
input x_4651;
input x_4652;
input x_4653;
input x_4654;
input x_4655;
input x_4656;
input x_4657;
input x_4658;
input x_4659;
input x_4660;
input x_4661;
input x_4662;
input x_4663;
input x_4664;
input x_4665;
input x_4666;
input x_4667;
input x_4668;
input x_4669;
input x_4670;
input x_4671;
input x_4672;
input x_4673;
input x_4674;
input x_4675;
input x_4676;
input x_4677;
input x_4678;
input x_4679;
input x_4680;
input x_4681;
input x_4682;
input x_4683;
input x_4684;
input x_4685;
input x_4686;
input x_4687;
input x_4688;
input x_4689;
input x_4690;
input x_4691;
input x_4692;
input x_4693;
input x_4694;
input x_4695;
input x_4696;
input x_4697;
input x_4698;
input x_4699;
input x_4700;
input x_4701;
input x_4702;
input x_4703;
input x_4704;
input x_4705;
input x_4706;
input x_4707;
input x_4708;
input x_4709;
input x_4710;
input x_4711;
input x_4712;
input x_4713;
input x_4714;
input x_4715;
input x_4716;
input x_4717;
input x_4718;
input x_4719;
input x_4720;
input x_4721;
input x_4722;
input x_4723;
input x_4724;
input x_4725;
input x_4726;
input x_4727;
input x_4728;
input x_4729;
input x_4730;
input x_4731;
input x_4732;
input x_4733;
input x_4734;
input x_4735;
input x_4736;
input x_4737;
input x_4738;
input x_4739;
input x_4740;
input x_4741;
input x_4742;
input x_4743;
input x_4744;
input x_4745;
input x_4746;
input x_4747;
input x_4748;
input x_4749;
input x_4750;
input x_4751;
input x_4752;
input x_4753;
input x_4754;
input x_4755;
input x_4756;
input x_4757;
input x_4758;
input x_4759;
input x_4760;
input x_4761;
input x_4762;
input x_4763;
input x_4764;
input x_4765;
input x_4766;
input x_4767;
input x_4768;
input x_4769;
input x_4770;
input x_4771;
input x_4772;
input x_4773;
input x_4774;
input x_4775;
input x_4776;
input x_4777;
input x_4778;
input x_4779;
input x_4780;
input x_4781;
input x_4782;
input x_4783;
input x_4784;
input x_4785;
input x_4786;
input x_4787;
input x_4788;
input x_4789;
input x_4790;
input x_4791;
input x_4792;
input x_4793;
input x_4794;
input x_4795;
input x_4796;
input x_4797;
input x_4798;
input x_4799;
input x_4800;
input x_4801;
input x_4802;
input x_4803;
input x_4804;
input x_4805;
input x_4806;
input x_4807;
input x_4808;
input x_4809;
input x_4810;
input x_4811;
input x_4812;
input x_4813;
input x_4814;
input x_4815;
input x_4816;
input x_4817;
input x_4818;
input x_4819;
input x_4820;
input x_4821;
input x_4822;
input x_4823;
input x_4824;
input x_4825;
input x_4826;
input x_4827;
input x_4828;
input x_4829;
input x_4830;
input x_4831;
input x_4832;
input x_4833;
input x_4834;
input x_4835;
input x_4836;
input x_4837;
input x_4838;
input x_4839;
input x_4840;
input x_4841;
input x_4842;
input x_4843;
input x_4844;
input x_4845;
input x_4846;
input x_4847;
input x_4848;
input x_4849;
input x_4850;
input x_4851;
input x_4852;
input x_4853;
input x_4854;
input x_4855;
input x_4856;
input x_4857;
input x_4858;
input x_4859;
input x_4860;
input x_4861;
input x_4862;
input x_4863;
input x_4864;
input x_4865;
input x_4866;
input x_4867;
input x_4868;
input x_4869;
input x_4870;
input x_4871;
input x_4872;
input x_4873;
input x_4874;
input x_4875;
input x_4876;
input x_4877;
input x_4878;
input x_4879;
input x_4880;
input x_4881;
input x_4882;
input x_4883;
input x_4884;
input x_4885;
input x_4886;
input x_4887;
input x_4888;
input x_4889;
input x_4890;
input x_4891;
input x_4892;
input x_4893;
input x_4894;
input x_4895;
input x_4896;
input x_4897;
input x_4898;
input x_4899;
input x_4900;
input x_4901;
input x_4902;
input x_4903;
input x_4904;
input x_4905;
input x_4906;
input x_4907;
input x_4908;
input x_4909;
input x_4910;
input x_4911;
input x_4912;
input x_4913;
input x_4914;
input x_4915;
input x_4916;
input x_4917;
input x_4918;
input x_4919;
input x_4920;
input x_4921;
input x_4922;
input x_4923;
input x_4924;
input x_4925;
input x_4926;
input x_4927;
input x_4928;
input x_4929;
input x_4930;
input x_4931;
input x_4932;
input x_4933;
input x_4934;
input x_4935;
input x_4936;
input x_4937;
input x_4938;
input x_4939;
input x_4940;
input x_4941;
input x_4942;
input x_4943;
input x_4944;
input x_4945;
input x_4946;
input x_4947;
input x_4948;
input x_4949;
input x_4950;
input x_4951;
input x_4952;
input x_4953;
input x_4954;
input x_4955;
input x_4956;
input x_4957;
input x_4958;
input x_4959;
input x_4960;
input x_4961;
input x_4962;
input x_4963;
input x_4964;
input x_4965;
input x_4966;
input x_4967;
input x_4968;
input x_4969;
input x_4970;
input x_4971;
input x_4972;
input x_4973;
input x_4974;
input x_4975;
input x_4976;
input x_4977;
input x_4978;
input x_4979;
input x_4980;
input x_4981;
input x_4982;
input x_4983;
input x_4984;
input x_4985;
input x_4986;
input x_4987;
input x_4988;
input x_4989;
input x_4990;
input x_4991;
input x_4992;
input x_4993;
input x_4994;
input x_4995;
input x_4996;
input x_4997;
input x_4998;
input x_4999;
input x_5000;
input x_5001;
input x_5002;
input x_5003;
input x_5004;
input x_5005;
input x_5006;
input x_5007;
input x_5008;
input x_5009;
input x_5010;
input x_5011;
input x_5012;
input x_5013;
input x_5014;
input x_5015;
input x_5016;
input x_5017;
input x_5018;
input x_5019;
input x_5020;
input x_5021;
input x_5022;
input x_5023;
input x_5024;
input x_5025;
input x_5026;
input x_5027;
input x_5028;
input x_5029;
input x_5030;
input x_5031;
input x_5032;
input x_5033;
input x_5034;
input x_5035;
input x_5036;
input x_5037;
input x_5038;
input x_5039;
input x_5040;
input x_5041;
input x_5042;
input x_5043;
input x_5044;
input x_5045;
input x_5046;
input x_5047;
input x_5048;
input x_5049;
input x_5050;
input x_5051;
input x_5052;
input x_5053;
input x_5054;
input x_5055;
input x_5056;
input x_5057;
input x_5058;
input x_5059;
input x_5060;
input x_5061;
input x_5062;
input x_5063;
input x_5064;
input x_5065;
input x_5066;
input x_5067;
input x_5068;
input x_5069;
input x_5070;
input x_5071;
input x_5072;
input x_5073;
input x_5074;
input x_5075;
input x_5076;
input x_5077;
input x_5078;
input x_5079;
input x_5080;
input x_5081;
input x_5082;
input x_5083;
input x_5084;
input x_5085;
input x_5086;
input x_5087;
input x_5088;
input x_5089;
input x_5090;
input x_5091;
input x_5092;
input x_5093;
input x_5094;
input x_5095;
input x_5096;
input x_5097;
input x_5098;
input x_5099;
input x_5100;
input x_5101;
input x_5102;
input x_5103;
input x_5104;
input x_5105;
input x_5106;
input x_5107;
input x_5108;
input x_5109;
input x_5110;
input x_5111;
input x_5112;
input x_5113;
input x_5114;
input x_5115;
input x_5116;
input x_5117;
input x_5118;
input x_5119;
input x_5120;
input x_5121;
input x_5122;
input x_5123;
input x_5124;
input x_5125;
input x_5126;
input x_5127;
input x_5128;
input x_5129;
input x_5130;
input x_5131;
input x_5132;
input x_5133;
input x_5134;
input x_5135;
input x_5136;
input x_5137;
input x_5138;
input x_5139;
input x_5140;
input x_5141;
input x_5142;
input x_5143;
input x_5144;
input x_5145;
input x_5146;
input x_5147;
input x_5148;
input x_5149;
input x_5150;
input x_5151;
input x_5152;
input x_5153;
input x_5154;
input x_5155;
input x_5156;
input x_5157;
input x_5158;
input x_5159;
input x_5160;
input x_5161;
input x_5162;
input x_5163;
input x_5164;
input x_5165;
input x_5166;
input x_5167;
input x_5168;
input x_5169;
input x_5170;
input x_5171;
input x_5172;
input x_5173;
input x_5174;
input x_5175;
input x_5176;
input x_5177;
input x_5178;
input x_5179;
input x_5180;
input x_5181;
input x_5182;
input x_5183;
input x_5184;
input x_5185;
input x_5186;
input x_5187;
input x_5188;
input x_5189;
input x_5190;
input x_5191;
input x_5192;
input x_5193;
input x_5194;
input x_5195;
input x_5196;
input x_5197;
input x_5198;
input x_5199;
input x_5200;
input x_5201;
input x_5202;
input x_5203;
input x_5204;
input x_5205;
input x_5206;
input x_5207;
input x_5208;
input x_5209;
input x_5210;
input x_5211;
input x_5212;
input x_5213;
input x_5214;
input x_5215;
input x_5216;
input x_5217;
input x_5218;
input x_5219;
input x_5220;
input x_5221;
input x_5222;
input x_5223;
input x_5224;
input x_5225;
input x_5226;
input x_5227;
input x_5228;
input x_5229;
input x_5230;
input x_5231;
input x_5232;
input x_5233;
input x_5234;
input x_5235;
input x_5236;
input x_5237;
input x_5238;
input x_5239;
input x_5240;
input x_5241;
input x_5242;
input x_5243;
input x_5244;
input x_5245;
input x_5246;
input x_5247;
input x_5248;
input x_5249;
input x_5250;
input x_5251;
input x_5252;
input x_5253;
input x_5254;
input x_5255;
input x_5256;
input x_5257;
input x_5258;
input x_5259;
input x_5260;
input x_5261;
input x_5262;
input x_5263;
input x_5264;
input x_5265;
input x_5266;
input x_5267;
input x_5268;
input x_5269;
input x_5270;
input x_5271;
input x_5272;
input x_5273;
input x_5274;
input x_5275;
input x_5276;
input x_5277;
input x_5278;
input x_5279;
input x_5280;
input x_5281;
input x_5282;
input x_5283;
input x_5284;
input x_5285;
input x_5286;
input x_5287;
input x_5288;
input x_5289;
input x_5290;
input x_5291;
input x_5292;
input x_5293;
input x_5294;
input x_5295;
input x_5296;
input x_5297;
input x_5298;
input x_5299;
input x_5300;
input x_5301;
input x_5302;
input x_5303;
input x_5304;
input x_5305;
input x_5306;
input x_5307;
input x_5308;
input x_5309;
input x_5310;
input x_5311;
input x_5312;
input x_5313;
input x_5314;
input x_5315;
input x_5316;
input x_5317;
input x_5318;
input x_5319;
input x_5320;
input x_5321;
input x_5322;
input x_5323;
input x_5324;
input x_5325;
input x_5326;
input x_5327;
input x_5328;
input x_5329;
input x_5330;
input x_5331;
input x_5332;
input x_5333;
input x_5334;
input x_5335;
input x_5336;
input x_5337;
input x_5338;
input x_5339;
input x_5340;
input x_5341;
input x_5342;
input x_5343;
input x_5344;
input x_5345;
input x_5346;
input x_5347;
input x_5348;
input x_5349;
input x_5350;
input x_5351;
input x_5352;
input x_5353;
input x_5354;
input x_5355;
input x_5356;
input x_5357;
input x_5358;
input x_5359;
input x_5360;
input x_5361;
input x_5362;
input x_5363;
input x_5364;
input x_5365;
input x_5366;
input x_5367;
input x_5368;
input x_5369;
input x_5370;
input x_5371;
input x_5372;
input x_5373;
input x_5374;
input x_5375;
input x_5376;
input x_5377;
input x_5378;
input x_5379;
input x_5380;
input x_5381;
input x_5382;
input x_5383;
input x_5384;
input x_5385;
input x_5386;
input x_5387;
input x_5388;
input x_5389;
input x_5390;
input x_5391;
input x_5392;
input x_5393;
input x_5394;
input x_5395;
input x_5396;
input x_5397;
input x_5398;
input x_5399;
input x_5400;
input x_5401;
input x_5402;
input x_5403;
input x_5404;
input x_5405;
input x_5406;
input x_5407;
input x_5408;
input x_5409;
input x_5410;
input x_5411;
input x_5412;
input x_5413;
input x_5414;
input x_5415;
input x_5416;
input x_5417;
input x_5418;
input x_5419;
input x_5420;
input x_5421;
input x_5422;
input x_5423;
input x_5424;
input x_5425;
input x_5426;
input x_5427;
input x_5428;
input x_5429;
input x_5430;
input x_5431;
input x_5432;
input x_5433;
input x_5434;
input x_5435;
input x_5436;
input x_5437;
input x_5438;
input x_5439;
input x_5440;
input x_5441;
input x_5442;
input x_5443;
input x_5444;
input x_5445;
input x_5446;
input x_5447;
input x_5448;
input x_5449;
input x_5450;
input x_5451;
input x_5452;
input x_5453;
input x_5454;
input x_5455;
input x_5456;
input x_5457;
input x_5458;
input x_5459;
input x_5460;
input x_5461;
input x_5462;
input x_5463;
input x_5464;
input x_5465;
input x_5466;
input x_5467;
input x_5468;
input x_5469;
input x_5470;
input x_5471;
input x_5472;
input x_5473;
input x_5474;
input x_5475;
input x_5476;
input x_5477;
input x_5478;
input x_5479;
input x_5480;
input x_5481;
input x_5482;
input x_5483;
input x_5484;
input x_5485;
input x_5486;
input x_5487;
input x_5488;
input x_5489;
input x_5490;
input x_5491;
input x_5492;
input x_5493;
input x_5494;
input x_5495;
input x_5496;
input x_5497;
input x_5498;
input x_5499;
input x_5500;
input x_5501;
input x_5502;
input x_5503;
input x_5504;
input x_5505;
input x_5506;
input x_5507;
input x_5508;
input x_5509;
input x_5510;
input x_5511;
input x_5512;
input x_5513;
input x_5514;
input x_5515;
input x_5516;
input x_5517;
input x_5518;
input x_5519;
input x_5520;
input x_5521;
input x_5522;
input x_5523;
input x_5524;
input x_5525;
input x_5526;
input x_5527;
input x_5528;
input x_5529;
input x_5530;
input x_5531;
input x_5532;
input x_5533;
input x_5534;
input x_5535;
input x_5536;
input x_5537;
input x_5538;
input x_5539;
input x_5540;
input x_5541;
input x_5542;
input x_5543;
input x_5544;
input x_5545;
input x_5546;
input x_5547;
input x_5548;
input x_5549;
input x_5550;
input x_5551;
input x_5552;
input x_5553;
input x_5554;
input x_5555;
input x_5556;
input x_5557;
input x_5558;
input x_5559;
input x_5560;
input x_5561;
input x_5562;
input x_5563;
input x_5564;
input x_5565;
input x_5566;
input x_5567;
input x_5568;
input x_5569;
input x_5570;
input x_5571;
input x_5572;
input x_5573;
input x_5574;
input x_5575;
input x_5576;
input x_5577;
input x_5578;
input x_5579;
input x_5580;
input x_5581;
input x_5582;
input x_5583;
input x_5584;
input x_5585;
input x_5586;
input x_5587;
input x_5588;
input x_5589;
input x_5590;
input x_5591;
input x_5592;
input x_5593;
input x_5594;
input x_5595;
input x_5596;
input x_5597;
input x_5598;
input x_5599;
input x_5600;
input x_5601;
input x_5602;
input x_5603;
input x_5604;
input x_5605;
input x_5606;
input x_5607;
input x_5608;
input x_5609;
input x_5610;
input x_5611;
input x_5612;
input x_5613;
input x_5614;
input x_5615;
input x_5616;
input x_5617;
input x_5618;
input x_5619;
input x_5620;
input x_5621;
input x_5622;
input x_5623;
input x_5624;
input x_5625;
input x_5626;
input x_5627;
input x_5628;
input x_5629;
input x_5630;
input x_5631;
input x_5632;
input x_5633;
input x_5634;
input x_5635;
input x_5636;
input x_5637;
input x_5638;
input x_5639;
input x_5640;
input x_5641;
input x_5642;
input x_5643;
input x_5644;
input x_5645;
input x_5646;
input x_5647;
input x_5648;
input x_5649;
input x_5650;
input x_5651;
input x_5652;
input x_5653;
input x_5654;
input x_5655;
input x_5656;
input x_5657;
input x_5658;
input x_5659;
input x_5660;
input x_5661;
input x_5662;
input x_5663;
input x_5664;
input x_5665;
input x_5666;
input x_5667;
input x_5668;
input x_5669;
input x_5670;
input x_5671;
input x_5672;
input x_5673;
input x_5674;
input x_5675;
input x_5676;
input x_5677;
input x_5678;
input x_5679;
input x_5680;
input x_5681;
input x_5682;
input x_5683;
input x_5684;
input x_5685;
input x_5686;
input x_5687;
input x_5688;
input x_5689;
input x_5690;
input x_5691;
input x_5692;
input x_5693;
input x_5694;
input x_5695;
input x_5696;
input x_5697;
input x_5698;
input x_5699;
input x_5700;
input x_5701;
input x_5702;
input x_5703;
input x_5704;
input x_5705;
input x_5706;
input x_5707;
input x_5708;
input x_5709;
input x_5710;
input x_5711;
input x_5712;
input x_5713;
input x_5714;
input x_5715;
input x_5716;
input x_5717;
input x_5718;
input x_5719;
input x_5720;
input x_5721;
input x_5722;
input x_5723;
input x_5724;
input x_5725;
input x_5726;
input x_5727;
input x_5728;
input x_5729;
input x_5730;
input x_5731;
input x_5732;
input x_5733;
input x_5734;
input x_5735;
input x_5736;
input x_5737;
input x_5738;
input x_5739;
input x_5740;
input x_5741;
input x_5742;
input x_5743;
input x_5744;
input x_5745;
input x_5746;
input x_5747;
input x_5748;
input x_5749;
input x_5750;
input x_5751;
input x_5752;
input x_5753;
input x_5754;
input x_5755;
input x_5756;
input x_5757;
input x_5758;
input x_5759;
input x_5760;
input x_5761;
input x_5762;
input x_5763;
input x_5764;
input x_5765;
input x_5766;
input x_5767;
input x_5768;
input x_5769;
input x_5770;
input x_5771;
input x_5772;
input x_5773;
input x_5774;
input x_5775;
input x_5776;
input x_5777;
input x_5778;
input x_5779;
input x_5780;
input x_5781;
input x_5782;
input x_5783;
input x_5784;
input x_5785;
input x_5786;
input x_5787;
input x_5788;
input x_5789;
input x_5790;
input x_5791;
input x_5792;
input x_5793;
input x_5794;
input x_5795;
input x_5796;
input x_5797;
input x_5798;
input x_5799;
input x_5800;
input x_5801;
input x_5802;
input x_5803;
input x_5804;
input x_5805;
input x_5806;
input x_5807;
input x_5808;
input x_5809;
input x_5810;
input x_5811;
input x_5812;
input x_5813;
input x_5814;
input x_5815;
input x_5816;
input x_5817;
input x_5818;
input x_5819;
input x_5820;
input x_5821;
input x_5822;
input x_5823;
input x_5824;
input x_5825;
input x_5826;
input x_5827;
input x_5828;
input x_5829;
input x_5830;
input x_5831;
input x_5832;
input x_5833;
input x_5834;
input x_5835;
input x_5836;
input x_5837;
input x_5838;
input x_5839;
input x_5840;
input x_5841;
input x_5842;
input x_5843;
input x_5844;
input x_5845;
input x_5846;
input x_5847;
input x_5848;
input x_5849;
input x_5850;
input x_5851;
input x_5852;
input x_5853;
input x_5854;
input x_5855;
input x_5856;
input x_5857;
input x_5858;
input x_5859;
input x_5860;
input x_5861;
input x_5862;
input x_5863;
input x_5864;
input x_5865;
input x_5866;
input x_5867;
input x_5868;
input x_5869;
input x_5870;
input x_5871;
input x_5872;
input x_5873;
input x_5874;
input x_5875;
input x_5876;
input x_5877;
input x_5878;
input x_5879;
input x_5880;
input x_5881;
input x_5882;
input x_5883;
input x_5884;
input x_5885;
input x_5886;
input x_5887;
input x_5888;
input x_5889;
input x_5890;
input x_5891;
input x_5892;
input x_5893;
input x_5894;
input x_5895;
input x_5896;
input x_5897;
input x_5898;
input x_5899;
input x_5900;
input x_5901;
input x_5902;
input x_5903;
input x_5904;
input x_5905;
input x_5906;
input x_5907;
input x_5908;
input x_5909;
input x_5910;
input x_5911;
input x_5912;
input x_5913;
input x_5914;
input x_5915;
input x_5916;
input x_5917;
input x_5918;
input x_5919;
input x_5920;
input x_5921;
input x_5922;
input x_5923;
input x_5924;
input x_5925;
input x_5926;
input x_5927;
input x_5928;
input x_5929;
input x_5930;
input x_5931;
input x_5932;
input x_5933;
input x_5934;
input x_5935;
input x_5936;
input x_5937;
input x_5938;
input x_5939;
input x_5940;
input x_5941;
input x_5942;
input x_5943;
input x_5944;
input x_5945;
input x_5946;
input x_5947;
input x_5948;
input x_5949;
input x_5950;
input x_5951;
input x_5952;
input x_5953;
input x_5954;
input x_5955;
input x_5956;
input x_5957;
input x_5958;
input x_5959;
input x_5960;
input x_5961;
input x_5962;
input x_5963;
input x_5964;
input x_5965;
input x_5966;
input x_5967;
input x_5968;
input x_5969;
input x_5970;
input x_5971;
input x_5972;
input x_5973;
input x_5974;
input x_5975;
input x_5976;
input x_5977;
input x_5978;
input x_5979;
input x_5980;
input x_5981;
input x_5982;
input x_5983;
input x_5984;
input x_5985;
input x_5986;
input x_5987;
input x_5988;
input x_5989;
input x_5990;
input x_5991;
input x_5992;
input x_5993;
input x_5994;
input x_5995;
input x_5996;
input x_5997;
input x_5998;
input x_5999;
input x_6000;
input x_6001;
input x_6002;
input x_6003;
input x_6004;
input x_6005;
input x_6006;
input x_6007;
input x_6008;
input x_6009;
input x_6010;
input x_6011;
input x_6012;
input x_6013;
input x_6014;
input x_6015;
input x_6016;
input x_6017;
input x_6018;
input x_6019;
input x_6020;
input x_6021;
input x_6022;
input x_6023;
input x_6024;
input x_6025;
input x_6026;
input x_6027;
input x_6028;
input x_6029;
input x_6030;
input x_6031;
input x_6032;
input x_6033;
input x_6034;
input x_6035;
input x_6036;
input x_6037;
input x_6038;
input x_6039;
input x_6040;
input x_6041;
input x_6042;
input x_6043;
input x_6044;
input x_6045;
input x_6046;
input x_6047;
input x_6048;
input x_6049;
input x_6050;
input x_6051;
input x_6052;
input x_6053;
input x_6054;
input x_6055;
input x_6056;
input x_6057;
input x_6058;
input x_6059;
input x_6060;
input x_6061;
input x_6062;
input x_6063;
input x_6064;
input x_6065;
input x_6066;
input x_6067;
input x_6068;
input x_6069;
input x_6070;
input x_6071;
input x_6072;
input x_6073;
input x_6074;
input x_6075;
input x_6076;
input x_6077;
input x_6078;
input x_6079;
input x_6080;
input x_6081;
input x_6082;
input x_6083;
input x_6084;
input x_6085;
input x_6086;
input x_6087;
input x_6088;
input x_6089;
input x_6090;
input x_6091;
input x_6092;
input x_6093;
input x_6094;
input x_6095;
input x_6096;
input x_6097;
input x_6098;
input x_6099;
input x_6100;
input x_6101;
input x_6102;
input x_6103;
input x_6104;
input x_6105;
input x_6106;
input x_6107;
input x_6108;
input x_6109;
input x_6110;
input x_6111;
input x_6112;
input x_6113;
input x_6114;
input x_6115;
input x_6116;
input x_6117;
input x_6118;
input x_6119;
input x_6120;
input x_6121;
input x_6122;
input x_6123;
input x_6124;
input x_6125;
input x_6126;
input x_6127;
input x_6128;
input x_6129;
input x_6130;
input x_6131;
input x_6132;
input x_6133;
input x_6134;
input x_6135;
input x_6136;
input x_6137;
input x_6138;
input x_6139;
input x_6140;
input x_6141;
input x_6142;
input x_6143;
input x_6144;
input x_6145;
input x_6146;
input x_6147;
input x_6148;
input x_6149;
input x_6150;
input x_6151;
input x_6152;
input x_6153;
input x_6154;
input x_6155;
input x_6156;
input x_6157;
input x_6158;
input x_6159;
input x_6160;
input x_6161;
input x_6162;
input x_6163;
input x_6164;
input x_6165;
input x_6166;
input x_6167;
input x_6168;
input x_6169;
input x_6170;
input x_6171;
input x_6172;
input x_6173;
input x_6174;
input x_6175;
input x_6176;
input x_6177;
input x_6178;
input x_6179;
input x_6180;
input x_6181;
input x_6182;
input x_6183;
input x_6184;
input x_6185;
input x_6186;
input x_6187;
input x_6188;
input x_6189;
input x_6190;
input x_6191;
input x_6192;
input x_6193;
input x_6194;
input x_6195;
input x_6196;
input x_6197;
input x_6198;
input x_6199;
input x_6200;
input x_6201;
input x_6202;
input x_6203;
input x_6204;
input x_6205;
input x_6206;
input x_6207;
input x_6208;
input x_6209;
input x_6210;
input x_6211;
input x_6212;
input x_6213;
input x_6214;
input x_6215;
input x_6216;
input x_6217;
input x_6218;
input x_6219;
input x_6220;
input x_6221;
input x_6222;
input x_6223;
input x_6224;
input x_6225;
input x_6226;
input x_6227;
input x_6228;
input x_6229;
input x_6230;
input x_6231;
input x_6232;
input x_6233;
input x_6234;
input x_6235;
input x_6236;
input x_6237;
input x_6238;
input x_6239;
input x_6240;
input x_6241;
input x_6242;
input x_6243;
input x_6244;
input x_6245;
input x_6246;
input x_6247;
input x_6248;
input x_6249;
input x_6250;
input x_6251;
input x_6252;
input x_6253;
input x_6254;
input x_6255;
input x_6256;
input x_6257;
input x_6258;
input x_6259;
input x_6260;
input x_6261;
input x_6262;
input x_6263;
input x_6264;
input x_6265;
input x_6266;
input x_6267;
input x_6268;
input x_6269;
input x_6270;
input x_6271;
input x_6272;
input x_6273;
input x_6274;
input x_6275;
input x_6276;
input x_6277;
input x_6278;
input x_6279;
input x_6280;
input x_6281;
input x_6282;
input x_6283;
input x_6284;
input x_6285;
input x_6286;
input x_6287;
input x_6288;
input x_6289;
input x_6290;
input x_6291;
input x_6292;
input x_6293;
input x_6294;
input x_6295;
input x_6296;
input x_6297;
input x_6298;
input x_6299;
input x_6300;
input x_6301;
input x_6302;
input x_6303;
input x_6304;
input x_6305;
input x_6306;
input x_6307;
input x_6308;
input x_6309;
input x_6310;
input x_6311;
input x_6312;
input x_6313;
input x_6314;
input x_6315;
input x_6316;
input x_6317;
input x_6318;
input x_6319;
input x_6320;
input x_6321;
input x_6322;
input x_6323;
input x_6324;
input x_6325;
input x_6326;
input x_6327;
input x_6328;
input x_6329;
input x_6330;
input x_6331;
input x_6332;
input x_6333;
input x_6334;
input x_6335;
input x_6336;
input x_6337;
input x_6338;
input x_6339;
input x_6340;
input x_6341;
input x_6342;
input x_6343;
input x_6344;
input x_6345;
input x_6346;
input x_6347;
input x_6348;
input x_6349;
input x_6350;
input x_6351;
input x_6352;
input x_6353;
input x_6354;
input x_6355;
input x_6356;
input x_6357;
input x_6358;
input x_6359;
input x_6360;
input x_6361;
input x_6362;
input x_6363;
input x_6364;
input x_6365;
input x_6366;
input x_6367;
input x_6368;
input x_6369;
input x_6370;
input x_6371;
input x_6372;
input x_6373;
input x_6374;
input x_6375;
input x_6376;
input x_6377;
input x_6378;
input x_6379;
input x_6380;
input x_6381;
input x_6382;
input x_6383;
input x_6384;
input x_6385;
input x_6386;
input x_6387;
input x_6388;
input x_6389;
input x_6390;
input x_6391;
input x_6392;
input x_6393;
input x_6394;
input x_6395;
input x_6396;
input x_6397;
input x_6398;
input x_6399;
input x_6400;
input x_6401;
input x_6402;
input x_6403;
input x_6404;
input x_6405;
input x_6406;
input x_6407;
input x_6408;
input x_6409;
input x_6410;
input x_6411;
input x_6412;
input x_6413;
input x_6414;
input x_6415;
input x_6416;
input x_6417;
input x_6418;
input x_6419;
input x_6420;
input x_6421;
input x_6422;
input x_6423;
input x_6424;
input x_6425;
input x_6426;
input x_6427;
input x_6428;
input x_6429;
input x_6430;
input x_6431;
input x_6432;
input x_6433;
input x_6434;
input x_6435;
input x_6436;
input x_6437;
input x_6438;
input x_6439;
input x_6440;
input x_6441;
input x_6442;
input x_6443;
input x_6444;
input x_6445;
input x_6446;
input x_6447;
input x_6448;
input x_6449;
input x_6450;
input x_6451;
input x_6452;
input x_6453;
input x_6454;
input x_6455;
input x_6456;
input x_6457;
input x_6458;
input x_6459;
input x_6460;
input x_6461;
input x_6462;
input x_6463;
input x_6464;
input x_6465;
input x_6466;
input x_6467;
input x_6468;
input x_6469;
input x_6470;
input x_6471;
input x_6472;
input x_6473;
input x_6474;
input x_6475;
input x_6476;
input x_6477;
input x_6478;
input x_6479;
input x_6480;
input x_6481;
input x_6482;
input x_6483;
input x_6484;
input x_6485;
input x_6486;
input x_6487;
input x_6488;
input x_6489;
input x_6490;
input x_6491;
input x_6492;
input x_6493;
input x_6494;
input x_6495;
input x_6496;
input x_6497;
input x_6498;
input x_6499;
input x_6500;
input x_6501;
input x_6502;
input x_6503;
input x_6504;
input x_6505;
input x_6506;
input x_6507;
input x_6508;
input x_6509;
input x_6510;
input x_6511;
input x_6512;
input x_6513;
input x_6514;
input x_6515;
input x_6516;
input x_6517;
input x_6518;
input x_6519;
input x_6520;
input x_6521;
input x_6522;
input x_6523;
input x_6524;
input x_6525;
input x_6526;
input x_6527;
input x_6528;
input x_6529;
input x_6530;
input x_6531;
input x_6532;
input x_6533;
input x_6534;
input x_6535;
input x_6536;
input x_6537;
input x_6538;
input x_6539;
input x_6540;
input x_6541;
input x_6542;
input x_6543;
input x_6544;
input x_6545;
input x_6546;
input x_6547;
input x_6548;
input x_6549;
input x_6550;
input x_6551;
input x_6552;
input x_6553;
input x_6554;
input x_6555;
input x_6556;
input x_6557;
input x_6558;
input x_6559;
input x_6560;
input x_6561;
input x_6562;
input x_6563;
input x_6564;
input x_6565;
input x_6566;
input x_6567;
input x_6568;
input x_6569;
input x_6570;
input x_6571;
input x_6572;
input x_6573;
input x_6574;
input x_6575;
input x_6576;
input x_6577;
input x_6578;
input x_6579;
input x_6580;
input x_6581;
input x_6582;
input x_6583;
input x_6584;
input x_6585;
input x_6586;
input x_6587;
input x_6588;
input x_6589;
input x_6590;
input x_6591;
input x_6592;
input x_6593;
input x_6594;
input x_6595;
input x_6596;
input x_6597;
input x_6598;
input x_6599;
input x_6600;
input x_6601;
input x_6602;
input x_6603;
input x_6604;
input x_6605;
input x_6606;
input x_6607;
input x_6608;
input x_6609;
input x_6610;
input x_6611;
input x_6612;
input x_6613;
input x_6614;
input x_6615;
input x_6616;
input x_6617;
input x_6618;
input x_6619;
input x_6620;
input x_6621;
input x_6622;
input x_6623;
input x_6624;
input x_6625;
input x_6626;
input x_6627;
input x_6628;
input x_6629;
input x_6630;
input x_6631;
input x_6632;
input x_6633;
input x_6634;
input x_6635;
input x_6636;
input x_6637;
input x_6638;
input x_6639;
input x_6640;
input x_6641;
input x_6642;
input x_6643;
input x_6644;
input x_6645;
input x_6646;
input x_6647;
input x_6648;
input x_6649;
input x_6650;
input x_6651;
input x_6652;
input x_6653;
input x_6654;
input x_6655;
input x_6656;
input x_6657;
input x_6658;
input x_6659;
input x_6660;
input x_6661;
input x_6662;
input x_6663;
input x_6664;
input x_6665;
input x_6666;
input x_6667;
input x_6668;
input x_6669;
input x_6670;
input x_6671;
input x_6672;
input x_6673;
input x_6674;
input x_6675;
input x_6676;
input x_6677;
input x_6678;
input x_6679;
input x_6680;
input x_6681;
input x_6682;
input x_6683;
input x_6684;
input x_6685;
input x_6686;
input x_6687;
input x_6688;
input x_6689;
input x_6690;
input x_6691;
input x_6692;
input x_6693;
input x_6694;
input x_6695;
input x_6696;
input x_6697;
input x_6698;
input x_6699;
input x_6700;
input x_6701;
input x_6702;
input x_6703;
input x_6704;
input x_6705;
input x_6706;
input x_6707;
input x_6708;
input x_6709;
input x_6710;
input x_6711;
input x_6712;
input x_6713;
input x_6714;
input x_6715;
input x_6716;
input x_6717;
input x_6718;
input x_6719;
input x_6720;
input x_6721;
input x_6722;
input x_6723;
input x_6724;
input x_6725;
input x_6726;
input x_6727;
input x_6728;
input x_6729;
input x_6730;
input x_6731;
input x_6732;
input x_6733;
input x_6734;
input x_6735;
input x_6736;
input x_6737;
input x_6738;
input x_6739;
input x_6740;
input x_6741;
input x_6742;
input x_6743;
input x_6744;
input x_6745;
input x_6746;
input x_6747;
input x_6748;
input x_6749;
input x_6750;
input x_6751;
input x_6752;
input x_6753;
input x_6754;
input x_6755;
input x_6756;
input x_6757;
input x_6758;
input x_6759;
input x_6760;
input x_6761;
input x_6762;
input x_6763;
input x_6764;
input x_6765;
input x_6766;
input x_6767;
input x_6768;
input x_6769;
input x_6770;
input x_6771;
input x_6772;
input x_6773;
input x_6774;
input x_6775;
input x_6776;
input x_6777;
input x_6778;
input x_6779;
input x_6780;
input x_6781;
input x_6782;
input x_6783;
input x_6784;
input x_6785;
input x_6786;
input x_6787;
input x_6788;
input x_6789;
input x_6790;
input x_6791;
input x_6792;
input x_6793;
input x_6794;
input x_6795;
input x_6796;
input x_6797;
input x_6798;
input x_6799;
input x_6800;
input x_6801;
input x_6802;
input x_6803;
input x_6804;
input x_6805;
input x_6806;
input x_6807;
input x_6808;
input x_6809;
input x_6810;
input x_6811;
input x_6812;
input x_6813;
input x_6814;
input x_6815;
input x_6816;
input x_6817;
input x_6818;
input x_6819;
input x_6820;
input x_6821;
input x_6822;
input x_6823;
input x_6824;
input x_6825;
input x_6826;
input x_6827;
input x_6828;
input x_6829;
input x_6830;
input x_6831;
input x_6832;
input x_6833;
input x_6834;
input x_6835;
input x_6836;
input x_6837;
input x_6838;
input x_6839;
input x_6840;
input x_6841;
input x_6842;
input x_6843;
input x_6844;
input x_6845;
input x_6846;
input x_6847;
input x_6848;
input x_6849;
input x_6850;
input x_6851;
input x_6852;
input x_6853;
input x_6854;
input x_6855;
input x_6856;
input x_6857;
input x_6858;
input x_6859;
input x_6860;
input x_6861;
input x_6862;
input x_6863;
input x_6864;
input x_6865;
input x_6866;
input x_6867;
input x_6868;
input x_6869;
input x_6870;
input x_6871;
input x_6872;
input x_6873;
input x_6874;
input x_6875;
input x_6876;
input x_6877;
input x_6878;
input x_6879;
input x_6880;
input x_6881;
input x_6882;
input x_6883;
input x_6884;
input x_6885;
input x_6886;
input x_6887;
input x_6888;
input x_6889;
input x_6890;
input x_6891;
input x_6892;
input x_6893;
input x_6894;
input x_6895;
input x_6896;
input x_6897;
input x_6898;
input x_6899;
input x_6900;
input x_6901;
input x_6902;
input x_6903;
input x_6904;
input x_6905;
input x_6906;
input x_6907;
input x_6908;
input x_6909;
input x_6910;
input x_6911;
input x_6912;
input x_6913;
input x_6914;
input x_6915;
input x_6916;
input x_6917;
input x_6918;
input x_6919;
input x_6920;
input x_6921;
input x_6922;
input x_6923;
input x_6924;
input x_6925;
input x_6926;
input x_6927;
input x_6928;
input x_6929;
input x_6930;
input x_6931;
input x_6932;
input x_6933;
input x_6934;
input x_6935;
input x_6936;
input x_6937;
input x_6938;
input x_6939;
input x_6940;
input x_6941;
input x_6942;
input x_6943;
input x_6944;
input x_6945;
input x_6946;
input x_6947;
input x_6948;
input x_6949;
input x_6950;
input x_6951;
input x_6952;
input x_6953;
input x_6954;
input x_6955;
input x_6956;
input x_6957;
input x_6958;
input x_6959;
input x_6960;
input x_6961;
input x_6962;
input x_6963;
input x_6964;
input x_6965;
input x_6966;
input x_6967;
input x_6968;
input x_6969;
input x_6970;
input x_6971;
input x_6972;
input x_6973;
input x_6974;
input x_6975;
input x_6976;
input x_6977;
input x_6978;
input x_6979;
input x_6980;
input x_6981;
input x_6982;
input x_6983;
input x_6984;
input x_6985;
input x_6986;
input x_6987;
input x_6988;
input x_6989;
input x_6990;
input x_6991;
input x_6992;
input x_6993;
input x_6994;
input x_6995;
input x_6996;
input x_6997;
input x_6998;
input x_6999;
input x_7000;
input x_7001;
input x_7002;
input x_7003;
input x_7004;
input x_7005;
input x_7006;
input x_7007;
input x_7008;
input x_7009;
input x_7010;
input x_7011;
input x_7012;
input x_7013;
input x_7014;
input x_7015;
input x_7016;
input x_7017;
input x_7018;
input x_7019;
input x_7020;
input x_7021;
input x_7022;
input x_7023;
input x_7024;
input x_7025;
input x_7026;
input x_7027;
input x_7028;
input x_7029;
input x_7030;
input x_7031;
input x_7032;
input x_7033;
input x_7034;
input x_7035;
input x_7036;
input x_7037;
input x_7038;
input x_7039;
input x_7040;
input x_7041;
input x_7042;
input x_7043;
input x_7044;
input x_7045;
input x_7046;
input x_7047;
input x_7048;
input x_7049;
input x_7050;
input x_7051;
input x_7052;
input x_7053;
input x_7054;
input x_7055;
input x_7056;
input x_7057;
input x_7058;
input x_7059;
input x_7060;
input x_7061;
input x_7062;
input x_7063;
input x_7064;
input x_7065;
input x_7066;
input x_7067;
input x_7068;
input x_7069;
input x_7070;
input x_7071;
input x_7072;
input x_7073;
input x_7074;
input x_7075;
input x_7076;
input x_7077;
input x_7078;
input x_7079;
input x_7080;
input x_7081;
input x_7082;
input x_7083;
input x_7084;
input x_7085;
input x_7086;
input x_7087;
input x_7088;
input x_7089;
input x_7090;
input x_7091;
input x_7092;
input x_7093;
input x_7094;
input x_7095;
input x_7096;
input x_7097;
input x_7098;
input x_7099;
input x_7100;
input x_7101;
input x_7102;
input x_7103;
input x_7104;
input x_7105;
input x_7106;
input x_7107;
input x_7108;
input x_7109;
input x_7110;
input x_7111;
input x_7112;
input x_7113;
input x_7114;
input x_7115;
input x_7116;
input x_7117;
input x_7118;
input x_7119;
input x_7120;
input x_7121;
input x_7122;
input x_7123;
input x_7124;
input x_7125;
input x_7126;
input x_7127;
input x_7128;
input x_7129;
input x_7130;
input x_7131;
input x_7132;
input x_7133;
input x_7134;
input x_7135;
input x_7136;
input x_7137;
input x_7138;
input x_7139;
input x_7140;
input x_7141;
input x_7142;
input x_7143;
input x_7144;
input x_7145;
input x_7146;
input x_7147;
input x_7148;
input x_7149;
input x_7150;
input x_7151;
input x_7152;
input x_7153;
input x_7154;
input x_7155;
input x_7156;
input x_7157;
input x_7158;
input x_7159;
input x_7160;
input x_7161;
input x_7162;
input x_7163;
input x_7164;
input x_7165;
input x_7166;
input x_7167;
input x_7168;
input x_7169;
input x_7170;
input x_7171;
input x_7172;
input x_7173;
input x_7174;
input x_7175;
input x_7176;
input x_7177;
input x_7178;
input x_7179;
input x_7180;
input x_7181;
input x_7182;
input x_7183;
input x_7184;
input x_7185;
input x_7186;
input x_7187;
input x_7188;
input x_7189;
input x_7190;
input x_7191;
input x_7192;
input x_7193;
input x_7194;
input x_7195;
input x_7196;
input x_7197;
input x_7198;
input x_7199;
input x_7200;
input x_7201;
input x_7202;
input x_7203;
input x_7204;
input x_7205;
input x_7206;
input x_7207;
input x_7208;
input x_7209;
input x_7210;
input x_7211;
input x_7212;
input x_7213;
input x_7214;
input x_7215;
input x_7216;
input x_7217;
input x_7218;
input x_7219;
input x_7220;
input x_7221;
input x_7222;
input x_7223;
input x_7224;
input x_7225;
input x_7226;
input x_7227;
input x_7228;
input x_7229;
input x_7230;
input x_7231;
input x_7232;
input x_7233;
input x_7234;
input x_7235;
input x_7236;
input x_7237;
input x_7238;
input x_7239;
input x_7240;
input x_7241;
input x_7242;
input x_7243;
input x_7244;
input x_7245;
input x_7246;
input x_7247;
input x_7248;
input x_7249;
input x_7250;
input x_7251;
input x_7252;
input x_7253;
input x_7254;
input x_7255;
input x_7256;
input x_7257;
input x_7258;
input x_7259;
input x_7260;
input x_7261;
input x_7262;
input x_7263;
input x_7264;
input x_7265;
input x_7266;
input x_7267;
input x_7268;
input x_7269;
input x_7270;
input x_7271;
input x_7272;
input x_7273;
input x_7274;
input x_7275;
input x_7276;
input x_7277;
input x_7278;
input x_7279;
input x_7280;
input x_7281;
input x_7282;
input x_7283;
input x_7284;
input x_7285;
input x_7286;
input x_7287;
input x_7288;
input x_7289;
input x_7290;
input x_7291;
input x_7292;
input x_7293;
input x_7294;
input x_7295;
input x_7296;
input x_7297;
input x_7298;
input x_7299;
input x_7300;
input x_7301;
input x_7302;
input x_7303;
input x_7304;
input x_7305;
input x_7306;
input x_7307;
input x_7308;
input x_7309;
input x_7310;
input x_7311;
input x_7312;
input x_7313;
input x_7314;
input x_7315;
input x_7316;
input x_7317;
input x_7318;
input x_7319;
input x_7320;
input x_7321;
input x_7322;
input x_7323;
input x_7324;
input x_7325;
input x_7326;
input x_7327;
input x_7328;
input x_7329;
input x_7330;
input x_7331;
input x_7332;
input x_7333;
input x_7334;
input x_7335;
input x_7336;
input x_7337;
input x_7338;
input x_7339;
input x_7340;
input x_7341;
input x_7342;
input x_7343;
input x_7344;
input x_7345;
input x_7346;
input x_7347;
input x_7348;
input x_7349;
input x_7350;
input x_7351;
input x_7352;
input x_7353;
input x_7354;
input x_7355;
input x_7356;
input x_7357;
input x_7358;
input x_7359;
input x_7360;
input x_7361;
input x_7362;
input x_7363;
input x_7364;
input x_7365;
input x_7366;
input x_7367;
input x_7368;
input x_7369;
input x_7370;
input x_7371;
input x_7372;
input x_7373;
input x_7374;
input x_7375;
input x_7376;
input x_7377;
input x_7378;
input x_7379;
input x_7380;
input x_7381;
input x_7382;
input x_7383;
input x_7384;
input x_7385;
input x_7386;
input x_7387;
input x_7388;
input x_7389;
input x_7390;
input x_7391;
input x_7392;
input x_7393;
input x_7394;
input x_7395;
input x_7396;
input x_7397;
input x_7398;
input x_7399;
input x_7400;
input x_7401;
input x_7402;
input x_7403;
input x_7404;
input x_7405;
input x_7406;
input x_7407;
input x_7408;
input x_7409;
input x_7410;
input x_7411;
input x_7412;
input x_7413;
input x_7414;
input x_7415;
input x_7416;
input x_7417;
input x_7418;
input x_7419;
input x_7420;
input x_7421;
input x_7422;
input x_7423;
input x_7424;
input x_7425;
input x_7426;
input x_7427;
input x_7428;
input x_7429;
input x_7430;
input x_7431;
input x_7432;
input x_7433;
input x_7434;
input x_7435;
input x_7436;
input x_7437;
input x_7438;
input x_7439;
input x_7440;
input x_7441;
input x_7442;
input x_7443;
input x_7444;
input x_7445;
input x_7446;
input x_7447;
input x_7448;
input x_7449;
input x_7450;
input x_7451;
input x_7452;
input x_7453;
input x_7454;
input x_7455;
input x_7456;
input x_7457;
input x_7458;
input x_7459;
input x_7460;
input x_7461;
input x_7462;
input x_7463;
input x_7464;
input x_7465;
input x_7466;
input x_7467;
input x_7468;
input x_7469;
input x_7470;
input x_7471;
input x_7472;
input x_7473;
input x_7474;
input x_7475;
input x_7476;
input x_7477;
input x_7478;
input x_7479;
input x_7480;
input x_7481;
input x_7482;
input x_7483;
input x_7484;
input x_7485;
input x_7486;
input x_7487;
input x_7488;
input x_7489;
input x_7490;
input x_7491;
input x_7492;
input x_7493;
input x_7494;
input x_7495;
input x_7496;
input x_7497;
input x_7498;
input x_7499;
input x_7500;
input x_7501;
input x_7502;
input x_7503;
input x_7504;
input x_7505;
input x_7506;
input x_7507;
input x_7508;
input x_7509;
input x_7510;
input x_7511;
input x_7512;
input x_7513;
input x_7514;
input x_7515;
input x_7516;
input x_7517;
input x_7518;
input x_7519;
input x_7520;
input x_7521;
input x_7522;
input x_7523;
input x_7524;
input x_7525;
input x_7526;
input x_7527;
input x_7528;
input x_7529;
input x_7530;
input x_7531;
input x_7532;
input x_7533;
input x_7534;
input x_7535;
input x_7536;
input x_7537;
input x_7538;
input x_7539;
input x_7540;
input x_7541;
input x_7542;
input x_7543;
input x_7544;
input x_7545;
input x_7546;
input x_7547;
input x_7548;
input x_7549;
input x_7550;
input x_7551;
input x_7552;
input x_7553;
input x_7554;
input x_7555;
input x_7556;
input x_7557;
input x_7558;
input x_7559;
input x_7560;
input x_7561;
input x_7562;
input x_7563;
input x_7564;
input x_7565;
input x_7566;
input x_7567;
input x_7568;
input x_7569;
input x_7570;
input x_7571;
input x_7572;
input x_7573;
input x_7574;
input x_7575;
input x_7576;
input x_7577;
input x_7578;
input x_7579;
input x_7580;
input x_7581;
input x_7582;
input x_7583;
input x_7584;
input x_7585;
input x_7586;
input x_7587;
input x_7588;
input x_7589;
input x_7590;
input x_7591;
input x_7592;
input x_7593;
input x_7594;
input x_7595;
input x_7596;
input x_7597;
input x_7598;
input x_7599;
input x_7600;
input x_7601;
input x_7602;
input x_7603;
input x_7604;
input x_7605;
input x_7606;
input x_7607;
input x_7608;
input x_7609;
input x_7610;
input x_7611;
input x_7612;
input x_7613;
input x_7614;
input x_7615;
input x_7616;
input x_7617;
input x_7618;
input x_7619;
input x_7620;
input x_7621;
input x_7622;
input x_7623;
input x_7624;
input x_7625;
input x_7626;
input x_7627;
input x_7628;
input x_7629;
input x_7630;
input x_7631;
input x_7632;
input x_7633;
input x_7634;
input x_7635;
input x_7636;
input x_7637;
input x_7638;
input x_7639;
input x_7640;
input x_7641;
input x_7642;
input x_7643;
input x_7644;
input x_7645;
input x_7646;
input x_7647;
input x_7648;
input x_7649;
input x_7650;
input x_7651;
input x_7652;
input x_7653;
input x_7654;
input x_7655;
input x_7656;
input x_7657;
input x_7658;
input x_7659;
input x_7660;
input x_7661;
input x_7662;
input x_7663;
input x_7664;
input x_7665;
input x_7666;
input x_7667;
input x_7668;
input x_7669;
input x_7670;
input x_7671;
input x_7672;
input x_7673;
input x_7674;
input x_7675;
input x_7676;
input x_7677;
input x_7678;
input x_7679;
input x_7680;
input x_7681;
input x_7682;
input x_7683;
input x_7684;
input x_7685;
input x_7686;
input x_7687;
input x_7688;
input x_7689;
input x_7690;
input x_7691;
input x_7692;
input x_7693;
input x_7694;
input x_7695;
input x_7696;
input x_7697;
input x_7698;
input x_7699;
input x_7700;
input x_7701;
input x_7702;
input x_7703;
input x_7704;
input x_7705;
input x_7706;
input x_7707;
input x_7708;
input x_7709;
input x_7710;
input x_7711;
input x_7712;
input x_7713;
input x_7714;
input x_7715;
input x_7716;
input x_7717;
input x_7718;
input x_7719;
input x_7720;
input x_7721;
input x_7722;
input x_7723;
input x_7724;
input x_7725;
input x_7726;
input x_7727;
input x_7728;
input x_7729;
input x_7730;
input x_7731;
input x_7732;
input x_7733;
input x_7734;
input x_7735;
input x_7736;
input x_7737;
input x_7738;
input x_7739;
input x_7740;
input x_7741;
input x_7742;
input x_7743;
input x_7744;
input x_7745;
input x_7746;
input x_7747;
input x_7748;
input x_7749;
input x_7750;
input x_7751;
input x_7752;
input x_7753;
input x_7754;
input x_7755;
input x_7756;
input x_7757;
input x_7758;
input x_7759;
input x_7760;
input x_7761;
input x_7762;
input x_7763;
input x_7764;
input x_7765;
input x_7766;
input x_7767;
input x_7768;
input x_7769;
input x_7770;
input x_7771;
input x_7772;
input x_7773;
input x_7774;
input x_7775;
input x_7776;
input x_7777;
input x_7778;
input x_7779;
input x_7780;
input x_7781;
input x_7782;
input x_7783;
input x_7784;
input x_7785;
input x_7786;
input x_7787;
input x_7788;
input x_7789;
input x_7790;
input x_7791;
input x_7792;
input x_7793;
input x_7794;
input x_7795;
input x_7796;
input x_7797;
input x_7798;
input x_7799;
input x_7800;
input x_7801;
input x_7802;
input x_7803;
input x_7804;
input x_7805;
input x_7806;
input x_7807;
input x_7808;
input x_7809;
input x_7810;
input x_7811;
input x_7812;
input x_7813;
input x_7814;
input x_7815;
input x_7816;
input x_7817;
input x_7818;
input x_7819;
input x_7820;
input x_7821;
input x_7822;
input x_7823;
input x_7824;
input x_7825;
input x_7826;
input x_7827;
input x_7828;
input x_7829;
input x_7830;
input x_7831;
input x_7832;
input x_7833;
input x_7834;
input x_7835;
input x_7836;
input x_7837;
input x_7838;
input x_7839;
input x_7840;
input x_7841;
input x_7842;
input x_7843;
input x_7844;
input x_7845;
input x_7846;
input x_7847;
input x_7848;
input x_7849;
input x_7850;
input x_7851;
input x_7852;
input x_7853;
input x_7854;
input x_7855;
input x_7856;
input x_7857;
input x_7858;
input x_7859;
input x_7860;
input x_7861;
input x_7862;
input x_7863;
input x_7864;
input x_7865;
input x_7866;
input x_7867;
input x_7868;
input x_7869;
input x_7870;
input x_7871;
input x_7872;
input x_7873;
input x_7874;
input x_7875;
input x_7876;
input x_7877;
input x_7878;
input x_7879;
input x_7880;
input x_7881;
input x_7882;
input x_7883;
input x_7884;
input x_7885;
input x_7886;
input x_7887;
input x_7888;
input x_7889;
input x_7890;
input x_7891;
input x_7892;
input x_7893;
input x_7894;
input x_7895;
input x_7896;
input x_7897;
input x_7898;
input x_7899;
input x_7900;
input x_7901;
input x_7902;
input x_7903;
input x_7904;
input x_7905;
input x_7906;
input x_7907;
input x_7908;
input x_7909;
input x_7910;
input x_7911;
input x_7912;
input x_7913;
input x_7914;
input x_7915;
input x_7916;
input x_7917;
input x_7918;
input x_7919;
input x_7920;
input x_7921;
input x_7922;
input x_7923;
input x_7924;
input x_7925;
input x_7926;
input x_7927;
input x_7928;
input x_7929;
input x_7930;
input x_7931;
input x_7932;
input x_7933;
input x_7934;
input x_7935;
input x_7936;
input x_7937;
input x_7938;
input x_7939;
input x_7940;
input x_7941;
input x_7942;
input x_7943;
input x_7944;
input x_7945;
input x_7946;
input x_7947;
input x_7948;
input x_7949;
input x_7950;
input x_7951;
input x_7952;
input x_7953;
input x_7954;
input x_7955;
input x_7956;
input x_7957;
input x_7958;
input x_7959;
input x_7960;
input x_7961;
input x_7962;
input x_7963;
input x_7964;
input x_7965;
input x_7966;
input x_7967;
input x_7968;
input x_7969;
input x_7970;
input x_7971;
input x_7972;
input x_7973;
input x_7974;
input x_7975;
input x_7976;
input x_7977;
input x_7978;
input x_7979;
input x_7980;
input x_7981;
input x_7982;
input x_7983;
input x_7984;
input x_7985;
input x_7986;
input x_7987;
input x_7988;
input x_7989;
input x_7990;
input x_7991;
input x_7992;
input x_7993;
input x_7994;
input x_7995;
input x_7996;
input x_7997;
input x_7998;
input x_7999;
input x_8000;
input x_8001;
input x_8002;
input x_8003;
input x_8004;
input x_8005;
input x_8006;
input x_8007;
input x_8008;
input x_8009;
input x_8010;
input x_8011;
input x_8012;
input x_8013;
input x_8014;
input x_8015;
input x_8016;
input x_8017;
input x_8018;
input x_8019;
input x_8020;
input x_8021;
input x_8022;
input x_8023;
input x_8024;
input x_8025;
input x_8026;
input x_8027;
input x_8028;
input x_8029;
input x_8030;
input x_8031;
input x_8032;
input x_8033;
input x_8034;
input x_8035;
input x_8036;
input x_8037;
input x_8038;
input x_8039;
input x_8040;
input x_8041;
input x_8042;
input x_8043;
input x_8044;
input x_8045;
input x_8046;
input x_8047;
input x_8048;
input x_8049;
input x_8050;
input x_8051;
input x_8052;
input x_8053;
input x_8054;
input x_8055;
input x_8056;
input x_8057;
input x_8058;
input x_8059;
input x_8060;
input x_8061;
input x_8062;
input x_8063;
input x_8064;
input x_8065;
input x_8066;
input x_8067;
input x_8068;
input x_8069;
input x_8070;
input x_8071;
input x_8072;
input x_8073;
input x_8074;
input x_8075;
input x_8076;
input x_8077;
input x_8078;
input x_8079;
input x_8080;
input x_8081;
input x_8082;
input x_8083;
input x_8084;
input x_8085;
input x_8086;
input x_8087;
input x_8088;
input x_8089;
input x_8090;
input x_8091;
input x_8092;
input x_8093;
input x_8094;
input x_8095;
input x_8096;
input x_8097;
input x_8098;
input x_8099;
input x_8100;
input x_8101;
input x_8102;
input x_8103;
input x_8104;
input x_8105;
input x_8106;
input x_8107;
input x_8108;
input x_8109;
input x_8110;
input x_8111;
input x_8112;
input x_8113;
input x_8114;
input x_8115;
input x_8116;
input x_8117;
input x_8118;
input x_8119;
input x_8120;
input x_8121;
input x_8122;
input x_8123;
input x_8124;
input x_8125;
input x_8126;
input x_8127;
input x_8128;
input x_8129;
input x_8130;
input x_8131;
input x_8132;
input x_8133;
input x_8134;
input x_8135;
input x_8136;
input x_8137;
input x_8138;
input x_8139;
input x_8140;
input x_8141;
input x_8142;
input x_8143;
input x_8144;
input x_8145;
input x_8146;
input x_8147;
input x_8148;
input x_8149;
input x_8150;
input x_8151;
input x_8152;
input x_8153;
input x_8154;
input x_8155;
input x_8156;
input x_8157;
input x_8158;
input x_8159;
input x_8160;
input x_8161;
input x_8162;
input x_8163;
input x_8164;
input x_8165;
input x_8166;
input x_8167;
input x_8168;
input x_8169;
input x_8170;
input x_8171;
input x_8172;
input x_8173;
input x_8174;
input x_8175;
input x_8176;
input x_8177;
input x_8178;
input x_8179;
input x_8180;
input x_8181;
input x_8182;
input x_8183;
input x_8184;
input x_8185;
input x_8186;
input x_8187;
input x_8188;
input x_8189;
input x_8190;
input x_8191;
input x_8192;
input x_8193;
input x_8194;
input x_8195;
input x_8196;
input x_8197;
input x_8198;
input x_8199;
input x_8200;
input x_8201;
input x_8202;
input x_8203;
input x_8204;
input x_8205;
input x_8206;
input x_8207;
input x_8208;
input x_8209;
input x_8210;
input x_8211;
input x_8212;
input x_8213;
input x_8214;
input x_8215;
input x_8216;
input x_8217;
input x_8218;
input x_8219;
input x_8220;
input x_8221;
input x_8222;
input x_8223;
input x_8224;
input x_8225;
input x_8226;
input x_8227;
input x_8228;
input x_8229;
input x_8230;
input x_8231;
input x_8232;
input x_8233;
input x_8234;
input x_8235;
input x_8236;
input x_8237;
input x_8238;
input x_8239;
input x_8240;
input x_8241;
input x_8242;
input x_8243;
input x_8244;
input x_8245;
input x_8246;
input x_8247;
input x_8248;
input x_8249;
input x_8250;
input x_8251;
input x_8252;
input x_8253;
input x_8254;
input x_8255;
input x_8256;
input x_8257;
input x_8258;
input x_8259;
input x_8260;
input x_8261;
input x_8262;
input x_8263;
input x_8264;
input x_8265;
input x_8266;
input x_8267;
input x_8268;
input x_8269;
input x_8270;
input x_8271;
input x_8272;
input x_8273;
input x_8274;
input x_8275;
input x_8276;
input x_8277;
input x_8278;
input x_8279;
input x_8280;
input x_8281;
input x_8282;
input x_8283;
input x_8284;
input x_8285;
input x_8286;
input x_8287;
input x_8288;
input x_8289;
input x_8290;
input x_8291;
input x_8292;
input x_8293;
input x_8294;
input x_8295;
input x_8296;
input x_8297;
input x_8298;
input x_8299;
input x_8300;
input x_8301;
input x_8302;
input x_8303;
input x_8304;
input x_8305;
input x_8306;
input x_8307;
input x_8308;
input x_8309;
input x_8310;
input x_8311;
input x_8312;
input x_8313;
input x_8314;
input x_8315;
input x_8316;
input x_8317;
input x_8318;
input x_8319;
input x_8320;
input x_8321;
input x_8322;
input x_8323;
input x_8324;
input x_8325;
input x_8326;
input x_8327;
input x_8328;
input x_8329;
input x_8330;
input x_8331;
input x_8332;
input x_8333;
input x_8334;
input x_8335;
input x_8336;
input x_8337;
input x_8338;
input x_8339;
input x_8340;
input x_8341;
input x_8342;
input x_8343;
input x_8344;
input x_8345;
input x_8346;
input x_8347;
input x_8348;
input x_8349;
input x_8350;
input x_8351;
input x_8352;
input x_8353;
input x_8354;
input x_8355;
input x_8356;
input x_8357;
input x_8358;
input x_8359;
input x_8360;
input x_8361;
input x_8362;
input x_8363;
input x_8364;
input x_8365;
input x_8366;
input x_8367;
input x_8368;
input x_8369;
input x_8370;
input x_8371;
input x_8372;
input x_8373;
input x_8374;
input x_8375;
input x_8376;
input x_8377;
input x_8378;
input x_8379;
input x_8380;
input x_8381;
input x_8382;
input x_8383;
input x_8384;
input x_8385;
input x_8386;
input x_8387;
input x_8388;
input x_8389;
input x_8390;
input x_8391;
input x_8392;
input x_8393;
input x_8394;
input x_8395;
input x_8396;
input x_8397;
input x_8398;
input x_8399;
input x_8400;
input x_8401;
input x_8402;
input x_8403;
input x_8404;
input x_8405;
input x_8406;
input x_8407;
input x_8408;
input x_8409;
input x_8410;
input x_8411;
input x_8412;
input x_8413;
input x_8414;
input x_8415;
input x_8416;
input x_8417;
input x_8418;
input x_8419;
input x_8420;
input x_8421;
input x_8422;
input x_8423;
input x_8424;
input x_8425;
input x_8426;
input x_8427;
input x_8428;
input x_8429;
input x_8430;
input x_8431;
input x_8432;
input x_8433;
input x_8434;
input x_8435;
input x_8436;
input x_8437;
input x_8438;
input x_8439;
input x_8440;
input x_8441;
input x_8442;
input x_8443;
input x_8444;
input x_8445;
input x_8446;
input x_8447;
input x_8448;
input x_8449;
input x_8450;
input x_8451;
input x_8452;
input x_8453;
input x_8454;
input x_8455;
input x_8456;
input x_8457;
input x_8458;
input x_8459;
input x_8460;
input x_8461;
input x_8462;
input x_8463;
input x_8464;
input x_8465;
input x_8466;
input x_8467;
input x_8468;
input x_8469;
input x_8470;
input x_8471;
input x_8472;
input x_8473;
input x_8474;
input x_8475;
input x_8476;
input x_8477;
input x_8478;
input x_8479;
input x_8480;
input x_8481;
input x_8482;
input x_8483;
input x_8484;
input x_8485;
input x_8486;
input x_8487;
input x_8488;
input x_8489;
input x_8490;
input x_8491;
input x_8492;
input x_8493;
input x_8494;
input x_8495;
input x_8496;
input x_8497;
input x_8498;
input x_8499;
input x_8500;
input x_8501;
input x_8502;
input x_8503;
input x_8504;
input x_8505;
input x_8506;
input x_8507;
input x_8508;
input x_8509;
input x_8510;
input x_8511;
input x_8512;
input x_8513;
input x_8514;
input x_8515;
input x_8516;
input x_8517;
input x_8518;
input x_8519;
input x_8520;
input x_8521;
input x_8522;
input x_8523;
input x_8524;
input x_8525;
input x_8526;
input x_8527;
input x_8528;
input x_8529;
input x_8530;
input x_8531;
input x_8532;
input x_8533;
input x_8534;
input x_8535;
input x_8536;
input x_8537;
input x_8538;
input x_8539;
input x_8540;
input x_8541;
input x_8542;
input x_8543;
input x_8544;
input x_8545;
input x_8546;
input x_8547;
input x_8548;
input x_8549;
input x_8550;
input x_8551;
input x_8552;
input x_8553;
input x_8554;
input x_8555;
input x_8556;
input x_8557;
input x_8558;
input x_8559;
input x_8560;
input x_8561;
input x_8562;
input x_8563;
input x_8564;
input x_8565;
input x_8566;
input x_8567;
input x_8568;
input x_8569;
input x_8570;
input x_8571;
input x_8572;
input x_8573;
input x_8574;
input x_8575;
input x_8576;
input x_8577;
input x_8578;
input x_8579;
input x_8580;
input x_8581;
input x_8582;
input x_8583;
input x_8584;
input x_8585;
input x_8586;
input x_8587;
input x_8588;
input x_8589;
input x_8590;
input x_8591;
input x_8592;
input x_8593;
input x_8594;
input x_8595;
input x_8596;
input x_8597;
input x_8598;
input x_8599;
input x_8600;
input x_8601;
input x_8602;
input x_8603;
input x_8604;
input x_8605;
input x_8606;
input x_8607;
input x_8608;
input x_8609;
input x_8610;
input x_8611;
input x_8612;
input x_8613;
input x_8614;
input x_8615;
input x_8616;
input x_8617;
input x_8618;
input x_8619;
input x_8620;
input x_8621;
input x_8622;
input x_8623;
input x_8624;
input x_8625;
input x_8626;
input x_8627;
input x_8628;
input x_8629;
input x_8630;
input x_8631;
input x_8632;
input x_8633;
input x_8634;
input x_8635;
input x_8636;
input x_8637;
input x_8638;
input x_8639;
input x_8640;
input x_8641;
input x_8642;
input x_8643;
input x_8644;
input x_8645;
input x_8646;
input x_8647;
input x_8648;
input x_8649;
input x_8650;
input x_8651;
input x_8652;
input x_8653;
input x_8654;
input x_8655;
input x_8656;
input x_8657;
input x_8658;
input x_8659;
input x_8660;
input x_8661;
input x_8662;
input x_8663;
input x_8664;
input x_8665;
input x_8666;
input x_8667;
input x_8668;
input x_8669;
input x_8670;
input x_8671;
input x_8672;
input x_8673;
input x_8674;
input x_8675;
input x_8676;
input x_8677;
input x_8678;
input x_8679;
input x_8680;
input x_8681;
input x_8682;
input x_8683;
input x_8684;
input x_8685;
input x_8686;
input x_8687;
input x_8688;
input x_8689;
input x_8690;
input x_8691;
input x_8692;
input x_8693;
input x_8694;
input x_8695;
input x_8696;
input x_8697;
input x_8698;
input x_8699;
input x_8700;
input x_8701;
input x_8702;
input x_8703;
input x_8704;
input x_8705;
input x_8706;
input x_8707;
input x_8708;
input x_8709;
input x_8710;
input x_8711;
input x_8712;
input x_8713;
input x_8714;
input x_8715;
input x_8716;
input x_8717;
input x_8718;
input x_8719;
input x_8720;
input x_8721;
input x_8722;
input x_8723;
input x_8724;
input x_8725;
input x_8726;
input x_8727;
input x_8728;
input x_8729;
input x_8730;
input x_8731;
input x_8732;
input x_8733;
input x_8734;
input x_8735;
input x_8736;
input x_8737;
input x_8738;
input x_8739;
input x_8740;
input x_8741;
input x_8742;
input x_8743;
input x_8744;
input x_8745;
input x_8746;
input x_8747;
input x_8748;
input x_8749;
input x_8750;
input x_8751;
input x_8752;
input x_8753;
input x_8754;
input x_8755;
input x_8756;
input x_8757;
input x_8758;
input x_8759;
input x_8760;
input x_8761;
input x_8762;
input x_8763;
input x_8764;
input x_8765;
input x_8766;
input x_8767;
input x_8768;
input x_8769;
input x_8770;
input x_8771;
input x_8772;
input x_8773;
input x_8774;
input x_8775;
input x_8776;
input x_8777;
input x_8778;
input x_8779;
input x_8780;
input x_8781;
input x_8782;
input x_8783;
input x_8784;
input x_8785;
input x_8786;
input x_8787;
input x_8788;
input x_8789;
input x_8790;
input x_8791;
input x_8792;
input x_8793;
input x_8794;
input x_8795;
input x_8796;
input x_8797;
input x_8798;
input x_8799;
input x_8800;
input x_8801;
input x_8802;
input x_8803;
input x_8804;
input x_8805;
input x_8806;
input x_8807;
input x_8808;
input x_8809;
input x_8810;
input x_8811;
input x_8812;
input x_8813;
input x_8814;
input x_8815;
input x_8816;
input x_8817;
input x_8818;
input x_8819;
input x_8820;
input x_8821;
input x_8822;
input x_8823;
input x_8824;
input x_8825;
input x_8826;
input x_8827;
input x_8828;
input x_8829;
input x_8830;
input x_8831;
input x_8832;
input x_8833;
input x_8834;
input x_8835;
input x_8836;
input x_8837;
input x_8838;
input x_8839;
input x_8840;
input x_8841;
input x_8842;
input x_8843;
input x_8844;
input x_8845;
input x_8846;
input x_8847;
input x_8848;
input x_8849;
input x_8850;
input x_8851;
input x_8852;
input x_8853;
input x_8854;
input x_8855;
input x_8856;
input x_8857;
input x_8858;
input x_8859;
input x_8860;
input x_8861;
input x_8862;
input x_8863;
input x_8864;
input x_8865;
input x_8866;
input x_8867;
input x_8868;
input x_8869;
input x_8870;
input x_8871;
input x_8872;
input x_8873;
input x_8874;
input x_8875;
input x_8876;
input x_8877;
input x_8878;
input x_8879;
input x_8880;
input x_8881;
input x_8882;
input x_8883;
input x_8884;
input x_8885;
input x_8886;
input x_8887;
input x_8888;
input x_8889;
input x_8890;
input x_8891;
input x_8892;
input x_8893;
input x_8894;
input x_8895;
input x_8896;
input x_8897;
input x_8898;
input x_8899;
input x_8900;
input x_8901;
input x_8902;
input x_8903;
input x_8904;
input x_8905;
input x_8906;
input x_8907;
input x_8908;
input x_8909;
input x_8910;
input x_8911;
input x_8912;
input x_8913;
input x_8914;
input x_8915;
input x_8916;
input x_8917;
input x_8918;
input x_8919;
input x_8920;
input x_8921;
input x_8922;
input x_8923;
input x_8924;
input x_8925;
input x_8926;
input x_8927;
input x_8928;
input x_8929;
input x_8930;
input x_8931;
input x_8932;
input x_8933;
input x_8934;
input x_8935;
input x_8936;
input x_8937;
input x_8938;
input x_8939;
input x_8940;
input x_8941;
input x_8942;
input x_8943;
input x_8944;
input x_8945;
input x_8946;
input x_8947;
input x_8948;
input x_8949;
input x_8950;
input x_8951;
input x_8952;
input x_8953;
input x_8954;
input x_8955;
input x_8956;
input x_8957;
input x_8958;
input x_8959;
input x_8960;
input x_8961;
input x_8962;
input x_8963;
input x_8964;
input x_8965;
input x_8966;
input x_8967;
input x_8968;
input x_8969;
input x_8970;
input x_8971;
input x_8972;
input x_8973;
input x_8974;
input x_8975;
input x_8976;
input x_8977;
input x_8978;
input x_8979;
input x_8980;
input x_8981;
input x_8982;
input x_8983;
input x_8984;
input x_8985;
input x_8986;
input x_8987;
input x_8988;
input x_8989;
input x_8990;
input x_8991;
input x_8992;
input x_8993;
input x_8994;
input x_8995;
input x_8996;
input x_8997;
input x_8998;
input x_8999;
input x_9000;
input x_9001;
input x_9002;
input x_9003;
input x_9004;
input x_9005;
input x_9006;
input x_9007;
input x_9008;
input x_9009;
input x_9010;
input x_9011;
input x_9012;
input x_9013;
input x_9014;
input x_9015;
input x_9016;
input x_9017;
input x_9018;
input x_9019;
input x_9020;
input x_9021;
input x_9022;
input x_9023;
input x_9024;
input x_9025;
input x_9026;
input x_9027;
input x_9028;
input x_9029;
input x_9030;
input x_9031;
input x_9032;
input x_9033;
input x_9034;
input x_9035;
input x_9036;
input x_9037;
input x_9038;
input x_9039;
input x_9040;
input x_9041;
input x_9042;
input x_9043;
input x_9044;
input x_9045;
input x_9046;
input x_9047;
input x_9048;
input x_9049;
input x_9050;
input x_9051;
input x_9052;
input x_9053;
input x_9054;
input x_9055;
input x_9056;
input x_9057;
input x_9058;
input x_9059;
input x_9060;
input x_9061;
input x_9062;
input x_9063;
input x_9064;
input x_9065;
input x_9066;
input x_9067;
input x_9068;
input x_9069;
input x_9070;
input x_9071;
input x_9072;
input x_9073;
input x_9074;
input x_9075;
input x_9076;
input x_9077;
input x_9078;
input x_9079;
input x_9080;
input x_9081;
input x_9082;
input x_9083;
input x_9084;
input x_9085;
input x_9086;
input x_9087;
input x_9088;
input x_9089;
input x_9090;
input x_9091;
input x_9092;
input x_9093;
input x_9094;
input x_9095;
input x_9096;
input x_9097;
input x_9098;
input x_9099;
input x_9100;
input x_9101;
input x_9102;
input x_9103;
input x_9104;
input x_9105;
input x_9106;
input x_9107;
input x_9108;
input x_9109;
input x_9110;
input x_9111;
input x_9112;
input x_9113;
input x_9114;
input x_9115;
input x_9116;
input x_9117;
input x_9118;
input x_9119;
input x_9120;
input x_9121;
input x_9122;
input x_9123;
input x_9124;
input x_9125;
input x_9126;
input x_9127;
input x_9128;
input x_9129;
input x_9130;
input x_9131;
input x_9132;
input x_9133;
input x_9134;
input x_9135;
input x_9136;
input x_9137;
input x_9138;
input x_9139;
input x_9140;
input x_9141;
input x_9142;
input x_9143;
input x_9144;
input x_9145;
input x_9146;
input x_9147;
input x_9148;
input x_9149;
input x_9150;
input x_9151;
input x_9152;
input x_9153;
input x_9154;
input x_9155;
input x_9156;
input x_9157;
input x_9158;
input x_9159;
input x_9160;
input x_9161;
input x_9162;
input x_9163;
input x_9164;
input x_9165;
input x_9166;
input x_9167;
input x_9168;
input x_9169;
input x_9170;
input x_9171;
input x_9172;
input x_9173;
input x_9174;
input x_9175;
input x_9176;
input x_9177;
input x_9178;
input x_9179;
input x_9180;
input x_9181;
input x_9182;
input x_9183;
input x_9184;
input x_9185;
input x_9186;
input x_9187;
input x_9188;
input x_9189;
input x_9190;
input x_9191;
input x_9192;
input x_9193;
input x_9194;
input x_9195;
input x_9196;
input x_9197;
input x_9198;
input x_9199;
input x_9200;
input x_9201;
input x_9202;
input x_9203;
input x_9204;
input x_9205;
input x_9206;
input x_9207;
input x_9208;
input x_9209;
input x_9210;
input x_9211;
input x_9212;
input x_9213;
input x_9214;
input x_9215;
input x_9216;
input x_9217;
input x_9218;
input x_9219;
input x_9220;
input x_9221;
input x_9222;
input x_9223;
input x_9224;
input x_9225;
input x_9226;
input x_9227;
input x_9228;
input x_9229;
input x_9230;
input x_9231;
input x_9232;
input x_9233;
input x_9234;
input x_9235;
input x_9236;
input x_9237;
input x_9238;
input x_9239;
input x_9240;
input x_9241;
input x_9242;
input x_9243;
input x_9244;
input x_9245;
input x_9246;
input x_9247;
input x_9248;
input x_9249;
input x_9250;
input x_9251;
input x_9252;
input x_9253;
input x_9254;
input x_9255;
input x_9256;
input x_9257;
input x_9258;
input x_9259;
input x_9260;
input x_9261;
input x_9262;
input x_9263;
input x_9264;
input x_9265;
input x_9266;
input x_9267;
input x_9268;
input x_9269;
input x_9270;
input x_9271;
input x_9272;
input x_9273;
input x_9274;
input x_9275;
input x_9276;
input x_9277;
input x_9278;
input x_9279;
input x_9280;
input x_9281;
input x_9282;
input x_9283;
input x_9284;
input x_9285;
input x_9286;
input x_9287;
input x_9288;
input x_9289;
input x_9290;
input x_9291;
input x_9292;
input x_9293;
input x_9294;
input x_9295;
input x_9296;
input x_9297;
input x_9298;
input x_9299;
input x_9300;
input x_9301;
input x_9302;
input x_9303;
input x_9304;
input x_9305;
input x_9306;
input x_9307;
input x_9308;
input x_9309;
input x_9310;
input x_9311;
input x_9312;
input x_9313;
input x_9314;
input x_9315;
input x_9316;
input x_9317;
input x_9318;
input x_9319;
input x_9320;
input x_9321;
input x_9322;
input x_9323;
input x_9324;
input x_9325;
input x_9326;
input x_9327;
input x_9328;
input x_9329;
input x_9330;
input x_9331;
input x_9332;
input x_9333;
input x_9334;
input x_9335;
input x_9336;
input x_9337;
input x_9338;
input x_9339;
input x_9340;
input x_9341;
input x_9342;
input x_9343;
input x_9344;
input x_9345;
input x_9346;
input x_9347;
input x_9348;
input x_9349;
input x_9350;
input x_9351;
input x_9352;
input x_9353;
input x_9354;
input x_9355;
input x_9356;
input x_9357;
input x_9358;
input x_9359;
input x_9360;
input x_9361;
input x_9362;
input x_9363;
input x_9364;
input x_9365;
input x_9366;
input x_9367;
input x_9368;
input x_9369;
input x_9370;
input x_9371;
input x_9372;
input x_9373;
input x_9374;
input x_9375;
input x_9376;
input x_9377;
input x_9378;
input x_9379;
input x_9380;
input x_9381;
input x_9382;
input x_9383;
input x_9384;
input x_9385;
input x_9386;
input x_9387;
input x_9388;
input x_9389;
input x_9390;
input x_9391;
input x_9392;
input x_9393;
input x_9394;
input x_9395;
input x_9396;
input x_9397;
input x_9398;
input x_9399;
input x_9400;
input x_9401;
input x_9402;
input x_9403;
input x_9404;
input x_9405;
input x_9406;
input x_9407;
input x_9408;
input x_9409;
input x_9410;
input x_9411;
input x_9412;
input x_9413;
input x_9414;
input x_9415;
input x_9416;
input x_9417;
input x_9418;
input x_9419;
input x_9420;
input x_9421;
input x_9422;
input x_9423;
input x_9424;
input x_9425;
input x_9426;
input x_9427;
input x_9428;
input x_9429;
input x_9430;
input x_9431;
input x_9432;
input x_9433;
input x_9434;
input x_9435;
input x_9436;
input x_9437;
input x_9438;
input x_9439;
input x_9440;
input x_9441;
input x_9442;
input x_9443;
input x_9444;
input x_9445;
input x_9446;
input x_9447;
input x_9448;
input x_9449;
input x_9450;
input x_9451;
input x_9452;
input x_9453;
input x_9454;
input x_9455;
input x_9456;
input x_9457;
input x_9458;
input x_9459;
input x_9460;
input x_9461;
input x_9462;
input x_9463;
input x_9464;
input x_9465;
input x_9466;
input x_9467;
input x_9468;
input x_9469;
input x_9470;
input x_9471;
input x_9472;
input x_9473;
input x_9474;
input x_9475;
input x_9476;
input x_9477;
input x_9478;
input x_9479;
input x_9480;
input x_9481;
input x_9482;
input x_9483;
input x_9484;
input x_9485;
input x_9486;
input x_9487;
input x_9488;
input x_9489;
input x_9490;
input x_9491;
input x_9492;
input x_9493;
input x_9494;
input x_9495;
input x_9496;
input x_9497;
input x_9498;
input x_9499;
input x_9500;
input x_9501;
input x_9502;
input x_9503;
input x_9504;
input x_9505;
input x_9506;
input x_9507;
input x_9508;
input x_9509;
input x_9510;
input x_9511;
input x_9512;
input x_9513;
input x_9514;
input x_9515;
input x_9516;
input x_9517;
input x_9518;
input x_9519;
input x_9520;
input x_9521;
input x_9522;
input x_9523;
input x_9524;
input x_9525;
input x_9526;
input x_9527;
input x_9528;
input x_9529;
input x_9530;
input x_9531;
input x_9532;
input x_9533;
input x_9534;
input x_9535;
input x_9536;
input x_9537;
input x_9538;
input x_9539;
input x_9540;
input x_9541;
input x_9542;
input x_9543;
input x_9544;
input x_9545;
input x_9546;
input x_9547;
input x_9548;
input x_9549;
input x_9550;
input x_9551;
input x_9552;
input x_9553;
input x_9554;
input x_9555;
input x_9556;
input x_9557;
input x_9558;
input x_9559;
input x_9560;
input x_9561;
input x_9562;
input x_9563;
input x_9564;
input x_9565;
input x_9566;
input x_9567;
input x_9568;
input x_9569;
input x_9570;
input x_9571;
input x_9572;
input x_9573;
input x_9574;
input x_9575;
input x_9576;
input x_9577;
input x_9578;
input x_9579;
input x_9580;
input x_9581;
input x_9582;
input x_9583;
input x_9584;
input x_9585;
input x_9586;
input x_9587;
input x_9588;
input x_9589;
input x_9590;
input x_9591;
input x_9592;
input x_9593;
input x_9594;
input x_9595;
input x_9596;
input x_9597;
input x_9598;
input x_9599;
input x_9600;
input x_9601;
input x_9602;
input x_9603;
input x_9604;
input x_9605;
input x_9606;
input x_9607;
input x_9608;
input x_9609;
input x_9610;
input x_9611;
input x_9612;
input x_9613;
input x_9614;
input x_9615;
input x_9616;
input x_9617;
input x_9618;
input x_9619;
input x_9620;
input x_9621;
input x_9622;
input x_9623;
input x_9624;
input x_9625;
input x_9626;
input x_9627;
input x_9628;
input x_9629;
input x_9630;
input x_9631;
input x_9632;
input x_9633;
input x_9634;
input x_9635;
input x_9636;
input x_9637;
input x_9638;
input x_9639;
input x_9640;
input x_9641;
input x_9642;
input x_9643;
input x_9644;
input x_9645;
input x_9646;
input x_9647;
input x_9648;
input x_9649;
input x_9650;
input x_9651;
input x_9652;
input x_9653;
input x_9654;
input x_9655;
input x_9656;
input x_9657;
input x_9658;
input x_9659;
input x_9660;
input x_9661;
input x_9662;
input x_9663;
input x_9664;
input x_9665;
input x_9666;
input x_9667;
input x_9668;
input x_9669;
input x_9670;
input x_9671;
input x_9672;
input x_9673;
input x_9674;
input x_9675;
input x_9676;
input x_9677;
input x_9678;
input x_9679;
input x_9680;
input x_9681;
input x_9682;
input x_9683;
input x_9684;
input x_9685;
input x_9686;
input x_9687;
input x_9688;
input x_9689;
input x_9690;
input x_9691;
input x_9692;
input x_9693;
input x_9694;
input x_9695;
input x_9696;
input x_9697;
input x_9698;
input x_9699;
input x_9700;
input x_9701;
input x_9702;
input x_9703;
input x_9704;
input x_9705;
input x_9706;
input x_9707;
input x_9708;
input x_9709;
input x_9710;
input x_9711;
input x_9712;
input x_9713;
input x_9714;
input x_9715;
input x_9716;
input x_9717;
input x_9718;
input x_9719;
input x_9720;
input x_9721;
input x_9722;
input x_9723;
input x_9724;
input x_9725;
input x_9726;
input x_9727;
input x_9728;
input x_9729;
input x_9730;
input x_9731;
input x_9732;
input x_9733;
input x_9734;
input x_9735;
input x_9736;
input x_9737;
input x_9738;
input x_9739;
input x_9740;
input x_9741;
input x_9742;
input x_9743;
input x_9744;
input x_9745;
input x_9746;
input x_9747;
input x_9748;
input x_9749;
input x_9750;
input x_9751;
input x_9752;
input x_9753;
input x_9754;
input x_9755;
input x_9756;
input x_9757;
input x_9758;
input x_9759;
input x_9760;
input x_9761;
input x_9762;
input x_9763;
input x_9764;
input x_9765;
input x_9766;
input x_9767;
input x_9768;
input x_9769;
input x_9770;
input x_9771;
input x_9772;
input x_9773;
input x_9774;
input x_9775;
input x_9776;
input x_9777;
input x_9778;
input x_9779;
input x_9780;
input x_9781;
input x_9782;
input x_9783;
input x_9784;
input x_9785;
input x_9786;
input x_9787;
input x_9788;
input x_9789;
input x_9790;
input x_9791;
input x_9792;
input x_9793;
input x_9794;
input x_9795;
input x_9796;
input x_9797;
input x_9798;
input x_9799;
input x_9800;
input x_9801;
input x_9802;
input x_9803;
input x_9804;
input x_9805;
input x_9806;
input x_9807;
input x_9808;
input x_9809;
input x_9810;
input x_9811;
input x_9812;
input x_9813;
input x_9814;
input x_9815;
input x_9816;
input x_9817;
input x_9818;
input x_9819;
input x_9820;
input x_9821;
input x_9822;
input x_9823;
input x_9824;
input x_9825;
input x_9826;
input x_9827;
input x_9828;
input x_9829;
input x_9830;
input x_9831;
input x_9832;
input x_9833;
input x_9834;
input x_9835;
input x_9836;
input x_9837;
input x_9838;
input x_9839;
input x_9840;
input x_9841;
input x_9842;
input x_9843;
input x_9844;
input x_9845;
input x_9846;
input x_9847;
input x_9848;
input x_9849;
input x_9850;
input x_9851;
input x_9852;
input x_9853;
input x_9854;
input x_9855;
input x_9856;
input x_9857;
input x_9858;
input x_9859;
input x_9860;
input x_9861;
input x_9862;
input x_9863;
input x_9864;
input x_9865;
input x_9866;
input x_9867;
input x_9868;
input x_9869;
input x_9870;
input x_9871;
input x_9872;
input x_9873;
input x_9874;
input x_9875;
input x_9876;
input x_9877;
input x_9878;
input x_9879;
input x_9880;
input x_9881;
input x_9882;
input x_9883;
input x_9884;
input x_9885;
input x_9886;
input x_9887;
input x_9888;
input x_9889;
input x_9890;
input x_9891;
input x_9892;
input x_9893;
input x_9894;
input x_9895;
input x_9896;
input x_9897;
input x_9898;
input x_9899;
input x_9900;
input x_9901;
input x_9902;
input x_9903;
input x_9904;
input x_9905;
input x_9906;
input x_9907;
input x_9908;
input x_9909;
input x_9910;
input x_9911;
input x_9912;
input x_9913;
input x_9914;
input x_9915;
input x_9916;
input x_9917;
input x_9918;
input x_9919;
input x_9920;
input x_9921;
input x_9922;
input x_9923;
input x_9924;
input x_9925;
input x_9926;
input x_9927;
input x_9928;
input x_9929;
input x_9930;
input x_9931;
input x_9932;
input x_9933;
input x_9934;
input x_9935;
input x_9936;
input x_9937;
input x_9938;
input x_9939;
input x_9940;
input x_9941;
input x_9942;
input x_9943;
input x_9944;
input x_9945;
input x_9946;
input x_9947;
input x_9948;
input x_9949;
input x_9950;
input x_9951;
input x_9952;
input x_9953;
input x_9954;
input x_9955;
input x_9956;
input x_9957;
input x_9958;
input x_9959;
input x_9960;
input x_9961;
input x_9962;
input x_9963;
input x_9964;
input x_9965;
input x_9966;
input x_9967;
input x_9968;
input x_9969;
input x_9970;
input x_9971;
input x_9972;
input x_9973;
input x_9974;
input x_9975;
input x_9976;
input x_9977;
input x_9978;
input x_9979;
input x_9980;
input x_9981;
input x_9982;
input x_9983;
input x_9984;
input x_9985;
input x_9986;
input x_9987;
input x_9988;
input x_9989;
input x_9990;
input x_9991;
input x_9992;
input x_9993;
input x_9994;
input x_9995;
input x_9996;
input x_9997;
input x_9998;
input x_9999;
input x_10000;
input x_10001;
input x_10002;
input x_10003;
input x_10004;
input x_10005;
input x_10006;
input x_10007;
input x_10008;
input x_10009;
input x_10010;
input x_10011;
input x_10012;
input x_10013;
input x_10014;
input x_10015;
input x_10016;
input x_10017;
input x_10018;
input x_10019;
input x_10020;
input x_10021;
input x_10022;
input x_10023;
input x_10024;
input x_10025;
input x_10026;
input x_10027;
input x_10028;
input x_10029;
input x_10030;
input x_10031;
input x_10032;
input x_10033;
input x_10034;
input x_10035;
input x_10036;
input x_10037;
input x_10038;
input x_10039;
input x_10040;
input x_10041;
input x_10042;
input x_10043;
input x_10044;
input x_10045;
input x_10046;
input x_10047;
input x_10048;
input x_10049;
input x_10050;
input x_10051;
input x_10052;
input x_10053;
input x_10054;
input x_10055;
input x_10056;
input x_10057;
input x_10058;
input x_10059;
input x_10060;
input x_10061;
input x_10062;
input x_10063;
input x_10064;
input x_10065;
input x_10066;
input x_10067;
input x_10068;
input x_10069;
input x_10070;
input x_10071;
input x_10072;
input x_10073;
input x_10074;
input x_10075;
input x_10076;
input x_10077;
input x_10078;
input x_10079;
input x_10080;
input x_10081;
input x_10082;
input x_10083;
input x_10084;
input x_10085;
input x_10086;
input x_10087;
input x_10088;
input x_10089;
input x_10090;
input x_10091;
input x_10092;
input x_10093;
input x_10094;
output o_1;
wire n_1;
wire n_2;
wire n_3;
wire n_4;
wire n_5;
wire n_6;
wire n_7;
wire n_8;
wire n_9;
wire n_10;
wire n_11;
wire n_12;
wire n_13;
wire n_14;
wire n_15;
wire n_16;
wire n_17;
wire n_18;
wire n_19;
wire n_20;
wire n_21;
wire n_22;
wire n_23;
wire n_24;
wire n_25;
wire n_26;
wire n_27;
wire n_28;
wire n_29;
wire n_30;
wire n_31;
wire n_32;
wire n_33;
wire n_34;
wire n_35;
wire n_36;
wire n_37;
wire n_38;
wire n_39;
wire n_40;
wire n_41;
wire n_42;
wire n_43;
wire n_44;
wire n_45;
wire n_46;
wire n_47;
wire n_48;
wire n_49;
wire n_50;
wire n_51;
wire n_52;
wire n_53;
wire n_54;
wire n_55;
wire n_56;
wire n_57;
wire n_58;
wire n_59;
wire n_60;
wire n_61;
wire n_62;
wire n_63;
wire n_64;
wire n_65;
wire n_66;
wire n_67;
wire n_68;
wire n_69;
wire n_70;
wire n_71;
wire n_72;
wire n_73;
wire n_74;
wire n_75;
wire n_76;
wire n_77;
wire n_78;
wire n_79;
wire n_80;
wire n_81;
wire n_82;
wire n_83;
wire n_84;
wire n_85;
wire n_86;
wire n_87;
wire n_88;
wire n_89;
wire n_90;
wire n_91;
wire n_92;
wire n_93;
wire n_94;
wire n_95;
wire n_96;
wire n_97;
wire n_98;
wire n_99;
wire n_100;
wire n_101;
wire n_102;
wire n_103;
wire n_104;
wire n_105;
wire n_106;
wire n_107;
wire n_108;
wire n_109;
wire n_110;
wire n_111;
wire n_112;
wire n_113;
wire n_114;
wire n_115;
wire n_116;
wire n_117;
wire n_118;
wire n_119;
wire n_120;
wire n_121;
wire n_122;
wire n_123;
wire n_124;
wire n_125;
wire n_126;
wire n_127;
wire n_128;
wire n_129;
wire n_130;
wire n_131;
wire n_132;
wire n_133;
wire n_134;
wire n_135;
wire n_136;
wire n_137;
wire n_138;
wire n_139;
wire n_140;
wire n_141;
wire n_142;
wire n_143;
wire n_144;
wire n_145;
wire n_146;
wire n_147;
wire n_148;
wire n_149;
wire n_150;
wire n_151;
wire n_152;
wire n_153;
wire n_154;
wire n_155;
wire n_156;
wire n_157;
wire n_158;
wire n_159;
wire n_160;
wire n_161;
wire n_162;
wire n_163;
wire n_164;
wire n_165;
wire n_166;
wire n_167;
wire n_168;
wire n_169;
wire n_170;
wire n_171;
wire n_172;
wire n_173;
wire n_174;
wire n_175;
wire n_176;
wire n_177;
wire n_178;
wire n_179;
wire n_180;
wire n_181;
wire n_182;
wire n_183;
wire n_184;
wire n_185;
wire n_186;
wire n_187;
wire n_188;
wire n_189;
wire n_190;
wire n_191;
wire n_192;
wire n_193;
wire n_194;
wire n_195;
wire n_196;
wire n_197;
wire n_198;
wire n_199;
wire n_200;
wire n_201;
wire n_202;
wire n_203;
wire n_204;
wire n_205;
wire n_206;
wire n_207;
wire n_208;
wire n_209;
wire n_210;
wire n_211;
wire n_212;
wire n_213;
wire n_214;
wire n_215;
wire n_216;
wire n_217;
wire n_218;
wire n_219;
wire n_220;
wire n_221;
wire n_222;
wire n_223;
wire n_224;
wire n_225;
wire n_226;
wire n_227;
wire n_228;
wire n_229;
wire n_230;
wire n_231;
wire n_232;
wire n_233;
wire n_234;
wire n_235;
wire n_236;
wire n_237;
wire n_238;
wire n_239;
wire n_240;
wire n_241;
wire n_242;
wire n_243;
wire n_244;
wire n_245;
wire n_246;
wire n_247;
wire n_248;
wire n_249;
wire n_250;
wire n_251;
wire n_252;
wire n_253;
wire n_254;
wire n_255;
wire n_256;
wire n_257;
wire n_258;
wire n_259;
wire n_260;
wire n_261;
wire n_262;
wire n_263;
wire n_264;
wire n_265;
wire n_266;
wire n_267;
wire n_268;
wire n_269;
wire n_270;
wire n_271;
wire n_272;
wire n_273;
wire n_274;
wire n_275;
wire n_276;
wire n_277;
wire n_278;
wire n_279;
wire n_280;
wire n_281;
wire n_282;
wire n_283;
wire n_284;
wire n_285;
wire n_286;
wire n_287;
wire n_288;
wire n_289;
wire n_290;
wire n_291;
wire n_292;
wire n_293;
wire n_294;
wire n_295;
wire n_296;
wire n_297;
wire n_298;
wire n_299;
wire n_300;
wire n_301;
wire n_302;
wire n_303;
wire n_304;
wire n_305;
wire n_306;
wire n_307;
wire n_308;
wire n_309;
wire n_310;
wire n_311;
wire n_312;
wire n_313;
wire n_314;
wire n_315;
wire n_316;
wire n_317;
wire n_318;
wire n_319;
wire n_320;
wire n_321;
wire n_322;
wire n_323;
wire n_324;
wire n_325;
wire n_326;
wire n_327;
wire n_328;
wire n_329;
wire n_330;
wire n_331;
wire n_332;
wire n_333;
wire n_334;
wire n_335;
wire n_336;
wire n_337;
wire n_338;
wire n_339;
wire n_340;
wire n_341;
wire n_342;
wire n_343;
wire n_344;
wire n_345;
wire n_346;
wire n_347;
wire n_348;
wire n_349;
wire n_350;
wire n_351;
wire n_352;
wire n_353;
wire n_354;
wire n_355;
wire n_356;
wire n_357;
wire n_358;
wire n_359;
wire n_360;
wire n_361;
wire n_362;
wire n_363;
wire n_364;
wire n_365;
wire n_366;
wire n_367;
wire n_368;
wire n_369;
wire n_370;
wire n_371;
wire n_372;
wire n_373;
wire n_374;
wire n_375;
wire n_376;
wire n_377;
wire n_378;
wire n_379;
wire n_380;
wire n_381;
wire n_382;
wire n_383;
wire n_384;
wire n_385;
wire n_386;
wire n_387;
wire n_388;
wire n_389;
wire n_390;
wire n_391;
wire n_392;
wire n_393;
wire n_394;
wire n_395;
wire n_396;
wire n_397;
wire n_398;
wire n_399;
wire n_400;
wire n_401;
wire n_402;
wire n_403;
wire n_404;
wire n_405;
wire n_406;
wire n_407;
wire n_408;
wire n_409;
wire n_410;
wire n_411;
wire n_412;
wire n_413;
wire n_414;
wire n_415;
wire n_416;
wire n_417;
wire n_418;
wire n_419;
wire n_420;
wire n_421;
wire n_422;
wire n_423;
wire n_424;
wire n_425;
wire n_426;
wire n_427;
wire n_428;
wire n_429;
wire n_430;
wire n_431;
wire n_432;
wire n_433;
wire n_434;
wire n_435;
wire n_436;
wire n_437;
wire n_438;
wire n_439;
wire n_440;
wire n_441;
wire n_442;
wire n_443;
wire n_444;
wire n_445;
wire n_446;
wire n_447;
wire n_448;
wire n_449;
wire n_450;
wire n_451;
wire n_452;
wire n_453;
wire n_454;
wire n_455;
wire n_456;
wire n_457;
wire n_458;
wire n_459;
wire n_460;
wire n_461;
wire n_462;
wire n_463;
wire n_464;
wire n_465;
wire n_466;
wire n_467;
wire n_468;
wire n_469;
wire n_470;
wire n_471;
wire n_472;
wire n_473;
wire n_474;
wire n_475;
wire n_476;
wire n_477;
wire n_478;
wire n_479;
wire n_480;
wire n_481;
wire n_482;
wire n_483;
wire n_484;
wire n_485;
wire n_486;
wire n_487;
wire n_488;
wire n_489;
wire n_490;
wire n_491;
wire n_492;
wire n_493;
wire n_494;
wire n_495;
wire n_496;
wire n_497;
wire n_498;
wire n_499;
wire n_500;
wire n_501;
wire n_502;
wire n_503;
wire n_504;
wire n_505;
wire n_506;
wire n_507;
wire n_508;
wire n_509;
wire n_510;
wire n_511;
wire n_512;
wire n_513;
wire n_514;
wire n_515;
wire n_516;
wire n_517;
wire n_518;
wire n_519;
wire n_520;
wire n_521;
wire n_522;
wire n_523;
wire n_524;
wire n_525;
wire n_526;
wire n_527;
wire n_528;
wire n_529;
wire n_530;
wire n_531;
wire n_532;
wire n_533;
wire n_534;
wire n_535;
wire n_536;
wire n_537;
wire n_538;
wire n_539;
wire n_540;
wire n_541;
wire n_542;
wire n_543;
wire n_544;
wire n_545;
wire n_546;
wire n_547;
wire n_548;
wire n_549;
wire n_550;
wire n_551;
wire n_552;
wire n_553;
wire n_554;
wire n_555;
wire n_556;
wire n_557;
wire n_558;
wire n_559;
wire n_560;
wire n_561;
wire n_562;
wire n_563;
wire n_564;
wire n_565;
wire n_566;
wire n_567;
wire n_568;
wire n_569;
wire n_570;
wire n_571;
wire n_572;
wire n_573;
wire n_574;
wire n_575;
wire n_576;
wire n_577;
wire n_578;
wire n_579;
wire n_580;
wire n_581;
wire n_582;
wire n_583;
wire n_584;
wire n_585;
wire n_586;
wire n_587;
wire n_588;
wire n_589;
wire n_590;
wire n_591;
wire n_592;
wire n_593;
wire n_594;
wire n_595;
wire n_596;
wire n_597;
wire n_598;
wire n_599;
wire n_600;
wire n_601;
wire n_602;
wire n_603;
wire n_604;
wire n_605;
wire n_606;
wire n_607;
wire n_608;
wire n_609;
wire n_610;
wire n_611;
wire n_612;
wire n_613;
wire n_614;
wire n_615;
wire n_616;
wire n_617;
wire n_618;
wire n_619;
wire n_620;
wire n_621;
wire n_622;
wire n_623;
wire n_624;
wire n_625;
wire n_626;
wire n_627;
wire n_628;
wire n_629;
wire n_630;
wire n_631;
wire n_632;
wire n_633;
wire n_634;
wire n_635;
wire n_636;
wire n_637;
wire n_638;
wire n_639;
wire n_640;
wire n_641;
wire n_642;
wire n_643;
wire n_644;
wire n_645;
wire n_646;
wire n_647;
wire n_648;
wire n_649;
wire n_650;
wire n_651;
wire n_652;
wire n_653;
wire n_654;
wire n_655;
wire n_656;
wire n_657;
wire n_658;
wire n_659;
wire n_660;
wire n_661;
wire n_662;
wire n_663;
wire n_664;
wire n_665;
wire n_666;
wire n_667;
wire n_668;
wire n_669;
wire n_670;
wire n_671;
wire n_672;
wire n_673;
wire n_674;
wire n_675;
wire n_676;
wire n_677;
wire n_678;
wire n_679;
wire n_680;
wire n_681;
wire n_682;
wire n_683;
wire n_684;
wire n_685;
wire n_686;
wire n_687;
wire n_688;
wire n_689;
wire n_690;
wire n_691;
wire n_692;
wire n_693;
wire n_694;
wire n_695;
wire n_696;
wire n_697;
wire n_698;
wire n_699;
wire n_700;
wire n_701;
wire n_702;
wire n_703;
wire n_704;
wire n_705;
wire n_706;
wire n_707;
wire n_708;
wire n_709;
wire n_710;
wire n_711;
wire n_712;
wire n_713;
wire n_714;
wire n_715;
wire n_716;
wire n_717;
wire n_718;
wire n_719;
wire n_720;
wire n_721;
wire n_722;
wire n_723;
wire n_724;
wire n_725;
wire n_726;
wire n_727;
wire n_728;
wire n_729;
wire n_730;
wire n_731;
wire n_732;
wire n_733;
wire n_734;
wire n_735;
wire n_736;
wire n_737;
wire n_738;
wire n_739;
wire n_740;
wire n_741;
wire n_742;
wire n_743;
wire n_744;
wire n_745;
wire n_746;
wire n_747;
wire n_748;
wire n_749;
wire n_750;
wire n_751;
wire n_752;
wire n_753;
wire n_754;
wire n_755;
wire n_756;
wire n_757;
wire n_758;
wire n_759;
wire n_760;
wire n_761;
wire n_762;
wire n_763;
wire n_764;
wire n_765;
wire n_766;
wire n_767;
wire n_768;
wire n_769;
wire n_770;
wire n_771;
wire n_772;
wire n_773;
wire n_774;
wire n_775;
wire n_776;
wire n_777;
wire n_778;
wire n_779;
wire n_780;
wire n_781;
wire n_782;
wire n_783;
wire n_784;
wire n_785;
wire n_786;
wire n_787;
wire n_788;
wire n_789;
wire n_790;
wire n_791;
wire n_792;
wire n_793;
wire n_794;
wire n_795;
wire n_796;
wire n_797;
wire n_798;
wire n_799;
wire n_800;
wire n_801;
wire n_802;
wire n_803;
wire n_804;
wire n_805;
wire n_806;
wire n_807;
wire n_808;
wire n_809;
wire n_810;
wire n_811;
wire n_812;
wire n_813;
wire n_814;
wire n_815;
wire n_816;
wire n_817;
wire n_818;
wire n_819;
wire n_820;
wire n_821;
wire n_822;
wire n_823;
wire n_824;
wire n_825;
wire n_826;
wire n_827;
wire n_828;
wire n_829;
wire n_830;
wire n_831;
wire n_832;
wire n_833;
wire n_834;
wire n_835;
wire n_836;
wire n_837;
wire n_838;
wire n_839;
wire n_840;
wire n_841;
wire n_842;
wire n_843;
wire n_844;
wire n_845;
wire n_846;
wire n_847;
wire n_848;
wire n_849;
wire n_850;
wire n_851;
wire n_852;
wire n_853;
wire n_854;
wire n_855;
wire n_856;
wire n_857;
wire n_858;
wire n_859;
wire n_860;
wire n_861;
wire n_862;
wire n_863;
wire n_864;
wire n_865;
wire n_866;
wire n_867;
wire n_868;
wire n_869;
wire n_870;
wire n_871;
wire n_872;
wire n_873;
wire n_874;
wire n_875;
wire n_876;
wire n_877;
wire n_878;
wire n_879;
wire n_880;
wire n_881;
wire n_882;
wire n_883;
wire n_884;
wire n_885;
wire n_886;
wire n_887;
wire n_888;
wire n_889;
wire n_890;
wire n_891;
wire n_892;
wire n_893;
wire n_894;
wire n_895;
wire n_896;
wire n_897;
wire n_898;
wire n_899;
wire n_900;
wire n_901;
wire n_902;
wire n_903;
wire n_904;
wire n_905;
wire n_906;
wire n_907;
wire n_908;
wire n_909;
wire n_910;
wire n_911;
wire n_912;
wire n_913;
wire n_914;
wire n_915;
wire n_916;
wire n_917;
wire n_918;
wire n_919;
wire n_920;
wire n_921;
wire n_922;
wire n_923;
wire n_924;
wire n_925;
wire n_926;
wire n_927;
wire n_928;
wire n_929;
wire n_930;
wire n_931;
wire n_932;
wire n_933;
wire n_934;
wire n_935;
wire n_936;
wire n_937;
wire n_938;
wire n_939;
wire n_940;
wire n_941;
wire n_942;
wire n_943;
wire n_944;
wire n_945;
wire n_946;
wire n_947;
wire n_948;
wire n_949;
wire n_950;
wire n_951;
wire n_952;
wire n_953;
wire n_954;
wire n_955;
wire n_956;
wire n_957;
wire n_958;
wire n_959;
wire n_960;
wire n_961;
wire n_962;
wire n_963;
wire n_964;
wire n_965;
wire n_966;
wire n_967;
wire n_968;
wire n_969;
wire n_970;
wire n_971;
wire n_972;
wire n_973;
wire n_974;
wire n_975;
wire n_976;
wire n_977;
wire n_978;
wire n_979;
wire n_980;
wire n_981;
wire n_982;
wire n_983;
wire n_984;
wire n_985;
wire n_986;
wire n_987;
wire n_988;
wire n_989;
wire n_990;
wire n_991;
wire n_992;
wire n_993;
wire n_994;
wire n_995;
wire n_996;
wire n_997;
wire n_998;
wire n_999;
wire n_1000;
wire n_1001;
wire n_1002;
wire n_1003;
wire n_1004;
wire n_1005;
wire n_1006;
wire n_1007;
wire n_1008;
wire n_1009;
wire n_1010;
wire n_1011;
wire n_1012;
wire n_1013;
wire n_1014;
wire n_1015;
wire n_1016;
wire n_1017;
wire n_1018;
wire n_1019;
wire n_1020;
wire n_1021;
wire n_1022;
wire n_1023;
wire n_1024;
wire n_1025;
wire n_1026;
wire n_1027;
wire n_1028;
wire n_1029;
wire n_1030;
wire n_1031;
wire n_1032;
wire n_1033;
wire n_1034;
wire n_1035;
wire n_1036;
wire n_1037;
wire n_1038;
wire n_1039;
wire n_1040;
wire n_1041;
wire n_1042;
wire n_1043;
wire n_1044;
wire n_1045;
wire n_1046;
wire n_1047;
wire n_1048;
wire n_1049;
wire n_1050;
wire n_1051;
wire n_1052;
wire n_1053;
wire n_1054;
wire n_1055;
wire n_1056;
wire n_1057;
wire n_1058;
wire n_1059;
wire n_1060;
wire n_1061;
wire n_1062;
wire n_1063;
wire n_1064;
wire n_1065;
wire n_1066;
wire n_1067;
wire n_1068;
wire n_1069;
wire n_1070;
wire n_1071;
wire n_1072;
wire n_1073;
wire n_1074;
wire n_1075;
wire n_1076;
wire n_1077;
wire n_1078;
wire n_1079;
wire n_1080;
wire n_1081;
wire n_1082;
wire n_1083;
wire n_1084;
wire n_1085;
wire n_1086;
wire n_1087;
wire n_1088;
wire n_1089;
wire n_1090;
wire n_1091;
wire n_1092;
wire n_1093;
wire n_1094;
wire n_1095;
wire n_1096;
wire n_1097;
wire n_1098;
wire n_1099;
wire n_1100;
wire n_1101;
wire n_1102;
wire n_1103;
wire n_1104;
wire n_1105;
wire n_1106;
wire n_1107;
wire n_1108;
wire n_1109;
wire n_1110;
wire n_1111;
wire n_1112;
wire n_1113;
wire n_1114;
wire n_1115;
wire n_1116;
wire n_1117;
wire n_1118;
wire n_1119;
wire n_1120;
wire n_1121;
wire n_1122;
wire n_1123;
wire n_1124;
wire n_1125;
wire n_1126;
wire n_1127;
wire n_1128;
wire n_1129;
wire n_1130;
wire n_1131;
wire n_1132;
wire n_1133;
wire n_1134;
wire n_1135;
wire n_1136;
wire n_1137;
wire n_1138;
wire n_1139;
wire n_1140;
wire n_1141;
wire n_1142;
wire n_1143;
wire n_1144;
wire n_1145;
wire n_1146;
wire n_1147;
wire n_1148;
wire n_1149;
wire n_1150;
wire n_1151;
wire n_1152;
wire n_1153;
wire n_1154;
wire n_1155;
wire n_1156;
wire n_1157;
wire n_1158;
wire n_1159;
wire n_1160;
wire n_1161;
wire n_1162;
wire n_1163;
wire n_1164;
wire n_1165;
wire n_1166;
wire n_1167;
wire n_1168;
wire n_1169;
wire n_1170;
wire n_1171;
wire n_1172;
wire n_1173;
wire n_1174;
wire n_1175;
wire n_1176;
wire n_1177;
wire n_1178;
wire n_1179;
wire n_1180;
wire n_1181;
wire n_1182;
wire n_1183;
wire n_1184;
wire n_1185;
wire n_1186;
wire n_1187;
wire n_1188;
wire n_1189;
wire n_1190;
wire n_1191;
wire n_1192;
wire n_1193;
wire n_1194;
wire n_1195;
wire n_1196;
wire n_1197;
wire n_1198;
wire n_1199;
wire n_1200;
wire n_1201;
wire n_1202;
wire n_1203;
wire n_1204;
wire n_1205;
wire n_1206;
wire n_1207;
wire n_1208;
wire n_1209;
wire n_1210;
wire n_1211;
wire n_1212;
wire n_1213;
wire n_1214;
wire n_1215;
wire n_1216;
wire n_1217;
wire n_1218;
wire n_1219;
wire n_1220;
wire n_1221;
wire n_1222;
wire n_1223;
wire n_1224;
wire n_1225;
wire n_1226;
wire n_1227;
wire n_1228;
wire n_1229;
wire n_1230;
wire n_1231;
wire n_1232;
wire n_1233;
wire n_1234;
wire n_1235;
wire n_1236;
wire n_1237;
wire n_1238;
wire n_1239;
wire n_1240;
wire n_1241;
wire n_1242;
wire n_1243;
wire n_1244;
wire n_1245;
wire n_1246;
wire n_1247;
wire n_1248;
wire n_1249;
wire n_1250;
wire n_1251;
wire n_1252;
wire n_1253;
wire n_1254;
wire n_1255;
wire n_1256;
wire n_1257;
wire n_1258;
wire n_1259;
wire n_1260;
wire n_1261;
wire n_1262;
wire n_1263;
wire n_1264;
wire n_1265;
wire n_1266;
wire n_1267;
wire n_1268;
wire n_1269;
wire n_1270;
wire n_1271;
wire n_1272;
wire n_1273;
wire n_1274;
wire n_1275;
wire n_1276;
wire n_1277;
wire n_1278;
wire n_1279;
wire n_1280;
wire n_1281;
wire n_1282;
wire n_1283;
wire n_1284;
wire n_1285;
wire n_1286;
wire n_1287;
wire n_1288;
wire n_1289;
wire n_1290;
wire n_1291;
wire n_1292;
wire n_1293;
wire n_1294;
wire n_1295;
wire n_1296;
wire n_1297;
wire n_1298;
wire n_1299;
wire n_1300;
wire n_1301;
wire n_1302;
wire n_1303;
wire n_1304;
wire n_1305;
wire n_1306;
wire n_1307;
wire n_1308;
wire n_1309;
wire n_1310;
wire n_1311;
wire n_1312;
wire n_1313;
wire n_1314;
wire n_1315;
wire n_1316;
wire n_1317;
wire n_1318;
wire n_1319;
wire n_1320;
wire n_1321;
wire n_1322;
wire n_1323;
wire n_1324;
wire n_1325;
wire n_1326;
wire n_1327;
wire n_1328;
wire n_1329;
wire n_1330;
wire n_1331;
wire n_1332;
wire n_1333;
wire n_1334;
wire n_1335;
wire n_1336;
wire n_1337;
wire n_1338;
wire n_1339;
wire n_1340;
wire n_1341;
wire n_1342;
wire n_1343;
wire n_1344;
wire n_1345;
wire n_1346;
wire n_1347;
wire n_1348;
wire n_1349;
wire n_1350;
wire n_1351;
wire n_1352;
wire n_1353;
wire n_1354;
wire n_1355;
wire n_1356;
wire n_1357;
wire n_1358;
wire n_1359;
wire n_1360;
wire n_1361;
wire n_1362;
wire n_1363;
wire n_1364;
wire n_1365;
wire n_1366;
wire n_1367;
wire n_1368;
wire n_1369;
wire n_1370;
wire n_1371;
wire n_1372;
wire n_1373;
wire n_1374;
wire n_1375;
wire n_1376;
wire n_1377;
wire n_1378;
wire n_1379;
wire n_1380;
wire n_1381;
wire n_1382;
wire n_1383;
wire n_1384;
wire n_1385;
wire n_1386;
wire n_1387;
wire n_1388;
wire n_1389;
wire n_1390;
wire n_1391;
wire n_1392;
wire n_1393;
wire n_1394;
wire n_1395;
wire n_1396;
wire n_1397;
wire n_1398;
wire n_1399;
wire n_1400;
wire n_1401;
wire n_1402;
wire n_1403;
wire n_1404;
wire n_1405;
wire n_1406;
wire n_1407;
wire n_1408;
wire n_1409;
wire n_1410;
wire n_1411;
wire n_1412;
wire n_1413;
wire n_1414;
wire n_1415;
wire n_1416;
wire n_1417;
wire n_1418;
wire n_1419;
wire n_1420;
wire n_1421;
wire n_1422;
wire n_1423;
wire n_1424;
wire n_1425;
wire n_1426;
wire n_1427;
wire n_1428;
wire n_1429;
wire n_1430;
wire n_1431;
wire n_1432;
wire n_1433;
wire n_1434;
wire n_1435;
wire n_1436;
wire n_1437;
wire n_1438;
wire n_1439;
wire n_1440;
wire n_1441;
wire n_1442;
wire n_1443;
wire n_1444;
wire n_1445;
wire n_1446;
wire n_1447;
wire n_1448;
wire n_1449;
wire n_1450;
wire n_1451;
wire n_1452;
wire n_1453;
wire n_1454;
wire n_1455;
wire n_1456;
wire n_1457;
wire n_1458;
wire n_1459;
wire n_1460;
wire n_1461;
wire n_1462;
wire n_1463;
wire n_1464;
wire n_1465;
wire n_1466;
wire n_1467;
wire n_1468;
wire n_1469;
wire n_1470;
wire n_1471;
wire n_1472;
wire n_1473;
wire n_1474;
wire n_1475;
wire n_1476;
wire n_1477;
wire n_1478;
wire n_1479;
wire n_1480;
wire n_1481;
wire n_1482;
wire n_1483;
wire n_1484;
wire n_1485;
wire n_1486;
wire n_1487;
wire n_1488;
wire n_1489;
wire n_1490;
wire n_1491;
wire n_1492;
wire n_1493;
wire n_1494;
wire n_1495;
wire n_1496;
wire n_1497;
wire n_1498;
wire n_1499;
wire n_1500;
wire n_1501;
wire n_1502;
wire n_1503;
wire n_1504;
wire n_1505;
wire n_1506;
wire n_1507;
wire n_1508;
wire n_1509;
wire n_1510;
wire n_1511;
wire n_1512;
wire n_1513;
wire n_1514;
wire n_1515;
wire n_1516;
wire n_1517;
wire n_1518;
wire n_1519;
wire n_1520;
wire n_1521;
wire n_1522;
wire n_1523;
wire n_1524;
wire n_1525;
wire n_1526;
wire n_1527;
wire n_1528;
wire n_1529;
wire n_1530;
wire n_1531;
wire n_1532;
wire n_1533;
wire n_1534;
wire n_1535;
wire n_1536;
wire n_1537;
wire n_1538;
wire n_1539;
wire n_1540;
wire n_1541;
wire n_1542;
wire n_1543;
wire n_1544;
wire n_1545;
wire n_1546;
wire n_1547;
wire n_1548;
wire n_1549;
wire n_1550;
wire n_1551;
wire n_1552;
wire n_1553;
wire n_1554;
wire n_1555;
wire n_1556;
wire n_1557;
wire n_1558;
wire n_1559;
wire n_1560;
wire n_1561;
wire n_1562;
wire n_1563;
wire n_1564;
wire n_1565;
wire n_1566;
wire n_1567;
wire n_1568;
wire n_1569;
wire n_1570;
wire n_1571;
wire n_1572;
wire n_1573;
wire n_1574;
wire n_1575;
wire n_1576;
wire n_1577;
wire n_1578;
wire n_1579;
wire n_1580;
wire n_1581;
wire n_1582;
wire n_1583;
wire n_1584;
wire n_1585;
wire n_1586;
wire n_1587;
wire n_1588;
wire n_1589;
wire n_1590;
wire n_1591;
wire n_1592;
wire n_1593;
wire n_1594;
wire n_1595;
wire n_1596;
wire n_1597;
wire n_1598;
wire n_1599;
wire n_1600;
wire n_1601;
wire n_1602;
wire n_1603;
wire n_1604;
wire n_1605;
wire n_1606;
wire n_1607;
wire n_1608;
wire n_1609;
wire n_1610;
wire n_1611;
wire n_1612;
wire n_1613;
wire n_1614;
wire n_1615;
wire n_1616;
wire n_1617;
wire n_1618;
wire n_1619;
wire n_1620;
wire n_1621;
wire n_1622;
wire n_1623;
wire n_1624;
wire n_1625;
wire n_1626;
wire n_1627;
wire n_1628;
wire n_1629;
wire n_1630;
wire n_1631;
wire n_1632;
wire n_1633;
wire n_1634;
wire n_1635;
wire n_1636;
wire n_1637;
wire n_1638;
wire n_1639;
wire n_1640;
wire n_1641;
wire n_1642;
wire n_1643;
wire n_1644;
wire n_1645;
wire n_1646;
wire n_1647;
wire n_1648;
wire n_1649;
wire n_1650;
wire n_1651;
wire n_1652;
wire n_1653;
wire n_1654;
wire n_1655;
wire n_1656;
wire n_1657;
wire n_1658;
wire n_1659;
wire n_1660;
wire n_1661;
wire n_1662;
wire n_1663;
wire n_1664;
wire n_1665;
wire n_1666;
wire n_1667;
wire n_1668;
wire n_1669;
wire n_1670;
wire n_1671;
wire n_1672;
wire n_1673;
wire n_1674;
wire n_1675;
wire n_1676;
wire n_1677;
wire n_1678;
wire n_1679;
wire n_1680;
wire n_1681;
wire n_1682;
wire n_1683;
wire n_1684;
wire n_1685;
wire n_1686;
wire n_1687;
wire n_1688;
wire n_1689;
wire n_1690;
wire n_1691;
wire n_1692;
wire n_1693;
wire n_1694;
wire n_1695;
wire n_1696;
wire n_1697;
wire n_1698;
wire n_1699;
wire n_1700;
wire n_1701;
wire n_1702;
wire n_1703;
wire n_1704;
wire n_1705;
wire n_1706;
wire n_1707;
wire n_1708;
wire n_1709;
wire n_1710;
wire n_1711;
wire n_1712;
wire n_1713;
wire n_1714;
wire n_1715;
wire n_1716;
wire n_1717;
wire n_1718;
wire n_1719;
wire n_1720;
wire n_1721;
wire n_1722;
wire n_1723;
wire n_1724;
wire n_1725;
wire n_1726;
wire n_1727;
wire n_1728;
wire n_1729;
wire n_1730;
wire n_1731;
wire n_1732;
wire n_1733;
wire n_1734;
wire n_1735;
wire n_1736;
wire n_1737;
wire n_1738;
wire n_1739;
wire n_1740;
wire n_1741;
wire n_1742;
wire n_1743;
wire n_1744;
wire n_1745;
wire n_1746;
wire n_1747;
wire n_1748;
wire n_1749;
wire n_1750;
wire n_1751;
wire n_1752;
wire n_1753;
wire n_1754;
wire n_1755;
wire n_1756;
wire n_1757;
wire n_1758;
wire n_1759;
wire n_1760;
wire n_1761;
wire n_1762;
wire n_1763;
wire n_1764;
wire n_1765;
wire n_1766;
wire n_1767;
wire n_1768;
wire n_1769;
wire n_1770;
wire n_1771;
wire n_1772;
wire n_1773;
wire n_1774;
wire n_1775;
wire n_1776;
wire n_1777;
wire n_1778;
wire n_1779;
wire n_1780;
wire n_1781;
wire n_1782;
wire n_1783;
wire n_1784;
wire n_1785;
wire n_1786;
wire n_1787;
wire n_1788;
wire n_1789;
wire n_1790;
wire n_1791;
wire n_1792;
wire n_1793;
wire n_1794;
wire n_1795;
wire n_1796;
wire n_1797;
wire n_1798;
wire n_1799;
wire n_1800;
wire n_1801;
wire n_1802;
wire n_1803;
wire n_1804;
wire n_1805;
wire n_1806;
wire n_1807;
wire n_1808;
wire n_1809;
wire n_1810;
wire n_1811;
wire n_1812;
wire n_1813;
wire n_1814;
wire n_1815;
wire n_1816;
wire n_1817;
wire n_1818;
wire n_1819;
wire n_1820;
wire n_1821;
wire n_1822;
wire n_1823;
wire n_1824;
wire n_1825;
wire n_1826;
wire n_1827;
wire n_1828;
wire n_1829;
wire n_1830;
wire n_1831;
wire n_1832;
wire n_1833;
wire n_1834;
wire n_1835;
wire n_1836;
wire n_1837;
wire n_1838;
wire n_1839;
wire n_1840;
wire n_1841;
wire n_1842;
wire n_1843;
wire n_1844;
wire n_1845;
wire n_1846;
wire n_1847;
wire n_1848;
wire n_1849;
wire n_1850;
wire n_1851;
wire n_1852;
wire n_1853;
wire n_1854;
wire n_1855;
wire n_1856;
wire n_1857;
wire n_1858;
wire n_1859;
wire n_1860;
wire n_1861;
wire n_1862;
wire n_1863;
wire n_1864;
wire n_1865;
wire n_1866;
wire n_1867;
wire n_1868;
wire n_1869;
wire n_1870;
wire n_1871;
wire n_1872;
wire n_1873;
wire n_1874;
wire n_1875;
wire n_1876;
wire n_1877;
wire n_1878;
wire n_1879;
wire n_1880;
wire n_1881;
wire n_1882;
wire n_1883;
wire n_1884;
wire n_1885;
wire n_1886;
wire n_1887;
wire n_1888;
wire n_1889;
wire n_1890;
wire n_1891;
wire n_1892;
wire n_1893;
wire n_1894;
wire n_1895;
wire n_1896;
wire n_1897;
wire n_1898;
wire n_1899;
wire n_1900;
wire n_1901;
wire n_1902;
wire n_1903;
wire n_1904;
wire n_1905;
wire n_1906;
wire n_1907;
wire n_1908;
wire n_1909;
wire n_1910;
wire n_1911;
wire n_1912;
wire n_1913;
wire n_1914;
wire n_1915;
wire n_1916;
wire n_1917;
wire n_1918;
wire n_1919;
wire n_1920;
wire n_1921;
wire n_1922;
wire n_1923;
wire n_1924;
wire n_1925;
wire n_1926;
wire n_1927;
wire n_1928;
wire n_1929;
wire n_1930;
wire n_1931;
wire n_1932;
wire n_1933;
wire n_1934;
wire n_1935;
wire n_1936;
wire n_1937;
wire n_1938;
wire n_1939;
wire n_1940;
wire n_1941;
wire n_1942;
wire n_1943;
wire n_1944;
wire n_1945;
wire n_1946;
wire n_1947;
wire n_1948;
wire n_1949;
wire n_1950;
wire n_1951;
wire n_1952;
wire n_1953;
wire n_1954;
wire n_1955;
wire n_1956;
wire n_1957;
wire n_1958;
wire n_1959;
wire n_1960;
wire n_1961;
wire n_1962;
wire n_1963;
wire n_1964;
wire n_1965;
wire n_1966;
wire n_1967;
wire n_1968;
wire n_1969;
wire n_1970;
wire n_1971;
wire n_1972;
wire n_1973;
wire n_1974;
wire n_1975;
wire n_1976;
wire n_1977;
wire n_1978;
wire n_1979;
wire n_1980;
wire n_1981;
wire n_1982;
wire n_1983;
wire n_1984;
wire n_1985;
wire n_1986;
wire n_1987;
wire n_1988;
wire n_1989;
wire n_1990;
wire n_1991;
wire n_1992;
wire n_1993;
wire n_1994;
wire n_1995;
wire n_1996;
wire n_1997;
wire n_1998;
wire n_1999;
wire n_2000;
wire n_2001;
wire n_2002;
wire n_2003;
wire n_2004;
wire n_2005;
wire n_2006;
wire n_2007;
wire n_2008;
wire n_2009;
wire n_2010;
wire n_2011;
wire n_2012;
wire n_2013;
wire n_2014;
wire n_2015;
wire n_2016;
wire n_2017;
wire n_2018;
wire n_2019;
wire n_2020;
wire n_2021;
wire n_2022;
wire n_2023;
wire n_2024;
wire n_2025;
wire n_2026;
wire n_2027;
wire n_2028;
wire n_2029;
wire n_2030;
wire n_2031;
wire n_2032;
wire n_2033;
wire n_2034;
wire n_2035;
wire n_2036;
wire n_2037;
wire n_2038;
wire n_2039;
wire n_2040;
wire n_2041;
wire n_2042;
wire n_2043;
wire n_2044;
wire n_2045;
wire n_2046;
wire n_2047;
wire n_2048;
wire n_2049;
wire n_2050;
wire n_2051;
wire n_2052;
wire n_2053;
wire n_2054;
wire n_2055;
wire n_2056;
wire n_2057;
wire n_2058;
wire n_2059;
wire n_2060;
wire n_2061;
wire n_2062;
wire n_2063;
wire n_2064;
wire n_2065;
wire n_2066;
wire n_2067;
wire n_2068;
wire n_2069;
wire n_2070;
wire n_2071;
wire n_2072;
wire n_2073;
wire n_2074;
wire n_2075;
wire n_2076;
wire n_2077;
wire n_2078;
wire n_2079;
wire n_2080;
wire n_2081;
wire n_2082;
wire n_2083;
wire n_2084;
wire n_2085;
wire n_2086;
wire n_2087;
wire n_2088;
wire n_2089;
wire n_2090;
wire n_2091;
wire n_2092;
wire n_2093;
wire n_2094;
wire n_2095;
wire n_2096;
wire n_2097;
wire n_2098;
wire n_2099;
wire n_2100;
wire n_2101;
wire n_2102;
wire n_2103;
wire n_2104;
wire n_2105;
wire n_2106;
wire n_2107;
wire n_2108;
wire n_2109;
wire n_2110;
wire n_2111;
wire n_2112;
wire n_2113;
wire n_2114;
wire n_2115;
wire n_2116;
wire n_2117;
wire n_2118;
wire n_2119;
wire n_2120;
wire n_2121;
wire n_2122;
wire n_2123;
wire n_2124;
wire n_2125;
wire n_2126;
wire n_2127;
wire n_2128;
wire n_2129;
wire n_2130;
wire n_2131;
wire n_2132;
wire n_2133;
wire n_2134;
wire n_2135;
wire n_2136;
wire n_2137;
wire n_2138;
wire n_2139;
wire n_2140;
wire n_2141;
wire n_2142;
wire n_2143;
wire n_2144;
wire n_2145;
wire n_2146;
wire n_2147;
wire n_2148;
wire n_2149;
wire n_2150;
wire n_2151;
wire n_2152;
wire n_2153;
wire n_2154;
wire n_2155;
wire n_2156;
wire n_2157;
wire n_2158;
wire n_2159;
wire n_2160;
wire n_2161;
wire n_2162;
wire n_2163;
wire n_2164;
wire n_2165;
wire n_2166;
wire n_2167;
wire n_2168;
wire n_2169;
wire n_2170;
wire n_2171;
wire n_2172;
wire n_2173;
wire n_2174;
wire n_2175;
wire n_2176;
wire n_2177;
wire n_2178;
wire n_2179;
wire n_2180;
wire n_2181;
wire n_2182;
wire n_2183;
wire n_2184;
wire n_2185;
wire n_2186;
wire n_2187;
wire n_2188;
wire n_2189;
wire n_2190;
wire n_2191;
wire n_2192;
wire n_2193;
wire n_2194;
wire n_2195;
wire n_2196;
wire n_2197;
wire n_2198;
wire n_2199;
wire n_2200;
wire n_2201;
wire n_2202;
wire n_2203;
wire n_2204;
wire n_2205;
wire n_2206;
wire n_2207;
wire n_2208;
wire n_2209;
wire n_2210;
wire n_2211;
wire n_2212;
wire n_2213;
wire n_2214;
wire n_2215;
wire n_2216;
wire n_2217;
wire n_2218;
wire n_2219;
wire n_2220;
wire n_2221;
wire n_2222;
wire n_2223;
wire n_2224;
wire n_2225;
wire n_2226;
wire n_2227;
wire n_2228;
wire n_2229;
wire n_2230;
wire n_2231;
wire n_2232;
wire n_2233;
wire n_2234;
wire n_2235;
wire n_2236;
wire n_2237;
wire n_2238;
wire n_2239;
wire n_2240;
wire n_2241;
wire n_2242;
wire n_2243;
wire n_2244;
wire n_2245;
wire n_2246;
wire n_2247;
wire n_2248;
wire n_2249;
wire n_2250;
wire n_2251;
wire n_2252;
wire n_2253;
wire n_2254;
wire n_2255;
wire n_2256;
wire n_2257;
wire n_2258;
wire n_2259;
wire n_2260;
wire n_2261;
wire n_2262;
wire n_2263;
wire n_2264;
wire n_2265;
wire n_2266;
wire n_2267;
wire n_2268;
wire n_2269;
wire n_2270;
wire n_2271;
wire n_2272;
wire n_2273;
wire n_2274;
wire n_2275;
wire n_2276;
wire n_2277;
wire n_2278;
wire n_2279;
wire n_2280;
wire n_2281;
wire n_2282;
wire n_2283;
wire n_2284;
wire n_2285;
wire n_2286;
wire n_2287;
wire n_2288;
wire n_2289;
wire n_2290;
wire n_2291;
wire n_2292;
wire n_2293;
wire n_2294;
wire n_2295;
wire n_2296;
wire n_2297;
wire n_2298;
wire n_2299;
wire n_2300;
wire n_2301;
wire n_2302;
wire n_2303;
wire n_2304;
wire n_2305;
wire n_2306;
wire n_2307;
wire n_2308;
wire n_2309;
wire n_2310;
wire n_2311;
wire n_2312;
wire n_2313;
wire n_2314;
wire n_2315;
wire n_2316;
wire n_2317;
wire n_2318;
wire n_2319;
wire n_2320;
wire n_2321;
wire n_2322;
wire n_2323;
wire n_2324;
wire n_2325;
wire n_2326;
wire n_2327;
wire n_2328;
wire n_2329;
wire n_2330;
wire n_2331;
wire n_2332;
wire n_2333;
wire n_2334;
wire n_2335;
wire n_2336;
wire n_2337;
wire n_2338;
wire n_2339;
wire n_2340;
wire n_2341;
wire n_2342;
wire n_2343;
wire n_2344;
wire n_2345;
wire n_2346;
wire n_2347;
wire n_2348;
wire n_2349;
wire n_2350;
wire n_2351;
wire n_2352;
wire n_2353;
wire n_2354;
wire n_2355;
wire n_2356;
wire n_2357;
wire n_2358;
wire n_2359;
wire n_2360;
wire n_2361;
wire n_2362;
wire n_2363;
wire n_2364;
wire n_2365;
wire n_2366;
wire n_2367;
wire n_2368;
wire n_2369;
wire n_2370;
wire n_2371;
wire n_2372;
wire n_2373;
wire n_2374;
wire n_2375;
wire n_2376;
wire n_2377;
wire n_2378;
wire n_2379;
wire n_2380;
wire n_2381;
wire n_2382;
wire n_2383;
wire n_2384;
wire n_2385;
wire n_2386;
wire n_2387;
wire n_2388;
wire n_2389;
wire n_2390;
wire n_2391;
wire n_2392;
wire n_2393;
wire n_2394;
wire n_2395;
wire n_2396;
wire n_2397;
wire n_2398;
wire n_2399;
wire n_2400;
wire n_2401;
wire n_2402;
wire n_2403;
wire n_2404;
wire n_2405;
wire n_2406;
wire n_2407;
wire n_2408;
wire n_2409;
wire n_2410;
wire n_2411;
wire n_2412;
wire n_2413;
wire n_2414;
wire n_2415;
wire n_2416;
wire n_2417;
wire n_2418;
wire n_2419;
wire n_2420;
wire n_2421;
wire n_2422;
wire n_2423;
wire n_2424;
wire n_2425;
wire n_2426;
wire n_2427;
wire n_2428;
wire n_2429;
wire n_2430;
wire n_2431;
wire n_2432;
wire n_2433;
wire n_2434;
wire n_2435;
wire n_2436;
wire n_2437;
wire n_2438;
wire n_2439;
wire n_2440;
wire n_2441;
wire n_2442;
wire n_2443;
wire n_2444;
wire n_2445;
wire n_2446;
wire n_2447;
wire n_2448;
wire n_2449;
wire n_2450;
wire n_2451;
wire n_2452;
wire n_2453;
wire n_2454;
wire n_2455;
wire n_2456;
wire n_2457;
wire n_2458;
wire n_2459;
wire n_2460;
wire n_2461;
wire n_2462;
wire n_2463;
wire n_2464;
wire n_2465;
wire n_2466;
wire n_2467;
wire n_2468;
wire n_2469;
wire n_2470;
wire n_2471;
wire n_2472;
wire n_2473;
wire n_2474;
wire n_2475;
wire n_2476;
wire n_2477;
wire n_2478;
wire n_2479;
wire n_2480;
wire n_2481;
wire n_2482;
wire n_2483;
wire n_2484;
wire n_2485;
wire n_2486;
wire n_2487;
wire n_2488;
wire n_2489;
wire n_2490;
wire n_2491;
wire n_2492;
wire n_2493;
wire n_2494;
wire n_2495;
wire n_2496;
wire n_2497;
wire n_2498;
wire n_2499;
wire n_2500;
wire n_2501;
wire n_2502;
wire n_2503;
wire n_2504;
wire n_2505;
wire n_2506;
wire n_2507;
wire n_2508;
wire n_2509;
wire n_2510;
wire n_2511;
wire n_2512;
wire n_2513;
wire n_2514;
wire n_2515;
wire n_2516;
wire n_2517;
wire n_2518;
wire n_2519;
wire n_2520;
wire n_2521;
wire n_2522;
wire n_2523;
wire n_2524;
wire n_2525;
wire n_2526;
wire n_2527;
wire n_2528;
wire n_2529;
wire n_2530;
wire n_2531;
wire n_2532;
wire n_2533;
wire n_2534;
wire n_2535;
wire n_2536;
wire n_2537;
wire n_2538;
wire n_2539;
wire n_2540;
wire n_2541;
wire n_2542;
wire n_2543;
wire n_2544;
wire n_2545;
wire n_2546;
wire n_2547;
wire n_2548;
wire n_2549;
wire n_2550;
wire n_2551;
wire n_2552;
wire n_2553;
wire n_2554;
wire n_2555;
wire n_2556;
wire n_2557;
wire n_2558;
wire n_2559;
wire n_2560;
wire n_2561;
wire n_2562;
wire n_2563;
wire n_2564;
wire n_2565;
wire n_2566;
wire n_2567;
wire n_2568;
wire n_2569;
wire n_2570;
wire n_2571;
wire n_2572;
wire n_2573;
wire n_2574;
wire n_2575;
wire n_2576;
wire n_2577;
wire n_2578;
wire n_2579;
wire n_2580;
wire n_2581;
wire n_2582;
wire n_2583;
wire n_2584;
wire n_2585;
wire n_2586;
wire n_2587;
wire n_2588;
wire n_2589;
wire n_2590;
wire n_2591;
wire n_2592;
wire n_2593;
wire n_2594;
wire n_2595;
wire n_2596;
wire n_2597;
wire n_2598;
wire n_2599;
wire n_2600;
wire n_2601;
wire n_2602;
wire n_2603;
wire n_2604;
wire n_2605;
wire n_2606;
wire n_2607;
wire n_2608;
wire n_2609;
wire n_2610;
wire n_2611;
wire n_2612;
wire n_2613;
wire n_2614;
wire n_2615;
wire n_2616;
wire n_2617;
wire n_2618;
wire n_2619;
wire n_2620;
wire n_2621;
wire n_2622;
wire n_2623;
wire n_2624;
wire n_2625;
wire n_2626;
wire n_2627;
wire n_2628;
wire n_2629;
wire n_2630;
wire n_2631;
wire n_2632;
wire n_2633;
wire n_2634;
wire n_2635;
wire n_2636;
wire n_2637;
wire n_2638;
wire n_2639;
wire n_2640;
wire n_2641;
wire n_2642;
wire n_2643;
wire n_2644;
wire n_2645;
wire n_2646;
wire n_2647;
wire n_2648;
wire n_2649;
wire n_2650;
wire n_2651;
wire n_2652;
wire n_2653;
wire n_2654;
wire n_2655;
wire n_2656;
wire n_2657;
wire n_2658;
wire n_2659;
wire n_2660;
wire n_2661;
wire n_2662;
wire n_2663;
wire n_2664;
wire n_2665;
wire n_2666;
wire n_2667;
wire n_2668;
wire n_2669;
wire n_2670;
wire n_2671;
wire n_2672;
wire n_2673;
wire n_2674;
wire n_2675;
wire n_2676;
wire n_2677;
wire n_2678;
wire n_2679;
wire n_2680;
wire n_2681;
wire n_2682;
wire n_2683;
wire n_2684;
wire n_2685;
wire n_2686;
wire n_2687;
wire n_2688;
wire n_2689;
wire n_2690;
wire n_2691;
wire n_2692;
wire n_2693;
wire n_2694;
wire n_2695;
wire n_2696;
wire n_2697;
wire n_2698;
wire n_2699;
wire n_2700;
wire n_2701;
wire n_2702;
wire n_2703;
wire n_2704;
wire n_2705;
wire n_2706;
wire n_2707;
wire n_2708;
wire n_2709;
wire n_2710;
wire n_2711;
wire n_2712;
wire n_2713;
wire n_2714;
wire n_2715;
wire n_2716;
wire n_2717;
wire n_2718;
wire n_2719;
wire n_2720;
wire n_2721;
wire n_2722;
wire n_2723;
wire n_2724;
wire n_2725;
wire n_2726;
wire n_2727;
wire n_2728;
wire n_2729;
wire n_2730;
wire n_2731;
wire n_2732;
wire n_2733;
wire n_2734;
wire n_2735;
wire n_2736;
wire n_2737;
wire n_2738;
wire n_2739;
wire n_2740;
wire n_2741;
wire n_2742;
wire n_2743;
wire n_2744;
wire n_2745;
wire n_2746;
wire n_2747;
wire n_2748;
wire n_2749;
wire n_2750;
wire n_2751;
wire n_2752;
wire n_2753;
wire n_2754;
wire n_2755;
wire n_2756;
wire n_2757;
wire n_2758;
wire n_2759;
wire n_2760;
wire n_2761;
wire n_2762;
wire n_2763;
wire n_2764;
wire n_2765;
wire n_2766;
wire n_2767;
wire n_2768;
wire n_2769;
wire n_2770;
wire n_2771;
wire n_2772;
wire n_2773;
wire n_2774;
wire n_2775;
wire n_2776;
wire n_2777;
wire n_2778;
wire n_2779;
wire n_2780;
wire n_2781;
wire n_2782;
wire n_2783;
wire n_2784;
wire n_2785;
wire n_2786;
wire n_2787;
wire n_2788;
wire n_2789;
wire n_2790;
wire n_2791;
wire n_2792;
wire n_2793;
wire n_2794;
wire n_2795;
wire n_2796;
wire n_2797;
wire n_2798;
wire n_2799;
wire n_2800;
wire n_2801;
wire n_2802;
wire n_2803;
wire n_2804;
wire n_2805;
wire n_2806;
wire n_2807;
wire n_2808;
wire n_2809;
wire n_2810;
wire n_2811;
wire n_2812;
wire n_2813;
wire n_2814;
wire n_2815;
wire n_2816;
wire n_2817;
wire n_2818;
wire n_2819;
wire n_2820;
wire n_2821;
wire n_2822;
wire n_2823;
wire n_2824;
wire n_2825;
wire n_2826;
wire n_2827;
wire n_2828;
wire n_2829;
wire n_2830;
wire n_2831;
wire n_2832;
wire n_2833;
wire n_2834;
wire n_2835;
wire n_2836;
wire n_2837;
wire n_2838;
wire n_2839;
wire n_2840;
wire n_2841;
wire n_2842;
wire n_2843;
wire n_2844;
wire n_2845;
wire n_2846;
wire n_2847;
wire n_2848;
wire n_2849;
wire n_2850;
wire n_2851;
wire n_2852;
wire n_2853;
wire n_2854;
wire n_2855;
wire n_2856;
wire n_2857;
wire n_2858;
wire n_2859;
wire n_2860;
wire n_2861;
wire n_2862;
wire n_2863;
wire n_2864;
wire n_2865;
wire n_2866;
wire n_2867;
wire n_2868;
wire n_2869;
wire n_2870;
wire n_2871;
wire n_2872;
wire n_2873;
wire n_2874;
wire n_2875;
wire n_2876;
wire n_2877;
wire n_2878;
wire n_2879;
wire n_2880;
wire n_2881;
wire n_2882;
wire n_2883;
wire n_2884;
wire n_2885;
wire n_2886;
wire n_2887;
wire n_2888;
wire n_2889;
wire n_2890;
wire n_2891;
wire n_2892;
wire n_2893;
wire n_2894;
wire n_2895;
wire n_2896;
wire n_2897;
wire n_2898;
wire n_2899;
wire n_2900;
wire n_2901;
wire n_2902;
wire n_2903;
wire n_2904;
wire n_2905;
wire n_2906;
wire n_2907;
wire n_2908;
wire n_2909;
wire n_2910;
wire n_2911;
wire n_2912;
wire n_2913;
wire n_2914;
wire n_2915;
wire n_2916;
wire n_2917;
wire n_2918;
wire n_2919;
wire n_2920;
wire n_2921;
wire n_2922;
wire n_2923;
wire n_2924;
wire n_2925;
wire n_2926;
wire n_2927;
wire n_2928;
wire n_2929;
wire n_2930;
wire n_2931;
wire n_2932;
wire n_2933;
wire n_2934;
wire n_2935;
wire n_2936;
wire n_2937;
wire n_2938;
wire n_2939;
wire n_2940;
wire n_2941;
wire n_2942;
wire n_2943;
wire n_2944;
wire n_2945;
wire n_2946;
wire n_2947;
wire n_2948;
wire n_2949;
wire n_2950;
wire n_2951;
wire n_2952;
wire n_2953;
wire n_2954;
wire n_2955;
wire n_2956;
wire n_2957;
wire n_2958;
wire n_2959;
wire n_2960;
wire n_2961;
wire n_2962;
wire n_2963;
wire n_2964;
wire n_2965;
wire n_2966;
wire n_2967;
wire n_2968;
wire n_2969;
wire n_2970;
wire n_2971;
wire n_2972;
wire n_2973;
wire n_2974;
wire n_2975;
wire n_2976;
wire n_2977;
wire n_2978;
wire n_2979;
wire n_2980;
wire n_2981;
wire n_2982;
wire n_2983;
wire n_2984;
wire n_2985;
wire n_2986;
wire n_2987;
wire n_2988;
wire n_2989;
wire n_2990;
wire n_2991;
wire n_2992;
wire n_2993;
wire n_2994;
wire n_2995;
wire n_2996;
wire n_2997;
wire n_2998;
wire n_2999;
wire n_3000;
wire n_3001;
wire n_3002;
wire n_3003;
wire n_3004;
wire n_3005;
wire n_3006;
wire n_3007;
wire n_3008;
wire n_3009;
wire n_3010;
wire n_3011;
wire n_3012;
wire n_3013;
wire n_3014;
wire n_3015;
wire n_3016;
wire n_3017;
wire n_3018;
wire n_3019;
wire n_3020;
wire n_3021;
wire n_3022;
wire n_3023;
wire n_3024;
wire n_3025;
wire n_3026;
wire n_3027;
wire n_3028;
wire n_3029;
wire n_3030;
wire n_3031;
wire n_3032;
wire n_3033;
wire n_3034;
wire n_3035;
wire n_3036;
wire n_3037;
wire n_3038;
wire n_3039;
wire n_3040;
wire n_3041;
wire n_3042;
wire n_3043;
wire n_3044;
wire n_3045;
wire n_3046;
wire n_3047;
wire n_3048;
wire n_3049;
wire n_3050;
wire n_3051;
wire n_3052;
wire n_3053;
wire n_3054;
wire n_3055;
wire n_3056;
wire n_3057;
wire n_3058;
wire n_3059;
wire n_3060;
wire n_3061;
wire n_3062;
wire n_3063;
wire n_3064;
wire n_3065;
wire n_3066;
wire n_3067;
wire n_3068;
wire n_3069;
wire n_3070;
wire n_3071;
wire n_3072;
wire n_3073;
wire n_3074;
wire n_3075;
wire n_3076;
wire n_3077;
wire n_3078;
wire n_3079;
wire n_3080;
wire n_3081;
wire n_3082;
wire n_3083;
wire n_3084;
wire n_3085;
wire n_3086;
wire n_3087;
wire n_3088;
wire n_3089;
wire n_3090;
wire n_3091;
wire n_3092;
wire n_3093;
wire n_3094;
wire n_3095;
wire n_3096;
wire n_3097;
wire n_3098;
wire n_3099;
wire n_3100;
wire n_3101;
wire n_3102;
wire n_3103;
wire n_3104;
wire n_3105;
wire n_3106;
wire n_3107;
wire n_3108;
wire n_3109;
wire n_3110;
wire n_3111;
wire n_3112;
wire n_3113;
wire n_3114;
wire n_3115;
wire n_3116;
wire n_3117;
wire n_3118;
wire n_3119;
wire n_3120;
wire n_3121;
wire n_3122;
wire n_3123;
wire n_3124;
wire n_3125;
wire n_3126;
wire n_3127;
wire n_3128;
wire n_3129;
wire n_3130;
wire n_3131;
wire n_3132;
wire n_3133;
wire n_3134;
wire n_3135;
wire n_3136;
wire n_3137;
wire n_3138;
wire n_3139;
wire n_3140;
wire n_3141;
wire n_3142;
wire n_3143;
wire n_3144;
wire n_3145;
wire n_3146;
wire n_3147;
wire n_3148;
wire n_3149;
wire n_3150;
wire n_3151;
wire n_3152;
wire n_3153;
wire n_3154;
wire n_3155;
wire n_3156;
wire n_3157;
wire n_3158;
wire n_3159;
wire n_3160;
wire n_3161;
wire n_3162;
wire n_3163;
wire n_3164;
wire n_3165;
wire n_3166;
wire n_3167;
wire n_3168;
wire n_3169;
wire n_3170;
wire n_3171;
wire n_3172;
wire n_3173;
wire n_3174;
wire n_3175;
wire n_3176;
wire n_3177;
wire n_3178;
wire n_3179;
wire n_3180;
wire n_3181;
wire n_3182;
wire n_3183;
wire n_3184;
wire n_3185;
wire n_3186;
wire n_3187;
wire n_3188;
wire n_3189;
wire n_3190;
wire n_3191;
wire n_3192;
wire n_3193;
wire n_3194;
wire n_3195;
wire n_3196;
wire n_3197;
wire n_3198;
wire n_3199;
wire n_3200;
wire n_3201;
wire n_3202;
wire n_3203;
wire n_3204;
wire n_3205;
wire n_3206;
wire n_3207;
wire n_3208;
wire n_3209;
wire n_3210;
wire n_3211;
wire n_3212;
wire n_3213;
wire n_3214;
wire n_3215;
wire n_3216;
wire n_3217;
wire n_3218;
wire n_3219;
wire n_3220;
wire n_3221;
wire n_3222;
wire n_3223;
wire n_3224;
wire n_3225;
wire n_3226;
wire n_3227;
wire n_3228;
wire n_3229;
wire n_3230;
wire n_3231;
wire n_3232;
wire n_3233;
wire n_3234;
wire n_3235;
wire n_3236;
wire n_3237;
wire n_3238;
wire n_3239;
wire n_3240;
wire n_3241;
wire n_3242;
wire n_3243;
wire n_3244;
wire n_3245;
wire n_3246;
wire n_3247;
wire n_3248;
wire n_3249;
wire n_3250;
wire n_3251;
wire n_3252;
wire n_3253;
wire n_3254;
wire n_3255;
wire n_3256;
wire n_3257;
wire n_3258;
wire n_3259;
wire n_3260;
wire n_3261;
wire n_3262;
wire n_3263;
wire n_3264;
wire n_3265;
wire n_3266;
wire n_3267;
wire n_3268;
wire n_3269;
wire n_3270;
wire n_3271;
wire n_3272;
wire n_3273;
wire n_3274;
wire n_3275;
wire n_3276;
wire n_3277;
wire n_3278;
wire n_3279;
wire n_3280;
wire n_3281;
wire n_3282;
wire n_3283;
wire n_3284;
wire n_3285;
wire n_3286;
wire n_3287;
wire n_3288;
wire n_3289;
wire n_3290;
wire n_3291;
wire n_3292;
wire n_3293;
wire n_3294;
wire n_3295;
wire n_3296;
wire n_3297;
wire n_3298;
wire n_3299;
wire n_3300;
wire n_3301;
wire n_3302;
wire n_3303;
wire n_3304;
wire n_3305;
wire n_3306;
wire n_3307;
wire n_3308;
wire n_3309;
wire n_3310;
wire n_3311;
wire n_3312;
wire n_3313;
wire n_3314;
wire n_3315;
wire n_3316;
wire n_3317;
wire n_3318;
wire n_3319;
wire n_3320;
wire n_3321;
wire n_3322;
wire n_3323;
wire n_3324;
wire n_3325;
wire n_3326;
wire n_3327;
wire n_3328;
wire n_3329;
wire n_3330;
wire n_3331;
wire n_3332;
wire n_3333;
wire n_3334;
wire n_3335;
wire n_3336;
wire n_3337;
wire n_3338;
wire n_3339;
wire n_3340;
wire n_3341;
wire n_3342;
wire n_3343;
wire n_3344;
wire n_3345;
wire n_3346;
wire n_3347;
wire n_3348;
wire n_3349;
wire n_3350;
wire n_3351;
wire n_3352;
wire n_3353;
wire n_3354;
wire n_3355;
wire n_3356;
wire n_3357;
wire n_3358;
wire n_3359;
wire n_3360;
wire n_3361;
wire n_3362;
wire n_3363;
wire n_3364;
wire n_3365;
wire n_3366;
wire n_3367;
wire n_3368;
wire n_3369;
wire n_3370;
wire n_3371;
wire n_3372;
wire n_3373;
wire n_3374;
wire n_3375;
wire n_3376;
wire n_3377;
wire n_3378;
wire n_3379;
wire n_3380;
wire n_3381;
wire n_3382;
wire n_3383;
wire n_3384;
wire n_3385;
wire n_3386;
wire n_3387;
wire n_3388;
wire n_3389;
wire n_3390;
wire n_3391;
wire n_3392;
wire n_3393;
wire n_3394;
wire n_3395;
wire n_3396;
wire n_3397;
wire n_3398;
wire n_3399;
wire n_3400;
wire n_3401;
wire n_3402;
wire n_3403;
wire n_3404;
wire n_3405;
wire n_3406;
wire n_3407;
wire n_3408;
wire n_3409;
wire n_3410;
wire n_3411;
wire n_3412;
wire n_3413;
wire n_3414;
wire n_3415;
wire n_3416;
wire n_3417;
wire n_3418;
wire n_3419;
wire n_3420;
wire n_3421;
wire n_3422;
wire n_3423;
wire n_3424;
wire n_3425;
wire n_3426;
wire n_3427;
wire n_3428;
wire n_3429;
wire n_3430;
wire n_3431;
wire n_3432;
wire n_3433;
wire n_3434;
wire n_3435;
wire n_3436;
wire n_3437;
wire n_3438;
wire n_3439;
wire n_3440;
wire n_3441;
wire n_3442;
wire n_3443;
wire n_3444;
wire n_3445;
wire n_3446;
wire n_3447;
wire n_3448;
wire n_3449;
wire n_3450;
wire n_3451;
wire n_3452;
wire n_3453;
wire n_3454;
wire n_3455;
wire n_3456;
wire n_3457;
wire n_3458;
wire n_3459;
wire n_3460;
wire n_3461;
wire n_3462;
wire n_3463;
wire n_3464;
wire n_3465;
wire n_3466;
wire n_3467;
wire n_3468;
wire n_3469;
wire n_3470;
wire n_3471;
wire n_3472;
wire n_3473;
wire n_3474;
wire n_3475;
wire n_3476;
wire n_3477;
wire n_3478;
wire n_3479;
wire n_3480;
wire n_3481;
wire n_3482;
wire n_3483;
wire n_3484;
wire n_3485;
wire n_3486;
wire n_3487;
wire n_3488;
wire n_3489;
wire n_3490;
wire n_3491;
wire n_3492;
wire n_3493;
wire n_3494;
wire n_3495;
wire n_3496;
wire n_3497;
wire n_3498;
wire n_3499;
wire n_3500;
wire n_3501;
wire n_3502;
wire n_3503;
wire n_3504;
wire n_3505;
wire n_3506;
wire n_3507;
wire n_3508;
wire n_3509;
wire n_3510;
wire n_3511;
wire n_3512;
wire n_3513;
wire n_3514;
wire n_3515;
wire n_3516;
wire n_3517;
wire n_3518;
wire n_3519;
wire n_3520;
wire n_3521;
wire n_3522;
wire n_3523;
wire n_3524;
wire n_3525;
wire n_3526;
wire n_3527;
wire n_3528;
wire n_3529;
wire n_3530;
wire n_3531;
wire n_3532;
wire n_3533;
wire n_3534;
wire n_3535;
wire n_3536;
wire n_3537;
wire n_3538;
wire n_3539;
wire n_3540;
wire n_3541;
wire n_3542;
wire n_3543;
wire n_3544;
wire n_3545;
wire n_3546;
wire n_3547;
wire n_3548;
wire n_3549;
wire n_3550;
wire n_3551;
wire n_3552;
wire n_3553;
wire n_3554;
wire n_3555;
wire n_3556;
wire n_3557;
wire n_3558;
wire n_3559;
wire n_3560;
wire n_3561;
wire n_3562;
wire n_3563;
wire n_3564;
wire n_3565;
wire n_3566;
wire n_3567;
wire n_3568;
wire n_3569;
wire n_3570;
wire n_3571;
wire n_3572;
wire n_3573;
wire n_3574;
wire n_3575;
wire n_3576;
wire n_3577;
wire n_3578;
wire n_3579;
wire n_3580;
wire n_3581;
wire n_3582;
wire n_3583;
wire n_3584;
wire n_3585;
wire n_3586;
wire n_3587;
wire n_3588;
wire n_3589;
wire n_3590;
wire n_3591;
wire n_3592;
wire n_3593;
wire n_3594;
wire n_3595;
wire n_3596;
wire n_3597;
wire n_3598;
wire n_3599;
wire n_3600;
wire n_3601;
wire n_3602;
wire n_3603;
wire n_3604;
wire n_3605;
wire n_3606;
wire n_3607;
wire n_3608;
wire n_3609;
wire n_3610;
wire n_3611;
wire n_3612;
wire n_3613;
wire n_3614;
wire n_3615;
wire n_3616;
wire n_3617;
wire n_3618;
wire n_3619;
wire n_3620;
wire n_3621;
wire n_3622;
wire n_3623;
wire n_3624;
wire n_3625;
wire n_3626;
wire n_3627;
wire n_3628;
wire n_3629;
wire n_3630;
wire n_3631;
wire n_3632;
wire n_3633;
wire n_3634;
wire n_3635;
wire n_3636;
wire n_3637;
wire n_3638;
wire n_3639;
wire n_3640;
wire n_3641;
wire n_3642;
wire n_3643;
wire n_3644;
wire n_3645;
wire n_3646;
wire n_3647;
wire n_3648;
wire n_3649;
wire n_3650;
wire n_3651;
wire n_3652;
wire n_3653;
wire n_3654;
wire n_3655;
wire n_3656;
wire n_3657;
wire n_3658;
wire n_3659;
wire n_3660;
wire n_3661;
wire n_3662;
wire n_3663;
wire n_3664;
wire n_3665;
wire n_3666;
wire n_3667;
wire n_3668;
wire n_3669;
wire n_3670;
wire n_3671;
wire n_3672;
wire n_3673;
wire n_3674;
wire n_3675;
wire n_3676;
wire n_3677;
wire n_3678;
wire n_3679;
wire n_3680;
wire n_3681;
wire n_3682;
wire n_3683;
wire n_3684;
wire n_3685;
wire n_3686;
wire n_3687;
wire n_3688;
wire n_3689;
wire n_3690;
wire n_3691;
wire n_3692;
wire n_3693;
wire n_3694;
wire n_3695;
wire n_3696;
wire n_3697;
wire n_3698;
wire n_3699;
wire n_3700;
wire n_3701;
wire n_3702;
wire n_3703;
wire n_3704;
wire n_3705;
wire n_3706;
wire n_3707;
wire n_3708;
wire n_3709;
wire n_3710;
wire n_3711;
wire n_3712;
wire n_3713;
wire n_3714;
wire n_3715;
wire n_3716;
wire n_3717;
wire n_3718;
wire n_3719;
wire n_3720;
wire n_3721;
wire n_3722;
wire n_3723;
wire n_3724;
wire n_3725;
wire n_3726;
wire n_3727;
wire n_3728;
wire n_3729;
wire n_3730;
wire n_3731;
wire n_3732;
wire n_3733;
wire n_3734;
wire n_3735;
wire n_3736;
wire n_3737;
wire n_3738;
wire n_3739;
wire n_3740;
wire n_3741;
wire n_3742;
wire n_3743;
wire n_3744;
wire n_3745;
wire n_3746;
wire n_3747;
wire n_3748;
wire n_3749;
wire n_3750;
wire n_3751;
wire n_3752;
wire n_3753;
wire n_3754;
wire n_3755;
wire n_3756;
wire n_3757;
wire n_3758;
wire n_3759;
wire n_3760;
wire n_3761;
wire n_3762;
wire n_3763;
wire n_3764;
wire n_3765;
wire n_3766;
wire n_3767;
wire n_3768;
wire n_3769;
wire n_3770;
wire n_3771;
wire n_3772;
wire n_3773;
wire n_3774;
wire n_3775;
wire n_3776;
wire n_3777;
wire n_3778;
wire n_3779;
wire n_3780;
wire n_3781;
wire n_3782;
wire n_3783;
wire n_3784;
wire n_3785;
wire n_3786;
wire n_3787;
wire n_3788;
wire n_3789;
wire n_3790;
wire n_3791;
wire n_3792;
wire n_3793;
wire n_3794;
wire n_3795;
wire n_3796;
wire n_3797;
wire n_3798;
wire n_3799;
wire n_3800;
wire n_3801;
wire n_3802;
wire n_3803;
wire n_3804;
wire n_3805;
wire n_3806;
wire n_3807;
wire n_3808;
wire n_3809;
wire n_3810;
wire n_3811;
wire n_3812;
wire n_3813;
wire n_3814;
wire n_3815;
wire n_3816;
wire n_3817;
wire n_3818;
wire n_3819;
wire n_3820;
wire n_3821;
wire n_3822;
wire n_3823;
wire n_3824;
wire n_3825;
wire n_3826;
wire n_3827;
wire n_3828;
wire n_3829;
wire n_3830;
wire n_3831;
wire n_3832;
wire n_3833;
wire n_3834;
wire n_3835;
wire n_3836;
wire n_3837;
wire n_3838;
wire n_3839;
wire n_3840;
wire n_3841;
wire n_3842;
wire n_3843;
wire n_3844;
wire n_3845;
wire n_3846;
wire n_3847;
wire n_3848;
wire n_3849;
wire n_3850;
wire n_3851;
wire n_3852;
wire n_3853;
wire n_3854;
wire n_3855;
wire n_3856;
wire n_3857;
wire n_3858;
wire n_3859;
wire n_3860;
wire n_3861;
wire n_3862;
wire n_3863;
wire n_3864;
wire n_3865;
wire n_3866;
wire n_3867;
wire n_3868;
wire n_3869;
wire n_3870;
wire n_3871;
wire n_3872;
wire n_3873;
wire n_3874;
wire n_3875;
wire n_3876;
wire n_3877;
wire n_3878;
wire n_3879;
wire n_3880;
wire n_3881;
wire n_3882;
wire n_3883;
wire n_3884;
wire n_3885;
wire n_3886;
wire n_3887;
wire n_3888;
wire n_3889;
wire n_3890;
wire n_3891;
wire n_3892;
wire n_3893;
wire n_3894;
wire n_3895;
wire n_3896;
wire n_3897;
wire n_3898;
wire n_3899;
wire n_3900;
wire n_3901;
wire n_3902;
wire n_3903;
wire n_3904;
wire n_3905;
wire n_3906;
wire n_3907;
wire n_3908;
wire n_3909;
wire n_3910;
wire n_3911;
wire n_3912;
wire n_3913;
wire n_3914;
wire n_3915;
wire n_3916;
wire n_3917;
wire n_3918;
wire n_3919;
wire n_3920;
wire n_3921;
wire n_3922;
wire n_3923;
wire n_3924;
wire n_3925;
wire n_3926;
wire n_3927;
wire n_3928;
wire n_3929;
wire n_3930;
wire n_3931;
wire n_3932;
wire n_3933;
wire n_3934;
wire n_3935;
wire n_3936;
wire n_3937;
wire n_3938;
wire n_3939;
wire n_3940;
wire n_3941;
wire n_3942;
wire n_3943;
wire n_3944;
wire n_3945;
wire n_3946;
wire n_3947;
wire n_3948;
wire n_3949;
wire n_3950;
wire n_3951;
wire n_3952;
wire n_3953;
wire n_3954;
wire n_3955;
wire n_3956;
wire n_3957;
wire n_3958;
wire n_3959;
wire n_3960;
wire n_3961;
wire n_3962;
wire n_3963;
wire n_3964;
wire n_3965;
wire n_3966;
wire n_3967;
wire n_3968;
wire n_3969;
wire n_3970;
wire n_3971;
wire n_3972;
wire n_3973;
wire n_3974;
wire n_3975;
wire n_3976;
wire n_3977;
wire n_3978;
wire n_3979;
wire n_3980;
wire n_3981;
wire n_3982;
wire n_3983;
wire n_3984;
wire n_3985;
wire n_3986;
wire n_3987;
wire n_3988;
wire n_3989;
wire n_3990;
wire n_3991;
wire n_3992;
wire n_3993;
wire n_3994;
wire n_3995;
wire n_3996;
wire n_3997;
wire n_3998;
wire n_3999;
wire n_4000;
wire n_4001;
wire n_4002;
wire n_4003;
wire n_4004;
wire n_4005;
wire n_4006;
wire n_4007;
wire n_4008;
wire n_4009;
wire n_4010;
wire n_4011;
wire n_4012;
wire n_4013;
wire n_4014;
wire n_4015;
wire n_4016;
wire n_4017;
wire n_4018;
wire n_4019;
wire n_4020;
wire n_4021;
wire n_4022;
wire n_4023;
wire n_4024;
wire n_4025;
wire n_4026;
wire n_4027;
wire n_4028;
wire n_4029;
wire n_4030;
wire n_4031;
wire n_4032;
wire n_4033;
wire n_4034;
wire n_4035;
wire n_4036;
wire n_4037;
wire n_4038;
wire n_4039;
wire n_4040;
wire n_4041;
wire n_4042;
wire n_4043;
wire n_4044;
wire n_4045;
wire n_4046;
wire n_4047;
wire n_4048;
wire n_4049;
wire n_4050;
wire n_4051;
wire n_4052;
wire n_4053;
wire n_4054;
wire n_4055;
wire n_4056;
wire n_4057;
wire n_4058;
wire n_4059;
wire n_4060;
wire n_4061;
wire n_4062;
wire n_4063;
wire n_4064;
wire n_4065;
wire n_4066;
wire n_4067;
wire n_4068;
wire n_4069;
wire n_4070;
wire n_4071;
wire n_4072;
wire n_4073;
wire n_4074;
wire n_4075;
wire n_4076;
wire n_4077;
wire n_4078;
wire n_4079;
wire n_4080;
wire n_4081;
wire n_4082;
wire n_4083;
wire n_4084;
wire n_4085;
wire n_4086;
wire n_4087;
wire n_4088;
wire n_4089;
wire n_4090;
wire n_4091;
wire n_4092;
wire n_4093;
wire n_4094;
wire n_4095;
wire n_4096;
wire n_4097;
wire n_4098;
wire n_4099;
wire n_4100;
wire n_4101;
wire n_4102;
wire n_4103;
wire n_4104;
wire n_4105;
wire n_4106;
wire n_4107;
wire n_4108;
wire n_4109;
wire n_4110;
wire n_4111;
wire n_4112;
wire n_4113;
wire n_4114;
wire n_4115;
wire n_4116;
wire n_4117;
wire n_4118;
wire n_4119;
wire n_4120;
wire n_4121;
wire n_4122;
wire n_4123;
wire n_4124;
wire n_4125;
wire n_4126;
wire n_4127;
wire n_4128;
wire n_4129;
wire n_4130;
wire n_4131;
wire n_4132;
wire n_4133;
wire n_4134;
wire n_4135;
wire n_4136;
wire n_4137;
wire n_4138;
wire n_4139;
wire n_4140;
wire n_4141;
wire n_4142;
wire n_4143;
wire n_4144;
wire n_4145;
wire n_4146;
wire n_4147;
wire n_4148;
wire n_4149;
wire n_4150;
wire n_4151;
wire n_4152;
wire n_4153;
wire n_4154;
wire n_4155;
wire n_4156;
wire n_4157;
wire n_4158;
wire n_4159;
wire n_4160;
wire n_4161;
wire n_4162;
wire n_4163;
wire n_4164;
wire n_4165;
wire n_4166;
wire n_4167;
wire n_4168;
wire n_4169;
wire n_4170;
wire n_4171;
wire n_4172;
wire n_4173;
wire n_4174;
wire n_4175;
wire n_4176;
wire n_4177;
wire n_4178;
wire n_4179;
wire n_4180;
wire n_4181;
wire n_4182;
wire n_4183;
wire n_4184;
wire n_4185;
wire n_4186;
wire n_4187;
wire n_4188;
wire n_4189;
wire n_4190;
wire n_4191;
wire n_4192;
wire n_4193;
wire n_4194;
wire n_4195;
wire n_4196;
wire n_4197;
wire n_4198;
wire n_4199;
wire n_4200;
wire n_4201;
wire n_4202;
wire n_4203;
wire n_4204;
wire n_4205;
wire n_4206;
wire n_4207;
wire n_4208;
wire n_4209;
wire n_4210;
wire n_4211;
wire n_4212;
wire n_4213;
wire n_4214;
wire n_4215;
wire n_4216;
wire n_4217;
wire n_4218;
wire n_4219;
wire n_4220;
wire n_4221;
wire n_4222;
wire n_4223;
wire n_4224;
wire n_4225;
wire n_4226;
wire n_4227;
wire n_4228;
wire n_4229;
wire n_4230;
wire n_4231;
wire n_4232;
wire n_4233;
wire n_4234;
wire n_4235;
wire n_4236;
wire n_4237;
wire n_4238;
wire n_4239;
wire n_4240;
wire n_4241;
wire n_4242;
wire n_4243;
wire n_4244;
wire n_4245;
wire n_4246;
wire n_4247;
wire n_4248;
wire n_4249;
wire n_4250;
wire n_4251;
wire n_4252;
wire n_4253;
wire n_4254;
wire n_4255;
wire n_4256;
wire n_4257;
wire n_4258;
wire n_4259;
wire n_4260;
wire n_4261;
wire n_4262;
wire n_4263;
wire n_4264;
wire n_4265;
wire n_4266;
wire n_4267;
wire n_4268;
wire n_4269;
wire n_4270;
wire n_4271;
wire n_4272;
wire n_4273;
wire n_4274;
wire n_4275;
wire n_4276;
wire n_4277;
wire n_4278;
wire n_4279;
wire n_4280;
wire n_4281;
wire n_4282;
wire n_4283;
wire n_4284;
wire n_4285;
wire n_4286;
wire n_4287;
wire n_4288;
wire n_4289;
wire n_4290;
wire n_4291;
wire n_4292;
wire n_4293;
wire n_4294;
wire n_4295;
wire n_4296;
wire n_4297;
wire n_4298;
wire n_4299;
wire n_4300;
wire n_4301;
wire n_4302;
wire n_4303;
wire n_4304;
wire n_4305;
wire n_4306;
wire n_4307;
wire n_4308;
wire n_4309;
wire n_4310;
wire n_4311;
wire n_4312;
wire n_4313;
wire n_4314;
wire n_4315;
wire n_4316;
wire n_4317;
wire n_4318;
wire n_4319;
wire n_4320;
wire n_4321;
wire n_4322;
wire n_4323;
wire n_4324;
wire n_4325;
wire n_4326;
wire n_4327;
wire n_4328;
wire n_4329;
wire n_4330;
wire n_4331;
wire n_4332;
wire n_4333;
wire n_4334;
wire n_4335;
wire n_4336;
wire n_4337;
wire n_4338;
wire n_4339;
wire n_4340;
wire n_4341;
wire n_4342;
wire n_4343;
wire n_4344;
wire n_4345;
wire n_4346;
wire n_4347;
wire n_4348;
wire n_4349;
wire n_4350;
wire n_4351;
wire n_4352;
wire n_4353;
wire n_4354;
wire n_4355;
wire n_4356;
wire n_4357;
wire n_4358;
wire n_4359;
wire n_4360;
wire n_4361;
wire n_4362;
wire n_4363;
wire n_4364;
wire n_4365;
wire n_4366;
wire n_4367;
wire n_4368;
wire n_4369;
wire n_4370;
wire n_4371;
wire n_4372;
wire n_4373;
wire n_4374;
wire n_4375;
wire n_4376;
wire n_4377;
wire n_4378;
wire n_4379;
wire n_4380;
wire n_4381;
wire n_4382;
wire n_4383;
wire n_4384;
wire n_4385;
wire n_4386;
wire n_4387;
wire n_4388;
wire n_4389;
wire n_4390;
wire n_4391;
wire n_4392;
wire n_4393;
wire n_4394;
wire n_4395;
wire n_4396;
wire n_4397;
wire n_4398;
wire n_4399;
wire n_4400;
wire n_4401;
wire n_4402;
wire n_4403;
wire n_4404;
wire n_4405;
wire n_4406;
wire n_4407;
wire n_4408;
wire n_4409;
wire n_4410;
wire n_4411;
wire n_4412;
wire n_4413;
wire n_4414;
wire n_4415;
wire n_4416;
wire n_4417;
wire n_4418;
wire n_4419;
wire n_4420;
wire n_4421;
wire n_4422;
wire n_4423;
wire n_4424;
wire n_4425;
wire n_4426;
wire n_4427;
wire n_4428;
wire n_4429;
wire n_4430;
wire n_4431;
wire n_4432;
wire n_4433;
wire n_4434;
wire n_4435;
wire n_4436;
wire n_4437;
wire n_4438;
wire n_4439;
wire n_4440;
wire n_4441;
wire n_4442;
wire n_4443;
wire n_4444;
wire n_4445;
wire n_4446;
wire n_4447;
wire n_4448;
wire n_4449;
wire n_4450;
wire n_4451;
wire n_4452;
wire n_4453;
wire n_4454;
wire n_4455;
wire n_4456;
wire n_4457;
wire n_4458;
wire n_4459;
wire n_4460;
wire n_4461;
wire n_4462;
wire n_4463;
wire n_4464;
wire n_4465;
wire n_4466;
wire n_4467;
wire n_4468;
wire n_4469;
wire n_4470;
wire n_4471;
wire n_4472;
wire n_4473;
wire n_4474;
wire n_4475;
wire n_4476;
wire n_4477;
wire n_4478;
wire n_4479;
wire n_4480;
wire n_4481;
wire n_4482;
wire n_4483;
wire n_4484;
wire n_4485;
wire n_4486;
wire n_4487;
wire n_4488;
wire n_4489;
wire n_4490;
wire n_4491;
wire n_4492;
wire n_4493;
wire n_4494;
wire n_4495;
wire n_4496;
wire n_4497;
wire n_4498;
wire n_4499;
wire n_4500;
wire n_4501;
wire n_4502;
wire n_4503;
wire n_4504;
wire n_4505;
wire n_4506;
wire n_4507;
wire n_4508;
wire n_4509;
wire n_4510;
wire n_4511;
wire n_4512;
wire n_4513;
wire n_4514;
wire n_4515;
wire n_4516;
wire n_4517;
wire n_4518;
wire n_4519;
wire n_4520;
wire n_4521;
wire n_4522;
wire n_4523;
wire n_4524;
wire n_4525;
wire n_4526;
wire n_4527;
wire n_4528;
wire n_4529;
wire n_4530;
wire n_4531;
wire n_4532;
wire n_4533;
wire n_4534;
wire n_4535;
wire n_4536;
wire n_4537;
wire n_4538;
wire n_4539;
wire n_4540;
wire n_4541;
wire n_4542;
wire n_4543;
wire n_4544;
wire n_4545;
wire n_4546;
wire n_4547;
wire n_4548;
wire n_4549;
wire n_4550;
wire n_4551;
wire n_4552;
wire n_4553;
wire n_4554;
wire n_4555;
wire n_4556;
wire n_4557;
wire n_4558;
wire n_4559;
wire n_4560;
wire n_4561;
wire n_4562;
wire n_4563;
wire n_4564;
wire n_4565;
wire n_4566;
wire n_4567;
wire n_4568;
wire n_4569;
wire n_4570;
wire n_4571;
wire n_4572;
wire n_4573;
wire n_4574;
wire n_4575;
wire n_4576;
wire n_4577;
wire n_4578;
wire n_4579;
wire n_4580;
wire n_4581;
wire n_4582;
wire n_4583;
wire n_4584;
wire n_4585;
wire n_4586;
wire n_4587;
wire n_4588;
wire n_4589;
wire n_4590;
wire n_4591;
wire n_4592;
wire n_4593;
wire n_4594;
wire n_4595;
wire n_4596;
wire n_4597;
wire n_4598;
wire n_4599;
wire n_4600;
wire n_4601;
wire n_4602;
wire n_4603;
wire n_4604;
wire n_4605;
wire n_4606;
wire n_4607;
wire n_4608;
wire n_4609;
wire n_4610;
wire n_4611;
wire n_4612;
wire n_4613;
wire n_4614;
wire n_4615;
wire n_4616;
wire n_4617;
wire n_4618;
wire n_4619;
wire n_4620;
wire n_4621;
wire n_4622;
wire n_4623;
wire n_4624;
wire n_4625;
wire n_4626;
wire n_4627;
wire n_4628;
wire n_4629;
wire n_4630;
wire n_4631;
wire n_4632;
wire n_4633;
wire n_4634;
wire n_4635;
wire n_4636;
wire n_4637;
wire n_4638;
wire n_4639;
wire n_4640;
wire n_4641;
wire n_4642;
wire n_4643;
wire n_4644;
wire n_4645;
wire n_4646;
wire n_4647;
wire n_4648;
wire n_4649;
wire n_4650;
wire n_4651;
wire n_4652;
wire n_4653;
wire n_4654;
wire n_4655;
wire n_4656;
wire n_4657;
wire n_4658;
wire n_4659;
wire n_4660;
wire n_4661;
wire n_4662;
wire n_4663;
wire n_4664;
wire n_4665;
wire n_4666;
wire n_4667;
wire n_4668;
wire n_4669;
wire n_4670;
wire n_4671;
wire n_4672;
wire n_4673;
wire n_4674;
wire n_4675;
wire n_4676;
wire n_4677;
wire n_4678;
wire n_4679;
wire n_4680;
wire n_4681;
wire n_4682;
wire n_4683;
wire n_4684;
wire n_4685;
wire n_4686;
wire n_4687;
wire n_4688;
wire n_4689;
wire n_4690;
wire n_4691;
wire n_4692;
wire n_4693;
wire n_4694;
wire n_4695;
wire n_4696;
wire n_4697;
wire n_4698;
wire n_4699;
wire n_4700;
wire n_4701;
wire n_4702;
wire n_4703;
wire n_4704;
wire n_4705;
wire n_4706;
wire n_4707;
wire n_4708;
wire n_4709;
wire n_4710;
wire n_4711;
wire n_4712;
wire n_4713;
wire n_4714;
wire n_4715;
wire n_4716;
wire n_4717;
wire n_4718;
wire n_4719;
wire n_4720;
wire n_4721;
wire n_4722;
wire n_4723;
wire n_4724;
wire n_4725;
wire n_4726;
wire n_4727;
wire n_4728;
wire n_4729;
wire n_4730;
wire n_4731;
wire n_4732;
wire n_4733;
wire n_4734;
wire n_4735;
wire n_4736;
wire n_4737;
wire n_4738;
wire n_4739;
wire n_4740;
wire n_4741;
wire n_4742;
wire n_4743;
wire n_4744;
wire n_4745;
wire n_4746;
wire n_4747;
wire n_4748;
wire n_4749;
wire n_4750;
wire n_4751;
wire n_4752;
wire n_4753;
wire n_4754;
wire n_4755;
wire n_4756;
wire n_4757;
wire n_4758;
wire n_4759;
wire n_4760;
wire n_4761;
wire n_4762;
wire n_4763;
wire n_4764;
wire n_4765;
wire n_4766;
wire n_4767;
wire n_4768;
wire n_4769;
wire n_4770;
wire n_4771;
wire n_4772;
wire n_4773;
wire n_4774;
wire n_4775;
wire n_4776;
wire n_4777;
wire n_4778;
wire n_4779;
wire n_4780;
wire n_4781;
wire n_4782;
wire n_4783;
wire n_4784;
wire n_4785;
wire n_4786;
wire n_4787;
wire n_4788;
wire n_4789;
wire n_4790;
wire n_4791;
wire n_4792;
wire n_4793;
wire n_4794;
wire n_4795;
wire n_4796;
wire n_4797;
wire n_4798;
wire n_4799;
wire n_4800;
wire n_4801;
wire n_4802;
wire n_4803;
wire n_4804;
wire n_4805;
wire n_4806;
wire n_4807;
wire n_4808;
wire n_4809;
wire n_4810;
wire n_4811;
wire n_4812;
wire n_4813;
wire n_4814;
wire n_4815;
wire n_4816;
wire n_4817;
wire n_4818;
wire n_4819;
wire n_4820;
wire n_4821;
wire n_4822;
wire n_4823;
wire n_4824;
wire n_4825;
wire n_4826;
wire n_4827;
wire n_4828;
wire n_4829;
wire n_4830;
wire n_4831;
wire n_4832;
wire n_4833;
wire n_4834;
wire n_4835;
wire n_4836;
wire n_4837;
wire n_4838;
wire n_4839;
wire n_4840;
wire n_4841;
wire n_4842;
wire n_4843;
wire n_4844;
wire n_4845;
wire n_4846;
wire n_4847;
wire n_4848;
wire n_4849;
wire n_4850;
wire n_4851;
wire n_4852;
wire n_4853;
wire n_4854;
wire n_4855;
wire n_4856;
wire n_4857;
wire n_4858;
wire n_4859;
wire n_4860;
wire n_4861;
wire n_4862;
wire n_4863;
wire n_4864;
wire n_4865;
wire n_4866;
wire n_4867;
wire n_4868;
wire n_4869;
wire n_4870;
wire n_4871;
wire n_4872;
wire n_4873;
wire n_4874;
wire n_4875;
wire n_4876;
wire n_4877;
wire n_4878;
wire n_4879;
wire n_4880;
wire n_4881;
wire n_4882;
wire n_4883;
wire n_4884;
wire n_4885;
wire n_4886;
wire n_4887;
wire n_4888;
wire n_4889;
wire n_4890;
wire n_4891;
wire n_4892;
wire n_4893;
wire n_4894;
wire n_4895;
wire n_4896;
wire n_4897;
wire n_4898;
wire n_4899;
wire n_4900;
wire n_4901;
wire n_4902;
wire n_4903;
wire n_4904;
wire n_4905;
wire n_4906;
wire n_4907;
wire n_4908;
wire n_4909;
wire n_4910;
wire n_4911;
wire n_4912;
wire n_4913;
wire n_4914;
wire n_4915;
wire n_4916;
wire n_4917;
wire n_4918;
wire n_4919;
wire n_4920;
wire n_4921;
wire n_4922;
wire n_4923;
wire n_4924;
wire n_4925;
wire n_4926;
wire n_4927;
wire n_4928;
wire n_4929;
wire n_4930;
wire n_4931;
wire n_4932;
wire n_4933;
wire n_4934;
wire n_4935;
wire n_4936;
wire n_4937;
wire n_4938;
wire n_4939;
wire n_4940;
wire n_4941;
wire n_4942;
wire n_4943;
wire n_4944;
wire n_4945;
wire n_4946;
wire n_4947;
wire n_4948;
wire n_4949;
wire n_4950;
wire n_4951;
wire n_4952;
wire n_4953;
wire n_4954;
wire n_4955;
wire n_4956;
wire n_4957;
wire n_4958;
wire n_4959;
wire n_4960;
wire n_4961;
wire n_4962;
wire n_4963;
wire n_4964;
wire n_4965;
wire n_4966;
wire n_4967;
wire n_4968;
wire n_4969;
wire n_4970;
wire n_4971;
wire n_4972;
wire n_4973;
wire n_4974;
wire n_4975;
wire n_4976;
wire n_4977;
wire n_4978;
wire n_4979;
wire n_4980;
wire n_4981;
wire n_4982;
wire n_4983;
wire n_4984;
wire n_4985;
wire n_4986;
wire n_4987;
wire n_4988;
wire n_4989;
wire n_4990;
wire n_4991;
wire n_4992;
wire n_4993;
wire n_4994;
wire n_4995;
wire n_4996;
wire n_4997;
wire n_4998;
wire n_4999;
wire n_5000;
wire n_5001;
wire n_5002;
wire n_5003;
wire n_5004;
wire n_5005;
wire n_5006;
wire n_5007;
wire n_5008;
wire n_5009;
wire n_5010;
wire n_5011;
wire n_5012;
wire n_5013;
wire n_5014;
wire n_5015;
wire n_5016;
wire n_5017;
wire n_5018;
wire n_5019;
wire n_5020;
wire n_5021;
wire n_5022;
wire n_5023;
wire n_5024;
wire n_5025;
wire n_5026;
wire n_5027;
wire n_5028;
wire n_5029;
wire n_5030;
wire n_5031;
wire n_5032;
wire n_5033;
wire n_5034;
wire n_5035;
wire n_5036;
wire n_5037;
wire n_5038;
wire n_5039;
wire n_5040;
wire n_5041;
wire n_5042;
wire n_5043;
wire n_5044;
wire n_5045;
wire n_5046;
wire n_5047;
wire n_5048;
wire n_5049;
wire n_5050;
wire n_5051;
wire n_5052;
wire n_5053;
wire n_5054;
wire n_5055;
wire n_5056;
wire n_5057;
wire n_5058;
wire n_5059;
wire n_5060;
wire n_5061;
wire n_5062;
wire n_5063;
wire n_5064;
wire n_5065;
wire n_5066;
wire n_5067;
wire n_5068;
wire n_5069;
wire n_5070;
wire n_5071;
wire n_5072;
wire n_5073;
wire n_5074;
wire n_5075;
wire n_5076;
wire n_5077;
wire n_5078;
wire n_5079;
wire n_5080;
wire n_5081;
wire n_5082;
wire n_5083;
wire n_5084;
wire n_5085;
wire n_5086;
wire n_5087;
wire n_5088;
wire n_5089;
wire n_5090;
wire n_5091;
wire n_5092;
wire n_5093;
wire n_5094;
wire n_5095;
wire n_5096;
wire n_5097;
wire n_5098;
wire n_5099;
wire n_5100;
wire n_5101;
wire n_5102;
wire n_5103;
wire n_5104;
wire n_5105;
wire n_5106;
wire n_5107;
wire n_5108;
wire n_5109;
wire n_5110;
wire n_5111;
wire n_5112;
wire n_5113;
wire n_5114;
wire n_5115;
wire n_5116;
wire n_5117;
wire n_5118;
wire n_5119;
wire n_5120;
wire n_5121;
wire n_5122;
wire n_5123;
wire n_5124;
wire n_5125;
wire n_5126;
wire n_5127;
wire n_5128;
wire n_5129;
wire n_5130;
wire n_5131;
wire n_5132;
wire n_5133;
wire n_5134;
wire n_5135;
wire n_5136;
wire n_5137;
wire n_5138;
wire n_5139;
wire n_5140;
wire n_5141;
wire n_5142;
wire n_5143;
wire n_5144;
wire n_5145;
wire n_5146;
wire n_5147;
wire n_5148;
wire n_5149;
wire n_5150;
wire n_5151;
wire n_5152;
wire n_5153;
wire n_5154;
wire n_5155;
wire n_5156;
wire n_5157;
wire n_5158;
wire n_5159;
wire n_5160;
wire n_5161;
wire n_5162;
wire n_5163;
wire n_5164;
wire n_5165;
wire n_5166;
wire n_5167;
wire n_5168;
wire n_5169;
wire n_5170;
wire n_5171;
wire n_5172;
wire n_5173;
wire n_5174;
wire n_5175;
wire n_5176;
wire n_5177;
wire n_5178;
wire n_5179;
wire n_5180;
wire n_5181;
wire n_5182;
wire n_5183;
wire n_5184;
wire n_5185;
wire n_5186;
wire n_5187;
wire n_5188;
wire n_5189;
wire n_5190;
wire n_5191;
wire n_5192;
wire n_5193;
wire n_5194;
wire n_5195;
wire n_5196;
wire n_5197;
wire n_5198;
wire n_5199;
wire n_5200;
wire n_5201;
wire n_5202;
wire n_5203;
wire n_5204;
wire n_5205;
wire n_5206;
wire n_5207;
wire n_5208;
wire n_5209;
wire n_5210;
wire n_5211;
wire n_5212;
wire n_5213;
wire n_5214;
wire n_5215;
wire n_5216;
wire n_5217;
wire n_5218;
wire n_5219;
wire n_5220;
wire n_5221;
wire n_5222;
wire n_5223;
wire n_5224;
wire n_5225;
wire n_5226;
wire n_5227;
wire n_5228;
wire n_5229;
wire n_5230;
wire n_5231;
wire n_5232;
wire n_5233;
wire n_5234;
wire n_5235;
wire n_5236;
wire n_5237;
wire n_5238;
wire n_5239;
wire n_5240;
wire n_5241;
wire n_5242;
wire n_5243;
wire n_5244;
wire n_5245;
wire n_5246;
wire n_5247;
wire n_5248;
wire n_5249;
wire n_5250;
wire n_5251;
wire n_5252;
wire n_5253;
wire n_5254;
wire n_5255;
wire n_5256;
wire n_5257;
wire n_5258;
wire n_5259;
wire n_5260;
wire n_5261;
wire n_5262;
wire n_5263;
wire n_5264;
wire n_5265;
wire n_5266;
wire n_5267;
wire n_5268;
wire n_5269;
wire n_5270;
wire n_5271;
wire n_5272;
wire n_5273;
wire n_5274;
wire n_5275;
wire n_5276;
wire n_5277;
wire n_5278;
wire n_5279;
wire n_5280;
wire n_5281;
wire n_5282;
wire n_5283;
wire n_5284;
wire n_5285;
wire n_5286;
wire n_5287;
wire n_5288;
wire n_5289;
wire n_5290;
wire n_5291;
wire n_5292;
wire n_5293;
wire n_5294;
wire n_5295;
wire n_5296;
wire n_5297;
wire n_5298;
wire n_5299;
wire n_5300;
wire n_5301;
wire n_5302;
wire n_5303;
wire n_5304;
wire n_5305;
wire n_5306;
wire n_5307;
wire n_5308;
wire n_5309;
wire n_5310;
wire n_5311;
wire n_5312;
wire n_5313;
wire n_5314;
wire n_5315;
wire n_5316;
wire n_5317;
wire n_5318;
wire n_5319;
wire n_5320;
wire n_5321;
wire n_5322;
wire n_5323;
wire n_5324;
wire n_5325;
wire n_5326;
wire n_5327;
wire n_5328;
wire n_5329;
wire n_5330;
wire n_5331;
wire n_5332;
wire n_5333;
wire n_5334;
wire n_5335;
wire n_5336;
wire n_5337;
wire n_5338;
wire n_5339;
wire n_5340;
wire n_5341;
wire n_5342;
wire n_5343;
wire n_5344;
wire n_5345;
wire n_5346;
wire n_5347;
wire n_5348;
wire n_5349;
wire n_5350;
wire n_5351;
wire n_5352;
wire n_5353;
wire n_5354;
wire n_5355;
wire n_5356;
wire n_5357;
wire n_5358;
wire n_5359;
wire n_5360;
wire n_5361;
wire n_5362;
wire n_5363;
wire n_5364;
wire n_5365;
wire n_5366;
wire n_5367;
wire n_5368;
wire n_5369;
wire n_5370;
wire n_5371;
wire n_5372;
wire n_5373;
wire n_5374;
wire n_5375;
wire n_5376;
wire n_5377;
wire n_5378;
wire n_5379;
wire n_5380;
wire n_5381;
wire n_5382;
wire n_5383;
wire n_5384;
wire n_5385;
wire n_5386;
wire n_5387;
wire n_5388;
wire n_5389;
wire n_5390;
wire n_5391;
wire n_5392;
wire n_5393;
wire n_5394;
wire n_5395;
wire n_5396;
wire n_5397;
wire n_5398;
wire n_5399;
wire n_5400;
wire n_5401;
wire n_5402;
wire n_5403;
wire n_5404;
wire n_5405;
wire n_5406;
wire n_5407;
wire n_5408;
wire n_5409;
wire n_5410;
wire n_5411;
wire n_5412;
wire n_5413;
wire n_5414;
wire n_5415;
wire n_5416;
wire n_5417;
wire n_5418;
wire n_5419;
wire n_5420;
wire n_5421;
wire n_5422;
wire n_5423;
wire n_5424;
wire n_5425;
wire n_5426;
wire n_5427;
wire n_5428;
wire n_5429;
wire n_5430;
wire n_5431;
wire n_5432;
wire n_5433;
wire n_5434;
wire n_5435;
wire n_5436;
wire n_5437;
wire n_5438;
wire n_5439;
wire n_5440;
wire n_5441;
wire n_5442;
wire n_5443;
wire n_5444;
wire n_5445;
wire n_5446;
wire n_5447;
wire n_5448;
wire n_5449;
wire n_5450;
wire n_5451;
wire n_5452;
wire n_5453;
wire n_5454;
wire n_5455;
wire n_5456;
wire n_5457;
wire n_5458;
wire n_5459;
wire n_5460;
wire n_5461;
wire n_5462;
wire n_5463;
wire n_5464;
wire n_5465;
wire n_5466;
wire n_5467;
wire n_5468;
wire n_5469;
wire n_5470;
wire n_5471;
wire n_5472;
wire n_5473;
wire n_5474;
wire n_5475;
wire n_5476;
wire n_5477;
wire n_5478;
wire n_5479;
wire n_5480;
wire n_5481;
wire n_5482;
wire n_5483;
wire n_5484;
wire n_5485;
wire n_5486;
wire n_5487;
wire n_5488;
wire n_5489;
wire n_5490;
wire n_5491;
wire n_5492;
wire n_5493;
wire n_5494;
wire n_5495;
wire n_5496;
wire n_5497;
wire n_5498;
wire n_5499;
wire n_5500;
wire n_5501;
wire n_5502;
wire n_5503;
wire n_5504;
wire n_5505;
wire n_5506;
wire n_5507;
wire n_5508;
wire n_5509;
wire n_5510;
wire n_5511;
wire n_5512;
wire n_5513;
wire n_5514;
wire n_5515;
wire n_5516;
wire n_5517;
wire n_5518;
wire n_5519;
wire n_5520;
wire n_5521;
wire n_5522;
wire n_5523;
wire n_5524;
wire n_5525;
wire n_5526;
wire n_5527;
wire n_5528;
wire n_5529;
wire n_5530;
wire n_5531;
wire n_5532;
wire n_5533;
wire n_5534;
wire n_5535;
wire n_5536;
wire n_5537;
wire n_5538;
wire n_5539;
wire n_5540;
wire n_5541;
wire n_5542;
wire n_5543;
wire n_5544;
wire n_5545;
wire n_5546;
wire n_5547;
wire n_5548;
wire n_5549;
wire n_5550;
wire n_5551;
wire n_5552;
wire n_5553;
wire n_5554;
wire n_5555;
wire n_5556;
wire n_5557;
wire n_5558;
wire n_5559;
wire n_5560;
wire n_5561;
wire n_5562;
wire n_5563;
wire n_5564;
wire n_5565;
wire n_5566;
wire n_5567;
wire n_5568;
wire n_5569;
wire n_5570;
wire n_5571;
wire n_5572;
wire n_5573;
wire n_5574;
wire n_5575;
wire n_5576;
wire n_5577;
wire n_5578;
wire n_5579;
wire n_5580;
wire n_5581;
wire n_5582;
wire n_5583;
wire n_5584;
wire n_5585;
wire n_5586;
wire n_5587;
wire n_5588;
wire n_5589;
wire n_5590;
wire n_5591;
wire n_5592;
wire n_5593;
wire n_5594;
wire n_5595;
wire n_5596;
wire n_5597;
wire n_5598;
wire n_5599;
wire n_5600;
wire n_5601;
wire n_5602;
wire n_5603;
wire n_5604;
wire n_5605;
wire n_5606;
wire n_5607;
wire n_5608;
wire n_5609;
wire n_5610;
wire n_5611;
wire n_5612;
wire n_5613;
wire n_5614;
wire n_5615;
wire n_5616;
wire n_5617;
wire n_5618;
wire n_5619;
wire n_5620;
wire n_5621;
wire n_5622;
wire n_5623;
wire n_5624;
wire n_5625;
wire n_5626;
wire n_5627;
wire n_5628;
wire n_5629;
wire n_5630;
wire n_5631;
wire n_5632;
wire n_5633;
wire n_5634;
wire n_5635;
wire n_5636;
wire n_5637;
wire n_5638;
wire n_5639;
wire n_5640;
wire n_5641;
wire n_5642;
wire n_5643;
wire n_5644;
wire n_5645;
wire n_5646;
wire n_5647;
wire n_5648;
wire n_5649;
wire n_5650;
wire n_5651;
wire n_5652;
wire n_5653;
wire n_5654;
wire n_5655;
wire n_5656;
wire n_5657;
wire n_5658;
wire n_5659;
wire n_5660;
wire n_5661;
wire n_5662;
wire n_5663;
wire n_5664;
wire n_5665;
wire n_5666;
wire n_5667;
wire n_5668;
wire n_5669;
wire n_5670;
wire n_5671;
wire n_5672;
wire n_5673;
wire n_5674;
wire n_5675;
wire n_5676;
wire n_5677;
wire n_5678;
wire n_5679;
wire n_5680;
wire n_5681;
wire n_5682;
wire n_5683;
wire n_5684;
wire n_5685;
wire n_5686;
wire n_5687;
wire n_5688;
wire n_5689;
wire n_5690;
wire n_5691;
wire n_5692;
wire n_5693;
wire n_5694;
wire n_5695;
wire n_5696;
wire n_5697;
wire n_5698;
wire n_5699;
wire n_5700;
wire n_5701;
wire n_5702;
wire n_5703;
wire n_5704;
wire n_5705;
wire n_5706;
wire n_5707;
wire n_5708;
wire n_5709;
wire n_5710;
wire n_5711;
wire n_5712;
wire n_5713;
wire n_5714;
wire n_5715;
wire n_5716;
wire n_5717;
wire n_5718;
wire n_5719;
wire n_5720;
wire n_5721;
wire n_5722;
wire n_5723;
wire n_5724;
wire n_5725;
wire n_5726;
wire n_5727;
wire n_5728;
wire n_5729;
wire n_5730;
wire n_5731;
wire n_5732;
wire n_5733;
wire n_5734;
wire n_5735;
wire n_5736;
wire n_5737;
wire n_5738;
wire n_5739;
wire n_5740;
wire n_5741;
wire n_5742;
wire n_5743;
wire n_5744;
wire n_5745;
wire n_5746;
wire n_5747;
wire n_5748;
wire n_5749;
wire n_5750;
wire n_5751;
wire n_5752;
wire n_5753;
wire n_5754;
wire n_5755;
wire n_5756;
wire n_5757;
wire n_5758;
wire n_5759;
wire n_5760;
wire n_5761;
wire n_5762;
wire n_5763;
wire n_5764;
wire n_5765;
wire n_5766;
wire n_5767;
wire n_5768;
wire n_5769;
wire n_5770;
wire n_5771;
wire n_5772;
wire n_5773;
wire n_5774;
wire n_5775;
wire n_5776;
wire n_5777;
wire n_5778;
wire n_5779;
wire n_5780;
wire n_5781;
wire n_5782;
wire n_5783;
wire n_5784;
wire n_5785;
wire n_5786;
wire n_5787;
wire n_5788;
wire n_5789;
wire n_5790;
wire n_5791;
wire n_5792;
wire n_5793;
wire n_5794;
wire n_5795;
wire n_5796;
wire n_5797;
wire n_5798;
wire n_5799;
wire n_5800;
wire n_5801;
wire n_5802;
wire n_5803;
wire n_5804;
wire n_5805;
wire n_5806;
wire n_5807;
wire n_5808;
wire n_5809;
wire n_5810;
wire n_5811;
wire n_5812;
wire n_5813;
wire n_5814;
wire n_5815;
wire n_5816;
wire n_5817;
wire n_5818;
wire n_5819;
wire n_5820;
wire n_5821;
wire n_5822;
wire n_5823;
wire n_5824;
wire n_5825;
wire n_5826;
wire n_5827;
wire n_5828;
wire n_5829;
wire n_5830;
wire n_5831;
wire n_5832;
wire n_5833;
wire n_5834;
wire n_5835;
wire n_5836;
wire n_5837;
wire n_5838;
wire n_5839;
wire n_5840;
wire n_5841;
wire n_5842;
wire n_5843;
wire n_5844;
wire n_5845;
wire n_5846;
wire n_5847;
wire n_5848;
wire n_5849;
wire n_5850;
wire n_5851;
wire n_5852;
wire n_5853;
wire n_5854;
wire n_5855;
wire n_5856;
wire n_5857;
wire n_5858;
wire n_5859;
wire n_5860;
wire n_5861;
wire n_5862;
wire n_5863;
wire n_5864;
wire n_5865;
wire n_5866;
wire n_5867;
wire n_5868;
wire n_5869;
wire n_5870;
wire n_5871;
wire n_5872;
wire n_5873;
wire n_5874;
wire n_5875;
wire n_5876;
wire n_5877;
wire n_5878;
wire n_5879;
wire n_5880;
wire n_5881;
wire n_5882;
wire n_5883;
wire n_5884;
wire n_5885;
wire n_5886;
wire n_5887;
wire n_5888;
wire n_5889;
wire n_5890;
wire n_5891;
wire n_5892;
wire n_5893;
wire n_5894;
wire n_5895;
wire n_5896;
wire n_5897;
wire n_5898;
wire n_5899;
wire n_5900;
wire n_5901;
wire n_5902;
wire n_5903;
wire n_5904;
wire n_5905;
wire n_5906;
wire n_5907;
wire n_5908;
wire n_5909;
wire n_5910;
wire n_5911;
wire n_5912;
wire n_5913;
wire n_5914;
wire n_5915;
wire n_5916;
wire n_5917;
wire n_5918;
wire n_5919;
wire n_5920;
wire n_5921;
wire n_5922;
wire n_5923;
wire n_5924;
wire n_5925;
wire n_5926;
wire n_5927;
wire n_5928;
wire n_5929;
wire n_5930;
wire n_5931;
wire n_5932;
wire n_5933;
wire n_5934;
wire n_5935;
wire n_5936;
wire n_5937;
wire n_5938;
wire n_5939;
wire n_5940;
wire n_5941;
wire n_5942;
wire n_5943;
wire n_5944;
wire n_5945;
wire n_5946;
wire n_5947;
wire n_5948;
wire n_5949;
wire n_5950;
wire n_5951;
wire n_5952;
wire n_5953;
wire n_5954;
wire n_5955;
wire n_5956;
wire n_5957;
wire n_5958;
wire n_5959;
wire n_5960;
wire n_5961;
wire n_5962;
wire n_5963;
wire n_5964;
wire n_5965;
wire n_5966;
wire n_5967;
wire n_5968;
wire n_5969;
wire n_5970;
wire n_5971;
wire n_5972;
wire n_5973;
wire n_5974;
wire n_5975;
wire n_5976;
wire n_5977;
wire n_5978;
wire n_5979;
wire n_5980;
wire n_5981;
wire n_5982;
wire n_5983;
wire n_5984;
wire n_5985;
wire n_5986;
wire n_5987;
wire n_5988;
wire n_5989;
wire n_5990;
wire n_5991;
wire n_5992;
wire n_5993;
wire n_5994;
wire n_5995;
wire n_5996;
wire n_5997;
wire n_5998;
wire n_5999;
wire n_6000;
wire n_6001;
wire n_6002;
wire n_6003;
wire n_6004;
wire n_6005;
wire n_6006;
wire n_6007;
wire n_6008;
wire n_6009;
wire n_6010;
wire n_6011;
wire n_6012;
wire n_6013;
wire n_6014;
wire n_6015;
wire n_6016;
wire n_6017;
wire n_6018;
wire n_6019;
wire n_6020;
wire n_6021;
wire n_6022;
wire n_6023;
wire n_6024;
wire n_6025;
wire n_6026;
wire n_6027;
wire n_6028;
wire n_6029;
wire n_6030;
wire n_6031;
wire n_6032;
wire n_6033;
wire n_6034;
wire n_6035;
wire n_6036;
wire n_6037;
wire n_6038;
wire n_6039;
wire n_6040;
wire n_6041;
wire n_6042;
wire n_6043;
wire n_6044;
wire n_6045;
wire n_6046;
wire n_6047;
wire n_6048;
wire n_6049;
wire n_6050;
wire n_6051;
wire n_6052;
wire n_6053;
wire n_6054;
wire n_6055;
wire n_6056;
wire n_6057;
wire n_6058;
wire n_6059;
wire n_6060;
wire n_6061;
wire n_6062;
wire n_6063;
wire n_6064;
wire n_6065;
wire n_6066;
wire n_6067;
wire n_6068;
wire n_6069;
wire n_6070;
wire n_6071;
wire n_6072;
wire n_6073;
wire n_6074;
wire n_6075;
wire n_6076;
wire n_6077;
wire n_6078;
wire n_6079;
wire n_6080;
wire n_6081;
wire n_6082;
wire n_6083;
wire n_6084;
wire n_6085;
wire n_6086;
wire n_6087;
wire n_6088;
wire n_6089;
wire n_6090;
wire n_6091;
wire n_6092;
wire n_6093;
wire n_6094;
wire n_6095;
wire n_6096;
wire n_6097;
wire n_6098;
wire n_6099;
wire n_6100;
wire n_6101;
wire n_6102;
wire n_6103;
wire n_6104;
wire n_6105;
wire n_6106;
wire n_6107;
wire n_6108;
wire n_6109;
wire n_6110;
wire n_6111;
wire n_6112;
wire n_6113;
wire n_6114;
wire n_6115;
wire n_6116;
wire n_6117;
wire n_6118;
wire n_6119;
wire n_6120;
wire n_6121;
wire n_6122;
wire n_6123;
wire n_6124;
wire n_6125;
wire n_6126;
wire n_6127;
wire n_6128;
wire n_6129;
wire n_6130;
wire n_6131;
wire n_6132;
wire n_6133;
wire n_6134;
wire n_6135;
wire n_6136;
wire n_6137;
wire n_6138;
wire n_6139;
wire n_6140;
wire n_6141;
wire n_6142;
wire n_6143;
wire n_6144;
wire n_6145;
wire n_6146;
wire n_6147;
wire n_6148;
wire n_6149;
wire n_6150;
wire n_6151;
wire n_6152;
wire n_6153;
wire n_6154;
wire n_6155;
wire n_6156;
wire n_6157;
wire n_6158;
wire n_6159;
wire n_6160;
wire n_6161;
wire n_6162;
wire n_6163;
wire n_6164;
wire n_6165;
wire n_6166;
wire n_6167;
wire n_6168;
wire n_6169;
wire n_6170;
wire n_6171;
wire n_6172;
wire n_6173;
wire n_6174;
wire n_6175;
wire n_6176;
wire n_6177;
wire n_6178;
wire n_6179;
wire n_6180;
wire n_6181;
wire n_6182;
wire n_6183;
wire n_6184;
wire n_6185;
wire n_6186;
wire n_6187;
wire n_6188;
wire n_6189;
wire n_6190;
wire n_6191;
wire n_6192;
wire n_6193;
wire n_6194;
wire n_6195;
wire n_6196;
wire n_6197;
wire n_6198;
wire n_6199;
wire n_6200;
wire n_6201;
wire n_6202;
wire n_6203;
wire n_6204;
wire n_6205;
wire n_6206;
wire n_6207;
wire n_6208;
wire n_6209;
wire n_6210;
wire n_6211;
wire n_6212;
wire n_6213;
wire n_6214;
wire n_6215;
wire n_6216;
wire n_6217;
wire n_6218;
wire n_6219;
wire n_6220;
wire n_6221;
wire n_6222;
wire n_6223;
wire n_6224;
wire n_6225;
wire n_6226;
wire n_6227;
wire n_6228;
wire n_6229;
wire n_6230;
wire n_6231;
wire n_6232;
wire n_6233;
wire n_6234;
wire n_6235;
wire n_6236;
wire n_6237;
wire n_6238;
wire n_6239;
wire n_6240;
wire n_6241;
wire n_6242;
wire n_6243;
wire n_6244;
wire n_6245;
wire n_6246;
wire n_6247;
wire n_6248;
wire n_6249;
wire n_6250;
wire n_6251;
wire n_6252;
wire n_6253;
wire n_6254;
wire n_6255;
wire n_6256;
wire n_6257;
wire n_6258;
wire n_6259;
wire n_6260;
wire n_6261;
wire n_6262;
wire n_6263;
wire n_6264;
wire n_6265;
wire n_6266;
wire n_6267;
wire n_6268;
wire n_6269;
wire n_6270;
wire n_6271;
wire n_6272;
wire n_6273;
wire n_6274;
wire n_6275;
wire n_6276;
wire n_6277;
wire n_6278;
wire n_6279;
wire n_6280;
wire n_6281;
wire n_6282;
wire n_6283;
wire n_6284;
wire n_6285;
wire n_6286;
wire n_6287;
wire n_6288;
wire n_6289;
wire n_6290;
wire n_6291;
wire n_6292;
wire n_6293;
wire n_6294;
wire n_6295;
wire n_6296;
wire n_6297;
wire n_6298;
wire n_6299;
wire n_6300;
wire n_6301;
wire n_6302;
wire n_6303;
wire n_6304;
wire n_6305;
wire n_6306;
wire n_6307;
wire n_6308;
wire n_6309;
wire n_6310;
wire n_6311;
wire n_6312;
wire n_6313;
wire n_6314;
wire n_6315;
wire n_6316;
wire n_6317;
wire n_6318;
wire n_6319;
wire n_6320;
wire n_6321;
wire n_6322;
wire n_6323;
wire n_6324;
wire n_6325;
wire n_6326;
wire n_6327;
wire n_6328;
wire n_6329;
wire n_6330;
wire n_6331;
wire n_6332;
wire n_6333;
wire n_6334;
wire n_6335;
wire n_6336;
wire n_6337;
wire n_6338;
wire n_6339;
wire n_6340;
wire n_6341;
wire n_6342;
wire n_6343;
wire n_6344;
wire n_6345;
wire n_6346;
wire n_6347;
wire n_6348;
wire n_6349;
wire n_6350;
wire n_6351;
wire n_6352;
wire n_6353;
wire n_6354;
wire n_6355;
wire n_6356;
wire n_6357;
wire n_6358;
wire n_6359;
wire n_6360;
wire n_6361;
wire n_6362;
wire n_6363;
wire n_6364;
wire n_6365;
wire n_6366;
wire n_6367;
wire n_6368;
wire n_6369;
wire n_6370;
wire n_6371;
wire n_6372;
wire n_6373;
wire n_6374;
wire n_6375;
wire n_6376;
wire n_6377;
wire n_6378;
wire n_6379;
wire n_6380;
wire n_6381;
wire n_6382;
wire n_6383;
wire n_6384;
wire n_6385;
wire n_6386;
wire n_6387;
wire n_6388;
wire n_6389;
wire n_6390;
wire n_6391;
wire n_6392;
wire n_6393;
wire n_6394;
wire n_6395;
wire n_6396;
wire n_6397;
wire n_6398;
wire n_6399;
wire n_6400;
wire n_6401;
wire n_6402;
wire n_6403;
wire n_6404;
wire n_6405;
wire n_6406;
wire n_6407;
wire n_6408;
wire n_6409;
wire n_6410;
wire n_6411;
wire n_6412;
wire n_6413;
wire n_6414;
wire n_6415;
wire n_6416;
wire n_6417;
wire n_6418;
wire n_6419;
wire n_6420;
wire n_6421;
wire n_6422;
wire n_6423;
wire n_6424;
wire n_6425;
wire n_6426;
wire n_6427;
wire n_6428;
wire n_6429;
wire n_6430;
wire n_6431;
wire n_6432;
wire n_6433;
wire n_6434;
wire n_6435;
wire n_6436;
wire n_6437;
wire n_6438;
wire n_6439;
wire n_6440;
wire n_6441;
wire n_6442;
wire n_6443;
wire n_6444;
wire n_6445;
wire n_6446;
wire n_6447;
wire n_6448;
wire n_6449;
wire n_6450;
wire n_6451;
wire n_6452;
wire n_6453;
wire n_6454;
wire n_6455;
wire n_6456;
wire n_6457;
wire n_6458;
wire n_6459;
wire n_6460;
wire n_6461;
wire n_6462;
wire n_6463;
wire n_6464;
wire n_6465;
wire n_6466;
wire n_6467;
wire n_6468;
wire n_6469;
wire n_6470;
wire n_6471;
wire n_6472;
wire n_6473;
wire n_6474;
wire n_6475;
wire n_6476;
wire n_6477;
wire n_6478;
wire n_6479;
wire n_6480;
wire n_6481;
wire n_6482;
wire n_6483;
wire n_6484;
wire n_6485;
wire n_6486;
wire n_6487;
wire n_6488;
wire n_6489;
wire n_6490;
wire n_6491;
wire n_6492;
wire n_6493;
wire n_6494;
wire n_6495;
wire n_6496;
wire n_6497;
wire n_6498;
wire n_6499;
wire n_6500;
wire n_6501;
wire n_6502;
wire n_6503;
wire n_6504;
wire n_6505;
wire n_6506;
wire n_6507;
wire n_6508;
wire n_6509;
wire n_6510;
wire n_6511;
wire n_6512;
wire n_6513;
wire n_6514;
wire n_6515;
wire n_6516;
wire n_6517;
wire n_6518;
wire n_6519;
wire n_6520;
wire n_6521;
wire n_6522;
wire n_6523;
wire n_6524;
wire n_6525;
wire n_6526;
wire n_6527;
wire n_6528;
wire n_6529;
wire n_6530;
wire n_6531;
wire n_6532;
wire n_6533;
wire n_6534;
wire n_6535;
wire n_6536;
wire n_6537;
wire n_6538;
wire n_6539;
wire n_6540;
wire n_6541;
wire n_6542;
wire n_6543;
wire n_6544;
wire n_6545;
wire n_6546;
wire n_6547;
wire n_6548;
wire n_6549;
wire n_6550;
wire n_6551;
wire n_6552;
wire n_6553;
wire n_6554;
wire n_6555;
wire n_6556;
wire n_6557;
wire n_6558;
wire n_6559;
wire n_6560;
wire n_6561;
wire n_6562;
wire n_6563;
wire n_6564;
wire n_6565;
wire n_6566;
wire n_6567;
wire n_6568;
wire n_6569;
wire n_6570;
wire n_6571;
wire n_6572;
wire n_6573;
wire n_6574;
wire n_6575;
wire n_6576;
wire n_6577;
wire n_6578;
wire n_6579;
wire n_6580;
wire n_6581;
wire n_6582;
wire n_6583;
wire n_6584;
wire n_6585;
wire n_6586;
wire n_6587;
wire n_6588;
wire n_6589;
wire n_6590;
wire n_6591;
wire n_6592;
wire n_6593;
wire n_6594;
wire n_6595;
wire n_6596;
wire n_6597;
wire n_6598;
wire n_6599;
wire n_6600;
wire n_6601;
wire n_6602;
wire n_6603;
wire n_6604;
wire n_6605;
wire n_6606;
wire n_6607;
wire n_6608;
wire n_6609;
wire n_6610;
wire n_6611;
wire n_6612;
wire n_6613;
wire n_6614;
wire n_6615;
wire n_6616;
wire n_6617;
wire n_6618;
wire n_6619;
wire n_6620;
wire n_6621;
wire n_6622;
wire n_6623;
wire n_6624;
wire n_6625;
wire n_6626;
wire n_6627;
wire n_6628;
wire n_6629;
wire n_6630;
wire n_6631;
wire n_6632;
wire n_6633;
wire n_6634;
wire n_6635;
wire n_6636;
wire n_6637;
wire n_6638;
wire n_6639;
wire n_6640;
wire n_6641;
wire n_6642;
wire n_6643;
wire n_6644;
wire n_6645;
wire n_6646;
wire n_6647;
wire n_6648;
wire n_6649;
wire n_6650;
wire n_6651;
wire n_6652;
wire n_6653;
wire n_6654;
wire n_6655;
wire n_6656;
wire n_6657;
wire n_6658;
wire n_6659;
wire n_6660;
wire n_6661;
wire n_6662;
wire n_6663;
wire n_6664;
wire n_6665;
wire n_6666;
wire n_6667;
wire n_6668;
wire n_6669;
wire n_6670;
wire n_6671;
wire n_6672;
wire n_6673;
wire n_6674;
wire n_6675;
wire n_6676;
wire n_6677;
wire n_6678;
wire n_6679;
wire n_6680;
wire n_6681;
wire n_6682;
wire n_6683;
wire n_6684;
wire n_6685;
wire n_6686;
wire n_6687;
wire n_6688;
wire n_6689;
wire n_6690;
wire n_6691;
wire n_6692;
wire n_6693;
wire n_6694;
wire n_6695;
wire n_6696;
wire n_6697;
wire n_6698;
wire n_6699;
wire n_6700;
wire n_6701;
wire n_6702;
wire n_6703;
wire n_6704;
wire n_6705;
wire n_6706;
wire n_6707;
wire n_6708;
wire n_6709;
wire n_6710;
wire n_6711;
wire n_6712;
wire n_6713;
wire n_6714;
wire n_6715;
wire n_6716;
wire n_6717;
wire n_6718;
wire n_6719;
wire n_6720;
wire n_6721;
wire n_6722;
wire n_6723;
wire n_6724;
wire n_6725;
wire n_6726;
wire n_6727;
wire n_6728;
wire n_6729;
wire n_6730;
wire n_6731;
wire n_6732;
wire n_6733;
wire n_6734;
wire n_6735;
wire n_6736;
wire n_6737;
wire n_6738;
wire n_6739;
wire n_6740;
wire n_6741;
wire n_6742;
wire n_6743;
wire n_6744;
wire n_6745;
wire n_6746;
wire n_6747;
wire n_6748;
wire n_6749;
wire n_6750;
wire n_6751;
wire n_6752;
wire n_6753;
wire n_6754;
wire n_6755;
wire n_6756;
wire n_6757;
wire n_6758;
wire n_6759;
wire n_6760;
wire n_6761;
wire n_6762;
wire n_6763;
wire n_6764;
wire n_6765;
wire n_6766;
wire n_6767;
wire n_6768;
wire n_6769;
wire n_6770;
wire n_6771;
wire n_6772;
wire n_6773;
wire n_6774;
wire n_6775;
wire n_6776;
wire n_6777;
wire n_6778;
wire n_6779;
wire n_6780;
wire n_6781;
wire n_6782;
wire n_6783;
wire n_6784;
wire n_6785;
wire n_6786;
wire n_6787;
wire n_6788;
wire n_6789;
wire n_6790;
wire n_6791;
wire n_6792;
wire n_6793;
wire n_6794;
wire n_6795;
wire n_6796;
wire n_6797;
wire n_6798;
wire n_6799;
wire n_6800;
wire n_6801;
wire n_6802;
wire n_6803;
wire n_6804;
wire n_6805;
wire n_6806;
wire n_6807;
wire n_6808;
wire n_6809;
wire n_6810;
wire n_6811;
wire n_6812;
wire n_6813;
wire n_6814;
wire n_6815;
wire n_6816;
wire n_6817;
wire n_6818;
wire n_6819;
wire n_6820;
wire n_6821;
wire n_6822;
wire n_6823;
wire n_6824;
wire n_6825;
wire n_6826;
wire n_6827;
wire n_6828;
wire n_6829;
wire n_6830;
wire n_6831;
wire n_6832;
wire n_6833;
wire n_6834;
wire n_6835;
wire n_6836;
wire n_6837;
wire n_6838;
wire n_6839;
wire n_6840;
wire n_6841;
wire n_6842;
wire n_6843;
wire n_6844;
wire n_6845;
wire n_6846;
wire n_6847;
wire n_6848;
wire n_6849;
wire n_6850;
wire n_6851;
wire n_6852;
wire n_6853;
wire n_6854;
wire n_6855;
wire n_6856;
wire n_6857;
wire n_6858;
wire n_6859;
wire n_6860;
wire n_6861;
wire n_6862;
wire n_6863;
wire n_6864;
wire n_6865;
wire n_6866;
wire n_6867;
wire n_6868;
wire n_6869;
wire n_6870;
wire n_6871;
wire n_6872;
wire n_6873;
wire n_6874;
wire n_6875;
wire n_6876;
wire n_6877;
wire n_6878;
wire n_6879;
wire n_6880;
wire n_6881;
wire n_6882;
wire n_6883;
wire n_6884;
wire n_6885;
wire n_6886;
wire n_6887;
wire n_6888;
wire n_6889;
wire n_6890;
wire n_6891;
wire n_6892;
wire n_6893;
wire n_6894;
wire n_6895;
wire n_6896;
wire n_6897;
wire n_6898;
wire n_6899;
wire n_6900;
wire n_6901;
wire n_6902;
wire n_6903;
wire n_6904;
wire n_6905;
wire n_6906;
wire n_6907;
wire n_6908;
wire n_6909;
wire n_6910;
wire n_6911;
wire n_6912;
wire n_6913;
wire n_6914;
wire n_6915;
wire n_6916;
wire n_6917;
wire n_6918;
wire n_6919;
wire n_6920;
wire n_6921;
wire n_6922;
wire n_6923;
wire n_6924;
wire n_6925;
wire n_6926;
wire n_6927;
wire n_6928;
wire n_6929;
wire n_6930;
wire n_6931;
wire n_6932;
wire n_6933;
wire n_6934;
wire n_6935;
wire n_6936;
wire n_6937;
wire n_6938;
wire n_6939;
wire n_6940;
wire n_6941;
wire n_6942;
wire n_6943;
wire n_6944;
wire n_6945;
wire n_6946;
wire n_6947;
wire n_6948;
wire n_6949;
wire n_6950;
wire n_6951;
wire n_6952;
wire n_6953;
wire n_6954;
wire n_6955;
wire n_6956;
wire n_6957;
wire n_6958;
wire n_6959;
wire n_6960;
wire n_6961;
wire n_6962;
wire n_6963;
wire n_6964;
wire n_6965;
wire n_6966;
wire n_6967;
wire n_6968;
wire n_6969;
wire n_6970;
wire n_6971;
wire n_6972;
wire n_6973;
wire n_6974;
wire n_6975;
wire n_6976;
wire n_6977;
wire n_6978;
wire n_6979;
wire n_6980;
wire n_6981;
wire n_6982;
wire n_6983;
wire n_6984;
wire n_6985;
wire n_6986;
wire n_6987;
wire n_6988;
wire n_6989;
wire n_6990;
wire n_6991;
wire n_6992;
wire n_6993;
wire n_6994;
wire n_6995;
wire n_6996;
wire n_6997;
wire n_6998;
wire n_6999;
wire n_7000;
wire n_7001;
wire n_7002;
wire n_7003;
wire n_7004;
wire n_7005;
wire n_7006;
wire n_7007;
wire n_7008;
wire n_7009;
wire n_7010;
wire n_7011;
wire n_7012;
wire n_7013;
wire n_7014;
wire n_7015;
wire n_7016;
wire n_7017;
wire n_7018;
wire n_7019;
wire n_7020;
wire n_7021;
wire n_7022;
wire n_7023;
wire n_7024;
wire n_7025;
wire n_7026;
wire n_7027;
wire n_7028;
wire n_7029;
wire n_7030;
wire n_7031;
wire n_7032;
wire n_7033;
wire n_7034;
wire n_7035;
wire n_7036;
wire n_7037;
wire n_7038;
wire n_7039;
wire n_7040;
wire n_7041;
wire n_7042;
wire n_7043;
wire n_7044;
wire n_7045;
wire n_7046;
wire n_7047;
wire n_7048;
wire n_7049;
wire n_7050;
wire n_7051;
wire n_7052;
wire n_7053;
wire n_7054;
wire n_7055;
wire n_7056;
wire n_7057;
wire n_7058;
wire n_7059;
wire n_7060;
wire n_7061;
wire n_7062;
wire n_7063;
wire n_7064;
wire n_7065;
wire n_7066;
wire n_7067;
wire n_7068;
wire n_7069;
wire n_7070;
wire n_7071;
wire n_7072;
wire n_7073;
wire n_7074;
wire n_7075;
wire n_7076;
wire n_7077;
wire n_7078;
wire n_7079;
wire n_7080;
wire n_7081;
wire n_7082;
wire n_7083;
wire n_7084;
wire n_7085;
wire n_7086;
wire n_7087;
wire n_7088;
wire n_7089;
wire n_7090;
wire n_7091;
wire n_7092;
wire n_7093;
wire n_7094;
wire n_7095;
wire n_7096;
wire n_7097;
wire n_7098;
wire n_7099;
wire n_7100;
wire n_7101;
wire n_7102;
wire n_7103;
wire n_7104;
wire n_7105;
wire n_7106;
wire n_7107;
wire n_7108;
wire n_7109;
wire n_7110;
wire n_7111;
wire n_7112;
wire n_7113;
wire n_7114;
wire n_7115;
wire n_7116;
wire n_7117;
wire n_7118;
wire n_7119;
wire n_7120;
wire n_7121;
wire n_7122;
wire n_7123;
wire n_7124;
wire n_7125;
wire n_7126;
wire n_7127;
wire n_7128;
wire n_7129;
wire n_7130;
wire n_7131;
wire n_7132;
wire n_7133;
wire n_7134;
wire n_7135;
wire n_7136;
wire n_7137;
wire n_7138;
wire n_7139;
wire n_7140;
wire n_7141;
wire n_7142;
wire n_7143;
wire n_7144;
wire n_7145;
wire n_7146;
wire n_7147;
wire n_7148;
wire n_7149;
wire n_7150;
wire n_7151;
wire n_7152;
wire n_7153;
wire n_7154;
wire n_7155;
wire n_7156;
wire n_7157;
wire n_7158;
wire n_7159;
wire n_7160;
wire n_7161;
wire n_7162;
wire n_7163;
wire n_7164;
wire n_7165;
wire n_7166;
wire n_7167;
wire n_7168;
wire n_7169;
wire n_7170;
wire n_7171;
wire n_7172;
wire n_7173;
wire n_7174;
wire n_7175;
wire n_7176;
wire n_7177;
wire n_7178;
wire n_7179;
wire n_7180;
wire n_7181;
wire n_7182;
wire n_7183;
wire n_7184;
wire n_7185;
wire n_7186;
wire n_7187;
wire n_7188;
wire n_7189;
wire n_7190;
wire n_7191;
wire n_7192;
wire n_7193;
wire n_7194;
wire n_7195;
wire n_7196;
wire n_7197;
wire n_7198;
wire n_7199;
wire n_7200;
wire n_7201;
wire n_7202;
wire n_7203;
wire n_7204;
wire n_7205;
wire n_7206;
wire n_7207;
wire n_7208;
wire n_7209;
wire n_7210;
wire n_7211;
wire n_7212;
wire n_7213;
wire n_7214;
wire n_7215;
wire n_7216;
wire n_7217;
wire n_7218;
wire n_7219;
wire n_7220;
wire n_7221;
wire n_7222;
wire n_7223;
wire n_7224;
wire n_7225;
wire n_7226;
wire n_7227;
wire n_7228;
wire n_7229;
wire n_7230;
wire n_7231;
wire n_7232;
wire n_7233;
wire n_7234;
wire n_7235;
wire n_7236;
wire n_7237;
wire n_7238;
wire n_7239;
wire n_7240;
wire n_7241;
wire n_7242;
wire n_7243;
wire n_7244;
wire n_7245;
wire n_7246;
wire n_7247;
wire n_7248;
wire n_7249;
wire n_7250;
wire n_7251;
wire n_7252;
wire n_7253;
wire n_7254;
wire n_7255;
wire n_7256;
wire n_7257;
wire n_7258;
wire n_7259;
wire n_7260;
wire n_7261;
wire n_7262;
wire n_7263;
wire n_7264;
wire n_7265;
wire n_7266;
wire n_7267;
wire n_7268;
wire n_7269;
wire n_7270;
wire n_7271;
wire n_7272;
wire n_7273;
wire n_7274;
wire n_7275;
wire n_7276;
wire n_7277;
wire n_7278;
wire n_7279;
wire n_7280;
wire n_7281;
wire n_7282;
wire n_7283;
wire n_7284;
wire n_7285;
wire n_7286;
wire n_7287;
wire n_7288;
wire n_7289;
wire n_7290;
wire n_7291;
wire n_7292;
wire n_7293;
wire n_7294;
wire n_7295;
wire n_7296;
wire n_7297;
wire n_7298;
wire n_7299;
wire n_7300;
wire n_7301;
wire n_7302;
wire n_7303;
wire n_7304;
wire n_7305;
wire n_7306;
wire n_7307;
wire n_7308;
wire n_7309;
wire n_7310;
wire n_7311;
wire n_7312;
wire n_7313;
wire n_7314;
wire n_7315;
wire n_7316;
wire n_7317;
wire n_7318;
wire n_7319;
wire n_7320;
wire n_7321;
wire n_7322;
wire n_7323;
wire n_7324;
wire n_7325;
wire n_7326;
wire n_7327;
wire n_7328;
wire n_7329;
wire n_7330;
wire n_7331;
wire n_7332;
wire n_7333;
wire n_7334;
wire n_7335;
wire n_7336;
wire n_7337;
wire n_7338;
wire n_7339;
wire n_7340;
wire n_7341;
wire n_7342;
wire n_7343;
wire n_7344;
wire n_7345;
wire n_7346;
wire n_7347;
wire n_7348;
wire n_7349;
wire n_7350;
wire n_7351;
wire n_7352;
wire n_7353;
wire n_7354;
wire n_7355;
wire n_7356;
wire n_7357;
wire n_7358;
wire n_7359;
wire n_7360;
wire n_7361;
wire n_7362;
wire n_7363;
wire n_7364;
wire n_7365;
wire n_7366;
wire n_7367;
wire n_7368;
wire n_7369;
wire n_7370;
wire n_7371;
wire n_7372;
wire n_7373;
wire n_7374;
wire n_7375;
wire n_7376;
wire n_7377;
wire n_7378;
wire n_7379;
wire n_7380;
wire n_7381;
wire n_7382;
wire n_7383;
wire n_7384;
wire n_7385;
wire n_7386;
wire n_7387;
wire n_7388;
wire n_7389;
wire n_7390;
wire n_7391;
wire n_7392;
wire n_7393;
wire n_7394;
wire n_7395;
wire n_7396;
wire n_7397;
wire n_7398;
wire n_7399;
wire n_7400;
wire n_7401;
wire n_7402;
wire n_7403;
wire n_7404;
wire n_7405;
wire n_7406;
wire n_7407;
wire n_7408;
wire n_7409;
wire n_7410;
wire n_7411;
wire n_7412;
wire n_7413;
wire n_7414;
wire n_7415;
wire n_7416;
wire n_7417;
wire n_7418;
wire n_7419;
wire n_7420;
wire n_7421;
wire n_7422;
wire n_7423;
wire n_7424;
wire n_7425;
wire n_7426;
wire n_7427;
wire n_7428;
wire n_7429;
wire n_7430;
wire n_7431;
wire n_7432;
wire n_7433;
wire n_7434;
wire n_7435;
wire n_7436;
wire n_7437;
wire n_7438;
wire n_7439;
wire n_7440;
wire n_7441;
wire n_7442;
wire n_7443;
wire n_7444;
wire n_7445;
wire n_7446;
wire n_7447;
wire n_7448;
wire n_7449;
wire n_7450;
wire n_7451;
wire n_7452;
wire n_7453;
wire n_7454;
wire n_7455;
wire n_7456;
wire n_7457;
wire n_7458;
wire n_7459;
wire n_7460;
wire n_7461;
wire n_7462;
wire n_7463;
wire n_7464;
wire n_7465;
wire n_7466;
wire n_7467;
wire n_7468;
wire n_7469;
wire n_7470;
wire n_7471;
wire n_7472;
wire n_7473;
wire n_7474;
wire n_7475;
wire n_7476;
wire n_7477;
wire n_7478;
wire n_7479;
wire n_7480;
wire n_7481;
wire n_7482;
wire n_7483;
wire n_7484;
wire n_7485;
wire n_7486;
wire n_7487;
wire n_7488;
wire n_7489;
wire n_7490;
wire n_7491;
wire n_7492;
wire n_7493;
wire n_7494;
wire n_7495;
wire n_7496;
wire n_7497;
wire n_7498;
wire n_7499;
wire n_7500;
wire n_7501;
wire n_7502;
wire n_7503;
wire n_7504;
wire n_7505;
wire n_7506;
wire n_7507;
wire n_7508;
wire n_7509;
wire n_7510;
wire n_7511;
wire n_7512;
wire n_7513;
wire n_7514;
wire n_7515;
wire n_7516;
wire n_7517;
wire n_7518;
wire n_7519;
wire n_7520;
wire n_7521;
wire n_7522;
wire n_7523;
wire n_7524;
wire n_7525;
wire n_7526;
wire n_7527;
wire n_7528;
wire n_7529;
wire n_7530;
wire n_7531;
wire n_7532;
wire n_7533;
wire n_7534;
wire n_7535;
wire n_7536;
wire n_7537;
wire n_7538;
wire n_7539;
wire n_7540;
wire n_7541;
wire n_7542;
wire n_7543;
wire n_7544;
wire n_7545;
wire n_7546;
wire n_7547;
wire n_7548;
wire n_7549;
wire n_7550;
wire n_7551;
wire n_7552;
wire n_7553;
wire n_7554;
wire n_7555;
wire n_7556;
wire n_7557;
wire n_7558;
wire n_7559;
wire n_7560;
wire n_7561;
wire n_7562;
wire n_7563;
wire n_7564;
wire n_7565;
wire n_7566;
wire n_7567;
wire n_7568;
wire n_7569;
wire n_7570;
wire n_7571;
wire n_7572;
wire n_7573;
wire n_7574;
wire n_7575;
wire n_7576;
wire n_7577;
wire n_7578;
wire n_7579;
wire n_7580;
wire n_7581;
wire n_7582;
wire n_7583;
wire n_7584;
wire n_7585;
wire n_7586;
wire n_7587;
wire n_7588;
wire n_7589;
wire n_7590;
wire n_7591;
wire n_7592;
wire n_7593;
wire n_7594;
wire n_7595;
wire n_7596;
wire n_7597;
wire n_7598;
wire n_7599;
wire n_7600;
wire n_7601;
wire n_7602;
wire n_7603;
wire n_7604;
wire n_7605;
wire n_7606;
wire n_7607;
wire n_7608;
wire n_7609;
wire n_7610;
wire n_7611;
wire n_7612;
wire n_7613;
wire n_7614;
wire n_7615;
wire n_7616;
wire n_7617;
wire n_7618;
wire n_7619;
wire n_7620;
wire n_7621;
wire n_7622;
wire n_7623;
wire n_7624;
wire n_7625;
wire n_7626;
wire n_7627;
wire n_7628;
wire n_7629;
wire n_7630;
wire n_7631;
wire n_7632;
wire n_7633;
wire n_7634;
wire n_7635;
wire n_7636;
wire n_7637;
wire n_7638;
wire n_7639;
wire n_7640;
wire n_7641;
wire n_7642;
wire n_7643;
wire n_7644;
wire n_7645;
wire n_7646;
wire n_7647;
wire n_7648;
wire n_7649;
wire n_7650;
wire n_7651;
wire n_7652;
wire n_7653;
wire n_7654;
wire n_7655;
wire n_7656;
wire n_7657;
wire n_7658;
wire n_7659;
wire n_7660;
wire n_7661;
wire n_7662;
wire n_7663;
wire n_7664;
wire n_7665;
wire n_7666;
wire n_7667;
wire n_7668;
wire n_7669;
wire n_7670;
wire n_7671;
wire n_7672;
wire n_7673;
wire n_7674;
wire n_7675;
wire n_7676;
wire n_7677;
wire n_7678;
wire n_7679;
wire n_7680;
wire n_7681;
wire n_7682;
wire n_7683;
wire n_7684;
wire n_7685;
wire n_7686;
wire n_7687;
wire n_7688;
wire n_7689;
wire n_7690;
wire n_7691;
wire n_7692;
wire n_7693;
wire n_7694;
wire n_7695;
wire n_7696;
wire n_7697;
wire n_7698;
wire n_7699;
wire n_7700;
wire n_7701;
wire n_7702;
wire n_7703;
wire n_7704;
wire n_7705;
wire n_7706;
wire n_7707;
wire n_7708;
wire n_7709;
wire n_7710;
wire n_7711;
wire n_7712;
wire n_7713;
wire n_7714;
wire n_7715;
wire n_7716;
wire n_7717;
wire n_7718;
wire n_7719;
wire n_7720;
wire n_7721;
wire n_7722;
wire n_7723;
wire n_7724;
wire n_7725;
wire n_7726;
wire n_7727;
wire n_7728;
wire n_7729;
wire n_7730;
wire n_7731;
wire n_7732;
wire n_7733;
wire n_7734;
wire n_7735;
wire n_7736;
wire n_7737;
wire n_7738;
wire n_7739;
wire n_7740;
wire n_7741;
wire n_7742;
wire n_7743;
wire n_7744;
wire n_7745;
wire n_7746;
wire n_7747;
wire n_7748;
wire n_7749;
wire n_7750;
wire n_7751;
wire n_7752;
wire n_7753;
wire n_7754;
wire n_7755;
wire n_7756;
wire n_7757;
wire n_7758;
wire n_7759;
wire n_7760;
wire n_7761;
wire n_7762;
wire n_7763;
wire n_7764;
wire n_7765;
wire n_7766;
wire n_7767;
wire n_7768;
wire n_7769;
wire n_7770;
wire n_7771;
wire n_7772;
wire n_7773;
wire n_7774;
wire n_7775;
wire n_7776;
wire n_7777;
wire n_7778;
wire n_7779;
wire n_7780;
wire n_7781;
wire n_7782;
wire n_7783;
wire n_7784;
wire n_7785;
wire n_7786;
wire n_7787;
wire n_7788;
wire n_7789;
wire n_7790;
wire n_7791;
wire n_7792;
wire n_7793;
wire n_7794;
wire n_7795;
wire n_7796;
wire n_7797;
wire n_7798;
wire n_7799;
wire n_7800;
wire n_7801;
wire n_7802;
wire n_7803;
wire n_7804;
wire n_7805;
wire n_7806;
wire n_7807;
wire n_7808;
wire n_7809;
wire n_7810;
wire n_7811;
wire n_7812;
wire n_7813;
wire n_7814;
wire n_7815;
wire n_7816;
wire n_7817;
wire n_7818;
wire n_7819;
wire n_7820;
wire n_7821;
wire n_7822;
wire n_7823;
wire n_7824;
wire n_7825;
wire n_7826;
wire n_7827;
wire n_7828;
wire n_7829;
wire n_7830;
wire n_7831;
wire n_7832;
wire n_7833;
wire n_7834;
wire n_7835;
wire n_7836;
wire n_7837;
wire n_7838;
wire n_7839;
wire n_7840;
wire n_7841;
wire n_7842;
wire n_7843;
wire n_7844;
wire n_7845;
wire n_7846;
wire n_7847;
wire n_7848;
wire n_7849;
wire n_7850;
wire n_7851;
wire n_7852;
wire n_7853;
wire n_7854;
wire n_7855;
wire n_7856;
wire n_7857;
wire n_7858;
wire n_7859;
wire n_7860;
wire n_7861;
wire n_7862;
wire n_7863;
wire n_7864;
wire n_7865;
wire n_7866;
wire n_7867;
wire n_7868;
wire n_7869;
wire n_7870;
wire n_7871;
wire n_7872;
wire n_7873;
wire n_7874;
wire n_7875;
wire n_7876;
wire n_7877;
wire n_7878;
wire n_7879;
wire n_7880;
wire n_7881;
wire n_7882;
wire n_7883;
wire n_7884;
wire n_7885;
wire n_7886;
wire n_7887;
wire n_7888;
wire n_7889;
wire n_7890;
wire n_7891;
wire n_7892;
wire n_7893;
wire n_7894;
wire n_7895;
wire n_7896;
wire n_7897;
wire n_7898;
wire n_7899;
wire n_7900;
wire n_7901;
wire n_7902;
wire n_7903;
wire n_7904;
wire n_7905;
wire n_7906;
wire n_7907;
wire n_7908;
wire n_7909;
wire n_7910;
wire n_7911;
wire n_7912;
wire n_7913;
wire n_7914;
wire n_7915;
wire n_7916;
wire n_7917;
wire n_7918;
wire n_7919;
wire n_7920;
wire n_7921;
wire n_7922;
wire n_7923;
wire n_7924;
wire n_7925;
wire n_7926;
wire n_7927;
wire n_7928;
wire n_7929;
wire n_7930;
wire n_7931;
wire n_7932;
wire n_7933;
wire n_7934;
wire n_7935;
wire n_7936;
wire n_7937;
wire n_7938;
wire n_7939;
wire n_7940;
wire n_7941;
wire n_7942;
wire n_7943;
wire n_7944;
wire n_7945;
wire n_7946;
wire n_7947;
wire n_7948;
wire n_7949;
wire n_7950;
wire n_7951;
wire n_7952;
wire n_7953;
wire n_7954;
wire n_7955;
wire n_7956;
wire n_7957;
wire n_7958;
wire n_7959;
wire n_7960;
wire n_7961;
wire n_7962;
wire n_7963;
wire n_7964;
wire n_7965;
wire n_7966;
wire n_7967;
wire n_7968;
wire n_7969;
wire n_7970;
wire n_7971;
wire n_7972;
wire n_7973;
wire n_7974;
wire n_7975;
wire n_7976;
wire n_7977;
wire n_7978;
wire n_7979;
wire n_7980;
wire n_7981;
wire n_7982;
wire n_7983;
wire n_7984;
wire n_7985;
wire n_7986;
wire n_7987;
wire n_7988;
wire n_7989;
wire n_7990;
wire n_7991;
wire n_7992;
wire n_7993;
wire n_7994;
wire n_7995;
wire n_7996;
wire n_7997;
wire n_7998;
wire n_7999;
wire n_8000;
wire n_8001;
wire n_8002;
wire n_8003;
wire n_8004;
wire n_8005;
wire n_8006;
wire n_8007;
wire n_8008;
wire n_8009;
wire n_8010;
wire n_8011;
wire n_8012;
wire n_8013;
wire n_8014;
wire n_8015;
wire n_8016;
wire n_8017;
wire n_8018;
wire n_8019;
wire n_8020;
wire n_8021;
wire n_8022;
wire n_8023;
wire n_8024;
wire n_8025;
wire n_8026;
wire n_8027;
wire n_8028;
wire n_8029;
wire n_8030;
wire n_8031;
wire n_8032;
wire n_8033;
wire n_8034;
wire n_8035;
wire n_8036;
wire n_8037;
wire n_8038;
wire n_8039;
wire n_8040;
wire n_8041;
wire n_8042;
wire n_8043;
wire n_8044;
wire n_8045;
wire n_8046;
wire n_8047;
wire n_8048;
wire n_8049;
wire n_8050;
wire n_8051;
wire n_8052;
wire n_8053;
wire n_8054;
wire n_8055;
wire n_8056;
wire n_8057;
wire n_8058;
wire n_8059;
wire n_8060;
wire n_8061;
wire n_8062;
wire n_8063;
wire n_8064;
wire n_8065;
wire n_8066;
wire n_8067;
wire n_8068;
wire n_8069;
wire n_8070;
wire n_8071;
wire n_8072;
wire n_8073;
wire n_8074;
wire n_8075;
wire n_8076;
wire n_8077;
wire n_8078;
wire n_8079;
wire n_8080;
wire n_8081;
wire n_8082;
wire n_8083;
wire n_8084;
wire n_8085;
wire n_8086;
wire n_8087;
wire n_8088;
wire n_8089;
wire n_8090;
wire n_8091;
wire n_8092;
wire n_8093;
wire n_8094;
wire n_8095;
wire n_8096;
wire n_8097;
wire n_8098;
wire n_8099;
wire n_8100;
wire n_8101;
wire n_8102;
wire n_8103;
wire n_8104;
wire n_8105;
wire n_8106;
wire n_8107;
wire n_8108;
wire n_8109;
wire n_8110;
wire n_8111;
wire n_8112;
wire n_8113;
wire n_8114;
wire n_8115;
wire n_8116;
wire n_8117;
wire n_8118;
wire n_8119;
wire n_8120;
wire n_8121;
wire n_8122;
wire n_8123;
wire n_8124;
wire n_8125;
wire n_8126;
wire n_8127;
wire n_8128;
wire n_8129;
wire n_8130;
wire n_8131;
wire n_8132;
wire n_8133;
wire n_8134;
wire n_8135;
wire n_8136;
wire n_8137;
wire n_8138;
wire n_8139;
wire n_8140;
wire n_8141;
wire n_8142;
wire n_8143;
wire n_8144;
wire n_8145;
wire n_8146;
wire n_8147;
wire n_8148;
wire n_8149;
wire n_8150;
wire n_8151;
wire n_8152;
wire n_8153;
wire n_8154;
wire n_8155;
wire n_8156;
wire n_8157;
wire n_8158;
wire n_8159;
wire n_8160;
wire n_8161;
wire n_8162;
wire n_8163;
wire n_8164;
wire n_8165;
wire n_8166;
wire n_8167;
wire n_8168;
wire n_8169;
wire n_8170;
wire n_8171;
wire n_8172;
wire n_8173;
wire n_8174;
wire n_8175;
wire n_8176;
wire n_8177;
wire n_8178;
wire n_8179;
wire n_8180;
wire n_8181;
wire n_8182;
wire n_8183;
wire n_8184;
wire n_8185;
wire n_8186;
wire n_8187;
wire n_8188;
wire n_8189;
wire n_8190;
wire n_8191;
wire n_8192;
wire n_8193;
wire n_8194;
wire n_8195;
wire n_8196;
wire n_8197;
wire n_8198;
wire n_8199;
wire n_8200;
wire n_8201;
wire n_8202;
wire n_8203;
wire n_8204;
wire n_8205;
wire n_8206;
wire n_8207;
wire n_8208;
wire n_8209;
wire n_8210;
wire n_8211;
wire n_8212;
wire n_8213;
wire n_8214;
wire n_8215;
wire n_8216;
wire n_8217;
wire n_8218;
wire n_8219;
wire n_8220;
wire n_8221;
wire n_8222;
wire n_8223;
wire n_8224;
wire n_8225;
wire n_8226;
wire n_8227;
wire n_8228;
wire n_8229;
wire n_8230;
wire n_8231;
wire n_8232;
wire n_8233;
wire n_8234;
wire n_8235;
wire n_8236;
wire n_8237;
wire n_8238;
wire n_8239;
wire n_8240;
wire n_8241;
wire n_8242;
wire n_8243;
wire n_8244;
wire n_8245;
wire n_8246;
wire n_8247;
wire n_8248;
wire n_8249;
wire n_8250;
wire n_8251;
wire n_8252;
wire n_8253;
wire n_8254;
wire n_8255;
wire n_8256;
wire n_8257;
wire n_8258;
wire n_8259;
wire n_8260;
wire n_8261;
wire n_8262;
wire n_8263;
wire n_8264;
wire n_8265;
wire n_8266;
wire n_8267;
wire n_8268;
wire n_8269;
wire n_8270;
wire n_8271;
wire n_8272;
wire n_8273;
wire n_8274;
wire n_8275;
wire n_8276;
wire n_8277;
wire n_8278;
wire n_8279;
wire n_8280;
wire n_8281;
wire n_8282;
wire n_8283;
wire n_8284;
wire n_8285;
wire n_8286;
wire n_8287;
wire n_8288;
wire n_8289;
wire n_8290;
wire n_8291;
wire n_8292;
wire n_8293;
wire n_8294;
wire n_8295;
wire n_8296;
wire n_8297;
wire n_8298;
wire n_8299;
wire n_8300;
wire n_8301;
wire n_8302;
wire n_8303;
wire n_8304;
wire n_8305;
wire n_8306;
wire n_8307;
wire n_8308;
wire n_8309;
wire n_8310;
wire n_8311;
wire n_8312;
wire n_8313;
wire n_8314;
wire n_8315;
wire n_8316;
wire n_8317;
wire n_8318;
wire n_8319;
wire n_8320;
wire n_8321;
wire n_8322;
wire n_8323;
wire n_8324;
wire n_8325;
wire n_8326;
wire n_8327;
wire n_8328;
wire n_8329;
wire n_8330;
wire n_8331;
wire n_8332;
wire n_8333;
wire n_8334;
wire n_8335;
wire n_8336;
wire n_8337;
wire n_8338;
wire n_8339;
wire n_8340;
wire n_8341;
wire n_8342;
wire n_8343;
wire n_8344;
wire n_8345;
wire n_8346;
wire n_8347;
wire n_8348;
wire n_8349;
wire n_8350;
wire n_8351;
wire n_8352;
wire n_8353;
wire n_8354;
wire n_8355;
wire n_8356;
wire n_8357;
wire n_8358;
wire n_8359;
wire n_8360;
wire n_8361;
wire n_8362;
wire n_8363;
wire n_8364;
wire n_8365;
wire n_8366;
wire n_8367;
wire n_8368;
wire n_8369;
wire n_8370;
wire n_8371;
wire n_8372;
wire n_8373;
wire n_8374;
wire n_8375;
wire n_8376;
wire n_8377;
wire n_8378;
wire n_8379;
wire n_8380;
wire n_8381;
wire n_8382;
wire n_8383;
wire n_8384;
wire n_8385;
wire n_8386;
wire n_8387;
wire n_8388;
wire n_8389;
wire n_8390;
wire n_8391;
wire n_8392;
wire n_8393;
wire n_8394;
wire n_8395;
wire n_8396;
wire n_8397;
wire n_8398;
wire n_8399;
wire n_8400;
wire n_8401;
wire n_8402;
wire n_8403;
wire n_8404;
wire n_8405;
wire n_8406;
wire n_8407;
wire n_8408;
wire n_8409;
wire n_8410;
wire n_8411;
wire n_8412;
wire n_8413;
wire n_8414;
wire n_8415;
wire n_8416;
wire n_8417;
wire n_8418;
wire n_8419;
wire n_8420;
wire n_8421;
wire n_8422;
wire n_8423;
wire n_8424;
wire n_8425;
wire n_8426;
wire n_8427;
wire n_8428;
wire n_8429;
wire n_8430;
wire n_8431;
wire n_8432;
wire n_8433;
wire n_8434;
wire n_8435;
wire n_8436;
wire n_8437;
wire n_8438;
wire n_8439;
wire n_8440;
wire n_8441;
wire n_8442;
wire n_8443;
wire n_8444;
wire n_8445;
wire n_8446;
wire n_8447;
wire n_8448;
wire n_8449;
wire n_8450;
wire n_8451;
wire n_8452;
wire n_8453;
wire n_8454;
wire n_8455;
wire n_8456;
wire n_8457;
wire n_8458;
wire n_8459;
wire n_8460;
wire n_8461;
wire n_8462;
wire n_8463;
wire n_8464;
wire n_8465;
wire n_8466;
wire n_8467;
wire n_8468;
wire n_8469;
wire n_8470;
wire n_8471;
wire n_8472;
wire n_8473;
wire n_8474;
wire n_8475;
wire n_8476;
wire n_8477;
wire n_8478;
wire n_8479;
wire n_8480;
wire n_8481;
wire n_8482;
wire n_8483;
wire n_8484;
wire n_8485;
wire n_8486;
wire n_8487;
wire n_8488;
wire n_8489;
wire n_8490;
wire n_8491;
wire n_8492;
wire n_8493;
wire n_8494;
wire n_8495;
wire n_8496;
wire n_8497;
wire n_8498;
wire n_8499;
wire n_8500;
wire n_8501;
wire n_8502;
wire n_8503;
wire n_8504;
wire n_8505;
wire n_8506;
wire n_8507;
wire n_8508;
wire n_8509;
wire n_8510;
wire n_8511;
wire n_8512;
wire n_8513;
wire n_8514;
wire n_8515;
wire n_8516;
wire n_8517;
wire n_8518;
wire n_8519;
wire n_8520;
wire n_8521;
wire n_8522;
wire n_8523;
wire n_8524;
wire n_8525;
wire n_8526;
wire n_8527;
wire n_8528;
wire n_8529;
wire n_8530;
wire n_8531;
wire n_8532;
wire n_8533;
wire n_8534;
wire n_8535;
wire n_8536;
wire n_8537;
wire n_8538;
wire n_8539;
wire n_8540;
wire n_8541;
wire n_8542;
wire n_8543;
wire n_8544;
wire n_8545;
wire n_8546;
wire n_8547;
wire n_8548;
wire n_8549;
wire n_8550;
wire n_8551;
wire n_8552;
wire n_8553;
wire n_8554;
wire n_8555;
wire n_8556;
wire n_8557;
wire n_8558;
wire n_8559;
wire n_8560;
wire n_8561;
wire n_8562;
wire n_8563;
wire n_8564;
wire n_8565;
wire n_8566;
wire n_8567;
wire n_8568;
wire n_8569;
wire n_8570;
wire n_8571;
wire n_8572;
wire n_8573;
wire n_8574;
wire n_8575;
wire n_8576;
wire n_8577;
wire n_8578;
wire n_8579;
wire n_8580;
wire n_8581;
wire n_8582;
wire n_8583;
wire n_8584;
wire n_8585;
wire n_8586;
wire n_8587;
wire n_8588;
wire n_8589;
wire n_8590;
wire n_8591;
wire n_8592;
wire n_8593;
wire n_8594;
wire n_8595;
wire n_8596;
wire n_8597;
wire n_8598;
wire n_8599;
wire n_8600;
wire n_8601;
wire n_8602;
wire n_8603;
wire n_8604;
wire n_8605;
wire n_8606;
wire n_8607;
wire n_8608;
wire n_8609;
wire n_8610;
wire n_8611;
wire n_8612;
wire n_8613;
wire n_8614;
wire n_8615;
wire n_8616;
wire n_8617;
wire n_8618;
wire n_8619;
wire n_8620;
wire n_8621;
wire n_8622;
wire n_8623;
wire n_8624;
wire n_8625;
wire n_8626;
wire n_8627;
wire n_8628;
wire n_8629;
wire n_8630;
wire n_8631;
wire n_8632;
wire n_8633;
wire n_8634;
wire n_8635;
wire n_8636;
wire n_8637;
wire n_8638;
wire n_8639;
wire n_8640;
wire n_8641;
wire n_8642;
wire n_8643;
wire n_8644;
wire n_8645;
wire n_8646;
wire n_8647;
wire n_8648;
wire n_8649;
wire n_8650;
wire n_8651;
wire n_8652;
wire n_8653;
wire n_8654;
wire n_8655;
wire n_8656;
wire n_8657;
wire n_8658;
wire n_8659;
wire n_8660;
wire n_8661;
wire n_8662;
wire n_8663;
wire n_8664;
wire n_8665;
wire n_8666;
wire n_8667;
wire n_8668;
wire n_8669;
wire n_8670;
wire n_8671;
wire n_8672;
wire n_8673;
wire n_8674;
wire n_8675;
wire n_8676;
wire n_8677;
wire n_8678;
wire n_8679;
wire n_8680;
wire n_8681;
wire n_8682;
wire n_8683;
wire n_8684;
wire n_8685;
wire n_8686;
wire n_8687;
wire n_8688;
wire n_8689;
wire n_8690;
wire n_8691;
wire n_8692;
wire n_8693;
wire n_8694;
wire n_8695;
wire n_8696;
wire n_8697;
wire n_8698;
wire n_8699;
wire n_8700;
wire n_8701;
wire n_8702;
wire n_8703;
wire n_8704;
wire n_8705;
wire n_8706;
wire n_8707;
wire n_8708;
wire n_8709;
wire n_8710;
wire n_8711;
wire n_8712;
wire n_8713;
wire n_8714;
wire n_8715;
wire n_8716;
wire n_8717;
wire n_8718;
wire n_8719;
wire n_8720;
wire n_8721;
wire n_8722;
wire n_8723;
wire n_8724;
wire n_8725;
wire n_8726;
wire n_8727;
wire n_8728;
wire n_8729;
wire n_8730;
wire n_8731;
wire n_8732;
wire n_8733;
wire n_8734;
wire n_8735;
wire n_8736;
wire n_8737;
wire n_8738;
wire n_8739;
wire n_8740;
wire n_8741;
wire n_8742;
wire n_8743;
wire n_8744;
wire n_8745;
wire n_8746;
wire n_8747;
wire n_8748;
wire n_8749;
wire n_8750;
wire n_8751;
wire n_8752;
wire n_8753;
wire n_8754;
wire n_8755;
wire n_8756;
wire n_8757;
wire n_8758;
wire n_8759;
wire n_8760;
wire n_8761;
wire n_8762;
wire n_8763;
wire n_8764;
wire n_8765;
wire n_8766;
wire n_8767;
wire n_8768;
wire n_8769;
wire n_8770;
wire n_8771;
wire n_8772;
wire n_8773;
wire n_8774;
wire n_8775;
wire n_8776;
wire n_8777;
wire n_8778;
wire n_8779;
wire n_8780;
wire n_8781;
wire n_8782;
wire n_8783;
wire n_8784;
wire n_8785;
wire n_8786;
wire n_8787;
wire n_8788;
wire n_8789;
wire n_8790;
wire n_8791;
wire n_8792;
wire n_8793;
wire n_8794;
wire n_8795;
wire n_8796;
wire n_8797;
wire n_8798;
wire n_8799;
wire n_8800;
wire n_8801;
wire n_8802;
wire n_8803;
wire n_8804;
wire n_8805;
wire n_8806;
wire n_8807;
wire n_8808;
wire n_8809;
wire n_8810;
wire n_8811;
wire n_8812;
wire n_8813;
wire n_8814;
wire n_8815;
wire n_8816;
wire n_8817;
wire n_8818;
wire n_8819;
wire n_8820;
wire n_8821;
wire n_8822;
wire n_8823;
wire n_8824;
wire n_8825;
wire n_8826;
wire n_8827;
wire n_8828;
wire n_8829;
wire n_8830;
wire n_8831;
wire n_8832;
wire n_8833;
wire n_8834;
wire n_8835;
wire n_8836;
wire n_8837;
wire n_8838;
wire n_8839;
wire n_8840;
wire n_8841;
wire n_8842;
wire n_8843;
wire n_8844;
wire n_8845;
wire n_8846;
wire n_8847;
wire n_8848;
wire n_8849;
wire n_8850;
wire n_8851;
wire n_8852;
wire n_8853;
wire n_8854;
wire n_8855;
wire n_8856;
wire n_8857;
wire n_8858;
wire n_8859;
wire n_8860;
wire n_8861;
wire n_8862;
wire n_8863;
wire n_8864;
wire n_8865;
wire n_8866;
wire n_8867;
wire n_8868;
wire n_8869;
wire n_8870;
wire n_8871;
wire n_8872;
wire n_8873;
wire n_8874;
wire n_8875;
wire n_8876;
wire n_8877;
wire n_8878;
wire n_8879;
wire n_8880;
wire n_8881;
wire n_8882;
wire n_8883;
wire n_8884;
wire n_8885;
wire n_8886;
wire n_8887;
wire n_8888;
wire n_8889;
wire n_8890;
wire n_8891;
wire n_8892;
wire n_8893;
wire n_8894;
wire n_8895;
wire n_8896;
wire n_8897;
wire n_8898;
wire n_8899;
wire n_8900;
wire n_8901;
wire n_8902;
wire n_8903;
wire n_8904;
wire n_8905;
wire n_8906;
wire n_8907;
wire n_8908;
wire n_8909;
wire n_8910;
wire n_8911;
wire n_8912;
wire n_8913;
wire n_8914;
wire n_8915;
wire n_8916;
wire n_8917;
wire n_8918;
wire n_8919;
wire n_8920;
wire n_8921;
wire n_8922;
wire n_8923;
wire n_8924;
wire n_8925;
wire n_8926;
wire n_8927;
wire n_8928;
wire n_8929;
wire n_8930;
wire n_8931;
wire n_8932;
wire n_8933;
wire n_8934;
wire n_8935;
wire n_8936;
wire n_8937;
wire n_8938;
wire n_8939;
wire n_8940;
wire n_8941;
wire n_8942;
wire n_8943;
wire n_8944;
wire n_8945;
wire n_8946;
wire n_8947;
wire n_8948;
wire n_8949;
wire n_8950;
wire n_8951;
wire n_8952;
wire n_8953;
wire n_8954;
wire n_8955;
wire n_8956;
wire n_8957;
wire n_8958;
wire n_8959;
wire n_8960;
wire n_8961;
wire n_8962;
wire n_8963;
wire n_8964;
wire n_8965;
wire n_8966;
wire n_8967;
wire n_8968;
wire n_8969;
wire n_8970;
wire n_8971;
wire n_8972;
wire n_8973;
wire n_8974;
wire n_8975;
wire n_8976;
wire n_8977;
wire n_8978;
wire n_8979;
wire n_8980;
wire n_8981;
wire n_8982;
wire n_8983;
wire n_8984;
wire n_8985;
wire n_8986;
wire n_8987;
wire n_8988;
wire n_8989;
wire n_8990;
wire n_8991;
wire n_8992;
wire n_8993;
wire n_8994;
wire n_8995;
wire n_8996;
wire n_8997;
wire n_8998;
wire n_8999;
wire n_9000;
wire n_9001;
wire n_9002;
wire n_9003;
wire n_9004;
wire n_9005;
wire n_9006;
wire n_9007;
wire n_9008;
wire n_9009;
wire n_9010;
wire n_9011;
wire n_9012;
wire n_9013;
wire n_9014;
wire n_9015;
wire n_9016;
wire n_9017;
wire n_9018;
wire n_9019;
wire n_9020;
wire n_9021;
wire n_9022;
wire n_9023;
wire n_9024;
wire n_9025;
wire n_9026;
wire n_9027;
wire n_9028;
wire n_9029;
wire n_9030;
wire n_9031;
wire n_9032;
wire n_9033;
wire n_9034;
wire n_9035;
wire n_9036;
wire n_9037;
wire n_9038;
wire n_9039;
wire n_9040;
wire n_9041;
wire n_9042;
wire n_9043;
wire n_9044;
wire n_9045;
wire n_9046;
wire n_9047;
wire n_9048;
wire n_9049;
wire n_9050;
wire n_9051;
wire n_9052;
wire n_9053;
wire n_9054;
wire n_9055;
wire n_9056;
wire n_9057;
wire n_9058;
wire n_9059;
wire n_9060;
wire n_9061;
wire n_9062;
wire n_9063;
wire n_9064;
wire n_9065;
wire n_9066;
wire n_9067;
wire n_9068;
wire n_9069;
wire n_9070;
wire n_9071;
wire n_9072;
wire n_9073;
wire n_9074;
wire n_9075;
wire n_9076;
wire n_9077;
wire n_9078;
wire n_9079;
wire n_9080;
wire n_9081;
wire n_9082;
wire n_9083;
wire n_9084;
wire n_9085;
wire n_9086;
wire n_9087;
wire n_9088;
wire n_9089;
wire n_9090;
wire n_9091;
wire n_9092;
wire n_9093;
wire n_9094;
wire n_9095;
wire n_9096;
wire n_9097;
wire n_9098;
wire n_9099;
wire n_9100;
wire n_9101;
wire n_9102;
wire n_9103;
wire n_9104;
wire n_9105;
wire n_9106;
wire n_9107;
wire n_9108;
wire n_9109;
wire n_9110;
wire n_9111;
wire n_9112;
wire n_9113;
wire n_9114;
wire n_9115;
wire n_9116;
wire n_9117;
wire n_9118;
wire n_9119;
wire n_9120;
wire n_9121;
wire n_9122;
wire n_9123;
wire n_9124;
wire n_9125;
wire n_9126;
wire n_9127;
wire n_9128;
wire n_9129;
wire n_9130;
wire n_9131;
wire n_9132;
wire n_9133;
wire n_9134;
wire n_9135;
wire n_9136;
wire n_9137;
wire n_9138;
wire n_9139;
wire n_9140;
wire n_9141;
wire n_9142;
wire n_9143;
wire n_9144;
wire n_9145;
wire n_9146;
wire n_9147;
wire n_9148;
wire n_9149;
wire n_9150;
wire n_9151;
wire n_9152;
wire n_9153;
wire n_9154;
wire n_9155;
wire n_9156;
wire n_9157;
wire n_9158;
wire n_9159;
wire n_9160;
wire n_9161;
wire n_9162;
wire n_9163;
wire n_9164;
wire n_9165;
wire n_9166;
wire n_9167;
wire n_9168;
wire n_9169;
wire n_9170;
wire n_9171;
wire n_9172;
wire n_9173;
wire n_9174;
wire n_9175;
wire n_9176;
wire n_9177;
wire n_9178;
wire n_9179;
wire n_9180;
wire n_9181;
wire n_9182;
wire n_9183;
wire n_9184;
wire n_9185;
wire n_9186;
wire n_9187;
wire n_9188;
wire n_9189;
wire n_9190;
wire n_9191;
wire n_9192;
wire n_9193;
wire n_9194;
wire n_9195;
wire n_9196;
wire n_9197;
wire n_9198;
wire n_9199;
wire n_9200;
wire n_9201;
wire n_9202;
wire n_9203;
wire n_9204;
wire n_9205;
wire n_9206;
wire n_9207;
wire n_9208;
wire n_9209;
wire n_9210;
wire n_9211;
wire n_9212;
wire n_9213;
wire n_9214;
wire n_9215;
wire n_9216;
wire n_9217;
wire n_9218;
wire n_9219;
wire n_9220;
wire n_9221;
wire n_9222;
wire n_9223;
wire n_9224;
wire n_9225;
wire n_9226;
wire n_9227;
wire n_9228;
wire n_9229;
wire n_9230;
wire n_9231;
wire n_9232;
wire n_9233;
wire n_9234;
wire n_9235;
wire n_9236;
wire n_9237;
wire n_9238;
wire n_9239;
wire n_9240;
wire n_9241;
wire n_9242;
wire n_9243;
wire n_9244;
wire n_9245;
wire n_9246;
wire n_9247;
wire n_9248;
wire n_9249;
wire n_9250;
wire n_9251;
wire n_9252;
wire n_9253;
wire n_9254;
wire n_9255;
wire n_9256;
wire n_9257;
wire n_9258;
wire n_9259;
wire n_9260;
wire n_9261;
wire n_9262;
wire n_9263;
wire n_9264;
wire n_9265;
wire n_9266;
wire n_9267;
wire n_9268;
wire n_9269;
wire n_9270;
wire n_9271;
wire n_9272;
wire n_9273;
wire n_9274;
wire n_9275;
wire n_9276;
wire n_9277;
wire n_9278;
wire n_9279;
wire n_9280;
wire n_9281;
wire n_9282;
wire n_9283;
wire n_9284;
wire n_9285;
wire n_9286;
wire n_9287;
wire n_9288;
wire n_9289;
wire n_9290;
wire n_9291;
wire n_9292;
wire n_9293;
wire n_9294;
wire n_9295;
wire n_9296;
wire n_9297;
wire n_9298;
wire n_9299;
wire n_9300;
wire n_9301;
wire n_9302;
wire n_9303;
wire n_9304;
wire n_9305;
wire n_9306;
wire n_9307;
wire n_9308;
wire n_9309;
wire n_9310;
wire n_9311;
wire n_9312;
wire n_9313;
wire n_9314;
wire n_9315;
wire n_9316;
wire n_9317;
wire n_9318;
wire n_9319;
wire n_9320;
wire n_9321;
wire n_9322;
wire n_9323;
wire n_9324;
wire n_9325;
wire n_9326;
wire n_9327;
wire n_9328;
wire n_9329;
wire n_9330;
wire n_9331;
wire n_9332;
wire n_9333;
wire n_9334;
wire n_9335;
wire n_9336;
wire n_9337;
wire n_9338;
wire n_9339;
wire n_9340;
wire n_9341;
wire n_9342;
wire n_9343;
wire n_9344;
wire n_9345;
wire n_9346;
wire n_9347;
wire n_9348;
wire n_9349;
wire n_9350;
wire n_9351;
wire n_9352;
wire n_9353;
wire n_9354;
wire n_9355;
wire n_9356;
wire n_9357;
wire n_9358;
wire n_9359;
wire n_9360;
wire n_9361;
wire n_9362;
wire n_9363;
wire n_9364;
wire n_9365;
wire n_9366;
wire n_9367;
wire n_9368;
wire n_9369;
wire n_9370;
wire n_9371;
wire n_9372;
wire n_9373;
wire n_9374;
wire n_9375;
wire n_9376;
wire n_9377;
wire n_9378;
wire n_9379;
wire n_9380;
wire n_9381;
wire n_9382;
wire n_9383;
wire n_9384;
wire n_9385;
wire n_9386;
wire n_9387;
wire n_9388;
wire n_9389;
wire n_9390;
wire n_9391;
wire n_9392;
wire n_9393;
wire n_9394;
wire n_9395;
wire n_9396;
wire n_9397;
wire n_9398;
wire n_9399;
wire n_9400;
wire n_9401;
wire n_9402;
wire n_9403;
wire n_9404;
wire n_9405;
wire n_9406;
wire n_9407;
wire n_9408;
wire n_9409;
wire n_9410;
wire n_9411;
wire n_9412;
wire n_9413;
wire n_9414;
wire n_9415;
wire n_9416;
wire n_9417;
wire n_9418;
wire n_9419;
wire n_9420;
wire n_9421;
wire n_9422;
wire n_9423;
wire n_9424;
wire n_9425;
wire n_9426;
wire n_9427;
wire n_9428;
wire n_9429;
wire n_9430;
wire n_9431;
wire n_9432;
wire n_9433;
wire n_9434;
wire n_9435;
wire n_9436;
wire n_9437;
wire n_9438;
wire n_9439;
wire n_9440;
wire n_9441;
wire n_9442;
wire n_9443;
wire n_9444;
wire n_9445;
wire n_9446;
wire n_9447;
wire n_9448;
wire n_9449;
wire n_9450;
wire n_9451;
wire n_9452;
wire n_9453;
wire n_9454;
wire n_9455;
wire n_9456;
wire n_9457;
wire n_9458;
wire n_9459;
wire n_9460;
wire n_9461;
wire n_9462;
wire n_9463;
wire n_9464;
wire n_9465;
wire n_9466;
wire n_9467;
wire n_9468;
wire n_9469;
wire n_9470;
wire n_9471;
wire n_9472;
wire n_9473;
wire n_9474;
wire n_9475;
wire n_9476;
wire n_9477;
wire n_9478;
wire n_9479;
wire n_9480;
wire n_9481;
wire n_9482;
wire n_9483;
wire n_9484;
wire n_9485;
wire n_9486;
wire n_9487;
wire n_9488;
wire n_9489;
wire n_9490;
wire n_9491;
wire n_9492;
wire n_9493;
wire n_9494;
wire n_9495;
wire n_9496;
wire n_9497;
wire n_9498;
wire n_9499;
wire n_9500;
wire n_9501;
wire n_9502;
wire n_9503;
wire n_9504;
wire n_9505;
wire n_9506;
wire n_9507;
wire n_9508;
wire n_9509;
wire n_9510;
wire n_9511;
wire n_9512;
wire n_9513;
wire n_9514;
wire n_9515;
wire n_9516;
wire n_9517;
wire n_9518;
wire n_9519;
wire n_9520;
wire n_9521;
wire n_9522;
wire n_9523;
wire n_9524;
wire n_9525;
wire n_9526;
wire n_9527;
wire n_9528;
wire n_9529;
wire n_9530;
wire n_9531;
wire n_9532;
wire n_9533;
wire n_9534;
wire n_9535;
wire n_9536;
wire n_9537;
wire n_9538;
wire n_9539;
wire n_9540;
wire n_9541;
wire n_9542;
wire n_9543;
wire n_9544;
wire n_9545;
wire n_9546;
wire n_9547;
wire n_9548;
wire n_9549;
wire n_9550;
wire n_9551;
wire n_9552;
wire n_9553;
wire n_9554;
wire n_9555;
wire n_9556;
wire n_9557;
wire n_9558;
wire n_9559;
wire n_9560;
wire n_9561;
wire n_9562;
wire n_9563;
wire n_9564;
wire n_9565;
wire n_9566;
wire n_9567;
wire n_9568;
wire n_9569;
wire n_9570;
wire n_9571;
wire n_9572;
wire n_9573;
wire n_9574;
wire n_9575;
wire n_9576;
wire n_9577;
wire n_9578;
wire n_9579;
wire n_9580;
wire n_9581;
wire n_9582;
wire n_9583;
wire n_9584;
wire n_9585;
wire n_9586;
wire n_9587;
wire n_9588;
wire n_9589;
wire n_9590;
wire n_9591;
wire n_9592;
wire n_9593;
wire n_9594;
wire n_9595;
wire n_9596;
wire n_9597;
wire n_9598;
wire n_9599;
wire n_9600;
wire n_9601;
wire n_9602;
wire n_9603;
wire n_9604;
wire n_9605;
wire n_9606;
wire n_9607;
wire n_9608;
wire n_9609;
wire n_9610;
wire n_9611;
wire n_9612;
wire n_9613;
wire n_9614;
wire n_9615;
wire n_9616;
wire n_9617;
wire n_9618;
wire n_9619;
wire n_9620;
wire n_9621;
wire n_9622;
wire n_9623;
wire n_9624;
wire n_9625;
wire n_9626;
wire n_9627;
wire n_9628;
wire n_9629;
wire n_9630;
wire n_9631;
wire n_9632;
wire n_9633;
wire n_9634;
wire n_9635;
wire n_9636;
wire n_9637;
wire n_9638;
wire n_9639;
wire n_9640;
wire n_9641;
wire n_9642;
wire n_9643;
wire n_9644;
wire n_9645;
wire n_9646;
wire n_9647;
wire n_9648;
wire n_9649;
wire n_9650;
wire n_9651;
wire n_9652;
wire n_9653;
wire n_9654;
wire n_9655;
wire n_9656;
wire n_9657;
wire n_9658;
wire n_9659;
wire n_9660;
wire n_9661;
wire n_9662;
wire n_9663;
wire n_9664;
wire n_9665;
wire n_9666;
wire n_9667;
wire n_9668;
wire n_9669;
wire n_9670;
wire n_9671;
wire n_9672;
wire n_9673;
wire n_9674;
wire n_9675;
wire n_9676;
wire n_9677;
wire n_9678;
wire n_9679;
wire n_9680;
wire n_9681;
wire n_9682;
wire n_9683;
wire n_9684;
wire n_9685;
wire n_9686;
wire n_9687;
wire n_9688;
wire n_9689;
wire n_9690;
wire n_9691;
wire n_9692;
wire n_9693;
wire n_9694;
wire n_9695;
wire n_9696;
wire n_9697;
wire n_9698;
wire n_9699;
wire n_9700;
wire n_9701;
wire n_9702;
wire n_9703;
wire n_9704;
wire n_9705;
wire n_9706;
wire n_9707;
wire n_9708;
wire n_9709;
wire n_9710;
wire n_9711;
wire n_9712;
wire n_9713;
wire n_9714;
wire n_9715;
wire n_9716;
wire n_9717;
wire n_9718;
wire n_9719;
wire n_9720;
wire n_9721;
wire n_9722;
wire n_9723;
wire n_9724;
wire n_9725;
wire n_9726;
wire n_9727;
wire n_9728;
wire n_9729;
wire n_9730;
wire n_9731;
wire n_9732;
wire n_9733;
wire n_9734;
wire n_9735;
wire n_9736;
wire n_9737;
wire n_9738;
wire n_9739;
wire n_9740;
wire n_9741;
wire n_9742;
wire n_9743;
wire n_9744;
wire n_9745;
wire n_9746;
wire n_9747;
wire n_9748;
wire n_9749;
wire n_9750;
wire n_9751;
wire n_9752;
wire n_9753;
wire n_9754;
wire n_9755;
wire n_9756;
wire n_9757;
wire n_9758;
wire n_9759;
wire n_9760;
wire n_9761;
wire n_9762;
wire n_9763;
wire n_9764;
wire n_9765;
wire n_9766;
wire n_9767;
wire n_9768;
wire n_9769;
wire n_9770;
wire n_9771;
wire n_9772;
wire n_9773;
wire n_9774;
wire n_9775;
wire n_9776;
wire n_9777;
wire n_9778;
wire n_9779;
wire n_9780;
wire n_9781;
wire n_9782;
wire n_9783;
wire n_9784;
wire n_9785;
wire n_9786;
wire n_9787;
wire n_9788;
wire n_9789;
wire n_9790;
wire n_9791;
wire n_9792;
wire n_9793;
wire n_9794;
wire n_9795;
wire n_9796;
wire n_9797;
wire n_9798;
wire n_9799;
wire n_9800;
wire n_9801;
wire n_9802;
wire n_9803;
wire n_9804;
wire n_9805;
wire n_9806;
wire n_9807;
wire n_9808;
wire n_9809;
wire n_9810;
wire n_9811;
wire n_9812;
wire n_9813;
wire n_9814;
wire n_9815;
wire n_9816;
wire n_9817;
wire n_9818;
wire n_9819;
wire n_9820;
wire n_9821;
wire n_9822;
wire n_9823;
wire n_9824;
wire n_9825;
wire n_9826;
wire n_9827;
wire n_9828;
wire n_9829;
wire n_9830;
wire n_9831;
wire n_9832;
wire n_9833;
wire n_9834;
wire n_9835;
wire n_9836;
wire n_9837;
wire n_9838;
wire n_9839;
wire n_9840;
wire n_9841;
wire n_9842;
wire n_9843;
wire n_9844;
wire n_9845;
wire n_9846;
wire n_9847;
wire n_9848;
wire n_9849;
wire n_9850;
wire n_9851;
wire n_9852;
wire n_9853;
wire n_9854;
wire n_9855;
wire n_9856;
wire n_9857;
wire n_9858;
wire n_9859;
wire n_9860;
wire n_9861;
wire n_9862;
wire n_9863;
wire n_9864;
wire n_9865;
wire n_9866;
wire n_9867;
wire n_9868;
wire n_9869;
wire n_9870;
wire n_9871;
wire n_9872;
wire n_9873;
wire n_9874;
wire n_9875;
wire n_9876;
wire n_9877;
wire n_9878;
wire n_9879;
wire n_9880;
wire n_9881;
wire n_9882;
wire n_9883;
wire n_9884;
wire n_9885;
wire n_9886;
wire n_9887;
wire n_9888;
wire n_9889;
wire n_9890;
wire n_9891;
wire n_9892;
wire n_9893;
wire n_9894;
wire n_9895;
wire n_9896;
wire n_9897;
wire n_9898;
wire n_9899;
wire n_9900;
wire n_9901;
wire n_9902;
wire n_9903;
wire n_9904;
wire n_9905;
wire n_9906;
wire n_9907;
wire n_9908;
wire n_9909;
wire n_9910;
wire n_9911;
wire n_9912;
wire n_9913;
wire n_9914;
wire n_9915;
wire n_9916;
wire n_9917;
wire n_9918;
wire n_9919;
wire n_9920;
wire n_9921;
wire n_9922;
wire n_9923;
wire n_9924;
wire n_9925;
wire n_9926;
wire n_9927;
wire n_9928;
wire n_9929;
wire n_9930;
wire n_9931;
wire n_9932;
wire n_9933;
wire n_9934;
wire n_9935;
wire n_9936;
wire n_9937;
wire n_9938;
wire n_9939;
wire n_9940;
wire n_9941;
wire n_9942;
wire n_9943;
wire n_9944;
wire n_9945;
wire n_9946;
wire n_9947;
wire n_9948;
wire n_9949;
wire n_9950;
wire n_9951;
wire n_9952;
wire n_9953;
wire n_9954;
wire n_9955;
wire n_9956;
wire n_9957;
wire n_9958;
wire n_9959;
wire n_9960;
wire n_9961;
wire n_9962;
wire n_9963;
wire n_9964;
wire n_9965;
wire n_9966;
wire n_9967;
wire n_9968;
wire n_9969;
wire n_9970;
wire n_9971;
wire n_9972;
wire n_9973;
wire n_9974;
wire n_9975;
wire n_9976;
wire n_9977;
wire n_9978;
wire n_9979;
wire n_9980;
wire n_9981;
wire n_9982;
wire n_9983;
wire n_9984;
wire n_9985;
wire n_9986;
wire n_9987;
wire n_9988;
wire n_9989;
wire n_9990;
wire n_9991;
wire n_9992;
wire n_9993;
wire n_9994;
wire n_9995;
wire n_9996;
wire n_9997;
wire n_9998;
wire n_9999;
wire n_10000;
wire n_10001;
wire n_10002;
wire n_10003;
wire n_10004;
wire n_10005;
wire n_10006;
wire n_10007;
wire n_10008;
wire n_10009;
wire n_10010;
wire n_10011;
wire n_10012;
wire n_10013;
wire n_10014;
wire n_10015;
wire n_10016;
wire n_10017;
wire n_10018;
wire n_10019;
wire n_10020;
wire n_10021;
wire n_10022;
wire n_10023;
wire n_10024;
wire n_10025;
wire n_10026;
wire n_10027;
wire n_10028;
wire n_10029;
wire n_10030;
wire n_10031;
wire n_10032;
wire n_10033;
wire n_10034;
wire n_10035;
wire n_10036;
wire n_10037;
wire n_10038;
wire n_10039;
wire n_10040;
wire n_10041;
wire n_10042;
wire n_10043;
wire n_10044;
wire n_10045;
wire n_10046;
wire n_10047;
wire n_10048;
wire n_10049;
wire n_10050;
wire n_10051;
wire n_10052;
wire n_10053;
wire n_10054;
wire n_10055;
wire n_10056;
wire n_10057;
wire n_10058;
wire n_10059;
wire n_10060;
wire n_10061;
wire n_10062;
wire n_10063;
wire n_10064;
wire n_10065;
wire n_10066;
wire n_10067;
wire n_10068;
wire n_10069;
wire n_10070;
wire n_10071;
wire n_10072;
wire n_10073;
wire n_10074;
wire n_10075;
wire n_10076;
wire n_10077;
wire n_10078;
wire n_10079;
wire n_10080;
wire n_10081;
wire n_10082;
wire n_10083;
wire n_10084;
wire n_10085;
wire n_10086;
wire n_10087;
wire n_10088;
wire n_10089;
wire n_10090;
wire n_10091;
wire n_10092;
wire n_10093;
wire n_10094;
wire n_10095;
wire n_10096;
wire n_10097;
wire n_10098;
wire n_10099;
wire n_10100;
wire n_10101;
wire n_10102;
wire n_10103;
wire n_10104;
wire n_10105;
wire n_10106;
wire n_10107;
wire n_10108;
wire n_10109;
wire n_10110;
wire n_10111;
wire n_10112;
wire n_10113;
wire n_10114;
wire n_10115;
wire n_10116;
wire n_10117;
wire n_10118;
wire n_10119;
wire n_10120;
wire n_10121;
wire n_10122;
wire n_10123;
wire n_10124;
wire n_10125;
wire n_10126;
wire n_10127;
wire n_10128;
wire n_10129;
wire n_10130;
wire n_10131;
wire n_10132;
wire n_10133;
wire n_10134;
wire n_10135;
wire n_10136;
wire n_10137;
wire n_10138;
wire n_10139;
wire n_10140;
wire n_10141;
wire n_10142;
wire n_10143;
wire n_10144;
wire n_10145;
wire n_10146;
wire n_10147;
wire n_10148;
wire n_10149;
wire n_10150;
wire n_10151;
wire n_10152;
wire n_10153;
wire n_10154;
wire n_10155;
wire n_10156;
wire n_10157;
wire n_10158;
wire n_10159;
wire n_10160;
wire n_10161;
wire n_10162;
wire n_10163;
wire n_10164;
wire n_10165;
wire n_10166;
wire n_10167;
wire n_10168;
wire n_10169;
wire n_10170;
wire n_10171;
wire n_10172;
wire n_10173;
wire n_10174;
wire n_10175;
wire n_10176;
wire n_10177;
wire n_10178;
wire n_10179;
wire n_10180;
wire n_10181;
wire n_10182;
wire n_10183;
wire n_10184;
wire n_10185;
wire n_10186;
wire n_10187;
wire n_10188;
wire n_10189;
wire n_10190;
wire n_10191;
wire n_10192;
wire n_10193;
wire n_10194;
wire n_10195;
wire n_10196;
wire n_10197;
wire n_10198;
wire n_10199;
wire n_10200;
wire n_10201;
wire n_10202;
wire n_10203;
wire n_10204;
wire n_10205;
wire n_10206;
wire n_10207;
wire n_10208;
wire n_10209;
wire n_10210;
wire n_10211;
wire n_10212;
wire n_10213;
wire n_10214;
wire n_10215;
wire n_10216;
wire n_10217;
wire n_10218;
wire n_10219;
wire n_10220;
wire n_10221;
wire n_10222;
wire n_10223;
wire n_10224;
wire n_10225;
wire n_10226;
wire n_10227;
wire n_10228;
wire n_10229;
wire n_10230;
wire n_10231;
wire n_10232;
wire n_10233;
wire n_10234;
wire n_10235;
wire n_10236;
wire n_10237;
wire n_10238;
wire n_10239;
wire n_10240;
wire n_10241;
wire n_10242;
wire n_10243;
wire n_10244;
wire n_10245;
wire n_10246;
wire n_10247;
wire n_10248;
wire n_10249;
wire n_10250;
wire n_10251;
wire n_10252;
wire n_10253;
wire n_10254;
wire n_10255;
wire n_10256;
wire n_10257;
wire n_10258;
wire n_10259;
wire n_10260;
wire n_10261;
wire n_10262;
wire n_10263;
wire n_10264;
wire n_10265;
wire n_10266;
wire n_10267;
wire n_10268;
wire n_10269;
wire n_10270;
wire n_10271;
wire n_10272;
wire n_10273;
wire n_10274;
wire n_10275;
wire n_10276;
wire n_10277;
wire n_10278;
wire n_10279;
wire n_10280;
wire n_10281;
wire n_10282;
wire n_10283;
wire n_10284;
wire n_10285;
wire n_10286;
wire n_10287;
wire n_10288;
wire n_10289;
wire n_10290;
wire n_10291;
wire n_10292;
wire n_10293;
wire n_10294;
wire n_10295;
wire n_10296;
wire n_10297;
wire n_10298;
wire n_10299;
wire n_10300;
wire n_10301;
wire n_10302;
wire n_10303;
wire n_10304;
wire n_10305;
wire n_10306;
wire n_10307;
wire n_10308;
wire n_10309;
wire n_10310;
wire n_10311;
wire n_10312;
wire n_10313;
wire n_10314;
wire n_10315;
wire n_10316;
wire n_10317;
wire n_10318;
wire n_10319;
wire n_10320;
wire n_10321;
wire n_10322;
wire n_10323;
wire n_10324;
wire n_10325;
wire n_10326;
wire n_10327;
wire n_10328;
wire n_10329;
wire n_10330;
wire n_10331;
wire n_10332;
wire n_10333;
wire n_10334;
wire n_10335;
wire n_10336;
wire n_10337;
wire n_10338;
wire n_10339;
wire n_10340;
wire n_10341;
wire n_10342;
wire n_10343;
wire n_10344;
wire n_10345;
wire n_10346;
wire n_10347;
wire n_10348;
wire n_10349;
wire n_10350;
wire n_10351;
wire n_10352;
wire n_10353;
wire n_10354;
wire n_10355;
wire n_10356;
wire n_10357;
wire n_10358;
wire n_10359;
wire n_10360;
wire n_10361;
wire n_10362;
wire n_10363;
wire n_10364;
wire n_10365;
wire n_10366;
wire n_10367;
wire n_10368;
wire n_10369;
wire n_10370;
wire n_10371;
wire n_10372;
wire n_10373;
wire n_10374;
wire n_10375;
wire n_10376;
wire n_10377;
wire n_10378;
wire n_10379;
wire n_10380;
wire n_10381;
wire n_10382;
wire n_10383;
wire n_10384;
wire n_10385;
wire n_10386;
wire n_10387;
wire n_10388;
wire n_10389;
wire n_10390;
wire n_10391;
wire n_10392;
wire n_10393;
wire n_10394;
wire n_10395;
wire n_10396;
wire n_10397;
wire n_10398;
wire n_10399;
wire n_10400;
wire n_10401;
wire n_10402;
wire n_10403;
wire n_10404;
wire n_10405;
wire n_10406;
wire n_10407;
wire n_10408;
wire n_10409;
wire n_10410;
wire n_10411;
wire n_10412;
wire n_10413;
wire n_10414;
wire n_10415;
wire n_10416;
wire n_10417;
wire n_10418;
wire n_10419;
wire n_10420;
wire n_10421;
wire n_10422;
wire n_10423;
wire n_10424;
wire n_10425;
wire n_10426;
wire n_10427;
wire n_10428;
wire n_10429;
wire n_10430;
wire n_10431;
wire n_10432;
wire n_10433;
wire n_10434;
wire n_10435;
wire n_10436;
wire n_10437;
wire n_10438;
wire n_10439;
wire n_10440;
wire n_10441;
wire n_10442;
wire n_10443;
wire n_10444;
wire n_10445;
wire n_10446;
wire n_10447;
wire n_10448;
wire n_10449;
wire n_10450;
wire n_10451;
wire n_10452;
wire n_10453;
wire n_10454;
wire n_10455;
wire n_10456;
wire n_10457;
wire n_10458;
wire n_10459;
wire n_10460;
wire n_10461;
wire n_10462;
wire n_10463;
wire n_10464;
wire n_10465;
wire n_10466;
wire n_10467;
wire n_10468;
wire n_10469;
wire n_10470;
wire n_10471;
wire n_10472;
wire n_10473;
wire n_10474;
wire n_10475;
wire n_10476;
wire n_10477;
wire n_10478;
wire n_10479;
wire n_10480;
wire n_10481;
wire n_10482;
wire n_10483;
wire n_10484;
wire n_10485;
wire n_10486;
wire n_10487;
wire n_10488;
wire n_10489;
wire n_10490;
wire n_10491;
wire n_10492;
wire n_10493;
wire n_10494;
wire n_10495;
wire n_10496;
wire n_10497;
wire n_10498;
wire n_10499;
wire n_10500;
wire n_10501;
wire n_10502;
wire n_10503;
wire n_10504;
wire n_10505;
wire n_10506;
wire n_10507;
wire n_10508;
wire n_10509;
wire n_10510;
wire n_10511;
wire n_10512;
wire n_10513;
wire n_10514;
wire n_10515;
wire n_10516;
wire n_10517;
wire n_10518;
wire n_10519;
wire n_10520;
wire n_10521;
wire n_10522;
wire n_10523;
wire n_10524;
wire n_10525;
wire n_10526;
wire n_10527;
wire n_10528;
wire n_10529;
wire n_10530;
wire n_10531;
wire n_10532;
wire n_10533;
wire n_10534;
wire n_10535;
wire n_10536;
wire n_10537;
wire n_10538;
wire n_10539;
wire n_10540;
wire n_10541;
wire n_10542;
wire n_10543;
wire n_10544;
wire n_10545;
wire n_10546;
wire n_10547;
wire n_10548;
wire n_10549;
wire n_10550;
wire n_10551;
wire n_10552;
wire n_10553;
wire n_10554;
wire n_10555;
wire n_10556;
wire n_10557;
wire n_10558;
wire n_10559;
wire n_10560;
wire n_10561;
wire n_10562;
wire n_10563;
wire n_10564;
wire n_10565;
wire n_10566;
wire n_10567;
wire n_10568;
wire n_10569;
wire n_10570;
wire n_10571;
wire n_10572;
wire n_10573;
wire n_10574;
wire n_10575;
wire n_10576;
wire n_10577;
wire n_10578;
wire n_10579;
wire n_10580;
wire n_10581;
wire n_10582;
wire n_10583;
wire n_10584;
wire n_10585;
wire n_10586;
wire n_10587;
wire n_10588;
wire n_10589;
wire n_10590;
wire n_10591;
wire n_10592;
wire n_10593;
wire n_10594;
wire n_10595;
wire n_10596;
wire n_10597;
wire n_10598;
wire n_10599;
wire n_10600;
wire n_10601;
wire n_10602;
wire n_10603;
wire n_10604;
wire n_10605;
wire n_10606;
wire n_10607;
wire n_10608;
wire n_10609;
wire n_10610;
wire n_10611;
wire n_10612;
wire n_10613;
wire n_10614;
wire n_10615;
wire n_10616;
wire n_10617;
wire n_10618;
wire n_10619;
wire n_10620;
wire n_10621;
wire n_10622;
wire n_10623;
wire n_10624;
wire n_10625;
wire n_10626;
wire n_10627;
wire n_10628;
wire n_10629;
wire n_10630;
wire n_10631;
wire n_10632;
wire n_10633;
wire n_10634;
wire n_10635;
wire n_10636;
wire n_10637;
wire n_10638;
wire n_10639;
wire n_10640;
wire n_10641;
wire n_10642;
wire n_10643;
wire n_10644;
wire n_10645;
wire n_10646;
wire n_10647;
wire n_10648;
wire n_10649;
wire n_10650;
wire n_10651;
wire n_10652;
wire n_10653;
wire n_10654;
wire n_10655;
wire n_10656;
wire n_10657;
wire n_10658;
wire n_10659;
wire n_10660;
wire n_10661;
wire n_10662;
wire n_10663;
wire n_10664;
wire n_10665;
wire n_10666;
wire n_10667;
wire n_10668;
wire n_10669;
wire n_10670;
wire n_10671;
wire n_10672;
wire n_10673;
wire n_10674;
wire n_10675;
wire n_10676;
wire n_10677;
wire n_10678;
wire n_10679;
wire n_10680;
wire n_10681;
wire n_10682;
wire n_10683;
wire n_10684;
wire n_10685;
wire n_10686;
wire n_10687;
wire n_10688;
wire n_10689;
wire n_10690;
wire n_10691;
wire n_10692;
wire n_10693;
wire n_10694;
wire n_10695;
wire n_10696;
wire n_10697;
wire n_10698;
wire n_10699;
wire n_10700;
wire n_10701;
wire n_10702;
wire n_10703;
wire n_10704;
wire n_10705;
wire n_10706;
wire n_10707;
wire n_10708;
wire n_10709;
wire n_10710;
wire n_10711;
wire n_10712;
wire n_10713;
wire n_10714;
wire n_10715;
wire n_10716;
wire n_10717;
wire n_10718;
wire n_10719;
wire n_10720;
wire n_10721;
wire n_10722;
wire n_10723;
wire n_10724;
wire n_10725;
wire n_10726;
wire n_10727;
wire n_10728;
wire n_10729;
wire n_10730;
wire n_10731;
wire n_10732;
wire n_10733;
wire n_10734;
wire n_10735;
wire n_10736;
wire n_10737;
wire n_10738;
wire n_10739;
wire n_10740;
wire n_10741;
wire n_10742;
wire n_10743;
wire n_10744;
wire n_10745;
wire n_10746;
wire n_10747;
wire n_10748;
wire n_10749;
wire n_10750;
wire n_10751;
wire n_10752;
wire n_10753;
wire n_10754;
wire n_10755;
wire n_10756;
wire n_10757;
wire n_10758;
wire n_10759;
wire n_10760;
wire n_10761;
wire n_10762;
wire n_10763;
wire n_10764;
wire n_10765;
wire n_10766;
wire n_10767;
wire n_10768;
wire n_10769;
wire n_10770;
wire n_10771;
wire n_10772;
wire n_10773;
wire n_10774;
wire n_10775;
wire n_10776;
wire n_10777;
wire n_10778;
wire n_10779;
wire n_10780;
wire n_10781;
wire n_10782;
wire n_10783;
wire n_10784;
wire n_10785;
wire n_10786;
wire n_10787;
wire n_10788;
wire n_10789;
wire n_10790;
wire n_10791;
wire n_10792;
wire n_10793;
wire n_10794;
wire n_10795;
wire n_10796;
wire n_10797;
wire n_10798;
wire n_10799;
wire n_10800;
wire n_10801;
wire n_10802;
wire n_10803;
wire n_10804;
wire n_10805;
wire n_10806;
wire n_10807;
wire n_10808;
wire n_10809;
wire n_10810;
wire n_10811;
wire n_10812;
wire n_10813;
wire n_10814;
wire n_10815;
wire n_10816;
wire n_10817;
wire n_10818;
wire n_10819;
wire n_10820;
wire n_10821;
wire n_10822;
wire n_10823;
wire n_10824;
wire n_10825;
wire n_10826;
wire n_10827;
wire n_10828;
wire n_10829;
wire n_10830;
wire n_10831;
wire n_10832;
wire n_10833;
wire n_10834;
wire n_10835;
wire n_10836;
wire n_10837;
wire n_10838;
wire n_10839;
wire n_10840;
wire n_10841;
wire n_10842;
wire n_10843;
wire n_10844;
wire n_10845;
wire n_10846;
wire n_10847;
wire n_10848;
wire n_10849;
wire n_10850;
wire n_10851;
wire n_10852;
wire n_10853;
wire n_10854;
wire n_10855;
wire n_10856;
wire n_10857;
wire n_10858;
wire n_10859;
wire n_10860;
wire n_10861;
wire n_10862;
wire n_10863;
wire n_10864;
wire n_10865;
wire n_10866;
wire n_10867;
wire n_10868;
wire n_10869;
wire n_10870;
wire n_10871;
wire n_10872;
wire n_10873;
wire n_10874;
wire n_10875;
wire n_10876;
wire n_10877;
wire n_10878;
wire n_10879;
wire n_10880;
wire n_10881;
wire n_10882;
wire n_10883;
wire n_10884;
wire n_10885;
wire n_10886;
wire n_10887;
wire n_10888;
wire n_10889;
wire n_10890;
wire n_10891;
wire n_10892;
wire n_10893;
wire n_10894;
wire n_10895;
wire n_10896;
wire n_10897;
wire n_10898;
wire n_10899;
wire n_10900;
wire n_10901;
wire n_10902;
wire n_10903;
wire n_10904;
wire n_10905;
wire n_10906;
wire n_10907;
wire n_10908;
wire n_10909;
wire n_10910;
wire n_10911;
wire n_10912;
wire n_10913;
wire n_10914;
wire n_10915;
wire n_10916;
wire n_10917;
wire n_10918;
wire n_10919;
wire n_10920;
wire n_10921;
wire n_10922;
wire n_10923;
wire n_10924;
wire n_10925;
wire n_10926;
wire n_10927;
wire n_10928;
wire n_10929;
wire n_10930;
wire n_10931;
wire n_10932;
wire n_10933;
wire n_10934;
wire n_10935;
wire n_10936;
wire n_10937;
wire n_10938;
wire n_10939;
wire n_10940;
wire n_10941;
wire n_10942;
wire n_10943;
wire n_10944;
wire n_10945;
wire n_10946;
wire n_10947;
wire n_10948;
wire n_10949;
wire n_10950;
wire n_10951;
wire n_10952;
wire n_10953;
wire n_10954;
wire n_10955;
wire n_10956;
wire n_10957;
wire n_10958;
wire n_10959;
wire n_10960;
wire n_10961;
wire n_10962;
wire n_10963;
wire n_10964;
wire n_10965;
wire n_10966;
wire n_10967;
wire n_10968;
wire n_10969;
wire n_10970;
wire n_10971;
wire n_10972;
wire n_10973;
wire n_10974;
wire n_10975;
wire n_10976;
wire n_10977;
wire n_10978;
wire n_10979;
wire n_10980;
wire n_10981;
wire n_10982;
wire n_10983;
wire n_10984;
wire n_10985;
wire n_10986;
wire n_10987;
wire n_10988;
wire n_10989;
wire n_10990;
wire n_10991;
wire n_10992;
wire n_10993;
wire n_10994;
wire n_10995;
wire n_10996;
wire n_10997;
wire n_10998;
wire n_10999;
wire n_11000;
wire n_11001;
wire n_11002;
wire n_11003;
wire n_11004;
wire n_11005;
wire n_11006;
wire n_11007;
wire n_11008;
wire n_11009;
wire n_11010;
wire n_11011;
wire n_11012;
wire n_11013;
wire n_11014;
wire n_11015;
wire n_11016;
wire n_11017;
wire n_11018;
wire n_11019;
wire n_11020;
wire n_11021;
wire n_11022;
wire n_11023;
wire n_11024;
wire n_11025;
wire n_11026;
wire n_11027;
wire n_11028;
wire n_11029;
wire n_11030;
wire n_11031;
wire n_11032;
wire n_11033;
wire n_11034;
wire n_11035;
wire n_11036;
wire n_11037;
wire n_11038;
wire n_11039;
wire n_11040;
wire n_11041;
wire n_11042;
wire n_11043;
wire n_11044;
wire n_11045;
wire n_11046;
wire n_11047;
wire n_11048;
wire n_11049;
wire n_11050;
wire n_11051;
wire n_11052;
wire n_11053;
wire n_11054;
wire n_11055;
wire n_11056;
wire n_11057;
wire n_11058;
wire n_11059;
wire n_11060;
wire n_11061;
wire n_11062;
wire n_11063;
wire n_11064;
wire n_11065;
wire n_11066;
wire n_11067;
wire n_11068;
wire n_11069;
wire n_11070;
wire n_11071;
wire n_11072;
wire n_11073;
wire n_11074;
wire n_11075;
wire n_11076;
wire n_11077;
wire n_11078;
wire n_11079;
wire n_11080;
wire n_11081;
wire n_11082;
wire n_11083;
wire n_11084;
wire n_11085;
wire n_11086;
wire n_11087;
wire n_11088;
wire n_11089;
wire n_11090;
wire n_11091;
wire n_11092;
wire n_11093;
wire n_11094;
wire n_11095;
wire n_11096;
wire n_11097;
wire n_11098;
wire n_11099;
wire n_11100;
wire n_11101;
wire n_11102;
wire n_11103;
wire n_11104;
wire n_11105;
wire n_11106;
wire n_11107;
wire n_11108;
wire n_11109;
wire n_11110;
wire n_11111;
wire n_11112;
wire n_11113;
wire n_11114;
wire n_11115;
wire n_11116;
wire n_11117;
wire n_11118;
wire n_11119;
wire n_11120;
wire n_11121;
wire n_11122;
wire n_11123;
wire n_11124;
wire n_11125;
wire n_11126;
wire n_11127;
wire n_11128;
wire n_11129;
wire n_11130;
wire n_11131;
wire n_11132;
wire n_11133;
wire n_11134;
wire n_11135;
wire n_11136;
wire n_11137;
wire n_11138;
wire n_11139;
wire n_11140;
wire n_11141;
wire n_11142;
wire n_11143;
wire n_11144;
wire n_11145;
wire n_11146;
wire n_11147;
wire n_11148;
wire n_11149;
wire n_11150;
wire n_11151;
wire n_11152;
wire n_11153;
wire n_11154;
wire n_11155;
wire n_11156;
wire n_11157;
wire n_11158;
wire n_11159;
wire n_11160;
wire n_11161;
wire n_11162;
wire n_11163;
wire n_11164;
wire n_11165;
wire n_11166;
wire n_11167;
wire n_11168;
wire n_11169;
wire n_11170;
wire n_11171;
wire n_11172;
wire n_11173;
wire n_11174;
wire n_11175;
wire n_11176;
wire n_11177;
wire n_11178;
wire n_11179;
wire n_11180;
wire n_11181;
wire n_11182;
wire n_11183;
wire n_11184;
wire n_11185;
wire n_11186;
wire n_11187;
wire n_11188;
wire n_11189;
wire n_11190;
wire n_11191;
wire n_11192;
wire n_11193;
wire n_11194;
wire n_11195;
wire n_11196;
wire n_11197;
wire n_11198;
wire n_11199;
wire n_11200;
wire n_11201;
wire n_11202;
wire n_11203;
wire n_11204;
wire n_11205;
wire n_11206;
wire n_11207;
wire n_11208;
wire n_11209;
wire n_11210;
wire n_11211;
wire n_11212;
wire n_11213;
wire n_11214;
wire n_11215;
wire n_11216;
wire n_11217;
wire n_11218;
wire n_11219;
wire n_11220;
wire n_11221;
wire n_11222;
wire n_11223;
wire n_11224;
wire n_11225;
wire n_11226;
wire n_11227;
wire n_11228;
wire n_11229;
wire n_11230;
wire n_11231;
wire n_11232;
wire n_11233;
wire n_11234;
wire n_11235;
wire n_11236;
wire n_11237;
wire n_11238;
wire n_11239;
wire n_11240;
wire n_11241;
wire n_11242;
wire n_11243;
wire n_11244;
wire n_11245;
wire n_11246;
wire n_11247;
wire n_11248;
wire n_11249;
wire n_11250;
wire n_11251;
wire n_11252;
wire n_11253;
wire n_11254;
wire n_11255;
wire n_11256;
wire n_11257;
wire n_11258;
wire n_11259;
wire n_11260;
wire n_11261;
wire n_11262;
wire n_11263;
wire n_11264;
wire n_11265;
wire n_11266;
wire n_11267;
wire n_11268;
wire n_11269;
wire n_11270;
wire n_11271;
wire n_11272;
wire n_11273;
wire n_11274;
wire n_11275;
wire n_11276;
wire n_11277;
wire n_11278;
wire n_11279;
wire n_11280;
wire n_11281;
wire n_11282;
wire n_11283;
wire n_11284;
wire n_11285;
wire n_11286;
wire n_11287;
wire n_11288;
wire n_11289;
wire n_11290;
wire n_11291;
wire n_11292;
wire n_11293;
wire n_11294;
wire n_11295;
wire n_11296;
wire n_11297;
wire n_11298;
wire n_11299;
wire n_11300;
wire n_11301;
wire n_11302;
wire n_11303;
wire n_11304;
wire n_11305;
wire n_11306;
wire n_11307;
wire n_11308;
wire n_11309;
wire n_11310;
wire n_11311;
wire n_11312;
wire n_11313;
wire n_11314;
wire n_11315;
wire n_11316;
wire n_11317;
wire n_11318;
wire n_11319;
wire n_11320;
wire n_11321;
wire n_11322;
wire n_11323;
wire n_11324;
wire n_11325;
wire n_11326;
wire n_11327;
wire n_11328;
wire n_11329;
wire n_11330;
wire n_11331;
wire n_11332;
wire n_11333;
wire n_11334;
wire n_11335;
wire n_11336;
wire n_11337;
wire n_11338;
wire n_11339;
wire n_11340;
wire n_11341;
wire n_11342;
wire n_11343;
wire n_11344;
wire n_11345;
wire n_11346;
wire n_11347;
wire n_11348;
wire n_11349;
wire n_11350;
wire n_11351;
wire n_11352;
wire n_11353;
wire n_11354;
wire n_11355;
wire n_11356;
wire n_11357;
wire n_11358;
wire n_11359;
wire n_11360;
wire n_11361;
wire n_11362;
wire n_11363;
wire n_11364;
wire n_11365;
wire n_11366;
wire n_11367;
wire n_11368;
wire n_11369;
wire n_11370;
wire n_11371;
wire n_11372;
wire n_11373;
wire n_11374;
wire n_11375;
wire n_11376;
wire n_11377;
wire n_11378;
wire n_11379;
wire n_11380;
wire n_11381;
wire n_11382;
wire n_11383;
wire n_11384;
wire n_11385;
wire n_11386;
wire n_11387;
wire n_11388;
wire n_11389;
wire n_11390;
wire n_11391;
wire n_11392;
wire n_11393;
wire n_11394;
wire n_11395;
wire n_11396;
wire n_11397;
wire n_11398;
wire n_11399;
wire n_11400;
wire n_11401;
wire n_11402;
wire n_11403;
wire n_11404;
wire n_11405;
wire n_11406;
wire n_11407;
wire n_11408;
wire n_11409;
wire n_11410;
wire n_11411;
wire n_11412;
wire n_11413;
wire n_11414;
wire n_11415;
wire n_11416;
wire n_11417;
wire n_11418;
wire n_11419;
wire n_11420;
wire n_11421;
wire n_11422;
wire n_11423;
wire n_11424;
wire n_11425;
wire n_11426;
wire n_11427;
wire n_11428;
wire n_11429;
wire n_11430;
wire n_11431;
wire n_11432;
wire n_11433;
wire n_11434;
wire n_11435;
wire n_11436;
wire n_11437;
wire n_11438;
wire n_11439;
wire n_11440;
wire n_11441;
wire n_11442;
wire n_11443;
wire n_11444;
wire n_11445;
wire n_11446;
wire n_11447;
wire n_11448;
wire n_11449;
wire n_11450;
wire n_11451;
wire n_11452;
wire n_11453;
wire n_11454;
wire n_11455;
wire n_11456;
wire n_11457;
wire n_11458;
wire n_11459;
wire n_11460;
wire n_11461;
wire n_11462;
wire n_11463;
wire n_11464;
wire n_11465;
wire n_11466;
wire n_11467;
wire n_11468;
wire n_11469;
wire n_11470;
wire n_11471;
wire n_11472;
wire n_11473;
wire n_11474;
wire n_11475;
wire n_11476;
wire n_11477;
wire n_11478;
wire n_11479;
wire n_11480;
wire n_11481;
wire n_11482;
wire n_11483;
wire n_11484;
wire n_11485;
wire n_11486;
wire n_11487;
wire n_11488;
wire n_11489;
wire n_11490;
wire n_11491;
wire n_11492;
wire n_11493;
wire n_11494;
wire n_11495;
wire n_11496;
wire n_11497;
wire n_11498;
wire n_11499;
wire n_11500;
wire n_11501;
wire n_11502;
wire n_11503;
wire n_11504;
wire n_11505;
wire n_11506;
wire n_11507;
wire n_11508;
wire n_11509;
wire n_11510;
wire n_11511;
wire n_11512;
wire n_11513;
wire n_11514;
wire n_11515;
wire n_11516;
wire n_11517;
wire n_11518;
wire n_11519;
wire n_11520;
wire n_11521;
wire n_11522;
wire n_11523;
wire n_11524;
wire n_11525;
wire n_11526;
wire n_11527;
wire n_11528;
wire n_11529;
wire n_11530;
wire n_11531;
wire n_11532;
wire n_11533;
wire n_11534;
wire n_11535;
wire n_11536;
wire n_11537;
wire n_11538;
wire n_11539;
wire n_11540;
wire n_11541;
wire n_11542;
wire n_11543;
wire n_11544;
wire n_11545;
wire n_11546;
wire n_11547;
wire n_11548;
wire n_11549;
wire n_11550;
wire n_11551;
wire n_11552;
wire n_11553;
wire n_11554;
wire n_11555;
wire n_11556;
wire n_11557;
wire n_11558;
wire n_11559;
wire n_11560;
wire n_11561;
wire n_11562;
wire n_11563;
wire n_11564;
wire n_11565;
wire n_11566;
wire n_11567;
wire n_11568;
wire n_11569;
wire n_11570;
wire n_11571;
wire n_11572;
wire n_11573;
wire n_11574;
wire n_11575;
wire n_11576;
wire n_11577;
wire n_11578;
wire n_11579;
wire n_11580;
wire n_11581;
wire n_11582;
wire n_11583;
wire n_11584;
wire n_11585;
wire n_11586;
wire n_11587;
wire n_11588;
wire n_11589;
wire n_11590;
wire n_11591;
wire n_11592;
wire n_11593;
wire n_11594;
wire n_11595;
wire n_11596;
wire n_11597;
wire n_11598;
wire n_11599;
wire n_11600;
wire n_11601;
wire n_11602;
wire n_11603;
wire n_11604;
wire n_11605;
wire n_11606;
wire n_11607;
wire n_11608;
wire n_11609;
wire n_11610;
wire n_11611;
wire n_11612;
wire n_11613;
wire n_11614;
wire n_11615;
wire n_11616;
wire n_11617;
wire n_11618;
wire n_11619;
wire n_11620;
wire n_11621;
wire n_11622;
wire n_11623;
wire n_11624;
wire n_11625;
wire n_11626;
wire n_11627;
wire n_11628;
wire n_11629;
wire n_11630;
wire n_11631;
wire n_11632;
wire n_11633;
wire n_11634;
wire n_11635;
wire n_11636;
wire n_11637;
wire n_11638;
wire n_11639;
wire n_11640;
wire n_11641;
wire n_11642;
wire n_11643;
wire n_11644;
wire n_11645;
wire n_11646;
wire n_11647;
wire n_11648;
wire n_11649;
wire n_11650;
wire n_11651;
wire n_11652;
wire n_11653;
wire n_11654;
wire n_11655;
wire n_11656;
wire n_11657;
wire n_11658;
wire n_11659;
wire n_11660;
wire n_11661;
wire n_11662;
wire n_11663;
wire n_11664;
wire n_11665;
wire n_11666;
wire n_11667;
wire n_11668;
wire n_11669;
wire n_11670;
wire n_11671;
wire n_11672;
wire n_11673;
wire n_11674;
wire n_11675;
wire n_11676;
wire n_11677;
wire n_11678;
wire n_11679;
wire n_11680;
wire n_11681;
wire n_11682;
wire n_11683;
wire n_11684;
wire n_11685;
wire n_11686;
wire n_11687;
wire n_11688;
wire n_11689;
wire n_11690;
wire n_11691;
wire n_11692;
wire n_11693;
wire n_11694;
wire n_11695;
wire n_11696;
wire n_11697;
wire n_11698;
wire n_11699;
wire n_11700;
wire n_11701;
wire n_11702;
wire n_11703;
wire n_11704;
wire n_11705;
wire n_11706;
wire n_11707;
wire n_11708;
wire n_11709;
wire n_11710;
wire n_11711;
wire n_11712;
wire n_11713;
wire n_11714;
wire n_11715;
wire n_11716;
wire n_11717;
wire n_11718;
wire n_11719;
wire n_11720;
wire n_11721;
wire n_11722;
wire n_11723;
wire n_11724;
wire n_11725;
wire n_11726;
wire n_11727;
wire n_11728;
wire n_11729;
wire n_11730;
wire n_11731;
wire n_11732;
wire n_11733;
wire n_11734;
wire n_11735;
wire n_11736;
wire n_11737;
wire n_11738;
wire n_11739;
wire n_11740;
wire n_11741;
wire n_11742;
wire n_11743;
wire n_11744;
wire n_11745;
wire n_11746;
wire n_11747;
wire n_11748;
wire n_11749;
wire n_11750;
wire n_11751;
wire n_11752;
wire n_11753;
wire n_11754;
wire n_11755;
wire n_11756;
wire n_11757;
wire n_11758;
wire n_11759;
wire n_11760;
wire n_11761;
wire n_11762;
wire n_11763;
wire n_11764;
wire n_11765;
wire n_11766;
wire n_11767;
wire n_11768;
wire n_11769;
wire n_11770;
wire n_11771;
wire n_11772;
wire n_11773;
wire n_11774;
wire n_11775;
wire n_11776;
wire n_11777;
wire n_11778;
wire n_11779;
wire n_11780;
wire n_11781;
wire n_11782;
wire n_11783;
wire n_11784;
wire n_11785;
wire n_11786;
wire n_11787;
wire n_11788;
wire n_11789;
wire n_11790;
wire n_11791;
wire n_11792;
wire n_11793;
wire n_11794;
wire n_11795;
wire n_11796;
wire n_11797;
wire n_11798;
wire n_11799;
wire n_11800;
wire n_11801;
wire n_11802;
wire n_11803;
wire n_11804;
wire n_11805;
wire n_11806;
wire n_11807;
wire n_11808;
wire n_11809;
wire n_11810;
wire n_11811;
wire n_11812;
wire n_11813;
wire n_11814;
wire n_11815;
wire n_11816;
wire n_11817;
wire n_11818;
wire n_11819;
wire n_11820;
wire n_11821;
wire n_11822;
wire n_11823;
wire n_11824;
wire n_11825;
wire n_11826;
wire n_11827;
wire n_11828;
wire n_11829;
wire n_11830;
wire n_11831;
wire n_11832;
wire n_11833;
wire n_11834;
wire n_11835;
wire n_11836;
wire n_11837;
wire n_11838;
wire n_11839;
wire n_11840;
wire n_11841;
wire n_11842;
wire n_11843;
wire n_11844;
wire n_11845;
wire n_11846;
wire n_11847;
wire n_11848;
wire n_11849;
wire n_11850;
wire n_11851;
wire n_11852;
wire n_11853;
wire n_11854;
wire n_11855;
wire n_11856;
wire n_11857;
wire n_11858;
wire n_11859;
wire n_11860;
wire n_11861;
wire n_11862;
wire n_11863;
wire n_11864;
wire n_11865;
wire n_11866;
wire n_11867;
wire n_11868;
wire n_11869;
wire n_11870;
wire n_11871;
wire n_11872;
wire n_11873;
wire n_11874;
wire n_11875;
wire n_11876;
wire n_11877;
wire n_11878;
wire n_11879;
wire n_11880;
wire n_11881;
wire n_11882;
wire n_11883;
wire n_11884;
wire n_11885;
wire n_11886;
wire n_11887;
wire n_11888;
wire n_11889;
wire n_11890;
wire n_11891;
wire n_11892;
wire n_11893;
wire n_11894;
wire n_11895;
wire n_11896;
wire n_11897;
wire n_11898;
wire n_11899;
wire n_11900;
wire n_11901;
wire n_11902;
wire n_11903;
wire n_11904;
wire n_11905;
wire n_11906;
wire n_11907;
wire n_11908;
wire n_11909;
wire n_11910;
wire n_11911;
wire n_11912;
wire n_11913;
wire n_11914;
wire n_11915;
wire n_11916;
wire n_11917;
wire n_11918;
wire n_11919;
wire n_11920;
wire n_11921;
wire n_11922;
wire n_11923;
wire n_11924;
wire n_11925;
wire n_11926;
wire n_11927;
wire n_11928;
wire n_11929;
wire n_11930;
wire n_11931;
wire n_11932;
wire n_11933;
wire n_11934;
wire n_11935;
wire n_11936;
wire n_11937;
wire n_11938;
wire n_11939;
wire n_11940;
wire n_11941;
wire n_11942;
wire n_11943;
wire n_11944;
wire n_11945;
wire n_11946;
wire n_11947;
wire n_11948;
wire n_11949;
wire n_11950;
wire n_11951;
wire n_11952;
wire n_11953;
wire n_11954;
wire n_11955;
wire n_11956;
wire n_11957;
wire n_11958;
wire n_11959;
wire n_11960;
wire n_11961;
wire n_11962;
wire n_11963;
wire n_11964;
wire n_11965;
wire n_11966;
wire n_11967;
wire n_11968;
wire n_11969;
wire n_11970;
wire n_11971;
wire n_11972;
wire n_11973;
wire n_11974;
wire n_11975;
wire n_11976;
wire n_11977;
wire n_11978;
wire n_11979;
wire n_11980;
wire n_11981;
wire n_11982;
wire n_11983;
wire n_11984;
wire n_11985;
wire n_11986;
wire n_11987;
wire n_11988;
wire n_11989;
wire n_11990;
wire n_11991;
wire n_11992;
wire n_11993;
wire n_11994;
wire n_11995;
wire n_11996;
wire n_11997;
wire n_11998;
wire n_11999;
wire n_12000;
wire n_12001;
wire n_12002;
wire n_12003;
wire n_12004;
wire n_12005;
wire n_12006;
wire n_12007;
wire n_12008;
wire n_12009;
wire n_12010;
wire n_12011;
wire n_12012;
wire n_12013;
wire n_12014;
wire n_12015;
wire n_12016;
wire n_12017;
wire n_12018;
wire n_12019;
wire n_12020;
wire n_12021;
wire n_12022;
wire n_12023;
wire n_12024;
wire n_12025;
wire n_12026;
wire n_12027;
wire n_12028;
wire n_12029;
wire n_12030;
wire n_12031;
wire n_12032;
wire n_12033;
wire n_12034;
wire n_12035;
wire n_12036;
wire n_12037;
wire n_12038;
wire n_12039;
wire n_12040;
wire n_12041;
wire n_12042;
wire n_12043;
wire n_12044;
wire n_12045;
wire n_12046;
wire n_12047;
wire n_12048;
wire n_12049;
wire n_12050;
wire n_12051;
wire n_12052;
wire n_12053;
wire n_12054;
wire n_12055;
wire n_12056;
wire n_12057;
wire n_12058;
wire n_12059;
wire n_12060;
wire n_12061;
wire n_12062;
wire n_12063;
wire n_12064;
wire n_12065;
wire n_12066;
wire n_12067;
wire n_12068;
wire n_12069;
wire n_12070;
wire n_12071;
wire n_12072;
wire n_12073;
wire n_12074;
wire n_12075;
wire n_12076;
wire n_12077;
wire n_12078;
wire n_12079;
wire n_12080;
wire n_12081;
wire n_12082;
wire n_12083;
wire n_12084;
wire n_12085;
wire n_12086;
wire n_12087;
wire n_12088;
wire n_12089;
wire n_12090;
wire n_12091;
wire n_12092;
wire n_12093;
wire n_12094;
wire n_12095;
wire n_12096;
wire n_12097;
wire n_12098;
wire n_12099;
wire n_12100;
wire n_12101;
wire n_12102;
wire n_12103;
wire n_12104;
wire n_12105;
wire n_12106;
wire n_12107;
wire n_12108;
wire n_12109;
wire n_12110;
wire n_12111;
wire n_12112;
wire n_12113;
wire n_12114;
wire n_12115;
wire n_12116;
wire n_12117;
wire n_12118;
wire n_12119;
wire n_12120;
wire n_12121;
wire n_12122;
wire n_12123;
wire n_12124;
wire n_12125;
wire n_12126;
wire n_12127;
wire n_12128;
wire n_12129;
wire n_12130;
wire n_12131;
wire n_12132;
wire n_12133;
wire n_12134;
wire n_12135;
wire n_12136;
wire n_12137;
wire n_12138;
wire n_12139;
wire n_12140;
wire n_12141;
wire n_12142;
wire n_12143;
wire n_12144;
wire n_12145;
wire n_12146;
wire n_12147;
wire n_12148;
wire n_12149;
wire n_12150;
wire n_12151;
wire n_12152;
wire n_12153;
wire n_12154;
wire n_12155;
wire n_12156;
wire n_12157;
wire n_12158;
wire n_12159;
wire n_12160;
wire n_12161;
wire n_12162;
wire n_12163;
wire n_12164;
wire n_12165;
wire n_12166;
wire n_12167;
wire n_12168;
wire n_12169;
wire n_12170;
wire n_12171;
wire n_12172;
wire n_12173;
wire n_12174;
wire n_12175;
wire n_12176;
wire n_12177;
wire n_12178;
wire n_12179;
wire n_12180;
wire n_12181;
wire n_12182;
wire n_12183;
wire n_12184;
wire n_12185;
wire n_12186;
wire n_12187;
wire n_12188;
wire n_12189;
wire n_12190;
wire n_12191;
wire n_12192;
wire n_12193;
wire n_12194;
wire n_12195;
wire n_12196;
wire n_12197;
wire n_12198;
wire n_12199;
wire n_12200;
wire n_12201;
wire n_12202;
wire n_12203;
wire n_12204;
wire n_12205;
wire n_12206;
wire n_12207;
wire n_12208;
wire n_12209;
wire n_12210;
wire n_12211;
wire n_12212;
wire n_12213;
wire n_12214;
wire n_12215;
wire n_12216;
wire n_12217;
wire n_12218;
wire n_12219;
wire n_12220;
wire n_12221;
wire n_12222;
wire n_12223;
wire n_12224;
wire n_12225;
wire n_12226;
wire n_12227;
wire n_12228;
wire n_12229;
wire n_12230;
wire n_12231;
wire n_12232;
wire n_12233;
wire n_12234;
wire n_12235;
wire n_12236;
wire n_12237;
wire n_12238;
wire n_12239;
wire n_12240;
wire n_12241;
wire n_12242;
wire n_12243;
wire n_12244;
wire n_12245;
wire n_12246;
wire n_12247;
wire n_12248;
wire n_12249;
wire n_12250;
wire n_12251;
wire n_12252;
wire n_12253;
wire n_12254;
wire n_12255;
wire n_12256;
wire n_12257;
wire n_12258;
wire n_12259;
wire n_12260;
wire n_12261;
wire n_12262;
wire n_12263;
wire n_12264;
wire n_12265;
wire n_12266;
wire n_12267;
wire n_12268;
wire n_12269;
wire n_12270;
wire n_12271;
wire n_12272;
wire n_12273;
wire n_12274;
wire n_12275;
wire n_12276;
wire n_12277;
wire n_12278;
wire n_12279;
wire n_12280;
wire n_12281;
wire n_12282;
wire n_12283;
wire n_12284;
wire n_12285;
wire n_12286;
wire n_12287;
wire n_12288;
wire n_12289;
wire n_12290;
wire n_12291;
wire n_12292;
wire n_12293;
wire n_12294;
wire n_12295;
wire n_12296;
wire n_12297;
wire n_12298;
wire n_12299;
wire n_12300;
wire n_12301;
wire n_12302;
wire n_12303;
wire n_12304;
wire n_12305;
wire n_12306;
wire n_12307;
wire n_12308;
wire n_12309;
wire n_12310;
wire n_12311;
wire n_12312;
wire n_12313;
wire n_12314;
wire n_12315;
wire n_12316;
wire n_12317;
wire n_12318;
wire n_12319;
wire n_12320;
wire n_12321;
wire n_12322;
wire n_12323;
wire n_12324;
wire n_12325;
wire n_12326;
wire n_12327;
wire n_12328;
wire n_12329;
wire n_12330;
wire n_12331;
wire n_12332;
wire n_12333;
wire n_12334;
wire n_12335;
wire n_12336;
wire n_12337;
wire n_12338;
wire n_12339;
wire n_12340;
wire n_12341;
wire n_12342;
wire n_12343;
wire n_12344;
wire n_12345;
wire n_12346;
wire n_12347;
wire n_12348;
wire n_12349;
wire n_12350;
wire n_12351;
wire n_12352;
wire n_12353;
wire n_12354;
wire n_12355;
wire n_12356;
wire n_12357;
wire n_12358;
wire n_12359;
wire n_12360;
wire n_12361;
wire n_12362;
wire n_12363;
wire n_12364;
wire n_12365;
wire n_12366;
wire n_12367;
wire n_12368;
wire n_12369;
wire n_12370;
wire n_12371;
wire n_12372;
wire n_12373;
wire n_12374;
wire n_12375;
wire n_12376;
wire n_12377;
wire n_12378;
wire n_12379;
wire n_12380;
wire n_12381;
wire n_12382;
wire n_12383;
wire n_12384;
wire n_12385;
wire n_12386;
wire n_12387;
wire n_12388;
wire n_12389;
wire n_12390;
wire n_12391;
wire n_12392;
wire n_12393;
wire n_12394;
wire n_12395;
wire n_12396;
wire n_12397;
wire n_12398;
wire n_12399;
wire n_12400;
wire n_12401;
wire n_12402;
wire n_12403;
wire n_12404;
wire n_12405;
wire n_12406;
wire n_12407;
wire n_12408;
wire n_12409;
wire n_12410;
wire n_12411;
wire n_12412;
wire n_12413;
wire n_12414;
wire n_12415;
wire n_12416;
wire n_12417;
wire n_12418;
wire n_12419;
wire n_12420;
wire n_12421;
wire n_12422;
wire n_12423;
wire n_12424;
wire n_12425;
wire n_12426;
wire n_12427;
wire n_12428;
wire n_12429;
wire n_12430;
wire n_12431;
wire n_12432;
wire n_12433;
wire n_12434;
wire n_12435;
wire n_12436;
wire n_12437;
wire n_12438;
wire n_12439;
wire n_12440;
wire n_12441;
wire n_12442;
wire n_12443;
wire n_12444;
wire n_12445;
wire n_12446;
wire n_12447;
wire n_12448;
wire n_12449;
wire n_12450;
wire n_12451;
wire n_12452;
wire n_12453;
wire n_12454;
wire n_12455;
wire n_12456;
wire n_12457;
wire n_12458;
wire n_12459;
wire n_12460;
wire n_12461;
wire n_12462;
wire n_12463;
wire n_12464;
wire n_12465;
wire n_12466;
wire n_12467;
wire n_12468;
wire n_12469;
wire n_12470;
wire n_12471;
wire n_12472;
wire n_12473;
wire n_12474;
wire n_12475;
wire n_12476;
wire n_12477;
wire n_12478;
wire n_12479;
wire n_12480;
wire n_12481;
wire n_12482;
wire n_12483;
wire n_12484;
wire n_12485;
wire n_12486;
wire n_12487;
wire n_12488;
wire n_12489;
wire n_12490;
wire n_12491;
wire n_12492;
wire n_12493;
wire n_12494;
wire n_12495;
wire n_12496;
wire n_12497;
wire n_12498;
wire n_12499;
wire n_12500;
wire n_12501;
wire n_12502;
wire n_12503;
wire n_12504;
wire n_12505;
wire n_12506;
wire n_12507;
wire n_12508;
wire n_12509;
wire n_12510;
wire n_12511;
wire n_12512;
wire n_12513;
wire n_12514;
wire n_12515;
wire n_12516;
wire n_12517;
wire n_12518;
wire n_12519;
wire n_12520;
wire n_12521;
wire n_12522;
wire n_12523;
wire n_12524;
wire n_12525;
wire n_12526;
wire n_12527;
wire n_12528;
wire n_12529;
wire n_12530;
wire n_12531;
wire n_12532;
wire n_12533;
wire n_12534;
wire n_12535;
wire n_12536;
wire n_12537;
wire n_12538;
wire n_12539;
wire n_12540;
wire n_12541;
wire n_12542;
wire n_12543;
wire n_12544;
wire n_12545;
wire n_12546;
wire n_12547;
wire n_12548;
wire n_12549;
wire n_12550;
wire n_12551;
wire n_12552;
wire n_12553;
wire n_12554;
wire n_12555;
wire n_12556;
wire n_12557;
wire n_12558;
wire n_12559;
wire n_12560;
wire n_12561;
wire n_12562;
wire n_12563;
wire n_12564;
wire n_12565;
wire n_12566;
wire n_12567;
wire n_12568;
wire n_12569;
wire n_12570;
wire n_12571;
wire n_12572;
wire n_12573;
wire n_12574;
wire n_12575;
wire n_12576;
wire n_12577;
wire n_12578;
wire n_12579;
wire n_12580;
wire n_12581;
wire n_12582;
wire n_12583;
wire n_12584;
wire n_12585;
wire n_12586;
wire n_12587;
wire n_12588;
wire n_12589;
wire n_12590;
wire n_12591;
wire n_12592;
wire n_12593;
wire n_12594;
wire n_12595;
wire n_12596;
wire n_12597;
wire n_12598;
wire n_12599;
wire n_12600;
wire n_12601;
wire n_12602;
wire n_12603;
wire n_12604;
wire n_12605;
wire n_12606;
wire n_12607;
wire n_12608;
wire n_12609;
wire n_12610;
wire n_12611;
wire n_12612;
wire n_12613;
wire n_12614;
wire n_12615;
wire n_12616;
wire n_12617;
wire n_12618;
wire n_12619;
wire n_12620;
wire n_12621;
wire n_12622;
wire n_12623;
wire n_12624;
wire n_12625;
wire n_12626;
wire n_12627;
wire n_12628;
wire n_12629;
wire n_12630;
wire n_12631;
wire n_12632;
wire n_12633;
wire n_12634;
wire n_12635;
wire n_12636;
wire n_12637;
wire n_12638;
wire n_12639;
wire n_12640;
wire n_12641;
wire n_12642;
wire n_12643;
wire n_12644;
wire n_12645;
wire n_12646;
wire n_12647;
wire n_12648;
wire n_12649;
wire n_12650;
wire n_12651;
wire n_12652;
wire n_12653;
wire n_12654;
wire n_12655;
wire n_12656;
wire n_12657;
wire n_12658;
wire n_12659;
wire n_12660;
wire n_12661;
wire n_12662;
wire n_12663;
wire n_12664;
wire n_12665;
wire n_12666;
wire n_12667;
wire n_12668;
wire n_12669;
wire n_12670;
wire n_12671;
wire n_12672;
wire n_12673;
wire n_12674;
wire n_12675;
wire n_12676;
wire n_12677;
wire n_12678;
wire n_12679;
wire n_12680;
wire n_12681;
wire n_12682;
wire n_12683;
wire n_12684;
wire n_12685;
wire n_12686;
wire n_12687;
wire n_12688;
wire n_12689;
wire n_12690;
wire n_12691;
wire n_12692;
wire n_12693;
wire n_12694;
wire n_12695;
wire n_12696;
wire n_12697;
wire n_12698;
wire n_12699;
wire n_12700;
wire n_12701;
wire n_12702;
wire n_12703;
wire n_12704;
wire n_12705;
wire n_12706;
wire n_12707;
wire n_12708;
wire n_12709;
wire n_12710;
wire n_12711;
wire n_12712;
wire n_12713;
wire n_12714;
wire n_12715;
wire n_12716;
wire n_12717;
wire n_12718;
wire n_12719;
wire n_12720;
wire n_12721;
wire n_12722;
wire n_12723;
wire n_12724;
wire n_12725;
wire n_12726;
wire n_12727;
wire n_12728;
wire n_12729;
wire n_12730;
wire n_12731;
wire n_12732;
wire n_12733;
wire n_12734;
wire n_12735;
wire n_12736;
wire n_12737;
wire n_12738;
wire n_12739;
wire n_12740;
wire n_12741;
wire n_12742;
wire n_12743;
wire n_12744;
wire n_12745;
wire n_12746;
wire n_12747;
wire n_12748;
wire n_12749;
wire n_12750;
wire n_12751;
wire n_12752;
wire n_12753;
wire n_12754;
wire n_12755;
wire n_12756;
wire n_12757;
wire n_12758;
wire n_12759;
wire n_12760;
wire n_12761;
wire n_12762;
wire n_12763;
wire n_12764;
wire n_12765;
wire n_12766;
wire n_12767;
wire n_12768;
wire n_12769;
wire n_12770;
wire n_12771;
wire n_12772;
wire n_12773;
wire n_12774;
wire n_12775;
wire n_12776;
wire n_12777;
wire n_12778;
wire n_12779;
wire n_12780;
wire n_12781;
wire n_12782;
wire n_12783;
wire n_12784;
wire n_12785;
wire n_12786;
wire n_12787;
wire n_12788;
wire n_12789;
wire n_12790;
wire n_12791;
wire n_12792;
wire n_12793;
wire n_12794;
wire n_12795;
wire n_12796;
wire n_12797;
wire n_12798;
wire n_12799;
wire n_12800;
wire n_12801;
wire n_12802;
wire n_12803;
wire n_12804;
wire n_12805;
wire n_12806;
wire n_12807;
wire n_12808;
wire n_12809;
wire n_12810;
wire n_12811;
wire n_12812;
wire n_12813;
wire n_12814;
wire n_12815;
wire n_12816;
wire n_12817;
wire n_12818;
wire n_12819;
wire n_12820;
wire n_12821;
wire n_12822;
wire n_12823;
wire n_12824;
wire n_12825;
wire n_12826;
wire n_12827;
wire n_12828;
wire n_12829;
wire n_12830;
wire n_12831;
wire n_12832;
wire n_12833;
wire n_12834;
wire n_12835;
wire n_12836;
wire n_12837;
wire n_12838;
wire n_12839;
wire n_12840;
wire n_12841;
wire n_12842;
wire n_12843;
wire n_12844;
wire n_12845;
wire n_12846;
wire n_12847;
wire n_12848;
wire n_12849;
wire n_12850;
wire n_12851;
wire n_12852;
wire n_12853;
wire n_12854;
wire n_12855;
wire n_12856;
wire n_12857;
wire n_12858;
wire n_12859;
wire n_12860;
wire n_12861;
wire n_12862;
wire n_12863;
wire n_12864;
wire n_12865;
wire n_12866;
wire n_12867;
wire n_12868;
wire n_12869;
wire n_12870;
wire n_12871;
wire n_12872;
wire n_12873;
wire n_12874;
wire n_12875;
wire n_12876;
wire n_12877;
wire n_12878;
wire n_12879;
wire n_12880;
wire n_12881;
wire n_12882;
wire n_12883;
wire n_12884;
wire n_12885;
wire n_12886;
wire n_12887;
wire n_12888;
wire n_12889;
wire n_12890;
wire n_12891;
wire n_12892;
wire n_12893;
wire n_12894;
wire n_12895;
wire n_12896;
wire n_12897;
wire n_12898;
wire n_12899;
wire n_12900;
wire n_12901;
wire n_12902;
wire n_12903;
wire n_12904;
wire n_12905;
wire n_12906;
wire n_12907;
wire n_12908;
wire n_12909;
wire n_12910;
wire n_12911;
wire n_12912;
wire n_12913;
wire n_12914;
wire n_12915;
wire n_12916;
wire n_12917;
wire n_12918;
wire n_12919;
wire n_12920;
wire n_12921;
wire n_12922;
wire n_12923;
wire n_12924;
wire n_12925;
wire n_12926;
wire n_12927;
wire n_12928;
wire n_12929;
wire n_12930;
wire n_12931;
wire n_12932;
wire n_12933;
wire n_12934;
wire n_12935;
wire n_12936;
wire n_12937;
wire n_12938;
wire n_12939;
wire n_12940;
wire n_12941;
wire n_12942;
wire n_12943;
wire n_12944;
wire n_12945;
wire n_12946;
wire n_12947;
wire n_12948;
wire n_12949;
wire n_12950;
wire n_12951;
wire n_12952;
wire n_12953;
wire n_12954;
wire n_12955;
wire n_12956;
wire n_12957;
wire n_12958;
wire n_12959;
wire n_12960;
wire n_12961;
wire n_12962;
wire n_12963;
wire n_12964;
wire n_12965;
wire n_12966;
wire n_12967;
wire n_12968;
wire n_12969;
wire n_12970;
wire n_12971;
wire n_12972;
wire n_12973;
wire n_12974;
wire n_12975;
wire n_12976;
wire n_12977;
wire n_12978;
wire n_12979;
wire n_12980;
wire n_12981;
wire n_12982;
wire n_12983;
wire n_12984;
wire n_12985;
wire n_12986;
wire n_12987;
wire n_12988;
wire n_12989;
wire n_12990;
wire n_12991;
wire n_12992;
wire n_12993;
wire n_12994;
wire n_12995;
wire n_12996;
wire n_12997;
wire n_12998;
wire n_12999;
wire n_13000;
wire n_13001;
wire n_13002;
wire n_13003;
wire n_13004;
wire n_13005;
wire n_13006;
wire n_13007;
wire n_13008;
wire n_13009;
wire n_13010;
wire n_13011;
wire n_13012;
wire n_13013;
wire n_13014;
wire n_13015;
wire n_13016;
wire n_13017;
wire n_13018;
wire n_13019;
wire n_13020;
wire n_13021;
wire n_13022;
wire n_13023;
wire n_13024;
wire n_13025;
wire n_13026;
wire n_13027;
wire n_13028;
wire n_13029;
wire n_13030;
wire n_13031;
wire n_13032;
wire n_13033;
wire n_13034;
wire n_13035;
wire n_13036;
wire n_13037;
wire n_13038;
wire n_13039;
wire n_13040;
wire n_13041;
wire n_13042;
wire n_13043;
wire n_13044;
wire n_13045;
wire n_13046;
wire n_13047;
wire n_13048;
wire n_13049;
wire n_13050;
wire n_13051;
wire n_13052;
wire n_13053;
wire n_13054;
wire n_13055;
wire n_13056;
wire n_13057;
wire n_13058;
wire n_13059;
wire n_13060;
wire n_13061;
wire n_13062;
wire n_13063;
wire n_13064;
wire n_13065;
wire n_13066;
wire n_13067;
wire n_13068;
wire n_13069;
wire n_13070;
wire n_13071;
wire n_13072;
wire n_13073;
wire n_13074;
wire n_13075;
wire n_13076;
wire n_13077;
wire n_13078;
wire n_13079;
wire n_13080;
wire n_13081;
wire n_13082;
wire n_13083;
wire n_13084;
wire n_13085;
wire n_13086;
wire n_13087;
wire n_13088;
wire n_13089;
wire n_13090;
wire n_13091;
wire n_13092;
wire n_13093;
wire n_13094;
wire n_13095;
wire n_13096;
wire n_13097;
wire n_13098;
wire n_13099;
wire n_13100;
wire n_13101;
wire n_13102;
wire n_13103;
wire n_13104;
wire n_13105;
wire n_13106;
wire n_13107;
wire n_13108;
wire n_13109;
wire n_13110;
wire n_13111;
wire n_13112;
wire n_13113;
wire n_13114;
wire n_13115;
wire n_13116;
wire n_13117;
wire n_13118;
wire n_13119;
wire n_13120;
wire n_13121;
wire n_13122;
wire n_13123;
wire n_13124;
wire n_13125;
wire n_13126;
wire n_13127;
wire n_13128;
wire n_13129;
wire n_13130;
wire n_13131;
wire n_13132;
wire n_13133;
wire n_13134;
wire n_13135;
wire n_13136;
wire n_13137;
wire n_13138;
wire n_13139;
wire n_13140;
wire n_13141;
wire n_13142;
wire n_13143;
wire n_13144;
wire n_13145;
wire n_13146;
wire n_13147;
wire n_13148;
wire n_13149;
wire n_13150;
wire n_13151;
wire n_13152;
wire n_13153;
wire n_13154;
wire n_13155;
wire n_13156;
wire n_13157;
wire n_13158;
wire n_13159;
wire n_13160;
wire n_13161;
wire n_13162;
wire n_13163;
wire n_13164;
wire n_13165;
wire n_13166;
wire n_13167;
wire n_13168;
wire n_13169;
wire n_13170;
wire n_13171;
wire n_13172;
wire n_13173;
wire n_13174;
wire n_13175;
wire n_13176;
wire n_13177;
wire n_13178;
wire n_13179;
wire n_13180;
wire n_13181;
wire n_13182;
wire n_13183;
wire n_13184;
wire n_13185;
wire n_13186;
wire n_13187;
wire n_13188;
wire n_13189;
wire n_13190;
wire n_13191;
wire n_13192;
wire n_13193;
wire n_13194;
wire n_13195;
wire n_13196;
wire n_13197;
wire n_13198;
wire n_13199;
wire n_13200;
wire n_13201;
wire n_13202;
wire n_13203;
wire n_13204;
wire n_13205;
wire n_13206;
wire n_13207;
wire n_13208;
wire n_13209;
wire n_13210;
wire n_13211;
wire n_13212;
wire n_13213;
wire n_13214;
wire n_13215;
wire n_13216;
wire n_13217;
wire n_13218;
wire n_13219;
wire n_13220;
wire n_13221;
wire n_13222;
wire n_13223;
wire n_13224;
wire n_13225;
wire n_13226;
wire n_13227;
wire n_13228;
wire n_13229;
wire n_13230;
wire n_13231;
wire n_13232;
wire n_13233;
wire n_13234;
wire n_13235;
wire n_13236;
wire n_13237;
wire n_13238;
wire n_13239;
wire n_13240;
wire n_13241;
wire n_13242;
wire n_13243;
wire n_13244;
wire n_13245;
wire n_13246;
wire n_13247;
wire n_13248;
wire n_13249;
wire n_13250;
wire n_13251;
wire n_13252;
wire n_13253;
wire n_13254;
wire n_13255;
wire n_13256;
wire n_13257;
wire n_13258;
wire n_13259;
wire n_13260;
wire n_13261;
wire n_13262;
wire n_13263;
wire n_13264;
wire n_13265;
wire n_13266;
wire n_13267;
wire n_13268;
wire n_13269;
wire n_13270;
wire n_13271;
wire n_13272;
wire n_13273;
wire n_13274;
wire n_13275;
wire n_13276;
wire n_13277;
wire n_13278;
wire n_13279;
wire n_13280;
wire n_13281;
wire n_13282;
wire n_13283;
wire n_13284;
wire n_13285;
wire n_13286;
wire n_13287;
wire n_13288;
wire n_13289;
wire n_13290;
wire n_13291;
wire n_13292;
wire n_13293;
wire n_13294;
wire n_13295;
wire n_13296;
wire n_13297;
wire n_13298;
wire n_13299;
wire n_13300;
wire n_13301;
wire n_13302;
wire n_13303;
wire n_13304;
wire n_13305;
wire n_13306;
wire n_13307;
wire n_13308;
wire n_13309;
wire n_13310;
wire n_13311;
wire n_13312;
wire n_13313;
wire n_13314;
wire n_13315;
wire n_13316;
wire n_13317;
wire n_13318;
wire n_13319;
wire n_13320;
wire n_13321;
wire n_13322;
wire n_13323;
wire n_13324;
wire n_13325;
wire n_13326;
wire n_13327;
wire n_13328;
wire n_13329;
wire n_13330;
wire n_13331;
wire n_13332;
wire n_13333;
wire n_13334;
wire n_13335;
wire n_13336;
wire n_13337;
wire n_13338;
wire n_13339;
wire n_13340;
wire n_13341;
wire n_13342;
wire n_13343;
wire n_13344;
wire n_13345;
wire n_13346;
wire n_13347;
wire n_13348;
wire n_13349;
wire n_13350;
wire n_13351;
wire n_13352;
wire n_13353;
wire n_13354;
wire n_13355;
wire n_13356;
wire n_13357;
wire n_13358;
wire n_13359;
wire n_13360;
wire n_13361;
wire n_13362;
wire n_13363;
wire n_13364;
wire n_13365;
wire n_13366;
wire n_13367;
wire n_13368;
wire n_13369;
wire n_13370;
wire n_13371;
wire n_13372;
wire n_13373;
wire n_13374;
wire n_13375;
wire n_13376;
wire n_13377;
wire n_13378;
wire n_13379;
wire n_13380;
wire n_13381;
wire n_13382;
wire n_13383;
wire n_13384;
wire n_13385;
wire n_13386;
wire n_13387;
wire n_13388;
wire n_13389;
wire n_13390;
wire n_13391;
wire n_13392;
wire n_13393;
wire n_13394;
wire n_13395;
wire n_13396;
wire n_13397;
wire n_13398;
wire n_13399;
wire n_13400;
wire n_13401;
wire n_13402;
wire n_13403;
wire n_13404;
wire n_13405;
wire n_13406;
wire n_13407;
wire n_13408;
wire n_13409;
wire n_13410;
wire n_13411;
wire n_13412;
wire n_13413;
wire n_13414;
wire n_13415;
wire n_13416;
wire n_13417;
wire n_13418;
wire n_13419;
wire n_13420;
wire n_13421;
wire n_13422;
wire n_13423;
wire n_13424;
wire n_13425;
wire n_13426;
wire n_13427;
wire n_13428;
wire n_13429;
wire n_13430;
wire n_13431;
wire n_13432;
wire n_13433;
wire n_13434;
wire n_13435;
wire n_13436;
wire n_13437;
wire n_13438;
wire n_13439;
wire n_13440;
wire n_13441;
wire n_13442;
wire n_13443;
wire n_13444;
wire n_13445;
wire n_13446;
wire n_13447;
wire n_13448;
wire n_13449;
wire n_13450;
wire n_13451;
wire n_13452;
wire n_13453;
wire n_13454;
wire n_13455;
wire n_13456;
wire n_13457;
wire n_13458;
wire n_13459;
wire n_13460;
wire n_13461;
wire n_13462;
wire n_13463;
wire n_13464;
wire n_13465;
wire n_13466;
wire n_13467;
wire n_13468;
wire n_13469;
wire n_13470;
wire n_13471;
wire n_13472;
wire n_13473;
wire n_13474;
wire n_13475;
wire n_13476;
wire n_13477;
wire n_13478;
wire n_13479;
wire n_13480;
wire n_13481;
wire n_13482;
wire n_13483;
wire n_13484;
wire n_13485;
wire n_13486;
wire n_13487;
wire n_13488;
wire n_13489;
wire n_13490;
wire n_13491;
wire n_13492;
wire n_13493;
wire n_13494;
wire n_13495;
wire n_13496;
wire n_13497;
wire n_13498;
wire n_13499;
wire n_13500;
wire n_13501;
wire n_13502;
wire n_13503;
wire n_13504;
wire n_13505;
wire n_13506;
wire n_13507;
wire n_13508;
wire n_13509;
wire n_13510;
wire n_13511;
wire n_13512;
wire n_13513;
wire n_13514;
wire n_13515;
wire n_13516;
wire n_13517;
wire n_13518;
wire n_13519;
wire n_13520;
wire n_13521;
wire n_13522;
wire n_13523;
wire n_13524;
wire n_13525;
wire n_13526;
wire n_13527;
wire n_13528;
wire n_13529;
wire n_13530;
wire n_13531;
wire n_13532;
wire n_13533;
wire n_13534;
wire n_13535;
wire n_13536;
wire n_13537;
wire n_13538;
wire n_13539;
wire n_13540;
wire n_13541;
wire n_13542;
wire n_13543;
wire n_13544;
wire n_13545;
wire n_13546;
wire n_13547;
wire n_13548;
wire n_13549;
wire n_13550;
wire n_13551;
wire n_13552;
wire n_13553;
wire n_13554;
wire n_13555;
wire n_13556;
wire n_13557;
wire n_13558;
wire n_13559;
wire n_13560;
wire n_13561;
wire n_13562;
wire n_13563;
wire n_13564;
wire n_13565;
wire n_13566;
wire n_13567;
wire n_13568;
wire n_13569;
wire n_13570;
wire n_13571;
wire n_13572;
wire n_13573;
wire n_13574;
wire n_13575;
wire n_13576;
wire n_13577;
wire n_13578;
wire n_13579;
wire n_13580;
wire n_13581;
wire n_13582;
wire n_13583;
wire n_13584;
wire n_13585;
wire n_13586;
wire n_13587;
wire n_13588;
wire n_13589;
wire n_13590;
wire n_13591;
wire n_13592;
wire n_13593;
wire n_13594;
wire n_13595;
wire n_13596;
wire n_13597;
wire n_13598;
wire n_13599;
wire n_13600;
wire n_13601;
wire n_13602;
wire n_13603;
wire n_13604;
wire n_13605;
wire n_13606;
wire n_13607;
wire n_13608;
wire n_13609;
wire n_13610;
wire n_13611;
wire n_13612;
wire n_13613;
wire n_13614;
wire n_13615;
wire n_13616;
wire n_13617;
wire n_13618;
wire n_13619;
wire n_13620;
wire n_13621;
wire n_13622;
wire n_13623;
wire n_13624;
wire n_13625;
wire n_13626;
wire n_13627;
wire n_13628;
wire n_13629;
wire n_13630;
wire n_13631;
wire n_13632;
wire n_13633;
wire n_13634;
wire n_13635;
wire n_13636;
wire n_13637;
wire n_13638;
wire n_13639;
wire n_13640;
wire n_13641;
wire n_13642;
wire n_13643;
wire n_13644;
wire n_13645;
wire n_13646;
wire n_13647;
wire n_13648;
wire n_13649;
wire n_13650;
wire n_13651;
wire n_13652;
wire n_13653;
wire n_13654;
wire n_13655;
wire n_13656;
wire n_13657;
wire n_13658;
wire n_13659;
wire n_13660;
wire n_13661;
wire n_13662;
wire n_13663;
wire n_13664;
wire n_13665;
wire n_13666;
wire n_13667;
wire n_13668;
wire n_13669;
wire n_13670;
wire n_13671;
wire n_13672;
wire n_13673;
wire n_13674;
wire n_13675;
wire n_13676;
wire n_13677;
wire n_13678;
wire n_13679;
wire n_13680;
wire n_13681;
wire n_13682;
wire n_13683;
wire n_13684;
wire n_13685;
wire n_13686;
wire n_13687;
wire n_13688;
wire n_13689;
wire n_13690;
wire n_13691;
wire n_13692;
wire n_13693;
wire n_13694;
wire n_13695;
wire n_13696;
wire n_13697;
wire n_13698;
wire n_13699;
wire n_13700;
wire n_13701;
wire n_13702;
wire n_13703;
wire n_13704;
wire n_13705;
wire n_13706;
wire n_13707;
wire n_13708;
wire n_13709;
wire n_13710;
wire n_13711;
wire n_13712;
wire n_13713;
wire n_13714;
wire n_13715;
wire n_13716;
wire n_13717;
wire n_13718;
wire n_13719;
wire n_13720;
wire n_13721;
wire n_13722;
wire n_13723;
wire n_13724;
wire n_13725;
wire n_13726;
wire n_13727;
wire n_13728;
wire n_13729;
wire n_13730;
wire n_13731;
wire n_13732;
wire n_13733;
wire n_13734;
wire n_13735;
wire n_13736;
wire n_13737;
wire n_13738;
wire n_13739;
wire n_13740;
wire n_13741;
wire n_13742;
wire n_13743;
wire n_13744;
wire n_13745;
wire n_13746;
wire n_13747;
wire n_13748;
wire n_13749;
wire n_13750;
wire n_13751;
wire n_13752;
wire n_13753;
wire n_13754;
wire n_13755;
wire n_13756;
wire n_13757;
wire n_13758;
wire n_13759;
wire n_13760;
wire n_13761;
wire n_13762;
wire n_13763;
wire n_13764;
wire n_13765;
wire n_13766;
wire n_13767;
wire n_13768;
wire n_13769;
wire n_13770;
wire n_13771;
wire n_13772;
wire n_13773;
wire n_13774;
wire n_13775;
wire n_13776;
wire n_13777;
wire n_13778;
wire n_13779;
wire n_13780;
wire n_13781;
wire n_13782;
wire n_13783;
wire n_13784;
wire n_13785;
wire n_13786;
wire n_13787;
wire n_13788;
wire n_13789;
wire n_13790;
wire n_13791;
wire n_13792;
wire n_13793;
wire n_13794;
wire n_13795;
wire n_13796;
wire n_13797;
wire n_13798;
wire n_13799;
wire n_13800;
wire n_13801;
wire n_13802;
wire n_13803;
wire n_13804;
wire n_13805;
wire n_13806;
wire n_13807;
wire n_13808;
wire n_13809;
wire n_13810;
wire n_13811;
wire n_13812;
wire n_13813;
wire n_13814;
wire n_13815;
wire n_13816;
wire n_13817;
wire n_13818;
wire n_13819;
wire n_13820;
wire n_13821;
wire n_13822;
wire n_13823;
wire n_13824;
wire n_13825;
wire n_13826;
wire n_13827;
wire n_13828;
wire n_13829;
wire n_13830;
wire n_13831;
wire n_13832;
wire n_13833;
wire n_13834;
wire n_13835;
wire n_13836;
wire n_13837;
wire n_13838;
wire n_13839;
wire n_13840;
wire n_13841;
wire n_13842;
wire n_13843;
wire n_13844;
wire n_13845;
wire n_13846;
wire n_13847;
wire n_13848;
wire n_13849;
wire n_13850;
wire n_13851;
wire n_13852;
wire n_13853;
wire n_13854;
wire n_13855;
wire n_13856;
wire n_13857;
wire n_13858;
wire n_13859;
wire n_13860;
wire n_13861;
wire n_13862;
wire n_13863;
wire n_13864;
wire n_13865;
wire n_13866;
wire n_13867;
wire n_13868;
wire n_13869;
wire n_13870;
wire n_13871;
wire n_13872;
wire n_13873;
wire n_13874;
wire n_13875;
wire n_13876;
wire n_13877;
wire n_13878;
wire n_13879;
wire n_13880;
wire n_13881;
wire n_13882;
wire n_13883;
wire n_13884;
wire n_13885;
wire n_13886;
wire n_13887;
wire n_13888;
wire n_13889;
wire n_13890;
wire n_13891;
wire n_13892;
wire n_13893;
wire n_13894;
wire n_13895;
wire n_13896;
wire n_13897;
wire n_13898;
wire n_13899;
wire n_13900;
wire n_13901;
wire n_13902;
wire n_13903;
wire n_13904;
wire n_13905;
wire n_13906;
wire n_13907;
wire n_13908;
wire n_13909;
wire n_13910;
wire n_13911;
wire n_13912;
wire n_13913;
wire n_13914;
wire n_13915;
wire n_13916;
wire n_13917;
wire n_13918;
wire n_13919;
wire n_13920;
wire n_13921;
wire n_13922;
wire n_13923;
wire n_13924;
wire n_13925;
wire n_13926;
wire n_13927;
wire n_13928;
wire n_13929;
wire n_13930;
wire n_13931;
wire n_13932;
wire n_13933;
wire n_13934;
wire n_13935;
wire n_13936;
wire n_13937;
wire n_13938;
wire n_13939;
wire n_13940;
wire n_13941;
wire n_13942;
wire n_13943;
wire n_13944;
wire n_13945;
wire n_13946;
wire n_13947;
wire n_13948;
wire n_13949;
wire n_13950;
wire n_13951;
wire n_13952;
wire n_13953;
wire n_13954;
wire n_13955;
wire n_13956;
wire n_13957;
wire n_13958;
wire n_13959;
wire n_13960;
wire n_13961;
wire n_13962;
wire n_13963;
wire n_13964;
wire n_13965;
wire n_13966;
wire n_13967;
wire n_13968;
wire n_13969;
wire n_13970;
wire n_13971;
wire n_13972;
wire n_13973;
wire n_13974;
wire n_13975;
wire n_13976;
wire n_13977;
wire n_13978;
wire n_13979;
wire n_13980;
wire n_13981;
wire n_13982;
wire n_13983;
wire n_13984;
wire n_13985;
wire n_13986;
wire n_13987;
wire n_13988;
wire n_13989;
wire n_13990;
wire n_13991;
wire n_13992;
wire n_13993;
wire n_13994;
wire n_13995;
wire n_13996;
wire n_13997;
wire n_13998;
wire n_13999;
wire n_14000;
wire n_14001;
wire n_14002;
wire n_14003;
wire n_14004;
wire n_14005;
wire n_14006;
wire n_14007;
wire n_14008;
wire n_14009;
wire n_14010;
wire n_14011;
wire n_14012;
wire n_14013;
wire n_14014;
wire n_14015;
wire n_14016;
wire n_14017;
wire n_14018;
wire n_14019;
wire n_14020;
wire n_14021;
wire n_14022;
wire n_14023;
wire n_14024;
wire n_14025;
wire n_14026;
wire n_14027;
wire n_14028;
wire n_14029;
wire n_14030;
wire n_14031;
wire n_14032;
wire n_14033;
wire n_14034;
wire n_14035;
wire n_14036;
wire n_14037;
wire n_14038;
wire n_14039;
wire n_14040;
wire n_14041;
wire n_14042;
wire n_14043;
wire n_14044;
wire n_14045;
wire n_14046;
wire n_14047;
wire n_14048;
wire n_14049;
wire n_14050;
wire n_14051;
wire n_14052;
wire n_14053;
wire n_14054;
wire n_14055;
wire n_14056;
wire n_14057;
wire n_14058;
wire n_14059;
wire n_14060;
wire n_14061;
wire n_14062;
wire n_14063;
wire n_14064;
wire n_14065;
wire n_14066;
wire n_14067;
wire n_14068;
wire n_14069;
wire n_14070;
wire n_14071;
wire n_14072;
wire n_14073;
wire n_14074;
wire n_14075;
wire n_14076;
wire n_14077;
wire n_14078;
wire n_14079;
wire n_14080;
wire n_14081;
wire n_14082;
wire n_14083;
wire n_14084;
wire n_14085;
wire n_14086;
wire n_14087;
wire n_14088;
wire n_14089;
wire n_14090;
wire n_14091;
wire n_14092;
wire n_14093;
wire n_14094;
wire n_14095;
wire n_14096;
wire n_14097;
wire n_14098;
wire n_14099;
wire n_14100;
wire n_14101;
wire n_14102;
wire n_14103;
wire n_14104;
wire n_14105;
wire n_14106;
wire n_14107;
wire n_14108;
wire n_14109;
wire n_14110;
wire n_14111;
wire n_14112;
wire n_14113;
wire n_14114;
wire n_14115;
wire n_14116;
wire n_14117;
wire n_14118;
wire n_14119;
wire n_14120;
wire n_14121;
wire n_14122;
wire n_14123;
wire n_14124;
wire n_14125;
wire n_14126;
wire n_14127;
wire n_14128;
wire n_14129;
wire n_14130;
wire n_14131;
wire n_14132;
wire n_14133;
wire n_14134;
wire n_14135;
wire n_14136;
wire n_14137;
wire n_14138;
wire n_14139;
wire n_14140;
wire n_14141;
wire n_14142;
wire n_14143;
wire n_14144;
wire n_14145;
wire n_14146;
wire n_14147;
wire n_14148;
wire n_14149;
wire n_14150;
wire n_14151;
wire n_14152;
wire n_14153;
wire n_14154;
wire n_14155;
wire n_14156;
wire n_14157;
wire n_14158;
wire n_14159;
wire n_14160;
wire n_14161;
wire n_14162;
wire n_14163;
wire n_14164;
wire n_14165;
wire n_14166;
wire n_14167;
wire n_14168;
wire n_14169;
wire n_14170;
wire n_14171;
wire n_14172;
wire n_14173;
wire n_14174;
wire n_14175;
wire n_14176;
wire n_14177;
wire n_14178;
wire n_14179;
wire n_14180;
wire n_14181;
wire n_14182;
wire n_14183;
wire n_14184;
wire n_14185;
wire n_14186;
wire n_14187;
wire n_14188;
wire n_14189;
wire n_14190;
wire n_14191;
wire n_14192;
wire n_14193;
wire n_14194;
wire n_14195;
wire n_14196;
wire n_14197;
wire n_14198;
wire n_14199;
wire n_14200;
wire n_14201;
wire n_14202;
wire n_14203;
wire n_14204;
wire n_14205;
wire n_14206;
wire n_14207;
wire n_14208;
wire n_14209;
wire n_14210;
wire n_14211;
wire n_14212;
wire n_14213;
wire n_14214;
wire n_14215;
wire n_14216;
wire n_14217;
wire n_14218;
wire n_14219;
wire n_14220;
wire n_14221;
wire n_14222;
wire n_14223;
wire n_14224;
wire n_14225;
wire n_14226;
wire n_14227;
wire n_14228;
wire n_14229;
wire n_14230;
wire n_14231;
wire n_14232;
wire n_14233;
wire n_14234;
wire n_14235;
wire n_14236;
wire n_14237;
wire n_14238;
wire n_14239;
wire n_14240;
wire n_14241;
wire n_14242;
wire n_14243;
wire n_14244;
wire n_14245;
wire n_14246;
wire n_14247;
wire n_14248;
wire n_14249;
wire n_14250;
wire n_14251;
wire n_14252;
wire n_14253;
wire n_14254;
wire n_14255;
wire n_14256;
wire n_14257;
wire n_14258;
wire n_14259;
wire n_14260;
wire n_14261;
wire n_14262;
wire n_14263;
wire n_14264;
wire n_14265;
wire n_14266;
wire n_14267;
wire n_14268;
wire n_14269;
wire n_14270;
wire n_14271;
wire n_14272;
wire n_14273;
wire n_14274;
wire n_14275;
wire n_14276;
wire n_14277;
wire n_14278;
wire n_14279;
wire n_14280;
wire n_14281;
wire n_14282;
wire n_14283;
wire n_14284;
wire n_14285;
wire n_14286;
wire n_14287;
wire n_14288;
wire n_14289;
wire n_14290;
wire n_14291;
wire n_14292;
wire n_14293;
wire n_14294;
wire n_14295;
wire n_14296;
wire n_14297;
wire n_14298;
wire n_14299;
wire n_14300;
wire n_14301;
wire n_14302;
wire n_14303;
wire n_14304;
wire n_14305;
wire n_14306;
wire n_14307;
wire n_14308;
wire n_14309;
wire n_14310;
wire n_14311;
wire n_14312;
wire n_14313;
wire n_14314;
wire n_14315;
wire n_14316;
wire n_14317;
wire n_14318;
wire n_14319;
wire n_14320;
wire n_14321;
wire n_14322;
wire n_14323;
wire n_14324;
wire n_14325;
wire n_14326;
wire n_14327;
wire n_14328;
wire n_14329;
wire n_14330;
wire n_14331;
wire n_14332;
wire n_14333;
wire n_14334;
wire n_14335;
wire n_14336;
wire n_14337;
wire n_14338;
wire n_14339;
wire n_14340;
wire n_14341;
wire n_14342;
wire n_14343;
wire n_14344;
wire n_14345;
wire n_14346;
wire n_14347;
wire n_14348;
wire n_14349;
wire n_14350;
wire n_14351;
wire n_14352;
wire n_14353;
wire n_14354;
wire n_14355;
wire n_14356;
wire n_14357;
wire n_14358;
wire n_14359;
wire n_14360;
wire n_14361;
wire n_14362;
wire n_14363;
wire n_14364;
wire n_14365;
wire n_14366;
wire n_14367;
wire n_14368;
wire n_14369;
wire n_14370;
wire n_14371;
wire n_14372;
wire n_14373;
wire n_14374;
wire n_14375;
wire n_14376;
wire n_14377;
wire n_14378;
wire n_14379;
wire n_14380;
wire n_14381;
wire n_14382;
wire n_14383;
wire n_14384;
wire n_14385;
wire n_14386;
wire n_14387;
wire n_14388;
wire n_14389;
wire n_14390;
wire n_14391;
wire n_14392;
wire n_14393;
wire n_14394;
wire n_14395;
wire n_14396;
wire n_14397;
wire n_14398;
wire n_14399;
wire n_14400;
wire n_14401;
wire n_14402;
wire n_14403;
wire n_14404;
wire n_14405;
wire n_14406;
wire n_14407;
wire n_14408;
wire n_14409;
wire n_14410;
wire n_14411;
wire n_14412;
wire n_14413;
wire n_14414;
wire n_14415;
wire n_14416;
wire n_14417;
wire n_14418;
wire n_14419;
wire n_14420;
wire n_14421;
wire n_14422;
wire n_14423;
wire n_14424;
wire n_14425;
wire n_14426;
wire n_14427;
wire n_14428;
wire n_14429;
wire n_14430;
wire n_14431;
wire n_14432;
wire n_14433;
wire n_14434;
wire n_14435;
wire n_14436;
wire n_14437;
wire n_14438;
wire n_14439;
wire n_14440;
wire n_14441;
wire n_14442;
wire n_14443;
wire n_14444;
wire n_14445;
wire n_14446;
wire n_14447;
wire n_14448;
wire n_14449;
wire n_14450;
wire n_14451;
wire n_14452;
wire n_14453;
wire n_14454;
wire n_14455;
wire n_14456;
wire n_14457;
wire n_14458;
wire n_14459;
wire n_14460;
wire n_14461;
wire n_14462;
wire n_14463;
wire n_14464;
wire n_14465;
wire n_14466;
wire n_14467;
wire n_14468;
wire n_14469;
wire n_14470;
wire n_14471;
wire n_14472;
wire n_14473;
wire n_14474;
wire n_14475;
wire n_14476;
wire n_14477;
wire n_14478;
wire n_14479;
wire n_14480;
wire n_14481;
wire n_14482;
wire n_14483;
wire n_14484;
wire n_14485;
wire n_14486;
wire n_14487;
wire n_14488;
wire n_14489;
wire n_14490;
wire n_14491;
wire n_14492;
wire n_14493;
wire n_14494;
wire n_14495;
wire n_14496;
wire n_14497;
wire n_14498;
wire n_14499;
wire n_14500;
wire n_14501;
wire n_14502;
wire n_14503;
wire n_14504;
wire n_14505;
wire n_14506;
wire n_14507;
wire n_14508;
wire n_14509;
wire n_14510;
wire n_14511;
wire n_14512;
wire n_14513;
wire n_14514;
wire n_14515;
wire n_14516;
wire n_14517;
wire n_14518;
wire n_14519;
wire n_14520;
wire n_14521;
wire n_14522;
wire n_14523;
wire n_14524;
wire n_14525;
wire n_14526;
wire n_14527;
wire n_14528;
wire n_14529;
wire n_14530;
wire n_14531;
wire n_14532;
wire n_14533;
wire n_14534;
wire n_14535;
wire n_14536;
wire n_14537;
wire n_14538;
wire n_14539;
wire n_14540;
wire n_14541;
wire n_14542;
wire n_14543;
wire n_14544;
wire n_14545;
wire n_14546;
wire n_14547;
wire n_14548;
wire n_14549;
wire n_14550;
wire n_14551;
wire n_14552;
wire n_14553;
wire n_14554;
wire n_14555;
wire n_14556;
wire n_14557;
wire n_14558;
wire n_14559;
wire n_14560;
wire n_14561;
wire n_14562;
wire n_14563;
wire n_14564;
wire n_14565;
wire n_14566;
wire n_14567;
wire n_14568;
wire n_14569;
wire n_14570;
wire n_14571;
wire n_14572;
wire n_14573;
wire n_14574;
wire n_14575;
wire n_14576;
wire n_14577;
wire n_14578;
wire n_14579;
wire n_14580;
wire n_14581;
wire n_14582;
wire n_14583;
wire n_14584;
wire n_14585;
wire n_14586;
wire n_14587;
wire n_14588;
wire n_14589;
wire n_14590;
wire n_14591;
wire n_14592;
wire n_14593;
wire n_14594;
wire n_14595;
wire n_14596;
wire n_14597;
wire n_14598;
wire n_14599;
wire n_14600;
wire n_14601;
wire n_14602;
wire n_14603;
wire n_14604;
wire n_14605;
wire n_14606;
wire n_14607;
wire n_14608;
wire n_14609;
wire n_14610;
wire n_14611;
wire n_14612;
wire n_14613;
wire n_14614;
wire n_14615;
wire n_14616;
wire n_14617;
wire n_14618;
wire n_14619;
wire n_14620;
wire n_14621;
wire n_14622;
wire n_14623;
wire n_14624;
wire n_14625;
wire n_14626;
wire n_14627;
wire n_14628;
wire n_14629;
wire n_14630;
wire n_14631;
wire n_14632;
wire n_14633;
wire n_14634;
wire n_14635;
wire n_14636;
wire n_14637;
wire n_14638;
wire n_14639;
wire n_14640;
wire n_14641;
wire n_14642;
wire n_14643;
wire n_14644;
wire n_14645;
wire n_14646;
wire n_14647;
wire n_14648;
wire n_14649;
wire n_14650;
wire n_14651;
wire n_14652;
wire n_14653;
wire n_14654;
wire n_14655;
wire n_14656;
wire n_14657;
wire n_14658;
wire n_14659;
wire n_14660;
wire n_14661;
wire n_14662;
wire n_14663;
wire n_14664;
wire n_14665;
wire n_14666;
wire n_14667;
wire n_14668;
wire n_14669;
wire n_14670;
wire n_14671;
wire n_14672;
wire n_14673;
wire n_14674;
wire n_14675;
wire n_14676;
wire n_14677;
wire n_14678;
wire n_14679;
wire n_14680;
wire n_14681;
wire n_14682;
wire n_14683;
wire n_14684;
wire n_14685;
wire n_14686;
wire n_14687;
wire n_14688;
wire n_14689;
wire n_14690;
wire n_14691;
wire n_14692;
wire n_14693;
wire n_14694;
wire n_14695;
wire n_14696;
wire n_14697;
wire n_14698;
wire n_14699;
wire n_14700;
wire n_14701;
wire n_14702;
wire n_14703;
wire n_14704;
wire n_14705;
wire n_14706;
wire n_14707;
wire n_14708;
wire n_14709;
wire n_14710;
wire n_14711;
wire n_14712;
wire n_14713;
wire n_14714;
wire n_14715;
wire n_14716;
wire n_14717;
wire n_14718;
wire n_14719;
wire n_14720;
wire n_14721;
wire n_14722;
wire n_14723;
wire n_14724;
wire n_14725;
wire n_14726;
wire n_14727;
wire n_14728;
wire n_14729;
wire n_14730;
wire n_14731;
wire n_14732;
wire n_14733;
wire n_14734;
wire n_14735;
wire n_14736;
wire n_14737;
wire n_14738;
wire n_14739;
wire n_14740;
wire n_14741;
wire n_14742;
wire n_14743;
wire n_14744;
wire n_14745;
wire n_14746;
wire n_14747;
wire n_14748;
wire n_14749;
wire n_14750;
wire n_14751;
wire n_14752;
wire n_14753;
wire n_14754;
wire n_14755;
wire n_14756;
wire n_14757;
wire n_14758;
wire n_14759;
wire n_14760;
wire n_14761;
wire n_14762;
wire n_14763;
wire n_14764;
wire n_14765;
wire n_14766;
wire n_14767;
wire n_14768;
wire n_14769;
wire n_14770;
wire n_14771;
wire n_14772;
wire n_14773;
wire n_14774;
wire n_14775;
wire n_14776;
wire n_14777;
wire n_14778;
wire n_14779;
wire n_14780;
wire n_14781;
wire n_14782;
wire n_14783;
wire n_14784;
wire n_14785;
wire n_14786;
wire n_14787;
wire n_14788;
wire n_14789;
wire n_14790;
wire n_14791;
wire n_14792;
wire n_14793;
wire n_14794;
wire n_14795;
wire n_14796;
wire n_14797;
wire n_14798;
wire n_14799;
wire n_14800;
wire n_14801;
wire n_14802;
wire n_14803;
wire n_14804;
wire n_14805;
wire n_14806;
wire n_14807;
wire n_14808;
wire n_14809;
wire n_14810;
wire n_14811;
wire n_14812;
wire n_14813;
wire n_14814;
wire n_14815;
wire n_14816;
wire n_14817;
wire n_14818;
wire n_14819;
wire n_14820;
wire n_14821;
wire n_14822;
wire n_14823;
wire n_14824;
wire n_14825;
wire n_14826;
wire n_14827;
wire n_14828;
wire n_14829;
wire n_14830;
wire n_14831;
wire n_14832;
wire n_14833;
wire n_14834;
wire n_14835;
wire n_14836;
wire n_14837;
wire n_14838;
wire n_14839;
wire n_14840;
wire n_14841;
wire n_14842;
wire n_14843;
wire n_14844;
wire n_14845;
wire n_14846;
wire n_14847;
wire n_14848;
wire n_14849;
wire n_14850;
wire n_14851;
wire n_14852;
wire n_14853;
wire n_14854;
wire n_14855;
wire n_14856;
wire n_14857;
wire n_14858;
wire n_14859;
wire n_14860;
wire n_14861;
wire n_14862;
wire n_14863;
wire n_14864;
wire n_14865;
wire n_14866;
wire n_14867;
wire n_14868;
wire n_14869;
wire n_14870;
wire n_14871;
wire n_14872;
wire n_14873;
wire n_14874;
wire n_14875;
wire n_14876;
wire n_14877;
wire n_14878;
wire n_14879;
wire n_14880;
wire n_14881;
wire n_14882;
wire n_14883;
wire n_14884;
wire n_14885;
wire n_14886;
wire n_14887;
wire n_14888;
wire n_14889;
wire n_14890;
wire n_14891;
wire n_14892;
wire n_14893;
wire n_14894;
wire n_14895;
wire n_14896;
wire n_14897;
wire n_14898;
wire n_14899;
wire n_14900;
wire n_14901;
wire n_14902;
wire n_14903;
wire n_14904;
wire n_14905;
wire n_14906;
wire n_14907;
wire n_14908;
wire n_14909;
wire n_14910;
wire n_14911;
wire n_14912;
wire n_14913;
wire n_14914;
wire n_14915;
wire n_14916;
wire n_14917;
wire n_14918;
wire n_14919;
wire n_14920;
wire n_14921;
wire n_14922;
wire n_14923;
wire n_14924;
wire n_14925;
wire n_14926;
wire n_14927;
wire n_14928;
wire n_14929;
wire n_14930;
wire n_14931;
wire n_14932;
wire n_14933;
wire n_14934;
wire n_14935;
wire n_14936;
wire n_14937;
wire n_14938;
wire n_14939;
wire n_14940;
wire n_14941;
wire n_14942;
wire n_14943;
wire n_14944;
wire n_14945;
wire n_14946;
wire n_14947;
wire n_14948;
wire n_14949;
wire n_14950;
wire n_14951;
wire n_14952;
wire n_14953;
wire n_14954;
wire n_14955;
wire n_14956;
wire n_14957;
wire n_14958;
wire n_14959;
wire n_14960;
wire n_14961;
wire n_14962;
wire n_14963;
wire n_14964;
wire n_14965;
wire n_14966;
wire n_14967;
wire n_14968;
wire n_14969;
wire n_14970;
wire n_14971;
wire n_14972;
wire n_14973;
wire n_14974;
wire n_14975;
wire n_14976;
wire n_14977;
wire n_14978;
wire n_14979;
wire n_14980;
wire n_14981;
wire n_14982;
wire n_14983;
wire n_14984;
wire n_14985;
wire n_14986;
wire n_14987;
wire n_14988;
wire n_14989;
wire n_14990;
wire n_14991;
wire n_14992;
wire n_14993;
wire n_14994;
wire n_14995;
wire n_14996;
wire n_14997;
wire n_14998;
wire n_14999;
wire n_15000;
wire n_15001;
wire n_15002;
wire n_15003;
wire n_15004;
wire n_15005;
wire n_15006;
wire n_15007;
wire n_15008;
wire n_15009;
wire n_15010;
wire n_15011;
wire n_15012;
wire n_15013;
wire n_15014;
wire n_15015;
wire n_15016;
wire n_15017;
wire n_15018;
wire n_15019;
wire n_15020;
wire n_15021;
wire n_15022;
wire n_15023;
wire n_15024;
wire n_15025;
wire n_15026;
wire n_15027;
wire n_15028;
wire n_15029;
wire n_15030;
wire n_15031;
wire n_15032;
wire n_15033;
wire n_15034;
wire n_15035;
wire n_15036;
wire n_15037;
wire n_15038;
wire n_15039;
wire n_15040;
wire n_15041;
wire n_15042;
wire n_15043;
wire n_15044;
wire n_15045;
wire n_15046;
wire n_15047;
wire n_15048;
wire n_15049;
wire n_15050;
wire n_15051;
wire n_15052;
wire n_15053;
wire n_15054;
wire n_15055;
wire n_15056;
wire n_15057;
wire n_15058;
wire n_15059;
wire n_15060;
wire n_15061;
wire n_15062;
wire n_15063;
wire n_15064;
wire n_15065;
wire n_15066;
wire n_15067;
wire n_15068;
wire n_15069;
wire n_15070;
wire n_15071;
wire n_15072;
wire n_15073;
wire n_15074;
wire n_15075;
wire n_15076;
wire n_15077;
wire n_15078;
wire n_15079;
wire n_15080;
wire n_15081;
wire n_15082;
wire n_15083;
wire n_15084;
wire n_15085;
wire n_15086;
wire n_15087;
wire n_15088;
wire n_15089;
wire n_15090;
wire n_15091;
wire n_15092;
wire n_15093;
wire n_15094;
wire n_15095;
wire n_15096;
wire n_15097;
wire n_15098;
wire n_15099;
wire n_15100;
wire n_15101;
wire n_15102;
wire n_15103;
wire n_15104;
wire n_15105;
wire n_15106;
wire n_15107;
wire n_15108;
wire n_15109;
wire n_15110;
wire n_15111;
wire n_15112;
wire n_15113;
wire n_15114;
wire n_15115;
wire n_15116;
wire n_15117;
wire n_15118;
wire n_15119;
wire n_15120;
wire n_15121;
wire n_15122;
wire n_15123;
wire n_15124;
wire n_15125;
wire n_15126;
wire n_15127;
wire n_15128;
wire n_15129;
wire n_15130;
wire n_15131;
wire n_15132;
wire n_15133;
wire n_15134;
wire n_15135;
wire n_15136;
wire n_15137;
wire n_15138;
wire n_15139;
wire n_15140;
wire n_15141;
wire n_15142;
wire n_15143;
wire n_15144;
wire n_15145;
wire n_15146;
wire n_15147;
wire n_15148;
wire n_15149;
wire n_15150;
wire n_15151;
wire n_15152;
wire n_15153;
wire n_15154;
wire n_15155;
wire n_15156;
wire n_15157;
wire n_15158;
wire n_15159;
wire n_15160;
wire n_15161;
wire n_15162;
wire n_15163;
wire n_15164;
wire n_15165;
wire n_15166;
wire n_15167;
wire n_15168;
wire n_15169;
wire n_15170;
wire n_15171;
wire n_15172;
wire n_15173;
wire n_15174;
wire n_15175;
wire n_15176;
wire n_15177;
wire n_15178;
wire n_15179;
wire n_15180;
wire n_15181;
wire n_15182;
wire n_15183;
wire n_15184;
wire n_15185;
wire n_15186;
wire n_15187;
wire n_15188;
wire n_15189;
wire n_15190;
wire n_15191;
wire n_15192;
wire n_15193;
wire n_15194;
wire n_15195;
wire n_15196;
wire n_15197;
wire n_15198;
wire n_15199;
wire n_15200;
wire n_15201;
wire n_15202;
wire n_15203;
wire n_15204;
wire n_15205;
wire n_15206;
wire n_15207;
wire n_15208;
wire n_15209;
wire n_15210;
wire n_15211;
wire n_15212;
wire n_15213;
wire n_15214;
wire n_15215;
wire n_15216;
wire n_15217;
wire n_15218;
wire n_15219;
wire n_15220;
wire n_15221;
wire n_15222;
wire n_15223;
wire n_15224;
wire n_15225;
wire n_15226;
wire n_15227;
wire n_15228;
wire n_15229;
wire n_15230;
wire n_15231;
wire n_15232;
wire n_15233;
wire n_15234;
wire n_15235;
wire n_15236;
wire n_15237;
wire n_15238;
wire n_15239;
wire n_15240;
wire n_15241;
wire n_15242;
wire n_15243;
wire n_15244;
wire n_15245;
wire n_15246;
wire n_15247;
wire n_15248;
wire n_15249;
wire n_15250;
wire n_15251;
wire n_15252;
wire n_15253;
wire n_15254;
wire n_15255;
wire n_15256;
wire n_15257;
wire n_15258;
wire n_15259;
wire n_15260;
wire n_15261;
wire n_15262;
wire n_15263;
wire n_15264;
wire n_15265;
wire n_15266;
wire n_15267;
wire n_15268;
wire n_15269;
wire n_15270;
wire n_15271;
wire n_15272;
wire n_15273;
wire n_15274;
wire n_15275;
wire n_15276;
wire n_15277;
wire n_15278;
wire n_15279;
wire n_15280;
wire n_15281;
wire n_15282;
wire n_15283;
wire n_15284;
wire n_15285;
wire n_15286;
wire n_15287;
wire n_15288;
wire n_15289;
wire n_15290;
wire n_15291;
wire n_15292;
wire n_15293;
wire n_15294;
wire n_15295;
wire n_15296;
wire n_15297;
wire n_15298;
wire n_15299;
wire n_15300;
wire n_15301;
wire n_15302;
wire n_15303;
wire n_15304;
wire n_15305;
wire n_15306;
wire n_15307;
wire n_15308;
wire n_15309;
wire n_15310;
wire n_15311;
wire n_15312;
wire n_15313;
wire n_15314;
wire n_15315;
wire n_15316;
wire n_15317;
wire n_15318;
wire n_15319;
wire n_15320;
wire n_15321;
wire n_15322;
wire n_15323;
wire n_15324;
wire n_15325;
wire n_15326;
wire n_15327;
wire n_15328;
wire n_15329;
wire n_15330;
wire n_15331;
wire n_15332;
wire n_15333;
wire n_15334;
wire n_15335;
wire n_15336;
wire n_15337;
wire n_15338;
wire n_15339;
wire n_15340;
wire n_15341;
wire n_15342;
wire n_15343;
wire n_15344;
wire n_15345;
wire n_15346;
wire n_15347;
wire n_15348;
wire n_15349;
wire n_15350;
wire n_15351;
wire n_15352;
wire n_15353;
wire n_15354;
wire n_15355;
wire n_15356;
wire n_15357;
wire n_15358;
wire n_15359;
wire n_15360;
wire n_15361;
wire n_15362;
wire n_15363;
wire n_15364;
wire n_15365;
wire n_15366;
wire n_15367;
wire n_15368;
wire n_15369;
wire n_15370;
wire n_15371;
wire n_15372;
wire n_15373;
wire n_15374;
wire n_15375;
wire n_15376;
wire n_15377;
wire n_15378;
wire n_15379;
wire n_15380;
wire n_15381;
wire n_15382;
wire n_15383;
wire n_15384;
wire n_15385;
wire n_15386;
wire n_15387;
wire n_15388;
wire n_15389;
wire n_15390;
wire n_15391;
wire n_15392;
wire n_15393;
wire n_15394;
wire n_15395;
wire n_15396;
wire n_15397;
wire n_15398;
wire n_15399;
wire n_15400;
wire n_15401;
wire n_15402;
wire n_15403;
wire n_15404;
wire n_15405;
wire n_15406;
wire n_15407;
wire n_15408;
wire n_15409;
wire n_15410;
wire n_15411;
wire n_15412;
wire n_15413;
wire n_15414;
wire n_15415;
wire n_15416;
wire n_15417;
wire n_15418;
wire n_15419;
wire n_15420;
wire n_15421;
wire n_15422;
wire n_15423;
wire n_15424;
wire n_15425;
wire n_15426;
wire n_15427;
wire n_15428;
wire n_15429;
wire n_15430;
wire n_15431;
wire n_15432;
wire n_15433;
wire n_15434;
wire n_15435;
wire n_15436;
wire n_15437;
wire n_15438;
wire n_15439;
wire n_15440;
wire n_15441;
wire n_15442;
wire n_15443;
wire n_15444;
wire n_15445;
wire n_15446;
wire n_15447;
wire n_15448;
wire n_15449;
wire n_15450;
wire n_15451;
wire n_15452;
wire n_15453;
wire n_15454;
wire n_15455;
wire n_15456;
wire n_15457;
wire n_15458;
wire n_15459;
wire n_15460;
wire n_15461;
wire n_15462;
wire n_15463;
wire n_15464;
wire n_15465;
wire n_15466;
wire n_15467;
wire n_15468;
wire n_15469;
wire n_15470;
wire n_15471;
wire n_15472;
wire n_15473;
wire n_15474;
wire n_15475;
wire n_15476;
wire n_15477;
wire n_15478;
wire n_15479;
wire n_15480;
wire n_15481;
wire n_15482;
wire n_15483;
wire n_15484;
wire n_15485;
wire n_15486;
wire n_15487;
wire n_15488;
wire n_15489;
wire n_15490;
wire n_15491;
wire n_15492;
wire n_15493;
wire n_15494;
wire n_15495;
wire n_15496;
wire n_15497;
wire n_15498;
wire n_15499;
wire n_15500;
wire n_15501;
wire n_15502;
wire n_15503;
wire n_15504;
wire n_15505;
wire n_15506;
wire n_15507;
wire n_15508;
wire n_15509;
wire n_15510;
wire n_15511;
wire n_15512;
wire n_15513;
wire n_15514;
wire n_15515;
wire n_15516;
wire n_15517;
wire n_15518;
wire n_15519;
wire n_15520;
wire n_15521;
wire n_15522;
wire n_15523;
wire n_15524;
wire n_15525;
wire n_15526;
wire n_15527;
wire n_15528;
wire n_15529;
wire n_15530;
wire n_15531;
wire n_15532;
wire n_15533;
wire n_15534;
wire n_15535;
wire n_15536;
wire n_15537;
wire n_15538;
wire n_15539;
wire n_15540;
wire n_15541;
wire n_15542;
wire n_15543;
wire n_15544;
wire n_15545;
wire n_15546;
wire n_15547;
wire n_15548;
wire n_15549;
wire n_15550;
wire n_15551;
wire n_15552;
wire n_15553;
wire n_15554;
wire n_15555;
wire n_15556;
wire n_15557;
wire n_15558;
wire n_15559;
wire n_15560;
wire n_15561;
wire n_15562;
wire n_15563;
wire n_15564;
wire n_15565;
wire n_15566;
wire n_15567;
wire n_15568;
wire n_15569;
wire n_15570;
wire n_15571;
wire n_15572;
wire n_15573;
wire n_15574;
wire n_15575;
wire n_15576;
wire n_15577;
wire n_15578;
wire n_15579;
wire n_15580;
wire n_15581;
wire n_15582;
wire n_15583;
wire n_15584;
wire n_15585;
wire n_15586;
wire n_15587;
wire n_15588;
wire n_15589;
wire n_15590;
wire n_15591;
wire n_15592;
wire n_15593;
wire n_15594;
wire n_15595;
wire n_15596;
wire n_15597;
wire n_15598;
wire n_15599;
wire n_15600;
wire n_15601;
wire n_15602;
wire n_15603;
wire n_15604;
wire n_15605;
wire n_15606;
wire n_15607;
wire n_15608;
wire n_15609;
wire n_15610;
wire n_15611;
wire n_15612;
wire n_15613;
wire n_15614;
wire n_15615;
wire n_15616;
wire n_15617;
wire n_15618;
wire n_15619;
wire n_15620;
wire n_15621;
wire n_15622;
wire n_15623;
wire n_15624;
wire n_15625;
wire n_15626;
wire n_15627;
wire n_15628;
wire n_15629;
wire n_15630;
wire n_15631;
wire n_15632;
wire n_15633;
wire n_15634;
wire n_15635;
wire n_15636;
wire n_15637;
wire n_15638;
wire n_15639;
wire n_15640;
wire n_15641;
wire n_15642;
wire n_15643;
wire n_15644;
wire n_15645;
wire n_15646;
wire n_15647;
wire n_15648;
wire n_15649;
wire n_15650;
wire n_15651;
wire n_15652;
wire n_15653;
wire n_15654;
wire n_15655;
wire n_15656;
wire n_15657;
wire n_15658;
wire n_15659;
wire n_15660;
wire n_15661;
wire n_15662;
wire n_15663;
wire n_15664;
wire n_15665;
wire n_15666;
wire n_15667;
wire n_15668;
wire n_15669;
wire n_15670;
wire n_15671;
wire n_15672;
wire n_15673;
wire n_15674;
wire n_15675;
wire n_15676;
wire n_15677;
wire n_15678;
wire n_15679;
wire n_15680;
wire n_15681;
wire n_15682;
wire n_15683;
wire n_15684;
wire n_15685;
wire n_15686;
wire n_15687;
wire n_15688;
wire n_15689;
wire n_15690;
wire n_15691;
wire n_15692;
wire n_15693;
wire n_15694;
wire n_15695;
wire n_15696;
wire n_15697;
wire n_15698;
wire n_15699;
wire n_15700;
wire n_15701;
wire n_15702;
wire n_15703;
wire n_15704;
wire n_15705;
wire n_15706;
wire n_15707;
wire n_15708;
wire n_15709;
wire n_15710;
wire n_15711;
wire n_15712;
wire n_15713;
wire n_15714;
wire n_15715;
wire n_15716;
wire n_15717;
wire n_15718;
wire n_15719;
wire n_15720;
wire n_15721;
wire n_15722;
wire n_15723;
wire n_15724;
wire n_15725;
wire n_15726;
wire n_15727;
wire n_15728;
wire n_15729;
wire n_15730;
wire n_15731;
wire n_15732;
wire n_15733;
wire n_15734;
wire n_15735;
wire n_15736;
wire n_15737;
wire n_15738;
wire n_15739;
wire n_15740;
wire n_15741;
wire n_15742;
wire n_15743;
wire n_15744;
wire n_15745;
wire n_15746;
wire n_15747;
wire n_15748;
wire n_15749;
wire n_15750;
wire n_15751;
wire n_15752;
wire n_15753;
wire n_15754;
wire n_15755;
wire n_15756;
wire n_15757;
wire n_15758;
wire n_15759;
wire n_15760;
wire n_15761;
wire n_15762;
wire n_15763;
wire n_15764;
wire n_15765;
wire n_15766;
wire n_15767;
wire n_15768;
wire n_15769;
wire n_15770;
wire n_15771;
wire n_15772;
wire n_15773;
wire n_15774;
wire n_15775;
wire n_15776;
wire n_15777;
wire n_15778;
wire n_15779;
wire n_15780;
wire n_15781;
wire n_15782;
wire n_15783;
wire n_15784;
wire n_15785;
wire n_15786;
wire n_15787;
wire n_15788;
wire n_15789;
wire n_15790;
wire n_15791;
wire n_15792;
wire n_15793;
wire n_15794;
wire n_15795;
wire n_15796;
wire n_15797;
wire n_15798;
wire n_15799;
wire n_15800;
wire n_15801;
wire n_15802;
wire n_15803;
wire n_15804;
wire n_15805;
wire n_15806;
wire n_15807;
wire n_15808;
wire n_15809;
wire n_15810;
wire n_15811;
wire n_15812;
wire n_15813;
wire n_15814;
wire n_15815;
wire n_15816;
wire n_15817;
wire n_15818;
wire n_15819;
wire n_15820;
wire n_15821;
wire n_15822;
wire n_15823;
wire n_15824;
wire n_15825;
wire n_15826;
wire n_15827;
wire n_15828;
wire n_15829;
wire n_15830;
wire n_15831;
wire n_15832;
wire n_15833;
wire n_15834;
wire n_15835;
wire n_15836;
wire n_15837;
wire n_15838;
wire n_15839;
wire n_15840;
wire n_15841;
wire n_15842;
wire n_15843;
wire n_15844;
wire n_15845;
wire n_15846;
wire n_15847;
wire n_15848;
wire n_15849;
wire n_15850;
wire n_15851;
wire n_15852;
wire n_15853;
wire n_15854;
wire n_15855;
wire n_15856;
wire n_15857;
wire n_15858;
wire n_15859;
wire n_15860;
wire n_15861;
wire n_15862;
wire n_15863;
wire n_15864;
wire n_15865;
wire n_15866;
wire n_15867;
wire n_15868;
wire n_15869;
wire n_15870;
wire n_15871;
wire n_15872;
wire n_15873;
wire n_15874;
wire n_15875;
wire n_15876;
wire n_15877;
wire n_15878;
wire n_15879;
wire n_15880;
wire n_15881;
wire n_15882;
wire n_15883;
wire n_15884;
wire n_15885;
wire n_15886;
wire n_15887;
wire n_15888;
wire n_15889;
wire n_15890;
wire n_15891;
wire n_15892;
wire n_15893;
wire n_15894;
wire n_15895;
wire n_15896;
wire n_15897;
wire n_15898;
wire n_15899;
wire n_15900;
wire n_15901;
wire n_15902;
wire n_15903;
wire n_15904;
wire n_15905;
wire n_15906;
wire n_15907;
wire n_15908;
wire n_15909;
wire n_15910;
wire n_15911;
wire n_15912;
wire n_15913;
wire n_15914;
wire n_15915;
wire n_15916;
wire n_15917;
wire n_15918;
wire n_15919;
wire n_15920;
wire n_15921;
wire n_15922;
wire n_15923;
wire n_15924;
wire n_15925;
wire n_15926;
wire n_15927;
wire n_15928;
wire n_15929;
wire n_15930;
wire n_15931;
wire n_15932;
wire n_15933;
wire n_15934;
wire n_15935;
wire n_15936;
wire n_15937;
wire n_15938;
wire n_15939;
wire n_15940;
wire n_15941;
wire n_15942;
wire n_15943;
wire n_15944;
wire n_15945;
wire n_15946;
wire n_15947;
wire n_15948;
wire n_15949;
wire n_15950;
wire n_15951;
wire n_15952;
wire n_15953;
wire n_15954;
wire n_15955;
wire n_15956;
wire n_15957;
wire n_15958;
wire n_15959;
wire n_15960;
wire n_15961;
wire n_15962;
wire n_15963;
wire n_15964;
wire n_15965;
wire n_15966;
wire n_15967;
wire n_15968;
wire n_15969;
wire n_15970;
wire n_15971;
wire n_15972;
wire n_15973;
wire n_15974;
wire n_15975;
wire n_15976;
wire n_15977;
wire n_15978;
wire n_15979;
wire n_15980;
wire n_15981;
wire n_15982;
wire n_15983;
wire n_15984;
wire n_15985;
wire n_15986;
wire n_15987;
wire n_15988;
wire n_15989;
wire n_15990;
wire n_15991;
wire n_15992;
wire n_15993;
wire n_15994;
wire n_15995;
wire n_15996;
wire n_15997;
wire n_15998;
wire n_15999;
wire n_16000;
wire n_16001;
wire n_16002;
wire n_16003;
wire n_16004;
wire n_16005;
wire n_16006;
wire n_16007;
wire n_16008;
wire n_16009;
wire n_16010;
wire n_16011;
wire n_16012;
wire n_16013;
wire n_16014;
wire n_16015;
wire n_16016;
wire n_16017;
wire n_16018;
wire n_16019;
wire n_16020;
wire n_16021;
wire n_16022;
wire n_16023;
wire n_16024;
wire n_16025;
wire n_16026;
wire n_16027;
wire n_16028;
wire n_16029;
wire n_16030;
wire n_16031;
wire n_16032;
wire n_16033;
wire n_16034;
wire n_16035;
wire n_16036;
wire n_16037;
wire n_16038;
wire n_16039;
wire n_16040;
wire n_16041;
wire n_16042;
wire n_16043;
wire n_16044;
wire n_16045;
wire n_16046;
wire n_16047;
wire n_16048;
wire n_16049;
wire n_16050;
wire n_16051;
wire n_16052;
wire n_16053;
wire n_16054;
wire n_16055;
wire n_16056;
wire n_16057;
wire n_16058;
wire n_16059;
wire n_16060;
wire n_16061;
wire n_16062;
wire n_16063;
wire n_16064;
wire n_16065;
wire n_16066;
wire n_16067;
wire n_16068;
wire n_16069;
wire n_16070;
wire n_16071;
wire n_16072;
wire n_16073;
wire n_16074;
wire n_16075;
wire n_16076;
wire n_16077;
wire n_16078;
wire n_16079;
wire n_16080;
wire n_16081;
wire n_16082;
wire n_16083;
wire n_16084;
wire n_16085;
wire n_16086;
wire n_16087;
wire n_16088;
wire n_16089;
wire n_16090;
wire n_16091;
wire n_16092;
wire n_16093;
wire n_16094;
wire n_16095;
wire n_16096;
wire n_16097;
wire n_16098;
wire n_16099;
wire n_16100;
wire n_16101;
wire n_16102;
wire n_16103;
wire n_16104;
wire n_16105;
wire n_16106;
wire n_16107;
wire n_16108;
wire n_16109;
wire n_16110;
wire n_16111;
wire n_16112;
wire n_16113;
wire n_16114;
wire n_16115;
wire n_16116;
wire n_16117;
wire n_16118;
wire n_16119;
wire n_16120;
wire n_16121;
wire n_16122;
wire n_16123;
wire n_16124;
wire n_16125;
wire n_16126;
wire n_16127;
wire n_16128;
wire n_16129;
wire n_16130;
wire n_16131;
wire n_16132;
wire n_16133;
wire n_16134;
wire n_16135;
wire n_16136;
wire n_16137;
wire n_16138;
wire n_16139;
wire n_16140;
wire n_16141;
wire n_16142;
wire n_16143;
wire n_16144;
wire n_16145;
wire n_16146;
wire n_16147;
wire n_16148;
wire n_16149;
wire n_16150;
wire n_16151;
wire n_16152;
wire n_16153;
wire n_16154;
wire n_16155;
wire n_16156;
wire n_16157;
wire n_16158;
wire n_16159;
wire n_16160;
wire n_16161;
wire n_16162;
wire n_16163;
wire n_16164;
wire n_16165;
wire n_16166;
wire n_16167;
wire n_16168;
wire n_16169;
wire n_16170;
wire n_16171;
wire n_16172;
wire n_16173;
wire n_16174;
wire n_16175;
wire n_16176;
wire n_16177;
wire n_16178;
wire n_16179;
wire n_16180;
wire n_16181;
wire n_16182;
wire n_16183;
wire n_16184;
wire n_16185;
wire n_16186;
wire n_16187;
wire n_16188;
wire n_16189;
wire n_16190;
wire n_16191;
wire n_16192;
wire n_16193;
wire n_16194;
wire n_16195;
wire n_16196;
wire n_16197;
wire n_16198;
wire n_16199;
wire n_16200;
wire n_16201;
wire n_16202;
wire n_16203;
wire n_16204;
wire n_16205;
wire n_16206;
wire n_16207;
wire n_16208;
wire n_16209;
wire n_16210;
wire n_16211;
wire n_16212;
wire n_16213;
wire n_16214;
wire n_16215;
wire n_16216;
wire n_16217;
wire n_16218;
wire n_16219;
wire n_16220;
wire n_16221;
wire n_16222;
wire n_16223;
wire n_16224;
wire n_16225;
wire n_16226;
wire n_16227;
wire n_16228;
wire n_16229;
wire n_16230;
wire n_16231;
wire n_16232;
wire n_16233;
wire n_16234;
wire n_16235;
wire n_16236;
wire n_16237;
wire n_16238;
wire n_16239;
wire n_16240;
wire n_16241;
wire n_16242;
wire n_16243;
wire n_16244;
wire n_16245;
wire n_16246;
wire n_16247;
wire n_16248;
wire n_16249;
wire n_16250;
wire n_16251;
wire n_16252;
wire n_16253;
wire n_16254;
wire n_16255;
wire n_16256;
wire n_16257;
wire n_16258;
wire n_16259;
wire n_16260;
wire n_16261;
wire n_16262;
wire n_16263;
wire n_16264;
wire n_16265;
wire n_16266;
wire n_16267;
wire n_16268;
wire n_16269;
wire n_16270;
wire n_16271;
wire n_16272;
wire n_16273;
wire n_16274;
wire n_16275;
wire n_16276;
wire n_16277;
wire n_16278;
wire n_16279;
wire n_16280;
wire n_16281;
wire n_16282;
wire n_16283;
wire n_16284;
wire n_16285;
wire n_16286;
wire n_16287;
wire n_16288;
wire n_16289;
wire n_16290;
wire n_16291;
wire n_16292;
wire n_16293;
wire n_16294;
wire n_16295;
wire n_16296;
wire n_16297;
wire n_16298;
wire n_16299;
wire n_16300;
wire n_16301;
wire n_16302;
wire n_16303;
wire n_16304;
wire n_16305;
wire n_16306;
wire n_16307;
wire n_16308;
wire n_16309;
wire n_16310;
wire n_16311;
wire n_16312;
wire n_16313;
wire n_16314;
wire n_16315;
wire n_16316;
wire n_16317;
wire n_16318;
wire n_16319;
wire n_16320;
wire n_16321;
wire n_16322;
wire n_16323;
wire n_16324;
wire n_16325;
wire n_16326;
wire n_16327;
wire n_16328;
wire n_16329;
wire n_16330;
wire n_16331;
wire n_16332;
wire n_16333;
wire n_16334;
wire n_16335;
wire n_16336;
wire n_16337;
wire n_16338;
wire n_16339;
wire n_16340;
wire n_16341;
wire n_16342;
wire n_16343;
wire n_16344;
wire n_16345;
wire n_16346;
wire n_16347;
wire n_16348;
wire n_16349;
wire n_16350;
wire n_16351;
wire n_16352;
wire n_16353;
wire n_16354;
wire n_16355;
wire n_16356;
wire n_16357;
wire n_16358;
wire n_16359;
wire n_16360;
wire n_16361;
wire n_16362;
wire n_16363;
wire n_16364;
wire n_16365;
wire n_16366;
wire n_16367;
wire n_16368;
wire n_16369;
wire n_16370;
wire n_16371;
wire n_16372;
wire n_16373;
wire n_16374;
wire n_16375;
wire n_16376;
wire n_16377;
wire n_16378;
wire n_16379;
wire n_16380;
wire n_16381;
wire n_16382;
wire n_16383;
wire n_16384;
wire n_16385;
wire n_16386;
wire n_16387;
wire n_16388;
wire n_16389;
wire n_16390;
wire n_16391;
wire n_16392;
wire n_16393;
wire n_16394;
wire n_16395;
wire n_16396;
wire n_16397;
wire n_16398;
wire n_16399;
wire n_16400;
wire n_16401;
wire n_16402;
wire n_16403;
wire n_16404;
wire n_16405;
wire n_16406;
wire n_16407;
wire n_16408;
wire n_16409;
wire n_16410;
wire n_16411;
wire n_16412;
wire n_16413;
wire n_16414;
wire n_16415;
wire n_16416;
wire n_16417;
wire n_16418;
wire n_16419;
wire n_16420;
wire n_16421;
wire n_16422;
wire n_16423;
wire n_16424;
wire n_16425;
wire n_16426;
wire n_16427;
wire n_16428;
wire n_16429;
wire n_16430;
wire n_16431;
wire n_16432;
wire n_16433;
wire n_16434;
wire n_16435;
wire n_16436;
wire n_16437;
wire n_16438;
wire n_16439;
wire n_16440;
wire n_16441;
wire n_16442;
wire n_16443;
wire n_16444;
wire n_16445;
wire n_16446;
wire n_16447;
wire n_16448;
wire n_16449;
wire n_16450;
wire n_16451;
wire n_16452;
wire n_16453;
wire n_16454;
wire n_16455;
wire n_16456;
wire n_16457;
wire n_16458;
wire n_16459;
wire n_16460;
wire n_16461;
wire n_16462;
wire n_16463;
wire n_16464;
wire n_16465;
wire n_16466;
wire n_16467;
wire n_16468;
wire n_16469;
wire n_16470;
wire n_16471;
wire n_16472;
wire n_16473;
wire n_16474;
wire n_16475;
wire n_16476;
wire n_16477;
wire n_16478;
wire n_16479;
wire n_16480;
wire n_16481;
wire n_16482;
wire n_16483;
wire n_16484;
wire n_16485;
wire n_16486;
wire n_16487;
wire n_16488;
wire n_16489;
wire n_16490;
wire n_16491;
wire n_16492;
wire n_16493;
wire n_16494;
wire n_16495;
wire n_16496;
wire n_16497;
wire n_16498;
wire n_16499;
wire n_16500;
wire n_16501;
wire n_16502;
wire n_16503;
wire n_16504;
wire n_16505;
wire n_16506;
wire n_16507;
wire n_16508;
wire n_16509;
wire n_16510;
wire n_16511;
wire n_16512;
wire n_16513;
wire n_16514;
wire n_16515;
wire n_16516;
wire n_16517;
wire n_16518;
wire n_16519;
wire n_16520;
wire n_16521;
wire n_16522;
wire n_16523;
wire n_16524;
wire n_16525;
wire n_16526;
wire n_16527;
wire n_16528;
wire n_16529;
wire n_16530;
wire n_16531;
wire n_16532;
wire n_16533;
wire n_16534;
wire n_16535;
wire n_16536;
wire n_16537;
wire n_16538;
wire n_16539;
wire n_16540;
wire n_16541;
wire n_16542;
wire n_16543;
wire n_16544;
wire n_16545;
wire n_16546;
wire n_16547;
wire n_16548;
wire n_16549;
wire n_16550;
wire n_16551;
wire n_16552;
wire n_16553;
wire n_16554;
wire n_16555;
wire n_16556;
wire n_16557;
wire n_16558;
wire n_16559;
wire n_16560;
wire n_16561;
wire n_16562;
wire n_16563;
wire n_16564;
wire n_16565;
wire n_16566;
wire n_16567;
wire n_16568;
wire n_16569;
wire n_16570;
wire n_16571;
wire n_16572;
wire n_16573;
wire n_16574;
wire n_16575;
wire n_16576;
wire n_16577;
wire n_16578;
wire n_16579;
wire n_16580;
wire n_16581;
wire n_16582;
wire n_16583;
wire n_16584;
wire n_16585;
wire n_16586;
wire n_16587;
wire n_16588;
wire n_16589;
wire n_16590;
wire n_16591;
wire n_16592;
wire n_16593;
wire n_16594;
wire n_16595;
wire n_16596;
wire n_16597;
wire n_16598;
wire n_16599;
wire n_16600;
wire n_16601;
wire n_16602;
wire n_16603;
wire n_16604;
wire n_16605;
wire n_16606;
wire n_16607;
wire n_16608;
wire n_16609;
wire n_16610;
wire n_16611;
wire n_16612;
wire n_16613;
wire n_16614;
wire n_16615;
wire n_16616;
wire n_16617;
wire n_16618;
wire n_16619;
wire n_16620;
wire n_16621;
wire n_16622;
wire n_16623;
wire n_16624;
wire n_16625;
wire n_16626;
wire n_16627;
wire n_16628;
wire n_16629;
wire n_16630;
wire n_16631;
wire n_16632;
wire n_16633;
wire n_16634;
wire n_16635;
wire n_16636;
wire n_16637;
wire n_16638;
wire n_16639;
wire n_16640;
wire n_16641;
wire n_16642;
wire n_16643;
wire n_16644;
wire n_16645;
wire n_16646;
wire n_16647;
wire n_16648;
wire n_16649;
wire n_16650;
wire n_16651;
wire n_16652;
wire n_16653;
wire n_16654;
wire n_16655;
wire n_16656;
wire n_16657;
wire n_16658;
wire n_16659;
wire n_16660;
wire n_16661;
wire n_16662;
wire n_16663;
wire n_16664;
wire n_16665;
wire n_16666;
wire n_16667;
wire n_16668;
wire n_16669;
wire n_16670;
wire n_16671;
wire n_16672;
wire n_16673;
wire n_16674;
wire n_16675;
wire n_16676;
wire n_16677;
wire n_16678;
wire n_16679;
wire n_16680;
wire n_16681;
wire n_16682;
wire n_16683;
wire n_16684;
wire n_16685;
wire n_16686;
wire n_16687;
wire n_16688;
wire n_16689;
wire n_16690;
wire n_16691;
wire n_16692;
wire n_16693;
wire n_16694;
wire n_16695;
wire n_16696;
wire n_16697;
wire n_16698;
wire n_16699;
wire n_16700;
wire n_16701;
wire n_16702;
wire n_16703;
wire n_16704;
wire n_16705;
wire n_16706;
wire n_16707;
wire n_16708;
wire n_16709;
wire n_16710;
wire n_16711;
wire n_16712;
wire n_16713;
wire n_16714;
wire n_16715;
wire n_16716;
wire n_16717;
wire n_16718;
wire n_16719;
wire n_16720;
wire n_16721;
wire n_16722;
wire n_16723;
wire n_16724;
wire n_16725;
wire n_16726;
wire n_16727;
wire n_16728;
wire n_16729;
wire n_16730;
wire n_16731;
wire n_16732;
wire n_16733;
wire n_16734;
wire n_16735;
wire n_16736;
wire n_16737;
wire n_16738;
wire n_16739;
wire n_16740;
wire n_16741;
wire n_16742;
wire n_16743;
wire n_16744;
wire n_16745;
wire n_16746;
wire n_16747;
wire n_16748;
wire n_16749;
wire n_16750;
wire n_16751;
wire n_16752;
wire n_16753;
wire n_16754;
wire n_16755;
wire n_16756;
wire n_16757;
wire n_16758;
wire n_16759;
wire n_16760;
wire n_16761;
wire n_16762;
wire n_16763;
wire n_16764;
wire n_16765;
wire n_16766;
wire n_16767;
wire n_16768;
wire n_16769;
wire n_16770;
wire n_16771;
wire n_16772;
wire n_16773;
wire n_16774;
wire n_16775;
wire n_16776;
wire n_16777;
wire n_16778;
wire n_16779;
wire n_16780;
wire n_16781;
wire n_16782;
wire n_16783;
wire n_16784;
wire n_16785;
wire n_16786;
wire n_16787;
wire n_16788;
wire n_16789;
wire n_16790;
wire n_16791;
wire n_16792;
wire n_16793;
wire n_16794;
wire n_16795;
wire n_16796;
wire n_16797;
wire n_16798;
wire n_16799;
wire n_16800;
wire n_16801;
wire n_16802;
wire n_16803;
wire n_16804;
wire n_16805;
wire n_16806;
wire n_16807;
wire n_16808;
wire n_16809;
wire n_16810;
wire n_16811;
wire n_16812;
wire n_16813;
wire n_16814;
wire n_16815;
wire n_16816;
wire n_16817;
wire n_16818;
wire n_16819;
wire n_16820;
wire n_16821;
wire n_16822;
wire n_16823;
wire n_16824;
wire n_16825;
wire n_16826;
wire n_16827;
wire n_16828;
wire n_16829;
wire n_16830;
wire n_16831;
wire n_16832;
wire n_16833;
wire n_16834;
wire n_16835;
wire n_16836;
wire n_16837;
wire n_16838;
wire n_16839;
wire n_16840;
wire n_16841;
wire n_16842;
wire n_16843;
wire n_16844;
wire n_16845;
wire n_16846;
wire n_16847;
wire n_16848;
wire n_16849;
wire n_16850;
wire n_16851;
wire n_16852;
wire n_16853;
wire n_16854;
wire n_16855;
wire n_16856;
wire n_16857;
wire n_16858;
wire n_16859;
wire n_16860;
wire n_16861;
wire n_16862;
wire n_16863;
wire n_16864;
wire n_16865;
wire n_16866;
wire n_16867;
wire n_16868;
wire n_16869;
wire n_16870;
wire n_16871;
wire n_16872;
wire n_16873;
wire n_16874;
wire n_16875;
wire n_16876;
wire n_16877;
wire n_16878;
wire n_16879;
wire n_16880;
wire n_16881;
wire n_16882;
wire n_16883;
wire n_16884;
wire n_16885;
wire n_16886;
wire n_16887;
wire n_16888;
wire n_16889;
wire n_16890;
wire n_16891;
wire n_16892;
wire n_16893;
wire n_16894;
wire n_16895;
wire n_16896;
wire n_16897;
wire n_16898;
wire n_16899;
wire n_16900;
wire n_16901;
wire n_16902;
wire n_16903;
wire n_16904;
wire n_16905;
wire n_16906;
wire n_16907;
wire n_16908;
wire n_16909;
wire n_16910;
wire n_16911;
wire n_16912;
wire n_16913;
wire n_16914;
wire n_16915;
wire n_16916;
wire n_16917;
wire n_16918;
wire n_16919;
wire n_16920;
wire n_16921;
wire n_16922;
wire n_16923;
wire n_16924;
wire n_16925;
wire n_16926;
wire n_16927;
wire n_16928;
wire n_16929;
wire n_16930;
wire n_16931;
wire n_16932;
wire n_16933;
wire n_16934;
wire n_16935;
wire n_16936;
wire n_16937;
wire n_16938;
wire n_16939;
wire n_16940;
wire n_16941;
wire n_16942;
wire n_16943;
wire n_16944;
wire n_16945;
wire n_16946;
wire n_16947;
wire n_16948;
wire n_16949;
wire n_16950;
wire n_16951;
wire n_16952;
wire n_16953;
wire n_16954;
wire n_16955;
wire n_16956;
wire n_16957;
wire n_16958;
wire n_16959;
wire n_16960;
wire n_16961;
wire n_16962;
wire n_16963;
wire n_16964;
wire n_16965;
wire n_16966;
wire n_16967;
wire n_16968;
wire n_16969;
wire n_16970;
wire n_16971;
wire n_16972;
wire n_16973;
wire n_16974;
wire n_16975;
wire n_16976;
wire n_16977;
wire n_16978;
wire n_16979;
wire n_16980;
wire n_16981;
wire n_16982;
wire n_16983;
wire n_16984;
wire n_16985;
wire n_16986;
wire n_16987;
wire n_16988;
wire n_16989;
wire n_16990;
wire n_16991;
wire n_16992;
wire n_16993;
wire n_16994;
wire n_16995;
wire n_16996;
wire n_16997;
wire n_16998;
wire n_16999;
wire n_17000;
wire n_17001;
wire n_17002;
wire n_17003;
wire n_17004;
wire n_17005;
wire n_17006;
wire n_17007;
wire n_17008;
wire n_17009;
wire n_17010;
wire n_17011;
wire n_17012;
wire n_17013;
wire n_17014;
wire n_17015;
wire n_17016;
wire n_17017;
wire n_17018;
wire n_17019;
wire n_17020;
wire n_17021;
wire n_17022;
wire n_17023;
wire n_17024;
wire n_17025;
wire n_17026;
wire n_17027;
wire n_17028;
wire n_17029;
wire n_17030;
wire n_17031;
wire n_17032;
wire n_17033;
wire n_17034;
wire n_17035;
wire n_17036;
wire n_17037;
wire n_17038;
wire n_17039;
wire n_17040;
wire n_17041;
wire n_17042;
wire n_17043;
wire n_17044;
wire n_17045;
wire n_17046;
wire n_17047;
wire n_17048;
wire n_17049;
wire n_17050;
wire n_17051;
wire n_17052;
wire n_17053;
wire n_17054;
wire n_17055;
wire n_17056;
wire n_17057;
wire n_17058;
wire n_17059;
wire n_17060;
wire n_17061;
wire n_17062;
wire n_17063;
wire n_17064;
wire n_17065;
wire n_17066;
wire n_17067;
wire n_17068;
wire n_17069;
wire n_17070;
wire n_17071;
wire n_17072;
wire n_17073;
wire n_17074;
wire n_17075;
wire n_17076;
wire n_17077;
wire n_17078;
wire n_17079;
wire n_17080;
wire n_17081;
wire n_17082;
wire n_17083;
wire n_17084;
wire n_17085;
wire n_17086;
wire n_17087;
wire n_17088;
wire n_17089;
wire n_17090;
wire n_17091;
wire n_17092;
wire n_17093;
wire n_17094;
wire n_17095;
wire n_17096;
wire n_17097;
wire n_17098;
wire n_17099;
wire n_17100;
wire n_17101;
wire n_17102;
wire n_17103;
wire n_17104;
wire n_17105;
wire n_17106;
wire n_17107;
wire n_17108;
wire n_17109;
wire n_17110;
wire n_17111;
wire n_17112;
wire n_17113;
wire n_17114;
wire n_17115;
wire n_17116;
wire n_17117;
wire n_17118;
wire n_17119;
wire n_17120;
wire n_17121;
wire n_17122;
wire n_17123;
wire n_17124;
wire n_17125;
wire n_17126;
wire n_17127;
wire n_17128;
wire n_17129;
wire n_17130;
wire n_17131;
wire n_17132;
wire n_17133;
wire n_17134;
wire n_17135;
wire n_17136;
wire n_17137;
wire n_17138;
wire n_17139;
wire n_17140;
wire n_17141;
wire n_17142;
wire n_17143;
wire n_17144;
wire n_17145;
wire n_17146;
wire n_17147;
wire n_17148;
wire n_17149;
wire n_17150;
wire n_17151;
wire n_17152;
wire n_17153;
wire n_17154;
wire n_17155;
wire n_17156;
wire n_17157;
wire n_17158;
wire n_17159;
wire n_17160;
wire n_17161;
wire n_17162;
wire n_17163;
wire n_17164;
wire n_17165;
wire n_17166;
wire n_17167;
wire n_17168;
wire n_17169;
wire n_17170;
wire n_17171;
wire n_17172;
wire n_17173;
wire n_17174;
wire n_17175;
wire n_17176;
wire n_17177;
wire n_17178;
wire n_17179;
wire n_17180;
wire n_17181;
wire n_17182;
wire n_17183;
wire n_17184;
wire n_17185;
wire n_17186;
wire n_17187;
wire n_17188;
wire n_17189;
wire n_17190;
wire n_17191;
wire n_17192;
wire n_17193;
wire n_17194;
wire n_17195;
wire n_17196;
wire n_17197;
wire n_17198;
wire n_17199;
wire n_17200;
wire n_17201;
wire n_17202;
wire n_17203;
wire n_17204;
wire n_17205;
wire n_17206;
wire n_17207;
wire n_17208;
wire n_17209;
wire n_17210;
wire n_17211;
wire n_17212;
wire n_17213;
wire n_17214;
wire n_17215;
wire n_17216;
wire n_17217;
wire n_17218;
wire n_17219;
wire n_17220;
wire n_17221;
wire n_17222;
wire n_17223;
wire n_17224;
wire n_17225;
wire n_17226;
wire n_17227;
wire n_17228;
wire n_17229;
wire n_17230;
wire n_17231;
wire n_17232;
wire n_17233;
wire n_17234;
wire n_17235;
wire n_17236;
wire n_17237;
wire n_17238;
wire n_17239;
wire n_17240;
wire n_17241;
wire n_17242;
wire n_17243;
wire n_17244;
wire n_17245;
wire n_17246;
wire n_17247;
wire n_17248;
wire n_17249;
wire n_17250;
wire n_17251;
wire n_17252;
wire n_17253;
wire n_17254;
wire n_17255;
wire n_17256;
wire n_17257;
wire n_17258;
wire n_17259;
wire n_17260;
wire n_17261;
wire n_17262;
wire n_17263;
wire n_17264;
wire n_17265;
wire n_17266;
wire n_17267;
wire n_17268;
wire n_17269;
wire n_17270;
wire n_17271;
wire n_17272;
wire n_17273;
wire n_17274;
wire n_17275;
wire n_17276;
wire n_17277;
wire n_17278;
wire n_17279;
wire n_17280;
wire n_17281;
wire n_17282;
wire n_17283;
wire n_17284;
wire n_17285;
wire n_17286;
wire n_17287;
wire n_17288;
wire n_17289;
wire n_17290;
wire n_17291;
wire n_17292;
wire n_17293;
wire n_17294;
wire n_17295;
wire n_17296;
wire n_17297;
wire n_17298;
wire n_17299;
wire n_17300;
wire n_17301;
wire n_17302;
wire n_17303;
wire n_17304;
wire n_17305;
wire n_17306;
wire n_17307;
wire n_17308;
wire n_17309;
wire n_17310;
wire n_17311;
wire n_17312;
wire n_17313;
wire n_17314;
wire n_17315;
wire n_17316;
wire n_17317;
wire n_17318;
wire n_17319;
wire n_17320;
wire n_17321;
wire n_17322;
wire n_17323;
wire n_17324;
wire n_17325;
wire n_17326;
wire n_17327;
wire n_17328;
wire n_17329;
wire n_17330;
wire n_17331;
wire n_17332;
wire n_17333;
wire n_17334;
wire n_17335;
wire n_17336;
wire n_17337;
wire n_17338;
wire n_17339;
wire n_17340;
wire n_17341;
wire n_17342;
wire n_17343;
wire n_17344;
wire n_17345;
wire n_17346;
wire n_17347;
wire n_17348;
wire n_17349;
wire n_17350;
wire n_17351;
wire n_17352;
wire n_17353;
wire n_17354;
wire n_17355;
wire n_17356;
wire n_17357;
wire n_17358;
wire n_17359;
wire n_17360;
wire n_17361;
wire n_17362;
wire n_17363;
wire n_17364;
wire n_17365;
wire n_17366;
wire n_17367;
wire n_17368;
wire n_17369;
wire n_17370;
wire n_17371;
wire n_17372;
wire n_17373;
wire n_17374;
wire n_17375;
wire n_17376;
wire n_17377;
wire n_17378;
wire n_17379;
wire n_17380;
wire n_17381;
wire n_17382;
wire n_17383;
wire n_17384;
wire n_17385;
wire n_17386;
wire n_17387;
wire n_17388;
wire n_17389;
wire n_17390;
wire n_17391;
wire n_17392;
wire n_17393;
wire n_17394;
wire n_17395;
wire n_17396;
wire n_17397;
wire n_17398;
wire n_17399;
wire n_17400;
wire n_17401;
wire n_17402;
wire n_17403;
wire n_17404;
wire n_17405;
wire n_17406;
wire n_17407;
wire n_17408;
wire n_17409;
wire n_17410;
wire n_17411;
wire n_17412;
wire n_17413;
wire n_17414;
wire n_17415;
wire n_17416;
wire n_17417;
wire n_17418;
wire n_17419;
wire n_17420;
wire n_17421;
wire n_17422;
wire n_17423;
wire n_17424;
wire n_17425;
wire n_17426;
wire n_17427;
wire n_17428;
wire n_17429;
wire n_17430;
wire n_17431;
wire n_17432;
wire n_17433;
wire n_17434;
wire n_17435;
wire n_17436;
wire n_17437;
wire n_17438;
wire n_17439;
wire n_17440;
wire n_17441;
wire n_17442;
wire n_17443;
wire n_17444;
wire n_17445;
wire n_17446;
wire n_17447;
wire n_17448;
wire n_17449;
wire n_17450;
wire n_17451;
wire n_17452;
wire n_17453;
wire n_17454;
wire n_17455;
wire n_17456;
wire n_17457;
wire n_17458;
wire n_17459;
wire n_17460;
wire n_17461;
wire n_17462;
wire n_17463;
wire n_17464;
wire n_17465;
wire n_17466;
wire n_17467;
wire n_17468;
wire n_17469;
wire n_17470;
wire n_17471;
wire n_17472;
wire n_17473;
wire n_17474;
wire n_17475;
wire n_17476;
wire n_17477;
wire n_17478;
wire n_17479;
wire n_17480;
wire n_17481;
wire n_17482;
wire n_17483;
wire n_17484;
wire n_17485;
wire n_17486;
wire n_17487;
wire n_17488;
wire n_17489;
wire n_17490;
wire n_17491;
wire n_17492;
wire n_17493;
wire n_17494;
wire n_17495;
wire n_17496;
wire n_17497;
wire n_17498;
wire n_17499;
wire n_17500;
wire n_17501;
wire n_17502;
wire n_17503;
wire n_17504;
wire n_17505;
wire n_17506;
wire n_17507;
wire n_17508;
wire n_17509;
wire n_17510;
wire n_17511;
wire n_17512;
wire n_17513;
wire n_17514;
wire n_17515;
wire n_17516;
wire n_17517;
wire n_17518;
wire n_17519;
wire n_17520;
wire n_17521;
wire n_17522;
wire n_17523;
wire n_17524;
wire n_17525;
wire n_17526;
wire n_17527;
wire n_17528;
wire n_17529;
wire n_17530;
wire n_17531;
wire n_17532;
wire n_17533;
wire n_17534;
wire n_17535;
wire n_17536;
wire n_17537;
wire n_17538;
wire n_17539;
wire n_17540;
wire n_17541;
wire n_17542;
wire n_17543;
wire n_17544;
wire n_17545;
wire n_17546;
wire n_17547;
wire n_17548;
wire n_17549;
wire n_17550;
wire n_17551;
wire n_17552;
wire n_17553;
wire n_17554;
wire n_17555;
wire n_17556;
wire n_17557;
wire n_17558;
wire n_17559;
wire n_17560;
wire n_17561;
wire n_17562;
wire n_17563;
wire n_17564;
wire n_17565;
wire n_17566;
wire n_17567;
wire n_17568;
wire n_17569;
wire n_17570;
wire n_17571;
wire n_17572;
wire n_17573;
wire n_17574;
wire n_17575;
wire n_17576;
wire n_17577;
wire n_17578;
wire n_17579;
wire n_17580;
wire n_17581;
wire n_17582;
wire n_17583;
wire n_17584;
wire n_17585;
wire n_17586;
wire n_17587;
wire n_17588;
wire n_17589;
wire n_17590;
wire n_17591;
wire n_17592;
wire n_17593;
wire n_17594;
wire n_17595;
wire n_17596;
wire n_17597;
wire n_17598;
wire n_17599;
wire n_17600;
wire n_17601;
wire n_17602;
wire n_17603;
wire n_17604;
wire n_17605;
wire n_17606;
wire n_17607;
wire n_17608;
wire n_17609;
wire n_17610;
wire n_17611;
wire n_17612;
wire n_17613;
wire n_17614;
wire n_17615;
wire n_17616;
wire n_17617;
wire n_17618;
wire n_17619;
wire n_17620;
wire n_17621;
wire n_17622;
wire n_17623;
wire n_17624;
wire n_17625;
wire n_17626;
wire n_17627;
wire n_17628;
wire n_17629;
wire n_17630;
wire n_17631;
wire n_17632;
wire n_17633;
wire n_17634;
wire n_17635;
wire n_17636;
wire n_17637;
wire n_17638;
wire n_17639;
wire n_17640;
wire n_17641;
wire n_17642;
wire n_17643;
wire n_17644;
wire n_17645;
wire n_17646;
wire n_17647;
wire n_17648;
wire n_17649;
wire n_17650;
wire n_17651;
wire n_17652;
wire n_17653;
wire n_17654;
wire n_17655;
wire n_17656;
wire n_17657;
wire n_17658;
wire n_17659;
wire n_17660;
wire n_17661;
wire n_17662;
wire n_17663;
wire n_17664;
wire n_17665;
wire n_17666;
wire n_17667;
wire n_17668;
wire n_17669;
wire n_17670;
wire n_17671;
wire n_17672;
wire n_17673;
wire n_17674;
wire n_17675;
wire n_17676;
wire n_17677;
wire n_17678;
wire n_17679;
wire n_17680;
wire n_17681;
wire n_17682;
wire n_17683;
wire n_17684;
wire n_17685;
wire n_17686;
wire n_17687;
wire n_17688;
wire n_17689;
wire n_17690;
wire n_17691;
wire n_17692;
wire n_17693;
wire n_17694;
wire n_17695;
wire n_17696;
wire n_17697;
wire n_17698;
wire n_17699;
wire n_17700;
wire n_17701;
wire n_17702;
wire n_17703;
wire n_17704;
wire n_17705;
wire n_17706;
wire n_17707;
wire n_17708;
wire n_17709;
wire n_17710;
wire n_17711;
wire n_17712;
wire n_17713;
wire n_17714;
wire n_17715;
wire n_17716;
wire n_17717;
wire n_17718;
wire n_17719;
wire n_17720;
wire n_17721;
wire n_17722;
wire n_17723;
wire n_17724;
wire n_17725;
wire n_17726;
wire n_17727;
wire n_17728;
wire n_17729;
wire n_17730;
wire n_17731;
wire n_17732;
wire n_17733;
wire n_17734;
wire n_17735;
wire n_17736;
wire n_17737;
wire n_17738;
wire n_17739;
wire n_17740;
wire n_17741;
wire n_17742;
wire n_17743;
wire n_17744;
wire n_17745;
wire n_17746;
wire n_17747;
wire n_17748;
wire n_17749;
wire n_17750;
wire n_17751;
wire n_17752;
wire n_17753;
wire n_17754;
wire n_17755;
wire n_17756;
wire n_17757;
wire n_17758;
wire n_17759;
wire n_17760;
wire n_17761;
wire n_17762;
wire n_17763;
wire n_17764;
wire n_17765;
wire n_17766;
wire n_17767;
wire n_17768;
wire n_17769;
wire n_17770;
wire n_17771;
wire n_17772;
wire n_17773;
wire n_17774;
wire n_17775;
wire n_17776;
wire n_17777;
wire n_17778;
wire n_17779;
wire n_17780;
wire n_17781;
wire n_17782;
wire n_17783;
wire n_17784;
wire n_17785;
wire n_17786;
wire n_17787;
wire n_17788;
wire n_17789;
wire n_17790;
wire n_17791;
wire n_17792;
wire n_17793;
wire n_17794;
wire n_17795;
wire n_17796;
wire n_17797;
wire n_17798;
wire n_17799;
wire n_17800;
wire n_17801;
wire n_17802;
wire n_17803;
wire n_17804;
wire n_17805;
wire n_17806;
wire n_17807;
wire n_17808;
wire n_17809;
wire n_17810;
wire n_17811;
wire n_17812;
wire n_17813;
wire n_17814;
wire n_17815;
wire n_17816;
wire n_17817;
wire n_17818;
wire n_17819;
wire n_17820;
wire n_17821;
wire n_17822;
wire n_17823;
wire n_17824;
wire n_17825;
wire n_17826;
wire n_17827;
wire n_17828;
wire n_17829;
wire n_17830;
wire n_17831;
wire n_17832;
wire n_17833;
wire n_17834;
wire n_17835;
wire n_17836;
wire n_17837;
wire n_17838;
wire n_17839;
wire n_17840;
wire n_17841;
wire n_17842;
wire n_17843;
wire n_17844;
wire n_17845;
wire n_17846;
wire n_17847;
wire n_17848;
wire n_17849;
wire n_17850;
wire n_17851;
wire n_17852;
wire n_17853;
wire n_17854;
wire n_17855;
wire n_17856;
wire n_17857;
wire n_17858;
wire n_17859;
wire n_17860;
wire n_17861;
wire n_17862;
wire n_17863;
wire n_17864;
wire n_17865;
wire n_17866;
wire n_17867;
wire n_17868;
wire n_17869;
wire n_17870;
wire n_17871;
wire n_17872;
wire n_17873;
wire n_17874;
wire n_17875;
wire n_17876;
wire n_17877;
wire n_17878;
wire n_17879;
wire n_17880;
wire n_17881;
wire n_17882;
wire n_17883;
wire n_17884;
wire n_17885;
wire n_17886;
wire n_17887;
wire n_17888;
wire n_17889;
wire n_17890;
wire n_17891;
wire n_17892;
wire n_17893;
wire n_17894;
wire n_17895;
wire n_17896;
wire n_17897;
wire n_17898;
wire n_17899;
wire n_17900;
wire n_17901;
wire n_17902;
wire n_17903;
wire n_17904;
wire n_17905;
wire n_17906;
wire n_17907;
wire n_17908;
wire n_17909;
wire n_17910;
wire n_17911;
wire n_17912;
wire n_17913;
wire n_17914;
wire n_17915;
wire n_17916;
wire n_17917;
wire n_17918;
wire n_17919;
wire n_17920;
wire n_17921;
wire n_17922;
wire n_17923;
wire n_17924;
wire n_17925;
wire n_17926;
wire n_17927;
wire n_17928;
wire n_17929;
wire n_17930;
wire n_17931;
wire n_17932;
wire n_17933;
wire n_17934;
wire n_17935;
wire n_17936;
wire n_17937;
wire n_17938;
wire n_17939;
wire n_17940;
wire n_17941;
wire n_17942;
wire n_17943;
wire n_17944;
wire n_17945;
wire n_17946;
wire n_17947;
wire n_17948;
wire n_17949;
wire n_17950;
wire n_17951;
wire n_17952;
wire n_17953;
wire n_17954;
wire n_17955;
wire n_17956;
wire n_17957;
wire n_17958;
wire n_17959;
wire n_17960;
wire n_17961;
wire n_17962;
wire n_17963;
wire n_17964;
wire n_17965;
wire n_17966;
wire n_17967;
wire n_17968;
wire n_17969;
wire n_17970;
wire n_17971;
wire n_17972;
wire n_17973;
wire n_17974;
wire n_17975;
wire n_17976;
wire n_17977;
wire n_17978;
wire n_17979;
wire n_17980;
wire n_17981;
wire n_17982;
wire n_17983;
wire n_17984;
wire n_17985;
wire n_17986;
wire n_17987;
wire n_17988;
wire n_17989;
wire n_17990;
wire n_17991;
wire n_17992;
wire n_17993;
wire n_17994;
wire n_17995;
wire n_17996;
wire n_17997;
wire n_17998;
wire n_17999;
wire n_18000;
wire n_18001;
wire n_18002;
wire n_18003;
wire n_18004;
wire n_18005;
wire n_18006;
wire n_18007;
wire n_18008;
wire n_18009;
wire n_18010;
wire n_18011;
wire n_18012;
wire n_18013;
wire n_18014;
wire n_18015;
wire n_18016;
wire n_18017;
wire n_18018;
wire n_18019;
wire n_18020;
wire n_18021;
wire n_18022;
wire n_18023;
wire n_18024;
wire n_18025;
wire n_18026;
wire n_18027;
wire n_18028;
wire n_18029;
wire n_18030;
wire n_18031;
wire n_18032;
wire n_18033;
wire n_18034;
wire n_18035;
wire n_18036;
wire n_18037;
wire n_18038;
wire n_18039;
wire n_18040;
wire n_18041;
wire n_18042;
wire n_18043;
wire n_18044;
wire n_18045;
wire n_18046;
wire n_18047;
wire n_18048;
wire n_18049;
wire n_18050;
wire n_18051;
wire n_18052;
wire n_18053;
wire n_18054;
wire n_18055;
wire n_18056;
wire n_18057;
wire n_18058;
wire n_18059;
wire n_18060;
wire n_18061;
wire n_18062;
wire n_18063;
wire n_18064;
wire n_18065;
wire n_18066;
wire n_18067;
wire n_18068;
wire n_18069;
wire n_18070;
wire n_18071;
wire n_18072;
wire n_18073;
wire n_18074;
wire n_18075;
wire n_18076;
wire n_18077;
wire n_18078;
wire n_18079;
wire n_18080;
wire n_18081;
wire n_18082;
wire n_18083;
wire n_18084;
wire n_18085;
wire n_18086;
wire n_18087;
wire n_18088;
wire n_18089;
wire n_18090;
wire n_18091;
wire n_18092;
wire n_18093;
wire n_18094;
wire n_18095;
wire n_18096;
wire n_18097;
wire n_18098;
wire n_18099;
wire n_18100;
wire n_18101;
wire n_18102;
wire n_18103;
wire n_18104;
wire n_18105;
wire n_18106;
wire n_18107;
wire n_18108;
wire n_18109;
wire n_18110;
wire n_18111;
wire n_18112;
wire n_18113;
wire n_18114;
wire n_18115;
wire n_18116;
wire n_18117;
wire n_18118;
wire n_18119;
wire n_18120;
wire n_18121;
wire n_18122;
wire n_18123;
wire n_18124;
wire n_18125;
wire n_18126;
wire n_18127;
wire n_18128;
wire n_18129;
wire n_18130;
wire n_18131;
wire n_18132;
wire n_18133;
wire n_18134;
wire n_18135;
wire n_18136;
wire n_18137;
wire n_18138;
wire n_18139;
wire n_18140;
wire n_18141;
wire n_18142;
wire n_18143;
wire n_18144;
wire n_18145;
wire n_18146;
wire n_18147;
wire n_18148;
wire n_18149;
wire n_18150;
wire n_18151;
wire n_18152;
wire n_18153;
wire n_18154;
wire n_18155;
wire n_18156;
wire n_18157;
wire n_18158;
wire n_18159;
wire n_18160;
wire n_18161;
wire n_18162;
wire n_18163;
wire n_18164;
wire n_18165;
wire n_18166;
wire n_18167;
wire n_18168;
wire n_18169;
wire n_18170;
wire n_18171;
wire n_18172;
wire n_18173;
wire n_18174;
wire n_18175;
wire n_18176;
wire n_18177;
wire n_18178;
wire n_18179;
wire n_18180;
wire n_18181;
wire n_18182;
wire n_18183;
wire n_18184;
wire n_18185;
wire n_18186;
wire n_18187;
wire n_18188;
wire n_18189;
wire n_18190;
wire n_18191;
wire n_18192;
wire n_18193;
wire n_18194;
wire n_18195;
wire n_18196;
wire n_18197;
wire n_18198;
wire n_18199;
wire n_18200;
wire n_18201;
wire n_18202;
wire n_18203;
wire n_18204;
wire n_18205;
wire n_18206;
wire n_18207;
wire n_18208;
wire n_18209;
wire n_18210;
wire n_18211;
wire n_18212;
wire n_18213;
wire n_18214;
wire n_18215;
wire n_18216;
wire n_18217;
wire n_18218;
wire n_18219;
wire n_18220;
wire n_18221;
wire n_18222;
wire n_18223;
wire n_18224;
wire n_18225;
wire n_18226;
wire n_18227;
wire n_18228;
wire n_18229;
wire n_18230;
wire n_18231;
wire n_18232;
wire n_18233;
wire n_18234;
wire n_18235;
wire n_18236;
wire n_18237;
wire n_18238;
wire n_18239;
wire n_18240;
wire n_18241;
wire n_18242;
wire n_18243;
wire n_18244;
wire n_18245;
wire n_18246;
wire n_18247;
wire n_18248;
wire n_18249;
wire n_18250;
wire n_18251;
wire n_18252;
wire n_18253;
wire n_18254;
wire n_18255;
wire n_18256;
wire n_18257;
wire n_18258;
wire n_18259;
wire n_18260;
wire n_18261;
wire n_18262;
wire n_18263;
wire n_18264;
wire n_18265;
wire n_18266;
wire n_18267;
wire n_18268;
wire n_18269;
wire n_18270;
wire n_18271;
wire n_18272;
wire n_18273;
wire n_18274;
wire n_18275;
wire n_18276;
wire n_18277;
wire n_18278;
wire n_18279;
wire n_18280;
wire n_18281;
wire n_18282;
wire n_18283;
wire n_18284;
wire n_18285;
wire n_18286;
wire n_18287;
wire n_18288;
wire n_18289;
wire n_18290;
wire n_18291;
wire n_18292;
wire n_18293;
wire n_18294;
wire n_18295;
wire n_18296;
wire n_18297;
wire n_18298;
wire n_18299;
wire n_18300;
wire n_18301;
wire n_18302;
wire n_18303;
wire n_18304;
wire n_18305;
wire n_18306;
wire n_18307;
wire n_18308;
wire n_18309;
wire n_18310;
wire n_18311;
wire n_18312;
wire n_18313;
wire n_18314;
wire n_18315;
wire n_18316;
wire n_18317;
wire n_18318;
wire n_18319;
wire n_18320;
wire n_18321;
wire n_18322;
wire n_18323;
wire n_18324;
wire n_18325;
wire n_18326;
wire n_18327;
wire n_18328;
wire n_18329;
wire n_18330;
wire n_18331;
wire n_18332;
wire n_18333;
wire n_18334;
wire n_18335;
wire n_18336;
wire n_18337;
wire n_18338;
wire n_18339;
wire n_18340;
wire n_18341;
wire n_18342;
wire n_18343;
wire n_18344;
wire n_18345;
wire n_18346;
wire n_18347;
wire n_18348;
wire n_18349;
wire n_18350;
wire n_18351;
wire n_18352;
wire n_18353;
wire n_18354;
wire n_18355;
wire n_18356;
wire n_18357;
wire n_18358;
wire n_18359;
wire n_18360;
wire n_18361;
wire n_18362;
wire n_18363;
wire n_18364;
wire n_18365;
wire n_18366;
wire n_18367;
wire n_18368;
wire n_18369;
wire n_18370;
wire n_18371;
wire n_18372;
wire n_18373;
wire n_18374;
wire n_18375;
wire n_18376;
wire n_18377;
wire n_18378;
wire n_18379;
wire n_18380;
wire n_18381;
wire n_18382;
wire n_18383;
wire n_18384;
wire n_18385;
wire n_18386;
wire n_18387;
wire n_18388;
wire n_18389;
wire n_18390;
wire n_18391;
wire n_18392;
wire n_18393;
wire n_18394;
wire n_18395;
wire n_18396;
wire n_18397;
wire n_18398;
wire n_18399;
wire n_18400;
wire n_18401;
wire n_18402;
wire n_18403;
wire n_18404;
wire n_18405;
wire n_18406;
wire n_18407;
wire n_18408;
wire n_18409;
wire n_18410;
wire n_18411;
wire n_18412;
wire n_18413;
wire n_18414;
wire n_18415;
wire n_18416;
wire n_18417;
wire n_18418;
wire n_18419;
wire n_18420;
wire n_18421;
wire n_18422;
wire n_18423;
wire n_18424;
wire n_18425;
wire n_18426;
wire n_18427;
wire n_18428;
wire n_18429;
wire n_18430;
wire n_18431;
wire n_18432;
wire n_18433;
wire n_18434;
wire n_18435;
wire n_18436;
wire n_18437;
wire n_18438;
wire n_18439;
wire n_18440;
wire n_18441;
wire n_18442;
wire n_18443;
wire n_18444;
wire n_18445;
wire n_18446;
wire n_18447;
wire n_18448;
wire n_18449;
wire n_18450;
wire n_18451;
wire n_18452;
wire n_18453;
wire n_18454;
wire n_18455;
wire n_18456;
wire n_18457;
wire n_18458;
wire n_18459;
wire n_18460;
wire n_18461;
wire n_18462;
wire n_18463;
wire n_18464;
wire n_18465;
wire n_18466;
wire n_18467;
wire n_18468;
wire n_18469;
wire n_18470;
wire n_18471;
wire n_18472;
wire n_18473;
wire n_18474;
wire n_18475;
wire n_18476;
wire n_18477;
wire n_18478;
wire n_18479;
wire n_18480;
wire n_18481;
wire n_18482;
wire n_18483;
wire n_18484;
wire n_18485;
wire n_18486;
wire n_18487;
wire n_18488;
wire n_18489;
wire n_18490;
wire n_18491;
wire n_18492;
wire n_18493;
wire n_18494;
wire n_18495;
wire n_18496;
wire n_18497;
wire n_18498;
wire n_18499;
wire n_18500;
wire n_18501;
wire n_18502;
wire n_18503;
wire n_18504;
wire n_18505;
wire n_18506;
wire n_18507;
wire n_18508;
wire n_18509;
wire n_18510;
wire n_18511;
wire n_18512;
wire n_18513;
wire n_18514;
wire n_18515;
wire n_18516;
wire n_18517;
wire n_18518;
wire n_18519;
wire n_18520;
wire n_18521;
wire n_18522;
wire n_18523;
wire n_18524;
wire n_18525;
wire n_18526;
wire n_18527;
wire n_18528;
wire n_18529;
wire n_18530;
wire n_18531;
wire n_18532;
wire n_18533;
wire n_18534;
wire n_18535;
wire n_18536;
wire n_18537;
wire n_18538;
wire n_18539;
wire n_18540;
wire n_18541;
wire n_18542;
wire n_18543;
wire n_18544;
wire n_18545;
wire n_18546;
wire n_18547;
wire n_18548;
wire n_18549;
wire n_18550;
wire n_18551;
wire n_18552;
wire n_18553;
wire n_18554;
wire n_18555;
wire n_18556;
wire n_18557;
wire n_18558;
wire n_18559;
wire n_18560;
wire n_18561;
wire n_18562;
wire n_18563;
wire n_18564;
wire n_18565;
wire n_18566;
wire n_18567;
wire n_18568;
wire n_18569;
wire n_18570;
wire n_18571;
wire n_18572;
wire n_18573;
wire n_18574;
wire n_18575;
wire n_18576;
wire n_18577;
wire n_18578;
wire n_18579;
wire n_18580;
wire n_18581;
wire n_18582;
wire n_18583;
wire n_18584;
wire n_18585;
wire n_18586;
wire n_18587;
wire n_18588;
wire n_18589;
wire n_18590;
wire n_18591;
wire n_18592;
wire n_18593;
wire n_18594;
wire n_18595;
wire n_18596;
wire n_18597;
wire n_18598;
wire n_18599;
wire n_18600;
wire n_18601;
wire n_18602;
wire n_18603;
wire n_18604;
wire n_18605;
wire n_18606;
wire n_18607;
wire n_18608;
wire n_18609;
wire n_18610;
wire n_18611;
wire n_18612;
wire n_18613;
wire n_18614;
wire n_18615;
wire n_18616;
wire n_18617;
wire n_18618;
wire n_18619;
wire n_18620;
wire n_18621;
wire n_18622;
wire n_18623;
wire n_18624;
wire n_18625;
wire n_18626;
wire n_18627;
wire n_18628;
wire n_18629;
wire n_18630;
wire n_18631;
wire n_18632;
wire n_18633;
wire n_18634;
wire n_18635;
wire n_18636;
wire n_18637;
wire n_18638;
wire n_18639;
wire n_18640;
wire n_18641;
wire n_18642;
wire n_18643;
wire n_18644;
wire n_18645;
wire n_18646;
wire n_18647;
wire n_18648;
wire n_18649;
wire n_18650;
wire n_18651;
wire n_18652;
wire n_18653;
wire n_18654;
wire n_18655;
wire n_18656;
wire n_18657;
wire n_18658;
wire n_18659;
wire n_18660;
wire n_18661;
wire n_18662;
wire n_18663;
wire n_18664;
wire n_18665;
wire n_18666;
wire n_18667;
wire n_18668;
wire n_18669;
wire n_18670;
wire n_18671;
wire n_18672;
wire n_18673;
wire n_18674;
wire n_18675;
wire n_18676;
wire n_18677;
wire n_18678;
wire n_18679;
wire n_18680;
wire n_18681;
wire n_18682;
wire n_18683;
wire n_18684;
wire n_18685;
wire n_18686;
wire n_18687;
wire n_18688;
wire n_18689;
wire n_18690;
wire n_18691;
wire n_18692;
wire n_18693;
wire n_18694;
wire n_18695;
wire n_18696;
wire n_18697;
wire n_18698;
wire n_18699;
wire n_18700;
wire n_18701;
wire n_18702;
wire n_18703;
wire n_18704;
wire n_18705;
wire n_18706;
wire n_18707;
wire n_18708;
wire n_18709;
wire n_18710;
wire n_18711;
wire n_18712;
wire n_18713;
wire n_18714;
wire n_18715;
wire n_18716;
wire n_18717;
wire n_18718;
wire n_18719;
wire n_18720;
wire n_18721;
wire n_18722;
wire n_18723;
wire n_18724;
wire n_18725;
wire n_18726;
wire n_18727;
wire n_18728;
wire n_18729;
wire n_18730;
wire n_18731;
wire n_18732;
wire n_18733;
wire n_18734;
wire n_18735;
wire n_18736;
wire n_18737;
wire n_18738;
wire n_18739;
wire n_18740;
wire n_18741;
wire n_18742;
wire n_18743;
wire n_18744;
wire n_18745;
wire n_18746;
wire n_18747;
wire n_18748;
wire n_18749;
wire n_18750;
wire n_18751;
wire n_18752;
wire n_18753;
wire n_18754;
wire n_18755;
wire n_18756;
wire n_18757;
wire n_18758;
wire n_18759;
wire n_18760;
wire n_18761;
wire n_18762;
wire n_18763;
wire n_18764;
wire n_18765;
wire n_18766;
wire n_18767;
wire n_18768;
wire n_18769;
wire n_18770;
wire n_18771;
wire n_18772;
wire n_18773;
wire n_18774;
wire n_18775;
wire n_18776;
wire n_18777;
wire n_18778;
wire n_18779;
wire n_18780;
wire n_18781;
wire n_18782;
wire n_18783;
wire n_18784;
wire n_18785;
wire n_18786;
wire n_18787;
wire n_18788;
wire n_18789;
wire n_18790;
wire n_18791;
wire n_18792;
wire n_18793;
wire n_18794;
wire n_18795;
wire n_18796;
wire n_18797;
wire n_18798;
wire n_18799;
wire n_18800;
wire n_18801;
wire n_18802;
wire n_18803;
wire n_18804;
wire n_18805;
wire n_18806;
wire n_18807;
wire n_18808;
wire n_18809;
wire n_18810;
wire n_18811;
wire n_18812;
wire n_18813;
wire n_18814;
wire n_18815;
wire n_18816;
wire n_18817;
wire n_18818;
wire n_18819;
wire n_18820;
wire n_18821;
wire n_18822;
wire n_18823;
wire n_18824;
wire n_18825;
wire n_18826;
wire n_18827;
wire n_18828;
wire n_18829;
wire n_18830;
wire n_18831;
wire n_18832;
wire n_18833;
wire n_18834;
wire n_18835;
wire n_18836;
wire n_18837;
wire n_18838;
wire n_18839;
wire n_18840;
wire n_18841;
wire n_18842;
wire n_18843;
wire n_18844;
wire n_18845;
wire n_18846;
wire n_18847;
wire n_18848;
wire n_18849;
wire n_18850;
wire n_18851;
wire n_18852;
wire n_18853;
wire n_18854;
wire n_18855;
wire n_18856;
wire n_18857;
wire n_18858;
wire n_18859;
wire n_18860;
wire n_18861;
wire n_18862;
wire n_18863;
wire n_18864;
wire n_18865;
wire n_18866;
wire n_18867;
wire n_18868;
wire n_18869;
wire n_18870;
wire n_18871;
wire n_18872;
wire n_18873;
wire n_18874;
wire n_18875;
wire n_18876;
wire n_18877;
wire n_18878;
wire n_18879;
wire n_18880;
wire n_18881;
wire n_18882;
wire n_18883;
wire n_18884;
wire n_18885;
wire n_18886;
wire n_18887;
wire n_18888;
wire n_18889;
wire n_18890;
wire n_18891;
wire n_18892;
wire n_18893;
wire n_18894;
wire n_18895;
wire n_18896;
wire n_18897;
wire n_18898;
wire n_18899;
wire n_18900;
wire n_18901;
wire n_18902;
wire n_18903;
wire n_18904;
wire n_18905;
wire n_18906;
wire n_18907;
wire n_18908;
wire n_18909;
wire n_18910;
wire n_18911;
wire n_18912;
wire n_18913;
wire n_18914;
wire n_18915;
wire n_18916;
wire n_18917;
wire n_18918;
wire n_18919;
wire n_18920;
wire n_18921;
wire n_18922;
wire n_18923;
wire n_18924;
wire n_18925;
wire n_18926;
wire n_18927;
wire n_18928;
wire n_18929;
wire n_18930;
wire n_18931;
wire n_18932;
wire n_18933;
wire n_18934;
wire n_18935;
wire n_18936;
wire n_18937;
wire n_18938;
wire n_18939;
wire n_18940;
wire n_18941;
wire n_18942;
wire n_18943;
wire n_18944;
wire n_18945;
wire n_18946;
wire n_18947;
wire n_18948;
wire n_18949;
wire n_18950;
wire n_18951;
wire n_18952;
wire n_18953;
wire n_18954;
wire n_18955;
wire n_18956;
wire n_18957;
wire n_18958;
wire n_18959;
wire n_18960;
wire n_18961;
wire n_18962;
wire n_18963;
wire n_18964;
wire n_18965;
wire n_18966;
wire n_18967;
wire n_18968;
wire n_18969;
wire n_18970;
wire n_18971;
wire n_18972;
wire n_18973;
wire n_18974;
wire n_18975;
wire n_18976;
wire n_18977;
wire n_18978;
wire n_18979;
wire n_18980;
wire n_18981;
wire n_18982;
wire n_18983;
wire n_18984;
wire n_18985;
wire n_18986;
wire n_18987;
wire n_18988;
wire n_18989;
wire n_18990;
wire n_18991;
wire n_18992;
wire n_18993;
wire n_18994;
wire n_18995;
wire n_18996;
wire n_18997;
wire n_18998;
wire n_18999;
wire n_19000;
wire n_19001;
wire n_19002;
wire n_19003;
wire n_19004;
wire n_19005;
wire n_19006;
wire n_19007;
wire n_19008;
wire n_19009;
wire n_19010;
wire n_19011;
wire n_19012;
wire n_19013;
wire n_19014;
wire n_19015;
wire n_19016;
wire n_19017;
wire n_19018;
wire n_19019;
wire n_19020;
wire n_19021;
wire n_19022;
wire n_19023;
wire n_19024;
wire n_19025;
wire n_19026;
wire n_19027;
wire n_19028;
wire n_19029;
wire n_19030;
wire n_19031;
wire n_19032;
wire n_19033;
wire n_19034;
wire n_19035;
wire n_19036;
wire n_19037;
wire n_19038;
wire n_19039;
wire n_19040;
wire n_19041;
wire n_19042;
wire n_19043;
wire n_19044;
wire n_19045;
wire n_19046;
wire n_19047;
wire n_19048;
wire n_19049;
wire n_19050;
wire n_19051;
wire n_19052;
wire n_19053;
wire n_19054;
wire n_19055;
wire n_19056;
wire n_19057;
wire n_19058;
wire n_19059;
wire n_19060;
wire n_19061;
wire n_19062;
wire n_19063;
wire n_19064;
wire n_19065;
wire n_19066;
wire n_19067;
wire n_19068;
wire n_19069;
wire n_19070;
wire n_19071;
wire n_19072;
wire n_19073;
wire n_19074;
wire n_19075;
wire n_19076;
wire n_19077;
wire n_19078;
wire n_19079;
wire n_19080;
wire n_19081;
wire n_19082;
wire n_19083;
wire n_19084;
wire n_19085;
wire n_19086;
wire n_19087;
wire n_19088;
wire n_19089;
wire n_19090;
wire n_19091;
wire n_19092;
wire n_19093;
wire n_19094;
wire n_19095;
wire n_19096;
wire n_19097;
wire n_19098;
wire n_19099;
wire n_19100;
wire n_19101;
wire n_19102;
wire n_19103;
wire n_19104;
wire n_19105;
wire n_19106;
wire n_19107;
wire n_19108;
wire n_19109;
wire n_19110;
wire n_19111;
wire n_19112;
wire n_19113;
wire n_19114;
wire n_19115;
wire n_19116;
wire n_19117;
wire n_19118;
wire n_19119;
wire n_19120;
wire n_19121;
wire n_19122;
wire n_19123;
wire n_19124;
wire n_19125;
wire n_19126;
wire n_19127;
wire n_19128;
wire n_19129;
wire n_19130;
wire n_19131;
wire n_19132;
wire n_19133;
wire n_19134;
wire n_19135;
wire n_19136;
wire n_19137;
wire n_19138;
wire n_19139;
wire n_19140;
wire n_19141;
wire n_19142;
wire n_19143;
wire n_19144;
wire n_19145;
wire n_19146;
wire n_19147;
wire n_19148;
wire n_19149;
wire n_19150;
wire n_19151;
wire n_19152;
wire n_19153;
wire n_19154;
wire n_19155;
wire n_19156;
wire n_19157;
wire n_19158;
wire n_19159;
wire n_19160;
wire n_19161;
wire n_19162;
wire n_19163;
wire n_19164;
wire n_19165;
wire n_19166;
wire n_19167;
wire n_19168;
wire n_19169;
wire n_19170;
wire n_19171;
wire n_19172;
wire n_19173;
wire n_19174;
wire n_19175;
wire n_19176;
wire n_19177;
wire n_19178;
wire n_19179;
wire n_19180;
wire n_19181;
wire n_19182;
wire n_19183;
wire n_19184;
wire n_19185;
wire n_19186;
wire n_19187;
wire n_19188;
wire n_19189;
wire n_19190;
wire n_19191;
wire n_19192;
wire n_19193;
wire n_19194;
wire n_19195;
wire n_19196;
wire n_19197;
wire n_19198;
wire n_19199;
wire n_19200;
wire n_19201;
wire n_19202;
wire n_19203;
wire n_19204;
wire n_19205;
wire n_19206;
wire n_19207;
wire n_19208;
wire n_19209;
wire n_19210;
wire n_19211;
wire n_19212;
wire n_19213;
wire n_19214;
wire n_19215;
wire n_19216;
wire n_19217;
wire n_19218;
wire n_19219;
wire n_19220;
wire n_19221;
wire n_19222;
wire n_19223;
wire n_19224;
wire n_19225;
wire n_19226;
wire n_19227;
wire n_19228;
wire n_19229;
wire n_19230;
wire n_19231;
wire n_19232;
wire n_19233;
wire n_19234;
wire n_19235;
wire n_19236;
wire n_19237;
wire n_19238;
wire n_19239;
wire n_19240;
wire n_19241;
wire n_19242;
wire n_19243;
wire n_19244;
wire n_19245;
wire n_19246;
wire n_19247;
wire n_19248;
wire n_19249;
wire n_19250;
wire n_19251;
wire n_19252;
wire n_19253;
wire n_19254;
wire n_19255;
wire n_19256;
wire n_19257;
wire n_19258;
wire n_19259;
wire n_19260;
wire n_19261;
wire n_19262;
wire n_19263;
wire n_19264;
wire n_19265;
wire n_19266;
wire n_19267;
wire n_19268;
wire n_19269;
wire n_19270;
wire n_19271;
wire n_19272;
wire n_19273;
wire n_19274;
wire n_19275;
wire n_19276;
wire n_19277;
wire n_19278;
wire n_19279;
wire n_19280;
wire n_19281;
wire n_19282;
wire n_19283;
wire n_19284;
wire n_19285;
wire n_19286;
wire n_19287;
wire n_19288;
wire n_19289;
wire n_19290;
wire n_19291;
wire n_19292;
wire n_19293;
wire n_19294;
wire n_19295;
wire n_19296;
wire n_19297;
wire n_19298;
wire n_19299;
wire n_19300;
wire n_19301;
wire n_19302;
wire n_19303;
wire n_19304;
wire n_19305;
wire n_19306;
wire n_19307;
wire n_19308;
wire n_19309;
wire n_19310;
wire n_19311;
wire n_19312;
wire n_19313;
wire n_19314;
wire n_19315;
wire n_19316;
wire n_19317;
wire n_19318;
wire n_19319;
wire n_19320;
wire n_19321;
wire n_19322;
wire n_19323;
wire n_19324;
wire n_19325;
wire n_19326;
wire n_19327;
wire n_19328;
wire n_19329;
wire n_19330;
wire n_19331;
wire n_19332;
wire n_19333;
wire n_19334;
wire n_19335;
wire n_19336;
wire n_19337;
wire n_19338;
wire n_19339;
wire n_19340;
wire n_19341;
wire n_19342;
wire n_19343;
wire n_19344;
wire n_19345;
wire n_19346;
wire n_19347;
wire n_19348;
wire n_19349;
wire n_19350;
wire n_19351;
wire n_19352;
wire n_19353;
wire n_19354;
wire n_19355;
wire n_19356;
wire n_19357;
wire n_19358;
wire n_19359;
wire n_19360;
wire n_19361;
wire n_19362;
wire n_19363;
wire n_19364;
wire n_19365;
wire n_19366;
wire n_19367;
wire n_19368;
wire n_19369;
wire n_19370;
wire n_19371;
wire n_19372;
wire n_19373;
wire n_19374;
wire n_19375;
wire n_19376;
wire n_19377;
wire n_19378;
wire n_19379;
wire n_19380;
wire n_19381;
wire n_19382;
wire n_19383;
wire n_19384;
wire n_19385;
wire n_19386;
wire n_19387;
wire n_19388;
wire n_19389;
wire n_19390;
wire n_19391;
wire n_19392;
wire n_19393;
wire n_19394;
wire n_19395;
wire n_19396;
wire n_19397;
wire n_19398;
wire n_19399;
wire n_19400;
wire n_19401;
wire n_19402;
wire n_19403;
wire n_19404;
wire n_19405;
wire n_19406;
wire n_19407;
wire n_19408;
wire n_19409;
wire n_19410;
wire n_19411;
wire n_19412;
wire n_19413;
wire n_19414;
wire n_19415;
wire n_19416;
wire n_19417;
wire n_19418;
wire n_19419;
wire n_19420;
wire n_19421;
wire n_19422;
wire n_19423;
wire n_19424;
wire n_19425;
wire n_19426;
wire n_19427;
wire n_19428;
wire n_19429;
wire n_19430;
wire n_19431;
wire n_19432;
wire n_19433;
wire n_19434;
wire n_19435;
wire n_19436;
wire n_19437;
wire n_19438;
wire n_19439;
wire n_19440;
wire n_19441;
wire n_19442;
wire n_19443;
wire n_19444;
wire n_19445;
wire n_19446;
wire n_19447;
wire n_19448;
wire n_19449;
wire n_19450;
wire n_19451;
wire n_19452;
wire n_19453;
wire n_19454;
wire n_19455;
wire n_19456;
wire n_19457;
wire n_19458;
wire n_19459;
wire n_19460;
wire n_19461;
wire n_19462;
wire n_19463;
wire n_19464;
wire n_19465;
wire n_19466;
wire n_19467;
wire n_19468;
wire n_19469;
wire n_19470;
wire n_19471;
wire n_19472;
wire n_19473;
wire n_19474;
wire n_19475;
wire n_19476;
wire n_19477;
wire n_19478;
wire n_19479;
wire n_19480;
wire n_19481;
wire n_19482;
wire n_19483;
wire n_19484;
wire n_19485;
wire n_19486;
wire n_19487;
wire n_19488;
wire n_19489;
wire n_19490;
wire n_19491;
wire n_19492;
wire n_19493;
wire n_19494;
wire n_19495;
wire n_19496;
wire n_19497;
wire n_19498;
wire n_19499;
wire n_19500;
wire n_19501;
wire n_19502;
wire n_19503;
wire n_19504;
wire n_19505;
wire n_19506;
wire n_19507;
wire n_19508;
wire n_19509;
wire n_19510;
wire n_19511;
wire n_19512;
wire n_19513;
wire n_19514;
wire n_19515;
wire n_19516;
wire n_19517;
wire n_19518;
wire n_19519;
wire n_19520;
wire n_19521;
wire n_19522;
wire n_19523;
wire n_19524;
wire n_19525;
wire n_19526;
wire n_19527;
wire n_19528;
wire n_19529;
wire n_19530;
wire n_19531;
wire n_19532;
wire n_19533;
wire n_19534;
wire n_19535;
wire n_19536;
wire n_19537;
wire n_19538;
wire n_19539;
wire n_19540;
wire n_19541;
wire n_19542;
wire n_19543;
wire n_19544;
wire n_19545;
wire n_19546;
wire n_19547;
wire n_19548;
wire n_19549;
wire n_19550;
wire n_19551;
wire n_19552;
wire n_19553;
wire n_19554;
wire n_19555;
wire n_19556;
wire n_19557;
wire n_19558;
wire n_19559;
wire n_19560;
wire n_19561;
wire n_19562;
wire n_19563;
wire n_19564;
wire n_19565;
wire n_19566;
wire n_19567;
wire n_19568;
wire n_19569;
wire n_19570;
wire n_19571;
wire n_19572;
wire n_19573;
wire n_19574;
wire n_19575;
wire n_19576;
wire n_19577;
wire n_19578;
wire n_19579;
wire n_19580;
wire n_19581;
wire n_19582;
wire n_19583;
wire n_19584;
wire n_19585;
wire n_19586;
wire n_19587;
wire n_19588;
wire n_19589;
wire n_19590;
wire n_19591;
wire n_19592;
wire n_19593;
wire n_19594;
wire n_19595;
wire n_19596;
wire n_19597;
wire n_19598;
wire n_19599;
wire n_19600;
wire n_19601;
wire n_19602;
wire n_19603;
wire n_19604;
wire n_19605;
wire n_19606;
wire n_19607;
wire n_19608;
wire n_19609;
wire n_19610;
wire n_19611;
wire n_19612;
wire n_19613;
wire n_19614;
wire n_19615;
wire n_19616;
wire n_19617;
wire n_19618;
wire n_19619;
wire n_19620;
wire n_19621;
wire n_19622;
wire n_19623;
wire n_19624;
wire n_19625;
wire n_19626;
wire n_19627;
wire n_19628;
wire n_19629;
wire n_19630;
wire n_19631;
wire n_19632;
wire n_19633;
wire n_19634;
wire n_19635;
wire n_19636;
wire n_19637;
wire n_19638;
wire n_19639;
wire n_19640;
wire n_19641;
wire n_19642;
wire n_19643;
wire n_19644;
wire n_19645;
wire n_19646;
wire n_19647;
wire n_19648;
wire n_19649;
wire n_19650;
wire n_19651;
wire n_19652;
wire n_19653;
wire n_19654;
wire n_19655;
wire n_19656;
wire n_19657;
wire n_19658;
wire n_19659;
wire n_19660;
wire n_19661;
wire n_19662;
wire n_19663;
wire n_19664;
wire n_19665;
wire n_19666;
wire n_19667;
wire n_19668;
wire n_19669;
wire n_19670;
wire n_19671;
wire n_19672;
wire n_19673;
wire n_19674;
wire n_19675;
wire n_19676;
wire n_19677;
wire n_19678;
wire n_19679;
wire n_19680;
wire n_19681;
wire n_19682;
wire n_19683;
wire n_19684;
wire n_19685;
wire n_19686;
wire n_19687;
wire n_19688;
wire n_19689;
wire n_19690;
wire n_19691;
wire n_19692;
wire n_19693;
wire n_19694;
wire n_19695;
wire n_19696;
wire n_19697;
wire n_19698;
wire n_19699;
wire n_19700;
wire n_19701;
wire n_19702;
wire n_19703;
wire n_19704;
wire n_19705;
wire n_19706;
wire n_19707;
wire n_19708;
wire n_19709;
wire n_19710;
wire n_19711;
wire n_19712;
wire n_19713;
wire n_19714;
wire n_19715;
wire n_19716;
wire n_19717;
wire n_19718;
wire n_19719;
wire n_19720;
wire n_19721;
wire n_19722;
wire n_19723;
wire n_19724;
wire n_19725;
wire n_19726;
wire n_19727;
wire n_19728;
wire n_19729;
wire n_19730;
wire n_19731;
wire n_19732;
wire n_19733;
wire n_19734;
wire n_19735;
wire n_19736;
wire n_19737;
wire n_19738;
wire n_19739;
wire n_19740;
wire n_19741;
wire n_19742;
wire n_19743;
wire n_19744;
wire n_19745;
wire n_19746;
wire n_19747;
wire n_19748;
wire n_19749;
wire n_19750;
wire n_19751;
wire n_19752;
wire n_19753;
wire n_19754;
wire n_19755;
wire n_19756;
wire n_19757;
wire n_19758;
wire n_19759;
wire n_19760;
wire n_19761;
wire n_19762;
wire n_19763;
wire n_19764;
wire n_19765;
wire n_19766;
wire n_19767;
wire n_19768;
wire n_19769;
wire n_19770;
wire n_19771;
wire n_19772;
wire n_19773;
wire n_19774;
wire n_19775;
wire n_19776;
wire n_19777;
wire n_19778;
wire n_19779;
wire n_19780;
wire n_19781;
wire n_19782;
wire n_19783;
wire n_19784;
wire n_19785;
wire n_19786;
wire n_19787;
wire n_19788;
wire n_19789;
wire n_19790;
wire n_19791;
wire n_19792;
wire n_19793;
wire n_19794;
wire n_19795;
wire n_19796;
wire n_19797;
wire n_19798;
wire n_19799;
wire n_19800;
wire n_19801;
wire n_19802;
wire n_19803;
wire n_19804;
wire n_19805;
wire n_19806;
wire n_19807;
wire n_19808;
wire n_19809;
wire n_19810;
wire n_19811;
wire n_19812;
wire n_19813;
wire n_19814;
wire n_19815;
wire n_19816;
wire n_19817;
wire n_19818;
wire n_19819;
wire n_19820;
wire n_19821;
wire n_19822;
wire n_19823;
wire n_19824;
wire n_19825;
wire n_19826;
wire n_19827;
wire n_19828;
wire n_19829;
wire n_19830;
wire n_19831;
wire n_19832;
wire n_19833;
wire n_19834;
wire n_19835;
wire n_19836;
wire n_19837;
wire n_19838;
wire n_19839;
wire n_19840;
wire n_19841;
wire n_19842;
wire n_19843;
wire n_19844;
wire n_19845;
wire n_19846;
wire n_19847;
wire n_19848;
wire n_19849;
wire n_19850;
wire n_19851;
wire n_19852;
wire n_19853;
wire n_19854;
wire n_19855;
wire n_19856;
wire n_19857;
wire n_19858;
wire n_19859;
wire n_19860;
wire n_19861;
wire n_19862;
wire n_19863;
wire n_19864;
wire n_19865;
wire n_19866;
wire n_19867;
wire n_19868;
wire n_19869;
wire n_19870;
wire n_19871;
wire n_19872;
wire n_19873;
wire n_19874;
wire n_19875;
wire n_19876;
wire n_19877;
wire n_19878;
wire n_19879;
wire n_19880;
wire n_19881;
wire n_19882;
wire n_19883;
wire n_19884;
wire n_19885;
wire n_19886;
wire n_19887;
wire n_19888;
wire n_19889;
wire n_19890;
wire n_19891;
wire n_19892;
wire n_19893;
wire n_19894;
wire n_19895;
wire n_19896;
wire n_19897;
wire n_19898;
wire n_19899;
wire n_19900;
wire n_19901;
wire n_19902;
wire n_19903;
wire n_19904;
wire n_19905;
wire n_19906;
wire n_19907;
wire n_19908;
wire n_19909;
wire n_19910;
wire n_19911;
wire n_19912;
wire n_19913;
wire n_19914;
wire n_19915;
wire n_19916;
wire n_19917;
wire n_19918;
wire n_19919;
wire n_19920;
wire n_19921;
wire n_19922;
wire n_19923;
wire n_19924;
wire n_19925;
wire n_19926;
wire n_19927;
wire n_19928;
wire n_19929;
wire n_19930;
wire n_19931;
wire n_19932;
wire n_19933;
wire n_19934;
wire n_19935;
wire n_19936;
wire n_19937;
wire n_19938;
wire n_19939;
wire n_19940;
wire n_19941;
wire n_19942;
wire n_19943;
wire n_19944;
wire n_19945;
wire n_19946;
wire n_19947;
wire n_19948;
wire n_19949;
wire n_19950;
wire n_19951;
wire n_19952;
wire n_19953;
wire n_19954;
wire n_19955;
wire n_19956;
wire n_19957;
wire n_19958;
wire n_19959;
wire n_19960;
wire n_19961;
wire n_19962;
wire n_19963;
wire n_19964;
wire n_19965;
wire n_19966;
wire n_19967;
wire n_19968;
wire n_19969;
wire n_19970;
wire n_19971;
wire n_19972;
wire n_19973;
wire n_19974;
wire n_19975;
wire n_19976;
wire n_19977;
wire n_19978;
wire n_19979;
wire n_19980;
wire n_19981;
wire n_19982;
wire n_19983;
wire n_19984;
wire n_19985;
wire n_19986;
wire n_19987;
wire n_19988;
wire n_19989;
wire n_19990;
wire n_19991;
wire n_19992;
wire n_19993;
wire n_19994;
wire n_19995;
wire n_19996;
wire n_19997;
wire n_19998;
wire n_19999;
wire n_20000;
wire n_20001;
wire n_20002;
wire n_20003;
wire n_20004;
wire n_20005;
wire n_20006;
wire n_20007;
wire n_20008;
wire n_20009;
wire n_20010;
wire n_20011;
wire n_20012;
wire n_20013;
wire n_20014;
wire n_20015;
wire n_20016;
wire n_20017;
wire n_20018;
wire n_20019;
wire n_20020;
wire n_20021;
wire n_20022;
wire n_20023;
wire n_20024;
wire n_20025;
wire n_20026;
wire n_20027;
wire n_20028;
wire n_20029;
wire n_20030;
wire n_20031;
wire n_20032;
wire n_20033;
wire n_20034;
wire n_20035;
wire n_20036;
wire n_20037;
wire n_20038;
wire n_20039;
wire n_20040;
wire n_20041;
wire n_20042;
wire n_20043;
wire n_20044;
wire n_20045;
wire n_20046;
wire n_20047;
wire n_20048;
wire n_20049;
wire n_20050;
wire n_20051;
wire n_20052;
wire n_20053;
wire n_20054;
wire n_20055;
wire n_20056;
wire n_20057;
wire n_20058;
wire n_20059;
wire n_20060;
wire n_20061;
wire n_20062;
wire n_20063;
wire n_20064;
wire n_20065;
wire n_20066;
wire n_20067;
wire n_20068;
wire n_20069;
wire n_20070;
wire n_20071;
wire n_20072;
wire n_20073;
wire n_20074;
wire n_20075;
wire n_20076;
wire n_20077;
wire n_20078;
wire n_20079;
wire n_20080;
wire n_20081;
wire n_20082;
wire n_20083;
wire n_20084;
wire n_20085;
wire n_20086;
wire n_20087;
wire n_20088;
wire n_20089;
wire n_20090;
wire n_20091;
wire n_20092;
wire n_20093;
wire n_20094;
wire n_20095;
wire n_20096;
wire n_20097;
wire n_20098;
wire n_20099;
wire n_20100;
wire n_20101;
wire n_20102;
wire n_20103;
wire n_20104;
wire n_20105;
wire n_20106;
wire n_20107;
wire n_20108;
wire n_20109;
wire n_20110;
wire n_20111;
wire n_20112;
wire n_20113;
wire n_20114;
wire n_20115;
wire n_20116;
wire n_20117;
wire n_20118;
wire n_20119;
wire n_20120;
wire n_20121;
wire n_20122;
wire n_20123;
wire n_20124;
wire n_20125;
wire n_20126;
wire n_20127;
wire n_20128;
wire n_20129;
wire n_20130;
wire n_20131;
wire n_20132;
wire n_20133;
wire n_20134;
wire n_20135;
wire n_20136;
wire n_20137;
wire n_20138;
wire n_20139;
wire n_20140;
wire n_20141;
wire n_20142;
wire n_20143;
wire n_20144;
wire n_20145;
wire n_20146;
wire n_20147;
wire n_20148;
wire n_20149;
wire n_20150;
wire n_20151;
wire n_20152;
wire n_20153;
wire n_20154;
wire n_20155;
wire n_20156;
wire n_20157;
wire n_20158;
wire n_20159;
wire n_20160;
wire n_20161;
wire n_20162;
wire n_20163;
wire n_20164;
wire n_20165;
wire n_20166;
wire n_20167;
wire n_20168;
wire n_20169;
wire n_20170;
wire n_20171;
wire n_20172;
wire n_20173;
wire n_20174;
wire n_20175;
wire n_20176;
wire n_20177;
wire n_20178;
wire n_20179;
wire n_20180;
wire n_20181;
wire n_20182;
wire n_20183;
wire n_20184;
wire n_20185;
wire n_20186;
wire n_20187;
wire n_20188;
wire n_20189;
wire n_20190;
wire n_20191;
wire n_20192;
wire n_20193;
wire n_20194;
wire n_20195;
wire n_20196;
wire n_20197;
wire n_20198;
wire n_20199;
wire n_20200;
wire n_20201;
wire n_20202;
wire n_20203;
wire n_20204;
wire n_20205;
wire n_20206;
wire n_20207;
wire n_20208;
wire n_20209;
wire n_20210;
wire n_20211;
wire n_20212;
wire n_20213;
wire n_20214;
wire n_20215;
wire n_20216;
wire n_20217;
wire n_20218;
wire n_20219;
wire n_20220;
wire n_20221;
wire n_20222;
wire n_20223;
wire n_20224;
wire n_20225;
wire n_20226;
wire n_20227;
wire n_20228;
wire n_20229;
wire n_20230;
wire n_20231;
wire n_20232;
wire n_20233;
wire n_20234;
wire n_20235;
wire n_20236;
wire n_20237;
wire n_20238;
wire n_20239;
wire n_20240;
wire n_20241;
wire n_20242;
wire n_20243;
wire n_20244;
wire n_20245;
wire n_20246;
wire n_20247;
wire n_20248;
wire n_20249;
wire n_20250;
wire n_20251;
wire n_20252;
wire n_20253;
wire n_20254;
wire n_20255;
wire n_20256;
wire n_20257;
wire n_20258;
wire n_20259;
wire n_20260;
wire n_20261;
wire n_20262;
wire n_20263;
wire n_20264;
wire n_20265;
wire n_20266;
wire n_20267;
wire n_20268;
wire n_20269;
wire n_20270;
wire n_20271;
wire n_20272;
wire n_20273;
wire n_20274;
wire n_20275;
wire n_20276;
wire n_20277;
wire n_20278;
wire n_20279;
wire n_20280;
wire n_20281;
wire n_20282;
wire n_20283;
wire n_20284;
wire n_20285;
wire n_20286;
wire n_20287;
wire n_20288;
wire n_20289;
wire n_20290;
wire n_20291;
wire n_20292;
wire n_20293;
wire n_20294;
wire n_20295;
wire n_20296;
wire n_20297;
wire n_20298;
wire n_20299;
wire n_20300;
wire n_20301;
wire n_20302;
wire n_20303;
wire n_20304;
wire n_20305;
wire n_20306;
wire n_20307;
wire n_20308;
wire n_20309;
wire n_20310;
wire n_20311;
wire n_20312;
wire n_20313;
wire n_20314;
wire n_20315;
wire n_20316;
wire n_20317;
wire n_20318;
wire n_20319;
wire n_20320;
wire n_20321;
wire n_20322;
wire n_20323;
wire n_20324;
wire n_20325;
wire n_20326;
wire n_20327;
wire n_20328;
wire n_20329;
wire n_20330;
wire n_20331;
wire n_20332;
wire n_20333;
wire n_20334;
wire n_20335;
wire n_20336;
wire n_20337;
wire n_20338;
wire n_20339;
wire n_20340;
wire n_20341;
wire n_20342;
wire n_20343;
wire n_20344;
wire n_20345;
wire n_20346;
wire n_20347;
wire n_20348;
wire n_20349;
wire n_20350;
wire n_20351;
wire n_20352;
wire n_20353;
wire n_20354;
wire n_20355;
wire n_20356;
wire n_20357;
wire n_20358;
wire n_20359;
wire n_20360;
wire n_20361;
wire n_20362;
wire n_20363;
wire n_20364;
wire n_20365;
wire n_20366;
wire n_20367;
wire n_20368;
wire n_20369;
wire n_20370;
wire n_20371;
wire n_20372;
wire n_20373;
wire n_20374;
wire n_20375;
wire n_20376;
wire n_20377;
wire n_20378;
wire n_20379;
wire n_20380;
wire n_20381;
wire n_20382;
wire n_20383;
wire n_20384;
wire n_20385;
wire n_20386;
wire n_20387;
wire n_20388;
wire n_20389;
wire n_20390;
wire n_20391;
wire n_20392;
wire n_20393;
wire n_20394;
wire n_20395;
wire n_20396;
wire n_20397;
wire n_20398;
wire n_20399;
wire n_20400;
wire n_20401;
wire n_20402;
wire n_20403;
wire n_20404;
wire n_20405;
wire n_20406;
wire n_20407;
wire n_20408;
wire n_20409;
wire n_20410;
wire n_20411;
wire n_20412;
wire n_20413;
wire n_20414;
wire n_20415;
wire n_20416;
wire n_20417;
wire n_20418;
wire n_20419;
wire n_20420;
wire n_20421;
wire n_20422;
wire n_20423;
wire n_20424;
wire n_20425;
wire n_20426;
wire n_20427;
wire n_20428;
wire n_20429;
wire n_20430;
wire n_20431;
wire n_20432;
wire n_20433;
wire n_20434;
wire n_20435;
wire n_20436;
wire n_20437;
wire n_20438;
wire n_20439;
wire n_20440;
wire n_20441;
wire n_20442;
wire n_20443;
wire n_20444;
wire n_20445;
wire n_20446;
wire n_20447;
wire n_20448;
wire n_20449;
wire n_20450;
wire n_20451;
wire n_20452;
wire n_20453;
wire n_20454;
wire n_20455;
wire n_20456;
wire n_20457;
wire n_20458;
wire n_20459;
wire n_20460;
wire n_20461;
wire n_20462;
wire n_20463;
wire n_20464;
wire n_20465;
wire n_20466;
wire n_20467;
wire n_20468;
wire n_20469;
wire n_20470;
wire n_20471;
wire n_20472;
wire n_20473;
wire n_20474;
wire n_20475;
wire n_20476;
wire n_20477;
wire n_20478;
wire n_20479;
wire n_20480;
wire n_20481;
wire n_20482;
wire n_20483;
wire n_20484;
wire n_20485;
wire n_20486;
wire n_20487;
wire n_20488;
wire n_20489;
wire n_20490;
wire n_20491;
wire n_20492;
wire n_20493;
wire n_20494;
wire n_20495;
wire n_20496;
wire n_20497;
wire n_20498;
wire n_20499;
wire n_20500;
wire n_20501;
wire n_20502;
wire n_20503;
wire n_20504;
wire n_20505;
wire n_20506;
wire n_20507;
wire n_20508;
wire n_20509;
wire n_20510;
wire n_20511;
wire n_20512;
wire n_20513;
wire n_20514;
wire n_20515;
wire n_20516;
wire n_20517;
wire n_20518;
wire n_20519;
wire n_20520;
wire n_20521;
wire n_20522;
wire n_20523;
wire n_20524;
wire n_20525;
wire n_20526;
wire n_20527;
wire n_20528;
wire n_20529;
wire n_20530;
wire n_20531;
wire n_20532;
wire n_20533;
wire n_20534;
wire n_20535;
wire n_20536;
wire n_20537;
wire n_20538;
wire n_20539;
wire n_20540;
wire n_20541;
wire n_20542;
wire n_20543;
wire n_20544;
wire n_20545;
wire n_20546;
wire n_20547;
wire n_20548;
wire n_20549;
wire n_20550;
wire n_20551;
wire n_20552;
wire n_20553;
wire n_20554;
wire n_20555;
wire n_20556;
wire n_20557;
wire n_20558;
wire n_20559;
wire n_20560;
wire n_20561;
wire n_20562;
wire n_20563;
wire n_20564;
wire n_20565;
wire n_20566;
wire n_20567;
wire n_20568;
wire n_20569;
wire n_20570;
wire n_20571;
wire n_20572;
wire n_20573;
wire n_20574;
wire n_20575;
wire n_20576;
wire n_20577;
wire n_20578;
wire n_20579;
wire n_20580;
wire n_20581;
wire n_20582;
wire n_20583;
wire n_20584;
wire n_20585;
wire n_20586;
wire n_20587;
wire n_20588;
wire n_20589;
wire n_20590;
wire n_20591;
wire n_20592;
wire n_20593;
wire n_20594;
wire n_20595;
wire n_20596;
wire n_20597;
wire n_20598;
wire n_20599;
wire n_20600;
wire n_20601;
wire n_20602;
wire n_20603;
wire n_20604;
wire n_20605;
wire n_20606;
wire n_20607;
wire n_20608;
wire n_20609;
wire n_20610;
wire n_20611;
wire n_20612;
wire n_20613;
wire n_20614;
wire n_20615;
wire n_20616;
wire n_20617;
wire n_20618;
wire n_20619;
wire n_20620;
wire n_20621;
wire n_20622;
wire n_20623;
wire n_20624;
wire n_20625;
wire n_20626;
wire n_20627;
wire n_20628;
wire n_20629;
wire n_20630;
wire n_20631;
wire n_20632;
wire n_20633;
wire n_20634;
wire n_20635;
wire n_20636;
wire n_20637;
wire n_20638;
wire n_20639;
wire n_20640;
wire n_20641;
wire n_20642;
wire n_20643;
wire n_20644;
wire n_20645;
wire n_20646;
wire n_20647;
wire n_20648;
wire n_20649;
wire n_20650;
wire n_20651;
wire n_20652;
wire n_20653;
wire n_20654;
wire n_20655;
wire n_20656;
wire n_20657;
wire n_20658;
wire n_20659;
wire n_20660;
wire n_20661;
wire n_20662;
wire n_20663;
wire n_20664;
wire n_20665;
wire n_20666;
wire n_20667;
wire n_20668;
wire n_20669;
wire n_20670;
wire n_20671;
wire n_20672;
wire n_20673;
wire n_20674;
wire n_20675;
wire n_20676;
wire n_20677;
wire n_20678;
wire n_20679;
wire n_20680;
wire n_20681;
wire n_20682;
wire n_20683;
wire n_20684;
wire n_20685;
wire n_20686;
wire n_20687;
wire n_20688;
wire n_20689;
wire n_20690;
wire n_20691;
wire n_20692;
wire n_20693;
wire n_20694;
wire n_20695;
wire n_20696;
wire n_20697;
wire n_20698;
wire n_20699;
wire n_20700;
wire n_20701;
wire n_20702;
wire n_20703;
wire n_20704;
wire n_20705;
wire n_20706;
wire n_20707;
wire n_20708;
wire n_20709;
wire n_20710;
wire n_20711;
wire n_20712;
wire n_20713;
wire n_20714;
wire n_20715;
wire n_20716;
wire n_20717;
wire n_20718;
wire n_20719;
wire n_20720;
wire n_20721;
wire n_20722;
wire n_20723;
wire n_20724;
wire n_20725;
wire n_20726;
wire n_20727;
wire n_20728;
wire n_20729;
wire n_20730;
wire n_20731;
wire n_20732;
wire n_20733;
wire n_20734;
wire n_20735;
wire n_20736;
wire n_20737;
wire n_20738;
wire n_20739;
wire n_20740;
wire n_20741;
wire n_20742;
wire n_20743;
wire n_20744;
wire n_20745;
wire n_20746;
wire n_20747;
wire n_20748;
wire n_20749;
wire n_20750;
wire n_20751;
wire n_20752;
wire n_20753;
wire n_20754;
wire n_20755;
wire n_20756;
wire n_20757;
wire n_20758;
wire n_20759;
wire n_20760;
wire n_20761;
wire n_20762;
wire n_20763;
wire n_20764;
wire n_20765;
wire n_20766;
wire n_20767;
wire n_20768;
wire n_20769;
wire n_20770;
wire n_20771;
wire n_20772;
wire n_20773;
wire n_20774;
wire n_20775;
wire n_20776;
wire n_20777;
wire n_20778;
wire n_20779;
wire n_20780;
wire n_20781;
wire n_20782;
wire n_20783;
wire n_20784;
wire n_20785;
wire n_20786;
wire n_20787;
wire n_20788;
wire n_20789;
wire n_20790;
wire n_20791;
wire n_20792;
wire n_20793;
wire n_20794;
wire n_20795;
wire n_20796;
wire n_20797;
wire n_20798;
wire n_20799;
wire n_20800;
wire n_20801;
wire n_20802;
wire n_20803;
wire n_20804;
wire n_20805;
wire n_20806;
wire n_20807;
wire n_20808;
wire n_20809;
wire n_20810;
wire n_20811;
wire n_20812;
wire n_20813;
wire n_20814;
wire n_20815;
wire n_20816;
wire n_20817;
wire n_20818;
wire n_20819;
wire n_20820;
wire n_20821;
wire n_20822;
wire n_20823;
wire n_20824;
wire n_20825;
wire n_20826;
wire n_20827;
wire n_20828;
wire n_20829;
wire n_20830;
wire n_20831;
wire n_20832;
wire n_20833;
wire n_20834;
wire n_20835;
wire n_20836;
wire n_20837;
wire n_20838;
wire n_20839;
wire n_20840;
wire n_20841;
wire n_20842;
wire n_20843;
wire n_20844;
wire n_20845;
wire n_20846;
wire n_20847;
wire n_20848;
wire n_20849;
wire n_20850;
wire n_20851;
wire n_20852;
wire n_20853;
wire n_20854;
wire n_20855;
wire n_20856;
wire n_20857;
wire n_20858;
wire n_20859;
wire n_20860;
wire n_20861;
wire n_20862;
wire n_20863;
wire n_20864;
wire n_20865;
wire n_20866;
wire n_20867;
wire n_20868;
wire n_20869;
wire n_20870;
wire n_20871;
wire n_20872;
wire n_20873;
wire n_20874;
wire n_20875;
wire n_20876;
wire n_20877;
wire n_20878;
wire n_20879;
wire n_20880;
wire n_20881;
wire n_20882;
wire n_20883;
wire n_20884;
wire n_20885;
wire n_20886;
wire n_20887;
wire n_20888;
wire n_20889;
wire n_20890;
wire n_20891;
wire n_20892;
wire n_20893;
wire n_20894;
wire n_20895;
wire n_20896;
wire n_20897;
wire n_20898;
wire n_20899;
wire n_20900;
wire n_20901;
wire n_20902;
wire n_20903;
wire n_20904;
wire n_20905;
wire n_20906;
wire n_20907;
wire n_20908;
wire n_20909;
wire n_20910;
wire n_20911;
wire n_20912;
wire n_20913;
wire n_20914;
wire n_20915;
wire n_20916;
wire n_20917;
wire n_20918;
wire n_20919;
wire n_20920;
wire n_20921;
wire n_20922;
wire n_20923;
wire n_20924;
wire n_20925;
wire n_20926;
wire n_20927;
wire n_20928;
wire n_20929;
wire n_20930;
wire n_20931;
wire n_20932;
wire n_20933;
wire n_20934;
wire n_20935;
wire n_20936;
wire n_20937;
wire n_20938;
wire n_20939;
wire n_20940;
wire n_20941;
wire n_20942;
wire n_20943;
wire n_20944;
wire n_20945;
wire n_20946;
wire n_20947;
wire n_20948;
wire n_20949;
wire n_20950;
wire n_20951;
wire n_20952;
wire n_20953;
wire n_20954;
wire n_20955;
wire n_20956;
wire n_20957;
wire n_20958;
wire n_20959;
wire n_20960;
wire n_20961;
wire n_20962;
wire n_20963;
wire n_20964;
wire n_20965;
wire n_20966;
wire n_20967;
wire n_20968;
wire n_20969;
wire n_20970;
wire n_20971;
wire n_20972;
wire n_20973;
wire n_20974;
wire n_20975;
wire n_20976;
wire n_20977;
wire n_20978;
wire n_20979;
wire n_20980;
wire n_20981;
wire n_20982;
wire n_20983;
wire n_20984;
wire n_20985;
wire n_20986;
wire n_20987;
wire n_20988;
wire n_20989;
wire n_20990;
wire n_20991;
wire n_20992;
wire n_20993;
wire n_20994;
wire n_20995;
wire n_20996;
wire n_20997;
wire n_20998;
wire n_20999;
wire n_21000;
wire n_21001;
wire n_21002;
wire n_21003;
wire n_21004;
wire n_21005;
wire n_21006;
wire n_21007;
wire n_21008;
wire n_21009;
wire n_21010;
wire n_21011;
wire n_21012;
wire n_21013;
wire n_21014;
wire n_21015;
wire n_21016;
wire n_21017;
wire n_21018;
wire n_21019;
wire n_21020;
wire n_21021;
wire n_21022;
wire n_21023;
wire n_21024;
wire n_21025;
wire n_21026;
wire n_21027;
wire n_21028;
wire n_21029;
wire n_21030;
wire n_21031;
wire n_21032;
wire n_21033;
wire n_21034;
wire n_21035;
wire n_21036;
wire n_21037;
wire n_21038;
wire n_21039;
wire n_21040;
wire n_21041;
wire n_21042;
wire n_21043;
wire n_21044;
wire n_21045;
wire n_21046;
wire n_21047;
wire n_21048;
wire n_21049;
wire n_21050;
wire n_21051;
wire n_21052;
wire n_21053;
wire n_21054;
wire n_21055;
wire n_21056;
wire n_21057;
wire n_21058;
wire n_21059;
wire n_21060;
wire n_21061;
wire n_21062;
wire n_21063;
wire n_21064;
wire n_21065;
wire n_21066;
wire n_21067;
wire n_21068;
wire n_21069;
wire n_21070;
wire n_21071;
wire n_21072;
wire n_21073;
wire n_21074;
wire n_21075;
wire n_21076;
wire n_21077;
wire n_21078;
wire n_21079;
wire n_21080;
wire n_21081;
wire n_21082;
wire n_21083;
wire n_21084;
wire n_21085;
wire n_21086;
wire n_21087;
wire n_21088;
wire n_21089;
wire n_21090;
wire n_21091;
wire n_21092;
wire n_21093;
wire n_21094;
wire n_21095;
wire n_21096;
wire n_21097;
wire n_21098;
wire n_21099;
wire n_21100;
wire n_21101;
wire n_21102;
wire n_21103;
wire n_21104;
wire n_21105;
wire n_21106;
wire n_21107;
wire n_21108;
wire n_21109;
wire n_21110;
wire n_21111;
wire n_21112;
wire n_21113;
wire n_21114;
wire n_21115;
wire n_21116;
wire n_21117;
wire n_21118;
wire n_21119;
wire n_21120;
wire n_21121;
wire n_21122;
wire n_21123;
wire n_21124;
wire n_21125;
wire n_21126;
wire n_21127;
wire n_21128;
wire n_21129;
wire n_21130;
wire n_21131;
wire n_21132;
wire n_21133;
wire n_21134;
wire n_21135;
wire n_21136;
wire n_21137;
wire n_21138;
wire n_21139;
wire n_21140;
wire n_21141;
wire n_21142;
wire n_21143;
wire n_21144;
wire n_21145;
wire n_21146;
wire n_21147;
wire n_21148;
wire n_21149;
wire n_21150;
wire n_21151;
wire n_21152;
wire n_21153;
wire n_21154;
wire n_21155;
wire n_21156;
wire n_21157;
wire n_21158;
wire n_21159;
wire n_21160;
wire n_21161;
wire n_21162;
wire n_21163;
wire n_21164;
wire n_21165;
wire n_21166;
wire n_21167;
wire n_21168;
wire n_21169;
wire n_21170;
wire n_21171;
wire n_21172;
wire n_21173;
wire n_21174;
wire n_21175;
wire n_21176;
wire n_21177;
wire n_21178;
wire n_21179;
wire n_21180;
wire n_21181;
wire n_21182;
wire n_21183;
wire n_21184;
wire n_21185;
wire n_21186;
wire n_21187;
wire n_21188;
wire n_21189;
wire n_21190;
wire n_21191;
wire n_21192;
wire n_21193;
wire n_21194;
wire n_21195;
wire n_21196;
wire n_21197;
wire n_21198;
wire n_21199;
wire n_21200;
wire n_21201;
wire n_21202;
wire n_21203;
wire n_21204;
wire n_21205;
wire n_21206;
wire n_21207;
wire n_21208;
wire n_21209;
wire n_21210;
wire n_21211;
wire n_21212;
wire n_21213;
wire n_21214;
wire n_21215;
wire n_21216;
wire n_21217;
wire n_21218;
wire n_21219;
wire n_21220;
wire n_21221;
wire n_21222;
wire n_21223;
wire n_21224;
wire n_21225;
wire n_21226;
wire n_21227;
wire n_21228;
wire n_21229;
wire n_21230;
wire n_21231;
wire n_21232;
wire n_21233;
wire n_21234;
wire n_21235;
wire n_21236;
wire n_21237;
wire n_21238;
wire n_21239;
wire n_21240;
wire n_21241;
wire n_21242;
wire n_21243;
wire n_21244;
wire n_21245;
wire n_21246;
wire n_21247;
wire n_21248;
wire n_21249;
wire n_21250;
wire n_21251;
wire n_21252;
wire n_21253;
wire n_21254;
wire n_21255;
wire n_21256;
wire n_21257;
wire n_21258;
wire n_21259;
wire n_21260;
wire n_21261;
wire n_21262;
wire n_21263;
wire n_21264;
wire n_21265;
wire n_21266;
wire n_21267;
wire n_21268;
wire n_21269;
wire n_21270;
wire n_21271;
wire n_21272;
wire n_21273;
wire n_21274;
wire n_21275;
wire n_21276;
wire n_21277;
wire n_21278;
wire n_21279;
wire n_21280;
wire n_21281;
wire n_21282;
wire n_21283;
wire n_21284;
wire n_21285;
wire n_21286;
wire n_21287;
wire n_21288;
wire n_21289;
wire n_21290;
wire n_21291;
wire n_21292;
wire n_21293;
wire n_21294;
wire n_21295;
wire n_21296;
wire n_21297;
wire n_21298;
wire n_21299;
wire n_21300;
wire n_21301;
wire n_21302;
wire n_21303;
wire n_21304;
wire n_21305;
wire n_21306;
wire n_21307;
wire n_21308;
wire n_21309;
wire n_21310;
wire n_21311;
wire n_21312;
wire n_21313;
wire n_21314;
wire n_21315;
wire n_21316;
wire n_21317;
wire n_21318;
wire n_21319;
wire n_21320;
wire n_21321;
wire n_21322;
wire n_21323;
wire n_21324;
wire n_21325;
wire n_21326;
wire n_21327;
wire n_21328;
wire n_21329;
wire n_21330;
wire n_21331;
wire n_21332;
wire n_21333;
wire n_21334;
wire n_21335;
wire n_21336;
wire n_21337;
wire n_21338;
wire n_21339;
wire n_21340;
wire n_21341;
wire n_21342;
wire n_21343;
wire n_21344;
wire n_21345;
wire n_21346;
wire n_21347;
wire n_21348;
wire n_21349;
wire n_21350;
wire n_21351;
wire n_21352;
wire n_21353;
wire n_21354;
wire n_21355;
wire n_21356;
wire n_21357;
wire n_21358;
wire n_21359;
wire n_21360;
wire n_21361;
wire n_21362;
wire n_21363;
wire n_21364;
wire n_21365;
wire n_21366;
wire n_21367;
wire n_21368;
wire n_21369;
wire n_21370;
wire n_21371;
wire n_21372;
wire n_21373;
wire n_21374;
wire n_21375;
wire n_21376;
wire n_21377;
wire n_21378;
wire n_21379;
wire n_21380;
wire n_21381;
wire n_21382;
wire n_21383;
wire n_21384;
wire n_21385;
wire n_21386;
wire n_21387;
wire n_21388;
wire n_21389;
wire n_21390;
wire n_21391;
wire n_21392;
wire n_21393;
wire n_21394;
wire n_21395;
wire n_21396;
wire n_21397;
wire n_21398;
wire n_21399;
wire n_21400;
wire n_21401;
wire n_21402;
wire n_21403;
wire n_21404;
wire n_21405;
wire n_21406;
wire n_21407;
wire n_21408;
wire n_21409;
wire n_21410;
wire n_21411;
wire n_21412;
wire n_21413;
wire n_21414;
wire n_21415;
wire n_21416;
wire n_21417;
wire n_21418;
wire n_21419;
wire n_21420;
wire n_21421;
wire n_21422;
wire n_21423;
wire n_21424;
wire n_21425;
wire n_21426;
wire n_21427;
wire n_21428;
wire n_21429;
wire n_21430;
wire n_21431;
wire n_21432;
wire n_21433;
wire n_21434;
wire n_21435;
wire n_21436;
wire n_21437;
wire n_21438;
wire n_21439;
wire n_21440;
wire n_21441;
wire n_21442;
wire n_21443;
wire n_21444;
wire n_21445;
wire n_21446;
wire n_21447;
wire n_21448;
wire n_21449;
wire n_21450;
wire n_21451;
wire n_21452;
wire n_21453;
wire n_21454;
wire n_21455;
wire n_21456;
wire n_21457;
wire n_21458;
wire n_21459;
wire n_21460;
wire n_21461;
wire n_21462;
wire n_21463;
wire n_21464;
wire n_21465;
wire n_21466;
wire n_21467;
wire n_21468;
wire n_21469;
wire n_21470;
wire n_21471;
wire n_21472;
wire n_21473;
wire n_21474;
wire n_21475;
wire n_21476;
wire n_21477;
wire n_21478;
wire n_21479;
wire n_21480;
wire n_21481;
wire n_21482;
wire n_21483;
wire n_21484;
wire n_21485;
wire n_21486;
wire n_21487;
wire n_21488;
wire n_21489;
wire n_21490;
wire n_21491;
wire n_21492;
wire n_21493;
wire n_21494;
wire n_21495;
wire n_21496;
wire n_21497;
wire n_21498;
wire n_21499;
wire n_21500;
wire n_21501;
wire n_21502;
wire n_21503;
wire n_21504;
wire n_21505;
wire n_21506;
wire n_21507;
wire n_21508;
wire n_21509;
wire n_21510;
wire n_21511;
wire n_21512;
wire n_21513;
wire n_21514;
wire n_21515;
wire n_21516;
wire n_21517;
wire n_21518;
wire n_21519;
wire n_21520;
wire n_21521;
wire n_21522;
wire n_21523;
wire n_21524;
wire n_21525;
wire n_21526;
wire n_21527;
wire n_21528;
wire n_21529;
wire n_21530;
wire n_21531;
wire n_21532;
wire n_21533;
wire n_21534;
wire n_21535;
wire n_21536;
wire n_21537;
wire n_21538;
wire n_21539;
wire n_21540;
wire n_21541;
wire n_21542;
wire n_21543;
wire n_21544;
wire n_21545;
wire n_21546;
wire n_21547;
wire n_21548;
wire n_21549;
wire n_21550;
wire n_21551;
wire n_21552;
wire n_21553;
wire n_21554;
wire n_21555;
wire n_21556;
wire n_21557;
wire n_21558;
wire n_21559;
wire n_21560;
wire n_21561;
wire n_21562;
wire n_21563;
wire n_21564;
wire n_21565;
wire n_21566;
wire n_21567;
wire n_21568;
wire n_21569;
wire n_21570;
wire n_21571;
wire n_21572;
wire n_21573;
wire n_21574;
wire n_21575;
wire n_21576;
wire n_21577;
wire n_21578;
wire n_21579;
wire n_21580;
wire n_21581;
wire n_21582;
wire n_21583;
wire n_21584;
wire n_21585;
wire n_21586;
wire n_21587;
wire n_21588;
wire n_21589;
wire n_21590;
wire n_21591;
wire n_21592;
wire n_21593;
wire n_21594;
wire n_21595;
wire n_21596;
wire n_21597;
wire n_21598;
wire n_21599;
wire n_21600;
wire n_21601;
wire n_21602;
wire n_21603;
wire n_21604;
wire n_21605;
wire n_21606;
wire n_21607;
wire n_21608;
wire n_21609;
wire n_21610;
wire n_21611;
wire n_21612;
wire n_21613;
wire n_21614;
wire n_21615;
wire n_21616;
wire n_21617;
wire n_21618;
wire n_21619;
wire n_21620;
wire n_21621;
wire n_21622;
wire n_21623;
wire n_21624;
wire n_21625;
wire n_21626;
wire n_21627;
wire n_21628;
wire n_21629;
wire n_21630;
wire n_21631;
wire n_21632;
wire n_21633;
wire n_21634;
wire n_21635;
wire n_21636;
wire n_21637;
wire n_21638;
wire n_21639;
wire n_21640;
wire n_21641;
wire n_21642;
wire n_21643;
wire n_21644;
wire n_21645;
wire n_21646;
wire n_21647;
wire n_21648;
wire n_21649;
wire n_21650;
wire n_21651;
wire n_21652;
wire n_21653;
wire n_21654;
wire n_21655;
wire n_21656;
wire n_21657;
wire n_21658;
wire n_21659;
wire n_21660;
wire n_21661;
wire n_21662;
wire n_21663;
wire n_21664;
wire n_21665;
wire n_21666;
wire n_21667;
wire n_21668;
wire n_21669;
wire n_21670;
wire n_21671;
wire n_21672;
wire n_21673;
wire n_21674;
wire n_21675;
wire n_21676;
wire n_21677;
wire n_21678;
wire n_21679;
wire n_21680;
wire n_21681;
wire n_21682;
wire n_21683;
wire n_21684;
wire n_21685;
wire n_21686;
wire n_21687;
wire n_21688;
wire n_21689;
wire n_21690;
wire n_21691;
wire n_21692;
wire n_21693;
wire n_21694;
wire n_21695;
wire n_21696;
wire n_21697;
wire n_21698;
wire n_21699;
wire n_21700;
wire n_21701;
wire n_21702;
wire n_21703;
wire n_21704;
wire n_21705;
wire n_21706;
wire n_21707;
wire n_21708;
wire n_21709;
wire n_21710;
wire n_21711;
wire n_21712;
wire n_21713;
wire n_21714;
wire n_21715;
wire n_21716;
wire n_21717;
wire n_21718;
wire n_21719;
wire n_21720;
wire n_21721;
wire n_21722;
wire n_21723;
wire n_21724;
wire n_21725;
wire n_21726;
wire n_21727;
wire n_21728;
wire n_21729;
wire n_21730;
wire n_21731;
wire n_21732;
wire n_21733;
wire n_21734;
wire n_21735;
wire n_21736;
wire n_21737;
wire n_21738;
wire n_21739;
wire n_21740;
wire n_21741;
wire n_21742;
wire n_21743;
wire n_21744;
wire n_21745;
wire n_21746;
wire n_21747;
wire n_21748;
wire n_21749;
wire n_21750;
wire n_21751;
wire n_21752;
wire n_21753;
wire n_21754;
wire n_21755;
wire n_21756;
wire n_21757;
wire n_21758;
wire n_21759;
wire n_21760;
wire n_21761;
wire n_21762;
wire n_21763;
wire n_21764;
wire n_21765;
wire n_21766;
wire n_21767;
wire n_21768;
wire n_21769;
wire n_21770;
wire n_21771;
wire n_21772;
wire n_21773;
wire n_21774;
wire n_21775;
wire n_21776;
wire n_21777;
wire n_21778;
wire n_21779;
wire n_21780;
wire n_21781;
wire n_21782;
wire n_21783;
wire n_21784;
wire n_21785;
wire n_21786;
wire n_21787;
wire n_21788;
wire n_21789;
wire n_21790;
wire n_21791;
wire n_21792;
wire n_21793;
wire n_21794;
wire n_21795;
wire n_21796;
wire n_21797;
wire n_21798;
wire n_21799;
wire n_21800;
wire n_21801;
wire n_21802;
wire n_21803;
wire n_21804;
wire n_21805;
wire n_21806;
wire n_21807;
wire n_21808;
wire n_21809;
wire n_21810;
wire n_21811;
wire n_21812;
wire n_21813;
wire n_21814;
wire n_21815;
wire n_21816;
wire n_21817;
wire n_21818;
wire n_21819;
wire n_21820;
wire n_21821;
wire n_21822;
wire n_21823;
wire n_21824;
wire n_21825;
wire n_21826;
wire n_21827;
wire n_21828;
wire n_21829;
wire n_21830;
wire n_21831;
wire n_21832;
wire n_21833;
wire n_21834;
wire n_21835;
wire n_21836;
wire n_21837;
wire n_21838;
wire n_21839;
wire n_21840;
wire n_21841;
wire n_21842;
wire n_21843;
wire n_21844;
wire n_21845;
wire n_21846;
wire n_21847;
wire n_21848;
wire n_21849;
wire n_21850;
wire n_21851;
wire n_21852;
wire n_21853;
wire n_21854;
wire n_21855;
wire n_21856;
wire n_21857;
wire n_21858;
wire n_21859;
wire n_21860;
wire n_21861;
wire n_21862;
wire n_21863;
wire n_21864;
wire n_21865;
wire n_21866;
wire n_21867;
wire n_21868;
wire n_21869;
wire n_21870;
wire n_21871;
wire n_21872;
wire n_21873;
wire n_21874;
wire n_21875;
wire n_21876;
wire n_21877;
wire n_21878;
wire n_21879;
wire n_21880;
wire n_21881;
wire n_21882;
wire n_21883;
wire n_21884;
wire n_21885;
wire n_21886;
wire n_21887;
wire n_21888;
wire n_21889;
wire n_21890;
wire n_21891;
wire n_21892;
wire n_21893;
wire n_21894;
wire n_21895;
wire n_21896;
wire n_21897;
wire n_21898;
wire n_21899;
wire n_21900;
wire n_21901;
wire n_21902;
wire n_21903;
wire n_21904;
wire n_21905;
wire n_21906;
wire n_21907;
wire n_21908;
wire n_21909;
wire n_21910;
wire n_21911;
wire n_21912;
wire n_21913;
wire n_21914;
wire n_21915;
wire n_21916;
wire n_21917;
wire n_21918;
wire n_21919;
wire n_21920;
wire n_21921;
wire n_21922;
wire n_21923;
wire n_21924;
wire n_21925;
wire n_21926;
wire n_21927;
wire n_21928;
wire n_21929;
wire n_21930;
wire n_21931;
wire n_21932;
wire n_21933;
wire n_21934;
wire n_21935;
wire n_21936;
wire n_21937;
wire n_21938;
wire n_21939;
wire n_21940;
wire n_21941;
wire n_21942;
wire n_21943;
wire n_21944;
wire n_21945;
wire n_21946;
wire n_21947;
wire n_21948;
wire n_21949;
wire n_21950;
wire n_21951;
wire n_21952;
wire n_21953;
wire n_21954;
wire n_21955;
wire n_21956;
wire n_21957;
wire n_21958;
wire n_21959;
wire n_21960;
wire n_21961;
wire n_21962;
wire n_21963;
wire n_21964;
wire n_21965;
wire n_21966;
wire n_21967;
wire n_21968;
wire n_21969;
wire n_21970;
wire n_21971;
wire n_21972;
wire n_21973;
wire n_21974;
wire n_21975;
wire n_21976;
wire n_21977;
wire n_21978;
wire n_21979;
wire n_21980;
wire n_21981;
wire n_21982;
wire n_21983;
wire n_21984;
wire n_21985;
wire n_21986;
wire n_21987;
wire n_21988;
wire n_21989;
wire n_21990;
wire n_21991;
wire n_21992;
wire n_21993;
wire n_21994;
wire n_21995;
wire n_21996;
wire n_21997;
wire n_21998;
wire n_21999;
wire n_22000;
wire n_22001;
wire n_22002;
wire n_22003;
wire n_22004;
wire n_22005;
wire n_22006;
wire n_22007;
wire n_22008;
wire n_22009;
wire n_22010;
wire n_22011;
wire n_22012;
wire n_22013;
wire n_22014;
wire n_22015;
wire n_22016;
wire n_22017;
wire n_22018;
wire n_22019;
wire n_22020;
wire n_22021;
wire n_22022;
wire n_22023;
wire n_22024;
wire n_22025;
wire n_22026;
wire n_22027;
wire n_22028;
wire n_22029;
wire n_22030;
wire n_22031;
wire n_22032;
wire n_22033;
wire n_22034;
wire n_22035;
wire n_22036;
wire n_22037;
wire n_22038;
wire n_22039;
wire n_22040;
wire n_22041;
wire n_22042;
wire n_22043;
wire n_22044;
wire n_22045;
wire n_22046;
wire n_22047;
wire n_22048;
wire n_22049;
wire n_22050;
wire n_22051;
wire n_22052;
wire n_22053;
wire n_22054;
wire n_22055;
wire n_22056;
wire n_22057;
wire n_22058;
wire n_22059;
wire n_22060;
wire n_22061;
wire n_22062;
wire n_22063;
wire n_22064;
wire n_22065;
wire n_22066;
wire n_22067;
wire n_22068;
wire n_22069;
wire n_22070;
wire n_22071;
wire n_22072;
wire n_22073;
wire n_22074;
wire n_22075;
wire n_22076;
wire n_22077;
wire n_22078;
wire n_22079;
wire n_22080;
wire n_22081;
wire n_22082;
wire n_22083;
wire n_22084;
wire n_22085;
wire n_22086;
wire n_22087;
wire n_22088;
wire n_22089;
wire n_22090;
wire n_22091;
wire n_22092;
wire n_22093;
wire n_22094;
wire n_22095;
wire n_22096;
wire n_22097;
wire n_22098;
wire n_22099;
wire n_22100;
wire n_22101;
wire n_22102;
wire n_22103;
wire n_22104;
wire n_22105;
wire n_22106;
wire n_22107;
wire n_22108;
wire n_22109;
wire n_22110;
wire n_22111;
wire n_22112;
wire n_22113;
wire n_22114;
wire n_22115;
wire n_22116;
wire n_22117;
wire n_22118;
wire n_22119;
wire n_22120;
wire n_22121;
wire n_22122;
wire n_22123;
wire n_22124;
wire n_22125;
wire n_22126;
wire n_22127;
wire n_22128;
wire n_22129;
wire n_22130;
wire n_22131;
wire n_22132;
wire n_22133;
wire n_22134;
wire n_22135;
wire n_22136;
wire n_22137;
wire n_22138;
wire n_22139;
wire n_22140;
wire n_22141;
wire n_22142;
wire n_22143;
wire n_22144;
wire n_22145;
wire n_22146;
wire n_22147;
wire n_22148;
wire n_22149;
wire n_22150;
wire n_22151;
wire n_22152;
wire n_22153;
wire n_22154;
wire n_22155;
wire n_22156;
wire n_22157;
wire n_22158;
wire n_22159;
wire n_22160;
wire n_22161;
wire n_22162;
wire n_22163;
wire n_22164;
wire n_22165;
wire n_22166;
wire n_22167;
wire n_22168;
wire n_22169;
wire n_22170;
wire n_22171;
wire n_22172;
wire n_22173;
wire n_22174;
wire n_22175;
wire n_22176;
wire n_22177;
wire n_22178;
wire n_22179;
wire n_22180;
wire n_22181;
wire n_22182;
wire n_22183;
wire n_22184;
wire n_22185;
wire n_22186;
wire n_22187;
wire n_22188;
wire n_22189;
wire n_22190;
wire n_22191;
wire n_22192;
wire n_22193;
wire n_22194;
wire n_22195;
wire n_22196;
wire n_22197;
wire n_22198;
wire n_22199;
wire n_22200;
wire n_22201;
wire n_22202;
wire n_22203;
wire n_22204;
wire n_22205;
wire n_22206;
wire n_22207;
wire n_22208;
wire n_22209;
wire n_22210;
wire n_22211;
wire n_22212;
wire n_22213;
wire n_22214;
wire n_22215;
wire n_22216;
wire n_22217;
wire n_22218;
wire n_22219;
wire n_22220;
wire n_22221;
wire n_22222;
wire n_22223;
wire n_22224;
wire n_22225;
wire n_22226;
wire n_22227;
wire n_22228;
wire n_22229;
wire n_22230;
wire n_22231;
wire n_22232;
wire n_22233;
wire n_22234;
wire n_22235;
wire n_22236;
wire n_22237;
wire n_22238;
wire n_22239;
wire n_22240;
wire n_22241;
wire n_22242;
wire n_22243;
wire n_22244;
wire n_22245;
wire n_22246;
wire n_22247;
wire n_22248;
wire n_22249;
wire n_22250;
wire n_22251;
wire n_22252;
wire n_22253;
wire n_22254;
wire n_22255;
wire n_22256;
wire n_22257;
wire n_22258;
wire n_22259;
wire n_22260;
wire n_22261;
wire n_22262;
wire n_22263;
wire n_22264;
wire n_22265;
wire n_22266;
wire n_22267;
wire n_22268;
wire n_22269;
wire n_22270;
wire n_22271;
wire n_22272;
wire n_22273;
wire n_22274;
wire n_22275;
wire n_22276;
wire n_22277;
wire n_22278;
wire n_22279;
wire n_22280;
wire n_22281;
wire n_22282;
wire n_22283;
wire n_22284;
wire n_22285;
wire n_22286;
wire n_22287;
wire n_22288;
wire n_22289;
wire n_22290;
wire n_22291;
wire n_22292;
wire n_22293;
wire n_22294;
wire n_22295;
wire n_22296;
wire n_22297;
wire n_22298;
wire n_22299;
wire n_22300;
wire n_22301;
wire n_22302;
wire n_22303;
wire n_22304;
wire n_22305;
wire n_22306;
wire n_22307;
wire n_22308;
wire n_22309;
wire n_22310;
wire n_22311;
wire n_22312;
wire n_22313;
wire n_22314;
wire n_22315;
wire n_22316;
wire n_22317;
wire n_22318;
wire n_22319;
wire n_22320;
wire n_22321;
wire n_22322;
wire n_22323;
wire n_22324;
wire n_22325;
wire n_22326;
wire n_22327;
wire n_22328;
wire n_22329;
wire n_22330;
wire n_22331;
wire n_22332;
wire n_22333;
wire n_22334;
wire n_22335;
wire n_22336;
wire n_22337;
wire n_22338;
wire n_22339;
wire n_22340;
wire n_22341;
wire n_22342;
wire n_22343;
wire n_22344;
wire n_22345;
wire n_22346;
wire n_22347;
wire n_22348;
wire n_22349;
wire n_22350;
wire n_22351;
wire n_22352;
wire n_22353;
wire n_22354;
wire n_22355;
wire n_22356;
wire n_22357;
wire n_22358;
wire n_22359;
wire n_22360;
wire n_22361;
wire n_22362;
wire n_22363;
wire n_22364;
wire n_22365;
wire n_22366;
wire n_22367;
wire n_22368;
wire n_22369;
wire n_22370;
wire n_22371;
wire n_22372;
wire n_22373;
wire n_22374;
wire n_22375;
wire n_22376;
wire n_22377;
wire n_22378;
wire n_22379;
wire n_22380;
wire n_22381;
wire n_22382;
wire n_22383;
wire n_22384;
wire n_22385;
wire n_22386;
wire n_22387;
wire n_22388;
wire n_22389;
wire n_22390;
wire n_22391;
wire n_22392;
wire n_22393;
wire n_22394;
wire n_22395;
wire n_22396;
wire n_22397;
wire n_22398;
wire n_22399;
wire n_22400;
wire n_22401;
wire n_22402;
wire n_22403;
wire n_22404;
wire n_22405;
wire n_22406;
wire n_22407;
wire n_22408;
wire n_22409;
wire n_22410;
wire n_22411;
wire n_22412;
wire n_22413;
wire n_22414;
wire n_22415;
wire n_22416;
wire n_22417;
wire n_22418;
wire n_22419;
wire n_22420;
wire n_22421;
wire n_22422;
wire n_22423;
wire n_22424;
wire n_22425;
wire n_22426;
wire n_22427;
wire n_22428;
wire n_22429;
wire n_22430;
wire n_22431;
wire n_22432;
wire n_22433;
wire n_22434;
wire n_22435;
wire n_22436;
wire n_22437;
wire n_22438;
wire n_22439;
wire n_22440;
wire n_22441;
wire n_22442;
wire n_22443;
wire n_22444;
wire n_22445;
wire n_22446;
wire n_22447;
wire n_22448;
wire n_22449;
wire n_22450;
wire n_22451;
wire n_22452;
wire n_22453;
wire n_22454;
wire n_22455;
wire n_22456;
wire n_22457;
wire n_22458;
wire n_22459;
wire n_22460;
wire n_22461;
wire n_22462;
wire n_22463;
wire n_22464;
wire n_22465;
wire n_22466;
wire n_22467;
wire n_22468;
wire n_22469;
wire n_22470;
wire n_22471;
wire n_22472;
wire n_22473;
wire n_22474;
wire n_22475;
wire n_22476;
wire n_22477;
wire n_22478;
wire n_22479;
wire n_22480;
wire n_22481;
wire n_22482;
wire n_22483;
wire n_22484;
wire n_22485;
wire n_22486;
wire n_22487;
wire n_22488;
wire n_22489;
wire n_22490;
wire n_22491;
wire n_22492;
wire n_22493;
wire n_22494;
wire n_22495;
wire n_22496;
wire n_22497;
wire n_22498;
wire n_22499;
wire n_22500;
wire n_22501;
wire n_22502;
wire n_22503;
wire n_22504;
wire n_22505;
wire n_22506;
wire n_22507;
wire n_22508;
wire n_22509;
wire n_22510;
wire n_22511;
wire n_22512;
wire n_22513;
wire n_22514;
wire n_22515;
wire n_22516;
wire n_22517;
wire n_22518;
wire n_22519;
wire n_22520;
wire n_22521;
wire n_22522;
wire n_22523;
wire n_22524;
wire n_22525;
wire n_22526;
wire n_22527;
wire n_22528;
wire n_22529;
wire n_22530;
wire n_22531;
wire n_22532;
wire n_22533;
wire n_22534;
wire n_22535;
wire n_22536;
wire n_22537;
wire n_22538;
wire n_22539;
wire n_22540;
wire n_22541;
wire n_22542;
wire n_22543;
wire n_22544;
wire n_22545;
wire n_22546;
wire n_22547;
wire n_22548;
wire n_22549;
wire n_22550;
wire n_22551;
wire n_22552;
wire n_22553;
wire n_22554;
wire n_22555;
wire n_22556;
wire n_22557;
wire n_22558;
wire n_22559;
wire n_22560;
wire n_22561;
wire n_22562;
wire n_22563;
wire n_22564;
wire n_22565;
wire n_22566;
wire n_22567;
wire n_22568;
wire n_22569;
wire n_22570;
wire n_22571;
wire n_22572;
wire n_22573;
wire n_22574;
wire n_22575;
wire n_22576;
wire n_22577;
wire n_22578;
wire n_22579;
wire n_22580;
wire n_22581;
wire n_22582;
wire n_22583;
wire n_22584;
wire n_22585;
wire n_22586;
wire n_22587;
wire n_22588;
wire n_22589;
wire n_22590;
wire n_22591;
wire n_22592;
wire n_22593;
wire n_22594;
wire n_22595;
wire n_22596;
wire n_22597;
wire n_22598;
wire n_22599;
wire n_22600;
wire n_22601;
wire n_22602;
wire n_22603;
wire n_22604;
wire n_22605;
wire n_22606;
wire n_22607;
wire n_22608;
wire n_22609;
wire n_22610;
wire n_22611;
wire n_22612;
wire n_22613;
wire n_22614;
wire n_22615;
wire n_22616;
wire n_22617;
wire n_22618;
wire n_22619;
wire n_22620;
wire n_22621;
wire n_22622;
wire n_22623;
wire n_22624;
wire n_22625;
wire n_22626;
wire n_22627;
wire n_22628;
wire n_22629;
wire n_22630;
wire n_22631;
wire n_22632;
wire n_22633;
wire n_22634;
wire n_22635;
wire n_22636;
wire n_22637;
wire n_22638;
wire n_22639;
wire n_22640;
wire n_22641;
wire n_22642;
wire n_22643;
wire n_22644;
wire n_22645;
wire n_22646;
wire n_22647;
wire n_22648;
wire n_22649;
wire n_22650;
wire n_22651;
wire n_22652;
wire n_22653;
wire n_22654;
wire n_22655;
wire n_22656;
wire n_22657;
wire n_22658;
wire n_22659;
wire n_22660;
wire n_22661;
wire n_22662;
wire n_22663;
wire n_22664;
wire n_22665;
wire n_22666;
wire n_22667;
wire n_22668;
wire n_22669;
wire n_22670;
wire n_22671;
wire n_22672;
wire n_22673;
wire n_22674;
wire n_22675;
wire n_22676;
wire n_22677;
wire n_22678;
wire n_22679;
wire n_22680;
wire n_22681;
wire n_22682;
wire n_22683;
wire n_22684;
wire n_22685;
wire n_22686;
wire n_22687;
wire n_22688;
wire n_22689;
wire n_22690;
wire n_22691;
wire n_22692;
wire n_22693;
wire n_22694;
wire n_22695;
wire n_22696;
wire n_22697;
wire n_22698;
wire n_22699;
wire n_22700;
wire n_22701;
wire n_22702;
wire n_22703;
wire n_22704;
wire n_22705;
wire n_22706;
wire n_22707;
wire n_22708;
wire n_22709;
wire n_22710;
wire n_22711;
wire n_22712;
wire n_22713;
wire n_22714;
wire n_22715;
wire n_22716;
wire n_22717;
wire n_22718;
wire n_22719;
wire n_22720;
wire n_22721;
wire n_22722;
wire n_22723;
wire n_22724;
wire n_22725;
wire n_22726;
wire n_22727;
wire n_22728;
wire n_22729;
wire n_22730;
wire n_22731;
wire n_22732;
wire n_22733;
wire n_22734;
wire n_22735;
wire n_22736;
wire n_22737;
wire n_22738;
wire n_22739;
wire n_22740;
wire n_22741;
wire n_22742;
wire n_22743;
wire n_22744;
wire n_22745;
wire n_22746;
wire n_22747;
wire n_22748;
wire n_22749;
wire n_22750;
wire n_22751;
wire n_22752;
wire n_22753;
wire n_22754;
wire n_22755;
wire n_22756;
wire n_22757;
wire n_22758;
wire n_22759;
wire n_22760;
wire n_22761;
wire n_22762;
wire n_22763;
wire n_22764;
wire n_22765;
wire n_22766;
wire n_22767;
wire n_22768;
wire n_22769;
wire n_22770;
wire n_22771;
wire n_22772;
wire n_22773;
wire n_22774;
wire n_22775;
wire n_22776;
wire n_22777;
wire n_22778;
wire n_22779;
wire n_22780;
wire n_22781;
wire n_22782;
wire n_22783;
wire n_22784;
wire n_22785;
wire n_22786;
wire n_22787;
wire n_22788;
wire n_22789;
wire n_22790;
wire n_22791;
wire n_22792;
wire n_22793;
wire n_22794;
wire n_22795;
wire n_22796;
wire n_22797;
wire n_22798;
wire n_22799;
wire n_22800;
wire n_22801;
wire n_22802;
wire n_22803;
wire n_22804;
wire n_22805;
wire n_22806;
wire n_22807;
wire n_22808;
wire n_22809;
wire n_22810;
wire n_22811;
wire n_22812;
wire n_22813;
wire n_22814;
wire n_22815;
wire n_22816;
wire n_22817;
wire n_22818;
wire n_22819;
wire n_22820;
wire n_22821;
wire n_22822;
wire n_22823;
wire n_22824;
wire n_22825;
wire n_22826;
wire n_22827;
wire n_22828;
wire n_22829;
wire n_22830;
wire n_22831;
wire n_22832;
wire n_22833;
wire n_22834;
wire n_22835;
wire n_22836;
wire n_22837;
wire n_22838;
wire n_22839;
wire n_22840;
wire n_22841;
wire n_22842;
wire n_22843;
wire n_22844;
wire n_22845;
wire n_22846;
wire n_22847;
wire n_22848;
wire n_22849;
wire n_22850;
wire n_22851;
wire n_22852;
wire n_22853;
wire n_22854;
wire n_22855;
wire n_22856;
wire n_22857;
wire n_22858;
wire n_22859;
wire n_22860;
wire n_22861;
wire n_22862;
wire n_22863;
wire n_22864;
wire n_22865;
wire n_22866;
wire n_22867;
wire n_22868;
wire n_22869;
wire n_22870;
wire n_22871;
wire n_22872;
wire n_22873;
wire n_22874;
wire n_22875;
wire n_22876;
wire n_22877;
wire n_22878;
wire n_22879;
wire n_22880;
wire n_22881;
wire n_22882;
wire n_22883;
wire n_22884;
wire n_22885;
wire n_22886;
wire n_22887;
wire n_22888;
wire n_22889;
wire n_22890;
wire n_22891;
wire n_22892;
wire n_22893;
wire n_22894;
wire n_22895;
wire n_22896;
wire n_22897;
wire n_22898;
wire n_22899;
wire n_22900;
wire n_22901;
wire n_22902;
wire n_22903;
wire n_22904;
wire n_22905;
wire n_22906;
wire n_22907;
wire n_22908;
wire n_22909;
wire n_22910;
wire n_22911;
wire n_22912;
wire n_22913;
wire n_22914;
wire n_22915;
wire n_22916;
wire n_22917;
wire n_22918;
wire n_22919;
wire n_22920;
wire n_22921;
wire n_22922;
wire n_22923;
wire n_22924;
wire n_22925;
wire n_22926;
wire n_22927;
wire n_22928;
wire n_22929;
wire n_22930;
wire n_22931;
wire n_22932;
wire n_22933;
wire n_22934;
wire n_22935;
wire n_22936;
wire n_22937;
wire n_22938;
wire n_22939;
wire n_22940;
wire n_22941;
wire n_22942;
wire n_22943;
wire n_22944;
wire n_22945;
wire n_22946;
wire n_22947;
wire n_22948;
wire n_22949;
wire n_22950;
wire n_22951;
wire n_22952;
wire n_22953;
wire n_22954;
wire n_22955;
wire n_22956;
wire n_22957;
wire n_22958;
wire n_22959;
wire n_22960;
wire n_22961;
wire n_22962;
wire n_22963;
wire n_22964;
wire n_22965;
wire n_22966;
wire n_22967;
wire n_22968;
wire n_22969;
wire n_22970;
wire n_22971;
wire n_22972;
wire n_22973;
wire n_22974;
wire n_22975;
wire n_22976;
wire n_22977;
wire n_22978;
wire n_22979;
wire n_22980;
wire n_22981;
wire n_22982;
wire n_22983;
wire n_22984;
wire n_22985;
wire n_22986;
wire n_22987;
wire n_22988;
wire n_22989;
wire n_22990;
wire n_22991;
wire n_22992;
wire n_22993;
wire n_22994;
wire n_22995;
wire n_22996;
wire n_22997;
wire n_22998;
wire n_22999;
wire n_23000;
wire n_23001;
wire n_23002;
wire n_23003;
wire n_23004;
wire n_23005;
wire n_23006;
wire n_23007;
wire n_23008;
wire n_23009;
wire n_23010;
wire n_23011;
wire n_23012;
wire n_23013;
wire n_23014;
wire n_23015;
wire n_23016;
wire n_23017;
wire n_23018;
wire n_23019;
wire n_23020;
wire n_23021;
wire n_23022;
wire n_23023;
wire n_23024;
wire n_23025;
wire n_23026;
wire n_23027;
wire n_23028;
wire n_23029;
wire n_23030;
wire n_23031;
wire n_23032;
wire n_23033;
wire n_23034;
wire n_23035;
wire n_23036;
wire n_23037;
wire n_23038;
wire n_23039;
wire n_23040;
wire n_23041;
wire n_23042;
wire n_23043;
wire n_23044;
wire n_23045;
wire n_23046;
wire n_23047;
wire n_23048;
wire n_23049;
wire n_23050;
wire n_23051;
wire n_23052;
wire n_23053;
wire n_23054;
wire n_23055;
wire n_23056;
wire n_23057;
wire n_23058;
wire n_23059;
wire n_23060;
wire n_23061;
wire n_23062;
wire n_23063;
wire n_23064;
wire n_23065;
wire n_23066;
wire n_23067;
wire n_23068;
wire n_23069;
wire n_23070;
wire n_23071;
wire n_23072;
wire n_23073;
wire n_23074;
wire n_23075;
wire n_23076;
wire n_23077;
wire n_23078;
wire n_23079;
wire n_23080;
wire n_23081;
wire n_23082;
wire n_23083;
wire n_23084;
wire n_23085;
wire n_23086;
wire n_23087;
wire n_23088;
wire n_23089;
wire n_23090;
wire n_23091;
wire n_23092;
wire n_23093;
wire n_23094;
wire n_23095;
wire n_23096;
wire n_23097;
wire n_23098;
wire n_23099;
wire n_23100;
wire n_23101;
wire n_23102;
wire n_23103;
wire n_23104;
wire n_23105;
wire n_23106;
wire n_23107;
wire n_23108;
wire n_23109;
wire n_23110;
wire n_23111;
wire n_23112;
wire n_23113;
wire n_23114;
wire n_23115;
wire n_23116;
wire n_23117;
wire n_23118;
wire n_23119;
wire n_23120;
wire n_23121;
wire n_23122;
wire n_23123;
wire n_23124;
wire n_23125;
wire n_23126;
wire n_23127;
wire n_23128;
wire n_23129;
wire n_23130;
wire n_23131;
wire n_23132;
wire n_23133;
wire n_23134;
wire n_23135;
wire n_23136;
wire n_23137;
wire n_23138;
wire n_23139;
wire n_23140;
wire n_23141;
wire n_23142;
wire n_23143;
wire n_23144;
wire n_23145;
wire n_23146;
wire n_23147;
wire n_23148;
wire n_23149;
wire n_23150;
wire n_23151;
wire n_23152;
wire n_23153;
wire n_23154;
wire n_23155;
wire n_23156;
wire n_23157;
wire n_23158;
wire n_23159;
wire n_23160;
wire n_23161;
wire n_23162;
wire n_23163;
wire n_23164;
wire n_23165;
wire n_23166;
wire n_23167;
wire n_23168;
wire n_23169;
wire n_23170;
wire n_23171;
wire n_23172;
wire n_23173;
wire n_23174;
wire n_23175;
wire n_23176;
wire n_23177;
wire n_23178;
wire n_23179;
wire n_23180;
wire n_23181;
wire n_23182;
wire n_23183;
wire n_23184;
wire n_23185;
wire n_23186;
wire n_23187;
wire n_23188;
wire n_23189;
wire n_23190;
wire n_23191;
wire n_23192;
wire n_23193;
wire n_23194;
wire n_23195;
wire n_23196;
wire n_23197;
wire n_23198;
wire n_23199;
wire n_23200;
wire n_23201;
wire n_23202;
wire n_23203;
wire n_23204;
wire n_23205;
wire n_23206;
wire n_23207;
wire n_23208;
wire n_23209;
wire n_23210;
wire n_23211;
wire n_23212;
wire n_23213;
wire n_23214;
wire n_23215;
wire n_23216;
wire n_23217;
wire n_23218;
wire n_23219;
wire n_23220;
wire n_23221;
wire n_23222;
wire n_23223;
wire n_23224;
wire n_23225;
wire n_23226;
wire n_23227;
wire n_23228;
wire n_23229;
wire n_23230;
wire n_23231;
wire n_23232;
wire n_23233;
wire n_23234;
wire n_23235;
wire n_23236;
wire n_23237;
wire n_23238;
wire n_23239;
wire n_23240;
wire n_23241;
wire n_23242;
wire n_23243;
wire n_23244;
wire n_23245;
wire n_23246;
wire n_23247;
wire n_23248;
wire n_23249;
wire n_23250;
wire n_23251;
wire n_23252;
wire n_23253;
wire n_23254;
wire n_23255;
wire n_23256;
wire n_23257;
wire n_23258;
wire n_23259;
wire n_23260;
wire n_23261;
wire n_23262;
wire n_23263;
wire n_23264;
wire n_23265;
wire n_23266;
wire n_23267;
wire n_23268;
wire n_23269;
wire n_23270;
wire n_23271;
wire n_23272;
wire n_23273;
wire n_23274;
wire n_23275;
wire n_23276;
wire n_23277;
wire n_23278;
wire n_23279;
wire n_23280;
wire n_23281;
wire n_23282;
wire n_23283;
wire n_23284;
wire n_23285;
wire n_23286;
wire n_23287;
wire n_23288;
wire n_23289;
wire n_23290;
wire n_23291;
wire n_23292;
wire n_23293;
wire n_23294;
wire n_23295;
wire n_23296;
wire n_23297;
wire n_23298;
wire n_23299;
wire n_23300;
wire n_23301;
wire n_23302;
wire n_23303;
wire n_23304;
wire n_23305;
wire n_23306;
wire n_23307;
wire n_23308;
wire n_23309;
wire n_23310;
wire n_23311;
wire n_23312;
wire n_23313;
wire n_23314;
wire n_23315;
wire n_23316;
wire n_23317;
wire n_23318;
wire n_23319;
wire n_23320;
wire n_23321;
wire n_23322;
wire n_23323;
wire n_23324;
wire n_23325;
wire n_23326;
wire n_23327;
wire n_23328;
wire n_23329;
wire n_23330;
wire n_23331;
wire n_23332;
wire n_23333;
wire n_23334;
wire n_23335;
wire n_23336;
wire n_23337;
wire n_23338;
wire n_23339;
wire n_23340;
wire n_23341;
wire n_23342;
wire n_23343;
wire n_23344;
wire n_23345;
wire n_23346;
wire n_23347;
wire n_23348;
wire n_23349;
wire n_23350;
wire n_23351;
wire n_23352;
wire n_23353;
wire n_23354;
wire n_23355;
wire n_23356;
wire n_23357;
wire n_23358;
wire n_23359;
wire n_23360;
wire n_23361;
wire n_23362;
wire n_23363;
wire n_23364;
wire n_23365;
wire n_23366;
wire n_23367;
wire n_23368;
wire n_23369;
wire n_23370;
wire n_23371;
wire n_23372;
wire n_23373;
wire n_23374;
wire n_23375;
wire n_23376;
wire n_23377;
wire n_23378;
wire n_23379;
wire n_23380;
wire n_23381;
wire n_23382;
wire n_23383;
wire n_23384;
wire n_23385;
wire n_23386;
wire n_23387;
wire n_23388;
wire n_23389;
wire n_23390;
wire n_23391;
wire n_23392;
wire n_23393;
wire n_23394;
wire n_23395;
wire n_23396;
wire n_23397;
wire n_23398;
wire n_23399;
wire n_23400;
wire n_23401;
wire n_23402;
wire n_23403;
wire n_23404;
wire n_23405;
wire n_23406;
wire n_23407;
wire n_23408;
wire n_23409;
wire n_23410;
wire n_23411;
wire n_23412;
wire n_23413;
wire n_23414;
wire n_23415;
wire n_23416;
wire n_23417;
wire n_23418;
wire n_23419;
wire n_23420;
wire n_23421;
wire n_23422;
wire n_23423;
wire n_23424;
wire n_23425;
wire n_23426;
wire n_23427;
wire n_23428;
wire n_23429;
wire n_23430;
wire n_23431;
wire n_23432;
wire n_23433;
wire n_23434;
wire n_23435;
wire n_23436;
wire n_23437;
wire n_23438;
wire n_23439;
wire n_23440;
wire n_23441;
wire n_23442;
wire n_23443;
wire n_23444;
wire n_23445;
wire n_23446;
wire n_23447;
wire n_23448;
wire n_23449;
wire n_23450;
wire n_23451;
wire n_23452;
wire n_23453;
wire n_23454;
wire n_23455;
wire n_23456;
wire n_23457;
wire n_23458;
wire n_23459;
wire n_23460;
wire n_23461;
wire n_23462;
wire n_23463;
wire n_23464;
wire n_23465;
wire n_23466;
wire n_23467;
wire n_23468;
wire n_23469;
wire n_23470;
wire n_23471;
wire n_23472;
wire n_23473;
wire n_23474;
wire n_23475;
wire n_23476;
wire n_23477;
wire n_23478;
wire n_23479;
wire n_23480;
wire n_23481;
wire n_23482;
wire n_23483;
wire n_23484;
wire n_23485;
wire n_23486;
wire n_23487;
wire n_23488;
wire n_23489;
wire n_23490;
wire n_23491;
wire n_23492;
wire n_23493;
wire n_23494;
wire n_23495;
wire n_23496;
wire n_23497;
wire n_23498;
wire n_23499;
wire n_23500;
wire n_23501;
wire n_23502;
wire n_23503;
wire n_23504;
wire n_23505;
wire n_23506;
wire n_23507;
wire n_23508;
wire n_23509;
wire n_23510;
wire n_23511;
wire n_23512;
wire n_23513;
wire n_23514;
wire n_23515;
wire n_23516;
wire n_23517;
wire n_23518;
wire n_23519;
wire n_23520;
wire n_23521;
wire n_23522;
wire n_23523;
wire n_23524;
wire n_23525;
wire n_23526;
wire n_23527;
wire n_23528;
wire n_23529;
wire n_23530;
wire n_23531;
wire n_23532;
wire n_23533;
wire n_23534;
wire n_23535;
wire n_23536;
wire n_23537;
wire n_23538;
wire n_23539;
wire n_23540;
wire n_23541;
wire n_23542;
wire n_23543;
wire n_23544;
wire n_23545;
wire n_23546;
wire n_23547;
wire n_23548;
wire n_23549;
wire n_23550;
wire n_23551;
wire n_23552;
wire n_23553;
wire n_23554;
wire n_23555;
wire n_23556;
wire n_23557;
wire n_23558;
wire n_23559;
wire n_23560;
wire n_23561;
wire n_23562;
wire n_23563;
wire n_23564;
wire n_23565;
wire n_23566;
wire n_23567;
wire n_23568;
wire n_23569;
wire n_23570;
wire n_23571;
wire n_23572;
wire n_23573;
wire n_23574;
wire n_23575;
wire n_23576;
wire n_23577;
wire n_23578;
wire n_23579;
wire n_23580;
wire n_23581;
wire n_23582;
wire n_23583;
wire n_23584;
wire n_23585;
wire n_23586;
wire n_23587;
wire n_23588;
wire n_23589;
wire n_23590;
wire n_23591;
wire n_23592;
wire n_23593;
wire n_23594;
wire n_23595;
wire n_23596;
wire n_23597;
wire n_23598;
wire n_23599;
wire n_23600;
wire n_23601;
wire n_23602;
wire n_23603;
wire n_23604;
wire n_23605;
wire n_23606;
wire n_23607;
wire n_23608;
wire n_23609;
wire n_23610;
wire n_23611;
wire n_23612;
wire n_23613;
wire n_23614;
wire n_23615;
wire n_23616;
wire n_23617;
wire n_23618;
wire n_23619;
wire n_23620;
wire n_23621;
wire n_23622;
wire n_23623;
wire n_23624;
wire n_23625;
wire n_23626;
wire n_23627;
wire n_23628;
wire n_23629;
wire n_23630;
wire n_23631;
wire n_23632;
wire n_23633;
wire n_23634;
wire n_23635;
wire n_23636;
wire n_23637;
wire n_23638;
wire n_23639;
wire n_23640;
wire n_23641;
wire n_23642;
wire n_23643;
wire n_23644;
wire n_23645;
wire n_23646;
wire n_23647;
wire n_23648;
wire n_23649;
wire n_23650;
wire n_23651;
wire n_23652;
wire n_23653;
wire n_23654;
wire n_23655;
wire n_23656;
wire n_23657;
wire n_23658;
wire n_23659;
wire n_23660;
wire n_23661;
wire n_23662;
wire n_23663;
wire n_23664;
wire n_23665;
wire n_23666;
wire n_23667;
wire n_23668;
wire n_23669;
wire n_23670;
wire n_23671;
wire n_23672;
wire n_23673;
wire n_23674;
wire n_23675;
wire n_23676;
wire n_23677;
wire n_23678;
wire n_23679;
wire n_23680;
wire n_23681;
wire n_23682;
wire n_23683;
wire n_23684;
wire n_23685;
wire n_23686;
wire n_23687;
wire n_23688;
wire n_23689;
wire n_23690;
wire n_23691;
wire n_23692;
wire n_23693;
wire n_23694;
wire n_23695;
wire n_23696;
wire n_23697;
wire n_23698;
wire n_23699;
wire n_23700;
wire n_23701;
wire n_23702;
wire n_23703;
wire n_23704;
wire n_23705;
wire n_23706;
wire n_23707;
wire n_23708;
wire n_23709;
wire n_23710;
wire n_23711;
wire n_23712;
wire n_23713;
wire n_23714;
wire n_23715;
wire n_23716;
wire n_23717;
wire n_23718;
wire n_23719;
wire n_23720;
wire n_23721;
wire n_23722;
wire n_23723;
wire n_23724;
wire n_23725;
wire n_23726;
wire n_23727;
wire n_23728;
wire n_23729;
wire n_23730;
wire n_23731;
wire n_23732;
wire n_23733;
wire n_23734;
wire n_23735;
wire n_23736;
wire n_23737;
wire n_23738;
wire n_23739;
wire n_23740;
wire n_23741;
wire n_23742;
wire n_23743;
wire n_23744;
wire n_23745;
wire n_23746;
wire n_23747;
wire n_23748;
wire n_23749;
wire n_23750;
wire n_23751;
wire n_23752;
wire n_23753;
wire n_23754;
wire n_23755;
wire n_23756;
wire n_23757;
wire n_23758;
wire n_23759;
wire n_23760;
wire n_23761;
wire n_23762;
wire n_23763;
wire n_23764;
wire n_23765;
wire n_23766;
wire n_23767;
wire n_23768;
wire n_23769;
wire n_23770;
wire n_23771;
wire n_23772;
wire n_23773;
wire n_23774;
wire n_23775;
wire n_23776;
wire n_23777;
wire n_23778;
wire n_23779;
wire n_23780;
wire n_23781;
wire n_23782;
wire n_23783;
wire n_23784;
wire n_23785;
wire n_23786;
wire n_23787;
wire n_23788;
wire n_23789;
wire n_23790;
wire n_23791;
wire n_23792;
wire n_23793;
wire n_23794;
wire n_23795;
wire n_23796;
wire n_23797;
wire n_23798;
wire n_23799;
wire n_23800;
wire n_23801;
wire n_23802;
wire n_23803;
wire n_23804;
wire n_23805;
wire n_23806;
wire n_23807;
wire n_23808;
wire n_23809;
wire n_23810;
wire n_23811;
wire n_23812;
wire n_23813;
wire n_23814;
wire n_23815;
wire n_23816;
wire n_23817;
wire n_23818;
wire n_23819;
wire n_23820;
wire n_23821;
wire n_23822;
wire n_23823;
wire n_23824;
wire n_23825;
wire n_23826;
wire n_23827;
wire n_23828;
wire n_23829;
wire n_23830;
wire n_23831;
wire n_23832;
wire n_23833;
wire n_23834;
wire n_23835;
wire n_23836;
wire n_23837;
wire n_23838;
wire n_23839;
wire n_23840;
wire n_23841;
wire n_23842;
wire n_23843;
wire n_23844;
wire n_23845;
wire n_23846;
wire n_23847;
wire n_23848;
wire n_23849;
wire n_23850;
wire n_23851;
wire n_23852;
wire n_23853;
wire n_23854;
wire n_23855;
wire n_23856;
wire n_23857;
wire n_23858;
wire n_23859;
wire n_23860;
wire n_23861;
wire n_23862;
wire n_23863;
wire n_23864;
wire n_23865;
wire n_23866;
wire n_23867;
wire n_23868;
wire n_23869;
wire n_23870;
wire n_23871;
wire n_23872;
wire n_23873;
wire n_23874;
wire n_23875;
wire n_23876;
wire n_23877;
wire n_23878;
wire n_23879;
wire n_23880;
wire n_23881;
wire n_23882;
wire n_23883;
wire n_23884;
wire n_23885;
wire n_23886;
wire n_23887;
wire n_23888;
wire n_23889;
wire n_23890;
wire n_23891;
wire n_23892;
wire n_23893;
wire n_23894;
wire n_23895;
wire n_23896;
wire n_23897;
wire n_23898;
wire n_23899;
wire n_23900;
wire n_23901;
wire n_23902;
wire n_23903;
wire n_23904;
wire n_23905;
wire n_23906;
wire n_23907;
wire n_23908;
wire n_23909;
wire n_23910;
wire n_23911;
wire n_23912;
wire n_23913;
wire n_23914;
wire n_23915;
wire n_23916;
wire n_23917;
wire n_23918;
wire n_23919;
wire n_23920;
wire n_23921;
wire n_23922;
wire n_23923;
wire n_23924;
wire n_23925;
wire n_23926;
wire n_23927;
wire n_23928;
wire n_23929;
wire n_23930;
wire n_23931;
wire n_23932;
wire n_23933;
wire n_23934;
wire n_23935;
wire n_23936;
wire n_23937;
wire n_23938;
wire n_23939;
wire n_23940;
wire n_23941;
wire n_23942;
wire n_23943;
wire n_23944;
wire n_23945;
wire n_23946;
wire n_23947;
wire n_23948;
wire n_23949;
wire n_23950;
wire n_23951;
wire n_23952;
wire n_23953;
wire n_23954;
wire n_23955;
wire n_23956;
wire n_23957;
wire n_23958;
wire n_23959;
wire n_23960;
wire n_23961;
wire n_23962;
wire n_23963;
wire n_23964;
wire n_23965;
wire n_23966;
wire n_23967;
wire n_23968;
wire n_23969;
wire n_23970;
wire n_23971;
wire n_23972;
wire n_23973;
wire n_23974;
wire n_23975;
wire n_23976;
wire n_23977;
wire n_23978;
wire n_23979;
wire n_23980;
wire n_23981;
wire n_23982;
wire n_23983;
wire n_23984;
wire n_23985;
wire n_23986;
wire n_23987;
wire n_23988;
wire n_23989;
wire n_23990;
wire n_23991;
wire n_23992;
wire n_23993;
wire n_23994;
wire n_23995;
wire n_23996;
wire n_23997;
wire n_23998;
wire n_23999;
wire n_24000;
wire n_24001;
wire n_24002;
wire n_24003;
wire n_24004;
wire n_24005;
wire n_24006;
wire n_24007;
wire n_24008;
wire n_24009;
wire n_24010;
wire n_24011;
wire n_24012;
wire n_24013;
wire n_24014;
wire n_24015;
wire n_24016;
wire n_24017;
wire n_24018;
wire n_24019;
wire n_24020;
wire n_24021;
wire n_24022;
wire n_24023;
wire n_24024;
wire n_24025;
wire n_24026;
wire n_24027;
wire n_24028;
wire n_24029;
wire n_24030;
wire n_24031;
wire n_24032;
wire n_24033;
wire n_24034;
wire n_24035;
wire n_24036;
wire n_24037;
wire n_24038;
wire n_24039;
wire n_24040;
wire n_24041;
wire n_24042;
wire n_24043;
wire n_24044;
wire n_24045;
wire n_24046;
wire n_24047;
wire n_24048;
wire n_24049;
wire n_24050;
wire n_24051;
wire n_24052;
wire n_24053;
wire n_24054;
wire n_24055;
wire n_24056;
wire n_24057;
wire n_24058;
wire n_24059;
wire n_24060;
wire n_24061;
wire n_24062;
wire n_24063;
wire n_24064;
wire n_24065;
wire n_24066;
wire n_24067;
wire n_24068;
wire n_24069;
wire n_24070;
wire n_24071;
wire n_24072;
wire n_24073;
wire n_24074;
wire n_24075;
wire n_24076;
wire n_24077;
wire n_24078;
wire n_24079;
wire n_24080;
wire n_24081;
wire n_24082;
wire n_24083;
wire n_24084;
wire n_24085;
wire n_24086;
wire n_24087;
wire n_24088;
wire n_24089;
wire n_24090;
wire n_24091;
wire n_24092;
wire n_24093;
wire n_24094;
wire n_24095;
wire n_24096;
wire n_24097;
wire n_24098;
wire n_24099;
wire n_24100;
wire n_24101;
wire n_24102;
wire n_24103;
wire n_24104;
wire n_24105;
wire n_24106;
wire n_24107;
wire n_24108;
wire n_24109;
wire n_24110;
wire n_24111;
wire n_24112;
wire n_24113;
wire n_24114;
wire n_24115;
wire n_24116;
wire n_24117;
wire n_24118;
wire n_24119;
wire n_24120;
wire n_24121;
wire n_24122;
wire n_24123;
wire n_24124;
wire n_24125;
wire n_24126;
wire n_24127;
wire n_24128;
wire n_24129;
wire n_24130;
wire n_24131;
wire n_24132;
wire n_24133;
wire n_24134;
wire n_24135;
wire n_24136;
wire n_24137;
wire n_24138;
wire n_24139;
wire n_24140;
wire n_24141;
wire n_24142;
wire n_24143;
wire n_24144;
wire n_24145;
wire n_24146;
wire n_24147;
wire n_24148;
wire n_24149;
wire n_24150;
wire n_24151;
wire n_24152;
wire n_24153;
wire n_24154;
wire n_24155;
wire n_24156;
wire n_24157;
wire n_24158;
wire n_24159;
wire n_24160;
wire n_24161;
wire n_24162;
wire n_24163;
wire n_24164;
wire n_24165;
wire n_24166;
wire n_24167;
wire n_24168;
wire n_24169;
wire n_24170;
wire n_24171;
wire n_24172;
wire n_24173;
wire n_24174;
wire n_24175;
wire n_24176;
wire n_24177;
wire n_24178;
wire n_24179;
wire n_24180;
wire n_24181;
wire n_24182;
wire n_24183;
wire n_24184;
wire n_24185;
wire n_24186;
wire n_24187;
wire n_24188;
wire n_24189;
wire n_24190;
wire n_24191;
wire n_24192;
wire n_24193;
wire n_24194;
wire n_24195;
wire n_24196;
wire n_24197;
wire n_24198;
wire n_24199;
wire n_24200;
wire n_24201;
wire n_24202;
wire n_24203;
wire n_24204;
wire n_24205;
wire n_24206;
wire n_24207;
wire n_24208;
wire n_24209;
wire n_24210;
wire n_24211;
wire n_24212;
wire n_24213;
wire n_24214;
wire n_24215;
wire n_24216;
wire n_24217;
wire n_24218;
wire n_24219;
wire n_24220;
wire n_24221;
wire n_24222;
wire n_24223;
wire n_24224;
wire n_24225;
wire n_24226;
wire n_24227;
wire n_24228;
wire n_24229;
wire n_24230;
wire n_24231;
wire n_24232;
wire n_24233;
wire n_24234;
wire n_24235;
wire n_24236;
wire n_24237;
wire n_24238;
wire n_24239;
wire n_24240;
wire n_24241;
wire n_24242;
wire n_24243;
wire n_24244;
wire n_24245;
wire n_24246;
wire n_24247;
wire n_24248;
wire n_24249;
wire n_24250;
wire n_24251;
wire n_24252;
wire n_24253;
wire n_24254;
wire n_24255;
wire n_24256;
wire n_24257;
wire n_24258;
wire n_24259;
wire n_24260;
wire n_24261;
wire n_24262;
wire n_24263;
wire n_24264;
wire n_24265;
wire n_24266;
wire n_24267;
wire n_24268;
wire n_24269;
wire n_24270;
wire n_24271;
wire n_24272;
wire n_24273;
wire n_24274;
wire n_24275;
wire n_24276;
wire n_24277;
wire n_24278;
wire n_24279;
wire n_24280;
wire n_24281;
wire n_24282;
wire n_24283;
wire n_24284;
wire n_24285;
wire n_24286;
wire n_24287;
wire n_24288;
wire n_24289;
wire n_24290;
wire n_24291;
wire n_24292;
wire n_24293;
wire n_24294;
wire n_24295;
wire n_24296;
wire n_24297;
wire n_24298;
wire n_24299;
wire n_24300;
wire n_24301;
wire n_24302;
wire n_24303;
wire n_24304;
wire n_24305;
wire n_24306;
wire n_24307;
wire n_24308;
wire n_24309;
wire n_24310;
wire n_24311;
wire n_24312;
wire n_24313;
wire n_24314;
wire n_24315;
wire n_24316;
wire n_24317;
wire n_24318;
wire n_24319;
wire n_24320;
wire n_24321;
wire n_24322;
wire n_24323;
wire n_24324;
wire n_24325;
wire n_24326;
wire n_24327;
wire n_24328;
wire n_24329;
wire n_24330;
wire n_24331;
wire n_24332;
wire n_24333;
wire n_24334;
wire n_24335;
wire n_24336;
wire n_24337;
wire n_24338;
wire n_24339;
wire n_24340;
wire n_24341;
wire n_24342;
wire n_24343;
wire n_24344;
wire n_24345;
wire n_24346;
wire n_24347;
wire n_24348;
wire n_24349;
wire n_24350;
wire n_24351;
wire n_24352;
wire n_24353;
wire n_24354;
wire n_24355;
wire n_24356;
wire n_24357;
wire n_24358;
wire n_24359;
wire n_24360;
wire n_24361;
wire n_24362;
wire n_24363;
wire n_24364;
wire n_24365;
wire n_24366;
wire n_24367;
wire n_24368;
wire n_24369;
wire n_24370;
wire n_24371;
wire n_24372;
wire n_24373;
wire n_24374;
wire n_24375;
wire n_24376;
wire n_24377;
wire n_24378;
wire n_24379;
wire n_24380;
wire n_24381;
wire n_24382;
wire n_24383;
wire n_24384;
wire n_24385;
wire n_24386;
wire n_24387;
wire n_24388;
wire n_24389;
wire n_24390;
wire n_24391;
wire n_24392;
wire n_24393;
wire n_24394;
wire n_24395;
wire n_24396;
wire n_24397;
wire n_24398;
wire n_24399;
wire n_24400;
wire n_24401;
wire n_24402;
wire n_24403;
wire n_24404;
wire n_24405;
wire n_24406;
wire n_24407;
wire n_24408;
wire n_24409;
wire n_24410;
wire n_24411;
wire n_24412;
wire n_24413;
wire n_24414;
wire n_24415;
wire n_24416;
wire n_24417;
wire n_24418;
wire n_24419;
wire n_24420;
wire n_24421;
wire n_24422;
wire n_24423;
wire n_24424;
wire n_24425;
wire n_24426;
wire n_24427;
wire n_24428;
wire n_24429;
wire n_24430;
wire n_24431;
wire n_24432;
wire n_24433;
wire n_24434;
wire n_24435;
wire n_24436;
wire n_24437;
wire n_24438;
wire n_24439;
wire n_24440;
wire n_24441;
wire n_24442;
wire n_24443;
wire n_24444;
wire n_24445;
wire n_24446;
wire n_24447;
wire n_24448;
wire n_24449;
wire n_24450;
wire n_24451;
wire n_24452;
wire n_24453;
wire n_24454;
wire n_24455;
wire n_24456;
wire n_24457;
wire n_24458;
wire n_24459;
wire n_24460;
wire n_24461;
wire n_24462;
wire n_24463;
wire n_24464;
wire n_24465;
wire n_24466;
wire n_24467;
wire n_24468;
wire n_24469;
wire n_24470;
wire n_24471;
wire n_24472;
wire n_24473;
wire n_24474;
wire n_24475;
wire n_24476;
wire n_24477;
wire n_24478;
wire n_24479;
wire n_24480;
wire n_24481;
wire n_24482;
wire n_24483;
wire n_24484;
wire n_24485;
wire n_24486;
wire n_24487;
wire n_24488;
wire n_24489;
wire n_24490;
wire n_24491;
wire n_24492;
wire n_24493;
wire n_24494;
wire n_24495;
wire n_24496;
wire n_24497;
wire n_24498;
wire n_24499;
wire n_24500;
wire n_24501;
wire n_24502;
wire n_24503;
wire n_24504;
wire n_24505;
wire n_24506;
wire n_24507;
wire n_24508;
wire n_24509;
wire n_24510;
wire n_24511;
wire n_24512;
wire n_24513;
wire n_24514;
wire n_24515;
wire n_24516;
wire n_24517;
wire n_24518;
wire n_24519;
wire n_24520;
wire n_24521;
wire n_24522;
wire n_24523;
wire n_24524;
wire n_24525;
wire n_24526;
wire n_24527;
wire n_24528;
wire n_24529;
wire n_24530;
wire n_24531;
wire n_24532;
wire n_24533;
wire n_24534;
wire n_24535;
wire n_24536;
wire n_24537;
wire n_24538;
wire n_24539;
wire n_24540;
wire n_24541;
wire n_24542;
wire n_24543;
wire n_24544;
wire n_24545;
wire n_24546;
wire n_24547;
wire n_24548;
wire n_24549;
wire n_24550;
wire n_24551;
wire n_24552;
wire n_24553;
wire n_24554;
wire n_24555;
wire n_24556;
wire n_24557;
wire n_24558;
wire n_24559;
wire n_24560;
wire n_24561;
wire n_24562;
wire n_24563;
wire n_24564;
wire n_24565;
wire n_24566;
wire n_24567;
wire n_24568;
wire n_24569;
wire n_24570;
wire n_24571;
wire n_24572;
wire n_24573;
wire n_24574;
wire n_24575;
wire n_24576;
wire n_24577;
wire n_24578;
wire n_24579;
wire n_24580;
wire n_24581;
wire n_24582;
wire n_24583;
wire n_24584;
wire n_24585;
wire n_24586;
wire n_24587;
wire n_24588;
wire n_24589;
wire n_24590;
wire n_24591;
wire n_24592;
wire n_24593;
wire n_24594;
wire n_24595;
wire n_24596;
wire n_24597;
wire n_24598;
wire n_24599;
wire n_24600;
wire n_24601;
wire n_24602;
wire n_24603;
wire n_24604;
wire n_24605;
wire n_24606;
wire n_24607;
wire n_24608;
wire n_24609;
wire n_24610;
wire n_24611;
wire n_24612;
wire n_24613;
wire n_24614;
wire n_24615;
wire n_24616;
wire n_24617;
wire n_24618;
wire n_24619;
wire n_24620;
wire n_24621;
wire n_24622;
wire n_24623;
wire n_24624;
wire n_24625;
wire n_24626;
wire n_24627;
wire n_24628;
wire n_24629;
wire n_24630;
wire n_24631;
wire n_24632;
wire n_24633;
wire n_24634;
wire n_24635;
wire n_24636;
wire n_24637;
wire n_24638;
wire n_24639;
wire n_24640;
wire n_24641;
wire n_24642;
wire n_24643;
wire n_24644;
wire n_24645;
wire n_24646;
wire n_24647;
wire n_24648;
wire n_24649;
wire n_24650;
wire n_24651;
wire n_24652;
wire n_24653;
wire n_24654;
wire n_24655;
wire n_24656;
wire n_24657;
wire n_24658;
wire n_24659;
wire n_24660;
wire n_24661;
wire n_24662;
wire n_24663;
wire n_24664;
wire n_24665;
wire n_24666;
wire n_24667;
wire n_24668;
wire n_24669;
wire n_24670;
wire n_24671;
wire n_24672;
wire n_24673;
wire n_24674;
wire n_24675;
wire n_24676;
wire n_24677;
wire n_24678;
wire n_24679;
wire n_24680;
wire n_24681;
wire n_24682;
wire n_24683;
wire n_24684;
wire n_24685;
wire n_24686;
wire n_24687;
wire n_24688;
wire n_24689;
wire n_24690;
wire n_24691;
wire n_24692;
wire n_24693;
wire n_24694;
wire n_24695;
wire n_24696;
wire n_24697;
wire n_24698;
wire n_24699;
wire n_24700;
wire n_24701;
wire n_24702;
wire n_24703;
wire n_24704;
wire n_24705;
wire n_24706;
wire n_24707;
wire n_24708;
wire n_24709;
wire n_24710;
wire n_24711;
wire n_24712;
wire n_24713;
wire n_24714;
wire n_24715;
wire n_24716;
wire n_24717;
wire n_24718;
wire n_24719;
wire n_24720;
wire n_24721;
wire n_24722;
wire n_24723;
wire n_24724;
wire n_24725;
wire n_24726;
wire n_24727;
wire n_24728;
wire n_24729;
wire n_24730;
wire n_24731;
wire n_24732;
wire n_24733;
wire n_24734;
wire n_24735;
wire n_24736;
wire n_24737;
wire n_24738;
wire n_24739;
wire n_24740;
wire n_24741;
wire n_24742;
wire n_24743;
wire n_24744;
wire n_24745;
wire n_24746;
wire n_24747;
wire n_24748;
wire n_24749;
wire n_24750;
wire n_24751;
wire n_24752;
wire n_24753;
wire n_24754;
wire n_24755;
wire n_24756;
wire n_24757;
wire n_24758;
wire n_24759;
wire n_24760;
wire n_24761;
wire n_24762;
wire n_24763;
wire n_24764;
wire n_24765;
wire n_24766;
wire n_24767;
wire n_24768;
wire n_24769;
wire n_24770;
wire n_24771;
wire n_24772;
wire n_24773;
wire n_24774;
wire n_24775;
wire n_24776;
wire n_24777;
wire n_24778;
wire n_24779;
wire n_24780;
wire n_24781;
wire n_24782;
wire n_24783;
wire n_24784;
wire n_24785;
wire n_24786;
wire n_24787;
wire n_24788;
wire n_24789;
wire n_24790;
wire n_24791;
wire n_24792;
wire n_24793;
wire n_24794;
wire n_24795;
wire n_24796;
wire n_24797;
wire n_24798;
wire n_24799;
wire n_24800;
wire n_24801;
wire n_24802;
wire n_24803;
wire n_24804;
wire n_24805;
wire n_24806;
wire n_24807;
wire n_24808;
wire n_24809;
wire n_24810;
wire n_24811;
wire n_24812;
wire n_24813;
wire n_24814;
wire n_24815;
wire n_24816;
wire n_24817;
wire n_24818;
wire n_24819;
wire n_24820;
wire n_24821;
wire n_24822;
wire n_24823;
wire n_24824;
wire n_24825;
wire n_24826;
wire n_24827;
wire n_24828;
wire n_24829;
wire n_24830;
wire n_24831;
wire n_24832;
wire n_24833;
wire n_24834;
wire n_24835;
wire n_24836;
wire n_24837;
wire n_24838;
wire n_24839;
wire n_24840;
wire n_24841;
wire n_24842;
wire n_24843;
wire n_24844;
wire n_24845;
wire n_24846;
wire n_24847;
wire n_24848;
wire n_24849;
wire n_24850;
wire n_24851;
wire n_24852;
wire n_24853;
wire n_24854;
wire n_24855;
wire n_24856;
wire n_24857;
wire n_24858;
wire n_24859;
wire n_24860;
wire n_24861;
wire n_24862;
wire n_24863;
wire n_24864;
wire n_24865;
wire n_24866;
wire n_24867;
wire n_24868;
wire n_24869;
wire n_24870;
wire n_24871;
wire n_24872;
wire n_24873;
wire n_24874;
wire n_24875;
wire n_24876;
wire n_24877;
wire n_24878;
wire n_24879;
wire n_24880;
wire n_24881;
wire n_24882;
wire n_24883;
wire n_24884;
wire n_24885;
wire n_24886;
wire n_24887;
wire n_24888;
wire n_24889;
wire n_24890;
wire n_24891;
wire n_24892;
wire n_24893;
wire n_24894;
wire n_24895;
wire n_24896;
wire n_24897;
wire n_24898;
wire n_24899;
wire n_24900;
wire n_24901;
wire n_24902;
wire n_24903;
wire n_24904;
wire n_24905;
wire n_24906;
wire n_24907;
wire n_24908;
wire n_24909;
wire n_24910;
wire n_24911;
wire n_24912;
wire n_24913;
wire n_24914;
wire n_24915;
wire n_24916;
wire n_24917;
wire n_24918;
wire n_24919;
wire n_24920;
wire n_24921;
wire n_24922;
wire n_24923;
wire n_24924;
wire n_24925;
wire n_24926;
wire n_24927;
wire n_24928;
wire n_24929;
wire n_24930;
wire n_24931;
wire n_24932;
wire n_24933;
wire n_24934;
wire n_24935;
wire n_24936;
wire n_24937;
wire n_24938;
wire n_24939;
wire n_24940;
wire n_24941;
wire n_24942;
wire n_24943;
wire n_24944;
wire n_24945;
wire n_24946;
wire n_24947;
wire n_24948;
wire n_24949;
wire n_24950;
wire n_24951;
wire n_24952;
wire n_24953;
wire n_24954;
wire n_24955;
wire n_24956;
wire n_24957;
wire n_24958;
wire n_24959;
wire n_24960;
wire n_24961;
wire n_24962;
wire n_24963;
wire n_24964;
wire n_24965;
wire n_24966;
wire n_24967;
wire n_24968;
wire n_24969;
wire n_24970;
wire n_24971;
wire n_24972;
wire n_24973;
wire n_24974;
wire n_24975;
wire n_24976;
wire n_24977;
wire n_24978;
wire n_24979;
wire n_24980;
wire n_24981;
wire n_24982;
wire n_24983;
wire n_24984;
wire n_24985;
wire n_24986;
wire n_24987;
wire n_24988;
wire n_24989;
wire n_24990;
wire n_24991;
wire n_24992;
wire n_24993;
wire n_24994;
wire n_24995;
wire n_24996;
wire n_24997;
wire n_24998;
wire n_24999;
wire n_25000;
wire n_25001;
wire n_25002;
wire n_25003;
wire n_25004;
wire n_25005;
wire n_25006;
wire n_25007;
wire n_25008;
wire n_25009;
wire n_25010;
wire n_25011;
wire n_25012;
wire n_25013;
wire n_25014;
wire n_25015;
wire n_25016;
wire n_25017;
wire n_25018;
wire n_25019;
wire n_25020;
wire n_25021;
wire n_25022;
wire n_25023;
wire n_25024;
wire n_25025;
wire n_25026;
wire n_25027;
wire n_25028;
wire n_25029;
wire n_25030;
wire n_25031;
wire n_25032;
wire n_25033;
wire n_25034;
wire n_25035;
wire n_25036;
wire n_25037;
wire n_25038;
wire n_25039;
wire n_25040;
wire n_25041;
wire n_25042;
wire n_25043;
wire n_25044;
wire n_25045;
wire n_25046;
wire n_25047;
wire n_25048;
wire n_25049;
wire n_25050;
wire n_25051;
wire n_25052;
wire n_25053;
wire n_25054;
wire n_25055;
wire n_25056;
wire n_25057;
wire n_25058;
wire n_25059;
wire n_25060;
wire n_25061;
wire n_25062;
wire n_25063;
wire n_25064;
wire n_25065;
wire n_25066;
wire n_25067;
wire n_25068;
wire n_25069;
wire n_25070;
wire n_25071;
wire n_25072;
wire n_25073;
wire n_25074;
wire n_25075;
wire n_25076;
wire n_25077;
wire n_25078;
wire n_25079;
wire n_25080;
wire n_25081;
wire n_25082;
wire n_25083;
wire n_25084;
wire n_25085;
wire n_25086;
wire n_25087;
wire n_25088;
wire n_25089;
wire n_25090;
wire n_25091;
wire n_25092;
wire n_25093;
wire n_25094;
wire n_25095;
wire n_25096;
wire n_25097;
wire n_25098;
wire n_25099;
wire n_25100;
wire n_25101;
wire n_25102;
wire n_25103;
wire n_25104;
wire n_25105;
wire n_25106;
wire n_25107;
wire n_25108;
wire n_25109;
wire n_25110;
wire n_25111;
wire n_25112;
wire n_25113;
wire n_25114;
wire n_25115;
wire n_25116;
wire n_25117;
wire n_25118;
wire n_25119;
wire n_25120;
wire n_25121;
wire n_25122;
wire n_25123;
wire n_25124;
wire n_25125;
wire n_25126;
wire n_25127;
wire n_25128;
wire n_25129;
wire n_25130;
wire n_25131;
wire n_25132;
wire n_25133;
wire n_25134;
wire n_25135;
wire n_25136;
wire n_25137;
wire n_25138;
wire n_25139;
wire n_25140;
wire n_25141;
wire n_25142;
wire n_25143;
wire n_25144;
wire n_25145;
wire n_25146;
wire n_25147;
wire n_25148;
wire n_25149;
wire n_25150;
wire n_25151;
wire n_25152;
wire n_25153;
wire n_25154;
wire n_25155;
wire n_25156;
wire n_25157;
wire n_25158;
wire n_25159;
wire n_25160;
wire n_25161;
wire n_25162;
wire n_25163;
wire n_25164;
wire n_25165;
wire n_25166;
wire n_25167;
wire n_25168;
wire n_25169;
wire n_25170;
wire n_25171;
wire n_25172;
wire n_25173;
wire n_25174;
wire n_25175;
wire n_25176;
wire n_25177;
wire n_25178;
wire n_25179;
wire n_25180;
wire n_25181;
wire n_25182;
wire n_25183;
wire n_25184;
wire n_25185;
wire n_25186;
wire n_25187;
wire n_25188;
wire n_25189;
wire n_25190;
wire n_25191;
wire n_25192;
wire n_25193;
wire n_25194;
wire n_25195;
wire n_25196;
wire n_25197;
wire n_25198;
wire n_25199;
wire n_25200;
wire n_25201;
wire n_25202;
wire n_25203;
wire n_25204;
wire n_25205;
wire n_25206;
wire n_25207;
wire n_25208;
wire n_25209;
wire n_25210;
wire n_25211;
wire n_25212;
wire n_25213;
wire n_25214;
wire n_25215;
wire n_25216;
wire n_25217;
wire n_25218;
wire n_25219;
wire n_25220;
wire n_25221;
wire n_25222;
wire n_25223;
wire n_25224;
wire n_25225;
wire n_25226;
wire n_25227;
wire n_25228;
wire n_25229;
wire n_25230;
wire n_25231;
wire n_25232;
wire n_25233;
wire n_25234;
wire n_25235;
wire n_25236;
wire n_25237;
wire n_25238;
wire n_25239;
wire n_25240;
wire n_25241;
wire n_25242;
wire n_25243;
wire n_25244;
wire n_25245;
wire n_25246;
wire n_25247;
wire n_25248;
wire n_25249;
wire n_25250;
wire n_25251;
wire n_25252;
wire n_25253;
wire n_25254;
wire n_25255;
wire n_25256;
wire n_25257;
wire n_25258;
wire n_25259;
wire n_25260;
wire n_25261;
wire n_25262;
wire n_25263;
wire n_25264;
wire n_25265;
wire n_25266;
wire n_25267;
wire n_25268;
wire n_25269;
wire n_25270;
wire n_25271;
wire n_25272;
wire n_25273;
wire n_25274;
wire n_25275;
wire n_25276;
wire n_25277;
wire n_25278;
wire n_25279;
wire n_25280;
wire n_25281;
wire n_25282;
wire n_25283;
wire n_25284;
wire n_25285;
wire n_25286;
wire n_25287;
wire n_25288;
wire n_25289;
wire n_25290;
wire n_25291;
wire n_25292;
wire n_25293;
wire n_25294;
wire n_25295;
wire n_25296;
wire n_25297;
wire n_25298;
wire n_25299;
wire n_25300;
wire n_25301;
wire n_25302;
wire n_25303;
wire n_25304;
wire n_25305;
wire n_25306;
wire n_25307;
wire n_25308;
wire n_25309;
wire n_25310;
wire n_25311;
wire n_25312;
wire n_25313;
wire n_25314;
wire n_25315;
wire n_25316;
wire n_25317;
wire n_25318;
wire n_25319;
wire n_25320;
wire n_25321;
wire n_25322;
wire n_25323;
wire n_25324;
wire n_25325;
wire n_25326;
wire n_25327;
wire n_25328;
wire n_25329;
wire n_25330;
wire n_25331;
wire n_25332;
wire n_25333;
wire n_25334;
wire n_25335;
wire n_25336;
wire n_25337;
wire n_25338;
wire n_25339;
wire n_25340;
wire n_25341;
wire n_25342;
wire n_25343;
wire n_25344;
wire n_25345;
wire n_25346;
wire n_25347;
wire n_25348;
wire n_25349;
wire n_25350;
wire n_25351;
wire n_25352;
wire n_25353;
wire n_25354;
wire n_25355;
wire n_25356;
wire n_25357;
wire n_25358;
wire n_25359;
wire n_25360;
wire n_25361;
wire n_25362;
wire n_25363;
wire n_25364;
wire n_25365;
wire n_25366;
wire n_25367;
wire n_25368;
wire n_25369;
wire n_25370;
wire n_25371;
wire n_25372;
wire n_25373;
wire n_25374;
wire n_25375;
wire n_25376;
wire n_25377;
wire n_25378;
wire n_25379;
wire n_25380;
wire n_25381;
wire n_25382;
wire n_25383;
wire n_25384;
wire n_25385;
wire n_25386;
wire n_25387;
wire n_25388;
wire n_25389;
wire n_25390;
wire n_25391;
wire n_25392;
wire n_25393;
wire n_25394;
wire n_25395;
wire n_25396;
wire n_25397;
wire n_25398;
wire n_25399;
wire n_25400;
wire n_25401;
wire n_25402;
wire n_25403;
wire n_25404;
wire n_25405;
wire n_25406;
wire n_25407;
wire n_25408;
wire n_25409;
wire n_25410;
wire n_25411;
wire n_25412;
wire n_25413;
wire n_25414;
wire n_25415;
wire n_25416;
wire n_25417;
wire n_25418;
wire n_25419;
wire n_25420;
wire n_25421;
wire n_25422;
wire n_25423;
wire n_25424;
wire n_25425;
wire n_25426;
wire n_25427;
wire n_25428;
wire n_25429;
wire n_25430;
wire n_25431;
wire n_25432;
wire n_25433;
wire n_25434;
wire n_25435;
wire n_25436;
wire n_25437;
wire n_25438;
wire n_25439;
wire n_25440;
wire n_25441;
wire n_25442;
wire n_25443;
wire n_25444;
wire n_25445;
wire n_25446;
wire n_25447;
wire n_25448;
wire n_25449;
wire n_25450;
wire n_25451;
wire n_25452;
wire n_25453;
wire n_25454;
wire n_25455;
wire n_25456;
wire n_25457;
wire n_25458;
wire n_25459;
wire n_25460;
wire n_25461;
wire n_25462;
wire n_25463;
wire n_25464;
wire n_25465;
wire n_25466;
wire n_25467;
wire n_25468;
wire n_25469;
wire n_25470;
wire n_25471;
wire n_25472;
wire n_25473;
wire n_25474;
wire n_25475;
wire n_25476;
wire n_25477;
wire n_25478;
wire n_25479;
wire n_25480;
wire n_25481;
wire n_25482;
wire n_25483;
wire n_25484;
wire n_25485;
wire n_25486;
wire n_25487;
wire n_25488;
wire n_25489;
wire n_25490;
wire n_25491;
wire n_25492;
wire n_25493;
wire n_25494;
wire n_25495;
wire n_25496;
wire n_25497;
wire n_25498;
wire n_25499;
wire n_25500;
wire n_25501;
wire n_25502;
wire n_25503;
wire n_25504;
wire n_25505;
wire n_25506;
wire n_25507;
wire n_25508;
wire n_25509;
wire n_25510;
wire n_25511;
wire n_25512;
wire n_25513;
wire n_25514;
wire n_25515;
wire n_25516;
wire n_25517;
wire n_25518;
wire n_25519;
wire n_25520;
wire n_25521;
wire n_25522;
wire n_25523;
wire n_25524;
wire n_25525;
wire n_25526;
wire n_25527;
wire n_25528;
wire n_25529;
wire n_25530;
wire n_25531;
wire n_25532;
wire n_25533;
wire n_25534;
wire n_25535;
wire n_25536;
wire n_25537;
wire n_25538;
wire n_25539;
wire n_25540;
wire n_25541;
wire n_25542;
wire n_25543;
wire n_25544;
wire n_25545;
wire n_25546;
wire n_25547;
wire n_25548;
wire n_25549;
wire n_25550;
wire n_25551;
wire n_25552;
wire n_25553;
wire n_25554;
wire n_25555;
wire n_25556;
wire n_25557;
wire n_25558;
wire n_25559;
wire n_25560;
wire n_25561;
wire n_25562;
wire n_25563;
wire n_25564;
wire n_25565;
wire n_25566;
wire n_25567;
wire n_25568;
wire n_25569;
wire n_25570;
wire n_25571;
wire n_25572;
wire n_25573;
wire n_25574;
wire n_25575;
wire n_25576;
wire n_25577;
wire n_25578;
wire n_25579;
wire n_25580;
wire n_25581;
wire n_25582;
wire n_25583;
wire n_25584;
wire n_25585;
wire n_25586;
wire n_25587;
wire n_25588;
wire n_25589;
wire n_25590;
wire n_25591;
wire n_25592;
wire n_25593;
wire n_25594;
wire n_25595;
wire n_25596;
wire n_25597;
wire n_25598;
wire n_25599;
wire n_25600;
wire n_25601;
wire n_25602;
wire n_25603;
wire n_25604;
wire n_25605;
wire n_25606;
wire n_25607;
wire n_25608;
wire n_25609;
wire n_25610;
wire n_25611;
wire n_25612;
wire n_25613;
wire n_25614;
wire n_25615;
wire n_25616;
wire n_25617;
wire n_25618;
wire n_25619;
wire n_25620;
wire n_25621;
wire n_25622;
wire n_25623;
wire n_25624;
wire n_25625;
wire n_25626;
wire n_25627;
wire n_25628;
wire n_25629;
wire n_25630;
wire n_25631;
wire n_25632;
wire n_25633;
wire n_25634;
wire n_25635;
wire n_25636;
wire n_25637;
wire n_25638;
wire n_25639;
wire n_25640;
wire n_25641;
wire n_25642;
wire n_25643;
wire n_25644;
wire n_25645;
wire n_25646;
wire n_25647;
wire n_25648;
wire n_25649;
wire n_25650;
wire n_25651;
wire n_25652;
wire n_25653;
wire n_25654;
wire n_25655;
wire n_25656;
wire n_25657;
wire n_25658;
wire n_25659;
wire n_25660;
wire n_25661;
wire n_25662;
wire n_25663;
wire n_25664;
wire n_25665;
wire n_25666;
wire n_25667;
wire n_25668;
wire n_25669;
wire n_25670;
wire n_25671;
wire n_25672;
wire n_25673;
wire n_25674;
wire n_25675;
wire n_25676;
wire n_25677;
wire n_25678;
wire n_25679;
wire n_25680;
wire n_25681;
wire n_25682;
wire n_25683;
wire n_25684;
wire n_25685;
wire n_25686;
wire n_25687;
wire n_25688;
wire n_25689;
wire n_25690;
wire n_25691;
wire n_25692;
wire n_25693;
wire n_25694;
wire n_25695;
wire n_25696;
wire n_25697;
wire n_25698;
wire n_25699;
wire n_25700;
wire n_25701;
wire n_25702;
wire n_25703;
wire n_25704;
wire n_25705;
wire n_25706;
wire n_25707;
wire n_25708;
wire n_25709;
wire n_25710;
wire n_25711;
wire n_25712;
wire n_25713;
wire n_25714;
wire n_25715;
wire n_25716;
wire n_25717;
wire n_25718;
wire n_25719;
wire n_25720;
wire n_25721;
wire n_25722;
wire n_25723;
wire n_25724;
wire n_25725;
wire n_25726;
wire n_25727;
wire n_25728;
wire n_25729;
wire n_25730;
wire n_25731;
wire n_25732;
wire n_25733;
wire n_25734;
wire n_25735;
wire n_25736;
wire n_25737;
wire n_25738;
wire n_25739;
wire n_25740;
wire n_25741;
wire n_25742;
wire n_25743;
wire n_25744;
wire n_25745;
wire n_25746;
wire n_25747;
wire n_25748;
wire n_25749;
wire n_25750;
wire n_25751;
wire n_25752;
wire n_25753;
wire n_25754;
wire n_25755;
wire n_25756;
wire n_25757;
wire n_25758;
wire n_25759;
wire n_25760;
wire n_25761;
wire n_25762;
wire n_25763;
wire n_25764;
wire n_25765;
wire n_25766;
wire n_25767;
wire n_25768;
wire n_25769;
wire n_25770;
wire n_25771;
wire n_25772;
wire n_25773;
wire n_25774;
wire n_25775;
wire n_25776;
wire n_25777;
wire n_25778;
wire n_25779;
wire n_25780;
wire n_25781;
wire n_25782;
wire n_25783;
wire n_25784;
wire n_25785;
wire n_25786;
wire n_25787;
wire n_25788;
wire n_25789;
wire n_25790;
wire n_25791;
wire n_25792;
wire n_25793;
wire n_25794;
wire n_25795;
wire n_25796;
wire n_25797;
wire n_25798;
wire n_25799;
wire n_25800;
wire n_25801;
wire n_25802;
wire n_25803;
wire n_25804;
wire n_25805;
wire n_25806;
wire n_25807;
wire n_25808;
wire n_25809;
wire n_25810;
wire n_25811;
wire n_25812;
wire n_25813;
wire n_25814;
wire n_25815;
wire n_25816;
wire n_25817;
wire n_25818;
wire n_25819;
wire n_25820;
wire n_25821;
wire n_25822;
wire n_25823;
wire n_25824;
wire n_25825;
wire n_25826;
wire n_25827;
wire n_25828;
wire n_25829;
wire n_25830;
wire n_25831;
wire n_25832;
wire n_25833;
wire n_25834;
wire n_25835;
wire n_25836;
wire n_25837;
wire n_25838;
wire n_25839;
wire n_25840;
wire n_25841;
wire n_25842;
wire n_25843;
wire n_25844;
wire n_25845;
wire n_25846;
wire n_25847;
wire n_25848;
wire n_25849;
wire n_25850;
wire n_25851;
wire n_25852;
wire n_25853;
wire n_25854;
wire n_25855;
wire n_25856;
wire n_25857;
wire n_25858;
wire n_25859;
wire n_25860;
wire n_25861;
wire n_25862;
wire n_25863;
wire n_25864;
wire n_25865;
wire n_25866;
wire n_25867;
wire n_25868;
wire n_25869;
wire n_25870;
wire n_25871;
wire n_25872;
wire n_25873;
wire n_25874;
wire n_25875;
wire n_25876;
wire n_25877;
wire n_25878;
wire n_25879;
wire n_25880;
wire n_25881;
wire n_25882;
wire n_25883;
wire n_25884;
wire n_25885;
wire n_25886;
wire n_25887;
wire n_25888;
wire n_25889;
wire n_25890;
wire n_25891;
wire n_25892;
wire n_25893;
wire n_25894;
wire n_25895;
wire n_25896;
wire n_25897;
wire n_25898;
wire n_25899;
wire n_25900;
wire n_25901;
wire n_25902;
wire n_25903;
wire n_25904;
wire n_25905;
wire n_25906;
wire n_25907;
wire n_25908;
wire n_25909;
wire n_25910;
wire n_25911;
wire n_25912;
wire n_25913;
wire n_25914;
wire n_25915;
wire n_25916;
wire n_25917;
wire n_25918;
wire n_25919;
wire n_25920;
wire n_25921;
wire n_25922;
wire n_25923;
wire n_25924;
wire n_25925;
wire n_25926;
wire n_25927;
wire n_25928;
wire n_25929;
wire n_25930;
wire n_25931;
wire n_25932;
wire n_25933;
wire n_25934;
wire n_25935;
wire n_25936;
wire n_25937;
wire n_25938;
wire n_25939;
wire n_25940;
wire n_25941;
wire n_25942;
wire n_25943;
wire n_25944;
wire n_25945;
wire n_25946;
wire n_25947;
wire n_25948;
wire n_25949;
wire n_25950;
wire n_25951;
wire n_25952;
wire n_25953;
wire n_25954;
wire n_25955;
wire n_25956;
wire n_25957;
wire n_25958;
wire n_25959;
wire n_25960;
wire n_25961;
wire n_25962;
wire n_25963;
wire n_25964;
wire n_25965;
wire n_25966;
wire n_25967;
wire n_25968;
wire n_25969;
wire n_25970;
wire n_25971;
wire n_25972;
wire n_25973;
wire n_25974;
wire n_25975;
wire n_25976;
wire n_25977;
wire n_25978;
wire n_25979;
wire n_25980;
wire n_25981;
wire n_25982;
wire n_25983;
wire n_25984;
wire n_25985;
wire n_25986;
wire n_25987;
wire n_25988;
wire n_25989;
wire n_25990;
wire n_25991;
wire n_25992;
wire n_25993;
wire n_25994;
wire n_25995;
wire n_25996;
wire n_25997;
wire n_25998;
wire n_25999;
wire n_26000;
wire n_26001;
wire n_26002;
wire n_26003;
wire n_26004;
wire n_26005;
wire n_26006;
wire n_26007;
wire n_26008;
wire n_26009;
wire n_26010;
wire n_26011;
wire n_26012;
wire n_26013;
wire n_26014;
wire n_26015;
wire n_26016;
wire n_26017;
wire n_26018;
wire n_26019;
wire n_26020;
wire n_26021;
wire n_26022;
wire n_26023;
wire n_26024;
wire n_26025;
wire n_26026;
wire n_26027;
wire n_26028;
wire n_26029;
wire n_26030;
wire n_26031;
wire n_26032;
wire n_26033;
wire n_26034;
wire n_26035;
wire n_26036;
wire n_26037;
wire n_26038;
wire n_26039;
wire n_26040;
wire n_26041;
wire n_26042;
wire n_26043;
wire n_26044;
wire n_26045;
wire n_26046;
wire n_26047;
wire n_26048;
wire n_26049;
wire n_26050;
wire n_26051;
wire n_26052;
wire n_26053;
wire n_26054;
wire n_26055;
wire n_26056;
wire n_26057;
wire n_26058;
wire n_26059;
wire n_26060;
wire n_26061;
wire n_26062;
wire n_26063;
wire n_26064;
wire n_26065;
wire n_26066;
wire n_26067;
wire n_26068;
wire n_26069;
wire n_26070;
wire n_26071;
wire n_26072;
wire n_26073;
wire n_26074;
wire n_26075;
wire n_26076;
wire n_26077;
wire n_26078;
wire n_26079;
wire n_26080;
wire n_26081;
wire n_26082;
wire n_26083;
wire n_26084;
wire n_26085;
wire n_26086;
wire n_26087;
wire n_26088;
wire n_26089;
wire n_26090;
wire n_26091;
wire n_26092;
wire n_26093;
wire n_26094;
wire n_26095;
wire n_26096;
wire n_26097;
wire n_26098;
wire n_26099;
wire n_26100;
wire n_26101;
wire n_26102;
wire n_26103;
wire n_26104;
wire n_26105;
wire n_26106;
wire n_26107;
wire n_26108;
wire n_26109;
wire n_26110;
wire n_26111;
wire n_26112;
wire n_26113;
wire n_26114;
wire n_26115;
wire n_26116;
wire n_26117;
wire n_26118;
wire n_26119;
wire n_26120;
wire n_26121;
wire n_26122;
wire n_26123;
wire n_26124;
wire n_26125;
wire n_26126;
wire n_26127;
wire n_26128;
wire n_26129;
wire n_26130;
wire n_26131;
wire n_26132;
wire n_26133;
wire n_26134;
wire n_26135;
wire n_26136;
wire n_26137;
wire n_26138;
wire n_26139;
wire n_26140;
wire n_26141;
wire n_26142;
wire n_26143;
wire n_26144;
wire n_26145;
wire n_26146;
wire n_26147;
wire n_26148;
wire n_26149;
wire n_26150;
wire n_26151;
wire n_26152;
wire n_26153;
wire n_26154;
wire n_26155;
wire n_26156;
wire n_26157;
wire n_26158;
wire n_26159;
wire n_26160;
wire n_26161;
wire n_26162;
wire n_26163;
wire n_26164;
wire n_26165;
wire n_26166;
wire n_26167;
wire n_26168;
wire n_26169;
wire n_26170;
wire n_26171;
wire n_26172;
wire n_26173;
wire n_26174;
wire n_26175;
wire n_26176;
wire n_26177;
wire n_26178;
wire n_26179;
wire n_26180;
wire n_26181;
wire n_26182;
wire n_26183;
wire n_26184;
wire n_26185;
wire n_26186;
wire n_26187;
wire n_26188;
wire n_26189;
wire n_26190;
wire n_26191;
wire n_26192;
wire n_26193;
wire n_26194;
wire n_26195;
wire n_26196;
wire n_26197;
wire n_26198;
wire n_26199;
wire n_26200;
wire n_26201;
wire n_26202;
wire n_26203;
wire n_26204;
wire n_26205;
wire n_26206;
wire n_26207;
wire n_26208;
wire n_26209;
wire n_26210;
wire n_26211;
wire n_26212;
wire n_26213;
wire n_26214;
wire n_26215;
wire n_26216;
wire n_26217;
wire n_26218;
wire n_26219;
wire n_26220;
wire n_26221;
wire n_26222;
wire n_26223;
wire n_26224;
wire n_26225;
wire n_26226;
wire n_26227;
wire n_26228;
wire n_26229;
wire n_26230;
wire n_26231;
wire n_26232;
wire n_26233;
wire n_26234;
wire n_26235;
wire n_26236;
wire n_26237;
wire n_26238;
wire n_26239;
wire n_26240;
wire n_26241;
wire n_26242;
wire n_26243;
wire n_26244;
wire n_26245;
wire n_26246;
wire n_26247;
wire n_26248;
wire n_26249;
wire n_26250;
wire n_26251;
wire n_26252;
wire n_26253;
wire n_26254;
wire n_26255;
wire n_26256;
wire n_26257;
wire n_26258;
wire n_26259;
wire n_26260;
wire n_26261;
wire n_26262;
wire n_26263;
wire n_26264;
wire n_26265;
wire n_26266;
wire n_26267;
wire n_26268;
wire n_26269;
wire n_26270;
wire n_26271;
wire n_26272;
wire n_26273;
wire n_26274;
wire n_26275;
wire n_26276;
wire n_26277;
wire n_26278;
wire n_26279;
wire n_26280;
wire n_26281;
wire n_26282;
wire n_26283;
wire n_26284;
wire n_26285;
wire n_26286;
wire n_26287;
wire n_26288;
wire n_26289;
wire n_26290;
wire n_26291;
wire n_26292;
wire n_26293;
wire n_26294;
wire n_26295;
wire n_26296;
wire n_26297;
wire n_26298;
wire n_26299;
wire n_26300;
wire n_26301;
wire n_26302;
wire n_26303;
wire n_26304;
wire n_26305;
wire n_26306;
wire n_26307;
wire n_26308;
wire n_26309;
wire n_26310;
wire n_26311;
wire n_26312;
wire n_26313;
wire n_26314;
wire n_26315;
wire n_26316;
wire n_26317;
wire n_26318;
wire n_26319;
wire n_26320;
wire n_26321;
wire n_26322;
wire n_26323;
wire n_26324;
wire n_26325;
wire n_26326;
wire n_26327;
wire n_26328;
wire n_26329;
wire n_26330;
wire n_26331;
wire n_26332;
wire n_26333;
wire n_26334;
wire n_26335;
wire n_26336;
wire n_26337;
wire n_26338;
wire n_26339;
wire n_26340;
wire n_26341;
wire n_26342;
wire n_26343;
wire n_26344;
wire n_26345;
wire n_26346;
wire n_26347;
wire n_26348;
wire n_26349;
wire n_26350;
wire n_26351;
wire n_26352;
wire n_26353;
wire n_26354;
wire n_26355;
wire n_26356;
wire n_26357;
wire n_26358;
wire n_26359;
wire n_26360;
wire n_26361;
wire n_26362;
wire n_26363;
wire n_26364;
wire n_26365;
wire n_26366;
wire n_26367;
wire n_26368;
wire n_26369;
wire n_26370;
wire n_26371;
wire n_26372;
wire n_26373;
wire n_26374;
wire n_26375;
wire n_26376;
wire n_26377;
wire n_26378;
wire n_26379;
wire n_26380;
wire n_26381;
wire n_26382;
wire n_26383;
wire n_26384;
wire n_26385;
wire n_26386;
wire n_26387;
wire n_26388;
wire n_26389;
wire n_26390;
wire n_26391;
wire n_26392;
wire n_26393;
wire n_26394;
wire n_26395;
wire n_26396;
wire n_26397;
wire n_26398;
wire n_26399;
wire n_26400;
wire n_26401;
wire n_26402;
wire n_26403;
wire n_26404;
wire n_26405;
wire n_26406;
wire n_26407;
wire n_26408;
wire n_26409;
wire n_26410;
wire n_26411;
wire n_26412;
wire n_26413;
wire n_26414;
wire n_26415;
wire n_26416;
wire n_26417;
wire n_26418;
wire n_26419;
wire n_26420;
wire n_26421;
wire n_26422;
wire n_26423;
wire n_26424;
wire n_26425;
wire n_26426;
wire n_26427;
wire n_26428;
wire n_26429;
wire n_26430;
wire n_26431;
wire n_26432;
wire n_26433;
wire n_26434;
wire n_26435;
wire n_26436;
wire n_26437;
wire n_26438;
wire n_26439;
wire n_26440;
wire n_26441;
wire n_26442;
wire n_26443;
wire n_26444;
wire n_26445;
wire n_26446;
wire n_26447;
wire n_26448;
wire n_26449;
wire n_26450;
wire n_26451;
wire n_26452;
wire n_26453;
wire n_26454;
wire n_26455;
wire n_26456;
wire n_26457;
wire n_26458;
wire n_26459;
wire n_26460;
wire n_26461;
wire n_26462;
wire n_26463;
wire n_26464;
wire n_26465;
wire n_26466;
wire n_26467;
wire n_26468;
wire n_26469;
wire n_26470;
wire n_26471;
wire n_26472;
wire n_26473;
wire n_26474;
wire n_26475;
wire n_26476;
wire n_26477;
wire n_26478;
wire n_26479;
wire n_26480;
wire n_26481;
wire n_26482;
wire n_26483;
wire n_26484;
wire n_26485;
wire n_26486;
wire n_26487;
wire n_26488;
wire n_26489;
wire n_26490;
wire n_26491;
wire n_26492;
wire n_26493;
wire n_26494;
wire n_26495;
wire n_26496;
wire n_26497;
wire n_26498;
wire n_26499;
wire n_26500;
wire n_26501;
wire n_26502;
wire n_26503;
wire n_26504;
wire n_26505;
wire n_26506;
wire n_26507;
wire n_26508;
wire n_26509;
wire n_26510;
wire n_26511;
wire n_26512;
wire n_26513;
wire n_26514;
wire n_26515;
wire n_26516;
wire n_26517;
wire n_26518;
wire n_26519;
wire n_26520;
wire n_26521;
wire n_26522;
wire n_26523;
wire n_26524;
wire n_26525;
wire n_26526;
wire n_26527;
wire n_26528;
wire n_26529;
wire n_26530;
wire n_26531;
wire n_26532;
wire n_26533;
wire n_26534;
wire n_26535;
wire n_26536;
wire n_26537;
wire n_26538;
wire n_26539;
wire n_26540;
wire n_26541;
wire n_26542;
wire n_26543;
wire n_26544;
wire n_26545;
wire n_26546;
wire n_26547;
wire n_26548;
wire n_26549;
wire n_26550;
wire n_26551;
wire n_26552;
wire n_26553;
wire n_26554;
wire n_26555;
wire n_26556;
wire n_26557;
wire n_26558;
wire n_26559;
wire n_26560;
wire n_26561;
wire n_26562;
wire n_26563;
wire n_26564;
wire n_26565;
wire n_26566;
wire n_26567;
wire n_26568;
wire n_26569;
wire n_26570;
wire n_26571;
wire n_26572;
wire n_26573;
wire n_26574;
wire n_26575;
wire n_26576;
wire n_26577;
wire n_26578;
wire n_26579;
wire n_26580;
wire n_26581;
wire n_26582;
wire n_26583;
wire n_26584;
wire n_26585;
wire n_26586;
wire n_26587;
wire n_26588;
wire n_26589;
wire n_26590;
wire n_26591;
wire n_26592;
wire n_26593;
wire n_26594;
wire n_26595;
wire n_26596;
wire n_26597;
wire n_26598;
wire n_26599;
wire n_26600;
wire n_26601;
wire n_26602;
wire n_26603;
wire n_26604;
wire n_26605;
wire n_26606;
wire n_26607;
wire n_26608;
wire n_26609;
wire n_26610;
wire n_26611;
wire n_26612;
wire n_26613;
wire n_26614;
wire n_26615;
wire n_26616;
wire n_26617;
wire n_26618;
wire n_26619;
wire n_26620;
wire n_26621;
wire n_26622;
wire n_26623;
wire n_26624;
wire n_26625;
wire n_26626;
wire n_26627;
wire n_26628;
wire n_26629;
wire n_26630;
wire n_26631;
wire n_26632;
wire n_26633;
wire n_26634;
wire n_26635;
wire n_26636;
wire n_26637;
wire n_26638;
wire n_26639;
wire n_26640;
wire n_26641;
wire n_26642;
wire n_26643;
wire n_26644;
wire n_26645;
wire n_26646;
wire n_26647;
wire n_26648;
wire n_26649;
wire n_26650;
wire n_26651;
wire n_26652;
wire n_26653;
wire n_26654;
wire n_26655;
wire n_26656;
wire n_26657;
wire n_26658;
wire n_26659;
wire n_26660;
wire n_26661;
wire n_26662;
wire n_26663;
wire n_26664;
wire n_26665;
wire n_26666;
wire n_26667;
wire n_26668;
wire n_26669;
wire n_26670;
wire n_26671;
wire n_26672;
wire n_26673;
wire n_26674;
wire n_26675;
wire n_26676;
wire n_26677;
wire n_26678;
wire n_26679;
wire n_26680;
wire n_26681;
wire n_26682;
wire n_26683;
wire n_26684;
wire n_26685;
wire n_26686;
wire n_26687;
wire n_26688;
wire n_26689;
wire n_26690;
wire n_26691;
wire n_26692;
wire n_26693;
wire n_26694;
wire n_26695;
wire n_26696;
wire n_26697;
wire n_26698;
wire n_26699;
wire n_26700;
wire n_26701;
wire n_26702;
wire n_26703;
wire n_26704;
wire n_26705;
wire n_26706;
wire n_26707;
wire n_26708;
wire n_26709;
wire n_26710;
wire n_26711;
wire n_26712;
wire n_26713;
wire n_26714;
wire n_26715;
wire n_26716;
wire n_26717;
wire n_26718;
wire n_26719;
wire n_26720;
wire n_26721;
wire n_26722;
wire n_26723;
wire n_26724;
wire n_26725;
wire n_26726;
wire n_26727;
wire n_26728;
wire n_26729;
wire n_26730;
wire n_26731;
wire n_26732;
wire n_26733;
wire n_26734;
wire n_26735;
wire n_26736;
wire n_26737;
wire n_26738;
wire n_26739;
wire n_26740;
wire n_26741;
wire n_26742;
wire n_26743;
wire n_26744;
wire n_26745;
wire n_26746;
wire n_26747;
wire n_26748;
wire n_26749;
wire n_26750;
wire n_26751;
wire n_26752;
wire n_26753;
wire n_26754;
wire n_26755;
wire n_26756;
wire n_26757;
wire n_26758;
wire n_26759;
wire n_26760;
wire n_26761;
wire n_26762;
wire n_26763;
wire n_26764;
wire n_26765;
wire n_26766;
wire n_26767;
wire n_26768;
wire n_26769;
wire n_26770;
wire n_26771;
wire n_26772;
wire n_26773;
wire n_26774;
wire n_26775;
wire n_26776;
wire n_26777;
wire n_26778;
wire n_26779;
wire n_26780;
wire n_26781;
wire n_26782;
wire n_26783;
wire n_26784;
wire n_26785;
wire n_26786;
wire n_26787;
wire n_26788;
wire n_26789;
wire n_26790;
wire n_26791;
wire n_26792;
wire n_26793;
wire n_26794;
wire n_26795;
wire n_26796;
wire n_26797;
wire n_26798;
wire n_26799;
wire n_26800;
wire n_26801;
wire n_26802;
wire n_26803;
wire n_26804;
wire n_26805;
wire n_26806;
wire n_26807;
wire n_26808;
wire n_26809;
wire n_26810;
wire n_26811;
wire n_26812;
wire n_26813;
wire n_26814;
wire n_26815;
wire n_26816;
wire n_26817;
wire n_26818;
wire n_26819;
wire n_26820;
wire n_26821;
wire n_26822;
wire n_26823;
wire n_26824;
wire n_26825;
wire n_26826;
wire n_26827;
wire n_26828;
wire n_26829;
wire n_26830;
wire n_26831;
wire n_26832;
wire n_26833;
wire n_26834;
wire n_26835;
wire n_26836;
wire n_26837;
wire n_26838;
wire n_26839;
wire n_26840;
wire n_26841;
wire n_26842;
wire n_26843;
wire n_26844;
wire n_26845;
wire n_26846;
wire n_26847;
wire n_26848;
wire n_26849;
wire n_26850;
wire n_26851;
wire n_26852;
wire n_26853;
wire n_26854;
wire n_26855;
wire n_26856;
wire n_26857;
wire n_26858;
wire n_26859;
wire n_26860;
wire n_26861;
wire n_26862;
wire n_26863;
wire n_26864;
wire n_26865;
wire n_26866;
wire n_26867;
wire n_26868;
wire n_26869;
wire n_26870;
wire n_26871;
wire n_26872;
wire n_26873;
wire n_26874;
wire n_26875;
wire n_26876;
wire n_26877;
wire n_26878;
wire n_26879;
wire n_26880;
wire n_26881;
wire n_26882;
wire n_26883;
wire n_26884;
wire n_26885;
wire n_26886;
wire n_26887;
wire n_26888;
wire n_26889;
wire n_26890;
wire n_26891;
wire n_26892;
wire n_26893;
wire n_26894;
wire n_26895;
wire n_26896;
wire n_26897;
wire n_26898;
wire n_26899;
wire n_26900;
wire n_26901;
wire n_26902;
wire n_26903;
wire n_26904;
wire n_26905;
wire n_26906;
wire n_26907;
wire n_26908;
wire n_26909;
wire n_26910;
wire n_26911;
wire n_26912;
wire n_26913;
wire n_26914;
wire n_26915;
wire n_26916;
wire n_26917;
wire n_26918;
wire n_26919;
wire n_26920;
wire n_26921;
wire n_26922;
wire n_26923;
wire n_26924;
wire n_26925;
wire n_26926;
wire n_26927;
wire n_26928;
wire n_26929;
wire n_26930;
wire n_26931;
wire n_26932;
wire n_26933;
wire n_26934;
wire n_26935;
wire n_26936;
wire n_26937;
wire n_26938;
wire n_26939;
wire n_26940;
wire n_26941;
wire n_26942;
wire n_26943;
wire n_26944;
wire n_26945;
wire n_26946;
wire n_26947;
wire n_26948;
wire n_26949;
wire n_26950;
wire n_26951;
wire n_26952;
wire n_26953;
wire n_26954;
wire n_26955;
wire n_26956;
wire n_26957;
wire n_26958;
wire n_26959;
wire n_26960;
wire n_26961;
wire n_26962;
wire n_26963;
wire n_26964;
wire n_26965;
wire n_26966;
wire n_26967;
wire n_26968;
wire n_26969;
wire n_26970;
wire n_26971;
wire n_26972;
wire n_26973;
wire n_26974;
wire n_26975;
wire n_26976;
wire n_26977;
wire n_26978;
wire n_26979;
wire n_26980;
wire n_26981;
wire n_26982;
wire n_26983;
wire n_26984;
wire n_26985;
wire n_26986;
wire n_26987;
wire n_26988;
wire n_26989;
wire n_26990;
wire n_26991;
wire n_26992;
wire n_26993;
wire n_26994;
wire n_26995;
wire n_26996;
wire n_26997;
wire n_26998;
wire n_26999;
wire n_27000;
wire n_27001;
wire n_27002;
wire n_27003;
wire n_27004;
wire n_27005;
wire n_27006;
wire n_27007;
wire n_27008;
wire n_27009;
wire n_27010;
wire n_27011;
wire n_27012;
wire n_27013;
wire n_27014;
wire n_27015;
wire n_27016;
wire n_27017;
wire n_27018;
wire n_27019;
wire n_27020;
wire n_27021;
wire n_27022;
wire n_27023;
wire n_27024;
wire n_27025;
wire n_27026;
wire n_27027;
wire n_27028;
wire n_27029;
wire n_27030;
wire n_27031;
wire n_27032;
wire n_27033;
wire n_27034;
wire n_27035;
wire n_27036;
wire n_27037;
wire n_27038;
wire n_27039;
wire n_27040;
wire n_27041;
wire n_27042;
wire n_27043;
wire n_27044;
wire n_27045;
wire n_27046;
wire n_27047;
wire n_27048;
wire n_27049;
wire n_27050;
wire n_27051;
wire n_27052;
wire n_27053;
wire n_27054;
wire n_27055;
wire n_27056;
wire n_27057;
wire n_27058;
wire n_27059;
wire n_27060;
wire n_27061;
wire n_27062;
wire n_27063;
wire n_27064;
wire n_27065;
wire n_27066;
wire n_27067;
wire n_27068;
wire n_27069;
wire n_27070;
wire n_27071;
wire n_27072;
wire n_27073;
wire n_27074;
wire n_27075;
wire n_27076;
wire n_27077;
wire n_27078;
wire n_27079;
wire n_27080;
wire n_27081;
wire n_27082;
wire n_27083;
wire n_27084;
wire n_27085;
wire n_27086;
wire n_27087;
wire n_27088;
wire n_27089;
wire n_27090;
wire n_27091;
wire n_27092;
wire n_27093;
wire n_27094;
wire n_27095;
wire n_27096;
wire n_27097;
wire n_27098;
wire n_27099;
wire n_27100;
wire n_27101;
wire n_27102;
wire n_27103;
wire n_27104;
wire n_27105;
wire n_27106;
wire n_27107;
wire n_27108;
wire n_27109;
wire n_27110;
wire n_27111;
wire n_27112;
wire n_27113;
wire n_27114;
wire n_27115;
wire n_27116;
wire n_27117;
wire n_27118;
wire n_27119;
wire n_27120;
wire n_27121;
wire n_27122;
wire n_27123;
wire n_27124;
wire n_27125;
wire n_27126;
wire n_27127;
wire n_27128;
wire n_27129;
wire n_27130;
wire n_27131;
wire n_27132;
wire n_27133;
wire n_27134;
wire n_27135;
wire n_27136;
wire n_27137;
wire n_27138;
wire n_27139;
wire n_27140;
wire n_27141;
wire n_27142;
wire n_27143;
wire n_27144;
wire n_27145;
wire n_27146;
wire n_27147;
wire n_27148;
wire n_27149;
wire n_27150;
wire n_27151;
wire n_27152;
wire n_27153;
wire n_27154;
wire n_27155;
wire n_27156;
wire n_27157;
wire n_27158;
wire n_27159;
wire n_27160;
wire n_27161;
wire n_27162;
wire n_27163;
wire n_27164;
wire n_27165;
wire n_27166;
wire n_27167;
wire n_27168;
wire n_27169;
wire n_27170;
wire n_27171;
wire n_27172;
wire n_27173;
wire n_27174;
wire n_27175;
wire n_27176;
wire n_27177;
wire n_27178;
wire n_27179;
wire n_27180;
wire n_27181;
wire n_27182;
wire n_27183;
wire n_27184;
wire n_27185;
wire n_27186;
wire n_27187;
wire n_27188;
wire n_27189;
wire n_27190;
wire n_27191;
wire n_27192;
wire n_27193;
wire n_27194;
wire n_27195;
wire n_27196;
wire n_27197;
wire n_27198;
wire n_27199;
wire n_27200;
wire n_27201;
wire n_27202;
wire n_27203;
wire n_27204;
wire n_27205;
wire n_27206;
wire n_27207;
wire n_27208;
wire n_27209;
wire n_27210;
wire n_27211;
wire n_27212;
wire n_27213;
wire n_27214;
wire n_27215;
wire n_27216;
wire n_27217;
wire n_27218;
wire n_27219;
wire n_27220;
wire n_27221;
wire n_27222;
wire n_27223;
wire n_27224;
wire n_27225;
wire n_27226;
wire n_27227;
wire n_27228;
wire n_27229;
wire n_27230;
wire n_27231;
wire n_27232;
wire n_27233;
wire n_27234;
wire n_27235;
wire n_27236;
wire n_27237;
wire n_27238;
wire n_27239;
wire n_27240;
wire n_27241;
wire n_27242;
wire n_27243;
wire n_27244;
wire n_27245;
wire n_27246;
wire n_27247;
wire n_27248;
wire n_27249;
wire n_27250;
wire n_27251;
wire n_27252;
wire n_27253;
wire n_27254;
wire n_27255;
wire n_27256;
wire n_27257;
wire n_27258;
wire n_27259;
wire n_27260;
wire n_27261;
wire n_27262;
wire n_27263;
wire n_27264;
wire n_27265;
wire n_27266;
wire n_27267;
wire n_27268;
wire n_27269;
wire n_27270;
wire n_27271;
wire n_27272;
wire n_27273;
wire n_27274;
wire n_27275;
wire n_27276;
wire n_27277;
wire n_27278;
wire n_27279;
wire n_27280;
wire n_27281;
wire n_27282;
wire n_27283;
wire n_27284;
wire n_27285;
wire n_27286;
wire n_27287;
wire n_27288;
wire n_27289;
wire n_27290;
wire n_27291;
wire n_27292;
wire n_27293;
wire n_27294;
wire n_27295;
wire n_27296;
wire n_27297;
wire n_27298;
wire n_27299;
wire n_27300;
wire n_27301;
wire n_27302;
wire n_27303;
wire n_27304;
wire n_27305;
wire n_27306;
wire n_27307;
wire n_27308;
wire n_27309;
wire n_27310;
wire n_27311;
wire n_27312;
wire n_27313;
wire n_27314;
wire n_27315;
wire n_27316;
wire n_27317;
wire n_27318;
wire n_27319;
wire n_27320;
wire n_27321;
wire n_27322;
wire n_27323;
wire n_27324;
wire n_27325;
wire n_27326;
wire n_27327;
wire n_27328;
wire n_27329;
wire n_27330;
wire n_27331;
wire n_27332;
wire n_27333;
wire n_27334;
wire n_27335;
wire n_27336;
wire n_27337;
wire n_27338;
wire n_27339;
wire n_27340;
wire n_27341;
wire n_27342;
wire n_27343;
wire n_27344;
wire n_27345;
wire n_27346;
wire n_27347;
wire n_27348;
wire n_27349;
wire n_27350;
wire n_27351;
wire n_27352;
wire n_27353;
wire n_27354;
wire n_27355;
wire n_27356;
wire n_27357;
wire n_27358;
wire n_27359;
wire n_27360;
wire n_27361;
wire n_27362;
wire n_27363;
wire n_27364;
wire n_27365;
wire n_27366;
wire n_27367;
wire n_27368;
wire n_27369;
wire n_27370;
wire n_27371;
wire n_27372;
wire n_27373;
wire n_27374;
wire n_27375;
wire n_27376;
wire n_27377;
wire n_27378;
wire n_27379;
wire n_27380;
wire n_27381;
wire n_27382;
wire n_27383;
wire n_27384;
wire n_27385;
wire n_27386;
wire n_27387;
wire n_27388;
wire n_27389;
wire n_27390;
wire n_27391;
wire n_27392;
wire n_27393;
wire n_27394;
wire n_27395;
wire n_27396;
wire n_27397;
wire n_27398;
wire n_27399;
wire n_27400;
wire n_27401;
wire n_27402;
wire n_27403;
wire n_27404;
wire n_27405;
wire n_27406;
wire n_27407;
wire n_27408;
wire n_27409;
wire n_27410;
wire n_27411;
wire n_27412;
wire n_27413;
wire n_27414;
wire n_27415;
wire n_27416;
wire n_27417;
wire n_27418;
wire n_27419;
wire n_27420;
wire n_27421;
wire n_27422;
wire n_27423;
wire n_27424;
wire n_27425;
wire n_27426;
wire n_27427;
wire n_27428;
wire n_27429;
wire n_27430;
wire n_27431;
wire n_27432;
wire n_27433;
wire n_27434;
wire n_27435;
wire n_27436;
wire n_27437;
wire n_27438;
wire n_27439;
wire n_27440;
wire n_27441;
wire n_27442;
wire n_27443;
wire n_27444;
wire n_27445;
wire n_27446;
wire n_27447;
wire n_27448;
wire n_27449;
wire n_27450;
wire n_27451;
wire n_27452;
wire n_27453;
wire n_27454;
wire n_27455;
wire n_27456;
wire n_27457;
wire n_27458;
wire n_27459;
wire n_27460;
wire n_27461;
wire n_27462;
wire n_27463;
wire n_27464;
wire n_27465;
wire n_27466;
wire n_27467;
wire n_27468;
wire n_27469;
wire n_27470;
wire n_27471;
wire n_27472;
wire n_27473;
wire n_27474;
wire n_27475;
wire n_27476;
wire n_27477;
wire n_27478;
wire n_27479;
wire n_27480;
wire n_27481;
wire n_27482;
wire n_27483;
wire n_27484;
wire n_27485;
wire n_27486;
wire n_27487;
wire n_27488;
wire n_27489;
wire n_27490;
wire n_27491;
wire n_27492;
wire n_27493;
wire n_27494;
wire n_27495;
wire n_27496;
wire n_27497;
wire n_27498;
wire n_27499;
wire n_27500;
wire n_27501;
wire n_27502;
wire n_27503;
wire n_27504;
wire n_27505;
wire n_27506;
wire n_27507;
wire n_27508;
wire n_27509;
wire n_27510;
wire n_27511;
wire n_27512;
wire n_27513;
wire n_27514;
wire n_27515;
wire n_27516;
wire n_27517;
wire n_27518;
wire n_27519;
wire n_27520;
wire n_27521;
wire n_27522;
wire n_27523;
wire n_27524;
wire n_27525;
wire n_27526;
wire n_27527;
wire n_27528;
wire n_27529;
wire n_27530;
wire n_27531;
wire n_27532;
wire n_27533;
wire n_27534;
wire n_27535;
wire n_27536;
wire n_27537;
wire n_27538;
wire n_27539;
wire n_27540;
wire n_27541;
wire n_27542;
wire n_27543;
wire n_27544;
wire n_27545;
wire n_27546;
wire n_27547;
wire n_27548;
wire n_27549;
wire n_27550;
wire n_27551;
wire n_27552;
wire n_27553;
wire n_27554;
wire n_27555;
wire n_27556;
wire n_27557;
wire n_27558;
wire n_27559;
wire n_27560;
wire n_27561;
wire n_27562;
wire n_27563;
wire n_27564;
wire n_27565;
wire n_27566;
wire n_27567;
wire n_27568;
wire n_27569;
wire n_27570;
wire n_27571;
wire n_27572;
wire n_27573;
wire n_27574;
wire n_27575;
wire n_27576;
wire n_27577;
wire n_27578;
wire n_27579;
wire n_27580;
wire n_27581;
wire n_27582;
wire n_27583;
wire n_27584;
wire n_27585;
wire n_27586;
wire n_27587;
wire n_27588;
wire n_27589;
wire n_27590;
wire n_27591;
wire n_27592;
wire n_27593;
wire n_27594;
wire n_27595;
wire n_27596;
wire n_27597;
wire n_27598;
wire n_27599;
wire n_27600;
wire n_27601;
wire n_27602;
wire n_27603;
wire n_27604;
wire n_27605;
wire n_27606;
wire n_27607;
wire n_27608;
wire n_27609;
wire n_27610;
wire n_27611;
wire n_27612;
wire n_27613;
wire n_27614;
wire n_27615;
wire n_27616;
wire n_27617;
wire n_27618;
wire n_27619;
wire n_27620;
wire n_27621;
wire n_27622;
wire n_27623;
wire n_27624;
wire n_27625;
wire n_27626;
wire n_27627;
wire n_27628;
wire n_27629;
wire n_27630;
wire n_27631;
wire n_27632;
wire n_27633;
wire n_27634;
wire n_27635;
wire n_27636;
wire n_27637;
wire n_27638;
wire n_27639;
wire n_27640;
wire n_27641;
wire n_27642;
wire n_27643;
wire n_27644;
wire n_27645;
wire n_27646;
wire n_27647;
wire n_27648;
wire n_27649;
wire n_27650;
wire n_27651;
wire n_27652;
wire n_27653;
wire n_27654;
wire n_27655;
wire n_27656;
wire n_27657;
wire n_27658;
wire n_27659;
wire n_27660;
wire n_27661;
wire n_27662;
wire n_27663;
wire n_27664;
wire n_27665;
wire n_27666;
wire n_27667;
wire n_27668;
wire n_27669;
wire n_27670;
wire n_27671;
wire n_27672;
wire n_27673;
wire n_27674;
wire n_27675;
wire n_27676;
wire n_27677;
wire n_27678;
wire n_27679;
wire n_27680;
wire n_27681;
wire n_27682;
wire n_27683;
wire n_27684;
wire n_27685;
wire n_27686;
wire n_27687;
wire n_27688;
wire n_27689;
wire n_27690;
wire n_27691;
wire n_27692;
wire n_27693;
wire n_27694;
wire n_27695;
wire n_27696;
wire n_27697;
wire n_27698;
wire n_27699;
wire n_27700;
wire n_27701;
wire n_27702;
wire n_27703;
wire n_27704;
wire n_27705;
wire n_27706;
wire n_27707;
wire n_27708;
wire n_27709;
wire n_27710;
wire n_27711;
wire n_27712;
wire n_27713;
wire n_27714;
wire n_27715;
wire n_27716;
wire n_27717;
wire n_27718;
wire n_27719;
wire n_27720;
wire n_27721;
wire n_27722;
wire n_27723;
wire n_27724;
wire n_27725;
wire n_27726;
wire n_27727;
wire n_27728;
wire n_27729;
wire n_27730;
wire n_27731;
wire n_27732;
wire n_27733;
wire n_27734;
wire n_27735;
wire n_27736;
wire n_27737;
wire n_27738;
wire n_27739;
wire n_27740;
wire n_27741;
wire n_27742;
wire n_27743;
wire n_27744;
wire n_27745;
wire n_27746;
wire n_27747;
wire n_27748;
wire n_27749;
wire n_27750;
wire n_27751;
wire n_27752;
wire n_27753;
wire n_27754;
wire n_27755;
wire n_27756;
wire n_27757;
wire n_27758;
wire n_27759;
wire n_27760;
wire n_27761;
wire n_27762;
wire n_27763;
wire n_27764;
wire n_27765;
wire n_27766;
wire n_27767;
wire n_27768;
wire n_27769;
wire n_27770;
wire n_27771;
wire n_27772;
wire n_27773;
wire n_27774;
wire n_27775;
wire n_27776;
wire n_27777;
wire n_27778;
wire n_27779;
wire n_27780;
wire n_27781;
wire n_27782;
wire n_27783;
wire n_27784;
wire n_27785;
wire n_27786;
wire n_27787;
wire n_27788;
wire n_27789;
wire n_27790;
wire n_27791;
wire n_27792;
wire n_27793;
wire n_27794;
wire n_27795;
wire n_27796;
wire n_27797;
wire n_27798;
wire n_27799;
wire n_27800;
wire n_27801;
wire n_27802;
wire n_27803;
wire n_27804;
wire n_27805;
wire n_27806;
wire n_27807;
wire n_27808;
wire n_27809;
wire n_27810;
wire n_27811;
wire n_27812;
wire n_27813;
wire n_27814;
wire n_27815;
wire n_27816;
wire n_27817;
wire n_27818;
wire n_27819;
wire n_27820;
wire n_27821;
wire n_27822;
wire n_27823;
wire n_27824;
wire n_27825;
wire n_27826;
wire n_27827;
wire n_27828;
wire n_27829;
wire n_27830;
wire n_27831;
wire n_27832;
wire n_27833;
wire n_27834;
wire n_27835;
wire n_27836;
wire n_27837;
wire n_27838;
wire n_27839;
wire n_27840;
wire n_27841;
wire n_27842;
wire n_27843;
wire n_27844;
wire n_27845;
wire n_27846;
wire n_27847;
wire n_27848;
wire n_27849;
wire n_27850;
wire n_27851;
wire n_27852;
wire n_27853;
wire n_27854;
wire n_27855;
wire n_27856;
wire n_27857;
wire n_27858;
wire n_27859;
wire n_27860;
wire n_27861;
wire n_27862;
wire n_27863;
wire n_27864;
wire n_27865;
wire n_27866;
wire n_27867;
wire n_27868;
wire n_27869;
wire n_27870;
wire n_27871;
wire n_27872;
wire n_27873;
wire n_27874;
wire n_27875;
wire n_27876;
wire n_27877;
wire n_27878;
wire n_27879;
wire n_27880;
wire n_27881;
wire n_27882;
wire n_27883;
wire n_27884;
wire n_27885;
wire n_27886;
wire n_27887;
wire n_27888;
wire n_27889;
wire n_27890;
wire n_27891;
wire n_27892;
wire n_27893;
wire n_27894;
wire n_27895;
wire n_27896;
wire n_27897;
wire n_27898;
wire n_27899;
wire n_27900;
wire n_27901;
wire n_27902;
wire n_27903;
wire n_27904;
wire n_27905;
wire n_27906;
wire n_27907;
wire n_27908;
wire n_27909;
wire n_27910;
wire n_27911;
wire n_27912;
wire n_27913;
wire n_27914;
wire n_27915;
wire n_27916;
wire n_27917;
wire n_27918;
wire n_27919;
wire n_27920;
wire n_27921;
wire n_27922;
wire n_27923;
wire n_27924;
wire n_27925;
wire n_27926;
wire n_27927;
wire n_27928;
wire n_27929;
wire n_27930;
wire n_27931;
wire n_27932;
wire n_27933;
wire n_27934;
wire n_27935;
wire n_27936;
wire n_27937;
wire n_27938;
wire n_27939;
wire n_27940;
wire n_27941;
wire n_27942;
wire n_27943;
wire n_27944;
wire n_27945;
wire n_27946;
wire n_27947;
wire n_27948;
wire n_27949;
wire n_27950;
wire n_27951;
wire n_27952;
wire n_27953;
wire n_27954;
wire n_27955;
wire n_27956;
wire n_27957;
wire n_27958;
wire n_27959;
wire n_27960;
wire n_27961;
wire n_27962;
wire n_27963;
wire n_27964;
wire n_27965;
wire n_27966;
wire n_27967;
wire n_27968;
wire n_27969;
wire n_27970;
wire n_27971;
wire n_27972;
wire n_27973;
wire n_27974;
wire n_27975;
wire n_27976;
wire n_27977;
wire n_27978;
wire n_27979;
wire n_27980;
wire n_27981;
wire n_27982;
wire n_27983;
wire n_27984;
wire n_27985;
wire n_27986;
wire n_27987;
wire n_27988;
wire n_27989;
wire n_27990;
wire n_27991;
wire n_27992;
wire n_27993;
wire n_27994;
wire n_27995;
wire n_27996;
wire n_27997;
wire n_27998;
wire n_27999;
wire n_28000;
wire n_28001;
wire n_28002;
wire n_28003;
wire n_28004;
wire n_28005;
wire n_28006;
wire n_28007;
wire n_28008;
wire n_28009;
wire n_28010;
wire n_28011;
wire n_28012;
wire n_28013;
wire n_28014;
wire n_28015;
wire n_28016;
wire n_28017;
wire n_28018;
wire n_28019;
wire n_28020;
wire n_28021;
wire n_28022;
wire n_28023;
wire n_28024;
wire n_28025;
wire n_28026;
wire n_28027;
wire n_28028;
wire n_28029;
wire n_28030;
wire n_28031;
wire n_28032;
wire n_28033;
wire n_28034;
wire n_28035;
wire n_28036;
wire n_28037;
wire n_28038;
wire n_28039;
wire n_28040;
wire n_28041;
wire n_28042;
wire n_28043;
wire n_28044;
wire n_28045;
wire n_28046;
wire n_28047;
wire n_28048;
wire n_28049;
wire n_28050;
wire n_28051;
wire n_28052;
wire n_28053;
wire n_28054;
wire n_28055;
wire n_28056;
wire n_28057;
wire n_28058;
wire n_28059;
wire n_28060;
wire n_28061;
wire n_28062;
wire n_28063;
wire n_28064;
wire n_28065;
wire n_28066;
wire n_28067;
wire n_28068;
wire n_28069;
wire n_28070;
wire n_28071;
wire n_28072;
wire n_28073;
wire n_28074;
wire n_28075;
wire n_28076;
wire n_28077;
wire n_28078;
wire n_28079;
wire n_28080;
wire n_28081;
wire n_28082;
wire n_28083;
wire n_28084;
wire n_28085;
wire n_28086;
wire n_28087;
wire n_28088;
wire n_28089;
wire n_28090;
wire n_28091;
wire n_28092;
wire n_28093;
wire n_28094;
wire n_28095;
wire n_28096;
wire n_28097;
wire n_28098;
wire n_28099;
wire n_28100;
wire n_28101;
wire n_28102;
wire n_28103;
wire n_28104;
wire n_28105;
wire n_28106;
wire n_28107;
wire n_28108;
wire n_28109;
wire n_28110;
wire n_28111;
wire n_28112;
wire n_28113;
wire n_28114;
wire n_28115;
wire n_28116;
wire n_28117;
wire n_28118;
wire n_28119;
wire n_28120;
wire n_28121;
wire n_28122;
wire n_28123;
wire n_28124;
wire n_28125;
wire n_28126;
wire n_28127;
wire n_28128;
wire n_28129;
wire n_28130;
wire n_28131;
wire n_28132;
wire n_28133;
wire n_28134;
wire n_28135;
wire n_28136;
wire n_28137;
wire n_28138;
wire n_28139;
wire n_28140;
wire n_28141;
wire n_28142;
wire n_28143;
wire n_28144;
wire n_28145;
wire n_28146;
wire n_28147;
wire n_28148;
wire n_28149;
wire n_28150;
wire n_28151;
wire n_28152;
wire n_28153;
wire n_28154;
wire n_28155;
wire n_28156;
wire n_28157;
wire n_28158;
wire n_28159;
wire n_28160;
wire n_28161;
wire n_28162;
wire n_28163;
wire n_28164;
wire n_28165;
wire n_28166;
wire n_28167;
wire n_28168;
wire n_28169;
wire n_28170;
wire n_28171;
wire n_28172;
wire n_28173;
wire n_28174;
wire n_28175;
wire n_28176;
wire n_28177;
wire n_28178;
wire n_28179;
wire n_28180;
wire n_28181;
wire n_28182;
wire n_28183;
wire n_28184;
wire n_28185;
wire n_28186;
wire n_28187;
wire n_28188;
wire n_28189;
wire n_28190;
wire n_28191;
wire n_28192;
wire n_28193;
wire n_28194;
wire n_28195;
wire n_28196;
wire n_28197;
wire n_28198;
wire n_28199;
wire n_28200;
wire n_28201;
wire n_28202;
wire n_28203;
wire n_28204;
wire n_28205;
wire n_28206;
wire n_28207;
wire n_28208;
wire n_28209;
wire n_28210;
wire n_28211;
wire n_28212;
wire n_28213;
wire n_28214;
wire n_28215;
wire n_28216;
wire n_28217;
wire n_28218;
wire n_28219;
wire n_28220;
wire n_28221;
wire n_28222;
wire n_28223;
wire n_28224;
wire n_28225;
wire n_28226;
wire n_28227;
wire n_28228;
wire n_28229;
wire n_28230;
wire n_28231;
wire n_28232;
wire n_28233;
wire n_28234;
wire n_28235;
wire n_28236;
wire n_28237;
wire n_28238;
wire n_28239;
wire n_28240;
wire n_28241;
wire n_28242;
wire n_28243;
wire n_28244;
wire n_28245;
wire n_28246;
wire n_28247;
wire n_28248;
wire n_28249;
wire n_28250;
wire n_28251;
wire n_28252;
wire n_28253;
wire n_28254;
wire n_28255;
wire n_28256;
wire n_28257;
wire n_28258;
wire n_28259;
wire n_28260;
wire n_28261;
wire n_28262;
wire n_28263;
wire n_28264;
wire n_28265;
wire n_28266;
wire n_28267;
wire n_28268;
wire n_28269;
wire n_28270;
wire n_28271;
wire n_28272;
wire n_28273;
wire n_28274;
wire n_28275;
wire n_28276;
wire n_28277;
wire n_28278;
wire n_28279;
wire n_28280;
wire n_28281;
wire n_28282;
wire n_28283;
wire n_28284;
wire n_28285;
wire n_28286;
wire n_28287;
wire n_28288;
wire n_28289;
wire n_28290;
wire n_28291;
wire n_28292;
wire n_28293;
wire n_28294;
wire n_28295;
wire n_28296;
wire n_28297;
wire n_28298;
wire n_28299;
wire n_28300;
wire n_28301;
wire n_28302;
wire n_28303;
wire n_28304;
wire n_28305;
wire n_28306;
wire n_28307;
wire n_28308;
wire n_28309;
wire n_28310;
wire n_28311;
wire n_28312;
wire n_28313;
wire n_28314;
wire n_28315;
wire n_28316;
wire n_28317;
wire n_28318;
wire n_28319;
wire n_28320;
wire n_28321;
wire n_28322;
wire n_28323;
wire n_28324;
wire n_28325;
wire n_28326;
wire n_28327;
wire n_28328;
wire n_28329;
wire n_28330;
wire n_28331;
wire n_28332;
wire n_28333;
wire n_28334;
wire n_28335;
wire n_28336;
wire n_28337;
wire n_28338;
wire n_28339;
wire n_28340;
wire n_28341;
wire n_28342;
wire n_28343;
wire n_28344;
wire n_28345;
wire n_28346;
wire n_28347;
wire n_28348;
wire n_28349;
wire n_28350;
wire n_28351;
wire n_28352;
wire n_28353;
wire n_28354;
wire n_28355;
wire n_28356;
wire n_28357;
wire n_28358;
wire n_28359;
wire n_28360;
wire n_28361;
wire n_28362;
wire n_28363;
wire n_28364;
wire n_28365;
wire n_28366;
wire n_28367;
wire n_28368;
wire n_28369;
wire n_28370;
wire n_28371;
wire n_28372;
wire n_28373;
wire n_28374;
wire n_28375;
wire n_28376;
wire n_28377;
wire n_28378;
wire n_28379;
wire n_28380;
wire n_28381;
wire n_28382;
wire n_28383;
wire n_28384;
wire n_28385;
wire n_28386;
wire n_28387;
wire n_28388;
wire n_28389;
wire n_28390;
wire n_28391;
wire n_28392;
wire n_28393;
wire n_28394;
wire n_28395;
wire n_28396;
wire n_28397;
wire n_28398;
wire n_28399;
wire n_28400;
wire n_28401;
wire n_28402;
wire n_28403;
wire n_28404;
wire n_28405;
wire n_28406;
wire n_28407;
wire n_28408;
wire n_28409;
wire n_28410;
wire n_28411;
wire n_28412;
wire n_28413;
wire n_28414;
wire n_28415;
wire n_28416;
wire n_28417;
wire n_28418;
wire n_28419;
wire n_28420;
wire n_28421;
wire n_28422;
wire n_28423;
wire n_28424;
wire n_28425;
wire n_28426;
wire n_28427;
wire n_28428;
wire n_28429;
wire n_28430;
wire n_28431;
wire n_28432;
wire n_28433;
wire n_28434;
wire n_28435;
wire n_28436;
wire n_28437;
wire n_28438;
wire n_28439;
wire n_28440;
wire n_28441;
wire n_28442;
wire n_28443;
wire n_28444;
wire n_28445;
wire n_28446;
wire n_28447;
wire n_28448;
wire n_28449;
wire n_28450;
wire n_28451;
wire n_28452;
wire n_28453;
wire n_28454;
wire n_28455;
wire n_28456;
wire n_28457;
wire n_28458;
wire n_28459;
wire n_28460;
wire n_28461;
wire n_28462;
wire n_28463;
wire n_28464;
wire n_28465;
wire n_28466;
wire n_28467;
wire n_28468;
wire n_28469;
wire n_28470;
wire n_28471;
wire n_28472;
wire n_28473;
wire n_28474;
wire n_28475;
wire n_28476;
wire n_28477;
wire n_28478;
wire n_28479;
wire n_28480;
wire n_28481;
wire n_28482;
wire n_28483;
wire n_28484;
wire n_28485;
wire n_28486;
wire n_28487;
wire n_28488;
wire n_28489;
wire n_28490;
wire n_28491;
wire n_28492;
wire n_28493;
wire n_28494;
wire n_28495;
wire n_28496;
wire n_28497;
wire n_28498;
wire n_28499;
wire n_28500;
wire n_28501;
wire n_28502;
wire n_28503;
wire n_28504;
wire n_28505;
wire n_28506;
wire n_28507;
wire n_28508;
wire n_28509;
wire n_28510;
wire n_28511;
wire n_28512;
wire n_28513;
wire n_28514;
wire n_28515;
wire n_28516;
wire n_28517;
wire n_28518;
wire n_28519;
wire n_28520;
wire n_28521;
wire n_28522;
wire n_28523;
wire n_28524;
wire n_28525;
wire n_28526;
wire n_28527;
wire n_28528;
wire n_28529;
wire n_28530;
wire n_28531;
wire n_28532;
wire n_28533;
wire n_28534;
wire n_28535;
wire n_28536;
wire n_28537;
wire n_28538;
wire n_28539;
wire n_28540;
wire n_28541;
wire n_28542;
wire n_28543;
wire n_28544;
wire n_28545;
wire n_28546;
wire n_28547;
wire n_28548;
wire n_28549;
wire n_28550;
wire n_28551;
wire n_28552;
wire n_28553;
wire n_28554;
wire n_28555;
wire n_28556;
wire n_28557;
wire n_28558;
wire n_28559;
wire n_28560;
wire n_28561;
wire n_28562;
wire n_28563;
wire n_28564;
wire n_28565;
wire n_28566;
wire n_28567;
wire n_28568;
wire n_28569;
wire n_28570;
wire n_28571;
wire n_28572;
wire n_28573;
wire n_28574;
wire n_28575;
wire n_28576;
wire n_28577;
wire n_28578;
wire n_28579;
wire n_28580;
wire n_28581;
wire n_28582;
wire n_28583;
wire n_28584;
wire n_28585;
wire n_28586;
wire n_28587;
wire n_28588;
wire n_28589;
wire n_28590;
wire n_28591;
wire n_28592;
wire n_28593;
wire n_28594;
wire n_28595;
wire n_28596;
wire n_28597;
wire n_28598;
wire n_28599;
wire n_28600;
wire n_28601;
wire n_28602;
wire n_28603;
wire n_28604;
wire n_28605;
wire n_28606;
wire n_28607;
wire n_28608;
wire n_28609;
wire n_28610;
wire n_28611;
wire n_28612;
wire n_28613;
wire n_28614;
wire n_28615;
wire n_28616;
wire n_28617;
wire n_28618;
wire n_28619;
wire n_28620;
wire n_28621;
wire n_28622;
wire n_28623;
wire n_28624;
wire n_28625;
wire n_28626;
wire n_28627;
wire n_28628;
wire n_28629;
wire n_28630;
wire n_28631;
wire n_28632;
wire n_28633;
wire n_28634;
wire n_28635;
wire n_28636;
wire n_28637;
wire n_28638;
wire n_28639;
wire n_28640;
wire n_28641;
wire n_28642;
wire n_28643;
wire n_28644;
wire n_28645;
wire n_28646;
wire n_28647;
wire n_28648;
wire n_28649;
wire n_28650;
wire n_28651;
wire n_28652;
wire n_28653;
wire n_28654;
wire n_28655;
wire n_28656;
wire n_28657;
wire n_28658;
wire n_28659;
wire n_28660;
wire n_28661;
wire n_28662;
wire n_28663;
wire n_28664;
wire n_28665;
wire n_28666;
wire n_28667;
wire n_28668;
wire n_28669;
wire n_28670;
wire n_28671;
wire n_28672;
wire n_28673;
wire n_28674;
wire n_28675;
wire n_28676;
wire n_28677;
wire n_28678;
wire n_28679;
wire n_28680;
wire n_28681;
wire n_28682;
wire n_28683;
wire n_28684;
wire n_28685;
wire n_28686;
wire n_28687;
wire n_28688;
wire n_28689;
wire n_28690;
wire n_28691;
wire n_28692;
wire n_28693;
wire n_28694;
wire n_28695;
wire n_28696;
wire n_28697;
wire n_28698;
wire n_28699;
wire n_28700;
wire n_28701;
wire n_28702;
wire n_28703;
wire n_28704;
wire n_28705;
wire n_28706;
wire n_28707;
wire n_28708;
wire n_28709;
wire n_28710;
wire n_28711;
wire n_28712;
wire n_28713;
wire n_28714;
wire n_28715;
wire n_28716;
wire n_28717;
wire n_28718;
wire n_28719;
wire n_28720;
wire n_28721;
wire n_28722;
wire n_28723;
wire n_28724;
wire n_28725;
wire n_28726;
wire n_28727;
wire n_28728;
wire n_28729;
wire n_28730;
wire n_28731;
wire n_28732;
wire n_28733;
wire n_28734;
wire n_28735;
wire n_28736;
wire n_28737;
wire n_28738;
wire n_28739;
wire n_28740;
wire n_28741;
wire n_28742;
wire n_28743;
wire n_28744;
wire n_28745;
wire n_28746;
wire n_28747;
wire n_28748;
wire n_28749;
wire n_28750;
wire n_28751;
wire n_28752;
wire n_28753;
wire n_28754;
wire n_28755;
wire n_28756;
wire n_28757;
wire n_28758;
wire n_28759;
wire n_28760;
wire n_28761;
wire n_28762;
wire n_28763;
wire n_28764;
wire n_28765;
wire n_28766;
wire n_28767;
wire n_28768;
wire n_28769;
wire n_28770;
wire n_28771;
wire n_28772;
wire n_28773;
wire n_28774;
wire n_28775;
wire n_28776;
wire n_28777;
wire n_28778;
wire n_28779;
wire n_28780;
wire n_28781;
wire n_28782;
wire n_28783;
wire n_28784;
wire n_28785;
wire n_28786;
wire n_28787;
wire n_28788;
wire n_28789;
wire n_28790;
wire n_28791;
wire n_28792;
wire n_28793;
wire n_28794;
wire n_28795;
wire n_28796;
wire n_28797;
wire n_28798;
wire n_28799;
wire n_28800;
wire n_28801;
wire n_28802;
wire n_28803;
wire n_28804;
wire n_28805;
wire n_28806;
wire n_28807;
wire n_28808;
wire n_28809;
wire n_28810;
wire n_28811;
wire n_28812;
wire n_28813;
wire n_28814;
wire n_28815;
wire n_28816;
wire n_28817;
wire n_28818;
wire n_28819;
wire n_28820;
wire n_28821;
wire n_28822;
wire n_28823;
wire n_28824;
wire n_28825;
wire n_28826;
wire n_28827;
wire n_28828;
wire n_28829;
wire n_28830;
wire n_28831;
wire n_28832;
wire n_28833;
wire n_28834;
wire n_28835;
wire n_28836;
wire n_28837;
wire n_28838;
wire n_28839;
wire n_28840;
wire n_28841;
wire n_28842;
wire n_28843;
wire n_28844;
wire n_28845;
wire n_28846;
wire n_28847;
wire n_28848;
wire n_28849;
wire n_28850;
wire n_28851;
wire n_28852;
wire n_28853;
wire n_28854;
wire n_28855;
wire n_28856;
wire n_28857;
wire n_28858;
wire n_28859;
wire n_28860;
wire n_28861;
wire n_28862;
wire n_28863;
wire n_28864;
wire n_28865;
wire n_28866;
wire n_28867;
wire n_28868;
wire n_28869;
wire n_28870;
wire n_28871;
wire n_28872;
wire n_28873;
wire n_28874;
wire n_28875;
wire n_28876;
wire n_28877;
wire n_28878;
wire n_28879;
wire n_28880;
wire n_28881;
wire n_28882;
wire n_28883;
wire n_28884;
wire n_28885;
wire n_28886;
wire n_28887;
wire n_28888;
wire n_28889;
wire n_28890;
wire n_28891;
wire n_28892;
wire n_28893;
wire n_28894;
wire n_28895;
wire n_28896;
wire n_28897;
wire n_28898;
wire n_28899;
wire n_28900;
wire n_28901;
wire n_28902;
wire n_28903;
wire n_28904;
wire n_28905;
wire n_28906;
wire n_28907;
wire n_28908;
wire n_28909;
wire n_28910;
wire n_28911;
wire n_28912;
wire n_28913;
wire n_28914;
wire n_28915;
wire n_28916;
wire n_28917;
wire n_28918;
wire n_28919;
wire n_28920;
wire n_28921;
wire n_28922;
wire n_28923;
wire n_28924;
wire n_28925;
wire n_28926;
wire n_28927;
wire n_28928;
wire n_28929;
wire n_28930;
wire n_28931;
wire n_28932;
wire n_28933;
wire n_28934;
wire n_28935;
wire n_28936;
wire n_28937;
wire n_28938;
wire n_28939;
wire n_28940;
wire n_28941;
wire n_28942;
wire n_28943;
wire n_28944;
wire n_28945;
wire n_28946;
wire n_28947;
wire n_28948;
wire n_28949;
wire n_28950;
wire n_28951;
wire n_28952;
wire n_28953;
wire n_28954;
wire n_28955;
wire n_28956;
wire n_28957;
wire n_28958;
wire n_28959;
wire n_28960;
wire n_28961;
wire n_28962;
wire n_28963;
wire n_28964;
wire n_28965;
wire n_28966;
wire n_28967;
wire n_28968;
wire n_28969;
wire n_28970;
wire n_28971;
wire n_28972;
wire n_28973;
wire n_28974;
wire n_28975;
wire n_28976;
wire n_28977;
wire n_28978;
wire n_28979;
wire n_28980;
wire n_28981;
wire n_28982;
wire n_28983;
wire n_28984;
wire n_28985;
wire n_28986;
wire n_28987;
wire n_28988;
wire n_28989;
wire n_28990;
wire n_28991;
wire n_28992;
wire n_28993;
wire n_28994;
wire n_28995;
wire n_28996;
wire n_28997;
wire n_28998;
wire n_28999;
wire n_29000;
wire n_29001;
wire n_29002;
wire n_29003;
wire n_29004;
wire n_29005;
wire n_29006;
wire n_29007;
wire n_29008;
wire n_29009;
wire n_29010;
wire n_29011;
wire n_29012;
wire n_29013;
wire n_29014;
wire n_29015;
wire n_29016;
wire n_29017;
wire n_29018;
wire n_29019;
wire n_29020;
wire n_29021;
wire n_29022;
wire n_29023;
wire n_29024;
wire n_29025;
wire n_29026;
wire n_29027;
wire n_29028;
wire n_29029;
wire n_29030;
wire n_29031;
wire n_29032;
wire n_29033;
wire n_29034;
wire n_29035;
wire n_29036;
wire n_29037;
wire n_29038;
wire n_29039;
wire n_29040;
wire n_29041;
wire n_29042;
wire n_29043;
wire n_29044;
wire n_29045;
wire n_29046;
wire n_29047;
wire n_29048;
wire n_29049;
wire n_29050;
wire n_29051;
wire n_29052;
wire n_29053;
wire n_29054;
wire n_29055;
wire n_29056;
wire n_29057;
wire n_29058;
wire n_29059;
wire n_29060;
wire n_29061;
wire n_29062;
wire n_29063;
wire n_29064;
wire n_29065;
wire n_29066;
wire n_29067;
wire n_29068;
wire n_29069;
wire n_29070;
wire n_29071;
wire n_29072;
wire n_29073;
wire n_29074;
wire n_29075;
wire n_29076;
wire n_29077;
wire n_29078;
wire n_29079;
wire n_29080;
wire n_29081;
wire n_29082;
wire n_29083;
wire n_29084;
wire n_29085;
wire n_29086;
wire n_29087;
wire n_29088;
wire n_29089;
wire n_29090;
wire n_29091;
wire n_29092;
wire n_29093;
wire n_29094;
wire n_29095;
wire n_29096;
wire n_29097;
wire n_29098;
wire n_29099;
wire n_29100;
wire n_29101;
wire n_29102;
wire n_29103;
wire n_29104;
wire n_29105;
wire n_29106;
wire n_29107;
wire n_29108;
wire n_29109;
wire n_29110;
wire n_29111;
wire n_29112;
wire n_29113;
wire n_29114;
wire n_29115;
wire n_29116;
wire n_29117;
wire n_29118;
wire n_29119;
wire n_29120;
wire n_29121;
wire n_29122;
wire n_29123;
wire n_29124;
wire n_29125;
wire n_29126;
wire n_29127;
wire n_29128;
wire n_29129;
wire n_29130;
wire n_29131;
wire n_29132;
wire n_29133;
wire n_29134;
wire n_29135;
wire n_29136;
wire n_29137;
wire n_29138;
wire n_29139;
wire n_29140;
wire n_29141;
wire n_29142;
wire n_29143;
wire n_29144;
wire n_29145;
wire n_29146;
wire n_29147;
wire n_29148;
wire n_29149;
wire n_29150;
wire n_29151;
wire n_29152;
wire n_29153;
wire n_29154;
wire n_29155;
wire n_29156;
wire n_29157;
wire n_29158;
wire n_29159;
wire n_29160;
wire n_29161;
wire n_29162;
wire n_29163;
wire n_29164;
wire n_29165;
wire n_29166;
wire n_29167;
wire n_29168;
wire n_29169;
wire n_29170;
wire n_29171;
wire n_29172;
wire n_29173;
wire n_29174;
wire n_29175;
wire n_29176;
wire n_29177;
wire n_29178;
wire n_29179;
wire n_29180;
wire n_29181;
wire n_29182;
wire n_29183;
wire n_29184;
wire n_29185;
wire n_29186;
wire n_29187;
wire n_29188;
wire n_29189;
wire n_29190;
wire n_29191;
wire n_29192;
wire n_29193;
wire n_29194;
wire n_29195;
wire n_29196;
wire n_29197;
wire n_29198;
wire n_29199;
wire n_29200;
wire n_29201;
wire n_29202;
wire n_29203;
wire n_29204;
wire n_29205;
wire n_29206;
wire n_29207;
wire n_29208;
wire n_29209;
wire n_29210;
wire n_29211;
wire n_29212;
wire n_29213;
wire n_29214;
wire n_29215;
wire n_29216;
wire n_29217;
wire n_29218;
wire n_29219;
wire n_29220;
wire n_29221;
wire n_29222;
wire n_29223;
wire n_29224;
wire n_29225;
wire n_29226;
wire n_29227;
wire n_29228;
wire n_29229;
wire n_29230;
wire n_29231;
wire n_29232;
wire n_29233;
wire n_29234;
wire n_29235;
wire n_29236;
wire n_29237;
wire n_29238;
wire n_29239;
wire n_29240;
wire n_29241;
wire n_29242;
wire n_29243;
wire n_29244;
wire n_29245;
wire n_29246;
wire n_29247;
wire n_29248;
wire n_29249;
wire n_29250;
wire n_29251;
wire n_29252;
wire n_29253;
wire n_29254;
wire n_29255;
wire n_29256;
wire n_29257;
wire n_29258;
wire n_29259;
wire n_29260;
wire n_29261;
wire n_29262;
wire n_29263;
wire n_29264;
wire n_29265;
wire n_29266;
wire n_29267;
wire n_29268;
wire n_29269;
wire n_29270;
wire n_29271;
wire n_29272;
wire n_29273;
wire n_29274;
wire n_29275;
wire n_29276;
wire n_29277;
wire n_29278;
wire n_29279;
wire n_29280;
wire n_29281;
wire n_29282;
wire n_29283;
wire n_29284;
wire n_29285;
wire n_29286;
wire n_29287;
wire n_29288;
wire n_29289;
wire n_29290;
wire n_29291;
wire n_29292;
wire n_29293;
wire n_29294;
wire n_29295;
wire n_29296;
wire n_29297;
wire n_29298;
wire n_29299;
wire n_29300;
wire n_29301;
wire n_29302;
wire n_29303;
wire n_29304;
wire n_29305;
wire n_29306;
wire n_29307;
wire n_29308;
wire n_29309;
wire n_29310;
wire n_29311;
wire n_29312;
wire n_29313;
wire n_29314;
wire n_29315;
wire n_29316;
wire n_29317;
wire n_29318;
wire n_29319;
wire n_29320;
wire n_29321;
wire n_29322;
wire n_29323;
wire n_29324;
wire n_29325;
wire n_29326;
wire n_29327;
wire n_29328;
wire n_29329;
wire n_29330;
wire n_29331;
wire n_29332;
wire n_29333;
wire n_29334;
wire n_29335;
wire n_29336;
wire n_29337;
wire n_29338;
wire n_29339;
wire n_29340;
wire n_29341;
wire n_29342;
wire n_29343;
wire n_29344;
wire n_29345;
wire n_29346;
wire n_29347;
wire n_29348;
wire n_29349;
wire n_29350;
wire n_29351;
wire n_29352;
wire n_29353;
wire n_29354;
wire n_29355;
wire n_29356;
wire n_29357;
wire n_29358;
wire n_29359;
wire n_29360;
wire n_29361;
wire n_29362;
wire n_29363;
wire n_29364;
wire n_29365;
wire n_29366;
wire n_29367;
wire n_29368;
wire n_29369;
wire n_29370;
wire n_29371;
wire n_29372;
wire n_29373;
wire n_29374;
wire n_29375;
wire n_29376;
wire n_29377;
wire n_29378;
wire n_29379;
wire n_29380;
wire n_29381;
wire n_29382;
wire n_29383;
wire n_29384;
wire n_29385;
wire n_29386;
wire n_29387;
wire n_29388;
wire n_29389;
wire n_29390;
wire n_29391;
wire n_29392;
wire n_29393;
wire n_29394;
wire n_29395;
wire n_29396;
wire n_29397;
wire n_29398;
wire n_29399;
wire n_29400;
wire n_29401;
wire n_29402;
wire n_29403;
wire n_29404;
wire n_29405;
wire n_29406;
wire n_29407;
wire n_29408;
wire n_29409;
wire n_29410;
wire n_29411;
wire n_29412;
wire n_29413;
wire n_29414;
wire n_29415;
wire n_29416;
wire n_29417;
wire n_29418;
wire n_29419;
wire n_29420;
wire n_29421;
wire n_29422;
wire n_29423;
wire n_29424;
wire n_29425;
wire n_29426;
wire n_29427;
wire n_29428;
wire n_29429;
wire n_29430;
wire n_29431;
wire n_29432;
wire n_29433;
wire n_29434;
wire n_29435;
wire n_29436;
wire n_29437;
wire n_29438;
wire n_29439;
wire n_29440;
wire n_29441;
wire n_29442;
wire n_29443;
wire n_29444;
wire n_29445;
wire n_29446;
wire n_29447;
wire n_29448;
wire n_29449;
wire n_29450;
wire n_29451;
wire n_29452;
wire n_29453;
wire n_29454;
wire n_29455;
wire n_29456;
wire n_29457;
wire n_29458;
wire n_29459;
wire n_29460;
wire n_29461;
wire n_29462;
wire n_29463;
wire n_29464;
wire n_29465;
wire n_29466;
wire n_29467;
wire n_29468;
wire n_29469;
wire n_29470;
wire n_29471;
wire n_29472;
wire n_29473;
wire n_29474;
wire n_29475;
wire n_29476;
wire n_29477;
wire n_29478;
wire n_29479;
wire n_29480;
wire n_29481;
wire n_29482;
wire n_29483;
wire n_29484;
wire n_29485;
wire n_29486;
wire n_29487;
wire n_29488;
wire n_29489;
wire n_29490;
wire n_29491;
wire n_29492;
wire n_29493;
wire n_29494;
wire n_29495;
wire n_29496;
wire n_29497;
wire n_29498;
wire n_29499;
wire n_29500;
wire n_29501;
wire n_29502;
wire n_29503;
wire n_29504;
wire n_29505;
wire n_29506;
wire n_29507;
wire n_29508;
wire n_29509;
wire n_29510;
wire n_29511;
wire n_29512;
wire n_29513;
wire n_29514;
wire n_29515;
wire n_29516;
wire n_29517;
wire n_29518;
wire n_29519;
wire n_29520;
wire n_29521;
wire n_29522;
wire n_29523;
wire n_29524;
wire n_29525;
wire n_29526;
wire n_29527;
wire n_29528;
wire n_29529;
wire n_29530;
wire n_29531;
wire n_29532;
wire n_29533;
wire n_29534;
wire n_29535;
wire n_29536;
wire n_29537;
wire n_29538;
wire n_29539;
wire n_29540;
wire n_29541;
wire n_29542;
wire n_29543;
wire n_29544;
wire n_29545;
wire n_29546;
wire n_29547;
wire n_29548;
wire n_29549;
wire n_29550;
wire n_29551;
wire n_29552;
wire n_29553;
wire n_29554;
wire n_29555;
wire n_29556;
wire n_29557;
wire n_29558;
wire n_29559;
wire n_29560;
wire n_29561;
wire n_29562;
wire n_29563;
wire n_29564;
wire n_29565;
wire n_29566;
wire n_29567;
wire n_29568;
wire n_29569;
wire n_29570;
wire n_29571;
wire n_29572;
wire n_29573;
wire n_29574;
wire n_29575;
wire n_29576;
wire n_29577;
wire n_29578;
wire n_29579;
wire n_29580;
wire n_29581;
wire n_29582;
wire n_29583;
wire n_29584;
wire n_29585;
wire n_29586;
wire n_29587;
wire n_29588;
wire n_29589;
wire n_29590;
wire n_29591;
wire n_29592;
wire n_29593;
wire n_29594;
wire n_29595;
wire n_29596;
wire n_29597;
wire n_29598;
wire n_29599;
wire n_29600;
wire n_29601;
wire n_29602;
wire n_29603;
wire n_29604;
wire n_29605;
wire n_29606;
wire n_29607;
wire n_29608;
wire n_29609;
wire n_29610;
wire n_29611;
wire n_29612;
wire n_29613;
wire n_29614;
wire n_29615;
wire n_29616;
wire n_29617;
wire n_29618;
wire n_29619;
wire n_29620;
wire n_29621;
wire n_29622;
wire n_29623;
wire n_29624;
wire n_29625;
wire n_29626;
wire n_29627;
wire n_29628;
wire n_29629;
wire n_29630;
wire n_29631;
wire n_29632;
wire n_29633;
wire n_29634;
wire n_29635;
wire n_29636;
wire n_29637;
wire n_29638;
wire n_29639;
wire n_29640;
wire n_29641;
wire n_29642;
wire n_29643;
wire n_29644;
wire n_29645;
wire n_29646;
wire n_29647;
wire n_29648;
wire n_29649;
wire n_29650;
wire n_29651;
wire n_29652;
wire n_29653;
wire n_29654;
wire n_29655;
wire n_29656;
wire n_29657;
wire n_29658;
wire n_29659;
wire n_29660;
wire n_29661;
wire n_29662;
wire n_29663;
wire n_29664;
wire n_29665;
wire n_29666;
wire n_29667;
wire n_29668;
wire n_29669;
wire n_29670;
wire n_29671;
wire n_29672;
wire n_29673;
wire n_29674;
wire n_29675;
wire n_29676;
wire n_29677;
wire n_29678;
wire n_29679;
wire n_29680;
wire n_29681;
wire n_29682;
wire n_29683;
wire n_29684;
wire n_29685;
wire n_29686;
wire n_29687;
wire n_29688;
wire n_29689;
wire n_29690;
wire n_29691;
wire n_29692;
wire n_29693;
wire n_29694;
wire n_29695;
wire n_29696;
wire n_29697;
wire n_29698;
wire n_29699;
wire n_29700;
wire n_29701;
wire n_29702;
wire n_29703;
wire n_29704;
wire n_29705;
wire n_29706;
wire n_29707;
wire n_29708;
wire n_29709;
wire n_29710;
wire n_29711;
wire n_29712;
wire n_29713;
wire n_29714;
wire n_29715;
wire n_29716;
wire n_29717;
wire n_29718;
wire n_29719;
wire n_29720;
wire n_29721;
wire n_29722;
wire n_29723;
wire n_29724;
wire n_29725;
wire n_29726;
wire n_29727;
wire n_29728;
wire n_29729;
wire n_29730;
wire n_29731;
wire n_29732;
wire n_29733;
wire n_29734;
wire n_29735;
wire n_29736;
wire n_29737;
wire n_29738;
wire n_29739;
wire n_29740;
wire n_29741;
wire n_29742;
wire n_29743;
wire n_29744;
wire n_29745;
wire n_29746;
wire n_29747;
wire n_29748;
wire n_29749;
wire n_29750;
wire n_29751;
wire n_29752;
wire n_29753;
wire n_29754;
wire n_29755;
wire n_29756;
wire n_29757;
wire n_29758;
wire n_29759;
wire n_29760;
wire n_29761;
wire n_29762;
wire n_29763;
wire n_29764;
wire n_29765;
wire n_29766;
wire n_29767;
wire n_29768;
wire n_29769;
wire n_29770;
wire n_29771;
wire n_29772;
wire n_29773;
wire n_29774;
wire n_29775;
wire n_29776;
wire n_29777;
wire n_29778;
wire n_29779;
wire n_29780;
wire n_29781;
wire n_29782;
wire n_29783;
wire n_29784;
wire n_29785;
wire n_29786;
wire n_29787;
wire n_29788;
wire n_29789;
wire n_29790;
wire n_29791;
wire n_29792;
wire n_29793;
wire n_29794;
wire n_29795;
wire n_29796;
wire n_29797;
wire n_29798;
wire n_29799;
wire n_29800;
wire n_29801;
wire n_29802;
wire n_29803;
wire n_29804;
wire n_29805;
wire n_29806;
wire n_29807;
wire n_29808;
wire n_29809;
wire n_29810;
wire n_29811;
wire n_29812;
wire n_29813;
wire n_29814;
wire n_29815;
wire n_29816;
wire n_29817;
wire n_29818;
wire n_29819;
wire n_29820;
wire n_29821;
wire n_29822;
wire n_29823;
wire n_29824;
wire n_29825;
wire n_29826;
wire n_29827;
wire n_29828;
wire n_29829;
wire n_29830;
wire n_29831;
wire n_29832;
wire n_29833;
wire n_29834;
wire n_29835;
wire n_29836;
wire n_29837;
wire n_29838;
wire n_29839;
wire n_29840;
wire n_29841;
wire n_29842;
wire n_29843;
wire n_29844;
wire n_29845;
wire n_29846;
wire n_29847;
wire n_29848;
wire n_29849;
wire n_29850;
wire n_29851;
wire n_29852;
wire n_29853;
wire n_29854;
wire n_29855;
wire n_29856;
wire n_29857;
wire n_29858;
wire n_29859;
wire n_29860;
wire n_29861;
wire n_29862;
wire n_29863;
wire n_29864;
wire n_29865;
wire n_29866;
wire n_29867;
wire n_29868;
wire n_29869;
wire n_29870;
wire n_29871;
wire n_29872;
wire n_29873;
wire n_29874;
wire n_29875;
wire n_29876;
wire n_29877;
wire n_29878;
wire n_29879;
wire n_29880;
wire n_29881;
wire n_29882;
wire n_29883;
wire n_29884;
wire n_29885;
wire n_29886;
wire n_29887;
wire n_29888;
wire n_29889;
wire n_29890;
wire n_29891;
wire n_29892;
wire n_29893;
wire n_29894;
wire n_29895;
wire n_29896;
wire n_29897;
wire n_29898;
wire n_29899;
wire n_29900;
wire n_29901;
wire n_29902;
wire n_29903;
wire n_29904;
wire n_29905;
wire n_29906;
wire n_29907;
wire n_29908;
wire n_29909;
wire n_29910;
wire n_29911;
wire n_29912;
wire n_29913;
wire n_29914;
wire n_29915;
wire n_29916;
wire n_29917;
wire n_29918;
wire n_29919;
wire n_29920;
wire n_29921;
wire n_29922;
wire n_29923;
wire n_29924;
wire n_29925;
wire n_29926;
wire n_29927;
wire n_29928;
wire n_29929;
wire n_29930;
wire n_29931;
wire n_29932;
wire n_29933;
wire n_29934;
wire n_29935;
wire n_29936;
wire n_29937;
wire n_29938;
wire n_29939;
wire n_29940;
wire n_29941;
wire n_29942;
wire n_29943;
wire n_29944;
wire n_29945;
wire n_29946;
wire n_29947;
wire n_29948;
wire n_29949;
wire n_29950;
wire n_29951;
wire n_29952;
wire n_29953;
wire n_29954;
wire n_29955;
wire n_29956;
wire n_29957;
wire n_29958;
wire n_29959;
wire n_29960;
wire n_29961;
wire n_29962;
wire n_29963;
wire n_29964;
wire n_29965;
wire n_29966;
wire n_29967;
wire n_29968;
wire n_29969;
wire n_29970;
wire n_29971;
wire n_29972;
wire n_29973;
wire n_29974;
wire n_29975;
wire n_29976;
wire n_29977;
wire n_29978;
wire n_29979;
wire n_29980;
wire n_29981;
wire n_29982;
wire n_29983;
wire n_29984;
wire n_29985;
wire n_29986;
wire n_29987;
wire n_29988;
wire n_29989;
wire n_29990;
wire n_29991;
wire n_29992;
wire n_29993;
wire n_29994;
wire n_29995;
wire n_29996;
wire n_29997;
wire n_29998;
wire n_29999;
wire n_30000;
wire n_30001;
wire n_30002;
wire n_30003;
wire n_30004;
wire n_30005;
wire n_30006;
wire n_30007;
wire n_30008;
wire n_30009;
wire n_30010;
wire n_30011;
wire n_30012;
wire n_30013;
wire n_30014;
wire n_30015;
wire n_30016;
wire n_30017;
wire n_30018;
wire n_30019;
wire n_30020;
wire n_30021;
wire n_30022;
wire n_30023;
wire n_30024;
wire n_30025;
wire n_30026;
wire n_30027;
wire n_30028;
wire n_30029;
wire n_30030;
wire n_30031;
wire n_30032;
wire n_30033;
wire n_30034;
wire n_30035;
wire n_30036;
wire n_30037;
wire n_30038;
wire n_30039;
wire n_30040;
wire n_30041;
wire n_30042;
wire n_30043;
wire n_30044;
wire n_30045;
wire n_30046;
wire n_30047;
wire n_30048;
wire n_30049;
wire n_30050;
wire n_30051;
wire n_30052;
wire n_30053;
wire n_30054;
wire n_30055;
wire n_30056;
wire n_30057;
wire n_30058;
wire n_30059;
wire n_30060;
wire n_30061;
wire n_30062;
wire n_30063;
wire n_30064;
wire n_30065;
wire n_30066;
wire n_30067;
wire n_30068;
wire n_30069;
wire n_30070;
wire n_30071;
wire n_30072;
wire n_30073;
wire n_30074;
wire n_30075;
wire n_30076;
wire n_30077;
wire n_30078;
wire n_30079;
wire n_30080;
wire n_30081;
wire n_30082;
wire n_30083;
wire n_30084;
wire n_30085;
wire n_30086;
wire n_30087;
wire n_30088;
wire n_30089;
wire n_30090;
wire n_30091;
wire n_30092;
wire n_30093;
wire n_30094;
wire n_30095;
wire n_30096;
wire n_30097;
wire n_30098;
wire n_30099;
wire n_30100;
wire n_30101;
wire n_30102;
wire n_30103;
wire n_30104;
wire n_30105;
wire n_30106;
wire n_30107;
wire n_30108;
wire n_30109;
wire n_30110;
wire n_30111;
wire n_30112;
wire n_30113;
wire n_30114;
wire n_30115;
wire n_30116;
wire n_30117;
wire n_30118;
wire n_30119;
wire n_30120;
wire n_30121;
wire n_30122;
wire n_30123;
wire n_30124;
wire n_30125;
wire n_30126;
wire n_30127;
wire n_30128;
wire n_30129;
wire n_30130;
wire n_30131;
wire n_30132;
wire n_30133;
wire n_30134;
wire n_30135;
wire n_30136;
wire n_30137;
wire n_30138;
wire n_30139;
wire n_30140;
wire n_30141;
wire n_30142;
wire n_30143;
wire n_30144;
wire n_30145;
wire n_30146;
wire n_30147;
wire n_30148;
wire n_30149;
wire n_30150;
wire n_30151;
wire n_30152;
wire n_30153;
wire n_30154;
wire n_30155;
wire n_30156;
wire n_30157;
wire n_30158;
wire n_30159;
wire n_30160;
wire n_30161;
wire n_30162;
wire n_30163;
wire n_30164;
wire n_30165;
wire n_30166;
wire n_30167;
wire n_30168;
wire n_30169;
wire n_30170;
wire n_30171;
wire n_30172;
wire n_30173;
wire n_30174;
wire n_30175;
wire n_30176;
wire n_30177;
wire n_30178;
wire n_30179;
wire n_30180;
wire n_30181;
wire n_30182;
wire n_30183;
wire n_30184;
wire n_30185;
wire n_30186;
wire n_30187;
wire n_30188;
wire n_30189;
wire n_30190;
wire n_30191;
wire n_30192;
wire n_30193;
wire n_30194;
wire n_30195;
wire n_30196;
wire n_30197;
wire n_30198;
wire n_30199;
wire n_30200;
wire n_30201;
wire n_30202;
wire n_30203;
wire n_30204;
wire n_30205;
wire n_30206;
wire n_30207;
wire n_30208;
wire n_30209;
wire n_30210;
wire n_30211;
wire n_30212;
wire n_30213;
wire n_30214;
wire n_30215;
wire n_30216;
wire n_30217;
wire n_30218;
wire n_30219;
wire n_30220;
wire n_30221;
wire n_30222;
wire n_30223;
wire n_30224;
wire n_30225;
wire n_30226;
wire n_30227;
wire n_30228;
wire n_30229;
wire n_30230;
wire n_30231;
wire n_30232;
wire n_30233;
wire n_30234;
wire n_30235;
wire n_30236;
wire n_30237;
wire n_30238;
wire n_30239;
wire n_30240;
wire n_30241;
wire n_30242;
wire n_30243;
wire n_30244;
wire n_30245;
wire n_30246;
wire n_30247;
wire n_30248;
wire n_30249;
wire n_30250;
wire n_30251;
wire n_30252;
wire n_30253;
wire n_30254;
wire n_30255;
wire n_30256;
wire n_30257;
wire n_30258;
wire n_30259;
wire n_30260;
wire n_30261;
wire n_30262;
wire n_30263;
wire n_30264;
wire n_30265;
wire n_30266;
wire n_30267;
wire n_30268;
wire n_30269;
wire n_30270;
wire n_30271;
wire n_30272;
wire n_30273;
wire n_30274;
wire n_30275;
wire n_30276;
wire n_30277;
wire n_30278;
wire n_30279;
wire n_30280;
wire n_30281;
wire n_30282;
wire n_30283;
wire n_30284;
wire n_30285;
wire n_30286;
wire n_30287;
wire n_30288;
wire n_30289;
wire n_30290;
wire n_30291;
wire n_30292;
wire n_30293;
wire n_30294;
wire n_30295;
wire n_30296;
wire n_30297;
wire n_30298;
wire n_30299;
wire n_30300;
wire n_30301;
wire n_30302;
wire n_30303;
wire n_30304;
wire n_30305;
wire n_30306;
wire n_30307;
wire n_30308;
wire n_30309;
wire n_30310;
wire n_30311;
wire n_30312;
wire n_30313;
wire n_30314;
wire n_30315;
wire n_30316;
wire n_30317;
wire n_30318;
wire n_30319;
wire n_30320;
wire n_30321;
wire n_30322;
wire n_30323;
wire n_30324;
wire n_30325;
wire n_30326;
wire n_30327;
wire n_30328;
wire n_30329;
wire n_30330;
wire n_30331;
wire n_30332;
wire n_30333;
wire n_30334;
wire n_30335;
wire n_30336;
wire n_30337;
wire n_30338;
wire n_30339;
wire n_30340;
wire n_30341;
wire n_30342;
wire n_30343;
wire n_30344;
wire n_30345;
wire n_30346;
wire n_30347;
wire n_30348;
wire n_30349;
wire n_30350;
wire n_30351;
wire n_30352;
wire n_30353;
wire n_30354;
wire n_30355;
wire n_30356;
wire n_30357;
wire n_30358;
wire n_30359;
wire n_30360;
wire n_30361;
wire n_30362;
wire n_30363;
wire n_30364;
wire n_30365;
wire n_30366;
wire n_30367;
wire n_30368;
wire n_30369;
wire n_30370;
wire n_30371;
wire n_30372;
wire n_30373;
wire n_30374;
wire n_30375;
wire n_30376;
wire n_30377;
wire n_30378;
wire n_30379;
wire n_30380;
wire n_30381;
wire n_30382;
wire n_30383;
wire n_30384;
wire n_30385;
wire n_30386;
wire n_30387;
wire n_30388;
wire n_30389;
wire n_30390;
wire n_30391;
wire n_30392;
wire n_30393;
wire n_30394;
wire n_30395;
wire n_30396;
wire n_30397;
wire n_30398;
wire n_30399;
wire n_30400;
wire n_30401;
wire n_30402;
wire n_30403;
wire n_30404;
wire n_30405;
wire n_30406;
wire n_30407;
wire n_30408;
wire n_30409;
wire n_30410;
wire n_30411;
wire n_30412;
wire n_30413;
wire n_30414;
wire n_30415;
wire n_30416;
wire n_30417;
wire n_30418;
wire n_30419;
wire n_30420;
wire n_30421;
wire n_30422;
wire n_30423;
wire n_30424;
wire n_30425;
wire n_30426;
wire n_30427;
wire n_30428;
wire n_30429;
wire n_30430;
wire n_30431;
wire n_30432;
wire n_30433;
wire n_30434;
wire n_30435;
wire n_30436;
wire n_30437;
wire n_30438;
wire n_30439;
wire n_30440;
wire n_30441;
wire n_30442;
wire n_30443;
wire n_30444;
wire n_30445;
wire n_30446;
wire n_30447;
wire n_30448;
wire n_30449;
wire n_30450;
wire n_30451;
wire n_30452;
wire n_30453;
wire n_30454;
wire n_30455;
wire n_30456;
wire n_30457;
wire n_30458;
wire n_30459;
wire n_30460;
wire n_30461;
wire n_30462;
wire n_30463;
wire n_30464;
wire n_30465;
wire n_30466;
wire n_30467;
wire n_30468;
wire n_30469;
wire n_30470;
wire n_30471;
wire n_30472;
wire n_30473;
wire n_30474;
wire n_30475;
wire n_30476;
wire n_30477;
wire n_30478;
wire n_30479;
wire n_30480;
wire n_30481;
wire n_30482;
wire n_30483;
wire n_30484;
wire n_30485;
wire n_30486;
wire n_30487;
wire n_30488;
wire n_30489;
wire n_30490;
wire n_30491;
wire n_30492;
wire n_30493;
wire n_30494;
wire n_30495;
wire n_30496;
wire n_30497;
wire n_30498;
wire n_30499;
wire n_30500;
wire n_30501;
wire n_30502;
wire n_30503;
wire n_30504;
wire n_30505;
wire n_30506;
wire n_30507;
wire n_30508;
wire n_30509;
wire n_30510;
wire n_30511;
wire n_30512;
wire n_30513;
wire n_30514;
wire n_30515;
wire n_30516;
wire n_30517;
wire n_30518;
wire n_30519;
wire n_30520;
wire n_30521;
wire n_30522;
wire n_30523;
wire n_30524;
wire n_30525;
wire n_30526;
wire n_30527;
wire n_30528;
wire n_30529;
wire n_30530;
wire n_30531;
wire n_30532;
wire n_30533;
wire n_30534;
wire n_30535;
wire n_30536;
wire n_30537;
wire n_30538;
wire n_30539;
wire n_30540;
wire n_30541;
wire n_30542;
wire n_30543;
wire n_30544;
wire n_30545;
wire n_30546;
wire n_30547;
wire n_30548;
wire n_30549;
wire n_30550;
wire n_30551;
wire n_30552;
wire n_30553;
wire n_30554;
wire n_30555;
wire n_30556;
wire n_30557;
wire n_30558;
wire n_30559;
wire n_30560;
wire n_30561;
wire n_30562;
wire n_30563;
wire n_30564;
wire n_30565;
wire n_30566;
wire n_30567;
wire n_30568;
wire n_30569;
wire n_30570;
wire n_30571;
wire n_30572;
wire n_30573;
wire n_30574;
wire n_30575;
wire n_30576;
wire n_30577;
wire n_30578;
wire n_30579;
wire n_30580;
wire n_30581;
wire n_30582;
wire n_30583;
wire n_30584;
wire n_30585;
wire n_30586;
wire n_30587;
wire n_30588;
wire n_30589;
wire n_30590;
wire n_30591;
wire n_30592;
wire n_30593;
wire n_30594;
wire n_30595;
wire n_30596;
wire n_30597;
wire n_30598;
wire n_30599;
wire n_30600;
wire n_30601;
wire n_30602;
wire n_30603;
wire n_30604;
wire n_30605;
wire n_30606;
wire n_30607;
wire n_30608;
wire n_30609;
wire n_30610;
wire n_30611;
wire n_30612;
wire n_30613;
wire n_30614;
wire n_30615;
wire n_30616;
wire n_30617;
wire n_30618;
wire n_30619;
wire n_30620;
wire n_30621;
wire n_30622;
wire n_30623;
wire n_30624;
wire n_30625;
wire n_30626;
wire n_30627;
wire n_30628;
wire n_30629;
wire n_30630;
wire n_30631;
wire n_30632;
wire n_30633;
wire n_30634;
wire n_30635;
wire n_30636;
wire n_30637;
wire n_30638;
wire n_30639;
wire n_30640;
wire n_30641;
wire n_30642;
wire n_30643;
wire n_30644;
wire n_30645;
wire n_30646;
wire n_30647;
wire n_30648;
wire n_30649;
wire n_30650;
wire n_30651;
wire n_30652;
wire n_30653;
wire n_30654;
wire n_30655;
wire n_30656;
wire n_30657;
wire n_30658;
wire n_30659;
wire n_30660;
wire n_30661;
wire n_30662;
wire n_30663;
wire n_30664;
wire n_30665;
wire n_30666;
wire n_30667;
wire n_30668;
wire n_30669;
wire n_30670;
wire n_30671;
wire n_30672;
wire n_30673;
wire n_30674;
wire n_30675;
wire n_30676;
wire n_30677;
wire n_30678;
wire n_30679;
wire n_30680;
wire n_30681;
wire n_30682;
wire n_30683;
wire n_30684;
wire n_30685;
wire n_30686;
wire n_30687;
wire n_30688;
wire n_30689;
wire n_30690;
wire n_30691;
wire n_30692;
wire n_30693;
wire n_30694;
wire n_30695;
wire n_30696;
wire n_30697;
wire n_30698;
wire n_30699;
wire n_30700;
wire n_30701;
wire n_30702;
wire n_30703;
wire n_30704;
wire n_30705;
wire n_30706;
wire n_30707;
wire n_30708;
wire n_30709;
wire n_30710;
wire n_30711;
wire n_30712;
wire n_30713;
wire n_30714;
wire n_30715;
wire n_30716;
wire n_30717;
wire n_30718;
wire n_30719;
wire n_30720;
wire n_30721;
wire n_30722;
wire n_30723;
wire n_30724;
wire n_30725;
wire n_30726;
wire n_30727;
wire n_30728;
wire n_30729;
wire n_30730;
wire n_30731;
wire n_30732;
wire n_30733;
wire n_30734;
wire n_30735;
wire n_30736;
wire n_30737;
wire n_30738;
wire n_30739;
wire n_30740;
wire n_30741;
wire n_30742;
wire n_30743;
wire n_30744;
wire n_30745;
wire n_30746;
wire n_30747;
wire n_30748;
wire n_30749;
wire n_30750;
wire n_30751;
wire n_30752;
wire n_30753;
wire n_30754;
wire n_30755;
wire n_30756;
wire n_30757;
wire n_30758;
wire n_30759;
wire n_30760;
wire n_30761;
wire n_30762;
wire n_30763;
wire n_30764;
wire n_30765;
wire n_30766;
wire n_30767;
wire n_30768;
wire n_30769;
wire n_30770;
wire n_30771;
wire n_30772;
wire n_30773;
wire n_30774;
wire n_30775;
wire n_30776;
wire n_30777;
wire n_30778;
wire n_30779;
wire n_30780;
wire n_30781;
wire n_30782;
wire n_30783;
wire n_30784;
wire n_30785;
wire n_30786;
wire n_30787;
wire n_30788;
wire n_30789;
wire n_30790;
wire n_30791;
wire n_30792;
wire n_30793;
wire n_30794;
wire n_30795;
wire n_30796;
wire n_30797;
wire n_30798;
wire n_30799;
wire n_30800;
wire n_30801;
wire n_30802;
wire n_30803;
wire n_30804;
wire n_30805;
wire n_30806;
wire n_30807;
wire n_30808;
wire n_30809;
wire n_30810;
wire n_30811;
wire n_30812;
wire n_30813;
wire n_30814;
wire n_30815;
wire n_30816;
wire n_30817;
wire n_30818;
wire n_30819;
wire n_30820;
wire n_30821;
wire n_30822;
wire n_30823;
wire n_30824;
wire n_30825;
wire n_30826;
wire n_30827;
wire n_30828;
wire n_30829;
wire n_30830;
wire n_30831;
wire n_30832;
wire n_30833;
wire n_30834;
wire n_30835;
wire n_30836;
wire n_30837;
wire n_30838;
wire n_30839;
wire n_30840;
wire n_30841;
wire n_30842;
wire n_30843;
wire n_30844;
wire n_30845;
wire n_30846;
wire n_30847;
wire n_30848;
wire n_30849;
wire n_30850;
wire n_30851;
wire n_30852;
wire n_30853;
wire n_30854;
wire n_30855;
wire n_30856;
wire n_30857;
wire n_30858;
wire n_30859;
wire n_30860;
wire n_30861;
wire n_30862;
wire n_30863;
wire n_30864;
wire n_30865;
wire n_30866;
wire n_30867;
wire n_30868;
wire n_30869;
wire n_30870;
wire n_30871;
wire n_30872;
wire n_30873;
wire n_30874;
wire n_30875;
wire n_30876;
wire n_30877;
wire n_30878;
wire n_30879;
wire n_30880;
wire n_30881;
wire n_30882;
wire n_30883;
wire n_30884;
wire n_30885;
wire n_30886;
wire n_30887;
wire n_30888;
wire n_30889;
wire n_30890;
wire n_30891;
wire n_30892;
wire n_30893;
wire n_30894;
wire n_30895;
wire n_30896;
wire n_30897;
wire n_30898;
wire n_30899;
wire n_30900;
wire n_30901;
wire n_30902;
wire n_30903;
wire n_30904;
wire n_30905;
wire n_30906;
wire n_30907;
wire n_30908;
wire n_30909;
wire n_30910;
wire n_30911;
wire n_30912;
wire n_30913;
wire n_30914;
wire n_30915;
wire n_30916;
wire n_30917;
wire n_30918;
wire n_30919;
wire n_30920;
wire n_30921;
wire n_30922;
wire n_30923;
wire n_30924;
wire n_30925;
wire n_30926;
wire n_30927;
wire n_30928;
wire n_30929;
wire n_30930;
wire n_30931;
wire n_30932;
wire n_30933;
wire n_30934;
wire n_30935;
wire n_30936;
wire n_30937;
wire n_30938;
wire n_30939;
wire n_30940;
wire n_30941;
wire n_30942;
wire n_30943;
wire n_30944;
wire n_30945;
wire n_30946;
wire n_30947;
wire n_30948;
wire n_30949;
wire n_30950;
wire n_30951;
wire n_30952;
wire n_30953;
wire n_30954;
wire n_30955;
wire n_30956;
wire n_30957;
wire n_30958;
wire n_30959;
wire n_30960;
wire n_30961;
wire n_30962;
wire n_30963;
wire n_30964;
wire n_30965;
wire n_30966;
wire n_30967;
wire n_30968;
wire n_30969;
wire n_30970;
wire n_30971;
wire n_30972;
wire n_30973;
wire n_30974;
wire n_30975;
wire n_30976;
wire n_30977;
wire n_30978;
wire n_30979;
wire n_30980;
wire n_30981;
wire n_30982;
wire n_30983;
wire n_30984;
wire n_30985;
wire n_30986;
wire n_30987;
wire n_30988;
wire n_30989;
wire n_30990;
wire n_30991;
wire n_30992;
wire n_30993;
wire n_30994;
wire n_30995;
wire n_30996;
wire n_30997;
wire n_30998;
wire n_30999;
wire n_31000;
wire n_31001;
wire n_31002;
wire n_31003;
wire n_31004;
wire n_31005;
wire n_31006;
wire n_31007;
wire n_31008;
wire n_31009;
wire n_31010;
wire n_31011;
wire n_31012;
wire n_31013;
wire n_31014;
wire n_31015;
wire n_31016;
wire n_31017;
wire n_31018;
wire n_31019;
wire n_31020;
wire n_31021;
wire n_31022;
wire n_31023;
wire n_31024;
wire n_31025;
wire n_31026;
wire n_31027;
wire n_31028;
wire n_31029;
wire n_31030;
wire n_31031;
wire n_31032;
wire n_31033;
wire n_31034;
wire n_31035;
wire n_31036;
wire n_31037;
wire n_31038;
wire n_31039;
wire n_31040;
wire n_31041;
wire n_31042;
wire n_31043;
wire n_31044;
wire n_31045;
wire n_31046;
wire n_31047;
wire n_31048;
wire n_31049;
wire n_31050;
wire n_31051;
wire n_31052;
wire n_31053;
wire n_31054;
wire n_31055;
wire n_31056;
wire n_31057;
wire n_31058;
wire n_31059;
wire n_31060;
wire n_31061;
wire n_31062;
wire n_31063;
wire n_31064;
wire n_31065;
wire n_31066;
wire n_31067;
wire n_31068;
wire n_31069;
wire n_31070;
wire n_31071;
wire n_31072;
wire n_31073;
wire n_31074;
wire n_31075;
wire n_31076;
wire n_31077;
wire n_31078;
wire n_31079;
wire n_31080;
wire n_31081;
wire n_31082;
wire n_31083;
wire n_31084;
wire n_31085;
wire n_31086;
wire n_31087;
wire n_31088;
wire n_31089;
wire n_31090;
wire n_31091;
wire n_31092;
wire n_31093;
wire n_31094;
wire n_31095;
wire n_31096;
wire n_31097;
wire n_31098;
wire n_31099;
wire n_31100;
wire n_31101;
wire n_31102;
wire n_31103;
wire n_31104;
wire n_31105;
wire n_31106;
wire n_31107;
wire n_31108;
wire n_31109;
wire n_31110;
wire n_31111;
wire n_31112;
wire n_31113;
wire n_31114;
wire n_31115;
wire n_31116;
wire n_31117;
wire n_31118;
wire n_31119;
wire n_31120;
wire n_31121;
wire n_31122;
wire n_31123;
wire n_31124;
wire n_31125;
wire n_31126;
wire n_31127;
wire n_31128;
wire n_31129;
wire n_31130;
wire n_31131;
wire n_31132;
wire n_31133;
wire n_31134;
wire n_31135;
wire n_31136;
wire n_31137;
wire n_31138;
wire n_31139;
wire n_31140;
wire n_31141;
wire n_31142;
wire n_31143;
wire n_31144;
wire n_31145;
wire n_31146;
wire n_31147;
wire n_31148;
wire n_31149;
wire n_31150;
wire n_31151;
wire n_31152;
wire n_31153;
wire n_31154;
wire n_31155;
wire n_31156;
wire n_31157;
wire n_31158;
wire n_31159;
wire n_31160;
wire n_31161;
wire n_31162;
wire n_31163;
wire n_31164;
wire n_31165;
wire n_31166;
wire n_31167;
wire n_31168;
wire n_31169;
wire n_31170;
wire n_31171;
wire n_31172;
wire n_31173;
wire n_31174;
wire n_31175;
wire n_31176;
wire n_31177;
wire n_31178;
wire n_31179;
wire n_31180;
wire n_31181;
wire n_31182;
wire n_31183;
wire n_31184;
wire n_31185;
wire n_31186;
wire n_31187;
wire n_31188;
wire n_31189;
wire n_31190;
wire n_31191;
wire n_31192;
wire n_31193;
wire n_31194;
wire n_31195;
wire n_31196;
wire n_31197;
wire n_31198;
wire n_31199;
wire n_31200;
wire n_31201;
wire n_31202;
wire n_31203;
wire n_31204;
wire n_31205;
wire n_31206;
wire n_31207;
wire n_31208;
wire n_31209;
wire n_31210;
wire n_31211;
wire n_31212;
wire n_31213;
wire n_31214;
wire n_31215;
wire n_31216;
wire n_31217;
wire n_31218;
wire n_31219;
wire n_31220;
wire n_31221;
wire n_31222;
wire n_31223;
wire n_31224;
wire n_31225;
wire n_31226;
wire n_31227;
wire n_31228;
wire n_31229;
wire n_31230;
wire n_31231;
wire n_31232;
wire n_31233;
wire n_31234;
wire n_31235;
wire n_31236;
wire n_31237;
wire n_31238;
wire n_31239;
wire n_31240;
wire n_31241;
wire n_31242;
wire n_31243;
wire n_31244;
wire n_31245;
wire n_31246;
wire n_31247;
wire n_31248;
wire n_31249;
wire n_31250;
wire n_31251;
wire n_31252;
wire n_31253;
wire n_31254;
wire n_31255;
wire n_31256;
wire n_31257;
wire n_31258;
wire n_31259;
wire n_31260;
wire n_31261;
wire n_31262;
wire n_31263;
wire n_31264;
wire n_31265;
wire n_31266;
wire n_31267;
wire n_31268;
wire n_31269;
wire n_31270;
wire n_31271;
wire n_31272;
wire n_31273;
wire n_31274;
wire n_31275;
wire n_31276;
wire n_31277;
wire n_31278;
wire n_31279;
wire n_31280;
wire n_31281;
wire n_31282;
wire n_31283;
wire n_31284;
wire n_31285;
wire n_31286;
wire n_31287;
wire n_31288;
wire n_31289;
wire n_31290;
wire n_31291;
wire n_31292;
wire n_31293;
wire n_31294;
wire n_31295;
wire n_31296;
wire n_31297;
wire n_31298;
wire n_31299;
wire n_31300;
wire n_31301;
wire n_31302;
wire n_31303;
wire n_31304;
wire n_31305;
wire n_31306;
wire n_31307;
wire n_31308;
wire n_31309;
wire n_31310;
wire n_31311;
wire n_31312;
wire n_31313;
wire n_31314;
wire n_31315;
wire n_31316;
wire n_31317;
wire n_31318;
wire n_31319;
wire n_31320;
wire n_31321;
wire n_31322;
wire n_31323;
wire n_31324;
wire n_31325;
wire n_31326;
wire n_31327;
wire n_31328;
wire n_31329;
wire n_31330;
wire n_31331;
wire n_31332;
wire n_31333;
wire n_31334;
wire n_31335;
wire n_31336;
wire n_31337;
wire n_31338;
wire n_31339;
wire n_31340;
wire n_31341;
wire n_31342;
wire n_31343;
wire n_31344;
wire n_31345;
wire n_31346;
wire n_31347;
wire n_31348;
wire n_31349;
wire n_31350;
wire n_31351;
wire n_31352;
wire n_31353;
wire n_31354;
wire n_31355;
wire n_31356;
wire n_31357;
wire n_31358;
wire n_31359;
wire n_31360;
wire n_31361;
wire n_31362;
wire n_31363;
wire n_31364;
wire n_31365;
wire n_31366;
wire n_31367;
wire n_31368;
wire n_31369;
wire n_31370;
wire n_31371;
wire n_31372;
wire n_31373;
wire n_31374;
wire n_31375;
wire n_31376;
wire n_31377;
wire n_31378;
wire n_31379;
wire n_31380;
wire n_31381;
wire n_31382;
wire n_31383;
wire n_31384;
wire n_31385;
wire n_31386;
wire n_31387;
wire n_31388;
wire n_31389;
wire n_31390;
wire n_31391;
wire n_31392;
wire n_31393;
wire n_31394;
wire n_31395;
wire n_31396;
wire n_31397;
wire n_31398;
wire n_31399;
wire n_31400;
wire n_31401;
wire n_31402;
wire n_31403;
wire n_31404;
wire n_31405;
wire n_31406;
wire n_31407;
wire n_31408;
wire n_31409;
wire n_31410;
wire n_31411;
wire n_31412;
wire n_31413;
wire n_31414;
wire n_31415;
wire n_31416;
wire n_31417;
wire n_31418;
wire n_31419;
wire n_31420;
wire n_31421;
wire n_31422;
wire n_31423;
wire n_31424;
wire n_31425;
wire n_31426;
wire n_31427;
wire n_31428;
wire n_31429;
wire n_31430;
wire n_31431;
wire n_31432;
wire n_31433;
wire n_31434;
wire n_31435;
wire n_31436;
wire n_31437;
wire n_31438;
wire n_31439;
wire n_31440;
wire n_31441;
wire n_31442;
wire n_31443;
wire n_31444;
wire n_31445;
wire n_31446;
wire n_31447;
wire n_31448;
wire n_31449;
wire n_31450;
wire n_31451;
wire n_31452;
wire n_31453;
wire n_31454;
wire n_31455;
wire n_31456;
wire n_31457;
wire n_31458;
wire n_31459;
wire n_31460;
wire n_31461;
wire n_31462;
wire n_31463;
wire n_31464;
wire n_31465;
wire n_31466;
wire n_31467;
wire n_31468;
wire n_31469;
wire n_31470;
wire n_31471;
wire n_31472;
wire n_31473;
wire n_31474;
wire n_31475;
wire n_31476;
wire n_31477;
wire n_31478;
wire n_31479;
wire n_31480;
wire n_31481;
wire n_31482;
wire n_31483;
wire n_31484;
wire n_31485;
wire n_31486;
wire n_31487;
wire n_31488;
wire n_31489;
wire n_31490;
wire n_31491;
wire n_31492;
wire n_31493;
wire n_31494;
wire n_31495;
wire n_31496;
wire n_31497;
wire n_31498;
wire n_31499;
wire n_31500;
wire n_31501;
wire n_31502;
wire n_31503;
wire n_31504;
wire n_31505;
wire n_31506;
wire n_31507;
wire n_31508;
wire n_31509;
wire n_31510;
wire n_31511;
wire n_31512;
wire n_31513;
wire n_31514;
wire n_31515;
wire n_31516;
wire n_31517;
wire n_31518;
wire n_31519;
wire n_31520;
wire n_31521;
wire n_31522;
wire n_31523;
wire n_31524;
wire n_31525;
wire n_31526;
wire n_31527;
wire n_31528;
wire n_31529;
wire n_31530;
wire n_31531;
wire n_31532;
wire n_31533;
wire n_31534;
wire n_31535;
wire n_31536;
wire n_31537;
wire n_31538;
wire n_31539;
wire n_31540;
wire n_31541;
wire n_31542;
wire n_31543;
wire n_31544;
wire n_31545;
wire n_31546;
wire n_31547;
wire n_31548;
wire n_31549;
wire n_31550;
wire n_31551;
wire n_31552;
wire n_31553;
wire n_31554;
wire n_31555;
wire n_31556;
wire n_31557;
wire n_31558;
wire n_31559;
wire n_31560;
wire n_31561;
wire n_31562;
wire n_31563;
wire n_31564;
wire n_31565;
wire n_31566;
wire n_31567;
wire n_31568;
wire n_31569;
wire n_31570;
wire n_31571;
wire n_31572;
wire n_31573;
wire n_31574;
wire n_31575;
wire n_31576;
wire n_31577;
wire n_31578;
wire n_31579;
wire n_31580;
wire n_31581;
wire n_31582;
wire n_31583;
wire n_31584;
wire n_31585;
wire n_31586;
wire n_31587;
wire n_31588;
wire n_31589;
wire n_31590;
wire n_31591;
wire n_31592;
wire n_31593;
wire n_31594;
wire n_31595;
wire n_31596;
wire n_31597;
wire n_31598;
wire n_31599;
wire n_31600;
wire n_31601;
wire n_31602;
wire n_31603;
wire n_31604;
wire n_31605;
wire n_31606;
wire n_31607;
wire n_31608;
wire n_31609;
wire n_31610;
wire n_31611;
wire n_31612;
wire n_31613;
wire n_31614;
wire n_31615;
wire n_31616;
wire n_31617;
wire n_31618;
wire n_31619;
wire n_31620;
wire n_31621;
wire n_31622;
wire n_31623;
wire n_31624;
wire n_31625;
wire n_31626;
wire n_31627;
wire n_31628;
wire n_31629;
wire n_31630;
wire n_31631;
wire n_31632;
wire n_31633;
wire n_31634;
wire n_31635;
wire n_31636;
wire n_31637;
wire n_31638;
wire n_31639;
wire n_31640;
wire n_31641;
wire n_31642;
wire n_31643;
wire n_31644;
wire n_31645;
wire n_31646;
wire n_31647;
wire n_31648;
wire n_31649;
wire n_31650;
wire n_31651;
wire n_31652;
wire n_31653;
wire n_31654;
wire n_31655;
wire n_31656;
wire n_31657;
wire n_31658;
wire n_31659;
wire n_31660;
wire n_31661;
wire n_31662;
wire n_31663;
wire n_31664;
wire n_31665;
wire n_31666;
wire n_31667;
wire n_31668;
wire n_31669;
wire n_31670;
wire n_31671;
wire n_31672;
wire n_31673;
wire n_31674;
wire n_31675;
wire n_31676;
wire n_31677;
wire n_31678;
wire n_31679;
wire n_31680;
wire n_31681;
wire n_31682;
wire n_31683;
wire n_31684;
wire n_31685;
wire n_31686;
wire n_31687;
wire n_31688;
wire n_31689;
wire n_31690;
wire n_31691;
wire n_31692;
wire n_31693;
wire n_31694;
wire n_31695;
wire n_31696;
wire n_31697;
wire n_31698;
wire n_31699;
wire n_31700;
wire n_31701;
wire n_31702;
wire n_31703;
wire n_31704;
wire n_31705;
wire n_31706;
wire n_31707;
wire n_31708;
wire n_31709;
wire n_31710;
wire n_31711;
wire n_31712;
wire n_31713;
wire n_31714;
wire n_31715;
wire n_31716;
wire n_31717;
wire n_31718;
wire n_31719;
wire n_31720;
wire n_31721;
wire n_31722;
wire n_31723;
wire n_31724;
wire n_31725;
wire n_31726;
wire n_31727;
wire n_31728;
wire n_31729;
wire n_31730;
wire n_31731;
wire n_31732;
wire n_31733;
wire n_31734;
wire n_31735;
wire n_31736;
wire n_31737;
wire n_31738;
wire n_31739;
wire n_31740;
wire n_31741;
wire n_31742;
wire n_31743;
wire n_31744;
wire n_31745;
wire n_31746;
wire n_31747;
wire n_31748;
wire n_31749;
wire n_31750;
wire n_31751;
wire n_31752;
wire n_31753;
wire n_31754;
wire n_31755;
wire n_31756;
wire n_31757;
wire n_31758;
wire n_31759;
wire n_31760;
wire n_31761;
wire n_31762;
wire n_31763;
wire n_31764;
wire n_31765;
wire n_31766;
wire n_31767;
wire n_31768;
wire n_31769;
wire n_31770;
wire n_31771;
wire n_31772;
wire n_31773;
wire n_31774;
wire n_31775;
wire n_31776;
wire n_31777;
wire n_31778;
wire n_31779;
wire n_31780;
wire n_31781;
wire n_31782;
wire n_31783;
wire n_31784;
wire n_31785;
wire n_31786;
wire n_31787;
wire n_31788;
wire n_31789;
wire n_31790;
wire n_31791;
wire n_31792;
wire n_31793;
wire n_31794;
wire n_31795;
wire n_31796;
wire n_31797;
wire n_31798;
wire n_31799;
wire n_31800;
wire n_31801;
wire n_31802;
wire n_31803;
wire n_31804;
wire n_31805;
wire n_31806;
wire n_31807;
wire n_31808;
wire n_31809;
wire n_31810;
wire n_31811;
wire n_31812;
wire n_31813;
wire n_31814;
wire n_31815;
wire n_31816;
wire n_31817;
wire n_31818;
wire n_31819;
wire n_31820;
wire n_31821;
wire n_31822;
wire n_31823;
wire n_31824;
wire n_31825;
wire n_31826;
wire n_31827;
wire n_31828;
wire n_31829;
wire n_31830;
wire n_31831;
wire n_31832;
wire n_31833;
wire n_31834;
wire n_31835;
wire n_31836;
wire n_31837;
wire n_31838;
wire n_31839;
wire n_31840;
wire n_31841;
wire n_31842;
wire n_31843;
wire n_31844;
wire n_31845;
wire n_31846;
wire n_31847;
wire n_31848;
wire n_31849;
wire n_31850;
wire n_31851;
wire n_31852;
wire n_31853;
wire n_31854;
wire n_31855;
wire n_31856;
wire n_31857;
wire n_31858;
wire n_31859;
wire n_31860;
wire n_31861;
wire n_31862;
wire n_31863;
wire n_31864;
wire n_31865;
wire n_31866;
wire n_31867;
wire n_31868;
wire n_31869;
wire n_31870;
wire n_31871;
wire n_31872;
wire n_31873;
wire n_31874;
wire n_31875;
wire n_31876;
wire n_31877;
wire n_31878;
wire n_31879;
wire n_31880;
wire n_31881;
wire n_31882;
wire n_31883;
wire n_31884;
wire n_31885;
wire n_31886;
wire n_31887;
wire n_31888;
wire n_31889;
wire n_31890;
wire n_31891;
wire n_31892;
wire n_31893;
wire n_31894;
wire n_31895;
wire n_31896;
wire n_31897;
wire n_31898;
wire n_31899;
wire n_31900;
wire n_31901;
wire n_31902;
wire n_31903;
wire n_31904;
wire n_31905;
wire n_31906;
wire n_31907;
wire n_31908;
wire n_31909;
wire n_31910;
wire n_31911;
wire n_31912;
wire n_31913;
wire n_31914;
wire n_31915;
wire n_31916;
wire n_31917;
wire n_31918;
wire n_31919;
wire n_31920;
wire n_31921;
wire n_31922;
wire n_31923;
wire n_31924;
wire n_31925;
wire n_31926;
wire n_31927;
wire n_31928;
wire n_31929;
wire n_31930;
wire n_31931;
wire n_31932;
wire n_31933;
wire n_31934;
wire n_31935;
wire n_31936;
wire n_31937;
wire n_31938;
wire n_31939;
wire n_31940;
wire n_31941;
wire n_31942;
wire n_31943;
wire n_31944;
wire n_31945;
wire n_31946;
wire n_31947;
wire n_31948;
wire n_31949;
wire n_31950;
wire n_31951;
wire n_31952;
wire n_31953;
wire n_31954;
wire n_31955;
wire n_31956;
wire n_31957;
wire n_31958;
wire n_31959;
wire n_31960;
wire n_31961;
wire n_31962;
wire n_31963;
wire n_31964;
wire n_31965;
wire n_31966;
wire n_31967;
wire n_31968;
wire n_31969;
wire n_31970;
wire n_31971;
wire n_31972;
wire n_31973;
wire n_31974;
wire n_31975;
wire n_31976;
wire n_31977;
wire n_31978;
wire n_31979;
wire n_31980;
wire n_31981;
wire n_31982;
wire n_31983;
wire n_31984;
wire n_31985;
wire n_31986;
wire n_31987;
wire n_31988;
wire n_31989;
wire n_31990;
wire n_31991;
wire n_31992;
wire n_31993;
wire n_31994;
wire n_31995;
wire n_31996;
wire n_31997;
wire n_31998;
wire n_31999;
wire n_32000;
wire n_32001;
wire n_32002;
wire n_32003;
wire n_32004;
wire n_32005;
wire n_32006;
wire n_32007;
wire n_32008;
wire n_32009;
wire n_32010;
wire n_32011;
wire n_32012;
wire n_32013;
wire n_32014;
wire n_32015;
wire n_32016;
wire n_32017;
wire n_32018;
wire n_32019;
wire n_32020;
wire n_32021;
wire n_32022;
wire n_32023;
wire n_32024;
wire n_32025;
wire n_32026;
wire n_32027;
wire n_32028;
wire n_32029;
wire n_32030;
wire n_32031;
wire n_32032;
wire n_32033;
wire n_32034;
wire n_32035;
wire n_32036;
wire n_32037;
wire n_32038;
wire n_32039;
wire n_32040;
wire n_32041;
wire n_32042;
wire n_32043;
wire n_32044;
wire n_32045;
wire n_32046;
wire n_32047;
wire n_32048;
wire n_32049;
wire n_32050;
wire n_32051;
wire n_32052;
wire n_32053;
wire n_32054;
wire n_32055;
wire n_32056;
wire n_32057;
wire n_32058;
wire n_32059;
wire n_32060;
wire n_32061;
wire n_32062;
wire n_32063;
wire n_32064;
wire n_32065;
wire n_32066;
wire n_32067;
wire n_32068;
wire n_32069;
wire n_32070;
wire n_32071;
wire n_32072;
wire n_32073;
wire n_32074;
wire n_32075;
wire n_32076;
wire n_32077;
wire n_32078;
wire n_32079;
wire n_32080;
wire n_32081;
wire n_32082;
wire n_32083;
wire n_32084;
wire n_32085;
wire n_32086;
wire n_32087;
wire n_32088;
wire n_32089;
wire n_32090;
wire n_32091;
wire n_32092;
wire n_32093;
wire n_32094;
wire n_32095;
wire n_32096;
wire n_32097;
wire n_32098;
wire n_32099;
wire n_32100;
wire n_32101;
wire n_32102;
wire n_32103;
wire n_32104;
wire n_32105;
wire n_32106;
wire n_32107;
wire n_32108;
wire n_32109;
wire n_32110;
wire n_32111;
wire n_32112;
wire n_32113;
wire n_32114;
wire n_32115;
wire n_32116;
wire n_32117;
wire n_32118;
wire n_32119;
wire n_32120;
wire n_32121;
wire n_32122;
wire n_32123;
wire n_32124;
wire n_32125;
wire n_32126;
wire n_32127;
wire n_32128;
wire n_32129;
wire n_32130;
wire n_32131;
wire n_32132;
wire n_32133;
wire n_32134;
wire n_32135;
wire n_32136;
wire n_32137;
wire n_32138;
wire n_32139;
wire n_32140;
wire n_32141;
wire n_32142;
wire n_32143;
wire n_32144;
wire n_32145;
wire n_32146;
wire n_32147;
wire n_32148;
wire n_32149;
wire n_32150;
wire n_32151;
wire n_32152;
wire n_32153;
wire n_32154;
wire n_32155;
wire n_32156;
wire n_32157;
wire n_32158;
wire n_32159;
wire n_32160;
wire n_32161;
wire n_32162;
wire n_32163;
wire n_32164;
wire n_32165;
wire n_32166;
wire n_32167;
wire n_32168;
wire n_32169;
wire n_32170;
wire n_32171;
wire n_32172;
wire n_32173;
wire n_32174;
wire n_32175;
wire n_32176;
wire n_32177;
wire n_32178;
wire n_32179;
wire n_32180;
wire n_32181;
wire n_32182;
wire n_32183;
wire n_32184;
wire n_32185;
wire n_32186;
wire n_32187;
wire n_32188;
wire n_32189;
wire n_32190;
wire n_32191;
wire n_32192;
wire n_32193;
wire n_32194;
wire n_32195;
wire n_32196;
wire n_32197;
wire n_32198;
wire n_32199;
wire n_32200;
wire n_32201;
wire n_32202;
wire n_32203;
wire n_32204;
wire n_32205;
wire n_32206;
wire n_32207;
wire n_32208;
wire n_32209;
wire n_32210;
wire n_32211;
wire n_32212;
wire n_32213;
wire n_32214;
wire n_32215;
wire n_32216;
wire n_32217;
wire n_32218;
wire n_32219;
wire n_32220;
wire n_32221;
wire n_32222;
wire n_32223;
wire n_32224;
wire n_32225;
wire n_32226;
wire n_32227;
wire n_32228;
wire n_32229;
wire n_32230;
wire n_32231;
wire n_32232;
wire n_32233;
wire n_32234;
wire n_32235;
wire n_32236;
wire n_32237;
wire n_32238;
wire n_32239;
wire n_32240;
wire n_32241;
wire n_32242;
wire n_32243;
wire n_32244;
wire n_32245;
wire n_32246;
wire n_32247;
wire n_32248;
wire n_32249;
wire n_32250;
wire n_32251;
wire n_32252;
wire n_32253;
wire n_32254;
wire n_32255;
wire n_32256;
wire n_32257;
wire n_32258;
wire n_32259;
wire n_32260;
wire n_32261;
wire n_32262;
wire n_32263;
wire n_32264;
wire n_32265;
wire n_32266;
wire n_32267;
wire n_32268;
wire n_32269;
wire n_32270;
wire n_32271;
wire n_32272;
wire n_32273;
wire n_32274;
wire n_32275;
wire n_32276;
wire n_32277;
wire n_32278;
wire n_32279;
wire n_32280;
wire n_32281;
wire n_32282;
wire n_32283;
wire n_32284;
wire n_32285;
wire n_32286;
wire n_32287;
wire n_32288;
wire n_32289;
wire n_32290;
wire n_32291;
wire n_32292;
wire n_32293;
wire n_32294;
wire n_32295;
wire n_32296;
wire n_32297;
wire n_32298;
wire n_32299;
wire n_32300;
wire n_32301;
wire n_32302;
wire n_32303;
wire n_32304;
wire n_32305;
wire n_32306;
wire n_32307;
wire n_32308;
wire n_32309;
wire n_32310;
wire n_32311;
wire n_32312;
wire n_32313;
wire n_32314;
wire n_32315;
wire n_32316;
wire n_32317;
wire n_32318;
wire n_32319;
wire n_32320;
wire n_32321;
wire n_32322;
wire n_32323;
wire n_32324;
wire n_32325;
wire n_32326;
wire n_32327;
wire n_32328;
wire n_32329;
wire n_32330;
wire n_32331;
wire n_32332;
wire n_32333;
wire n_32334;
wire n_32335;
wire n_32336;
wire n_32337;
wire n_32338;
wire n_32339;
wire n_32340;
wire n_32341;
wire n_32342;
wire n_32343;
wire n_32344;
wire n_32345;
wire n_32346;
wire n_32347;
wire n_32348;
wire n_32349;
wire n_32350;
wire n_32351;
wire n_32352;
wire n_32353;
wire n_32354;
wire n_32355;
wire n_32356;
wire n_32357;
wire n_32358;
wire n_32359;
wire n_32360;
wire n_32361;
wire n_32362;
wire n_32363;
wire n_32364;
wire n_32365;
wire n_32366;
wire n_32367;
wire n_32368;
wire n_32369;
wire n_32370;
wire n_32371;
wire n_32372;
wire n_32373;
wire n_32374;
wire n_32375;
wire n_32376;
wire n_32377;
wire n_32378;
wire n_32379;
wire n_32380;
wire n_32381;
wire n_32382;
wire n_32383;
wire n_32384;
wire n_32385;
wire n_32386;
wire n_32387;
wire n_32388;
wire n_32389;
wire n_32390;
wire n_32391;
wire n_32392;
wire n_32393;
wire n_32394;
wire n_32395;
wire n_32396;
wire n_32397;
wire n_32398;
wire n_32399;
wire n_32400;
wire n_32401;
wire n_32402;
wire n_32403;
wire n_32404;
wire n_32405;
wire n_32406;
wire n_32407;
wire n_32408;
wire n_32409;
wire n_32410;
wire n_32411;
wire n_32412;
wire n_32413;
wire n_32414;
wire n_32415;
wire n_32416;
wire n_32417;
wire n_32418;
wire n_32419;
wire n_32420;
wire n_32421;
wire n_32422;
wire n_32423;
wire n_32424;
wire n_32425;
wire n_32426;
wire n_32427;
wire n_32428;
wire n_32429;
wire n_32430;
wire n_32431;
wire n_32432;
wire n_32433;
wire n_32434;
wire n_32435;
wire n_32436;
wire n_32437;
wire n_32438;
wire n_32439;
wire n_32440;
wire n_32441;
wire n_32442;
wire n_32443;
wire n_32444;
wire n_32445;
wire n_32446;
wire n_32447;
wire n_32448;
wire n_32449;
wire n_32450;
wire n_32451;
wire n_32452;
wire n_32453;
wire n_32454;
wire n_32455;
wire n_32456;
wire n_32457;
wire n_32458;
wire n_32459;
wire n_32460;
wire n_32461;
wire n_32462;
wire n_32463;
wire n_32464;
wire n_32465;
wire n_32466;
wire n_32467;
wire n_32468;
wire n_32469;
wire n_32470;
wire n_32471;
wire n_32472;
wire n_32473;
wire n_32474;
wire n_32475;
wire n_32476;
wire n_32477;
wire n_32478;
wire n_32479;
wire n_32480;
wire n_32481;
wire n_32482;
wire n_32483;
wire n_32484;
wire n_32485;
wire n_32486;
wire n_32487;
wire n_32488;
wire n_32489;
wire n_32490;
wire n_32491;
wire n_32492;
wire n_32493;
wire n_32494;
wire n_32495;
wire n_32496;
wire n_32497;
wire n_32498;
wire n_32499;
wire n_32500;
wire n_32501;
wire n_32502;
wire n_32503;
wire n_32504;
wire n_32505;
wire n_32506;
wire n_32507;
wire n_32508;
wire n_32509;
wire n_32510;
wire n_32511;
wire n_32512;
wire n_32513;
wire n_32514;
wire n_32515;
wire n_32516;
wire n_32517;
wire n_32518;
wire n_32519;
wire n_32520;
wire n_32521;
wire n_32522;
wire n_32523;
wire n_32524;
wire n_32525;
wire n_32526;
wire n_32527;
wire n_32528;
wire n_32529;
wire n_32530;
wire n_32531;
wire n_32532;
wire n_32533;
wire n_32534;
wire n_32535;
wire n_32536;
wire n_32537;
wire n_32538;
wire n_32539;
wire n_32540;
wire n_32541;
wire n_32542;
wire n_32543;
wire n_32544;
wire n_32545;
wire n_32546;
wire n_32547;
wire n_32548;
wire n_32549;
wire n_32550;
wire n_32551;
wire n_32552;
wire n_32553;
wire n_32554;
wire n_32555;
wire n_32556;
wire n_32557;
wire n_32558;
wire n_32559;
wire n_32560;
wire n_32561;
wire n_32562;
wire n_32563;
wire n_32564;
wire n_32565;
wire n_32566;
wire n_32567;
wire n_32568;
wire n_32569;
wire n_32570;
wire n_32571;
wire n_32572;
wire n_32573;
wire n_32574;
wire n_32575;
wire n_32576;
wire n_32577;
wire n_32578;
wire n_32579;
wire n_32580;
wire n_32581;
wire n_32582;
wire n_32583;
wire n_32584;
wire n_32585;
wire n_32586;
wire n_32587;
wire n_32588;
wire n_32589;
wire n_32590;
wire n_32591;
wire n_32592;
wire n_32593;
wire n_32594;
wire n_32595;
wire n_32596;
wire n_32597;
wire n_32598;
wire n_32599;
wire n_32600;
wire n_32601;
wire n_32602;
wire n_32603;
wire n_32604;
wire n_32605;
wire n_32606;
wire n_32607;
wire n_32608;
wire n_32609;
wire n_32610;
wire n_32611;
wire n_32612;
wire n_32613;
wire n_32614;
wire n_32615;
wire n_32616;
wire n_32617;
wire n_32618;
wire n_32619;
wire n_32620;
wire n_32621;
wire n_32622;
wire n_32623;
wire n_32624;
wire n_32625;
wire n_32626;
wire n_32627;
wire n_32628;
wire n_32629;
wire n_32630;
wire n_32631;
wire n_32632;
wire n_32633;
wire n_32634;
wire n_32635;
wire n_32636;
wire n_32637;
wire n_32638;
wire n_32639;
wire n_32640;
wire n_32641;
wire n_32642;
wire n_32643;
wire n_32644;
wire n_32645;
wire n_32646;
wire n_32647;
wire n_32648;
wire n_32649;
wire n_32650;
wire n_32651;
wire n_32652;
wire n_32653;
wire n_32654;
wire n_32655;
wire n_32656;
wire n_32657;
wire n_32658;
wire n_32659;
wire n_32660;
wire n_32661;
wire n_32662;
wire n_32663;
wire n_32664;
wire n_32665;
wire n_32666;
wire n_32667;
wire n_32668;
wire n_32669;
wire n_32670;
wire n_32671;
wire n_32672;
wire n_32673;
wire n_32674;
wire n_32675;
wire n_32676;
wire n_32677;
wire n_32678;
wire n_32679;
wire n_32680;
wire n_32681;
wire n_32682;
wire n_32683;
wire n_32684;
wire n_32685;
wire n_32686;
wire n_32687;
wire n_32688;
wire n_32689;
wire n_32690;
wire n_32691;
wire n_32692;
wire n_32693;
wire n_32694;
wire n_32695;
wire n_32696;
wire n_32697;
wire n_32698;
wire n_32699;
wire n_32700;
wire n_32701;
wire n_32702;
wire n_32703;
wire n_32704;
wire n_32705;
wire n_32706;
wire n_32707;
wire n_32708;
wire n_32709;
wire n_32710;
wire n_32711;
wire n_32712;
wire n_32713;
wire n_32714;
wire n_32715;
wire n_32716;
wire n_32717;
wire n_32718;
wire n_32719;
wire n_32720;
wire n_32721;
wire n_32722;
wire n_32723;
wire n_32724;
wire n_32725;
wire n_32726;
wire n_32727;
wire n_32728;
wire n_32729;
wire n_32730;
wire n_32731;
wire n_32732;
wire n_32733;
wire n_32734;
wire n_32735;
wire n_32736;
wire n_32737;
wire n_32738;
wire n_32739;
wire n_32740;
wire n_32741;
wire n_32742;
wire n_32743;
wire n_32744;
wire n_32745;
wire n_32746;
wire n_32747;
wire n_32748;
wire n_32749;
wire n_32750;
wire n_32751;
wire n_32752;
wire n_32753;
wire n_32754;
wire n_32755;
wire n_32756;
wire n_32757;
wire n_32758;
wire n_32759;
wire n_32760;
wire n_32761;
wire n_32762;
wire n_32763;
wire n_32764;
wire n_32765;
wire n_32766;
wire n_32767;
wire n_32768;
wire n_32769;
wire n_32770;
wire n_32771;
wire n_32772;
wire n_32773;
wire n_32774;
wire n_32775;
wire n_32776;
wire n_32777;
wire n_32778;
wire n_32779;
wire n_32780;
wire n_32781;
wire n_32782;
wire n_32783;
wire n_32784;
wire n_32785;
wire n_32786;
wire n_32787;
wire n_32788;
wire n_32789;
wire n_32790;
wire n_32791;
wire n_32792;
wire n_32793;
wire n_32794;
wire n_32795;
wire n_32796;
wire n_32797;
wire n_32798;
wire n_32799;
wire n_32800;
wire n_32801;
wire n_32802;
wire n_32803;
wire n_32804;
wire n_32805;
wire n_32806;
wire n_32807;
wire n_32808;
wire n_32809;
wire n_32810;
wire n_32811;
wire n_32812;
wire n_32813;
wire n_32814;
wire n_32815;
wire n_32816;
wire n_32817;
wire n_32818;
wire n_32819;
wire n_32820;
wire n_32821;
wire n_32822;
wire n_32823;
wire n_32824;
wire n_32825;
wire n_32826;
wire n_32827;
wire n_32828;
wire n_32829;
wire n_32830;
wire n_32831;
wire n_32832;
wire n_32833;
wire n_32834;
wire n_32835;
wire n_32836;
wire n_32837;
wire n_32838;
wire n_32839;
wire n_32840;
wire n_32841;
wire n_32842;
wire n_32843;
wire n_32844;
wire n_32845;
wire n_32846;
wire n_32847;
wire n_32848;
wire n_32849;
wire n_32850;
wire n_32851;
wire n_32852;
wire n_32853;
wire n_32854;
wire n_32855;
wire n_32856;
wire n_32857;
wire n_32858;
wire n_32859;
wire n_32860;
wire n_32861;
wire n_32862;
wire n_32863;
wire n_32864;
wire n_32865;
wire n_32866;
wire n_32867;
wire n_32868;
wire n_32869;
wire n_32870;
wire n_32871;
wire n_32872;
wire n_32873;
wire n_32874;
wire n_32875;
wire n_32876;
wire n_32877;
wire n_32878;
wire n_32879;
wire n_32880;
wire n_32881;
wire n_32882;
wire n_32883;
wire n_32884;
wire n_32885;
wire n_32886;
wire n_32887;
wire n_32888;
wire n_32889;
wire n_32890;
wire n_32891;
wire n_32892;
wire n_32893;
wire n_32894;
wire n_32895;
wire n_32896;
wire n_32897;
wire n_32898;
wire n_32899;
wire n_32900;
wire n_32901;
wire n_32902;
wire n_32903;
wire n_32904;
wire n_32905;
wire n_32906;
wire n_32907;
wire n_32908;
wire n_32909;
wire n_32910;
wire n_32911;
wire n_32912;
wire n_32913;
wire n_32914;
wire n_32915;
wire n_32916;
wire n_32917;
wire n_32918;
wire n_32919;
wire n_32920;
wire n_32921;
wire n_32922;
wire n_32923;
wire n_32924;
wire n_32925;
wire n_32926;
wire n_32927;
wire n_32928;
wire n_32929;
wire n_32930;
wire n_32931;
wire n_32932;
wire n_32933;
wire n_32934;
wire n_32935;
wire n_32936;
wire n_32937;
wire n_32938;
wire n_32939;
wire n_32940;
wire n_32941;
wire n_32942;
wire n_32943;
wire n_32944;
wire n_32945;
wire n_32946;
wire n_32947;
wire n_32948;
wire n_32949;
wire n_32950;
wire n_32951;
wire n_32952;
wire n_32953;
wire n_32954;
wire n_32955;
wire n_32956;
wire n_32957;
wire n_32958;
wire n_32959;
wire n_32960;
wire n_32961;
wire n_32962;
wire n_32963;
wire n_32964;
wire n_32965;
wire n_32966;
wire n_32967;
wire n_32968;
wire n_32969;
wire n_32970;
wire n_32971;
wire n_32972;
wire n_32973;
wire n_32974;
wire n_32975;
wire n_32976;
wire n_32977;
wire n_32978;
wire n_32979;
wire n_32980;
wire n_32981;
wire n_32982;
wire n_32983;
wire n_32984;
wire n_32985;
wire n_32986;
wire n_32987;
wire n_32988;
wire n_32989;
wire n_32990;
wire n_32991;
wire n_32992;
wire n_32993;
wire n_32994;
wire n_32995;
wire n_32996;
wire n_32997;
wire n_32998;
wire n_32999;
wire n_33000;
wire n_33001;
wire n_33002;
wire n_33003;
wire n_33004;
wire n_33005;
wire n_33006;
wire n_33007;
wire n_33008;
wire n_33009;
wire n_33010;
wire n_33011;
wire n_33012;
wire n_33013;
wire n_33014;
wire n_33015;
wire n_33016;
wire n_33017;
wire n_33018;
wire n_33019;
wire n_33020;
wire n_33021;
wire n_33022;
wire n_33023;
wire n_33024;
wire n_33025;
wire n_33026;
wire n_33027;
wire n_33028;
wire n_33029;
wire n_33030;
wire n_33031;
wire n_33032;
wire n_33033;
wire n_33034;
wire n_33035;
wire n_33036;
wire n_33037;
wire n_33038;
wire n_33039;
wire n_33040;
wire n_33041;
wire n_33042;
wire n_33043;
wire n_33044;
wire n_33045;
wire n_33046;
wire n_33047;
wire n_33048;
wire n_33049;
wire n_33050;
wire n_33051;
wire n_33052;
wire n_33053;
wire n_33054;
wire n_33055;
wire n_33056;
wire n_33057;
wire n_33058;
wire n_33059;
wire n_33060;
wire n_33061;
wire n_33062;
wire n_33063;
wire n_33064;
wire n_33065;
wire n_33066;
wire n_33067;
wire n_33068;
wire n_33069;
wire n_33070;
wire n_33071;
wire n_33072;
wire n_33073;
wire n_33074;
wire n_33075;
wire n_33076;
wire n_33077;
wire n_33078;
wire n_33079;
wire n_33080;
wire n_33081;
wire n_33082;
wire n_33083;
wire n_33084;
wire n_33085;
wire n_33086;
wire n_33087;
wire n_33088;
wire n_33089;
wire n_33090;
wire n_33091;
wire n_33092;
wire n_33093;
wire n_33094;
wire n_33095;
wire n_33096;
wire n_33097;
wire n_33098;
wire n_33099;
wire n_33100;
wire n_33101;
wire n_33102;
wire n_33103;
wire n_33104;
wire n_33105;
wire n_33106;
wire n_33107;
wire n_33108;
wire n_33109;
wire n_33110;
wire n_33111;
wire n_33112;
wire n_33113;
wire n_33114;
wire n_33115;
wire n_33116;
wire n_33117;
wire n_33118;
wire n_33119;
wire n_33120;
wire n_33121;
wire n_33122;
wire n_33123;
wire n_33124;
wire n_33125;
wire n_33126;
wire n_33127;
wire n_33128;
wire n_33129;
wire n_33130;
wire n_33131;
wire n_33132;
wire n_33133;
wire n_33134;
wire n_33135;
wire n_33136;
wire n_33137;
wire n_33138;
wire n_33139;
wire n_33140;
wire n_33141;
wire n_33142;
wire n_33143;
wire n_33144;
wire n_33145;
wire n_33146;
wire n_33147;
wire n_33148;
wire n_33149;
wire n_33150;
wire n_33151;
wire n_33152;
wire n_33153;
wire n_33154;
wire n_33155;
wire n_33156;
wire n_33157;
wire n_33158;
wire n_33159;
wire n_33160;
wire n_33161;
wire n_33162;
wire n_33163;
wire n_33164;
wire n_33165;
wire n_33166;
wire n_33167;
wire n_33168;
wire n_33169;
wire n_33170;
wire n_33171;
wire n_33172;
wire n_33173;
wire n_33174;
wire n_33175;
wire n_33176;
wire n_33177;
wire n_33178;
wire n_33179;
wire n_33180;
wire n_33181;
wire n_33182;
wire n_33183;
wire n_33184;
wire n_33185;
wire n_33186;
wire n_33187;
wire n_33188;
wire n_33189;
wire n_33190;
wire n_33191;
wire n_33192;
wire n_33193;
wire n_33194;
wire n_33195;
wire n_33196;
wire n_33197;
wire n_33198;
wire n_33199;
wire n_33200;
wire n_33201;
wire n_33202;
wire n_33203;
wire n_33204;
wire n_33205;
wire n_33206;
wire n_33207;
wire n_33208;
wire n_33209;
wire n_33210;
wire n_33211;
wire n_33212;
wire n_33213;
wire n_33214;
wire n_33215;
wire n_33216;
wire n_33217;
wire n_33218;
wire n_33219;
wire n_33220;
wire n_33221;
wire n_33222;
wire n_33223;
wire n_33224;
wire n_33225;
wire n_33226;
wire n_33227;
wire n_33228;
wire n_33229;
wire n_33230;
wire n_33231;
wire n_33232;
wire n_33233;
wire n_33234;
wire n_33235;
wire n_33236;
wire n_33237;
wire n_33238;
wire n_33239;
wire n_33240;
wire n_33241;
wire n_33242;
wire n_33243;
wire n_33244;
wire n_33245;
wire n_33246;
wire n_33247;
wire n_33248;
wire n_33249;
wire n_33250;
wire n_33251;
wire n_33252;
wire n_33253;
wire n_33254;
wire n_33255;
wire n_33256;
wire n_33257;
wire n_33258;
wire n_33259;
wire n_33260;
wire n_33261;
wire n_33262;
wire n_33263;
wire n_33264;
wire n_33265;
wire n_33266;
wire n_33267;
wire n_33268;
wire n_33269;
wire n_33270;
wire n_33271;
wire n_33272;
wire n_33273;
wire n_33274;
wire n_33275;
wire n_33276;
wire n_33277;
wire n_33278;
wire n_33279;
wire n_33280;
wire n_33281;
wire n_33282;
wire n_33283;
wire n_33284;
wire n_33285;
wire n_33286;
wire n_33287;
wire n_33288;
wire n_33289;
wire n_33290;
wire n_33291;
wire n_33292;
wire n_33293;
wire n_33294;
wire n_33295;
wire n_33296;
wire n_33297;
wire n_33298;
wire n_33299;
wire n_33300;
wire n_33301;
wire n_33302;
wire n_33303;
wire n_33304;
wire n_33305;
wire n_33306;
wire n_33307;
wire n_33308;
wire n_33309;
wire n_33310;
wire n_33311;
wire n_33312;
wire n_33313;
wire n_33314;
wire n_33315;
wire n_33316;
wire n_33317;
wire n_33318;
wire n_33319;
wire n_33320;
wire n_33321;
wire n_33322;
wire n_33323;
wire n_33324;
wire n_33325;
wire n_33326;
wire n_33327;
wire n_33328;
wire n_33329;
wire n_33330;
wire n_33331;
wire n_33332;
wire n_33333;
wire n_33334;
wire n_33335;
wire n_33336;
wire n_33337;
wire n_33338;
wire n_33339;
wire n_33340;
wire n_33341;
wire n_33342;
wire n_33343;
wire n_33344;
wire n_33345;
wire n_33346;
wire n_33347;
wire n_33348;
wire n_33349;
wire n_33350;
wire n_33351;
wire n_33352;
wire n_33353;
wire n_33354;
wire n_33355;
wire n_33356;
wire n_33357;
wire n_33358;
wire n_33359;
wire n_33360;
wire n_33361;
wire n_33362;
wire n_33363;
wire n_33364;
wire n_33365;
wire n_33366;
wire n_33367;
wire n_33368;
wire n_33369;
wire n_33370;
wire n_33371;
wire n_33372;
wire n_33373;
wire n_33374;
wire n_33375;
wire n_33376;
wire n_33377;
wire n_33378;
wire n_33379;
wire n_33380;
wire n_33381;
wire n_33382;
wire n_33383;
wire n_33384;
wire n_33385;
wire n_33386;
wire n_33387;
wire n_33388;
wire n_33389;
wire n_33390;
wire n_33391;
wire n_33392;
wire n_33393;
wire n_33394;
wire n_33395;
wire n_33396;
wire n_33397;
wire n_33398;
wire n_33399;
wire n_33400;
wire n_33401;
wire n_33402;
wire n_33403;
wire n_33404;
wire n_33405;
wire n_33406;
wire n_33407;
wire n_33408;
wire n_33409;
wire n_33410;
wire n_33411;
wire n_33412;
wire n_33413;
wire n_33414;
wire n_33415;
wire n_33416;
wire n_33417;
wire n_33418;
wire n_33419;
wire n_33420;
wire n_33421;
wire n_33422;
wire n_33423;
wire n_33424;
wire n_33425;
wire n_33426;
wire n_33427;
wire n_33428;
wire n_33429;
wire n_33430;
wire n_33431;
wire n_33432;
wire n_33433;
wire n_33434;
wire n_33435;
wire n_33436;
wire n_33437;
wire n_33438;
wire n_33439;
wire n_33440;
wire n_33441;
wire n_33442;
wire n_33443;
wire n_33444;
wire n_33445;
wire n_33446;
wire n_33447;
wire n_33448;
wire n_33449;
wire n_33450;
wire n_33451;
wire n_33452;
wire n_33453;
wire n_33454;
wire n_33455;
wire n_33456;
wire n_33457;
wire n_33458;
wire n_33459;
wire n_33460;
wire n_33461;
wire n_33462;
wire n_33463;
wire n_33464;
wire n_33465;
wire n_33466;
wire n_33467;
wire n_33468;
wire n_33469;
wire n_33470;
wire n_33471;
wire n_33472;
wire n_33473;
wire n_33474;
wire n_33475;
wire n_33476;
wire n_33477;
wire n_33478;
wire n_33479;
wire n_33480;
wire n_33481;
wire n_33482;
wire n_33483;
wire n_33484;
wire n_33485;
wire n_33486;
wire n_33487;
wire n_33488;
wire n_33489;
wire n_33490;
wire n_33491;
wire n_33492;
wire n_33493;
wire n_33494;
wire n_33495;
wire n_33496;
wire n_33497;
wire n_33498;
wire n_33499;
wire n_33500;
wire n_33501;
wire n_33502;
wire n_33503;
wire n_33504;
wire n_33505;
wire n_33506;
wire n_33507;
wire n_33508;
wire n_33509;
wire n_33510;
wire n_33511;
wire n_33512;
wire n_33513;
wire n_33514;
wire n_33515;
wire n_33516;
wire n_33517;
wire n_33518;
wire n_33519;
wire n_33520;
wire n_33521;
wire n_33522;
wire n_33523;
wire n_33524;
wire n_33525;
wire n_33526;
wire n_33527;
wire n_33528;
wire n_33529;
wire n_33530;
wire n_33531;
wire n_33532;
wire n_33533;
wire n_33534;
wire n_33535;
wire n_33536;
wire n_33537;
wire n_33538;
wire n_33539;
wire n_33540;
wire n_33541;
wire n_33542;
wire n_33543;
wire n_33544;
wire n_33545;
wire n_33546;
wire n_33547;
wire n_33548;
wire n_33549;
wire n_33550;
wire n_33551;
wire n_33552;
wire n_33553;
wire n_33554;
wire n_33555;
wire n_33556;
wire n_33557;
wire n_33558;
wire n_33559;
wire n_33560;
wire n_33561;
wire n_33562;
wire n_33563;
wire n_33564;
wire n_33565;
wire n_33566;
wire n_33567;
wire n_33568;
wire n_33569;
wire n_33570;
wire n_33571;
wire n_33572;
wire n_33573;
wire n_33574;
wire n_33575;
wire n_33576;
wire n_33577;
wire n_33578;
wire n_33579;
wire n_33580;
wire n_33581;
wire n_33582;
wire n_33583;
wire n_33584;
wire n_33585;
wire n_33586;
wire n_33587;
wire n_33588;
wire n_33589;
wire n_33590;
wire n_33591;
wire n_33592;
wire n_33593;
wire n_33594;
wire n_33595;
wire n_33596;
wire n_33597;
wire n_33598;
wire n_33599;
wire n_33600;
wire n_33601;
wire n_33602;
wire n_33603;
wire n_33604;
wire n_33605;
wire n_33606;
wire n_33607;
wire n_33608;
wire n_33609;
wire n_33610;
wire n_33611;
wire n_33612;
wire n_33613;
wire n_33614;
wire n_33615;
wire n_33616;
wire n_33617;
wire n_33618;
wire n_33619;
wire n_33620;
wire n_33621;
wire n_33622;
wire n_33623;
wire n_33624;
wire n_33625;
wire n_33626;
wire n_33627;
wire n_33628;
wire n_33629;
wire n_33630;
wire n_33631;
wire n_33632;
wire n_33633;
wire n_33634;
wire n_33635;
wire n_33636;
wire n_33637;
wire n_33638;
wire n_33639;
wire n_33640;
wire n_33641;
wire n_33642;
wire n_33643;
wire n_33644;
wire n_33645;
wire n_33646;
wire n_33647;
wire n_33648;
wire n_33649;
wire n_33650;
wire n_33651;
wire n_33652;
wire n_33653;
wire n_33654;
wire n_33655;
wire n_33656;
wire n_33657;
wire n_33658;
wire n_33659;
wire n_33660;
wire n_33661;
wire n_33662;
wire n_33663;
wire n_33664;
wire n_33665;
wire n_33666;
wire n_33667;
wire n_33668;
wire n_33669;
wire n_33670;
wire n_33671;
wire n_33672;
wire n_33673;
wire n_33674;
wire n_33675;
wire n_33676;
wire n_33677;
wire n_33678;
wire n_33679;
wire n_33680;
wire n_33681;
wire n_33682;
wire n_33683;
wire n_33684;
wire n_33685;
wire n_33686;
wire n_33687;
wire n_33688;
wire n_33689;
wire n_33690;
wire n_33691;
wire n_33692;
wire n_33693;
wire n_33694;
wire n_33695;
wire n_33696;
wire n_33697;
wire n_33698;
wire n_33699;
wire n_33700;
wire n_33701;
wire n_33702;
wire n_33703;
wire n_33704;
wire n_33705;
wire n_33706;
wire n_33707;
wire n_33708;
wire n_33709;
wire n_33710;
wire n_33711;
wire n_33712;
wire n_33713;
wire n_33714;
wire n_33715;
wire n_33716;
wire n_33717;
wire n_33718;
wire n_33719;
wire n_33720;
wire n_33721;
wire n_33722;
wire n_33723;
wire n_33724;
wire n_33725;
wire n_33726;
wire n_33727;
wire n_33728;
wire n_33729;
wire n_33730;
wire n_33731;
wire n_33732;
wire n_33733;
wire n_33734;
wire n_33735;
wire n_33736;
wire n_33737;
wire n_33738;
wire n_33739;
wire n_33740;
wire n_33741;
wire n_33742;
wire n_33743;
wire n_33744;
wire n_33745;
wire n_33746;
wire n_33747;
wire n_33748;
wire n_33749;
wire n_33750;
wire n_33751;
wire n_33752;
wire n_33753;
wire n_33754;
wire n_33755;
wire n_33756;
wire n_33757;
wire n_33758;
wire n_33759;
wire n_33760;
wire n_33761;
wire n_33762;
wire n_33763;
wire n_33764;
wire n_33765;
wire n_33766;
wire n_33767;
wire n_33768;
wire n_33769;
wire n_33770;
wire n_33771;
wire n_33772;
wire n_33773;
wire n_33774;
wire n_33775;
wire n_33776;
wire n_33777;
wire n_33778;
wire n_33779;
wire n_33780;
wire n_33781;
wire n_33782;
wire n_33783;
wire n_33784;
wire n_33785;
wire n_33786;
wire n_33787;
wire n_33788;
wire n_33789;
wire n_33790;
wire n_33791;
wire n_33792;
wire n_33793;
wire n_33794;
wire n_33795;
wire n_33796;
wire n_33797;
wire n_33798;
wire n_33799;
wire n_33800;
wire n_33801;
wire n_33802;
wire n_33803;
wire n_33804;
wire n_33805;
wire n_33806;
wire n_33807;
wire n_33808;
wire n_33809;
wire n_33810;
wire n_33811;
wire n_33812;
wire n_33813;
wire n_33814;
wire n_33815;
wire n_33816;
wire n_33817;
wire n_33818;
wire n_33819;
wire n_33820;
wire n_33821;
wire n_33822;
wire n_33823;
wire n_33824;
wire n_33825;
wire n_33826;
wire n_33827;
wire n_33828;
wire n_33829;
wire n_33830;
wire n_33831;
wire n_33832;
wire n_33833;
wire n_33834;
wire n_33835;
wire n_33836;
wire n_33837;
wire n_33838;
wire n_33839;
wire n_33840;
wire n_33841;
wire n_33842;
wire n_33843;
wire n_33844;
wire n_33845;
wire n_33846;
wire n_33847;
wire n_33848;
wire n_33849;
wire n_33850;
wire n_33851;
wire n_33852;
wire n_33853;
wire n_33854;
wire n_33855;
wire n_33856;
wire n_33857;
wire n_33858;
wire n_33859;
wire n_33860;
wire n_33861;
wire n_33862;
wire n_33863;
wire n_33864;
wire n_33865;
wire n_33866;
wire n_33867;
wire n_33868;
wire n_33869;
wire n_33870;
wire n_33871;
wire n_33872;
wire n_33873;
wire n_33874;
wire n_33875;
wire n_33876;
wire n_33877;
wire n_33878;
wire n_33879;
wire n_33880;
wire n_33881;
wire n_33882;
wire n_33883;
wire n_33884;
wire n_33885;
wire n_33886;
wire n_33887;
wire n_33888;
wire n_33889;
wire n_33890;
wire n_33891;
wire n_33892;
wire n_33893;
wire n_33894;
wire n_33895;
wire n_33896;
wire n_33897;
wire n_33898;
wire n_33899;
wire n_33900;
wire n_33901;
wire n_33902;
wire n_33903;
wire n_33904;
wire n_33905;
wire n_33906;
wire n_33907;
wire n_33908;
wire n_33909;
wire n_33910;
wire n_33911;
wire n_33912;
wire n_33913;
wire n_33914;
wire n_33915;
wire n_33916;
wire n_33917;
wire n_33918;
wire n_33919;
wire n_33920;
wire n_33921;
wire n_33922;
wire n_33923;
wire n_33924;
wire n_33925;
wire n_33926;
wire n_33927;
wire n_33928;
wire n_33929;
wire n_33930;
wire n_33931;
wire n_33932;
wire n_33933;
wire n_33934;
wire n_33935;
wire n_33936;
wire n_33937;
wire n_33938;
wire n_33939;
wire n_33940;
wire n_33941;
wire n_33942;
wire n_33943;
wire n_33944;
wire n_33945;
wire n_33946;
wire n_33947;
wire n_33948;
wire n_33949;
wire n_33950;
wire n_33951;
wire n_33952;
wire n_33953;
wire n_33954;
wire n_33955;
wire n_33956;
wire n_33957;
wire n_33958;
wire n_33959;
wire n_33960;
wire n_33961;
wire n_33962;
wire n_33963;
wire n_33964;
wire n_33965;
wire n_33966;
wire n_33967;
wire n_33968;
wire n_33969;
wire n_33970;
wire n_33971;
wire n_33972;
wire n_33973;
wire n_33974;
wire n_33975;
wire n_33976;
wire n_33977;
wire n_33978;
wire n_33979;
wire n_33980;
wire n_33981;
wire n_33982;
wire n_33983;
wire n_33984;
wire n_33985;
wire n_33986;
wire n_33987;
wire n_33988;
wire n_33989;
wire n_33990;
wire n_33991;
wire n_33992;
wire n_33993;
wire n_33994;
wire n_33995;
wire n_33996;
wire n_33997;
wire n_33998;
wire n_33999;
wire n_34000;
wire n_34001;
wire n_34002;
wire n_34003;
wire n_34004;
wire n_34005;
wire n_34006;
wire n_34007;
wire n_34008;
wire n_34009;
wire n_34010;
wire n_34011;
wire n_34012;
wire n_34013;
wire n_34014;
wire n_34015;
wire n_34016;
wire n_34017;
wire n_34018;
wire n_34019;
wire n_34020;
wire n_34021;
wire n_34022;
wire n_34023;
wire n_34024;
wire n_34025;
wire n_34026;
wire n_34027;
wire n_34028;
wire n_34029;
wire n_34030;
wire n_34031;
wire n_34032;
wire n_34033;
wire n_34034;
wire n_34035;
wire n_34036;
wire n_34037;
wire n_34038;
wire n_34039;
wire n_34040;
wire n_34041;
wire n_34042;
wire n_34043;
wire n_34044;
wire n_34045;
wire n_34046;
wire n_34047;
wire n_34048;
wire n_34049;
wire n_34050;
wire n_34051;
wire n_34052;
wire n_34053;
wire n_34054;
wire n_34055;
wire n_34056;
wire n_34057;
wire n_34058;
wire n_34059;
wire n_34060;
wire n_34061;
wire n_34062;
wire n_34063;
wire n_34064;
wire n_34065;
wire n_34066;
wire n_34067;
wire n_34068;
wire n_34069;
wire n_34070;
wire n_34071;
wire n_34072;
wire n_34073;
wire n_34074;
wire n_34075;
wire n_34076;
wire n_34077;
wire n_34078;
wire n_34079;
wire n_34080;
wire n_34081;
wire n_34082;
wire n_34083;
wire n_34084;
wire n_34085;
wire n_34086;
wire n_34087;
wire n_34088;
wire n_34089;
wire n_34090;
wire n_34091;
wire n_34092;
wire n_34093;
wire n_34094;
wire n_34095;
wire n_34096;
wire n_34097;
wire n_34098;
wire n_34099;
wire n_34100;
wire n_34101;
wire n_34102;
wire n_34103;
wire n_34104;
wire n_34105;
wire n_34106;
wire n_34107;
wire n_34108;
wire n_34109;
wire n_34110;
wire n_34111;
wire n_34112;
wire n_34113;
wire n_34114;
wire n_34115;
wire n_34116;
wire n_34117;
wire n_34118;
wire n_34119;
wire n_34120;
wire n_34121;
wire n_34122;
wire n_34123;
wire n_34124;
wire n_34125;
wire n_34126;
wire n_34127;
wire n_34128;
wire n_34129;
wire n_34130;
wire n_34131;
wire n_34132;
wire n_34133;
wire n_34134;
wire n_34135;
wire n_34136;
wire n_34137;
wire n_34138;
wire n_34139;
wire n_34140;
wire n_34141;
wire n_34142;
wire n_34143;
wire n_34144;
wire n_34145;
wire n_34146;
wire n_34147;
wire n_34148;
wire n_34149;
wire n_34150;
wire n_34151;
wire n_34152;
wire n_34153;
wire n_34154;
wire n_34155;
wire n_34156;
wire n_34157;
wire n_34158;
wire n_34159;
wire n_34160;
wire n_34161;
wire n_34162;
wire n_34163;
wire n_34164;
wire n_34165;
wire n_34166;
wire n_34167;
wire n_34168;
wire n_34169;
wire n_34170;
wire n_34171;
wire n_34172;
wire n_34173;
wire n_34174;
wire n_34175;
wire n_34176;
wire n_34177;
wire n_34178;
wire n_34179;
wire n_34180;
wire n_34181;
wire n_34182;
wire n_34183;
wire n_34184;
wire n_34185;
wire n_34186;
wire n_34187;
wire n_34188;
wire n_34189;
wire n_34190;
wire n_34191;
wire n_34192;
wire n_34193;
wire n_34194;
wire n_34195;
wire n_34196;
wire n_34197;
wire n_34198;
wire n_34199;
wire n_34200;
wire n_34201;
wire n_34202;
wire n_34203;
wire n_34204;
wire n_34205;
wire n_34206;
wire n_34207;
wire n_34208;
wire n_34209;
wire n_34210;
wire n_34211;
wire n_34212;
wire n_34213;
wire n_34214;
wire n_34215;
wire n_34216;
wire n_34217;
wire n_34218;
wire n_34219;
wire n_34220;
wire n_34221;
wire n_34222;
wire n_34223;
wire n_34224;
wire n_34225;
wire n_34226;
wire n_34227;
wire n_34228;
wire n_34229;
wire n_34230;
wire n_34231;
wire n_34232;
wire n_34233;
wire n_34234;
wire n_34235;
wire n_34236;
wire n_34237;
wire n_34238;
wire n_34239;
wire n_34240;
wire n_34241;
wire n_34242;
wire n_34243;
wire n_34244;
wire n_34245;
wire n_34246;
wire n_34247;
wire n_34248;
wire n_34249;
wire n_34250;
wire n_34251;
wire n_34252;
wire n_34253;
wire n_34254;
wire n_34255;
wire n_34256;
wire n_34257;
wire n_34258;
wire n_34259;
wire n_34260;
wire n_34261;
wire n_34262;
wire n_34263;
wire n_34264;
wire n_34265;
wire n_34266;
wire n_34267;
wire n_34268;
wire n_34269;
wire n_34270;
wire n_34271;
wire n_34272;
wire n_34273;
wire n_34274;
wire n_34275;
wire n_34276;
wire n_34277;
wire n_34278;
wire n_34279;
wire n_34280;
wire n_34281;
wire n_34282;
wire n_34283;
wire n_34284;
wire n_34285;
wire n_34286;
wire n_34287;
wire n_34288;
wire n_34289;
wire n_34290;
wire n_34291;
wire n_34292;
wire n_34293;
wire n_34294;
wire n_34295;
wire n_34296;
wire n_34297;
wire n_34298;
wire n_34299;
wire n_34300;
wire n_34301;
wire n_34302;
wire n_34303;
wire n_34304;
wire n_34305;
wire n_34306;
wire n_34307;
wire n_34308;
wire n_34309;
wire n_34310;
wire n_34311;
wire n_34312;
wire n_34313;
wire n_34314;
wire n_34315;
wire n_34316;
wire n_34317;
wire n_34318;
wire n_34319;
wire n_34320;
wire n_34321;
wire n_34322;
wire n_34323;
wire n_34324;
wire n_34325;
wire n_34326;
wire n_34327;
wire n_34328;
wire n_34329;
wire n_34330;
wire n_34331;
wire n_34332;
wire n_34333;
wire n_34334;
wire n_34335;
wire n_34336;
wire n_34337;
wire n_34338;
wire n_34339;
wire n_34340;
wire n_34341;
wire n_34342;
wire n_34343;
wire n_34344;
wire n_34345;
wire n_34346;
wire n_34347;
wire n_34348;
wire n_34349;
wire n_34350;
wire n_34351;
wire n_34352;
wire n_34353;
wire n_34354;
wire n_34355;
wire n_34356;
wire n_34357;
wire n_34358;
wire n_34359;
wire n_34360;
wire n_34361;
wire n_34362;
wire n_34363;
wire n_34364;
wire n_34365;
wire n_34366;
wire n_34367;
wire n_34368;
wire n_34369;
wire n_34370;
wire n_34371;
wire n_34372;
wire n_34373;
wire n_34374;
wire n_34375;
wire n_34376;
wire n_34377;
wire n_34378;
wire n_34379;
wire n_34380;
wire n_34381;
wire n_34382;
wire n_34383;
wire n_34384;
wire n_34385;
wire n_34386;
wire n_34387;
wire n_34388;
wire n_34389;
wire n_34390;
wire n_34391;
wire n_34392;
wire n_34393;
wire n_34394;
wire n_34395;
wire n_34396;
wire n_34397;
wire n_34398;
wire n_34399;
wire n_34400;
wire n_34401;
wire n_34402;
wire n_34403;
wire n_34404;
wire n_34405;
wire n_34406;
wire n_34407;
wire n_34408;
wire n_34409;
wire n_34410;
wire n_34411;
wire n_34412;
wire n_34413;
wire n_34414;
wire n_34415;
wire n_34416;
wire n_34417;
wire n_34418;
wire n_34419;
wire n_34420;
wire n_34421;
wire n_34422;
wire n_34423;
wire n_34424;
wire n_34425;
wire n_34426;
wire n_34427;
wire n_34428;
wire n_34429;
wire n_34430;
wire n_34431;
wire n_34432;
wire n_34433;
wire n_34434;
wire n_34435;
wire n_34436;
wire n_34437;
wire n_34438;
wire n_34439;
wire n_34440;
wire n_34441;
wire n_34442;
wire n_34443;
wire n_34444;
wire n_34445;
wire n_34446;
wire n_34447;
wire n_34448;
wire n_34449;
wire n_34450;
wire n_34451;
wire n_34452;
wire n_34453;
wire n_34454;
wire n_34455;
wire n_34456;
wire n_34457;
wire n_34458;
wire n_34459;
wire n_34460;
wire n_34461;
wire n_34462;
wire n_34463;
wire n_34464;
wire n_34465;
wire n_34466;
wire n_34467;
wire n_34468;
wire n_34469;
wire n_34470;
wire n_34471;
wire n_34472;
wire n_34473;
wire n_34474;
wire n_34475;
wire n_34476;
wire n_34477;
wire n_34478;
wire n_34479;
wire n_34480;
wire n_34481;
wire n_34482;
wire n_34483;
wire n_34484;
wire n_34485;
wire n_34486;
wire n_34487;
wire n_34488;
wire n_34489;
wire n_34490;
wire n_34491;
wire n_34492;
wire n_34493;
wire n_34494;
wire n_34495;
wire n_34496;
wire n_34497;
wire n_34498;
wire n_34499;
wire n_34500;
wire n_34501;
wire n_34502;
wire n_34503;
wire n_34504;
wire n_34505;
wire n_34506;
wire n_34507;
wire n_34508;
wire n_34509;
wire n_34510;
wire n_34511;
wire n_34512;
wire n_34513;
wire n_34514;
wire n_34515;
wire n_34516;
wire n_34517;
wire n_34518;
wire n_34519;
wire n_34520;
wire n_34521;
wire n_34522;
wire n_34523;
wire n_34524;
wire n_34525;
wire n_34526;
wire n_34527;
wire n_34528;
wire n_34529;
wire n_34530;
wire n_34531;
wire n_34532;
wire n_34533;
wire n_34534;
wire n_34535;
wire n_34536;
wire n_34537;
wire n_34538;
wire n_34539;
wire n_34540;
wire n_34541;
wire n_34542;
wire n_34543;
wire n_34544;
wire n_34545;
wire n_34546;
wire n_34547;
wire n_34548;
wire n_34549;
wire n_34550;
wire n_34551;
wire n_34552;
wire n_34553;
wire n_34554;
wire n_34555;
wire n_34556;
wire n_34557;
wire n_34558;
wire n_34559;
wire n_34560;
wire n_34561;
wire n_34562;
wire n_34563;
wire n_34564;
wire n_34565;
wire n_34566;
wire n_34567;
wire n_34568;
wire n_34569;
wire n_34570;
wire n_34571;
wire n_34572;
wire n_34573;
wire n_34574;
wire n_34575;
wire n_34576;
wire n_34577;
wire n_34578;
wire n_34579;
wire n_34580;
wire n_34581;
wire n_34582;
wire n_34583;
wire n_34584;
wire n_34585;
wire n_34586;
wire n_34587;
wire n_34588;
wire n_34589;
wire n_34590;
wire n_34591;
wire n_34592;
wire n_34593;
wire n_34594;
wire n_34595;
wire n_34596;
wire n_34597;
wire n_34598;
wire n_34599;
wire n_34600;
wire n_34601;
wire n_34602;
wire n_34603;
wire n_34604;
wire n_34605;
wire n_34606;
wire n_34607;
wire n_34608;
wire n_34609;
wire n_34610;
wire n_34611;
wire n_34612;
wire n_34613;
wire n_34614;
wire n_34615;
wire n_34616;
wire n_34617;
wire n_34618;
wire n_34619;
wire n_34620;
wire n_34621;
wire n_34622;
wire n_34623;
wire n_34624;
wire n_34625;
wire n_34626;
wire n_34627;
wire n_34628;
wire n_34629;
wire n_34630;
wire n_34631;
wire n_34632;
wire n_34633;
wire n_34634;
wire n_34635;
wire n_34636;
wire n_34637;
wire n_34638;
wire n_34639;
wire n_34640;
wire n_34641;
wire n_34642;
wire n_34643;
wire n_34644;
wire n_34645;
wire n_34646;
wire n_34647;
wire n_34648;
wire n_34649;
wire n_34650;
wire n_34651;
wire n_34652;
wire n_34653;
wire n_34654;
wire n_34655;
wire n_34656;
wire n_34657;
wire n_34658;
wire n_34659;
wire n_34660;
wire n_34661;
wire n_34662;
wire n_34663;
wire n_34664;
wire n_34665;
wire n_34666;
wire n_34667;
wire n_34668;
wire n_34669;
wire n_34670;
wire n_34671;
wire n_34672;
wire n_34673;
wire n_34674;
wire n_34675;
wire n_34676;
wire n_34677;
wire n_34678;
wire n_34679;
wire n_34680;
wire n_34681;
wire n_34682;
wire n_34683;
wire n_34684;
wire n_34685;
wire n_34686;
wire n_34687;
wire n_34688;
wire n_34689;
wire n_34690;
wire n_34691;
wire n_34692;
wire n_34693;
wire n_34694;
wire n_34695;
wire n_34696;
wire n_34697;
wire n_34698;
wire n_34699;
wire n_34700;
wire n_34701;
wire n_34702;
wire n_34703;
wire n_34704;
wire n_34705;
wire n_34706;
wire n_34707;
wire n_34708;
wire n_34709;
wire n_34710;
wire n_34711;
wire n_34712;
wire n_34713;
wire n_34714;
wire n_34715;
wire n_34716;
wire n_34717;
wire n_34718;
wire n_34719;
wire n_34720;
wire n_34721;
wire n_34722;
wire n_34723;
wire n_34724;
wire n_34725;
wire n_34726;
wire n_34727;
wire n_34728;
wire n_34729;
wire n_34730;
wire n_34731;
wire n_34732;
wire n_34733;
wire n_34734;
wire n_34735;
wire n_34736;
wire n_34737;
wire n_34738;
wire n_34739;
wire n_34740;
wire n_34741;
wire n_34742;
wire n_34743;
wire n_34744;
wire n_34745;
wire n_34746;
wire n_34747;
wire n_34748;
wire n_34749;
wire n_34750;
wire n_34751;
wire n_34752;
wire n_34753;
wire n_34754;
wire n_34755;
wire n_34756;
wire n_34757;
wire n_34758;
wire n_34759;
wire n_34760;
wire n_34761;
wire n_34762;
wire n_34763;
wire n_34764;
wire n_34765;
wire n_34766;
wire n_34767;
wire n_34768;
wire n_34769;
wire n_34770;
wire n_34771;
wire n_34772;
wire n_34773;
wire n_34774;
wire n_34775;
wire n_34776;
wire n_34777;
wire n_34778;
wire n_34779;
wire n_34780;
wire n_34781;
wire n_34782;
wire n_34783;
wire n_34784;
wire n_34785;
wire n_34786;
wire n_34787;
wire n_34788;
wire n_34789;
wire n_34790;
wire n_34791;
wire n_34792;
wire n_34793;
wire n_34794;
wire n_34795;
wire n_34796;
wire n_34797;
wire n_34798;
wire n_34799;
wire n_34800;
wire n_34801;
wire n_34802;
wire n_34803;
wire n_34804;
wire n_34805;
wire n_34806;
wire n_34807;
wire n_34808;
wire n_34809;
wire n_34810;
wire n_34811;
wire n_34812;
wire n_34813;
wire n_34814;
wire n_34815;
wire n_34816;
wire n_34817;
wire n_34818;
wire n_34819;
wire n_34820;
wire n_34821;
wire n_34822;
wire n_34823;
wire n_34824;
wire n_34825;
wire n_34826;
wire n_34827;
wire n_34828;
wire n_34829;
wire n_34830;
wire n_34831;
wire n_34832;
wire n_34833;
wire n_34834;
wire n_34835;
wire n_34836;
wire n_34837;
wire n_34838;
wire n_34839;
wire n_34840;
wire n_34841;
wire n_34842;
wire n_34843;
wire n_34844;
wire n_34845;
wire n_34846;
wire n_34847;
wire n_34848;
wire n_34849;
wire n_34850;
wire n_34851;
wire n_34852;
wire n_34853;
wire n_34854;
wire n_34855;
wire n_34856;
wire n_34857;
wire n_34858;
wire n_34859;
wire n_34860;
wire n_34861;
wire n_34862;
wire n_34863;
wire n_34864;
wire n_34865;
wire n_34866;
wire n_34867;
wire n_34868;
wire n_34869;
wire n_34870;
wire n_34871;
wire n_34872;
wire n_34873;
wire n_34874;
wire n_34875;
wire n_34876;
wire n_34877;
wire n_34878;
wire n_34879;
wire n_34880;
wire n_34881;
wire n_34882;
wire n_34883;
wire n_34884;
wire n_34885;
wire n_34886;
wire n_34887;
wire n_34888;
wire n_34889;
wire n_34890;
wire n_34891;
wire n_34892;
wire n_34893;
wire n_34894;
wire n_34895;
wire n_34896;
wire n_34897;
wire n_34898;
wire n_34899;
wire n_34900;
wire n_34901;
wire n_34902;
wire n_34903;
wire n_34904;
wire n_34905;
wire n_34906;
wire n_34907;
wire n_34908;
wire n_34909;
wire n_34910;
wire n_34911;
wire n_34912;
wire n_34913;
wire n_34914;
wire n_34915;
wire n_34916;
wire n_34917;
wire n_34918;
wire n_34919;
wire n_34920;
wire n_34921;
wire n_34922;
wire n_34923;
wire n_34924;
wire n_34925;
wire n_34926;
wire n_34927;
wire n_34928;
wire n_34929;
wire n_34930;
wire n_34931;
wire n_34932;
wire n_34933;
wire n_34934;
wire n_34935;
wire n_34936;
wire n_34937;
wire n_34938;
wire n_34939;
wire n_34940;
wire n_34941;
wire n_34942;
wire n_34943;
wire n_34944;
wire n_34945;
wire n_34946;
wire n_34947;
wire n_34948;
wire n_34949;
wire n_34950;
wire n_34951;
wire n_34952;
wire n_34953;
wire n_34954;
wire n_34955;
wire n_34956;
wire n_34957;
wire n_34958;
wire n_34959;
wire n_34960;
wire n_34961;
wire n_34962;
wire n_34963;
wire n_34964;
wire n_34965;
wire n_34966;
wire n_34967;
wire n_34968;
wire n_34969;
wire n_34970;
wire n_34971;
wire n_34972;
wire n_34973;
wire n_34974;
wire n_34975;
wire n_34976;
wire n_34977;
wire n_34978;
wire n_34979;
wire n_34980;
wire n_34981;
wire n_34982;
wire n_34983;
wire n_34984;
wire n_34985;
wire n_34986;
wire n_34987;
wire n_34988;
wire n_34989;
wire n_34990;
wire n_34991;
wire n_34992;
wire n_34993;
wire n_34994;
wire n_34995;
wire n_34996;
wire n_34997;
wire n_34998;
wire n_34999;
wire n_35000;
wire n_35001;
wire n_35002;
wire n_35003;
wire n_35004;
wire n_35005;
wire n_35006;
wire n_35007;
wire n_35008;
wire n_35009;
wire n_35010;
wire n_35011;
wire n_35012;
wire n_35013;
wire n_35014;
wire n_35015;
wire n_35016;
wire n_35017;
wire n_35018;
wire n_35019;
wire n_35020;
wire n_35021;
wire n_35022;
wire n_35023;
wire n_35024;
wire n_35025;
wire n_35026;
wire n_35027;
wire n_35028;
wire n_35029;
wire n_35030;
wire n_35031;
wire n_35032;
wire n_35033;
wire n_35034;
wire n_35035;
wire n_35036;
wire n_35037;
wire n_35038;
wire n_35039;
wire n_35040;
wire n_35041;
wire n_35042;
wire n_35043;
wire n_35044;
wire n_35045;
wire n_35046;
wire n_35047;
wire n_35048;
wire n_35049;
wire n_35050;
wire n_35051;
wire n_35052;
wire n_35053;
wire n_35054;
wire n_35055;
wire n_35056;
wire n_35057;
wire n_35058;
wire n_35059;
wire n_35060;
wire n_35061;
wire n_35062;
wire n_35063;
wire n_35064;
wire n_35065;
wire n_35066;
wire n_35067;
wire n_35068;
wire n_35069;
wire n_35070;
wire n_35071;
wire n_35072;
wire n_35073;
wire n_35074;
wire n_35075;
wire n_35076;
wire n_35077;
wire n_35078;
wire n_35079;
wire n_35080;
wire n_35081;
wire n_35082;
wire n_35083;
wire n_35084;
wire n_35085;
wire n_35086;
wire n_35087;
wire n_35088;
wire n_35089;
wire n_35090;
wire n_35091;
wire n_35092;
wire n_35093;
wire n_35094;
wire n_35095;
wire n_35096;
wire n_35097;
wire n_35098;
wire n_35099;
wire n_35100;
wire n_35101;
wire n_35102;
wire n_35103;
wire n_35104;
wire n_35105;
wire n_35106;
wire n_35107;
wire n_35108;
wire n_35109;
wire n_35110;
wire n_35111;
wire n_35112;
wire n_35113;
wire n_35114;
wire n_35115;
wire n_35116;
wire n_35117;
wire n_35118;
wire n_35119;
wire n_35120;
wire n_35121;
wire n_35122;
wire n_35123;
wire n_35124;
wire n_35125;
wire n_35126;
wire n_35127;
wire n_35128;
wire n_35129;
wire n_35130;
wire n_35131;
wire n_35132;
wire n_35133;
wire n_35134;
wire n_35135;
wire n_35136;
wire n_35137;
wire n_35138;
wire n_35139;
wire n_35140;
wire n_35141;
wire n_35142;
wire n_35143;
wire n_35144;
wire n_35145;
wire n_35146;
wire n_35147;
wire n_35148;
wire n_35149;
wire n_35150;
wire n_35151;
wire n_35152;
wire n_35153;
wire n_35154;
wire n_35155;
wire n_35156;
wire n_35157;
wire n_35158;
wire n_35159;
wire n_35160;
wire n_35161;
wire n_35162;
wire n_35163;
wire n_35164;
wire n_35165;
wire n_35166;
wire n_35167;
wire n_35168;
wire n_35169;
wire n_35170;
wire n_35171;
wire n_35172;
wire n_35173;
wire n_35174;
wire n_35175;
wire n_35176;
wire n_35177;
wire n_35178;
wire n_35179;
wire n_35180;
wire n_35181;
wire n_35182;
wire n_35183;
wire n_35184;
wire n_35185;
wire n_35186;
wire n_35187;
wire n_35188;
wire n_35189;
wire n_35190;
wire n_35191;
wire n_35192;
wire n_35193;
wire n_35194;
wire n_35195;
wire n_35196;
wire n_35197;
wire n_35198;
wire n_35199;
wire n_35200;
wire n_35201;
wire n_35202;
wire n_35203;
wire n_35204;
wire n_35205;
wire n_35206;
wire n_35207;
wire n_35208;
wire n_35209;
wire n_35210;
wire n_35211;
wire n_35212;
wire n_35213;
wire n_35214;
wire n_35215;
wire n_35216;
wire n_35217;
wire n_35218;
wire n_35219;
wire n_35220;
wire n_35221;
wire n_35222;
wire n_35223;
wire n_35224;
wire n_35225;
wire n_35226;
wire n_35227;
wire n_35228;
wire n_35229;
wire n_35230;
wire n_35231;
wire n_35232;
wire n_35233;
wire n_35234;
wire n_35235;
wire n_35236;
wire n_35237;
wire n_35238;
wire n_35239;
wire n_35240;
wire n_35241;
wire n_35242;
wire n_35243;
wire n_35244;
wire n_35245;
wire n_35246;
wire n_35247;
wire n_35248;
wire n_35249;
wire n_35250;
wire n_35251;
wire n_35252;
wire n_35253;
wire n_35254;
wire n_35255;
wire n_35256;
wire n_35257;
wire n_35258;
wire n_35259;
wire n_35260;
wire n_35261;
wire n_35262;
wire n_35263;
wire n_35264;
wire n_35265;
wire n_35266;
wire n_35267;
wire n_35268;
wire n_35269;
wire n_35270;
wire n_35271;
wire n_35272;
wire n_35273;
wire n_35274;
wire n_35275;
wire n_35276;
wire n_35277;
wire n_35278;
wire n_35279;
wire n_35280;
wire n_35281;
wire n_35282;
wire n_35283;
wire n_35284;
wire n_35285;
wire n_35286;
wire n_35287;
wire n_35288;
wire n_35289;
wire n_35290;
wire n_35291;
wire n_35292;
wire n_35293;
wire n_35294;
wire n_35295;
wire n_35296;
wire n_35297;
wire n_35298;
wire n_35299;
wire n_35300;
wire n_35301;
wire n_35302;
wire n_35303;
wire n_35304;
wire n_35305;
wire n_35306;
wire n_35307;
wire n_35308;
wire n_35309;
wire n_35310;
wire n_35311;
wire n_35312;
wire n_35313;
wire n_35314;
wire n_35315;
wire n_35316;
wire n_35317;
wire n_35318;
wire n_35319;
wire n_35320;
wire n_35321;
wire n_35322;
wire n_35323;
wire n_35324;
wire n_35325;
wire n_35326;
wire n_35327;
wire n_35328;
wire n_35329;
wire n_35330;
wire n_35331;
wire n_35332;
wire n_35333;
wire n_35334;
wire n_35335;
wire n_35336;
wire n_35337;
wire n_35338;
wire n_35339;
wire n_35340;
wire n_35341;
wire n_35342;
wire n_35343;
wire n_35344;
wire n_35345;
wire n_35346;
wire n_35347;
wire n_35348;
wire n_35349;
wire n_35350;
wire n_35351;
wire n_35352;
wire n_35353;
wire n_35354;
wire n_35355;
wire n_35356;
wire n_35357;
wire n_35358;
wire n_35359;
wire n_35360;
wire n_35361;
wire n_35362;
wire n_35363;
wire n_35364;
wire n_35365;
wire n_35366;
wire n_35367;
wire n_35368;
wire n_35369;
wire n_35370;
wire n_35371;
wire n_35372;
wire n_35373;
wire n_35374;
wire n_35375;
wire n_35376;
wire n_35377;
wire n_35378;
wire n_35379;
wire n_35380;
wire n_35381;
wire n_35382;
wire n_35383;
wire n_35384;
wire n_35385;
wire n_35386;
wire n_35387;
wire n_35388;
wire n_35389;
wire n_35390;
wire n_35391;
wire n_35392;
wire n_35393;
wire n_35394;
wire n_35395;
wire n_35396;
wire n_35397;
wire n_35398;
wire n_35399;
wire n_35400;
wire n_35401;
wire n_35402;
wire n_35403;
wire n_35404;
wire n_35405;
wire n_35406;
wire n_35407;
wire n_35408;
wire n_35409;
wire n_35410;
wire n_35411;
wire n_35412;
wire n_35413;
wire n_35414;
wire n_35415;
wire n_35416;
wire n_35417;
wire n_35418;
wire n_35419;
wire n_35420;
wire n_35421;
wire n_35422;
wire n_35423;
wire n_35424;
wire n_35425;
wire n_35426;
wire n_35427;
wire n_35428;
wire n_35429;
wire n_35430;
wire n_35431;
wire n_35432;
wire n_35433;
wire n_35434;
wire n_35435;
wire n_35436;
wire n_35437;
wire n_35438;
wire n_35439;
wire n_35440;
wire n_35441;
wire n_35442;
wire n_35443;
wire n_35444;
wire n_35445;
wire n_35446;
wire n_35447;
wire n_35448;
wire n_35449;
wire n_35450;
wire n_35451;
wire n_35452;
wire n_35453;
wire n_35454;
wire n_35455;
wire n_35456;
wire n_35457;
wire n_35458;
wire n_35459;
wire n_35460;
wire n_35461;
wire n_35462;
wire n_35463;
wire n_35464;
wire n_35465;
wire n_35466;
wire n_35467;
wire n_35468;
wire n_35469;
wire n_35470;
wire n_35471;
wire n_35472;
wire n_35473;
wire n_35474;
wire n_35475;
wire n_35476;
wire n_35477;
wire n_35478;
wire n_35479;
wire n_35480;
wire n_35481;
wire n_35482;
wire n_35483;
wire n_35484;
wire n_35485;
wire n_35486;
wire n_35487;
wire n_35488;
wire n_35489;
wire n_35490;
wire n_35491;
wire n_35492;
wire n_35493;
wire n_35494;
wire n_35495;
wire n_35496;
wire n_35497;
wire n_35498;
wire n_35499;
wire n_35500;
wire n_35501;
wire n_35502;
wire n_35503;
wire n_35504;
wire n_35505;
wire n_35506;
wire n_35507;
wire n_35508;
wire n_35509;
wire n_35510;
wire n_35511;
wire n_35512;
wire n_35513;
wire n_35514;
wire n_35515;
wire n_35516;
wire n_35517;
wire n_35518;
wire n_35519;
wire n_35520;
wire n_35521;
wire n_35522;
wire n_35523;
wire n_35524;
wire n_35525;
wire n_35526;
wire n_35527;
wire n_35528;
wire n_35529;
wire n_35530;
wire n_35531;
wire n_35532;
wire n_35533;
wire n_35534;
wire n_35535;
wire n_35536;
wire n_35537;
wire n_35538;
wire n_35539;
wire n_35540;
wire n_35541;
wire n_35542;
wire n_35543;
wire n_35544;
wire n_35545;
wire n_35546;
wire n_35547;
wire n_35548;
wire n_35549;
wire n_35550;
wire n_35551;
wire n_35552;
wire n_35553;
wire n_35554;
wire n_35555;
wire n_35556;
wire n_35557;
wire n_35558;
wire n_35559;
wire n_35560;
wire n_35561;
wire n_35562;
wire n_35563;
wire n_35564;
wire n_35565;
wire n_35566;
wire n_35567;
wire n_35568;
wire n_35569;
wire n_35570;
wire n_35571;
wire n_35572;
wire n_35573;
wire n_35574;
wire n_35575;
wire n_35576;
wire n_35577;
wire n_35578;
wire n_35579;
wire n_35580;
wire n_35581;
wire n_35582;
wire n_35583;
wire n_35584;
wire n_35585;
wire n_35586;
wire n_35587;
wire n_35588;
wire n_35589;
wire n_35590;
wire n_35591;
wire n_35592;
wire n_35593;
wire n_35594;
wire n_35595;
wire n_35596;
wire n_35597;
wire n_35598;
wire n_35599;
wire n_35600;
wire n_35601;
wire n_35602;
wire n_35603;
wire n_35604;
wire n_35605;
wire n_35606;
wire n_35607;
wire n_35608;
wire n_35609;
wire n_35610;
wire n_35611;
wire n_35612;
wire n_35613;
wire n_35614;
wire n_35615;
wire n_35616;
wire n_35617;
wire n_35618;
wire n_35619;
wire n_35620;
wire n_35621;
wire n_35622;
wire n_35623;
wire n_35624;
wire n_35625;
wire n_35626;
wire n_35627;
wire n_35628;
wire n_35629;
wire n_35630;
wire n_35631;
wire n_35632;
wire n_35633;
wire n_35634;
wire n_35635;
wire n_35636;
wire n_35637;
wire n_35638;
wire n_35639;
wire n_35640;
wire n_35641;
wire n_35642;
wire n_35643;
wire n_35644;
wire n_35645;
wire n_35646;
wire n_35647;
wire n_35648;
wire n_35649;
wire n_35650;
wire n_35651;
wire n_35652;
wire n_35653;
wire n_35654;
wire n_35655;
wire n_35656;
wire n_35657;
wire n_35658;
wire n_35659;
wire n_35660;
wire n_35661;
wire n_35662;
wire n_35663;
wire n_35664;
wire n_35665;
wire n_35666;
wire n_35667;
wire n_35668;
wire n_35669;
wire n_35670;
wire n_35671;
wire n_35672;
wire n_35673;
wire n_35674;
wire n_35675;
wire n_35676;
wire n_35677;
wire n_35678;
wire n_35679;
wire n_35680;
wire n_35681;
wire n_35682;
wire n_35683;
wire n_35684;
wire n_35685;
wire n_35686;
wire n_35687;
wire n_35688;
wire n_35689;
wire n_35690;
wire n_35691;
wire n_35692;
wire n_35693;
wire n_35694;
wire n_35695;
wire n_35696;
wire n_35697;
wire n_35698;
wire n_35699;
wire n_35700;
wire n_35701;
wire n_35702;
wire n_35703;
wire n_35704;
wire n_35705;
wire n_35706;
wire n_35707;
wire n_35708;
wire n_35709;
wire n_35710;
wire n_35711;
wire n_35712;
wire n_35713;
wire n_35714;
wire n_35715;
wire n_35716;
wire n_35717;
wire n_35718;
wire n_35719;
wire n_35720;
wire n_35721;
wire n_35722;
wire n_35723;
wire n_35724;
wire n_35725;
wire n_35726;
wire n_35727;
wire n_35728;
wire n_35729;
wire n_35730;
wire n_35731;
wire n_35732;
wire n_35733;
wire n_35734;
wire n_35735;
wire n_35736;
wire n_35737;
wire n_35738;
wire n_35739;
wire n_35740;
wire n_35741;
wire n_35742;
wire n_35743;
wire n_35744;
wire n_35745;
wire n_35746;
wire n_35747;
wire n_35748;
wire n_35749;
wire n_35750;
wire n_35751;
wire n_35752;
wire n_35753;
wire n_35754;
wire n_35755;
wire n_35756;
wire n_35757;
wire n_35758;
wire n_35759;
wire n_35760;
wire n_35761;
wire n_35762;
wire n_35763;
wire n_35764;
wire n_35765;
wire n_35766;
wire n_35767;
wire n_35768;
wire n_35769;
wire n_35770;
wire n_35771;
wire n_35772;
wire n_35773;
wire n_35774;
wire n_35775;
wire n_35776;
wire n_35777;
wire n_35778;
wire n_35779;
wire n_35780;
wire n_35781;
wire n_35782;
wire n_35783;
wire n_35784;
wire n_35785;
wire n_35786;
wire n_35787;
wire n_35788;
wire n_35789;
wire n_35790;
wire n_35791;
wire n_35792;
wire n_35793;
wire n_35794;
wire n_35795;
wire n_35796;
wire n_35797;
wire n_35798;
wire n_35799;
wire n_35800;
wire n_35801;
wire n_35802;
wire n_35803;
wire n_35804;
wire n_35805;
wire n_35806;
wire n_35807;
wire n_35808;
wire n_35809;
wire n_35810;
wire n_35811;
wire n_35812;
wire n_35813;
wire n_35814;
wire n_35815;
wire n_35816;
wire n_35817;
wire n_35818;
wire n_35819;
wire n_35820;
wire n_35821;
wire n_35822;
wire n_35823;
wire n_35824;
wire n_35825;
wire n_35826;
wire n_35827;
wire n_35828;
wire n_35829;
wire n_35830;
wire n_35831;
wire n_35832;
wire n_35833;
wire n_35834;
wire n_35835;
wire n_35836;
wire n_35837;
wire n_35838;
wire n_35839;
wire n_35840;
wire n_35841;
wire n_35842;
wire n_35843;
wire n_35844;
wire n_35845;
wire n_35846;
wire n_35847;
wire n_35848;
wire n_35849;
wire n_35850;
wire n_35851;
wire n_35852;
wire n_35853;
wire n_35854;
wire n_35855;
wire n_35856;
wire n_35857;
wire n_35858;
wire n_35859;
wire n_35860;
wire n_35861;
wire n_35862;
wire n_35863;
wire n_35864;
wire n_35865;
wire n_35866;
wire n_35867;
wire n_35868;
wire n_35869;
wire n_35870;
wire n_35871;
wire n_35872;
wire n_35873;
wire n_35874;
wire n_35875;
wire n_35876;
wire n_35877;
wire n_35878;
wire n_35879;
wire n_35880;
wire n_35881;
wire n_35882;
wire n_35883;
wire n_35884;
wire n_35885;
wire n_35886;
wire n_35887;
wire n_35888;
wire n_35889;
wire n_35890;
wire n_35891;
wire n_35892;
wire n_35893;
wire n_35894;
wire n_35895;
wire n_35896;
wire n_35897;
wire n_35898;
wire n_35899;
wire n_35900;
wire n_35901;
wire n_35902;
wire n_35903;
wire n_35904;
wire n_35905;
wire n_35906;
wire n_35907;
wire n_35908;
wire n_35909;
wire n_35910;
wire n_35911;
wire n_35912;
wire n_35913;
wire n_35914;
wire n_35915;
wire n_35916;
wire n_35917;
wire n_35918;
wire n_35919;
wire n_35920;
wire n_35921;
wire n_35922;
wire n_35923;
wire n_35924;
wire n_35925;
wire n_35926;
wire n_35927;
wire n_35928;
wire n_35929;
wire n_35930;
wire n_35931;
wire n_35932;
wire n_35933;
wire n_35934;
wire n_35935;
wire n_35936;
wire n_35937;
wire n_35938;
wire n_35939;
wire n_35940;
wire n_35941;
wire n_35942;
wire n_35943;
wire n_35944;
wire n_35945;
wire n_35946;
wire n_35947;
wire n_35948;
wire n_35949;
wire n_35950;
wire n_35951;
wire n_35952;
wire n_35953;
wire n_35954;
wire n_35955;
wire n_35956;
wire n_35957;
wire n_35958;
wire n_35959;
wire n_35960;
wire n_35961;
wire n_35962;
wire n_35963;
wire n_35964;
wire n_35965;
wire n_35966;
wire n_35967;
wire n_35968;
wire n_35969;
wire n_35970;
wire n_35971;
wire n_35972;
wire n_35973;
wire n_35974;
wire n_35975;
wire n_35976;
wire n_35977;
wire n_35978;
wire n_35979;
wire n_35980;
wire n_35981;
wire n_35982;
wire n_35983;
wire n_35984;
wire n_35985;
wire n_35986;
wire n_35987;
wire n_35988;
wire n_35989;
wire n_35990;
wire n_35991;
wire n_35992;
wire n_35993;
wire n_35994;
wire n_35995;
wire n_35996;
wire n_35997;
wire n_35998;
wire n_35999;
wire n_36000;
wire n_36001;
wire n_36002;
wire n_36003;
wire n_36004;
wire n_36005;
wire n_36006;
wire n_36007;
wire n_36008;
wire n_36009;
wire n_36010;
wire n_36011;
wire n_36012;
wire n_36013;
wire n_36014;
wire n_36015;
wire n_36016;
wire n_36017;
wire n_36018;
wire n_36019;
wire n_36020;
wire n_36021;
wire n_36022;
wire n_36023;
wire n_36024;
wire n_36025;
wire n_36026;
wire n_36027;
wire n_36028;
wire n_36029;
wire n_36030;
wire n_36031;
wire n_36032;
wire n_36033;
wire n_36034;
wire n_36035;
wire n_36036;
wire n_36037;
wire n_36038;
wire n_36039;
wire n_36040;
wire n_36041;
wire n_36042;
wire n_36043;
wire n_36044;
wire n_36045;
wire n_36046;
wire n_36047;
wire n_36048;
wire n_36049;
wire n_36050;
wire n_36051;
wire n_36052;
wire n_36053;
wire n_36054;
wire n_36055;
wire n_36056;
wire n_36057;
wire n_36058;
wire n_36059;
wire n_36060;
wire n_36061;
wire n_36062;
wire n_36063;
wire n_36064;
wire n_36065;
wire n_36066;
wire n_36067;
wire n_36068;
wire n_36069;
wire n_36070;
wire n_36071;
wire n_36072;
wire n_36073;
wire n_36074;
wire n_36075;
wire n_36076;
wire n_36077;
wire n_36078;
wire n_36079;
wire n_36080;
wire n_36081;
wire n_36082;
wire n_36083;
wire n_36084;
wire n_36085;
wire n_36086;
wire n_36087;
wire n_36088;
wire n_36089;
wire n_36090;
wire n_36091;
wire n_36092;
wire n_36093;
wire n_36094;
wire n_36095;
wire n_36096;
wire n_36097;
wire n_36098;
wire n_36099;
wire n_36100;
wire n_36101;
wire n_36102;
wire n_36103;
wire n_36104;
wire n_36105;
wire n_36106;
wire n_36107;
wire n_36108;
wire n_36109;
wire n_36110;
wire n_36111;
wire n_36112;
wire n_36113;
wire n_36114;
wire n_36115;
wire n_36116;
wire n_36117;
wire n_36118;
wire n_36119;
wire n_36120;
wire n_36121;
wire n_36122;
wire n_36123;
wire n_36124;
wire n_36125;
wire n_36126;
wire n_36127;
wire n_36128;
wire n_36129;
wire n_36130;
wire n_36131;
wire n_36132;
wire n_36133;
wire n_36134;
wire n_36135;
wire n_36136;
wire n_36137;
wire n_36138;
wire n_36139;
wire n_36140;
wire n_36141;
wire n_36142;
wire n_36143;
wire n_36144;
wire n_36145;
wire n_36146;
wire n_36147;
wire n_36148;
wire n_36149;
wire n_36150;
wire n_36151;
wire n_36152;
wire n_36153;
wire n_36154;
wire n_36155;
wire n_36156;
wire n_36157;
wire n_36158;
wire n_36159;
wire n_36160;
wire n_36161;
wire n_36162;
wire n_36163;
wire n_36164;
wire n_36165;
wire n_36166;
wire n_36167;
wire n_36168;
wire n_36169;
wire n_36170;
wire n_36171;
wire n_36172;
wire n_36173;
wire n_36174;
wire n_36175;
wire n_36176;
wire n_36177;
wire n_36178;
wire n_36179;
wire n_36180;
wire n_36181;
wire n_36182;
wire n_36183;
wire n_36184;
wire n_36185;
wire n_36186;
wire n_36187;
wire n_36188;
wire n_36189;
wire n_36190;
wire n_36191;
wire n_36192;
wire n_36193;
wire n_36194;
wire n_36195;
wire n_36196;
wire n_36197;
wire n_36198;
wire n_36199;
wire n_36200;
wire n_36201;
wire n_36202;
wire n_36203;
wire n_36204;
wire n_36205;
wire n_36206;
wire n_36207;
wire n_36208;
wire n_36209;
wire n_36210;
wire n_36211;
wire n_36212;
wire n_36213;
wire n_36214;
wire n_36215;
wire n_36216;
wire n_36217;
wire n_36218;
wire n_36219;
wire n_36220;
wire n_36221;
wire n_36222;
wire n_36223;
wire n_36224;
wire n_36225;
wire n_36226;
wire n_36227;
wire n_36228;
wire n_36229;
wire n_36230;
wire n_36231;
wire n_36232;
wire n_36233;
wire n_36234;
wire n_36235;
wire n_36236;
wire n_36237;
wire n_36238;
wire n_36239;
wire n_36240;
wire n_36241;
wire n_36242;
wire n_36243;
wire n_36244;
wire n_36245;
wire n_36246;
wire n_36247;
wire n_36248;
wire n_36249;
wire n_36250;
wire n_36251;
wire n_36252;
wire n_36253;
wire n_36254;
wire n_36255;
wire n_36256;
wire n_36257;
wire n_36258;
wire n_36259;
wire n_36260;
wire n_36261;
wire n_36262;
wire n_36263;
wire n_36264;
wire n_36265;
wire n_36266;
wire n_36267;
wire n_36268;
wire n_36269;
wire n_36270;
wire n_36271;
wire n_36272;
wire n_36273;
wire n_36274;
wire n_36275;
wire n_36276;
wire n_36277;
wire n_36278;
wire n_36279;
wire n_36280;
wire n_36281;
wire n_36282;
wire n_36283;
wire n_36284;
wire n_36285;
wire n_36286;
wire n_36287;
wire n_36288;
wire n_36289;
wire n_36290;
wire n_36291;
wire n_36292;
wire n_36293;
wire n_36294;
wire n_36295;
wire n_36296;
wire n_36297;
wire n_36298;
wire n_36299;
wire n_36300;
wire n_36301;
wire n_36302;
wire n_36303;
wire n_36304;
wire n_36305;
wire n_36306;
wire n_36307;
wire n_36308;
wire n_36309;
wire n_36310;
wire n_36311;
wire n_36312;
wire n_36313;
wire n_36314;
wire n_36315;
wire n_36316;
wire n_36317;
wire n_36318;
wire n_36319;
wire n_36320;
wire n_36321;
wire n_36322;
wire n_36323;
wire n_36324;
wire n_36325;
wire n_36326;
wire n_36327;
wire n_36328;
wire n_36329;
wire n_36330;
wire n_36331;
wire n_36332;
wire n_36333;
wire n_36334;
wire n_36335;
wire n_36336;
wire n_36337;
wire n_36338;
wire n_36339;
wire n_36340;
wire n_36341;
wire n_36342;
wire n_36343;
wire n_36344;
wire n_36345;
wire n_36346;
wire n_36347;
wire n_36348;
wire n_36349;
wire n_36350;
wire n_36351;
wire n_36352;
wire n_36353;
wire n_36354;
wire n_36355;
wire n_36356;
wire n_36357;
wire n_36358;
wire n_36359;
wire n_36360;
wire n_36361;
wire n_36362;
wire n_36363;
wire n_36364;
wire n_36365;
wire n_36366;
wire n_36367;
wire n_36368;
wire n_36369;
wire n_36370;
wire n_36371;
wire n_36372;
wire n_36373;
wire n_36374;
wire n_36375;
wire n_36376;
wire n_36377;
wire n_36378;
wire n_36379;
wire n_36380;
wire n_36381;
wire n_36382;
wire n_36383;
wire n_36384;
wire n_36385;
wire n_36386;
wire n_36387;
wire n_36388;
wire n_36389;
wire n_36390;
wire n_36391;
wire n_36392;
wire n_36393;
wire n_36394;
wire n_36395;
wire n_36396;
wire n_36397;
wire n_36398;
wire n_36399;
wire n_36400;
wire n_36401;
wire n_36402;
wire n_36403;
wire n_36404;
wire n_36405;
wire n_36406;
wire n_36407;
wire n_36408;
wire n_36409;
wire n_36410;
wire n_36411;
wire n_36412;
wire n_36413;
wire n_36414;
wire n_36415;
wire n_36416;
wire n_36417;
wire n_36418;
wire n_36419;
wire n_36420;
wire n_36421;
wire n_36422;
wire n_36423;
wire n_36424;
wire n_36425;
wire n_36426;
wire n_36427;
wire n_36428;
wire n_36429;
wire n_36430;
wire n_36431;
wire n_36432;
wire n_36433;
wire n_36434;
wire n_36435;
wire n_36436;
wire n_36437;
wire n_36438;
wire n_36439;
wire n_36440;
wire n_36441;
wire n_36442;
wire n_36443;
wire n_36444;
wire n_36445;
wire n_36446;
wire n_36447;
wire n_36448;
wire n_36449;
wire n_36450;
wire n_36451;
wire n_36452;
wire n_36453;
wire n_36454;
wire n_36455;
wire n_36456;
wire n_36457;
wire n_36458;
wire n_36459;
wire n_36460;
wire n_36461;
wire n_36462;
wire n_36463;
wire n_36464;
wire n_36465;
wire n_36466;
wire n_36467;
wire n_36468;
wire n_36469;
wire n_36470;
wire n_36471;
wire n_36472;
wire n_36473;
wire n_36474;
wire n_36475;
wire n_36476;
wire n_36477;
wire n_36478;
wire n_36479;
wire n_36480;
wire n_36481;
wire n_36482;
wire n_36483;
wire n_36484;
wire n_36485;
wire n_36486;
wire n_36487;
wire n_36488;
wire n_36489;
wire n_36490;
wire n_36491;
wire n_36492;
wire n_36493;
wire n_36494;
wire n_36495;
wire n_36496;
wire n_36497;
wire n_36498;
wire n_36499;
wire n_36500;
wire n_36501;
wire n_36502;
wire n_36503;
wire n_36504;
wire n_36505;
wire n_36506;
wire n_36507;
wire n_36508;
wire n_36509;
wire n_36510;
wire n_36511;
wire n_36512;
wire n_36513;
wire n_36514;
wire n_36515;
wire n_36516;
wire n_36517;
wire n_36518;
wire n_36519;
wire n_36520;
wire n_36521;
wire n_36522;
wire n_36523;
wire n_36524;
wire n_36525;
wire n_36526;
wire n_36527;
wire n_36528;
wire n_36529;
wire n_36530;
wire n_36531;
wire n_36532;
wire n_36533;
wire n_36534;
wire n_36535;
wire n_36536;
wire n_36537;
wire n_36538;
wire n_36539;
wire n_36540;
wire n_36541;
wire n_36542;
wire n_36543;
wire n_36544;
wire n_36545;
wire n_36546;
wire n_36547;
wire n_36548;
wire n_36549;
wire n_36550;
wire n_36551;
wire n_36552;
wire n_36553;
wire n_36554;
wire n_36555;
wire n_36556;
wire n_36557;
wire n_36558;
wire n_36559;
wire n_36560;
wire n_36561;
wire n_36562;
wire n_36563;
wire n_36564;
wire n_36565;
wire n_36566;
wire n_36567;
wire n_36568;
wire n_36569;
wire n_36570;
wire n_36571;
wire n_36572;
wire n_36573;
wire n_36574;
wire n_36575;
wire n_36576;
wire n_36577;
wire n_36578;
wire n_36579;
wire n_36580;
wire n_36581;
wire n_36582;
wire n_36583;
wire n_36584;
wire n_36585;
wire n_36586;
wire n_36587;
wire n_36588;
wire n_36589;
wire n_36590;
wire n_36591;
wire n_36592;
wire n_36593;
wire n_36594;
wire n_36595;
wire n_36596;
wire n_36597;
wire n_36598;
wire n_36599;
wire n_36600;
wire n_36601;
wire n_36602;
wire n_36603;
wire n_36604;
wire n_36605;
wire n_36606;
wire n_36607;
wire n_36608;
wire n_36609;
wire n_36610;
wire n_36611;
wire n_36612;
wire n_36613;
wire n_36614;
wire n_36615;
wire n_36616;
wire n_36617;
wire n_36618;
wire n_36619;
wire n_36620;
wire n_36621;
wire n_36622;
wire n_36623;
wire n_36624;
wire n_36625;
wire n_36626;
wire n_36627;
wire n_36628;
wire n_36629;
wire n_36630;
wire n_36631;
wire n_36632;
wire n_36633;
wire n_36634;
wire n_36635;
wire n_36636;
wire n_36637;
wire n_36638;
wire n_36639;
wire n_36640;
wire n_36641;
wire n_36642;
wire n_36643;
wire n_36644;
wire n_36645;
wire n_36646;
wire n_36647;
wire n_36648;
wire n_36649;
wire n_36650;
wire n_36651;
wire n_36652;
wire n_36653;
wire n_36654;
wire n_36655;
wire n_36656;
wire n_36657;
wire n_36658;
wire n_36659;
wire n_36660;
wire n_36661;
wire n_36662;
wire n_36663;
wire n_36664;
wire n_36665;
wire n_36666;
wire n_36667;
wire n_36668;
wire n_36669;
wire n_36670;
wire n_36671;
wire n_36672;
wire n_36673;
wire n_36674;
wire n_36675;
wire n_36676;
wire n_36677;
wire n_36678;
wire n_36679;
wire n_36680;
wire n_36681;
wire n_36682;
wire n_36683;
wire n_36684;
wire n_36685;
wire n_36686;
wire n_36687;
wire n_36688;
wire n_36689;
wire n_36690;
wire n_36691;
wire n_36692;
wire n_36693;
wire n_36694;
wire n_36695;
wire n_36696;
wire n_36697;
wire n_36698;
wire n_36699;
wire n_36700;
wire n_36701;
wire n_36702;
wire n_36703;
wire n_36704;
wire n_36705;
wire n_36706;
wire n_36707;
wire n_36708;
wire n_36709;
wire n_36710;
wire n_36711;
wire n_36712;
wire n_36713;
wire n_36714;
wire n_36715;
wire n_36716;
wire n_36717;
wire n_36718;
wire n_36719;
wire n_36720;
wire n_36721;
wire n_36722;
wire n_36723;
wire n_36724;
wire n_36725;
wire n_36726;
wire n_36727;
wire n_36728;
wire n_36729;
wire n_36730;
wire n_36731;
wire n_36732;
wire n_36733;
wire n_36734;
wire n_36735;
wire n_36736;
wire n_36737;
wire n_36738;
wire n_36739;
wire n_36740;
wire n_36741;
wire n_36742;
wire n_36743;
wire n_36744;
wire n_36745;
wire n_36746;
wire n_36747;
wire n_36748;
wire n_36749;
wire n_36750;
wire n_36751;
wire n_36752;
wire n_36753;
wire n_36754;
wire n_36755;
wire n_36756;
wire n_36757;
wire n_36758;
wire n_36759;
wire n_36760;
wire n_36761;
wire n_36762;
wire n_36763;
wire n_36764;
wire n_36765;
wire n_36766;
wire n_36767;
wire n_36768;
wire n_36769;
wire n_36770;
wire n_36771;
wire n_36772;
wire n_36773;
wire n_36774;
wire n_36775;
wire n_36776;
wire n_36777;
wire n_36778;
wire n_36779;
wire n_36780;
wire n_36781;
wire n_36782;
wire n_36783;
wire n_36784;
wire n_36785;
wire n_36786;
wire n_36787;
wire n_36788;
wire n_36789;
wire n_36790;
wire n_36791;
wire n_36792;
wire n_36793;
wire n_36794;
wire n_36795;
wire n_36796;
wire n_36797;
wire n_36798;
wire n_36799;
wire n_36800;
wire n_36801;
wire n_36802;
wire n_36803;
wire n_36804;
wire n_36805;
wire n_36806;
wire n_36807;
wire n_36808;
wire n_36809;
wire n_36810;
wire n_36811;
wire n_36812;
wire n_36813;
wire n_36814;
wire n_36815;
wire n_36816;
wire n_36817;
wire n_36818;
wire n_36819;
wire n_36820;
wire n_36821;
wire n_36822;
wire n_36823;
wire n_36824;
wire n_36825;
wire n_36826;
wire n_36827;
wire n_36828;
wire n_36829;
wire n_36830;
wire n_36831;
wire n_36832;
wire n_36833;
wire n_36834;
wire n_36835;
wire n_36836;
wire n_36837;
wire n_36838;
wire n_36839;
wire n_36840;
wire n_36841;
wire n_36842;
wire n_36843;
wire n_36844;
wire n_36845;
wire n_36846;
wire n_36847;
wire n_36848;
wire n_36849;
wire n_36850;
wire n_36851;
wire n_36852;
wire n_36853;
wire n_36854;
wire n_36855;
wire n_36856;
wire n_36857;
wire n_36858;
wire n_36859;
wire n_36860;
wire n_36861;
wire n_36862;
wire n_36863;
wire n_36864;
wire n_36865;
wire n_36866;
wire n_36867;
wire n_36868;
wire n_36869;
wire n_36870;
wire n_36871;
wire n_36872;
wire n_36873;
wire n_36874;
wire n_36875;
wire n_36876;
wire n_36877;
wire n_36878;
wire n_36879;
wire n_36880;
wire n_36881;
wire n_36882;
wire n_36883;
wire n_36884;
wire n_36885;
wire n_36886;
wire n_36887;
wire n_36888;
wire n_36889;
wire n_36890;
wire n_36891;
wire n_36892;
wire n_36893;
wire n_36894;
wire n_36895;
wire n_36896;
wire n_36897;
wire n_36898;
wire n_36899;
wire n_36900;
wire n_36901;
wire n_36902;
wire n_36903;
wire n_36904;
wire n_36905;
wire n_36906;
wire n_36907;
wire n_36908;
wire n_36909;
wire n_36910;
wire n_36911;
wire n_36912;
wire n_36913;
wire n_36914;
wire n_36915;
wire n_36916;
wire n_36917;
wire n_36918;
wire n_36919;
wire n_36920;
wire n_36921;
wire n_36922;
wire n_36923;
wire n_36924;
wire n_36925;
wire n_36926;
wire n_36927;
wire n_36928;
wire n_36929;
wire n_36930;
wire n_36931;
wire n_36932;
wire n_36933;
wire n_36934;
wire n_36935;
wire n_36936;
wire n_36937;
wire n_36938;
wire n_36939;
wire n_36940;
wire n_36941;
wire n_36942;
wire n_36943;
wire n_36944;
wire n_36945;
wire n_36946;
wire n_36947;
wire n_36948;
wire n_36949;
wire n_36950;
wire n_36951;
wire n_36952;
wire n_36953;
wire n_36954;
wire n_36955;
wire n_36956;
wire n_36957;
wire n_36958;
wire n_36959;
wire n_36960;
wire n_36961;
wire n_36962;
wire n_36963;
wire n_36964;
wire n_36965;
wire n_36966;
wire n_36967;
wire n_36968;
wire n_36969;
wire n_36970;
wire n_36971;
wire n_36972;
wire n_36973;
wire n_36974;
wire n_36975;
wire n_36976;
wire n_36977;
wire n_36978;
wire n_36979;
wire n_36980;
wire n_36981;
wire n_36982;
wire n_36983;
wire n_36984;
wire n_36985;
wire n_36986;
wire n_36987;
wire n_36988;
wire n_36989;
wire n_36990;
wire n_36991;
wire n_36992;
wire n_36993;
wire n_36994;
wire n_36995;
wire n_36996;
wire n_36997;
wire n_36998;
wire n_36999;
wire n_37000;
wire n_37001;
wire n_37002;
wire n_37003;
wire n_37004;
wire n_37005;
wire n_37006;
wire n_37007;
wire n_37008;
wire n_37009;
wire n_37010;
wire n_37011;
wire n_37012;
wire n_37013;
wire n_37014;
wire n_37015;
wire n_37016;
wire n_37017;
wire n_37018;
wire n_37019;
wire n_37020;
wire n_37021;
wire n_37022;
wire n_37023;
wire n_37024;
wire n_37025;
wire n_37026;
wire n_37027;
wire n_37028;
wire n_37029;
wire n_37030;
wire n_37031;
wire n_37032;
wire n_37033;
wire n_37034;
wire n_37035;
wire n_37036;
wire n_37037;
wire n_37038;
wire n_37039;
wire n_37040;
wire n_37041;
wire n_37042;
wire n_37043;
wire n_37044;
wire n_37045;
wire n_37046;
wire n_37047;
wire n_37048;
wire n_37049;
wire n_37050;
wire n_37051;
wire n_37052;
wire n_37053;
wire n_37054;
wire n_37055;
wire n_37056;
wire n_37057;
wire n_37058;
wire n_37059;
wire n_37060;
wire n_37061;
wire n_37062;
wire n_37063;
wire n_37064;
wire n_37065;
wire n_37066;
wire n_37067;
wire n_37068;
wire n_37069;
wire n_37070;
wire n_37071;
wire n_37072;
wire n_37073;
wire n_37074;
wire n_37075;
wire n_37076;
wire n_37077;
wire n_37078;
wire n_37079;
wire n_37080;
wire n_37081;
wire n_37082;
wire n_37083;
wire n_37084;
wire n_37085;
wire n_37086;
wire n_37087;
wire n_37088;
wire n_37089;
wire n_37090;
wire n_37091;
wire n_37092;
wire n_37093;
wire n_37094;
wire n_37095;
wire n_37096;
wire n_37097;
wire n_37098;
wire n_37099;
wire n_37100;
wire n_37101;
wire n_37102;
wire n_37103;
wire n_37104;
wire n_37105;
wire n_37106;
wire n_37107;
wire n_37108;
wire n_37109;
wire n_37110;
wire n_37111;
wire n_37112;
wire n_37113;
wire n_37114;
wire n_37115;
wire n_37116;
wire n_37117;
wire n_37118;
wire n_37119;
wire n_37120;
wire n_37121;
wire n_37122;
wire n_37123;
wire n_37124;
wire n_37125;
wire n_37126;
wire n_37127;
wire n_37128;
wire n_37129;
wire n_37130;
wire n_37131;
wire n_37132;
wire n_37133;
wire n_37134;
wire n_37135;
wire n_37136;
wire n_37137;
wire n_37138;
wire n_37139;
wire n_37140;
wire n_37141;
wire n_37142;
wire n_37143;
wire n_37144;
wire n_37145;
wire n_37146;
wire n_37147;
wire n_37148;
wire n_37149;
wire n_37150;
wire n_37151;
wire n_37152;
wire n_37153;
wire n_37154;
wire n_37155;
wire n_37156;
wire n_37157;
wire n_37158;
wire n_37159;
wire n_37160;
wire n_37161;
wire n_37162;
wire n_37163;
wire n_37164;
wire n_37165;
wire n_37166;
wire n_37167;
wire n_37168;
wire n_37169;
wire n_37170;
wire n_37171;
wire n_37172;
wire n_37173;
wire n_37174;
wire n_37175;
wire n_37176;
wire n_37177;
wire n_37178;
wire n_37179;
wire n_37180;
wire n_37181;
wire n_37182;
wire n_37183;
wire n_37184;
wire n_37185;
wire n_37186;
wire n_37187;
wire n_37188;
wire n_37189;
wire n_37190;
wire n_37191;
wire n_37192;
wire n_37193;
wire n_37194;
wire n_37195;
wire n_37196;
wire n_37197;
wire n_37198;
wire n_37199;
wire n_37200;
wire n_37201;
wire n_37202;
wire n_37203;
wire n_37204;
wire n_37205;
wire n_37206;
wire n_37207;
wire n_37208;
wire n_37209;
wire n_37210;
wire n_37211;
wire n_37212;
wire n_37213;
wire n_37214;
wire n_37215;
wire n_37216;
wire n_37217;
wire n_37218;
wire n_37219;
wire n_37220;
wire n_37221;
wire n_37222;
wire n_37223;
wire n_37224;
wire n_37225;
wire n_37226;
wire n_37227;
wire n_37228;
wire n_37229;
wire n_37230;
wire n_37231;
wire n_37232;
wire n_37233;
wire n_37234;
wire n_37235;
wire n_37236;
wire n_37237;
wire n_37238;
wire n_37239;
wire n_37240;
wire n_37241;
wire n_37242;
wire n_37243;
wire n_37244;
wire n_37245;
wire n_37246;
wire n_37247;
wire n_37248;
wire n_37249;
wire n_37250;
wire n_37251;
wire n_37252;
wire n_37253;
wire n_37254;
wire n_37255;
wire n_37256;
wire n_37257;
wire n_37258;
wire n_37259;
wire n_37260;
wire n_37261;
wire n_37262;
wire n_37263;
wire n_37264;
wire n_37265;
wire n_37266;
wire n_37267;
wire n_37268;
wire n_37269;
wire n_37270;
wire n_37271;
wire n_37272;
wire n_37273;
wire n_37274;
wire n_37275;
wire n_37276;
wire n_37277;
wire n_37278;
wire n_37279;
wire n_37280;
wire n_37281;
wire n_37282;
wire n_37283;
wire n_37284;
wire n_37285;
wire n_37286;
wire n_37287;
wire n_37288;
wire n_37289;
wire n_37290;
wire n_37291;
wire n_37292;
wire n_37293;
wire n_37294;
wire n_37295;
wire n_37296;
wire n_37297;
wire n_37298;
wire n_37299;
wire n_37300;
wire n_37301;
wire n_37302;
wire n_37303;
wire n_37304;
wire n_37305;
wire n_37306;
wire n_37307;
wire n_37308;
wire n_37309;
wire n_37310;
wire n_37311;
wire n_37312;
wire n_37313;
wire n_37314;
wire n_37315;
wire n_37316;
wire n_37317;
wire n_37318;
wire n_37319;
wire n_37320;
wire n_37321;
wire n_37322;
wire n_37323;
wire n_37324;
wire n_37325;
wire n_37326;
wire n_37327;
wire n_37328;
wire n_37329;
wire n_37330;
wire n_37331;
wire n_37332;
wire n_37333;
wire n_37334;
wire n_37335;
wire n_37336;
wire n_37337;
wire n_37338;
wire n_37339;
wire n_37340;
wire n_37341;
wire n_37342;
wire n_37343;
wire n_37344;
wire n_37345;
wire n_37346;
wire n_37347;
wire n_37348;
wire n_37349;
wire n_37350;
wire n_37351;
wire n_37352;
wire n_37353;
wire n_37354;
wire n_37355;
wire n_37356;
wire n_37357;
wire n_37358;
wire n_37359;
wire n_37360;
wire n_37361;
wire n_37362;
wire n_37363;
wire n_37364;
wire n_37365;
wire n_37366;
wire n_37367;
wire n_37368;
wire n_37369;
wire n_37370;
wire n_37371;
wire n_37372;
wire n_37373;
wire n_37374;
wire n_37375;
wire n_37376;
wire n_37377;
wire n_37378;
wire n_37379;
wire n_37380;
wire n_37381;
wire n_37382;
wire n_37383;
wire n_37384;
wire n_37385;
wire n_37386;
wire n_37387;
wire n_37388;
wire n_37389;
wire n_37390;
wire n_37391;
wire n_37392;
wire n_37393;
wire n_37394;
wire n_37395;
wire n_37396;
wire n_37397;
wire n_37398;
wire n_37399;
wire n_37400;
wire n_37401;
wire n_37402;
wire n_37403;
wire n_37404;
wire n_37405;
wire n_37406;
wire n_37407;
wire n_37408;
wire n_37409;
wire n_37410;
wire n_37411;
wire n_37412;
wire n_37413;
wire n_37414;
wire n_37415;
wire n_37416;
wire n_37417;
wire n_37418;
wire n_37419;
wire n_37420;
wire n_37421;
wire n_37422;
wire n_37423;
wire n_37424;
wire n_37425;
wire n_37426;
wire n_37427;
wire n_37428;
wire n_37429;
wire n_37430;
wire n_37431;
wire n_37432;
wire n_37433;
wire n_37434;
wire n_37435;
wire n_37436;
wire n_37437;
wire n_37438;
wire n_37439;
wire n_37440;
wire n_37441;
wire n_37442;
wire n_37443;
wire n_37444;
wire n_37445;
wire n_37446;
wire n_37447;
wire n_37448;
wire n_37449;
wire n_37450;
wire n_37451;
wire n_37452;
wire n_37453;
wire n_37454;
wire n_37455;
wire n_37456;
wire n_37457;
wire n_37458;
wire n_37459;
wire n_37460;
wire n_37461;
wire n_37462;
wire n_37463;
wire n_37464;
wire n_37465;
wire n_37466;
wire n_37467;
wire n_37468;
wire n_37469;
wire n_37470;
wire n_37471;
wire n_37472;
wire n_37473;
wire n_37474;
wire n_37475;
wire n_37476;
wire n_37477;
wire n_37478;
wire n_37479;
wire n_37480;
wire n_37481;
wire n_37482;
wire n_37483;
wire n_37484;
wire n_37485;
wire n_37486;
wire n_37487;
wire n_37488;
wire n_37489;
wire n_37490;
wire n_37491;
wire n_37492;
wire n_37493;
wire n_37494;
wire n_37495;
wire n_37496;
wire n_37497;
wire n_37498;
wire n_37499;
wire n_37500;
wire n_37501;
wire n_37502;
wire n_37503;
wire n_37504;
wire n_37505;
wire n_37506;
wire n_37507;
wire n_37508;
wire n_37509;
wire n_37510;
wire n_37511;
wire n_37512;
wire n_37513;
wire n_37514;
wire n_37515;
wire n_37516;
wire n_37517;
wire n_37518;
wire n_37519;
wire n_37520;
wire n_37521;
wire n_37522;
wire n_37523;
wire n_37524;
wire n_37525;
wire n_37526;
wire n_37527;
wire n_37528;
wire n_37529;
wire n_37530;
wire n_37531;
wire n_37532;
wire n_37533;
wire n_37534;
wire n_37535;
wire n_37536;
wire n_37537;
wire n_37538;
wire n_37539;
wire n_37540;
wire n_37541;
wire n_37542;
wire n_37543;
wire n_37544;
wire n_37545;
wire n_37546;
wire n_37547;
wire n_37548;
wire n_37549;
wire n_37550;
wire n_37551;
wire n_37552;
wire n_37553;
wire n_37554;
wire n_37555;
wire n_37556;
wire n_37557;
wire n_37558;
wire n_37559;
wire n_37560;
wire n_37561;
wire n_37562;
wire n_37563;
wire n_37564;
wire n_37565;
wire n_37566;
wire n_37567;
wire n_37568;
wire n_37569;
wire n_37570;
wire n_37571;
wire n_37572;
wire n_37573;
wire n_37574;
wire n_37575;
wire n_37576;
wire n_37577;
wire n_37578;
wire n_37579;
wire n_37580;
wire n_37581;
wire n_37582;
wire n_37583;
wire n_37584;
wire n_37585;
wire n_37586;
wire n_37587;
wire n_37588;
wire n_37589;
wire n_37590;
wire n_37591;
wire n_37592;
wire n_37593;
wire n_37594;
wire n_37595;
wire n_37596;
wire n_37597;
wire n_37598;
wire n_37599;
wire n_37600;
wire n_37601;
wire n_37602;
wire n_37603;
wire n_37604;
wire n_37605;
wire n_37606;
wire n_37607;
wire n_37608;
wire n_37609;
wire n_37610;
wire n_37611;
wire n_37612;
wire n_37613;
wire n_37614;
wire n_37615;
wire n_37616;
wire n_37617;
wire n_37618;
wire n_37619;
wire n_37620;
wire n_37621;
wire n_37622;
wire n_37623;
wire n_37624;
wire n_37625;
wire n_37626;
wire n_37627;
wire n_37628;
wire n_37629;
wire n_37630;
wire n_37631;
wire n_37632;
wire n_37633;
wire n_37634;
wire n_37635;
wire n_37636;
wire n_37637;
wire n_37638;
wire n_37639;
wire n_37640;
wire n_37641;
wire n_37642;
wire n_37643;
wire n_37644;
wire n_37645;
wire n_37646;
wire n_37647;
wire n_37648;
wire n_37649;
wire n_37650;
wire n_37651;
wire n_37652;
wire n_37653;
wire n_37654;
wire n_37655;
wire n_37656;
wire n_37657;
wire n_37658;
wire n_37659;
wire n_37660;
wire n_37661;
wire n_37662;
wire n_37663;
wire n_37664;
wire n_37665;
wire n_37666;
wire n_37667;
wire n_37668;
wire n_37669;
wire n_37670;
wire n_37671;
wire n_37672;
wire n_37673;
wire n_37674;
wire n_37675;
wire n_37676;
wire n_37677;
wire n_37678;
wire n_37679;
wire n_37680;
wire n_37681;
wire n_37682;
wire n_37683;
wire n_37684;
wire n_37685;
wire n_37686;
wire n_37687;
wire n_37688;
wire n_37689;
wire n_37690;
wire n_37691;
wire n_37692;
wire n_37693;
wire n_37694;
wire n_37695;
wire n_37696;
wire n_37697;
wire n_37698;
wire n_37699;
wire n_37700;
wire n_37701;
wire n_37702;
wire n_37703;
wire n_37704;
wire n_37705;
wire n_37706;
wire n_37707;
wire n_37708;
wire n_37709;
wire n_37710;
wire n_37711;
wire n_37712;
wire n_37713;
wire n_37714;
wire n_37715;
wire n_37716;
wire n_37717;
wire n_37718;
wire n_37719;
wire n_37720;
wire n_37721;
wire n_37722;
wire n_37723;
wire n_37724;
wire n_37725;
wire n_37726;
wire n_37727;
wire n_37728;
wire n_37729;
wire n_37730;
wire n_37731;
wire n_37732;
wire n_37733;
wire n_37734;
wire n_37735;
wire n_37736;
wire n_37737;
wire n_37738;
wire n_37739;
wire n_37740;
wire n_37741;
wire n_37742;
wire n_37743;
wire n_37744;
wire n_37745;
wire n_37746;
wire n_37747;
wire n_37748;
wire n_37749;
wire n_37750;
wire n_37751;
wire n_37752;
wire n_37753;
wire n_37754;
wire n_37755;
wire n_37756;
wire n_37757;
wire n_37758;
wire n_37759;
wire n_37760;
wire n_37761;
wire n_37762;
wire n_37763;
wire n_37764;
wire n_37765;
wire n_37766;
wire n_37767;
wire n_37768;
wire n_37769;
wire n_37770;
wire n_37771;
wire n_37772;
wire n_37773;
wire n_37774;
wire n_37775;
wire n_37776;
wire n_37777;
wire n_37778;
wire n_37779;
wire n_37780;
wire n_37781;
wire n_37782;
wire n_37783;
wire n_37784;
wire n_37785;
wire n_37786;
wire n_37787;
wire n_37788;
wire n_37789;
wire n_37790;
wire n_37791;
wire n_37792;
wire n_37793;
wire n_37794;
wire n_37795;
wire n_37796;
wire n_37797;
wire n_37798;
wire n_37799;
wire n_37800;
wire n_37801;
wire n_37802;
wire n_37803;
wire n_37804;
wire n_37805;
wire n_37806;
wire n_37807;
wire n_37808;
wire n_37809;
wire n_37810;
wire n_37811;
wire n_37812;
wire n_37813;
wire n_37814;
wire n_37815;
wire n_37816;
wire n_37817;
wire n_37818;
wire n_37819;
wire n_37820;
wire n_37821;
wire n_37822;
wire n_37823;
wire n_37824;
wire n_37825;
wire n_37826;
wire n_37827;
wire n_37828;
wire n_37829;
wire n_37830;
wire n_37831;
wire n_37832;
wire n_37833;
wire n_37834;
wire n_37835;
wire n_37836;
wire n_37837;
wire n_37838;
wire n_37839;
wire n_37840;
wire n_37841;
wire n_37842;
wire n_37843;
wire n_37844;
wire n_37845;
wire n_37846;
wire n_37847;
wire n_37848;
wire n_37849;
wire n_37850;
wire n_37851;
wire n_37852;
wire n_37853;
wire n_37854;
wire n_37855;
wire n_37856;
wire n_37857;
wire n_37858;
wire n_37859;
wire n_37860;
wire n_37861;
wire n_37862;
wire n_37863;
wire n_37864;
wire n_37865;
wire n_37866;
wire n_37867;
wire n_37868;
wire n_37869;
wire n_37870;
wire n_37871;
wire n_37872;
wire n_37873;
wire n_37874;
wire n_37875;
wire n_37876;
wire n_37877;
wire n_37878;
wire n_37879;
wire n_37880;
wire n_37881;
wire n_37882;
wire n_37883;
wire n_37884;
wire n_37885;
wire n_37886;
wire n_37887;
wire n_37888;
wire n_37889;
wire n_37890;
wire n_37891;
wire n_37892;
wire n_37893;
wire n_37894;
wire n_37895;
wire n_37896;
wire n_37897;
wire n_37898;
wire n_37899;
wire n_37900;
wire n_37901;
wire n_37902;
wire n_37903;
wire n_37904;
wire n_37905;
wire n_37906;
wire n_37907;
wire n_37908;
wire n_37909;
wire n_37910;
wire n_37911;
wire n_37912;
wire n_37913;
wire n_37914;
wire n_37915;
wire n_37916;
wire n_37917;
wire n_37918;
wire n_37919;
wire n_37920;
wire n_37921;
wire n_37922;
wire n_37923;
wire n_37924;
wire n_37925;
wire n_37926;
wire n_37927;
wire n_37928;
wire n_37929;
wire n_37930;
wire n_37931;
wire n_37932;
wire n_37933;
wire n_37934;
wire n_37935;
wire n_37936;
wire n_37937;
wire n_37938;
wire n_37939;
wire n_37940;
wire n_37941;
wire n_37942;
wire n_37943;
wire n_37944;
wire n_37945;
wire n_37946;
wire n_37947;
wire n_37948;
wire n_37949;
wire n_37950;
wire n_37951;
wire n_37952;
wire n_37953;
wire n_37954;
wire n_37955;
wire n_37956;
wire n_37957;
wire n_37958;
wire n_37959;
wire n_37960;
wire n_37961;
wire n_37962;
wire n_37963;
wire n_37964;
wire n_37965;
wire n_37966;
wire n_37967;
wire n_37968;
wire n_37969;
wire n_37970;
wire n_37971;
wire n_37972;
wire n_37973;
wire n_37974;
wire n_37975;
wire n_37976;
wire n_37977;
wire n_37978;
wire n_37979;
wire n_37980;
wire n_37981;
wire n_37982;
wire n_37983;
wire n_37984;
wire n_37985;
wire n_37986;
wire n_37987;
wire n_37988;
wire n_37989;
wire n_37990;
wire n_37991;
wire n_37992;
wire n_37993;
wire n_37994;
wire n_37995;
wire n_37996;
wire n_37997;
wire n_37998;
wire n_37999;
wire n_38000;
wire n_38001;
wire n_38002;
wire n_38003;
wire n_38004;
wire n_38005;
wire n_38006;
wire n_38007;
wire n_38008;
wire n_38009;
wire n_38010;
wire n_38011;
wire n_38012;
wire n_38013;
wire n_38014;
wire n_38015;
wire n_38016;
wire n_38017;
wire n_38018;
wire n_38019;
wire n_38020;
wire n_38021;
wire n_38022;
wire n_38023;
wire n_38024;
wire n_38025;
wire n_38026;
wire n_38027;
wire n_38028;
wire n_38029;
wire n_38030;
wire n_38031;
wire n_38032;
wire n_38033;
wire n_38034;
wire n_38035;
wire n_38036;
wire n_38037;
wire n_38038;
wire n_38039;
wire n_38040;
wire n_38041;
wire n_38042;
wire n_38043;
wire n_38044;
wire n_38045;
wire n_38046;
wire n_38047;
wire n_38048;
wire n_38049;
wire n_38050;
wire n_38051;
wire n_38052;
wire n_38053;
wire n_38054;
wire n_38055;
wire n_38056;
wire n_38057;
wire n_38058;
wire n_38059;
wire n_38060;
wire n_38061;
wire n_38062;
wire n_38063;
wire n_38064;
wire n_38065;
wire n_38066;
wire n_38067;
wire n_38068;
wire n_38069;
wire n_38070;
wire n_38071;
wire n_38072;
wire n_38073;
wire n_38074;
wire n_38075;
wire n_38076;
wire n_38077;
wire n_38078;
wire n_38079;
wire n_38080;
wire n_38081;
wire n_38082;
wire n_38083;
wire n_38084;
wire n_38085;
wire n_38086;
wire n_38087;
wire n_38088;
wire n_38089;
wire n_38090;
wire n_38091;
wire n_38092;
wire n_38093;
wire n_38094;
wire n_38095;
wire n_38096;
wire n_38097;
wire n_38098;
wire n_38099;
wire n_38100;
wire n_38101;
wire n_38102;
wire n_38103;
wire n_38104;
wire n_38105;
wire n_38106;
wire n_38107;
wire n_38108;
wire n_38109;
wire n_38110;
wire n_38111;
wire n_38112;
wire n_38113;
wire n_38114;
wire n_38115;
wire n_38116;
wire n_38117;
wire n_38118;
wire n_38119;
wire n_38120;
wire n_38121;
wire n_38122;
wire n_38123;
wire n_38124;
wire n_38125;
wire n_38126;
wire n_38127;
wire n_38128;
wire n_38129;
wire n_38130;
wire n_38131;
wire n_38132;
wire n_38133;
wire n_38134;
wire n_38135;
wire n_38136;
wire n_38137;
wire n_38138;
wire n_38139;
wire n_38140;
wire n_38141;
wire n_38142;
wire n_38143;
wire n_38144;
wire n_38145;
wire n_38146;
wire n_38147;
wire n_38148;
wire n_38149;
wire n_38150;
wire n_38151;
wire n_38152;
wire n_38153;
wire n_38154;
wire n_38155;
wire n_38156;
wire n_38157;
wire n_38158;
wire n_38159;
wire n_38160;
wire n_38161;
wire n_38162;
wire n_38163;
wire n_38164;
wire n_38165;
wire n_38166;
wire n_38167;
wire n_38168;
wire n_38169;
wire n_38170;
wire n_38171;
wire n_38172;
wire n_38173;
wire n_38174;
wire n_38175;
wire n_38176;
wire n_38177;
wire n_38178;
wire n_38179;
wire n_38180;
wire n_38181;
wire n_38182;
wire n_38183;
wire n_38184;
wire n_38185;
wire n_38186;
wire n_38187;
wire n_38188;
wire n_38189;
wire n_38190;
wire n_38191;
wire n_38192;
wire n_38193;
wire n_38194;
wire n_38195;
wire n_38196;
wire n_38197;
wire n_38198;
wire n_38199;
wire n_38200;
wire n_38201;
wire n_38202;
wire n_38203;
wire n_38204;
wire n_38205;
wire n_38206;
wire n_38207;
wire n_38208;
wire n_38209;
wire n_38210;
wire n_38211;
wire n_38212;
wire n_38213;
wire n_38214;
wire n_38215;
wire n_38216;
wire n_38217;
wire n_38218;
wire n_38219;
wire n_38220;
wire n_38221;
wire n_38222;
wire n_38223;
wire n_38224;
wire n_38225;
wire n_38226;
wire n_38227;
wire n_38228;
wire n_38229;
wire n_38230;
wire n_38231;
wire n_38232;
wire n_38233;
wire n_38234;
wire n_38235;
wire n_38236;
wire n_38237;
wire n_38238;
wire n_38239;
wire n_38240;
wire n_38241;
wire n_38242;
wire n_38243;
wire n_38244;
wire n_38245;
wire n_38246;
wire n_38247;
wire n_38248;
wire n_38249;
wire n_38250;
wire n_38251;
wire n_38252;
wire n_38253;
wire n_38254;
wire n_38255;
wire n_38256;
wire n_38257;
wire n_38258;
wire n_38259;
wire n_38260;
wire n_38261;
wire n_38262;
wire n_38263;
wire n_38264;
wire n_38265;
wire n_38266;
wire n_38267;
wire n_38268;
wire n_38269;
wire n_38270;
wire n_38271;
wire n_38272;
wire n_38273;
wire n_38274;
wire n_38275;
wire n_38276;
wire n_38277;
wire n_38278;
wire n_38279;
wire n_38280;
wire n_38281;
wire n_38282;
wire n_38283;
wire n_38284;
wire n_38285;
wire n_38286;
wire n_38287;
wire n_38288;
wire n_38289;
wire n_38290;
wire n_38291;
wire n_38292;
wire n_38293;
wire n_38294;
wire n_38295;
wire n_38296;
wire n_38297;
wire n_38298;
wire n_38299;
wire n_38300;
wire n_38301;
wire n_38302;
wire n_38303;
wire n_38304;
wire n_38305;
wire n_38306;
wire n_38307;
wire n_38308;
wire n_38309;
wire n_38310;
wire n_38311;
wire n_38312;
wire n_38313;
wire n_38314;
wire n_38315;
wire n_38316;
wire n_38317;
wire n_38318;
wire n_38319;
wire n_38320;
wire n_38321;
wire n_38322;
wire n_38323;
wire n_38324;
wire n_38325;
wire n_38326;
wire n_38327;
wire n_38328;
wire n_38329;
wire n_38330;
wire n_38331;
wire n_38332;
wire n_38333;
wire n_38334;
wire n_38335;
wire n_38336;
wire n_38337;
wire n_38338;
wire n_38339;
wire n_38340;
wire n_38341;
wire n_38342;
wire n_38343;
wire n_38344;
wire n_38345;
wire n_38346;
wire n_38347;
wire n_38348;
wire n_38349;
wire n_38350;
wire n_38351;
wire n_38352;
wire n_38353;
wire n_38354;
wire n_38355;
wire n_38356;
wire n_38357;
wire n_38358;
wire n_38359;
wire n_38360;
wire n_38361;
wire n_38362;
wire n_38363;
wire n_38364;
wire n_38365;
wire n_38366;
wire n_38367;
wire n_38368;
wire n_38369;
wire n_38370;
wire n_38371;
wire n_38372;
wire n_38373;
wire n_38374;
wire n_38375;
wire n_38376;
wire n_38377;
wire n_38378;
wire n_38379;
wire n_38380;
wire n_38381;
wire n_38382;
wire n_38383;
wire n_38384;
wire n_38385;
wire n_38386;
wire n_38387;
wire n_38388;
wire n_38389;
wire n_38390;
wire n_38391;
wire n_38392;
wire n_38393;
wire n_38394;
wire n_38395;
wire n_38396;
wire n_38397;
wire n_38398;
wire n_38399;
wire n_38400;
wire n_38401;
wire n_38402;
wire n_38403;
wire n_38404;
wire n_38405;
wire n_38406;
wire n_38407;
wire n_38408;
wire n_38409;
wire n_38410;
wire n_38411;
wire n_38412;
wire n_38413;
wire n_38414;
wire n_38415;
wire n_38416;
wire n_38417;
wire n_38418;
wire n_38419;
wire n_38420;
wire n_38421;
wire n_38422;
wire n_38423;
wire n_38424;
wire n_38425;
wire n_38426;
wire n_38427;
wire n_38428;
wire n_38429;
wire n_38430;
wire n_38431;
wire n_38432;
wire n_38433;
wire n_38434;
wire n_38435;
wire n_38436;
wire n_38437;
wire n_38438;
wire n_38439;
wire n_38440;
wire n_38441;
wire n_38442;
wire n_38443;
wire n_38444;
wire n_38445;
wire n_38446;
wire n_38447;
wire n_38448;
wire n_38449;
wire n_38450;
wire n_38451;
wire n_38452;
wire n_38453;
wire n_38454;
wire n_38455;
wire n_38456;
wire n_38457;
wire n_38458;
wire n_38459;
wire n_38460;
wire n_38461;
wire n_38462;
wire n_38463;
wire n_38464;
wire n_38465;
wire n_38466;
wire n_38467;
wire n_38468;
wire n_38469;
wire n_38470;
wire n_38471;
wire n_38472;
wire n_38473;
wire n_38474;
wire n_38475;
wire n_38476;
wire n_38477;
wire n_38478;
wire n_38479;
wire n_38480;
wire n_38481;
wire n_38482;
wire n_38483;
wire n_38484;
wire n_38485;
wire n_38486;
wire n_38487;
wire n_38488;
wire n_38489;
wire n_38490;
wire n_38491;
wire n_38492;
wire n_38493;
wire n_38494;
wire n_38495;
wire n_38496;
wire n_38497;
wire n_38498;
wire n_38499;
wire n_38500;
wire n_38501;
wire n_38502;
wire n_38503;
wire n_38504;
wire n_38505;
wire n_38506;
wire n_38507;
wire n_38508;
wire n_38509;
wire n_38510;
wire n_38511;
wire n_38512;
wire n_38513;
wire n_38514;
wire n_38515;
wire n_38516;
wire n_38517;
wire n_38518;
wire n_38519;
wire n_38520;
wire n_38521;
wire n_38522;
wire n_38523;
wire n_38524;
wire n_38525;
wire n_38526;
wire n_38527;
wire n_38528;
wire n_38529;
wire n_38530;
wire n_38531;
wire n_38532;
wire n_38533;
wire n_38534;
wire n_38535;
wire n_38536;
wire n_38537;
wire n_38538;
wire n_38539;
wire n_38540;
wire n_38541;
wire n_38542;
wire n_38543;
wire n_38544;
wire n_38545;
wire n_38546;
wire n_38547;
wire n_38548;
wire n_38549;
wire n_38550;
wire n_38551;
wire n_38552;
wire n_38553;
wire n_38554;
wire n_38555;
wire n_38556;
wire n_38557;
wire n_38558;
wire n_38559;
wire n_38560;
wire n_38561;
wire n_38562;
wire n_38563;
wire n_38564;
wire n_38565;
wire n_38566;
wire n_38567;
wire n_38568;
wire n_38569;
wire n_38570;
wire n_38571;
wire n_38572;
wire n_38573;
wire n_38574;
wire n_38575;
wire n_38576;
wire n_38577;
wire n_38578;
wire n_38579;
wire n_38580;
wire n_38581;
wire n_38582;
wire n_38583;
wire n_38584;
wire n_38585;
wire n_38586;
wire n_38587;
wire n_38588;
wire n_38589;
wire n_38590;
wire n_38591;
wire n_38592;
wire n_38593;
wire n_38594;
wire n_38595;
wire n_38596;
wire n_38597;
wire n_38598;
wire n_38599;
wire n_38600;
wire n_38601;
wire n_38602;
wire n_38603;
wire n_38604;
wire n_38605;
wire n_38606;
wire n_38607;
wire n_38608;
wire n_38609;
wire n_38610;
wire n_38611;
wire n_38612;
wire n_38613;
wire n_38614;
wire n_38615;
wire n_38616;
wire n_38617;
wire n_38618;
wire n_38619;
wire n_38620;
wire n_38621;
wire n_38622;
wire n_38623;
wire n_38624;
wire n_38625;
wire n_38626;
wire n_38627;
wire n_38628;
wire n_38629;
wire n_38630;
wire n_38631;
wire n_38632;
wire n_38633;
wire n_38634;
wire n_38635;
wire n_38636;
wire n_38637;
wire n_38638;
wire n_38639;
wire n_38640;
wire n_38641;
wire n_38642;
wire n_38643;
wire n_38644;
wire n_38645;
wire n_38646;
wire n_38647;
wire n_38648;
wire n_38649;
wire n_38650;
wire n_38651;
wire n_38652;
wire n_38653;
wire n_38654;
wire n_38655;
wire n_38656;
wire n_38657;
wire n_38658;
wire n_38659;
wire n_38660;
wire n_38661;
wire n_38662;
wire n_38663;
wire n_38664;
wire n_38665;
wire n_38666;
wire n_38667;
wire n_38668;
wire n_38669;
wire n_38670;
wire n_38671;
wire n_38672;
wire n_38673;
wire n_38674;
wire n_38675;
wire n_38676;
wire n_38677;
wire n_38678;
wire n_38679;
wire n_38680;
wire n_38681;
wire n_38682;
wire n_38683;
wire n_38684;
wire n_38685;
wire n_38686;
wire n_38687;
wire n_38688;
wire n_38689;
wire n_38690;
wire n_38691;
wire n_38692;
wire n_38693;
wire n_38694;
wire n_38695;
wire n_38696;
wire n_38697;
wire n_38698;
wire n_38699;
wire n_38700;
wire n_38701;
wire n_38702;
wire n_38703;
wire n_38704;
wire n_38705;
wire n_38706;
wire n_38707;
wire n_38708;
wire n_38709;
wire n_38710;
wire n_38711;
wire n_38712;
wire n_38713;
wire n_38714;
wire n_38715;
wire n_38716;
wire n_38717;
wire n_38718;
wire n_38719;
wire n_38720;
wire n_38721;
wire n_38722;
wire n_38723;
wire n_38724;
wire n_38725;
wire n_38726;
wire n_38727;
wire n_38728;
wire n_38729;
wire n_38730;
wire n_38731;
wire n_38732;
wire n_38733;
wire n_38734;
wire n_38735;
wire n_38736;
wire n_38737;
wire n_38738;
wire n_38739;
wire n_38740;
wire n_38741;
wire n_38742;
wire n_38743;
wire n_38744;
wire n_38745;
wire n_38746;
wire n_38747;
wire n_38748;
wire n_38749;
wire n_38750;
wire n_38751;
wire n_38752;
wire n_38753;
wire n_38754;
wire n_38755;
wire n_38756;
wire n_38757;
wire n_38758;
wire n_38759;
wire n_38760;
wire n_38761;
wire n_38762;
wire n_38763;
wire n_38764;
wire n_38765;
wire n_38766;
wire n_38767;
wire n_38768;
wire n_38769;
wire n_38770;
wire n_38771;
wire n_38772;
wire n_38773;
wire n_38774;
wire n_38775;
wire n_38776;
wire n_38777;
wire n_38778;
wire n_38779;
wire n_38780;
wire n_38781;
wire n_38782;
wire n_38783;
wire n_38784;
wire n_38785;
wire n_38786;
wire n_38787;
wire n_38788;
wire n_38789;
wire n_38790;
wire n_38791;
wire n_38792;
wire n_38793;
wire n_38794;
wire n_38795;
wire n_38796;
wire n_38797;
wire n_38798;
wire n_38799;
wire n_38800;
wire n_38801;
wire n_38802;
wire n_38803;
wire n_38804;
wire n_38805;
wire n_38806;
wire n_38807;
wire n_38808;
wire n_38809;
wire n_38810;
wire n_38811;
wire n_38812;
wire n_38813;
wire n_38814;
wire n_38815;
wire n_38816;
wire n_38817;
wire n_38818;
wire n_38819;
wire n_38820;
wire n_38821;
wire n_38822;
wire n_38823;
wire n_38824;
wire n_38825;
wire n_38826;
wire n_38827;
wire n_38828;
wire n_38829;
wire n_38830;
wire n_38831;
wire n_38832;
wire n_38833;
wire n_38834;
wire n_38835;
wire n_38836;
wire n_38837;
wire n_38838;
wire n_38839;
wire n_38840;
wire n_38841;
wire n_38842;
wire n_38843;
wire n_38844;
wire n_38845;
wire n_38846;
wire n_38847;
wire n_38848;
wire n_38849;
wire n_38850;
wire n_38851;
wire n_38852;
wire n_38853;
wire n_38854;
wire n_38855;
wire n_38856;
wire n_38857;
wire n_38858;
wire n_38859;
wire n_38860;
wire n_38861;
wire n_38862;
wire n_38863;
wire n_38864;
wire n_38865;
wire n_38866;
wire n_38867;
wire n_38868;
wire n_38869;
wire n_38870;
wire n_38871;
wire n_38872;
wire n_38873;
wire n_38874;
wire n_38875;
wire n_38876;
wire n_38877;
wire n_38878;
wire n_38879;
wire n_38880;
wire n_38881;
wire n_38882;
wire n_38883;
wire n_38884;
wire n_38885;
wire n_38886;
wire n_38887;
wire n_38888;
wire n_38889;
wire n_38890;
wire n_38891;
wire n_38892;
wire n_38893;
wire n_38894;
wire n_38895;
wire n_38896;
wire n_38897;
wire n_38898;
wire n_38899;
wire n_38900;
wire n_38901;
wire n_38902;
wire n_38903;
wire n_38904;
wire n_38905;
wire n_38906;
wire n_38907;
wire n_38908;
wire n_38909;
wire n_38910;
wire n_38911;
wire n_38912;
wire n_38913;
wire n_38914;
wire n_38915;
wire n_38916;
wire n_38917;
wire n_38918;
wire n_38919;
wire n_38920;
wire n_38921;
wire n_38922;
wire n_38923;
wire n_38924;
wire n_38925;
wire n_38926;
wire n_38927;
wire n_38928;
wire n_38929;
wire n_38930;
wire n_38931;
wire n_38932;
wire n_38933;
wire n_38934;
wire n_38935;
wire n_38936;
wire n_38937;
wire n_38938;
wire n_38939;
wire n_38940;
wire n_38941;
wire n_38942;
wire n_38943;
wire n_38944;
wire n_38945;
wire n_38946;
wire n_38947;
wire n_38948;
wire n_38949;
wire n_38950;
wire n_38951;
wire n_38952;
wire n_38953;
wire n_38954;
wire n_38955;
wire n_38956;
wire n_38957;
wire n_38958;
wire n_38959;
wire n_38960;
wire n_38961;
wire n_38962;
wire n_38963;
wire n_38964;
wire n_38965;
wire n_38966;
wire n_38967;
wire n_38968;
wire n_38969;
wire n_38970;
wire n_38971;
wire n_38972;
wire n_38973;
wire n_38974;
wire n_38975;
wire n_38976;
wire n_38977;
wire n_38978;
wire n_38979;
wire n_38980;
wire n_38981;
wire n_38982;
wire n_38983;
wire n_38984;
wire n_38985;
wire n_38986;
wire n_38987;
wire n_38988;
wire n_38989;
wire n_38990;
wire n_38991;
wire n_38992;
wire n_38993;
wire n_38994;
wire n_38995;
wire n_38996;
wire n_38997;
wire n_38998;
wire n_38999;
wire n_39000;
wire n_39001;
wire n_39002;
wire n_39003;
wire n_39004;
wire n_39005;
wire n_39006;
wire n_39007;
wire n_39008;
wire n_39009;
wire n_39010;
wire n_39011;
wire n_39012;
wire n_39013;
wire n_39014;
wire n_39015;
wire n_39016;
wire n_39017;
wire n_39018;
wire n_39019;
wire n_39020;
wire n_39021;
wire n_39022;
wire n_39023;
wire n_39024;
wire n_39025;
wire n_39026;
wire n_39027;
wire n_39028;
wire n_39029;
wire n_39030;
wire n_39031;
wire n_39032;
wire n_39033;
wire n_39034;
wire n_39035;
wire n_39036;
wire n_39037;
wire n_39038;
wire n_39039;
wire n_39040;
wire n_39041;
wire n_39042;
wire n_39043;
wire n_39044;
wire n_39045;
wire n_39046;
wire n_39047;
wire n_39048;
wire n_39049;
wire n_39050;
wire n_39051;
wire n_39052;
wire n_39053;
wire n_39054;
wire n_39055;
wire n_39056;
wire n_39057;
wire n_39058;
wire n_39059;
wire n_39060;
wire n_39061;
wire n_39062;
wire n_39063;
wire n_39064;
wire n_39065;
wire n_39066;
wire n_39067;
wire n_39068;
wire n_39069;
wire n_39070;
wire n_39071;
wire n_39072;
wire n_39073;
wire n_39074;
wire n_39075;
wire n_39076;
wire n_39077;
wire n_39078;
wire n_39079;
wire n_39080;
wire n_39081;
wire n_39082;
wire n_39083;
wire n_39084;
wire n_39085;
wire n_39086;
wire n_39087;
wire n_39088;
wire n_39089;
wire n_39090;
wire n_39091;
wire n_39092;
wire n_39093;
wire n_39094;
wire n_39095;
wire n_39096;
wire n_39097;
wire n_39098;
wire n_39099;
wire n_39100;
wire n_39101;
wire n_39102;
wire n_39103;
wire n_39104;
wire n_39105;
wire n_39106;
wire n_39107;
wire n_39108;
wire n_39109;
wire n_39110;
wire n_39111;
wire n_39112;
wire n_39113;
wire n_39114;
wire n_39115;
wire n_39116;
wire n_39117;
wire n_39118;
wire n_39119;
wire n_39120;
wire n_39121;
wire n_39122;
wire n_39123;
wire n_39124;
wire n_39125;
wire n_39126;
wire n_39127;
wire n_39128;
wire n_39129;
wire n_39130;
wire n_39131;
wire n_39132;
wire n_39133;
wire n_39134;
wire n_39135;
wire n_39136;
wire n_39137;
wire n_39138;
wire n_39139;
wire n_39140;
wire n_39141;
wire n_39142;
wire n_39143;
wire n_39144;
wire n_39145;
wire n_39146;
wire n_39147;
wire n_39148;
wire n_39149;
wire n_39150;
wire n_39151;
wire n_39152;
wire n_39153;
wire n_39154;
wire n_39155;
wire n_39156;
wire n_39157;
wire n_39158;
wire n_39159;
wire n_39160;
wire n_39161;
wire n_39162;
wire n_39163;
wire n_39164;
wire n_39165;
wire n_39166;
wire n_39167;
wire n_39168;
wire n_39169;
wire n_39170;
wire n_39171;
wire n_39172;
wire n_39173;
wire n_39174;
wire n_39175;
wire n_39176;
wire n_39177;
wire n_39178;
wire n_39179;
wire n_39180;
wire n_39181;
wire n_39182;
wire n_39183;
wire n_39184;
wire n_39185;
wire n_39186;
wire n_39187;
wire n_39188;
wire n_39189;
wire n_39190;
wire n_39191;
wire n_39192;
wire n_39193;
wire n_39194;
wire n_39195;
wire n_39196;
wire n_39197;
wire n_39198;
wire n_39199;
wire n_39200;
wire n_39201;
wire n_39202;
wire n_39203;
wire n_39204;
wire n_39205;
wire n_39206;
wire n_39207;
wire n_39208;
wire n_39209;
wire n_39210;
wire n_39211;
wire n_39212;
wire n_39213;
wire n_39214;
wire n_39215;
wire n_39216;
wire n_39217;
wire n_39218;
wire n_39219;
wire n_39220;
wire n_39221;
wire n_39222;
wire n_39223;
wire n_39224;
wire n_39225;
wire n_39226;
wire n_39227;
wire n_39228;
wire n_39229;
wire n_39230;
wire n_39231;
wire n_39232;
wire n_39233;
wire n_39234;
wire n_39235;
wire n_39236;
wire n_39237;
wire n_39238;
wire n_39239;
wire n_39240;
wire n_39241;
wire n_39242;
wire n_39243;
wire n_39244;
wire n_39245;
wire n_39246;
wire n_39247;
wire n_39248;
wire n_39249;
wire n_39250;
wire n_39251;
wire n_39252;
wire n_39253;
wire n_39254;
wire n_39255;
wire n_39256;
wire n_39257;
wire n_39258;
wire n_39259;
wire n_39260;
wire n_39261;
wire n_39262;
wire n_39263;
wire n_39264;
wire n_39265;
wire n_39266;
wire n_39267;
wire n_39268;
wire n_39269;
wire n_39270;
wire n_39271;
wire n_39272;
wire n_39273;
wire n_39274;
wire n_39275;
wire n_39276;
wire n_39277;
wire n_39278;
wire n_39279;
wire n_39280;
wire n_39281;
wire n_39282;
wire n_39283;
wire n_39284;
wire n_39285;
wire n_39286;
wire n_39287;
wire n_39288;
wire n_39289;
wire n_39290;
wire n_39291;
wire n_39292;
wire n_39293;
wire n_39294;
wire n_39295;
wire n_39296;
wire n_39297;
wire n_39298;
wire n_39299;
wire n_39300;
wire n_39301;
wire n_39302;
wire n_39303;
wire n_39304;
wire n_39305;
wire n_39306;
wire n_39307;
wire n_39308;
wire n_39309;
wire n_39310;
wire n_39311;
wire n_39312;
wire n_39313;
wire n_39314;
wire n_39315;
wire n_39316;
wire n_39317;
wire n_39318;
wire n_39319;
wire n_39320;
wire n_39321;
wire n_39322;
wire n_39323;
wire n_39324;
wire n_39325;
wire n_39326;
wire n_39327;
wire n_39328;
wire n_39329;
wire n_39330;
wire n_39331;
wire n_39332;
wire n_39333;
wire n_39334;
wire n_39335;
wire n_39336;
wire n_39337;
wire n_39338;
wire n_39339;
wire n_39340;
wire n_39341;
wire n_39342;
wire n_39343;
wire n_39344;
wire n_39345;
wire n_39346;
wire n_39347;
wire n_39348;
wire n_39349;
wire n_39350;
wire n_39351;
wire n_39352;
wire n_39353;
wire n_39354;
wire n_39355;
wire n_39356;
wire n_39357;
wire n_39358;
wire n_39359;
wire n_39360;
wire n_39361;
wire n_39362;
wire n_39363;
wire n_39364;
wire n_39365;
wire n_39366;
wire n_39367;
wire n_39368;
wire n_39369;
wire n_39370;
wire n_39371;
wire n_39372;
wire n_39373;
wire n_39374;
wire n_39375;
wire n_39376;
wire n_39377;
wire n_39378;
wire n_39379;
wire n_39380;
wire n_39381;
wire n_39382;
wire n_39383;
wire n_39384;
wire n_39385;
wire n_39386;
wire n_39387;
wire n_39388;
wire n_39389;
wire n_39390;
wire n_39391;
wire n_39392;
wire n_39393;
wire n_39394;
wire n_39395;
wire n_39396;
wire n_39397;
wire n_39398;
wire n_39399;
wire n_39400;
wire n_39401;
wire n_39402;
wire n_39403;
wire n_39404;
wire n_39405;
wire n_39406;
wire n_39407;
wire n_39408;
wire n_39409;
wire n_39410;
wire n_39411;
wire n_39412;
wire n_39413;
wire n_39414;
wire n_39415;
wire n_39416;
wire n_39417;
wire n_39418;
wire n_39419;
wire n_39420;
wire n_39421;
wire n_39422;
wire n_39423;
wire n_39424;
wire n_39425;
wire n_39426;
wire n_39427;
wire n_39428;
wire n_39429;
wire n_39430;
wire n_39431;
wire n_39432;
wire n_39433;
wire n_39434;
wire n_39435;
wire n_39436;
wire n_39437;
wire n_39438;
wire n_39439;
wire n_39440;
wire n_39441;
wire n_39442;
wire n_39443;
wire n_39444;
wire n_39445;
wire n_39446;
wire n_39447;
wire n_39448;
wire n_39449;
wire n_39450;
wire n_39451;
wire n_39452;
wire n_39453;
wire n_39454;
wire n_39455;
wire n_39456;
wire n_39457;
wire n_39458;
wire n_39459;
wire n_39460;
wire n_39461;
wire n_39462;
wire n_39463;
wire n_39464;
wire n_39465;
wire n_39466;
wire n_39467;
wire n_39468;
wire n_39469;
wire n_39470;
wire n_39471;
wire n_39472;
wire n_39473;
wire n_39474;
wire n_39475;
wire n_39476;
wire n_39477;
wire n_39478;
wire n_39479;
wire n_39480;
wire n_39481;
wire n_39482;
wire n_39483;
wire n_39484;
wire n_39485;
wire n_39486;
wire n_39487;
wire n_39488;
wire n_39489;
wire n_39490;
wire n_39491;
wire n_39492;
wire n_39493;
wire n_39494;
wire n_39495;
wire n_39496;
wire n_39497;
wire n_39498;
wire n_39499;
wire n_39500;
wire n_39501;
wire n_39502;
wire n_39503;
wire n_39504;
wire n_39505;
wire n_39506;
wire n_39507;
wire n_39508;
wire n_39509;
wire n_39510;
wire n_39511;
wire n_39512;
wire n_39513;
wire n_39514;
wire n_39515;
wire n_39516;
wire n_39517;
wire n_39518;
wire n_39519;
wire n_39520;
wire n_39521;
wire n_39522;
wire n_39523;
wire n_39524;
wire n_39525;
wire n_39526;
wire n_39527;
wire n_39528;
wire n_39529;
wire n_39530;
wire n_39531;
wire n_39532;
wire n_39533;
wire n_39534;
wire n_39535;
wire n_39536;
wire n_39537;
wire n_39538;
wire n_39539;
wire n_39540;
wire n_39541;
wire n_39542;
wire n_39543;
wire n_39544;
wire n_39545;
wire n_39546;
wire n_39547;
wire n_39548;
wire n_39549;
wire n_39550;
wire n_39551;
wire n_39552;
wire n_39553;
wire n_39554;
wire n_39555;
wire n_39556;
wire n_39557;
wire n_39558;
wire n_39559;
wire n_39560;
wire n_39561;
wire n_39562;
wire n_39563;
wire n_39564;
wire n_39565;
wire n_39566;
wire n_39567;
wire n_39568;
wire n_39569;
wire n_39570;
wire n_39571;
wire n_39572;
wire n_39573;
wire n_39574;
wire n_39575;
wire n_39576;
wire n_39577;
wire n_39578;
wire n_39579;
wire n_39580;
wire n_39581;
wire n_39582;
wire n_39583;
wire n_39584;
wire n_39585;
wire n_39586;
wire n_39587;
wire n_39588;
wire n_39589;
wire n_39590;
wire n_39591;
wire n_39592;
wire n_39593;
wire n_39594;
wire n_39595;
wire n_39596;
wire n_39597;
wire n_39598;
wire n_39599;
wire n_39600;
wire n_39601;
wire n_39602;
wire n_39603;
wire n_39604;
wire n_39605;
wire n_39606;
wire n_39607;
wire n_39608;
wire n_39609;
wire n_39610;
wire n_39611;
wire n_39612;
wire n_39613;
wire n_39614;
wire n_39615;
wire n_39616;
wire n_39617;
wire n_39618;
wire n_39619;
wire n_39620;
wire n_39621;
wire n_39622;
wire n_39623;
wire n_39624;
wire n_39625;
wire n_39626;
wire n_39627;
wire n_39628;
wire n_39629;
wire n_39630;
wire n_39631;
wire n_39632;
wire n_39633;
wire n_39634;
wire n_39635;
wire n_39636;
wire n_39637;
wire n_39638;
wire n_39639;
wire n_39640;
wire n_39641;
wire n_39642;
wire n_39643;
wire n_39644;
wire n_39645;
wire n_39646;
wire n_39647;
wire n_39648;
wire n_39649;
wire n_39650;
wire n_39651;
wire n_39652;
wire n_39653;
wire n_39654;
wire n_39655;
wire n_39656;
wire n_39657;
wire n_39658;
wire n_39659;
wire n_39660;
wire n_39661;
wire n_39662;
wire n_39663;
wire n_39664;
wire n_39665;
wire n_39666;
wire n_39667;
wire n_39668;
wire n_39669;
wire n_39670;
wire n_39671;
wire n_39672;
wire n_39673;
wire n_39674;
wire n_39675;
wire n_39676;
wire n_39677;
wire n_39678;
wire n_39679;
wire n_39680;
wire n_39681;
wire n_39682;
wire n_39683;
wire n_39684;
wire n_39685;
wire n_39686;
wire n_39687;
wire n_39688;
wire n_39689;
wire n_39690;
wire n_39691;
wire n_39692;
wire n_39693;
wire n_39694;
wire n_39695;
wire n_39696;
wire n_39697;
wire n_39698;
wire n_39699;
wire n_39700;
wire n_39701;
wire n_39702;
wire n_39703;
wire n_39704;
wire n_39705;
wire n_39706;
wire n_39707;
wire n_39708;
wire n_39709;
wire n_39710;
wire n_39711;
wire n_39712;
wire n_39713;
wire n_39714;
wire n_39715;
wire n_39716;
wire n_39717;
wire n_39718;
wire n_39719;
wire n_39720;
wire n_39721;
wire n_39722;
wire n_39723;
wire n_39724;
wire n_39725;
wire n_39726;
wire n_39727;
wire n_39728;
wire n_39729;
wire n_39730;
wire n_39731;
wire n_39732;
wire n_39733;
wire n_39734;
wire n_39735;
wire n_39736;
wire n_39737;
wire n_39738;
wire n_39739;
wire n_39740;
wire n_39741;
wire n_39742;
wire n_39743;
wire n_39744;
wire n_39745;
wire n_39746;
wire n_39747;
wire n_39748;
wire n_39749;
wire n_39750;
wire n_39751;
wire n_39752;
wire n_39753;
wire n_39754;
wire n_39755;
wire n_39756;
wire n_39757;
wire n_39758;
wire n_39759;
wire n_39760;
wire n_39761;
wire n_39762;
wire n_39763;
wire n_39764;
wire n_39765;
wire n_39766;
wire n_39767;
wire n_39768;
wire n_39769;
wire n_39770;
wire n_39771;
wire n_39772;
wire n_39773;
wire n_39774;
wire n_39775;
wire n_39776;
wire n_39777;
wire n_39778;
wire n_39779;
wire n_39780;
wire n_39781;
wire n_39782;
wire n_39783;
wire n_39784;
wire n_39785;
wire n_39786;
wire n_39787;
wire n_39788;
wire n_39789;
wire n_39790;
wire n_39791;
wire n_39792;
wire n_39793;
wire n_39794;
wire n_39795;
wire n_39796;
wire n_39797;
wire n_39798;
wire n_39799;
wire n_39800;
wire n_39801;
wire n_39802;
wire n_39803;
wire n_39804;
wire n_39805;
wire n_39806;
wire n_39807;
wire n_39808;
wire n_39809;
wire n_39810;
wire n_39811;
wire n_39812;
wire n_39813;
wire n_39814;
wire n_39815;
wire n_39816;
wire n_39817;
wire n_39818;
wire n_39819;
wire n_39820;
wire n_39821;
wire n_39822;
wire n_39823;
wire n_39824;
wire n_39825;
wire n_39826;
wire n_39827;
wire n_39828;
wire n_39829;
wire n_39830;
wire n_39831;
wire n_39832;
wire n_39833;
wire n_39834;
wire n_39835;
wire n_39836;
wire n_39837;
wire n_39838;
wire n_39839;
wire n_39840;
wire n_39841;
wire n_39842;
wire n_39843;
wire n_39844;
wire n_39845;
wire n_39846;
wire n_39847;
wire n_39848;
wire n_39849;
wire n_39850;
wire n_39851;
wire n_39852;
wire n_39853;
wire n_39854;
wire n_39855;
wire n_39856;
wire n_39857;
wire n_39858;
wire n_39859;
wire n_39860;
wire n_39861;
wire n_39862;
wire n_39863;
wire n_39864;
wire n_39865;
wire n_39866;
wire n_39867;
wire n_39868;
wire n_39869;
wire n_39870;
wire n_39871;
wire n_39872;
wire n_39873;
wire n_39874;
wire n_39875;
wire n_39876;
wire n_39877;
wire n_39878;
wire n_39879;
wire n_39880;
wire n_39881;
wire n_39882;
wire n_39883;
wire n_39884;
wire n_39885;
wire n_39886;
wire n_39887;
wire n_39888;
wire n_39889;
wire n_39890;
wire n_39891;
wire n_39892;
wire n_39893;
wire n_39894;
wire n_39895;
wire n_39896;
wire n_39897;
wire n_39898;
wire n_39899;
wire n_39900;
wire n_39901;
wire n_39902;
wire n_39903;
wire n_39904;
wire n_39905;
wire n_39906;
wire n_39907;
wire n_39908;
wire n_39909;
wire n_39910;
wire n_39911;
wire n_39912;
wire n_39913;
wire n_39914;
wire n_39915;
wire n_39916;
wire n_39917;
wire n_39918;
wire n_39919;
wire n_39920;
wire n_39921;
wire n_39922;
wire n_39923;
wire n_39924;
wire n_39925;
wire n_39926;
wire n_39927;
wire n_39928;
wire n_39929;
wire n_39930;
wire n_39931;
wire n_39932;
wire n_39933;
wire n_39934;
wire n_39935;
wire n_39936;
wire n_39937;
wire n_39938;
wire n_39939;
wire n_39940;
wire n_39941;
wire n_39942;
wire n_39943;
wire n_39944;
wire n_39945;
wire n_39946;
wire n_39947;
wire n_39948;
wire n_39949;
wire n_39950;
wire n_39951;
wire n_39952;
wire n_39953;
wire n_39954;
wire n_39955;
wire n_39956;
wire n_39957;
wire n_39958;
wire n_39959;
wire n_39960;
wire n_39961;
wire n_39962;
wire n_39963;
wire n_39964;
wire n_39965;
wire n_39966;
wire n_39967;
wire n_39968;
wire n_39969;
wire n_39970;
wire n_39971;
wire n_39972;
wire n_39973;
wire n_39974;
wire n_39975;
wire n_39976;
wire n_39977;
wire n_39978;
wire n_39979;
wire n_39980;
wire n_39981;
wire n_39982;
wire n_39983;
wire n_39984;
wire n_39985;
wire n_39986;
wire n_39987;
wire n_39988;
wire n_39989;
wire n_39990;
wire n_39991;
wire n_39992;
wire n_39993;
wire n_39994;
wire n_39995;
wire n_39996;
wire n_39997;
wire n_39998;
wire n_39999;
wire n_40000;
wire n_40001;
wire n_40002;
wire n_40003;
wire n_40004;
wire n_40005;
wire n_40006;
wire n_40007;
wire n_40008;
wire n_40009;
wire n_40010;
wire n_40011;
wire n_40012;
wire n_40013;
wire n_40014;
wire n_40015;
wire n_40016;
wire n_40017;
wire n_40018;
wire n_40019;
wire n_40020;
wire n_40021;
wire n_40022;
wire n_40023;
wire n_40024;
wire n_40025;
wire n_40026;
wire n_40027;
wire n_40028;
wire n_40029;
wire n_40030;
wire n_40031;
wire n_40032;
wire n_40033;
wire n_40034;
wire n_40035;
wire n_40036;
wire n_40037;
wire n_40038;
wire n_40039;
wire n_40040;
wire n_40041;
wire n_40042;
wire n_40043;
wire n_40044;
wire n_40045;
wire n_40046;
wire n_40047;
wire n_40048;
wire n_40049;
wire n_40050;
wire n_40051;
wire n_40052;
wire n_40053;
wire n_40054;
wire n_40055;
wire n_40056;
wire n_40057;
wire n_40058;
wire n_40059;
wire n_40060;
wire n_40061;
wire n_40062;
wire n_40063;
wire n_40064;
wire n_40065;
wire n_40066;
wire n_40067;
wire n_40068;
wire n_40069;
wire n_40070;
wire n_40071;
wire n_40072;
wire n_40073;
wire n_40074;
wire n_40075;
wire n_40076;
wire n_40077;
wire n_40078;
wire n_40079;
wire n_40080;
wire n_40081;
wire n_40082;
wire n_40083;
wire n_40084;
wire n_40085;
wire n_40086;
wire n_40087;
wire n_40088;
wire n_40089;
wire n_40090;
wire n_40091;
wire n_40092;
wire n_40093;
wire n_40094;
wire n_40095;
wire n_40096;
wire n_40097;
wire n_40098;
wire n_40099;
wire n_40100;
wire n_40101;
wire n_40102;
wire n_40103;
wire n_40104;
wire n_40105;
wire n_40106;
wire n_40107;
wire n_40108;
wire n_40109;
wire n_40110;
wire n_40111;
wire n_40112;
wire n_40113;
wire n_40114;
wire n_40115;
wire n_40116;
wire n_40117;
wire n_40118;
wire n_40119;
wire n_40120;
wire n_40121;
wire n_40122;
wire n_40123;
wire n_40124;
wire n_40125;
wire n_40126;
wire n_40127;
wire n_40128;
wire n_40129;
wire n_40130;
wire n_40131;
wire n_40132;
wire n_40133;
wire n_40134;
wire n_40135;
wire n_40136;
wire n_40137;
wire n_40138;
wire n_40139;
wire n_40140;
wire n_40141;
wire n_40142;
wire n_40143;
wire n_40144;
wire n_40145;
wire n_40146;
wire n_40147;
wire n_40148;
wire n_40149;
wire n_40150;
wire n_40151;
wire n_40152;
wire n_40153;
wire n_40154;
wire n_40155;
wire n_40156;
wire n_40157;
wire n_40158;
wire n_40159;
wire n_40160;
wire n_40161;
wire n_40162;
wire n_40163;
wire n_40164;
wire n_40165;
wire n_40166;
wire n_40167;
wire n_40168;
wire n_40169;
wire n_40170;
wire n_40171;
wire n_40172;
wire n_40173;
wire n_40174;
wire n_40175;
wire n_40176;
wire n_40177;
wire n_40178;
wire n_40179;
wire n_40180;
wire n_40181;
wire n_40182;
wire n_40183;
wire n_40184;
wire n_40185;
wire n_40186;
wire n_40187;
wire n_40188;
wire n_40189;
wire n_40190;
wire n_40191;
wire n_40192;
wire n_40193;
wire n_40194;
wire n_40195;
wire n_40196;
wire n_40197;
wire n_40198;
wire n_40199;
wire n_40200;
wire n_40201;
wire n_40202;
wire n_40203;
wire n_40204;
wire n_40205;
wire n_40206;
wire n_40207;
wire n_40208;
wire n_40209;
wire n_40210;
wire n_40211;
wire n_40212;
wire n_40213;
wire n_40214;
wire n_40215;
wire n_40216;
wire n_40217;
wire n_40218;
wire n_40219;
wire n_40220;
wire n_40221;
wire n_40222;
wire n_40223;
wire n_40224;
wire n_40225;
wire n_40226;
wire n_40227;
wire n_40228;
wire n_40229;
wire n_40230;
wire n_40231;
wire n_40232;
wire n_40233;
wire n_40234;
wire n_40235;
wire n_40236;
wire n_40237;
wire n_40238;
wire n_40239;
wire n_40240;
wire n_40241;
wire n_40242;
wire n_40243;
wire n_40244;
wire n_40245;
wire n_40246;
wire n_40247;
wire n_40248;
wire n_40249;
wire n_40250;
wire n_40251;
wire n_40252;
wire n_40253;
wire n_40254;
wire n_40255;
wire n_40256;
wire n_40257;
wire n_40258;
wire n_40259;
wire n_40260;
wire n_40261;
wire n_40262;
wire n_40263;
wire n_40264;
wire n_40265;
wire n_40266;
wire n_40267;
wire n_40268;
wire n_40269;
wire n_40270;
wire n_40271;
wire n_40272;
wire n_40273;
wire n_40274;
wire n_40275;
wire n_40276;
wire n_40277;
wire n_40278;
wire n_40279;
wire n_40280;
wire n_40281;
wire n_40282;
wire n_40283;
wire n_40284;
wire n_40285;
wire n_40286;
wire n_40287;
wire n_40288;
wire n_40289;
wire n_40290;
wire n_40291;
wire n_40292;
wire n_40293;
wire n_40294;
wire n_40295;
wire n_40296;
wire n_40297;
wire n_40298;
wire n_40299;
wire n_40300;
wire n_40301;
wire n_40302;
wire n_40303;
wire n_40304;
wire n_40305;
wire n_40306;
wire n_40307;
wire n_40308;
wire n_40309;
wire n_40310;
wire n_40311;
wire n_40312;
wire n_40313;
wire n_40314;
wire n_40315;
wire n_40316;
wire n_40317;
wire n_40318;
wire n_40319;
wire n_40320;
wire n_40321;
wire n_40322;
wire n_40323;
wire n_40324;
wire n_40325;
wire n_40326;
wire n_40327;
wire n_40328;
wire n_40329;
wire n_40330;
wire n_40331;
wire n_40332;
wire n_40333;
wire n_40334;
wire n_40335;
wire n_40336;
wire n_40337;
wire n_40338;
wire n_40339;
wire n_40340;
wire n_40341;
wire n_40342;
wire n_40343;
wire n_40344;
wire n_40345;
wire n_40346;
wire n_40347;
wire n_40348;
wire n_40349;
wire n_40350;
wire n_40351;
wire n_40352;
wire n_40353;
wire n_40354;
wire n_40355;
wire n_40356;
wire n_40357;
wire n_40358;
wire n_40359;
wire n_40360;
wire n_40361;
wire n_40362;
wire n_40363;
wire n_40364;
wire n_40365;
wire n_40366;
wire n_40367;
wire n_40368;
wire n_40369;
wire n_40370;
wire n_40371;
wire n_40372;
wire n_40373;
wire n_40374;
wire n_40375;
wire n_40376;
wire n_40377;
wire n_40378;
wire n_40379;
wire n_40380;
wire n_40381;
wire n_40382;
wire n_40383;
wire n_40384;
wire n_40385;
wire n_40386;
wire n_40387;
wire n_40388;
wire n_40389;
wire n_40390;
wire n_40391;
wire n_40392;
wire n_40393;
wire n_40394;
wire n_40395;
wire n_40396;
wire n_40397;
wire n_40398;
wire n_40399;
wire n_40400;
wire n_40401;
wire n_40402;
wire n_40403;
wire n_40404;
wire n_40405;
wire n_40406;
wire n_40407;
wire n_40408;
wire n_40409;
wire n_40410;
wire n_40411;
wire n_40412;
wire n_40413;
wire n_40414;
wire n_40415;
wire n_40416;
wire n_40417;
wire n_40418;
wire n_40419;
wire n_40420;
wire n_40421;
wire n_40422;
wire n_40423;
wire n_40424;
wire n_40425;
wire n_40426;
wire n_40427;
wire n_40428;
wire n_40429;
wire n_40430;
wire n_40431;
wire n_40432;
wire n_40433;
wire n_40434;
wire n_40435;
wire n_40436;
wire n_40437;
wire n_40438;
wire n_40439;
wire n_40440;
wire n_40441;
wire n_40442;
wire n_40443;
wire n_40444;
wire n_40445;
wire n_40446;
wire n_40447;
wire n_40448;
wire n_40449;
wire n_40450;
wire n_40451;
wire n_40452;
wire n_40453;
wire n_40454;
wire n_40455;
wire n_40456;
wire n_40457;
wire n_40458;
wire n_40459;
wire n_40460;
wire n_40461;
wire n_40462;
wire n_40463;
wire n_40464;
wire n_40465;
wire n_40466;
wire n_40467;
wire n_40468;
wire n_40469;
wire n_40470;
wire n_40471;
wire n_40472;
wire n_40473;
wire n_40474;
wire n_40475;
wire n_40476;
wire n_40477;
wire n_40478;
wire n_40479;
wire n_40480;
wire n_40481;
wire n_40482;
wire n_40483;
wire n_40484;
wire n_40485;
wire n_40486;
wire n_40487;
wire n_40488;
wire n_40489;
wire n_40490;
wire n_40491;
wire n_40492;
wire n_40493;
wire n_40494;
wire n_40495;
wire n_40496;
wire n_40497;
wire n_40498;
wire n_40499;
wire n_40500;
wire n_40501;
wire n_40502;
wire n_40503;
wire n_40504;
wire n_40505;
wire n_40506;
wire n_40507;
wire n_40508;
wire n_40509;
wire n_40510;
wire n_40511;
wire n_40512;
wire n_40513;
wire n_40514;
wire n_40515;
wire n_40516;
wire n_40517;
wire n_40518;
wire n_40519;
wire n_40520;
wire n_40521;
wire n_40522;
wire n_40523;
wire n_40524;
wire n_40525;
wire n_40526;
wire n_40527;
wire n_40528;
wire n_40529;
wire n_40530;
wire n_40531;
wire n_40532;
wire n_40533;
wire n_40534;
wire n_40535;
wire n_40536;
wire n_40537;
wire n_40538;
wire n_40539;
wire n_40540;
wire n_40541;
wire n_40542;
wire n_40543;
wire n_40544;
wire n_40545;
wire n_40546;
wire n_40547;
wire n_40548;
wire n_40549;
wire n_40550;
wire n_40551;
wire n_40552;
wire n_40553;
wire n_40554;
wire n_40555;
wire n_40556;
wire n_40557;
wire n_40558;
wire n_40559;
wire n_40560;
wire n_40561;
wire n_40562;
wire n_40563;
wire n_40564;
wire n_40565;
wire n_40566;
wire n_40567;
wire n_40568;
wire n_40569;
wire n_40570;
wire n_40571;
wire n_40572;
wire n_40573;
wire n_40574;
wire n_40575;
wire n_40576;
wire n_40577;
wire n_40578;
wire n_40579;
wire n_40580;
wire n_40581;
wire n_40582;
wire n_40583;
wire n_40584;
wire n_40585;
wire n_40586;
wire n_40587;
wire n_40588;
wire n_40589;
wire n_40590;
wire n_40591;
wire n_40592;
wire n_40593;
wire n_40594;
wire n_40595;
wire n_40596;
wire n_40597;
wire n_40598;
wire n_40599;
wire n_40600;
wire n_40601;
wire n_40602;
wire n_40603;
wire n_40604;
wire n_40605;
wire n_40606;
wire n_40607;
wire n_40608;
wire n_40609;
wire n_40610;
wire n_40611;
wire n_40612;
wire n_40613;
wire n_40614;
wire n_40615;
wire n_40616;
wire n_40617;
wire n_40618;
wire n_40619;
wire n_40620;
wire n_40621;
wire n_40622;
wire n_40623;
wire n_40624;
wire n_40625;
wire n_40626;
wire n_40627;
wire n_40628;
wire n_40629;
wire n_40630;
wire n_40631;
wire n_40632;
wire n_40633;
wire n_40634;
wire n_40635;
wire n_40636;
wire n_40637;
wire n_40638;
wire n_40639;
wire n_40640;
wire n_40641;
wire n_40642;
wire n_40643;
wire n_40644;
wire n_40645;
wire n_40646;
wire n_40647;
wire n_40648;
wire n_40649;
wire n_40650;
wire n_40651;
wire n_40652;
wire n_40653;
wire n_40654;
wire n_40655;
wire n_40656;
wire n_40657;
wire n_40658;
wire n_40659;
wire n_40660;
wire n_40661;
wire n_40662;
wire n_40663;
wire n_40664;
wire n_40665;
wire n_40666;
wire n_40667;
wire n_40668;
wire n_40669;
wire n_40670;
wire n_40671;
wire n_40672;
wire n_40673;
wire n_40674;
wire n_40675;
wire n_40676;
wire n_40677;
wire n_40678;
wire n_40679;
wire n_40680;
wire n_40681;
wire n_40682;
wire n_40683;
wire n_40684;
wire n_40685;
wire n_40686;
wire n_40687;
wire n_40688;
wire n_40689;
wire n_40690;
wire n_40691;
wire n_40692;
wire n_40693;
wire n_40694;
wire n_40695;
wire n_40696;
wire n_40697;
wire n_40698;
wire n_40699;
wire n_40700;
wire n_40701;
wire n_40702;
wire n_40703;
wire n_40704;
wire n_40705;
wire n_40706;
wire n_40707;
wire n_40708;
wire n_40709;
wire n_40710;
wire n_40711;
wire n_40712;
wire n_40713;
wire n_40714;
wire n_40715;
wire n_40716;
wire n_40717;
wire n_40718;
wire n_40719;
wire n_40720;
wire n_40721;
wire n_40722;
wire n_40723;
wire n_40724;
wire n_40725;
wire n_40726;
wire n_40727;
wire n_40728;
wire n_40729;
wire n_40730;
wire n_40731;
wire n_40732;
wire n_40733;
wire n_40734;
wire n_40735;
wire n_40736;
wire n_40737;
wire n_40738;
wire n_40739;
wire n_40740;
wire n_40741;
wire n_40742;
wire n_40743;
wire n_40744;
wire n_40745;
wire n_40746;
wire n_40747;
wire n_40748;
wire n_40749;
wire n_40750;
wire n_40751;
wire n_40752;
wire n_40753;
wire n_40754;
wire n_40755;
wire n_40756;
wire n_40757;
wire n_40758;
wire n_40759;
wire n_40760;
wire n_40761;
wire n_40762;
wire n_40763;
wire n_40764;
wire n_40765;
wire n_40766;
wire n_40767;
wire n_40768;
wire n_40769;
wire n_40770;
wire n_40771;
wire n_40772;
wire n_40773;
wire n_40774;
wire n_40775;
wire n_40776;
wire n_40777;
wire n_40778;
wire n_40779;
wire n_40780;
wire n_40781;
wire n_40782;
wire n_40783;
wire n_40784;
wire n_40785;
wire n_40786;
wire n_40787;
wire n_40788;
wire n_40789;
wire n_40790;
wire n_40791;
wire n_40792;
wire n_40793;
wire n_40794;
wire n_40795;
wire n_40796;
wire n_40797;
wire n_40798;
wire n_40799;
wire n_40800;
wire n_40801;
wire n_40802;
wire n_40803;
wire n_40804;
wire n_40805;
wire n_40806;
wire n_40807;
wire n_40808;
wire n_40809;
wire n_40810;
wire n_40811;
wire n_40812;
wire n_40813;
wire n_40814;
wire n_40815;
wire n_40816;
wire n_40817;
wire n_40818;
wire n_40819;
wire n_40820;
wire n_40821;
wire n_40822;
wire n_40823;
wire n_40824;
wire n_40825;
wire n_40826;
wire n_40827;
wire n_40828;
wire n_40829;
wire n_40830;
wire n_40831;
wire n_40832;
wire n_40833;
wire n_40834;
wire n_40835;
wire n_40836;
wire n_40837;
wire n_40838;
wire n_40839;
wire n_40840;
wire n_40841;
wire n_40842;
wire n_40843;
wire n_40844;
wire n_40845;
wire n_40846;
wire n_40847;
wire n_40848;
wire n_40849;
wire n_40850;
wire n_40851;
wire n_40852;
wire n_40853;
wire n_40854;
wire n_40855;
wire n_40856;
wire n_40857;
wire n_40858;
wire n_40859;
wire n_40860;
wire n_40861;
wire n_40862;
wire n_40863;
wire n_40864;
wire n_40865;
wire n_40866;
wire n_40867;
wire n_40868;
wire n_40869;
wire n_40870;
wire n_40871;
wire n_40872;
wire n_40873;
wire n_40874;
wire n_40875;
wire n_40876;
wire n_40877;
wire n_40878;
wire n_40879;
wire n_40880;
wire n_40881;
wire n_40882;
wire n_40883;
wire n_40884;
wire n_40885;
wire n_40886;
wire n_40887;
wire n_40888;
wire n_40889;
wire n_40890;
wire n_40891;
wire n_40892;
wire n_40893;
wire n_40894;
wire n_40895;
wire n_40896;
wire n_40897;
wire n_40898;
wire n_40899;
wire n_40900;
wire n_40901;
wire n_40902;
wire n_40903;
wire n_40904;
wire n_40905;
wire n_40906;
wire n_40907;
wire n_40908;
wire n_40909;
wire n_40910;
wire n_40911;
wire n_40912;
wire n_40913;
wire n_40914;
wire n_40915;
wire n_40916;
wire n_40917;
wire n_40918;
wire n_40919;
wire n_40920;
wire n_40921;
wire n_40922;
wire n_40923;
wire n_40924;
wire n_40925;
wire n_40926;
wire n_40927;
wire n_40928;
wire n_40929;
wire n_40930;
wire n_40931;
wire n_40932;
wire n_40933;
wire n_40934;
wire n_40935;
wire n_40936;
wire n_40937;
wire n_40938;
wire n_40939;
wire n_40940;
wire n_40941;
wire n_40942;
wire n_40943;
wire n_40944;
wire n_40945;
wire n_40946;
wire n_40947;
wire n_40948;
wire n_40949;
wire n_40950;
wire n_40951;
wire n_40952;
wire n_40953;
wire n_40954;
wire n_40955;
wire n_40956;
wire n_40957;
wire n_40958;
wire n_40959;
wire n_40960;
wire n_40961;
wire n_40962;
wire n_40963;
wire n_40964;
wire n_40965;
wire n_40966;
wire n_40967;
wire n_40968;
wire n_40969;
wire n_40970;
wire n_40971;
wire n_40972;
wire n_40973;
wire n_40974;
wire n_40975;
wire n_40976;
wire n_40977;
wire n_40978;
wire n_40979;
wire n_40980;
wire n_40981;
wire n_40982;
wire n_40983;
wire n_40984;
wire n_40985;
wire n_40986;
wire n_40987;
wire n_40988;
wire n_40989;
wire n_40990;
wire n_40991;
wire n_40992;
wire n_40993;
wire n_40994;
wire n_40995;
wire n_40996;
wire n_40997;
wire n_40998;
wire n_40999;
wire n_41000;
wire n_41001;
wire n_41002;
wire n_41003;
wire n_41004;
wire n_41005;
wire n_41006;
wire n_41007;
wire n_41008;
wire n_41009;
wire n_41010;
wire n_41011;
wire n_41012;
wire n_41013;
wire n_41014;
wire n_41015;
wire n_41016;
wire n_41017;
wire n_41018;
wire n_41019;
wire n_41020;
wire n_41021;
wire n_41022;
wire n_41023;
wire n_41024;
wire n_41025;
wire n_41026;
wire n_41027;
wire n_41028;
wire n_41029;
wire n_41030;
wire n_41031;
wire n_41032;
wire n_41033;
wire n_41034;
wire n_41035;
wire n_41036;
wire n_41037;
wire n_41038;
wire n_41039;
wire n_41040;
wire n_41041;
wire n_41042;
wire n_41043;
wire n_41044;
wire n_41045;
wire n_41046;
wire n_41047;
wire n_41048;
wire n_41049;
wire n_41050;
wire n_41051;
wire n_41052;
wire n_41053;
wire n_41054;
wire n_41055;
wire n_41056;
wire n_41057;
wire n_41058;
wire n_41059;
wire n_41060;
wire n_41061;
wire n_41062;
wire n_41063;
wire n_41064;
wire n_41065;
wire n_41066;
wire n_41067;
wire n_41068;
wire n_41069;
wire n_41070;
wire n_41071;
wire n_41072;
wire n_41073;
wire n_41074;
wire n_41075;
wire n_41076;
wire n_41077;
wire n_41078;
wire n_41079;
wire n_41080;
wire n_41081;
wire n_41082;
wire n_41083;
wire n_41084;
wire n_41085;
wire n_41086;
wire n_41087;
wire n_41088;
wire n_41089;
wire n_41090;
wire n_41091;
wire n_41092;
wire n_41093;
wire n_41094;
wire n_41095;
wire n_41096;
wire n_41097;
wire n_41098;
wire n_41099;
wire n_41100;
wire n_41101;
wire n_41102;
wire n_41103;
wire n_41104;
wire n_41105;
wire n_41106;
wire n_41107;
wire n_41108;
wire n_41109;
wire n_41110;
wire n_41111;
wire n_41112;
wire n_41113;
wire n_41114;
wire n_41115;
wire n_41116;
wire n_41117;
wire n_41118;
wire n_41119;
wire n_41120;
wire n_41121;
wire n_41122;
wire n_41123;
wire n_41124;
wire n_41125;
wire n_41126;
wire n_41127;
wire n_41128;
wire n_41129;
wire n_41130;
wire n_41131;
wire n_41132;
wire n_41133;
wire n_41134;
wire n_41135;
wire n_41136;
wire n_41137;
wire n_41138;
wire n_41139;
wire n_41140;
wire n_41141;
wire n_41142;
wire n_41143;
wire n_41144;
wire n_41145;
wire n_41146;
wire n_41147;
wire n_41148;
wire n_41149;
wire n_41150;
wire n_41151;
wire n_41152;
wire n_41153;
wire n_41154;
wire n_41155;
wire n_41156;
wire n_41157;
wire n_41158;
wire n_41159;
wire n_41160;
wire n_41161;
wire n_41162;
wire n_41163;
wire n_41164;
wire n_41165;
wire n_41166;
wire n_41167;
wire n_41168;
wire n_41169;
wire n_41170;
wire n_41171;
wire n_41172;
wire n_41173;
wire n_41174;
wire n_41175;
wire n_41176;
wire n_41177;
wire n_41178;
wire n_41179;
wire n_41180;
wire n_41181;
wire n_41182;
wire n_41183;
wire n_41184;
wire n_41185;
wire n_41186;
wire n_41187;
wire n_41188;
wire n_41189;
wire n_41190;
wire n_41191;
wire n_41192;
wire n_41193;
wire n_41194;
wire n_41195;
wire n_41196;
wire n_41197;
wire n_41198;
wire n_41199;
wire n_41200;
wire n_41201;
wire n_41202;
wire n_41203;
wire n_41204;
wire n_41205;
wire n_41206;
wire n_41207;
wire n_41208;
wire n_41209;
wire n_41210;
wire n_41211;
wire n_41212;
wire n_41213;
wire n_41214;
wire n_41215;
wire n_41216;
wire n_41217;
wire n_41218;
wire n_41219;
wire n_41220;
wire n_41221;
wire n_41222;
wire n_41223;
wire n_41224;
wire n_41225;
wire n_41226;
wire n_41227;
wire n_41228;
wire n_41229;
wire n_41230;
wire n_41231;
wire n_41232;
wire n_41233;
wire n_41234;
wire n_41235;
wire n_41236;
wire n_41237;
wire n_41238;
wire n_41239;
wire n_41240;
wire n_41241;
wire n_41242;
wire n_41243;
wire n_41244;
wire n_41245;
wire n_41246;
wire n_41247;
wire n_41248;
wire n_41249;
wire n_41250;
wire n_41251;
wire n_41252;
wire n_41253;
wire n_41254;
wire n_41255;
wire n_41256;
wire n_41257;
wire n_41258;
wire n_41259;
wire n_41260;
wire n_41261;
wire n_41262;
wire n_41263;
wire n_41264;
wire n_41265;
wire n_41266;
wire n_41267;
wire n_41268;
wire n_41269;
wire n_41270;
wire n_41271;
wire n_41272;
wire n_41273;
wire n_41274;
wire n_41275;
wire n_41276;
wire n_41277;
wire n_41278;
wire n_41279;
wire n_41280;
wire n_41281;
wire n_41282;
wire n_41283;
wire n_41284;
wire n_41285;
wire n_41286;
wire n_41287;
wire n_41288;
wire n_41289;
wire n_41290;
wire n_41291;
wire n_41292;
wire n_41293;
wire n_41294;
wire n_41295;
wire n_41296;
wire n_41297;
wire n_41298;
wire n_41299;
wire n_41300;
wire n_41301;
wire n_41302;
wire n_41303;
wire n_41304;
wire n_41305;
wire n_41306;
wire n_41307;
wire n_41308;
wire n_41309;
wire n_41310;
wire n_41311;
wire n_41312;
wire n_41313;
wire n_41314;
wire n_41315;
wire n_41316;
wire n_41317;
wire n_41318;
wire n_41319;
wire n_41320;
wire n_41321;
wire n_41322;
wire n_41323;
wire n_41324;
wire n_41325;
wire n_41326;
wire n_41327;
wire n_41328;
wire n_41329;
wire n_41330;
wire n_41331;
wire n_41332;
wire n_41333;
wire n_41334;
wire n_41335;
wire n_41336;
wire n_41337;
wire n_41338;
wire n_41339;
wire n_41340;
wire n_41341;
wire n_41342;
wire n_41343;
wire n_41344;
wire n_41345;
wire n_41346;
wire n_41347;
wire n_41348;
wire n_41349;
wire n_41350;
wire n_41351;
wire n_41352;
wire n_41353;
wire n_41354;
wire n_41355;
wire n_41356;
wire n_41357;
wire n_41358;
wire n_41359;
wire n_41360;
wire n_41361;
wire n_41362;
wire n_41363;
wire n_41364;
wire n_41365;
wire n_41366;
wire n_41367;
wire n_41368;
wire n_41369;
wire n_41370;
wire n_41371;
wire n_41372;
wire n_41373;
wire n_41374;
wire n_41375;
wire n_41376;
wire n_41377;
wire n_41378;
wire n_41379;
wire n_41380;
wire n_41381;
wire n_41382;
wire n_41383;
wire n_41384;
wire n_41385;
wire n_41386;
wire n_41387;
wire n_41388;
wire n_41389;
wire n_41390;
wire n_41391;
wire n_41392;
wire n_41393;
wire n_41394;
wire n_41395;
wire n_41396;
wire n_41397;
wire n_41398;
wire n_41399;
wire n_41400;
wire n_41401;
wire n_41402;
wire n_41403;
wire n_41404;
wire n_41405;
wire n_41406;
wire n_41407;
wire n_41408;
wire n_41409;
wire n_41410;
wire n_41411;
wire n_41412;
wire n_41413;
wire n_41414;
wire n_41415;
wire n_41416;
wire n_41417;
wire n_41418;
wire n_41419;
wire n_41420;
wire n_41421;
wire n_41422;
wire n_41423;
wire n_41424;
wire n_41425;
wire n_41426;
wire n_41427;
wire n_41428;
wire n_41429;
wire n_41430;
wire n_41431;
wire n_41432;
wire n_41433;
wire n_41434;
wire n_41435;
wire n_41436;
wire n_41437;
wire n_41438;
wire n_41439;
wire n_41440;
wire n_41441;
wire n_41442;
wire n_41443;
wire n_41444;
wire n_41445;
wire n_41446;
wire n_41447;
wire n_41448;
wire n_41449;
wire n_41450;
wire n_41451;
wire n_41452;
wire n_41453;
wire n_41454;
wire n_41455;
wire n_41456;
wire n_41457;
wire n_41458;
wire n_41459;
wire n_41460;
wire n_41461;
wire n_41462;
wire n_41463;
wire n_41464;
wire n_41465;
wire n_41466;
wire n_41467;
wire n_41468;
wire n_41469;
wire n_41470;
wire n_41471;
wire n_41472;
wire n_41473;
wire n_41474;
wire n_41475;
wire n_41476;
wire n_41477;
wire n_41478;
wire n_41479;
wire n_41480;
wire n_41481;
wire n_41482;
wire n_41483;
wire n_41484;
wire n_41485;
wire n_41486;
wire n_41487;
wire n_41488;
wire n_41489;
wire n_41490;
wire n_41491;
wire n_41492;
wire n_41493;
wire n_41494;
wire n_41495;
wire n_41496;
wire n_41497;
wire n_41498;
wire n_41499;
wire n_41500;
wire n_41501;
wire n_41502;
wire n_41503;
wire n_41504;
wire n_41505;
wire n_41506;
wire n_41507;
wire n_41508;
wire n_41509;
wire n_41510;
wire n_41511;
wire n_41512;
wire n_41513;
wire n_41514;
wire n_41515;
wire n_41516;
wire n_41517;
wire n_41518;
wire n_41519;
wire n_41520;
wire n_41521;
wire n_41522;
wire n_41523;
wire n_41524;
wire n_41525;
wire n_41526;
wire n_41527;
wire n_41528;
wire n_41529;
wire n_41530;
wire n_41531;
wire n_41532;
wire n_41533;
wire n_41534;
wire n_41535;
wire n_41536;
wire n_41537;
wire n_41538;
wire n_41539;
wire n_41540;
wire n_41541;
wire n_41542;
wire n_41543;
wire n_41544;
wire n_41545;
wire n_41546;
wire n_41547;
wire n_41548;
wire n_41549;
wire n_41550;
wire n_41551;
wire n_41552;
wire n_41553;
wire n_41554;
wire n_41555;
wire n_41556;
wire n_41557;
wire n_41558;
wire n_41559;
wire n_41560;
wire n_41561;
wire n_41562;
wire n_41563;
wire n_41564;
wire n_41565;
wire n_41566;
wire n_41567;
wire n_41568;
wire n_41569;
wire n_41570;
wire n_41571;
wire n_41572;
wire n_41573;
wire n_41574;
wire n_41575;
wire n_41576;
wire n_41577;
wire n_41578;
wire n_41579;
wire n_41580;
wire n_41581;
wire n_41582;
wire n_41583;
wire n_41584;
wire n_41585;
wire n_41586;
wire n_41587;
wire n_41588;
wire n_41589;
wire n_41590;
wire n_41591;
wire n_41592;
wire n_41593;
wire n_41594;
wire n_41595;
wire n_41596;
wire n_41597;
wire n_41598;
wire n_41599;
wire n_41600;
wire n_41601;
wire n_41602;
wire n_41603;
wire n_41604;
wire n_41605;
wire n_41606;
wire n_41607;
wire n_41608;
wire n_41609;
wire n_41610;
wire n_41611;
wire n_41612;
wire n_41613;
wire n_41614;
wire n_41615;
wire n_41616;
wire n_41617;
wire n_41618;
wire n_41619;
wire n_41620;
wire n_41621;
wire n_41622;
wire n_41623;
wire n_41624;
wire n_41625;
wire n_41626;
wire n_41627;
wire n_41628;
wire n_41629;
wire n_41630;
wire n_41631;
wire n_41632;
wire n_41633;
wire n_41634;
wire n_41635;
wire n_41636;
wire n_41637;
wire n_41638;
wire n_41639;
wire n_41640;
wire n_41641;
wire n_41642;
wire n_41643;
wire n_41644;
wire n_41645;
wire n_41646;
wire n_41647;
wire n_41648;
wire n_41649;
wire n_41650;
wire n_41651;
wire n_41652;
wire n_41653;
wire n_41654;
wire n_41655;
wire n_41656;
wire n_41657;
wire n_41658;
wire n_41659;
wire n_41660;
wire n_41661;
wire n_41662;
wire n_41663;
wire n_41664;
wire n_41665;
wire n_41666;
wire n_41667;
wire n_41668;
wire n_41669;
wire n_41670;
wire n_41671;
wire n_41672;
wire n_41673;
wire n_41674;
wire n_41675;
wire n_41676;
wire n_41677;
wire n_41678;
wire n_41679;
wire n_41680;
wire n_41681;
wire n_41682;
wire n_41683;
wire n_41684;
wire n_41685;
wire n_41686;
wire n_41687;
wire n_41688;
wire n_41689;
wire n_41690;
wire n_41691;
wire n_41692;
wire n_41693;
wire n_41694;
wire n_41695;
wire n_41696;
wire n_41697;
wire n_41698;
wire n_41699;
wire n_41700;
wire n_41701;
wire n_41702;
wire n_41703;
wire n_41704;
wire n_41705;
wire n_41706;
wire n_41707;
wire n_41708;
wire n_41709;
wire n_41710;
wire n_41711;
wire n_41712;
wire n_41713;
wire n_41714;
wire n_41715;
wire n_41716;
wire n_41717;
wire n_41718;
wire n_41719;
wire n_41720;
wire n_41721;
wire n_41722;
wire n_41723;
wire n_41724;
wire n_41725;
wire n_41726;
wire n_41727;
wire n_41728;
wire n_41729;
wire n_41730;
wire n_41731;
wire n_41732;
wire n_41733;
wire n_41734;
wire n_41735;
wire n_41736;
wire n_41737;
wire n_41738;
wire n_41739;
wire n_41740;
wire n_41741;
wire n_41742;
wire n_41743;
wire n_41744;
wire n_41745;
wire n_41746;
wire n_41747;
wire n_41748;
wire n_41749;
wire n_41750;
wire n_41751;
wire n_41752;
wire n_41753;
wire n_41754;
wire n_41755;
wire n_41756;
wire n_41757;
wire n_41758;
wire n_41759;
wire n_41760;
wire n_41761;
wire n_41762;
wire n_41763;
wire n_41764;
wire n_41765;
wire n_41766;
wire n_41767;
wire n_41768;
wire n_41769;
wire n_41770;
wire n_41771;
wire n_41772;
wire n_41773;
wire n_41774;
wire n_41775;
wire n_41776;
wire n_41777;
wire n_41778;
wire n_41779;
wire n_41780;
wire n_41781;
wire n_41782;
wire n_41783;
wire n_41784;
wire n_41785;
wire n_41786;
wire n_41787;
wire n_41788;
wire n_41789;
wire n_41790;
wire n_41791;
wire n_41792;
wire n_41793;
wire n_41794;
wire n_41795;
wire n_41796;
wire n_41797;
wire n_41798;
wire n_41799;
wire n_41800;
wire n_41801;
wire n_41802;
wire n_41803;
wire n_41804;
wire n_41805;
wire n_41806;
wire n_41807;
wire n_41808;
wire n_41809;
wire n_41810;
wire n_41811;
wire n_41812;
wire n_41813;
wire n_41814;
wire n_41815;
wire n_41816;
wire n_41817;
wire n_41818;
wire n_41819;
wire n_41820;
wire n_41821;
wire n_41822;
wire n_41823;
wire n_41824;
wire n_41825;
wire n_41826;
wire n_41827;
wire n_41828;
wire n_41829;
wire n_41830;
wire n_41831;
wire n_41832;
wire n_41833;
wire n_41834;
wire n_41835;
wire n_41836;
wire n_41837;
wire n_41838;
wire n_41839;
wire n_41840;
wire n_41841;
wire n_41842;
wire n_41843;
wire n_41844;
wire n_41845;
wire n_41846;
wire n_41847;
wire n_41848;
wire n_41849;
wire n_41850;
wire n_41851;
wire n_41852;
wire n_41853;
wire n_41854;
wire n_41855;
wire n_41856;
wire n_41857;
wire n_41858;
wire n_41859;
wire n_41860;
wire n_41861;
wire n_41862;
wire n_41863;
wire n_41864;
wire n_41865;
wire n_41866;
wire n_41867;
wire n_41868;
wire n_41869;
wire n_41870;
wire n_41871;
wire n_41872;
wire n_41873;
wire n_41874;
wire n_41875;
wire n_41876;
wire n_41877;
wire n_41878;
wire n_41879;
wire n_41880;
wire n_41881;
wire n_41882;
wire n_41883;
wire n_41884;
wire n_41885;
wire n_41886;
wire n_41887;
wire n_41888;
wire n_41889;
wire n_41890;
wire n_41891;
wire n_41892;
wire n_41893;
wire n_41894;
wire n_41895;
wire n_41896;
wire n_41897;
wire n_41898;
wire n_41899;
wire n_41900;
wire n_41901;
wire n_41902;
wire n_41903;
wire n_41904;
wire n_41905;
wire n_41906;
wire n_41907;
wire n_41908;
wire n_41909;
wire n_41910;
wire n_41911;
wire n_41912;
wire n_41913;
wire n_41914;
wire n_41915;
wire n_41916;
wire n_41917;
wire n_41918;
wire n_41919;
wire n_41920;
wire n_41921;
wire n_41922;
wire n_41923;
wire n_41924;
wire n_41925;
wire n_41926;
wire n_41927;
wire n_41928;
wire n_41929;
wire n_41930;
wire n_41931;
wire n_41932;
wire n_41933;
wire n_41934;
wire n_41935;
wire n_41936;
wire n_41937;
wire n_41938;
wire n_41939;
wire n_41940;
wire n_41941;
wire n_41942;
wire n_41943;
wire n_41944;
wire n_41945;
wire n_41946;
wire n_41947;
wire n_41948;
wire n_41949;
wire n_41950;
wire n_41951;
wire n_41952;
wire n_41953;
wire n_41954;
wire n_41955;
wire n_41956;
wire n_41957;
wire n_41958;
wire n_41959;
wire n_41960;
wire n_41961;
wire n_41962;
wire n_41963;
wire n_41964;
wire n_41965;
wire n_41966;
wire n_41967;
wire n_41968;
wire n_41969;
wire n_41970;
wire n_41971;
wire n_41972;
wire n_41973;
wire n_41974;
wire n_41975;
wire n_41976;
wire n_41977;
wire n_41978;
wire n_41979;
wire n_41980;
wire n_41981;
wire n_41982;
wire n_41983;
wire n_41984;
wire n_41985;
wire n_41986;
wire n_41987;
wire n_41988;
wire n_41989;
wire n_41990;
wire n_41991;
wire n_41992;
wire n_41993;
wire n_41994;
wire n_41995;
wire n_41996;
wire n_41997;
wire n_41998;
wire n_41999;
wire n_42000;
wire n_42001;
wire n_42002;
wire n_42003;
wire n_42004;
wire n_42005;
wire n_42006;
wire n_42007;
wire n_42008;
wire n_42009;
wire n_42010;
wire n_42011;
wire n_42012;
wire n_42013;
wire n_42014;
wire n_42015;
wire n_42016;
wire n_42017;
wire n_42018;
wire n_42019;
wire n_42020;
wire n_42021;
wire n_42022;
wire n_42023;
wire n_42024;
wire n_42025;
wire n_42026;
wire n_42027;
wire n_42028;
wire n_42029;
wire n_42030;
wire n_42031;
wire n_42032;
wire n_42033;
wire n_42034;
wire n_42035;
wire n_42036;
wire n_42037;
wire n_42038;
wire n_42039;
wire n_42040;
wire n_42041;
wire n_42042;
wire n_42043;
wire n_42044;
wire n_42045;
wire n_42046;
wire n_42047;
wire n_42048;
wire n_42049;
wire n_42050;
wire n_42051;
wire n_42052;
wire n_42053;
wire n_42054;
wire n_42055;
wire n_42056;
wire n_42057;
wire n_42058;
wire n_42059;
wire n_42060;
wire n_42061;
wire n_42062;
wire n_42063;
wire n_42064;
wire n_42065;
wire n_42066;
wire n_42067;
wire n_42068;
wire n_42069;
wire n_42070;
wire n_42071;
wire n_42072;
wire n_42073;
wire n_42074;
wire n_42075;
wire n_42076;
wire n_42077;
wire n_42078;
wire n_42079;
wire n_42080;
wire n_42081;
wire n_42082;
wire n_42083;
wire n_42084;
wire n_42085;
wire n_42086;
wire n_42087;
wire n_42088;
wire n_42089;
wire n_42090;
wire n_42091;
wire n_42092;
wire n_42093;
wire n_42094;
wire n_42095;
wire n_42096;
wire n_42097;
wire n_42098;
wire n_42099;
wire n_42100;
wire n_42101;
wire n_42102;
wire n_42103;
wire n_42104;
wire n_42105;
wire n_42106;
wire n_42107;
wire n_42108;
wire n_42109;
wire n_42110;
wire n_42111;
wire n_42112;
wire n_42113;
wire n_42114;
wire n_42115;
wire n_42116;
wire n_42117;
wire n_42118;
wire n_42119;
wire n_42120;
wire n_42121;
wire n_42122;
wire n_42123;
wire n_42124;
wire n_42125;
wire n_42126;
wire n_42127;
wire n_42128;
wire n_42129;
wire n_42130;
wire n_42131;
wire n_42132;
wire n_42133;
wire n_42134;
wire n_42135;
wire n_42136;
wire n_42137;
wire n_42138;
wire n_42139;
wire n_42140;
wire n_42141;
wire n_42142;
wire n_42143;
wire n_42144;
wire n_42145;
wire n_42146;
wire n_42147;
wire n_42148;
wire n_42149;
wire n_42150;
wire n_42151;
wire n_42152;
wire n_42153;
wire n_42154;
wire n_42155;
wire n_42156;
wire n_42157;
wire n_42158;
wire n_42159;
wire n_42160;
wire n_42161;
wire n_42162;
wire n_42163;
wire n_42164;
wire n_42165;
wire n_42166;
wire n_42167;
wire n_42168;
wire n_42169;
wire n_42170;
wire n_42171;
wire n_42172;
wire n_42173;
wire n_42174;
wire n_42175;
wire n_42176;
wire n_42177;
wire n_42178;
wire n_42179;
wire n_42180;
wire n_42181;
wire n_42182;
wire n_42183;
wire n_42184;
wire n_42185;
wire n_42186;
wire n_42187;
wire n_42188;
wire n_42189;
wire n_42190;
wire n_42191;
wire n_42192;
wire n_42193;
wire n_42194;
wire n_42195;
wire n_42196;
wire n_42197;
wire n_42198;
wire n_42199;
wire n_42200;
wire n_42201;
wire n_42202;
wire n_42203;
wire n_42204;
wire n_42205;
wire n_42206;
wire n_42207;
wire n_42208;
wire n_42209;
wire n_42210;
wire n_42211;
wire n_42212;
wire n_42213;
wire n_42214;
wire n_42215;
wire n_42216;
wire n_42217;
wire n_42218;
wire n_42219;
wire n_42220;
wire n_42221;
wire n_42222;
wire n_42223;
wire n_42224;
wire n_42225;
wire n_42226;
wire n_42227;
wire n_42228;
wire n_42229;
wire n_42230;
wire n_42231;
wire n_42232;
wire n_42233;
wire n_42234;
wire n_42235;
wire n_42236;
wire n_42237;
wire n_42238;
wire n_42239;
wire n_42240;
wire n_42241;
wire n_42242;
wire n_42243;
wire n_42244;
wire n_42245;
wire n_42246;
wire n_42247;
wire n_42248;
wire n_42249;
wire n_42250;
wire n_42251;
wire n_42252;
wire n_42253;
wire n_42254;
wire n_42255;
wire n_42256;
wire n_42257;
wire n_42258;
wire n_42259;
wire n_42260;
wire n_42261;
wire n_42262;
wire n_42263;
wire n_42264;
wire n_42265;
wire n_42266;
wire n_42267;
wire n_42268;
wire n_42269;
wire n_42270;
wire n_42271;
wire n_42272;
wire n_42273;
wire n_42274;
wire n_42275;
wire n_42276;
wire n_42277;
wire n_42278;
wire n_42279;
wire n_42280;
wire n_42281;
wire n_42282;
wire n_42283;
wire n_42284;
wire n_42285;
wire n_42286;
wire n_42287;
wire n_42288;
wire n_42289;
wire n_42290;
wire n_42291;
wire n_42292;
wire n_42293;
wire n_42294;
wire n_42295;
wire n_42296;
wire n_42297;
wire n_42298;
wire n_42299;
wire n_42300;
wire n_42301;
wire n_42302;
wire n_42303;
wire n_42304;
wire n_42305;
wire n_42306;
wire n_42307;
wire n_42308;
wire n_42309;
wire n_42310;
wire n_42311;
wire n_42312;
wire n_42313;
wire n_42314;
wire n_42315;
wire n_42316;
wire n_42317;
wire n_42318;
wire n_42319;
wire n_42320;
wire n_42321;
wire n_42322;
wire n_42323;
wire n_42324;
wire n_42325;
wire n_42326;
wire n_42327;
wire n_42328;
wire n_42329;
wire n_42330;
wire n_42331;
wire n_42332;
wire n_42333;
wire n_42334;
wire n_42335;
wire n_42336;
wire n_42337;
wire n_42338;
wire n_42339;
wire n_42340;
wire n_42341;
wire n_42342;
wire n_42343;
wire n_42344;
wire n_42345;
wire n_42346;
wire n_42347;
wire n_42348;
wire n_42349;
wire n_42350;
wire n_42351;
wire n_42352;
wire n_42353;
wire n_42354;
wire n_42355;
wire n_42356;
wire n_42357;
wire n_42358;
wire n_42359;
wire n_42360;
wire n_42361;
wire n_42362;
wire n_42363;
wire n_42364;
wire n_42365;
wire n_42366;
wire n_42367;
wire n_42368;
wire n_42369;
wire n_42370;
wire n_42371;
wire n_42372;
wire n_42373;
wire n_42374;
wire n_42375;
wire n_42376;
wire n_42377;
wire n_42378;
wire n_42379;
wire n_42380;
wire n_42381;
wire n_42382;
wire n_42383;
wire n_42384;
wire n_42385;
wire n_42386;
wire n_42387;
wire n_42388;
wire n_42389;
wire n_42390;
wire n_42391;
wire n_42392;
wire n_42393;
wire n_42394;
wire n_42395;
wire n_42396;
wire n_42397;
wire n_42398;
wire n_42399;
wire n_42400;
wire n_42401;
wire n_42402;
wire n_42403;
wire n_42404;
wire n_42405;
wire n_42406;
wire n_42407;
wire n_42408;
wire n_42409;
wire n_42410;
wire n_42411;
wire n_42412;
wire n_42413;
wire n_42414;
wire n_42415;
wire n_42416;
wire n_42417;
wire n_42418;
wire n_42419;
wire n_42420;
wire n_42421;
wire n_42422;
wire n_42423;
wire n_42424;
wire n_42425;
wire n_42426;
wire n_42427;
wire n_42428;
wire n_42429;
wire n_42430;
wire n_42431;
wire n_42432;
wire n_42433;
wire n_42434;
wire n_42435;
wire n_42436;
wire n_42437;
wire n_42438;
wire n_42439;
wire n_42440;
wire n_42441;
wire n_42442;
wire n_42443;
wire n_42444;
wire n_42445;
wire n_42446;
wire n_42447;
wire n_42448;
wire n_42449;
wire n_42450;
wire n_42451;
wire n_42452;
wire n_42453;
wire n_42454;
wire n_42455;
wire n_42456;
wire n_42457;
wire n_42458;
wire n_42459;
wire n_42460;
wire n_42461;
wire n_42462;
wire n_42463;
wire n_42464;
wire n_42465;
wire n_42466;
wire n_42467;
wire n_42468;
wire n_42469;
wire n_42470;
wire n_42471;
wire n_42472;
wire n_42473;
wire n_42474;
wire n_42475;
wire n_42476;
wire n_42477;
wire n_42478;
wire n_42479;
wire n_42480;
wire n_42481;
wire n_42482;
wire n_42483;
wire n_42484;
wire n_42485;
wire n_42486;
wire n_42487;
wire n_42488;
wire n_42489;
wire n_42490;
wire n_42491;
wire n_42492;
wire n_42493;
wire n_42494;
wire n_42495;
wire n_42496;
wire n_42497;
wire n_42498;
wire n_42499;
wire n_42500;
wire n_42501;
wire n_42502;
wire n_42503;
wire n_42504;
wire n_42505;
wire n_42506;
wire n_42507;
wire n_42508;
wire n_42509;
wire n_42510;
wire n_42511;
wire n_42512;
wire n_42513;
wire n_42514;
wire n_42515;
wire n_42516;
wire n_42517;
wire n_42518;
wire n_42519;
wire n_42520;
wire n_42521;
wire n_42522;
wire n_42523;
wire n_42524;
wire n_42525;
wire n_42526;
wire n_42527;
wire n_42528;
wire n_42529;
wire n_42530;
wire n_42531;
wire n_42532;
wire n_42533;
wire n_42534;
wire n_42535;
wire n_42536;
wire n_42537;
wire n_42538;
wire n_42539;
wire n_42540;
wire n_42541;
wire n_42542;
wire n_42543;
wire n_42544;
wire n_42545;
wire n_42546;
wire n_42547;
wire n_42548;
wire n_42549;
wire n_42550;
wire n_42551;
wire n_42552;
wire n_42553;
wire n_42554;
wire n_42555;
wire n_42556;
wire n_42557;
wire n_42558;
wire n_42559;
wire n_42560;
wire n_42561;
wire n_42562;
wire n_42563;
wire n_42564;
wire n_42565;
wire n_42566;
wire n_42567;
wire n_42568;
wire n_42569;
wire n_42570;
wire n_42571;
wire n_42572;
wire n_42573;
wire n_42574;
wire n_42575;
wire n_42576;
wire n_42577;
wire n_42578;
wire n_42579;
wire n_42580;
wire n_42581;
wire n_42582;
wire n_42583;
wire n_42584;
wire n_42585;
wire n_42586;
wire n_42587;
wire n_42588;
wire n_42589;
wire n_42590;
wire n_42591;
wire n_42592;
wire n_42593;
wire n_42594;
wire n_42595;
wire n_42596;
wire n_42597;
wire n_42598;
wire n_42599;
wire n_42600;
wire n_42601;
wire n_42602;
wire n_42603;
wire n_42604;
wire n_42605;
wire n_42606;
wire n_42607;
wire n_42608;
wire n_42609;
wire n_42610;
wire n_42611;
wire n_42612;
wire n_42613;
wire n_42614;
wire n_42615;
wire n_42616;
wire n_42617;
wire n_42618;
wire n_42619;
wire n_42620;
wire n_42621;
wire n_42622;
wire n_42623;
wire n_42624;
wire n_42625;
wire n_42626;
wire n_42627;
wire n_42628;
wire n_42629;
wire n_42630;
wire n_42631;
wire n_42632;
wire n_42633;
wire n_42634;
wire n_42635;
wire n_42636;
wire n_42637;
wire n_42638;
wire n_42639;
wire n_42640;
wire n_42641;
wire n_42642;
wire n_42643;
wire n_42644;
wire n_42645;
wire n_42646;
wire n_42647;
wire n_42648;
wire n_42649;
wire n_42650;
wire n_42651;
wire n_42652;
wire n_42653;
wire n_42654;
wire n_42655;
wire n_42656;
wire n_42657;
wire n_42658;
wire n_42659;
wire n_42660;
wire n_42661;
wire n_42662;
wire n_42663;
wire n_42664;
wire n_42665;
wire n_42666;
wire n_42667;
wire n_42668;
wire n_42669;
wire n_42670;
wire n_42671;
wire n_42672;
wire n_42673;
wire n_42674;
wire n_42675;
wire n_42676;
wire n_42677;
wire n_42678;
wire n_42679;
wire n_42680;
wire n_42681;
wire n_42682;
wire n_42683;
wire n_42684;
wire n_42685;
wire n_42686;
wire n_42687;
wire n_42688;
wire n_42689;
wire n_42690;
wire n_42691;
wire n_42692;
wire n_42693;
wire n_42694;
wire n_42695;
wire n_42696;
wire n_42697;
wire n_42698;
wire n_42699;
wire n_42700;
wire n_42701;
wire n_42702;
wire n_42703;
wire n_42704;
wire n_42705;
wire n_42706;
wire n_42707;
wire n_42708;
wire n_42709;
wire n_42710;
wire n_42711;
wire n_42712;
wire n_42713;
wire n_42714;
wire n_42715;
wire n_42716;
wire n_42717;
wire n_42718;
wire n_42719;
wire n_42720;
wire n_42721;
wire n_42722;
wire n_42723;
wire n_42724;
wire n_42725;
wire n_42726;
wire n_42727;
wire n_42728;
wire n_42729;
wire n_42730;
wire n_42731;
wire n_42732;
wire n_42733;
wire n_42734;
wire n_42735;
wire n_42736;
wire n_42737;
wire n_42738;
wire n_42739;
wire n_42740;
wire n_42741;
wire n_42742;
wire n_42743;
wire n_42744;
wire n_42745;
wire n_42746;
wire n_42747;
wire n_42748;
wire n_42749;
wire n_42750;
wire n_42751;
wire n_42752;
wire n_42753;
wire n_42754;
wire n_42755;
wire n_42756;
wire n_42757;
wire n_42758;
wire n_42759;
wire n_42760;
wire n_42761;
wire n_42762;
wire n_42763;
wire n_42764;
wire n_42765;
wire n_42766;
wire n_42767;
wire n_42768;
wire n_42769;
wire n_42770;
wire n_42771;
wire n_42772;
wire n_42773;
wire n_42774;
wire n_42775;
wire n_42776;
wire n_42777;
wire n_42778;
wire n_42779;
wire n_42780;
wire n_42781;
wire n_42782;
wire n_42783;
wire n_42784;
wire n_42785;
wire n_42786;
wire n_42787;
wire n_42788;
wire n_42789;
wire n_42790;
wire n_42791;
wire n_42792;
wire n_42793;
wire n_42794;
wire n_42795;
wire n_42796;
wire n_42797;
wire n_42798;
wire n_42799;
wire n_42800;
wire n_42801;
wire n_42802;
wire n_42803;
wire n_42804;
wire n_42805;
wire n_42806;
wire n_42807;
wire n_42808;
wire n_42809;
wire n_42810;
wire n_42811;
wire n_42812;
wire n_42813;
wire n_42814;
wire n_42815;
wire n_42816;
wire n_42817;
wire n_42818;
wire n_42819;
wire n_42820;
wire n_42821;
wire n_42822;
wire n_42823;
wire n_42824;
wire n_42825;
wire n_42826;
wire n_42827;
wire n_42828;
wire n_42829;
wire n_42830;
wire n_42831;
wire n_42832;
wire n_42833;
wire n_42834;
wire n_42835;
wire n_42836;
wire n_42837;
wire n_42838;
wire n_42839;
wire n_42840;
wire n_42841;
wire n_42842;
wire n_42843;
wire n_42844;
wire n_42845;
wire n_42846;
wire n_42847;
wire n_42848;
wire n_42849;
wire n_42850;
wire n_42851;
wire n_42852;
wire n_42853;
wire n_42854;
wire n_42855;
wire n_42856;
wire n_42857;
wire n_42858;
wire n_42859;
wire n_42860;
wire n_42861;
wire n_42862;
wire n_42863;
wire n_42864;
wire n_42865;
wire n_42866;
wire n_42867;
wire n_42868;
wire n_42869;
wire n_42870;
wire n_42871;
wire n_42872;
wire n_42873;
wire n_42874;
wire n_42875;
wire n_42876;
wire n_42877;
wire n_42878;
wire n_42879;
wire n_42880;
wire n_42881;
wire n_42882;
wire n_42883;
wire n_42884;
wire n_42885;
wire n_42886;
wire n_42887;
wire n_42888;
wire n_42889;
wire n_42890;
wire n_42891;
wire n_42892;
wire n_42893;
wire n_42894;
wire n_42895;
wire n_42896;
wire n_42897;
wire n_42898;
wire n_42899;
wire n_42900;
wire n_42901;
wire n_42902;
wire n_42903;
wire n_42904;
wire n_42905;
wire n_42906;
wire n_42907;
wire n_42908;
wire n_42909;
wire n_42910;
wire n_42911;
wire n_42912;
wire n_42913;
wire n_42914;
wire n_42915;
wire n_42916;
wire n_42917;
wire n_42918;
wire n_42919;
wire n_42920;
wire n_42921;
wire n_42922;
wire n_42923;
wire n_42924;
wire n_42925;
wire n_42926;
wire n_42927;
wire n_42928;
wire n_42929;
wire n_42930;
wire n_42931;
wire n_42932;
wire n_42933;
wire n_42934;
wire n_42935;
wire n_42936;
wire n_42937;
wire n_42938;
wire n_42939;
wire n_42940;
wire n_42941;
wire n_42942;
wire n_42943;
wire n_42944;
wire n_42945;
wire n_42946;
wire n_42947;
wire n_42948;
wire n_42949;
wire n_42950;
wire n_42951;
wire n_42952;
wire n_42953;
wire n_42954;
wire n_42955;
wire n_42956;
wire n_42957;
wire n_42958;
wire n_42959;
wire n_42960;
wire n_42961;
wire n_42962;
wire n_42963;
wire n_42964;
wire n_42965;
wire n_42966;
wire n_42967;
wire n_42968;
wire n_42969;
wire n_42970;
wire n_42971;
wire n_42972;
wire n_42973;
wire n_42974;
wire n_42975;
wire n_42976;
wire n_42977;
wire n_42978;
wire n_42979;
wire n_42980;
wire n_42981;
wire n_42982;
wire n_42983;
wire n_42984;
wire n_42985;
wire n_42986;
wire n_42987;
wire n_42988;
wire n_42989;
wire n_42990;
wire n_42991;
wire n_42992;
wire n_42993;
wire n_42994;
wire n_42995;
wire n_42996;
wire n_42997;
wire n_42998;
wire n_42999;
wire n_43000;
wire n_43001;
wire n_43002;
wire n_43003;
wire n_43004;
wire n_43005;
wire n_43006;
wire n_43007;
wire n_43008;
wire n_43009;
wire n_43010;
wire n_43011;
wire n_43012;
wire n_43013;
wire n_43014;
wire n_43015;
wire n_43016;
wire n_43017;
wire n_43018;
wire n_43019;
wire n_43020;
wire n_43021;
wire n_43022;
wire n_43023;
wire n_43024;
wire n_43025;
wire n_43026;
wire n_43027;
wire n_43028;
wire n_43029;
wire n_43030;
wire n_43031;
wire n_43032;
wire n_43033;
wire n_43034;
wire n_43035;
wire n_43036;
wire n_43037;
wire n_43038;
wire n_43039;
wire n_43040;
wire n_43041;
wire n_43042;
wire n_43043;
wire n_43044;
wire n_43045;
wire n_43046;
wire n_43047;
wire n_43048;
wire n_43049;
wire n_43050;
wire n_43051;
wire n_43052;
wire n_43053;
wire n_43054;
wire n_43055;
wire n_43056;
wire n_43057;
wire n_43058;
wire n_43059;
wire n_43060;
wire n_43061;
wire n_43062;
wire n_43063;
wire n_43064;
wire n_43065;
wire n_43066;
wire n_43067;
wire n_43068;
wire n_43069;
wire n_43070;
wire n_43071;
wire n_43072;
wire n_43073;
wire n_43074;
wire n_43075;
wire n_43076;
wire n_43077;
wire n_43078;
wire n_43079;
wire n_43080;
wire n_43081;
wire n_43082;
wire n_43083;
wire n_43084;
wire n_43085;
wire n_43086;
wire n_43087;
wire n_43088;
wire n_43089;
wire n_43090;
wire n_43091;
wire n_43092;
wire n_43093;
wire n_43094;
wire n_43095;
wire n_43096;
wire n_43097;
wire n_43098;
wire n_43099;
wire n_43100;
wire n_43101;
wire n_43102;
wire n_43103;
wire n_43104;
wire n_43105;
wire n_43106;
wire n_43107;
wire n_43108;
wire n_43109;
wire n_43110;
wire n_43111;
wire n_43112;
wire n_43113;
wire n_43114;
wire n_43115;
wire n_43116;
wire n_43117;
wire n_43118;
wire n_43119;
wire n_43120;
wire n_43121;
wire n_43122;
wire n_43123;
wire n_43124;
wire n_43125;
wire n_43126;
wire n_43127;
wire n_43128;
wire n_43129;
wire n_43130;
wire n_43131;
wire n_43132;
wire n_43133;
wire n_43134;
wire n_43135;
wire n_43136;
wire n_43137;
wire n_43138;
wire n_43139;
wire n_43140;
wire n_43141;
wire n_43142;
wire n_43143;
wire n_43144;
wire n_43145;
wire n_43146;
wire n_43147;
wire n_43148;
wire n_43149;
wire n_43150;
wire n_43151;
wire n_43152;
wire n_43153;
wire n_43154;
wire n_43155;
wire n_43156;
wire n_43157;
wire n_43158;
wire n_43159;
wire n_43160;
wire n_43161;
wire n_43162;
wire n_43163;
wire n_43164;
wire n_43165;
wire n_43166;
wire n_43167;
wire n_43168;
wire n_43169;
wire n_43170;
wire n_43171;
wire n_43172;
wire n_43173;
wire n_43174;
wire n_43175;
wire n_43176;
wire n_43177;
wire n_43178;
wire n_43179;
wire n_43180;
wire n_43181;
wire n_43182;
wire n_43183;
wire n_43184;
wire n_43185;
wire n_43186;
wire n_43187;
wire n_43188;
wire n_43189;
wire n_43190;
wire n_43191;
wire n_43192;
wire n_43193;
wire n_43194;
wire n_43195;
wire n_43196;
wire n_43197;
wire n_43198;
wire n_43199;
wire n_43200;
wire n_43201;
wire n_43202;
wire n_43203;
wire n_43204;
wire n_43205;
wire n_43206;
wire n_43207;
wire n_43208;
wire n_43209;
wire n_43210;
wire n_43211;
wire n_43212;
wire n_43213;
wire n_43214;
wire n_43215;
wire n_43216;
wire n_43217;
wire n_43218;
wire n_43219;
wire n_43220;
wire n_43221;
wire n_43222;
wire n_43223;
wire n_43224;
wire n_43225;
wire n_43226;
wire n_43227;
wire n_43228;
wire n_43229;
wire n_43230;
wire n_43231;
wire n_43232;
wire n_43233;
wire n_43234;
wire n_43235;
wire n_43236;
wire n_43237;
wire n_43238;
wire n_43239;
wire n_43240;
wire n_43241;
wire n_43242;
wire n_43243;
wire n_43244;
wire n_43245;
wire n_43246;
wire n_43247;
wire n_43248;
wire n_43249;
wire n_43250;
wire n_43251;
wire n_43252;
wire n_43253;
wire n_43254;
wire n_43255;
wire n_43256;
wire n_43257;
wire n_43258;
wire n_43259;
wire n_43260;
wire n_43261;
wire n_43262;
wire n_43263;
wire n_43264;
wire n_43265;
wire n_43266;
wire n_43267;
wire n_43268;
wire n_43269;
wire n_43270;
wire n_43271;
wire n_43272;
wire n_43273;
wire n_43274;
wire n_43275;
wire n_43276;
wire n_43277;
wire n_43278;
wire n_43279;
wire n_43280;
wire n_43281;
wire n_43282;
wire n_43283;
wire n_43284;
wire n_43285;
wire n_43286;
wire n_43287;
wire n_43288;
wire n_43289;
wire n_43290;
wire n_43291;
wire n_43292;
wire n_43293;
wire n_43294;
wire n_43295;
wire n_43296;
wire n_43297;
wire n_43298;
wire n_43299;
wire n_43300;
wire n_43301;
wire n_43302;
wire n_43303;
wire n_43304;
wire n_43305;
wire n_43306;
wire n_43307;
wire n_43308;
wire n_43309;
wire n_43310;
wire n_43311;
wire n_43312;
wire n_43313;
wire n_43314;
wire n_43315;
wire n_43316;
wire n_43317;
wire n_43318;
wire n_43319;
wire n_43320;
wire n_43321;
wire n_43322;
wire n_43323;
wire n_43324;
wire n_43325;
wire n_43326;
wire n_43327;
wire n_43328;
wire n_43329;
wire n_43330;
wire n_43331;
wire n_43332;
wire n_43333;
wire n_43334;
wire n_43335;
wire n_43336;
wire n_43337;
wire n_43338;
wire n_43339;
wire n_43340;
wire n_43341;
wire n_43342;
wire n_43343;
wire n_43344;
wire n_43345;
wire n_43346;
wire n_43347;
wire n_43348;
wire n_43349;
wire n_43350;
wire n_43351;
wire n_43352;
wire n_43353;
wire n_43354;
wire n_43355;
wire n_43356;
wire n_43357;
wire n_43358;
wire n_43359;
wire n_43360;
wire n_43361;
wire n_43362;
wire n_43363;
wire n_43364;
wire n_43365;
wire n_43366;
wire n_43367;
wire n_43368;
wire n_43369;
wire n_43370;
wire n_43371;
wire n_43372;
wire n_43373;
wire n_43374;
wire n_43375;
wire n_43376;
wire n_43377;
wire n_43378;
wire n_43379;
wire n_43380;
wire n_43381;
wire n_43382;
wire n_43383;
wire n_43384;
wire n_43385;
wire n_43386;
wire n_43387;
wire n_43388;
wire n_43389;
wire n_43390;
wire n_43391;
wire n_43392;
wire n_43393;
wire n_43394;
wire n_43395;
wire n_43396;
wire n_43397;
wire n_43398;
wire n_43399;
wire n_43400;
wire n_43401;
wire n_43402;
wire n_43403;
wire n_43404;
wire n_43405;
wire n_43406;
wire n_43407;
wire n_43408;
wire n_43409;
wire n_43410;
wire n_43411;
wire n_43412;
wire n_43413;
wire n_43414;
wire n_43415;
wire n_43416;
wire n_43417;
wire n_43418;
wire n_43419;
wire n_43420;
wire n_43421;
wire n_43422;
wire n_43423;
wire n_43424;
wire n_43425;
wire n_43426;
wire n_43427;
wire n_43428;
wire n_43429;
wire n_43430;
wire n_43431;
wire n_43432;
wire n_43433;
wire n_43434;
wire n_43435;
wire n_43436;
wire n_43437;
wire n_43438;
wire n_43439;
wire n_43440;
wire n_43441;
wire n_43442;
wire n_43443;
wire n_43444;
wire n_43445;
wire n_43446;
wire n_43447;
wire n_43448;
wire n_43449;
wire n_43450;
wire n_43451;
wire n_43452;
wire n_43453;
wire n_43454;
wire n_43455;
wire n_43456;
wire n_43457;
wire n_43458;
wire n_43459;
wire n_43460;
wire n_43461;
wire n_43462;
wire n_43463;
wire n_43464;
wire n_43465;
wire n_43466;
wire n_43467;
wire n_43468;
wire n_43469;
wire n_43470;
wire n_43471;
wire n_43472;
wire n_43473;
wire n_43474;
wire n_43475;
wire n_43476;
wire n_43477;
wire n_43478;
wire n_43479;
wire n_43480;
wire n_43481;
wire n_43482;
wire n_43483;
wire n_43484;
wire n_43485;
wire n_43486;
wire n_43487;
wire n_43488;
wire n_43489;
wire n_43490;
wire n_43491;
wire n_43492;
wire n_43493;
wire n_43494;
wire n_43495;
wire n_43496;
wire n_43497;
wire n_43498;
wire n_43499;
wire n_43500;
wire n_43501;
wire n_43502;
wire n_43503;
wire n_43504;
wire n_43505;
wire n_43506;
wire n_43507;
wire n_43508;
wire n_43509;
wire n_43510;
wire n_43511;
wire n_43512;
wire n_43513;
wire n_43514;
wire n_43515;
wire n_43516;
wire n_43517;
wire n_43518;
wire n_43519;
wire n_43520;
wire n_43521;
wire n_43522;
wire n_43523;
wire n_43524;
wire n_43525;
wire n_43526;
wire n_43527;
wire n_43528;
wire n_43529;
wire n_43530;
wire n_43531;
wire n_43532;
wire n_43533;
wire n_43534;
wire n_43535;
wire n_43536;
wire n_43537;
wire n_43538;
wire n_43539;
wire n_43540;
wire n_43541;
wire n_43542;
wire n_43543;
wire n_43544;
wire n_43545;
wire n_43546;
wire n_43547;
wire n_43548;
wire n_43549;
wire n_43550;
wire n_43551;
wire n_43552;
wire n_43553;
wire n_43554;
wire n_43555;
wire n_43556;
wire n_43557;
wire n_43558;
wire n_43559;
wire n_43560;
wire n_43561;
wire n_43562;
wire n_43563;
wire n_43564;
wire n_43565;
wire n_43566;
wire n_43567;
wire n_43568;
wire n_43569;
wire n_43570;
wire n_43571;
wire n_43572;
wire n_43573;
wire n_43574;
wire n_43575;
wire n_43576;
wire n_43577;
wire n_43578;
wire n_43579;
wire n_43580;
wire n_43581;
wire n_43582;
wire n_43583;
wire n_43584;
wire n_43585;
wire n_43586;
wire n_43587;
wire n_43588;
wire n_43589;
wire n_43590;
wire n_43591;
wire n_43592;
wire n_43593;
wire n_43594;
wire n_43595;
wire n_43596;
wire n_43597;
wire n_43598;
wire n_43599;
wire n_43600;
wire n_43601;
wire n_43602;
wire n_43603;
wire n_43604;
wire n_43605;
wire n_43606;
wire n_43607;
wire n_43608;
wire n_43609;
wire n_43610;
wire n_43611;
wire n_43612;
wire n_43613;
wire n_43614;
wire n_43615;
wire n_43616;
wire n_43617;
wire n_43618;
wire n_43619;
wire n_43620;
wire n_43621;
wire n_43622;
wire n_43623;
wire n_43624;
wire n_43625;
wire n_43626;
wire n_43627;
wire n_43628;
wire n_43629;
wire n_43630;
wire n_43631;
wire n_43632;
wire n_43633;
wire n_43634;
wire n_43635;
wire n_43636;
wire n_43637;
wire n_43638;
wire n_43639;
wire n_43640;
wire n_43641;
wire n_43642;
wire n_43643;
wire n_43644;
wire n_43645;
wire n_43646;
wire n_43647;
wire n_43648;
wire n_43649;
wire n_43650;
wire n_43651;
wire n_43652;
wire n_43653;
wire n_43654;
wire n_43655;
wire n_43656;
wire n_43657;
wire n_43658;
wire n_43659;
wire n_43660;
wire n_43661;
wire n_43662;
wire n_43663;
wire n_43664;
wire n_43665;
wire n_43666;
wire n_43667;
wire n_43668;
wire n_43669;
wire n_43670;
wire n_43671;
wire n_43672;
wire n_43673;
wire n_43674;
wire n_43675;
wire n_43676;
wire n_43677;
wire n_43678;
wire n_43679;
wire n_43680;
wire n_43681;
wire n_43682;
wire n_43683;
wire n_43684;
wire n_43685;
wire n_43686;
wire n_43687;
wire n_43688;
wire n_43689;
wire n_43690;
wire n_43691;
wire n_43692;
wire n_43693;
wire n_43694;
wire n_43695;
wire n_43696;
wire n_43697;
wire n_43698;
wire n_43699;
wire n_43700;
wire n_43701;
wire n_43702;
wire n_43703;
wire n_43704;
wire n_43705;
wire n_43706;
wire n_43707;
wire n_43708;
wire n_43709;
wire n_43710;
wire n_43711;
wire n_43712;
wire n_43713;
wire n_43714;
wire n_43715;
wire n_43716;
wire n_43717;
wire n_43718;
wire n_43719;
wire n_43720;
wire n_43721;
wire n_43722;
wire n_43723;
wire n_43724;
wire n_43725;
wire n_43726;
wire n_43727;
wire n_43728;
wire n_43729;
wire n_43730;
wire n_43731;
wire n_43732;
wire n_43733;
wire n_43734;
wire n_43735;
wire n_43736;
wire n_43737;
wire n_43738;
wire n_43739;
wire n_43740;
wire n_43741;
wire n_43742;
wire n_43743;
wire n_43744;
wire n_43745;
wire n_43746;
wire n_43747;
wire n_43748;
wire n_43749;
wire n_43750;
wire n_43751;
wire n_43752;
wire n_43753;
wire n_43754;
wire n_43755;
wire n_43756;
wire n_43757;
wire n_43758;
wire n_43759;
wire n_43760;
wire n_43761;
wire n_43762;
wire n_43763;
wire n_43764;
wire n_43765;
wire n_43766;
wire n_43767;
wire n_43768;
wire n_43769;
wire n_43770;
wire n_43771;
wire n_43772;
wire n_43773;
wire n_43774;
wire n_43775;
wire n_43776;
wire n_43777;
wire n_43778;
wire n_43779;
wire n_43780;
wire n_43781;
wire n_43782;
wire n_43783;
wire n_43784;
wire n_43785;
wire n_43786;
wire n_43787;
wire n_43788;
wire n_43789;
wire n_43790;
wire n_43791;
wire n_43792;
wire n_43793;
wire n_43794;
wire n_43795;
wire n_43796;
wire n_43797;
wire n_43798;
wire n_43799;
wire n_43800;
wire n_43801;
wire n_43802;
wire n_43803;
wire n_43804;
wire n_43805;
wire n_43806;
wire n_43807;
wire n_43808;
wire n_43809;
wire n_43810;
wire n_43811;
wire n_43812;
wire n_43813;
wire n_43814;
wire n_43815;
wire n_43816;
wire n_43817;
wire n_43818;
wire n_43819;
wire n_43820;
wire n_43821;
wire n_43822;
wire n_43823;
wire n_43824;
wire n_43825;
wire n_43826;
wire n_43827;
wire n_43828;
wire n_43829;
wire n_43830;
wire n_43831;
wire n_43832;
wire n_43833;
wire n_43834;
wire n_43835;
wire n_43836;
wire n_43837;
wire n_43838;
wire n_43839;
wire n_43840;
wire n_43841;
wire n_43842;
wire n_43843;
wire n_43844;
wire n_43845;
wire n_43846;
wire n_43847;
wire n_43848;
wire n_43849;
wire n_43850;
wire n_43851;
wire n_43852;
wire n_43853;
wire n_43854;
wire n_43855;
wire n_43856;
wire n_43857;
wire n_43858;
wire n_43859;
wire n_43860;
wire n_43861;
wire n_43862;
wire n_43863;
wire n_43864;
wire n_43865;
wire n_43866;
wire n_43867;
wire n_43868;
wire n_43869;
wire n_43870;
wire n_43871;
wire n_43872;
wire n_43873;
wire n_43874;
wire n_43875;
wire n_43876;
wire n_43877;
wire n_43878;
wire n_43879;
wire n_43880;
wire n_43881;
wire n_43882;
wire n_43883;
wire n_43884;
wire n_43885;
wire n_43886;
wire n_43887;
wire n_43888;
wire n_43889;
wire n_43890;
wire n_43891;
wire n_43892;
wire n_43893;
wire n_43894;
wire n_43895;
wire n_43896;
wire n_43897;
wire n_43898;
wire n_43899;
wire n_43900;
wire n_43901;
wire n_43902;
wire n_43903;
wire n_43904;
wire n_43905;
wire n_43906;
wire n_43907;
wire n_43908;
wire n_43909;
wire n_43910;
wire n_43911;
wire n_43912;
wire n_43913;
wire n_43914;
wire n_43915;
wire n_43916;
wire n_43917;
wire n_43918;
wire n_43919;
wire n_43920;
wire n_43921;
wire n_43922;
wire n_43923;
wire n_43924;
wire n_43925;
wire n_43926;
wire n_43927;
wire n_43928;
wire n_43929;
wire n_43930;
wire n_43931;
wire n_43932;
wire n_43933;
wire n_43934;
wire n_43935;
wire n_43936;
wire n_43937;
wire n_43938;
wire n_43939;
wire n_43940;
wire n_43941;
wire n_43942;
wire n_43943;
wire n_43944;
wire n_43945;
wire n_43946;
wire n_43947;
wire n_43948;
wire n_43949;
wire n_43950;
wire n_43951;
wire n_43952;
wire n_43953;
wire n_43954;
wire n_43955;
wire n_43956;
wire n_43957;
wire n_43958;
wire n_43959;
wire n_43960;
wire n_43961;
wire n_43962;
wire n_43963;
wire n_43964;
wire n_43965;
wire n_43966;
wire n_43967;
wire n_43968;
wire n_43969;
wire n_43970;
wire n_43971;
wire n_43972;
wire n_43973;
wire n_43974;
wire n_43975;
wire n_43976;
wire n_43977;
wire n_43978;
wire n_43979;
wire n_43980;
wire n_43981;
wire n_43982;
wire n_43983;
wire n_43984;
wire n_43985;
wire n_43986;
wire n_43987;
wire n_43988;
wire n_43989;
wire n_43990;
wire n_43991;
wire n_43992;
wire n_43993;
wire n_43994;
wire n_43995;
wire n_43996;
wire n_43997;
wire n_43998;
wire n_43999;
wire n_44000;
wire n_44001;
wire n_44002;
wire n_44003;
wire n_44004;
wire n_44005;
wire n_44006;
wire n_44007;
wire n_44008;
wire n_44009;
wire n_44010;
wire n_44011;
wire n_44012;
wire n_44013;
wire n_44014;
wire n_44015;
wire n_44016;
wire n_44017;
wire n_44018;
wire n_44019;
wire n_44020;
wire n_44021;
wire n_44022;
wire n_44023;
wire n_44024;
wire n_44025;
wire n_44026;
wire n_44027;
wire n_44028;
wire n_44029;
wire n_44030;
wire n_44031;
wire n_44032;
wire n_44033;
wire n_44034;
wire n_44035;
wire n_44036;
wire n_44037;
wire n_44038;
wire n_44039;
wire n_44040;
wire n_44041;
wire n_44042;
wire n_44043;
wire n_44044;
wire n_44045;
wire n_44046;
wire n_44047;
wire n_44048;
wire n_44049;
wire n_44050;
wire n_44051;
wire n_44052;
wire n_44053;
wire n_44054;
wire n_44055;
wire n_44056;
wire n_44057;
wire n_44058;
wire n_44059;
wire n_44060;
wire n_44061;
wire n_44062;
wire n_44063;
wire n_44064;
wire n_44065;
wire n_44066;
wire n_44067;
wire n_44068;
wire n_44069;
wire n_44070;
wire n_44071;
wire n_44072;
wire n_44073;
wire n_44074;
wire n_44075;
wire n_44076;
wire n_44077;
wire n_44078;
wire n_44079;
wire n_44080;
wire n_44081;
wire n_44082;
wire n_44083;
wire n_44084;
wire n_44085;
wire n_44086;
wire n_44087;
wire n_44088;
wire n_44089;
wire n_44090;
wire n_44091;
wire n_44092;
wire n_44093;
wire n_44094;
wire n_44095;
wire n_44096;
wire n_44097;
wire n_44098;
wire n_44099;
wire n_44100;
wire n_44101;
wire n_44102;
wire n_44103;
wire n_44104;
wire n_44105;
wire n_44106;
wire n_44107;
wire n_44108;
wire n_44109;
wire n_44110;
wire n_44111;
wire n_44112;
wire n_44113;
wire n_44114;
wire n_44115;
wire n_44116;
wire n_44117;
wire n_44118;
wire n_44119;
wire n_44120;
wire n_44121;
wire n_44122;
wire n_44123;
wire n_44124;
wire n_44125;
wire n_44126;
wire n_44127;
wire n_44128;
wire n_44129;
wire n_44130;
wire n_44131;
wire n_44132;
wire n_44133;
wire n_44134;
wire n_44135;
wire n_44136;
wire n_44137;
wire n_44138;
wire n_44139;
wire n_44140;
wire n_44141;
wire n_44142;
wire n_44143;
wire n_44144;
wire n_44145;
wire n_44146;
wire n_44147;
wire n_44148;
wire n_44149;
wire n_44150;
wire n_44151;
wire n_44152;
wire n_44153;
wire n_44154;
wire n_44155;
wire n_44156;
wire n_44157;
wire n_44158;
wire n_44159;
wire n_44160;
wire n_44161;
wire n_44162;
wire n_44163;
wire n_44164;
wire n_44165;
wire n_44166;
wire n_44167;
wire n_44168;
wire n_44169;
wire n_44170;
wire n_44171;
wire n_44172;
wire n_44173;
wire n_44174;
wire n_44175;
wire n_44176;
wire n_44177;
wire n_44178;
wire n_44179;
wire n_44180;
wire n_44181;
wire n_44182;
wire n_44183;
wire n_44184;
wire n_44185;
wire n_44186;
wire n_44187;
wire n_44188;
wire n_44189;
wire n_44190;
wire n_44191;
wire n_44192;
wire n_44193;
wire n_44194;
wire n_44195;
wire n_44196;
wire n_44197;
wire n_44198;
wire n_44199;
wire n_44200;
wire n_44201;
wire n_44202;
wire n_44203;
wire n_44204;
wire n_44205;
wire n_44206;
wire n_44207;
wire n_44208;
wire n_44209;
wire n_44210;
wire n_44211;
wire n_44212;
wire n_44213;
wire n_44214;
wire n_44215;
wire n_44216;
wire n_44217;
wire n_44218;
wire n_44219;
wire n_44220;
wire n_44221;
wire n_44222;
wire n_44223;
wire n_44224;
wire n_44225;
wire n_44226;
wire n_44227;
wire n_44228;
wire n_44229;
wire n_44230;
wire n_44231;
wire n_44232;
wire n_44233;
wire n_44234;
wire n_44235;
wire n_44236;
wire n_44237;
wire n_44238;
wire n_44239;
wire n_44240;
wire n_44241;
wire n_44242;
wire n_44243;
wire n_44244;
wire n_44245;
wire n_44246;
wire n_44247;
wire n_44248;
wire n_44249;
wire n_44250;
wire n_44251;
wire n_44252;
wire n_44253;
wire n_44254;
wire n_44255;
wire n_44256;
wire n_44257;
wire n_44258;
wire n_44259;
wire n_44260;
wire n_44261;
wire n_44262;
wire n_44263;
wire n_44264;
wire n_44265;
wire n_44266;
wire n_44267;
wire n_44268;
wire n_44269;
wire n_44270;
wire n_44271;
wire n_44272;
wire n_44273;
wire n_44274;
wire n_44275;
wire n_44276;
wire n_44277;
wire n_44278;
wire n_44279;
wire n_44280;
wire n_44281;
wire n_44282;
wire n_44283;
wire n_44284;
wire n_44285;
wire n_44286;
wire n_44287;
wire n_44288;
wire n_44289;
wire n_44290;
wire n_44291;
wire n_44292;
wire n_44293;
wire n_44294;
wire n_44295;
wire n_44296;
wire n_44297;
wire n_44298;
wire n_44299;
wire n_44300;
wire n_44301;
wire n_44302;
wire n_44303;
wire n_44304;
wire n_44305;
wire n_44306;
wire n_44307;
wire n_44308;
wire n_44309;
wire n_44310;
wire n_44311;
wire n_44312;
wire n_44313;
wire n_44314;
wire n_44315;
wire n_44316;
wire n_44317;
wire n_44318;
wire n_44319;
wire n_44320;
wire n_44321;
wire n_44322;
wire n_44323;
wire n_44324;
wire n_44325;
wire n_44326;
wire n_44327;
wire n_44328;
wire n_44329;
wire n_44330;
wire n_44331;
wire n_44332;
wire n_44333;
wire n_44334;
wire n_44335;
wire n_44336;
wire n_44337;
wire n_44338;
wire n_44339;
wire n_44340;
wire n_44341;
wire n_44342;
wire n_44343;
wire n_44344;
wire n_44345;
wire n_44346;
wire n_44347;
wire n_44348;
wire n_44349;
wire n_44350;
wire n_44351;
wire n_44352;
wire n_44353;
wire n_44354;
wire n_44355;
wire n_44356;
wire n_44357;
wire n_44358;
wire n_44359;
wire n_44360;
wire n_44361;
wire n_44362;
wire n_44363;
wire n_44364;
wire n_44365;
wire n_44366;
wire n_44367;
wire n_44368;
wire n_44369;
wire n_44370;
wire n_44371;
wire n_44372;
wire n_44373;
wire n_44374;
wire n_44375;
wire n_44376;
wire n_44377;
wire n_44378;
wire n_44379;
wire n_44380;
wire n_44381;
wire n_44382;
wire n_44383;
wire n_44384;
wire n_44385;
wire n_44386;
wire n_44387;
wire n_44388;
wire n_44389;
wire n_44390;
wire n_44391;
wire n_44392;
wire n_44393;
wire n_44394;
wire n_44395;
wire n_44396;
wire n_44397;
wire n_44398;
wire n_44399;
wire n_44400;
wire n_44401;
wire n_44402;
wire n_44403;
wire n_44404;
wire n_44405;
wire n_44406;
wire n_44407;
wire n_44408;
wire n_44409;
wire n_44410;
wire n_44411;
wire n_44412;
wire n_44413;
wire n_44414;
wire n_44415;
wire n_44416;
wire n_44417;
wire n_44418;
wire n_44419;
wire n_44420;
wire n_44421;
wire n_44422;
wire n_44423;
wire n_44424;
wire n_44425;
wire n_44426;
wire n_44427;
wire n_44428;
wire n_44429;
wire n_44430;
wire n_44431;
wire n_44432;
wire n_44433;
wire n_44434;
wire n_44435;
wire n_44436;
wire n_44437;
wire n_44438;
wire n_44439;
wire n_44440;
wire n_44441;
wire n_44442;
wire n_44443;
wire n_44444;
wire n_44445;
wire n_44446;
wire n_44447;
wire n_44448;
wire n_44449;
wire n_44450;
wire n_44451;
wire n_44452;
wire n_44453;
wire n_44454;
wire n_44455;
wire n_44456;
wire n_44457;
wire n_44458;
wire n_44459;
wire n_44460;
wire n_44461;
wire n_44462;
wire n_44463;
wire n_44464;
wire n_44465;
wire n_44466;
wire n_44467;
wire n_44468;
wire n_44469;
wire n_44470;
wire n_44471;
wire n_44472;
wire n_44473;
wire n_44474;
wire n_44475;
wire n_44476;
wire n_44477;
wire n_44478;
wire n_44479;
wire n_44480;
wire n_44481;
wire n_44482;
wire n_44483;
wire n_44484;
wire n_44485;
wire n_44486;
wire n_44487;
wire n_44488;
wire n_44489;
wire n_44490;
wire n_44491;
wire n_44492;
wire n_44493;
wire n_44494;
wire n_44495;
wire n_44496;
wire n_44497;
wire n_44498;
wire n_44499;
wire n_44500;
wire n_44501;
wire n_44502;
wire n_44503;
wire n_44504;
wire n_44505;
wire n_44506;
wire n_44507;
wire n_44508;
wire n_44509;
wire n_44510;
wire n_44511;
wire n_44512;
wire n_44513;
wire n_44514;
wire n_44515;
wire n_44516;
wire n_44517;
wire n_44518;
wire n_44519;
wire n_44520;
wire n_44521;
wire n_44522;
wire n_44523;
wire n_44524;
wire n_44525;
wire n_44526;
wire n_44527;
wire n_44528;
wire n_44529;
wire n_44530;
wire n_44531;
wire n_44532;
wire n_44533;
wire n_44534;
wire n_44535;
wire n_44536;
wire n_44537;
wire n_44538;
wire n_44539;
wire n_44540;
wire n_44541;
wire n_44542;
wire n_44543;
wire n_44544;
wire n_44545;
wire n_44546;
wire n_44547;
wire n_44548;
wire n_44549;
wire n_44550;
wire n_44551;
wire n_44552;
wire n_44553;
wire n_44554;
wire n_44555;
wire n_44556;
wire n_44557;
wire n_44558;
wire n_44559;
wire n_44560;
wire n_44561;
wire n_44562;
wire n_44563;
wire n_44564;
wire n_44565;
wire n_44566;
wire n_44567;
wire n_44568;
wire n_44569;
wire n_44570;
wire n_44571;
wire n_44572;
wire n_44573;
wire n_44574;
wire n_44575;
wire n_44576;
wire n_44577;
wire n_44578;
wire n_44579;
wire n_44580;
wire n_44581;
wire n_44582;
wire n_44583;
wire n_44584;
wire n_44585;
wire n_44586;
wire n_44587;
wire n_44588;
wire n_44589;
wire n_44590;
wire n_44591;
wire n_44592;
wire n_44593;
wire n_44594;
wire n_44595;
wire n_44596;
wire n_44597;
wire n_44598;
wire n_44599;
wire n_44600;
wire n_44601;
wire n_44602;
wire n_44603;
wire n_44604;
wire n_44605;
wire n_44606;
wire n_44607;
wire n_44608;
wire n_44609;
wire n_44610;
wire n_44611;
wire n_44612;
wire n_44613;
wire n_44614;
wire n_44615;
wire n_44616;
wire n_44617;
wire n_44618;
wire n_44619;
wire n_44620;
wire n_44621;
wire n_44622;
wire n_44623;
wire n_44624;
wire n_44625;
wire n_44626;
wire n_44627;
wire n_44628;
wire n_44629;
wire n_44630;
wire n_44631;
wire n_44632;
wire n_44633;
wire n_44634;
wire n_44635;
wire n_44636;
wire n_44637;
wire n_44638;
wire n_44639;
wire n_44640;
wire n_44641;
wire n_44642;
wire n_44643;
wire n_44644;
wire n_44645;
wire n_44646;
wire n_44647;
wire n_44648;
wire n_44649;
wire n_44650;
wire n_44651;
wire n_44652;
wire n_44653;
wire n_44654;
wire n_44655;
wire n_44656;
wire n_44657;
wire n_44658;
wire n_44659;
wire n_44660;
wire n_44661;
wire n_44662;
wire n_44663;
wire n_44664;
wire n_44665;
wire n_44666;
wire n_44667;
wire n_44668;
wire n_44669;
wire n_44670;
wire n_44671;
wire n_44672;
wire n_44673;
wire n_44674;
wire n_44675;
wire n_44676;
wire n_44677;
wire n_44678;
wire n_44679;
wire n_44680;
wire n_44681;
wire n_44682;
wire n_44683;
wire n_44684;
wire n_44685;
wire n_44686;
wire n_44687;
wire n_44688;
wire n_44689;
wire n_44690;
wire n_44691;
wire n_44692;
wire n_44693;
wire n_44694;
wire n_44695;
wire n_44696;
wire n_44697;
wire n_44698;
wire n_44699;
wire n_44700;
wire n_44701;
wire n_44702;
wire n_44703;
wire n_44704;
wire n_44705;
wire n_44706;
wire n_44707;
wire n_44708;
wire n_44709;
wire n_44710;
wire n_44711;
wire n_44712;
wire n_44713;
wire n_44714;
wire n_44715;
wire n_44716;
wire n_44717;
wire n_44718;
wire n_44719;
wire n_44720;
wire n_44721;
wire n_44722;
wire n_44723;
wire n_44724;
wire n_44725;
wire n_44726;
wire n_44727;
wire n_44728;
wire n_44729;
wire n_44730;
wire n_44731;
wire n_44732;
wire n_44733;
wire n_44734;
wire n_44735;
wire n_44736;
wire n_44737;
wire n_44738;
wire n_44739;
wire n_44740;
wire n_44741;
wire n_44742;
wire n_44743;
wire n_44744;
wire n_44745;
wire n_44746;
wire n_44747;
wire n_44748;
wire n_44749;
wire n_44750;
wire n_44751;
wire n_44752;
wire n_44753;
wire n_44754;
wire n_44755;
wire n_44756;
wire n_44757;
wire n_44758;
wire n_44759;
wire n_44760;
wire n_44761;
wire n_44762;
wire n_44763;
wire n_44764;
wire n_44765;
wire n_44766;
wire n_44767;
wire n_44768;
wire n_44769;
wire n_44770;
wire n_44771;
wire n_44772;
wire n_44773;
wire n_44774;
wire n_44775;
wire n_44776;
wire n_44777;
wire n_44778;
wire n_44779;
wire n_44780;
wire n_44781;
wire n_44782;
wire n_44783;
wire n_44784;
wire n_44785;
wire n_44786;
wire n_44787;
wire n_44788;
wire n_44789;
wire n_44790;
wire n_44791;
wire n_44792;
wire n_44793;
wire n_44794;
wire n_44795;
wire n_44796;
wire n_44797;
wire n_44798;
wire n_44799;
wire n_44800;
wire n_44801;
wire n_44802;
wire n_44803;
wire n_44804;
wire n_44805;
wire n_44806;
wire n_44807;
wire n_44808;
wire n_44809;
wire n_44810;
wire n_44811;
wire n_44812;
wire n_44813;
wire n_44814;
wire n_44815;
wire n_44816;
wire n_44817;
wire n_44818;
wire n_44819;
wire n_44820;
wire n_44821;
wire n_44822;
wire n_44823;
wire n_44824;
wire n_44825;
wire n_44826;
wire n_44827;
wire n_44828;
wire n_44829;
wire n_44830;
wire n_44831;
wire n_44832;
wire n_44833;
wire n_44834;
wire n_44835;
wire n_44836;
wire n_44837;
wire n_44838;
wire n_44839;
wire n_44840;
wire n_44841;
wire n_44842;
wire n_44843;
wire n_44844;
wire n_44845;
wire n_44846;
wire n_44847;
wire n_44848;
wire n_44849;
wire n_44850;
wire n_44851;
wire n_44852;
wire n_44853;
wire n_44854;
wire n_44855;
wire n_44856;
wire n_44857;
wire n_44858;
wire n_44859;
wire n_44860;
wire n_44861;
wire n_44862;
wire n_44863;
wire n_44864;
wire n_44865;
wire n_44866;
wire n_44867;
wire n_44868;
wire n_44869;
wire n_44870;
wire n_44871;
wire n_44872;
wire n_44873;
wire n_44874;
wire n_44875;
wire n_44876;
wire n_44877;
wire n_44878;
wire n_44879;
wire n_44880;
wire n_44881;
wire n_44882;
wire n_44883;
wire n_44884;
wire n_44885;
wire n_44886;
wire n_44887;
wire n_44888;
wire n_44889;
wire n_44890;
wire n_44891;
wire n_44892;
wire n_44893;
wire n_44894;
wire n_44895;
wire n_44896;
wire n_44897;
wire n_44898;
wire n_44899;
wire n_44900;
wire n_44901;
wire n_44902;
wire n_44903;
wire n_44904;
wire n_44905;
wire n_44906;
wire n_44907;
wire n_44908;
wire n_44909;
wire n_44910;
wire n_44911;
wire n_44912;
wire n_44913;
wire n_44914;
wire n_44915;
wire n_44916;
wire n_44917;
wire n_44918;
wire n_44919;
wire n_44920;
wire n_44921;
wire n_44922;
wire n_44923;
wire n_44924;
wire n_44925;
wire n_44926;
wire n_44927;
wire n_44928;
wire n_44929;
wire n_44930;
wire n_44931;
wire n_44932;
wire n_44933;
wire n_44934;
wire n_44935;
wire n_44936;
wire n_44937;
wire n_44938;
wire n_44939;
wire n_44940;
wire n_44941;
wire n_44942;
wire n_44943;
wire n_44944;
wire n_44945;
wire n_44946;
wire n_44947;
wire n_44948;
wire n_44949;
wire n_44950;
wire n_44951;
wire n_44952;
wire n_44953;
wire n_44954;
wire n_44955;
wire n_44956;
wire n_44957;
wire n_44958;
wire n_44959;
wire n_44960;
wire n_44961;
wire n_44962;
wire n_44963;
wire n_44964;
wire n_44965;
wire n_44966;
wire n_44967;
wire n_44968;
wire n_44969;
wire n_44970;
wire n_44971;
wire n_44972;
wire n_44973;
wire n_44974;
wire n_44975;
wire n_44976;
wire n_44977;
wire n_44978;
wire n_44979;
wire n_44980;
wire n_44981;
wire n_44982;
wire n_44983;
wire n_44984;
wire n_44985;
wire n_44986;
wire n_44987;
wire n_44988;
wire n_44989;
wire n_44990;
wire n_44991;
wire n_44992;
wire n_44993;
wire n_44994;
wire n_44995;
wire n_44996;
wire n_44997;
wire n_44998;
wire n_44999;
wire n_45000;
wire n_45001;
wire n_45002;
wire n_45003;
wire n_45004;
wire n_45005;
wire n_45006;
wire n_45007;
wire n_45008;
wire n_45009;
wire n_45010;
wire n_45011;
wire n_45012;
wire n_45013;
wire n_45014;
wire n_45015;
wire n_45016;
wire n_45017;
wire n_45018;
wire n_45019;
wire n_45020;
wire n_45021;
wire n_45022;
wire n_45023;
wire n_45024;
wire n_45025;
wire n_45026;
wire n_45027;
wire n_45028;
wire n_45029;
wire n_45030;
wire n_45031;
wire n_45032;
wire n_45033;
wire n_45034;
wire n_45035;
wire n_45036;
wire n_45037;
wire n_45038;
wire n_45039;
wire n_45040;
wire n_45041;
wire n_45042;
wire n_45043;
wire n_45044;
wire n_45045;
wire n_45046;
wire n_45047;
wire n_45048;
wire n_45049;
wire n_45050;
wire n_45051;
wire n_45052;
wire n_45053;
wire n_45054;
wire n_45055;
wire n_45056;
wire n_45057;
wire n_45058;
wire n_45059;
wire n_45060;
wire n_45061;
wire n_45062;
wire n_45063;
wire n_45064;
wire n_45065;
wire n_45066;
wire n_45067;
wire n_45068;
wire n_45069;
wire n_45070;
wire n_45071;
wire n_45072;
wire n_45073;
wire n_45074;
wire n_45075;
wire n_45076;
wire n_45077;
wire n_45078;
wire n_45079;
wire n_45080;
wire n_45081;
wire n_45082;
wire n_45083;
wire n_45084;
wire n_45085;
wire n_45086;
wire n_45087;
wire n_45088;
wire n_45089;
wire n_45090;
wire n_45091;
wire n_45092;
wire n_45093;
wire n_45094;
wire n_45095;
wire n_45096;
wire n_45097;
wire n_45098;
wire n_45099;
wire n_45100;
wire n_45101;
wire n_45102;
wire n_45103;
wire n_45104;
wire n_45105;
wire n_45106;
wire n_45107;
wire n_45108;
wire n_45109;
wire n_45110;
wire n_45111;
wire n_45112;
wire n_45113;
wire n_45114;
wire n_45115;
wire n_45116;
wire n_45117;
wire n_45118;
wire n_45119;
wire n_45120;
wire n_45121;
wire n_45122;
wire n_45123;
wire n_45124;
wire n_45125;
wire n_45126;
wire n_45127;
wire n_45128;
wire n_45129;
wire n_45130;
wire n_45131;
wire n_45132;
wire n_45133;
wire n_45134;
wire n_45135;
wire n_45136;
wire n_45137;
wire n_45138;
wire n_45139;
wire n_45140;
wire n_45141;
wire n_45142;
wire n_45143;
wire n_45144;
wire n_45145;
wire n_45146;
wire n_45147;
wire n_45148;
wire n_45149;
wire n_45150;
wire n_45151;
wire n_45152;
wire n_45153;
wire n_45154;
wire n_45155;
wire n_45156;
wire n_45157;
wire n_45158;
wire n_45159;
wire n_45160;
wire n_45161;
wire n_45162;
wire n_45163;
wire n_45164;
wire n_45165;
wire n_45166;
wire n_45167;
wire n_45168;
wire n_45169;
wire n_45170;
wire n_45171;
wire n_45172;
wire n_45173;
wire n_45174;
wire n_45175;
wire n_45176;
wire n_45177;
wire n_45178;
wire n_45179;
wire n_45180;
wire n_45181;
wire n_45182;
wire n_45183;
wire n_45184;
wire n_45185;
wire n_45186;
wire n_45187;
wire n_45188;
wire n_45189;
wire n_45190;
wire n_45191;
wire n_45192;
wire n_45193;
wire n_45194;
wire n_45195;
wire n_45196;
wire n_45197;
wire n_45198;
wire n_45199;
wire n_45200;
wire n_45201;
wire n_45202;
wire n_45203;
wire n_45204;
wire n_45205;
wire n_45206;
wire n_45207;
wire n_45208;
wire n_45209;
wire n_45210;
wire n_45211;
wire n_45212;
wire n_45213;
wire n_45214;
wire n_45215;
wire n_45216;
wire n_45217;
wire n_45218;
wire n_45219;
wire n_45220;
wire n_45221;
wire n_45222;
wire n_45223;
wire n_45224;
wire n_45225;
wire n_45226;
wire n_45227;
wire n_45228;
wire n_45229;
wire n_45230;
wire n_45231;
wire n_45232;
wire n_45233;
wire n_45234;
wire n_45235;
wire n_45236;
wire n_45237;
wire n_45238;
wire n_45239;
wire n_45240;
wire n_45241;
wire n_45242;
wire n_45243;
wire n_45244;
wire n_45245;
wire n_45246;
wire n_45247;
wire n_45248;
wire n_45249;
wire n_45250;
wire n_45251;
wire n_45252;
wire n_45253;
wire n_45254;
wire n_45255;
wire n_45256;
wire n_45257;
wire n_45258;
wire n_45259;
wire n_45260;
wire n_45261;
wire n_45262;
wire n_45263;
wire n_45264;
wire n_45265;
wire n_45266;
wire n_45267;
wire n_45268;
wire n_45269;
wire n_45270;
wire n_45271;
wire n_45272;
wire n_45273;
wire n_45274;
wire n_45275;
wire n_45276;
wire n_45277;
wire n_45278;
wire n_45279;
wire n_45280;
wire n_45281;
wire n_45282;
wire n_45283;
wire n_45284;
wire n_45285;
wire n_45286;
wire n_45287;
wire n_45288;
wire n_45289;
wire n_45290;
wire n_45291;
wire n_45292;
wire n_45293;
wire n_45294;
wire n_45295;
wire n_45296;
wire n_45297;
wire n_45298;
wire n_45299;
wire n_45300;
wire n_45301;
wire n_45302;
wire n_45303;
wire n_45304;
wire n_45305;
wire n_45306;
wire n_45307;
wire n_45308;
wire n_45309;
wire n_45310;
wire n_45311;
wire n_45312;
wire n_45313;
wire n_45314;
wire n_45315;
wire n_45316;
wire n_45317;
wire n_45318;
wire n_45319;
wire n_45320;
wire n_45321;
wire n_45322;
wire n_45323;
wire n_45324;
wire n_45325;
wire n_45326;
wire n_45327;
wire n_45328;
wire n_45329;
wire n_45330;
wire n_45331;
wire n_45332;
wire n_45333;
wire n_45334;
wire n_45335;
wire n_45336;
wire n_45337;
wire n_45338;
wire n_45339;
wire n_45340;
wire n_45341;
wire n_45342;
wire n_45343;
wire n_45344;
wire n_45345;
wire n_45346;
wire n_45347;
wire n_45348;
wire n_45349;
wire n_45350;
wire n_45351;
wire n_45352;
wire n_45353;
wire n_45354;
wire n_45355;
wire n_45356;
wire n_45357;
wire n_45358;
wire n_45359;
wire n_45360;
wire n_45361;
wire n_45362;
wire n_45363;
wire n_45364;
wire n_45365;
wire n_45366;
wire n_45367;
wire n_45368;
wire n_45369;
wire n_45370;
wire n_45371;
wire n_45372;
wire n_45373;
wire n_45374;
wire n_45375;
wire n_45376;
wire n_45377;
wire n_45378;
wire n_45379;
wire n_45380;
wire n_45381;
wire n_45382;
wire n_45383;
wire n_45384;
wire n_45385;
wire n_45386;
wire n_45387;
wire n_45388;
wire n_45389;
wire n_45390;
wire n_45391;
wire n_45392;
wire n_45393;
wire n_45394;
wire n_45395;
wire n_45396;
wire n_45397;
wire n_45398;
wire n_45399;
wire n_45400;
wire n_45401;
wire n_45402;
wire n_45403;
wire n_45404;
wire n_45405;
wire n_45406;
wire n_45407;
wire n_45408;
wire n_45409;
wire n_45410;
wire n_45411;
wire n_45412;
wire n_45413;
wire n_45414;
wire n_45415;
wire n_45416;
wire n_45417;
wire n_45418;
wire n_45419;
wire n_45420;
wire n_45421;
wire n_45422;
wire n_45423;
wire n_45424;
wire n_45425;
wire n_45426;
wire n_45427;
wire n_45428;
wire n_45429;
wire n_45430;
wire n_45431;
wire n_45432;
wire n_45433;
wire n_45434;
wire n_45435;
wire n_45436;
wire n_45437;
wire n_45438;
wire n_45439;
wire n_45440;
wire n_45441;
wire n_45442;
wire n_45443;
wire n_45444;
wire n_45445;
wire n_45446;
wire n_45447;
wire n_45448;
wire n_45449;
wire n_45450;
wire n_45451;
wire n_45452;
wire n_45453;
wire n_45454;
wire n_45455;
wire n_45456;
wire n_45457;
wire n_45458;
wire n_45459;
wire n_45460;
wire n_45461;
wire n_45462;
wire n_45463;
wire n_45464;
wire n_45465;
wire n_45466;
wire n_45467;
wire n_45468;
wire n_45469;
wire n_45470;
wire n_45471;
wire n_45472;
wire n_45473;
wire n_45474;
wire n_45475;
wire n_45476;
wire n_45477;
wire n_45478;
wire n_45479;
wire n_45480;
wire n_45481;
wire n_45482;
wire n_45483;
wire n_45484;
wire n_45485;
wire n_45486;
wire n_45487;
wire n_45488;
wire n_45489;
wire n_45490;
wire n_45491;
wire n_45492;
wire n_45493;
wire n_45494;
wire n_45495;
wire n_45496;
wire n_45497;
wire n_45498;
wire n_45499;
wire n_45500;
wire n_45501;
wire n_45502;
wire n_45503;
wire n_45504;
wire n_45505;
wire n_45506;
wire n_45507;
wire n_45508;
wire n_45509;
wire n_45510;
wire n_45511;
wire n_45512;
wire n_45513;
wire n_45514;
wire n_45515;
wire n_45516;
wire n_45517;
wire n_45518;
wire n_45519;
wire n_45520;
wire n_45521;
wire n_45522;
wire n_45523;
wire n_45524;
wire n_45525;
wire n_45526;
wire n_45527;
wire n_45528;
wire n_45529;
wire n_45530;
wire n_45531;
wire n_45532;
wire n_45533;
wire n_45534;
wire n_45535;
wire n_45536;
wire n_45537;
wire n_45538;
wire n_45539;
wire n_45540;
wire n_45541;
wire n_45542;
wire n_45543;
wire n_45544;
wire n_45545;
wire n_45546;
wire n_45547;
wire n_45548;
wire n_45549;
wire n_45550;
wire n_45551;
wire n_45552;
wire n_45553;
wire n_45554;
wire n_45555;
wire n_45556;
wire n_45557;
wire n_45558;
wire n_45559;
wire n_45560;
wire n_45561;
wire n_45562;
wire n_45563;
wire n_45564;
wire n_45565;
wire n_45566;
wire n_45567;
wire n_45568;
wire n_45569;
wire n_45570;
wire n_45571;
wire n_45572;
wire n_45573;
wire n_45574;
wire n_45575;
wire n_45576;
wire n_45577;
wire n_45578;
wire n_45579;
wire n_45580;
wire n_45581;
wire n_45582;
wire n_45583;
wire n_45584;
wire n_45585;
wire n_45586;
wire n_45587;
wire n_45588;
wire n_45589;
wire n_45590;
wire n_45591;
wire n_45592;
wire n_45593;
wire n_45594;
wire n_45595;
wire n_45596;
wire n_45597;
wire n_45598;
wire n_45599;
wire n_45600;
wire n_45601;
wire n_45602;
wire n_45603;
wire n_45604;
wire n_45605;
wire n_45606;
wire n_45607;
wire n_45608;
wire n_45609;
wire n_45610;
wire n_45611;
wire n_45612;
wire n_45613;
wire n_45614;
wire n_45615;
wire n_45616;
wire n_45617;
wire n_45618;
wire n_45619;
wire n_45620;
wire n_45621;
wire n_45622;
wire n_45623;
wire n_45624;
wire n_45625;
wire n_45626;
wire n_45627;
wire n_45628;
wire n_45629;
wire n_45630;
wire n_45631;
wire n_45632;
wire n_45633;
wire n_45634;
wire n_45635;
wire n_45636;
wire n_45637;
wire n_45638;
wire n_45639;
wire n_45640;
wire n_45641;
wire n_45642;
wire n_45643;
wire n_45644;
wire n_45645;
wire n_45646;
wire n_45647;
wire n_45648;
wire n_45649;
wire n_45650;
wire n_45651;
wire n_45652;
wire n_45653;
wire n_45654;
wire n_45655;
wire n_45656;
wire n_45657;
wire n_45658;
wire n_45659;
wire n_45660;
wire n_45661;
wire n_45662;
wire n_45663;
wire n_45664;
wire n_45665;
wire n_45666;
wire n_45667;
wire n_45668;
wire n_45669;
wire n_45670;
wire n_45671;
wire n_45672;
wire n_45673;
wire n_45674;
wire n_45675;
wire n_45676;
wire n_45677;
wire n_45678;
wire n_45679;
wire n_45680;
wire n_45681;
wire n_45682;
wire n_45683;
wire n_45684;
wire n_45685;
wire n_45686;
wire n_45687;
wire n_45688;
wire n_45689;
wire n_45690;
wire n_45691;
wire n_45692;
wire n_45693;
wire n_45694;
wire n_45695;
wire n_45696;
wire n_45697;
wire n_45698;
wire n_45699;
wire n_45700;
wire n_45701;
wire n_45702;
wire n_45703;
wire n_45704;
wire n_45705;
wire n_45706;
wire n_45707;
wire n_45708;
wire n_45709;
wire n_45710;
wire n_45711;
wire n_45712;
wire n_45713;
wire n_45714;
wire n_45715;
wire n_45716;
wire n_45717;
wire n_45718;
wire n_45719;
wire n_45720;
wire n_45721;
wire n_45722;
wire n_45723;
wire n_45724;
wire n_45725;
wire n_45726;
wire n_45727;
wire n_45728;
wire n_45729;
wire n_45730;
wire n_45731;
wire n_45732;
wire n_45733;
wire n_45734;
wire n_45735;
wire n_45736;
wire n_45737;
wire n_45738;
wire n_45739;
wire n_45740;
wire n_45741;
wire n_45742;
wire n_45743;
wire n_45744;
wire n_45745;
wire n_45746;
wire n_45747;
wire n_45748;
wire n_45749;
wire n_45750;
wire n_45751;
wire n_45752;
wire n_45753;
wire n_45754;
wire n_45755;
wire n_45756;
wire n_45757;
wire n_45758;
wire n_45759;
wire n_45760;
wire n_45761;
wire n_45762;
wire n_45763;
wire n_45764;
wire n_45765;
wire n_45766;
wire n_45767;
wire n_45768;
wire n_45769;
wire n_45770;
wire n_45771;
wire n_45772;
wire n_45773;
wire n_45774;
wire n_45775;
wire n_45776;
wire n_45777;
wire n_45778;
wire n_45779;
wire n_45780;
wire n_45781;
wire n_45782;
wire n_45783;
wire n_45784;
wire n_45785;
wire n_45786;
wire n_45787;
wire n_45788;
wire n_45789;
wire n_45790;
wire n_45791;
wire n_45792;
wire n_45793;
wire n_45794;
wire n_45795;
wire n_45796;
wire n_45797;
wire n_45798;
wire n_45799;
wire n_45800;
wire n_45801;
wire n_45802;
wire n_45803;
wire n_45804;
wire n_45805;
wire n_45806;
wire n_45807;
wire n_45808;
wire n_45809;
wire n_45810;
wire n_45811;
wire n_45812;
wire n_45813;
wire n_45814;
wire n_45815;
wire n_45816;
wire n_45817;
wire n_45818;
wire n_45819;
wire n_45820;
wire n_45821;
wire n_45822;
wire n_45823;
wire n_45824;
wire n_45825;
wire n_45826;
wire n_45827;
wire n_45828;
wire n_45829;
wire n_45830;
wire n_45831;
wire n_45832;
wire n_45833;
wire n_45834;
wire n_45835;
wire n_45836;
wire n_45837;
wire n_45838;
wire n_45839;
wire n_45840;
wire n_45841;
wire n_45842;
wire n_45843;
wire n_45844;
wire n_45845;
wire n_45846;
wire n_45847;
wire n_45848;
wire n_45849;
wire n_45850;
wire n_45851;
wire n_45852;
wire n_45853;
wire n_45854;
wire n_45855;
wire n_45856;
wire n_45857;
wire n_45858;
wire n_45859;
wire n_45860;
wire n_45861;
wire n_45862;
wire n_45863;
wire n_45864;
wire n_45865;
wire n_45866;
wire n_45867;
wire n_45868;
wire n_45869;
wire n_45870;
wire n_45871;
wire n_45872;
wire n_45873;
wire n_45874;
wire n_45875;
wire n_45876;
wire n_45877;
wire n_45878;
wire n_45879;
wire n_45880;
wire n_45881;
wire n_45882;
wire n_45883;
wire n_45884;
wire n_45885;
wire n_45886;
wire n_45887;
wire n_45888;
wire n_45889;
wire n_45890;
wire n_45891;
wire n_45892;
wire n_45893;
wire n_45894;
wire n_45895;
wire n_45896;
wire n_45897;
wire n_45898;
wire n_45899;
wire n_45900;
wire n_45901;
wire n_45902;
wire n_45903;
wire n_45904;
wire n_45905;
wire n_45906;
wire n_45907;
wire n_45908;
wire n_45909;
wire n_45910;
wire n_45911;
wire n_45912;
wire n_45913;
wire n_45914;
wire n_45915;
wire n_45916;
wire n_45917;
wire n_45918;
wire n_45919;
wire n_45920;
wire n_45921;
wire n_45922;
wire n_45923;
wire n_45924;
wire n_45925;
wire n_45926;
wire n_45927;
wire n_45928;
wire n_45929;
wire n_45930;
wire n_45931;
wire n_45932;
wire n_45933;
wire n_45934;
wire n_45935;
wire n_45936;
wire n_45937;
wire n_45938;
wire n_45939;
wire n_45940;
wire n_45941;
wire n_45942;
wire n_45943;
wire n_45944;
wire n_45945;
wire n_45946;
wire n_45947;
wire n_45948;
wire n_45949;
wire n_45950;
wire n_45951;
wire n_45952;
wire n_45953;
wire n_45954;
wire n_45955;
wire n_45956;
wire n_45957;
wire n_45958;
wire n_45959;
wire n_45960;
wire n_45961;
wire n_45962;
wire n_45963;
wire n_45964;
wire n_45965;
wire n_45966;
wire n_45967;
wire n_45968;
wire n_45969;
wire n_45970;
wire n_45971;
wire n_45972;
wire n_45973;
wire n_45974;
wire n_45975;
wire n_45976;
wire n_45977;
wire n_45978;
wire n_45979;
wire n_45980;
wire n_45981;
wire n_45982;
wire n_45983;
wire n_45984;
wire n_45985;
wire n_45986;
wire n_45987;
wire n_45988;
wire n_45989;
wire n_45990;
wire n_45991;
wire n_45992;
wire n_45993;
wire n_45994;
wire n_45995;
wire n_45996;
wire n_45997;
wire n_45998;
wire n_45999;
wire n_46000;
wire n_46001;
wire n_46002;
wire n_46003;
wire n_46004;
wire n_46005;
wire n_46006;
wire n_46007;
wire n_46008;
wire n_46009;
wire n_46010;
wire n_46011;
wire n_46012;
wire n_46013;
wire n_46014;
wire n_46015;
wire n_46016;
wire n_46017;
wire n_46018;
wire n_46019;
wire n_46020;
wire n_46021;
wire n_46022;
wire n_46023;
wire n_46024;
wire n_46025;
wire n_46026;
wire n_46027;
wire n_46028;
wire n_46029;
wire n_46030;
wire n_46031;
wire n_46032;
wire n_46033;
wire n_46034;
wire n_46035;
wire n_46036;
wire n_46037;
wire n_46038;
wire n_46039;
wire n_46040;
wire n_46041;
wire n_46042;
wire n_46043;
wire n_46044;
wire n_46045;
wire n_46046;
wire n_46047;
wire n_46048;
wire n_46049;
wire n_46050;
wire n_46051;
wire n_46052;
wire n_46053;
wire n_46054;
wire n_46055;
wire n_46056;
wire n_46057;
wire n_46058;
wire n_46059;
wire n_46060;
wire n_46061;
wire n_46062;
wire n_46063;
wire n_46064;
wire n_46065;
wire n_46066;
wire n_46067;
wire n_46068;
wire n_46069;
wire n_46070;
wire n_46071;
wire n_46072;
wire n_46073;
wire n_46074;
wire n_46075;
wire n_46076;
wire n_46077;
wire n_46078;
wire n_46079;
wire n_46080;
wire n_46081;
wire n_46082;
wire n_46083;
wire n_46084;
wire n_46085;
wire n_46086;
wire n_46087;
wire n_46088;
wire n_46089;
wire n_46090;
wire n_46091;
wire n_46092;
wire n_46093;
wire n_46094;
wire n_46095;
wire n_46096;
wire n_46097;
wire n_46098;
wire n_46099;
wire n_46100;
wire n_46101;
wire n_46102;
wire n_46103;
wire n_46104;
wire n_46105;
wire n_46106;
wire n_46107;
wire n_46108;
wire n_46109;
wire n_46110;
wire n_46111;
wire n_46112;
wire n_46113;
wire n_46114;
wire n_46115;
wire n_46116;
wire n_46117;
wire n_46118;
wire n_46119;
wire n_46120;
wire n_46121;
wire n_46122;
wire n_46123;
wire n_46124;
wire n_46125;
wire n_46126;
wire n_46127;
wire n_46128;
wire n_46129;
wire n_46130;
wire n_46131;
wire n_46132;
wire n_46133;
wire n_46134;
wire n_46135;
wire n_46136;
wire n_46137;
wire n_46138;
wire n_46139;
wire n_46140;
wire n_46141;
wire n_46142;
wire n_46143;
wire n_46144;
wire n_46145;
wire n_46146;
wire n_46147;
wire n_46148;
wire n_46149;
wire n_46150;
wire n_46151;
wire n_46152;
wire n_46153;
wire n_46154;
wire n_46155;
wire n_46156;
wire n_46157;
wire n_46158;
wire n_46159;
wire n_46160;
wire n_46161;
wire n_46162;
wire n_46163;
wire n_46164;
wire n_46165;
wire n_46166;
wire n_46167;
wire n_46168;
wire n_46169;
wire n_46170;
wire n_46171;
wire n_46172;
wire n_46173;
wire n_46174;
wire n_46175;
wire n_46176;
wire n_46177;
wire n_46178;
wire n_46179;
wire n_46180;
wire n_46181;
wire n_46182;
wire n_46183;
wire n_46184;
wire n_46185;
wire n_46186;
wire n_46187;
wire n_46188;
wire n_46189;
wire n_46190;
wire n_46191;
wire n_46192;
wire n_46193;
wire n_46194;
wire n_46195;
wire n_46196;
wire n_46197;
wire n_46198;
wire n_46199;
wire n_46200;
wire n_46201;
wire n_46202;
wire n_46203;
wire n_46204;
wire n_46205;
wire n_46206;
wire n_46207;
wire n_46208;
wire n_46209;
wire n_46210;
wire n_46211;
wire n_46212;
wire n_46213;
wire n_46214;
wire n_46215;
wire n_46216;
wire n_46217;
wire n_46218;
wire n_46219;
wire n_46220;
wire n_46221;
wire n_46222;
wire n_46223;
wire n_46224;
wire n_46225;
wire n_46226;
wire n_46227;
wire n_46228;
wire n_46229;
wire n_46230;
wire n_46231;
wire n_46232;
wire n_46233;
wire n_46234;
wire n_46235;
wire n_46236;
wire n_46237;
wire n_46238;
wire n_46239;
wire n_46240;
wire n_46241;
wire n_46242;
wire n_46243;
wire n_46244;
wire n_46245;
wire n_46246;
wire n_46247;
wire n_46248;
wire n_46249;
wire n_46250;
wire n_46251;
wire n_46252;
wire n_46253;
wire n_46254;
wire n_46255;
wire n_46256;
wire n_46257;
wire n_46258;
wire n_46259;
wire n_46260;
wire n_46261;
wire n_46262;
wire n_46263;
wire n_46264;
wire n_46265;
wire n_46266;
wire n_46267;
wire n_46268;
wire n_46269;
wire n_46270;
wire n_46271;
wire n_46272;
wire n_46273;
wire n_46274;
wire n_46275;
wire n_46276;
wire n_46277;
wire n_46278;
wire n_46279;
wire n_46280;
wire n_46281;
wire n_46282;
wire n_46283;
wire n_46284;
wire n_46285;
wire n_46286;
wire n_46287;
wire n_46288;
wire n_46289;
wire n_46290;
wire n_46291;
wire n_46292;
wire n_46293;
wire n_46294;
wire n_46295;
wire n_46296;
wire n_46297;
wire n_46298;
wire n_46299;
wire n_46300;
wire n_46301;
wire n_46302;
wire n_46303;
wire n_46304;
wire n_46305;
wire n_46306;
wire n_46307;
wire n_46308;
wire n_46309;
wire n_46310;
wire n_46311;
wire n_46312;
wire n_46313;
wire n_46314;
wire n_46315;
wire n_46316;
wire n_46317;
wire n_46318;
wire n_46319;
wire n_46320;
wire n_46321;
wire n_46322;
wire n_46323;
wire n_46324;
wire n_46325;
wire n_46326;
wire n_46327;
wire n_46328;
wire n_46329;
wire n_46330;
wire n_46331;
wire n_46332;
wire n_46333;
wire n_46334;
wire n_46335;
wire n_46336;
wire n_46337;
wire n_46338;
wire n_46339;
wire n_46340;
wire n_46341;
wire n_46342;
wire n_46343;
wire n_46344;
wire n_46345;
wire n_46346;
wire n_46347;
wire n_46348;
wire n_46349;
wire n_46350;
wire n_46351;
wire n_46352;
wire n_46353;
wire n_46354;
wire n_46355;
wire n_46356;
wire n_46357;
wire n_46358;
wire n_46359;
wire n_46360;
wire n_46361;
wire n_46362;
wire n_46363;
wire n_46364;
wire n_46365;
wire n_46366;
wire n_46367;
wire n_46368;
wire n_46369;
wire n_46370;
wire n_46371;
wire n_46372;
wire n_46373;
wire n_46374;
wire n_46375;
wire n_46376;
wire n_46377;
wire n_46378;
wire n_46379;
wire n_46380;
wire n_46381;
wire n_46382;
wire n_46383;
wire n_46384;
wire n_46385;
wire n_46386;
wire n_46387;
wire n_46388;
wire n_46389;
wire n_46390;
wire n_46391;
wire n_46392;
wire n_46393;
wire n_46394;
wire n_46395;
wire n_46396;
wire n_46397;
wire n_46398;
wire n_46399;
wire n_46400;
wire n_46401;
wire n_46402;
wire n_46403;
wire n_46404;
wire n_46405;
wire n_46406;
wire n_46407;
wire n_46408;
wire n_46409;
wire n_46410;
wire n_46411;
wire n_46412;
wire n_46413;
wire n_46414;
wire n_46415;
wire n_46416;
wire n_46417;
wire n_46418;
wire n_46419;
wire n_46420;
wire n_46421;
wire n_46422;
wire n_46423;
wire n_46424;
wire n_46425;
wire n_46426;
wire n_46427;
wire n_46428;
wire n_46429;
wire n_46430;
wire n_46431;
wire n_46432;
wire n_46433;
wire n_46434;
wire n_46435;
wire n_46436;
wire n_46437;
wire n_46438;
wire n_46439;
wire n_46440;
wire n_46441;
wire n_46442;
wire n_46443;
wire n_46444;
wire n_46445;
wire n_46446;
wire n_46447;
wire n_46448;
wire n_46449;
wire n_46450;
wire n_46451;
wire n_46452;
wire n_46453;
wire n_46454;
wire n_46455;
wire n_46456;
wire n_46457;
wire n_46458;
wire n_46459;
wire n_46460;
wire n_46461;
wire n_46462;
wire n_46463;
wire n_46464;
wire n_46465;
wire n_46466;
wire n_46467;
wire n_46468;
wire n_46469;
wire n_46470;
wire n_46471;
wire n_46472;
wire n_46473;
wire n_46474;
wire n_46475;
wire n_46476;
wire n_46477;
wire n_46478;
wire n_46479;
wire n_46480;
wire n_46481;
wire n_46482;
wire n_46483;
wire n_46484;
wire n_46485;
wire n_46486;
wire n_46487;
wire n_46488;
wire n_46489;
wire n_46490;
wire n_46491;
wire n_46492;
wire n_46493;
wire n_46494;
wire n_46495;
wire n_46496;
wire n_46497;
wire n_46498;
wire n_46499;
wire n_46500;
wire n_46501;
wire n_46502;
wire n_46503;
wire n_46504;
wire n_46505;
wire n_46506;
wire n_46507;
wire n_46508;
wire n_46509;
wire n_46510;
wire n_46511;
wire n_46512;
wire n_46513;
wire n_46514;
wire n_46515;
wire n_46516;
wire n_46517;
wire n_46518;
wire n_46519;
wire n_46520;
wire n_46521;
wire n_46522;
wire n_46523;
wire n_46524;
wire n_46525;
wire n_46526;
wire n_46527;
wire n_46528;
wire n_46529;
wire n_46530;
wire n_46531;
wire n_46532;
wire n_46533;
wire n_46534;
wire n_46535;
wire n_46536;
wire n_46537;
wire n_46538;
wire n_46539;
wire n_46540;
wire n_46541;
wire n_46542;
wire n_46543;
wire n_46544;
wire n_46545;
wire n_46546;
wire n_46547;
wire n_46548;
wire n_46549;
wire n_46550;
wire n_46551;
wire n_46552;
wire n_46553;
wire n_46554;
wire n_46555;
wire n_46556;
wire n_46557;
wire n_46558;
wire n_46559;
wire n_46560;
wire n_46561;
wire n_46562;
wire n_46563;
wire n_46564;
wire n_46565;
wire n_46566;
wire n_46567;
wire n_46568;
wire n_46569;
wire n_46570;
wire n_46571;
wire n_46572;
wire n_46573;
wire n_46574;
wire n_46575;
wire n_46576;
wire n_46577;
wire n_46578;
wire n_46579;
wire n_46580;
wire n_46581;
wire n_46582;
wire n_46583;
wire n_46584;
wire n_46585;
wire n_46586;
wire n_46587;
wire n_46588;
wire n_46589;
wire n_46590;
wire n_46591;
wire n_46592;
wire n_46593;
wire n_46594;
wire n_46595;
wire n_46596;
wire n_46597;
wire n_46598;
wire n_46599;
wire n_46600;
wire n_46601;
wire n_46602;
wire n_46603;
wire n_46604;
wire n_46605;
wire n_46606;
wire n_46607;
wire n_46608;
wire n_46609;
wire n_46610;
wire n_46611;
wire n_46612;
wire n_46613;
wire n_46614;
wire n_46615;
wire n_46616;
wire n_46617;
wire n_46618;
wire n_46619;
wire n_46620;
wire n_46621;
wire n_46622;
wire n_46623;
wire n_46624;
wire n_46625;
wire n_46626;
wire n_46627;
wire n_46628;
wire n_46629;
wire n_46630;
wire n_46631;
wire n_46632;
wire n_46633;
wire n_46634;
wire n_46635;
wire n_46636;
wire n_46637;
wire n_46638;
wire n_46639;
wire n_46640;
wire n_46641;
wire n_46642;
wire n_46643;
wire n_46644;
wire n_46645;
wire n_46646;
wire n_46647;
wire n_46648;
wire n_46649;
wire n_46650;
wire n_46651;
wire n_46652;
wire n_46653;
wire n_46654;
wire n_46655;
wire n_46656;
wire n_46657;
wire n_46658;
wire n_46659;
wire n_46660;
wire n_46661;
wire n_46662;
wire n_46663;
wire n_46664;
wire n_46665;
wire n_46666;
wire n_46667;
wire n_46668;
wire n_46669;
wire n_46670;
wire n_46671;
wire n_46672;
wire n_46673;
wire n_46674;
wire n_46675;
wire n_46676;
wire n_46677;
wire n_46678;
wire n_46679;
wire n_46680;
wire n_46681;
wire n_46682;
wire n_46683;
wire n_46684;
wire n_46685;
wire n_46686;
wire n_46687;
wire n_46688;
wire n_46689;
wire n_46690;
wire n_46691;
wire n_46692;
wire n_46693;
wire n_46694;
wire n_46695;
wire n_46696;
wire n_46697;
wire n_46698;
wire n_46699;
wire n_46700;
wire n_46701;
wire n_46702;
wire n_46703;
wire n_46704;
wire n_46705;
wire n_46706;
wire n_46707;
wire n_46708;
wire n_46709;
wire n_46710;
wire n_46711;
wire n_46712;
wire n_46713;
wire n_46714;
wire n_46715;
wire n_46716;
wire n_46717;
wire n_46718;
wire n_46719;
wire n_46720;
wire n_46721;
wire n_46722;
wire n_46723;
wire n_46724;
wire n_46725;
wire n_46726;
wire n_46727;
wire n_46728;
wire n_46729;
wire n_46730;
wire n_46731;
wire n_46732;
wire n_46733;
wire n_46734;
wire n_46735;
wire n_46736;
wire n_46737;
wire n_46738;
wire n_46739;
wire n_46740;
wire n_46741;
wire n_46742;
wire n_46743;
wire n_46744;
wire n_46745;
wire n_46746;
wire n_46747;
wire n_46748;
wire n_46749;
wire n_46750;
wire n_46751;
wire n_46752;
wire n_46753;
wire n_46754;
wire n_46755;
wire n_46756;
wire n_46757;
wire n_46758;
wire n_46759;
wire n_46760;
wire n_46761;
wire n_46762;
wire n_46763;
wire n_46764;
wire n_46765;
wire n_46766;
wire n_46767;
wire n_46768;
wire n_46769;
wire n_46770;
wire n_46771;
wire n_46772;
wire n_46773;
wire n_46774;
wire n_46775;
wire n_46776;
wire n_46777;
wire n_46778;
wire n_46779;
wire n_46780;
wire n_46781;
wire n_46782;
wire n_46783;
wire n_46784;
wire n_46785;
wire n_46786;
wire n_46787;
wire n_46788;
wire n_46789;
wire n_46790;
wire n_46791;
wire n_46792;
wire n_46793;
wire n_46794;
wire n_46795;
wire n_46796;
wire n_46797;
wire n_46798;
wire n_46799;
wire n_46800;
wire n_46801;
wire n_46802;
wire n_46803;
wire n_46804;
wire n_46805;
wire n_46806;
wire n_46807;
wire n_46808;
wire n_46809;
wire n_46810;
wire n_46811;
wire n_46812;
wire n_46813;
wire n_46814;
wire n_46815;
wire n_46816;
wire n_46817;
wire n_46818;
wire n_46819;
wire n_46820;
wire n_46821;
wire n_46822;
wire n_46823;
wire n_46824;
wire n_46825;
wire n_46826;
wire n_46827;
wire n_46828;
wire n_46829;
wire n_46830;
wire n_46831;
wire n_46832;
wire n_46833;
wire n_46834;
wire n_46835;
wire n_46836;
wire n_46837;
wire n_46838;
wire n_46839;
wire n_46840;
wire n_46841;
wire n_46842;
wire n_46843;
wire n_46844;
wire n_46845;
wire n_46846;
wire n_46847;
wire n_46848;
wire n_46849;
wire n_46850;
wire n_46851;
wire n_46852;
wire n_46853;
wire n_46854;
wire n_46855;
wire n_46856;
wire n_46857;
wire n_46858;
wire n_46859;
wire n_46860;
wire n_46861;
wire n_46862;
wire n_46863;
wire n_46864;
wire n_46865;
wire n_46866;
wire n_46867;
wire n_46868;
wire n_46869;
wire n_46870;
wire n_46871;
wire n_46872;
wire n_46873;
wire n_46874;
wire n_46875;
wire n_46876;
wire n_46877;
wire n_46878;
wire n_46879;
wire n_46880;
wire n_46881;
wire n_46882;
wire n_46883;
wire n_46884;
wire n_46885;
wire n_46886;
wire n_46887;
wire n_46888;
wire n_46889;
wire n_46890;
wire n_46891;
wire n_46892;
wire n_46893;
wire n_46894;
wire n_46895;
wire n_46896;
wire n_46897;
wire n_46898;
wire n_46899;
wire n_46900;
wire n_46901;
wire n_46902;
wire n_46903;
wire n_46904;
wire n_46905;
wire n_46906;
wire n_46907;
wire n_46908;
wire n_46909;
wire n_46910;
wire n_46911;
wire n_46912;
wire n_46913;
wire n_46914;
wire n_46915;
wire n_46916;
wire n_46917;
wire n_46918;
wire n_46919;
wire n_46920;
wire n_46921;
wire n_46922;
wire n_46923;
wire n_46924;
wire n_46925;
wire n_46926;
wire n_46927;
wire n_46928;
wire n_46929;
wire n_46930;
wire n_46931;
wire n_46932;
wire n_46933;
wire n_46934;
wire n_46935;
wire n_46936;
wire n_46937;
wire n_46938;
wire n_46939;
wire n_46940;
wire n_46941;
wire n_46942;
wire n_46943;
wire n_46944;
wire n_46945;
wire n_46946;
wire n_46947;
wire n_46948;
wire n_46949;
wire n_46950;
wire n_46951;
wire n_46952;
wire n_46953;
wire n_46954;
wire n_46955;
wire n_46956;
wire n_46957;
wire n_46958;
wire n_46959;
wire n_46960;
wire n_46961;
wire n_46962;
wire n_46963;
wire n_46964;
wire n_46965;
wire n_46966;
wire n_46967;
wire n_46968;
wire n_46969;
wire n_46970;
wire n_46971;
wire n_46972;
wire n_46973;
wire n_46974;
wire n_46975;
wire n_46976;
wire n_46977;
wire n_46978;
wire n_46979;
wire n_46980;
wire n_46981;
wire n_46982;
wire n_46983;
wire n_46984;
wire n_46985;
wire n_46986;
wire n_46987;
wire n_46988;
wire n_46989;
wire n_46990;
wire n_46991;
wire n_46992;
wire n_46993;
wire n_46994;
wire n_46995;
wire n_46996;
wire n_46997;
wire n_46998;
wire n_46999;
wire n_47000;
wire n_47001;
wire n_47002;
wire n_47003;
wire n_47004;
wire n_47005;
wire n_47006;
wire n_47007;
wire n_47008;
wire n_47009;
wire n_47010;
wire n_47011;
wire n_47012;
wire n_47013;
wire n_47014;
wire n_47015;
wire n_47016;
wire n_47017;
wire n_47018;
wire n_47019;
wire n_47020;
wire n_47021;
wire n_47022;
wire n_47023;
wire n_47024;
wire n_47025;
wire n_47026;
wire n_47027;
wire n_47028;
wire n_47029;
wire n_47030;
wire n_47031;
wire n_47032;
wire n_47033;
wire n_47034;
wire n_47035;
wire n_47036;
wire n_47037;
wire n_47038;
wire n_47039;
wire n_47040;
wire n_47041;
wire n_47042;
wire n_47043;
wire n_47044;
wire n_47045;
wire n_47046;
wire n_47047;
wire n_47048;
wire n_47049;
wire n_47050;
wire n_47051;
wire n_47052;
wire n_47053;
wire n_47054;
wire n_47055;
wire n_47056;
wire n_47057;
wire n_47058;
wire n_47059;
wire n_47060;
wire n_47061;
wire n_47062;
wire n_47063;
wire n_47064;
wire n_47065;
wire n_47066;
wire n_47067;
wire n_47068;
wire n_47069;
wire n_47070;
wire n_47071;
wire n_47072;
wire n_47073;
wire n_47074;
wire n_47075;
wire n_47076;
wire n_47077;
wire n_47078;
wire n_47079;
wire n_47080;
wire n_47081;
wire n_47082;
wire n_47083;
wire n_47084;
wire n_47085;
wire n_47086;
wire n_47087;
wire n_47088;
wire n_47089;
wire n_47090;
wire n_47091;
wire n_47092;
wire n_47093;
wire n_47094;
wire n_47095;
wire n_47096;
wire n_47097;
wire n_47098;
wire n_47099;
wire n_47100;
wire n_47101;
wire n_47102;
wire n_47103;
wire n_47104;
wire n_47105;
wire n_47106;
wire n_47107;
wire n_47108;
wire n_47109;
wire n_47110;
wire n_47111;
wire n_47112;
wire n_47113;
wire n_47114;
wire n_47115;
wire n_47116;
wire n_47117;
wire n_47118;
wire n_47119;
wire n_47120;
wire n_47121;
wire n_47122;
wire n_47123;
wire n_47124;
wire n_47125;
wire n_47126;
wire n_47127;
wire n_47128;
wire n_47129;
wire n_47130;
wire n_47131;
wire n_47132;
wire n_47133;
wire n_47134;
wire n_47135;
wire n_47136;
wire n_47137;
wire n_47138;
wire n_47139;
wire n_47140;
wire n_47141;
wire n_47142;
wire n_47143;
wire n_47144;
wire n_47145;
wire n_47146;
wire n_47147;
wire n_47148;
wire n_47149;
wire n_47150;
wire n_47151;
wire n_47152;
wire n_47153;
wire n_47154;
wire n_47155;
wire n_47156;
wire n_47157;
wire n_47158;
wire n_47159;
wire n_47160;
wire n_47161;
wire n_47162;
wire n_47163;
wire n_47164;
wire n_47165;
wire n_47166;
wire n_47167;
wire n_47168;
wire n_47169;
wire n_47170;
wire n_47171;
wire n_47172;
wire n_47173;
wire n_47174;
wire n_47175;
wire n_47176;
wire n_47177;
wire n_47178;
wire n_47179;
wire n_47180;
wire n_47181;
wire n_47182;
wire n_47183;
wire n_47184;
wire n_47185;
wire n_47186;
wire n_47187;
wire n_47188;
wire n_47189;
wire n_47190;
wire n_47191;
wire n_47192;
wire n_47193;
wire n_47194;
wire n_47195;
wire n_47196;
wire n_47197;
wire n_47198;
wire n_47199;
wire n_47200;
wire n_47201;
wire n_47202;
wire n_47203;
wire n_47204;
wire n_47205;
wire n_47206;
wire n_47207;
wire n_47208;
wire n_47209;
wire n_47210;
wire n_47211;
wire n_47212;
wire n_47213;
wire n_47214;
wire n_47215;
wire n_47216;
wire n_47217;
wire n_47218;
wire n_47219;
wire n_47220;
wire n_47221;
wire n_47222;
wire n_47223;
wire n_47224;
wire n_47225;
wire n_47226;
wire n_47227;
wire n_47228;
wire n_47229;
wire n_47230;
wire n_47231;
wire n_47232;
wire n_47233;
wire n_47234;
wire n_47235;
wire n_47236;
wire n_47237;
wire n_47238;
wire n_47239;
wire n_47240;
wire n_47241;
wire n_47242;
wire n_47243;
wire n_47244;
wire n_47245;
wire n_47246;
wire n_47247;
wire n_47248;
wire n_47249;
wire n_47250;
wire n_47251;
wire n_47252;
wire n_47253;
wire n_47254;
wire n_47255;
wire n_47256;
wire n_47257;
wire n_47258;
wire n_47259;
wire n_47260;
wire n_47261;
wire n_47262;
wire n_47263;
wire n_47264;
wire n_47265;
wire n_47266;
wire n_47267;
wire n_47268;
wire n_47269;
wire n_47270;
wire n_47271;
wire n_47272;
wire n_47273;
wire n_47274;
wire n_47275;
wire n_47276;
wire n_47277;
wire n_47278;
wire n_47279;
wire n_47280;
wire n_47281;
wire n_47282;
wire n_47283;
wire n_47284;
wire n_47285;
wire n_47286;
wire n_47287;
wire n_47288;
wire n_47289;
wire n_47290;
wire n_47291;
wire n_47292;
wire n_47293;
wire n_47294;
wire n_47295;
wire n_47296;
wire n_47297;
wire n_47298;
wire n_47299;
wire n_47300;
wire n_47301;
wire n_47302;
wire n_47303;
wire n_47304;
wire n_47305;
wire n_47306;
wire n_47307;
wire n_47308;
wire n_47309;
wire n_47310;
wire n_47311;
wire n_47312;
wire n_47313;
wire n_47314;
wire n_47315;
wire n_47316;
wire n_47317;
wire n_47318;
wire n_47319;
wire n_47320;
wire n_47321;
wire n_47322;
wire n_47323;
wire n_47324;
wire n_47325;
wire n_47326;
wire n_47327;
wire n_47328;
wire n_47329;
wire n_47330;
wire n_47331;
wire n_47332;
wire n_47333;
wire n_47334;
wire n_47335;
wire n_47336;
wire n_47337;
wire n_47338;
wire n_47339;
wire n_47340;
wire n_47341;
wire n_47342;
wire n_47343;
wire n_47344;
wire n_47345;
wire n_47346;
wire n_47347;
wire n_47348;
wire n_47349;
wire n_47350;
wire n_47351;
wire n_47352;
wire n_47353;
wire n_47354;
wire n_47355;
wire n_47356;
wire n_47357;
wire n_47358;
wire n_47359;
wire n_47360;
wire n_47361;
wire n_47362;
wire n_47363;
wire n_47364;
wire n_47365;
wire n_47366;
wire n_47367;
wire n_47368;
wire n_47369;
wire n_47370;
wire n_47371;
wire n_47372;
wire n_47373;
wire n_47374;
wire n_47375;
wire n_47376;
wire n_47377;
wire n_47378;
wire n_47379;
wire n_47380;
wire n_47381;
wire n_47382;
wire n_47383;
wire n_47384;
wire n_47385;
wire n_47386;
wire n_47387;
wire n_47388;
wire n_47389;
wire n_47390;
wire n_47391;
wire n_47392;
wire n_47393;
wire n_47394;
wire n_47395;
wire n_47396;
wire n_47397;
wire n_47398;
wire n_47399;
wire n_47400;
wire n_47401;
wire n_47402;
wire n_47403;
wire n_47404;
wire n_47405;
wire n_47406;
wire n_47407;
wire n_47408;
wire n_47409;
wire n_47410;
wire n_47411;
wire n_47412;
wire n_47413;
wire n_47414;
wire n_47415;
wire n_47416;
wire n_47417;
wire n_47418;
wire n_47419;
wire n_47420;
wire n_47421;
wire n_47422;
wire n_47423;
wire n_47424;
wire n_47425;
wire n_47426;
wire n_47427;
wire n_47428;
wire n_47429;
wire n_47430;
wire n_47431;
wire n_47432;
wire n_47433;
wire n_47434;
wire n_47435;
wire n_47436;
wire n_47437;
wire n_47438;
wire n_47439;
wire n_47440;
wire n_47441;
wire n_47442;
wire n_47443;
wire n_47444;
wire n_47445;
wire n_47446;
wire n_47447;
wire n_47448;
wire n_47449;
wire n_47450;
wire n_47451;
wire n_47452;
wire n_47453;
wire n_47454;
wire n_47455;
wire n_47456;
wire n_47457;
wire n_47458;
wire n_47459;
wire n_47460;
wire n_47461;
wire n_47462;
wire n_47463;
wire n_47464;
wire n_47465;
wire n_47466;
wire n_47467;
wire n_47468;
wire n_47469;
wire n_47470;
wire n_47471;
wire n_47472;
wire n_47473;
wire n_47474;
wire n_47475;
wire n_47476;
wire n_47477;
wire n_47478;
wire n_47479;
wire n_47480;
wire n_47481;
wire n_47482;
wire n_47483;
wire n_47484;
wire n_47485;
wire n_47486;
wire n_47487;
wire n_47488;
wire n_47489;
wire n_47490;
wire n_47491;
wire n_47492;
wire n_47493;
wire n_47494;
wire n_47495;
wire n_47496;
wire n_47497;
wire n_47498;
wire n_47499;
wire n_47500;
wire n_47501;
wire n_47502;
wire n_47503;
wire n_47504;
wire n_47505;
wire n_47506;
wire n_47507;
wire n_47508;
wire n_47509;
wire n_47510;
wire n_47511;
wire n_47512;
wire n_47513;
wire n_47514;
wire n_47515;
wire n_47516;
wire n_47517;
wire n_47518;
wire n_47519;
wire n_47520;
wire n_47521;
wire n_47522;
wire n_47523;
wire n_47524;
wire n_47525;
wire n_47526;
wire n_47527;
wire n_47528;
wire n_47529;
wire n_47530;
wire n_47531;
wire n_47532;
wire n_47533;
wire n_47534;
wire n_47535;
wire n_47536;
wire n_47537;
wire n_47538;
wire n_47539;
wire n_47540;
wire n_47541;
wire n_47542;
wire n_47543;
wire n_47544;
wire n_47545;
wire n_47546;
wire n_47547;
wire n_47548;
wire n_47549;
wire n_47550;
wire n_47551;
wire n_47552;
wire n_47553;
wire n_47554;
wire n_47555;
wire n_47556;
wire n_47557;
wire n_47558;
wire n_47559;
wire n_47560;
wire n_47561;
wire n_47562;
wire n_47563;
wire n_47564;
wire n_47565;
wire n_47566;
wire n_47567;
wire n_47568;
wire n_47569;
wire n_47570;
wire n_47571;
wire n_47572;
wire n_47573;
wire n_47574;
wire n_47575;
wire n_47576;
wire n_47577;
wire n_47578;
wire n_47579;
wire n_47580;
wire n_47581;
wire n_47582;
wire n_47583;
wire n_47584;
wire n_47585;
wire n_47586;
wire n_47587;
wire n_47588;
wire n_47589;
wire n_47590;
wire n_47591;
wire n_47592;
wire n_47593;
wire n_47594;
wire n_47595;
wire n_47596;
wire n_47597;
wire n_47598;
wire n_47599;
wire n_47600;
wire n_47601;
wire n_47602;
wire n_47603;
wire n_47604;
wire n_47605;
wire n_47606;
wire n_47607;
wire n_47608;
wire n_47609;
wire n_47610;
wire n_47611;
wire n_47612;
wire n_47613;
wire n_47614;
wire n_47615;
wire n_47616;
wire n_47617;
wire n_47618;
wire n_47619;
wire n_47620;
wire n_47621;
wire n_47622;
wire n_47623;
wire n_47624;
wire n_47625;
wire n_47626;
wire n_47627;
wire n_47628;
wire n_47629;
wire n_47630;
wire n_47631;
wire n_47632;
wire n_47633;
wire n_47634;
wire n_47635;
wire n_47636;
wire n_47637;
wire n_47638;
wire n_47639;
wire n_47640;
wire n_47641;
wire n_47642;
wire n_47643;
wire n_47644;
wire n_47645;
wire n_47646;
wire n_47647;
wire n_47648;
wire n_47649;
wire n_47650;
wire n_47651;
wire n_47652;
wire n_47653;
wire n_47654;
wire n_47655;
wire n_47656;
wire n_47657;
wire n_47658;
wire n_47659;
wire n_47660;
wire n_47661;
wire n_47662;
wire n_47663;
wire n_47664;
wire n_47665;
wire n_47666;
wire n_47667;
wire n_47668;
wire n_47669;
wire n_47670;
wire n_47671;
wire n_47672;
wire n_47673;
wire n_47674;
wire n_47675;
wire n_47676;
wire n_47677;
wire n_47678;
wire n_47679;
wire n_47680;
wire n_47681;
wire n_47682;
wire n_47683;
wire n_47684;
wire n_47685;
wire n_47686;
wire n_47687;
wire n_47688;
wire n_47689;
wire n_47690;
wire n_47691;
wire n_47692;
wire n_47693;
wire n_47694;
wire n_47695;
wire n_47696;
wire n_47697;
wire n_47698;
wire n_47699;
wire n_47700;
wire n_47701;
wire n_47702;
wire n_47703;
wire n_47704;
wire n_47705;
wire n_47706;
wire n_47707;
wire n_47708;
wire n_47709;
wire n_47710;
wire n_47711;
wire n_47712;
wire n_47713;
wire n_47714;
wire n_47715;
wire n_47716;
wire n_47717;
wire n_47718;
wire n_47719;
wire n_47720;
wire n_47721;
wire n_47722;
wire n_47723;
wire n_47724;
wire n_47725;
wire n_47726;
wire n_47727;
wire n_47728;
wire n_47729;
wire n_47730;
wire n_47731;
wire n_47732;
wire n_47733;
wire n_47734;
wire n_47735;
wire n_47736;
wire n_47737;
wire n_47738;
wire n_47739;
wire n_47740;
wire n_47741;
wire n_47742;
wire n_47743;
wire n_47744;
wire n_47745;
wire n_47746;
wire n_47747;
wire n_47748;
wire n_47749;
wire n_47750;
wire n_47751;
wire n_47752;
wire n_47753;
wire n_47754;
wire n_47755;
wire n_47756;
wire n_47757;
wire n_47758;
wire n_47759;
wire n_47760;
wire n_47761;
wire n_47762;
wire n_47763;
wire n_47764;
wire n_47765;
wire n_47766;
wire n_47767;
wire n_47768;
wire n_47769;
wire n_47770;
wire n_47771;
wire n_47772;
wire n_47773;
wire n_47774;
wire n_47775;
wire n_47776;
wire n_47777;
wire n_47778;
wire n_47779;
wire n_47780;
wire n_47781;
wire n_47782;
wire n_47783;
wire n_47784;
wire n_47785;
wire n_47786;
wire n_47787;
wire n_47788;
wire n_47789;
wire n_47790;
wire n_47791;
wire n_47792;
wire n_47793;
wire n_47794;
wire n_47795;
wire n_47796;
wire n_47797;
wire n_47798;
wire n_47799;
wire n_47800;
wire n_47801;
wire n_47802;
wire n_47803;
wire n_47804;
wire n_47805;
wire n_47806;
wire n_47807;
wire n_47808;
wire n_47809;
wire n_47810;
wire n_47811;
wire n_47812;
wire n_47813;
wire n_47814;
wire n_47815;
wire n_47816;
wire n_47817;
wire n_47818;
wire n_47819;
wire n_47820;
wire n_47821;
wire n_47822;
wire n_47823;
wire n_47824;
wire n_47825;
wire n_47826;
wire n_47827;
wire n_47828;
wire n_47829;
wire n_47830;
wire n_47831;
wire n_47832;
wire n_47833;
wire n_47834;
wire n_47835;
wire n_47836;
wire n_47837;
wire n_47838;
wire n_47839;
wire n_47840;
wire n_47841;
wire n_47842;
wire n_47843;
wire n_47844;
wire n_47845;
wire n_47846;
wire n_47847;
wire n_47848;
wire n_47849;
wire n_47850;
wire n_47851;
wire n_47852;
wire n_47853;
wire n_47854;
wire n_47855;
wire n_47856;
wire n_47857;
wire n_47858;
wire n_47859;
wire n_47860;
wire n_47861;
wire n_47862;
wire n_47863;
wire n_47864;
wire n_47865;
wire n_47866;
wire n_47867;
wire n_47868;
wire n_47869;
wire n_47870;
wire n_47871;
wire n_47872;
wire n_47873;
wire n_47874;
wire n_47875;
wire n_47876;
wire n_47877;
wire n_47878;
wire n_47879;
wire n_47880;
wire n_47881;
wire n_47882;
wire n_47883;
wire n_47884;
wire n_47885;
wire n_47886;
wire n_47887;
wire n_47888;
wire n_47889;
wire n_47890;
wire n_47891;
wire n_47892;
wire n_47893;
wire n_47894;
wire n_47895;
wire n_47896;
wire n_47897;
wire n_47898;
wire n_47899;
wire n_47900;
wire n_47901;
wire n_47902;
wire n_47903;
wire n_47904;
wire n_47905;
wire n_47906;
wire n_47907;
wire n_47908;
wire n_47909;
wire n_47910;
wire n_47911;
wire n_47912;
wire n_47913;
wire n_47914;
wire n_47915;
wire n_47916;
wire n_47917;
wire n_47918;
wire n_47919;
wire n_47920;
wire n_47921;
wire n_47922;
wire n_47923;
wire n_47924;
wire n_47925;
wire n_47926;
wire n_47927;
wire n_47928;
wire n_47929;
wire n_47930;
wire n_47931;
wire n_47932;
wire n_47933;
wire n_47934;
wire n_47935;
wire n_47936;
wire n_47937;
wire n_47938;
wire n_47939;
wire n_47940;
wire n_47941;
wire n_47942;
wire n_47943;
wire n_47944;
wire n_47945;
wire n_47946;
wire n_47947;
wire n_47948;
wire n_47949;
wire n_47950;
wire n_47951;
wire n_47952;
wire n_47953;
wire n_47954;
wire n_47955;
wire n_47956;
wire n_47957;
wire n_47958;
wire n_47959;
wire n_47960;
wire n_47961;
wire n_47962;
wire n_47963;
wire n_47964;
wire n_47965;
wire n_47966;
wire n_47967;
wire n_47968;
wire n_47969;
wire n_47970;
wire n_47971;
wire n_47972;
wire n_47973;
wire n_47974;
wire n_47975;
wire n_47976;
wire n_47977;
wire n_47978;
wire n_47979;
wire n_47980;
wire n_47981;
wire n_47982;
wire n_47983;
wire n_47984;
wire n_47985;
wire n_47986;
wire n_47987;
wire n_47988;
wire n_47989;
wire n_47990;
wire n_47991;
wire n_47992;
wire n_47993;
wire n_47994;
wire n_47995;
wire n_47996;
wire n_47997;
wire n_47998;
wire n_47999;
wire n_48000;
wire n_48001;
wire n_48002;
wire n_48003;
wire n_48004;
wire n_48005;
wire n_48006;
wire n_48007;
wire n_48008;
wire n_48009;
wire n_48010;
wire n_48011;
wire n_48012;
wire n_48013;
wire n_48014;
wire n_48015;
wire n_48016;
wire n_48017;
wire n_48018;
wire n_48019;
wire n_48020;
wire n_48021;
wire n_48022;
wire n_48023;
wire n_48024;
wire n_48025;
wire n_48026;
wire n_48027;
wire n_48028;
wire n_48029;
wire n_48030;
wire n_48031;
wire n_48032;
wire n_48033;
wire n_48034;
wire n_48035;
wire n_48036;
wire n_48037;
wire n_48038;
wire n_48039;
wire n_48040;
wire n_48041;
wire n_48042;
wire n_48043;
wire n_48044;
wire n_48045;
wire n_48046;
wire n_48047;
wire n_48048;
wire n_48049;
wire n_48050;
wire n_48051;
wire n_48052;
wire n_48053;
wire n_48054;
wire n_48055;
wire n_48056;
wire n_48057;
wire n_48058;
wire n_48059;
wire n_48060;
wire n_48061;
wire n_48062;
wire n_48063;
wire n_48064;
wire n_48065;
wire n_48066;
wire n_48067;
wire n_48068;
wire n_48069;
wire n_48070;
wire n_48071;
wire n_48072;
wire n_48073;
wire n_48074;
wire n_48075;
wire n_48076;
wire n_48077;
wire n_48078;
wire n_48079;
wire n_48080;
wire n_48081;
wire n_48082;
wire n_48083;
wire n_48084;
wire n_48085;
wire n_48086;
wire n_48087;
wire n_48088;
wire n_48089;
wire n_48090;
wire n_48091;
wire n_48092;
wire n_48093;
wire n_48094;
wire n_48095;
wire n_48096;
wire n_48097;
wire n_48098;
wire n_48099;
wire n_48100;
wire n_48101;
wire n_48102;
wire n_48103;
wire n_48104;
wire n_48105;
wire n_48106;
wire n_48107;
wire n_48108;
wire n_48109;
wire n_48110;
wire n_48111;
wire n_48112;
wire n_48113;
wire n_48114;
wire n_48115;
wire n_48116;
wire n_48117;
wire n_48118;
wire n_48119;
wire n_48120;
wire n_48121;
wire n_48122;
wire n_48123;
wire n_48124;
wire n_48125;
wire n_48126;
wire n_48127;
wire n_48128;
wire n_48129;
wire n_48130;
wire n_48131;
wire n_48132;
wire n_48133;
wire n_48134;
wire n_48135;
wire n_48136;
wire n_48137;
wire n_48138;
wire n_48139;
wire n_48140;
wire n_48141;
wire n_48142;
wire n_48143;
wire n_48144;
wire n_48145;
wire n_48146;
wire n_48147;
wire n_48148;
wire n_48149;
wire n_48150;
wire n_48151;
wire n_48152;
wire n_48153;
wire n_48154;
wire n_48155;
wire n_48156;
wire n_48157;
wire n_48158;
wire n_48159;
wire n_48160;
wire n_48161;
wire n_48162;
wire n_48163;
wire n_48164;
wire n_48165;
wire n_48166;
wire n_48167;
wire n_48168;
wire n_48169;
wire n_48170;
wire n_48171;
wire n_48172;
wire n_48173;
wire n_48174;
wire n_48175;
wire n_48176;
wire n_48177;
wire n_48178;
wire n_48179;
wire n_48180;
wire n_48181;
wire n_48182;
wire n_48183;
wire n_48184;
wire n_48185;
wire n_48186;
wire n_48187;
wire n_48188;
wire n_48189;
wire n_48190;
wire n_48191;
wire n_48192;
wire n_48193;
wire n_48194;
wire n_48195;
wire n_48196;
wire n_48197;
wire n_48198;
wire n_48199;
wire n_48200;
wire n_48201;
wire n_48202;
wire n_48203;
wire n_48204;
wire n_48205;
wire n_48206;
wire n_48207;
wire n_48208;
wire n_48209;
wire n_48210;
wire n_48211;
wire n_48212;
wire n_48213;
wire n_48214;
wire n_48215;
wire n_48216;
wire n_48217;
wire n_48218;
wire n_48219;
wire n_48220;
wire n_48221;
wire n_48222;
wire n_48223;
wire n_48224;
wire n_48225;
wire n_48226;
wire n_48227;
wire n_48228;
wire n_48229;
wire n_48230;
wire n_48231;
wire n_48232;
wire n_48233;
wire n_48234;
wire n_48235;
wire n_48236;
wire n_48237;
wire n_48238;
wire n_48239;
wire n_48240;
wire n_48241;
wire n_48242;
wire n_48243;
wire n_48244;
wire n_48245;
wire n_48246;
wire n_48247;
wire n_48248;
wire n_48249;
wire n_48250;
wire n_48251;
wire n_48252;
wire n_48253;
wire n_48254;
wire n_48255;
wire n_48256;
wire n_48257;
wire n_48258;
wire n_48259;
wire n_48260;
wire n_48261;
wire n_48262;
wire n_48263;
wire n_48264;
wire n_48265;
wire n_48266;
wire n_48267;
wire n_48268;
wire n_48269;
wire n_48270;
wire n_48271;
wire n_48272;
wire n_48273;
wire n_48274;
wire n_48275;
wire n_48276;
wire n_48277;
wire n_48278;
wire n_48279;
wire n_48280;
wire n_48281;
wire n_48282;
wire n_48283;
wire n_48284;
wire n_48285;
wire n_48286;
wire n_48287;
wire n_48288;
wire n_48289;
wire n_48290;
wire n_48291;
wire n_48292;
wire n_48293;
wire n_48294;
wire n_48295;
wire n_48296;
wire n_48297;
wire n_48298;
wire n_48299;
wire n_48300;
wire n_48301;
wire n_48302;
wire n_48303;
wire n_48304;
wire n_48305;
wire n_48306;
wire n_48307;
wire n_48308;
wire n_48309;
wire n_48310;
wire n_48311;
wire n_48312;
wire n_48313;
wire n_48314;
wire n_48315;
wire n_48316;
wire n_48317;
wire n_48318;
wire n_48319;
wire n_48320;
wire n_48321;
wire n_48322;
wire n_48323;
wire n_48324;
wire n_48325;
wire n_48326;
wire n_48327;
wire n_48328;
wire n_48329;
wire n_48330;
wire n_48331;
wire n_48332;
wire n_48333;
wire n_48334;
wire n_48335;
wire n_48336;
wire n_48337;
wire n_48338;
wire n_48339;
wire n_48340;
wire n_48341;
wire n_48342;
wire n_48343;
wire n_48344;
wire n_48345;
wire n_48346;
wire n_48347;
wire n_48348;
wire n_48349;
wire n_48350;
wire n_48351;
wire n_48352;
wire n_48353;
wire n_48354;
wire n_48355;
wire n_48356;
wire n_48357;
wire n_48358;
wire n_48359;
wire n_48360;
wire n_48361;
wire n_48362;
wire n_48363;
wire n_48364;
wire n_48365;
wire n_48366;
wire n_48367;
wire n_48368;
wire n_48369;
wire n_48370;
wire n_48371;
wire n_48372;
wire n_48373;
wire n_48374;
wire n_48375;
wire n_48376;
wire n_48377;
wire n_48378;
wire n_48379;
wire n_48380;
wire n_48381;
wire n_48382;
wire n_48383;
wire n_48384;
wire n_48385;
wire n_48386;
wire n_48387;
wire n_48388;
wire n_48389;
wire n_48390;
wire n_48391;
wire n_48392;
wire n_48393;
wire n_48394;
wire n_48395;
wire n_48396;
wire n_48397;
wire n_48398;
wire n_48399;
wire n_48400;
wire n_48401;
wire n_48402;
wire n_48403;
wire n_48404;
wire n_48405;
wire n_48406;
wire n_48407;
wire n_48408;
wire n_48409;
wire n_48410;
wire n_48411;
wire n_48412;
wire n_48413;
wire n_48414;
wire n_48415;
wire n_48416;
wire n_48417;
wire n_48418;
wire n_48419;
wire n_48420;
wire n_48421;
wire n_48422;
wire n_48423;
wire n_48424;
wire n_48425;
wire n_48426;
wire n_48427;
wire n_48428;
wire n_48429;
wire n_48430;
wire n_48431;
wire n_48432;
wire n_48433;
wire n_48434;
wire n_48435;
wire n_48436;
wire n_48437;
wire n_48438;
wire n_48439;
wire n_48440;
wire n_48441;
wire n_48442;
wire n_48443;
wire n_48444;
wire n_48445;
wire n_48446;
wire n_48447;
wire n_48448;
wire n_48449;
wire n_48450;
wire n_48451;
wire n_48452;
wire n_48453;
wire n_48454;
wire n_48455;
wire n_48456;
wire n_48457;
wire n_48458;
wire n_48459;
wire n_48460;
wire n_48461;
wire n_48462;
wire n_48463;
wire n_48464;
wire n_48465;
wire n_48466;
wire n_48467;
wire n_48468;
wire n_48469;
wire n_48470;
wire n_48471;
wire n_48472;
wire n_48473;
wire n_48474;
wire n_48475;
wire n_48476;
wire n_48477;
wire n_48478;
wire n_48479;
wire n_48480;
wire n_48481;
wire n_48482;
wire n_48483;
wire n_48484;
wire n_48485;
wire n_48486;
wire n_48487;
wire n_48488;
wire n_48489;
wire n_48490;
wire n_48491;
wire n_48492;
wire n_48493;
wire n_48494;
wire n_48495;
wire n_48496;
wire n_48497;
wire n_48498;
wire n_48499;
wire n_48500;
wire n_48501;
wire n_48502;
wire n_48503;
wire n_48504;
wire n_48505;
wire n_48506;
wire n_48507;
wire n_48508;
wire n_48509;
wire n_48510;
wire n_48511;
wire n_48512;
wire n_48513;
wire n_48514;
wire n_48515;
wire n_48516;
wire n_48517;
wire n_48518;
wire n_48519;
wire n_48520;
wire n_48521;
wire n_48522;
wire n_48523;
wire n_48524;
wire n_48525;
wire n_48526;
wire n_48527;
wire n_48528;
wire n_48529;
wire n_48530;
wire n_48531;
wire n_48532;
wire n_48533;
wire n_48534;
wire n_48535;
wire n_48536;
wire n_48537;
wire n_48538;
wire n_48539;
wire n_48540;
wire n_48541;
wire n_48542;
wire n_48543;
wire n_48544;
wire n_48545;
wire n_48546;
wire n_48547;
wire n_48548;
wire n_48549;
wire n_48550;
wire n_48551;
wire n_48552;
wire n_48553;
wire n_48554;
wire n_48555;
wire n_48556;
wire n_48557;
wire n_48558;
wire n_48559;
wire n_48560;
wire n_48561;
wire n_48562;
wire n_48563;
wire n_48564;
wire n_48565;
wire n_48566;
wire n_48567;
wire n_48568;
wire n_48569;
wire n_48570;
wire n_48571;
wire n_48572;
wire n_48573;
wire n_48574;
wire n_48575;
wire n_48576;
wire n_48577;
wire n_48578;
wire n_48579;
wire n_48580;
wire n_48581;
wire n_48582;
wire n_48583;
wire n_48584;
wire n_48585;
wire n_48586;
wire n_48587;
wire n_48588;
wire n_48589;
wire n_48590;
wire n_48591;
wire n_48592;
wire n_48593;
wire n_48594;
wire n_48595;
wire n_48596;
wire n_48597;
wire n_48598;
wire n_48599;
wire n_48600;
wire n_48601;
wire n_48602;
wire n_48603;
wire n_48604;
wire n_48605;
wire n_48606;
wire n_48607;
wire n_48608;
wire n_48609;
wire n_48610;
wire n_48611;
wire n_48612;
wire n_48613;
wire n_48614;
wire n_48615;
wire n_48616;
wire n_48617;
wire n_48618;
wire n_48619;
wire n_48620;
wire n_48621;
wire n_48622;
wire n_48623;
wire n_48624;
wire n_48625;
wire n_48626;
wire n_48627;
wire n_48628;
wire n_48629;
wire n_48630;
wire n_48631;
wire n_48632;
wire n_48633;
wire n_48634;
wire n_48635;
wire n_48636;
wire n_48637;
wire n_48638;
wire n_48639;
wire n_48640;
wire n_48641;
wire n_48642;
wire n_48643;
wire n_48644;
wire n_48645;
wire n_48646;
wire n_48647;
wire n_48648;
wire n_48649;
wire n_48650;
wire n_48651;
wire n_48652;
wire n_48653;
wire n_48654;
wire n_48655;
wire n_48656;
wire n_48657;
wire n_48658;
assign n_1 = ~x_41 & ~x_42;
assign n_2 =  x_43 &  n_1;
assign n_3 = ~x_34 &  x_35;
assign n_4 = ~x_33 &  x_36;
assign n_5 =  n_3 &  n_4;
assign n_6 =  x_39 & ~x_40;
assign n_7 = ~x_37 &  x_38;
assign n_8 =  n_6 &  n_7;
assign n_9 =  n_5 &  n_8;
assign n_10 =  n_2 &  n_9;
assign n_11 =  x_42 & ~x_43;
assign n_12 = ~x_40 & ~x_41;
assign n_13 =  x_39 &  n_12;
assign n_14 = ~x_37 &  n_5;
assign n_15 =  x_38 &  n_14;
assign n_16 =  n_13 &  n_15;
assign n_17 = ~n_11 &  n_16;
assign n_18 =  x_5063 & ~n_17;
assign n_19 = ~n_10 & ~n_18;
assign n_20 =  x_5063 & ~n_19;
assign n_21 = ~x_5063 &  n_19;
assign n_22 = ~n_20 & ~n_21;
assign n_23 =  x_5062 & ~n_17;
assign n_24 =  x_5062 &  n_23;
assign n_25 = ~x_5062 & ~n_23;
assign n_26 = ~n_24 & ~n_25;
assign n_27 =  x_5061 & ~n_17;
assign n_28 =  x_5061 &  n_27;
assign n_29 = ~x_5061 & ~n_27;
assign n_30 = ~n_28 & ~n_29;
assign n_31 =  x_5060 & ~n_17;
assign n_32 =  x_5060 &  n_31;
assign n_33 = ~x_5060 & ~n_31;
assign n_34 = ~n_32 & ~n_33;
assign n_35 =  x_5059 & ~n_17;
assign n_36 =  x_5059 &  n_35;
assign n_37 = ~x_5059 & ~n_35;
assign n_38 = ~n_36 & ~n_37;
assign n_39 =  x_5058 & ~n_17;
assign n_40 =  x_5058 &  n_39;
assign n_41 = ~x_5058 & ~n_39;
assign n_42 = ~n_40 & ~n_41;
assign n_43 =  x_5057 & ~n_17;
assign n_44 =  x_5057 &  n_43;
assign n_45 = ~x_5057 & ~n_43;
assign n_46 = ~n_44 & ~n_45;
assign n_47 =  x_5056 & ~n_17;
assign n_48 =  x_5056 &  n_47;
assign n_49 = ~x_5056 & ~n_47;
assign n_50 = ~n_48 & ~n_49;
assign n_51 =  x_5055 & ~n_17;
assign n_52 =  x_5055 &  n_51;
assign n_53 = ~x_5055 & ~n_51;
assign n_54 = ~n_52 & ~n_53;
assign n_55 =  x_5054 & ~n_17;
assign n_56 =  x_5054 &  n_55;
assign n_57 = ~x_5054 & ~n_55;
assign n_58 = ~n_56 & ~n_57;
assign n_59 =  x_5053 & ~n_17;
assign n_60 =  x_5053 &  n_59;
assign n_61 = ~x_5053 & ~n_59;
assign n_62 = ~n_60 & ~n_61;
assign n_63 =  x_5052 & ~n_17;
assign n_64 =  x_5052 &  n_63;
assign n_65 = ~x_5052 & ~n_63;
assign n_66 = ~n_64 & ~n_65;
assign n_67 =  x_5051 & ~n_17;
assign n_68 =  x_5051 &  n_67;
assign n_69 = ~x_5051 & ~n_67;
assign n_70 = ~n_68 & ~n_69;
assign n_71 =  x_5050 & ~n_17;
assign n_72 =  x_5050 &  n_71;
assign n_73 = ~x_5050 & ~n_71;
assign n_74 = ~n_72 & ~n_73;
assign n_75 =  x_5049 & ~n_17;
assign n_76 =  x_5049 &  n_75;
assign n_77 = ~x_5049 & ~n_75;
assign n_78 = ~n_76 & ~n_77;
assign n_79 =  x_5048 & ~n_17;
assign n_80 =  x_5048 &  n_79;
assign n_81 = ~x_5048 & ~n_79;
assign n_82 = ~n_80 & ~n_81;
assign n_83 =  x_5047 & ~n_17;
assign n_84 =  x_5047 &  n_83;
assign n_85 = ~x_5047 & ~n_83;
assign n_86 = ~n_84 & ~n_85;
assign n_87 =  x_5046 & ~n_17;
assign n_88 =  x_5046 &  n_87;
assign n_89 = ~x_5046 & ~n_87;
assign n_90 = ~n_88 & ~n_89;
assign n_91 =  x_5045 & ~n_17;
assign n_92 =  x_5045 &  n_91;
assign n_93 = ~x_5045 & ~n_91;
assign n_94 = ~n_92 & ~n_93;
assign n_95 =  x_5044 & ~n_17;
assign n_96 =  x_5044 &  n_95;
assign n_97 = ~x_5044 & ~n_95;
assign n_98 = ~n_96 & ~n_97;
assign n_99 =  x_5043 & ~n_17;
assign n_100 =  x_5043 &  n_99;
assign n_101 = ~x_5043 & ~n_99;
assign n_102 = ~n_100 & ~n_101;
assign n_103 =  x_5042 & ~n_17;
assign n_104 =  x_5042 &  n_103;
assign n_105 = ~x_5042 & ~n_103;
assign n_106 = ~n_104 & ~n_105;
assign n_107 =  x_5041 & ~n_17;
assign n_108 =  x_5041 &  n_107;
assign n_109 = ~x_5041 & ~n_107;
assign n_110 = ~n_108 & ~n_109;
assign n_111 =  x_5040 & ~n_17;
assign n_112 =  x_5040 &  n_111;
assign n_113 = ~x_5040 & ~n_111;
assign n_114 = ~n_112 & ~n_113;
assign n_115 =  x_5039 & ~n_17;
assign n_116 =  x_5039 &  n_115;
assign n_117 = ~x_5039 & ~n_115;
assign n_118 = ~n_116 & ~n_117;
assign n_119 =  x_5038 & ~n_17;
assign n_120 =  x_5038 &  n_119;
assign n_121 = ~x_5038 & ~n_119;
assign n_122 = ~n_120 & ~n_121;
assign n_123 =  x_5037 & ~n_17;
assign n_124 =  x_5037 &  n_123;
assign n_125 = ~x_5037 & ~n_123;
assign n_126 = ~n_124 & ~n_125;
assign n_127 =  x_5036 & ~n_17;
assign n_128 =  x_5036 &  n_127;
assign n_129 = ~x_5036 & ~n_127;
assign n_130 = ~n_128 & ~n_129;
assign n_131 =  x_5035 & ~n_17;
assign n_132 =  x_5035 &  n_131;
assign n_133 = ~x_5035 & ~n_131;
assign n_134 = ~n_132 & ~n_133;
assign n_135 =  x_5034 & ~n_17;
assign n_136 =  x_5034 &  n_135;
assign n_137 = ~x_5034 & ~n_135;
assign n_138 = ~n_136 & ~n_137;
assign n_139 =  x_5033 & ~n_17;
assign n_140 =  x_5033 &  n_139;
assign n_141 = ~x_5033 & ~n_139;
assign n_142 = ~n_140 & ~n_141;
assign n_143 =  x_5032 & ~n_17;
assign n_144 =  x_5032 &  n_143;
assign n_145 = ~x_5032 & ~n_143;
assign n_146 = ~n_144 & ~n_145;
assign n_147 = ~x_33 &  x_34;
assign n_148 = ~x_35 & ~x_36;
assign n_149 = ~x_37 &  n_148;
assign n_150 =  n_147 &  n_149;
assign n_151 = ~x_38 &  x_39;
assign n_152 =  x_41 & ~x_42;
assign n_153 =  x_43 &  n_152;
assign n_154 =  x_40 &  n_153;
assign n_155 =  n_151 &  n_154;
assign n_156 =  n_150 &  n_155;
assign n_157 =  x_5031 & ~n_156;
assign n_158 =  i_32 &  n_156;
assign n_159 = ~n_157 & ~n_158;
assign n_160 =  x_5031 & ~n_159;
assign n_161 = ~x_5031 &  n_159;
assign n_162 = ~n_160 & ~n_161;
assign n_163 =  x_5030 & ~n_156;
assign n_164 =  i_31 &  n_156;
assign n_165 = ~n_163 & ~n_164;
assign n_166 =  x_5030 & ~n_165;
assign n_167 = ~x_5030 &  n_165;
assign n_168 = ~n_166 & ~n_167;
assign n_169 =  x_5029 & ~n_156;
assign n_170 =  i_30 &  n_156;
assign n_171 = ~n_169 & ~n_170;
assign n_172 =  x_5029 & ~n_171;
assign n_173 = ~x_5029 &  n_171;
assign n_174 = ~n_172 & ~n_173;
assign n_175 =  x_5028 & ~n_156;
assign n_176 =  i_29 &  n_156;
assign n_177 = ~n_175 & ~n_176;
assign n_178 =  x_5028 & ~n_177;
assign n_179 = ~x_5028 &  n_177;
assign n_180 = ~n_178 & ~n_179;
assign n_181 =  x_5027 & ~n_156;
assign n_182 =  i_28 &  n_156;
assign n_183 = ~n_181 & ~n_182;
assign n_184 =  x_5027 & ~n_183;
assign n_185 = ~x_5027 &  n_183;
assign n_186 = ~n_184 & ~n_185;
assign n_187 =  x_5026 & ~n_156;
assign n_188 =  i_27 &  n_156;
assign n_189 = ~n_187 & ~n_188;
assign n_190 =  x_5026 & ~n_189;
assign n_191 = ~x_5026 &  n_189;
assign n_192 = ~n_190 & ~n_191;
assign n_193 =  x_5025 & ~n_156;
assign n_194 =  i_26 &  n_156;
assign n_195 = ~n_193 & ~n_194;
assign n_196 =  x_5025 & ~n_195;
assign n_197 = ~x_5025 &  n_195;
assign n_198 = ~n_196 & ~n_197;
assign n_199 =  x_5024 & ~n_156;
assign n_200 =  i_25 &  n_156;
assign n_201 = ~n_199 & ~n_200;
assign n_202 =  x_5024 & ~n_201;
assign n_203 = ~x_5024 &  n_201;
assign n_204 = ~n_202 & ~n_203;
assign n_205 =  x_5023 & ~n_156;
assign n_206 =  i_24 &  n_156;
assign n_207 = ~n_205 & ~n_206;
assign n_208 =  x_5023 & ~n_207;
assign n_209 = ~x_5023 &  n_207;
assign n_210 = ~n_208 & ~n_209;
assign n_211 =  x_5022 & ~n_156;
assign n_212 =  i_23 &  n_156;
assign n_213 = ~n_211 & ~n_212;
assign n_214 =  x_5022 & ~n_213;
assign n_215 = ~x_5022 &  n_213;
assign n_216 = ~n_214 & ~n_215;
assign n_217 =  x_5021 & ~n_156;
assign n_218 =  i_22 &  n_156;
assign n_219 = ~n_217 & ~n_218;
assign n_220 =  x_5021 & ~n_219;
assign n_221 = ~x_5021 &  n_219;
assign n_222 = ~n_220 & ~n_221;
assign n_223 =  x_5020 & ~n_156;
assign n_224 =  i_21 &  n_156;
assign n_225 = ~n_223 & ~n_224;
assign n_226 =  x_5020 & ~n_225;
assign n_227 = ~x_5020 &  n_225;
assign n_228 = ~n_226 & ~n_227;
assign n_229 =  x_5019 & ~n_156;
assign n_230 =  i_20 &  n_156;
assign n_231 = ~n_229 & ~n_230;
assign n_232 =  x_5019 & ~n_231;
assign n_233 = ~x_5019 &  n_231;
assign n_234 = ~n_232 & ~n_233;
assign n_235 =  x_5018 & ~n_156;
assign n_236 =  i_19 &  n_156;
assign n_237 = ~n_235 & ~n_236;
assign n_238 =  x_5018 & ~n_237;
assign n_239 = ~x_5018 &  n_237;
assign n_240 = ~n_238 & ~n_239;
assign n_241 =  x_5017 & ~n_156;
assign n_242 =  i_18 &  n_156;
assign n_243 = ~n_241 & ~n_242;
assign n_244 =  x_5017 & ~n_243;
assign n_245 = ~x_5017 &  n_243;
assign n_246 = ~n_244 & ~n_245;
assign n_247 =  x_5016 & ~n_156;
assign n_248 =  i_17 &  n_156;
assign n_249 = ~n_247 & ~n_248;
assign n_250 =  x_5016 & ~n_249;
assign n_251 = ~x_5016 &  n_249;
assign n_252 = ~n_250 & ~n_251;
assign n_253 =  x_5015 & ~n_156;
assign n_254 =  i_16 &  n_156;
assign n_255 = ~n_253 & ~n_254;
assign n_256 =  x_5015 & ~n_255;
assign n_257 = ~x_5015 &  n_255;
assign n_258 = ~n_256 & ~n_257;
assign n_259 =  x_5014 & ~n_156;
assign n_260 =  i_15 &  n_156;
assign n_261 = ~n_259 & ~n_260;
assign n_262 =  x_5014 & ~n_261;
assign n_263 = ~x_5014 &  n_261;
assign n_264 = ~n_262 & ~n_263;
assign n_265 =  x_5013 & ~n_156;
assign n_266 =  i_14 &  n_156;
assign n_267 = ~n_265 & ~n_266;
assign n_268 =  x_5013 & ~n_267;
assign n_269 = ~x_5013 &  n_267;
assign n_270 = ~n_268 & ~n_269;
assign n_271 =  x_5012 & ~n_156;
assign n_272 =  i_13 &  n_156;
assign n_273 = ~n_271 & ~n_272;
assign n_274 =  x_5012 & ~n_273;
assign n_275 = ~x_5012 &  n_273;
assign n_276 = ~n_274 & ~n_275;
assign n_277 =  x_5011 & ~n_156;
assign n_278 =  i_12 &  n_156;
assign n_279 = ~n_277 & ~n_278;
assign n_280 =  x_5011 & ~n_279;
assign n_281 = ~x_5011 &  n_279;
assign n_282 = ~n_280 & ~n_281;
assign n_283 =  x_5010 & ~n_156;
assign n_284 =  i_11 &  n_156;
assign n_285 = ~n_283 & ~n_284;
assign n_286 =  x_5010 & ~n_285;
assign n_287 = ~x_5010 &  n_285;
assign n_288 = ~n_286 & ~n_287;
assign n_289 =  x_5009 & ~n_156;
assign n_290 =  i_10 &  n_156;
assign n_291 = ~n_289 & ~n_290;
assign n_292 =  x_5009 & ~n_291;
assign n_293 = ~x_5009 &  n_291;
assign n_294 = ~n_292 & ~n_293;
assign n_295 =  x_5008 & ~n_156;
assign n_296 =  i_9 &  n_156;
assign n_297 = ~n_295 & ~n_296;
assign n_298 =  x_5008 & ~n_297;
assign n_299 = ~x_5008 &  n_297;
assign n_300 = ~n_298 & ~n_299;
assign n_301 =  x_5007 & ~n_156;
assign n_302 =  i_8 &  n_156;
assign n_303 = ~n_301 & ~n_302;
assign n_304 =  x_5007 & ~n_303;
assign n_305 = ~x_5007 &  n_303;
assign n_306 = ~n_304 & ~n_305;
assign n_307 =  x_5006 & ~n_156;
assign n_308 =  i_7 &  n_156;
assign n_309 = ~n_307 & ~n_308;
assign n_310 =  x_5006 & ~n_309;
assign n_311 = ~x_5006 &  n_309;
assign n_312 = ~n_310 & ~n_311;
assign n_313 =  x_5005 & ~n_156;
assign n_314 =  i_6 &  n_156;
assign n_315 = ~n_313 & ~n_314;
assign n_316 =  x_5005 & ~n_315;
assign n_317 = ~x_5005 &  n_315;
assign n_318 = ~n_316 & ~n_317;
assign n_319 =  x_5004 & ~n_156;
assign n_320 =  i_5 &  n_156;
assign n_321 = ~n_319 & ~n_320;
assign n_322 =  x_5004 & ~n_321;
assign n_323 = ~x_5004 &  n_321;
assign n_324 = ~n_322 & ~n_323;
assign n_325 =  x_5003 & ~n_156;
assign n_326 =  i_4 &  n_156;
assign n_327 = ~n_325 & ~n_326;
assign n_328 =  x_5003 & ~n_327;
assign n_329 = ~x_5003 &  n_327;
assign n_330 = ~n_328 & ~n_329;
assign n_331 =  x_5002 & ~n_156;
assign n_332 =  i_3 &  n_156;
assign n_333 = ~n_331 & ~n_332;
assign n_334 =  x_5002 & ~n_333;
assign n_335 = ~x_5002 &  n_333;
assign n_336 = ~n_334 & ~n_335;
assign n_337 =  x_5001 & ~n_156;
assign n_338 =  i_2 &  n_156;
assign n_339 = ~n_337 & ~n_338;
assign n_340 =  x_5001 & ~n_339;
assign n_341 = ~x_5001 &  n_339;
assign n_342 = ~n_340 & ~n_341;
assign n_343 =  x_5000 & ~n_156;
assign n_344 =  i_1 &  n_156;
assign n_345 = ~n_343 & ~n_344;
assign n_346 =  x_5000 & ~n_345;
assign n_347 = ~x_5000 &  n_345;
assign n_348 = ~n_346 & ~n_347;
assign n_349 = ~x_42 & ~x_43;
assign n_350 =  x_40 & ~x_41;
assign n_351 =  n_349 &  n_350;
assign n_352 = ~x_33 & ~x_34;
assign n_353 = ~x_35 &  x_36;
assign n_354 =  n_352 &  n_353;
assign n_355 =  x_37 &  n_354;
assign n_356 = ~x_38 &  n_355;
assign n_357 = ~x_39 &  n_356;
assign n_358 =  n_351 &  n_357;
assign n_359 =  x_4999 & ~n_358;
assign n_360 =  x_2058 &  n_358;
assign n_361 = ~n_359 & ~n_360;
assign n_362 =  x_4999 & ~n_361;
assign n_363 = ~x_4999 &  n_361;
assign n_364 = ~n_362 & ~n_363;
assign n_365 =  x_4998 & ~n_358;
assign n_366 =  x_2057 &  n_358;
assign n_367 = ~n_365 & ~n_366;
assign n_368 =  x_4998 & ~n_367;
assign n_369 = ~x_4998 &  n_367;
assign n_370 = ~n_368 & ~n_369;
assign n_371 =  x_4997 & ~n_358;
assign n_372 =  x_2056 &  n_358;
assign n_373 = ~n_371 & ~n_372;
assign n_374 =  x_4997 & ~n_373;
assign n_375 = ~x_4997 &  n_373;
assign n_376 = ~n_374 & ~n_375;
assign n_377 =  x_4996 & ~n_358;
assign n_378 =  x_2055 &  n_358;
assign n_379 = ~n_377 & ~n_378;
assign n_380 =  x_4996 & ~n_379;
assign n_381 = ~x_4996 &  n_379;
assign n_382 = ~n_380 & ~n_381;
assign n_383 =  x_4995 & ~n_358;
assign n_384 =  x_2054 &  n_358;
assign n_385 = ~n_383 & ~n_384;
assign n_386 =  x_4995 & ~n_385;
assign n_387 = ~x_4995 &  n_385;
assign n_388 = ~n_386 & ~n_387;
assign n_389 =  x_4994 & ~n_358;
assign n_390 =  x_2053 &  n_358;
assign n_391 = ~n_389 & ~n_390;
assign n_392 =  x_4994 & ~n_391;
assign n_393 = ~x_4994 &  n_391;
assign n_394 = ~n_392 & ~n_393;
assign n_395 =  x_4993 & ~n_358;
assign n_396 =  x_2052 &  n_358;
assign n_397 = ~n_395 & ~n_396;
assign n_398 =  x_4993 & ~n_397;
assign n_399 = ~x_4993 &  n_397;
assign n_400 = ~n_398 & ~n_399;
assign n_401 =  x_4992 & ~n_358;
assign n_402 =  x_2051 &  n_358;
assign n_403 = ~n_401 & ~n_402;
assign n_404 =  x_4992 & ~n_403;
assign n_405 = ~x_4992 &  n_403;
assign n_406 = ~n_404 & ~n_405;
assign n_407 =  x_4991 & ~n_358;
assign n_408 =  x_2050 &  n_358;
assign n_409 = ~n_407 & ~n_408;
assign n_410 =  x_4991 & ~n_409;
assign n_411 = ~x_4991 &  n_409;
assign n_412 = ~n_410 & ~n_411;
assign n_413 =  x_4990 & ~n_358;
assign n_414 =  x_2049 &  n_358;
assign n_415 = ~n_413 & ~n_414;
assign n_416 =  x_4990 & ~n_415;
assign n_417 = ~x_4990 &  n_415;
assign n_418 = ~n_416 & ~n_417;
assign n_419 =  x_4989 & ~n_358;
assign n_420 =  x_2048 &  n_358;
assign n_421 = ~n_419 & ~n_420;
assign n_422 =  x_4989 & ~n_421;
assign n_423 = ~x_4989 &  n_421;
assign n_424 = ~n_422 & ~n_423;
assign n_425 =  x_4988 & ~n_358;
assign n_426 =  x_2047 &  n_358;
assign n_427 = ~n_425 & ~n_426;
assign n_428 =  x_4988 & ~n_427;
assign n_429 = ~x_4988 &  n_427;
assign n_430 = ~n_428 & ~n_429;
assign n_431 =  x_4987 & ~n_358;
assign n_432 =  x_2046 &  n_358;
assign n_433 = ~n_431 & ~n_432;
assign n_434 =  x_4987 & ~n_433;
assign n_435 = ~x_4987 &  n_433;
assign n_436 = ~n_434 & ~n_435;
assign n_437 =  x_4986 & ~n_358;
assign n_438 =  x_2045 &  n_358;
assign n_439 = ~n_437 & ~n_438;
assign n_440 =  x_4986 & ~n_439;
assign n_441 = ~x_4986 &  n_439;
assign n_442 = ~n_440 & ~n_441;
assign n_443 =  x_4985 & ~n_358;
assign n_444 =  x_2044 &  n_358;
assign n_445 = ~n_443 & ~n_444;
assign n_446 =  x_4985 & ~n_445;
assign n_447 = ~x_4985 &  n_445;
assign n_448 = ~n_446 & ~n_447;
assign n_449 =  x_4984 & ~n_358;
assign n_450 =  x_2043 &  n_358;
assign n_451 = ~n_449 & ~n_450;
assign n_452 =  x_4984 & ~n_451;
assign n_453 = ~x_4984 &  n_451;
assign n_454 = ~n_452 & ~n_453;
assign n_455 =  x_4983 & ~n_358;
assign n_456 =  x_2042 &  n_358;
assign n_457 = ~n_455 & ~n_456;
assign n_458 =  x_4983 & ~n_457;
assign n_459 = ~x_4983 &  n_457;
assign n_460 = ~n_458 & ~n_459;
assign n_461 =  x_4982 & ~n_358;
assign n_462 =  x_2041 &  n_358;
assign n_463 = ~n_461 & ~n_462;
assign n_464 =  x_4982 & ~n_463;
assign n_465 = ~x_4982 &  n_463;
assign n_466 = ~n_464 & ~n_465;
assign n_467 =  x_4981 & ~n_358;
assign n_468 =  x_2040 &  n_358;
assign n_469 = ~n_467 & ~n_468;
assign n_470 =  x_4981 & ~n_469;
assign n_471 = ~x_4981 &  n_469;
assign n_472 = ~n_470 & ~n_471;
assign n_473 =  x_4980 & ~n_358;
assign n_474 =  x_2039 &  n_358;
assign n_475 = ~n_473 & ~n_474;
assign n_476 =  x_4980 & ~n_475;
assign n_477 = ~x_4980 &  n_475;
assign n_478 = ~n_476 & ~n_477;
assign n_479 =  x_4979 & ~n_358;
assign n_480 =  x_2038 &  n_358;
assign n_481 = ~n_479 & ~n_480;
assign n_482 =  x_4979 & ~n_481;
assign n_483 = ~x_4979 &  n_481;
assign n_484 = ~n_482 & ~n_483;
assign n_485 =  x_4978 & ~n_358;
assign n_486 =  x_2037 &  n_358;
assign n_487 = ~n_485 & ~n_486;
assign n_488 =  x_4978 & ~n_487;
assign n_489 = ~x_4978 &  n_487;
assign n_490 = ~n_488 & ~n_489;
assign n_491 =  x_4977 & ~n_358;
assign n_492 =  x_2036 &  n_358;
assign n_493 = ~n_491 & ~n_492;
assign n_494 =  x_4977 & ~n_493;
assign n_495 = ~x_4977 &  n_493;
assign n_496 = ~n_494 & ~n_495;
assign n_497 =  x_4976 & ~n_358;
assign n_498 =  x_2035 &  n_358;
assign n_499 = ~n_497 & ~n_498;
assign n_500 =  x_4976 & ~n_499;
assign n_501 = ~x_4976 &  n_499;
assign n_502 = ~n_500 & ~n_501;
assign n_503 =  x_4975 & ~n_358;
assign n_504 =  x_2034 &  n_358;
assign n_505 = ~n_503 & ~n_504;
assign n_506 =  x_4975 & ~n_505;
assign n_507 = ~x_4975 &  n_505;
assign n_508 = ~n_506 & ~n_507;
assign n_509 =  x_4974 & ~n_358;
assign n_510 =  x_2033 &  n_358;
assign n_511 = ~n_509 & ~n_510;
assign n_512 =  x_4974 & ~n_511;
assign n_513 = ~x_4974 &  n_511;
assign n_514 = ~n_512 & ~n_513;
assign n_515 =  x_4973 & ~n_358;
assign n_516 =  x_2032 &  n_358;
assign n_517 = ~n_515 & ~n_516;
assign n_518 =  x_4973 & ~n_517;
assign n_519 = ~x_4973 &  n_517;
assign n_520 = ~n_518 & ~n_519;
assign n_521 =  x_4972 & ~n_358;
assign n_522 =  x_2031 &  n_358;
assign n_523 = ~n_521 & ~n_522;
assign n_524 =  x_4972 & ~n_523;
assign n_525 = ~x_4972 &  n_523;
assign n_526 = ~n_524 & ~n_525;
assign n_527 =  x_4971 & ~n_358;
assign n_528 =  x_2030 &  n_358;
assign n_529 = ~n_527 & ~n_528;
assign n_530 =  x_4971 & ~n_529;
assign n_531 = ~x_4971 &  n_529;
assign n_532 = ~n_530 & ~n_531;
assign n_533 =  x_4970 & ~n_358;
assign n_534 =  x_2029 &  n_358;
assign n_535 = ~n_533 & ~n_534;
assign n_536 =  x_4970 & ~n_535;
assign n_537 = ~x_4970 &  n_535;
assign n_538 = ~n_536 & ~n_537;
assign n_539 =  x_4969 & ~n_358;
assign n_540 =  x_2028 &  n_358;
assign n_541 = ~n_539 & ~n_540;
assign n_542 =  x_4969 & ~n_541;
assign n_543 = ~x_4969 &  n_541;
assign n_544 = ~n_542 & ~n_543;
assign n_545 =  x_4968 & ~n_358;
assign n_546 =  x_2027 &  n_358;
assign n_547 = ~n_545 & ~n_546;
assign n_548 =  x_4968 & ~n_547;
assign n_549 = ~x_4968 &  n_547;
assign n_550 = ~n_548 & ~n_549;
assign n_551 =  n_352 &  n_148;
assign n_552 =  x_37 &  n_551;
assign n_553 =  x_41 &  x_42;
assign n_554 = ~x_43 &  n_553;
assign n_555 = ~x_40 &  n_554;
assign n_556 =  x_38 &  x_39;
assign n_557 =  n_555 &  n_556;
assign n_558 =  n_552 &  n_557;
assign n_559 =  x_811 &  n_558;
assign n_560 =  n_556 &  n_552;
assign n_561 = ~x_40 &  x_41;
assign n_562 = ~n_561 & ~n_350;
assign n_563 =  n_11 & ~n_562;
assign n_564 =  n_560 &  n_563;
assign n_565 =  x_4967 & ~n_564;
assign n_566 = ~n_559 & ~n_565;
assign n_567 =  x_4967 & ~n_566;
assign n_568 = ~x_4967 &  n_566;
assign n_569 = ~n_567 & ~n_568;
assign n_570 =  x_810 &  n_558;
assign n_571 =  x_4966 & ~n_564;
assign n_572 = ~n_570 & ~n_571;
assign n_573 =  x_4966 & ~n_572;
assign n_574 = ~x_4966 &  n_572;
assign n_575 = ~n_573 & ~n_574;
assign n_576 =  x_809 &  n_558;
assign n_577 =  x_4965 & ~n_564;
assign n_578 = ~n_576 & ~n_577;
assign n_579 =  x_4965 & ~n_578;
assign n_580 = ~x_4965 &  n_578;
assign n_581 = ~n_579 & ~n_580;
assign n_582 =  x_808 &  n_558;
assign n_583 =  x_4964 & ~n_564;
assign n_584 = ~n_582 & ~n_583;
assign n_585 =  x_4964 & ~n_584;
assign n_586 = ~x_4964 &  n_584;
assign n_587 = ~n_585 & ~n_586;
assign n_588 =  x_807 &  n_558;
assign n_589 =  x_4963 & ~n_564;
assign n_590 = ~n_588 & ~n_589;
assign n_591 =  x_4963 & ~n_590;
assign n_592 = ~x_4963 &  n_590;
assign n_593 = ~n_591 & ~n_592;
assign n_594 =  x_806 &  n_558;
assign n_595 =  x_4962 & ~n_564;
assign n_596 = ~n_594 & ~n_595;
assign n_597 =  x_4962 & ~n_596;
assign n_598 = ~x_4962 &  n_596;
assign n_599 = ~n_597 & ~n_598;
assign n_600 =  x_805 &  n_558;
assign n_601 =  x_4961 & ~n_564;
assign n_602 = ~n_600 & ~n_601;
assign n_603 =  x_4961 & ~n_602;
assign n_604 = ~x_4961 &  n_602;
assign n_605 = ~n_603 & ~n_604;
assign n_606 =  x_804 &  n_558;
assign n_607 =  x_4960 & ~n_564;
assign n_608 = ~n_606 & ~n_607;
assign n_609 =  x_4960 & ~n_608;
assign n_610 = ~x_4960 &  n_608;
assign n_611 = ~n_609 & ~n_610;
assign n_612 =  x_803 &  n_558;
assign n_613 =  x_4959 & ~n_564;
assign n_614 = ~n_612 & ~n_613;
assign n_615 =  x_4959 & ~n_614;
assign n_616 = ~x_4959 &  n_614;
assign n_617 = ~n_615 & ~n_616;
assign n_618 =  x_802 &  n_558;
assign n_619 =  x_4958 & ~n_564;
assign n_620 = ~n_618 & ~n_619;
assign n_621 =  x_4958 & ~n_620;
assign n_622 = ~x_4958 &  n_620;
assign n_623 = ~n_621 & ~n_622;
assign n_624 =  x_801 &  n_558;
assign n_625 =  x_4957 & ~n_564;
assign n_626 = ~n_624 & ~n_625;
assign n_627 =  x_4957 & ~n_626;
assign n_628 = ~x_4957 &  n_626;
assign n_629 = ~n_627 & ~n_628;
assign n_630 =  x_800 &  n_558;
assign n_631 =  x_4956 & ~n_564;
assign n_632 = ~n_630 & ~n_631;
assign n_633 =  x_4956 & ~n_632;
assign n_634 = ~x_4956 &  n_632;
assign n_635 = ~n_633 & ~n_634;
assign n_636 =  x_799 &  n_558;
assign n_637 =  x_4955 & ~n_564;
assign n_638 = ~n_636 & ~n_637;
assign n_639 =  x_4955 & ~n_638;
assign n_640 = ~x_4955 &  n_638;
assign n_641 = ~n_639 & ~n_640;
assign n_642 =  x_798 &  n_558;
assign n_643 =  x_4954 & ~n_564;
assign n_644 = ~n_642 & ~n_643;
assign n_645 =  x_4954 & ~n_644;
assign n_646 = ~x_4954 &  n_644;
assign n_647 = ~n_645 & ~n_646;
assign n_648 =  x_797 &  n_558;
assign n_649 =  x_4953 & ~n_564;
assign n_650 = ~n_648 & ~n_649;
assign n_651 =  x_4953 & ~n_650;
assign n_652 = ~x_4953 &  n_650;
assign n_653 = ~n_651 & ~n_652;
assign n_654 =  x_796 &  n_558;
assign n_655 =  x_4952 & ~n_564;
assign n_656 = ~n_654 & ~n_655;
assign n_657 =  x_4952 & ~n_656;
assign n_658 = ~x_4952 &  n_656;
assign n_659 = ~n_657 & ~n_658;
assign n_660 =  x_795 &  n_558;
assign n_661 =  x_4951 & ~n_564;
assign n_662 = ~n_660 & ~n_661;
assign n_663 =  x_4951 & ~n_662;
assign n_664 = ~x_4951 &  n_662;
assign n_665 = ~n_663 & ~n_664;
assign n_666 =  x_794 &  n_558;
assign n_667 =  x_4950 & ~n_564;
assign n_668 = ~n_666 & ~n_667;
assign n_669 =  x_4950 & ~n_668;
assign n_670 = ~x_4950 &  n_668;
assign n_671 = ~n_669 & ~n_670;
assign n_672 =  x_793 &  n_558;
assign n_673 =  x_4949 & ~n_564;
assign n_674 = ~n_672 & ~n_673;
assign n_675 =  x_4949 & ~n_674;
assign n_676 = ~x_4949 &  n_674;
assign n_677 = ~n_675 & ~n_676;
assign n_678 =  x_792 &  n_558;
assign n_679 =  x_4948 & ~n_564;
assign n_680 = ~n_678 & ~n_679;
assign n_681 =  x_4948 & ~n_680;
assign n_682 = ~x_4948 &  n_680;
assign n_683 = ~n_681 & ~n_682;
assign n_684 =  x_791 &  n_558;
assign n_685 =  x_4947 & ~n_564;
assign n_686 = ~n_684 & ~n_685;
assign n_687 =  x_4947 & ~n_686;
assign n_688 = ~x_4947 &  n_686;
assign n_689 = ~n_687 & ~n_688;
assign n_690 =  x_790 &  n_558;
assign n_691 =  x_4946 & ~n_564;
assign n_692 = ~n_690 & ~n_691;
assign n_693 =  x_4946 & ~n_692;
assign n_694 = ~x_4946 &  n_692;
assign n_695 = ~n_693 & ~n_694;
assign n_696 =  x_789 &  n_558;
assign n_697 =  x_4945 & ~n_564;
assign n_698 = ~n_696 & ~n_697;
assign n_699 =  x_4945 & ~n_698;
assign n_700 = ~x_4945 &  n_698;
assign n_701 = ~n_699 & ~n_700;
assign n_702 =  x_788 &  n_558;
assign n_703 =  x_4944 & ~n_564;
assign n_704 = ~n_702 & ~n_703;
assign n_705 =  x_4944 & ~n_704;
assign n_706 = ~x_4944 &  n_704;
assign n_707 = ~n_705 & ~n_706;
assign n_708 =  x_787 &  n_558;
assign n_709 =  x_4943 & ~n_564;
assign n_710 = ~n_708 & ~n_709;
assign n_711 =  x_4943 & ~n_710;
assign n_712 = ~x_4943 &  n_710;
assign n_713 = ~n_711 & ~n_712;
assign n_714 =  x_786 &  n_558;
assign n_715 =  x_4942 & ~n_564;
assign n_716 = ~n_714 & ~n_715;
assign n_717 =  x_4942 & ~n_716;
assign n_718 = ~x_4942 &  n_716;
assign n_719 = ~n_717 & ~n_718;
assign n_720 =  x_785 &  n_558;
assign n_721 =  x_4941 & ~n_564;
assign n_722 = ~n_720 & ~n_721;
assign n_723 =  x_4941 & ~n_722;
assign n_724 = ~x_4941 &  n_722;
assign n_725 = ~n_723 & ~n_724;
assign n_726 =  x_784 &  n_558;
assign n_727 =  x_4940 & ~n_564;
assign n_728 = ~n_726 & ~n_727;
assign n_729 =  x_4940 & ~n_728;
assign n_730 = ~x_4940 &  n_728;
assign n_731 = ~n_729 & ~n_730;
assign n_732 =  x_783 &  n_558;
assign n_733 =  x_4939 & ~n_564;
assign n_734 = ~n_732 & ~n_733;
assign n_735 =  x_4939 & ~n_734;
assign n_736 = ~x_4939 &  n_734;
assign n_737 = ~n_735 & ~n_736;
assign n_738 =  x_782 &  n_558;
assign n_739 =  x_4938 & ~n_564;
assign n_740 = ~n_738 & ~n_739;
assign n_741 =  x_4938 & ~n_740;
assign n_742 = ~x_4938 &  n_740;
assign n_743 = ~n_741 & ~n_742;
assign n_744 =  x_781 &  n_558;
assign n_745 =  x_4937 & ~n_564;
assign n_746 = ~n_744 & ~n_745;
assign n_747 =  x_4937 & ~n_746;
assign n_748 = ~x_4937 &  n_746;
assign n_749 = ~n_747 & ~n_748;
assign n_750 =  x_780 &  n_558;
assign n_751 =  x_4936 & ~n_564;
assign n_752 = ~n_750 & ~n_751;
assign n_753 =  x_4936 & ~n_752;
assign n_754 = ~x_4936 &  n_752;
assign n_755 = ~n_753 & ~n_754;
assign n_756 = ~x_37 & ~x_38;
assign n_757 =  n_756 &  n_551;
assign n_758 = ~x_43 &  n_1;
assign n_759 = ~x_39 & ~x_40;
assign n_760 =  n_758 &  n_759;
assign n_761 =  n_757 &  n_760;
assign n_762 =  n_759 &  n_757;
assign n_763 = ~x_41 &  n_762;
assign n_764 =  x_35 & ~x_36;
assign n_765 =  n_764 &  n_352;
assign n_766 =  x_40 &  x_41;
assign n_767 =  x_37 &  x_38;
assign n_768 = ~x_39 &  n_767;
assign n_769 =  n_766 &  n_768;
assign n_770 =  n_765 &  n_769;
assign n_771 = ~x_1585 & ~x_3230;
assign n_772 =  x_1585 &  x_3230;
assign n_773 = ~n_771 & ~n_772;
assign n_774 = ~x_1598 & ~x_3243;
assign n_775 =  x_1598 &  x_3243;
assign n_776 = ~n_774 & ~n_775;
assign n_777 = ~n_773 & ~n_776;
assign n_778 = ~x_1603 & ~x_3248;
assign n_779 =  x_1603 &  x_3248;
assign n_780 = ~n_778 & ~n_779;
assign n_781 = ~x_1610 & ~x_3255;
assign n_782 =  x_1610 &  x_3255;
assign n_783 = ~n_781 & ~n_782;
assign n_784 = ~n_780 & ~n_783;
assign n_785 =  n_777 &  n_784;
assign n_786 = ~x_1583 & ~x_3228;
assign n_787 =  x_1583 &  x_3228;
assign n_788 = ~n_786 & ~n_787;
assign n_789 = ~x_1582 &  x_3227;
assign n_790 = ~x_1594 &  x_3239;
assign n_791 = ~n_789 & ~n_790;
assign n_792 = ~n_788 &  n_791;
assign n_793 = ~x_1604 & ~x_3249;
assign n_794 =  x_1604 &  x_3249;
assign n_795 = ~n_793 & ~n_794;
assign n_796 = ~x_1579 & ~x_3224;
assign n_797 =  x_1579 &  x_3224;
assign n_798 = ~n_796 & ~n_797;
assign n_799 = ~n_795 & ~n_798;
assign n_800 =  n_792 &  n_799;
assign n_801 =  n_785 &  n_800;
assign n_802 =  n_770 &  n_801;
assign n_803 = ~x_1596 &  x_3241;
assign n_804 =  x_1601 & ~x_3246;
assign n_805 = ~n_803 & ~n_804;
assign n_806 = ~x_1601 &  x_3246;
assign n_807 = ~x_1607 &  x_3252;
assign n_808 = ~n_806 & ~n_807;
assign n_809 =  n_805 &  n_808;
assign n_810 =  x_1591 & ~x_3236;
assign n_811 =  x_1606 & ~x_3251;
assign n_812 = ~n_810 & ~n_811;
assign n_813 = ~x_1606 &  x_3251;
assign n_814 =  x_1596 & ~x_3241;
assign n_815 = ~n_813 & ~n_814;
assign n_816 =  n_812 &  n_815;
assign n_817 =  n_809 &  n_816;
assign n_818 =  x_1609 & ~x_3254;
assign n_819 = ~x_1609 &  x_3254;
assign n_820 = ~n_818 & ~n_819;
assign n_821 =  x_1599 & ~x_3244;
assign n_822 = ~x_1599 &  x_3244;
assign n_823 = ~n_821 & ~n_822;
assign n_824 =  n_820 &  n_823;
assign n_825 =  x_1586 & ~x_3231;
assign n_826 =  x_1607 & ~x_3252;
assign n_827 = ~n_825 & ~n_826;
assign n_828 =  x_1595 & ~x_3240;
assign n_829 = ~x_1595 &  x_3240;
assign n_830 = ~n_828 & ~n_829;
assign n_831 =  n_827 &  n_830;
assign n_832 =  n_824 &  n_831;
assign n_833 =  n_817 &  n_832;
assign n_834 = ~x_1608 &  x_3253;
assign n_835 =  x_1587 & ~x_3232;
assign n_836 = ~n_834 & ~n_835;
assign n_837 = ~x_1587 &  x_3232;
assign n_838 =  x_1584 & ~x_3229;
assign n_839 = ~n_837 & ~n_838;
assign n_840 =  n_836 &  n_839;
assign n_841 = ~x_1590 &  x_3235;
assign n_842 = ~x_1597 &  x_3242;
assign n_843 = ~n_841 & ~n_842;
assign n_844 =  x_1602 & ~x_3247;
assign n_845 =  x_1608 & ~x_3253;
assign n_846 = ~n_844 & ~n_845;
assign n_847 =  n_843 &  n_846;
assign n_848 =  n_840 &  n_847;
assign n_849 = ~x_1592 &  x_3237;
assign n_850 = ~x_1586 &  x_3231;
assign n_851 = ~n_849 & ~n_850;
assign n_852 =  x_1592 & ~x_3237;
assign n_853 =  x_1605 & ~x_3250;
assign n_854 = ~n_852 & ~n_853;
assign n_855 =  n_851 &  n_854;
assign n_856 = ~x_1584 &  x_3229;
assign n_857 = ~x_1605 &  x_3250;
assign n_858 = ~n_856 & ~n_857;
assign n_859 =  x_1582 & ~x_3227;
assign n_860 = ~x_1591 &  x_3236;
assign n_861 = ~n_859 & ~n_860;
assign n_862 =  n_858 &  n_861;
assign n_863 =  n_855 &  n_862;
assign n_864 =  n_848 &  n_863;
assign n_865 =  x_1593 & ~x_3238;
assign n_866 = ~x_1593 &  x_3238;
assign n_867 = ~n_865 & ~n_866;
assign n_868 = ~x_1589 &  x_3234;
assign n_869 =  x_1600 & ~x_3245;
assign n_870 = ~n_868 & ~n_869;
assign n_871 =  n_867 &  n_870;
assign n_872 =  x_1580 & ~x_3225;
assign n_873 = ~x_1580 &  x_3225;
assign n_874 = ~n_872 & ~n_873;
assign n_875 =  x_1588 & ~x_3233;
assign n_876 = ~x_1588 &  x_3233;
assign n_877 = ~n_875 & ~n_876;
assign n_878 =  n_874 &  n_877;
assign n_879 =  n_871 &  n_878;
assign n_880 =  x_1597 & ~x_3242;
assign n_881 =  x_1594 & ~x_3239;
assign n_882 = ~n_880 & ~n_881;
assign n_883 = ~x_1602 &  x_3247;
assign n_884 =  x_1590 & ~x_3235;
assign n_885 = ~n_883 & ~n_884;
assign n_886 =  n_882 &  n_885;
assign n_887 =  x_1589 & ~x_3234;
assign n_888 = ~x_1581 &  x_3226;
assign n_889 = ~n_887 & ~n_888;
assign n_890 = ~x_1600 &  x_3245;
assign n_891 =  x_1581 & ~x_3226;
assign n_892 = ~n_890 & ~n_891;
assign n_893 =  n_889 &  n_892;
assign n_894 =  n_886 &  n_893;
assign n_895 =  n_879 &  n_894;
assign n_896 =  n_864 &  n_895;
assign n_897 =  n_833 &  n_896;
assign n_898 =  n_802 &  n_897;
assign n_899 = ~n_763 & ~n_898;
assign n_900 =  n_349 & ~n_899;
assign n_901 =  x_4935 & ~n_900;
assign n_902 = ~n_761 & ~n_901;
assign n_903 =  x_4935 & ~n_902;
assign n_904 = ~x_4935 &  n_902;
assign n_905 = ~n_903 & ~n_904;
assign n_906 =  x_4934 & ~n_900;
assign n_907 = ~n_761 & ~n_906;
assign n_908 =  x_4934 & ~n_907;
assign n_909 = ~x_4934 &  n_907;
assign n_910 = ~n_908 & ~n_909;
assign n_911 =  x_4933 & ~n_900;
assign n_912 =  x_4933 &  n_911;
assign n_913 = ~x_4933 & ~n_911;
assign n_914 = ~n_912 & ~n_913;
assign n_915 =  x_4932 & ~n_900;
assign n_916 = ~n_761 & ~n_915;
assign n_917 =  x_4932 & ~n_916;
assign n_918 = ~x_4932 &  n_916;
assign n_919 = ~n_917 & ~n_918;
assign n_920 =  x_4931 & ~n_900;
assign n_921 = ~n_761 & ~n_920;
assign n_922 =  x_4931 & ~n_921;
assign n_923 = ~x_4931 &  n_921;
assign n_924 = ~n_922 & ~n_923;
assign n_925 =  x_4930 & ~n_900;
assign n_926 = ~n_761 & ~n_925;
assign n_927 =  x_4930 & ~n_926;
assign n_928 = ~x_4930 &  n_926;
assign n_929 = ~n_927 & ~n_928;
assign n_930 =  x_4929 & ~n_900;
assign n_931 = ~n_761 & ~n_930;
assign n_932 =  x_4929 & ~n_931;
assign n_933 = ~x_4929 &  n_931;
assign n_934 = ~n_932 & ~n_933;
assign n_935 =  x_4928 & ~n_900;
assign n_936 =  x_4928 &  n_935;
assign n_937 = ~x_4928 & ~n_935;
assign n_938 = ~n_936 & ~n_937;
assign n_939 =  x_4927 & ~n_900;
assign n_940 = ~n_761 & ~n_939;
assign n_941 =  x_4927 & ~n_940;
assign n_942 = ~x_4927 &  n_940;
assign n_943 = ~n_941 & ~n_942;
assign n_944 =  x_4926 & ~n_900;
assign n_945 =  x_4926 &  n_944;
assign n_946 = ~x_4926 & ~n_944;
assign n_947 = ~n_945 & ~n_946;
assign n_948 =  x_4925 & ~n_900;
assign n_949 = ~n_761 & ~n_948;
assign n_950 =  x_4925 & ~n_949;
assign n_951 = ~x_4925 &  n_949;
assign n_952 = ~n_950 & ~n_951;
assign n_953 =  x_4924 & ~n_900;
assign n_954 =  x_4924 &  n_953;
assign n_955 = ~x_4924 & ~n_953;
assign n_956 = ~n_954 & ~n_955;
assign n_957 =  x_4923 & ~n_900;
assign n_958 =  x_4923 &  n_957;
assign n_959 = ~x_4923 & ~n_957;
assign n_960 = ~n_958 & ~n_959;
assign n_961 =  x_4922 & ~n_900;
assign n_962 =  x_4922 &  n_961;
assign n_963 = ~x_4922 & ~n_961;
assign n_964 = ~n_962 & ~n_963;
assign n_965 =  x_4921 & ~n_900;
assign n_966 =  x_4921 &  n_965;
assign n_967 = ~x_4921 & ~n_965;
assign n_968 = ~n_966 & ~n_967;
assign n_969 =  x_4920 & ~n_900;
assign n_970 =  x_4920 &  n_969;
assign n_971 = ~x_4920 & ~n_969;
assign n_972 = ~n_970 & ~n_971;
assign n_973 =  x_4919 & ~n_900;
assign n_974 =  x_4919 &  n_973;
assign n_975 = ~x_4919 & ~n_973;
assign n_976 = ~n_974 & ~n_975;
assign n_977 =  x_4918 & ~n_900;
assign n_978 =  x_4918 &  n_977;
assign n_979 = ~x_4918 & ~n_977;
assign n_980 = ~n_978 & ~n_979;
assign n_981 =  x_4917 & ~n_900;
assign n_982 =  x_4917 &  n_981;
assign n_983 = ~x_4917 & ~n_981;
assign n_984 = ~n_982 & ~n_983;
assign n_985 =  x_4916 & ~n_900;
assign n_986 =  x_4916 &  n_985;
assign n_987 = ~x_4916 & ~n_985;
assign n_988 = ~n_986 & ~n_987;
assign n_989 =  x_4915 & ~n_900;
assign n_990 =  x_4915 &  n_989;
assign n_991 = ~x_4915 & ~n_989;
assign n_992 = ~n_990 & ~n_991;
assign n_993 =  x_4914 & ~n_900;
assign n_994 =  x_4914 &  n_993;
assign n_995 = ~x_4914 & ~n_993;
assign n_996 = ~n_994 & ~n_995;
assign n_997 =  x_4913 & ~n_900;
assign n_998 =  x_4913 &  n_997;
assign n_999 = ~x_4913 & ~n_997;
assign n_1000 = ~n_998 & ~n_999;
assign n_1001 =  x_4912 & ~n_900;
assign n_1002 =  x_4912 &  n_1001;
assign n_1003 = ~x_4912 & ~n_1001;
assign n_1004 = ~n_1002 & ~n_1003;
assign n_1005 =  x_4911 & ~n_900;
assign n_1006 =  x_4911 &  n_1005;
assign n_1007 = ~x_4911 & ~n_1005;
assign n_1008 = ~n_1006 & ~n_1007;
assign n_1009 =  x_4910 & ~n_900;
assign n_1010 =  x_4910 &  n_1009;
assign n_1011 = ~x_4910 & ~n_1009;
assign n_1012 = ~n_1010 & ~n_1011;
assign n_1013 =  x_4909 & ~n_900;
assign n_1014 =  x_4909 &  n_1013;
assign n_1015 = ~x_4909 & ~n_1013;
assign n_1016 = ~n_1014 & ~n_1015;
assign n_1017 =  x_4908 & ~n_900;
assign n_1018 =  x_4908 &  n_1017;
assign n_1019 = ~x_4908 & ~n_1017;
assign n_1020 = ~n_1018 & ~n_1019;
assign n_1021 =  x_4907 & ~n_900;
assign n_1022 =  x_4907 &  n_1021;
assign n_1023 = ~x_4907 & ~n_1021;
assign n_1024 = ~n_1022 & ~n_1023;
assign n_1025 =  x_4906 & ~n_900;
assign n_1026 =  x_4906 &  n_1025;
assign n_1027 = ~x_4906 & ~n_1025;
assign n_1028 = ~n_1026 & ~n_1027;
assign n_1029 =  x_4905 & ~n_900;
assign n_1030 =  x_4905 &  n_1029;
assign n_1031 = ~x_4905 & ~n_1029;
assign n_1032 = ~n_1030 & ~n_1031;
assign n_1033 =  x_4904 & ~n_900;
assign n_1034 =  x_4904 &  n_1033;
assign n_1035 = ~x_4904 & ~n_1033;
assign n_1036 = ~n_1034 & ~n_1035;
assign n_1037 =  x_42 &  x_43;
assign n_1038 =  x_41 &  n_1037;
assign n_1039 =  x_33 & ~x_34;
assign n_1040 =  n_148 &  n_1039;
assign n_1041 =  x_39 &  n_7;
assign n_1042 =  n_1040 &  n_1041;
assign n_1043 =  x_40 &  n_1042;
assign n_1044 =  n_1038 &  n_1043;
assign n_1045 =  x_4903 & ~n_1044;
assign n_1046 =  x_4903 &  n_1045;
assign n_1047 = ~x_4903 & ~n_1045;
assign n_1048 = ~n_1046 & ~n_1047;
assign n_1049 =  x_4902 & ~n_1044;
assign n_1050 =  x_4902 &  n_1049;
assign n_1051 = ~x_4902 & ~n_1049;
assign n_1052 = ~n_1050 & ~n_1051;
assign n_1053 =  x_4901 & ~n_1044;
assign n_1054 =  x_4901 &  n_1053;
assign n_1055 = ~x_4901 & ~n_1053;
assign n_1056 = ~n_1054 & ~n_1055;
assign n_1057 =  x_4900 & ~n_1044;
assign n_1058 =  x_4900 &  n_1057;
assign n_1059 = ~x_4900 & ~n_1057;
assign n_1060 = ~n_1058 & ~n_1059;
assign n_1061 =  x_4899 & ~n_1044;
assign n_1062 =  x_4899 &  n_1061;
assign n_1063 = ~x_4899 & ~n_1061;
assign n_1064 = ~n_1062 & ~n_1063;
assign n_1065 =  x_4898 & ~n_1044;
assign n_1066 =  x_4898 &  n_1065;
assign n_1067 = ~x_4898 & ~n_1065;
assign n_1068 = ~n_1066 & ~n_1067;
assign n_1069 =  x_4897 & ~n_1044;
assign n_1070 =  x_4897 &  n_1069;
assign n_1071 = ~x_4897 & ~n_1069;
assign n_1072 = ~n_1070 & ~n_1071;
assign n_1073 =  x_4896 & ~n_1044;
assign n_1074 =  x_4896 &  n_1073;
assign n_1075 = ~x_4896 & ~n_1073;
assign n_1076 = ~n_1074 & ~n_1075;
assign n_1077 =  x_4895 & ~n_1044;
assign n_1078 =  x_4895 &  n_1077;
assign n_1079 = ~x_4895 & ~n_1077;
assign n_1080 = ~n_1078 & ~n_1079;
assign n_1081 =  x_4894 & ~n_1044;
assign n_1082 =  x_4894 &  n_1081;
assign n_1083 = ~x_4894 & ~n_1081;
assign n_1084 = ~n_1082 & ~n_1083;
assign n_1085 =  x_4893 & ~n_1044;
assign n_1086 =  x_4893 &  n_1085;
assign n_1087 = ~x_4893 & ~n_1085;
assign n_1088 = ~n_1086 & ~n_1087;
assign n_1089 =  x_4892 & ~n_1044;
assign n_1090 =  x_4892 &  n_1089;
assign n_1091 = ~x_4892 & ~n_1089;
assign n_1092 = ~n_1090 & ~n_1091;
assign n_1093 =  x_4891 & ~n_1044;
assign n_1094 =  x_4891 &  n_1093;
assign n_1095 = ~x_4891 & ~n_1093;
assign n_1096 = ~n_1094 & ~n_1095;
assign n_1097 =  x_4890 & ~n_1044;
assign n_1098 =  x_4890 &  n_1097;
assign n_1099 = ~x_4890 & ~n_1097;
assign n_1100 = ~n_1098 & ~n_1099;
assign n_1101 =  x_4889 & ~n_1044;
assign n_1102 =  x_4889 &  n_1101;
assign n_1103 = ~x_4889 & ~n_1101;
assign n_1104 = ~n_1102 & ~n_1103;
assign n_1105 =  x_4888 & ~n_1044;
assign n_1106 =  x_4888 &  n_1105;
assign n_1107 = ~x_4888 & ~n_1105;
assign n_1108 = ~n_1106 & ~n_1107;
assign n_1109 =  x_4887 & ~n_1044;
assign n_1110 =  x_4887 &  n_1109;
assign n_1111 = ~x_4887 & ~n_1109;
assign n_1112 = ~n_1110 & ~n_1111;
assign n_1113 =  x_4886 & ~n_1044;
assign n_1114 =  x_4886 &  n_1113;
assign n_1115 = ~x_4886 & ~n_1113;
assign n_1116 = ~n_1114 & ~n_1115;
assign n_1117 =  x_4885 & ~n_1044;
assign n_1118 =  x_4885 &  n_1117;
assign n_1119 = ~x_4885 & ~n_1117;
assign n_1120 = ~n_1118 & ~n_1119;
assign n_1121 =  x_4884 & ~n_1044;
assign n_1122 =  x_4884 &  n_1121;
assign n_1123 = ~x_4884 & ~n_1121;
assign n_1124 = ~n_1122 & ~n_1123;
assign n_1125 =  x_4883 & ~n_1044;
assign n_1126 =  x_4883 &  n_1125;
assign n_1127 = ~x_4883 & ~n_1125;
assign n_1128 = ~n_1126 & ~n_1127;
assign n_1129 =  x_4882 & ~n_1044;
assign n_1130 =  x_4882 &  n_1129;
assign n_1131 = ~x_4882 & ~n_1129;
assign n_1132 = ~n_1130 & ~n_1131;
assign n_1133 =  x_4881 & ~n_1044;
assign n_1134 =  x_4881 &  n_1133;
assign n_1135 = ~x_4881 & ~n_1133;
assign n_1136 = ~n_1134 & ~n_1135;
assign n_1137 =  x_4880 & ~n_1044;
assign n_1138 =  x_4880 &  n_1137;
assign n_1139 = ~x_4880 & ~n_1137;
assign n_1140 = ~n_1138 & ~n_1139;
assign n_1141 =  x_4879 & ~n_1044;
assign n_1142 =  x_4879 &  n_1141;
assign n_1143 = ~x_4879 & ~n_1141;
assign n_1144 = ~n_1142 & ~n_1143;
assign n_1145 =  x_4878 & ~n_1044;
assign n_1146 =  x_4878 &  n_1145;
assign n_1147 = ~x_4878 & ~n_1145;
assign n_1148 = ~n_1146 & ~n_1147;
assign n_1149 =  x_4877 & ~n_1044;
assign n_1150 =  x_4877 &  n_1149;
assign n_1151 = ~x_4877 & ~n_1149;
assign n_1152 = ~n_1150 & ~n_1151;
assign n_1153 =  x_4876 & ~n_1044;
assign n_1154 =  x_4876 &  n_1153;
assign n_1155 = ~x_4876 & ~n_1153;
assign n_1156 = ~n_1154 & ~n_1155;
assign n_1157 =  x_4875 & ~n_1044;
assign n_1158 =  x_4875 &  n_1157;
assign n_1159 = ~x_4875 & ~n_1157;
assign n_1160 = ~n_1158 & ~n_1159;
assign n_1161 =  x_4874 & ~n_1044;
assign n_1162 =  x_4874 &  n_1161;
assign n_1163 = ~x_4874 & ~n_1161;
assign n_1164 = ~n_1162 & ~n_1163;
assign n_1165 =  x_4873 & ~n_1044;
assign n_1166 =  x_4873 &  n_1165;
assign n_1167 = ~x_4873 & ~n_1165;
assign n_1168 = ~n_1166 & ~n_1167;
assign n_1169 =  x_4872 & ~n_1044;
assign n_1170 =  x_4872 &  n_1169;
assign n_1171 = ~x_4872 & ~n_1169;
assign n_1172 = ~n_1170 & ~n_1171;
assign n_1173 =  x_38 &  n_150;
assign n_1174 =  x_39 &  x_40;
assign n_1175 =  n_554 &  n_1174;
assign n_1176 =  n_1173 &  n_1175;
assign n_1177 =  x_4871 & ~n_1176;
assign n_1178 =  x_4871 &  n_1177;
assign n_1179 = ~x_4871 & ~n_1177;
assign n_1180 = ~n_1178 & ~n_1179;
assign n_1181 =  x_4870 & ~n_1176;
assign n_1182 =  x_4870 &  n_1181;
assign n_1183 = ~x_4870 & ~n_1181;
assign n_1184 = ~n_1182 & ~n_1183;
assign n_1185 =  x_4869 & ~n_1176;
assign n_1186 =  x_4869 &  n_1185;
assign n_1187 = ~x_4869 & ~n_1185;
assign n_1188 = ~n_1186 & ~n_1187;
assign n_1189 =  x_4868 & ~n_1176;
assign n_1190 =  x_4868 &  n_1189;
assign n_1191 = ~x_4868 & ~n_1189;
assign n_1192 = ~n_1190 & ~n_1191;
assign n_1193 =  x_4867 & ~n_1176;
assign n_1194 =  x_4867 &  n_1193;
assign n_1195 = ~x_4867 & ~n_1193;
assign n_1196 = ~n_1194 & ~n_1195;
assign n_1197 =  x_4866 & ~n_1176;
assign n_1198 =  x_4866 &  n_1197;
assign n_1199 = ~x_4866 & ~n_1197;
assign n_1200 = ~n_1198 & ~n_1199;
assign n_1201 =  x_4865 & ~n_1176;
assign n_1202 =  x_4865 &  n_1201;
assign n_1203 = ~x_4865 & ~n_1201;
assign n_1204 = ~n_1202 & ~n_1203;
assign n_1205 =  x_4864 & ~n_1176;
assign n_1206 =  x_4864 &  n_1205;
assign n_1207 = ~x_4864 & ~n_1205;
assign n_1208 = ~n_1206 & ~n_1207;
assign n_1209 =  x_4863 & ~n_1176;
assign n_1210 =  x_4863 &  n_1209;
assign n_1211 = ~x_4863 & ~n_1209;
assign n_1212 = ~n_1210 & ~n_1211;
assign n_1213 =  x_4862 & ~n_1176;
assign n_1214 =  x_4862 &  n_1213;
assign n_1215 = ~x_4862 & ~n_1213;
assign n_1216 = ~n_1214 & ~n_1215;
assign n_1217 =  x_4861 & ~n_1176;
assign n_1218 =  x_4861 &  n_1217;
assign n_1219 = ~x_4861 & ~n_1217;
assign n_1220 = ~n_1218 & ~n_1219;
assign n_1221 =  x_4860 & ~n_1176;
assign n_1222 =  x_4860 &  n_1221;
assign n_1223 = ~x_4860 & ~n_1221;
assign n_1224 = ~n_1222 & ~n_1223;
assign n_1225 =  x_4859 & ~n_1176;
assign n_1226 =  x_4859 &  n_1225;
assign n_1227 = ~x_4859 & ~n_1225;
assign n_1228 = ~n_1226 & ~n_1227;
assign n_1229 =  x_4858 & ~n_1176;
assign n_1230 =  x_4858 &  n_1229;
assign n_1231 = ~x_4858 & ~n_1229;
assign n_1232 = ~n_1230 & ~n_1231;
assign n_1233 =  x_4857 & ~n_1176;
assign n_1234 =  x_4857 &  n_1233;
assign n_1235 = ~x_4857 & ~n_1233;
assign n_1236 = ~n_1234 & ~n_1235;
assign n_1237 =  x_4856 & ~n_1176;
assign n_1238 =  x_4856 &  n_1237;
assign n_1239 = ~x_4856 & ~n_1237;
assign n_1240 = ~n_1238 & ~n_1239;
assign n_1241 =  x_4855 & ~n_1176;
assign n_1242 =  x_4855 &  n_1241;
assign n_1243 = ~x_4855 & ~n_1241;
assign n_1244 = ~n_1242 & ~n_1243;
assign n_1245 =  x_4854 & ~n_1176;
assign n_1246 =  x_4854 &  n_1245;
assign n_1247 = ~x_4854 & ~n_1245;
assign n_1248 = ~n_1246 & ~n_1247;
assign n_1249 =  x_4853 & ~n_1176;
assign n_1250 =  x_4853 &  n_1249;
assign n_1251 = ~x_4853 & ~n_1249;
assign n_1252 = ~n_1250 & ~n_1251;
assign n_1253 =  x_4852 & ~n_1176;
assign n_1254 =  x_4852 &  n_1253;
assign n_1255 = ~x_4852 & ~n_1253;
assign n_1256 = ~n_1254 & ~n_1255;
assign n_1257 =  x_4851 & ~n_1176;
assign n_1258 =  x_4851 &  n_1257;
assign n_1259 = ~x_4851 & ~n_1257;
assign n_1260 = ~n_1258 & ~n_1259;
assign n_1261 =  x_4850 & ~n_1176;
assign n_1262 =  x_4850 &  n_1261;
assign n_1263 = ~x_4850 & ~n_1261;
assign n_1264 = ~n_1262 & ~n_1263;
assign n_1265 =  x_4849 & ~n_1176;
assign n_1266 =  x_4849 &  n_1265;
assign n_1267 = ~x_4849 & ~n_1265;
assign n_1268 = ~n_1266 & ~n_1267;
assign n_1269 =  x_4848 & ~n_1176;
assign n_1270 =  x_4848 &  n_1269;
assign n_1271 = ~x_4848 & ~n_1269;
assign n_1272 = ~n_1270 & ~n_1271;
assign n_1273 =  x_4847 & ~n_1176;
assign n_1274 =  x_4847 &  n_1273;
assign n_1275 = ~x_4847 & ~n_1273;
assign n_1276 = ~n_1274 & ~n_1275;
assign n_1277 =  x_4846 & ~n_1176;
assign n_1278 =  x_4846 &  n_1277;
assign n_1279 = ~x_4846 & ~n_1277;
assign n_1280 = ~n_1278 & ~n_1279;
assign n_1281 =  x_4845 & ~n_1176;
assign n_1282 =  x_4845 &  n_1281;
assign n_1283 = ~x_4845 & ~n_1281;
assign n_1284 = ~n_1282 & ~n_1283;
assign n_1285 =  x_4844 & ~n_1176;
assign n_1286 =  x_4844 &  n_1285;
assign n_1287 = ~x_4844 & ~n_1285;
assign n_1288 = ~n_1286 & ~n_1287;
assign n_1289 =  x_4843 & ~n_1176;
assign n_1290 =  x_4843 &  n_1289;
assign n_1291 = ~x_4843 & ~n_1289;
assign n_1292 = ~n_1290 & ~n_1291;
assign n_1293 =  x_4842 & ~n_1176;
assign n_1294 =  x_4842 &  n_1293;
assign n_1295 = ~x_4842 & ~n_1293;
assign n_1296 = ~n_1294 & ~n_1295;
assign n_1297 =  x_4841 & ~n_1176;
assign n_1298 =  x_4841 &  n_1297;
assign n_1299 = ~x_4841 & ~n_1297;
assign n_1300 = ~n_1298 & ~n_1299;
assign n_1301 =  x_4840 & ~n_1176;
assign n_1302 =  x_4840 &  n_1301;
assign n_1303 = ~x_4840 & ~n_1301;
assign n_1304 = ~n_1302 & ~n_1303;
assign n_1305 = ~x_39 &  x_40;
assign n_1306 =  n_7 &  n_765;
assign n_1307 =  n_1305 &  n_1306;
assign n_1308 =  n_1038 &  n_1307;
assign n_1309 =  x_4839 & ~n_1308;
assign n_1310 =  x_2058 &  n_1308;
assign n_1311 = ~n_1309 & ~n_1310;
assign n_1312 =  x_4839 & ~n_1311;
assign n_1313 = ~x_4839 &  n_1311;
assign n_1314 = ~n_1312 & ~n_1313;
assign n_1315 =  x_4838 & ~n_1308;
assign n_1316 =  x_2057 &  n_1308;
assign n_1317 = ~n_1315 & ~n_1316;
assign n_1318 =  x_4838 & ~n_1317;
assign n_1319 = ~x_4838 &  n_1317;
assign n_1320 = ~n_1318 & ~n_1319;
assign n_1321 =  x_4837 & ~n_1308;
assign n_1322 =  x_2056 &  n_1308;
assign n_1323 = ~n_1321 & ~n_1322;
assign n_1324 =  x_4837 & ~n_1323;
assign n_1325 = ~x_4837 &  n_1323;
assign n_1326 = ~n_1324 & ~n_1325;
assign n_1327 =  x_4836 & ~n_1308;
assign n_1328 =  x_2055 &  n_1308;
assign n_1329 = ~n_1327 & ~n_1328;
assign n_1330 =  x_4836 & ~n_1329;
assign n_1331 = ~x_4836 &  n_1329;
assign n_1332 = ~n_1330 & ~n_1331;
assign n_1333 =  x_4835 & ~n_1308;
assign n_1334 =  x_2054 &  n_1308;
assign n_1335 = ~n_1333 & ~n_1334;
assign n_1336 =  x_4835 & ~n_1335;
assign n_1337 = ~x_4835 &  n_1335;
assign n_1338 = ~n_1336 & ~n_1337;
assign n_1339 =  x_4834 & ~n_1308;
assign n_1340 =  x_2053 &  n_1308;
assign n_1341 = ~n_1339 & ~n_1340;
assign n_1342 =  x_4834 & ~n_1341;
assign n_1343 = ~x_4834 &  n_1341;
assign n_1344 = ~n_1342 & ~n_1343;
assign n_1345 =  x_4833 & ~n_1308;
assign n_1346 =  x_2052 &  n_1308;
assign n_1347 = ~n_1345 & ~n_1346;
assign n_1348 =  x_4833 & ~n_1347;
assign n_1349 = ~x_4833 &  n_1347;
assign n_1350 = ~n_1348 & ~n_1349;
assign n_1351 =  x_4832 & ~n_1308;
assign n_1352 =  x_2051 &  n_1308;
assign n_1353 = ~n_1351 & ~n_1352;
assign n_1354 =  x_4832 & ~n_1353;
assign n_1355 = ~x_4832 &  n_1353;
assign n_1356 = ~n_1354 & ~n_1355;
assign n_1357 =  x_4831 & ~n_1308;
assign n_1358 =  x_2050 &  n_1308;
assign n_1359 = ~n_1357 & ~n_1358;
assign n_1360 =  x_4831 & ~n_1359;
assign n_1361 = ~x_4831 &  n_1359;
assign n_1362 = ~n_1360 & ~n_1361;
assign n_1363 =  x_4830 & ~n_1308;
assign n_1364 =  x_2049 &  n_1308;
assign n_1365 = ~n_1363 & ~n_1364;
assign n_1366 =  x_4830 & ~n_1365;
assign n_1367 = ~x_4830 &  n_1365;
assign n_1368 = ~n_1366 & ~n_1367;
assign n_1369 =  x_4829 & ~n_1308;
assign n_1370 =  x_2048 &  n_1308;
assign n_1371 = ~n_1369 & ~n_1370;
assign n_1372 =  x_4829 & ~n_1371;
assign n_1373 = ~x_4829 &  n_1371;
assign n_1374 = ~n_1372 & ~n_1373;
assign n_1375 =  x_4828 & ~n_1308;
assign n_1376 =  x_2047 &  n_1308;
assign n_1377 = ~n_1375 & ~n_1376;
assign n_1378 =  x_4828 & ~n_1377;
assign n_1379 = ~x_4828 &  n_1377;
assign n_1380 = ~n_1378 & ~n_1379;
assign n_1381 =  x_4827 & ~n_1308;
assign n_1382 =  x_2046 &  n_1308;
assign n_1383 = ~n_1381 & ~n_1382;
assign n_1384 =  x_4827 & ~n_1383;
assign n_1385 = ~x_4827 &  n_1383;
assign n_1386 = ~n_1384 & ~n_1385;
assign n_1387 =  x_4826 & ~n_1308;
assign n_1388 =  x_2045 &  n_1308;
assign n_1389 = ~n_1387 & ~n_1388;
assign n_1390 =  x_4826 & ~n_1389;
assign n_1391 = ~x_4826 &  n_1389;
assign n_1392 = ~n_1390 & ~n_1391;
assign n_1393 =  x_4825 & ~n_1308;
assign n_1394 =  x_2044 &  n_1308;
assign n_1395 = ~n_1393 & ~n_1394;
assign n_1396 =  x_4825 & ~n_1395;
assign n_1397 = ~x_4825 &  n_1395;
assign n_1398 = ~n_1396 & ~n_1397;
assign n_1399 =  x_4824 & ~n_1308;
assign n_1400 =  x_2043 &  n_1308;
assign n_1401 = ~n_1399 & ~n_1400;
assign n_1402 =  x_4824 & ~n_1401;
assign n_1403 = ~x_4824 &  n_1401;
assign n_1404 = ~n_1402 & ~n_1403;
assign n_1405 =  x_4823 & ~n_1308;
assign n_1406 =  x_2042 &  n_1308;
assign n_1407 = ~n_1405 & ~n_1406;
assign n_1408 =  x_4823 & ~n_1407;
assign n_1409 = ~x_4823 &  n_1407;
assign n_1410 = ~n_1408 & ~n_1409;
assign n_1411 =  x_4822 & ~n_1308;
assign n_1412 =  x_2041 &  n_1308;
assign n_1413 = ~n_1411 & ~n_1412;
assign n_1414 =  x_4822 & ~n_1413;
assign n_1415 = ~x_4822 &  n_1413;
assign n_1416 = ~n_1414 & ~n_1415;
assign n_1417 =  x_4821 & ~n_1308;
assign n_1418 =  x_2040 &  n_1308;
assign n_1419 = ~n_1417 & ~n_1418;
assign n_1420 =  x_4821 & ~n_1419;
assign n_1421 = ~x_4821 &  n_1419;
assign n_1422 = ~n_1420 & ~n_1421;
assign n_1423 =  x_4820 & ~n_1308;
assign n_1424 =  x_2039 &  n_1308;
assign n_1425 = ~n_1423 & ~n_1424;
assign n_1426 =  x_4820 & ~n_1425;
assign n_1427 = ~x_4820 &  n_1425;
assign n_1428 = ~n_1426 & ~n_1427;
assign n_1429 =  x_4819 & ~n_1308;
assign n_1430 =  x_2038 &  n_1308;
assign n_1431 = ~n_1429 & ~n_1430;
assign n_1432 =  x_4819 & ~n_1431;
assign n_1433 = ~x_4819 &  n_1431;
assign n_1434 = ~n_1432 & ~n_1433;
assign n_1435 =  x_4818 & ~n_1308;
assign n_1436 =  x_2037 &  n_1308;
assign n_1437 = ~n_1435 & ~n_1436;
assign n_1438 =  x_4818 & ~n_1437;
assign n_1439 = ~x_4818 &  n_1437;
assign n_1440 = ~n_1438 & ~n_1439;
assign n_1441 =  x_4817 & ~n_1308;
assign n_1442 =  x_2036 &  n_1308;
assign n_1443 = ~n_1441 & ~n_1442;
assign n_1444 =  x_4817 & ~n_1443;
assign n_1445 = ~x_4817 &  n_1443;
assign n_1446 = ~n_1444 & ~n_1445;
assign n_1447 =  x_4816 & ~n_1308;
assign n_1448 =  x_2035 &  n_1308;
assign n_1449 = ~n_1447 & ~n_1448;
assign n_1450 =  x_4816 & ~n_1449;
assign n_1451 = ~x_4816 &  n_1449;
assign n_1452 = ~n_1450 & ~n_1451;
assign n_1453 =  x_4815 & ~n_1308;
assign n_1454 =  x_2034 &  n_1308;
assign n_1455 = ~n_1453 & ~n_1454;
assign n_1456 =  x_4815 & ~n_1455;
assign n_1457 = ~x_4815 &  n_1455;
assign n_1458 = ~n_1456 & ~n_1457;
assign n_1459 =  x_4814 & ~n_1308;
assign n_1460 =  x_2033 &  n_1308;
assign n_1461 = ~n_1459 & ~n_1460;
assign n_1462 =  x_4814 & ~n_1461;
assign n_1463 = ~x_4814 &  n_1461;
assign n_1464 = ~n_1462 & ~n_1463;
assign n_1465 =  x_4813 & ~n_1308;
assign n_1466 =  x_2032 &  n_1308;
assign n_1467 = ~n_1465 & ~n_1466;
assign n_1468 =  x_4813 & ~n_1467;
assign n_1469 = ~x_4813 &  n_1467;
assign n_1470 = ~n_1468 & ~n_1469;
assign n_1471 =  x_4812 & ~n_1308;
assign n_1472 =  x_2031 &  n_1308;
assign n_1473 = ~n_1471 & ~n_1472;
assign n_1474 =  x_4812 & ~n_1473;
assign n_1475 = ~x_4812 &  n_1473;
assign n_1476 = ~n_1474 & ~n_1475;
assign n_1477 =  x_4811 & ~n_1308;
assign n_1478 =  x_2030 &  n_1308;
assign n_1479 = ~n_1477 & ~n_1478;
assign n_1480 =  x_4811 & ~n_1479;
assign n_1481 = ~x_4811 &  n_1479;
assign n_1482 = ~n_1480 & ~n_1481;
assign n_1483 =  x_4810 & ~n_1308;
assign n_1484 =  x_2029 &  n_1308;
assign n_1485 = ~n_1483 & ~n_1484;
assign n_1486 =  x_4810 & ~n_1485;
assign n_1487 = ~x_4810 &  n_1485;
assign n_1488 = ~n_1486 & ~n_1487;
assign n_1489 =  x_4809 & ~n_1308;
assign n_1490 =  x_2028 &  n_1308;
assign n_1491 = ~n_1489 & ~n_1490;
assign n_1492 =  x_4809 & ~n_1491;
assign n_1493 = ~x_4809 &  n_1491;
assign n_1494 = ~n_1492 & ~n_1493;
assign n_1495 =  x_4808 & ~n_1308;
assign n_1496 =  x_2027 &  n_1308;
assign n_1497 = ~n_1495 & ~n_1496;
assign n_1498 =  x_4808 & ~n_1497;
assign n_1499 = ~x_4808 &  n_1497;
assign n_1500 = ~n_1498 & ~n_1499;
assign n_1501 = ~x_37 &  n_764;
assign n_1502 =  n_352 &  n_1501;
assign n_1503 = ~x_38 &  n_1502;
assign n_1504 =  n_6 &  n_1503;
assign n_1505 =  n_758 &  n_1504;
assign n_1506 =  x_4807 & ~n_1505;
assign n_1507 =  x_2058 &  n_1505;
assign n_1508 = ~n_1506 & ~n_1507;
assign n_1509 =  x_4807 & ~n_1508;
assign n_1510 = ~x_4807 &  n_1508;
assign n_1511 = ~n_1509 & ~n_1510;
assign n_1512 =  x_4806 & ~n_1505;
assign n_1513 =  x_2057 &  n_1505;
assign n_1514 = ~n_1512 & ~n_1513;
assign n_1515 =  x_4806 & ~n_1514;
assign n_1516 = ~x_4806 &  n_1514;
assign n_1517 = ~n_1515 & ~n_1516;
assign n_1518 =  x_4805 & ~n_1505;
assign n_1519 =  x_2056 &  n_1505;
assign n_1520 = ~n_1518 & ~n_1519;
assign n_1521 =  x_4805 & ~n_1520;
assign n_1522 = ~x_4805 &  n_1520;
assign n_1523 = ~n_1521 & ~n_1522;
assign n_1524 =  x_4804 & ~n_1505;
assign n_1525 =  x_2055 &  n_1505;
assign n_1526 = ~n_1524 & ~n_1525;
assign n_1527 =  x_4804 & ~n_1526;
assign n_1528 = ~x_4804 &  n_1526;
assign n_1529 = ~n_1527 & ~n_1528;
assign n_1530 =  x_4803 & ~n_1505;
assign n_1531 =  x_2054 &  n_1505;
assign n_1532 = ~n_1530 & ~n_1531;
assign n_1533 =  x_4803 & ~n_1532;
assign n_1534 = ~x_4803 &  n_1532;
assign n_1535 = ~n_1533 & ~n_1534;
assign n_1536 =  x_4802 & ~n_1505;
assign n_1537 =  x_2053 &  n_1505;
assign n_1538 = ~n_1536 & ~n_1537;
assign n_1539 =  x_4802 & ~n_1538;
assign n_1540 = ~x_4802 &  n_1538;
assign n_1541 = ~n_1539 & ~n_1540;
assign n_1542 =  x_4801 & ~n_1505;
assign n_1543 =  x_2052 &  n_1505;
assign n_1544 = ~n_1542 & ~n_1543;
assign n_1545 =  x_4801 & ~n_1544;
assign n_1546 = ~x_4801 &  n_1544;
assign n_1547 = ~n_1545 & ~n_1546;
assign n_1548 =  x_4800 & ~n_1505;
assign n_1549 =  x_2051 &  n_1505;
assign n_1550 = ~n_1548 & ~n_1549;
assign n_1551 =  x_4800 & ~n_1550;
assign n_1552 = ~x_4800 &  n_1550;
assign n_1553 = ~n_1551 & ~n_1552;
assign n_1554 =  x_4799 & ~n_1505;
assign n_1555 =  x_2050 &  n_1505;
assign n_1556 = ~n_1554 & ~n_1555;
assign n_1557 =  x_4799 & ~n_1556;
assign n_1558 = ~x_4799 &  n_1556;
assign n_1559 = ~n_1557 & ~n_1558;
assign n_1560 =  x_4798 & ~n_1505;
assign n_1561 =  x_2049 &  n_1505;
assign n_1562 = ~n_1560 & ~n_1561;
assign n_1563 =  x_4798 & ~n_1562;
assign n_1564 = ~x_4798 &  n_1562;
assign n_1565 = ~n_1563 & ~n_1564;
assign n_1566 =  x_4797 & ~n_1505;
assign n_1567 =  x_2048 &  n_1505;
assign n_1568 = ~n_1566 & ~n_1567;
assign n_1569 =  x_4797 & ~n_1568;
assign n_1570 = ~x_4797 &  n_1568;
assign n_1571 = ~n_1569 & ~n_1570;
assign n_1572 =  x_4796 & ~n_1505;
assign n_1573 =  x_2047 &  n_1505;
assign n_1574 = ~n_1572 & ~n_1573;
assign n_1575 =  x_4796 & ~n_1574;
assign n_1576 = ~x_4796 &  n_1574;
assign n_1577 = ~n_1575 & ~n_1576;
assign n_1578 =  x_4795 & ~n_1505;
assign n_1579 =  x_2046 &  n_1505;
assign n_1580 = ~n_1578 & ~n_1579;
assign n_1581 =  x_4795 & ~n_1580;
assign n_1582 = ~x_4795 &  n_1580;
assign n_1583 = ~n_1581 & ~n_1582;
assign n_1584 =  x_4794 & ~n_1505;
assign n_1585 =  x_2045 &  n_1505;
assign n_1586 = ~n_1584 & ~n_1585;
assign n_1587 =  x_4794 & ~n_1586;
assign n_1588 = ~x_4794 &  n_1586;
assign n_1589 = ~n_1587 & ~n_1588;
assign n_1590 =  x_4793 & ~n_1505;
assign n_1591 =  x_2044 &  n_1505;
assign n_1592 = ~n_1590 & ~n_1591;
assign n_1593 =  x_4793 & ~n_1592;
assign n_1594 = ~x_4793 &  n_1592;
assign n_1595 = ~n_1593 & ~n_1594;
assign n_1596 =  x_4792 & ~n_1505;
assign n_1597 =  x_2043 &  n_1505;
assign n_1598 = ~n_1596 & ~n_1597;
assign n_1599 =  x_4792 & ~n_1598;
assign n_1600 = ~x_4792 &  n_1598;
assign n_1601 = ~n_1599 & ~n_1600;
assign n_1602 =  x_4791 & ~n_1505;
assign n_1603 =  x_2042 &  n_1505;
assign n_1604 = ~n_1602 & ~n_1603;
assign n_1605 =  x_4791 & ~n_1604;
assign n_1606 = ~x_4791 &  n_1604;
assign n_1607 = ~n_1605 & ~n_1606;
assign n_1608 =  x_4790 & ~n_1505;
assign n_1609 =  x_2041 &  n_1505;
assign n_1610 = ~n_1608 & ~n_1609;
assign n_1611 =  x_4790 & ~n_1610;
assign n_1612 = ~x_4790 &  n_1610;
assign n_1613 = ~n_1611 & ~n_1612;
assign n_1614 =  x_4789 & ~n_1505;
assign n_1615 =  x_2040 &  n_1505;
assign n_1616 = ~n_1614 & ~n_1615;
assign n_1617 =  x_4789 & ~n_1616;
assign n_1618 = ~x_4789 &  n_1616;
assign n_1619 = ~n_1617 & ~n_1618;
assign n_1620 =  x_4788 & ~n_1505;
assign n_1621 =  x_2039 &  n_1505;
assign n_1622 = ~n_1620 & ~n_1621;
assign n_1623 =  x_4788 & ~n_1622;
assign n_1624 = ~x_4788 &  n_1622;
assign n_1625 = ~n_1623 & ~n_1624;
assign n_1626 =  x_4787 & ~n_1505;
assign n_1627 =  x_2038 &  n_1505;
assign n_1628 = ~n_1626 & ~n_1627;
assign n_1629 =  x_4787 & ~n_1628;
assign n_1630 = ~x_4787 &  n_1628;
assign n_1631 = ~n_1629 & ~n_1630;
assign n_1632 =  x_4786 & ~n_1505;
assign n_1633 =  x_2037 &  n_1505;
assign n_1634 = ~n_1632 & ~n_1633;
assign n_1635 =  x_4786 & ~n_1634;
assign n_1636 = ~x_4786 &  n_1634;
assign n_1637 = ~n_1635 & ~n_1636;
assign n_1638 =  x_4785 & ~n_1505;
assign n_1639 =  x_2036 &  n_1505;
assign n_1640 = ~n_1638 & ~n_1639;
assign n_1641 =  x_4785 & ~n_1640;
assign n_1642 = ~x_4785 &  n_1640;
assign n_1643 = ~n_1641 & ~n_1642;
assign n_1644 =  x_4784 & ~n_1505;
assign n_1645 =  x_2035 &  n_1505;
assign n_1646 = ~n_1644 & ~n_1645;
assign n_1647 =  x_4784 & ~n_1646;
assign n_1648 = ~x_4784 &  n_1646;
assign n_1649 = ~n_1647 & ~n_1648;
assign n_1650 =  x_4783 & ~n_1505;
assign n_1651 =  x_2034 &  n_1505;
assign n_1652 = ~n_1650 & ~n_1651;
assign n_1653 =  x_4783 & ~n_1652;
assign n_1654 = ~x_4783 &  n_1652;
assign n_1655 = ~n_1653 & ~n_1654;
assign n_1656 =  x_4782 & ~n_1505;
assign n_1657 =  x_2033 &  n_1505;
assign n_1658 = ~n_1656 & ~n_1657;
assign n_1659 =  x_4782 & ~n_1658;
assign n_1660 = ~x_4782 &  n_1658;
assign n_1661 = ~n_1659 & ~n_1660;
assign n_1662 =  x_4781 & ~n_1505;
assign n_1663 =  x_2032 &  n_1505;
assign n_1664 = ~n_1662 & ~n_1663;
assign n_1665 =  x_4781 & ~n_1664;
assign n_1666 = ~x_4781 &  n_1664;
assign n_1667 = ~n_1665 & ~n_1666;
assign n_1668 =  x_4780 & ~n_1505;
assign n_1669 =  x_2031 &  n_1505;
assign n_1670 = ~n_1668 & ~n_1669;
assign n_1671 =  x_4780 & ~n_1670;
assign n_1672 = ~x_4780 &  n_1670;
assign n_1673 = ~n_1671 & ~n_1672;
assign n_1674 =  x_4779 & ~n_1505;
assign n_1675 =  x_2030 &  n_1505;
assign n_1676 = ~n_1674 & ~n_1675;
assign n_1677 =  x_4779 & ~n_1676;
assign n_1678 = ~x_4779 &  n_1676;
assign n_1679 = ~n_1677 & ~n_1678;
assign n_1680 =  x_4778 & ~n_1505;
assign n_1681 =  x_2029 &  n_1505;
assign n_1682 = ~n_1680 & ~n_1681;
assign n_1683 =  x_4778 & ~n_1682;
assign n_1684 = ~x_4778 &  n_1682;
assign n_1685 = ~n_1683 & ~n_1684;
assign n_1686 =  x_4777 & ~n_1505;
assign n_1687 =  x_2028 &  n_1505;
assign n_1688 = ~n_1686 & ~n_1687;
assign n_1689 =  x_4777 & ~n_1688;
assign n_1690 = ~x_4777 &  n_1688;
assign n_1691 = ~n_1689 & ~n_1690;
assign n_1692 =  x_4776 & ~n_1505;
assign n_1693 =  x_2027 &  n_1505;
assign n_1694 = ~n_1692 & ~n_1693;
assign n_1695 =  x_4776 & ~n_1694;
assign n_1696 = ~x_4776 &  n_1694;
assign n_1697 = ~n_1695 & ~n_1696;
assign n_1698 =  x_38 &  n_355;
assign n_1699 =  n_759 &  n_1698;
assign n_1700 =  n_152 &  n_1699;
assign n_1701 =  x_43 &  n_1700;
assign n_1702 =  x_4775 & ~n_1701;
assign n_1703 =  x_1610 &  n_1701;
assign n_1704 = ~n_1702 & ~n_1703;
assign n_1705 =  x_4775 & ~n_1704;
assign n_1706 = ~x_4775 &  n_1704;
assign n_1707 = ~n_1705 & ~n_1706;
assign n_1708 =  x_4774 & ~n_1701;
assign n_1709 =  x_1609 &  n_1701;
assign n_1710 = ~n_1708 & ~n_1709;
assign n_1711 =  x_4774 & ~n_1710;
assign n_1712 = ~x_4774 &  n_1710;
assign n_1713 = ~n_1711 & ~n_1712;
assign n_1714 =  x_4773 & ~n_1701;
assign n_1715 =  x_1608 &  n_1701;
assign n_1716 = ~n_1714 & ~n_1715;
assign n_1717 =  x_4773 & ~n_1716;
assign n_1718 = ~x_4773 &  n_1716;
assign n_1719 = ~n_1717 & ~n_1718;
assign n_1720 =  x_4772 & ~n_1701;
assign n_1721 =  x_1607 &  n_1701;
assign n_1722 = ~n_1720 & ~n_1721;
assign n_1723 =  x_4772 & ~n_1722;
assign n_1724 = ~x_4772 &  n_1722;
assign n_1725 = ~n_1723 & ~n_1724;
assign n_1726 =  x_4771 & ~n_1701;
assign n_1727 =  x_1606 &  n_1701;
assign n_1728 = ~n_1726 & ~n_1727;
assign n_1729 =  x_4771 & ~n_1728;
assign n_1730 = ~x_4771 &  n_1728;
assign n_1731 = ~n_1729 & ~n_1730;
assign n_1732 =  x_4770 & ~n_1701;
assign n_1733 =  x_1605 &  n_1701;
assign n_1734 = ~n_1732 & ~n_1733;
assign n_1735 =  x_4770 & ~n_1734;
assign n_1736 = ~x_4770 &  n_1734;
assign n_1737 = ~n_1735 & ~n_1736;
assign n_1738 =  x_4769 & ~n_1701;
assign n_1739 =  x_1604 &  n_1701;
assign n_1740 = ~n_1738 & ~n_1739;
assign n_1741 =  x_4769 & ~n_1740;
assign n_1742 = ~x_4769 &  n_1740;
assign n_1743 = ~n_1741 & ~n_1742;
assign n_1744 =  x_4768 & ~n_1701;
assign n_1745 =  x_1603 &  n_1701;
assign n_1746 = ~n_1744 & ~n_1745;
assign n_1747 =  x_4768 & ~n_1746;
assign n_1748 = ~x_4768 &  n_1746;
assign n_1749 = ~n_1747 & ~n_1748;
assign n_1750 =  x_4767 & ~n_1701;
assign n_1751 =  x_1602 &  n_1701;
assign n_1752 = ~n_1750 & ~n_1751;
assign n_1753 =  x_4767 & ~n_1752;
assign n_1754 = ~x_4767 &  n_1752;
assign n_1755 = ~n_1753 & ~n_1754;
assign n_1756 =  x_4766 & ~n_1701;
assign n_1757 =  x_1601 &  n_1701;
assign n_1758 = ~n_1756 & ~n_1757;
assign n_1759 =  x_4766 & ~n_1758;
assign n_1760 = ~x_4766 &  n_1758;
assign n_1761 = ~n_1759 & ~n_1760;
assign n_1762 =  x_4765 & ~n_1701;
assign n_1763 =  x_1600 &  n_1701;
assign n_1764 = ~n_1762 & ~n_1763;
assign n_1765 =  x_4765 & ~n_1764;
assign n_1766 = ~x_4765 &  n_1764;
assign n_1767 = ~n_1765 & ~n_1766;
assign n_1768 =  x_4764 & ~n_1701;
assign n_1769 =  x_1599 &  n_1701;
assign n_1770 = ~n_1768 & ~n_1769;
assign n_1771 =  x_4764 & ~n_1770;
assign n_1772 = ~x_4764 &  n_1770;
assign n_1773 = ~n_1771 & ~n_1772;
assign n_1774 =  x_4763 & ~n_1701;
assign n_1775 =  x_1598 &  n_1701;
assign n_1776 = ~n_1774 & ~n_1775;
assign n_1777 =  x_4763 & ~n_1776;
assign n_1778 = ~x_4763 &  n_1776;
assign n_1779 = ~n_1777 & ~n_1778;
assign n_1780 =  x_4762 & ~n_1701;
assign n_1781 =  x_1597 &  n_1701;
assign n_1782 = ~n_1780 & ~n_1781;
assign n_1783 =  x_4762 & ~n_1782;
assign n_1784 = ~x_4762 &  n_1782;
assign n_1785 = ~n_1783 & ~n_1784;
assign n_1786 =  x_4761 & ~n_1701;
assign n_1787 =  x_1596 &  n_1701;
assign n_1788 = ~n_1786 & ~n_1787;
assign n_1789 =  x_4761 & ~n_1788;
assign n_1790 = ~x_4761 &  n_1788;
assign n_1791 = ~n_1789 & ~n_1790;
assign n_1792 =  x_4760 & ~n_1701;
assign n_1793 =  x_1595 &  n_1701;
assign n_1794 = ~n_1792 & ~n_1793;
assign n_1795 =  x_4760 & ~n_1794;
assign n_1796 = ~x_4760 &  n_1794;
assign n_1797 = ~n_1795 & ~n_1796;
assign n_1798 =  x_4759 & ~n_1701;
assign n_1799 =  x_1594 &  n_1701;
assign n_1800 = ~n_1798 & ~n_1799;
assign n_1801 =  x_4759 & ~n_1800;
assign n_1802 = ~x_4759 &  n_1800;
assign n_1803 = ~n_1801 & ~n_1802;
assign n_1804 =  x_4758 & ~n_1701;
assign n_1805 =  x_1593 &  n_1701;
assign n_1806 = ~n_1804 & ~n_1805;
assign n_1807 =  x_4758 & ~n_1806;
assign n_1808 = ~x_4758 &  n_1806;
assign n_1809 = ~n_1807 & ~n_1808;
assign n_1810 =  x_4757 & ~n_1701;
assign n_1811 =  x_1592 &  n_1701;
assign n_1812 = ~n_1810 & ~n_1811;
assign n_1813 =  x_4757 & ~n_1812;
assign n_1814 = ~x_4757 &  n_1812;
assign n_1815 = ~n_1813 & ~n_1814;
assign n_1816 =  x_4756 & ~n_1701;
assign n_1817 =  x_1591 &  n_1701;
assign n_1818 = ~n_1816 & ~n_1817;
assign n_1819 =  x_4756 & ~n_1818;
assign n_1820 = ~x_4756 &  n_1818;
assign n_1821 = ~n_1819 & ~n_1820;
assign n_1822 =  x_4755 & ~n_1701;
assign n_1823 =  x_1590 &  n_1701;
assign n_1824 = ~n_1822 & ~n_1823;
assign n_1825 =  x_4755 & ~n_1824;
assign n_1826 = ~x_4755 &  n_1824;
assign n_1827 = ~n_1825 & ~n_1826;
assign n_1828 =  x_4754 & ~n_1701;
assign n_1829 =  x_1589 &  n_1701;
assign n_1830 = ~n_1828 & ~n_1829;
assign n_1831 =  x_4754 & ~n_1830;
assign n_1832 = ~x_4754 &  n_1830;
assign n_1833 = ~n_1831 & ~n_1832;
assign n_1834 =  x_4753 & ~n_1701;
assign n_1835 =  x_1588 &  n_1701;
assign n_1836 = ~n_1834 & ~n_1835;
assign n_1837 =  x_4753 & ~n_1836;
assign n_1838 = ~x_4753 &  n_1836;
assign n_1839 = ~n_1837 & ~n_1838;
assign n_1840 =  x_4752 & ~n_1701;
assign n_1841 =  x_1587 &  n_1701;
assign n_1842 = ~n_1840 & ~n_1841;
assign n_1843 =  x_4752 & ~n_1842;
assign n_1844 = ~x_4752 &  n_1842;
assign n_1845 = ~n_1843 & ~n_1844;
assign n_1846 =  x_4751 & ~n_1701;
assign n_1847 =  x_1586 &  n_1701;
assign n_1848 = ~n_1846 & ~n_1847;
assign n_1849 =  x_4751 & ~n_1848;
assign n_1850 = ~x_4751 &  n_1848;
assign n_1851 = ~n_1849 & ~n_1850;
assign n_1852 =  x_4750 & ~n_1701;
assign n_1853 =  x_1585 &  n_1701;
assign n_1854 = ~n_1852 & ~n_1853;
assign n_1855 =  x_4750 & ~n_1854;
assign n_1856 = ~x_4750 &  n_1854;
assign n_1857 = ~n_1855 & ~n_1856;
assign n_1858 =  x_4749 & ~n_1701;
assign n_1859 =  x_1584 &  n_1701;
assign n_1860 = ~n_1858 & ~n_1859;
assign n_1861 =  x_4749 & ~n_1860;
assign n_1862 = ~x_4749 &  n_1860;
assign n_1863 = ~n_1861 & ~n_1862;
assign n_1864 =  x_4748 & ~n_1701;
assign n_1865 =  x_1583 &  n_1701;
assign n_1866 = ~n_1864 & ~n_1865;
assign n_1867 =  x_4748 & ~n_1866;
assign n_1868 = ~x_4748 &  n_1866;
assign n_1869 = ~n_1867 & ~n_1868;
assign n_1870 =  x_4747 & ~n_1701;
assign n_1871 =  x_1582 &  n_1701;
assign n_1872 = ~n_1870 & ~n_1871;
assign n_1873 =  x_4747 & ~n_1872;
assign n_1874 = ~x_4747 &  n_1872;
assign n_1875 = ~n_1873 & ~n_1874;
assign n_1876 =  x_4746 & ~n_1701;
assign n_1877 =  x_1581 &  n_1701;
assign n_1878 = ~n_1876 & ~n_1877;
assign n_1879 =  x_4746 & ~n_1878;
assign n_1880 = ~x_4746 &  n_1878;
assign n_1881 = ~n_1879 & ~n_1880;
assign n_1882 =  x_4745 & ~n_1701;
assign n_1883 =  x_1580 &  n_1701;
assign n_1884 = ~n_1882 & ~n_1883;
assign n_1885 =  x_4745 & ~n_1884;
assign n_1886 = ~x_4745 &  n_1884;
assign n_1887 = ~n_1885 & ~n_1886;
assign n_1888 =  x_4744 & ~n_1701;
assign n_1889 =  x_1579 &  n_1701;
assign n_1890 = ~n_1888 & ~n_1889;
assign n_1891 =  x_4744 & ~n_1890;
assign n_1892 = ~x_4744 &  n_1890;
assign n_1893 = ~n_1891 & ~n_1892;
assign n_1894 = ~x_43 &  n_766;
assign n_1895 = ~x_42 &  n_1894;
assign n_1896 =  x_38 & ~x_39;
assign n_1897 =  x_35 &  n_147;
assign n_1898 = ~x_36 &  x_37;
assign n_1899 =  n_1897 &  n_1898;
assign n_1900 =  n_1896 &  n_1899;
assign n_1901 =  n_1895 &  n_1900;
assign n_1902 =  x_4743 & ~n_1901;
assign n_1903 =  x_427 &  n_1901;
assign n_1904 = ~n_1902 & ~n_1903;
assign n_1905 =  x_4743 & ~n_1904;
assign n_1906 = ~x_4743 &  n_1904;
assign n_1907 = ~n_1905 & ~n_1906;
assign n_1908 =  x_4742 & ~n_1901;
assign n_1909 =  x_426 &  n_1901;
assign n_1910 = ~n_1908 & ~n_1909;
assign n_1911 =  x_4742 & ~n_1910;
assign n_1912 = ~x_4742 &  n_1910;
assign n_1913 = ~n_1911 & ~n_1912;
assign n_1914 =  x_4741 & ~n_1901;
assign n_1915 =  x_425 &  n_1901;
assign n_1916 = ~n_1914 & ~n_1915;
assign n_1917 =  x_4741 & ~n_1916;
assign n_1918 = ~x_4741 &  n_1916;
assign n_1919 = ~n_1917 & ~n_1918;
assign n_1920 =  x_4740 & ~n_1901;
assign n_1921 =  x_424 &  n_1901;
assign n_1922 = ~n_1920 & ~n_1921;
assign n_1923 =  x_4740 & ~n_1922;
assign n_1924 = ~x_4740 &  n_1922;
assign n_1925 = ~n_1923 & ~n_1924;
assign n_1926 =  x_4739 & ~n_1901;
assign n_1927 =  x_423 &  n_1901;
assign n_1928 = ~n_1926 & ~n_1927;
assign n_1929 =  x_4739 & ~n_1928;
assign n_1930 = ~x_4739 &  n_1928;
assign n_1931 = ~n_1929 & ~n_1930;
assign n_1932 =  x_4738 & ~n_1901;
assign n_1933 =  x_422 &  n_1901;
assign n_1934 = ~n_1932 & ~n_1933;
assign n_1935 =  x_4738 & ~n_1934;
assign n_1936 = ~x_4738 &  n_1934;
assign n_1937 = ~n_1935 & ~n_1936;
assign n_1938 =  x_4737 & ~n_1901;
assign n_1939 =  x_421 &  n_1901;
assign n_1940 = ~n_1938 & ~n_1939;
assign n_1941 =  x_4737 & ~n_1940;
assign n_1942 = ~x_4737 &  n_1940;
assign n_1943 = ~n_1941 & ~n_1942;
assign n_1944 =  x_4736 & ~n_1901;
assign n_1945 =  x_420 &  n_1901;
assign n_1946 = ~n_1944 & ~n_1945;
assign n_1947 =  x_4736 & ~n_1946;
assign n_1948 = ~x_4736 &  n_1946;
assign n_1949 = ~n_1947 & ~n_1948;
assign n_1950 =  x_4735 & ~n_1901;
assign n_1951 =  x_419 &  n_1901;
assign n_1952 = ~n_1950 & ~n_1951;
assign n_1953 =  x_4735 & ~n_1952;
assign n_1954 = ~x_4735 &  n_1952;
assign n_1955 = ~n_1953 & ~n_1954;
assign n_1956 =  x_4734 & ~n_1901;
assign n_1957 =  x_418 &  n_1901;
assign n_1958 = ~n_1956 & ~n_1957;
assign n_1959 =  x_4734 & ~n_1958;
assign n_1960 = ~x_4734 &  n_1958;
assign n_1961 = ~n_1959 & ~n_1960;
assign n_1962 =  x_4733 & ~n_1901;
assign n_1963 =  x_417 &  n_1901;
assign n_1964 = ~n_1962 & ~n_1963;
assign n_1965 =  x_4733 & ~n_1964;
assign n_1966 = ~x_4733 &  n_1964;
assign n_1967 = ~n_1965 & ~n_1966;
assign n_1968 =  x_4732 & ~n_1901;
assign n_1969 =  x_416 &  n_1901;
assign n_1970 = ~n_1968 & ~n_1969;
assign n_1971 =  x_4732 & ~n_1970;
assign n_1972 = ~x_4732 &  n_1970;
assign n_1973 = ~n_1971 & ~n_1972;
assign n_1974 =  x_4731 & ~n_1901;
assign n_1975 =  x_415 &  n_1901;
assign n_1976 = ~n_1974 & ~n_1975;
assign n_1977 =  x_4731 & ~n_1976;
assign n_1978 = ~x_4731 &  n_1976;
assign n_1979 = ~n_1977 & ~n_1978;
assign n_1980 =  x_4730 & ~n_1901;
assign n_1981 =  x_414 &  n_1901;
assign n_1982 = ~n_1980 & ~n_1981;
assign n_1983 =  x_4730 & ~n_1982;
assign n_1984 = ~x_4730 &  n_1982;
assign n_1985 = ~n_1983 & ~n_1984;
assign n_1986 =  x_4729 & ~n_1901;
assign n_1987 =  x_413 &  n_1901;
assign n_1988 = ~n_1986 & ~n_1987;
assign n_1989 =  x_4729 & ~n_1988;
assign n_1990 = ~x_4729 &  n_1988;
assign n_1991 = ~n_1989 & ~n_1990;
assign n_1992 =  x_4728 & ~n_1901;
assign n_1993 =  x_412 &  n_1901;
assign n_1994 = ~n_1992 & ~n_1993;
assign n_1995 =  x_4728 & ~n_1994;
assign n_1996 = ~x_4728 &  n_1994;
assign n_1997 = ~n_1995 & ~n_1996;
assign n_1998 =  x_4727 & ~n_1901;
assign n_1999 =  x_411 &  n_1901;
assign n_2000 = ~n_1998 & ~n_1999;
assign n_2001 =  x_4727 & ~n_2000;
assign n_2002 = ~x_4727 &  n_2000;
assign n_2003 = ~n_2001 & ~n_2002;
assign n_2004 =  x_4726 & ~n_1901;
assign n_2005 =  x_410 &  n_1901;
assign n_2006 = ~n_2004 & ~n_2005;
assign n_2007 =  x_4726 & ~n_2006;
assign n_2008 = ~x_4726 &  n_2006;
assign n_2009 = ~n_2007 & ~n_2008;
assign n_2010 =  x_4725 & ~n_1901;
assign n_2011 =  x_409 &  n_1901;
assign n_2012 = ~n_2010 & ~n_2011;
assign n_2013 =  x_4725 & ~n_2012;
assign n_2014 = ~x_4725 &  n_2012;
assign n_2015 = ~n_2013 & ~n_2014;
assign n_2016 =  x_4724 & ~n_1901;
assign n_2017 =  x_408 &  n_1901;
assign n_2018 = ~n_2016 & ~n_2017;
assign n_2019 =  x_4724 & ~n_2018;
assign n_2020 = ~x_4724 &  n_2018;
assign n_2021 = ~n_2019 & ~n_2020;
assign n_2022 =  x_4723 & ~n_1901;
assign n_2023 =  x_407 &  n_1901;
assign n_2024 = ~n_2022 & ~n_2023;
assign n_2025 =  x_4723 & ~n_2024;
assign n_2026 = ~x_4723 &  n_2024;
assign n_2027 = ~n_2025 & ~n_2026;
assign n_2028 =  x_4722 & ~n_1901;
assign n_2029 =  x_406 &  n_1901;
assign n_2030 = ~n_2028 & ~n_2029;
assign n_2031 =  x_4722 & ~n_2030;
assign n_2032 = ~x_4722 &  n_2030;
assign n_2033 = ~n_2031 & ~n_2032;
assign n_2034 =  x_4721 & ~n_1901;
assign n_2035 =  x_405 &  n_1901;
assign n_2036 = ~n_2034 & ~n_2035;
assign n_2037 =  x_4721 & ~n_2036;
assign n_2038 = ~x_4721 &  n_2036;
assign n_2039 = ~n_2037 & ~n_2038;
assign n_2040 =  x_4720 & ~n_1901;
assign n_2041 =  x_404 &  n_1901;
assign n_2042 = ~n_2040 & ~n_2041;
assign n_2043 =  x_4720 & ~n_2042;
assign n_2044 = ~x_4720 &  n_2042;
assign n_2045 = ~n_2043 & ~n_2044;
assign n_2046 =  x_4719 & ~n_1901;
assign n_2047 =  x_403 &  n_1901;
assign n_2048 = ~n_2046 & ~n_2047;
assign n_2049 =  x_4719 & ~n_2048;
assign n_2050 = ~x_4719 &  n_2048;
assign n_2051 = ~n_2049 & ~n_2050;
assign n_2052 =  x_4718 & ~n_1901;
assign n_2053 =  x_402 &  n_1901;
assign n_2054 = ~n_2052 & ~n_2053;
assign n_2055 =  x_4718 & ~n_2054;
assign n_2056 = ~x_4718 &  n_2054;
assign n_2057 = ~n_2055 & ~n_2056;
assign n_2058 =  x_4717 & ~n_1901;
assign n_2059 =  x_401 &  n_1901;
assign n_2060 = ~n_2058 & ~n_2059;
assign n_2061 =  x_4717 & ~n_2060;
assign n_2062 = ~x_4717 &  n_2060;
assign n_2063 = ~n_2061 & ~n_2062;
assign n_2064 =  x_4716 & ~n_1901;
assign n_2065 =  x_400 &  n_1901;
assign n_2066 = ~n_2064 & ~n_2065;
assign n_2067 =  x_4716 & ~n_2066;
assign n_2068 = ~x_4716 &  n_2066;
assign n_2069 = ~n_2067 & ~n_2068;
assign n_2070 =  x_4715 & ~n_1901;
assign n_2071 =  x_399 &  n_1901;
assign n_2072 = ~n_2070 & ~n_2071;
assign n_2073 =  x_4715 & ~n_2072;
assign n_2074 = ~x_4715 &  n_2072;
assign n_2075 = ~n_2073 & ~n_2074;
assign n_2076 =  x_4714 & ~n_1901;
assign n_2077 =  x_398 &  n_1901;
assign n_2078 = ~n_2076 & ~n_2077;
assign n_2079 =  x_4714 & ~n_2078;
assign n_2080 = ~x_4714 &  n_2078;
assign n_2081 = ~n_2079 & ~n_2080;
assign n_2082 =  x_4713 & ~n_1901;
assign n_2083 =  x_397 &  n_1901;
assign n_2084 = ~n_2082 & ~n_2083;
assign n_2085 =  x_4713 & ~n_2084;
assign n_2086 = ~x_4713 &  n_2084;
assign n_2087 = ~n_2085 & ~n_2086;
assign n_2088 =  x_4712 & ~n_1901;
assign n_2089 =  x_396 &  n_1901;
assign n_2090 = ~n_2088 & ~n_2089;
assign n_2091 =  x_4712 & ~n_2090;
assign n_2092 = ~x_4712 &  n_2090;
assign n_2093 = ~n_2091 & ~n_2092;
assign n_2094 =  n_349 &  n_561;
assign n_2095 =  n_1039 &  n_149;
assign n_2096 =  n_2095 &  n_151;
assign n_2097 =  n_2094 &  n_2096;
assign n_2098 =  x_4711 & ~n_2097;
assign n_2099 =  i_32 &  n_2097;
assign n_2100 = ~n_2098 & ~n_2099;
assign n_2101 =  x_4711 & ~n_2100;
assign n_2102 = ~x_4711 &  n_2100;
assign n_2103 = ~n_2101 & ~n_2102;
assign n_2104 =  x_4710 & ~n_2097;
assign n_2105 =  i_31 &  n_2097;
assign n_2106 = ~n_2104 & ~n_2105;
assign n_2107 =  x_4710 & ~n_2106;
assign n_2108 = ~x_4710 &  n_2106;
assign n_2109 = ~n_2107 & ~n_2108;
assign n_2110 =  x_4709 & ~n_2097;
assign n_2111 =  i_30 &  n_2097;
assign n_2112 = ~n_2110 & ~n_2111;
assign n_2113 =  x_4709 & ~n_2112;
assign n_2114 = ~x_4709 &  n_2112;
assign n_2115 = ~n_2113 & ~n_2114;
assign n_2116 =  x_4708 & ~n_2097;
assign n_2117 =  i_29 &  n_2097;
assign n_2118 = ~n_2116 & ~n_2117;
assign n_2119 =  x_4708 & ~n_2118;
assign n_2120 = ~x_4708 &  n_2118;
assign n_2121 = ~n_2119 & ~n_2120;
assign n_2122 =  x_4707 & ~n_2097;
assign n_2123 =  i_28 &  n_2097;
assign n_2124 = ~n_2122 & ~n_2123;
assign n_2125 =  x_4707 & ~n_2124;
assign n_2126 = ~x_4707 &  n_2124;
assign n_2127 = ~n_2125 & ~n_2126;
assign n_2128 =  x_4706 & ~n_2097;
assign n_2129 =  i_27 &  n_2097;
assign n_2130 = ~n_2128 & ~n_2129;
assign n_2131 =  x_4706 & ~n_2130;
assign n_2132 = ~x_4706 &  n_2130;
assign n_2133 = ~n_2131 & ~n_2132;
assign n_2134 =  x_4705 & ~n_2097;
assign n_2135 =  i_26 &  n_2097;
assign n_2136 = ~n_2134 & ~n_2135;
assign n_2137 =  x_4705 & ~n_2136;
assign n_2138 = ~x_4705 &  n_2136;
assign n_2139 = ~n_2137 & ~n_2138;
assign n_2140 =  x_4704 & ~n_2097;
assign n_2141 =  i_25 &  n_2097;
assign n_2142 = ~n_2140 & ~n_2141;
assign n_2143 =  x_4704 & ~n_2142;
assign n_2144 = ~x_4704 &  n_2142;
assign n_2145 = ~n_2143 & ~n_2144;
assign n_2146 =  x_4703 & ~n_2097;
assign n_2147 =  i_24 &  n_2097;
assign n_2148 = ~n_2146 & ~n_2147;
assign n_2149 =  x_4703 & ~n_2148;
assign n_2150 = ~x_4703 &  n_2148;
assign n_2151 = ~n_2149 & ~n_2150;
assign n_2152 =  x_4702 & ~n_2097;
assign n_2153 =  i_23 &  n_2097;
assign n_2154 = ~n_2152 & ~n_2153;
assign n_2155 =  x_4702 & ~n_2154;
assign n_2156 = ~x_4702 &  n_2154;
assign n_2157 = ~n_2155 & ~n_2156;
assign n_2158 =  x_4701 & ~n_2097;
assign n_2159 =  i_22 &  n_2097;
assign n_2160 = ~n_2158 & ~n_2159;
assign n_2161 =  x_4701 & ~n_2160;
assign n_2162 = ~x_4701 &  n_2160;
assign n_2163 = ~n_2161 & ~n_2162;
assign n_2164 =  x_4700 & ~n_2097;
assign n_2165 =  i_21 &  n_2097;
assign n_2166 = ~n_2164 & ~n_2165;
assign n_2167 =  x_4700 & ~n_2166;
assign n_2168 = ~x_4700 &  n_2166;
assign n_2169 = ~n_2167 & ~n_2168;
assign n_2170 =  x_4699 & ~n_2097;
assign n_2171 =  i_20 &  n_2097;
assign n_2172 = ~n_2170 & ~n_2171;
assign n_2173 =  x_4699 & ~n_2172;
assign n_2174 = ~x_4699 &  n_2172;
assign n_2175 = ~n_2173 & ~n_2174;
assign n_2176 =  x_4698 & ~n_2097;
assign n_2177 =  i_19 &  n_2097;
assign n_2178 = ~n_2176 & ~n_2177;
assign n_2179 =  x_4698 & ~n_2178;
assign n_2180 = ~x_4698 &  n_2178;
assign n_2181 = ~n_2179 & ~n_2180;
assign n_2182 =  x_4697 & ~n_2097;
assign n_2183 =  i_18 &  n_2097;
assign n_2184 = ~n_2182 & ~n_2183;
assign n_2185 =  x_4697 & ~n_2184;
assign n_2186 = ~x_4697 &  n_2184;
assign n_2187 = ~n_2185 & ~n_2186;
assign n_2188 =  x_4696 & ~n_2097;
assign n_2189 =  i_17 &  n_2097;
assign n_2190 = ~n_2188 & ~n_2189;
assign n_2191 =  x_4696 & ~n_2190;
assign n_2192 = ~x_4696 &  n_2190;
assign n_2193 = ~n_2191 & ~n_2192;
assign n_2194 =  x_4695 & ~n_2097;
assign n_2195 =  i_16 &  n_2097;
assign n_2196 = ~n_2194 & ~n_2195;
assign n_2197 =  x_4695 & ~n_2196;
assign n_2198 = ~x_4695 &  n_2196;
assign n_2199 = ~n_2197 & ~n_2198;
assign n_2200 =  x_4694 & ~n_2097;
assign n_2201 =  i_15 &  n_2097;
assign n_2202 = ~n_2200 & ~n_2201;
assign n_2203 =  x_4694 & ~n_2202;
assign n_2204 = ~x_4694 &  n_2202;
assign n_2205 = ~n_2203 & ~n_2204;
assign n_2206 =  x_4693 & ~n_2097;
assign n_2207 =  i_14 &  n_2097;
assign n_2208 = ~n_2206 & ~n_2207;
assign n_2209 =  x_4693 & ~n_2208;
assign n_2210 = ~x_4693 &  n_2208;
assign n_2211 = ~n_2209 & ~n_2210;
assign n_2212 =  x_4692 & ~n_2097;
assign n_2213 =  i_13 &  n_2097;
assign n_2214 = ~n_2212 & ~n_2213;
assign n_2215 =  x_4692 & ~n_2214;
assign n_2216 = ~x_4692 &  n_2214;
assign n_2217 = ~n_2215 & ~n_2216;
assign n_2218 =  x_4691 & ~n_2097;
assign n_2219 =  i_12 &  n_2097;
assign n_2220 = ~n_2218 & ~n_2219;
assign n_2221 =  x_4691 & ~n_2220;
assign n_2222 = ~x_4691 &  n_2220;
assign n_2223 = ~n_2221 & ~n_2222;
assign n_2224 =  x_4690 & ~n_2097;
assign n_2225 =  i_11 &  n_2097;
assign n_2226 = ~n_2224 & ~n_2225;
assign n_2227 =  x_4690 & ~n_2226;
assign n_2228 = ~x_4690 &  n_2226;
assign n_2229 = ~n_2227 & ~n_2228;
assign n_2230 =  x_4689 & ~n_2097;
assign n_2231 =  i_10 &  n_2097;
assign n_2232 = ~n_2230 & ~n_2231;
assign n_2233 =  x_4689 & ~n_2232;
assign n_2234 = ~x_4689 &  n_2232;
assign n_2235 = ~n_2233 & ~n_2234;
assign n_2236 =  x_4688 & ~n_2097;
assign n_2237 =  i_9 &  n_2097;
assign n_2238 = ~n_2236 & ~n_2237;
assign n_2239 =  x_4688 & ~n_2238;
assign n_2240 = ~x_4688 &  n_2238;
assign n_2241 = ~n_2239 & ~n_2240;
assign n_2242 =  x_4687 & ~n_2097;
assign n_2243 =  i_8 &  n_2097;
assign n_2244 = ~n_2242 & ~n_2243;
assign n_2245 =  x_4687 & ~n_2244;
assign n_2246 = ~x_4687 &  n_2244;
assign n_2247 = ~n_2245 & ~n_2246;
assign n_2248 =  x_4686 & ~n_2097;
assign n_2249 =  i_7 &  n_2097;
assign n_2250 = ~n_2248 & ~n_2249;
assign n_2251 =  x_4686 & ~n_2250;
assign n_2252 = ~x_4686 &  n_2250;
assign n_2253 = ~n_2251 & ~n_2252;
assign n_2254 =  x_4685 & ~n_2097;
assign n_2255 =  i_6 &  n_2097;
assign n_2256 = ~n_2254 & ~n_2255;
assign n_2257 =  x_4685 & ~n_2256;
assign n_2258 = ~x_4685 &  n_2256;
assign n_2259 = ~n_2257 & ~n_2258;
assign n_2260 =  x_4684 & ~n_2097;
assign n_2261 =  i_5 &  n_2097;
assign n_2262 = ~n_2260 & ~n_2261;
assign n_2263 =  x_4684 & ~n_2262;
assign n_2264 = ~x_4684 &  n_2262;
assign n_2265 = ~n_2263 & ~n_2264;
assign n_2266 =  x_4683 & ~n_2097;
assign n_2267 =  i_4 &  n_2097;
assign n_2268 = ~n_2266 & ~n_2267;
assign n_2269 =  x_4683 & ~n_2268;
assign n_2270 = ~x_4683 &  n_2268;
assign n_2271 = ~n_2269 & ~n_2270;
assign n_2272 =  x_4682 & ~n_2097;
assign n_2273 =  i_3 &  n_2097;
assign n_2274 = ~n_2272 & ~n_2273;
assign n_2275 =  x_4682 & ~n_2274;
assign n_2276 = ~x_4682 &  n_2274;
assign n_2277 = ~n_2275 & ~n_2276;
assign n_2278 =  x_4681 & ~n_2097;
assign n_2279 =  i_2 &  n_2097;
assign n_2280 = ~n_2278 & ~n_2279;
assign n_2281 =  x_4681 & ~n_2280;
assign n_2282 = ~x_4681 &  n_2280;
assign n_2283 = ~n_2281 & ~n_2282;
assign n_2284 =  x_4680 & ~n_2097;
assign n_2285 =  i_1 &  n_2097;
assign n_2286 = ~n_2284 & ~n_2285;
assign n_2287 =  x_4680 & ~n_2286;
assign n_2288 = ~x_4680 &  n_2286;
assign n_2289 = ~n_2287 & ~n_2288;
assign n_2290 = ~x_38 & ~x_39;
assign n_2291 =  n_2095 &  n_2290;
assign n_2292 =  n_1895 &  n_2291;
assign n_2293 =  x_4679 & ~n_2292;
assign n_2294 =  i_32 &  n_2292;
assign n_2295 = ~n_2293 & ~n_2294;
assign n_2296 =  x_4679 & ~n_2295;
assign n_2297 = ~x_4679 &  n_2295;
assign n_2298 = ~n_2296 & ~n_2297;
assign n_2299 =  x_4678 & ~n_2292;
assign n_2300 =  i_31 &  n_2292;
assign n_2301 = ~n_2299 & ~n_2300;
assign n_2302 =  x_4678 & ~n_2301;
assign n_2303 = ~x_4678 &  n_2301;
assign n_2304 = ~n_2302 & ~n_2303;
assign n_2305 =  x_4677 & ~n_2292;
assign n_2306 =  i_30 &  n_2292;
assign n_2307 = ~n_2305 & ~n_2306;
assign n_2308 =  x_4677 & ~n_2307;
assign n_2309 = ~x_4677 &  n_2307;
assign n_2310 = ~n_2308 & ~n_2309;
assign n_2311 =  x_4676 & ~n_2292;
assign n_2312 =  i_29 &  n_2292;
assign n_2313 = ~n_2311 & ~n_2312;
assign n_2314 =  x_4676 & ~n_2313;
assign n_2315 = ~x_4676 &  n_2313;
assign n_2316 = ~n_2314 & ~n_2315;
assign n_2317 =  x_4675 & ~n_2292;
assign n_2318 =  i_28 &  n_2292;
assign n_2319 = ~n_2317 & ~n_2318;
assign n_2320 =  x_4675 & ~n_2319;
assign n_2321 = ~x_4675 &  n_2319;
assign n_2322 = ~n_2320 & ~n_2321;
assign n_2323 =  x_4674 & ~n_2292;
assign n_2324 =  i_27 &  n_2292;
assign n_2325 = ~n_2323 & ~n_2324;
assign n_2326 =  x_4674 & ~n_2325;
assign n_2327 = ~x_4674 &  n_2325;
assign n_2328 = ~n_2326 & ~n_2327;
assign n_2329 =  x_4673 & ~n_2292;
assign n_2330 =  i_26 &  n_2292;
assign n_2331 = ~n_2329 & ~n_2330;
assign n_2332 =  x_4673 & ~n_2331;
assign n_2333 = ~x_4673 &  n_2331;
assign n_2334 = ~n_2332 & ~n_2333;
assign n_2335 =  x_4672 & ~n_2292;
assign n_2336 =  i_25 &  n_2292;
assign n_2337 = ~n_2335 & ~n_2336;
assign n_2338 =  x_4672 & ~n_2337;
assign n_2339 = ~x_4672 &  n_2337;
assign n_2340 = ~n_2338 & ~n_2339;
assign n_2341 =  x_4671 & ~n_2292;
assign n_2342 =  i_24 &  n_2292;
assign n_2343 = ~n_2341 & ~n_2342;
assign n_2344 =  x_4671 & ~n_2343;
assign n_2345 = ~x_4671 &  n_2343;
assign n_2346 = ~n_2344 & ~n_2345;
assign n_2347 =  x_4670 & ~n_2292;
assign n_2348 =  i_23 &  n_2292;
assign n_2349 = ~n_2347 & ~n_2348;
assign n_2350 =  x_4670 & ~n_2349;
assign n_2351 = ~x_4670 &  n_2349;
assign n_2352 = ~n_2350 & ~n_2351;
assign n_2353 =  x_4669 & ~n_2292;
assign n_2354 =  i_22 &  n_2292;
assign n_2355 = ~n_2353 & ~n_2354;
assign n_2356 =  x_4669 & ~n_2355;
assign n_2357 = ~x_4669 &  n_2355;
assign n_2358 = ~n_2356 & ~n_2357;
assign n_2359 =  x_4668 & ~n_2292;
assign n_2360 =  i_21 &  n_2292;
assign n_2361 = ~n_2359 & ~n_2360;
assign n_2362 =  x_4668 & ~n_2361;
assign n_2363 = ~x_4668 &  n_2361;
assign n_2364 = ~n_2362 & ~n_2363;
assign n_2365 =  x_4667 & ~n_2292;
assign n_2366 =  i_20 &  n_2292;
assign n_2367 = ~n_2365 & ~n_2366;
assign n_2368 =  x_4667 & ~n_2367;
assign n_2369 = ~x_4667 &  n_2367;
assign n_2370 = ~n_2368 & ~n_2369;
assign n_2371 =  x_4666 & ~n_2292;
assign n_2372 =  i_19 &  n_2292;
assign n_2373 = ~n_2371 & ~n_2372;
assign n_2374 =  x_4666 & ~n_2373;
assign n_2375 = ~x_4666 &  n_2373;
assign n_2376 = ~n_2374 & ~n_2375;
assign n_2377 =  x_4665 & ~n_2292;
assign n_2378 =  i_18 &  n_2292;
assign n_2379 = ~n_2377 & ~n_2378;
assign n_2380 =  x_4665 & ~n_2379;
assign n_2381 = ~x_4665 &  n_2379;
assign n_2382 = ~n_2380 & ~n_2381;
assign n_2383 =  x_4664 & ~n_2292;
assign n_2384 =  i_17 &  n_2292;
assign n_2385 = ~n_2383 & ~n_2384;
assign n_2386 =  x_4664 & ~n_2385;
assign n_2387 = ~x_4664 &  n_2385;
assign n_2388 = ~n_2386 & ~n_2387;
assign n_2389 =  x_4663 & ~n_2292;
assign n_2390 =  i_16 &  n_2292;
assign n_2391 = ~n_2389 & ~n_2390;
assign n_2392 =  x_4663 & ~n_2391;
assign n_2393 = ~x_4663 &  n_2391;
assign n_2394 = ~n_2392 & ~n_2393;
assign n_2395 =  x_4662 & ~n_2292;
assign n_2396 =  i_15 &  n_2292;
assign n_2397 = ~n_2395 & ~n_2396;
assign n_2398 =  x_4662 & ~n_2397;
assign n_2399 = ~x_4662 &  n_2397;
assign n_2400 = ~n_2398 & ~n_2399;
assign n_2401 =  x_4661 & ~n_2292;
assign n_2402 =  i_14 &  n_2292;
assign n_2403 = ~n_2401 & ~n_2402;
assign n_2404 =  x_4661 & ~n_2403;
assign n_2405 = ~x_4661 &  n_2403;
assign n_2406 = ~n_2404 & ~n_2405;
assign n_2407 =  x_4660 & ~n_2292;
assign n_2408 =  i_13 &  n_2292;
assign n_2409 = ~n_2407 & ~n_2408;
assign n_2410 =  x_4660 & ~n_2409;
assign n_2411 = ~x_4660 &  n_2409;
assign n_2412 = ~n_2410 & ~n_2411;
assign n_2413 =  x_4659 & ~n_2292;
assign n_2414 =  i_12 &  n_2292;
assign n_2415 = ~n_2413 & ~n_2414;
assign n_2416 =  x_4659 & ~n_2415;
assign n_2417 = ~x_4659 &  n_2415;
assign n_2418 = ~n_2416 & ~n_2417;
assign n_2419 =  x_4658 & ~n_2292;
assign n_2420 =  i_11 &  n_2292;
assign n_2421 = ~n_2419 & ~n_2420;
assign n_2422 =  x_4658 & ~n_2421;
assign n_2423 = ~x_4658 &  n_2421;
assign n_2424 = ~n_2422 & ~n_2423;
assign n_2425 =  x_4657 & ~n_2292;
assign n_2426 =  i_10 &  n_2292;
assign n_2427 = ~n_2425 & ~n_2426;
assign n_2428 =  x_4657 & ~n_2427;
assign n_2429 = ~x_4657 &  n_2427;
assign n_2430 = ~n_2428 & ~n_2429;
assign n_2431 =  x_4656 & ~n_2292;
assign n_2432 =  i_9 &  n_2292;
assign n_2433 = ~n_2431 & ~n_2432;
assign n_2434 =  x_4656 & ~n_2433;
assign n_2435 = ~x_4656 &  n_2433;
assign n_2436 = ~n_2434 & ~n_2435;
assign n_2437 =  x_4655 & ~n_2292;
assign n_2438 =  i_8 &  n_2292;
assign n_2439 = ~n_2437 & ~n_2438;
assign n_2440 =  x_4655 & ~n_2439;
assign n_2441 = ~x_4655 &  n_2439;
assign n_2442 = ~n_2440 & ~n_2441;
assign n_2443 =  x_4654 & ~n_2292;
assign n_2444 =  i_7 &  n_2292;
assign n_2445 = ~n_2443 & ~n_2444;
assign n_2446 =  x_4654 & ~n_2445;
assign n_2447 = ~x_4654 &  n_2445;
assign n_2448 = ~n_2446 & ~n_2447;
assign n_2449 =  x_4653 & ~n_2292;
assign n_2450 =  i_6 &  n_2292;
assign n_2451 = ~n_2449 & ~n_2450;
assign n_2452 =  x_4653 & ~n_2451;
assign n_2453 = ~x_4653 &  n_2451;
assign n_2454 = ~n_2452 & ~n_2453;
assign n_2455 =  x_4652 & ~n_2292;
assign n_2456 =  i_5 &  n_2292;
assign n_2457 = ~n_2455 & ~n_2456;
assign n_2458 =  x_4652 & ~n_2457;
assign n_2459 = ~x_4652 &  n_2457;
assign n_2460 = ~n_2458 & ~n_2459;
assign n_2461 =  x_4651 & ~n_2292;
assign n_2462 =  i_4 &  n_2292;
assign n_2463 = ~n_2461 & ~n_2462;
assign n_2464 =  x_4651 & ~n_2463;
assign n_2465 = ~x_4651 &  n_2463;
assign n_2466 = ~n_2464 & ~n_2465;
assign n_2467 =  x_4650 & ~n_2292;
assign n_2468 =  i_3 &  n_2292;
assign n_2469 = ~n_2467 & ~n_2468;
assign n_2470 =  x_4650 & ~n_2469;
assign n_2471 = ~x_4650 &  n_2469;
assign n_2472 = ~n_2470 & ~n_2471;
assign n_2473 =  x_4649 & ~n_2292;
assign n_2474 =  i_2 &  n_2292;
assign n_2475 = ~n_2473 & ~n_2474;
assign n_2476 =  x_4649 & ~n_2475;
assign n_2477 = ~x_4649 &  n_2475;
assign n_2478 = ~n_2476 & ~n_2477;
assign n_2479 =  x_4648 & ~n_2292;
assign n_2480 =  i_1 &  n_2292;
assign n_2481 = ~n_2479 & ~n_2480;
assign n_2482 =  x_4648 & ~n_2481;
assign n_2483 = ~x_4648 &  n_2481;
assign n_2484 = ~n_2482 & ~n_2483;
assign n_2485 =  x_36 &  x_37;
assign n_2486 =  n_1897 &  n_2485;
assign n_2487 =  n_2290 &  n_2486;
assign n_2488 =  n_2094 &  n_2487;
assign n_2489 =  x_4647 & ~n_2488;
assign n_2490 =  i_32 &  n_2488;
assign n_2491 = ~n_2489 & ~n_2490;
assign n_2492 =  x_4647 & ~n_2491;
assign n_2493 = ~x_4647 &  n_2491;
assign n_2494 = ~n_2492 & ~n_2493;
assign n_2495 =  x_4646 & ~n_2488;
assign n_2496 =  i_31 &  n_2488;
assign n_2497 = ~n_2495 & ~n_2496;
assign n_2498 =  x_4646 & ~n_2497;
assign n_2499 = ~x_4646 &  n_2497;
assign n_2500 = ~n_2498 & ~n_2499;
assign n_2501 =  x_4645 & ~n_2488;
assign n_2502 =  i_30 &  n_2488;
assign n_2503 = ~n_2501 & ~n_2502;
assign n_2504 =  x_4645 & ~n_2503;
assign n_2505 = ~x_4645 &  n_2503;
assign n_2506 = ~n_2504 & ~n_2505;
assign n_2507 =  x_4644 & ~n_2488;
assign n_2508 =  i_29 &  n_2488;
assign n_2509 = ~n_2507 & ~n_2508;
assign n_2510 =  x_4644 & ~n_2509;
assign n_2511 = ~x_4644 &  n_2509;
assign n_2512 = ~n_2510 & ~n_2511;
assign n_2513 =  x_4643 & ~n_2488;
assign n_2514 =  i_28 &  n_2488;
assign n_2515 = ~n_2513 & ~n_2514;
assign n_2516 =  x_4643 & ~n_2515;
assign n_2517 = ~x_4643 &  n_2515;
assign n_2518 = ~n_2516 & ~n_2517;
assign n_2519 =  x_4642 & ~n_2488;
assign n_2520 =  i_27 &  n_2488;
assign n_2521 = ~n_2519 & ~n_2520;
assign n_2522 =  x_4642 & ~n_2521;
assign n_2523 = ~x_4642 &  n_2521;
assign n_2524 = ~n_2522 & ~n_2523;
assign n_2525 =  x_4641 & ~n_2488;
assign n_2526 =  i_26 &  n_2488;
assign n_2527 = ~n_2525 & ~n_2526;
assign n_2528 =  x_4641 & ~n_2527;
assign n_2529 = ~x_4641 &  n_2527;
assign n_2530 = ~n_2528 & ~n_2529;
assign n_2531 =  x_4640 & ~n_2488;
assign n_2532 =  i_25 &  n_2488;
assign n_2533 = ~n_2531 & ~n_2532;
assign n_2534 =  x_4640 & ~n_2533;
assign n_2535 = ~x_4640 &  n_2533;
assign n_2536 = ~n_2534 & ~n_2535;
assign n_2537 =  x_4639 & ~n_2488;
assign n_2538 =  i_24 &  n_2488;
assign n_2539 = ~n_2537 & ~n_2538;
assign n_2540 =  x_4639 & ~n_2539;
assign n_2541 = ~x_4639 &  n_2539;
assign n_2542 = ~n_2540 & ~n_2541;
assign n_2543 =  x_4638 & ~n_2488;
assign n_2544 =  i_23 &  n_2488;
assign n_2545 = ~n_2543 & ~n_2544;
assign n_2546 =  x_4638 & ~n_2545;
assign n_2547 = ~x_4638 &  n_2545;
assign n_2548 = ~n_2546 & ~n_2547;
assign n_2549 =  x_4637 & ~n_2488;
assign n_2550 =  i_22 &  n_2488;
assign n_2551 = ~n_2549 & ~n_2550;
assign n_2552 =  x_4637 & ~n_2551;
assign n_2553 = ~x_4637 &  n_2551;
assign n_2554 = ~n_2552 & ~n_2553;
assign n_2555 =  x_4636 & ~n_2488;
assign n_2556 =  i_21 &  n_2488;
assign n_2557 = ~n_2555 & ~n_2556;
assign n_2558 =  x_4636 & ~n_2557;
assign n_2559 = ~x_4636 &  n_2557;
assign n_2560 = ~n_2558 & ~n_2559;
assign n_2561 =  x_4635 & ~n_2488;
assign n_2562 =  i_20 &  n_2488;
assign n_2563 = ~n_2561 & ~n_2562;
assign n_2564 =  x_4635 & ~n_2563;
assign n_2565 = ~x_4635 &  n_2563;
assign n_2566 = ~n_2564 & ~n_2565;
assign n_2567 =  x_4634 & ~n_2488;
assign n_2568 =  i_19 &  n_2488;
assign n_2569 = ~n_2567 & ~n_2568;
assign n_2570 =  x_4634 & ~n_2569;
assign n_2571 = ~x_4634 &  n_2569;
assign n_2572 = ~n_2570 & ~n_2571;
assign n_2573 =  x_4633 & ~n_2488;
assign n_2574 =  i_18 &  n_2488;
assign n_2575 = ~n_2573 & ~n_2574;
assign n_2576 =  x_4633 & ~n_2575;
assign n_2577 = ~x_4633 &  n_2575;
assign n_2578 = ~n_2576 & ~n_2577;
assign n_2579 =  x_4632 & ~n_2488;
assign n_2580 =  i_17 &  n_2488;
assign n_2581 = ~n_2579 & ~n_2580;
assign n_2582 =  x_4632 & ~n_2581;
assign n_2583 = ~x_4632 &  n_2581;
assign n_2584 = ~n_2582 & ~n_2583;
assign n_2585 =  x_4631 & ~n_2488;
assign n_2586 =  i_16 &  n_2488;
assign n_2587 = ~n_2585 & ~n_2586;
assign n_2588 =  x_4631 & ~n_2587;
assign n_2589 = ~x_4631 &  n_2587;
assign n_2590 = ~n_2588 & ~n_2589;
assign n_2591 =  x_4630 & ~n_2488;
assign n_2592 =  i_15 &  n_2488;
assign n_2593 = ~n_2591 & ~n_2592;
assign n_2594 =  x_4630 & ~n_2593;
assign n_2595 = ~x_4630 &  n_2593;
assign n_2596 = ~n_2594 & ~n_2595;
assign n_2597 =  x_4629 & ~n_2488;
assign n_2598 =  i_14 &  n_2488;
assign n_2599 = ~n_2597 & ~n_2598;
assign n_2600 =  x_4629 & ~n_2599;
assign n_2601 = ~x_4629 &  n_2599;
assign n_2602 = ~n_2600 & ~n_2601;
assign n_2603 =  x_4628 & ~n_2488;
assign n_2604 =  i_13 &  n_2488;
assign n_2605 = ~n_2603 & ~n_2604;
assign n_2606 =  x_4628 & ~n_2605;
assign n_2607 = ~x_4628 &  n_2605;
assign n_2608 = ~n_2606 & ~n_2607;
assign n_2609 =  x_4627 & ~n_2488;
assign n_2610 =  i_12 &  n_2488;
assign n_2611 = ~n_2609 & ~n_2610;
assign n_2612 =  x_4627 & ~n_2611;
assign n_2613 = ~x_4627 &  n_2611;
assign n_2614 = ~n_2612 & ~n_2613;
assign n_2615 =  x_4626 & ~n_2488;
assign n_2616 =  i_11 &  n_2488;
assign n_2617 = ~n_2615 & ~n_2616;
assign n_2618 =  x_4626 & ~n_2617;
assign n_2619 = ~x_4626 &  n_2617;
assign n_2620 = ~n_2618 & ~n_2619;
assign n_2621 =  x_4625 & ~n_2488;
assign n_2622 =  i_10 &  n_2488;
assign n_2623 = ~n_2621 & ~n_2622;
assign n_2624 =  x_4625 & ~n_2623;
assign n_2625 = ~x_4625 &  n_2623;
assign n_2626 = ~n_2624 & ~n_2625;
assign n_2627 =  x_4624 & ~n_2488;
assign n_2628 =  i_9 &  n_2488;
assign n_2629 = ~n_2627 & ~n_2628;
assign n_2630 =  x_4624 & ~n_2629;
assign n_2631 = ~x_4624 &  n_2629;
assign n_2632 = ~n_2630 & ~n_2631;
assign n_2633 =  x_4623 & ~n_2488;
assign n_2634 =  i_8 &  n_2488;
assign n_2635 = ~n_2633 & ~n_2634;
assign n_2636 =  x_4623 & ~n_2635;
assign n_2637 = ~x_4623 &  n_2635;
assign n_2638 = ~n_2636 & ~n_2637;
assign n_2639 =  x_4622 & ~n_2488;
assign n_2640 =  i_7 &  n_2488;
assign n_2641 = ~n_2639 & ~n_2640;
assign n_2642 =  x_4622 & ~n_2641;
assign n_2643 = ~x_4622 &  n_2641;
assign n_2644 = ~n_2642 & ~n_2643;
assign n_2645 =  x_4621 & ~n_2488;
assign n_2646 =  i_6 &  n_2488;
assign n_2647 = ~n_2645 & ~n_2646;
assign n_2648 =  x_4621 & ~n_2647;
assign n_2649 = ~x_4621 &  n_2647;
assign n_2650 = ~n_2648 & ~n_2649;
assign n_2651 =  x_4620 & ~n_2488;
assign n_2652 =  i_5 &  n_2488;
assign n_2653 = ~n_2651 & ~n_2652;
assign n_2654 =  x_4620 & ~n_2653;
assign n_2655 = ~x_4620 &  n_2653;
assign n_2656 = ~n_2654 & ~n_2655;
assign n_2657 =  x_4619 & ~n_2488;
assign n_2658 =  i_4 &  n_2488;
assign n_2659 = ~n_2657 & ~n_2658;
assign n_2660 =  x_4619 & ~n_2659;
assign n_2661 = ~x_4619 &  n_2659;
assign n_2662 = ~n_2660 & ~n_2661;
assign n_2663 =  x_4618 & ~n_2488;
assign n_2664 =  i_3 &  n_2488;
assign n_2665 = ~n_2663 & ~n_2664;
assign n_2666 =  x_4618 & ~n_2665;
assign n_2667 = ~x_4618 &  n_2665;
assign n_2668 = ~n_2666 & ~n_2667;
assign n_2669 =  x_4617 & ~n_2488;
assign n_2670 =  i_2 &  n_2488;
assign n_2671 = ~n_2669 & ~n_2670;
assign n_2672 =  x_4617 & ~n_2671;
assign n_2673 = ~x_4617 &  n_2671;
assign n_2674 = ~n_2672 & ~n_2673;
assign n_2675 =  x_4616 & ~n_2488;
assign n_2676 =  i_1 &  n_2488;
assign n_2677 = ~n_2675 & ~n_2676;
assign n_2678 =  x_4616 & ~n_2677;
assign n_2679 = ~x_4616 &  n_2677;
assign n_2680 = ~n_2678 & ~n_2679;
assign n_2681 = ~x_41 &  n_759;
assign n_2682 =  n_1037 &  n_2681;
assign n_2683 =  x_36 & ~x_37;
assign n_2684 =  n_1897 &  n_2683;
assign n_2685 =  x_38 &  n_2684;
assign n_2686 =  n_2682 &  n_2685;
assign n_2687 =  x_4615 & ~n_2686;
assign n_2688 =  i_32 &  n_2686;
assign n_2689 = ~n_2687 & ~n_2688;
assign n_2690 =  x_4615 & ~n_2689;
assign n_2691 = ~x_4615 &  n_2689;
assign n_2692 = ~n_2690 & ~n_2691;
assign n_2693 =  x_4614 & ~n_2686;
assign n_2694 =  i_31 &  n_2686;
assign n_2695 = ~n_2693 & ~n_2694;
assign n_2696 =  x_4614 & ~n_2695;
assign n_2697 = ~x_4614 &  n_2695;
assign n_2698 = ~n_2696 & ~n_2697;
assign n_2699 =  x_4613 & ~n_2686;
assign n_2700 =  i_30 &  n_2686;
assign n_2701 = ~n_2699 & ~n_2700;
assign n_2702 =  x_4613 & ~n_2701;
assign n_2703 = ~x_4613 &  n_2701;
assign n_2704 = ~n_2702 & ~n_2703;
assign n_2705 =  x_4612 & ~n_2686;
assign n_2706 =  i_29 &  n_2686;
assign n_2707 = ~n_2705 & ~n_2706;
assign n_2708 =  x_4612 & ~n_2707;
assign n_2709 = ~x_4612 &  n_2707;
assign n_2710 = ~n_2708 & ~n_2709;
assign n_2711 =  x_4611 & ~n_2686;
assign n_2712 =  i_28 &  n_2686;
assign n_2713 = ~n_2711 & ~n_2712;
assign n_2714 =  x_4611 & ~n_2713;
assign n_2715 = ~x_4611 &  n_2713;
assign n_2716 = ~n_2714 & ~n_2715;
assign n_2717 =  x_4610 & ~n_2686;
assign n_2718 =  i_27 &  n_2686;
assign n_2719 = ~n_2717 & ~n_2718;
assign n_2720 =  x_4610 & ~n_2719;
assign n_2721 = ~x_4610 &  n_2719;
assign n_2722 = ~n_2720 & ~n_2721;
assign n_2723 =  x_4609 & ~n_2686;
assign n_2724 =  i_26 &  n_2686;
assign n_2725 = ~n_2723 & ~n_2724;
assign n_2726 =  x_4609 & ~n_2725;
assign n_2727 = ~x_4609 &  n_2725;
assign n_2728 = ~n_2726 & ~n_2727;
assign n_2729 =  x_4608 & ~n_2686;
assign n_2730 =  i_25 &  n_2686;
assign n_2731 = ~n_2729 & ~n_2730;
assign n_2732 =  x_4608 & ~n_2731;
assign n_2733 = ~x_4608 &  n_2731;
assign n_2734 = ~n_2732 & ~n_2733;
assign n_2735 =  x_4607 & ~n_2686;
assign n_2736 =  i_24 &  n_2686;
assign n_2737 = ~n_2735 & ~n_2736;
assign n_2738 =  x_4607 & ~n_2737;
assign n_2739 = ~x_4607 &  n_2737;
assign n_2740 = ~n_2738 & ~n_2739;
assign n_2741 =  x_4606 & ~n_2686;
assign n_2742 =  i_23 &  n_2686;
assign n_2743 = ~n_2741 & ~n_2742;
assign n_2744 =  x_4606 & ~n_2743;
assign n_2745 = ~x_4606 &  n_2743;
assign n_2746 = ~n_2744 & ~n_2745;
assign n_2747 =  x_4605 & ~n_2686;
assign n_2748 =  i_22 &  n_2686;
assign n_2749 = ~n_2747 & ~n_2748;
assign n_2750 =  x_4605 & ~n_2749;
assign n_2751 = ~x_4605 &  n_2749;
assign n_2752 = ~n_2750 & ~n_2751;
assign n_2753 =  x_4604 & ~n_2686;
assign n_2754 =  i_21 &  n_2686;
assign n_2755 = ~n_2753 & ~n_2754;
assign n_2756 =  x_4604 & ~n_2755;
assign n_2757 = ~x_4604 &  n_2755;
assign n_2758 = ~n_2756 & ~n_2757;
assign n_2759 =  x_4603 & ~n_2686;
assign n_2760 =  i_20 &  n_2686;
assign n_2761 = ~n_2759 & ~n_2760;
assign n_2762 =  x_4603 & ~n_2761;
assign n_2763 = ~x_4603 &  n_2761;
assign n_2764 = ~n_2762 & ~n_2763;
assign n_2765 =  x_4602 & ~n_2686;
assign n_2766 =  i_19 &  n_2686;
assign n_2767 = ~n_2765 & ~n_2766;
assign n_2768 =  x_4602 & ~n_2767;
assign n_2769 = ~x_4602 &  n_2767;
assign n_2770 = ~n_2768 & ~n_2769;
assign n_2771 =  x_4601 & ~n_2686;
assign n_2772 =  i_18 &  n_2686;
assign n_2773 = ~n_2771 & ~n_2772;
assign n_2774 =  x_4601 & ~n_2773;
assign n_2775 = ~x_4601 &  n_2773;
assign n_2776 = ~n_2774 & ~n_2775;
assign n_2777 =  x_4600 & ~n_2686;
assign n_2778 =  i_17 &  n_2686;
assign n_2779 = ~n_2777 & ~n_2778;
assign n_2780 =  x_4600 & ~n_2779;
assign n_2781 = ~x_4600 &  n_2779;
assign n_2782 = ~n_2780 & ~n_2781;
assign n_2783 =  x_4599 & ~n_2686;
assign n_2784 =  i_16 &  n_2686;
assign n_2785 = ~n_2783 & ~n_2784;
assign n_2786 =  x_4599 & ~n_2785;
assign n_2787 = ~x_4599 &  n_2785;
assign n_2788 = ~n_2786 & ~n_2787;
assign n_2789 =  x_4598 & ~n_2686;
assign n_2790 =  i_15 &  n_2686;
assign n_2791 = ~n_2789 & ~n_2790;
assign n_2792 =  x_4598 & ~n_2791;
assign n_2793 = ~x_4598 &  n_2791;
assign n_2794 = ~n_2792 & ~n_2793;
assign n_2795 =  x_4597 & ~n_2686;
assign n_2796 =  i_14 &  n_2686;
assign n_2797 = ~n_2795 & ~n_2796;
assign n_2798 =  x_4597 & ~n_2797;
assign n_2799 = ~x_4597 &  n_2797;
assign n_2800 = ~n_2798 & ~n_2799;
assign n_2801 =  x_4596 & ~n_2686;
assign n_2802 =  i_13 &  n_2686;
assign n_2803 = ~n_2801 & ~n_2802;
assign n_2804 =  x_4596 & ~n_2803;
assign n_2805 = ~x_4596 &  n_2803;
assign n_2806 = ~n_2804 & ~n_2805;
assign n_2807 =  x_4595 & ~n_2686;
assign n_2808 =  i_12 &  n_2686;
assign n_2809 = ~n_2807 & ~n_2808;
assign n_2810 =  x_4595 & ~n_2809;
assign n_2811 = ~x_4595 &  n_2809;
assign n_2812 = ~n_2810 & ~n_2811;
assign n_2813 =  x_4594 & ~n_2686;
assign n_2814 =  i_11 &  n_2686;
assign n_2815 = ~n_2813 & ~n_2814;
assign n_2816 =  x_4594 & ~n_2815;
assign n_2817 = ~x_4594 &  n_2815;
assign n_2818 = ~n_2816 & ~n_2817;
assign n_2819 =  x_4593 & ~n_2686;
assign n_2820 =  i_10 &  n_2686;
assign n_2821 = ~n_2819 & ~n_2820;
assign n_2822 =  x_4593 & ~n_2821;
assign n_2823 = ~x_4593 &  n_2821;
assign n_2824 = ~n_2822 & ~n_2823;
assign n_2825 =  x_4592 & ~n_2686;
assign n_2826 =  i_9 &  n_2686;
assign n_2827 = ~n_2825 & ~n_2826;
assign n_2828 =  x_4592 & ~n_2827;
assign n_2829 = ~x_4592 &  n_2827;
assign n_2830 = ~n_2828 & ~n_2829;
assign n_2831 =  x_4591 & ~n_2686;
assign n_2832 =  i_8 &  n_2686;
assign n_2833 = ~n_2831 & ~n_2832;
assign n_2834 =  x_4591 & ~n_2833;
assign n_2835 = ~x_4591 &  n_2833;
assign n_2836 = ~n_2834 & ~n_2835;
assign n_2837 =  x_4590 & ~n_2686;
assign n_2838 =  i_7 &  n_2686;
assign n_2839 = ~n_2837 & ~n_2838;
assign n_2840 =  x_4590 & ~n_2839;
assign n_2841 = ~x_4590 &  n_2839;
assign n_2842 = ~n_2840 & ~n_2841;
assign n_2843 =  x_4589 & ~n_2686;
assign n_2844 =  i_6 &  n_2686;
assign n_2845 = ~n_2843 & ~n_2844;
assign n_2846 =  x_4589 & ~n_2845;
assign n_2847 = ~x_4589 &  n_2845;
assign n_2848 = ~n_2846 & ~n_2847;
assign n_2849 =  x_4588 & ~n_2686;
assign n_2850 =  i_5 &  n_2686;
assign n_2851 = ~n_2849 & ~n_2850;
assign n_2852 =  x_4588 & ~n_2851;
assign n_2853 = ~x_4588 &  n_2851;
assign n_2854 = ~n_2852 & ~n_2853;
assign n_2855 =  x_4587 & ~n_2686;
assign n_2856 =  i_4 &  n_2686;
assign n_2857 = ~n_2855 & ~n_2856;
assign n_2858 =  x_4587 & ~n_2857;
assign n_2859 = ~x_4587 &  n_2857;
assign n_2860 = ~n_2858 & ~n_2859;
assign n_2861 =  x_4586 & ~n_2686;
assign n_2862 =  i_3 &  n_2686;
assign n_2863 = ~n_2861 & ~n_2862;
assign n_2864 =  x_4586 & ~n_2863;
assign n_2865 = ~x_4586 &  n_2863;
assign n_2866 = ~n_2864 & ~n_2865;
assign n_2867 =  x_4585 & ~n_2686;
assign n_2868 =  i_2 &  n_2686;
assign n_2869 = ~n_2867 & ~n_2868;
assign n_2870 =  x_4585 & ~n_2869;
assign n_2871 = ~x_4585 &  n_2869;
assign n_2872 = ~n_2870 & ~n_2871;
assign n_2873 =  x_4584 & ~n_2686;
assign n_2874 =  i_1 &  n_2686;
assign n_2875 = ~n_2873 & ~n_2874;
assign n_2876 =  x_4584 & ~n_2875;
assign n_2877 = ~x_4584 &  n_2875;
assign n_2878 = ~n_2876 & ~n_2877;
assign n_2879 =  x_37 & ~x_38;
assign n_2880 =  n_1305 &  n_2879;
assign n_2881 =  n_765 &  n_2880;
assign n_2882 = ~x_43 &  n_2881;
assign n_2883 =  n_1 &  n_2882;
assign n_2884 =  x_4424 &  n_2883;
assign n_2885 = ~n_1 &  n_2882;
assign n_2886 =  i_32 &  n_2885;
assign n_2887 =  x_4583 & ~n_2882;
assign n_2888 = ~n_2886 & ~n_2887;
assign n_2889 = ~n_2884 &  n_2888;
assign n_2890 =  x_4583 & ~n_2889;
assign n_2891 = ~x_4583 &  n_2889;
assign n_2892 = ~n_2890 & ~n_2891;
assign n_2893 =  x_4423 &  n_2883;
assign n_2894 =  i_31 &  n_2885;
assign n_2895 =  x_4582 & ~n_2882;
assign n_2896 = ~n_2894 & ~n_2895;
assign n_2897 = ~n_2893 &  n_2896;
assign n_2898 =  x_4582 & ~n_2897;
assign n_2899 = ~x_4582 &  n_2897;
assign n_2900 = ~n_2898 & ~n_2899;
assign n_2901 =  x_4422 &  n_2883;
assign n_2902 =  i_30 &  n_2885;
assign n_2903 =  x_4581 & ~n_2882;
assign n_2904 = ~n_2902 & ~n_2903;
assign n_2905 = ~n_2901 &  n_2904;
assign n_2906 =  x_4581 & ~n_2905;
assign n_2907 = ~x_4581 &  n_2905;
assign n_2908 = ~n_2906 & ~n_2907;
assign n_2909 =  x_4421 &  n_2883;
assign n_2910 =  i_29 &  n_2885;
assign n_2911 =  x_4580 & ~n_2882;
assign n_2912 = ~n_2910 & ~n_2911;
assign n_2913 = ~n_2909 &  n_2912;
assign n_2914 =  x_4580 & ~n_2913;
assign n_2915 = ~x_4580 &  n_2913;
assign n_2916 = ~n_2914 & ~n_2915;
assign n_2917 =  x_4420 &  n_2883;
assign n_2918 =  i_28 &  n_2885;
assign n_2919 =  x_4579 & ~n_2882;
assign n_2920 = ~n_2918 & ~n_2919;
assign n_2921 = ~n_2917 &  n_2920;
assign n_2922 =  x_4579 & ~n_2921;
assign n_2923 = ~x_4579 &  n_2921;
assign n_2924 = ~n_2922 & ~n_2923;
assign n_2925 =  x_4419 &  n_2883;
assign n_2926 =  i_27 &  n_2885;
assign n_2927 =  x_4578 & ~n_2882;
assign n_2928 = ~n_2926 & ~n_2927;
assign n_2929 = ~n_2925 &  n_2928;
assign n_2930 =  x_4578 & ~n_2929;
assign n_2931 = ~x_4578 &  n_2929;
assign n_2932 = ~n_2930 & ~n_2931;
assign n_2933 =  x_4418 &  n_2883;
assign n_2934 =  i_26 &  n_2885;
assign n_2935 =  x_4577 & ~n_2882;
assign n_2936 = ~n_2934 & ~n_2935;
assign n_2937 = ~n_2933 &  n_2936;
assign n_2938 =  x_4577 & ~n_2937;
assign n_2939 = ~x_4577 &  n_2937;
assign n_2940 = ~n_2938 & ~n_2939;
assign n_2941 =  x_4417 &  n_2883;
assign n_2942 =  i_25 &  n_2885;
assign n_2943 =  x_4576 & ~n_2882;
assign n_2944 = ~n_2942 & ~n_2943;
assign n_2945 = ~n_2941 &  n_2944;
assign n_2946 =  x_4576 & ~n_2945;
assign n_2947 = ~x_4576 &  n_2945;
assign n_2948 = ~n_2946 & ~n_2947;
assign n_2949 =  x_4416 &  n_2883;
assign n_2950 =  i_24 &  n_2885;
assign n_2951 =  x_4575 & ~n_2882;
assign n_2952 = ~n_2950 & ~n_2951;
assign n_2953 = ~n_2949 &  n_2952;
assign n_2954 =  x_4575 & ~n_2953;
assign n_2955 = ~x_4575 &  n_2953;
assign n_2956 = ~n_2954 & ~n_2955;
assign n_2957 =  x_4415 &  n_2883;
assign n_2958 =  i_23 &  n_2885;
assign n_2959 =  x_4574 & ~n_2882;
assign n_2960 = ~n_2958 & ~n_2959;
assign n_2961 = ~n_2957 &  n_2960;
assign n_2962 =  x_4574 & ~n_2961;
assign n_2963 = ~x_4574 &  n_2961;
assign n_2964 = ~n_2962 & ~n_2963;
assign n_2965 =  x_4414 &  n_2883;
assign n_2966 =  i_22 &  n_2885;
assign n_2967 =  x_4573 & ~n_2882;
assign n_2968 = ~n_2966 & ~n_2967;
assign n_2969 = ~n_2965 &  n_2968;
assign n_2970 =  x_4573 & ~n_2969;
assign n_2971 = ~x_4573 &  n_2969;
assign n_2972 = ~n_2970 & ~n_2971;
assign n_2973 =  x_4413 &  n_2883;
assign n_2974 =  i_21 &  n_2885;
assign n_2975 =  x_4572 & ~n_2882;
assign n_2976 = ~n_2974 & ~n_2975;
assign n_2977 = ~n_2973 &  n_2976;
assign n_2978 =  x_4572 & ~n_2977;
assign n_2979 = ~x_4572 &  n_2977;
assign n_2980 = ~n_2978 & ~n_2979;
assign n_2981 =  x_4412 &  n_2883;
assign n_2982 =  i_20 &  n_2885;
assign n_2983 =  x_4571 & ~n_2882;
assign n_2984 = ~n_2982 & ~n_2983;
assign n_2985 = ~n_2981 &  n_2984;
assign n_2986 =  x_4571 & ~n_2985;
assign n_2987 = ~x_4571 &  n_2985;
assign n_2988 = ~n_2986 & ~n_2987;
assign n_2989 =  x_4411 &  n_2883;
assign n_2990 =  i_19 &  n_2885;
assign n_2991 =  x_4570 & ~n_2882;
assign n_2992 = ~n_2990 & ~n_2991;
assign n_2993 = ~n_2989 &  n_2992;
assign n_2994 =  x_4570 & ~n_2993;
assign n_2995 = ~x_4570 &  n_2993;
assign n_2996 = ~n_2994 & ~n_2995;
assign n_2997 =  x_4410 &  n_2883;
assign n_2998 =  i_18 &  n_2885;
assign n_2999 =  x_4569 & ~n_2882;
assign n_3000 = ~n_2998 & ~n_2999;
assign n_3001 = ~n_2997 &  n_3000;
assign n_3002 =  x_4569 & ~n_3001;
assign n_3003 = ~x_4569 &  n_3001;
assign n_3004 = ~n_3002 & ~n_3003;
assign n_3005 =  x_4409 &  n_2883;
assign n_3006 =  i_17 &  n_2885;
assign n_3007 =  x_4568 & ~n_2882;
assign n_3008 = ~n_3006 & ~n_3007;
assign n_3009 = ~n_3005 &  n_3008;
assign n_3010 =  x_4568 & ~n_3009;
assign n_3011 = ~x_4568 &  n_3009;
assign n_3012 = ~n_3010 & ~n_3011;
assign n_3013 =  x_4408 &  n_2883;
assign n_3014 =  i_16 &  n_2885;
assign n_3015 =  x_4567 & ~n_2882;
assign n_3016 = ~n_3014 & ~n_3015;
assign n_3017 = ~n_3013 &  n_3016;
assign n_3018 =  x_4567 & ~n_3017;
assign n_3019 = ~x_4567 &  n_3017;
assign n_3020 = ~n_3018 & ~n_3019;
assign n_3021 =  x_4407 &  n_2883;
assign n_3022 =  i_15 &  n_2885;
assign n_3023 =  x_4566 & ~n_2882;
assign n_3024 = ~n_3022 & ~n_3023;
assign n_3025 = ~n_3021 &  n_3024;
assign n_3026 =  x_4566 & ~n_3025;
assign n_3027 = ~x_4566 &  n_3025;
assign n_3028 = ~n_3026 & ~n_3027;
assign n_3029 =  x_4406 &  n_2883;
assign n_3030 =  i_14 &  n_2885;
assign n_3031 =  x_4565 & ~n_2882;
assign n_3032 = ~n_3030 & ~n_3031;
assign n_3033 = ~n_3029 &  n_3032;
assign n_3034 =  x_4565 & ~n_3033;
assign n_3035 = ~x_4565 &  n_3033;
assign n_3036 = ~n_3034 & ~n_3035;
assign n_3037 =  x_4405 &  n_2883;
assign n_3038 =  i_13 &  n_2885;
assign n_3039 =  x_4564 & ~n_2882;
assign n_3040 = ~n_3038 & ~n_3039;
assign n_3041 = ~n_3037 &  n_3040;
assign n_3042 =  x_4564 & ~n_3041;
assign n_3043 = ~x_4564 &  n_3041;
assign n_3044 = ~n_3042 & ~n_3043;
assign n_3045 =  x_4404 &  n_2883;
assign n_3046 =  i_12 &  n_2885;
assign n_3047 =  x_4563 & ~n_2882;
assign n_3048 = ~n_3046 & ~n_3047;
assign n_3049 = ~n_3045 &  n_3048;
assign n_3050 =  x_4563 & ~n_3049;
assign n_3051 = ~x_4563 &  n_3049;
assign n_3052 = ~n_3050 & ~n_3051;
assign n_3053 =  x_4403 &  n_2883;
assign n_3054 =  i_11 &  n_2885;
assign n_3055 =  x_4562 & ~n_2882;
assign n_3056 = ~n_3054 & ~n_3055;
assign n_3057 = ~n_3053 &  n_3056;
assign n_3058 =  x_4562 & ~n_3057;
assign n_3059 = ~x_4562 &  n_3057;
assign n_3060 = ~n_3058 & ~n_3059;
assign n_3061 =  x_4402 &  n_2883;
assign n_3062 =  i_10 &  n_2885;
assign n_3063 =  x_4561 & ~n_2882;
assign n_3064 = ~n_3062 & ~n_3063;
assign n_3065 = ~n_3061 &  n_3064;
assign n_3066 =  x_4561 & ~n_3065;
assign n_3067 = ~x_4561 &  n_3065;
assign n_3068 = ~n_3066 & ~n_3067;
assign n_3069 =  x_4401 &  n_2883;
assign n_3070 =  i_9 &  n_2885;
assign n_3071 =  x_4560 & ~n_2882;
assign n_3072 = ~n_3070 & ~n_3071;
assign n_3073 = ~n_3069 &  n_3072;
assign n_3074 =  x_4560 & ~n_3073;
assign n_3075 = ~x_4560 &  n_3073;
assign n_3076 = ~n_3074 & ~n_3075;
assign n_3077 =  x_4400 &  n_2883;
assign n_3078 =  i_8 &  n_2885;
assign n_3079 =  x_4559 & ~n_2882;
assign n_3080 = ~n_3078 & ~n_3079;
assign n_3081 = ~n_3077 &  n_3080;
assign n_3082 =  x_4559 & ~n_3081;
assign n_3083 = ~x_4559 &  n_3081;
assign n_3084 = ~n_3082 & ~n_3083;
assign n_3085 =  x_4399 &  n_2883;
assign n_3086 =  i_7 &  n_2885;
assign n_3087 =  x_4558 & ~n_2882;
assign n_3088 = ~n_3086 & ~n_3087;
assign n_3089 = ~n_3085 &  n_3088;
assign n_3090 =  x_4558 & ~n_3089;
assign n_3091 = ~x_4558 &  n_3089;
assign n_3092 = ~n_3090 & ~n_3091;
assign n_3093 =  x_4398 &  n_2883;
assign n_3094 =  i_6 &  n_2885;
assign n_3095 =  x_4557 & ~n_2882;
assign n_3096 = ~n_3094 & ~n_3095;
assign n_3097 = ~n_3093 &  n_3096;
assign n_3098 =  x_4557 & ~n_3097;
assign n_3099 = ~x_4557 &  n_3097;
assign n_3100 = ~n_3098 & ~n_3099;
assign n_3101 =  x_4397 &  n_2883;
assign n_3102 =  i_5 &  n_2885;
assign n_3103 =  x_4556 & ~n_2882;
assign n_3104 = ~n_3102 & ~n_3103;
assign n_3105 = ~n_3101 &  n_3104;
assign n_3106 =  x_4556 & ~n_3105;
assign n_3107 = ~x_4556 &  n_3105;
assign n_3108 = ~n_3106 & ~n_3107;
assign n_3109 =  x_4396 &  n_2883;
assign n_3110 =  i_4 &  n_2885;
assign n_3111 =  x_4555 & ~n_2882;
assign n_3112 = ~n_3110 & ~n_3111;
assign n_3113 = ~n_3109 &  n_3112;
assign n_3114 =  x_4555 & ~n_3113;
assign n_3115 = ~x_4555 &  n_3113;
assign n_3116 = ~n_3114 & ~n_3115;
assign n_3117 =  x_4395 &  n_2883;
assign n_3118 =  i_3 &  n_2885;
assign n_3119 =  x_4554 & ~n_2882;
assign n_3120 = ~n_3118 & ~n_3119;
assign n_3121 = ~n_3117 &  n_3120;
assign n_3122 =  x_4554 & ~n_3121;
assign n_3123 = ~x_4554 &  n_3121;
assign n_3124 = ~n_3122 & ~n_3123;
assign n_3125 =  x_4394 &  n_2883;
assign n_3126 =  i_2 &  n_2885;
assign n_3127 =  x_4553 & ~n_2882;
assign n_3128 = ~n_3126 & ~n_3127;
assign n_3129 = ~n_3125 &  n_3128;
assign n_3130 =  x_4553 & ~n_3129;
assign n_3131 = ~x_4553 &  n_3129;
assign n_3132 = ~n_3130 & ~n_3131;
assign n_3133 =  x_4393 &  n_2883;
assign n_3134 =  i_1 &  n_2885;
assign n_3135 =  x_4552 & ~n_2882;
assign n_3136 = ~n_3134 & ~n_3135;
assign n_3137 = ~n_3133 &  n_3136;
assign n_3138 =  x_4552 & ~n_3137;
assign n_3139 = ~x_4552 &  n_3137;
assign n_3140 = ~n_3138 & ~n_3139;
assign n_3141 =  x_36 &  n_1897;
assign n_3142 =  n_759 &  n_7;
assign n_3143 =  x_41 &  n_349;
assign n_3144 =  n_3142 &  n_3143;
assign n_3145 =  n_3141 &  n_3144;
assign n_3146 =  x_4551 & ~n_3145;
assign n_3147 =  i_32 &  n_3145;
assign n_3148 = ~n_3146 & ~n_3147;
assign n_3149 =  x_4551 & ~n_3148;
assign n_3150 = ~x_4551 &  n_3148;
assign n_3151 = ~n_3149 & ~n_3150;
assign n_3152 =  x_4550 & ~n_3145;
assign n_3153 =  i_31 &  n_3145;
assign n_3154 = ~n_3152 & ~n_3153;
assign n_3155 =  x_4550 & ~n_3154;
assign n_3156 = ~x_4550 &  n_3154;
assign n_3157 = ~n_3155 & ~n_3156;
assign n_3158 =  x_4549 & ~n_3145;
assign n_3159 =  i_30 &  n_3145;
assign n_3160 = ~n_3158 & ~n_3159;
assign n_3161 =  x_4549 & ~n_3160;
assign n_3162 = ~x_4549 &  n_3160;
assign n_3163 = ~n_3161 & ~n_3162;
assign n_3164 =  x_4548 & ~n_3145;
assign n_3165 =  i_29 &  n_3145;
assign n_3166 = ~n_3164 & ~n_3165;
assign n_3167 =  x_4548 & ~n_3166;
assign n_3168 = ~x_4548 &  n_3166;
assign n_3169 = ~n_3167 & ~n_3168;
assign n_3170 =  x_4547 & ~n_3145;
assign n_3171 =  i_28 &  n_3145;
assign n_3172 = ~n_3170 & ~n_3171;
assign n_3173 =  x_4547 & ~n_3172;
assign n_3174 = ~x_4547 &  n_3172;
assign n_3175 = ~n_3173 & ~n_3174;
assign n_3176 =  x_4546 & ~n_3145;
assign n_3177 =  i_27 &  n_3145;
assign n_3178 = ~n_3176 & ~n_3177;
assign n_3179 =  x_4546 & ~n_3178;
assign n_3180 = ~x_4546 &  n_3178;
assign n_3181 = ~n_3179 & ~n_3180;
assign n_3182 =  x_4545 & ~n_3145;
assign n_3183 =  i_26 &  n_3145;
assign n_3184 = ~n_3182 & ~n_3183;
assign n_3185 =  x_4545 & ~n_3184;
assign n_3186 = ~x_4545 &  n_3184;
assign n_3187 = ~n_3185 & ~n_3186;
assign n_3188 =  x_4544 & ~n_3145;
assign n_3189 =  i_25 &  n_3145;
assign n_3190 = ~n_3188 & ~n_3189;
assign n_3191 =  x_4544 & ~n_3190;
assign n_3192 = ~x_4544 &  n_3190;
assign n_3193 = ~n_3191 & ~n_3192;
assign n_3194 =  x_4543 & ~n_3145;
assign n_3195 =  i_24 &  n_3145;
assign n_3196 = ~n_3194 & ~n_3195;
assign n_3197 =  x_4543 & ~n_3196;
assign n_3198 = ~x_4543 &  n_3196;
assign n_3199 = ~n_3197 & ~n_3198;
assign n_3200 =  x_4542 & ~n_3145;
assign n_3201 =  i_23 &  n_3145;
assign n_3202 = ~n_3200 & ~n_3201;
assign n_3203 =  x_4542 & ~n_3202;
assign n_3204 = ~x_4542 &  n_3202;
assign n_3205 = ~n_3203 & ~n_3204;
assign n_3206 =  x_4541 & ~n_3145;
assign n_3207 =  i_22 &  n_3145;
assign n_3208 = ~n_3206 & ~n_3207;
assign n_3209 =  x_4541 & ~n_3208;
assign n_3210 = ~x_4541 &  n_3208;
assign n_3211 = ~n_3209 & ~n_3210;
assign n_3212 =  x_4540 & ~n_3145;
assign n_3213 =  i_21 &  n_3145;
assign n_3214 = ~n_3212 & ~n_3213;
assign n_3215 =  x_4540 & ~n_3214;
assign n_3216 = ~x_4540 &  n_3214;
assign n_3217 = ~n_3215 & ~n_3216;
assign n_3218 =  x_4539 & ~n_3145;
assign n_3219 =  i_20 &  n_3145;
assign n_3220 = ~n_3218 & ~n_3219;
assign n_3221 =  x_4539 & ~n_3220;
assign n_3222 = ~x_4539 &  n_3220;
assign n_3223 = ~n_3221 & ~n_3222;
assign n_3224 =  x_4538 & ~n_3145;
assign n_3225 =  i_19 &  n_3145;
assign n_3226 = ~n_3224 & ~n_3225;
assign n_3227 =  x_4538 & ~n_3226;
assign n_3228 = ~x_4538 &  n_3226;
assign n_3229 = ~n_3227 & ~n_3228;
assign n_3230 =  x_4537 & ~n_3145;
assign n_3231 =  i_18 &  n_3145;
assign n_3232 = ~n_3230 & ~n_3231;
assign n_3233 =  x_4537 & ~n_3232;
assign n_3234 = ~x_4537 &  n_3232;
assign n_3235 = ~n_3233 & ~n_3234;
assign n_3236 =  x_4536 & ~n_3145;
assign n_3237 =  i_17 &  n_3145;
assign n_3238 = ~n_3236 & ~n_3237;
assign n_3239 =  x_4536 & ~n_3238;
assign n_3240 = ~x_4536 &  n_3238;
assign n_3241 = ~n_3239 & ~n_3240;
assign n_3242 =  x_4535 & ~n_3145;
assign n_3243 =  i_16 &  n_3145;
assign n_3244 = ~n_3242 & ~n_3243;
assign n_3245 =  x_4535 & ~n_3244;
assign n_3246 = ~x_4535 &  n_3244;
assign n_3247 = ~n_3245 & ~n_3246;
assign n_3248 =  x_4534 & ~n_3145;
assign n_3249 =  i_15 &  n_3145;
assign n_3250 = ~n_3248 & ~n_3249;
assign n_3251 =  x_4534 & ~n_3250;
assign n_3252 = ~x_4534 &  n_3250;
assign n_3253 = ~n_3251 & ~n_3252;
assign n_3254 =  x_4533 & ~n_3145;
assign n_3255 =  i_14 &  n_3145;
assign n_3256 = ~n_3254 & ~n_3255;
assign n_3257 =  x_4533 & ~n_3256;
assign n_3258 = ~x_4533 &  n_3256;
assign n_3259 = ~n_3257 & ~n_3258;
assign n_3260 =  x_4532 & ~n_3145;
assign n_3261 =  i_13 &  n_3145;
assign n_3262 = ~n_3260 & ~n_3261;
assign n_3263 =  x_4532 & ~n_3262;
assign n_3264 = ~x_4532 &  n_3262;
assign n_3265 = ~n_3263 & ~n_3264;
assign n_3266 =  x_4531 & ~n_3145;
assign n_3267 =  i_12 &  n_3145;
assign n_3268 = ~n_3266 & ~n_3267;
assign n_3269 =  x_4531 & ~n_3268;
assign n_3270 = ~x_4531 &  n_3268;
assign n_3271 = ~n_3269 & ~n_3270;
assign n_3272 =  x_4530 & ~n_3145;
assign n_3273 =  i_11 &  n_3145;
assign n_3274 = ~n_3272 & ~n_3273;
assign n_3275 =  x_4530 & ~n_3274;
assign n_3276 = ~x_4530 &  n_3274;
assign n_3277 = ~n_3275 & ~n_3276;
assign n_3278 =  x_4529 & ~n_3145;
assign n_3279 =  i_10 &  n_3145;
assign n_3280 = ~n_3278 & ~n_3279;
assign n_3281 =  x_4529 & ~n_3280;
assign n_3282 = ~x_4529 &  n_3280;
assign n_3283 = ~n_3281 & ~n_3282;
assign n_3284 =  x_4528 & ~n_3145;
assign n_3285 =  i_9 &  n_3145;
assign n_3286 = ~n_3284 & ~n_3285;
assign n_3287 =  x_4528 & ~n_3286;
assign n_3288 = ~x_4528 &  n_3286;
assign n_3289 = ~n_3287 & ~n_3288;
assign n_3290 =  x_4527 & ~n_3145;
assign n_3291 =  i_8 &  n_3145;
assign n_3292 = ~n_3290 & ~n_3291;
assign n_3293 =  x_4527 & ~n_3292;
assign n_3294 = ~x_4527 &  n_3292;
assign n_3295 = ~n_3293 & ~n_3294;
assign n_3296 =  x_4526 & ~n_3145;
assign n_3297 =  i_7 &  n_3145;
assign n_3298 = ~n_3296 & ~n_3297;
assign n_3299 =  x_4526 & ~n_3298;
assign n_3300 = ~x_4526 &  n_3298;
assign n_3301 = ~n_3299 & ~n_3300;
assign n_3302 =  x_4525 & ~n_3145;
assign n_3303 =  i_6 &  n_3145;
assign n_3304 = ~n_3302 & ~n_3303;
assign n_3305 =  x_4525 & ~n_3304;
assign n_3306 = ~x_4525 &  n_3304;
assign n_3307 = ~n_3305 & ~n_3306;
assign n_3308 =  x_4524 & ~n_3145;
assign n_3309 =  i_5 &  n_3145;
assign n_3310 = ~n_3308 & ~n_3309;
assign n_3311 =  x_4524 & ~n_3310;
assign n_3312 = ~x_4524 &  n_3310;
assign n_3313 = ~n_3311 & ~n_3312;
assign n_3314 =  x_4523 & ~n_3145;
assign n_3315 =  i_4 &  n_3145;
assign n_3316 = ~n_3314 & ~n_3315;
assign n_3317 =  x_4523 & ~n_3316;
assign n_3318 = ~x_4523 &  n_3316;
assign n_3319 = ~n_3317 & ~n_3318;
assign n_3320 =  x_4522 & ~n_3145;
assign n_3321 =  i_3 &  n_3145;
assign n_3322 = ~n_3320 & ~n_3321;
assign n_3323 =  x_4522 & ~n_3322;
assign n_3324 = ~x_4522 &  n_3322;
assign n_3325 = ~n_3323 & ~n_3324;
assign n_3326 =  x_4521 & ~n_3145;
assign n_3327 =  i_2 &  n_3145;
assign n_3328 = ~n_3326 & ~n_3327;
assign n_3329 =  x_4521 & ~n_3328;
assign n_3330 = ~x_4521 &  n_3328;
assign n_3331 = ~n_3329 & ~n_3330;
assign n_3332 =  x_4520 & ~n_3145;
assign n_3333 =  i_1 &  n_3145;
assign n_3334 = ~n_3332 & ~n_3333;
assign n_3335 =  x_4520 & ~n_3334;
assign n_3336 = ~x_4520 &  n_3334;
assign n_3337 = ~n_3335 & ~n_3336;
assign n_3338 =  x_41 &  n_6;
assign n_3339 =  n_1037 &  n_3338;
assign n_3340 =  n_3339 &  n_2685;
assign n_3341 = ~x_41 &  x_42;
assign n_3342 =  n_3141 &  n_8;
assign n_3343 =  n_3341 &  n_3342;
assign n_3344 = ~x_43 &  n_3343;
assign n_3345 = ~n_3340 & ~n_3344;
assign n_3346 =  n_1174 &  n_2685;
assign n_3347 =  n_2 &  n_3346;
assign n_3348 =  n_553 &  n_3342;
assign n_3349 = ~x_43 &  n_3348;
assign n_3350 = ~n_3347 & ~n_3349;
assign n_3351 =  x_4519 &  n_3350;
assign n_3352 =  n_3345 & ~n_3351;
assign n_3353 =  x_4519 & ~n_3352;
assign n_3354 = ~x_4519 &  n_3352;
assign n_3355 = ~n_3353 & ~n_3354;
assign n_3356 =  n_3345 &  n_3350;
assign n_3357 =  x_4518 &  n_3356;
assign n_3358 =  x_4518 &  n_3357;
assign n_3359 = ~x_4518 & ~n_3357;
assign n_3360 = ~n_3358 & ~n_3359;
assign n_3361 =  x_4517 &  n_3356;
assign n_3362 =  x_4517 &  n_3361;
assign n_3363 = ~x_4517 & ~n_3361;
assign n_3364 = ~n_3362 & ~n_3363;
assign n_3365 =  x_4516 &  n_3356;
assign n_3366 =  x_4516 &  n_3365;
assign n_3367 = ~x_4516 & ~n_3365;
assign n_3368 = ~n_3366 & ~n_3367;
assign n_3369 =  x_4515 &  n_3356;
assign n_3370 =  x_4515 &  n_3369;
assign n_3371 = ~x_4515 & ~n_3369;
assign n_3372 = ~n_3370 & ~n_3371;
assign n_3373 =  x_4514 &  n_3356;
assign n_3374 =  x_4514 &  n_3373;
assign n_3375 = ~x_4514 & ~n_3373;
assign n_3376 = ~n_3374 & ~n_3375;
assign n_3377 =  x_4513 &  n_3356;
assign n_3378 =  x_4513 &  n_3377;
assign n_3379 = ~x_4513 & ~n_3377;
assign n_3380 = ~n_3378 & ~n_3379;
assign n_3381 =  x_4512 &  n_3356;
assign n_3382 =  x_4512 &  n_3381;
assign n_3383 = ~x_4512 & ~n_3381;
assign n_3384 = ~n_3382 & ~n_3383;
assign n_3385 =  x_4511 &  n_3356;
assign n_3386 =  x_4511 &  n_3385;
assign n_3387 = ~x_4511 & ~n_3385;
assign n_3388 = ~n_3386 & ~n_3387;
assign n_3389 =  x_4510 &  n_3356;
assign n_3390 =  x_4510 &  n_3389;
assign n_3391 = ~x_4510 & ~n_3389;
assign n_3392 = ~n_3390 & ~n_3391;
assign n_3393 =  x_4509 &  n_3356;
assign n_3394 =  x_4509 &  n_3393;
assign n_3395 = ~x_4509 & ~n_3393;
assign n_3396 = ~n_3394 & ~n_3395;
assign n_3397 =  x_4508 &  n_3356;
assign n_3398 =  x_4508 &  n_3397;
assign n_3399 = ~x_4508 & ~n_3397;
assign n_3400 = ~n_3398 & ~n_3399;
assign n_3401 =  x_4507 &  n_3356;
assign n_3402 =  x_4507 &  n_3401;
assign n_3403 = ~x_4507 & ~n_3401;
assign n_3404 = ~n_3402 & ~n_3403;
assign n_3405 =  x_4506 &  n_3356;
assign n_3406 =  x_4506 &  n_3405;
assign n_3407 = ~x_4506 & ~n_3405;
assign n_3408 = ~n_3406 & ~n_3407;
assign n_3409 =  x_4505 &  n_3356;
assign n_3410 =  x_4505 &  n_3409;
assign n_3411 = ~x_4505 & ~n_3409;
assign n_3412 = ~n_3410 & ~n_3411;
assign n_3413 =  x_4504 &  n_3356;
assign n_3414 =  x_4504 &  n_3413;
assign n_3415 = ~x_4504 & ~n_3413;
assign n_3416 = ~n_3414 & ~n_3415;
assign n_3417 =  x_4503 &  n_3356;
assign n_3418 =  x_4503 &  n_3417;
assign n_3419 = ~x_4503 & ~n_3417;
assign n_3420 = ~n_3418 & ~n_3419;
assign n_3421 =  x_4502 &  n_3356;
assign n_3422 =  x_4502 &  n_3421;
assign n_3423 = ~x_4502 & ~n_3421;
assign n_3424 = ~n_3422 & ~n_3423;
assign n_3425 =  x_4501 &  n_3356;
assign n_3426 =  x_4501 &  n_3425;
assign n_3427 = ~x_4501 & ~n_3425;
assign n_3428 = ~n_3426 & ~n_3427;
assign n_3429 =  x_4500 &  n_3356;
assign n_3430 =  x_4500 &  n_3429;
assign n_3431 = ~x_4500 & ~n_3429;
assign n_3432 = ~n_3430 & ~n_3431;
assign n_3433 =  x_4499 &  n_3356;
assign n_3434 =  x_4499 &  n_3433;
assign n_3435 = ~x_4499 & ~n_3433;
assign n_3436 = ~n_3434 & ~n_3435;
assign n_3437 =  x_4498 &  n_3356;
assign n_3438 =  x_4498 &  n_3437;
assign n_3439 = ~x_4498 & ~n_3437;
assign n_3440 = ~n_3438 & ~n_3439;
assign n_3441 =  x_4497 &  n_3356;
assign n_3442 =  x_4497 &  n_3441;
assign n_3443 = ~x_4497 & ~n_3441;
assign n_3444 = ~n_3442 & ~n_3443;
assign n_3445 =  x_4496 &  n_3356;
assign n_3446 =  x_4496 &  n_3445;
assign n_3447 = ~x_4496 & ~n_3445;
assign n_3448 = ~n_3446 & ~n_3447;
assign n_3449 =  x_4495 &  n_3356;
assign n_3450 =  x_4495 &  n_3449;
assign n_3451 = ~x_4495 & ~n_3449;
assign n_3452 = ~n_3450 & ~n_3451;
assign n_3453 =  x_4494 &  n_3356;
assign n_3454 =  x_4494 &  n_3453;
assign n_3455 = ~x_4494 & ~n_3453;
assign n_3456 = ~n_3454 & ~n_3455;
assign n_3457 =  x_4493 &  n_3356;
assign n_3458 =  x_4493 &  n_3457;
assign n_3459 = ~x_4493 & ~n_3457;
assign n_3460 = ~n_3458 & ~n_3459;
assign n_3461 =  x_4492 &  n_3356;
assign n_3462 =  x_4492 &  n_3461;
assign n_3463 = ~x_4492 & ~n_3461;
assign n_3464 = ~n_3462 & ~n_3463;
assign n_3465 =  x_4491 &  n_3356;
assign n_3466 =  x_4491 &  n_3465;
assign n_3467 = ~x_4491 & ~n_3465;
assign n_3468 = ~n_3466 & ~n_3467;
assign n_3469 =  x_4490 &  n_3356;
assign n_3470 =  x_4490 &  n_3469;
assign n_3471 = ~x_4490 & ~n_3469;
assign n_3472 = ~n_3470 & ~n_3471;
assign n_3473 =  x_4489 &  n_3356;
assign n_3474 =  x_4489 &  n_3473;
assign n_3475 = ~x_4489 & ~n_3473;
assign n_3476 = ~n_3474 & ~n_3475;
assign n_3477 =  x_4488 &  n_3356;
assign n_3478 =  x_4488 &  n_3477;
assign n_3479 = ~x_4488 & ~n_3477;
assign n_3480 = ~n_3478 & ~n_3479;
assign n_3481 =  x_4487 & ~n_900;
assign n_3482 = ~n_761 & ~n_3481;
assign n_3483 =  x_4487 & ~n_3482;
assign n_3484 = ~x_4487 &  n_3482;
assign n_3485 = ~n_3483 & ~n_3484;
assign n_3486 =  x_4486 & ~n_900;
assign n_3487 =  x_4486 &  n_3486;
assign n_3488 = ~x_4486 & ~n_3486;
assign n_3489 = ~n_3487 & ~n_3488;
assign n_3490 =  x_4485 & ~n_900;
assign n_3491 =  x_4485 &  n_3490;
assign n_3492 = ~x_4485 & ~n_3490;
assign n_3493 = ~n_3491 & ~n_3492;
assign n_3494 =  x_4484 & ~n_900;
assign n_3495 =  x_4484 &  n_3494;
assign n_3496 = ~x_4484 & ~n_3494;
assign n_3497 = ~n_3495 & ~n_3496;
assign n_3498 =  x_4483 & ~n_900;
assign n_3499 = ~n_761 & ~n_3498;
assign n_3500 =  x_4483 & ~n_3499;
assign n_3501 = ~x_4483 &  n_3499;
assign n_3502 = ~n_3500 & ~n_3501;
assign n_3503 =  x_4482 & ~n_900;
assign n_3504 = ~n_761 & ~n_3503;
assign n_3505 =  x_4482 & ~n_3504;
assign n_3506 = ~x_4482 &  n_3504;
assign n_3507 = ~n_3505 & ~n_3506;
assign n_3508 =  x_4481 & ~n_900;
assign n_3509 = ~n_761 & ~n_3508;
assign n_3510 =  x_4481 & ~n_3509;
assign n_3511 = ~x_4481 &  n_3509;
assign n_3512 = ~n_3510 & ~n_3511;
assign n_3513 =  x_4480 & ~n_900;
assign n_3514 =  x_4480 &  n_3513;
assign n_3515 = ~x_4480 & ~n_3513;
assign n_3516 = ~n_3514 & ~n_3515;
assign n_3517 =  x_4479 & ~n_900;
assign n_3518 = ~n_761 & ~n_3517;
assign n_3519 =  x_4479 & ~n_3518;
assign n_3520 = ~x_4479 &  n_3518;
assign n_3521 = ~n_3519 & ~n_3520;
assign n_3522 =  x_4478 & ~n_900;
assign n_3523 =  x_4478 &  n_3522;
assign n_3524 = ~x_4478 & ~n_3522;
assign n_3525 = ~n_3523 & ~n_3524;
assign n_3526 =  x_4477 & ~n_900;
assign n_3527 = ~n_761 & ~n_3526;
assign n_3528 =  x_4477 & ~n_3527;
assign n_3529 = ~x_4477 &  n_3527;
assign n_3530 = ~n_3528 & ~n_3529;
assign n_3531 =  x_4476 & ~n_900;
assign n_3532 =  x_4476 &  n_3531;
assign n_3533 = ~x_4476 & ~n_3531;
assign n_3534 = ~n_3532 & ~n_3533;
assign n_3535 =  x_4475 & ~n_900;
assign n_3536 =  x_4475 &  n_3535;
assign n_3537 = ~x_4475 & ~n_3535;
assign n_3538 = ~n_3536 & ~n_3537;
assign n_3539 =  x_4474 & ~n_900;
assign n_3540 =  x_4474 &  n_3539;
assign n_3541 = ~x_4474 & ~n_3539;
assign n_3542 = ~n_3540 & ~n_3541;
assign n_3543 =  x_4473 & ~n_900;
assign n_3544 =  x_4473 &  n_3543;
assign n_3545 = ~x_4473 & ~n_3543;
assign n_3546 = ~n_3544 & ~n_3545;
assign n_3547 =  x_4472 & ~n_900;
assign n_3548 =  x_4472 &  n_3547;
assign n_3549 = ~x_4472 & ~n_3547;
assign n_3550 = ~n_3548 & ~n_3549;
assign n_3551 =  x_4471 & ~n_900;
assign n_3552 =  x_4471 &  n_3551;
assign n_3553 = ~x_4471 & ~n_3551;
assign n_3554 = ~n_3552 & ~n_3553;
assign n_3555 =  x_4470 & ~n_900;
assign n_3556 =  x_4470 &  n_3555;
assign n_3557 = ~x_4470 & ~n_3555;
assign n_3558 = ~n_3556 & ~n_3557;
assign n_3559 =  x_4469 & ~n_900;
assign n_3560 =  x_4469 &  n_3559;
assign n_3561 = ~x_4469 & ~n_3559;
assign n_3562 = ~n_3560 & ~n_3561;
assign n_3563 =  x_4468 & ~n_900;
assign n_3564 =  x_4468 &  n_3563;
assign n_3565 = ~x_4468 & ~n_3563;
assign n_3566 = ~n_3564 & ~n_3565;
assign n_3567 =  x_4467 & ~n_900;
assign n_3568 =  x_4467 &  n_3567;
assign n_3569 = ~x_4467 & ~n_3567;
assign n_3570 = ~n_3568 & ~n_3569;
assign n_3571 =  x_4466 & ~n_900;
assign n_3572 =  x_4466 &  n_3571;
assign n_3573 = ~x_4466 & ~n_3571;
assign n_3574 = ~n_3572 & ~n_3573;
assign n_3575 =  x_4465 & ~n_900;
assign n_3576 =  x_4465 &  n_3575;
assign n_3577 = ~x_4465 & ~n_3575;
assign n_3578 = ~n_3576 & ~n_3577;
assign n_3579 =  x_4464 & ~n_900;
assign n_3580 =  x_4464 &  n_3579;
assign n_3581 = ~x_4464 & ~n_3579;
assign n_3582 = ~n_3580 & ~n_3581;
assign n_3583 =  x_4463 & ~n_900;
assign n_3584 =  x_4463 &  n_3583;
assign n_3585 = ~x_4463 & ~n_3583;
assign n_3586 = ~n_3584 & ~n_3585;
assign n_3587 =  x_4462 & ~n_900;
assign n_3588 =  x_4462 &  n_3587;
assign n_3589 = ~x_4462 & ~n_3587;
assign n_3590 = ~n_3588 & ~n_3589;
assign n_3591 =  x_4461 & ~n_900;
assign n_3592 =  x_4461 &  n_3591;
assign n_3593 = ~x_4461 & ~n_3591;
assign n_3594 = ~n_3592 & ~n_3593;
assign n_3595 =  x_4460 & ~n_900;
assign n_3596 =  x_4460 &  n_3595;
assign n_3597 = ~x_4460 & ~n_3595;
assign n_3598 = ~n_3596 & ~n_3597;
assign n_3599 =  x_4459 & ~n_900;
assign n_3600 =  x_4459 &  n_3599;
assign n_3601 = ~x_4459 & ~n_3599;
assign n_3602 = ~n_3600 & ~n_3601;
assign n_3603 =  x_4458 & ~n_900;
assign n_3604 =  x_4458 &  n_3603;
assign n_3605 = ~x_4458 & ~n_3603;
assign n_3606 = ~n_3604 & ~n_3605;
assign n_3607 =  x_4457 & ~n_900;
assign n_3608 =  x_4457 &  n_3607;
assign n_3609 = ~x_4457 & ~n_3607;
assign n_3610 = ~n_3608 & ~n_3609;
assign n_3611 =  x_4456 & ~n_900;
assign n_3612 =  x_4456 &  n_3611;
assign n_3613 = ~x_4456 & ~n_3611;
assign n_3614 = ~n_3612 & ~n_3613;
assign n_3615 = ~x_37 &  n_354;
assign n_3616 =  n_556 &  n_3615;
assign n_3617 = ~x_40 &  n_3616;
assign n_3618 =  n_3143 &  n_3617;
assign n_3619 =  n_556 &  n_355;
assign n_3620 =  x_40 &  n_3619;
assign n_3621 =  n_3143 &  n_3620;
assign n_3622 = ~n_3618 & ~n_3621;
assign n_3623 =  n_1305 &  n_2;
assign n_3624 =  n_3623 &  n_1306;
assign n_3625 =  n_759 &  n_2;
assign n_3626 =  n_3625 &  n_1698;
assign n_3627 = ~n_3624 & ~n_3626;
assign n_3628 =  n_759 &  n_2879;
assign n_3629 =  n_765 &  n_3628;
assign n_3630 =  n_152 &  n_3629;
assign n_3631 = ~x_43 &  n_3630;
assign n_3632 =  n_553 &  n_765;
assign n_3633 =  n_3628 &  n_3632;
assign n_3634 =  n_2 &  n_2881;
assign n_3635 = ~n_3633 & ~n_3634;
assign n_3636 = ~n_3631 &  n_3635;
assign n_3637 =  n_3627 &  n_3636;
assign n_3638 =  n_3622 &  n_3637;
assign n_3639 =  x_4424 &  n_3638;
assign n_3640 = ~n_3618 &  n_3635;
assign n_3641 =  i_32 & ~n_3640;
assign n_3642 =  x_3703 &  n_3621;
assign n_3643 =  x_2682 &  n_3631;
assign n_3644 =  x_3799 &  n_3626;
assign n_3645 =  x_2714 &  n_3624;
assign n_3646 = ~n_3644 & ~n_3645;
assign n_3647 = ~n_3643 &  n_3646;
assign n_3648 = ~n_3642 &  n_3647;
assign n_3649 = ~n_3641 &  n_3648;
assign n_3650 = ~n_3639 &  n_3649;
assign n_3651 =  x_4424 & ~n_3650;
assign n_3652 = ~x_4424 &  n_3650;
assign n_3653 = ~n_3651 & ~n_3652;
assign n_3654 =  x_4423 &  n_3638;
assign n_3655 =  i_31 & ~n_3640;
assign n_3656 =  x_3702 &  n_3621;
assign n_3657 =  x_2681 &  n_3631;
assign n_3658 =  x_3798 &  n_3626;
assign n_3659 =  x_2713 &  n_3624;
assign n_3660 = ~n_3658 & ~n_3659;
assign n_3661 = ~n_3657 &  n_3660;
assign n_3662 = ~n_3656 &  n_3661;
assign n_3663 = ~n_3655 &  n_3662;
assign n_3664 = ~n_3654 &  n_3663;
assign n_3665 =  x_4423 & ~n_3664;
assign n_3666 = ~x_4423 &  n_3664;
assign n_3667 = ~n_3665 & ~n_3666;
assign n_3668 =  x_4422 &  n_3638;
assign n_3669 =  i_30 & ~n_3640;
assign n_3670 =  x_3701 &  n_3621;
assign n_3671 =  x_2680 &  n_3631;
assign n_3672 =  x_3797 &  n_3626;
assign n_3673 =  x_2712 &  n_3624;
assign n_3674 = ~n_3672 & ~n_3673;
assign n_3675 = ~n_3671 &  n_3674;
assign n_3676 = ~n_3670 &  n_3675;
assign n_3677 = ~n_3669 &  n_3676;
assign n_3678 = ~n_3668 &  n_3677;
assign n_3679 =  x_4422 & ~n_3678;
assign n_3680 = ~x_4422 &  n_3678;
assign n_3681 = ~n_3679 & ~n_3680;
assign n_3682 =  x_4421 &  n_3638;
assign n_3683 =  i_29 & ~n_3640;
assign n_3684 =  x_3700 &  n_3621;
assign n_3685 =  x_2679 &  n_3631;
assign n_3686 =  x_3796 &  n_3626;
assign n_3687 =  x_2711 &  n_3624;
assign n_3688 = ~n_3686 & ~n_3687;
assign n_3689 = ~n_3685 &  n_3688;
assign n_3690 = ~n_3684 &  n_3689;
assign n_3691 = ~n_3683 &  n_3690;
assign n_3692 = ~n_3682 &  n_3691;
assign n_3693 =  x_4421 & ~n_3692;
assign n_3694 = ~x_4421 &  n_3692;
assign n_3695 = ~n_3693 & ~n_3694;
assign n_3696 =  x_4420 &  n_3638;
assign n_3697 =  i_28 & ~n_3640;
assign n_3698 =  x_3699 &  n_3621;
assign n_3699 =  x_2678 &  n_3631;
assign n_3700 =  x_3795 &  n_3626;
assign n_3701 =  x_2710 &  n_3624;
assign n_3702 = ~n_3700 & ~n_3701;
assign n_3703 = ~n_3699 &  n_3702;
assign n_3704 = ~n_3698 &  n_3703;
assign n_3705 = ~n_3697 &  n_3704;
assign n_3706 = ~n_3696 &  n_3705;
assign n_3707 =  x_4420 & ~n_3706;
assign n_3708 = ~x_4420 &  n_3706;
assign n_3709 = ~n_3707 & ~n_3708;
assign n_3710 =  x_4419 &  n_3638;
assign n_3711 =  i_27 & ~n_3640;
assign n_3712 =  x_3698 &  n_3621;
assign n_3713 =  x_2677 &  n_3631;
assign n_3714 =  x_3794 &  n_3626;
assign n_3715 =  x_2709 &  n_3624;
assign n_3716 = ~n_3714 & ~n_3715;
assign n_3717 = ~n_3713 &  n_3716;
assign n_3718 = ~n_3712 &  n_3717;
assign n_3719 = ~n_3711 &  n_3718;
assign n_3720 = ~n_3710 &  n_3719;
assign n_3721 =  x_4419 & ~n_3720;
assign n_3722 = ~x_4419 &  n_3720;
assign n_3723 = ~n_3721 & ~n_3722;
assign n_3724 =  x_4418 &  n_3638;
assign n_3725 =  i_26 & ~n_3640;
assign n_3726 =  x_3697 &  n_3621;
assign n_3727 =  x_2676 &  n_3631;
assign n_3728 =  x_3793 &  n_3626;
assign n_3729 =  x_2708 &  n_3624;
assign n_3730 = ~n_3728 & ~n_3729;
assign n_3731 = ~n_3727 &  n_3730;
assign n_3732 = ~n_3726 &  n_3731;
assign n_3733 = ~n_3725 &  n_3732;
assign n_3734 = ~n_3724 &  n_3733;
assign n_3735 =  x_4418 & ~n_3734;
assign n_3736 = ~x_4418 &  n_3734;
assign n_3737 = ~n_3735 & ~n_3736;
assign n_3738 =  x_4417 &  n_3638;
assign n_3739 =  i_25 & ~n_3640;
assign n_3740 =  x_3696 &  n_3621;
assign n_3741 =  x_2675 &  n_3631;
assign n_3742 =  x_3792 &  n_3626;
assign n_3743 =  x_2707 &  n_3624;
assign n_3744 = ~n_3742 & ~n_3743;
assign n_3745 = ~n_3741 &  n_3744;
assign n_3746 = ~n_3740 &  n_3745;
assign n_3747 = ~n_3739 &  n_3746;
assign n_3748 = ~n_3738 &  n_3747;
assign n_3749 =  x_4417 & ~n_3748;
assign n_3750 = ~x_4417 &  n_3748;
assign n_3751 = ~n_3749 & ~n_3750;
assign n_3752 =  x_4416 &  n_3638;
assign n_3753 =  i_24 & ~n_3640;
assign n_3754 =  x_3695 &  n_3621;
assign n_3755 =  x_2674 &  n_3631;
assign n_3756 =  x_3791 &  n_3626;
assign n_3757 =  x_2706 &  n_3624;
assign n_3758 = ~n_3756 & ~n_3757;
assign n_3759 = ~n_3755 &  n_3758;
assign n_3760 = ~n_3754 &  n_3759;
assign n_3761 = ~n_3753 &  n_3760;
assign n_3762 = ~n_3752 &  n_3761;
assign n_3763 =  x_4416 & ~n_3762;
assign n_3764 = ~x_4416 &  n_3762;
assign n_3765 = ~n_3763 & ~n_3764;
assign n_3766 =  x_4415 &  n_3638;
assign n_3767 =  i_23 & ~n_3640;
assign n_3768 =  x_3694 &  n_3621;
assign n_3769 =  x_2673 &  n_3631;
assign n_3770 =  x_3790 &  n_3626;
assign n_3771 =  x_2705 &  n_3624;
assign n_3772 = ~n_3770 & ~n_3771;
assign n_3773 = ~n_3769 &  n_3772;
assign n_3774 = ~n_3768 &  n_3773;
assign n_3775 = ~n_3767 &  n_3774;
assign n_3776 = ~n_3766 &  n_3775;
assign n_3777 =  x_4415 & ~n_3776;
assign n_3778 = ~x_4415 &  n_3776;
assign n_3779 = ~n_3777 & ~n_3778;
assign n_3780 =  x_4414 &  n_3638;
assign n_3781 =  i_22 & ~n_3640;
assign n_3782 =  x_3693 &  n_3621;
assign n_3783 =  x_2672 &  n_3631;
assign n_3784 =  x_3789 &  n_3626;
assign n_3785 =  x_2704 &  n_3624;
assign n_3786 = ~n_3784 & ~n_3785;
assign n_3787 = ~n_3783 &  n_3786;
assign n_3788 = ~n_3782 &  n_3787;
assign n_3789 = ~n_3781 &  n_3788;
assign n_3790 = ~n_3780 &  n_3789;
assign n_3791 =  x_4414 & ~n_3790;
assign n_3792 = ~x_4414 &  n_3790;
assign n_3793 = ~n_3791 & ~n_3792;
assign n_3794 =  x_4413 &  n_3638;
assign n_3795 =  i_21 & ~n_3640;
assign n_3796 =  x_3692 &  n_3621;
assign n_3797 =  x_2671 &  n_3631;
assign n_3798 =  x_3788 &  n_3626;
assign n_3799 =  x_2703 &  n_3624;
assign n_3800 = ~n_3798 & ~n_3799;
assign n_3801 = ~n_3797 &  n_3800;
assign n_3802 = ~n_3796 &  n_3801;
assign n_3803 = ~n_3795 &  n_3802;
assign n_3804 = ~n_3794 &  n_3803;
assign n_3805 =  x_4413 & ~n_3804;
assign n_3806 = ~x_4413 &  n_3804;
assign n_3807 = ~n_3805 & ~n_3806;
assign n_3808 =  x_4412 &  n_3638;
assign n_3809 =  i_20 & ~n_3640;
assign n_3810 =  x_3691 &  n_3621;
assign n_3811 =  x_2670 &  n_3631;
assign n_3812 =  x_3787 &  n_3626;
assign n_3813 =  x_2702 &  n_3624;
assign n_3814 = ~n_3812 & ~n_3813;
assign n_3815 = ~n_3811 &  n_3814;
assign n_3816 = ~n_3810 &  n_3815;
assign n_3817 = ~n_3809 &  n_3816;
assign n_3818 = ~n_3808 &  n_3817;
assign n_3819 =  x_4412 & ~n_3818;
assign n_3820 = ~x_4412 &  n_3818;
assign n_3821 = ~n_3819 & ~n_3820;
assign n_3822 =  x_4411 &  n_3638;
assign n_3823 =  i_19 & ~n_3640;
assign n_3824 =  x_3690 &  n_3621;
assign n_3825 =  x_2669 &  n_3631;
assign n_3826 =  x_3786 &  n_3626;
assign n_3827 =  x_2701 &  n_3624;
assign n_3828 = ~n_3826 & ~n_3827;
assign n_3829 = ~n_3825 &  n_3828;
assign n_3830 = ~n_3824 &  n_3829;
assign n_3831 = ~n_3823 &  n_3830;
assign n_3832 = ~n_3822 &  n_3831;
assign n_3833 =  x_4411 & ~n_3832;
assign n_3834 = ~x_4411 &  n_3832;
assign n_3835 = ~n_3833 & ~n_3834;
assign n_3836 =  x_4410 &  n_3638;
assign n_3837 =  i_18 & ~n_3640;
assign n_3838 =  x_3689 &  n_3621;
assign n_3839 =  x_2668 &  n_3631;
assign n_3840 =  x_3785 &  n_3626;
assign n_3841 =  x_2700 &  n_3624;
assign n_3842 = ~n_3840 & ~n_3841;
assign n_3843 = ~n_3839 &  n_3842;
assign n_3844 = ~n_3838 &  n_3843;
assign n_3845 = ~n_3837 &  n_3844;
assign n_3846 = ~n_3836 &  n_3845;
assign n_3847 =  x_4410 & ~n_3846;
assign n_3848 = ~x_4410 &  n_3846;
assign n_3849 = ~n_3847 & ~n_3848;
assign n_3850 =  x_4409 &  n_3638;
assign n_3851 =  i_17 & ~n_3640;
assign n_3852 =  x_3688 &  n_3621;
assign n_3853 =  x_2667 &  n_3631;
assign n_3854 =  x_3784 &  n_3626;
assign n_3855 =  x_2699 &  n_3624;
assign n_3856 = ~n_3854 & ~n_3855;
assign n_3857 = ~n_3853 &  n_3856;
assign n_3858 = ~n_3852 &  n_3857;
assign n_3859 = ~n_3851 &  n_3858;
assign n_3860 = ~n_3850 &  n_3859;
assign n_3861 =  x_4409 & ~n_3860;
assign n_3862 = ~x_4409 &  n_3860;
assign n_3863 = ~n_3861 & ~n_3862;
assign n_3864 =  x_4408 &  n_3638;
assign n_3865 =  i_16 & ~n_3640;
assign n_3866 =  x_3687 &  n_3621;
assign n_3867 =  x_2666 &  n_3631;
assign n_3868 =  x_3783 &  n_3626;
assign n_3869 =  x_2698 &  n_3624;
assign n_3870 = ~n_3868 & ~n_3869;
assign n_3871 = ~n_3867 &  n_3870;
assign n_3872 = ~n_3866 &  n_3871;
assign n_3873 = ~n_3865 &  n_3872;
assign n_3874 = ~n_3864 &  n_3873;
assign n_3875 =  x_4408 & ~n_3874;
assign n_3876 = ~x_4408 &  n_3874;
assign n_3877 = ~n_3875 & ~n_3876;
assign n_3878 =  x_4407 &  n_3638;
assign n_3879 =  i_15 & ~n_3640;
assign n_3880 =  x_3686 &  n_3621;
assign n_3881 =  x_2665 &  n_3631;
assign n_3882 =  x_3782 &  n_3626;
assign n_3883 =  x_2697 &  n_3624;
assign n_3884 = ~n_3882 & ~n_3883;
assign n_3885 = ~n_3881 &  n_3884;
assign n_3886 = ~n_3880 &  n_3885;
assign n_3887 = ~n_3879 &  n_3886;
assign n_3888 = ~n_3878 &  n_3887;
assign n_3889 =  x_4407 & ~n_3888;
assign n_3890 = ~x_4407 &  n_3888;
assign n_3891 = ~n_3889 & ~n_3890;
assign n_3892 =  x_4406 &  n_3638;
assign n_3893 =  i_14 & ~n_3640;
assign n_3894 =  x_3685 &  n_3621;
assign n_3895 =  x_2664 &  n_3631;
assign n_3896 =  x_3781 &  n_3626;
assign n_3897 =  x_2696 &  n_3624;
assign n_3898 = ~n_3896 & ~n_3897;
assign n_3899 = ~n_3895 &  n_3898;
assign n_3900 = ~n_3894 &  n_3899;
assign n_3901 = ~n_3893 &  n_3900;
assign n_3902 = ~n_3892 &  n_3901;
assign n_3903 =  x_4406 & ~n_3902;
assign n_3904 = ~x_4406 &  n_3902;
assign n_3905 = ~n_3903 & ~n_3904;
assign n_3906 =  x_4405 &  n_3638;
assign n_3907 =  i_13 & ~n_3640;
assign n_3908 =  x_3684 &  n_3621;
assign n_3909 =  x_2663 &  n_3631;
assign n_3910 =  x_3780 &  n_3626;
assign n_3911 =  x_2695 &  n_3624;
assign n_3912 = ~n_3910 & ~n_3911;
assign n_3913 = ~n_3909 &  n_3912;
assign n_3914 = ~n_3908 &  n_3913;
assign n_3915 = ~n_3907 &  n_3914;
assign n_3916 = ~n_3906 &  n_3915;
assign n_3917 =  x_4405 & ~n_3916;
assign n_3918 = ~x_4405 &  n_3916;
assign n_3919 = ~n_3917 & ~n_3918;
assign n_3920 =  x_4404 &  n_3638;
assign n_3921 =  i_12 & ~n_3640;
assign n_3922 =  x_3683 &  n_3621;
assign n_3923 =  x_2662 &  n_3631;
assign n_3924 =  x_3779 &  n_3626;
assign n_3925 =  x_2694 &  n_3624;
assign n_3926 = ~n_3924 & ~n_3925;
assign n_3927 = ~n_3923 &  n_3926;
assign n_3928 = ~n_3922 &  n_3927;
assign n_3929 = ~n_3921 &  n_3928;
assign n_3930 = ~n_3920 &  n_3929;
assign n_3931 =  x_4404 & ~n_3930;
assign n_3932 = ~x_4404 &  n_3930;
assign n_3933 = ~n_3931 & ~n_3932;
assign n_3934 =  x_4403 &  n_3638;
assign n_3935 =  i_11 & ~n_3640;
assign n_3936 =  x_3682 &  n_3621;
assign n_3937 =  x_2661 &  n_3631;
assign n_3938 =  x_3778 &  n_3626;
assign n_3939 =  x_2693 &  n_3624;
assign n_3940 = ~n_3938 & ~n_3939;
assign n_3941 = ~n_3937 &  n_3940;
assign n_3942 = ~n_3936 &  n_3941;
assign n_3943 = ~n_3935 &  n_3942;
assign n_3944 = ~n_3934 &  n_3943;
assign n_3945 =  x_4403 & ~n_3944;
assign n_3946 = ~x_4403 &  n_3944;
assign n_3947 = ~n_3945 & ~n_3946;
assign n_3948 =  x_4402 &  n_3638;
assign n_3949 =  i_10 & ~n_3640;
assign n_3950 =  x_3681 &  n_3621;
assign n_3951 =  x_2660 &  n_3631;
assign n_3952 =  x_3777 &  n_3626;
assign n_3953 =  x_2692 &  n_3624;
assign n_3954 = ~n_3952 & ~n_3953;
assign n_3955 = ~n_3951 &  n_3954;
assign n_3956 = ~n_3950 &  n_3955;
assign n_3957 = ~n_3949 &  n_3956;
assign n_3958 = ~n_3948 &  n_3957;
assign n_3959 =  x_4402 & ~n_3958;
assign n_3960 = ~x_4402 &  n_3958;
assign n_3961 = ~n_3959 & ~n_3960;
assign n_3962 =  x_4401 &  n_3638;
assign n_3963 =  i_9 & ~n_3640;
assign n_3964 =  x_3680 &  n_3621;
assign n_3965 =  x_2659 &  n_3631;
assign n_3966 =  x_3776 &  n_3626;
assign n_3967 =  x_2691 &  n_3624;
assign n_3968 = ~n_3966 & ~n_3967;
assign n_3969 = ~n_3965 &  n_3968;
assign n_3970 = ~n_3964 &  n_3969;
assign n_3971 = ~n_3963 &  n_3970;
assign n_3972 = ~n_3962 &  n_3971;
assign n_3973 =  x_4401 & ~n_3972;
assign n_3974 = ~x_4401 &  n_3972;
assign n_3975 = ~n_3973 & ~n_3974;
assign n_3976 =  x_4400 &  n_3638;
assign n_3977 =  i_8 & ~n_3640;
assign n_3978 =  x_3679 &  n_3621;
assign n_3979 =  x_2658 &  n_3631;
assign n_3980 =  x_3775 &  n_3626;
assign n_3981 =  x_2690 &  n_3624;
assign n_3982 = ~n_3980 & ~n_3981;
assign n_3983 = ~n_3979 &  n_3982;
assign n_3984 = ~n_3978 &  n_3983;
assign n_3985 = ~n_3977 &  n_3984;
assign n_3986 = ~n_3976 &  n_3985;
assign n_3987 =  x_4400 & ~n_3986;
assign n_3988 = ~x_4400 &  n_3986;
assign n_3989 = ~n_3987 & ~n_3988;
assign n_3990 =  x_4399 &  n_3638;
assign n_3991 =  i_7 & ~n_3640;
assign n_3992 =  x_3678 &  n_3621;
assign n_3993 =  x_2657 &  n_3631;
assign n_3994 =  x_3774 &  n_3626;
assign n_3995 =  x_2689 &  n_3624;
assign n_3996 = ~n_3994 & ~n_3995;
assign n_3997 = ~n_3993 &  n_3996;
assign n_3998 = ~n_3992 &  n_3997;
assign n_3999 = ~n_3991 &  n_3998;
assign n_4000 = ~n_3990 &  n_3999;
assign n_4001 =  x_4399 & ~n_4000;
assign n_4002 = ~x_4399 &  n_4000;
assign n_4003 = ~n_4001 & ~n_4002;
assign n_4004 =  x_4398 &  n_3638;
assign n_4005 =  i_6 & ~n_3640;
assign n_4006 =  x_3677 &  n_3621;
assign n_4007 =  x_2656 &  n_3631;
assign n_4008 =  x_3773 &  n_3626;
assign n_4009 =  x_2688 &  n_3624;
assign n_4010 = ~n_4008 & ~n_4009;
assign n_4011 = ~n_4007 &  n_4010;
assign n_4012 = ~n_4006 &  n_4011;
assign n_4013 = ~n_4005 &  n_4012;
assign n_4014 = ~n_4004 &  n_4013;
assign n_4015 =  x_4398 & ~n_4014;
assign n_4016 = ~x_4398 &  n_4014;
assign n_4017 = ~n_4015 & ~n_4016;
assign n_4018 =  x_4397 &  n_3638;
assign n_4019 =  i_5 & ~n_3640;
assign n_4020 =  x_3676 &  n_3621;
assign n_4021 =  x_2655 &  n_3631;
assign n_4022 =  x_3772 &  n_3626;
assign n_4023 =  x_2687 &  n_3624;
assign n_4024 = ~n_4022 & ~n_4023;
assign n_4025 = ~n_4021 &  n_4024;
assign n_4026 = ~n_4020 &  n_4025;
assign n_4027 = ~n_4019 &  n_4026;
assign n_4028 = ~n_4018 &  n_4027;
assign n_4029 =  x_4397 & ~n_4028;
assign n_4030 = ~x_4397 &  n_4028;
assign n_4031 = ~n_4029 & ~n_4030;
assign n_4032 =  x_4396 &  n_3638;
assign n_4033 =  i_4 & ~n_3640;
assign n_4034 =  x_3675 &  n_3621;
assign n_4035 =  x_2654 &  n_3631;
assign n_4036 =  x_3771 &  n_3626;
assign n_4037 =  x_2686 &  n_3624;
assign n_4038 = ~n_4036 & ~n_4037;
assign n_4039 = ~n_4035 &  n_4038;
assign n_4040 = ~n_4034 &  n_4039;
assign n_4041 = ~n_4033 &  n_4040;
assign n_4042 = ~n_4032 &  n_4041;
assign n_4043 =  x_4396 & ~n_4042;
assign n_4044 = ~x_4396 &  n_4042;
assign n_4045 = ~n_4043 & ~n_4044;
assign n_4046 =  x_4395 &  n_3638;
assign n_4047 =  i_3 & ~n_3640;
assign n_4048 =  x_3674 &  n_3621;
assign n_4049 =  x_2653 &  n_3631;
assign n_4050 =  x_3770 &  n_3626;
assign n_4051 =  x_2685 &  n_3624;
assign n_4052 = ~n_4050 & ~n_4051;
assign n_4053 = ~n_4049 &  n_4052;
assign n_4054 = ~n_4048 &  n_4053;
assign n_4055 = ~n_4047 &  n_4054;
assign n_4056 = ~n_4046 &  n_4055;
assign n_4057 =  x_4395 & ~n_4056;
assign n_4058 = ~x_4395 &  n_4056;
assign n_4059 = ~n_4057 & ~n_4058;
assign n_4060 =  x_4394 &  n_3638;
assign n_4061 =  i_2 & ~n_3640;
assign n_4062 =  x_3673 &  n_3621;
assign n_4063 =  x_2652 &  n_3631;
assign n_4064 =  x_3769 &  n_3626;
assign n_4065 =  x_2684 &  n_3624;
assign n_4066 = ~n_4064 & ~n_4065;
assign n_4067 = ~n_4063 &  n_4066;
assign n_4068 = ~n_4062 &  n_4067;
assign n_4069 = ~n_4061 &  n_4068;
assign n_4070 = ~n_4060 &  n_4069;
assign n_4071 =  x_4394 & ~n_4070;
assign n_4072 = ~x_4394 &  n_4070;
assign n_4073 = ~n_4071 & ~n_4072;
assign n_4074 =  x_4393 &  n_3638;
assign n_4075 =  i_1 & ~n_3640;
assign n_4076 =  x_3672 &  n_3621;
assign n_4077 =  x_2651 &  n_3631;
assign n_4078 =  x_3768 &  n_3626;
assign n_4079 =  x_2683 &  n_3624;
assign n_4080 = ~n_4078 & ~n_4079;
assign n_4081 = ~n_4077 &  n_4080;
assign n_4082 = ~n_4076 &  n_4081;
assign n_4083 = ~n_4075 &  n_4082;
assign n_4084 = ~n_4074 &  n_4083;
assign n_4085 =  x_4393 & ~n_4084;
assign n_4086 = ~x_4393 &  n_4084;
assign n_4087 = ~n_4085 & ~n_4086;
assign n_4088 =  n_3341 &  n_759;
assign n_4089 = ~x_43 &  n_4088;
assign n_4090 =  n_4089 &  n_1173;
assign n_4091 =  x_4392 & ~n_4090;
assign n_4092 =  i_32 &  n_4090;
assign n_4093 = ~n_4091 & ~n_4092;
assign n_4094 =  x_4392 & ~n_4093;
assign n_4095 = ~x_4392 &  n_4093;
assign n_4096 = ~n_4094 & ~n_4095;
assign n_4097 =  x_4391 & ~n_4090;
assign n_4098 =  i_31 &  n_4090;
assign n_4099 = ~n_4097 & ~n_4098;
assign n_4100 =  x_4391 & ~n_4099;
assign n_4101 = ~x_4391 &  n_4099;
assign n_4102 = ~n_4100 & ~n_4101;
assign n_4103 =  x_4390 & ~n_4090;
assign n_4104 =  i_30 &  n_4090;
assign n_4105 = ~n_4103 & ~n_4104;
assign n_4106 =  x_4390 & ~n_4105;
assign n_4107 = ~x_4390 &  n_4105;
assign n_4108 = ~n_4106 & ~n_4107;
assign n_4109 =  x_4389 & ~n_4090;
assign n_4110 =  i_29 &  n_4090;
assign n_4111 = ~n_4109 & ~n_4110;
assign n_4112 =  x_4389 & ~n_4111;
assign n_4113 = ~x_4389 &  n_4111;
assign n_4114 = ~n_4112 & ~n_4113;
assign n_4115 =  x_4388 & ~n_4090;
assign n_4116 =  i_28 &  n_4090;
assign n_4117 = ~n_4115 & ~n_4116;
assign n_4118 =  x_4388 & ~n_4117;
assign n_4119 = ~x_4388 &  n_4117;
assign n_4120 = ~n_4118 & ~n_4119;
assign n_4121 =  x_4387 & ~n_4090;
assign n_4122 =  i_27 &  n_4090;
assign n_4123 = ~n_4121 & ~n_4122;
assign n_4124 =  x_4387 & ~n_4123;
assign n_4125 = ~x_4387 &  n_4123;
assign n_4126 = ~n_4124 & ~n_4125;
assign n_4127 =  x_4386 & ~n_4090;
assign n_4128 =  i_26 &  n_4090;
assign n_4129 = ~n_4127 & ~n_4128;
assign n_4130 =  x_4386 & ~n_4129;
assign n_4131 = ~x_4386 &  n_4129;
assign n_4132 = ~n_4130 & ~n_4131;
assign n_4133 =  x_4385 & ~n_4090;
assign n_4134 =  i_25 &  n_4090;
assign n_4135 = ~n_4133 & ~n_4134;
assign n_4136 =  x_4385 & ~n_4135;
assign n_4137 = ~x_4385 &  n_4135;
assign n_4138 = ~n_4136 & ~n_4137;
assign n_4139 =  x_4384 & ~n_4090;
assign n_4140 =  i_24 &  n_4090;
assign n_4141 = ~n_4139 & ~n_4140;
assign n_4142 =  x_4384 & ~n_4141;
assign n_4143 = ~x_4384 &  n_4141;
assign n_4144 = ~n_4142 & ~n_4143;
assign n_4145 =  x_4383 & ~n_4090;
assign n_4146 =  i_23 &  n_4090;
assign n_4147 = ~n_4145 & ~n_4146;
assign n_4148 =  x_4383 & ~n_4147;
assign n_4149 = ~x_4383 &  n_4147;
assign n_4150 = ~n_4148 & ~n_4149;
assign n_4151 =  x_4382 & ~n_4090;
assign n_4152 =  i_22 &  n_4090;
assign n_4153 = ~n_4151 & ~n_4152;
assign n_4154 =  x_4382 & ~n_4153;
assign n_4155 = ~x_4382 &  n_4153;
assign n_4156 = ~n_4154 & ~n_4155;
assign n_4157 =  x_4381 & ~n_4090;
assign n_4158 =  i_21 &  n_4090;
assign n_4159 = ~n_4157 & ~n_4158;
assign n_4160 =  x_4381 & ~n_4159;
assign n_4161 = ~x_4381 &  n_4159;
assign n_4162 = ~n_4160 & ~n_4161;
assign n_4163 =  x_4380 & ~n_4090;
assign n_4164 =  i_20 &  n_4090;
assign n_4165 = ~n_4163 & ~n_4164;
assign n_4166 =  x_4380 & ~n_4165;
assign n_4167 = ~x_4380 &  n_4165;
assign n_4168 = ~n_4166 & ~n_4167;
assign n_4169 =  x_4379 & ~n_4090;
assign n_4170 =  i_19 &  n_4090;
assign n_4171 = ~n_4169 & ~n_4170;
assign n_4172 =  x_4379 & ~n_4171;
assign n_4173 = ~x_4379 &  n_4171;
assign n_4174 = ~n_4172 & ~n_4173;
assign n_4175 =  x_4378 & ~n_4090;
assign n_4176 =  i_18 &  n_4090;
assign n_4177 = ~n_4175 & ~n_4176;
assign n_4178 =  x_4378 & ~n_4177;
assign n_4179 = ~x_4378 &  n_4177;
assign n_4180 = ~n_4178 & ~n_4179;
assign n_4181 =  x_4377 & ~n_4090;
assign n_4182 =  i_17 &  n_4090;
assign n_4183 = ~n_4181 & ~n_4182;
assign n_4184 =  x_4377 & ~n_4183;
assign n_4185 = ~x_4377 &  n_4183;
assign n_4186 = ~n_4184 & ~n_4185;
assign n_4187 =  x_4376 & ~n_4090;
assign n_4188 =  i_16 &  n_4090;
assign n_4189 = ~n_4187 & ~n_4188;
assign n_4190 =  x_4376 & ~n_4189;
assign n_4191 = ~x_4376 &  n_4189;
assign n_4192 = ~n_4190 & ~n_4191;
assign n_4193 =  x_4375 & ~n_4090;
assign n_4194 =  i_15 &  n_4090;
assign n_4195 = ~n_4193 & ~n_4194;
assign n_4196 =  x_4375 & ~n_4195;
assign n_4197 = ~x_4375 &  n_4195;
assign n_4198 = ~n_4196 & ~n_4197;
assign n_4199 =  x_4374 & ~n_4090;
assign n_4200 =  i_14 &  n_4090;
assign n_4201 = ~n_4199 & ~n_4200;
assign n_4202 =  x_4374 & ~n_4201;
assign n_4203 = ~x_4374 &  n_4201;
assign n_4204 = ~n_4202 & ~n_4203;
assign n_4205 =  x_4373 & ~n_4090;
assign n_4206 =  i_13 &  n_4090;
assign n_4207 = ~n_4205 & ~n_4206;
assign n_4208 =  x_4373 & ~n_4207;
assign n_4209 = ~x_4373 &  n_4207;
assign n_4210 = ~n_4208 & ~n_4209;
assign n_4211 =  x_4372 & ~n_4090;
assign n_4212 =  i_12 &  n_4090;
assign n_4213 = ~n_4211 & ~n_4212;
assign n_4214 =  x_4372 & ~n_4213;
assign n_4215 = ~x_4372 &  n_4213;
assign n_4216 = ~n_4214 & ~n_4215;
assign n_4217 =  x_4371 & ~n_4090;
assign n_4218 =  i_11 &  n_4090;
assign n_4219 = ~n_4217 & ~n_4218;
assign n_4220 =  x_4371 & ~n_4219;
assign n_4221 = ~x_4371 &  n_4219;
assign n_4222 = ~n_4220 & ~n_4221;
assign n_4223 =  x_4370 & ~n_4090;
assign n_4224 =  i_10 &  n_4090;
assign n_4225 = ~n_4223 & ~n_4224;
assign n_4226 =  x_4370 & ~n_4225;
assign n_4227 = ~x_4370 &  n_4225;
assign n_4228 = ~n_4226 & ~n_4227;
assign n_4229 =  x_4369 & ~n_4090;
assign n_4230 =  i_9 &  n_4090;
assign n_4231 = ~n_4229 & ~n_4230;
assign n_4232 =  x_4369 & ~n_4231;
assign n_4233 = ~x_4369 &  n_4231;
assign n_4234 = ~n_4232 & ~n_4233;
assign n_4235 =  x_4368 & ~n_4090;
assign n_4236 =  i_8 &  n_4090;
assign n_4237 = ~n_4235 & ~n_4236;
assign n_4238 =  x_4368 & ~n_4237;
assign n_4239 = ~x_4368 &  n_4237;
assign n_4240 = ~n_4238 & ~n_4239;
assign n_4241 =  x_4367 & ~n_4090;
assign n_4242 =  i_7 &  n_4090;
assign n_4243 = ~n_4241 & ~n_4242;
assign n_4244 =  x_4367 & ~n_4243;
assign n_4245 = ~x_4367 &  n_4243;
assign n_4246 = ~n_4244 & ~n_4245;
assign n_4247 =  x_4366 & ~n_4090;
assign n_4248 =  i_6 &  n_4090;
assign n_4249 = ~n_4247 & ~n_4248;
assign n_4250 =  x_4366 & ~n_4249;
assign n_4251 = ~x_4366 &  n_4249;
assign n_4252 = ~n_4250 & ~n_4251;
assign n_4253 =  x_4365 & ~n_4090;
assign n_4254 =  i_5 &  n_4090;
assign n_4255 = ~n_4253 & ~n_4254;
assign n_4256 =  x_4365 & ~n_4255;
assign n_4257 = ~x_4365 &  n_4255;
assign n_4258 = ~n_4256 & ~n_4257;
assign n_4259 =  x_4364 & ~n_4090;
assign n_4260 =  i_4 &  n_4090;
assign n_4261 = ~n_4259 & ~n_4260;
assign n_4262 =  x_4364 & ~n_4261;
assign n_4263 = ~x_4364 &  n_4261;
assign n_4264 = ~n_4262 & ~n_4263;
assign n_4265 =  x_4363 & ~n_4090;
assign n_4266 =  i_3 &  n_4090;
assign n_4267 = ~n_4265 & ~n_4266;
assign n_4268 =  x_4363 & ~n_4267;
assign n_4269 = ~x_4363 &  n_4267;
assign n_4270 = ~n_4268 & ~n_4269;
assign n_4271 =  x_4362 & ~n_4090;
assign n_4272 =  i_2 &  n_4090;
assign n_4273 = ~n_4271 & ~n_4272;
assign n_4274 =  x_4362 & ~n_4273;
assign n_4275 = ~x_4362 &  n_4273;
assign n_4276 = ~n_4274 & ~n_4275;
assign n_4277 =  x_4361 & ~n_4090;
assign n_4278 =  i_1 &  n_4090;
assign n_4279 = ~n_4277 & ~n_4278;
assign n_4280 =  x_4361 & ~n_4279;
assign n_4281 = ~x_4361 &  n_4279;
assign n_4282 = ~n_4280 & ~n_4281;
assign n_4283 =  n_13 &  n_1173;
assign n_4284 =  n_11 &  n_4283;
assign n_4285 = ~x_41 &  n_1174;
assign n_4286 =  n_1173 &  n_4285;
assign n_4287 =  n_1037 &  n_4286;
assign n_4288 =  n_148 &  n_147;
assign n_4289 =  x_37 &  n_4288;
assign n_4290 = ~x_38 &  n_4289;
assign n_4291 =  n_4290 &  n_3623;
assign n_4292 =  n_4290 &  n_760;
assign n_4293 = ~n_4291 & ~n_4292;
assign n_4294 = ~n_4287 &  n_4293;
assign n_4295 = ~n_4284 &  n_4294;
assign n_4296 =  x_4360 &  n_4295;
assign n_4297 =  x_4040 &  x_4136;
assign n_4298 = ~x_4040 & ~x_4136;
assign n_4299 = ~n_4297 & ~n_4298;
assign n_4300 =  n_4287 &  n_4299;
assign n_4301 =  x_715 &  x_4871;
assign n_4302 = ~x_715 & ~x_4871;
assign n_4303 = ~n_4301 & ~n_4302;
assign n_4304 =  n_4292 &  n_4303;
assign n_4305 =  x_1162 &  x_3287;
assign n_4306 = ~x_1162 & ~x_3287;
assign n_4307 = ~n_4305 & ~n_4306;
assign n_4308 =  n_4291 &  n_4307;
assign n_4309 = ~n_4304 & ~n_4308;
assign n_4310 = ~n_4300 &  n_4309;
assign n_4311 = ~n_4296 &  n_4310;
assign n_4312 =  x_4360 & ~n_4311;
assign n_4313 = ~x_4360 &  n_4311;
assign n_4314 = ~n_4312 & ~n_4313;
assign n_4315 =  x_4359 &  n_4295;
assign n_4316 = ~x_3286 & ~x_3287;
assign n_4317 =  x_3286 &  x_3287;
assign n_4318 = ~n_4316 & ~n_4317;
assign n_4319 =  x_1161 &  n_4318;
assign n_4320 = ~x_1161 & ~n_4318;
assign n_4321 = ~n_4319 & ~n_4320;
assign n_4322 = ~n_4305 & ~n_4321;
assign n_4323 =  n_4305 &  n_4321;
assign n_4324 =  n_4291 & ~n_4323;
assign n_4325 = ~n_4322 &  n_4324;
assign n_4326 = ~x_714 & ~x_715;
assign n_4327 =  x_714 &  x_715;
assign n_4328 = ~n_4326 & ~n_4327;
assign n_4329 =  x_4870 &  n_4328;
assign n_4330 = ~x_4870 & ~n_4328;
assign n_4331 = ~n_4329 & ~n_4330;
assign n_4332 = ~n_4301 & ~n_4331;
assign n_4333 =  n_4301 &  n_4331;
assign n_4334 =  n_4292 & ~n_4333;
assign n_4335 = ~n_4332 &  n_4334;
assign n_4336 = ~x_4135 & ~x_4136;
assign n_4337 =  x_4135 &  x_4136;
assign n_4338 = ~n_4336 & ~n_4337;
assign n_4339 =  x_4039 &  n_4338;
assign n_4340 = ~x_4039 & ~n_4338;
assign n_4341 = ~n_4339 & ~n_4340;
assign n_4342 =  n_4297 &  n_4341;
assign n_4343 = ~n_4297 & ~n_4341;
assign n_4344 = ~n_4342 & ~n_4343;
assign n_4345 =  n_4287 &  n_4344;
assign n_4346 = ~n_4335 & ~n_4345;
assign n_4347 = ~n_4325 &  n_4346;
assign n_4348 = ~n_4315 &  n_4347;
assign n_4349 =  x_4359 & ~n_4348;
assign n_4350 = ~x_4359 &  n_4348;
assign n_4351 = ~n_4349 & ~n_4350;
assign n_4352 =  x_4358 &  n_4295;
assign n_4353 = ~x_713 &  n_4326;
assign n_4354 =  x_713 & ~n_4326;
assign n_4355 = ~n_4353 & ~n_4354;
assign n_4356 =  x_714 & ~x_4870;
assign n_4357 =  n_4301 & ~n_4356;
assign n_4358 = ~n_4357 & ~n_4329;
assign n_4359 =  n_4355 & ~n_4358;
assign n_4360 = ~n_4355 &  n_4358;
assign n_4361 = ~n_4359 & ~n_4360;
assign n_4362 = ~x_4869 & ~n_4361;
assign n_4363 =  x_4869 & ~n_4360;
assign n_4364 = ~n_4359 &  n_4363;
assign n_4365 =  n_4292 & ~n_4364;
assign n_4366 = ~n_4362 &  n_4365;
assign n_4367 = ~n_4352 & ~n_4366;
assign n_4368 = ~x_3285 &  n_4316;
assign n_4369 =  x_3285 & ~n_4316;
assign n_4370 = ~n_4368 & ~n_4369;
assign n_4371 = ~x_1161 &  x_3286;
assign n_4372 =  n_4305 & ~n_4371;
assign n_4373 = ~n_4372 & ~n_4319;
assign n_4374 =  n_4370 & ~n_4373;
assign n_4375 = ~n_4370 &  n_4373;
assign n_4376 = ~n_4374 & ~n_4375;
assign n_4377 = ~x_1160 & ~n_4376;
assign n_4378 =  x_1160 & ~n_4375;
assign n_4379 = ~n_4374 &  n_4378;
assign n_4380 =  n_4291 & ~n_4379;
assign n_4381 = ~n_4377 &  n_4380;
assign n_4382 = ~x_4134 &  n_4336;
assign n_4383 =  x_4134 & ~n_4336;
assign n_4384 = ~n_4382 & ~n_4383;
assign n_4385 = ~x_4039 &  x_4135;
assign n_4386 =  n_4297 & ~n_4385;
assign n_4387 = ~n_4386 & ~n_4339;
assign n_4388 =  n_4384 & ~n_4387;
assign n_4389 = ~n_4384 &  n_4387;
assign n_4390 = ~n_4388 & ~n_4389;
assign n_4391 = ~x_4038 & ~n_4390;
assign n_4392 =  x_4038 & ~n_4389;
assign n_4393 = ~n_4388 &  n_4392;
assign n_4394 =  n_4287 & ~n_4393;
assign n_4395 = ~n_4391 &  n_4394;
assign n_4396 = ~n_4381 & ~n_4395;
assign n_4397 =  n_4367 &  n_4396;
assign n_4398 =  x_4358 & ~n_4397;
assign n_4399 = ~x_4358 &  n_4397;
assign n_4400 = ~n_4398 & ~n_4399;
assign n_4401 =  x_4357 &  n_4295;
assign n_4402 = ~x_712 &  n_4353;
assign n_4403 =  x_712 & ~n_4353;
assign n_4404 = ~n_4402 & ~n_4403;
assign n_4405 = ~n_4359 & ~n_4363;
assign n_4406 =  n_4404 & ~n_4405;
assign n_4407 = ~n_4404 &  n_4405;
assign n_4408 = ~n_4406 & ~n_4407;
assign n_4409 = ~x_4868 & ~n_4408;
assign n_4410 =  x_4868 & ~n_4407;
assign n_4411 = ~n_4406 &  n_4410;
assign n_4412 =  n_4292 & ~n_4411;
assign n_4413 = ~n_4409 &  n_4412;
assign n_4414 = ~n_4401 & ~n_4413;
assign n_4415 = ~x_3284 &  n_4368;
assign n_4416 =  x_3284 & ~n_4368;
assign n_4417 = ~n_4415 & ~n_4416;
assign n_4418 = ~n_4374 & ~n_4378;
assign n_4419 =  n_4417 & ~n_4418;
assign n_4420 = ~n_4417 &  n_4418;
assign n_4421 = ~n_4419 & ~n_4420;
assign n_4422 = ~x_1159 & ~n_4421;
assign n_4423 =  x_1159 & ~n_4420;
assign n_4424 = ~n_4419 &  n_4423;
assign n_4425 =  n_4291 & ~n_4424;
assign n_4426 = ~n_4422 &  n_4425;
assign n_4427 = ~x_4133 &  n_4382;
assign n_4428 =  x_4133 & ~n_4382;
assign n_4429 = ~n_4427 & ~n_4428;
assign n_4430 = ~n_4388 & ~n_4392;
assign n_4431 =  n_4429 & ~n_4430;
assign n_4432 = ~n_4429 &  n_4430;
assign n_4433 = ~n_4431 & ~n_4432;
assign n_4434 = ~x_4037 & ~n_4433;
assign n_4435 =  x_4037 & ~n_4432;
assign n_4436 = ~n_4431 &  n_4435;
assign n_4437 =  n_4287 & ~n_4436;
assign n_4438 = ~n_4434 &  n_4437;
assign n_4439 = ~n_4426 & ~n_4438;
assign n_4440 =  n_4414 &  n_4439;
assign n_4441 =  x_4357 & ~n_4440;
assign n_4442 = ~x_4357 &  n_4440;
assign n_4443 = ~n_4441 & ~n_4442;
assign n_4444 =  x_4356 &  n_4295;
assign n_4445 = ~x_3283 &  n_4415;
assign n_4446 =  x_3283 & ~n_4415;
assign n_4447 = ~n_4445 & ~n_4446;
assign n_4448 = ~n_4419 & ~n_4423;
assign n_4449 =  n_4447 & ~n_4448;
assign n_4450 = ~n_4447 &  n_4448;
assign n_4451 = ~n_4449 & ~n_4450;
assign n_4452 = ~x_1158 & ~n_4451;
assign n_4453 =  x_1158 & ~n_4450;
assign n_4454 = ~n_4449 &  n_4453;
assign n_4455 =  n_4291 & ~n_4454;
assign n_4456 = ~n_4452 &  n_4455;
assign n_4457 = ~n_4444 & ~n_4456;
assign n_4458 = ~x_4132 &  n_4427;
assign n_4459 =  x_4132 & ~n_4427;
assign n_4460 = ~n_4458 & ~n_4459;
assign n_4461 = ~n_4431 & ~n_4435;
assign n_4462 =  n_4460 & ~n_4461;
assign n_4463 = ~n_4460 &  n_4461;
assign n_4464 = ~n_4462 & ~n_4463;
assign n_4465 = ~x_4036 & ~n_4464;
assign n_4466 =  x_4036 & ~n_4463;
assign n_4467 = ~n_4462 &  n_4466;
assign n_4468 =  n_4287 & ~n_4467;
assign n_4469 = ~n_4465 &  n_4468;
assign n_4470 = ~x_711 &  n_4402;
assign n_4471 =  x_711 & ~n_4402;
assign n_4472 = ~n_4470 & ~n_4471;
assign n_4473 = ~n_4406 & ~n_4410;
assign n_4474 =  n_4472 & ~n_4473;
assign n_4475 = ~n_4472 &  n_4473;
assign n_4476 = ~n_4474 & ~n_4475;
assign n_4477 = ~x_4867 & ~n_4476;
assign n_4478 =  x_4867 & ~n_4475;
assign n_4479 = ~n_4474 &  n_4478;
assign n_4480 =  n_4292 & ~n_4479;
assign n_4481 = ~n_4477 &  n_4480;
assign n_4482 = ~n_4469 & ~n_4481;
assign n_4483 =  n_4457 &  n_4482;
assign n_4484 =  x_4356 & ~n_4483;
assign n_4485 = ~x_4356 &  n_4483;
assign n_4486 = ~n_4484 & ~n_4485;
assign n_4487 =  x_4355 &  n_4295;
assign n_4488 = ~x_3282 &  n_4445;
assign n_4489 =  x_3282 & ~n_4445;
assign n_4490 = ~n_4488 & ~n_4489;
assign n_4491 = ~n_4449 & ~n_4453;
assign n_4492 =  n_4490 & ~n_4491;
assign n_4493 = ~n_4490 &  n_4491;
assign n_4494 = ~n_4492 & ~n_4493;
assign n_4495 = ~x_1157 & ~n_4494;
assign n_4496 =  x_1157 & ~n_4493;
assign n_4497 = ~n_4492 &  n_4496;
assign n_4498 =  n_4291 & ~n_4497;
assign n_4499 = ~n_4495 &  n_4498;
assign n_4500 = ~n_4487 & ~n_4499;
assign n_4501 = ~x_4131 &  n_4458;
assign n_4502 =  x_4131 & ~n_4458;
assign n_4503 = ~n_4501 & ~n_4502;
assign n_4504 = ~n_4462 & ~n_4466;
assign n_4505 =  n_4503 & ~n_4504;
assign n_4506 = ~n_4503 &  n_4504;
assign n_4507 = ~n_4505 & ~n_4506;
assign n_4508 = ~x_4035 & ~n_4507;
assign n_4509 =  x_4035 & ~n_4506;
assign n_4510 = ~n_4505 &  n_4509;
assign n_4511 =  n_4287 & ~n_4510;
assign n_4512 = ~n_4508 &  n_4511;
assign n_4513 = ~x_710 &  n_4470;
assign n_4514 =  x_710 & ~n_4470;
assign n_4515 = ~n_4513 & ~n_4514;
assign n_4516 = ~n_4474 & ~n_4478;
assign n_4517 =  n_4515 & ~n_4516;
assign n_4518 = ~n_4515 &  n_4516;
assign n_4519 = ~n_4517 & ~n_4518;
assign n_4520 = ~x_4866 & ~n_4519;
assign n_4521 =  x_4866 & ~n_4518;
assign n_4522 = ~n_4517 &  n_4521;
assign n_4523 =  n_4292 & ~n_4522;
assign n_4524 = ~n_4520 &  n_4523;
assign n_4525 = ~n_4512 & ~n_4524;
assign n_4526 =  n_4500 &  n_4525;
assign n_4527 =  x_4355 & ~n_4526;
assign n_4528 = ~x_4355 &  n_4526;
assign n_4529 = ~n_4527 & ~n_4528;
assign n_4530 =  x_4354 &  n_4295;
assign n_4531 = ~x_3281 &  n_4488;
assign n_4532 =  x_3281 & ~n_4488;
assign n_4533 = ~n_4531 & ~n_4532;
assign n_4534 = ~n_4492 & ~n_4496;
assign n_4535 =  n_4533 & ~n_4534;
assign n_4536 = ~n_4533 &  n_4534;
assign n_4537 = ~n_4535 & ~n_4536;
assign n_4538 = ~x_1156 & ~n_4537;
assign n_4539 =  x_1156 & ~n_4536;
assign n_4540 = ~n_4535 &  n_4539;
assign n_4541 =  n_4291 & ~n_4540;
assign n_4542 = ~n_4538 &  n_4541;
assign n_4543 = ~n_4530 & ~n_4542;
assign n_4544 = ~x_4130 &  n_4501;
assign n_4545 =  x_4130 & ~n_4501;
assign n_4546 = ~n_4544 & ~n_4545;
assign n_4547 = ~n_4505 & ~n_4509;
assign n_4548 =  n_4546 & ~n_4547;
assign n_4549 = ~n_4546 &  n_4547;
assign n_4550 = ~n_4548 & ~n_4549;
assign n_4551 = ~x_4034 & ~n_4550;
assign n_4552 =  x_4034 & ~n_4549;
assign n_4553 = ~n_4548 &  n_4552;
assign n_4554 =  n_4287 & ~n_4553;
assign n_4555 = ~n_4551 &  n_4554;
assign n_4556 = ~x_709 &  n_4513;
assign n_4557 =  x_709 & ~n_4513;
assign n_4558 = ~n_4556 & ~n_4557;
assign n_4559 = ~n_4517 & ~n_4521;
assign n_4560 =  n_4558 & ~n_4559;
assign n_4561 = ~n_4558 &  n_4559;
assign n_4562 = ~n_4560 & ~n_4561;
assign n_4563 = ~x_4865 & ~n_4562;
assign n_4564 =  x_4865 & ~n_4561;
assign n_4565 = ~n_4560 &  n_4564;
assign n_4566 =  n_4292 & ~n_4565;
assign n_4567 = ~n_4563 &  n_4566;
assign n_4568 = ~n_4555 & ~n_4567;
assign n_4569 =  n_4543 &  n_4568;
assign n_4570 =  x_4354 & ~n_4569;
assign n_4571 = ~x_4354 &  n_4569;
assign n_4572 = ~n_4570 & ~n_4571;
assign n_4573 =  x_4353 &  n_4295;
assign n_4574 = ~x_3280 &  n_4531;
assign n_4575 =  x_3280 & ~n_4531;
assign n_4576 = ~n_4574 & ~n_4575;
assign n_4577 = ~n_4535 & ~n_4539;
assign n_4578 =  n_4576 & ~n_4577;
assign n_4579 = ~n_4576 &  n_4577;
assign n_4580 = ~n_4578 & ~n_4579;
assign n_4581 = ~x_1155 & ~n_4580;
assign n_4582 =  x_1155 & ~n_4579;
assign n_4583 = ~n_4578 &  n_4582;
assign n_4584 =  n_4291 & ~n_4583;
assign n_4585 = ~n_4581 &  n_4584;
assign n_4586 = ~n_4573 & ~n_4585;
assign n_4587 = ~x_4129 &  n_4544;
assign n_4588 =  x_4129 & ~n_4544;
assign n_4589 = ~n_4587 & ~n_4588;
assign n_4590 = ~n_4548 & ~n_4552;
assign n_4591 =  n_4589 & ~n_4590;
assign n_4592 = ~n_4589 &  n_4590;
assign n_4593 = ~n_4591 & ~n_4592;
assign n_4594 = ~x_4033 & ~n_4593;
assign n_4595 =  x_4033 & ~n_4592;
assign n_4596 = ~n_4591 &  n_4595;
assign n_4597 =  n_4287 & ~n_4596;
assign n_4598 = ~n_4594 &  n_4597;
assign n_4599 = ~x_708 &  n_4556;
assign n_4600 =  x_708 & ~n_4556;
assign n_4601 = ~n_4599 & ~n_4600;
assign n_4602 = ~n_4560 & ~n_4564;
assign n_4603 =  n_4601 & ~n_4602;
assign n_4604 = ~n_4601 &  n_4602;
assign n_4605 = ~n_4603 & ~n_4604;
assign n_4606 = ~x_4864 & ~n_4605;
assign n_4607 =  x_4864 & ~n_4604;
assign n_4608 = ~n_4603 &  n_4607;
assign n_4609 =  n_4292 & ~n_4608;
assign n_4610 = ~n_4606 &  n_4609;
assign n_4611 = ~n_4598 & ~n_4610;
assign n_4612 =  n_4586 &  n_4611;
assign n_4613 =  x_4353 & ~n_4612;
assign n_4614 = ~x_4353 &  n_4612;
assign n_4615 = ~n_4613 & ~n_4614;
assign n_4616 =  x_4352 &  n_4295;
assign n_4617 = ~x_3279 &  n_4574;
assign n_4618 =  x_3279 & ~n_4574;
assign n_4619 = ~n_4617 & ~n_4618;
assign n_4620 = ~n_4578 & ~n_4582;
assign n_4621 =  n_4619 & ~n_4620;
assign n_4622 = ~n_4619 &  n_4620;
assign n_4623 = ~n_4621 & ~n_4622;
assign n_4624 = ~x_1154 & ~n_4623;
assign n_4625 =  x_1154 & ~n_4622;
assign n_4626 = ~n_4621 &  n_4625;
assign n_4627 =  n_4291 & ~n_4626;
assign n_4628 = ~n_4624 &  n_4627;
assign n_4629 = ~n_4616 & ~n_4628;
assign n_4630 = ~x_4128 &  n_4587;
assign n_4631 =  x_4128 & ~n_4587;
assign n_4632 = ~n_4630 & ~n_4631;
assign n_4633 = ~n_4591 & ~n_4595;
assign n_4634 =  n_4632 & ~n_4633;
assign n_4635 = ~n_4632 &  n_4633;
assign n_4636 = ~n_4634 & ~n_4635;
assign n_4637 = ~x_4032 & ~n_4636;
assign n_4638 =  x_4032 & ~n_4635;
assign n_4639 = ~n_4634 &  n_4638;
assign n_4640 =  n_4287 & ~n_4639;
assign n_4641 = ~n_4637 &  n_4640;
assign n_4642 = ~x_707 &  n_4599;
assign n_4643 =  x_707 & ~n_4599;
assign n_4644 = ~n_4642 & ~n_4643;
assign n_4645 = ~n_4603 & ~n_4607;
assign n_4646 =  n_4644 & ~n_4645;
assign n_4647 = ~n_4644 &  n_4645;
assign n_4648 = ~n_4646 & ~n_4647;
assign n_4649 = ~x_4863 & ~n_4648;
assign n_4650 =  x_4863 & ~n_4647;
assign n_4651 = ~n_4646 &  n_4650;
assign n_4652 =  n_4292 & ~n_4651;
assign n_4653 = ~n_4649 &  n_4652;
assign n_4654 = ~n_4641 & ~n_4653;
assign n_4655 =  n_4629 &  n_4654;
assign n_4656 =  x_4352 & ~n_4655;
assign n_4657 = ~x_4352 &  n_4655;
assign n_4658 = ~n_4656 & ~n_4657;
assign n_4659 =  x_4351 &  n_4295;
assign n_4660 = ~x_3278 &  n_4617;
assign n_4661 =  x_3278 & ~n_4617;
assign n_4662 = ~n_4660 & ~n_4661;
assign n_4663 = ~n_4621 & ~n_4625;
assign n_4664 =  n_4662 & ~n_4663;
assign n_4665 = ~n_4662 &  n_4663;
assign n_4666 = ~n_4664 & ~n_4665;
assign n_4667 = ~x_1153 & ~n_4666;
assign n_4668 =  x_1153 & ~n_4665;
assign n_4669 = ~n_4664 &  n_4668;
assign n_4670 =  n_4291 & ~n_4669;
assign n_4671 = ~n_4667 &  n_4670;
assign n_4672 = ~n_4659 & ~n_4671;
assign n_4673 = ~x_4127 &  n_4630;
assign n_4674 =  x_4127 & ~n_4630;
assign n_4675 = ~n_4673 & ~n_4674;
assign n_4676 = ~n_4634 & ~n_4638;
assign n_4677 =  n_4675 & ~n_4676;
assign n_4678 = ~n_4675 &  n_4676;
assign n_4679 = ~n_4677 & ~n_4678;
assign n_4680 = ~x_4031 & ~n_4679;
assign n_4681 =  x_4031 & ~n_4678;
assign n_4682 = ~n_4677 &  n_4681;
assign n_4683 =  n_4287 & ~n_4682;
assign n_4684 = ~n_4680 &  n_4683;
assign n_4685 = ~x_706 &  n_4642;
assign n_4686 =  x_706 & ~n_4642;
assign n_4687 = ~n_4685 & ~n_4686;
assign n_4688 = ~n_4646 & ~n_4650;
assign n_4689 =  n_4687 & ~n_4688;
assign n_4690 = ~n_4687 &  n_4688;
assign n_4691 = ~n_4689 & ~n_4690;
assign n_4692 = ~x_4862 & ~n_4691;
assign n_4693 =  x_4862 & ~n_4690;
assign n_4694 = ~n_4689 &  n_4693;
assign n_4695 =  n_4292 & ~n_4694;
assign n_4696 = ~n_4692 &  n_4695;
assign n_4697 = ~n_4684 & ~n_4696;
assign n_4698 =  n_4672 &  n_4697;
assign n_4699 =  x_4351 & ~n_4698;
assign n_4700 = ~x_4351 &  n_4698;
assign n_4701 = ~n_4699 & ~n_4700;
assign n_4702 =  x_4350 &  n_4295;
assign n_4703 = ~x_3277 &  n_4660;
assign n_4704 =  x_3277 & ~n_4660;
assign n_4705 = ~n_4703 & ~n_4704;
assign n_4706 = ~n_4664 & ~n_4668;
assign n_4707 =  n_4705 & ~n_4706;
assign n_4708 = ~n_4705 &  n_4706;
assign n_4709 = ~n_4707 & ~n_4708;
assign n_4710 = ~x_1152 & ~n_4709;
assign n_4711 =  x_1152 & ~n_4708;
assign n_4712 = ~n_4707 &  n_4711;
assign n_4713 =  n_4291 & ~n_4712;
assign n_4714 = ~n_4710 &  n_4713;
assign n_4715 = ~n_4702 & ~n_4714;
assign n_4716 = ~x_4126 &  n_4673;
assign n_4717 =  x_4126 & ~n_4673;
assign n_4718 = ~n_4716 & ~n_4717;
assign n_4719 = ~n_4677 & ~n_4681;
assign n_4720 =  n_4718 & ~n_4719;
assign n_4721 = ~n_4718 &  n_4719;
assign n_4722 = ~n_4720 & ~n_4721;
assign n_4723 = ~x_4030 & ~n_4722;
assign n_4724 =  x_4030 & ~n_4721;
assign n_4725 = ~n_4720 &  n_4724;
assign n_4726 =  n_4287 & ~n_4725;
assign n_4727 = ~n_4723 &  n_4726;
assign n_4728 = ~x_705 &  n_4685;
assign n_4729 =  x_705 & ~n_4685;
assign n_4730 = ~n_4728 & ~n_4729;
assign n_4731 = ~n_4689 & ~n_4693;
assign n_4732 =  n_4730 & ~n_4731;
assign n_4733 = ~n_4730 &  n_4731;
assign n_4734 = ~n_4732 & ~n_4733;
assign n_4735 = ~x_4861 & ~n_4734;
assign n_4736 =  x_4861 & ~n_4733;
assign n_4737 = ~n_4732 &  n_4736;
assign n_4738 =  n_4292 & ~n_4737;
assign n_4739 = ~n_4735 &  n_4738;
assign n_4740 = ~n_4727 & ~n_4739;
assign n_4741 =  n_4715 &  n_4740;
assign n_4742 =  x_4350 & ~n_4741;
assign n_4743 = ~x_4350 &  n_4741;
assign n_4744 = ~n_4742 & ~n_4743;
assign n_4745 =  x_4349 &  n_4295;
assign n_4746 = ~x_3276 &  n_4703;
assign n_4747 =  x_3276 & ~n_4703;
assign n_4748 = ~n_4746 & ~n_4747;
assign n_4749 = ~n_4707 & ~n_4711;
assign n_4750 =  n_4748 & ~n_4749;
assign n_4751 = ~n_4748 &  n_4749;
assign n_4752 = ~n_4750 & ~n_4751;
assign n_4753 = ~x_1151 & ~n_4752;
assign n_4754 =  x_1151 & ~n_4751;
assign n_4755 = ~n_4750 &  n_4754;
assign n_4756 =  n_4291 & ~n_4755;
assign n_4757 = ~n_4753 &  n_4756;
assign n_4758 = ~n_4745 & ~n_4757;
assign n_4759 = ~x_4125 &  n_4716;
assign n_4760 =  x_4125 & ~n_4716;
assign n_4761 = ~n_4759 & ~n_4760;
assign n_4762 = ~n_4720 & ~n_4724;
assign n_4763 =  n_4761 & ~n_4762;
assign n_4764 = ~n_4761 &  n_4762;
assign n_4765 = ~n_4763 & ~n_4764;
assign n_4766 = ~x_4029 & ~n_4765;
assign n_4767 =  x_4029 & ~n_4764;
assign n_4768 = ~n_4763 &  n_4767;
assign n_4769 =  n_4287 & ~n_4768;
assign n_4770 = ~n_4766 &  n_4769;
assign n_4771 = ~x_704 &  n_4728;
assign n_4772 =  x_704 & ~n_4728;
assign n_4773 = ~n_4771 & ~n_4772;
assign n_4774 = ~n_4732 & ~n_4736;
assign n_4775 =  n_4773 & ~n_4774;
assign n_4776 = ~n_4773 &  n_4774;
assign n_4777 = ~n_4775 & ~n_4776;
assign n_4778 = ~x_4860 & ~n_4777;
assign n_4779 =  x_4860 & ~n_4776;
assign n_4780 = ~n_4775 &  n_4779;
assign n_4781 =  n_4292 & ~n_4780;
assign n_4782 = ~n_4778 &  n_4781;
assign n_4783 = ~n_4770 & ~n_4782;
assign n_4784 =  n_4758 &  n_4783;
assign n_4785 =  x_4349 & ~n_4784;
assign n_4786 = ~x_4349 &  n_4784;
assign n_4787 = ~n_4785 & ~n_4786;
assign n_4788 =  x_4348 &  n_4295;
assign n_4789 = ~x_3275 &  n_4746;
assign n_4790 =  x_3275 & ~n_4746;
assign n_4791 = ~n_4789 & ~n_4790;
assign n_4792 = ~n_4750 & ~n_4754;
assign n_4793 =  n_4791 & ~n_4792;
assign n_4794 = ~n_4791 &  n_4792;
assign n_4795 = ~n_4793 & ~n_4794;
assign n_4796 = ~x_1150 & ~n_4795;
assign n_4797 =  x_1150 & ~n_4794;
assign n_4798 = ~n_4793 &  n_4797;
assign n_4799 =  n_4291 & ~n_4798;
assign n_4800 = ~n_4796 &  n_4799;
assign n_4801 = ~n_4788 & ~n_4800;
assign n_4802 = ~x_4124 &  n_4759;
assign n_4803 =  x_4124 & ~n_4759;
assign n_4804 = ~n_4802 & ~n_4803;
assign n_4805 = ~n_4763 & ~n_4767;
assign n_4806 =  n_4804 & ~n_4805;
assign n_4807 = ~n_4804 &  n_4805;
assign n_4808 = ~n_4806 & ~n_4807;
assign n_4809 = ~x_4028 & ~n_4808;
assign n_4810 =  x_4028 & ~n_4807;
assign n_4811 = ~n_4806 &  n_4810;
assign n_4812 =  n_4287 & ~n_4811;
assign n_4813 = ~n_4809 &  n_4812;
assign n_4814 = ~x_703 &  n_4771;
assign n_4815 =  x_703 & ~n_4771;
assign n_4816 = ~n_4814 & ~n_4815;
assign n_4817 = ~n_4775 & ~n_4779;
assign n_4818 =  n_4816 & ~n_4817;
assign n_4819 = ~n_4816 &  n_4817;
assign n_4820 = ~n_4818 & ~n_4819;
assign n_4821 = ~x_4859 & ~n_4820;
assign n_4822 =  x_4859 & ~n_4819;
assign n_4823 = ~n_4818 &  n_4822;
assign n_4824 =  n_4292 & ~n_4823;
assign n_4825 = ~n_4821 &  n_4824;
assign n_4826 = ~n_4813 & ~n_4825;
assign n_4827 =  n_4801 &  n_4826;
assign n_4828 =  x_4348 & ~n_4827;
assign n_4829 = ~x_4348 &  n_4827;
assign n_4830 = ~n_4828 & ~n_4829;
assign n_4831 =  x_4347 &  n_4295;
assign n_4832 = ~x_3274 &  n_4789;
assign n_4833 =  x_3274 & ~n_4789;
assign n_4834 = ~n_4832 & ~n_4833;
assign n_4835 = ~n_4793 & ~n_4797;
assign n_4836 =  n_4834 & ~n_4835;
assign n_4837 = ~n_4834 &  n_4835;
assign n_4838 = ~n_4836 & ~n_4837;
assign n_4839 = ~x_1149 & ~n_4838;
assign n_4840 =  x_1149 & ~n_4837;
assign n_4841 = ~n_4836 &  n_4840;
assign n_4842 =  n_4291 & ~n_4841;
assign n_4843 = ~n_4839 &  n_4842;
assign n_4844 = ~n_4831 & ~n_4843;
assign n_4845 = ~x_4123 &  n_4802;
assign n_4846 =  x_4123 & ~n_4802;
assign n_4847 = ~n_4845 & ~n_4846;
assign n_4848 = ~n_4806 & ~n_4810;
assign n_4849 =  n_4847 & ~n_4848;
assign n_4850 = ~n_4847 &  n_4848;
assign n_4851 = ~n_4849 & ~n_4850;
assign n_4852 = ~x_4027 & ~n_4851;
assign n_4853 =  x_4027 & ~n_4850;
assign n_4854 = ~n_4849 &  n_4853;
assign n_4855 =  n_4287 & ~n_4854;
assign n_4856 = ~n_4852 &  n_4855;
assign n_4857 = ~x_702 &  n_4814;
assign n_4858 =  x_702 & ~n_4814;
assign n_4859 = ~n_4857 & ~n_4858;
assign n_4860 = ~n_4818 & ~n_4822;
assign n_4861 =  n_4859 & ~n_4860;
assign n_4862 = ~n_4859 &  n_4860;
assign n_4863 = ~n_4861 & ~n_4862;
assign n_4864 = ~x_4858 & ~n_4863;
assign n_4865 =  x_4858 & ~n_4862;
assign n_4866 = ~n_4861 &  n_4865;
assign n_4867 =  n_4292 & ~n_4866;
assign n_4868 = ~n_4864 &  n_4867;
assign n_4869 = ~n_4856 & ~n_4868;
assign n_4870 =  n_4844 &  n_4869;
assign n_4871 =  x_4347 & ~n_4870;
assign n_4872 = ~x_4347 &  n_4870;
assign n_4873 = ~n_4871 & ~n_4872;
assign n_4874 =  x_4346 &  n_4295;
assign n_4875 = ~x_3273 &  n_4832;
assign n_4876 =  x_3273 & ~n_4832;
assign n_4877 = ~n_4875 & ~n_4876;
assign n_4878 = ~n_4836 & ~n_4840;
assign n_4879 =  n_4877 & ~n_4878;
assign n_4880 = ~n_4877 &  n_4878;
assign n_4881 = ~n_4879 & ~n_4880;
assign n_4882 = ~x_1148 & ~n_4881;
assign n_4883 =  x_1148 & ~n_4880;
assign n_4884 = ~n_4879 &  n_4883;
assign n_4885 =  n_4291 & ~n_4884;
assign n_4886 = ~n_4882 &  n_4885;
assign n_4887 = ~n_4874 & ~n_4886;
assign n_4888 = ~x_4122 &  n_4845;
assign n_4889 =  x_4122 & ~n_4845;
assign n_4890 = ~n_4888 & ~n_4889;
assign n_4891 = ~n_4849 & ~n_4853;
assign n_4892 =  n_4890 & ~n_4891;
assign n_4893 = ~n_4890 &  n_4891;
assign n_4894 = ~n_4892 & ~n_4893;
assign n_4895 = ~x_4026 & ~n_4894;
assign n_4896 =  x_4026 & ~n_4893;
assign n_4897 = ~n_4892 &  n_4896;
assign n_4898 =  n_4287 & ~n_4897;
assign n_4899 = ~n_4895 &  n_4898;
assign n_4900 = ~x_701 &  n_4857;
assign n_4901 =  x_701 & ~n_4857;
assign n_4902 = ~n_4900 & ~n_4901;
assign n_4903 = ~n_4861 & ~n_4865;
assign n_4904 =  n_4902 & ~n_4903;
assign n_4905 = ~n_4902 &  n_4903;
assign n_4906 = ~n_4904 & ~n_4905;
assign n_4907 = ~x_4857 & ~n_4906;
assign n_4908 =  x_4857 & ~n_4905;
assign n_4909 = ~n_4904 &  n_4908;
assign n_4910 =  n_4292 & ~n_4909;
assign n_4911 = ~n_4907 &  n_4910;
assign n_4912 = ~n_4899 & ~n_4911;
assign n_4913 =  n_4887 &  n_4912;
assign n_4914 =  x_4346 & ~n_4913;
assign n_4915 = ~x_4346 &  n_4913;
assign n_4916 = ~n_4914 & ~n_4915;
assign n_4917 =  x_4345 &  n_4295;
assign n_4918 = ~x_3272 &  n_4875;
assign n_4919 =  x_3272 & ~n_4875;
assign n_4920 = ~n_4918 & ~n_4919;
assign n_4921 = ~n_4879 & ~n_4883;
assign n_4922 =  n_4920 & ~n_4921;
assign n_4923 = ~n_4920 &  n_4921;
assign n_4924 = ~n_4922 & ~n_4923;
assign n_4925 = ~x_1147 & ~n_4924;
assign n_4926 =  x_1147 & ~n_4923;
assign n_4927 = ~n_4922 &  n_4926;
assign n_4928 =  n_4291 & ~n_4927;
assign n_4929 = ~n_4925 &  n_4928;
assign n_4930 = ~n_4917 & ~n_4929;
assign n_4931 = ~x_4121 &  n_4888;
assign n_4932 =  x_4121 & ~n_4888;
assign n_4933 = ~n_4931 & ~n_4932;
assign n_4934 = ~n_4892 & ~n_4896;
assign n_4935 =  n_4933 & ~n_4934;
assign n_4936 = ~n_4933 &  n_4934;
assign n_4937 = ~n_4935 & ~n_4936;
assign n_4938 = ~x_4025 & ~n_4937;
assign n_4939 =  x_4025 & ~n_4936;
assign n_4940 = ~n_4935 &  n_4939;
assign n_4941 =  n_4287 & ~n_4940;
assign n_4942 = ~n_4938 &  n_4941;
assign n_4943 = ~x_700 &  n_4900;
assign n_4944 =  x_700 & ~n_4900;
assign n_4945 = ~n_4943 & ~n_4944;
assign n_4946 = ~n_4904 & ~n_4908;
assign n_4947 =  n_4945 & ~n_4946;
assign n_4948 = ~n_4945 &  n_4946;
assign n_4949 = ~n_4947 & ~n_4948;
assign n_4950 = ~x_4856 & ~n_4949;
assign n_4951 =  x_4856 & ~n_4948;
assign n_4952 = ~n_4947 &  n_4951;
assign n_4953 =  n_4292 & ~n_4952;
assign n_4954 = ~n_4950 &  n_4953;
assign n_4955 = ~n_4942 & ~n_4954;
assign n_4956 =  n_4930 &  n_4955;
assign n_4957 =  x_4345 & ~n_4956;
assign n_4958 = ~x_4345 &  n_4956;
assign n_4959 = ~n_4957 & ~n_4958;
assign n_4960 =  x_4344 &  n_4295;
assign n_4961 = ~x_3271 &  n_4918;
assign n_4962 =  x_3271 & ~n_4918;
assign n_4963 = ~n_4961 & ~n_4962;
assign n_4964 = ~n_4922 & ~n_4926;
assign n_4965 =  n_4963 & ~n_4964;
assign n_4966 = ~n_4963 &  n_4964;
assign n_4967 = ~n_4965 & ~n_4966;
assign n_4968 = ~x_1146 & ~n_4967;
assign n_4969 =  x_1146 & ~n_4966;
assign n_4970 = ~n_4965 &  n_4969;
assign n_4971 =  n_4291 & ~n_4970;
assign n_4972 = ~n_4968 &  n_4971;
assign n_4973 = ~n_4960 & ~n_4972;
assign n_4974 = ~x_4120 &  n_4931;
assign n_4975 =  x_4120 & ~n_4931;
assign n_4976 = ~n_4974 & ~n_4975;
assign n_4977 = ~n_4935 & ~n_4939;
assign n_4978 =  n_4976 & ~n_4977;
assign n_4979 = ~n_4976 &  n_4977;
assign n_4980 = ~n_4978 & ~n_4979;
assign n_4981 = ~x_4024 & ~n_4980;
assign n_4982 =  x_4024 & ~n_4979;
assign n_4983 = ~n_4978 &  n_4982;
assign n_4984 =  n_4287 & ~n_4983;
assign n_4985 = ~n_4981 &  n_4984;
assign n_4986 = ~x_699 &  n_4943;
assign n_4987 =  x_699 & ~n_4943;
assign n_4988 = ~n_4986 & ~n_4987;
assign n_4989 = ~n_4947 & ~n_4951;
assign n_4990 =  n_4988 & ~n_4989;
assign n_4991 = ~n_4988 &  n_4989;
assign n_4992 = ~n_4990 & ~n_4991;
assign n_4993 = ~x_4855 & ~n_4992;
assign n_4994 =  x_4855 & ~n_4991;
assign n_4995 = ~n_4990 &  n_4994;
assign n_4996 =  n_4292 & ~n_4995;
assign n_4997 = ~n_4993 &  n_4996;
assign n_4998 = ~n_4985 & ~n_4997;
assign n_4999 =  n_4973 &  n_4998;
assign n_5000 =  x_4344 & ~n_4999;
assign n_5001 = ~x_4344 &  n_4999;
assign n_5002 = ~n_5000 & ~n_5001;
assign n_5003 =  x_4343 &  n_4295;
assign n_5004 = ~x_3270 &  n_4961;
assign n_5005 =  x_3270 & ~n_4961;
assign n_5006 = ~n_5004 & ~n_5005;
assign n_5007 = ~n_4965 & ~n_4969;
assign n_5008 =  n_5006 & ~n_5007;
assign n_5009 = ~n_5006 &  n_5007;
assign n_5010 = ~n_5008 & ~n_5009;
assign n_5011 = ~x_1145 & ~n_5010;
assign n_5012 =  x_1145 & ~n_5009;
assign n_5013 = ~n_5008 &  n_5012;
assign n_5014 =  n_4291 & ~n_5013;
assign n_5015 = ~n_5011 &  n_5014;
assign n_5016 = ~n_5003 & ~n_5015;
assign n_5017 = ~x_4119 &  n_4974;
assign n_5018 =  x_4119 & ~n_4974;
assign n_5019 = ~n_5017 & ~n_5018;
assign n_5020 = ~n_4978 & ~n_4982;
assign n_5021 =  n_5019 & ~n_5020;
assign n_5022 = ~n_5019 &  n_5020;
assign n_5023 = ~n_5021 & ~n_5022;
assign n_5024 = ~x_4023 & ~n_5023;
assign n_5025 =  x_4023 & ~n_5022;
assign n_5026 = ~n_5021 &  n_5025;
assign n_5027 =  n_4287 & ~n_5026;
assign n_5028 = ~n_5024 &  n_5027;
assign n_5029 = ~x_698 &  n_4986;
assign n_5030 =  x_698 & ~n_4986;
assign n_5031 = ~n_5029 & ~n_5030;
assign n_5032 = ~n_4990 & ~n_4994;
assign n_5033 =  n_5031 & ~n_5032;
assign n_5034 = ~n_5031 &  n_5032;
assign n_5035 = ~n_5033 & ~n_5034;
assign n_5036 = ~x_4854 & ~n_5035;
assign n_5037 =  x_4854 & ~n_5034;
assign n_5038 = ~n_5033 &  n_5037;
assign n_5039 =  n_4292 & ~n_5038;
assign n_5040 = ~n_5036 &  n_5039;
assign n_5041 = ~n_5028 & ~n_5040;
assign n_5042 =  n_5016 &  n_5041;
assign n_5043 =  x_4343 & ~n_5042;
assign n_5044 = ~x_4343 &  n_5042;
assign n_5045 = ~n_5043 & ~n_5044;
assign n_5046 =  x_4342 &  n_4295;
assign n_5047 = ~x_3269 &  n_5004;
assign n_5048 =  x_3269 & ~n_5004;
assign n_5049 = ~n_5047 & ~n_5048;
assign n_5050 = ~n_5008 & ~n_5012;
assign n_5051 =  n_5049 & ~n_5050;
assign n_5052 = ~n_5049 &  n_5050;
assign n_5053 = ~n_5051 & ~n_5052;
assign n_5054 = ~x_1144 & ~n_5053;
assign n_5055 =  x_1144 & ~n_5052;
assign n_5056 = ~n_5051 &  n_5055;
assign n_5057 =  n_4291 & ~n_5056;
assign n_5058 = ~n_5054 &  n_5057;
assign n_5059 = ~n_5046 & ~n_5058;
assign n_5060 = ~x_4118 &  n_5017;
assign n_5061 =  x_4118 & ~n_5017;
assign n_5062 = ~n_5060 & ~n_5061;
assign n_5063 = ~n_5021 & ~n_5025;
assign n_5064 =  n_5062 & ~n_5063;
assign n_5065 = ~n_5062 &  n_5063;
assign n_5066 = ~n_5064 & ~n_5065;
assign n_5067 = ~x_4022 & ~n_5066;
assign n_5068 =  x_4022 & ~n_5065;
assign n_5069 = ~n_5064 &  n_5068;
assign n_5070 =  n_4287 & ~n_5069;
assign n_5071 = ~n_5067 &  n_5070;
assign n_5072 = ~x_697 &  n_5029;
assign n_5073 =  x_697 & ~n_5029;
assign n_5074 = ~n_5072 & ~n_5073;
assign n_5075 = ~n_5033 & ~n_5037;
assign n_5076 =  n_5074 & ~n_5075;
assign n_5077 = ~n_5074 &  n_5075;
assign n_5078 = ~n_5076 & ~n_5077;
assign n_5079 = ~x_4853 & ~n_5078;
assign n_5080 =  x_4853 & ~n_5077;
assign n_5081 = ~n_5076 &  n_5080;
assign n_5082 =  n_4292 & ~n_5081;
assign n_5083 = ~n_5079 &  n_5082;
assign n_5084 = ~n_5071 & ~n_5083;
assign n_5085 =  n_5059 &  n_5084;
assign n_5086 =  x_4342 & ~n_5085;
assign n_5087 = ~x_4342 &  n_5085;
assign n_5088 = ~n_5086 & ~n_5087;
assign n_5089 =  x_4341 &  n_4295;
assign n_5090 = ~x_3268 &  n_5047;
assign n_5091 =  x_3268 & ~n_5047;
assign n_5092 = ~n_5090 & ~n_5091;
assign n_5093 = ~n_5051 & ~n_5055;
assign n_5094 =  n_5092 & ~n_5093;
assign n_5095 = ~n_5092 &  n_5093;
assign n_5096 = ~n_5094 & ~n_5095;
assign n_5097 = ~x_1143 & ~n_5096;
assign n_5098 =  x_1143 & ~n_5095;
assign n_5099 = ~n_5094 &  n_5098;
assign n_5100 =  n_4291 & ~n_5099;
assign n_5101 = ~n_5097 &  n_5100;
assign n_5102 = ~n_5089 & ~n_5101;
assign n_5103 = ~x_4117 &  n_5060;
assign n_5104 =  x_4117 & ~n_5060;
assign n_5105 = ~n_5103 & ~n_5104;
assign n_5106 = ~n_5064 & ~n_5068;
assign n_5107 =  n_5105 & ~n_5106;
assign n_5108 = ~n_5105 &  n_5106;
assign n_5109 = ~n_5107 & ~n_5108;
assign n_5110 = ~x_4021 & ~n_5109;
assign n_5111 =  x_4021 & ~n_5108;
assign n_5112 = ~n_5107 &  n_5111;
assign n_5113 =  n_4287 & ~n_5112;
assign n_5114 = ~n_5110 &  n_5113;
assign n_5115 = ~x_696 &  n_5072;
assign n_5116 =  x_696 & ~n_5072;
assign n_5117 = ~n_5115 & ~n_5116;
assign n_5118 = ~n_5076 & ~n_5080;
assign n_5119 =  n_5117 & ~n_5118;
assign n_5120 = ~n_5117 &  n_5118;
assign n_5121 = ~n_5119 & ~n_5120;
assign n_5122 = ~x_4852 & ~n_5121;
assign n_5123 =  x_4852 & ~n_5120;
assign n_5124 = ~n_5119 &  n_5123;
assign n_5125 =  n_4292 & ~n_5124;
assign n_5126 = ~n_5122 &  n_5125;
assign n_5127 = ~n_5114 & ~n_5126;
assign n_5128 =  n_5102 &  n_5127;
assign n_5129 =  x_4341 & ~n_5128;
assign n_5130 = ~x_4341 &  n_5128;
assign n_5131 = ~n_5129 & ~n_5130;
assign n_5132 =  x_4340 &  n_4295;
assign n_5133 = ~x_3267 &  n_5090;
assign n_5134 =  x_3267 & ~n_5090;
assign n_5135 = ~n_5133 & ~n_5134;
assign n_5136 = ~n_5094 & ~n_5098;
assign n_5137 =  n_5135 & ~n_5136;
assign n_5138 = ~n_5135 &  n_5136;
assign n_5139 = ~n_5137 & ~n_5138;
assign n_5140 = ~x_1142 & ~n_5139;
assign n_5141 =  x_1142 & ~n_5138;
assign n_5142 = ~n_5137 &  n_5141;
assign n_5143 =  n_4291 & ~n_5142;
assign n_5144 = ~n_5140 &  n_5143;
assign n_5145 = ~n_5132 & ~n_5144;
assign n_5146 = ~x_4116 &  n_5103;
assign n_5147 =  x_4116 & ~n_5103;
assign n_5148 = ~n_5146 & ~n_5147;
assign n_5149 = ~n_5107 & ~n_5111;
assign n_5150 =  n_5148 & ~n_5149;
assign n_5151 = ~n_5148 &  n_5149;
assign n_5152 = ~n_5150 & ~n_5151;
assign n_5153 = ~x_4020 & ~n_5152;
assign n_5154 =  x_4020 & ~n_5151;
assign n_5155 = ~n_5150 &  n_5154;
assign n_5156 =  n_4287 & ~n_5155;
assign n_5157 = ~n_5153 &  n_5156;
assign n_5158 = ~x_695 &  n_5115;
assign n_5159 =  x_695 & ~n_5115;
assign n_5160 = ~n_5158 & ~n_5159;
assign n_5161 = ~n_5119 & ~n_5123;
assign n_5162 =  n_5160 & ~n_5161;
assign n_5163 = ~n_5160 &  n_5161;
assign n_5164 = ~n_5162 & ~n_5163;
assign n_5165 = ~x_4851 & ~n_5164;
assign n_5166 =  x_4851 & ~n_5163;
assign n_5167 = ~n_5162 &  n_5166;
assign n_5168 =  n_4292 & ~n_5167;
assign n_5169 = ~n_5165 &  n_5168;
assign n_5170 = ~n_5157 & ~n_5169;
assign n_5171 =  n_5145 &  n_5170;
assign n_5172 =  x_4340 & ~n_5171;
assign n_5173 = ~x_4340 &  n_5171;
assign n_5174 = ~n_5172 & ~n_5173;
assign n_5175 =  x_4339 &  n_4295;
assign n_5176 = ~x_3266 &  n_5133;
assign n_5177 =  x_3266 & ~n_5133;
assign n_5178 = ~n_5176 & ~n_5177;
assign n_5179 = ~n_5137 & ~n_5141;
assign n_5180 =  n_5178 & ~n_5179;
assign n_5181 = ~n_5178 &  n_5179;
assign n_5182 = ~n_5180 & ~n_5181;
assign n_5183 = ~x_1141 & ~n_5182;
assign n_5184 =  x_1141 & ~n_5181;
assign n_5185 = ~n_5180 &  n_5184;
assign n_5186 =  n_4291 & ~n_5185;
assign n_5187 = ~n_5183 &  n_5186;
assign n_5188 = ~n_5175 & ~n_5187;
assign n_5189 = ~x_4115 &  n_5146;
assign n_5190 =  x_4115 & ~n_5146;
assign n_5191 = ~n_5189 & ~n_5190;
assign n_5192 = ~n_5150 & ~n_5154;
assign n_5193 =  n_5191 & ~n_5192;
assign n_5194 = ~n_5191 &  n_5192;
assign n_5195 = ~n_5193 & ~n_5194;
assign n_5196 = ~x_4019 & ~n_5195;
assign n_5197 =  x_4019 & ~n_5194;
assign n_5198 = ~n_5193 &  n_5197;
assign n_5199 =  n_4287 & ~n_5198;
assign n_5200 = ~n_5196 &  n_5199;
assign n_5201 = ~x_694 &  n_5158;
assign n_5202 =  x_694 & ~n_5158;
assign n_5203 = ~n_5201 & ~n_5202;
assign n_5204 = ~n_5162 & ~n_5166;
assign n_5205 =  n_5203 & ~n_5204;
assign n_5206 = ~n_5203 &  n_5204;
assign n_5207 = ~n_5205 & ~n_5206;
assign n_5208 = ~x_4850 & ~n_5207;
assign n_5209 =  x_4850 & ~n_5206;
assign n_5210 = ~n_5205 &  n_5209;
assign n_5211 =  n_4292 & ~n_5210;
assign n_5212 = ~n_5208 &  n_5211;
assign n_5213 = ~n_5200 & ~n_5212;
assign n_5214 =  n_5188 &  n_5213;
assign n_5215 =  x_4339 & ~n_5214;
assign n_5216 = ~x_4339 &  n_5214;
assign n_5217 = ~n_5215 & ~n_5216;
assign n_5218 =  x_4338 &  n_4295;
assign n_5219 = ~x_3265 &  n_5176;
assign n_5220 =  x_3265 & ~n_5176;
assign n_5221 = ~n_5219 & ~n_5220;
assign n_5222 = ~n_5180 & ~n_5184;
assign n_5223 =  n_5221 & ~n_5222;
assign n_5224 = ~n_5221 &  n_5222;
assign n_5225 = ~n_5223 & ~n_5224;
assign n_5226 = ~x_1140 & ~n_5225;
assign n_5227 =  x_1140 & ~n_5224;
assign n_5228 = ~n_5223 &  n_5227;
assign n_5229 =  n_4291 & ~n_5228;
assign n_5230 = ~n_5226 &  n_5229;
assign n_5231 = ~n_5218 & ~n_5230;
assign n_5232 = ~x_4114 &  n_5189;
assign n_5233 =  x_4114 & ~n_5189;
assign n_5234 = ~n_5232 & ~n_5233;
assign n_5235 = ~n_5193 & ~n_5197;
assign n_5236 =  n_5234 & ~n_5235;
assign n_5237 = ~n_5234 &  n_5235;
assign n_5238 = ~n_5236 & ~n_5237;
assign n_5239 = ~x_4018 & ~n_5238;
assign n_5240 =  x_4018 & ~n_5237;
assign n_5241 = ~n_5236 &  n_5240;
assign n_5242 =  n_4287 & ~n_5241;
assign n_5243 = ~n_5239 &  n_5242;
assign n_5244 = ~x_693 &  n_5201;
assign n_5245 =  x_693 & ~n_5201;
assign n_5246 = ~n_5244 & ~n_5245;
assign n_5247 = ~n_5205 & ~n_5209;
assign n_5248 =  n_5246 & ~n_5247;
assign n_5249 = ~n_5246 &  n_5247;
assign n_5250 = ~n_5248 & ~n_5249;
assign n_5251 = ~x_4849 & ~n_5250;
assign n_5252 =  x_4849 & ~n_5249;
assign n_5253 = ~n_5248 &  n_5252;
assign n_5254 =  n_4292 & ~n_5253;
assign n_5255 = ~n_5251 &  n_5254;
assign n_5256 = ~n_5243 & ~n_5255;
assign n_5257 =  n_5231 &  n_5256;
assign n_5258 =  x_4338 & ~n_5257;
assign n_5259 = ~x_4338 &  n_5257;
assign n_5260 = ~n_5258 & ~n_5259;
assign n_5261 =  x_4337 &  n_4295;
assign n_5262 = ~x_3264 &  n_5219;
assign n_5263 =  x_3264 & ~n_5219;
assign n_5264 = ~n_5262 & ~n_5263;
assign n_5265 = ~n_5223 & ~n_5227;
assign n_5266 =  n_5264 & ~n_5265;
assign n_5267 = ~n_5264 &  n_5265;
assign n_5268 = ~n_5266 & ~n_5267;
assign n_5269 = ~x_1139 & ~n_5268;
assign n_5270 =  x_1139 & ~n_5267;
assign n_5271 = ~n_5266 &  n_5270;
assign n_5272 =  n_4291 & ~n_5271;
assign n_5273 = ~n_5269 &  n_5272;
assign n_5274 = ~n_5261 & ~n_5273;
assign n_5275 = ~x_4113 &  n_5232;
assign n_5276 =  x_4113 & ~n_5232;
assign n_5277 = ~n_5275 & ~n_5276;
assign n_5278 = ~n_5236 & ~n_5240;
assign n_5279 =  n_5277 & ~n_5278;
assign n_5280 = ~n_5277 &  n_5278;
assign n_5281 = ~n_5279 & ~n_5280;
assign n_5282 = ~x_4017 & ~n_5281;
assign n_5283 =  x_4017 & ~n_5280;
assign n_5284 = ~n_5279 &  n_5283;
assign n_5285 =  n_4287 & ~n_5284;
assign n_5286 = ~n_5282 &  n_5285;
assign n_5287 = ~x_692 &  n_5244;
assign n_5288 =  x_692 & ~n_5244;
assign n_5289 = ~n_5287 & ~n_5288;
assign n_5290 = ~n_5248 & ~n_5252;
assign n_5291 =  n_5289 & ~n_5290;
assign n_5292 = ~n_5289 &  n_5290;
assign n_5293 = ~n_5291 & ~n_5292;
assign n_5294 = ~x_4848 & ~n_5293;
assign n_5295 =  x_4848 & ~n_5292;
assign n_5296 = ~n_5291 &  n_5295;
assign n_5297 =  n_4292 & ~n_5296;
assign n_5298 = ~n_5294 &  n_5297;
assign n_5299 = ~n_5286 & ~n_5298;
assign n_5300 =  n_5274 &  n_5299;
assign n_5301 =  x_4337 & ~n_5300;
assign n_5302 = ~x_4337 &  n_5300;
assign n_5303 = ~n_5301 & ~n_5302;
assign n_5304 =  x_4336 &  n_4295;
assign n_5305 = ~x_3263 &  n_5262;
assign n_5306 =  x_3263 & ~n_5262;
assign n_5307 = ~n_5305 & ~n_5306;
assign n_5308 = ~n_5266 & ~n_5270;
assign n_5309 =  n_5307 & ~n_5308;
assign n_5310 = ~n_5307 &  n_5308;
assign n_5311 = ~n_5309 & ~n_5310;
assign n_5312 = ~x_1138 & ~n_5311;
assign n_5313 =  x_1138 & ~n_5310;
assign n_5314 = ~n_5309 &  n_5313;
assign n_5315 =  n_4291 & ~n_5314;
assign n_5316 = ~n_5312 &  n_5315;
assign n_5317 = ~n_5304 & ~n_5316;
assign n_5318 = ~x_4112 &  n_5275;
assign n_5319 =  x_4112 & ~n_5275;
assign n_5320 = ~n_5318 & ~n_5319;
assign n_5321 = ~n_5279 & ~n_5283;
assign n_5322 =  n_5320 & ~n_5321;
assign n_5323 = ~n_5320 &  n_5321;
assign n_5324 = ~n_5322 & ~n_5323;
assign n_5325 = ~x_4016 & ~n_5324;
assign n_5326 =  x_4016 & ~n_5323;
assign n_5327 = ~n_5322 &  n_5326;
assign n_5328 =  n_4287 & ~n_5327;
assign n_5329 = ~n_5325 &  n_5328;
assign n_5330 = ~x_691 &  n_5287;
assign n_5331 =  x_691 & ~n_5287;
assign n_5332 = ~n_5330 & ~n_5331;
assign n_5333 = ~n_5291 & ~n_5295;
assign n_5334 =  n_5332 & ~n_5333;
assign n_5335 = ~n_5332 &  n_5333;
assign n_5336 = ~n_5334 & ~n_5335;
assign n_5337 = ~x_4847 & ~n_5336;
assign n_5338 =  x_4847 & ~n_5335;
assign n_5339 = ~n_5334 &  n_5338;
assign n_5340 =  n_4292 & ~n_5339;
assign n_5341 = ~n_5337 &  n_5340;
assign n_5342 = ~n_5329 & ~n_5341;
assign n_5343 =  n_5317 &  n_5342;
assign n_5344 =  x_4336 & ~n_5343;
assign n_5345 = ~x_4336 &  n_5343;
assign n_5346 = ~n_5344 & ~n_5345;
assign n_5347 =  x_4335 &  n_4295;
assign n_5348 = ~x_3262 &  n_5305;
assign n_5349 =  x_3262 & ~n_5305;
assign n_5350 = ~n_5348 & ~n_5349;
assign n_5351 = ~n_5309 & ~n_5313;
assign n_5352 =  n_5350 & ~n_5351;
assign n_5353 = ~n_5350 &  n_5351;
assign n_5354 = ~n_5352 & ~n_5353;
assign n_5355 = ~x_1137 & ~n_5354;
assign n_5356 =  x_1137 & ~n_5353;
assign n_5357 = ~n_5352 &  n_5356;
assign n_5358 =  n_4291 & ~n_5357;
assign n_5359 = ~n_5355 &  n_5358;
assign n_5360 = ~n_5347 & ~n_5359;
assign n_5361 = ~x_4111 &  n_5318;
assign n_5362 =  x_4111 & ~n_5318;
assign n_5363 = ~n_5361 & ~n_5362;
assign n_5364 = ~n_5322 & ~n_5326;
assign n_5365 =  n_5363 & ~n_5364;
assign n_5366 = ~n_5363 &  n_5364;
assign n_5367 = ~n_5365 & ~n_5366;
assign n_5368 = ~x_4015 & ~n_5367;
assign n_5369 =  x_4015 & ~n_5366;
assign n_5370 = ~n_5365 &  n_5369;
assign n_5371 =  n_4287 & ~n_5370;
assign n_5372 = ~n_5368 &  n_5371;
assign n_5373 = ~x_690 &  n_5330;
assign n_5374 =  x_690 & ~n_5330;
assign n_5375 = ~n_5373 & ~n_5374;
assign n_5376 = ~n_5334 & ~n_5338;
assign n_5377 =  n_5375 & ~n_5376;
assign n_5378 = ~n_5375 &  n_5376;
assign n_5379 = ~n_5377 & ~n_5378;
assign n_5380 = ~x_4846 & ~n_5379;
assign n_5381 =  x_4846 & ~n_5378;
assign n_5382 = ~n_5377 &  n_5381;
assign n_5383 =  n_4292 & ~n_5382;
assign n_5384 = ~n_5380 &  n_5383;
assign n_5385 = ~n_5372 & ~n_5384;
assign n_5386 =  n_5360 &  n_5385;
assign n_5387 =  x_4335 & ~n_5386;
assign n_5388 = ~x_4335 &  n_5386;
assign n_5389 = ~n_5387 & ~n_5388;
assign n_5390 =  x_4334 &  n_4295;
assign n_5391 = ~x_3261 &  n_5348;
assign n_5392 =  x_3261 & ~n_5348;
assign n_5393 = ~n_5391 & ~n_5392;
assign n_5394 = ~n_5352 & ~n_5356;
assign n_5395 =  n_5393 & ~n_5394;
assign n_5396 = ~n_5393 &  n_5394;
assign n_5397 = ~n_5395 & ~n_5396;
assign n_5398 = ~x_1136 & ~n_5397;
assign n_5399 =  x_1136 & ~n_5396;
assign n_5400 = ~n_5395 &  n_5399;
assign n_5401 =  n_4291 & ~n_5400;
assign n_5402 = ~n_5398 &  n_5401;
assign n_5403 = ~n_5390 & ~n_5402;
assign n_5404 = ~x_4110 &  n_5361;
assign n_5405 =  x_4110 & ~n_5361;
assign n_5406 = ~n_5404 & ~n_5405;
assign n_5407 = ~n_5365 & ~n_5369;
assign n_5408 =  n_5406 & ~n_5407;
assign n_5409 = ~n_5406 &  n_5407;
assign n_5410 = ~n_5408 & ~n_5409;
assign n_5411 = ~x_4014 & ~n_5410;
assign n_5412 =  x_4014 & ~n_5409;
assign n_5413 = ~n_5408 &  n_5412;
assign n_5414 =  n_4287 & ~n_5413;
assign n_5415 = ~n_5411 &  n_5414;
assign n_5416 = ~x_689 &  n_5373;
assign n_5417 =  x_689 & ~n_5373;
assign n_5418 = ~n_5416 & ~n_5417;
assign n_5419 = ~n_5377 & ~n_5381;
assign n_5420 =  n_5418 & ~n_5419;
assign n_5421 = ~n_5418 &  n_5419;
assign n_5422 = ~n_5420 & ~n_5421;
assign n_5423 = ~x_4845 & ~n_5422;
assign n_5424 =  x_4845 & ~n_5421;
assign n_5425 = ~n_5420 &  n_5424;
assign n_5426 =  n_4292 & ~n_5425;
assign n_5427 = ~n_5423 &  n_5426;
assign n_5428 = ~n_5415 & ~n_5427;
assign n_5429 =  n_5403 &  n_5428;
assign n_5430 =  x_4334 & ~n_5429;
assign n_5431 = ~x_4334 &  n_5429;
assign n_5432 = ~n_5430 & ~n_5431;
assign n_5433 =  x_4333 &  n_4295;
assign n_5434 = ~x_3260 &  n_5391;
assign n_5435 =  x_3260 & ~n_5391;
assign n_5436 = ~n_5434 & ~n_5435;
assign n_5437 = ~n_5395 & ~n_5399;
assign n_5438 =  n_5436 & ~n_5437;
assign n_5439 = ~n_5436 &  n_5437;
assign n_5440 = ~n_5438 & ~n_5439;
assign n_5441 = ~x_1135 & ~n_5440;
assign n_5442 =  x_1135 & ~n_5439;
assign n_5443 = ~n_5438 &  n_5442;
assign n_5444 =  n_4291 & ~n_5443;
assign n_5445 = ~n_5441 &  n_5444;
assign n_5446 = ~n_5433 & ~n_5445;
assign n_5447 = ~x_4109 &  n_5404;
assign n_5448 =  x_4109 & ~n_5404;
assign n_5449 = ~n_5447 & ~n_5448;
assign n_5450 = ~n_5408 & ~n_5412;
assign n_5451 =  n_5449 & ~n_5450;
assign n_5452 = ~n_5449 &  n_5450;
assign n_5453 = ~n_5451 & ~n_5452;
assign n_5454 = ~x_4013 & ~n_5453;
assign n_5455 =  x_4013 & ~n_5452;
assign n_5456 = ~n_5451 &  n_5455;
assign n_5457 =  n_4287 & ~n_5456;
assign n_5458 = ~n_5454 &  n_5457;
assign n_5459 = ~x_688 &  n_5416;
assign n_5460 =  x_688 & ~n_5416;
assign n_5461 = ~n_5459 & ~n_5460;
assign n_5462 = ~n_5420 & ~n_5424;
assign n_5463 =  n_5461 & ~n_5462;
assign n_5464 = ~n_5461 &  n_5462;
assign n_5465 = ~n_5463 & ~n_5464;
assign n_5466 = ~x_4844 & ~n_5465;
assign n_5467 =  x_4844 & ~n_5464;
assign n_5468 = ~n_5463 &  n_5467;
assign n_5469 =  n_4292 & ~n_5468;
assign n_5470 = ~n_5466 &  n_5469;
assign n_5471 = ~n_5458 & ~n_5470;
assign n_5472 =  n_5446 &  n_5471;
assign n_5473 =  x_4333 & ~n_5472;
assign n_5474 = ~x_4333 &  n_5472;
assign n_5475 = ~n_5473 & ~n_5474;
assign n_5476 =  x_4332 &  n_4295;
assign n_5477 = ~x_3259 &  n_5434;
assign n_5478 =  x_3259 & ~n_5434;
assign n_5479 = ~n_5477 & ~n_5478;
assign n_5480 = ~n_5438 & ~n_5442;
assign n_5481 =  n_5479 & ~n_5480;
assign n_5482 = ~n_5479 &  n_5480;
assign n_5483 = ~n_5481 & ~n_5482;
assign n_5484 = ~x_1134 & ~n_5483;
assign n_5485 =  x_1134 & ~n_5482;
assign n_5486 = ~n_5481 &  n_5485;
assign n_5487 =  n_4291 & ~n_5486;
assign n_5488 = ~n_5484 &  n_5487;
assign n_5489 = ~n_5476 & ~n_5488;
assign n_5490 = ~x_4108 &  n_5447;
assign n_5491 =  x_4108 & ~n_5447;
assign n_5492 = ~n_5490 & ~n_5491;
assign n_5493 = ~n_5451 & ~n_5455;
assign n_5494 =  n_5492 & ~n_5493;
assign n_5495 = ~n_5492 &  n_5493;
assign n_5496 = ~n_5494 & ~n_5495;
assign n_5497 = ~x_4012 & ~n_5496;
assign n_5498 =  x_4012 & ~n_5495;
assign n_5499 = ~n_5494 &  n_5498;
assign n_5500 =  n_4287 & ~n_5499;
assign n_5501 = ~n_5497 &  n_5500;
assign n_5502 = ~x_687 &  n_5459;
assign n_5503 =  x_687 & ~n_5459;
assign n_5504 = ~n_5502 & ~n_5503;
assign n_5505 = ~n_5463 & ~n_5467;
assign n_5506 =  n_5504 & ~n_5505;
assign n_5507 = ~n_5504 &  n_5505;
assign n_5508 = ~n_5506 & ~n_5507;
assign n_5509 = ~x_4843 & ~n_5508;
assign n_5510 =  x_4843 & ~n_5507;
assign n_5511 = ~n_5506 &  n_5510;
assign n_5512 =  n_4292 & ~n_5511;
assign n_5513 = ~n_5509 &  n_5512;
assign n_5514 = ~n_5501 & ~n_5513;
assign n_5515 =  n_5489 &  n_5514;
assign n_5516 =  x_4332 & ~n_5515;
assign n_5517 = ~x_4332 &  n_5515;
assign n_5518 = ~n_5516 & ~n_5517;
assign n_5519 =  x_4331 &  n_4295;
assign n_5520 = ~x_3258 &  n_5477;
assign n_5521 =  x_3258 & ~n_5477;
assign n_5522 = ~n_5520 & ~n_5521;
assign n_5523 = ~n_5481 & ~n_5485;
assign n_5524 =  n_5522 & ~n_5523;
assign n_5525 = ~n_5522 &  n_5523;
assign n_5526 = ~n_5524 & ~n_5525;
assign n_5527 = ~x_1133 & ~n_5526;
assign n_5528 =  x_1133 & ~n_5525;
assign n_5529 = ~n_5524 &  n_5528;
assign n_5530 =  n_4291 & ~n_5529;
assign n_5531 = ~n_5527 &  n_5530;
assign n_5532 = ~n_5519 & ~n_5531;
assign n_5533 = ~x_4107 &  n_5490;
assign n_5534 =  x_4107 & ~n_5490;
assign n_5535 = ~n_5533 & ~n_5534;
assign n_5536 = ~n_5494 & ~n_5498;
assign n_5537 =  n_5535 & ~n_5536;
assign n_5538 = ~n_5535 &  n_5536;
assign n_5539 = ~n_5537 & ~n_5538;
assign n_5540 = ~x_4011 & ~n_5539;
assign n_5541 =  x_4011 & ~n_5538;
assign n_5542 = ~n_5537 &  n_5541;
assign n_5543 =  n_4287 & ~n_5542;
assign n_5544 = ~n_5540 &  n_5543;
assign n_5545 = ~x_686 &  n_5502;
assign n_5546 =  x_686 & ~n_5502;
assign n_5547 = ~n_5545 & ~n_5546;
assign n_5548 = ~n_5506 & ~n_5510;
assign n_5549 =  n_5547 & ~n_5548;
assign n_5550 = ~n_5547 &  n_5548;
assign n_5551 = ~n_5549 & ~n_5550;
assign n_5552 = ~x_4842 & ~n_5551;
assign n_5553 =  x_4842 & ~n_5550;
assign n_5554 = ~n_5549 &  n_5553;
assign n_5555 =  n_4292 & ~n_5554;
assign n_5556 = ~n_5552 &  n_5555;
assign n_5557 = ~n_5544 & ~n_5556;
assign n_5558 =  n_5532 &  n_5557;
assign n_5559 =  x_4331 & ~n_5558;
assign n_5560 = ~x_4331 &  n_5558;
assign n_5561 = ~n_5559 & ~n_5560;
assign n_5562 =  x_4330 &  n_4295;
assign n_5563 = ~x_3257 &  n_5520;
assign n_5564 =  x_3257 & ~n_5520;
assign n_5565 = ~n_5563 & ~n_5564;
assign n_5566 = ~n_5524 & ~n_5528;
assign n_5567 =  n_5565 & ~n_5566;
assign n_5568 = ~n_5565 &  n_5566;
assign n_5569 = ~n_5567 & ~n_5568;
assign n_5570 = ~x_1132 & ~n_5569;
assign n_5571 =  x_1132 & ~n_5568;
assign n_5572 = ~n_5567 &  n_5571;
assign n_5573 =  n_4291 & ~n_5572;
assign n_5574 = ~n_5570 &  n_5573;
assign n_5575 = ~n_5562 & ~n_5574;
assign n_5576 = ~x_4106 &  n_5533;
assign n_5577 =  x_4106 & ~n_5533;
assign n_5578 = ~n_5576 & ~n_5577;
assign n_5579 = ~n_5537 & ~n_5541;
assign n_5580 =  n_5578 & ~n_5579;
assign n_5581 = ~n_5578 &  n_5579;
assign n_5582 = ~n_5580 & ~n_5581;
assign n_5583 = ~x_4010 & ~n_5582;
assign n_5584 =  x_4010 & ~n_5581;
assign n_5585 = ~n_5580 &  n_5584;
assign n_5586 =  n_4287 & ~n_5585;
assign n_5587 = ~n_5583 &  n_5586;
assign n_5588 = ~x_685 &  n_5545;
assign n_5589 =  x_685 & ~n_5545;
assign n_5590 = ~n_5588 & ~n_5589;
assign n_5591 = ~n_5549 & ~n_5553;
assign n_5592 =  n_5590 & ~n_5591;
assign n_5593 = ~n_5590 &  n_5591;
assign n_5594 = ~n_5592 & ~n_5593;
assign n_5595 = ~x_4841 & ~n_5594;
assign n_5596 =  x_4841 & ~n_5593;
assign n_5597 = ~n_5592 &  n_5596;
assign n_5598 =  n_4292 & ~n_5597;
assign n_5599 = ~n_5595 &  n_5598;
assign n_5600 = ~n_5587 & ~n_5599;
assign n_5601 =  n_5575 &  n_5600;
assign n_5602 =  x_4330 & ~n_5601;
assign n_5603 = ~x_4330 &  n_5601;
assign n_5604 = ~n_5602 & ~n_5603;
assign n_5605 =  x_4329 &  n_4295;
assign n_5606 = ~n_5592 & ~n_5596;
assign n_5607 =  x_684 & ~x_4840;
assign n_5608 = ~x_684 &  x_4840;
assign n_5609 = ~n_5607 & ~n_5608;
assign n_5610 =  n_5588 &  n_5609;
assign n_5611 = ~n_5588 & ~n_5609;
assign n_5612 = ~n_5610 & ~n_5611;
assign n_5613 =  n_5606 & ~n_5612;
assign n_5614 = ~n_5606 &  n_5612;
assign n_5615 =  n_4292 & ~n_5614;
assign n_5616 = ~n_5613 &  n_5615;
assign n_5617 = ~n_5605 & ~n_5616;
assign n_5618 = ~n_5567 & ~n_5571;
assign n_5619 =  x_1131 & ~x_3256;
assign n_5620 = ~x_1131 &  x_3256;
assign n_5621 = ~n_5619 & ~n_5620;
assign n_5622 =  n_5563 &  n_5621;
assign n_5623 = ~n_5563 & ~n_5621;
assign n_5624 = ~n_5622 & ~n_5623;
assign n_5625 =  n_5618 & ~n_5624;
assign n_5626 = ~n_5618 &  n_5624;
assign n_5627 =  n_4291 & ~n_5626;
assign n_5628 = ~n_5625 &  n_5627;
assign n_5629 = ~n_5580 & ~n_5584;
assign n_5630 =  x_4009 & ~x_4105;
assign n_5631 = ~x_4009 &  x_4105;
assign n_5632 = ~n_5630 & ~n_5631;
assign n_5633 =  n_5576 &  n_5632;
assign n_5634 = ~n_5576 & ~n_5632;
assign n_5635 = ~n_5633 & ~n_5634;
assign n_5636 =  n_5629 & ~n_5635;
assign n_5637 = ~n_5629 &  n_5635;
assign n_5638 =  n_4287 & ~n_5637;
assign n_5639 = ~n_5636 &  n_5638;
assign n_5640 = ~n_5628 & ~n_5639;
assign n_5641 =  n_5617 &  n_5640;
assign n_5642 =  x_4329 & ~n_5641;
assign n_5643 = ~x_4329 &  n_5641;
assign n_5644 = ~n_5642 & ~n_5643;
assign n_5645 = ~x_43 &  n_3341;
assign n_5646 =  n_1305 &  n_1173;
assign n_5647 =  n_5645 &  n_5646;
assign n_5648 =  x_40 &  n_151;
assign n_5649 =  n_150 &  n_5648;
assign n_5650 =  n_3143 &  n_5649;
assign n_5651 = ~x_38 &  n_6;
assign n_5652 =  n_1038 &  n_5651;
assign n_5653 =  n_150 &  n_5652;
assign n_5654 = ~x_42 &  x_43;
assign n_5655 =  x_41 &  n_759;
assign n_5656 =  n_5654 &  n_5655;
assign n_5657 =  n_1173 &  n_5656;
assign n_5658 = ~n_5653 & ~n_5657;
assign n_5659 = ~n_5650 &  n_5658;
assign n_5660 = ~n_5647 &  n_5659;
assign n_5661 =  x_4328 &  n_5660;
assign n_5662 =  x_3319 &  n_5647;
assign n_5663 =  x_4392 &  n_5657;
assign n_5664 =  x_5031 &  n_5650;
assign n_5665 = ~n_5663 & ~n_5664;
assign n_5666 = ~n_5662 &  n_5665;
assign n_5667 = ~n_5661 &  n_5666;
assign n_5668 =  x_4328 & ~n_5667;
assign n_5669 = ~x_4328 &  n_5667;
assign n_5670 = ~n_5668 & ~n_5669;
assign n_5671 =  x_4327 &  n_5660;
assign n_5672 =  x_3318 &  n_5647;
assign n_5673 =  x_4391 &  n_5657;
assign n_5674 =  x_5030 &  n_5650;
assign n_5675 = ~n_5673 & ~n_5674;
assign n_5676 = ~n_5672 &  n_5675;
assign n_5677 = ~n_5671 &  n_5676;
assign n_5678 =  x_4327 & ~n_5677;
assign n_5679 = ~x_4327 &  n_5677;
assign n_5680 = ~n_5678 & ~n_5679;
assign n_5681 =  x_4326 &  n_5660;
assign n_5682 =  x_3317 &  n_5647;
assign n_5683 =  x_4390 &  n_5657;
assign n_5684 =  x_5029 &  n_5650;
assign n_5685 = ~n_5683 & ~n_5684;
assign n_5686 = ~n_5682 &  n_5685;
assign n_5687 = ~n_5681 &  n_5686;
assign n_5688 =  x_4326 & ~n_5687;
assign n_5689 = ~x_4326 &  n_5687;
assign n_5690 = ~n_5688 & ~n_5689;
assign n_5691 =  x_4325 &  n_5660;
assign n_5692 =  x_3316 &  n_5647;
assign n_5693 =  x_4389 &  n_5657;
assign n_5694 =  x_5028 &  n_5650;
assign n_5695 = ~n_5693 & ~n_5694;
assign n_5696 = ~n_5692 &  n_5695;
assign n_5697 = ~n_5691 &  n_5696;
assign n_5698 =  x_4325 & ~n_5697;
assign n_5699 = ~x_4325 &  n_5697;
assign n_5700 = ~n_5698 & ~n_5699;
assign n_5701 =  x_4324 &  n_5660;
assign n_5702 =  x_3315 &  n_5647;
assign n_5703 =  x_4388 &  n_5657;
assign n_5704 =  x_5027 &  n_5650;
assign n_5705 = ~n_5703 & ~n_5704;
assign n_5706 = ~n_5702 &  n_5705;
assign n_5707 = ~n_5701 &  n_5706;
assign n_5708 =  x_4324 & ~n_5707;
assign n_5709 = ~x_4324 &  n_5707;
assign n_5710 = ~n_5708 & ~n_5709;
assign n_5711 =  x_4323 &  n_5660;
assign n_5712 =  x_3314 &  n_5647;
assign n_5713 =  x_4387 &  n_5657;
assign n_5714 =  x_5026 &  n_5650;
assign n_5715 = ~n_5713 & ~n_5714;
assign n_5716 = ~n_5712 &  n_5715;
assign n_5717 = ~n_5711 &  n_5716;
assign n_5718 =  x_4323 & ~n_5717;
assign n_5719 = ~x_4323 &  n_5717;
assign n_5720 = ~n_5718 & ~n_5719;
assign n_5721 =  x_4322 &  n_5660;
assign n_5722 =  x_3313 &  n_5647;
assign n_5723 =  x_4386 &  n_5657;
assign n_5724 =  x_5025 &  n_5650;
assign n_5725 = ~n_5723 & ~n_5724;
assign n_5726 = ~n_5722 &  n_5725;
assign n_5727 = ~n_5721 &  n_5726;
assign n_5728 =  x_4322 & ~n_5727;
assign n_5729 = ~x_4322 &  n_5727;
assign n_5730 = ~n_5728 & ~n_5729;
assign n_5731 =  x_4321 &  n_5660;
assign n_5732 =  x_3312 &  n_5647;
assign n_5733 =  x_4385 &  n_5657;
assign n_5734 =  x_5024 &  n_5650;
assign n_5735 = ~n_5733 & ~n_5734;
assign n_5736 = ~n_5732 &  n_5735;
assign n_5737 = ~n_5731 &  n_5736;
assign n_5738 =  x_4321 & ~n_5737;
assign n_5739 = ~x_4321 &  n_5737;
assign n_5740 = ~n_5738 & ~n_5739;
assign n_5741 =  x_4320 &  n_5660;
assign n_5742 =  x_3311 &  n_5647;
assign n_5743 =  x_4384 &  n_5657;
assign n_5744 =  x_5023 &  n_5650;
assign n_5745 = ~n_5743 & ~n_5744;
assign n_5746 = ~n_5742 &  n_5745;
assign n_5747 = ~n_5741 &  n_5746;
assign n_5748 =  x_4320 & ~n_5747;
assign n_5749 = ~x_4320 &  n_5747;
assign n_5750 = ~n_5748 & ~n_5749;
assign n_5751 =  x_4319 &  n_5660;
assign n_5752 =  x_3310 &  n_5647;
assign n_5753 =  x_4383 &  n_5657;
assign n_5754 =  x_5022 &  n_5650;
assign n_5755 = ~n_5753 & ~n_5754;
assign n_5756 = ~n_5752 &  n_5755;
assign n_5757 = ~n_5751 &  n_5756;
assign n_5758 =  x_4319 & ~n_5757;
assign n_5759 = ~x_4319 &  n_5757;
assign n_5760 = ~n_5758 & ~n_5759;
assign n_5761 =  x_4318 &  n_5660;
assign n_5762 =  x_3309 &  n_5647;
assign n_5763 =  x_4382 &  n_5657;
assign n_5764 =  x_5021 &  n_5650;
assign n_5765 = ~n_5763 & ~n_5764;
assign n_5766 = ~n_5762 &  n_5765;
assign n_5767 = ~n_5761 &  n_5766;
assign n_5768 =  x_4318 & ~n_5767;
assign n_5769 = ~x_4318 &  n_5767;
assign n_5770 = ~n_5768 & ~n_5769;
assign n_5771 =  x_4317 &  n_5660;
assign n_5772 =  x_3308 &  n_5647;
assign n_5773 =  x_4381 &  n_5657;
assign n_5774 =  x_5020 &  n_5650;
assign n_5775 = ~n_5773 & ~n_5774;
assign n_5776 = ~n_5772 &  n_5775;
assign n_5777 = ~n_5771 &  n_5776;
assign n_5778 =  x_4317 & ~n_5777;
assign n_5779 = ~x_4317 &  n_5777;
assign n_5780 = ~n_5778 & ~n_5779;
assign n_5781 =  x_4316 &  n_5660;
assign n_5782 =  x_3307 &  n_5647;
assign n_5783 =  x_4380 &  n_5657;
assign n_5784 =  x_5019 &  n_5650;
assign n_5785 = ~n_5783 & ~n_5784;
assign n_5786 = ~n_5782 &  n_5785;
assign n_5787 = ~n_5781 &  n_5786;
assign n_5788 =  x_4316 & ~n_5787;
assign n_5789 = ~x_4316 &  n_5787;
assign n_5790 = ~n_5788 & ~n_5789;
assign n_5791 =  x_4315 &  n_5660;
assign n_5792 =  x_3306 &  n_5647;
assign n_5793 =  x_4379 &  n_5657;
assign n_5794 =  x_5018 &  n_5650;
assign n_5795 = ~n_5793 & ~n_5794;
assign n_5796 = ~n_5792 &  n_5795;
assign n_5797 = ~n_5791 &  n_5796;
assign n_5798 =  x_4315 & ~n_5797;
assign n_5799 = ~x_4315 &  n_5797;
assign n_5800 = ~n_5798 & ~n_5799;
assign n_5801 =  x_4314 &  n_5660;
assign n_5802 =  x_3305 &  n_5647;
assign n_5803 =  x_4378 &  n_5657;
assign n_5804 =  x_5017 &  n_5650;
assign n_5805 = ~n_5803 & ~n_5804;
assign n_5806 = ~n_5802 &  n_5805;
assign n_5807 = ~n_5801 &  n_5806;
assign n_5808 =  x_4314 & ~n_5807;
assign n_5809 = ~x_4314 &  n_5807;
assign n_5810 = ~n_5808 & ~n_5809;
assign n_5811 =  x_4313 &  n_5660;
assign n_5812 =  x_3304 &  n_5647;
assign n_5813 =  x_4377 &  n_5657;
assign n_5814 =  x_5016 &  n_5650;
assign n_5815 = ~n_5813 & ~n_5814;
assign n_5816 = ~n_5812 &  n_5815;
assign n_5817 = ~n_5811 &  n_5816;
assign n_5818 =  x_4313 & ~n_5817;
assign n_5819 = ~x_4313 &  n_5817;
assign n_5820 = ~n_5818 & ~n_5819;
assign n_5821 =  x_4312 &  n_5660;
assign n_5822 =  x_3303 &  n_5647;
assign n_5823 =  x_4376 &  n_5657;
assign n_5824 =  x_5015 &  n_5650;
assign n_5825 = ~n_5823 & ~n_5824;
assign n_5826 = ~n_5822 &  n_5825;
assign n_5827 = ~n_5821 &  n_5826;
assign n_5828 =  x_4312 & ~n_5827;
assign n_5829 = ~x_4312 &  n_5827;
assign n_5830 = ~n_5828 & ~n_5829;
assign n_5831 =  x_4311 &  n_5660;
assign n_5832 =  x_3302 &  n_5647;
assign n_5833 =  x_4375 &  n_5657;
assign n_5834 =  x_5014 &  n_5650;
assign n_5835 = ~n_5833 & ~n_5834;
assign n_5836 = ~n_5832 &  n_5835;
assign n_5837 = ~n_5831 &  n_5836;
assign n_5838 =  x_4311 & ~n_5837;
assign n_5839 = ~x_4311 &  n_5837;
assign n_5840 = ~n_5838 & ~n_5839;
assign n_5841 =  x_4310 &  n_5660;
assign n_5842 =  x_3301 &  n_5647;
assign n_5843 =  x_4374 &  n_5657;
assign n_5844 =  x_5013 &  n_5650;
assign n_5845 = ~n_5843 & ~n_5844;
assign n_5846 = ~n_5842 &  n_5845;
assign n_5847 = ~n_5841 &  n_5846;
assign n_5848 =  x_4310 & ~n_5847;
assign n_5849 = ~x_4310 &  n_5847;
assign n_5850 = ~n_5848 & ~n_5849;
assign n_5851 =  x_4309 &  n_5660;
assign n_5852 =  x_3300 &  n_5647;
assign n_5853 =  x_4373 &  n_5657;
assign n_5854 =  x_5012 &  n_5650;
assign n_5855 = ~n_5853 & ~n_5854;
assign n_5856 = ~n_5852 &  n_5855;
assign n_5857 = ~n_5851 &  n_5856;
assign n_5858 =  x_4309 & ~n_5857;
assign n_5859 = ~x_4309 &  n_5857;
assign n_5860 = ~n_5858 & ~n_5859;
assign n_5861 =  x_4308 &  n_5660;
assign n_5862 =  x_3299 &  n_5647;
assign n_5863 =  x_4372 &  n_5657;
assign n_5864 =  x_5011 &  n_5650;
assign n_5865 = ~n_5863 & ~n_5864;
assign n_5866 = ~n_5862 &  n_5865;
assign n_5867 = ~n_5861 &  n_5866;
assign n_5868 =  x_4308 & ~n_5867;
assign n_5869 = ~x_4308 &  n_5867;
assign n_5870 = ~n_5868 & ~n_5869;
assign n_5871 =  x_4307 &  n_5660;
assign n_5872 =  x_3298 &  n_5647;
assign n_5873 =  x_4371 &  n_5657;
assign n_5874 =  x_5010 &  n_5650;
assign n_5875 = ~n_5873 & ~n_5874;
assign n_5876 = ~n_5872 &  n_5875;
assign n_5877 = ~n_5871 &  n_5876;
assign n_5878 =  x_4307 & ~n_5877;
assign n_5879 = ~x_4307 &  n_5877;
assign n_5880 = ~n_5878 & ~n_5879;
assign n_5881 =  x_4306 &  n_5660;
assign n_5882 =  x_3297 &  n_5647;
assign n_5883 =  x_4370 &  n_5657;
assign n_5884 =  x_5009 &  n_5650;
assign n_5885 = ~n_5883 & ~n_5884;
assign n_5886 = ~n_5882 &  n_5885;
assign n_5887 = ~n_5881 &  n_5886;
assign n_5888 =  x_4306 & ~n_5887;
assign n_5889 = ~x_4306 &  n_5887;
assign n_5890 = ~n_5888 & ~n_5889;
assign n_5891 =  x_4305 &  n_5660;
assign n_5892 =  x_3296 &  n_5647;
assign n_5893 =  x_4369 &  n_5657;
assign n_5894 =  x_5008 &  n_5650;
assign n_5895 = ~n_5893 & ~n_5894;
assign n_5896 = ~n_5892 &  n_5895;
assign n_5897 = ~n_5891 &  n_5896;
assign n_5898 =  x_4305 & ~n_5897;
assign n_5899 = ~x_4305 &  n_5897;
assign n_5900 = ~n_5898 & ~n_5899;
assign n_5901 =  x_4304 &  n_5660;
assign n_5902 =  x_3295 &  n_5647;
assign n_5903 =  x_4368 &  n_5657;
assign n_5904 =  x_5007 &  n_5650;
assign n_5905 = ~n_5903 & ~n_5904;
assign n_5906 = ~n_5902 &  n_5905;
assign n_5907 = ~n_5901 &  n_5906;
assign n_5908 =  x_4304 & ~n_5907;
assign n_5909 = ~x_4304 &  n_5907;
assign n_5910 = ~n_5908 & ~n_5909;
assign n_5911 =  x_4303 &  n_5660;
assign n_5912 =  x_3294 &  n_5647;
assign n_5913 =  x_4367 &  n_5657;
assign n_5914 =  x_5006 &  n_5650;
assign n_5915 = ~n_5913 & ~n_5914;
assign n_5916 = ~n_5912 &  n_5915;
assign n_5917 = ~n_5911 &  n_5916;
assign n_5918 =  x_4303 & ~n_5917;
assign n_5919 = ~x_4303 &  n_5917;
assign n_5920 = ~n_5918 & ~n_5919;
assign n_5921 =  x_4302 &  n_5660;
assign n_5922 =  x_3293 &  n_5647;
assign n_5923 =  x_4366 &  n_5657;
assign n_5924 =  x_5005 &  n_5650;
assign n_5925 = ~n_5923 & ~n_5924;
assign n_5926 = ~n_5922 &  n_5925;
assign n_5927 = ~n_5921 &  n_5926;
assign n_5928 =  x_4302 & ~n_5927;
assign n_5929 = ~x_4302 &  n_5927;
assign n_5930 = ~n_5928 & ~n_5929;
assign n_5931 =  x_4301 &  n_5660;
assign n_5932 =  x_3292 &  n_5647;
assign n_5933 =  x_4365 &  n_5657;
assign n_5934 =  x_5004 &  n_5650;
assign n_5935 = ~n_5933 & ~n_5934;
assign n_5936 = ~n_5932 &  n_5935;
assign n_5937 = ~n_5931 &  n_5936;
assign n_5938 =  x_4301 & ~n_5937;
assign n_5939 = ~x_4301 &  n_5937;
assign n_5940 = ~n_5938 & ~n_5939;
assign n_5941 =  x_4300 &  n_5660;
assign n_5942 =  x_3291 &  n_5647;
assign n_5943 =  x_4364 &  n_5657;
assign n_5944 =  x_5003 &  n_5650;
assign n_5945 = ~n_5943 & ~n_5944;
assign n_5946 = ~n_5942 &  n_5945;
assign n_5947 = ~n_5941 &  n_5946;
assign n_5948 =  x_4300 & ~n_5947;
assign n_5949 = ~x_4300 &  n_5947;
assign n_5950 = ~n_5948 & ~n_5949;
assign n_5951 =  x_4299 &  n_5660;
assign n_5952 =  x_3290 &  n_5647;
assign n_5953 =  x_4363 &  n_5657;
assign n_5954 =  x_5002 &  n_5650;
assign n_5955 = ~n_5953 & ~n_5954;
assign n_5956 = ~n_5952 &  n_5955;
assign n_5957 = ~n_5951 &  n_5956;
assign n_5958 =  x_4299 & ~n_5957;
assign n_5959 = ~x_4299 &  n_5957;
assign n_5960 = ~n_5958 & ~n_5959;
assign n_5961 =  x_4298 &  n_5660;
assign n_5962 =  x_3289 &  n_5647;
assign n_5963 =  x_4362 &  n_5657;
assign n_5964 =  x_5001 &  n_5650;
assign n_5965 = ~n_5963 & ~n_5964;
assign n_5966 = ~n_5962 &  n_5965;
assign n_5967 = ~n_5961 &  n_5966;
assign n_5968 =  x_4298 & ~n_5967;
assign n_5969 = ~x_4298 &  n_5967;
assign n_5970 = ~n_5968 & ~n_5969;
assign n_5971 =  x_4297 &  n_5660;
assign n_5972 =  x_3288 &  n_5647;
assign n_5973 =  x_4361 &  n_5657;
assign n_5974 =  x_5000 &  n_5650;
assign n_5975 = ~n_5973 & ~n_5974;
assign n_5976 = ~n_5972 &  n_5975;
assign n_5977 = ~n_5971 &  n_5976;
assign n_5978 =  x_4297 & ~n_5977;
assign n_5979 = ~x_4297 &  n_5977;
assign n_5980 = ~n_5978 & ~n_5979;
assign n_5981 = ~x_42 &  n_350;
assign n_5982 =  n_1896 &  n_2684;
assign n_5983 =  n_5981 &  n_5982;
assign n_5984 =  x_40 &  n_2487;
assign n_5985 =  n_3341 &  n_5984;
assign n_5986 = ~n_5983 & ~n_5985;
assign n_5987 =  x_43 & ~n_5986;
assign n_5988 =  x_4296 & ~n_5987;
assign n_5989 =  i_32 &  n_5987;
assign n_5990 = ~n_5988 & ~n_5989;
assign n_5991 =  x_4296 & ~n_5990;
assign n_5992 = ~x_4296 &  n_5990;
assign n_5993 = ~n_5991 & ~n_5992;
assign n_5994 =  x_4295 & ~n_5987;
assign n_5995 =  i_31 &  n_5987;
assign n_5996 = ~n_5994 & ~n_5995;
assign n_5997 =  x_4295 & ~n_5996;
assign n_5998 = ~x_4295 &  n_5996;
assign n_5999 = ~n_5997 & ~n_5998;
assign n_6000 =  x_4294 & ~n_5987;
assign n_6001 =  i_30 &  n_5987;
assign n_6002 = ~n_6000 & ~n_6001;
assign n_6003 =  x_4294 & ~n_6002;
assign n_6004 = ~x_4294 &  n_6002;
assign n_6005 = ~n_6003 & ~n_6004;
assign n_6006 =  x_4293 & ~n_5987;
assign n_6007 =  i_29 &  n_5987;
assign n_6008 = ~n_6006 & ~n_6007;
assign n_6009 =  x_4293 & ~n_6008;
assign n_6010 = ~x_4293 &  n_6008;
assign n_6011 = ~n_6009 & ~n_6010;
assign n_6012 =  x_4292 & ~n_5987;
assign n_6013 =  i_28 &  n_5987;
assign n_6014 = ~n_6012 & ~n_6013;
assign n_6015 =  x_4292 & ~n_6014;
assign n_6016 = ~x_4292 &  n_6014;
assign n_6017 = ~n_6015 & ~n_6016;
assign n_6018 =  x_4291 & ~n_5987;
assign n_6019 =  i_27 &  n_5987;
assign n_6020 = ~n_6018 & ~n_6019;
assign n_6021 =  x_4291 & ~n_6020;
assign n_6022 = ~x_4291 &  n_6020;
assign n_6023 = ~n_6021 & ~n_6022;
assign n_6024 =  x_4290 & ~n_5987;
assign n_6025 =  i_26 &  n_5987;
assign n_6026 = ~n_6024 & ~n_6025;
assign n_6027 =  x_4290 & ~n_6026;
assign n_6028 = ~x_4290 &  n_6026;
assign n_6029 = ~n_6027 & ~n_6028;
assign n_6030 =  x_4289 & ~n_5987;
assign n_6031 =  i_25 &  n_5987;
assign n_6032 = ~n_6030 & ~n_6031;
assign n_6033 =  x_4289 & ~n_6032;
assign n_6034 = ~x_4289 &  n_6032;
assign n_6035 = ~n_6033 & ~n_6034;
assign n_6036 =  x_4288 & ~n_5987;
assign n_6037 =  i_24 &  n_5987;
assign n_6038 = ~n_6036 & ~n_6037;
assign n_6039 =  x_4288 & ~n_6038;
assign n_6040 = ~x_4288 &  n_6038;
assign n_6041 = ~n_6039 & ~n_6040;
assign n_6042 =  x_4287 & ~n_5987;
assign n_6043 =  i_23 &  n_5987;
assign n_6044 = ~n_6042 & ~n_6043;
assign n_6045 =  x_4287 & ~n_6044;
assign n_6046 = ~x_4287 &  n_6044;
assign n_6047 = ~n_6045 & ~n_6046;
assign n_6048 =  x_4286 & ~n_5987;
assign n_6049 =  i_22 &  n_5987;
assign n_6050 = ~n_6048 & ~n_6049;
assign n_6051 =  x_4286 & ~n_6050;
assign n_6052 = ~x_4286 &  n_6050;
assign n_6053 = ~n_6051 & ~n_6052;
assign n_6054 =  x_4285 & ~n_5987;
assign n_6055 =  i_21 &  n_5987;
assign n_6056 = ~n_6054 & ~n_6055;
assign n_6057 =  x_4285 & ~n_6056;
assign n_6058 = ~x_4285 &  n_6056;
assign n_6059 = ~n_6057 & ~n_6058;
assign n_6060 =  x_4284 & ~n_5987;
assign n_6061 =  i_20 &  n_5987;
assign n_6062 = ~n_6060 & ~n_6061;
assign n_6063 =  x_4284 & ~n_6062;
assign n_6064 = ~x_4284 &  n_6062;
assign n_6065 = ~n_6063 & ~n_6064;
assign n_6066 =  x_4283 & ~n_5987;
assign n_6067 =  i_19 &  n_5987;
assign n_6068 = ~n_6066 & ~n_6067;
assign n_6069 =  x_4283 & ~n_6068;
assign n_6070 = ~x_4283 &  n_6068;
assign n_6071 = ~n_6069 & ~n_6070;
assign n_6072 =  x_4282 & ~n_5987;
assign n_6073 =  i_18 &  n_5987;
assign n_6074 = ~n_6072 & ~n_6073;
assign n_6075 =  x_4282 & ~n_6074;
assign n_6076 = ~x_4282 &  n_6074;
assign n_6077 = ~n_6075 & ~n_6076;
assign n_6078 =  x_4281 & ~n_5987;
assign n_6079 =  i_17 &  n_5987;
assign n_6080 = ~n_6078 & ~n_6079;
assign n_6081 =  x_4281 & ~n_6080;
assign n_6082 = ~x_4281 &  n_6080;
assign n_6083 = ~n_6081 & ~n_6082;
assign n_6084 =  x_4280 & ~n_5987;
assign n_6085 =  i_16 &  n_5987;
assign n_6086 = ~n_6084 & ~n_6085;
assign n_6087 =  x_4280 & ~n_6086;
assign n_6088 = ~x_4280 &  n_6086;
assign n_6089 = ~n_6087 & ~n_6088;
assign n_6090 =  x_4279 & ~n_5987;
assign n_6091 =  i_15 &  n_5987;
assign n_6092 = ~n_6090 & ~n_6091;
assign n_6093 =  x_4279 & ~n_6092;
assign n_6094 = ~x_4279 &  n_6092;
assign n_6095 = ~n_6093 & ~n_6094;
assign n_6096 =  x_4278 & ~n_5987;
assign n_6097 =  i_14 &  n_5987;
assign n_6098 = ~n_6096 & ~n_6097;
assign n_6099 =  x_4278 & ~n_6098;
assign n_6100 = ~x_4278 &  n_6098;
assign n_6101 = ~n_6099 & ~n_6100;
assign n_6102 =  x_4277 & ~n_5987;
assign n_6103 =  i_13 &  n_5987;
assign n_6104 = ~n_6102 & ~n_6103;
assign n_6105 =  x_4277 & ~n_6104;
assign n_6106 = ~x_4277 &  n_6104;
assign n_6107 = ~n_6105 & ~n_6106;
assign n_6108 =  x_4276 & ~n_5987;
assign n_6109 =  i_12 &  n_5987;
assign n_6110 = ~n_6108 & ~n_6109;
assign n_6111 =  x_4276 & ~n_6110;
assign n_6112 = ~x_4276 &  n_6110;
assign n_6113 = ~n_6111 & ~n_6112;
assign n_6114 =  x_4275 & ~n_5987;
assign n_6115 =  i_11 &  n_5987;
assign n_6116 = ~n_6114 & ~n_6115;
assign n_6117 =  x_4275 & ~n_6116;
assign n_6118 = ~x_4275 &  n_6116;
assign n_6119 = ~n_6117 & ~n_6118;
assign n_6120 =  x_4274 & ~n_5987;
assign n_6121 =  i_10 &  n_5987;
assign n_6122 = ~n_6120 & ~n_6121;
assign n_6123 =  x_4274 & ~n_6122;
assign n_6124 = ~x_4274 &  n_6122;
assign n_6125 = ~n_6123 & ~n_6124;
assign n_6126 =  x_4273 & ~n_5987;
assign n_6127 =  i_9 &  n_5987;
assign n_6128 = ~n_6126 & ~n_6127;
assign n_6129 =  x_4273 & ~n_6128;
assign n_6130 = ~x_4273 &  n_6128;
assign n_6131 = ~n_6129 & ~n_6130;
assign n_6132 =  x_4272 & ~n_5987;
assign n_6133 =  i_8 &  n_5987;
assign n_6134 = ~n_6132 & ~n_6133;
assign n_6135 =  x_4272 & ~n_6134;
assign n_6136 = ~x_4272 &  n_6134;
assign n_6137 = ~n_6135 & ~n_6136;
assign n_6138 =  x_4271 & ~n_5987;
assign n_6139 =  i_7 &  n_5987;
assign n_6140 = ~n_6138 & ~n_6139;
assign n_6141 =  x_4271 & ~n_6140;
assign n_6142 = ~x_4271 &  n_6140;
assign n_6143 = ~n_6141 & ~n_6142;
assign n_6144 =  x_4270 & ~n_5987;
assign n_6145 =  i_6 &  n_5987;
assign n_6146 = ~n_6144 & ~n_6145;
assign n_6147 =  x_4270 & ~n_6146;
assign n_6148 = ~x_4270 &  n_6146;
assign n_6149 = ~n_6147 & ~n_6148;
assign n_6150 =  x_4269 & ~n_5987;
assign n_6151 =  i_5 &  n_5987;
assign n_6152 = ~n_6150 & ~n_6151;
assign n_6153 =  x_4269 & ~n_6152;
assign n_6154 = ~x_4269 &  n_6152;
assign n_6155 = ~n_6153 & ~n_6154;
assign n_6156 =  x_4268 & ~n_5987;
assign n_6157 =  i_4 &  n_5987;
assign n_6158 = ~n_6156 & ~n_6157;
assign n_6159 =  x_4268 & ~n_6158;
assign n_6160 = ~x_4268 &  n_6158;
assign n_6161 = ~n_6159 & ~n_6160;
assign n_6162 =  x_4267 & ~n_5987;
assign n_6163 =  i_3 &  n_5987;
assign n_6164 = ~n_6162 & ~n_6163;
assign n_6165 =  x_4267 & ~n_6164;
assign n_6166 = ~x_4267 &  n_6164;
assign n_6167 = ~n_6165 & ~n_6166;
assign n_6168 =  x_4266 & ~n_5987;
assign n_6169 =  i_2 &  n_5987;
assign n_6170 = ~n_6168 & ~n_6169;
assign n_6171 =  x_4266 & ~n_6170;
assign n_6172 = ~x_4266 &  n_6170;
assign n_6173 = ~n_6171 & ~n_6172;
assign n_6174 =  x_4265 & ~n_5987;
assign n_6175 =  i_1 &  n_5987;
assign n_6176 = ~n_6174 & ~n_6175;
assign n_6177 =  x_4265 & ~n_6176;
assign n_6178 = ~x_4265 &  n_6176;
assign n_6179 = ~n_6177 & ~n_6178;
assign n_6180 = ~x_42 &  n_12;
assign n_6181 =  x_39 &  n_767;
assign n_6182 =  n_5 &  n_6181;
assign n_6183 =  n_6180 &  n_6182;
assign n_6184 = ~x_43 &  n_6183;
assign n_6185 =  x_4264 & ~n_6184;
assign n_6186 =  i_32 &  n_6184;
assign n_6187 = ~n_6185 & ~n_6186;
assign n_6188 =  x_4264 & ~n_6187;
assign n_6189 = ~x_4264 &  n_6187;
assign n_6190 = ~n_6188 & ~n_6189;
assign n_6191 =  x_4263 & ~n_6184;
assign n_6192 =  i_31 &  n_6184;
assign n_6193 = ~n_6191 & ~n_6192;
assign n_6194 =  x_4263 & ~n_6193;
assign n_6195 = ~x_4263 &  n_6193;
assign n_6196 = ~n_6194 & ~n_6195;
assign n_6197 =  x_4262 & ~n_6184;
assign n_6198 =  i_30 &  n_6184;
assign n_6199 = ~n_6197 & ~n_6198;
assign n_6200 =  x_4262 & ~n_6199;
assign n_6201 = ~x_4262 &  n_6199;
assign n_6202 = ~n_6200 & ~n_6201;
assign n_6203 =  x_4261 & ~n_6184;
assign n_6204 =  i_29 &  n_6184;
assign n_6205 = ~n_6203 & ~n_6204;
assign n_6206 =  x_4261 & ~n_6205;
assign n_6207 = ~x_4261 &  n_6205;
assign n_6208 = ~n_6206 & ~n_6207;
assign n_6209 =  x_4260 & ~n_6184;
assign n_6210 =  i_28 &  n_6184;
assign n_6211 = ~n_6209 & ~n_6210;
assign n_6212 =  x_4260 & ~n_6211;
assign n_6213 = ~x_4260 &  n_6211;
assign n_6214 = ~n_6212 & ~n_6213;
assign n_6215 =  x_4259 & ~n_6184;
assign n_6216 =  i_27 &  n_6184;
assign n_6217 = ~n_6215 & ~n_6216;
assign n_6218 =  x_4259 & ~n_6217;
assign n_6219 = ~x_4259 &  n_6217;
assign n_6220 = ~n_6218 & ~n_6219;
assign n_6221 =  x_4258 & ~n_6184;
assign n_6222 =  i_26 &  n_6184;
assign n_6223 = ~n_6221 & ~n_6222;
assign n_6224 =  x_4258 & ~n_6223;
assign n_6225 = ~x_4258 &  n_6223;
assign n_6226 = ~n_6224 & ~n_6225;
assign n_6227 =  x_4257 & ~n_6184;
assign n_6228 =  i_25 &  n_6184;
assign n_6229 = ~n_6227 & ~n_6228;
assign n_6230 =  x_4257 & ~n_6229;
assign n_6231 = ~x_4257 &  n_6229;
assign n_6232 = ~n_6230 & ~n_6231;
assign n_6233 =  x_4256 & ~n_6184;
assign n_6234 =  i_24 &  n_6184;
assign n_6235 = ~n_6233 & ~n_6234;
assign n_6236 =  x_4256 & ~n_6235;
assign n_6237 = ~x_4256 &  n_6235;
assign n_6238 = ~n_6236 & ~n_6237;
assign n_6239 =  x_4255 & ~n_6184;
assign n_6240 =  i_23 &  n_6184;
assign n_6241 = ~n_6239 & ~n_6240;
assign n_6242 =  x_4255 & ~n_6241;
assign n_6243 = ~x_4255 &  n_6241;
assign n_6244 = ~n_6242 & ~n_6243;
assign n_6245 =  x_4254 & ~n_6184;
assign n_6246 =  i_22 &  n_6184;
assign n_6247 = ~n_6245 & ~n_6246;
assign n_6248 =  x_4254 & ~n_6247;
assign n_6249 = ~x_4254 &  n_6247;
assign n_6250 = ~n_6248 & ~n_6249;
assign n_6251 =  x_4253 & ~n_6184;
assign n_6252 =  i_21 &  n_6184;
assign n_6253 = ~n_6251 & ~n_6252;
assign n_6254 =  x_4253 & ~n_6253;
assign n_6255 = ~x_4253 &  n_6253;
assign n_6256 = ~n_6254 & ~n_6255;
assign n_6257 =  x_4252 & ~n_6184;
assign n_6258 =  i_20 &  n_6184;
assign n_6259 = ~n_6257 & ~n_6258;
assign n_6260 =  x_4252 & ~n_6259;
assign n_6261 = ~x_4252 &  n_6259;
assign n_6262 = ~n_6260 & ~n_6261;
assign n_6263 =  x_4251 & ~n_6184;
assign n_6264 =  i_19 &  n_6184;
assign n_6265 = ~n_6263 & ~n_6264;
assign n_6266 =  x_4251 & ~n_6265;
assign n_6267 = ~x_4251 &  n_6265;
assign n_6268 = ~n_6266 & ~n_6267;
assign n_6269 =  x_4250 & ~n_6184;
assign n_6270 =  i_18 &  n_6184;
assign n_6271 = ~n_6269 & ~n_6270;
assign n_6272 =  x_4250 & ~n_6271;
assign n_6273 = ~x_4250 &  n_6271;
assign n_6274 = ~n_6272 & ~n_6273;
assign n_6275 =  x_4249 & ~n_6184;
assign n_6276 =  i_17 &  n_6184;
assign n_6277 = ~n_6275 & ~n_6276;
assign n_6278 =  x_4249 & ~n_6277;
assign n_6279 = ~x_4249 &  n_6277;
assign n_6280 = ~n_6278 & ~n_6279;
assign n_6281 =  x_4248 & ~n_6184;
assign n_6282 =  i_16 &  n_6184;
assign n_6283 = ~n_6281 & ~n_6282;
assign n_6284 =  x_4248 & ~n_6283;
assign n_6285 = ~x_4248 &  n_6283;
assign n_6286 = ~n_6284 & ~n_6285;
assign n_6287 =  x_4247 & ~n_6184;
assign n_6288 =  i_15 &  n_6184;
assign n_6289 = ~n_6287 & ~n_6288;
assign n_6290 =  x_4247 & ~n_6289;
assign n_6291 = ~x_4247 &  n_6289;
assign n_6292 = ~n_6290 & ~n_6291;
assign n_6293 =  x_4246 & ~n_6184;
assign n_6294 =  i_14 &  n_6184;
assign n_6295 = ~n_6293 & ~n_6294;
assign n_6296 =  x_4246 & ~n_6295;
assign n_6297 = ~x_4246 &  n_6295;
assign n_6298 = ~n_6296 & ~n_6297;
assign n_6299 =  x_4245 & ~n_6184;
assign n_6300 =  i_13 &  n_6184;
assign n_6301 = ~n_6299 & ~n_6300;
assign n_6302 =  x_4245 & ~n_6301;
assign n_6303 = ~x_4245 &  n_6301;
assign n_6304 = ~n_6302 & ~n_6303;
assign n_6305 =  x_4244 & ~n_6184;
assign n_6306 =  i_12 &  n_6184;
assign n_6307 = ~n_6305 & ~n_6306;
assign n_6308 =  x_4244 & ~n_6307;
assign n_6309 = ~x_4244 &  n_6307;
assign n_6310 = ~n_6308 & ~n_6309;
assign n_6311 =  x_4243 & ~n_6184;
assign n_6312 =  i_11 &  n_6184;
assign n_6313 = ~n_6311 & ~n_6312;
assign n_6314 =  x_4243 & ~n_6313;
assign n_6315 = ~x_4243 &  n_6313;
assign n_6316 = ~n_6314 & ~n_6315;
assign n_6317 =  x_4242 & ~n_6184;
assign n_6318 =  i_10 &  n_6184;
assign n_6319 = ~n_6317 & ~n_6318;
assign n_6320 =  x_4242 & ~n_6319;
assign n_6321 = ~x_4242 &  n_6319;
assign n_6322 = ~n_6320 & ~n_6321;
assign n_6323 =  x_4241 & ~n_6184;
assign n_6324 =  i_9 &  n_6184;
assign n_6325 = ~n_6323 & ~n_6324;
assign n_6326 =  x_4241 & ~n_6325;
assign n_6327 = ~x_4241 &  n_6325;
assign n_6328 = ~n_6326 & ~n_6327;
assign n_6329 =  x_4240 & ~n_6184;
assign n_6330 =  i_8 &  n_6184;
assign n_6331 = ~n_6329 & ~n_6330;
assign n_6332 =  x_4240 & ~n_6331;
assign n_6333 = ~x_4240 &  n_6331;
assign n_6334 = ~n_6332 & ~n_6333;
assign n_6335 =  x_4239 & ~n_6184;
assign n_6336 =  i_7 &  n_6184;
assign n_6337 = ~n_6335 & ~n_6336;
assign n_6338 =  x_4239 & ~n_6337;
assign n_6339 = ~x_4239 &  n_6337;
assign n_6340 = ~n_6338 & ~n_6339;
assign n_6341 =  x_4238 & ~n_6184;
assign n_6342 =  i_6 &  n_6184;
assign n_6343 = ~n_6341 & ~n_6342;
assign n_6344 =  x_4238 & ~n_6343;
assign n_6345 = ~x_4238 &  n_6343;
assign n_6346 = ~n_6344 & ~n_6345;
assign n_6347 =  x_4237 & ~n_6184;
assign n_6348 =  i_5 &  n_6184;
assign n_6349 = ~n_6347 & ~n_6348;
assign n_6350 =  x_4237 & ~n_6349;
assign n_6351 = ~x_4237 &  n_6349;
assign n_6352 = ~n_6350 & ~n_6351;
assign n_6353 =  x_4236 & ~n_6184;
assign n_6354 =  i_4 &  n_6184;
assign n_6355 = ~n_6353 & ~n_6354;
assign n_6356 =  x_4236 & ~n_6355;
assign n_6357 = ~x_4236 &  n_6355;
assign n_6358 = ~n_6356 & ~n_6357;
assign n_6359 =  x_4235 & ~n_6184;
assign n_6360 =  i_3 &  n_6184;
assign n_6361 = ~n_6359 & ~n_6360;
assign n_6362 =  x_4235 & ~n_6361;
assign n_6363 = ~x_4235 &  n_6361;
assign n_6364 = ~n_6362 & ~n_6363;
assign n_6365 =  x_4234 & ~n_6184;
assign n_6366 =  i_2 &  n_6184;
assign n_6367 = ~n_6365 & ~n_6366;
assign n_6368 =  x_4234 & ~n_6367;
assign n_6369 = ~x_4234 &  n_6367;
assign n_6370 = ~n_6368 & ~n_6369;
assign n_6371 =  x_4233 & ~n_6184;
assign n_6372 =  i_1 &  n_6184;
assign n_6373 = ~n_6371 & ~n_6372;
assign n_6374 =  x_4233 & ~n_6373;
assign n_6375 = ~x_4233 &  n_6373;
assign n_6376 = ~n_6374 & ~n_6375;
assign n_6377 = ~x_38 &  n_3338;
assign n_6378 =  n_5654 &  n_6377;
assign n_6379 =  x_37 &  n_5;
assign n_6380 =  n_6378 &  n_6379;
assign n_6381 =  x_4232 & ~n_6380;
assign n_6382 =  i_32 &  n_6380;
assign n_6383 = ~n_6381 & ~n_6382;
assign n_6384 =  x_4232 & ~n_6383;
assign n_6385 = ~x_4232 &  n_6383;
assign n_6386 = ~n_6384 & ~n_6385;
assign n_6387 =  x_4231 & ~n_6380;
assign n_6388 =  i_31 &  n_6380;
assign n_6389 = ~n_6387 & ~n_6388;
assign n_6390 =  x_4231 & ~n_6389;
assign n_6391 = ~x_4231 &  n_6389;
assign n_6392 = ~n_6390 & ~n_6391;
assign n_6393 =  x_4230 & ~n_6380;
assign n_6394 =  i_30 &  n_6380;
assign n_6395 = ~n_6393 & ~n_6394;
assign n_6396 =  x_4230 & ~n_6395;
assign n_6397 = ~x_4230 &  n_6395;
assign n_6398 = ~n_6396 & ~n_6397;
assign n_6399 =  x_4229 & ~n_6380;
assign n_6400 =  i_29 &  n_6380;
assign n_6401 = ~n_6399 & ~n_6400;
assign n_6402 =  x_4229 & ~n_6401;
assign n_6403 = ~x_4229 &  n_6401;
assign n_6404 = ~n_6402 & ~n_6403;
assign n_6405 =  x_4228 & ~n_6380;
assign n_6406 =  i_28 &  n_6380;
assign n_6407 = ~n_6405 & ~n_6406;
assign n_6408 =  x_4228 & ~n_6407;
assign n_6409 = ~x_4228 &  n_6407;
assign n_6410 = ~n_6408 & ~n_6409;
assign n_6411 =  x_4227 & ~n_6380;
assign n_6412 =  i_27 &  n_6380;
assign n_6413 = ~n_6411 & ~n_6412;
assign n_6414 =  x_4227 & ~n_6413;
assign n_6415 = ~x_4227 &  n_6413;
assign n_6416 = ~n_6414 & ~n_6415;
assign n_6417 =  x_4226 & ~n_6380;
assign n_6418 =  i_26 &  n_6380;
assign n_6419 = ~n_6417 & ~n_6418;
assign n_6420 =  x_4226 & ~n_6419;
assign n_6421 = ~x_4226 &  n_6419;
assign n_6422 = ~n_6420 & ~n_6421;
assign n_6423 =  x_4225 & ~n_6380;
assign n_6424 =  i_25 &  n_6380;
assign n_6425 = ~n_6423 & ~n_6424;
assign n_6426 =  x_4225 & ~n_6425;
assign n_6427 = ~x_4225 &  n_6425;
assign n_6428 = ~n_6426 & ~n_6427;
assign n_6429 =  x_4224 & ~n_6380;
assign n_6430 =  i_24 &  n_6380;
assign n_6431 = ~n_6429 & ~n_6430;
assign n_6432 =  x_4224 & ~n_6431;
assign n_6433 = ~x_4224 &  n_6431;
assign n_6434 = ~n_6432 & ~n_6433;
assign n_6435 =  x_4223 & ~n_6380;
assign n_6436 =  i_23 &  n_6380;
assign n_6437 = ~n_6435 & ~n_6436;
assign n_6438 =  x_4223 & ~n_6437;
assign n_6439 = ~x_4223 &  n_6437;
assign n_6440 = ~n_6438 & ~n_6439;
assign n_6441 =  x_4222 & ~n_6380;
assign n_6442 =  i_22 &  n_6380;
assign n_6443 = ~n_6441 & ~n_6442;
assign n_6444 =  x_4222 & ~n_6443;
assign n_6445 = ~x_4222 &  n_6443;
assign n_6446 = ~n_6444 & ~n_6445;
assign n_6447 =  x_4221 & ~n_6380;
assign n_6448 =  i_21 &  n_6380;
assign n_6449 = ~n_6447 & ~n_6448;
assign n_6450 =  x_4221 & ~n_6449;
assign n_6451 = ~x_4221 &  n_6449;
assign n_6452 = ~n_6450 & ~n_6451;
assign n_6453 =  x_4220 & ~n_6380;
assign n_6454 =  i_20 &  n_6380;
assign n_6455 = ~n_6453 & ~n_6454;
assign n_6456 =  x_4220 & ~n_6455;
assign n_6457 = ~x_4220 &  n_6455;
assign n_6458 = ~n_6456 & ~n_6457;
assign n_6459 =  x_4219 & ~n_6380;
assign n_6460 =  i_19 &  n_6380;
assign n_6461 = ~n_6459 & ~n_6460;
assign n_6462 =  x_4219 & ~n_6461;
assign n_6463 = ~x_4219 &  n_6461;
assign n_6464 = ~n_6462 & ~n_6463;
assign n_6465 =  x_4218 & ~n_6380;
assign n_6466 =  i_18 &  n_6380;
assign n_6467 = ~n_6465 & ~n_6466;
assign n_6468 =  x_4218 & ~n_6467;
assign n_6469 = ~x_4218 &  n_6467;
assign n_6470 = ~n_6468 & ~n_6469;
assign n_6471 =  x_4217 & ~n_6380;
assign n_6472 =  i_17 &  n_6380;
assign n_6473 = ~n_6471 & ~n_6472;
assign n_6474 =  x_4217 & ~n_6473;
assign n_6475 = ~x_4217 &  n_6473;
assign n_6476 = ~n_6474 & ~n_6475;
assign n_6477 =  x_4216 & ~n_6380;
assign n_6478 =  i_16 &  n_6380;
assign n_6479 = ~n_6477 & ~n_6478;
assign n_6480 =  x_4216 & ~n_6479;
assign n_6481 = ~x_4216 &  n_6479;
assign n_6482 = ~n_6480 & ~n_6481;
assign n_6483 =  x_4215 & ~n_6380;
assign n_6484 =  i_15 &  n_6380;
assign n_6485 = ~n_6483 & ~n_6484;
assign n_6486 =  x_4215 & ~n_6485;
assign n_6487 = ~x_4215 &  n_6485;
assign n_6488 = ~n_6486 & ~n_6487;
assign n_6489 =  x_4214 & ~n_6380;
assign n_6490 =  i_14 &  n_6380;
assign n_6491 = ~n_6489 & ~n_6490;
assign n_6492 =  x_4214 & ~n_6491;
assign n_6493 = ~x_4214 &  n_6491;
assign n_6494 = ~n_6492 & ~n_6493;
assign n_6495 =  x_4213 & ~n_6380;
assign n_6496 =  i_13 &  n_6380;
assign n_6497 = ~n_6495 & ~n_6496;
assign n_6498 =  x_4213 & ~n_6497;
assign n_6499 = ~x_4213 &  n_6497;
assign n_6500 = ~n_6498 & ~n_6499;
assign n_6501 =  x_4212 & ~n_6380;
assign n_6502 =  i_12 &  n_6380;
assign n_6503 = ~n_6501 & ~n_6502;
assign n_6504 =  x_4212 & ~n_6503;
assign n_6505 = ~x_4212 &  n_6503;
assign n_6506 = ~n_6504 & ~n_6505;
assign n_6507 =  x_4211 & ~n_6380;
assign n_6508 =  i_11 &  n_6380;
assign n_6509 = ~n_6507 & ~n_6508;
assign n_6510 =  x_4211 & ~n_6509;
assign n_6511 = ~x_4211 &  n_6509;
assign n_6512 = ~n_6510 & ~n_6511;
assign n_6513 =  x_4210 & ~n_6380;
assign n_6514 =  i_10 &  n_6380;
assign n_6515 = ~n_6513 & ~n_6514;
assign n_6516 =  x_4210 & ~n_6515;
assign n_6517 = ~x_4210 &  n_6515;
assign n_6518 = ~n_6516 & ~n_6517;
assign n_6519 =  x_4209 & ~n_6380;
assign n_6520 =  i_9 &  n_6380;
assign n_6521 = ~n_6519 & ~n_6520;
assign n_6522 =  x_4209 & ~n_6521;
assign n_6523 = ~x_4209 &  n_6521;
assign n_6524 = ~n_6522 & ~n_6523;
assign n_6525 =  n_5654 &  n_350;
assign n_6526 =  n_3141 &  n_768;
assign n_6527 =  n_6525 &  n_6526;
assign n_6528 =  x_3505 & ~n_6527;
assign n_6529 =  i_26 &  n_6527;
assign n_6530 = ~n_6528 & ~n_6529;
assign n_6531 =  x_3505 & ~n_6530;
assign n_6532 = ~x_3505 &  n_6530;
assign n_6533 = ~n_6531 & ~n_6532;
assign n_6534 =  x_3504 & ~n_6527;
assign n_6535 =  i_25 &  n_6527;
assign n_6536 = ~n_6534 & ~n_6535;
assign n_6537 =  x_3504 & ~n_6536;
assign n_6538 = ~x_3504 &  n_6536;
assign n_6539 = ~n_6537 & ~n_6538;
assign n_6540 =  x_3503 & ~n_6527;
assign n_6541 =  i_24 &  n_6527;
assign n_6542 = ~n_6540 & ~n_6541;
assign n_6543 =  x_3503 & ~n_6542;
assign n_6544 = ~x_3503 &  n_6542;
assign n_6545 = ~n_6543 & ~n_6544;
assign n_6546 =  x_3502 & ~n_6527;
assign n_6547 =  i_23 &  n_6527;
assign n_6548 = ~n_6546 & ~n_6547;
assign n_6549 =  x_3502 & ~n_6548;
assign n_6550 = ~x_3502 &  n_6548;
assign n_6551 = ~n_6549 & ~n_6550;
assign n_6552 =  x_3501 & ~n_6527;
assign n_6553 =  i_22 &  n_6527;
assign n_6554 = ~n_6552 & ~n_6553;
assign n_6555 =  x_3501 & ~n_6554;
assign n_6556 = ~x_3501 &  n_6554;
assign n_6557 = ~n_6555 & ~n_6556;
assign n_6558 =  x_3500 & ~n_6527;
assign n_6559 =  i_21 &  n_6527;
assign n_6560 = ~n_6558 & ~n_6559;
assign n_6561 =  x_3500 & ~n_6560;
assign n_6562 = ~x_3500 &  n_6560;
assign n_6563 = ~n_6561 & ~n_6562;
assign n_6564 =  x_3499 & ~n_6527;
assign n_6565 =  i_20 &  n_6527;
assign n_6566 = ~n_6564 & ~n_6565;
assign n_6567 =  x_3499 & ~n_6566;
assign n_6568 = ~x_3499 &  n_6566;
assign n_6569 = ~n_6567 & ~n_6568;
assign n_6570 =  x_3498 & ~n_6527;
assign n_6571 =  i_19 &  n_6527;
assign n_6572 = ~n_6570 & ~n_6571;
assign n_6573 =  x_3498 & ~n_6572;
assign n_6574 = ~x_3498 &  n_6572;
assign n_6575 = ~n_6573 & ~n_6574;
assign n_6576 =  x_3497 & ~n_6527;
assign n_6577 =  i_18 &  n_6527;
assign n_6578 = ~n_6576 & ~n_6577;
assign n_6579 =  x_3497 & ~n_6578;
assign n_6580 = ~x_3497 &  n_6578;
assign n_6581 = ~n_6579 & ~n_6580;
assign n_6582 =  x_3496 & ~n_6527;
assign n_6583 =  i_17 &  n_6527;
assign n_6584 = ~n_6582 & ~n_6583;
assign n_6585 =  x_3496 & ~n_6584;
assign n_6586 = ~x_3496 &  n_6584;
assign n_6587 = ~n_6585 & ~n_6586;
assign n_6588 =  x_3495 & ~n_6527;
assign n_6589 =  i_16 &  n_6527;
assign n_6590 = ~n_6588 & ~n_6589;
assign n_6591 =  x_3495 & ~n_6590;
assign n_6592 = ~x_3495 &  n_6590;
assign n_6593 = ~n_6591 & ~n_6592;
assign n_6594 =  x_3494 & ~n_6527;
assign n_6595 =  i_15 &  n_6527;
assign n_6596 = ~n_6594 & ~n_6595;
assign n_6597 =  x_3494 & ~n_6596;
assign n_6598 = ~x_3494 &  n_6596;
assign n_6599 = ~n_6597 & ~n_6598;
assign n_6600 =  x_3493 & ~n_6527;
assign n_6601 =  i_14 &  n_6527;
assign n_6602 = ~n_6600 & ~n_6601;
assign n_6603 =  x_3493 & ~n_6602;
assign n_6604 = ~x_3493 &  n_6602;
assign n_6605 = ~n_6603 & ~n_6604;
assign n_6606 =  x_3492 & ~n_6527;
assign n_6607 =  i_13 &  n_6527;
assign n_6608 = ~n_6606 & ~n_6607;
assign n_6609 =  x_3492 & ~n_6608;
assign n_6610 = ~x_3492 &  n_6608;
assign n_6611 = ~n_6609 & ~n_6610;
assign n_6612 =  x_3491 & ~n_6527;
assign n_6613 =  i_12 &  n_6527;
assign n_6614 = ~n_6612 & ~n_6613;
assign n_6615 =  x_3491 & ~n_6614;
assign n_6616 = ~x_3491 &  n_6614;
assign n_6617 = ~n_6615 & ~n_6616;
assign n_6618 =  x_3490 & ~n_6527;
assign n_6619 =  i_11 &  n_6527;
assign n_6620 = ~n_6618 & ~n_6619;
assign n_6621 =  x_3490 & ~n_6620;
assign n_6622 = ~x_3490 &  n_6620;
assign n_6623 = ~n_6621 & ~n_6622;
assign n_6624 =  x_3489 & ~n_6527;
assign n_6625 =  i_10 &  n_6527;
assign n_6626 = ~n_6624 & ~n_6625;
assign n_6627 =  x_3489 & ~n_6626;
assign n_6628 = ~x_3489 &  n_6626;
assign n_6629 = ~n_6627 & ~n_6628;
assign n_6630 =  x_3488 & ~n_6527;
assign n_6631 =  i_9 &  n_6527;
assign n_6632 = ~n_6630 & ~n_6631;
assign n_6633 =  x_3488 & ~n_6632;
assign n_6634 = ~x_3488 &  n_6632;
assign n_6635 = ~n_6633 & ~n_6634;
assign n_6636 =  x_3487 & ~n_6527;
assign n_6637 =  i_8 &  n_6527;
assign n_6638 = ~n_6636 & ~n_6637;
assign n_6639 =  x_3487 & ~n_6638;
assign n_6640 = ~x_3487 &  n_6638;
assign n_6641 = ~n_6639 & ~n_6640;
assign n_6642 =  x_3486 & ~n_6527;
assign n_6643 =  i_7 &  n_6527;
assign n_6644 = ~n_6642 & ~n_6643;
assign n_6645 =  x_3486 & ~n_6644;
assign n_6646 = ~x_3486 &  n_6644;
assign n_6647 = ~n_6645 & ~n_6646;
assign n_6648 =  x_3485 & ~n_6527;
assign n_6649 =  i_6 &  n_6527;
assign n_6650 = ~n_6648 & ~n_6649;
assign n_6651 =  x_3485 & ~n_6650;
assign n_6652 = ~x_3485 &  n_6650;
assign n_6653 = ~n_6651 & ~n_6652;
assign n_6654 =  x_3484 & ~n_6527;
assign n_6655 =  i_5 &  n_6527;
assign n_6656 = ~n_6654 & ~n_6655;
assign n_6657 =  x_3484 & ~n_6656;
assign n_6658 = ~x_3484 &  n_6656;
assign n_6659 = ~n_6657 & ~n_6658;
assign n_6660 =  x_3483 & ~n_6527;
assign n_6661 =  i_4 &  n_6527;
assign n_6662 = ~n_6660 & ~n_6661;
assign n_6663 =  x_3483 & ~n_6662;
assign n_6664 = ~x_3483 &  n_6662;
assign n_6665 = ~n_6663 & ~n_6664;
assign n_6666 =  x_3482 & ~n_6527;
assign n_6667 =  i_3 &  n_6527;
assign n_6668 = ~n_6666 & ~n_6667;
assign n_6669 =  x_3482 & ~n_6668;
assign n_6670 = ~x_3482 &  n_6668;
assign n_6671 = ~n_6669 & ~n_6670;
assign n_6672 =  x_3481 & ~n_6527;
assign n_6673 =  i_2 &  n_6527;
assign n_6674 = ~n_6672 & ~n_6673;
assign n_6675 =  x_3481 & ~n_6674;
assign n_6676 = ~x_3481 &  n_6674;
assign n_6677 = ~n_6675 & ~n_6676;
assign n_6678 =  x_3480 & ~n_6527;
assign n_6679 =  i_1 &  n_6527;
assign n_6680 = ~n_6678 & ~n_6679;
assign n_6681 =  x_3480 & ~n_6680;
assign n_6682 = ~x_3480 &  n_6680;
assign n_6683 = ~n_6681 & ~n_6682;
assign n_6684 =  x_3479 & ~n_1901;
assign n_6685 =  x_1578 &  n_1901;
assign n_6686 = ~n_6684 & ~n_6685;
assign n_6687 =  x_3479 & ~n_6686;
assign n_6688 = ~x_3479 &  n_6686;
assign n_6689 = ~n_6687 & ~n_6688;
assign n_6690 =  x_3478 & ~n_1901;
assign n_6691 =  x_1577 &  n_1901;
assign n_6692 = ~n_6690 & ~n_6691;
assign n_6693 =  x_3478 & ~n_6692;
assign n_6694 = ~x_3478 &  n_6692;
assign n_6695 = ~n_6693 & ~n_6694;
assign n_6696 =  x_3477 & ~n_1901;
assign n_6697 =  x_1576 &  n_1901;
assign n_6698 = ~n_6696 & ~n_6697;
assign n_6699 =  x_3477 & ~n_6698;
assign n_6700 = ~x_3477 &  n_6698;
assign n_6701 = ~n_6699 & ~n_6700;
assign n_6702 =  x_3476 & ~n_1901;
assign n_6703 =  x_1575 &  n_1901;
assign n_6704 = ~n_6702 & ~n_6703;
assign n_6705 =  x_3476 & ~n_6704;
assign n_6706 = ~x_3476 &  n_6704;
assign n_6707 = ~n_6705 & ~n_6706;
assign n_6708 =  x_3475 & ~n_1901;
assign n_6709 =  x_1574 &  n_1901;
assign n_6710 = ~n_6708 & ~n_6709;
assign n_6711 =  x_3475 & ~n_6710;
assign n_6712 = ~x_3475 &  n_6710;
assign n_6713 = ~n_6711 & ~n_6712;
assign n_6714 =  x_3474 & ~n_1901;
assign n_6715 =  x_1573 &  n_1901;
assign n_6716 = ~n_6714 & ~n_6715;
assign n_6717 =  x_3474 & ~n_6716;
assign n_6718 = ~x_3474 &  n_6716;
assign n_6719 = ~n_6717 & ~n_6718;
assign n_6720 =  x_3473 & ~n_1901;
assign n_6721 =  x_1572 &  n_1901;
assign n_6722 = ~n_6720 & ~n_6721;
assign n_6723 =  x_3473 & ~n_6722;
assign n_6724 = ~x_3473 &  n_6722;
assign n_6725 = ~n_6723 & ~n_6724;
assign n_6726 =  x_3472 & ~n_1901;
assign n_6727 =  x_1571 &  n_1901;
assign n_6728 = ~n_6726 & ~n_6727;
assign n_6729 =  x_3472 & ~n_6728;
assign n_6730 = ~x_3472 &  n_6728;
assign n_6731 = ~n_6729 & ~n_6730;
assign n_6732 =  x_3471 & ~n_1901;
assign n_6733 =  x_1570 &  n_1901;
assign n_6734 = ~n_6732 & ~n_6733;
assign n_6735 =  x_3471 & ~n_6734;
assign n_6736 = ~x_3471 &  n_6734;
assign n_6737 = ~n_6735 & ~n_6736;
assign n_6738 =  x_3470 & ~n_1901;
assign n_6739 =  x_1569 &  n_1901;
assign n_6740 = ~n_6738 & ~n_6739;
assign n_6741 =  x_3470 & ~n_6740;
assign n_6742 = ~x_3470 &  n_6740;
assign n_6743 = ~n_6741 & ~n_6742;
assign n_6744 =  x_3469 & ~n_1901;
assign n_6745 =  x_1568 &  n_1901;
assign n_6746 = ~n_6744 & ~n_6745;
assign n_6747 =  x_3469 & ~n_6746;
assign n_6748 = ~x_3469 &  n_6746;
assign n_6749 = ~n_6747 & ~n_6748;
assign n_6750 =  x_3468 & ~n_1901;
assign n_6751 =  x_1567 &  n_1901;
assign n_6752 = ~n_6750 & ~n_6751;
assign n_6753 =  x_3468 & ~n_6752;
assign n_6754 = ~x_3468 &  n_6752;
assign n_6755 = ~n_6753 & ~n_6754;
assign n_6756 =  x_3467 & ~n_1901;
assign n_6757 =  x_1566 &  n_1901;
assign n_6758 = ~n_6756 & ~n_6757;
assign n_6759 =  x_3467 & ~n_6758;
assign n_6760 = ~x_3467 &  n_6758;
assign n_6761 = ~n_6759 & ~n_6760;
assign n_6762 =  x_3466 & ~n_1901;
assign n_6763 =  x_1565 &  n_1901;
assign n_6764 = ~n_6762 & ~n_6763;
assign n_6765 =  x_3466 & ~n_6764;
assign n_6766 = ~x_3466 &  n_6764;
assign n_6767 = ~n_6765 & ~n_6766;
assign n_6768 =  x_3465 & ~n_1901;
assign n_6769 =  x_1564 &  n_1901;
assign n_6770 = ~n_6768 & ~n_6769;
assign n_6771 =  x_3465 & ~n_6770;
assign n_6772 = ~x_3465 &  n_6770;
assign n_6773 = ~n_6771 & ~n_6772;
assign n_6774 =  x_3464 & ~n_1901;
assign n_6775 =  x_1563 &  n_1901;
assign n_6776 = ~n_6774 & ~n_6775;
assign n_6777 =  x_3464 & ~n_6776;
assign n_6778 = ~x_3464 &  n_6776;
assign n_6779 = ~n_6777 & ~n_6778;
assign n_6780 =  x_3463 & ~n_1901;
assign n_6781 =  x_1562 &  n_1901;
assign n_6782 = ~n_6780 & ~n_6781;
assign n_6783 =  x_3463 & ~n_6782;
assign n_6784 = ~x_3463 &  n_6782;
assign n_6785 = ~n_6783 & ~n_6784;
assign n_6786 =  x_3462 & ~n_1901;
assign n_6787 =  x_1561 &  n_1901;
assign n_6788 = ~n_6786 & ~n_6787;
assign n_6789 =  x_3462 & ~n_6788;
assign n_6790 = ~x_3462 &  n_6788;
assign n_6791 = ~n_6789 & ~n_6790;
assign n_6792 =  x_3461 & ~n_1901;
assign n_6793 =  x_1560 &  n_1901;
assign n_6794 = ~n_6792 & ~n_6793;
assign n_6795 =  x_3461 & ~n_6794;
assign n_6796 = ~x_3461 &  n_6794;
assign n_6797 = ~n_6795 & ~n_6796;
assign n_6798 =  x_3460 & ~n_1901;
assign n_6799 =  x_1559 &  n_1901;
assign n_6800 = ~n_6798 & ~n_6799;
assign n_6801 =  x_3460 & ~n_6800;
assign n_6802 = ~x_3460 &  n_6800;
assign n_6803 = ~n_6801 & ~n_6802;
assign n_6804 =  x_3459 & ~n_1901;
assign n_6805 =  x_1558 &  n_1901;
assign n_6806 = ~n_6804 & ~n_6805;
assign n_6807 =  x_3459 & ~n_6806;
assign n_6808 = ~x_3459 &  n_6806;
assign n_6809 = ~n_6807 & ~n_6808;
assign n_6810 =  x_3458 & ~n_1901;
assign n_6811 =  x_1557 &  n_1901;
assign n_6812 = ~n_6810 & ~n_6811;
assign n_6813 =  x_3458 & ~n_6812;
assign n_6814 = ~x_3458 &  n_6812;
assign n_6815 = ~n_6813 & ~n_6814;
assign n_6816 =  x_3457 & ~n_1901;
assign n_6817 =  x_1556 &  n_1901;
assign n_6818 = ~n_6816 & ~n_6817;
assign n_6819 =  x_3457 & ~n_6818;
assign n_6820 = ~x_3457 &  n_6818;
assign n_6821 = ~n_6819 & ~n_6820;
assign n_6822 =  x_3456 & ~n_1901;
assign n_6823 =  x_1555 &  n_1901;
assign n_6824 = ~n_6822 & ~n_6823;
assign n_6825 =  x_3456 & ~n_6824;
assign n_6826 = ~x_3456 &  n_6824;
assign n_6827 = ~n_6825 & ~n_6826;
assign n_6828 =  x_3455 & ~n_1901;
assign n_6829 =  x_1554 &  n_1901;
assign n_6830 = ~n_6828 & ~n_6829;
assign n_6831 =  x_3455 & ~n_6830;
assign n_6832 = ~x_3455 &  n_6830;
assign n_6833 = ~n_6831 & ~n_6832;
assign n_6834 =  x_3454 & ~n_1901;
assign n_6835 =  x_1553 &  n_1901;
assign n_6836 = ~n_6834 & ~n_6835;
assign n_6837 =  x_3454 & ~n_6836;
assign n_6838 = ~x_3454 &  n_6836;
assign n_6839 = ~n_6837 & ~n_6838;
assign n_6840 =  x_3453 & ~n_1901;
assign n_6841 =  x_1552 &  n_1901;
assign n_6842 = ~n_6840 & ~n_6841;
assign n_6843 =  x_3453 & ~n_6842;
assign n_6844 = ~x_3453 &  n_6842;
assign n_6845 = ~n_6843 & ~n_6844;
assign n_6846 =  x_3452 & ~n_1901;
assign n_6847 =  x_1551 &  n_1901;
assign n_6848 = ~n_6846 & ~n_6847;
assign n_6849 =  x_3452 & ~n_6848;
assign n_6850 = ~x_3452 &  n_6848;
assign n_6851 = ~n_6849 & ~n_6850;
assign n_6852 =  x_3451 & ~n_1901;
assign n_6853 =  x_1550 &  n_1901;
assign n_6854 = ~n_6852 & ~n_6853;
assign n_6855 =  x_3451 & ~n_6854;
assign n_6856 = ~x_3451 &  n_6854;
assign n_6857 = ~n_6855 & ~n_6856;
assign n_6858 =  x_3450 & ~n_1901;
assign n_6859 =  x_1549 &  n_1901;
assign n_6860 = ~n_6858 & ~n_6859;
assign n_6861 =  x_3450 & ~n_6860;
assign n_6862 = ~x_3450 &  n_6860;
assign n_6863 = ~n_6861 & ~n_6862;
assign n_6864 =  x_3449 & ~n_1901;
assign n_6865 =  x_1548 &  n_1901;
assign n_6866 = ~n_6864 & ~n_6865;
assign n_6867 =  x_3449 & ~n_6866;
assign n_6868 = ~x_3449 &  n_6866;
assign n_6869 = ~n_6867 & ~n_6868;
assign n_6870 =  x_3448 & ~n_1901;
assign n_6871 =  x_1547 &  n_1901;
assign n_6872 = ~n_6870 & ~n_6871;
assign n_6873 =  x_3448 & ~n_6872;
assign n_6874 = ~x_3448 &  n_6872;
assign n_6875 = ~n_6873 & ~n_6874;
assign n_6876 =  n_1305 &  n_153;
assign n_6877 = ~x_38 &  n_6876;
assign n_6878 =  n_6877 &  n_14;
assign n_6879 =  x_2314 &  n_6878;
assign n_6880 =  n_3341 &  n_5651;
assign n_6881 =  n_4289 &  n_6880;
assign n_6882 =  n_756 &  n_1305;
assign n_6883 =  n_5 &  n_6882;
assign n_6884 =  n_152 &  n_6883;
assign n_6885 = ~n_6881 & ~n_6884;
assign n_6886 =  x_43 & ~n_6885;
assign n_6887 =  x_3447 & ~n_6886;
assign n_6888 = ~n_6879 & ~n_6887;
assign n_6889 =  x_3447 & ~n_6888;
assign n_6890 = ~x_3447 &  n_6888;
assign n_6891 = ~n_6889 & ~n_6890;
assign n_6892 =  x_2313 &  n_6878;
assign n_6893 =  x_3446 & ~n_6886;
assign n_6894 = ~n_6892 & ~n_6893;
assign n_6895 =  x_3446 & ~n_6894;
assign n_6896 = ~x_3446 &  n_6894;
assign n_6897 = ~n_6895 & ~n_6896;
assign n_6898 =  x_2312 &  n_6878;
assign n_6899 =  x_3445 & ~n_6886;
assign n_6900 = ~n_6898 & ~n_6899;
assign n_6901 =  x_3445 & ~n_6900;
assign n_6902 = ~x_3445 &  n_6900;
assign n_6903 = ~n_6901 & ~n_6902;
assign n_6904 =  x_2311 &  n_6878;
assign n_6905 =  x_3444 & ~n_6886;
assign n_6906 = ~n_6904 & ~n_6905;
assign n_6907 =  x_3444 & ~n_6906;
assign n_6908 = ~x_3444 &  n_6906;
assign n_6909 = ~n_6907 & ~n_6908;
assign n_6910 =  x_2310 &  n_6878;
assign n_6911 =  x_3443 & ~n_6886;
assign n_6912 = ~n_6910 & ~n_6911;
assign n_6913 =  x_3443 & ~n_6912;
assign n_6914 = ~x_3443 &  n_6912;
assign n_6915 = ~n_6913 & ~n_6914;
assign n_6916 =  x_2309 &  n_6878;
assign n_6917 =  x_3442 & ~n_6886;
assign n_6918 = ~n_6916 & ~n_6917;
assign n_6919 =  x_3442 & ~n_6918;
assign n_6920 = ~x_3442 &  n_6918;
assign n_6921 = ~n_6919 & ~n_6920;
assign n_6922 =  x_2308 &  n_6878;
assign n_6923 =  x_3441 & ~n_6886;
assign n_6924 = ~n_6922 & ~n_6923;
assign n_6925 =  x_3441 & ~n_6924;
assign n_6926 = ~x_3441 &  n_6924;
assign n_6927 = ~n_6925 & ~n_6926;
assign n_6928 =  x_2307 &  n_6878;
assign n_6929 =  x_3440 & ~n_6886;
assign n_6930 = ~n_6928 & ~n_6929;
assign n_6931 =  x_3440 & ~n_6930;
assign n_6932 = ~x_3440 &  n_6930;
assign n_6933 = ~n_6931 & ~n_6932;
assign n_6934 =  x_2306 &  n_6878;
assign n_6935 =  x_3439 & ~n_6886;
assign n_6936 = ~n_6934 & ~n_6935;
assign n_6937 =  x_3439 & ~n_6936;
assign n_6938 = ~x_3439 &  n_6936;
assign n_6939 = ~n_6937 & ~n_6938;
assign n_6940 =  x_2305 &  n_6878;
assign n_6941 =  x_3438 & ~n_6886;
assign n_6942 = ~n_6940 & ~n_6941;
assign n_6943 =  x_3438 & ~n_6942;
assign n_6944 = ~x_3438 &  n_6942;
assign n_6945 = ~n_6943 & ~n_6944;
assign n_6946 =  x_2304 &  n_6878;
assign n_6947 =  x_3437 & ~n_6886;
assign n_6948 = ~n_6946 & ~n_6947;
assign n_6949 =  x_3437 & ~n_6948;
assign n_6950 = ~x_3437 &  n_6948;
assign n_6951 = ~n_6949 & ~n_6950;
assign n_6952 =  x_2303 &  n_6878;
assign n_6953 =  x_3436 & ~n_6886;
assign n_6954 = ~n_6952 & ~n_6953;
assign n_6955 =  x_3436 & ~n_6954;
assign n_6956 = ~x_3436 &  n_6954;
assign n_6957 = ~n_6955 & ~n_6956;
assign n_6958 =  x_2302 &  n_6878;
assign n_6959 =  x_3435 & ~n_6886;
assign n_6960 = ~n_6958 & ~n_6959;
assign n_6961 =  x_3435 & ~n_6960;
assign n_6962 = ~x_3435 &  n_6960;
assign n_6963 = ~n_6961 & ~n_6962;
assign n_6964 =  x_2301 &  n_6878;
assign n_6965 =  x_3434 & ~n_6886;
assign n_6966 = ~n_6964 & ~n_6965;
assign n_6967 =  x_3434 & ~n_6966;
assign n_6968 = ~x_3434 &  n_6966;
assign n_6969 = ~n_6967 & ~n_6968;
assign n_6970 =  x_2300 &  n_6878;
assign n_6971 =  x_3433 & ~n_6886;
assign n_6972 = ~n_6970 & ~n_6971;
assign n_6973 =  x_3433 & ~n_6972;
assign n_6974 = ~x_3433 &  n_6972;
assign n_6975 = ~n_6973 & ~n_6974;
assign n_6976 =  x_2299 &  n_6878;
assign n_6977 =  x_3432 & ~n_6886;
assign n_6978 = ~n_6976 & ~n_6977;
assign n_6979 =  x_3432 & ~n_6978;
assign n_6980 = ~x_3432 &  n_6978;
assign n_6981 = ~n_6979 & ~n_6980;
assign n_6982 =  x_2298 &  n_6878;
assign n_6983 =  x_3431 & ~n_6886;
assign n_6984 = ~n_6982 & ~n_6983;
assign n_6985 =  x_3431 & ~n_6984;
assign n_6986 = ~x_3431 &  n_6984;
assign n_6987 = ~n_6985 & ~n_6986;
assign n_6988 =  x_2297 &  n_6878;
assign n_6989 =  x_3430 & ~n_6886;
assign n_6990 = ~n_6988 & ~n_6989;
assign n_6991 =  x_3430 & ~n_6990;
assign n_6992 = ~x_3430 &  n_6990;
assign n_6993 = ~n_6991 & ~n_6992;
assign n_6994 =  x_2296 &  n_6878;
assign n_6995 =  x_3429 & ~n_6886;
assign n_6996 = ~n_6994 & ~n_6995;
assign n_6997 =  x_3429 & ~n_6996;
assign n_6998 = ~x_3429 &  n_6996;
assign n_6999 = ~n_6997 & ~n_6998;
assign n_7000 =  x_2295 &  n_6878;
assign n_7001 =  x_3428 & ~n_6886;
assign n_7002 = ~n_7000 & ~n_7001;
assign n_7003 =  x_3428 & ~n_7002;
assign n_7004 = ~x_3428 &  n_7002;
assign n_7005 = ~n_7003 & ~n_7004;
assign n_7006 =  x_2294 &  n_6878;
assign n_7007 =  x_3427 & ~n_6886;
assign n_7008 = ~n_7006 & ~n_7007;
assign n_7009 =  x_3427 & ~n_7008;
assign n_7010 = ~x_3427 &  n_7008;
assign n_7011 = ~n_7009 & ~n_7010;
assign n_7012 =  x_2293 &  n_6878;
assign n_7013 =  x_3426 & ~n_6886;
assign n_7014 = ~n_7012 & ~n_7013;
assign n_7015 =  x_3426 & ~n_7014;
assign n_7016 = ~x_3426 &  n_7014;
assign n_7017 = ~n_7015 & ~n_7016;
assign n_7018 =  x_2292 &  n_6878;
assign n_7019 =  x_3425 & ~n_6886;
assign n_7020 = ~n_7018 & ~n_7019;
assign n_7021 =  x_3425 & ~n_7020;
assign n_7022 = ~x_3425 &  n_7020;
assign n_7023 = ~n_7021 & ~n_7022;
assign n_7024 =  x_2291 &  n_6878;
assign n_7025 =  x_3424 & ~n_6886;
assign n_7026 = ~n_7024 & ~n_7025;
assign n_7027 =  x_3424 & ~n_7026;
assign n_7028 = ~x_3424 &  n_7026;
assign n_7029 = ~n_7027 & ~n_7028;
assign n_7030 =  x_2290 &  n_6878;
assign n_7031 =  x_3423 & ~n_6886;
assign n_7032 = ~n_7030 & ~n_7031;
assign n_7033 =  x_3423 & ~n_7032;
assign n_7034 = ~x_3423 &  n_7032;
assign n_7035 = ~n_7033 & ~n_7034;
assign n_7036 =  x_2289 &  n_6878;
assign n_7037 =  x_3422 & ~n_6886;
assign n_7038 = ~n_7036 & ~n_7037;
assign n_7039 =  x_3422 & ~n_7038;
assign n_7040 = ~x_3422 &  n_7038;
assign n_7041 = ~n_7039 & ~n_7040;
assign n_7042 =  x_2288 &  n_6878;
assign n_7043 =  x_3421 & ~n_6886;
assign n_7044 = ~n_7042 & ~n_7043;
assign n_7045 =  x_3421 & ~n_7044;
assign n_7046 = ~x_3421 &  n_7044;
assign n_7047 = ~n_7045 & ~n_7046;
assign n_7048 =  x_2287 &  n_6878;
assign n_7049 =  x_3420 & ~n_6886;
assign n_7050 = ~n_7048 & ~n_7049;
assign n_7051 =  x_3420 & ~n_7050;
assign n_7052 = ~x_3420 &  n_7050;
assign n_7053 = ~n_7051 & ~n_7052;
assign n_7054 =  x_2286 &  n_6878;
assign n_7055 =  x_3419 & ~n_6886;
assign n_7056 = ~n_7054 & ~n_7055;
assign n_7057 =  x_3419 & ~n_7056;
assign n_7058 = ~x_3419 &  n_7056;
assign n_7059 = ~n_7057 & ~n_7058;
assign n_7060 =  x_2285 &  n_6878;
assign n_7061 =  x_3418 & ~n_6886;
assign n_7062 = ~n_7060 & ~n_7061;
assign n_7063 =  x_3418 & ~n_7062;
assign n_7064 = ~x_3418 &  n_7062;
assign n_7065 = ~n_7063 & ~n_7064;
assign n_7066 =  x_2284 &  n_6878;
assign n_7067 =  x_3417 & ~n_6886;
assign n_7068 = ~n_7066 & ~n_7067;
assign n_7069 =  x_3417 & ~n_7068;
assign n_7070 = ~x_3417 &  n_7068;
assign n_7071 = ~n_7069 & ~n_7070;
assign n_7072 =  x_2283 &  n_6878;
assign n_7073 =  x_3416 & ~n_6886;
assign n_7074 = ~n_7072 & ~n_7073;
assign n_7075 =  x_3416 & ~n_7074;
assign n_7076 = ~x_3416 &  n_7074;
assign n_7077 = ~n_7075 & ~n_7076;
assign n_7078 =  n_759 &  n_3143;
assign n_7079 = ~x_38 &  n_14;
assign n_7080 =  n_7078 &  n_7079;
assign n_7081 =  x_3415 & ~n_7080;
assign n_7082 =  x_4743 &  n_7080;
assign n_7083 = ~n_7081 & ~n_7082;
assign n_7084 =  x_3415 & ~n_7083;
assign n_7085 = ~x_3415 &  n_7083;
assign n_7086 = ~n_7084 & ~n_7085;
assign n_7087 =  x_3414 & ~n_7080;
assign n_7088 =  x_4742 &  n_7080;
assign n_7089 = ~n_7087 & ~n_7088;
assign n_7090 =  x_3414 & ~n_7089;
assign n_7091 = ~x_3414 &  n_7089;
assign n_7092 = ~n_7090 & ~n_7091;
assign n_7093 =  x_3413 & ~n_7080;
assign n_7094 =  x_4741 &  n_7080;
assign n_7095 = ~n_7093 & ~n_7094;
assign n_7096 =  x_3413 & ~n_7095;
assign n_7097 = ~x_3413 &  n_7095;
assign n_7098 = ~n_7096 & ~n_7097;
assign n_7099 =  x_3412 & ~n_7080;
assign n_7100 =  x_4740 &  n_7080;
assign n_7101 = ~n_7099 & ~n_7100;
assign n_7102 =  x_3412 & ~n_7101;
assign n_7103 = ~x_3412 &  n_7101;
assign n_7104 = ~n_7102 & ~n_7103;
assign n_7105 =  x_3411 & ~n_7080;
assign n_7106 =  x_4739 &  n_7080;
assign n_7107 = ~n_7105 & ~n_7106;
assign n_7108 =  x_3411 & ~n_7107;
assign n_7109 = ~x_3411 &  n_7107;
assign n_7110 = ~n_7108 & ~n_7109;
assign n_7111 =  x_3410 & ~n_7080;
assign n_7112 =  x_4738 &  n_7080;
assign n_7113 = ~n_7111 & ~n_7112;
assign n_7114 =  x_3410 & ~n_7113;
assign n_7115 = ~x_3410 &  n_7113;
assign n_7116 = ~n_7114 & ~n_7115;
assign n_7117 =  x_3409 & ~n_7080;
assign n_7118 =  x_4737 &  n_7080;
assign n_7119 = ~n_7117 & ~n_7118;
assign n_7120 =  x_3409 & ~n_7119;
assign n_7121 = ~x_3409 &  n_7119;
assign n_7122 = ~n_7120 & ~n_7121;
assign n_7123 =  x_3408 & ~n_7080;
assign n_7124 =  x_4736 &  n_7080;
assign n_7125 = ~n_7123 & ~n_7124;
assign n_7126 =  x_3408 & ~n_7125;
assign n_7127 = ~x_3408 &  n_7125;
assign n_7128 = ~n_7126 & ~n_7127;
assign n_7129 =  x_3407 & ~n_7080;
assign n_7130 =  x_4735 &  n_7080;
assign n_7131 = ~n_7129 & ~n_7130;
assign n_7132 =  x_3407 & ~n_7131;
assign n_7133 = ~x_3407 &  n_7131;
assign n_7134 = ~n_7132 & ~n_7133;
assign n_7135 =  x_3406 & ~n_7080;
assign n_7136 =  x_4734 &  n_7080;
assign n_7137 = ~n_7135 & ~n_7136;
assign n_7138 =  x_3406 & ~n_7137;
assign n_7139 = ~x_3406 &  n_7137;
assign n_7140 = ~n_7138 & ~n_7139;
assign n_7141 =  x_3405 & ~n_7080;
assign n_7142 =  x_4733 &  n_7080;
assign n_7143 = ~n_7141 & ~n_7142;
assign n_7144 =  x_3405 & ~n_7143;
assign n_7145 = ~x_3405 &  n_7143;
assign n_7146 = ~n_7144 & ~n_7145;
assign n_7147 =  x_3404 & ~n_7080;
assign n_7148 =  x_4732 &  n_7080;
assign n_7149 = ~n_7147 & ~n_7148;
assign n_7150 =  x_3404 & ~n_7149;
assign n_7151 = ~x_3404 &  n_7149;
assign n_7152 = ~n_7150 & ~n_7151;
assign n_7153 =  x_3403 & ~n_7080;
assign n_7154 =  x_4731 &  n_7080;
assign n_7155 = ~n_7153 & ~n_7154;
assign n_7156 =  x_3403 & ~n_7155;
assign n_7157 = ~x_3403 &  n_7155;
assign n_7158 = ~n_7156 & ~n_7157;
assign n_7159 =  x_3402 & ~n_7080;
assign n_7160 =  x_4730 &  n_7080;
assign n_7161 = ~n_7159 & ~n_7160;
assign n_7162 =  x_3402 & ~n_7161;
assign n_7163 = ~x_3402 &  n_7161;
assign n_7164 = ~n_7162 & ~n_7163;
assign n_7165 =  x_3401 & ~n_7080;
assign n_7166 =  x_4729 &  n_7080;
assign n_7167 = ~n_7165 & ~n_7166;
assign n_7168 =  x_3401 & ~n_7167;
assign n_7169 = ~x_3401 &  n_7167;
assign n_7170 = ~n_7168 & ~n_7169;
assign n_7171 =  x_3400 & ~n_7080;
assign n_7172 =  x_4728 &  n_7080;
assign n_7173 = ~n_7171 & ~n_7172;
assign n_7174 =  x_3400 & ~n_7173;
assign n_7175 = ~x_3400 &  n_7173;
assign n_7176 = ~n_7174 & ~n_7175;
assign n_7177 =  x_3399 & ~n_7080;
assign n_7178 =  x_4727 &  n_7080;
assign n_7179 = ~n_7177 & ~n_7178;
assign n_7180 =  x_3399 & ~n_7179;
assign n_7181 = ~x_3399 &  n_7179;
assign n_7182 = ~n_7180 & ~n_7181;
assign n_7183 =  x_3398 & ~n_7080;
assign n_7184 =  x_4726 &  n_7080;
assign n_7185 = ~n_7183 & ~n_7184;
assign n_7186 =  x_3398 & ~n_7185;
assign n_7187 = ~x_3398 &  n_7185;
assign n_7188 = ~n_7186 & ~n_7187;
assign n_7189 =  x_3397 & ~n_7080;
assign n_7190 =  x_4725 &  n_7080;
assign n_7191 = ~n_7189 & ~n_7190;
assign n_7192 =  x_3397 & ~n_7191;
assign n_7193 = ~x_3397 &  n_7191;
assign n_7194 = ~n_7192 & ~n_7193;
assign n_7195 =  x_3396 & ~n_7080;
assign n_7196 =  x_4724 &  n_7080;
assign n_7197 = ~n_7195 & ~n_7196;
assign n_7198 =  x_3396 & ~n_7197;
assign n_7199 = ~x_3396 &  n_7197;
assign n_7200 = ~n_7198 & ~n_7199;
assign n_7201 =  x_3395 & ~n_7080;
assign n_7202 =  x_4723 &  n_7080;
assign n_7203 = ~n_7201 & ~n_7202;
assign n_7204 =  x_3395 & ~n_7203;
assign n_7205 = ~x_3395 &  n_7203;
assign n_7206 = ~n_7204 & ~n_7205;
assign n_7207 =  x_3394 & ~n_7080;
assign n_7208 =  x_4722 &  n_7080;
assign n_7209 = ~n_7207 & ~n_7208;
assign n_7210 =  x_3394 & ~n_7209;
assign n_7211 = ~x_3394 &  n_7209;
assign n_7212 = ~n_7210 & ~n_7211;
assign n_7213 =  x_3393 & ~n_7080;
assign n_7214 =  x_4721 &  n_7080;
assign n_7215 = ~n_7213 & ~n_7214;
assign n_7216 =  x_3393 & ~n_7215;
assign n_7217 = ~x_3393 &  n_7215;
assign n_7218 = ~n_7216 & ~n_7217;
assign n_7219 =  x_3392 & ~n_7080;
assign n_7220 =  x_4720 &  n_7080;
assign n_7221 = ~n_7219 & ~n_7220;
assign n_7222 =  x_3392 & ~n_7221;
assign n_7223 = ~x_3392 &  n_7221;
assign n_7224 = ~n_7222 & ~n_7223;
assign n_7225 =  x_3391 & ~n_7080;
assign n_7226 =  x_4719 &  n_7080;
assign n_7227 = ~n_7225 & ~n_7226;
assign n_7228 =  x_3391 & ~n_7227;
assign n_7229 = ~x_3391 &  n_7227;
assign n_7230 = ~n_7228 & ~n_7229;
assign n_7231 =  x_3390 & ~n_7080;
assign n_7232 =  x_4718 &  n_7080;
assign n_7233 = ~n_7231 & ~n_7232;
assign n_7234 =  x_3390 & ~n_7233;
assign n_7235 = ~x_3390 &  n_7233;
assign n_7236 = ~n_7234 & ~n_7235;
assign n_7237 =  x_3389 & ~n_7080;
assign n_7238 =  x_4717 &  n_7080;
assign n_7239 = ~n_7237 & ~n_7238;
assign n_7240 =  x_3389 & ~n_7239;
assign n_7241 = ~x_3389 &  n_7239;
assign n_7242 = ~n_7240 & ~n_7241;
assign n_7243 =  x_3388 & ~n_7080;
assign n_7244 =  x_4716 &  n_7080;
assign n_7245 = ~n_7243 & ~n_7244;
assign n_7246 =  x_3388 & ~n_7245;
assign n_7247 = ~x_3388 &  n_7245;
assign n_7248 = ~n_7246 & ~n_7247;
assign n_7249 =  x_3387 & ~n_7080;
assign n_7250 =  x_4715 &  n_7080;
assign n_7251 = ~n_7249 & ~n_7250;
assign n_7252 =  x_3387 & ~n_7251;
assign n_7253 = ~x_3387 &  n_7251;
assign n_7254 = ~n_7252 & ~n_7253;
assign n_7255 =  x_3386 & ~n_7080;
assign n_7256 =  x_4714 &  n_7080;
assign n_7257 = ~n_7255 & ~n_7256;
assign n_7258 =  x_3386 & ~n_7257;
assign n_7259 = ~x_3386 &  n_7257;
assign n_7260 = ~n_7258 & ~n_7259;
assign n_7261 =  x_3385 & ~n_7080;
assign n_7262 =  x_4713 &  n_7080;
assign n_7263 = ~n_7261 & ~n_7262;
assign n_7264 =  x_3385 & ~n_7263;
assign n_7265 = ~x_3385 &  n_7263;
assign n_7266 = ~n_7264 & ~n_7265;
assign n_7267 =  x_3384 & ~n_7080;
assign n_7268 =  x_4712 &  n_7080;
assign n_7269 = ~n_7267 & ~n_7268;
assign n_7270 =  x_3384 & ~n_7269;
assign n_7271 = ~x_3384 &  n_7269;
assign n_7272 = ~n_7270 & ~n_7271;
assign n_7273 =  n_551 &  n_8;
assign n_7274 =  n_1 &  n_7273;
assign n_7275 =  i_32 &  n_7274;
assign n_7276 =  x_3383 & ~n_7274;
assign n_7277 = ~n_7275 & ~n_7276;
assign n_7278 =  x_3383 & ~n_7277;
assign n_7279 = ~x_3383 &  n_7277;
assign n_7280 = ~n_7278 & ~n_7279;
assign n_7281 =  i_31 &  n_7274;
assign n_7282 =  x_3382 & ~n_7274;
assign n_7283 = ~n_7281 & ~n_7282;
assign n_7284 =  x_3382 & ~n_7283;
assign n_7285 = ~x_3382 &  n_7283;
assign n_7286 = ~n_7284 & ~n_7285;
assign n_7287 =  i_30 &  n_7274;
assign n_7288 =  x_3381 & ~n_7274;
assign n_7289 = ~n_7287 & ~n_7288;
assign n_7290 =  x_3381 & ~n_7289;
assign n_7291 = ~x_3381 &  n_7289;
assign n_7292 = ~n_7290 & ~n_7291;
assign n_7293 =  i_29 &  n_7274;
assign n_7294 =  x_3380 & ~n_7274;
assign n_7295 = ~n_7293 & ~n_7294;
assign n_7296 =  x_3380 & ~n_7295;
assign n_7297 = ~x_3380 &  n_7295;
assign n_7298 = ~n_7296 & ~n_7297;
assign n_7299 =  i_28 &  n_7274;
assign n_7300 =  x_3379 & ~n_7274;
assign n_7301 = ~n_7299 & ~n_7300;
assign n_7302 =  x_3379 & ~n_7301;
assign n_7303 = ~x_3379 &  n_7301;
assign n_7304 = ~n_7302 & ~n_7303;
assign n_7305 =  i_27 &  n_7274;
assign n_7306 =  x_3378 & ~n_7274;
assign n_7307 = ~n_7305 & ~n_7306;
assign n_7308 =  x_3378 & ~n_7307;
assign n_7309 = ~x_3378 &  n_7307;
assign n_7310 = ~n_7308 & ~n_7309;
assign n_7311 =  i_26 &  n_7274;
assign n_7312 =  x_3377 & ~n_7274;
assign n_7313 = ~n_7311 & ~n_7312;
assign n_7314 =  x_3377 & ~n_7313;
assign n_7315 = ~x_3377 &  n_7313;
assign n_7316 = ~n_7314 & ~n_7315;
assign n_7317 =  i_25 &  n_7274;
assign n_7318 =  x_3376 & ~n_7274;
assign n_7319 = ~n_7317 & ~n_7318;
assign n_7320 =  x_3376 & ~n_7319;
assign n_7321 = ~x_3376 &  n_7319;
assign n_7322 = ~n_7320 & ~n_7321;
assign n_7323 =  i_24 &  n_7274;
assign n_7324 =  x_3375 & ~n_7274;
assign n_7325 = ~n_7323 & ~n_7324;
assign n_7326 =  x_3375 & ~n_7325;
assign n_7327 = ~x_3375 &  n_7325;
assign n_7328 = ~n_7326 & ~n_7327;
assign n_7329 =  i_23 &  n_7274;
assign n_7330 =  x_3374 & ~n_7274;
assign n_7331 = ~n_7329 & ~n_7330;
assign n_7332 =  x_3374 & ~n_7331;
assign n_7333 = ~x_3374 &  n_7331;
assign n_7334 = ~n_7332 & ~n_7333;
assign n_7335 =  i_22 &  n_7274;
assign n_7336 =  x_3373 & ~n_7274;
assign n_7337 = ~n_7335 & ~n_7336;
assign n_7338 =  x_3373 & ~n_7337;
assign n_7339 = ~x_3373 &  n_7337;
assign n_7340 = ~n_7338 & ~n_7339;
assign n_7341 =  i_21 &  n_7274;
assign n_7342 =  x_3372 & ~n_7274;
assign n_7343 = ~n_7341 & ~n_7342;
assign n_7344 =  x_3372 & ~n_7343;
assign n_7345 = ~x_3372 &  n_7343;
assign n_7346 = ~n_7344 & ~n_7345;
assign n_7347 =  i_20 &  n_7274;
assign n_7348 =  x_3371 & ~n_7274;
assign n_7349 = ~n_7347 & ~n_7348;
assign n_7350 =  x_3371 & ~n_7349;
assign n_7351 = ~x_3371 &  n_7349;
assign n_7352 = ~n_7350 & ~n_7351;
assign n_7353 =  i_19 &  n_7274;
assign n_7354 =  x_3370 & ~n_7274;
assign n_7355 = ~n_7353 & ~n_7354;
assign n_7356 =  x_3370 & ~n_7355;
assign n_7357 = ~x_3370 &  n_7355;
assign n_7358 = ~n_7356 & ~n_7357;
assign n_7359 =  i_18 &  n_7274;
assign n_7360 =  x_3369 & ~n_7274;
assign n_7361 = ~n_7359 & ~n_7360;
assign n_7362 =  x_3369 & ~n_7361;
assign n_7363 = ~x_3369 &  n_7361;
assign n_7364 = ~n_7362 & ~n_7363;
assign n_7365 =  i_17 &  n_7274;
assign n_7366 =  x_3368 & ~n_7274;
assign n_7367 = ~n_7365 & ~n_7366;
assign n_7368 =  x_3368 & ~n_7367;
assign n_7369 = ~x_3368 &  n_7367;
assign n_7370 = ~n_7368 & ~n_7369;
assign n_7371 =  i_16 &  n_7274;
assign n_7372 =  x_3367 & ~n_7274;
assign n_7373 = ~n_7371 & ~n_7372;
assign n_7374 =  x_3367 & ~n_7373;
assign n_7375 = ~x_3367 &  n_7373;
assign n_7376 = ~n_7374 & ~n_7375;
assign n_7377 =  i_15 &  n_7274;
assign n_7378 =  x_3366 & ~n_7274;
assign n_7379 = ~n_7377 & ~n_7378;
assign n_7380 =  x_3366 & ~n_7379;
assign n_7381 = ~x_3366 &  n_7379;
assign n_7382 = ~n_7380 & ~n_7381;
assign n_7383 =  i_14 &  n_7274;
assign n_7384 =  x_3365 & ~n_7274;
assign n_7385 = ~n_7383 & ~n_7384;
assign n_7386 =  x_3365 & ~n_7385;
assign n_7387 = ~x_3365 &  n_7385;
assign n_7388 = ~n_7386 & ~n_7387;
assign n_7389 =  i_13 &  n_7274;
assign n_7390 =  x_3364 & ~n_7274;
assign n_7391 = ~n_7389 & ~n_7390;
assign n_7392 =  x_3364 & ~n_7391;
assign n_7393 = ~x_3364 &  n_7391;
assign n_7394 = ~n_7392 & ~n_7393;
assign n_7395 =  i_12 &  n_7274;
assign n_7396 =  x_3363 & ~n_7274;
assign n_7397 = ~n_7395 & ~n_7396;
assign n_7398 =  x_3363 & ~n_7397;
assign n_7399 = ~x_3363 &  n_7397;
assign n_7400 = ~n_7398 & ~n_7399;
assign n_7401 =  i_11 &  n_7274;
assign n_7402 =  x_3362 & ~n_7274;
assign n_7403 = ~n_7401 & ~n_7402;
assign n_7404 =  x_3362 & ~n_7403;
assign n_7405 = ~x_3362 &  n_7403;
assign n_7406 = ~n_7404 & ~n_7405;
assign n_7407 =  i_10 &  n_7274;
assign n_7408 =  x_3361 & ~n_7274;
assign n_7409 = ~n_7407 & ~n_7408;
assign n_7410 =  x_3361 & ~n_7409;
assign n_7411 = ~x_3361 &  n_7409;
assign n_7412 = ~n_7410 & ~n_7411;
assign n_7413 =  i_9 &  n_7274;
assign n_7414 =  x_3360 & ~n_7274;
assign n_7415 = ~n_7413 & ~n_7414;
assign n_7416 =  x_3360 & ~n_7415;
assign n_7417 = ~x_3360 &  n_7415;
assign n_7418 = ~n_7416 & ~n_7417;
assign n_7419 =  i_8 &  n_7274;
assign n_7420 =  x_3359 & ~n_7274;
assign n_7421 = ~n_7419 & ~n_7420;
assign n_7422 =  x_3359 & ~n_7421;
assign n_7423 = ~x_3359 &  n_7421;
assign n_7424 = ~n_7422 & ~n_7423;
assign n_7425 =  i_7 &  n_7274;
assign n_7426 =  x_3358 & ~n_7274;
assign n_7427 = ~n_7425 & ~n_7426;
assign n_7428 =  x_3358 & ~n_7427;
assign n_7429 = ~x_3358 &  n_7427;
assign n_7430 = ~n_7428 & ~n_7429;
assign n_7431 =  i_6 &  n_7274;
assign n_7432 =  x_3357 & ~n_7274;
assign n_7433 = ~n_7431 & ~n_7432;
assign n_7434 =  x_3357 & ~n_7433;
assign n_7435 = ~x_3357 &  n_7433;
assign n_7436 = ~n_7434 & ~n_7435;
assign n_7437 =  i_5 &  n_7274;
assign n_7438 =  x_3356 & ~n_7274;
assign n_7439 = ~n_7437 & ~n_7438;
assign n_7440 =  x_3356 & ~n_7439;
assign n_7441 = ~x_3356 &  n_7439;
assign n_7442 = ~n_7440 & ~n_7441;
assign n_7443 =  i_4 &  n_7274;
assign n_7444 =  x_3355 & ~n_7274;
assign n_7445 = ~n_7443 & ~n_7444;
assign n_7446 =  x_3355 & ~n_7445;
assign n_7447 = ~x_3355 &  n_7445;
assign n_7448 = ~n_7446 & ~n_7447;
assign n_7449 =  i_3 &  n_7274;
assign n_7450 =  x_3354 & ~n_7274;
assign n_7451 = ~n_7449 & ~n_7450;
assign n_7452 =  x_3354 & ~n_7451;
assign n_7453 = ~x_3354 &  n_7451;
assign n_7454 = ~n_7452 & ~n_7453;
assign n_7455 =  i_2 &  n_7274;
assign n_7456 =  x_3353 & ~n_7274;
assign n_7457 = ~n_7455 & ~n_7456;
assign n_7458 =  x_3353 & ~n_7457;
assign n_7459 = ~x_3353 &  n_7457;
assign n_7460 = ~n_7458 & ~n_7459;
assign n_7461 =  i_1 &  n_7274;
assign n_7462 =  x_3352 & ~n_7274;
assign n_7463 = ~n_7461 & ~n_7462;
assign n_7464 =  x_3352 & ~n_7463;
assign n_7465 = ~x_3352 &  n_7463;
assign n_7466 = ~n_7464 & ~n_7465;
assign n_7467 =  n_766 &  n_11;
assign n_7468 =  n_7467 &  n_6182;
assign n_7469 =  x_3351 & ~n_7468;
assign n_7470 =  i_32 &  n_7468;
assign n_7471 = ~n_7469 & ~n_7470;
assign n_7472 =  x_3351 & ~n_7471;
assign n_7473 = ~x_3351 &  n_7471;
assign n_7474 = ~n_7472 & ~n_7473;
assign n_7475 =  x_3350 & ~n_7468;
assign n_7476 =  i_31 &  n_7468;
assign n_7477 = ~n_7475 & ~n_7476;
assign n_7478 =  x_3350 & ~n_7477;
assign n_7479 = ~x_3350 &  n_7477;
assign n_7480 = ~n_7478 & ~n_7479;
assign n_7481 =  x_3349 & ~n_7468;
assign n_7482 =  i_30 &  n_7468;
assign n_7483 = ~n_7481 & ~n_7482;
assign n_7484 =  x_3349 & ~n_7483;
assign n_7485 = ~x_3349 &  n_7483;
assign n_7486 = ~n_7484 & ~n_7485;
assign n_7487 =  x_3348 & ~n_7468;
assign n_7488 =  i_29 &  n_7468;
assign n_7489 = ~n_7487 & ~n_7488;
assign n_7490 =  x_3348 & ~n_7489;
assign n_7491 = ~x_3348 &  n_7489;
assign n_7492 = ~n_7490 & ~n_7491;
assign n_7493 =  x_3347 & ~n_7468;
assign n_7494 =  i_28 &  n_7468;
assign n_7495 = ~n_7493 & ~n_7494;
assign n_7496 =  x_3347 & ~n_7495;
assign n_7497 = ~x_3347 &  n_7495;
assign n_7498 = ~n_7496 & ~n_7497;
assign n_7499 =  x_3346 & ~n_7468;
assign n_7500 =  i_27 &  n_7468;
assign n_7501 = ~n_7499 & ~n_7500;
assign n_7502 =  x_3346 & ~n_7501;
assign n_7503 = ~x_3346 &  n_7501;
assign n_7504 = ~n_7502 & ~n_7503;
assign n_7505 =  x_3345 & ~n_7468;
assign n_7506 =  i_26 &  n_7468;
assign n_7507 = ~n_7505 & ~n_7506;
assign n_7508 =  x_3345 & ~n_7507;
assign n_7509 = ~x_3345 &  n_7507;
assign n_7510 = ~n_7508 & ~n_7509;
assign n_7511 =  x_3344 & ~n_7468;
assign n_7512 =  i_25 &  n_7468;
assign n_7513 = ~n_7511 & ~n_7512;
assign n_7514 =  x_3344 & ~n_7513;
assign n_7515 = ~x_3344 &  n_7513;
assign n_7516 = ~n_7514 & ~n_7515;
assign n_7517 =  x_3343 & ~n_7468;
assign n_7518 =  i_24 &  n_7468;
assign n_7519 = ~n_7517 & ~n_7518;
assign n_7520 =  x_3343 & ~n_7519;
assign n_7521 = ~x_3343 &  n_7519;
assign n_7522 = ~n_7520 & ~n_7521;
assign n_7523 =  x_3342 & ~n_7468;
assign n_7524 =  i_23 &  n_7468;
assign n_7525 = ~n_7523 & ~n_7524;
assign n_7526 =  x_3342 & ~n_7525;
assign n_7527 = ~x_3342 &  n_7525;
assign n_7528 = ~n_7526 & ~n_7527;
assign n_7529 =  x_3341 & ~n_7468;
assign n_7530 =  i_22 &  n_7468;
assign n_7531 = ~n_7529 & ~n_7530;
assign n_7532 =  x_3341 & ~n_7531;
assign n_7533 = ~x_3341 &  n_7531;
assign n_7534 = ~n_7532 & ~n_7533;
assign n_7535 =  x_3340 & ~n_7468;
assign n_7536 =  i_21 &  n_7468;
assign n_7537 = ~n_7535 & ~n_7536;
assign n_7538 =  x_3340 & ~n_7537;
assign n_7539 = ~x_3340 &  n_7537;
assign n_7540 = ~n_7538 & ~n_7539;
assign n_7541 =  x_3339 & ~n_7468;
assign n_7542 =  i_20 &  n_7468;
assign n_7543 = ~n_7541 & ~n_7542;
assign n_7544 =  x_3339 & ~n_7543;
assign n_7545 = ~x_3339 &  n_7543;
assign n_7546 = ~n_7544 & ~n_7545;
assign n_7547 =  x_3338 & ~n_7468;
assign n_7548 =  i_19 &  n_7468;
assign n_7549 = ~n_7547 & ~n_7548;
assign n_7550 =  x_3338 & ~n_7549;
assign n_7551 = ~x_3338 &  n_7549;
assign n_7552 = ~n_7550 & ~n_7551;
assign n_7553 =  x_3337 & ~n_7468;
assign n_7554 =  i_18 &  n_7468;
assign n_7555 = ~n_7553 & ~n_7554;
assign n_7556 =  x_3337 & ~n_7555;
assign n_7557 = ~x_3337 &  n_7555;
assign n_7558 = ~n_7556 & ~n_7557;
assign n_7559 =  x_3336 & ~n_7468;
assign n_7560 =  i_17 &  n_7468;
assign n_7561 = ~n_7559 & ~n_7560;
assign n_7562 =  x_3336 & ~n_7561;
assign n_7563 = ~x_3336 &  n_7561;
assign n_7564 = ~n_7562 & ~n_7563;
assign n_7565 =  x_3335 & ~n_7468;
assign n_7566 =  i_16 &  n_7468;
assign n_7567 = ~n_7565 & ~n_7566;
assign n_7568 =  x_3335 & ~n_7567;
assign n_7569 = ~x_3335 &  n_7567;
assign n_7570 = ~n_7568 & ~n_7569;
assign n_7571 =  x_3334 & ~n_7468;
assign n_7572 =  i_15 &  n_7468;
assign n_7573 = ~n_7571 & ~n_7572;
assign n_7574 =  x_3334 & ~n_7573;
assign n_7575 = ~x_3334 &  n_7573;
assign n_7576 = ~n_7574 & ~n_7575;
assign n_7577 =  x_3333 & ~n_7468;
assign n_7578 =  i_14 &  n_7468;
assign n_7579 = ~n_7577 & ~n_7578;
assign n_7580 =  x_3333 & ~n_7579;
assign n_7581 = ~x_3333 &  n_7579;
assign n_7582 = ~n_7580 & ~n_7581;
assign n_7583 =  x_3332 & ~n_7468;
assign n_7584 =  i_13 &  n_7468;
assign n_7585 = ~n_7583 & ~n_7584;
assign n_7586 =  x_3332 & ~n_7585;
assign n_7587 = ~x_3332 &  n_7585;
assign n_7588 = ~n_7586 & ~n_7587;
assign n_7589 =  x_3331 & ~n_7468;
assign n_7590 =  i_12 &  n_7468;
assign n_7591 = ~n_7589 & ~n_7590;
assign n_7592 =  x_3331 & ~n_7591;
assign n_7593 = ~x_3331 &  n_7591;
assign n_7594 = ~n_7592 & ~n_7593;
assign n_7595 =  x_3330 & ~n_7468;
assign n_7596 =  i_11 &  n_7468;
assign n_7597 = ~n_7595 & ~n_7596;
assign n_7598 =  x_3330 & ~n_7597;
assign n_7599 = ~x_3330 &  n_7597;
assign n_7600 = ~n_7598 & ~n_7599;
assign n_7601 =  x_3329 & ~n_7468;
assign n_7602 =  i_10 &  n_7468;
assign n_7603 = ~n_7601 & ~n_7602;
assign n_7604 =  x_3329 & ~n_7603;
assign n_7605 = ~x_3329 &  n_7603;
assign n_7606 = ~n_7604 & ~n_7605;
assign n_7607 =  x_3328 & ~n_7468;
assign n_7608 =  i_9 &  n_7468;
assign n_7609 = ~n_7607 & ~n_7608;
assign n_7610 =  x_3328 & ~n_7609;
assign n_7611 = ~x_3328 &  n_7609;
assign n_7612 = ~n_7610 & ~n_7611;
assign n_7613 =  x_3327 & ~n_7468;
assign n_7614 =  i_8 &  n_7468;
assign n_7615 = ~n_7613 & ~n_7614;
assign n_7616 =  x_3327 & ~n_7615;
assign n_7617 = ~x_3327 &  n_7615;
assign n_7618 = ~n_7616 & ~n_7617;
assign n_7619 =  x_3326 & ~n_7468;
assign n_7620 =  i_7 &  n_7468;
assign n_7621 = ~n_7619 & ~n_7620;
assign n_7622 =  x_3326 & ~n_7621;
assign n_7623 = ~x_3326 &  n_7621;
assign n_7624 = ~n_7622 & ~n_7623;
assign n_7625 =  x_3325 & ~n_7468;
assign n_7626 =  i_6 &  n_7468;
assign n_7627 = ~n_7625 & ~n_7626;
assign n_7628 =  x_3325 & ~n_7627;
assign n_7629 = ~x_3325 &  n_7627;
assign n_7630 = ~n_7628 & ~n_7629;
assign n_7631 =  x_3324 & ~n_7468;
assign n_7632 =  i_5 &  n_7468;
assign n_7633 = ~n_7631 & ~n_7632;
assign n_7634 =  x_3324 & ~n_7633;
assign n_7635 = ~x_3324 &  n_7633;
assign n_7636 = ~n_7634 & ~n_7635;
assign n_7637 =  x_3323 & ~n_7468;
assign n_7638 =  i_4 &  n_7468;
assign n_7639 = ~n_7637 & ~n_7638;
assign n_7640 =  x_3323 & ~n_7639;
assign n_7641 = ~x_3323 &  n_7639;
assign n_7642 = ~n_7640 & ~n_7641;
assign n_7643 =  x_3322 & ~n_7468;
assign n_7644 =  i_3 &  n_7468;
assign n_7645 = ~n_7643 & ~n_7644;
assign n_7646 =  x_3322 & ~n_7645;
assign n_7647 = ~x_3322 &  n_7645;
assign n_7648 = ~n_7646 & ~n_7647;
assign n_7649 =  x_3321 & ~n_7468;
assign n_7650 =  i_2 &  n_7468;
assign n_7651 = ~n_7649 & ~n_7650;
assign n_7652 =  x_3321 & ~n_7651;
assign n_7653 = ~x_3321 &  n_7651;
assign n_7654 = ~n_7652 & ~n_7653;
assign n_7655 =  x_3320 & ~n_7468;
assign n_7656 =  i_1 &  n_7468;
assign n_7657 = ~n_7655 & ~n_7656;
assign n_7658 =  x_3320 & ~n_7657;
assign n_7659 = ~x_3320 &  n_7657;
assign n_7660 = ~n_7658 & ~n_7659;
assign n_7661 =  n_3341 &  n_5646;
assign n_7662 =  x_43 &  n_7661;
assign n_7663 =  x_3319 & ~n_7662;
assign n_7664 =  i_32 &  n_7662;
assign n_7665 = ~n_7663 & ~n_7664;
assign n_7666 =  x_3319 & ~n_7665;
assign n_7667 = ~x_3319 &  n_7665;
assign n_7668 = ~n_7666 & ~n_7667;
assign n_7669 =  x_3318 & ~n_7662;
assign n_7670 =  i_31 &  n_7662;
assign n_7671 = ~n_7669 & ~n_7670;
assign n_7672 =  x_3318 & ~n_7671;
assign n_7673 = ~x_3318 &  n_7671;
assign n_7674 = ~n_7672 & ~n_7673;
assign n_7675 =  x_3317 & ~n_7662;
assign n_7676 =  i_30 &  n_7662;
assign n_7677 = ~n_7675 & ~n_7676;
assign n_7678 =  x_3317 & ~n_7677;
assign n_7679 = ~x_3317 &  n_7677;
assign n_7680 = ~n_7678 & ~n_7679;
assign n_7681 =  x_3316 & ~n_7662;
assign n_7682 =  i_29 &  n_7662;
assign n_7683 = ~n_7681 & ~n_7682;
assign n_7684 =  x_3316 & ~n_7683;
assign n_7685 = ~x_3316 &  n_7683;
assign n_7686 = ~n_7684 & ~n_7685;
assign n_7687 =  x_3315 & ~n_7662;
assign n_7688 =  i_28 &  n_7662;
assign n_7689 = ~n_7687 & ~n_7688;
assign n_7690 =  x_3315 & ~n_7689;
assign n_7691 = ~x_3315 &  n_7689;
assign n_7692 = ~n_7690 & ~n_7691;
assign n_7693 =  x_3314 & ~n_7662;
assign n_7694 =  i_27 &  n_7662;
assign n_7695 = ~n_7693 & ~n_7694;
assign n_7696 =  x_3314 & ~n_7695;
assign n_7697 = ~x_3314 &  n_7695;
assign n_7698 = ~n_7696 & ~n_7697;
assign n_7699 =  x_3313 & ~n_7662;
assign n_7700 =  i_26 &  n_7662;
assign n_7701 = ~n_7699 & ~n_7700;
assign n_7702 =  x_3313 & ~n_7701;
assign n_7703 = ~x_3313 &  n_7701;
assign n_7704 = ~n_7702 & ~n_7703;
assign n_7705 =  x_3312 & ~n_7662;
assign n_7706 =  i_25 &  n_7662;
assign n_7707 = ~n_7705 & ~n_7706;
assign n_7708 =  x_3312 & ~n_7707;
assign n_7709 = ~x_3312 &  n_7707;
assign n_7710 = ~n_7708 & ~n_7709;
assign n_7711 =  x_3311 & ~n_7662;
assign n_7712 =  i_24 &  n_7662;
assign n_7713 = ~n_7711 & ~n_7712;
assign n_7714 =  x_3311 & ~n_7713;
assign n_7715 = ~x_3311 &  n_7713;
assign n_7716 = ~n_7714 & ~n_7715;
assign n_7717 =  x_3310 & ~n_7662;
assign n_7718 =  i_23 &  n_7662;
assign n_7719 = ~n_7717 & ~n_7718;
assign n_7720 =  x_3310 & ~n_7719;
assign n_7721 = ~x_3310 &  n_7719;
assign n_7722 = ~n_7720 & ~n_7721;
assign n_7723 =  x_3309 & ~n_7662;
assign n_7724 =  i_22 &  n_7662;
assign n_7725 = ~n_7723 & ~n_7724;
assign n_7726 =  x_3309 & ~n_7725;
assign n_7727 = ~x_3309 &  n_7725;
assign n_7728 = ~n_7726 & ~n_7727;
assign n_7729 =  x_3308 & ~n_7662;
assign n_7730 =  i_21 &  n_7662;
assign n_7731 = ~n_7729 & ~n_7730;
assign n_7732 =  x_3308 & ~n_7731;
assign n_7733 = ~x_3308 &  n_7731;
assign n_7734 = ~n_7732 & ~n_7733;
assign n_7735 =  x_3307 & ~n_7662;
assign n_7736 =  i_20 &  n_7662;
assign n_7737 = ~n_7735 & ~n_7736;
assign n_7738 =  x_3307 & ~n_7737;
assign n_7739 = ~x_3307 &  n_7737;
assign n_7740 = ~n_7738 & ~n_7739;
assign n_7741 =  x_3306 & ~n_7662;
assign n_7742 =  i_19 &  n_7662;
assign n_7743 = ~n_7741 & ~n_7742;
assign n_7744 =  x_3306 & ~n_7743;
assign n_7745 = ~x_3306 &  n_7743;
assign n_7746 = ~n_7744 & ~n_7745;
assign n_7747 =  x_3305 & ~n_7662;
assign n_7748 =  i_18 &  n_7662;
assign n_7749 = ~n_7747 & ~n_7748;
assign n_7750 =  x_3305 & ~n_7749;
assign n_7751 = ~x_3305 &  n_7749;
assign n_7752 = ~n_7750 & ~n_7751;
assign n_7753 =  x_3304 & ~n_7662;
assign n_7754 =  i_17 &  n_7662;
assign n_7755 = ~n_7753 & ~n_7754;
assign n_7756 =  x_3304 & ~n_7755;
assign n_7757 = ~x_3304 &  n_7755;
assign n_7758 = ~n_7756 & ~n_7757;
assign n_7759 =  x_3303 & ~n_7662;
assign n_7760 =  i_16 &  n_7662;
assign n_7761 = ~n_7759 & ~n_7760;
assign n_7762 =  x_3303 & ~n_7761;
assign n_7763 = ~x_3303 &  n_7761;
assign n_7764 = ~n_7762 & ~n_7763;
assign n_7765 =  x_3302 & ~n_7662;
assign n_7766 =  i_15 &  n_7662;
assign n_7767 = ~n_7765 & ~n_7766;
assign n_7768 =  x_3302 & ~n_7767;
assign n_7769 = ~x_3302 &  n_7767;
assign n_7770 = ~n_7768 & ~n_7769;
assign n_7771 =  x_3301 & ~n_7662;
assign n_7772 =  i_14 &  n_7662;
assign n_7773 = ~n_7771 & ~n_7772;
assign n_7774 =  x_3301 & ~n_7773;
assign n_7775 = ~x_3301 &  n_7773;
assign n_7776 = ~n_7774 & ~n_7775;
assign n_7777 =  x_3300 & ~n_7662;
assign n_7778 =  i_13 &  n_7662;
assign n_7779 = ~n_7777 & ~n_7778;
assign n_7780 =  x_3300 & ~n_7779;
assign n_7781 = ~x_3300 &  n_7779;
assign n_7782 = ~n_7780 & ~n_7781;
assign n_7783 =  x_3299 & ~n_7662;
assign n_7784 =  i_12 &  n_7662;
assign n_7785 = ~n_7783 & ~n_7784;
assign n_7786 =  x_3299 & ~n_7785;
assign n_7787 = ~x_3299 &  n_7785;
assign n_7788 = ~n_7786 & ~n_7787;
assign n_7789 =  x_3298 & ~n_7662;
assign n_7790 =  i_11 &  n_7662;
assign n_7791 = ~n_7789 & ~n_7790;
assign n_7792 =  x_3298 & ~n_7791;
assign n_7793 = ~x_3298 &  n_7791;
assign n_7794 = ~n_7792 & ~n_7793;
assign n_7795 =  x_3297 & ~n_7662;
assign n_7796 =  i_10 &  n_7662;
assign n_7797 = ~n_7795 & ~n_7796;
assign n_7798 =  x_3297 & ~n_7797;
assign n_7799 = ~x_3297 &  n_7797;
assign n_7800 = ~n_7798 & ~n_7799;
assign n_7801 =  x_3296 & ~n_7662;
assign n_7802 =  i_9 &  n_7662;
assign n_7803 = ~n_7801 & ~n_7802;
assign n_7804 =  x_3296 & ~n_7803;
assign n_7805 = ~x_3296 &  n_7803;
assign n_7806 = ~n_7804 & ~n_7805;
assign n_7807 =  x_3295 & ~n_7662;
assign n_7808 =  i_8 &  n_7662;
assign n_7809 = ~n_7807 & ~n_7808;
assign n_7810 =  x_3295 & ~n_7809;
assign n_7811 = ~x_3295 &  n_7809;
assign n_7812 = ~n_7810 & ~n_7811;
assign n_7813 =  x_3294 & ~n_7662;
assign n_7814 =  i_7 &  n_7662;
assign n_7815 = ~n_7813 & ~n_7814;
assign n_7816 =  x_3294 & ~n_7815;
assign n_7817 = ~x_3294 &  n_7815;
assign n_7818 = ~n_7816 & ~n_7817;
assign n_7819 =  x_3293 & ~n_7662;
assign n_7820 =  i_6 &  n_7662;
assign n_7821 = ~n_7819 & ~n_7820;
assign n_7822 =  x_3293 & ~n_7821;
assign n_7823 = ~x_3293 &  n_7821;
assign n_7824 = ~n_7822 & ~n_7823;
assign n_7825 =  x_3292 & ~n_7662;
assign n_7826 =  i_5 &  n_7662;
assign n_7827 = ~n_7825 & ~n_7826;
assign n_7828 =  x_3292 & ~n_7827;
assign n_7829 = ~x_3292 &  n_7827;
assign n_7830 = ~n_7828 & ~n_7829;
assign n_7831 =  x_3291 & ~n_7662;
assign n_7832 =  i_4 &  n_7662;
assign n_7833 = ~n_7831 & ~n_7832;
assign n_7834 =  x_3291 & ~n_7833;
assign n_7835 = ~x_3291 &  n_7833;
assign n_7836 = ~n_7834 & ~n_7835;
assign n_7837 =  x_3290 & ~n_7662;
assign n_7838 =  i_3 &  n_7662;
assign n_7839 = ~n_7837 & ~n_7838;
assign n_7840 =  x_3290 & ~n_7839;
assign n_7841 = ~x_3290 &  n_7839;
assign n_7842 = ~n_7840 & ~n_7841;
assign n_7843 =  x_3289 & ~n_7662;
assign n_7844 =  i_2 &  n_7662;
assign n_7845 = ~n_7843 & ~n_7844;
assign n_7846 =  x_3289 & ~n_7845;
assign n_7847 = ~x_3289 &  n_7845;
assign n_7848 = ~n_7846 & ~n_7847;
assign n_7849 =  x_3288 & ~n_7662;
assign n_7850 =  i_1 &  n_7662;
assign n_7851 = ~n_7849 & ~n_7850;
assign n_7852 =  x_3288 & ~n_7851;
assign n_7853 = ~x_3288 &  n_7851;
assign n_7854 = ~n_7852 & ~n_7853;
assign n_7855 =  n_11 &  n_5655;
assign n_7856 =  n_4290 &  n_7855;
assign n_7857 =  x_3287 & ~n_7856;
assign n_7858 =  i_32 &  n_7856;
assign n_7859 = ~n_7857 & ~n_7858;
assign n_7860 =  x_3287 & ~n_7859;
assign n_7861 = ~x_3287 &  n_7859;
assign n_7862 = ~n_7860 & ~n_7861;
assign n_7863 =  x_3286 & ~n_7856;
assign n_7864 =  i_31 &  n_7856;
assign n_7865 = ~n_7863 & ~n_7864;
assign n_7866 =  x_3286 & ~n_7865;
assign n_7867 = ~x_3286 &  n_7865;
assign n_7868 = ~n_7866 & ~n_7867;
assign n_7869 =  x_3285 & ~n_7856;
assign n_7870 =  i_30 &  n_7856;
assign n_7871 = ~n_7869 & ~n_7870;
assign n_7872 =  x_3285 & ~n_7871;
assign n_7873 = ~x_3285 &  n_7871;
assign n_7874 = ~n_7872 & ~n_7873;
assign n_7875 =  x_3284 & ~n_7856;
assign n_7876 =  i_29 &  n_7856;
assign n_7877 = ~n_7875 & ~n_7876;
assign n_7878 =  x_3284 & ~n_7877;
assign n_7879 = ~x_3284 &  n_7877;
assign n_7880 = ~n_7878 & ~n_7879;
assign n_7881 =  x_3283 & ~n_7856;
assign n_7882 =  i_28 &  n_7856;
assign n_7883 = ~n_7881 & ~n_7882;
assign n_7884 =  x_3283 & ~n_7883;
assign n_7885 = ~x_3283 &  n_7883;
assign n_7886 = ~n_7884 & ~n_7885;
assign n_7887 =  x_3282 & ~n_7856;
assign n_7888 =  i_27 &  n_7856;
assign n_7889 = ~n_7887 & ~n_7888;
assign n_7890 =  x_3282 & ~n_7889;
assign n_7891 = ~x_3282 &  n_7889;
assign n_7892 = ~n_7890 & ~n_7891;
assign n_7893 =  x_3281 & ~n_7856;
assign n_7894 =  i_26 &  n_7856;
assign n_7895 = ~n_7893 & ~n_7894;
assign n_7896 =  x_3281 & ~n_7895;
assign n_7897 = ~x_3281 &  n_7895;
assign n_7898 = ~n_7896 & ~n_7897;
assign n_7899 =  x_3280 & ~n_7856;
assign n_7900 =  i_25 &  n_7856;
assign n_7901 = ~n_7899 & ~n_7900;
assign n_7902 =  x_3280 & ~n_7901;
assign n_7903 = ~x_3280 &  n_7901;
assign n_7904 = ~n_7902 & ~n_7903;
assign n_7905 =  x_3279 & ~n_7856;
assign n_7906 =  i_24 &  n_7856;
assign n_7907 = ~n_7905 & ~n_7906;
assign n_7908 =  x_3279 & ~n_7907;
assign n_7909 = ~x_3279 &  n_7907;
assign n_7910 = ~n_7908 & ~n_7909;
assign n_7911 =  x_3278 & ~n_7856;
assign n_7912 =  i_23 &  n_7856;
assign n_7913 = ~n_7911 & ~n_7912;
assign n_7914 =  x_3278 & ~n_7913;
assign n_7915 = ~x_3278 &  n_7913;
assign n_7916 = ~n_7914 & ~n_7915;
assign n_7917 =  x_3277 & ~n_7856;
assign n_7918 =  i_22 &  n_7856;
assign n_7919 = ~n_7917 & ~n_7918;
assign n_7920 =  x_3277 & ~n_7919;
assign n_7921 = ~x_3277 &  n_7919;
assign n_7922 = ~n_7920 & ~n_7921;
assign n_7923 =  x_3276 & ~n_7856;
assign n_7924 =  i_21 &  n_7856;
assign n_7925 = ~n_7923 & ~n_7924;
assign n_7926 =  x_3276 & ~n_7925;
assign n_7927 = ~x_3276 &  n_7925;
assign n_7928 = ~n_7926 & ~n_7927;
assign n_7929 =  x_3275 & ~n_7856;
assign n_7930 =  i_20 &  n_7856;
assign n_7931 = ~n_7929 & ~n_7930;
assign n_7932 =  x_3275 & ~n_7931;
assign n_7933 = ~x_3275 &  n_7931;
assign n_7934 = ~n_7932 & ~n_7933;
assign n_7935 =  x_3274 & ~n_7856;
assign n_7936 =  i_19 &  n_7856;
assign n_7937 = ~n_7935 & ~n_7936;
assign n_7938 =  x_3274 & ~n_7937;
assign n_7939 = ~x_3274 &  n_7937;
assign n_7940 = ~n_7938 & ~n_7939;
assign n_7941 =  x_3273 & ~n_7856;
assign n_7942 =  i_18 &  n_7856;
assign n_7943 = ~n_7941 & ~n_7942;
assign n_7944 =  x_3273 & ~n_7943;
assign n_7945 = ~x_3273 &  n_7943;
assign n_7946 = ~n_7944 & ~n_7945;
assign n_7947 =  x_3272 & ~n_7856;
assign n_7948 =  i_17 &  n_7856;
assign n_7949 = ~n_7947 & ~n_7948;
assign n_7950 =  x_3272 & ~n_7949;
assign n_7951 = ~x_3272 &  n_7949;
assign n_7952 = ~n_7950 & ~n_7951;
assign n_7953 =  x_3271 & ~n_7856;
assign n_7954 =  i_16 &  n_7856;
assign n_7955 = ~n_7953 & ~n_7954;
assign n_7956 =  x_3271 & ~n_7955;
assign n_7957 = ~x_3271 &  n_7955;
assign n_7958 = ~n_7956 & ~n_7957;
assign n_7959 =  x_3270 & ~n_7856;
assign n_7960 =  i_15 &  n_7856;
assign n_7961 = ~n_7959 & ~n_7960;
assign n_7962 =  x_3270 & ~n_7961;
assign n_7963 = ~x_3270 &  n_7961;
assign n_7964 = ~n_7962 & ~n_7963;
assign n_7965 =  x_3269 & ~n_7856;
assign n_7966 =  i_14 &  n_7856;
assign n_7967 = ~n_7965 & ~n_7966;
assign n_7968 =  x_3269 & ~n_7967;
assign n_7969 = ~x_3269 &  n_7967;
assign n_7970 = ~n_7968 & ~n_7969;
assign n_7971 =  x_3268 & ~n_7856;
assign n_7972 =  i_13 &  n_7856;
assign n_7973 = ~n_7971 & ~n_7972;
assign n_7974 =  x_3268 & ~n_7973;
assign n_7975 = ~x_3268 &  n_7973;
assign n_7976 = ~n_7974 & ~n_7975;
assign n_7977 =  x_3267 & ~n_7856;
assign n_7978 =  i_12 &  n_7856;
assign n_7979 = ~n_7977 & ~n_7978;
assign n_7980 =  x_3267 & ~n_7979;
assign n_7981 = ~x_3267 &  n_7979;
assign n_7982 = ~n_7980 & ~n_7981;
assign n_7983 =  x_3266 & ~n_7856;
assign n_7984 =  i_11 &  n_7856;
assign n_7985 = ~n_7983 & ~n_7984;
assign n_7986 =  x_3266 & ~n_7985;
assign n_7987 = ~x_3266 &  n_7985;
assign n_7988 = ~n_7986 & ~n_7987;
assign n_7989 =  x_3265 & ~n_7856;
assign n_7990 =  i_10 &  n_7856;
assign n_7991 = ~n_7989 & ~n_7990;
assign n_7992 =  x_3265 & ~n_7991;
assign n_7993 = ~x_3265 &  n_7991;
assign n_7994 = ~n_7992 & ~n_7993;
assign n_7995 =  x_3264 & ~n_7856;
assign n_7996 =  i_9 &  n_7856;
assign n_7997 = ~n_7995 & ~n_7996;
assign n_7998 =  x_3264 & ~n_7997;
assign n_7999 = ~x_3264 &  n_7997;
assign n_8000 = ~n_7998 & ~n_7999;
assign n_8001 =  x_3263 & ~n_7856;
assign n_8002 =  i_8 &  n_7856;
assign n_8003 = ~n_8001 & ~n_8002;
assign n_8004 =  x_3263 & ~n_8003;
assign n_8005 = ~x_3263 &  n_8003;
assign n_8006 = ~n_8004 & ~n_8005;
assign n_8007 =  x_3262 & ~n_7856;
assign n_8008 =  i_7 &  n_7856;
assign n_8009 = ~n_8007 & ~n_8008;
assign n_8010 =  x_3262 & ~n_8009;
assign n_8011 = ~x_3262 &  n_8009;
assign n_8012 = ~n_8010 & ~n_8011;
assign n_8013 =  x_3261 & ~n_7856;
assign n_8014 =  i_6 &  n_7856;
assign n_8015 = ~n_8013 & ~n_8014;
assign n_8016 =  x_3261 & ~n_8015;
assign n_8017 = ~x_3261 &  n_8015;
assign n_8018 = ~n_8016 & ~n_8017;
assign n_8019 =  x_3260 & ~n_7856;
assign n_8020 =  i_5 &  n_7856;
assign n_8021 = ~n_8019 & ~n_8020;
assign n_8022 =  x_3260 & ~n_8021;
assign n_8023 = ~x_3260 &  n_8021;
assign n_8024 = ~n_8022 & ~n_8023;
assign n_8025 =  x_3259 & ~n_7856;
assign n_8026 =  i_4 &  n_7856;
assign n_8027 = ~n_8025 & ~n_8026;
assign n_8028 =  x_3259 & ~n_8027;
assign n_8029 = ~x_3259 &  n_8027;
assign n_8030 = ~n_8028 & ~n_8029;
assign n_8031 =  x_3258 & ~n_7856;
assign n_8032 =  i_3 &  n_7856;
assign n_8033 = ~n_8031 & ~n_8032;
assign n_8034 =  x_3258 & ~n_8033;
assign n_8035 = ~x_3258 &  n_8033;
assign n_8036 = ~n_8034 & ~n_8035;
assign n_8037 =  x_3257 & ~n_7856;
assign n_8038 =  i_2 &  n_7856;
assign n_8039 = ~n_8037 & ~n_8038;
assign n_8040 =  x_3257 & ~n_8039;
assign n_8041 = ~x_3257 &  n_8039;
assign n_8042 = ~n_8040 & ~n_8041;
assign n_8043 =  x_3256 & ~n_7856;
assign n_8044 =  i_1 &  n_7856;
assign n_8045 = ~n_8043 & ~n_8044;
assign n_8046 =  x_3256 & ~n_8045;
assign n_8047 = ~x_3256 &  n_8045;
assign n_8048 = ~n_8046 & ~n_8047;
assign n_8049 =  x_40 &  n_560;
assign n_8050 = ~n_762 & ~n_8049;
assign n_8051 =  n_758 & ~n_8050;
assign n_8052 =  x_3255 & ~n_8051;
assign n_8053 =  x_38 &  n_552;
assign n_8054 =  n_349 &  n_4285;
assign n_8055 =  n_8053 &  n_8054;
assign n_8056 = ~x_3255 &  n_8055;
assign n_8057 = ~n_761 & ~n_8056;
assign n_8058 = ~n_8052 &  n_8057;
assign n_8059 =  x_3255 & ~n_8058;
assign n_8060 = ~x_3255 &  n_8058;
assign n_8061 = ~n_8059 & ~n_8060;
assign n_8062 =  n_8051 & ~n_8056;
assign n_8063 =  x_3254 & ~n_8062;
assign n_8064 = ~x_3254 &  x_3255;
assign n_8065 =  n_8055 &  n_8064;
assign n_8066 = ~n_8063 & ~n_8065;
assign n_8067 =  x_3254 & ~n_8066;
assign n_8068 = ~x_3254 &  n_8066;
assign n_8069 = ~n_8067 & ~n_8068;
assign n_8070 =  x_3253 & ~n_8051;
assign n_8071 =  x_3254 &  x_3255;
assign n_8072 =  x_3253 &  n_8071;
assign n_8073 = ~x_3253 & ~n_8071;
assign n_8074 = ~n_8072 & ~n_8073;
assign n_8075 =  n_8055 &  n_8074;
assign n_8076 = ~n_8070 & ~n_8075;
assign n_8077 =  x_3253 & ~n_8076;
assign n_8078 = ~x_3253 &  n_8076;
assign n_8079 = ~n_8077 & ~n_8078;
assign n_8080 =  x_3252 & ~n_8051;
assign n_8081 =  x_3252 &  n_8072;
assign n_8082 = ~x_3252 & ~n_8072;
assign n_8083 = ~n_8081 & ~n_8082;
assign n_8084 =  n_8055 &  n_8083;
assign n_8085 = ~n_8080 & ~n_8084;
assign n_8086 =  x_3252 & ~n_8085;
assign n_8087 = ~x_3252 &  n_8085;
assign n_8088 = ~n_8086 & ~n_8087;
assign n_8089 =  n_8055 &  n_8081;
assign n_8090 = ~x_3251 & ~n_8089;
assign n_8091 =  x_3251 &  n_8081;
assign n_8092 =  n_8055 & ~n_8091;
assign n_8093 =  n_8051 & ~n_8092;
assign n_8094 = ~n_8090 & ~n_8093;
assign n_8095 = ~n_761 & ~n_8094;
assign n_8096 =  x_3251 & ~n_8095;
assign n_8097 = ~x_3251 &  n_8095;
assign n_8098 = ~n_8096 & ~n_8097;
assign n_8099 =  n_8055 &  n_8091;
assign n_8100 = ~x_3250 & ~n_8099;
assign n_8101 =  x_3250 & ~n_8092;
assign n_8102 =  n_8051 &  n_8101;
assign n_8103 = ~n_8100 & ~n_8102;
assign n_8104 = ~n_761 & ~n_8103;
assign n_8105 =  x_3250 & ~n_8104;
assign n_8106 = ~x_3250 &  n_8104;
assign n_8107 = ~n_8105 & ~n_8106;
assign n_8108 =  x_3250 &  n_8091;
assign n_8109 = ~x_3249 & ~n_8108;
assign n_8110 =  x_3249 &  n_8108;
assign n_8111 =  n_8055 & ~n_8110;
assign n_8112 = ~n_8109 &  n_8111;
assign n_8113 =  x_3249 & ~n_8051;
assign n_8114 = ~n_761 & ~n_8113;
assign n_8115 = ~n_8112 &  n_8114;
assign n_8116 =  x_3249 & ~n_8115;
assign n_8117 = ~x_3249 &  n_8115;
assign n_8118 = ~n_8116 & ~n_8117;
assign n_8119 =  x_3248 & ~n_8051;
assign n_8120 = ~x_3248 & ~n_8110;
assign n_8121 =  x_3248 &  n_8110;
assign n_8122 =  n_8055 & ~n_8121;
assign n_8123 = ~n_8120 &  n_8122;
assign n_8124 = ~n_8119 & ~n_8123;
assign n_8125 =  x_3248 & ~n_8124;
assign n_8126 = ~x_3248 &  n_8124;
assign n_8127 = ~n_8125 & ~n_8126;
assign n_8128 = ~x_3247 & ~n_8121;
assign n_8129 =  x_3247 &  n_8121;
assign n_8130 =  n_8055 & ~n_8129;
assign n_8131 = ~n_8128 &  n_8130;
assign n_8132 =  x_3247 & ~n_8051;
assign n_8133 = ~n_761 & ~n_8132;
assign n_8134 = ~n_8131 &  n_8133;
assign n_8135 =  x_3247 & ~n_8134;
assign n_8136 = ~x_3247 &  n_8134;
assign n_8137 = ~n_8135 & ~n_8136;
assign n_8138 =  x_3246 & ~n_8051;
assign n_8139 = ~x_3246 & ~n_8129;
assign n_8140 =  x_3246 &  n_8129;
assign n_8141 =  n_8055 & ~n_8140;
assign n_8142 = ~n_8139 &  n_8141;
assign n_8143 = ~n_8138 & ~n_8142;
assign n_8144 =  x_3246 & ~n_8143;
assign n_8145 = ~x_3246 &  n_8143;
assign n_8146 = ~n_8144 & ~n_8145;
assign n_8147 = ~x_3245 & ~n_8140;
assign n_8148 =  x_3245 &  n_8140;
assign n_8149 =  n_8055 & ~n_8148;
assign n_8150 = ~n_8147 &  n_8149;
assign n_8151 =  x_3245 & ~n_8051;
assign n_8152 = ~n_761 & ~n_8151;
assign n_8153 = ~n_8150 &  n_8152;
assign n_8154 =  x_3245 & ~n_8153;
assign n_8155 = ~x_3245 &  n_8153;
assign n_8156 = ~n_8154 & ~n_8155;
assign n_8157 =  x_3244 & ~n_8051;
assign n_8158 = ~x_3244 & ~n_8148;
assign n_8159 =  x_3244 &  n_8148;
assign n_8160 =  n_8055 & ~n_8159;
assign n_8161 = ~n_8158 &  n_8160;
assign n_8162 = ~n_8157 & ~n_8161;
assign n_8163 =  x_3244 & ~n_8162;
assign n_8164 = ~x_3244 &  n_8162;
assign n_8165 = ~n_8163 & ~n_8164;
assign n_8166 =  x_3243 & ~n_8051;
assign n_8167 = ~x_3243 & ~n_8159;
assign n_8168 =  x_3243 &  n_8159;
assign n_8169 =  n_8055 & ~n_8168;
assign n_8170 = ~n_8167 &  n_8169;
assign n_8171 = ~n_8166 & ~n_8170;
assign n_8172 =  x_3243 & ~n_8171;
assign n_8173 = ~x_3243 &  n_8171;
assign n_8174 = ~n_8172 & ~n_8173;
assign n_8175 =  x_3242 & ~n_8051;
assign n_8176 = ~x_3242 & ~n_8168;
assign n_8177 =  x_3242 &  n_8168;
assign n_8178 =  n_8055 & ~n_8177;
assign n_8179 = ~n_8176 &  n_8178;
assign n_8180 = ~n_8175 & ~n_8179;
assign n_8181 =  x_3242 & ~n_8180;
assign n_8182 = ~x_3242 &  n_8180;
assign n_8183 = ~n_8181 & ~n_8182;
assign n_8184 =  x_3241 & ~n_8051;
assign n_8185 = ~x_3241 & ~n_8177;
assign n_8186 =  x_3241 &  n_8177;
assign n_8187 =  n_8055 & ~n_8186;
assign n_8188 = ~n_8185 &  n_8187;
assign n_8189 = ~n_8184 & ~n_8188;
assign n_8190 =  x_3241 & ~n_8189;
assign n_8191 = ~x_3241 &  n_8189;
assign n_8192 = ~n_8190 & ~n_8191;
assign n_8193 =  x_3240 & ~n_8051;
assign n_8194 = ~x_3240 & ~n_8186;
assign n_8195 =  x_3240 &  n_8186;
assign n_8196 =  n_8055 & ~n_8195;
assign n_8197 = ~n_8194 &  n_8196;
assign n_8198 = ~n_8193 & ~n_8197;
assign n_8199 =  x_3240 & ~n_8198;
assign n_8200 = ~x_3240 &  n_8198;
assign n_8201 = ~n_8199 & ~n_8200;
assign n_8202 =  x_3239 & ~n_8051;
assign n_8203 = ~x_3239 & ~n_8195;
assign n_8204 =  x_3239 &  n_8195;
assign n_8205 =  n_8055 & ~n_8204;
assign n_8206 = ~n_8203 &  n_8205;
assign n_8207 = ~n_8202 & ~n_8206;
assign n_8208 =  x_3239 & ~n_8207;
assign n_8209 = ~x_3239 &  n_8207;
assign n_8210 = ~n_8208 & ~n_8209;
assign n_8211 =  x_3238 & ~n_8051;
assign n_8212 = ~x_3238 & ~n_8204;
assign n_8213 =  x_3238 &  n_8204;
assign n_8214 =  n_8055 & ~n_8213;
assign n_8215 = ~n_8212 &  n_8214;
assign n_8216 = ~n_8211 & ~n_8215;
assign n_8217 =  x_3238 & ~n_8216;
assign n_8218 = ~x_3238 &  n_8216;
assign n_8219 = ~n_8217 & ~n_8218;
assign n_8220 =  x_3237 & ~n_8051;
assign n_8221 = ~x_3237 & ~n_8213;
assign n_8222 =  x_3237 &  n_8213;
assign n_8223 =  n_8055 & ~n_8222;
assign n_8224 = ~n_8221 &  n_8223;
assign n_8225 = ~n_8220 & ~n_8224;
assign n_8226 =  x_3237 & ~n_8225;
assign n_8227 = ~x_3237 &  n_8225;
assign n_8228 = ~n_8226 & ~n_8227;
assign n_8229 =  x_3236 & ~n_8051;
assign n_8230 = ~x_3236 & ~n_8222;
assign n_8231 =  x_3236 &  n_8222;
assign n_8232 =  n_8055 & ~n_8231;
assign n_8233 = ~n_8230 &  n_8232;
assign n_8234 = ~n_8229 & ~n_8233;
assign n_8235 =  x_3236 & ~n_8234;
assign n_8236 = ~x_3236 &  n_8234;
assign n_8237 = ~n_8235 & ~n_8236;
assign n_8238 =  x_3235 & ~n_8051;
assign n_8239 = ~x_3235 & ~n_8231;
assign n_8240 =  x_3235 &  n_8231;
assign n_8241 =  n_8055 & ~n_8240;
assign n_8242 = ~n_8239 &  n_8241;
assign n_8243 = ~n_8238 & ~n_8242;
assign n_8244 =  x_3235 & ~n_8243;
assign n_8245 = ~x_3235 &  n_8243;
assign n_8246 = ~n_8244 & ~n_8245;
assign n_8247 =  x_3234 & ~n_8051;
assign n_8248 = ~x_3234 & ~n_8240;
assign n_8249 =  x_3234 &  n_8240;
assign n_8250 =  n_8055 & ~n_8249;
assign n_8251 = ~n_8248 &  n_8250;
assign n_8252 = ~n_8247 & ~n_8251;
assign n_8253 =  x_3234 & ~n_8252;
assign n_8254 = ~x_3234 &  n_8252;
assign n_8255 = ~n_8253 & ~n_8254;
assign n_8256 =  x_3233 & ~n_8051;
assign n_8257 = ~x_3233 & ~n_8249;
assign n_8258 =  x_3233 &  n_8249;
assign n_8259 =  n_8055 & ~n_8258;
assign n_8260 = ~n_8257 &  n_8259;
assign n_8261 = ~n_8256 & ~n_8260;
assign n_8262 =  x_3233 & ~n_8261;
assign n_8263 = ~x_3233 &  n_8261;
assign n_8264 = ~n_8262 & ~n_8263;
assign n_8265 =  x_3232 & ~n_8051;
assign n_8266 = ~x_3232 & ~n_8258;
assign n_8267 =  x_3232 &  n_8258;
assign n_8268 =  n_8055 & ~n_8267;
assign n_8269 = ~n_8266 &  n_8268;
assign n_8270 = ~n_8265 & ~n_8269;
assign n_8271 =  x_3232 & ~n_8270;
assign n_8272 = ~x_3232 &  n_8270;
assign n_8273 = ~n_8271 & ~n_8272;
assign n_8274 =  x_3231 & ~n_8051;
assign n_8275 = ~x_3231 & ~n_8267;
assign n_8276 =  x_3231 &  n_8267;
assign n_8277 =  n_8055 & ~n_8276;
assign n_8278 = ~n_8275 &  n_8277;
assign n_8279 = ~n_8274 & ~n_8278;
assign n_8280 =  x_3231 & ~n_8279;
assign n_8281 = ~x_3231 &  n_8279;
assign n_8282 = ~n_8280 & ~n_8281;
assign n_8283 =  x_3230 & ~n_8051;
assign n_8284 = ~x_3230 & ~n_8276;
assign n_8285 =  x_3230 &  n_8276;
assign n_8286 =  n_8055 & ~n_8285;
assign n_8287 = ~n_8284 &  n_8286;
assign n_8288 = ~n_8283 & ~n_8287;
assign n_8289 =  x_3230 & ~n_8288;
assign n_8290 = ~x_3230 &  n_8288;
assign n_8291 = ~n_8289 & ~n_8290;
assign n_8292 =  x_3229 & ~n_8051;
assign n_8293 = ~x_3229 & ~n_8285;
assign n_8294 =  x_3229 &  n_8285;
assign n_8295 =  n_8055 & ~n_8294;
assign n_8296 = ~n_8293 &  n_8295;
assign n_8297 = ~n_8292 & ~n_8296;
assign n_8298 =  x_3229 & ~n_8297;
assign n_8299 = ~x_3229 &  n_8297;
assign n_8300 = ~n_8298 & ~n_8299;
assign n_8301 =  x_3228 & ~n_8051;
assign n_8302 = ~x_3228 & ~n_8294;
assign n_8303 =  x_3228 &  n_8294;
assign n_8304 =  n_8055 & ~n_8303;
assign n_8305 = ~n_8302 &  n_8304;
assign n_8306 = ~n_8301 & ~n_8305;
assign n_8307 =  x_3228 & ~n_8306;
assign n_8308 = ~x_3228 &  n_8306;
assign n_8309 = ~n_8307 & ~n_8308;
assign n_8310 =  x_3227 & ~n_8051;
assign n_8311 = ~x_3227 & ~n_8303;
assign n_8312 =  x_3227 &  n_8303;
assign n_8313 =  n_8055 & ~n_8312;
assign n_8314 = ~n_8311 &  n_8313;
assign n_8315 = ~n_8310 & ~n_8314;
assign n_8316 =  x_3227 & ~n_8315;
assign n_8317 = ~x_3227 &  n_8315;
assign n_8318 = ~n_8316 & ~n_8317;
assign n_8319 =  x_3226 & ~n_8051;
assign n_8320 = ~x_3226 & ~n_8312;
assign n_8321 =  x_3226 &  n_8312;
assign n_8322 =  n_8055 & ~n_8321;
assign n_8323 = ~n_8320 &  n_8322;
assign n_8324 = ~n_8319 & ~n_8323;
assign n_8325 =  x_3226 & ~n_8324;
assign n_8326 = ~x_3226 &  n_8324;
assign n_8327 = ~n_8325 & ~n_8326;
assign n_8328 =  x_3225 &  n_8321;
assign n_8329 =  n_8055 & ~n_8328;
assign n_8330 =  n_8051 & ~n_8329;
assign n_8331 =  x_3225 & ~n_8330;
assign n_8332 =  n_8321 &  n_8329;
assign n_8333 = ~n_8331 & ~n_8332;
assign n_8334 =  x_3225 & ~n_8333;
assign n_8335 = ~x_3225 &  n_8333;
assign n_8336 = ~n_8334 & ~n_8335;
assign n_8337 =  x_3224 & ~n_8330;
assign n_8338 = ~x_3224 &  n_8055;
assign n_8339 =  n_8328 &  n_8338;
assign n_8340 = ~n_8337 & ~n_8339;
assign n_8341 =  x_3224 & ~n_8340;
assign n_8342 = ~x_3224 &  n_8340;
assign n_8343 = ~n_8341 & ~n_8342;
assign n_8344 =  n_1037 &  n_12;
assign n_8345 =  n_1041 &  n_8344;
assign n_8346 =  n_1040 &  n_8345;
assign n_8347 =  x_41 &  n_1040;
assign n_8348 =  n_2880 &  n_8347;
assign n_8349 =  n_11 &  n_8348;
assign n_8350 = ~n_8346 & ~n_8349;
assign n_8351 =  n_555 &  n_2291;
assign n_8352 = ~x_41 &  n_1305;
assign n_8353 =  n_1037 &  n_8352;
assign n_8354 =  x_38 &  n_2486;
assign n_8355 =  n_8353 &  n_8354;
assign n_8356 = ~n_8351 & ~n_8355;
assign n_8357 =  n_8350 &  n_8356;
assign n_8358 =  n_1175 &  n_2685;
assign n_8359 =  x_37 &  n_1040;
assign n_8360 =  n_151 &  n_8359;
assign n_8361 =  n_349 &  n_12;
assign n_8362 =  n_8360 &  n_8361;
assign n_8363 = ~n_8358 & ~n_8362;
assign n_8364 =  n_8360 &  n_8344;
assign n_8365 =  n_5654 &  n_12;
assign n_8366 =  n_8360 &  n_8365;
assign n_8367 = ~n_8364 & ~n_8366;
assign n_8368 =  n_8363 &  n_8367;
assign n_8369 =  n_8357 &  n_8368;
assign n_8370 =  x_3192 &  n_8369;
assign n_8371 =  i_32 & ~n_8368;
assign n_8372 =  x_2154 &  n_8346;
assign n_8373 =  x_1194 &  n_8355;
assign n_8374 = ~n_8372 & ~n_8373;
assign n_8375 =  x_2282 &  n_8349;
assign n_8376 =  x_1226 &  n_8351;
assign n_8377 = ~n_8375 & ~n_8376;
assign n_8378 =  n_8374 &  n_8377;
assign n_8379 = ~n_8371 &  n_8378;
assign n_8380 = ~n_8370 &  n_8379;
assign n_8381 =  x_3192 & ~n_8380;
assign n_8382 = ~x_3192 &  n_8380;
assign n_8383 = ~n_8381 & ~n_8382;
assign n_8384 =  x_3191 &  n_8369;
assign n_8385 =  i_31 & ~n_8368;
assign n_8386 =  x_2153 &  n_8346;
assign n_8387 =  x_1193 &  n_8355;
assign n_8388 = ~n_8386 & ~n_8387;
assign n_8389 =  x_2281 &  n_8349;
assign n_8390 =  x_1225 &  n_8351;
assign n_8391 = ~n_8389 & ~n_8390;
assign n_8392 =  n_8388 &  n_8391;
assign n_8393 = ~n_8385 &  n_8392;
assign n_8394 = ~n_8384 &  n_8393;
assign n_8395 =  x_3191 & ~n_8394;
assign n_8396 = ~x_3191 &  n_8394;
assign n_8397 = ~n_8395 & ~n_8396;
assign n_8398 =  x_3190 &  n_8369;
assign n_8399 =  i_30 & ~n_8368;
assign n_8400 =  x_2152 &  n_8346;
assign n_8401 =  x_1192 &  n_8355;
assign n_8402 = ~n_8400 & ~n_8401;
assign n_8403 =  x_2280 &  n_8349;
assign n_8404 =  x_1224 &  n_8351;
assign n_8405 = ~n_8403 & ~n_8404;
assign n_8406 =  n_8402 &  n_8405;
assign n_8407 = ~n_8399 &  n_8406;
assign n_8408 = ~n_8398 &  n_8407;
assign n_8409 =  x_3190 & ~n_8408;
assign n_8410 = ~x_3190 &  n_8408;
assign n_8411 = ~n_8409 & ~n_8410;
assign n_8412 =  x_3189 &  n_8369;
assign n_8413 =  i_29 & ~n_8368;
assign n_8414 =  x_2151 &  n_8346;
assign n_8415 =  x_1191 &  n_8355;
assign n_8416 = ~n_8414 & ~n_8415;
assign n_8417 =  x_2279 &  n_8349;
assign n_8418 =  x_1223 &  n_8351;
assign n_8419 = ~n_8417 & ~n_8418;
assign n_8420 =  n_8416 &  n_8419;
assign n_8421 = ~n_8413 &  n_8420;
assign n_8422 = ~n_8412 &  n_8421;
assign n_8423 =  x_3189 & ~n_8422;
assign n_8424 = ~x_3189 &  n_8422;
assign n_8425 = ~n_8423 & ~n_8424;
assign n_8426 =  x_3188 &  n_8369;
assign n_8427 =  i_28 & ~n_8368;
assign n_8428 =  x_2150 &  n_8346;
assign n_8429 =  x_1190 &  n_8355;
assign n_8430 = ~n_8428 & ~n_8429;
assign n_8431 =  x_2278 &  n_8349;
assign n_8432 =  x_1222 &  n_8351;
assign n_8433 = ~n_8431 & ~n_8432;
assign n_8434 =  n_8430 &  n_8433;
assign n_8435 = ~n_8427 &  n_8434;
assign n_8436 = ~n_8426 &  n_8435;
assign n_8437 =  x_3188 & ~n_8436;
assign n_8438 = ~x_3188 &  n_8436;
assign n_8439 = ~n_8437 & ~n_8438;
assign n_8440 =  x_3187 &  n_8369;
assign n_8441 =  i_27 & ~n_8368;
assign n_8442 =  x_2149 &  n_8346;
assign n_8443 =  x_1189 &  n_8355;
assign n_8444 = ~n_8442 & ~n_8443;
assign n_8445 =  x_2277 &  n_8349;
assign n_8446 =  x_1221 &  n_8351;
assign n_8447 = ~n_8445 & ~n_8446;
assign n_8448 =  n_8444 &  n_8447;
assign n_8449 = ~n_8441 &  n_8448;
assign n_8450 = ~n_8440 &  n_8449;
assign n_8451 =  x_3187 & ~n_8450;
assign n_8452 = ~x_3187 &  n_8450;
assign n_8453 = ~n_8451 & ~n_8452;
assign n_8454 =  x_3186 &  n_8369;
assign n_8455 =  i_26 & ~n_8368;
assign n_8456 =  x_2148 &  n_8346;
assign n_8457 =  x_1188 &  n_8355;
assign n_8458 = ~n_8456 & ~n_8457;
assign n_8459 =  x_2276 &  n_8349;
assign n_8460 =  x_1220 &  n_8351;
assign n_8461 = ~n_8459 & ~n_8460;
assign n_8462 =  n_8458 &  n_8461;
assign n_8463 = ~n_8455 &  n_8462;
assign n_8464 = ~n_8454 &  n_8463;
assign n_8465 =  x_3186 & ~n_8464;
assign n_8466 = ~x_3186 &  n_8464;
assign n_8467 = ~n_8465 & ~n_8466;
assign n_8468 =  x_3185 &  n_8369;
assign n_8469 =  i_25 & ~n_8368;
assign n_8470 =  x_2147 &  n_8346;
assign n_8471 =  x_1187 &  n_8355;
assign n_8472 = ~n_8470 & ~n_8471;
assign n_8473 =  x_2275 &  n_8349;
assign n_8474 =  x_1219 &  n_8351;
assign n_8475 = ~n_8473 & ~n_8474;
assign n_8476 =  n_8472 &  n_8475;
assign n_8477 = ~n_8469 &  n_8476;
assign n_8478 = ~n_8468 &  n_8477;
assign n_8479 =  x_3185 & ~n_8478;
assign n_8480 = ~x_3185 &  n_8478;
assign n_8481 = ~n_8479 & ~n_8480;
assign n_8482 =  x_3184 &  n_8369;
assign n_8483 =  i_24 & ~n_8368;
assign n_8484 =  x_2146 &  n_8346;
assign n_8485 =  x_1186 &  n_8355;
assign n_8486 = ~n_8484 & ~n_8485;
assign n_8487 =  x_2274 &  n_8349;
assign n_8488 =  x_1218 &  n_8351;
assign n_8489 = ~n_8487 & ~n_8488;
assign n_8490 =  n_8486 &  n_8489;
assign n_8491 = ~n_8483 &  n_8490;
assign n_8492 = ~n_8482 &  n_8491;
assign n_8493 =  x_3184 & ~n_8492;
assign n_8494 = ~x_3184 &  n_8492;
assign n_8495 = ~n_8493 & ~n_8494;
assign n_8496 =  x_3183 &  n_8369;
assign n_8497 =  i_23 & ~n_8368;
assign n_8498 =  x_2145 &  n_8346;
assign n_8499 =  x_1185 &  n_8355;
assign n_8500 = ~n_8498 & ~n_8499;
assign n_8501 =  x_2273 &  n_8349;
assign n_8502 =  x_1217 &  n_8351;
assign n_8503 = ~n_8501 & ~n_8502;
assign n_8504 =  n_8500 &  n_8503;
assign n_8505 = ~n_8497 &  n_8504;
assign n_8506 = ~n_8496 &  n_8505;
assign n_8507 =  x_3183 & ~n_8506;
assign n_8508 = ~x_3183 &  n_8506;
assign n_8509 = ~n_8507 & ~n_8508;
assign n_8510 =  x_3182 &  n_8369;
assign n_8511 =  i_22 & ~n_8368;
assign n_8512 =  x_2144 &  n_8346;
assign n_8513 =  x_1184 &  n_8355;
assign n_8514 = ~n_8512 & ~n_8513;
assign n_8515 =  x_2272 &  n_8349;
assign n_8516 =  x_1216 &  n_8351;
assign n_8517 = ~n_8515 & ~n_8516;
assign n_8518 =  n_8514 &  n_8517;
assign n_8519 = ~n_8511 &  n_8518;
assign n_8520 = ~n_8510 &  n_8519;
assign n_8521 =  x_3182 & ~n_8520;
assign n_8522 = ~x_3182 &  n_8520;
assign n_8523 = ~n_8521 & ~n_8522;
assign n_8524 =  x_3181 &  n_8369;
assign n_8525 =  i_21 & ~n_8368;
assign n_8526 =  x_2143 &  n_8346;
assign n_8527 =  x_1183 &  n_8355;
assign n_8528 = ~n_8526 & ~n_8527;
assign n_8529 =  x_2271 &  n_8349;
assign n_8530 =  x_1215 &  n_8351;
assign n_8531 = ~n_8529 & ~n_8530;
assign n_8532 =  n_8528 &  n_8531;
assign n_8533 = ~n_8525 &  n_8532;
assign n_8534 = ~n_8524 &  n_8533;
assign n_8535 =  x_3181 & ~n_8534;
assign n_8536 = ~x_3181 &  n_8534;
assign n_8537 = ~n_8535 & ~n_8536;
assign n_8538 =  x_3180 &  n_8369;
assign n_8539 =  i_20 & ~n_8368;
assign n_8540 =  x_2142 &  n_8346;
assign n_8541 =  x_1182 &  n_8355;
assign n_8542 = ~n_8540 & ~n_8541;
assign n_8543 =  x_2270 &  n_8349;
assign n_8544 =  x_1214 &  n_8351;
assign n_8545 = ~n_8543 & ~n_8544;
assign n_8546 =  n_8542 &  n_8545;
assign n_8547 = ~n_8539 &  n_8546;
assign n_8548 = ~n_8538 &  n_8547;
assign n_8549 =  x_3180 & ~n_8548;
assign n_8550 = ~x_3180 &  n_8548;
assign n_8551 = ~n_8549 & ~n_8550;
assign n_8552 =  x_3179 &  n_8369;
assign n_8553 =  i_19 & ~n_8368;
assign n_8554 =  x_2141 &  n_8346;
assign n_8555 =  x_1181 &  n_8355;
assign n_8556 = ~n_8554 & ~n_8555;
assign n_8557 =  x_2269 &  n_8349;
assign n_8558 =  x_1213 &  n_8351;
assign n_8559 = ~n_8557 & ~n_8558;
assign n_8560 =  n_8556 &  n_8559;
assign n_8561 = ~n_8553 &  n_8560;
assign n_8562 = ~n_8552 &  n_8561;
assign n_8563 =  x_3179 & ~n_8562;
assign n_8564 = ~x_3179 &  n_8562;
assign n_8565 = ~n_8563 & ~n_8564;
assign n_8566 =  x_3178 &  n_8369;
assign n_8567 =  i_18 & ~n_8368;
assign n_8568 =  x_2140 &  n_8346;
assign n_8569 =  x_1180 &  n_8355;
assign n_8570 = ~n_8568 & ~n_8569;
assign n_8571 =  x_2268 &  n_8349;
assign n_8572 =  x_1212 &  n_8351;
assign n_8573 = ~n_8571 & ~n_8572;
assign n_8574 =  n_8570 &  n_8573;
assign n_8575 = ~n_8567 &  n_8574;
assign n_8576 = ~n_8566 &  n_8575;
assign n_8577 =  x_3178 & ~n_8576;
assign n_8578 = ~x_3178 &  n_8576;
assign n_8579 = ~n_8577 & ~n_8578;
assign n_8580 =  x_3177 &  n_8369;
assign n_8581 =  i_17 & ~n_8368;
assign n_8582 =  x_2139 &  n_8346;
assign n_8583 =  x_1179 &  n_8355;
assign n_8584 = ~n_8582 & ~n_8583;
assign n_8585 =  x_2267 &  n_8349;
assign n_8586 =  x_1211 &  n_8351;
assign n_8587 = ~n_8585 & ~n_8586;
assign n_8588 =  n_8584 &  n_8587;
assign n_8589 = ~n_8581 &  n_8588;
assign n_8590 = ~n_8580 &  n_8589;
assign n_8591 =  x_3177 & ~n_8590;
assign n_8592 = ~x_3177 &  n_8590;
assign n_8593 = ~n_8591 & ~n_8592;
assign n_8594 =  x_3176 &  n_8369;
assign n_8595 =  i_16 & ~n_8368;
assign n_8596 =  x_2138 &  n_8346;
assign n_8597 =  x_1178 &  n_8355;
assign n_8598 = ~n_8596 & ~n_8597;
assign n_8599 =  x_2266 &  n_8349;
assign n_8600 =  x_1210 &  n_8351;
assign n_8601 = ~n_8599 & ~n_8600;
assign n_8602 =  n_8598 &  n_8601;
assign n_8603 = ~n_8595 &  n_8602;
assign n_8604 = ~n_8594 &  n_8603;
assign n_8605 =  x_3176 & ~n_8604;
assign n_8606 = ~x_3176 &  n_8604;
assign n_8607 = ~n_8605 & ~n_8606;
assign n_8608 =  x_3175 &  n_8369;
assign n_8609 =  i_15 & ~n_8368;
assign n_8610 =  x_2137 &  n_8346;
assign n_8611 =  x_1177 &  n_8355;
assign n_8612 = ~n_8610 & ~n_8611;
assign n_8613 =  x_2265 &  n_8349;
assign n_8614 =  x_1209 &  n_8351;
assign n_8615 = ~n_8613 & ~n_8614;
assign n_8616 =  n_8612 &  n_8615;
assign n_8617 = ~n_8609 &  n_8616;
assign n_8618 = ~n_8608 &  n_8617;
assign n_8619 =  x_3175 & ~n_8618;
assign n_8620 = ~x_3175 &  n_8618;
assign n_8621 = ~n_8619 & ~n_8620;
assign n_8622 =  x_3174 &  n_8369;
assign n_8623 =  i_14 & ~n_8368;
assign n_8624 =  x_2136 &  n_8346;
assign n_8625 =  x_1176 &  n_8355;
assign n_8626 = ~n_8624 & ~n_8625;
assign n_8627 =  x_2264 &  n_8349;
assign n_8628 =  x_1208 &  n_8351;
assign n_8629 = ~n_8627 & ~n_8628;
assign n_8630 =  n_8626 &  n_8629;
assign n_8631 = ~n_8623 &  n_8630;
assign n_8632 = ~n_8622 &  n_8631;
assign n_8633 =  x_3174 & ~n_8632;
assign n_8634 = ~x_3174 &  n_8632;
assign n_8635 = ~n_8633 & ~n_8634;
assign n_8636 =  x_3173 &  n_8369;
assign n_8637 =  i_13 & ~n_8368;
assign n_8638 =  x_2135 &  n_8346;
assign n_8639 =  x_1175 &  n_8355;
assign n_8640 = ~n_8638 & ~n_8639;
assign n_8641 =  x_2263 &  n_8349;
assign n_8642 =  x_1207 &  n_8351;
assign n_8643 = ~n_8641 & ~n_8642;
assign n_8644 =  n_8640 &  n_8643;
assign n_8645 = ~n_8637 &  n_8644;
assign n_8646 = ~n_8636 &  n_8645;
assign n_8647 =  x_3173 & ~n_8646;
assign n_8648 = ~x_3173 &  n_8646;
assign n_8649 = ~n_8647 & ~n_8648;
assign n_8650 =  x_3172 &  n_8369;
assign n_8651 =  i_12 & ~n_8368;
assign n_8652 =  x_2134 &  n_8346;
assign n_8653 =  x_1174 &  n_8355;
assign n_8654 = ~n_8652 & ~n_8653;
assign n_8655 =  x_2262 &  n_8349;
assign n_8656 =  x_1206 &  n_8351;
assign n_8657 = ~n_8655 & ~n_8656;
assign n_8658 =  n_8654 &  n_8657;
assign n_8659 = ~n_8651 &  n_8658;
assign n_8660 = ~n_8650 &  n_8659;
assign n_8661 =  x_3172 & ~n_8660;
assign n_8662 = ~x_3172 &  n_8660;
assign n_8663 = ~n_8661 & ~n_8662;
assign n_8664 =  x_3171 &  n_8369;
assign n_8665 =  i_11 & ~n_8368;
assign n_8666 =  x_2133 &  n_8346;
assign n_8667 =  x_1173 &  n_8355;
assign n_8668 = ~n_8666 & ~n_8667;
assign n_8669 =  x_2261 &  n_8349;
assign n_8670 =  x_1205 &  n_8351;
assign n_8671 = ~n_8669 & ~n_8670;
assign n_8672 =  n_8668 &  n_8671;
assign n_8673 = ~n_8665 &  n_8672;
assign n_8674 = ~n_8664 &  n_8673;
assign n_8675 =  x_3171 & ~n_8674;
assign n_8676 = ~x_3171 &  n_8674;
assign n_8677 = ~n_8675 & ~n_8676;
assign n_8678 =  x_3170 &  n_8369;
assign n_8679 =  i_10 & ~n_8368;
assign n_8680 =  x_2132 &  n_8346;
assign n_8681 =  x_1172 &  n_8355;
assign n_8682 = ~n_8680 & ~n_8681;
assign n_8683 =  x_2260 &  n_8349;
assign n_8684 =  x_1204 &  n_8351;
assign n_8685 = ~n_8683 & ~n_8684;
assign n_8686 =  n_8682 &  n_8685;
assign n_8687 = ~n_8679 &  n_8686;
assign n_8688 = ~n_8678 &  n_8687;
assign n_8689 =  x_3170 & ~n_8688;
assign n_8690 = ~x_3170 &  n_8688;
assign n_8691 = ~n_8689 & ~n_8690;
assign n_8692 =  x_3169 &  n_8369;
assign n_8693 =  i_9 & ~n_8368;
assign n_8694 =  x_2131 &  n_8346;
assign n_8695 =  x_1171 &  n_8355;
assign n_8696 = ~n_8694 & ~n_8695;
assign n_8697 =  x_2259 &  n_8349;
assign n_8698 =  x_1203 &  n_8351;
assign n_8699 = ~n_8697 & ~n_8698;
assign n_8700 =  n_8696 &  n_8699;
assign n_8701 = ~n_8693 &  n_8700;
assign n_8702 = ~n_8692 &  n_8701;
assign n_8703 =  x_3169 & ~n_8702;
assign n_8704 = ~x_3169 &  n_8702;
assign n_8705 = ~n_8703 & ~n_8704;
assign n_8706 =  x_3168 &  n_8369;
assign n_8707 =  i_8 & ~n_8368;
assign n_8708 =  x_2130 &  n_8346;
assign n_8709 =  x_1170 &  n_8355;
assign n_8710 = ~n_8708 & ~n_8709;
assign n_8711 =  x_2258 &  n_8349;
assign n_8712 =  x_1202 &  n_8351;
assign n_8713 = ~n_8711 & ~n_8712;
assign n_8714 =  n_8710 &  n_8713;
assign n_8715 = ~n_8707 &  n_8714;
assign n_8716 = ~n_8706 &  n_8715;
assign n_8717 =  x_3168 & ~n_8716;
assign n_8718 = ~x_3168 &  n_8716;
assign n_8719 = ~n_8717 & ~n_8718;
assign n_8720 =  x_3167 &  n_8369;
assign n_8721 =  i_7 & ~n_8368;
assign n_8722 =  x_2129 &  n_8346;
assign n_8723 =  x_1169 &  n_8355;
assign n_8724 = ~n_8722 & ~n_8723;
assign n_8725 =  x_2257 &  n_8349;
assign n_8726 =  x_1201 &  n_8351;
assign n_8727 = ~n_8725 & ~n_8726;
assign n_8728 =  n_8724 &  n_8727;
assign n_8729 = ~n_8721 &  n_8728;
assign n_8730 = ~n_8720 &  n_8729;
assign n_8731 =  x_3167 & ~n_8730;
assign n_8732 = ~x_3167 &  n_8730;
assign n_8733 = ~n_8731 & ~n_8732;
assign n_8734 =  x_3166 &  n_8369;
assign n_8735 =  i_6 & ~n_8368;
assign n_8736 =  x_2128 &  n_8346;
assign n_8737 =  x_1168 &  n_8355;
assign n_8738 = ~n_8736 & ~n_8737;
assign n_8739 =  x_2256 &  n_8349;
assign n_8740 =  x_1200 &  n_8351;
assign n_8741 = ~n_8739 & ~n_8740;
assign n_8742 =  n_8738 &  n_8741;
assign n_8743 = ~n_8735 &  n_8742;
assign n_8744 = ~n_8734 &  n_8743;
assign n_8745 =  x_3166 & ~n_8744;
assign n_8746 = ~x_3166 &  n_8744;
assign n_8747 = ~n_8745 & ~n_8746;
assign n_8748 =  x_3165 &  n_8369;
assign n_8749 =  i_5 & ~n_8368;
assign n_8750 =  x_2127 &  n_8346;
assign n_8751 =  x_1167 &  n_8355;
assign n_8752 = ~n_8750 & ~n_8751;
assign n_8753 =  x_2255 &  n_8349;
assign n_8754 =  x_1199 &  n_8351;
assign n_8755 = ~n_8753 & ~n_8754;
assign n_8756 =  n_8752 &  n_8755;
assign n_8757 = ~n_8749 &  n_8756;
assign n_8758 = ~n_8748 &  n_8757;
assign n_8759 =  x_3165 & ~n_8758;
assign n_8760 = ~x_3165 &  n_8758;
assign n_8761 = ~n_8759 & ~n_8760;
assign n_8762 =  x_3164 &  n_8369;
assign n_8763 =  i_4 & ~n_8368;
assign n_8764 =  x_2126 &  n_8346;
assign n_8765 =  x_1166 &  n_8355;
assign n_8766 = ~n_8764 & ~n_8765;
assign n_8767 =  x_2254 &  n_8349;
assign n_8768 =  x_1198 &  n_8351;
assign n_8769 = ~n_8767 & ~n_8768;
assign n_8770 =  n_8766 &  n_8769;
assign n_8771 = ~n_8763 &  n_8770;
assign n_8772 = ~n_8762 &  n_8771;
assign n_8773 =  x_3164 & ~n_8772;
assign n_8774 = ~x_3164 &  n_8772;
assign n_8775 = ~n_8773 & ~n_8774;
assign n_8776 =  x_3163 &  n_8369;
assign n_8777 =  i_3 & ~n_8368;
assign n_8778 =  x_2125 &  n_8346;
assign n_8779 =  x_1165 &  n_8355;
assign n_8780 = ~n_8778 & ~n_8779;
assign n_8781 =  x_2253 &  n_8349;
assign n_8782 =  x_1197 &  n_8351;
assign n_8783 = ~n_8781 & ~n_8782;
assign n_8784 =  n_8780 &  n_8783;
assign n_8785 = ~n_8777 &  n_8784;
assign n_8786 = ~n_8776 &  n_8785;
assign n_8787 =  x_3163 & ~n_8786;
assign n_8788 = ~x_3163 &  n_8786;
assign n_8789 = ~n_8787 & ~n_8788;
assign n_8790 =  x_3162 &  n_8369;
assign n_8791 =  i_2 & ~n_8368;
assign n_8792 =  x_2124 &  n_8346;
assign n_8793 =  x_1164 &  n_8355;
assign n_8794 = ~n_8792 & ~n_8793;
assign n_8795 =  x_2252 &  n_8349;
assign n_8796 =  x_1196 &  n_8351;
assign n_8797 = ~n_8795 & ~n_8796;
assign n_8798 =  n_8794 &  n_8797;
assign n_8799 = ~n_8791 &  n_8798;
assign n_8800 = ~n_8790 &  n_8799;
assign n_8801 =  x_3162 & ~n_8800;
assign n_8802 = ~x_3162 &  n_8800;
assign n_8803 = ~n_8801 & ~n_8802;
assign n_8804 =  x_3161 &  n_8369;
assign n_8805 =  i_1 & ~n_8368;
assign n_8806 =  x_2123 &  n_8346;
assign n_8807 =  x_1163 &  n_8355;
assign n_8808 = ~n_8806 & ~n_8807;
assign n_8809 =  x_2251 &  n_8349;
assign n_8810 =  x_1195 &  n_8351;
assign n_8811 = ~n_8809 & ~n_8810;
assign n_8812 =  n_8808 &  n_8811;
assign n_8813 = ~n_8805 &  n_8812;
assign n_8814 = ~n_8804 &  n_8813;
assign n_8815 =  x_3161 & ~n_8814;
assign n_8816 = ~x_3161 &  n_8814;
assign n_8817 = ~n_8815 & ~n_8816;
assign n_8818 =  n_1038 &  n_1305;
assign n_8819 =  n_8818 &  n_8354;
assign n_8820 =  x_3160 & ~n_8819;
assign n_8821 =  x_3160 &  n_8820;
assign n_8822 = ~x_3160 & ~n_8820;
assign n_8823 = ~n_8821 & ~n_8822;
assign n_8824 =  x_3159 & ~n_8819;
assign n_8825 =  x_3159 &  n_8824;
assign n_8826 = ~x_3159 & ~n_8824;
assign n_8827 = ~n_8825 & ~n_8826;
assign n_8828 =  x_3158 & ~n_8819;
assign n_8829 =  x_3158 &  n_8828;
assign n_8830 = ~x_3158 & ~n_8828;
assign n_8831 = ~n_8829 & ~n_8830;
assign n_8832 =  x_3157 & ~n_8819;
assign n_8833 =  x_3157 &  n_8832;
assign n_8834 = ~x_3157 & ~n_8832;
assign n_8835 = ~n_8833 & ~n_8834;
assign n_8836 =  x_3156 & ~n_8819;
assign n_8837 =  x_3156 &  n_8836;
assign n_8838 = ~x_3156 & ~n_8836;
assign n_8839 = ~n_8837 & ~n_8838;
assign n_8840 =  x_3155 & ~n_8819;
assign n_8841 =  x_3155 &  n_8840;
assign n_8842 = ~x_3155 & ~n_8840;
assign n_8843 = ~n_8841 & ~n_8842;
assign n_8844 =  x_3154 & ~n_8819;
assign n_8845 =  x_3154 &  n_8844;
assign n_8846 = ~x_3154 & ~n_8844;
assign n_8847 = ~n_8845 & ~n_8846;
assign n_8848 =  x_3153 & ~n_8819;
assign n_8849 =  x_3153 &  n_8848;
assign n_8850 = ~x_3153 & ~n_8848;
assign n_8851 = ~n_8849 & ~n_8850;
assign n_8852 =  x_3152 & ~n_8819;
assign n_8853 =  x_3152 &  n_8852;
assign n_8854 = ~x_3152 & ~n_8852;
assign n_8855 = ~n_8853 & ~n_8854;
assign n_8856 =  x_3151 & ~n_8819;
assign n_8857 =  x_3151 &  n_8856;
assign n_8858 = ~x_3151 & ~n_8856;
assign n_8859 = ~n_8857 & ~n_8858;
assign n_8860 =  x_3150 & ~n_8819;
assign n_8861 =  x_3150 &  n_8860;
assign n_8862 = ~x_3150 & ~n_8860;
assign n_8863 = ~n_8861 & ~n_8862;
assign n_8864 =  x_3149 & ~n_8819;
assign n_8865 =  x_3149 &  n_8864;
assign n_8866 = ~x_3149 & ~n_8864;
assign n_8867 = ~n_8865 & ~n_8866;
assign n_8868 =  x_3148 & ~n_8819;
assign n_8869 =  x_3148 &  n_8868;
assign n_8870 = ~x_3148 & ~n_8868;
assign n_8871 = ~n_8869 & ~n_8870;
assign n_8872 =  x_3147 & ~n_8819;
assign n_8873 =  x_3147 &  n_8872;
assign n_8874 = ~x_3147 & ~n_8872;
assign n_8875 = ~n_8873 & ~n_8874;
assign n_8876 =  x_3146 & ~n_8819;
assign n_8877 =  x_3146 &  n_8876;
assign n_8878 = ~x_3146 & ~n_8876;
assign n_8879 = ~n_8877 & ~n_8878;
assign n_8880 =  x_3145 & ~n_8819;
assign n_8881 =  x_3145 &  n_8880;
assign n_8882 = ~x_3145 & ~n_8880;
assign n_8883 = ~n_8881 & ~n_8882;
assign n_8884 =  x_3144 & ~n_8819;
assign n_8885 =  x_3144 &  n_8884;
assign n_8886 = ~x_3144 & ~n_8884;
assign n_8887 = ~n_8885 & ~n_8886;
assign n_8888 =  x_3143 & ~n_8819;
assign n_8889 =  x_3143 &  n_8888;
assign n_8890 = ~x_3143 & ~n_8888;
assign n_8891 = ~n_8889 & ~n_8890;
assign n_8892 =  x_3142 & ~n_8819;
assign n_8893 =  x_3142 &  n_8892;
assign n_8894 = ~x_3142 & ~n_8892;
assign n_8895 = ~n_8893 & ~n_8894;
assign n_8896 =  x_3141 & ~n_8819;
assign n_8897 =  x_3141 &  n_8896;
assign n_8898 = ~x_3141 & ~n_8896;
assign n_8899 = ~n_8897 & ~n_8898;
assign n_8900 =  x_3140 & ~n_8819;
assign n_8901 =  x_3140 &  n_8900;
assign n_8902 = ~x_3140 & ~n_8900;
assign n_8903 = ~n_8901 & ~n_8902;
assign n_8904 =  x_3139 & ~n_8819;
assign n_8905 =  x_3139 &  n_8904;
assign n_8906 = ~x_3139 & ~n_8904;
assign n_8907 = ~n_8905 & ~n_8906;
assign n_8908 =  x_3138 & ~n_8819;
assign n_8909 =  x_3138 &  n_8908;
assign n_8910 = ~x_3138 & ~n_8908;
assign n_8911 = ~n_8909 & ~n_8910;
assign n_8912 =  x_3137 & ~n_8819;
assign n_8913 =  x_3137 &  n_8912;
assign n_8914 = ~x_3137 & ~n_8912;
assign n_8915 = ~n_8913 & ~n_8914;
assign n_8916 =  x_3136 & ~n_8819;
assign n_8917 =  x_3136 &  n_8916;
assign n_8918 = ~x_3136 & ~n_8916;
assign n_8919 = ~n_8917 & ~n_8918;
assign n_8920 =  x_3135 & ~n_8819;
assign n_8921 =  x_3135 &  n_8920;
assign n_8922 = ~x_3135 & ~n_8920;
assign n_8923 = ~n_8921 & ~n_8922;
assign n_8924 =  x_3134 & ~n_8819;
assign n_8925 =  x_3134 &  n_8924;
assign n_8926 = ~x_3134 & ~n_8924;
assign n_8927 = ~n_8925 & ~n_8926;
assign n_8928 =  x_3133 & ~n_8819;
assign n_8929 =  x_3133 &  n_8928;
assign n_8930 = ~x_3133 & ~n_8928;
assign n_8931 = ~n_8929 & ~n_8930;
assign n_8932 =  x_3132 & ~n_8819;
assign n_8933 =  x_3132 &  n_8932;
assign n_8934 = ~x_3132 & ~n_8932;
assign n_8935 = ~n_8933 & ~n_8934;
assign n_8936 =  x_3131 & ~n_8819;
assign n_8937 =  x_3131 &  n_8936;
assign n_8938 = ~x_3131 & ~n_8936;
assign n_8939 = ~n_8937 & ~n_8938;
assign n_8940 =  x_3130 & ~n_8819;
assign n_8941 =  x_3130 &  n_8940;
assign n_8942 = ~x_3130 & ~n_8940;
assign n_8943 = ~n_8941 & ~n_8942;
assign n_8944 =  x_3129 & ~n_8819;
assign n_8945 =  x_3129 &  n_8944;
assign n_8946 = ~x_3129 & ~n_8944;
assign n_8947 = ~n_8945 & ~n_8946;
assign n_8948 =  x_3128 & ~n_7274;
assign n_8949 = ~n_7275 & ~n_8948;
assign n_8950 =  x_3128 & ~n_8949;
assign n_8951 = ~x_3128 &  n_8949;
assign n_8952 = ~n_8950 & ~n_8951;
assign n_8953 =  x_3127 & ~n_7274;
assign n_8954 = ~n_7281 & ~n_8953;
assign n_8955 =  x_3127 & ~n_8954;
assign n_8956 = ~x_3127 &  n_8954;
assign n_8957 = ~n_8955 & ~n_8956;
assign n_8958 =  x_3126 & ~n_7274;
assign n_8959 = ~n_7287 & ~n_8958;
assign n_8960 =  x_3126 & ~n_8959;
assign n_8961 = ~x_3126 &  n_8959;
assign n_8962 = ~n_8960 & ~n_8961;
assign n_8963 =  x_3125 & ~n_7274;
assign n_8964 = ~n_7293 & ~n_8963;
assign n_8965 =  x_3125 & ~n_8964;
assign n_8966 = ~x_3125 &  n_8964;
assign n_8967 = ~n_8965 & ~n_8966;
assign n_8968 =  x_3124 & ~n_7274;
assign n_8969 = ~n_7299 & ~n_8968;
assign n_8970 =  x_3124 & ~n_8969;
assign n_8971 = ~x_3124 &  n_8969;
assign n_8972 = ~n_8970 & ~n_8971;
assign n_8973 =  x_3123 & ~n_7274;
assign n_8974 = ~n_7305 & ~n_8973;
assign n_8975 =  x_3123 & ~n_8974;
assign n_8976 = ~x_3123 &  n_8974;
assign n_8977 = ~n_8975 & ~n_8976;
assign n_8978 =  x_3122 & ~n_7274;
assign n_8979 = ~n_7311 & ~n_8978;
assign n_8980 =  x_3122 & ~n_8979;
assign n_8981 = ~x_3122 &  n_8979;
assign n_8982 = ~n_8980 & ~n_8981;
assign n_8983 =  x_3121 & ~n_7274;
assign n_8984 = ~n_7317 & ~n_8983;
assign n_8985 =  x_3121 & ~n_8984;
assign n_8986 = ~x_3121 &  n_8984;
assign n_8987 = ~n_8985 & ~n_8986;
assign n_8988 =  x_3120 & ~n_7274;
assign n_8989 = ~n_7323 & ~n_8988;
assign n_8990 =  x_3120 & ~n_8989;
assign n_8991 = ~x_3120 &  n_8989;
assign n_8992 = ~n_8990 & ~n_8991;
assign n_8993 =  x_3119 & ~n_7274;
assign n_8994 = ~n_7329 & ~n_8993;
assign n_8995 =  x_3119 & ~n_8994;
assign n_8996 = ~x_3119 &  n_8994;
assign n_8997 = ~n_8995 & ~n_8996;
assign n_8998 =  x_3118 & ~n_7274;
assign n_8999 = ~n_7335 & ~n_8998;
assign n_9000 =  x_3118 & ~n_8999;
assign n_9001 = ~x_3118 &  n_8999;
assign n_9002 = ~n_9000 & ~n_9001;
assign n_9003 =  x_3117 & ~n_7274;
assign n_9004 = ~n_7341 & ~n_9003;
assign n_9005 =  x_3117 & ~n_9004;
assign n_9006 = ~x_3117 &  n_9004;
assign n_9007 = ~n_9005 & ~n_9006;
assign n_9008 =  x_3116 & ~n_7274;
assign n_9009 = ~n_7347 & ~n_9008;
assign n_9010 =  x_3116 & ~n_9009;
assign n_9011 = ~x_3116 &  n_9009;
assign n_9012 = ~n_9010 & ~n_9011;
assign n_9013 =  x_3115 & ~n_7274;
assign n_9014 = ~n_7353 & ~n_9013;
assign n_9015 =  x_3115 & ~n_9014;
assign n_9016 = ~x_3115 &  n_9014;
assign n_9017 = ~n_9015 & ~n_9016;
assign n_9018 =  x_3114 & ~n_7274;
assign n_9019 = ~n_7359 & ~n_9018;
assign n_9020 =  x_3114 & ~n_9019;
assign n_9021 = ~x_3114 &  n_9019;
assign n_9022 = ~n_9020 & ~n_9021;
assign n_9023 =  x_3113 & ~n_7274;
assign n_9024 = ~n_7365 & ~n_9023;
assign n_9025 =  x_3113 & ~n_9024;
assign n_9026 = ~x_3113 &  n_9024;
assign n_9027 = ~n_9025 & ~n_9026;
assign n_9028 =  x_3112 & ~n_7274;
assign n_9029 = ~n_7371 & ~n_9028;
assign n_9030 =  x_3112 & ~n_9029;
assign n_9031 = ~x_3112 &  n_9029;
assign n_9032 = ~n_9030 & ~n_9031;
assign n_9033 =  x_3111 & ~n_7274;
assign n_9034 = ~n_7377 & ~n_9033;
assign n_9035 =  x_3111 & ~n_9034;
assign n_9036 = ~x_3111 &  n_9034;
assign n_9037 = ~n_9035 & ~n_9036;
assign n_9038 =  x_3110 & ~n_7274;
assign n_9039 = ~n_7383 & ~n_9038;
assign n_9040 =  x_3110 & ~n_9039;
assign n_9041 = ~x_3110 &  n_9039;
assign n_9042 = ~n_9040 & ~n_9041;
assign n_9043 =  x_3109 & ~n_7274;
assign n_9044 = ~n_7389 & ~n_9043;
assign n_9045 =  x_3109 & ~n_9044;
assign n_9046 = ~x_3109 &  n_9044;
assign n_9047 = ~n_9045 & ~n_9046;
assign n_9048 =  x_3108 & ~n_7274;
assign n_9049 = ~n_7395 & ~n_9048;
assign n_9050 =  x_3108 & ~n_9049;
assign n_9051 = ~x_3108 &  n_9049;
assign n_9052 = ~n_9050 & ~n_9051;
assign n_9053 =  x_3107 & ~n_7274;
assign n_9054 = ~n_7401 & ~n_9053;
assign n_9055 =  x_3107 & ~n_9054;
assign n_9056 = ~x_3107 &  n_9054;
assign n_9057 = ~n_9055 & ~n_9056;
assign n_9058 =  x_3106 & ~n_7274;
assign n_9059 = ~n_7407 & ~n_9058;
assign n_9060 =  x_3106 & ~n_9059;
assign n_9061 = ~x_3106 &  n_9059;
assign n_9062 = ~n_9060 & ~n_9061;
assign n_9063 =  x_3105 & ~n_7274;
assign n_9064 = ~n_7413 & ~n_9063;
assign n_9065 =  x_3105 & ~n_9064;
assign n_9066 = ~x_3105 &  n_9064;
assign n_9067 = ~n_9065 & ~n_9066;
assign n_9068 =  x_3104 & ~n_7274;
assign n_9069 = ~n_7419 & ~n_9068;
assign n_9070 =  x_3104 & ~n_9069;
assign n_9071 = ~x_3104 &  n_9069;
assign n_9072 = ~n_9070 & ~n_9071;
assign n_9073 =  x_3103 & ~n_7274;
assign n_9074 = ~n_7425 & ~n_9073;
assign n_9075 =  x_3103 & ~n_9074;
assign n_9076 = ~x_3103 &  n_9074;
assign n_9077 = ~n_9075 & ~n_9076;
assign n_9078 =  x_3102 & ~n_7274;
assign n_9079 = ~n_7431 & ~n_9078;
assign n_9080 =  x_3102 & ~n_9079;
assign n_9081 = ~x_3102 &  n_9079;
assign n_9082 = ~n_9080 & ~n_9081;
assign n_9083 =  x_3101 & ~n_7274;
assign n_9084 = ~n_7437 & ~n_9083;
assign n_9085 =  x_3101 & ~n_9084;
assign n_9086 = ~x_3101 &  n_9084;
assign n_9087 = ~n_9085 & ~n_9086;
assign n_9088 =  x_3100 & ~n_7274;
assign n_9089 = ~n_7443 & ~n_9088;
assign n_9090 =  x_3100 & ~n_9089;
assign n_9091 = ~x_3100 &  n_9089;
assign n_9092 = ~n_9090 & ~n_9091;
assign n_9093 =  x_3099 & ~n_7274;
assign n_9094 = ~n_7449 & ~n_9093;
assign n_9095 =  x_3099 & ~n_9094;
assign n_9096 = ~x_3099 &  n_9094;
assign n_9097 = ~n_9095 & ~n_9096;
assign n_9098 =  x_3098 & ~n_7274;
assign n_9099 = ~n_7455 & ~n_9098;
assign n_9100 =  x_3098 & ~n_9099;
assign n_9101 = ~x_3098 &  n_9099;
assign n_9102 = ~n_9100 & ~n_9101;
assign n_9103 =  x_3097 & ~n_7274;
assign n_9104 = ~n_7461 & ~n_9103;
assign n_9105 =  x_3097 & ~n_9104;
assign n_9106 = ~x_3097 &  n_9104;
assign n_9107 = ~n_9105 & ~n_9106;
assign n_9108 =  x_3255 &  n_558;
assign n_9109 =  x_3096 & ~n_564;
assign n_9110 = ~n_9108 & ~n_9109;
assign n_9111 =  x_3096 & ~n_9110;
assign n_9112 = ~x_3096 &  n_9110;
assign n_9113 = ~n_9111 & ~n_9112;
assign n_9114 =  x_3254 &  n_558;
assign n_9115 =  x_3095 & ~n_564;
assign n_9116 = ~n_9114 & ~n_9115;
assign n_9117 =  x_3095 & ~n_9116;
assign n_9118 = ~x_3095 &  n_9116;
assign n_9119 = ~n_9117 & ~n_9118;
assign n_9120 =  x_3253 &  n_558;
assign n_9121 =  x_3094 & ~n_564;
assign n_9122 = ~n_9120 & ~n_9121;
assign n_9123 =  x_3094 & ~n_9122;
assign n_9124 = ~x_3094 &  n_9122;
assign n_9125 = ~n_9123 & ~n_9124;
assign n_9126 =  x_3252 &  n_558;
assign n_9127 =  x_3093 & ~n_564;
assign n_9128 = ~n_9126 & ~n_9127;
assign n_9129 =  x_3093 & ~n_9128;
assign n_9130 = ~x_3093 &  n_9128;
assign n_9131 = ~n_9129 & ~n_9130;
assign n_9132 =  x_3251 &  n_558;
assign n_9133 =  x_3092 & ~n_564;
assign n_9134 = ~n_9132 & ~n_9133;
assign n_9135 =  x_3092 & ~n_9134;
assign n_9136 = ~x_3092 &  n_9134;
assign n_9137 = ~n_9135 & ~n_9136;
assign n_9138 =  x_3250 &  n_558;
assign n_9139 =  x_3091 & ~n_564;
assign n_9140 = ~n_9138 & ~n_9139;
assign n_9141 =  x_3091 & ~n_9140;
assign n_9142 = ~x_3091 &  n_9140;
assign n_9143 = ~n_9141 & ~n_9142;
assign n_9144 =  x_3249 &  n_558;
assign n_9145 =  x_3090 & ~n_564;
assign n_9146 = ~n_9144 & ~n_9145;
assign n_9147 =  x_3090 & ~n_9146;
assign n_9148 = ~x_3090 &  n_9146;
assign n_9149 = ~n_9147 & ~n_9148;
assign n_9150 =  x_3248 &  n_558;
assign n_9151 =  x_3089 & ~n_564;
assign n_9152 = ~n_9150 & ~n_9151;
assign n_9153 =  x_3089 & ~n_9152;
assign n_9154 = ~x_3089 &  n_9152;
assign n_9155 = ~n_9153 & ~n_9154;
assign n_9156 =  x_3247 &  n_558;
assign n_9157 =  x_3088 & ~n_564;
assign n_9158 = ~n_9156 & ~n_9157;
assign n_9159 =  x_3088 & ~n_9158;
assign n_9160 = ~x_3088 &  n_9158;
assign n_9161 = ~n_9159 & ~n_9160;
assign n_9162 =  x_3246 &  n_558;
assign n_9163 =  x_3087 & ~n_564;
assign n_9164 = ~n_9162 & ~n_9163;
assign n_9165 =  x_3087 & ~n_9164;
assign n_9166 = ~x_3087 &  n_9164;
assign n_9167 = ~n_9165 & ~n_9166;
assign n_9168 =  x_3245 &  n_558;
assign n_9169 =  x_3086 & ~n_564;
assign n_9170 = ~n_9168 & ~n_9169;
assign n_9171 =  x_3086 & ~n_9170;
assign n_9172 = ~x_3086 &  n_9170;
assign n_9173 = ~n_9171 & ~n_9172;
assign n_9174 =  x_3244 &  n_558;
assign n_9175 =  x_3085 & ~n_564;
assign n_9176 = ~n_9174 & ~n_9175;
assign n_9177 =  x_3085 & ~n_9176;
assign n_9178 = ~x_3085 &  n_9176;
assign n_9179 = ~n_9177 & ~n_9178;
assign n_9180 =  x_3243 &  n_558;
assign n_9181 =  x_3084 & ~n_564;
assign n_9182 = ~n_9180 & ~n_9181;
assign n_9183 =  x_3084 & ~n_9182;
assign n_9184 = ~x_3084 &  n_9182;
assign n_9185 = ~n_9183 & ~n_9184;
assign n_9186 =  x_3242 &  n_558;
assign n_9187 =  x_3083 & ~n_564;
assign n_9188 = ~n_9186 & ~n_9187;
assign n_9189 =  x_3083 & ~n_9188;
assign n_9190 = ~x_3083 &  n_9188;
assign n_9191 = ~n_9189 & ~n_9190;
assign n_9192 =  x_3241 &  n_558;
assign n_9193 =  x_3082 & ~n_564;
assign n_9194 = ~n_9192 & ~n_9193;
assign n_9195 =  x_3082 & ~n_9194;
assign n_9196 = ~x_3082 &  n_9194;
assign n_9197 = ~n_9195 & ~n_9196;
assign n_9198 =  x_3240 &  n_558;
assign n_9199 =  x_3081 & ~n_564;
assign n_9200 = ~n_9198 & ~n_9199;
assign n_9201 =  x_3081 & ~n_9200;
assign n_9202 = ~x_3081 &  n_9200;
assign n_9203 = ~n_9201 & ~n_9202;
assign n_9204 =  x_3239 &  n_558;
assign n_9205 =  x_3080 & ~n_564;
assign n_9206 = ~n_9204 & ~n_9205;
assign n_9207 =  x_3080 & ~n_9206;
assign n_9208 = ~x_3080 &  n_9206;
assign n_9209 = ~n_9207 & ~n_9208;
assign n_9210 =  x_3238 &  n_558;
assign n_9211 =  x_3079 & ~n_564;
assign n_9212 = ~n_9210 & ~n_9211;
assign n_9213 =  x_3079 & ~n_9212;
assign n_9214 = ~x_3079 &  n_9212;
assign n_9215 = ~n_9213 & ~n_9214;
assign n_9216 =  x_3237 &  n_558;
assign n_9217 =  x_3078 & ~n_564;
assign n_9218 = ~n_9216 & ~n_9217;
assign n_9219 =  x_3078 & ~n_9218;
assign n_9220 = ~x_3078 &  n_9218;
assign n_9221 = ~n_9219 & ~n_9220;
assign n_9222 =  x_3236 &  n_558;
assign n_9223 =  x_3077 & ~n_564;
assign n_9224 = ~n_9222 & ~n_9223;
assign n_9225 =  x_3077 & ~n_9224;
assign n_9226 = ~x_3077 &  n_9224;
assign n_9227 = ~n_9225 & ~n_9226;
assign n_9228 =  x_3235 &  n_558;
assign n_9229 =  x_3076 & ~n_564;
assign n_9230 = ~n_9228 & ~n_9229;
assign n_9231 =  x_3076 & ~n_9230;
assign n_9232 = ~x_3076 &  n_9230;
assign n_9233 = ~n_9231 & ~n_9232;
assign n_9234 =  x_3234 &  n_558;
assign n_9235 =  x_3075 & ~n_564;
assign n_9236 = ~n_9234 & ~n_9235;
assign n_9237 =  x_3075 & ~n_9236;
assign n_9238 = ~x_3075 &  n_9236;
assign n_9239 = ~n_9237 & ~n_9238;
assign n_9240 =  x_3233 &  n_558;
assign n_9241 =  x_3074 & ~n_564;
assign n_9242 = ~n_9240 & ~n_9241;
assign n_9243 =  x_3074 & ~n_9242;
assign n_9244 = ~x_3074 &  n_9242;
assign n_9245 = ~n_9243 & ~n_9244;
assign n_9246 =  x_3232 &  n_558;
assign n_9247 =  x_3073 & ~n_564;
assign n_9248 = ~n_9246 & ~n_9247;
assign n_9249 =  x_3073 & ~n_9248;
assign n_9250 = ~x_3073 &  n_9248;
assign n_9251 = ~n_9249 & ~n_9250;
assign n_9252 =  x_3231 &  n_558;
assign n_9253 =  x_3072 & ~n_564;
assign n_9254 = ~n_9252 & ~n_9253;
assign n_9255 =  x_3072 & ~n_9254;
assign n_9256 = ~x_3072 &  n_9254;
assign n_9257 = ~n_9255 & ~n_9256;
assign n_9258 =  x_3230 &  n_558;
assign n_9259 =  x_3071 & ~n_564;
assign n_9260 = ~n_9258 & ~n_9259;
assign n_9261 =  x_3071 & ~n_9260;
assign n_9262 = ~x_3071 &  n_9260;
assign n_9263 = ~n_9261 & ~n_9262;
assign n_9264 =  x_3229 &  n_558;
assign n_9265 =  x_3070 & ~n_564;
assign n_9266 = ~n_9264 & ~n_9265;
assign n_9267 =  x_3070 & ~n_9266;
assign n_9268 = ~x_3070 &  n_9266;
assign n_9269 = ~n_9267 & ~n_9268;
assign n_9270 =  x_3228 &  n_558;
assign n_9271 =  x_3069 & ~n_564;
assign n_9272 = ~n_9270 & ~n_9271;
assign n_9273 =  x_3069 & ~n_9272;
assign n_9274 = ~x_3069 &  n_9272;
assign n_9275 = ~n_9273 & ~n_9274;
assign n_9276 =  x_3227 &  n_558;
assign n_9277 =  x_3068 & ~n_564;
assign n_9278 = ~n_9276 & ~n_9277;
assign n_9279 =  x_3068 & ~n_9278;
assign n_9280 = ~x_3068 &  n_9278;
assign n_9281 = ~n_9279 & ~n_9280;
assign n_9282 =  x_3226 &  n_558;
assign n_9283 =  x_3067 & ~n_564;
assign n_9284 = ~n_9282 & ~n_9283;
assign n_9285 =  x_3067 & ~n_9284;
assign n_9286 = ~x_3067 &  n_9284;
assign n_9287 = ~n_9285 & ~n_9286;
assign n_9288 =  x_3225 &  n_558;
assign n_9289 =  x_3066 & ~n_564;
assign n_9290 = ~n_9288 & ~n_9289;
assign n_9291 =  x_3066 & ~n_9290;
assign n_9292 = ~x_3066 &  n_9290;
assign n_9293 = ~n_9291 & ~n_9292;
assign n_9294 =  x_3224 &  n_558;
assign n_9295 =  x_3065 & ~n_564;
assign n_9296 = ~n_9294 & ~n_9295;
assign n_9297 =  x_3065 & ~n_9296;
assign n_9298 = ~x_3065 &  n_9296;
assign n_9299 = ~n_9297 & ~n_9298;
assign n_9300 =  n_349 &  n_770;
assign n_9301 =  x_1599 & ~x_3085;
assign n_9302 = ~x_1599 &  x_3085;
assign n_9303 = ~n_9301 & ~n_9302;
assign n_9304 =  x_1610 & ~x_3096;
assign n_9305 = ~x_1610 &  x_3096;
assign n_9306 = ~n_9304 & ~n_9305;
assign n_9307 =  n_9303 &  n_9306;
assign n_9308 = ~x_1589 &  x_3075;
assign n_9309 = ~x_1580 &  x_3066;
assign n_9310 = ~n_9308 & ~n_9309;
assign n_9311 =  x_1607 & ~x_3093;
assign n_9312 =  x_1580 & ~x_3066;
assign n_9313 = ~n_9311 & ~n_9312;
assign n_9314 =  n_9310 &  n_9313;
assign n_9315 =  n_9307 &  n_9314;
assign n_9316 =  x_1582 & ~x_3068;
assign n_9317 =  x_1581 & ~x_3067;
assign n_9318 = ~n_9316 & ~n_9317;
assign n_9319 =  x_1590 & ~x_3076;
assign n_9320 = ~x_1590 &  x_3076;
assign n_9321 = ~n_9319 & ~n_9320;
assign n_9322 =  n_9318 &  n_9321;
assign n_9323 = ~x_1581 &  x_3067;
assign n_9324 = ~x_1592 &  x_3078;
assign n_9325 = ~n_9323 & ~n_9324;
assign n_9326 = ~x_1607 &  x_3093;
assign n_9327 =  x_1592 & ~x_3078;
assign n_9328 = ~n_9326 & ~n_9327;
assign n_9329 =  n_9325 &  n_9328;
assign n_9330 =  n_9322 &  n_9329;
assign n_9331 =  n_9315 &  n_9330;
assign n_9332 = ~x_1583 & ~x_3069;
assign n_9333 =  x_1583 &  x_3069;
assign n_9334 = ~n_9332 & ~n_9333;
assign n_9335 = ~x_1603 & ~x_3089;
assign n_9336 =  x_1603 &  x_3089;
assign n_9337 = ~n_9335 & ~n_9336;
assign n_9338 = ~n_9334 & ~n_9337;
assign n_9339 = ~x_1585 & ~x_3071;
assign n_9340 =  x_1585 &  x_3071;
assign n_9341 = ~n_9339 & ~n_9340;
assign n_9342 = ~x_1605 & ~x_3091;
assign n_9343 =  x_1605 &  x_3091;
assign n_9344 = ~n_9342 & ~n_9343;
assign n_9345 = ~n_9341 & ~n_9344;
assign n_9346 =  n_9338 &  n_9345;
assign n_9347 = ~x_1602 & ~x_3088;
assign n_9348 =  x_1602 &  x_3088;
assign n_9349 = ~n_9347 & ~n_9348;
assign n_9350 = ~x_1600 & ~x_3086;
assign n_9351 =  x_1600 &  x_3086;
assign n_9352 = ~n_9350 & ~n_9351;
assign n_9353 = ~n_9349 & ~n_9352;
assign n_9354 = ~x_1596 & ~x_3082;
assign n_9355 =  x_1596 &  x_3082;
assign n_9356 = ~n_9354 & ~n_9355;
assign n_9357 = ~x_1608 & ~x_3094;
assign n_9358 =  x_1608 &  x_3094;
assign n_9359 = ~n_9357 & ~n_9358;
assign n_9360 = ~n_9356 & ~n_9359;
assign n_9361 =  n_9353 &  n_9360;
assign n_9362 =  n_9346 &  n_9361;
assign n_9363 =  n_9331 &  n_9362;
assign n_9364 =  x_1601 & ~x_3087;
assign n_9365 = ~x_1601 &  x_3087;
assign n_9366 = ~n_9364 & ~n_9365;
assign n_9367 = ~x_1606 &  x_3092;
assign n_9368 =  x_1604 & ~x_3090;
assign n_9369 = ~n_9367 & ~n_9368;
assign n_9370 =  n_9366 &  n_9369;
assign n_9371 =  x_1594 & ~x_3080;
assign n_9372 =  x_1606 & ~x_3092;
assign n_9373 = ~n_9371 & ~n_9372;
assign n_9374 =  x_1595 & ~x_3081;
assign n_9375 = ~x_1604 &  x_3090;
assign n_9376 = ~n_9374 & ~n_9375;
assign n_9377 =  n_9373 &  n_9376;
assign n_9378 =  n_9370 &  n_9377;
assign n_9379 =  x_1586 & ~x_3072;
assign n_9380 = ~x_1586 &  x_3072;
assign n_9381 = ~n_9379 & ~n_9380;
assign n_9382 = ~x_1582 &  x_3068;
assign n_9383 =  x_1589 & ~x_3075;
assign n_9384 = ~n_9382 & ~n_9383;
assign n_9385 =  n_9381 &  n_9384;
assign n_9386 =  x_1584 & ~x_3070;
assign n_9387 = ~x_1584 &  x_3070;
assign n_9388 = ~n_9386 & ~n_9387;
assign n_9389 =  x_1591 & ~x_3077;
assign n_9390 = ~x_1591 &  x_3077;
assign n_9391 = ~n_9389 & ~n_9390;
assign n_9392 =  n_9388 &  n_9391;
assign n_9393 =  n_9385 &  n_9392;
assign n_9394 =  n_9378 &  n_9393;
assign n_9395 = ~x_1595 &  x_3081;
assign n_9396 =  x_1579 & ~x_3065;
assign n_9397 = ~n_9395 & ~n_9396;
assign n_9398 = ~x_1579 &  x_3065;
assign n_9399 =  x_1593 & ~x_3079;
assign n_9400 = ~n_9398 & ~n_9399;
assign n_9401 =  n_9397 &  n_9400;
assign n_9402 =  x_1597 & ~x_3083;
assign n_9403 = ~x_1597 &  x_3083;
assign n_9404 = ~n_9402 & ~n_9403;
assign n_9405 =  x_1609 & ~x_3095;
assign n_9406 = ~x_1609 &  x_3095;
assign n_9407 = ~n_9405 & ~n_9406;
assign n_9408 =  n_9404 &  n_9407;
assign n_9409 =  n_9401 &  n_9408;
assign n_9410 =  x_1598 & ~x_3084;
assign n_9411 =  x_1588 & ~x_3074;
assign n_9412 = ~n_9410 & ~n_9411;
assign n_9413 = ~x_1594 &  x_3080;
assign n_9414 = ~x_1598 &  x_3084;
assign n_9415 = ~n_9413 & ~n_9414;
assign n_9416 =  n_9412 &  n_9415;
assign n_9417 = ~x_1593 &  x_3079;
assign n_9418 =  x_1587 & ~x_3073;
assign n_9419 = ~n_9417 & ~n_9418;
assign n_9420 = ~x_1587 &  x_3073;
assign n_9421 = ~x_1588 &  x_3074;
assign n_9422 = ~n_9420 & ~n_9421;
assign n_9423 =  n_9419 &  n_9422;
assign n_9424 =  n_9416 &  n_9423;
assign n_9425 =  n_9409 &  n_9424;
assign n_9426 =  n_9394 &  n_9425;
assign n_9427 =  n_9363 &  n_9426;
assign n_9428 =  n_9300 & ~n_9427;
assign n_9429 =  n_2 &  n_8049;
assign n_9430 = ~n_9300 & ~n_564;
assign n_9431 = ~n_9429 &  n_9430;
assign n_9432 = ~n_9428 & ~n_9431;
assign n_9433 =  x_2969 & ~n_9432;
assign n_9434 =  x_3255 &  n_9429;
assign n_9435 =  x_4487 &  n_558;
assign n_9436 = ~n_9434 & ~n_9435;
assign n_9437 = ~n_9433 &  n_9436;
assign n_9438 =  x_2969 & ~n_9437;
assign n_9439 = ~x_2969 &  n_9437;
assign n_9440 = ~n_9438 & ~n_9439;
assign n_9441 =  x_2968 & ~n_9432;
assign n_9442 =  x_3254 &  n_9429;
assign n_9443 =  x_4486 &  n_558;
assign n_9444 = ~n_9442 & ~n_9443;
assign n_9445 = ~n_9441 &  n_9444;
assign n_9446 =  x_2968 & ~n_9445;
assign n_9447 = ~x_2968 &  n_9445;
assign n_9448 = ~n_9446 & ~n_9447;
assign n_9449 =  x_2967 & ~n_9432;
assign n_9450 =  x_3253 &  n_9429;
assign n_9451 =  x_4485 &  n_558;
assign n_9452 = ~n_9450 & ~n_9451;
assign n_9453 = ~n_9449 &  n_9452;
assign n_9454 =  x_2967 & ~n_9453;
assign n_9455 = ~x_2967 &  n_9453;
assign n_9456 = ~n_9454 & ~n_9455;
assign n_9457 =  x_2966 & ~n_9432;
assign n_9458 =  x_3252 &  n_9429;
assign n_9459 =  x_4484 &  n_558;
assign n_9460 = ~n_9458 & ~n_9459;
assign n_9461 = ~n_9457 &  n_9460;
assign n_9462 =  x_2966 & ~n_9461;
assign n_9463 = ~x_2966 &  n_9461;
assign n_9464 = ~n_9462 & ~n_9463;
assign n_9465 =  x_2965 & ~n_9432;
assign n_9466 =  x_3251 &  n_9429;
assign n_9467 =  x_4483 &  n_558;
assign n_9468 = ~n_9466 & ~n_9467;
assign n_9469 = ~n_9465 &  n_9468;
assign n_9470 =  x_2965 & ~n_9469;
assign n_9471 = ~x_2965 &  n_9469;
assign n_9472 = ~n_9470 & ~n_9471;
assign n_9473 =  x_2964 & ~n_9432;
assign n_9474 =  x_3250 &  n_9429;
assign n_9475 =  x_4482 &  n_558;
assign n_9476 = ~n_9474 & ~n_9475;
assign n_9477 = ~n_9473 &  n_9476;
assign n_9478 =  x_2964 & ~n_9477;
assign n_9479 = ~x_2964 &  n_9477;
assign n_9480 = ~n_9478 & ~n_9479;
assign n_9481 =  x_2963 & ~n_9432;
assign n_9482 =  x_3249 &  n_9429;
assign n_9483 =  x_4481 &  n_558;
assign n_9484 = ~n_9482 & ~n_9483;
assign n_9485 = ~n_9481 &  n_9484;
assign n_9486 =  x_2963 & ~n_9485;
assign n_9487 = ~x_2963 &  n_9485;
assign n_9488 = ~n_9486 & ~n_9487;
assign n_9489 =  x_2962 & ~n_9432;
assign n_9490 =  x_3248 &  n_9429;
assign n_9491 =  x_4480 &  n_558;
assign n_9492 = ~n_9490 & ~n_9491;
assign n_9493 = ~n_9489 &  n_9492;
assign n_9494 =  x_2962 & ~n_9493;
assign n_9495 = ~x_2962 &  n_9493;
assign n_9496 = ~n_9494 & ~n_9495;
assign n_9497 =  x_2961 & ~n_9432;
assign n_9498 =  x_3247 &  n_9429;
assign n_9499 =  x_4479 &  n_558;
assign n_9500 = ~n_9498 & ~n_9499;
assign n_9501 = ~n_9497 &  n_9500;
assign n_9502 =  x_2961 & ~n_9501;
assign n_9503 = ~x_2961 &  n_9501;
assign n_9504 = ~n_9502 & ~n_9503;
assign n_9505 =  x_2960 & ~n_9432;
assign n_9506 =  x_3246 &  n_9429;
assign n_9507 =  x_4478 &  n_558;
assign n_9508 = ~n_9506 & ~n_9507;
assign n_9509 = ~n_9505 &  n_9508;
assign n_9510 =  x_2960 & ~n_9509;
assign n_9511 = ~x_2960 &  n_9509;
assign n_9512 = ~n_9510 & ~n_9511;
assign n_9513 =  x_2959 & ~n_9432;
assign n_9514 =  x_3245 &  n_9429;
assign n_9515 =  x_4477 &  n_558;
assign n_9516 = ~n_9514 & ~n_9515;
assign n_9517 = ~n_9513 &  n_9516;
assign n_9518 =  x_2959 & ~n_9517;
assign n_9519 = ~x_2959 &  n_9517;
assign n_9520 = ~n_9518 & ~n_9519;
assign n_9521 =  x_2958 & ~n_9432;
assign n_9522 =  x_3244 &  n_9429;
assign n_9523 =  x_4476 &  n_558;
assign n_9524 = ~n_9522 & ~n_9523;
assign n_9525 = ~n_9521 &  n_9524;
assign n_9526 =  x_2958 & ~n_9525;
assign n_9527 = ~x_2958 &  n_9525;
assign n_9528 = ~n_9526 & ~n_9527;
assign n_9529 =  x_2957 & ~n_9432;
assign n_9530 =  x_3243 &  n_9429;
assign n_9531 =  x_4475 &  n_558;
assign n_9532 = ~n_9530 & ~n_9531;
assign n_9533 = ~n_9529 &  n_9532;
assign n_9534 =  x_2957 & ~n_9533;
assign n_9535 = ~x_2957 &  n_9533;
assign n_9536 = ~n_9534 & ~n_9535;
assign n_9537 =  x_2956 & ~n_9432;
assign n_9538 =  x_3242 &  n_9429;
assign n_9539 =  x_4474 &  n_558;
assign n_9540 = ~n_9538 & ~n_9539;
assign n_9541 = ~n_9537 &  n_9540;
assign n_9542 =  x_2956 & ~n_9541;
assign n_9543 = ~x_2956 &  n_9541;
assign n_9544 = ~n_9542 & ~n_9543;
assign n_9545 =  x_2955 & ~n_9432;
assign n_9546 =  x_3241 &  n_9429;
assign n_9547 =  x_4473 &  n_558;
assign n_9548 = ~n_9546 & ~n_9547;
assign n_9549 = ~n_9545 &  n_9548;
assign n_9550 =  x_2955 & ~n_9549;
assign n_9551 = ~x_2955 &  n_9549;
assign n_9552 = ~n_9550 & ~n_9551;
assign n_9553 =  x_2954 & ~n_9432;
assign n_9554 =  x_3240 &  n_9429;
assign n_9555 =  x_4472 &  n_558;
assign n_9556 = ~n_9554 & ~n_9555;
assign n_9557 = ~n_9553 &  n_9556;
assign n_9558 =  x_2954 & ~n_9557;
assign n_9559 = ~x_2954 &  n_9557;
assign n_9560 = ~n_9558 & ~n_9559;
assign n_9561 =  x_2953 & ~n_9432;
assign n_9562 =  x_3239 &  n_9429;
assign n_9563 =  x_4471 &  n_558;
assign n_9564 = ~n_9562 & ~n_9563;
assign n_9565 = ~n_9561 &  n_9564;
assign n_9566 =  x_2953 & ~n_9565;
assign n_9567 = ~x_2953 &  n_9565;
assign n_9568 = ~n_9566 & ~n_9567;
assign n_9569 =  x_2952 & ~n_9432;
assign n_9570 =  x_3238 &  n_9429;
assign n_9571 =  x_4470 &  n_558;
assign n_9572 = ~n_9570 & ~n_9571;
assign n_9573 = ~n_9569 &  n_9572;
assign n_9574 =  x_2952 & ~n_9573;
assign n_9575 = ~x_2952 &  n_9573;
assign n_9576 = ~n_9574 & ~n_9575;
assign n_9577 =  x_2951 & ~n_9432;
assign n_9578 =  x_3237 &  n_9429;
assign n_9579 =  x_4469 &  n_558;
assign n_9580 = ~n_9578 & ~n_9579;
assign n_9581 = ~n_9577 &  n_9580;
assign n_9582 =  x_2951 & ~n_9581;
assign n_9583 = ~x_2951 &  n_9581;
assign n_9584 = ~n_9582 & ~n_9583;
assign n_9585 =  x_2950 & ~n_9432;
assign n_9586 =  x_3236 &  n_9429;
assign n_9587 =  x_4468 &  n_558;
assign n_9588 = ~n_9586 & ~n_9587;
assign n_9589 = ~n_9585 &  n_9588;
assign n_9590 =  x_2950 & ~n_9589;
assign n_9591 = ~x_2950 &  n_9589;
assign n_9592 = ~n_9590 & ~n_9591;
assign n_9593 =  x_2949 & ~n_9432;
assign n_9594 =  x_3235 &  n_9429;
assign n_9595 =  x_4467 &  n_558;
assign n_9596 = ~n_9594 & ~n_9595;
assign n_9597 = ~n_9593 &  n_9596;
assign n_9598 =  x_2949 & ~n_9597;
assign n_9599 = ~x_2949 &  n_9597;
assign n_9600 = ~n_9598 & ~n_9599;
assign n_9601 =  x_2948 & ~n_9432;
assign n_9602 =  x_3234 &  n_9429;
assign n_9603 =  x_4466 &  n_558;
assign n_9604 = ~n_9602 & ~n_9603;
assign n_9605 = ~n_9601 &  n_9604;
assign n_9606 =  x_2948 & ~n_9605;
assign n_9607 = ~x_2948 &  n_9605;
assign n_9608 = ~n_9606 & ~n_9607;
assign n_9609 =  x_2947 & ~n_9432;
assign n_9610 =  x_3233 &  n_9429;
assign n_9611 =  x_4465 &  n_558;
assign n_9612 = ~n_9610 & ~n_9611;
assign n_9613 = ~n_9609 &  n_9612;
assign n_9614 =  x_2947 & ~n_9613;
assign n_9615 = ~x_2947 &  n_9613;
assign n_9616 = ~n_9614 & ~n_9615;
assign n_9617 =  x_2946 & ~n_9432;
assign n_9618 =  x_3232 &  n_9429;
assign n_9619 =  x_4464 &  n_558;
assign n_9620 = ~n_9618 & ~n_9619;
assign n_9621 = ~n_9617 &  n_9620;
assign n_9622 =  x_2946 & ~n_9621;
assign n_9623 = ~x_2946 &  n_9621;
assign n_9624 = ~n_9622 & ~n_9623;
assign n_9625 =  x_2945 & ~n_9432;
assign n_9626 =  x_3231 &  n_9429;
assign n_9627 =  x_4463 &  n_558;
assign n_9628 = ~n_9626 & ~n_9627;
assign n_9629 = ~n_9625 &  n_9628;
assign n_9630 =  x_2945 & ~n_9629;
assign n_9631 = ~x_2945 &  n_9629;
assign n_9632 = ~n_9630 & ~n_9631;
assign n_9633 =  x_2944 & ~n_9432;
assign n_9634 =  x_3230 &  n_9429;
assign n_9635 =  x_4462 &  n_558;
assign n_9636 = ~n_9634 & ~n_9635;
assign n_9637 = ~n_9633 &  n_9636;
assign n_9638 =  x_2944 & ~n_9637;
assign n_9639 = ~x_2944 &  n_9637;
assign n_9640 = ~n_9638 & ~n_9639;
assign n_9641 =  x_2943 & ~n_9432;
assign n_9642 =  x_3229 &  n_9429;
assign n_9643 =  x_4461 &  n_558;
assign n_9644 = ~n_9642 & ~n_9643;
assign n_9645 = ~n_9641 &  n_9644;
assign n_9646 =  x_2943 & ~n_9645;
assign n_9647 = ~x_2943 &  n_9645;
assign n_9648 = ~n_9646 & ~n_9647;
assign n_9649 =  x_2942 & ~n_9432;
assign n_9650 =  x_3228 &  n_9429;
assign n_9651 =  x_4460 &  n_558;
assign n_9652 = ~n_9650 & ~n_9651;
assign n_9653 = ~n_9649 &  n_9652;
assign n_9654 =  x_2942 & ~n_9653;
assign n_9655 = ~x_2942 &  n_9653;
assign n_9656 = ~n_9654 & ~n_9655;
assign n_9657 =  x_2941 & ~n_9432;
assign n_9658 =  x_3227 &  n_9429;
assign n_9659 =  x_4459 &  n_558;
assign n_9660 = ~n_9658 & ~n_9659;
assign n_9661 = ~n_9657 &  n_9660;
assign n_9662 =  x_2941 & ~n_9661;
assign n_9663 = ~x_2941 &  n_9661;
assign n_9664 = ~n_9662 & ~n_9663;
assign n_9665 =  x_2940 & ~n_9432;
assign n_9666 =  x_3226 &  n_9429;
assign n_9667 =  x_4458 &  n_558;
assign n_9668 = ~n_9666 & ~n_9667;
assign n_9669 = ~n_9665 &  n_9668;
assign n_9670 =  x_2940 & ~n_9669;
assign n_9671 = ~x_2940 &  n_9669;
assign n_9672 = ~n_9670 & ~n_9671;
assign n_9673 =  x_2939 & ~n_9432;
assign n_9674 =  x_3225 &  n_9429;
assign n_9675 =  x_4457 &  n_558;
assign n_9676 = ~n_9674 & ~n_9675;
assign n_9677 = ~n_9673 &  n_9676;
assign n_9678 =  x_2939 & ~n_9677;
assign n_9679 = ~x_2939 &  n_9677;
assign n_9680 = ~n_9678 & ~n_9679;
assign n_9681 =  x_2938 & ~n_9432;
assign n_9682 =  x_3224 &  n_9429;
assign n_9683 =  x_4456 &  n_558;
assign n_9684 = ~n_9682 & ~n_9683;
assign n_9685 = ~n_9681 &  n_9684;
assign n_9686 =  x_2938 & ~n_9685;
assign n_9687 = ~x_2938 &  n_9685;
assign n_9688 = ~n_9686 & ~n_9687;
assign n_9689 =  x_42 &  n_766;
assign n_9690 =  x_43 &  n_9689;
assign n_9691 =  n_9690 &  n_1900;
assign n_9692 =  x_2874 & ~n_9691;
assign n_9693 =  x_1834 &  n_9691;
assign n_9694 = ~n_9692 & ~n_9693;
assign n_9695 =  x_2874 & ~n_9694;
assign n_9696 = ~x_2874 &  n_9694;
assign n_9697 = ~n_9695 & ~n_9696;
assign n_9698 =  x_2873 & ~n_9691;
assign n_9699 =  x_1833 &  n_9691;
assign n_9700 = ~n_9698 & ~n_9699;
assign n_9701 =  x_2873 & ~n_9700;
assign n_9702 = ~x_2873 &  n_9700;
assign n_9703 = ~n_9701 & ~n_9702;
assign n_9704 =  x_2872 & ~n_9691;
assign n_9705 =  x_1832 &  n_9691;
assign n_9706 = ~n_9704 & ~n_9705;
assign n_9707 =  x_2872 & ~n_9706;
assign n_9708 = ~x_2872 &  n_9706;
assign n_9709 = ~n_9707 & ~n_9708;
assign n_9710 =  x_2871 & ~n_9691;
assign n_9711 =  x_1831 &  n_9691;
assign n_9712 = ~n_9710 & ~n_9711;
assign n_9713 =  x_2871 & ~n_9712;
assign n_9714 = ~x_2871 &  n_9712;
assign n_9715 = ~n_9713 & ~n_9714;
assign n_9716 =  x_2870 & ~n_9691;
assign n_9717 =  x_1830 &  n_9691;
assign n_9718 = ~n_9716 & ~n_9717;
assign n_9719 =  x_2870 & ~n_9718;
assign n_9720 = ~x_2870 &  n_9718;
assign n_9721 = ~n_9719 & ~n_9720;
assign n_9722 =  x_2869 & ~n_9691;
assign n_9723 =  x_1829 &  n_9691;
assign n_9724 = ~n_9722 & ~n_9723;
assign n_9725 =  x_2869 & ~n_9724;
assign n_9726 = ~x_2869 &  n_9724;
assign n_9727 = ~n_9725 & ~n_9726;
assign n_9728 =  x_2868 & ~n_9691;
assign n_9729 =  x_1828 &  n_9691;
assign n_9730 = ~n_9728 & ~n_9729;
assign n_9731 =  x_2868 & ~n_9730;
assign n_9732 = ~x_2868 &  n_9730;
assign n_9733 = ~n_9731 & ~n_9732;
assign n_9734 =  x_2867 & ~n_9691;
assign n_9735 =  x_1827 &  n_9691;
assign n_9736 = ~n_9734 & ~n_9735;
assign n_9737 =  x_2867 & ~n_9736;
assign n_9738 = ~x_2867 &  n_9736;
assign n_9739 = ~n_9737 & ~n_9738;
assign n_9740 =  x_2866 & ~n_9691;
assign n_9741 =  x_1826 &  n_9691;
assign n_9742 = ~n_9740 & ~n_9741;
assign n_9743 =  x_2866 & ~n_9742;
assign n_9744 = ~x_2866 &  n_9742;
assign n_9745 = ~n_9743 & ~n_9744;
assign n_9746 =  x_2865 & ~n_9691;
assign n_9747 =  x_1825 &  n_9691;
assign n_9748 = ~n_9746 & ~n_9747;
assign n_9749 =  x_2865 & ~n_9748;
assign n_9750 = ~x_2865 &  n_9748;
assign n_9751 = ~n_9749 & ~n_9750;
assign n_9752 =  x_2864 & ~n_9691;
assign n_9753 =  x_1824 &  n_9691;
assign n_9754 = ~n_9752 & ~n_9753;
assign n_9755 =  x_2864 & ~n_9754;
assign n_9756 = ~x_2864 &  n_9754;
assign n_9757 = ~n_9755 & ~n_9756;
assign n_9758 =  x_2863 & ~n_9691;
assign n_9759 =  x_1823 &  n_9691;
assign n_9760 = ~n_9758 & ~n_9759;
assign n_9761 =  x_2863 & ~n_9760;
assign n_9762 = ~x_2863 &  n_9760;
assign n_9763 = ~n_9761 & ~n_9762;
assign n_9764 =  x_2862 & ~n_9691;
assign n_9765 =  x_1822 &  n_9691;
assign n_9766 = ~n_9764 & ~n_9765;
assign n_9767 =  x_2862 & ~n_9766;
assign n_9768 = ~x_2862 &  n_9766;
assign n_9769 = ~n_9767 & ~n_9768;
assign n_9770 =  x_2861 & ~n_9691;
assign n_9771 =  x_1821 &  n_9691;
assign n_9772 = ~n_9770 & ~n_9771;
assign n_9773 =  x_2861 & ~n_9772;
assign n_9774 = ~x_2861 &  n_9772;
assign n_9775 = ~n_9773 & ~n_9774;
assign n_9776 =  x_2860 & ~n_9691;
assign n_9777 =  x_1820 &  n_9691;
assign n_9778 = ~n_9776 & ~n_9777;
assign n_9779 =  x_2860 & ~n_9778;
assign n_9780 = ~x_2860 &  n_9778;
assign n_9781 = ~n_9779 & ~n_9780;
assign n_9782 =  x_2859 & ~n_9691;
assign n_9783 =  x_1819 &  n_9691;
assign n_9784 = ~n_9782 & ~n_9783;
assign n_9785 =  x_2859 & ~n_9784;
assign n_9786 = ~x_2859 &  n_9784;
assign n_9787 = ~n_9785 & ~n_9786;
assign n_9788 =  x_2858 & ~n_9691;
assign n_9789 =  x_1818 &  n_9691;
assign n_9790 = ~n_9788 & ~n_9789;
assign n_9791 =  x_2858 & ~n_9790;
assign n_9792 = ~x_2858 &  n_9790;
assign n_9793 = ~n_9791 & ~n_9792;
assign n_9794 =  x_2857 & ~n_9691;
assign n_9795 =  x_1817 &  n_9691;
assign n_9796 = ~n_9794 & ~n_9795;
assign n_9797 =  x_2857 & ~n_9796;
assign n_9798 = ~x_2857 &  n_9796;
assign n_9799 = ~n_9797 & ~n_9798;
assign n_9800 =  x_2856 & ~n_9691;
assign n_9801 =  x_1816 &  n_9691;
assign n_9802 = ~n_9800 & ~n_9801;
assign n_9803 =  x_2856 & ~n_9802;
assign n_9804 = ~x_2856 &  n_9802;
assign n_9805 = ~n_9803 & ~n_9804;
assign n_9806 =  x_2855 & ~n_9691;
assign n_9807 =  x_1815 &  n_9691;
assign n_9808 = ~n_9806 & ~n_9807;
assign n_9809 =  x_2855 & ~n_9808;
assign n_9810 = ~x_2855 &  n_9808;
assign n_9811 = ~n_9809 & ~n_9810;
assign n_9812 =  x_2854 & ~n_9691;
assign n_9813 =  x_1814 &  n_9691;
assign n_9814 = ~n_9812 & ~n_9813;
assign n_9815 =  x_2854 & ~n_9814;
assign n_9816 = ~x_2854 &  n_9814;
assign n_9817 = ~n_9815 & ~n_9816;
assign n_9818 =  x_2853 & ~n_9691;
assign n_9819 =  x_1813 &  n_9691;
assign n_9820 = ~n_9818 & ~n_9819;
assign n_9821 =  x_2853 & ~n_9820;
assign n_9822 = ~x_2853 &  n_9820;
assign n_9823 = ~n_9821 & ~n_9822;
assign n_9824 =  x_2852 & ~n_9691;
assign n_9825 =  x_1812 &  n_9691;
assign n_9826 = ~n_9824 & ~n_9825;
assign n_9827 =  x_2852 & ~n_9826;
assign n_9828 = ~x_2852 &  n_9826;
assign n_9829 = ~n_9827 & ~n_9828;
assign n_9830 =  x_2851 & ~n_9691;
assign n_9831 =  x_1811 &  n_9691;
assign n_9832 = ~n_9830 & ~n_9831;
assign n_9833 =  x_2851 & ~n_9832;
assign n_9834 = ~x_2851 &  n_9832;
assign n_9835 = ~n_9833 & ~n_9834;
assign n_9836 =  x_2850 & ~n_9691;
assign n_9837 =  x_1810 &  n_9691;
assign n_9838 = ~n_9836 & ~n_9837;
assign n_9839 =  x_2850 & ~n_9838;
assign n_9840 = ~x_2850 &  n_9838;
assign n_9841 = ~n_9839 & ~n_9840;
assign n_9842 =  x_2849 & ~n_9691;
assign n_9843 =  x_1809 &  n_9691;
assign n_9844 = ~n_9842 & ~n_9843;
assign n_9845 =  x_2849 & ~n_9844;
assign n_9846 = ~x_2849 &  n_9844;
assign n_9847 = ~n_9845 & ~n_9846;
assign n_9848 =  x_2848 & ~n_9691;
assign n_9849 =  x_1808 &  n_9691;
assign n_9850 = ~n_9848 & ~n_9849;
assign n_9851 =  x_2848 & ~n_9850;
assign n_9852 = ~x_2848 &  n_9850;
assign n_9853 = ~n_9851 & ~n_9852;
assign n_9854 =  x_2847 & ~n_9691;
assign n_9855 =  x_1807 &  n_9691;
assign n_9856 = ~n_9854 & ~n_9855;
assign n_9857 =  x_2847 & ~n_9856;
assign n_9858 = ~x_2847 &  n_9856;
assign n_9859 = ~n_9857 & ~n_9858;
assign n_9860 =  x_2846 & ~n_9691;
assign n_9861 =  x_1806 &  n_9691;
assign n_9862 = ~n_9860 & ~n_9861;
assign n_9863 =  x_2846 & ~n_9862;
assign n_9864 = ~x_2846 &  n_9862;
assign n_9865 = ~n_9863 & ~n_9864;
assign n_9866 =  x_2845 & ~n_9691;
assign n_9867 =  x_1805 &  n_9691;
assign n_9868 = ~n_9866 & ~n_9867;
assign n_9869 =  x_2845 & ~n_9868;
assign n_9870 = ~x_2845 &  n_9868;
assign n_9871 = ~n_9869 & ~n_9870;
assign n_9872 =  x_2844 & ~n_9691;
assign n_9873 =  x_1804 &  n_9691;
assign n_9874 = ~n_9872 & ~n_9873;
assign n_9875 =  x_2844 & ~n_9874;
assign n_9876 = ~x_2844 &  n_9874;
assign n_9877 = ~n_9875 & ~n_9876;
assign n_9878 =  x_2843 & ~n_9691;
assign n_9879 =  x_1803 &  n_9691;
assign n_9880 = ~n_9878 & ~n_9879;
assign n_9881 =  x_2843 & ~n_9880;
assign n_9882 = ~x_2843 &  n_9880;
assign n_9883 = ~n_9881 & ~n_9882;
assign n_9884 =  n_12 &  n_11;
assign n_9885 =  n_9884 &  n_357;
assign n_9886 =  x_2810 & ~n_9885;
assign n_9887 =  i_32 &  n_9885;
assign n_9888 = ~n_9886 & ~n_9887;
assign n_9889 =  x_2810 & ~n_9888;
assign n_9890 = ~x_2810 &  n_9888;
assign n_9891 = ~n_9889 & ~n_9890;
assign n_9892 =  x_2809 & ~n_9885;
assign n_9893 =  i_31 &  n_9885;
assign n_9894 = ~n_9892 & ~n_9893;
assign n_9895 =  x_2809 & ~n_9894;
assign n_9896 = ~x_2809 &  n_9894;
assign n_9897 = ~n_9895 & ~n_9896;
assign n_9898 =  x_2808 & ~n_9885;
assign n_9899 =  i_30 &  n_9885;
assign n_9900 = ~n_9898 & ~n_9899;
assign n_9901 =  x_2808 & ~n_9900;
assign n_9902 = ~x_2808 &  n_9900;
assign n_9903 = ~n_9901 & ~n_9902;
assign n_9904 =  x_2807 & ~n_9885;
assign n_9905 =  i_29 &  n_9885;
assign n_9906 = ~n_9904 & ~n_9905;
assign n_9907 =  x_2807 & ~n_9906;
assign n_9908 = ~x_2807 &  n_9906;
assign n_9909 = ~n_9907 & ~n_9908;
assign n_9910 =  x_2806 & ~n_9885;
assign n_9911 =  i_28 &  n_9885;
assign n_9912 = ~n_9910 & ~n_9911;
assign n_9913 =  x_2806 & ~n_9912;
assign n_9914 = ~x_2806 &  n_9912;
assign n_9915 = ~n_9913 & ~n_9914;
assign n_9916 =  x_2805 & ~n_9885;
assign n_9917 =  i_27 &  n_9885;
assign n_9918 = ~n_9916 & ~n_9917;
assign n_9919 =  x_2805 & ~n_9918;
assign n_9920 = ~x_2805 &  n_9918;
assign n_9921 = ~n_9919 & ~n_9920;
assign n_9922 =  x_2804 & ~n_9885;
assign n_9923 =  i_26 &  n_9885;
assign n_9924 = ~n_9922 & ~n_9923;
assign n_9925 =  x_2804 & ~n_9924;
assign n_9926 = ~x_2804 &  n_9924;
assign n_9927 = ~n_9925 & ~n_9926;
assign n_9928 =  x_2803 & ~n_9885;
assign n_9929 =  i_25 &  n_9885;
assign n_9930 = ~n_9928 & ~n_9929;
assign n_9931 =  x_2803 & ~n_9930;
assign n_9932 = ~x_2803 &  n_9930;
assign n_9933 = ~n_9931 & ~n_9932;
assign n_9934 =  x_2802 & ~n_9885;
assign n_9935 =  i_24 &  n_9885;
assign n_9936 = ~n_9934 & ~n_9935;
assign n_9937 =  x_2802 & ~n_9936;
assign n_9938 = ~x_2802 &  n_9936;
assign n_9939 = ~n_9937 & ~n_9938;
assign n_9940 =  x_2801 & ~n_9885;
assign n_9941 =  i_23 &  n_9885;
assign n_9942 = ~n_9940 & ~n_9941;
assign n_9943 =  x_2801 & ~n_9942;
assign n_9944 = ~x_2801 &  n_9942;
assign n_9945 = ~n_9943 & ~n_9944;
assign n_9946 =  x_2800 & ~n_9885;
assign n_9947 =  i_22 &  n_9885;
assign n_9948 = ~n_9946 & ~n_9947;
assign n_9949 =  x_2800 & ~n_9948;
assign n_9950 = ~x_2800 &  n_9948;
assign n_9951 = ~n_9949 & ~n_9950;
assign n_9952 =  x_2799 & ~n_9885;
assign n_9953 =  i_21 &  n_9885;
assign n_9954 = ~n_9952 & ~n_9953;
assign n_9955 =  x_2799 & ~n_9954;
assign n_9956 = ~x_2799 &  n_9954;
assign n_9957 = ~n_9955 & ~n_9956;
assign n_9958 =  x_2798 & ~n_9885;
assign n_9959 =  i_20 &  n_9885;
assign n_9960 = ~n_9958 & ~n_9959;
assign n_9961 =  x_2798 & ~n_9960;
assign n_9962 = ~x_2798 &  n_9960;
assign n_9963 = ~n_9961 & ~n_9962;
assign n_9964 =  x_2797 & ~n_9885;
assign n_9965 =  i_19 &  n_9885;
assign n_9966 = ~n_9964 & ~n_9965;
assign n_9967 =  x_2797 & ~n_9966;
assign n_9968 = ~x_2797 &  n_9966;
assign n_9969 = ~n_9967 & ~n_9968;
assign n_9970 =  x_2796 & ~n_9885;
assign n_9971 =  i_18 &  n_9885;
assign n_9972 = ~n_9970 & ~n_9971;
assign n_9973 =  x_2796 & ~n_9972;
assign n_9974 = ~x_2796 &  n_9972;
assign n_9975 = ~n_9973 & ~n_9974;
assign n_9976 =  x_2795 & ~n_9885;
assign n_9977 =  i_17 &  n_9885;
assign n_9978 = ~n_9976 & ~n_9977;
assign n_9979 =  x_2795 & ~n_9978;
assign n_9980 = ~x_2795 &  n_9978;
assign n_9981 = ~n_9979 & ~n_9980;
assign n_9982 =  x_2794 & ~n_9885;
assign n_9983 =  i_16 &  n_9885;
assign n_9984 = ~n_9982 & ~n_9983;
assign n_9985 =  x_2794 & ~n_9984;
assign n_9986 = ~x_2794 &  n_9984;
assign n_9987 = ~n_9985 & ~n_9986;
assign n_9988 =  x_2793 & ~n_9885;
assign n_9989 =  i_15 &  n_9885;
assign n_9990 = ~n_9988 & ~n_9989;
assign n_9991 =  x_2793 & ~n_9990;
assign n_9992 = ~x_2793 &  n_9990;
assign n_9993 = ~n_9991 & ~n_9992;
assign n_9994 =  x_2792 & ~n_9885;
assign n_9995 =  i_14 &  n_9885;
assign n_9996 = ~n_9994 & ~n_9995;
assign n_9997 =  x_2792 & ~n_9996;
assign n_9998 = ~x_2792 &  n_9996;
assign n_9999 = ~n_9997 & ~n_9998;
assign n_10000 =  x_2791 & ~n_9885;
assign n_10001 =  i_13 &  n_9885;
assign n_10002 = ~n_10000 & ~n_10001;
assign n_10003 =  x_2791 & ~n_10002;
assign n_10004 = ~x_2791 &  n_10002;
assign n_10005 = ~n_10003 & ~n_10004;
assign n_10006 =  x_2790 & ~n_9885;
assign n_10007 =  i_12 &  n_9885;
assign n_10008 = ~n_10006 & ~n_10007;
assign n_10009 =  x_2790 & ~n_10008;
assign n_10010 = ~x_2790 &  n_10008;
assign n_10011 = ~n_10009 & ~n_10010;
assign n_10012 =  x_2789 & ~n_9885;
assign n_10013 =  i_11 &  n_9885;
assign n_10014 = ~n_10012 & ~n_10013;
assign n_10015 =  x_2789 & ~n_10014;
assign n_10016 = ~x_2789 &  n_10014;
assign n_10017 = ~n_10015 & ~n_10016;
assign n_10018 =  x_2788 & ~n_9885;
assign n_10019 =  i_10 &  n_9885;
assign n_10020 = ~n_10018 & ~n_10019;
assign n_10021 =  x_2788 & ~n_10020;
assign n_10022 = ~x_2788 &  n_10020;
assign n_10023 = ~n_10021 & ~n_10022;
assign n_10024 =  x_2787 & ~n_9885;
assign n_10025 =  i_9 &  n_9885;
assign n_10026 = ~n_10024 & ~n_10025;
assign n_10027 =  x_2787 & ~n_10026;
assign n_10028 = ~x_2787 &  n_10026;
assign n_10029 = ~n_10027 & ~n_10028;
assign n_10030 =  x_2786 & ~n_9885;
assign n_10031 =  i_8 &  n_9885;
assign n_10032 = ~n_10030 & ~n_10031;
assign n_10033 =  x_2786 & ~n_10032;
assign n_10034 = ~x_2786 &  n_10032;
assign n_10035 = ~n_10033 & ~n_10034;
assign n_10036 =  x_2785 & ~n_9885;
assign n_10037 =  i_7 &  n_9885;
assign n_10038 = ~n_10036 & ~n_10037;
assign n_10039 =  x_2785 & ~n_10038;
assign n_10040 = ~x_2785 &  n_10038;
assign n_10041 = ~n_10039 & ~n_10040;
assign n_10042 =  x_2784 & ~n_9885;
assign n_10043 =  i_6 &  n_9885;
assign n_10044 = ~n_10042 & ~n_10043;
assign n_10045 =  x_2784 & ~n_10044;
assign n_10046 = ~x_2784 &  n_10044;
assign n_10047 = ~n_10045 & ~n_10046;
assign n_10048 =  x_2783 & ~n_9885;
assign n_10049 =  i_5 &  n_9885;
assign n_10050 = ~n_10048 & ~n_10049;
assign n_10051 =  x_2783 & ~n_10050;
assign n_10052 = ~x_2783 &  n_10050;
assign n_10053 = ~n_10051 & ~n_10052;
assign n_10054 =  x_2782 & ~n_9885;
assign n_10055 =  i_4 &  n_9885;
assign n_10056 = ~n_10054 & ~n_10055;
assign n_10057 =  x_2782 & ~n_10056;
assign n_10058 = ~x_2782 &  n_10056;
assign n_10059 = ~n_10057 & ~n_10058;
assign n_10060 =  x_2781 & ~n_9885;
assign n_10061 =  i_3 &  n_9885;
assign n_10062 = ~n_10060 & ~n_10061;
assign n_10063 =  x_2781 & ~n_10062;
assign n_10064 = ~x_2781 &  n_10062;
assign n_10065 = ~n_10063 & ~n_10064;
assign n_10066 =  x_2780 & ~n_9885;
assign n_10067 =  i_2 &  n_9885;
assign n_10068 = ~n_10066 & ~n_10067;
assign n_10069 =  x_2780 & ~n_10068;
assign n_10070 = ~x_2780 &  n_10068;
assign n_10071 = ~n_10069 & ~n_10070;
assign n_10072 =  x_2779 & ~n_9885;
assign n_10073 =  i_1 &  n_9885;
assign n_10074 = ~n_10072 & ~n_10073;
assign n_10075 =  x_2779 & ~n_10074;
assign n_10076 = ~x_2779 &  n_10074;
assign n_10077 = ~n_10075 & ~n_10076;
assign n_10078 =  n_7 &  n_1305;
assign n_10079 =  n_5654 &  n_551;
assign n_10080 = ~x_41 &  n_10079;
assign n_10081 =  n_10078 &  n_10080;
assign n_10082 =  x_2778 & ~n_10081;
assign n_10083 =  i_32 &  n_10081;
assign n_10084 = ~n_10082 & ~n_10083;
assign n_10085 =  x_2778 & ~n_10084;
assign n_10086 = ~x_2778 &  n_10084;
assign n_10087 = ~n_10085 & ~n_10086;
assign n_10088 =  x_2777 & ~n_10081;
assign n_10089 =  i_31 &  n_10081;
assign n_10090 = ~n_10088 & ~n_10089;
assign n_10091 =  x_2777 & ~n_10090;
assign n_10092 = ~x_2777 &  n_10090;
assign n_10093 = ~n_10091 & ~n_10092;
assign n_10094 =  x_2776 & ~n_10081;
assign n_10095 =  i_30 &  n_10081;
assign n_10096 = ~n_10094 & ~n_10095;
assign n_10097 =  x_2776 & ~n_10096;
assign n_10098 = ~x_2776 &  n_10096;
assign n_10099 = ~n_10097 & ~n_10098;
assign n_10100 =  x_2775 & ~n_10081;
assign n_10101 =  i_29 &  n_10081;
assign n_10102 = ~n_10100 & ~n_10101;
assign n_10103 =  x_2775 & ~n_10102;
assign n_10104 = ~x_2775 &  n_10102;
assign n_10105 = ~n_10103 & ~n_10104;
assign n_10106 =  x_2774 & ~n_10081;
assign n_10107 =  i_28 &  n_10081;
assign n_10108 = ~n_10106 & ~n_10107;
assign n_10109 =  x_2774 & ~n_10108;
assign n_10110 = ~x_2774 &  n_10108;
assign n_10111 = ~n_10109 & ~n_10110;
assign n_10112 =  x_2773 & ~n_10081;
assign n_10113 =  i_27 &  n_10081;
assign n_10114 = ~n_10112 & ~n_10113;
assign n_10115 =  x_2773 & ~n_10114;
assign n_10116 = ~x_2773 &  n_10114;
assign n_10117 = ~n_10115 & ~n_10116;
assign n_10118 =  x_2772 & ~n_10081;
assign n_10119 =  i_26 &  n_10081;
assign n_10120 = ~n_10118 & ~n_10119;
assign n_10121 =  x_2772 & ~n_10120;
assign n_10122 = ~x_2772 &  n_10120;
assign n_10123 = ~n_10121 & ~n_10122;
assign n_10124 =  x_2771 & ~n_10081;
assign n_10125 =  i_25 &  n_10081;
assign n_10126 = ~n_10124 & ~n_10125;
assign n_10127 =  x_2771 & ~n_10126;
assign n_10128 = ~x_2771 &  n_10126;
assign n_10129 = ~n_10127 & ~n_10128;
assign n_10130 =  x_2770 & ~n_10081;
assign n_10131 =  i_24 &  n_10081;
assign n_10132 = ~n_10130 & ~n_10131;
assign n_10133 =  x_2770 & ~n_10132;
assign n_10134 = ~x_2770 &  n_10132;
assign n_10135 = ~n_10133 & ~n_10134;
assign n_10136 =  x_2769 & ~n_10081;
assign n_10137 =  i_23 &  n_10081;
assign n_10138 = ~n_10136 & ~n_10137;
assign n_10139 =  x_2769 & ~n_10138;
assign n_10140 = ~x_2769 &  n_10138;
assign n_10141 = ~n_10139 & ~n_10140;
assign n_10142 =  x_2768 & ~n_10081;
assign n_10143 =  i_22 &  n_10081;
assign n_10144 = ~n_10142 & ~n_10143;
assign n_10145 =  x_2768 & ~n_10144;
assign n_10146 = ~x_2768 &  n_10144;
assign n_10147 = ~n_10145 & ~n_10146;
assign n_10148 =  x_2767 & ~n_10081;
assign n_10149 =  i_21 &  n_10081;
assign n_10150 = ~n_10148 & ~n_10149;
assign n_10151 =  x_2767 & ~n_10150;
assign n_10152 = ~x_2767 &  n_10150;
assign n_10153 = ~n_10151 & ~n_10152;
assign n_10154 =  x_2766 & ~n_10081;
assign n_10155 =  i_20 &  n_10081;
assign n_10156 = ~n_10154 & ~n_10155;
assign n_10157 =  x_2766 & ~n_10156;
assign n_10158 = ~x_2766 &  n_10156;
assign n_10159 = ~n_10157 & ~n_10158;
assign n_10160 =  x_2765 & ~n_10081;
assign n_10161 =  i_19 &  n_10081;
assign n_10162 = ~n_10160 & ~n_10161;
assign n_10163 =  x_2765 & ~n_10162;
assign n_10164 = ~x_2765 &  n_10162;
assign n_10165 = ~n_10163 & ~n_10164;
assign n_10166 =  x_2764 & ~n_10081;
assign n_10167 =  i_18 &  n_10081;
assign n_10168 = ~n_10166 & ~n_10167;
assign n_10169 =  x_2764 & ~n_10168;
assign n_10170 = ~x_2764 &  n_10168;
assign n_10171 = ~n_10169 & ~n_10170;
assign n_10172 =  x_2763 & ~n_10081;
assign n_10173 =  i_17 &  n_10081;
assign n_10174 = ~n_10172 & ~n_10173;
assign n_10175 =  x_2763 & ~n_10174;
assign n_10176 = ~x_2763 &  n_10174;
assign n_10177 = ~n_10175 & ~n_10176;
assign n_10178 =  x_2762 & ~n_10081;
assign n_10179 =  i_16 &  n_10081;
assign n_10180 = ~n_10178 & ~n_10179;
assign n_10181 =  x_2762 & ~n_10180;
assign n_10182 = ~x_2762 &  n_10180;
assign n_10183 = ~n_10181 & ~n_10182;
assign n_10184 =  x_2761 & ~n_10081;
assign n_10185 =  i_15 &  n_10081;
assign n_10186 = ~n_10184 & ~n_10185;
assign n_10187 =  x_2761 & ~n_10186;
assign n_10188 = ~x_2761 &  n_10186;
assign n_10189 = ~n_10187 & ~n_10188;
assign n_10190 =  x_2760 & ~n_10081;
assign n_10191 =  i_14 &  n_10081;
assign n_10192 = ~n_10190 & ~n_10191;
assign n_10193 =  x_2760 & ~n_10192;
assign n_10194 = ~x_2760 &  n_10192;
assign n_10195 = ~n_10193 & ~n_10194;
assign n_10196 =  x_2759 & ~n_10081;
assign n_10197 =  i_13 &  n_10081;
assign n_10198 = ~n_10196 & ~n_10197;
assign n_10199 =  x_2759 & ~n_10198;
assign n_10200 = ~x_2759 &  n_10198;
assign n_10201 = ~n_10199 & ~n_10200;
assign n_10202 =  x_2758 & ~n_10081;
assign n_10203 =  i_12 &  n_10081;
assign n_10204 = ~n_10202 & ~n_10203;
assign n_10205 =  x_2758 & ~n_10204;
assign n_10206 = ~x_2758 &  n_10204;
assign n_10207 = ~n_10205 & ~n_10206;
assign n_10208 =  x_2757 & ~n_10081;
assign n_10209 =  i_11 &  n_10081;
assign n_10210 = ~n_10208 & ~n_10209;
assign n_10211 =  x_2757 & ~n_10210;
assign n_10212 = ~x_2757 &  n_10210;
assign n_10213 = ~n_10211 & ~n_10212;
assign n_10214 =  x_2756 & ~n_10081;
assign n_10215 =  i_10 &  n_10081;
assign n_10216 = ~n_10214 & ~n_10215;
assign n_10217 =  x_2756 & ~n_10216;
assign n_10218 = ~x_2756 &  n_10216;
assign n_10219 = ~n_10217 & ~n_10218;
assign n_10220 =  x_2755 & ~n_10081;
assign n_10221 =  i_9 &  n_10081;
assign n_10222 = ~n_10220 & ~n_10221;
assign n_10223 =  x_2755 & ~n_10222;
assign n_10224 = ~x_2755 &  n_10222;
assign n_10225 = ~n_10223 & ~n_10224;
assign n_10226 =  x_2754 & ~n_10081;
assign n_10227 =  i_8 &  n_10081;
assign n_10228 = ~n_10226 & ~n_10227;
assign n_10229 =  x_2754 & ~n_10228;
assign n_10230 = ~x_2754 &  n_10228;
assign n_10231 = ~n_10229 & ~n_10230;
assign n_10232 =  x_2753 & ~n_10081;
assign n_10233 =  i_7 &  n_10081;
assign n_10234 = ~n_10232 & ~n_10233;
assign n_10235 =  x_2753 & ~n_10234;
assign n_10236 = ~x_2753 &  n_10234;
assign n_10237 = ~n_10235 & ~n_10236;
assign n_10238 =  x_2752 & ~n_10081;
assign n_10239 =  i_6 &  n_10081;
assign n_10240 = ~n_10238 & ~n_10239;
assign n_10241 =  x_2752 & ~n_10240;
assign n_10242 = ~x_2752 &  n_10240;
assign n_10243 = ~n_10241 & ~n_10242;
assign n_10244 =  x_2751 & ~n_10081;
assign n_10245 =  i_5 &  n_10081;
assign n_10246 = ~n_10244 & ~n_10245;
assign n_10247 =  x_2751 & ~n_10246;
assign n_10248 = ~x_2751 &  n_10246;
assign n_10249 = ~n_10247 & ~n_10248;
assign n_10250 =  x_2750 & ~n_10081;
assign n_10251 =  i_4 &  n_10081;
assign n_10252 = ~n_10250 & ~n_10251;
assign n_10253 =  x_2750 & ~n_10252;
assign n_10254 = ~x_2750 &  n_10252;
assign n_10255 = ~n_10253 & ~n_10254;
assign n_10256 =  x_2749 & ~n_10081;
assign n_10257 =  i_3 &  n_10081;
assign n_10258 = ~n_10256 & ~n_10257;
assign n_10259 =  x_2749 & ~n_10258;
assign n_10260 = ~x_2749 &  n_10258;
assign n_10261 = ~n_10259 & ~n_10260;
assign n_10262 =  x_2748 & ~n_10081;
assign n_10263 =  i_2 &  n_10081;
assign n_10264 = ~n_10262 & ~n_10263;
assign n_10265 =  x_2748 & ~n_10264;
assign n_10266 = ~x_2748 &  n_10264;
assign n_10267 = ~n_10265 & ~n_10266;
assign n_10268 =  x_2747 & ~n_10081;
assign n_10269 =  i_1 &  n_10081;
assign n_10270 = ~n_10268 & ~n_10269;
assign n_10271 =  x_2747 & ~n_10270;
assign n_10272 = ~x_2747 &  n_10270;
assign n_10273 = ~n_10271 & ~n_10272;
assign n_10274 =  x_41 &  n_1305;
assign n_10275 =  n_349 &  n_10274;
assign n_10276 =  n_7 &  n_551;
assign n_10277 =  n_10275 &  n_10276;
assign n_10278 =  x_2746 & ~n_10277;
assign n_10279 =  i_32 &  n_10277;
assign n_10280 = ~n_10278 & ~n_10279;
assign n_10281 =  x_2746 & ~n_10280;
assign n_10282 = ~x_2746 &  n_10280;
assign n_10283 = ~n_10281 & ~n_10282;
assign n_10284 =  x_2745 & ~n_10277;
assign n_10285 =  i_31 &  n_10277;
assign n_10286 = ~n_10284 & ~n_10285;
assign n_10287 =  x_2745 & ~n_10286;
assign n_10288 = ~x_2745 &  n_10286;
assign n_10289 = ~n_10287 & ~n_10288;
assign n_10290 =  x_2744 & ~n_10277;
assign n_10291 =  i_30 &  n_10277;
assign n_10292 = ~n_10290 & ~n_10291;
assign n_10293 =  x_2744 & ~n_10292;
assign n_10294 = ~x_2744 &  n_10292;
assign n_10295 = ~n_10293 & ~n_10294;
assign n_10296 =  x_2743 & ~n_10277;
assign n_10297 =  i_29 &  n_10277;
assign n_10298 = ~n_10296 & ~n_10297;
assign n_10299 =  x_2743 & ~n_10298;
assign n_10300 = ~x_2743 &  n_10298;
assign n_10301 = ~n_10299 & ~n_10300;
assign n_10302 =  x_2742 & ~n_10277;
assign n_10303 =  i_28 &  n_10277;
assign n_10304 = ~n_10302 & ~n_10303;
assign n_10305 =  x_2742 & ~n_10304;
assign n_10306 = ~x_2742 &  n_10304;
assign n_10307 = ~n_10305 & ~n_10306;
assign n_10308 =  x_2741 & ~n_10277;
assign n_10309 =  i_27 &  n_10277;
assign n_10310 = ~n_10308 & ~n_10309;
assign n_10311 =  x_2741 & ~n_10310;
assign n_10312 = ~x_2741 &  n_10310;
assign n_10313 = ~n_10311 & ~n_10312;
assign n_10314 =  x_2740 & ~n_10277;
assign n_10315 =  i_26 &  n_10277;
assign n_10316 = ~n_10314 & ~n_10315;
assign n_10317 =  x_2740 & ~n_10316;
assign n_10318 = ~x_2740 &  n_10316;
assign n_10319 = ~n_10317 & ~n_10318;
assign n_10320 =  x_2739 & ~n_10277;
assign n_10321 =  i_25 &  n_10277;
assign n_10322 = ~n_10320 & ~n_10321;
assign n_10323 =  x_2739 & ~n_10322;
assign n_10324 = ~x_2739 &  n_10322;
assign n_10325 = ~n_10323 & ~n_10324;
assign n_10326 =  x_2738 & ~n_10277;
assign n_10327 =  i_24 &  n_10277;
assign n_10328 = ~n_10326 & ~n_10327;
assign n_10329 =  x_2738 & ~n_10328;
assign n_10330 = ~x_2738 &  n_10328;
assign n_10331 = ~n_10329 & ~n_10330;
assign n_10332 =  x_2737 & ~n_10277;
assign n_10333 =  i_23 &  n_10277;
assign n_10334 = ~n_10332 & ~n_10333;
assign n_10335 =  x_2737 & ~n_10334;
assign n_10336 = ~x_2737 &  n_10334;
assign n_10337 = ~n_10335 & ~n_10336;
assign n_10338 =  x_2736 & ~n_10277;
assign n_10339 =  i_22 &  n_10277;
assign n_10340 = ~n_10338 & ~n_10339;
assign n_10341 =  x_2736 & ~n_10340;
assign n_10342 = ~x_2736 &  n_10340;
assign n_10343 = ~n_10341 & ~n_10342;
assign n_10344 =  x_2735 & ~n_10277;
assign n_10345 =  i_21 &  n_10277;
assign n_10346 = ~n_10344 & ~n_10345;
assign n_10347 =  x_2735 & ~n_10346;
assign n_10348 = ~x_2735 &  n_10346;
assign n_10349 = ~n_10347 & ~n_10348;
assign n_10350 =  x_2734 & ~n_10277;
assign n_10351 =  i_20 &  n_10277;
assign n_10352 = ~n_10350 & ~n_10351;
assign n_10353 =  x_2734 & ~n_10352;
assign n_10354 = ~x_2734 &  n_10352;
assign n_10355 = ~n_10353 & ~n_10354;
assign n_10356 =  x_2733 & ~n_10277;
assign n_10357 =  i_19 &  n_10277;
assign n_10358 = ~n_10356 & ~n_10357;
assign n_10359 =  x_2733 & ~n_10358;
assign n_10360 = ~x_2733 &  n_10358;
assign n_10361 = ~n_10359 & ~n_10360;
assign n_10362 =  x_2732 & ~n_10277;
assign n_10363 =  i_18 &  n_10277;
assign n_10364 = ~n_10362 & ~n_10363;
assign n_10365 =  x_2732 & ~n_10364;
assign n_10366 = ~x_2732 &  n_10364;
assign n_10367 = ~n_10365 & ~n_10366;
assign n_10368 =  x_2731 & ~n_10277;
assign n_10369 =  i_17 &  n_10277;
assign n_10370 = ~n_10368 & ~n_10369;
assign n_10371 =  x_2731 & ~n_10370;
assign n_10372 = ~x_2731 &  n_10370;
assign n_10373 = ~n_10371 & ~n_10372;
assign n_10374 =  x_2730 & ~n_10277;
assign n_10375 =  i_16 &  n_10277;
assign n_10376 = ~n_10374 & ~n_10375;
assign n_10377 =  x_2730 & ~n_10376;
assign n_10378 = ~x_2730 &  n_10376;
assign n_10379 = ~n_10377 & ~n_10378;
assign n_10380 =  x_2729 & ~n_10277;
assign n_10381 =  i_15 &  n_10277;
assign n_10382 = ~n_10380 & ~n_10381;
assign n_10383 =  x_2729 & ~n_10382;
assign n_10384 = ~x_2729 &  n_10382;
assign n_10385 = ~n_10383 & ~n_10384;
assign n_10386 =  x_2728 & ~n_10277;
assign n_10387 =  i_14 &  n_10277;
assign n_10388 = ~n_10386 & ~n_10387;
assign n_10389 =  x_2728 & ~n_10388;
assign n_10390 = ~x_2728 &  n_10388;
assign n_10391 = ~n_10389 & ~n_10390;
assign n_10392 =  x_2727 & ~n_10277;
assign n_10393 =  i_13 &  n_10277;
assign n_10394 = ~n_10392 & ~n_10393;
assign n_10395 =  x_2727 & ~n_10394;
assign n_10396 = ~x_2727 &  n_10394;
assign n_10397 = ~n_10395 & ~n_10396;
assign n_10398 =  x_2726 & ~n_10277;
assign n_10399 =  i_12 &  n_10277;
assign n_10400 = ~n_10398 & ~n_10399;
assign n_10401 =  x_2726 & ~n_10400;
assign n_10402 = ~x_2726 &  n_10400;
assign n_10403 = ~n_10401 & ~n_10402;
assign n_10404 =  x_2725 & ~n_10277;
assign n_10405 =  i_11 &  n_10277;
assign n_10406 = ~n_10404 & ~n_10405;
assign n_10407 =  x_2725 & ~n_10406;
assign n_10408 = ~x_2725 &  n_10406;
assign n_10409 = ~n_10407 & ~n_10408;
assign n_10410 =  x_2724 & ~n_10277;
assign n_10411 =  i_10 &  n_10277;
assign n_10412 = ~n_10410 & ~n_10411;
assign n_10413 =  x_2724 & ~n_10412;
assign n_10414 = ~x_2724 &  n_10412;
assign n_10415 = ~n_10413 & ~n_10414;
assign n_10416 =  x_2723 & ~n_10277;
assign n_10417 =  i_9 &  n_10277;
assign n_10418 = ~n_10416 & ~n_10417;
assign n_10419 =  x_2723 & ~n_10418;
assign n_10420 = ~x_2723 &  n_10418;
assign n_10421 = ~n_10419 & ~n_10420;
assign n_10422 =  x_2722 & ~n_10277;
assign n_10423 =  i_8 &  n_10277;
assign n_10424 = ~n_10422 & ~n_10423;
assign n_10425 =  x_2722 & ~n_10424;
assign n_10426 = ~x_2722 &  n_10424;
assign n_10427 = ~n_10425 & ~n_10426;
assign n_10428 =  x_2721 & ~n_10277;
assign n_10429 =  i_7 &  n_10277;
assign n_10430 = ~n_10428 & ~n_10429;
assign n_10431 =  x_2721 & ~n_10430;
assign n_10432 = ~x_2721 &  n_10430;
assign n_10433 = ~n_10431 & ~n_10432;
assign n_10434 =  x_2720 & ~n_10277;
assign n_10435 =  i_6 &  n_10277;
assign n_10436 = ~n_10434 & ~n_10435;
assign n_10437 =  x_2720 & ~n_10436;
assign n_10438 = ~x_2720 &  n_10436;
assign n_10439 = ~n_10437 & ~n_10438;
assign n_10440 =  x_2719 & ~n_10277;
assign n_10441 =  i_5 &  n_10277;
assign n_10442 = ~n_10440 & ~n_10441;
assign n_10443 =  x_2719 & ~n_10442;
assign n_10444 = ~x_2719 &  n_10442;
assign n_10445 = ~n_10443 & ~n_10444;
assign n_10446 =  x_2718 & ~n_10277;
assign n_10447 =  i_4 &  n_10277;
assign n_10448 = ~n_10446 & ~n_10447;
assign n_10449 =  x_2718 & ~n_10448;
assign n_10450 = ~x_2718 &  n_10448;
assign n_10451 = ~n_10449 & ~n_10450;
assign n_10452 =  x_2717 & ~n_10277;
assign n_10453 =  i_3 &  n_10277;
assign n_10454 = ~n_10452 & ~n_10453;
assign n_10455 =  x_2717 & ~n_10454;
assign n_10456 = ~x_2717 &  n_10454;
assign n_10457 = ~n_10455 & ~n_10456;
assign n_10458 =  x_2716 & ~n_10277;
assign n_10459 =  i_2 &  n_10277;
assign n_10460 = ~n_10458 & ~n_10459;
assign n_10461 =  x_2716 & ~n_10460;
assign n_10462 = ~x_2716 &  n_10460;
assign n_10463 = ~n_10461 & ~n_10462;
assign n_10464 =  x_2715 & ~n_10277;
assign n_10465 =  i_1 &  n_10277;
assign n_10466 = ~n_10464 & ~n_10465;
assign n_10467 =  x_2715 & ~n_10466;
assign n_10468 = ~x_2715 &  n_10466;
assign n_10469 = ~n_10467 & ~n_10468;
assign n_10470 =  n_151 &  n_1502;
assign n_10471 =  n_5981 &  n_10470;
assign n_10472 = ~x_43 &  n_10471;
assign n_10473 =  n_3142 &  n_3632;
assign n_10474 = ~x_43 &  n_10473;
assign n_10475 =  n_1896 &  n_8365;
assign n_10476 =  n_10475 &  n_1502;
assign n_10477 =  n_151 &  n_12;
assign n_10478 =  n_1037 &  n_10477;
assign n_10479 =  n_10478 &  n_1502;
assign n_10480 = ~n_10476 & ~n_10479;
assign n_10481 = ~n_10474 &  n_10480;
assign n_10482 = ~n_10472 &  n_10481;
assign n_10483 =  x_2714 &  n_10482;
assign n_10484 =  x_3863 &  n_10472;
assign n_10485 =  x_3639 &  n_10474;
assign n_10486 =  x_4807 &  n_10479;
assign n_10487 =  x_1962 &  n_10476;
assign n_10488 = ~n_10486 & ~n_10487;
assign n_10489 = ~n_10485 &  n_10488;
assign n_10490 = ~n_10484 &  n_10489;
assign n_10491 = ~n_10483 &  n_10490;
assign n_10492 =  x_2714 & ~n_10491;
assign n_10493 = ~x_2714 &  n_10491;
assign n_10494 = ~n_10492 & ~n_10493;
assign n_10495 =  x_2713 &  n_10482;
assign n_10496 =  x_3862 &  n_10472;
assign n_10497 =  x_3638 &  n_10474;
assign n_10498 =  x_4806 &  n_10479;
assign n_10499 =  x_1961 &  n_10476;
assign n_10500 = ~n_10498 & ~n_10499;
assign n_10501 = ~n_10497 &  n_10500;
assign n_10502 = ~n_10496 &  n_10501;
assign n_10503 = ~n_10495 &  n_10502;
assign n_10504 =  x_2713 & ~n_10503;
assign n_10505 = ~x_2713 &  n_10503;
assign n_10506 = ~n_10504 & ~n_10505;
assign n_10507 =  x_2712 &  n_10482;
assign n_10508 =  x_3861 &  n_10472;
assign n_10509 =  x_3637 &  n_10474;
assign n_10510 =  x_4805 &  n_10479;
assign n_10511 =  x_1960 &  n_10476;
assign n_10512 = ~n_10510 & ~n_10511;
assign n_10513 = ~n_10509 &  n_10512;
assign n_10514 = ~n_10508 &  n_10513;
assign n_10515 = ~n_10507 &  n_10514;
assign n_10516 =  x_2712 & ~n_10515;
assign n_10517 = ~x_2712 &  n_10515;
assign n_10518 = ~n_10516 & ~n_10517;
assign n_10519 =  x_2711 &  n_10482;
assign n_10520 =  x_3860 &  n_10472;
assign n_10521 =  x_3636 &  n_10474;
assign n_10522 =  x_4804 &  n_10479;
assign n_10523 =  x_1959 &  n_10476;
assign n_10524 = ~n_10522 & ~n_10523;
assign n_10525 = ~n_10521 &  n_10524;
assign n_10526 = ~n_10520 &  n_10525;
assign n_10527 = ~n_10519 &  n_10526;
assign n_10528 =  x_2711 & ~n_10527;
assign n_10529 = ~x_2711 &  n_10527;
assign n_10530 = ~n_10528 & ~n_10529;
assign n_10531 =  x_2710 &  n_10482;
assign n_10532 =  x_3859 &  n_10472;
assign n_10533 =  x_3635 &  n_10474;
assign n_10534 =  x_4803 &  n_10479;
assign n_10535 =  x_1958 &  n_10476;
assign n_10536 = ~n_10534 & ~n_10535;
assign n_10537 = ~n_10533 &  n_10536;
assign n_10538 = ~n_10532 &  n_10537;
assign n_10539 = ~n_10531 &  n_10538;
assign n_10540 =  x_2710 & ~n_10539;
assign n_10541 = ~x_2710 &  n_10539;
assign n_10542 = ~n_10540 & ~n_10541;
assign n_10543 =  x_2709 &  n_10482;
assign n_10544 =  x_3858 &  n_10472;
assign n_10545 =  x_3634 &  n_10474;
assign n_10546 =  x_4802 &  n_10479;
assign n_10547 =  x_1957 &  n_10476;
assign n_10548 = ~n_10546 & ~n_10547;
assign n_10549 = ~n_10545 &  n_10548;
assign n_10550 = ~n_10544 &  n_10549;
assign n_10551 = ~n_10543 &  n_10550;
assign n_10552 =  x_2709 & ~n_10551;
assign n_10553 = ~x_2709 &  n_10551;
assign n_10554 = ~n_10552 & ~n_10553;
assign n_10555 =  x_2708 &  n_10482;
assign n_10556 =  x_3857 &  n_10472;
assign n_10557 =  x_3633 &  n_10474;
assign n_10558 =  x_4801 &  n_10479;
assign n_10559 =  x_1956 &  n_10476;
assign n_10560 = ~n_10558 & ~n_10559;
assign n_10561 = ~n_10557 &  n_10560;
assign n_10562 = ~n_10556 &  n_10561;
assign n_10563 = ~n_10555 &  n_10562;
assign n_10564 =  x_2708 & ~n_10563;
assign n_10565 = ~x_2708 &  n_10563;
assign n_10566 = ~n_10564 & ~n_10565;
assign n_10567 =  x_2707 &  n_10482;
assign n_10568 =  x_3856 &  n_10472;
assign n_10569 =  x_3632 &  n_10474;
assign n_10570 =  x_4800 &  n_10479;
assign n_10571 =  x_1955 &  n_10476;
assign n_10572 = ~n_10570 & ~n_10571;
assign n_10573 = ~n_10569 &  n_10572;
assign n_10574 = ~n_10568 &  n_10573;
assign n_10575 = ~n_10567 &  n_10574;
assign n_10576 =  x_2707 & ~n_10575;
assign n_10577 = ~x_2707 &  n_10575;
assign n_10578 = ~n_10576 & ~n_10577;
assign n_10579 =  x_2706 &  n_10482;
assign n_10580 =  x_3855 &  n_10472;
assign n_10581 =  x_3631 &  n_10474;
assign n_10582 =  x_4799 &  n_10479;
assign n_10583 =  x_1954 &  n_10476;
assign n_10584 = ~n_10582 & ~n_10583;
assign n_10585 = ~n_10581 &  n_10584;
assign n_10586 = ~n_10580 &  n_10585;
assign n_10587 = ~n_10579 &  n_10586;
assign n_10588 =  x_2706 & ~n_10587;
assign n_10589 = ~x_2706 &  n_10587;
assign n_10590 = ~n_10588 & ~n_10589;
assign n_10591 =  x_2705 &  n_10482;
assign n_10592 =  x_3854 &  n_10472;
assign n_10593 =  x_3630 &  n_10474;
assign n_10594 =  x_4798 &  n_10479;
assign n_10595 =  x_1953 &  n_10476;
assign n_10596 = ~n_10594 & ~n_10595;
assign n_10597 = ~n_10593 &  n_10596;
assign n_10598 = ~n_10592 &  n_10597;
assign n_10599 = ~n_10591 &  n_10598;
assign n_10600 =  x_2705 & ~n_10599;
assign n_10601 = ~x_2705 &  n_10599;
assign n_10602 = ~n_10600 & ~n_10601;
assign n_10603 =  x_2704 &  n_10482;
assign n_10604 =  x_3853 &  n_10472;
assign n_10605 =  x_3629 &  n_10474;
assign n_10606 =  x_4797 &  n_10479;
assign n_10607 =  x_1952 &  n_10476;
assign n_10608 = ~n_10606 & ~n_10607;
assign n_10609 = ~n_10605 &  n_10608;
assign n_10610 = ~n_10604 &  n_10609;
assign n_10611 = ~n_10603 &  n_10610;
assign n_10612 =  x_2704 & ~n_10611;
assign n_10613 = ~x_2704 &  n_10611;
assign n_10614 = ~n_10612 & ~n_10613;
assign n_10615 =  x_2703 &  n_10482;
assign n_10616 =  x_3852 &  n_10472;
assign n_10617 =  x_3628 &  n_10474;
assign n_10618 =  x_4796 &  n_10479;
assign n_10619 =  x_1951 &  n_10476;
assign n_10620 = ~n_10618 & ~n_10619;
assign n_10621 = ~n_10617 &  n_10620;
assign n_10622 = ~n_10616 &  n_10621;
assign n_10623 = ~n_10615 &  n_10622;
assign n_10624 =  x_2703 & ~n_10623;
assign n_10625 = ~x_2703 &  n_10623;
assign n_10626 = ~n_10624 & ~n_10625;
assign n_10627 =  x_2702 &  n_10482;
assign n_10628 =  x_3851 &  n_10472;
assign n_10629 =  x_3627 &  n_10474;
assign n_10630 =  x_4795 &  n_10479;
assign n_10631 =  x_1950 &  n_10476;
assign n_10632 = ~n_10630 & ~n_10631;
assign n_10633 = ~n_10629 &  n_10632;
assign n_10634 = ~n_10628 &  n_10633;
assign n_10635 = ~n_10627 &  n_10634;
assign n_10636 =  x_2702 & ~n_10635;
assign n_10637 = ~x_2702 &  n_10635;
assign n_10638 = ~n_10636 & ~n_10637;
assign n_10639 =  x_2701 &  n_10482;
assign n_10640 =  x_3850 &  n_10472;
assign n_10641 =  x_3626 &  n_10474;
assign n_10642 =  x_4794 &  n_10479;
assign n_10643 =  x_1949 &  n_10476;
assign n_10644 = ~n_10642 & ~n_10643;
assign n_10645 = ~n_10641 &  n_10644;
assign n_10646 = ~n_10640 &  n_10645;
assign n_10647 = ~n_10639 &  n_10646;
assign n_10648 =  x_2701 & ~n_10647;
assign n_10649 = ~x_2701 &  n_10647;
assign n_10650 = ~n_10648 & ~n_10649;
assign n_10651 =  x_2700 &  n_10482;
assign n_10652 =  x_3849 &  n_10472;
assign n_10653 =  x_3625 &  n_10474;
assign n_10654 =  x_4793 &  n_10479;
assign n_10655 =  x_1948 &  n_10476;
assign n_10656 = ~n_10654 & ~n_10655;
assign n_10657 = ~n_10653 &  n_10656;
assign n_10658 = ~n_10652 &  n_10657;
assign n_10659 = ~n_10651 &  n_10658;
assign n_10660 =  x_2700 & ~n_10659;
assign n_10661 = ~x_2700 &  n_10659;
assign n_10662 = ~n_10660 & ~n_10661;
assign n_10663 =  x_2699 &  n_10482;
assign n_10664 =  x_3848 &  n_10472;
assign n_10665 =  x_3624 &  n_10474;
assign n_10666 =  x_4792 &  n_10479;
assign n_10667 =  x_1947 &  n_10476;
assign n_10668 = ~n_10666 & ~n_10667;
assign n_10669 = ~n_10665 &  n_10668;
assign n_10670 = ~n_10664 &  n_10669;
assign n_10671 = ~n_10663 &  n_10670;
assign n_10672 =  x_2699 & ~n_10671;
assign n_10673 = ~x_2699 &  n_10671;
assign n_10674 = ~n_10672 & ~n_10673;
assign n_10675 =  x_2698 &  n_10482;
assign n_10676 =  x_3847 &  n_10472;
assign n_10677 =  x_3623 &  n_10474;
assign n_10678 =  x_4791 &  n_10479;
assign n_10679 =  x_1946 &  n_10476;
assign n_10680 = ~n_10678 & ~n_10679;
assign n_10681 = ~n_10677 &  n_10680;
assign n_10682 = ~n_10676 &  n_10681;
assign n_10683 = ~n_10675 &  n_10682;
assign n_10684 =  x_2698 & ~n_10683;
assign n_10685 = ~x_2698 &  n_10683;
assign n_10686 = ~n_10684 & ~n_10685;
assign n_10687 =  x_2697 &  n_10482;
assign n_10688 =  x_3846 &  n_10472;
assign n_10689 =  x_3622 &  n_10474;
assign n_10690 =  x_4790 &  n_10479;
assign n_10691 =  x_1945 &  n_10476;
assign n_10692 = ~n_10690 & ~n_10691;
assign n_10693 = ~n_10689 &  n_10692;
assign n_10694 = ~n_10688 &  n_10693;
assign n_10695 = ~n_10687 &  n_10694;
assign n_10696 =  x_2697 & ~n_10695;
assign n_10697 = ~x_2697 &  n_10695;
assign n_10698 = ~n_10696 & ~n_10697;
assign n_10699 =  x_2696 &  n_10482;
assign n_10700 =  x_3845 &  n_10472;
assign n_10701 =  x_3621 &  n_10474;
assign n_10702 =  x_4789 &  n_10479;
assign n_10703 =  x_1944 &  n_10476;
assign n_10704 = ~n_10702 & ~n_10703;
assign n_10705 = ~n_10701 &  n_10704;
assign n_10706 = ~n_10700 &  n_10705;
assign n_10707 = ~n_10699 &  n_10706;
assign n_10708 =  x_2696 & ~n_10707;
assign n_10709 = ~x_2696 &  n_10707;
assign n_10710 = ~n_10708 & ~n_10709;
assign n_10711 =  x_2695 &  n_10482;
assign n_10712 =  x_3844 &  n_10472;
assign n_10713 =  x_3620 &  n_10474;
assign n_10714 =  x_4788 &  n_10479;
assign n_10715 =  x_1943 &  n_10476;
assign n_10716 = ~n_10714 & ~n_10715;
assign n_10717 = ~n_10713 &  n_10716;
assign n_10718 = ~n_10712 &  n_10717;
assign n_10719 = ~n_10711 &  n_10718;
assign n_10720 =  x_2695 & ~n_10719;
assign n_10721 = ~x_2695 &  n_10719;
assign n_10722 = ~n_10720 & ~n_10721;
assign n_10723 =  x_2694 &  n_10482;
assign n_10724 =  x_3843 &  n_10472;
assign n_10725 =  x_3619 &  n_10474;
assign n_10726 =  x_4787 &  n_10479;
assign n_10727 =  x_1942 &  n_10476;
assign n_10728 = ~n_10726 & ~n_10727;
assign n_10729 = ~n_10725 &  n_10728;
assign n_10730 = ~n_10724 &  n_10729;
assign n_10731 = ~n_10723 &  n_10730;
assign n_10732 =  x_2694 & ~n_10731;
assign n_10733 = ~x_2694 &  n_10731;
assign n_10734 = ~n_10732 & ~n_10733;
assign n_10735 =  x_2693 &  n_10482;
assign n_10736 =  x_3842 &  n_10472;
assign n_10737 =  x_3618 &  n_10474;
assign n_10738 =  x_4786 &  n_10479;
assign n_10739 =  x_1941 &  n_10476;
assign n_10740 = ~n_10738 & ~n_10739;
assign n_10741 = ~n_10737 &  n_10740;
assign n_10742 = ~n_10736 &  n_10741;
assign n_10743 = ~n_10735 &  n_10742;
assign n_10744 =  x_2693 & ~n_10743;
assign n_10745 = ~x_2693 &  n_10743;
assign n_10746 = ~n_10744 & ~n_10745;
assign n_10747 =  x_2692 &  n_10482;
assign n_10748 =  x_3841 &  n_10472;
assign n_10749 =  x_3617 &  n_10474;
assign n_10750 =  x_4785 &  n_10479;
assign n_10751 =  x_1940 &  n_10476;
assign n_10752 = ~n_10750 & ~n_10751;
assign n_10753 = ~n_10749 &  n_10752;
assign n_10754 = ~n_10748 &  n_10753;
assign n_10755 = ~n_10747 &  n_10754;
assign n_10756 =  x_2692 & ~n_10755;
assign n_10757 = ~x_2692 &  n_10755;
assign n_10758 = ~n_10756 & ~n_10757;
assign n_10759 =  x_2691 &  n_10482;
assign n_10760 =  x_3840 &  n_10472;
assign n_10761 =  x_3616 &  n_10474;
assign n_10762 =  x_4784 &  n_10479;
assign n_10763 =  x_1939 &  n_10476;
assign n_10764 = ~n_10762 & ~n_10763;
assign n_10765 = ~n_10761 &  n_10764;
assign n_10766 = ~n_10760 &  n_10765;
assign n_10767 = ~n_10759 &  n_10766;
assign n_10768 =  x_2691 & ~n_10767;
assign n_10769 = ~x_2691 &  n_10767;
assign n_10770 = ~n_10768 & ~n_10769;
assign n_10771 =  x_2690 &  n_10482;
assign n_10772 =  x_3839 &  n_10472;
assign n_10773 =  x_3615 &  n_10474;
assign n_10774 =  x_4783 &  n_10479;
assign n_10775 =  x_1938 &  n_10476;
assign n_10776 = ~n_10774 & ~n_10775;
assign n_10777 = ~n_10773 &  n_10776;
assign n_10778 = ~n_10772 &  n_10777;
assign n_10779 = ~n_10771 &  n_10778;
assign n_10780 =  x_2690 & ~n_10779;
assign n_10781 = ~x_2690 &  n_10779;
assign n_10782 = ~n_10780 & ~n_10781;
assign n_10783 =  x_2689 &  n_10482;
assign n_10784 =  x_3838 &  n_10472;
assign n_10785 =  x_3614 &  n_10474;
assign n_10786 =  x_4782 &  n_10479;
assign n_10787 =  x_1937 &  n_10476;
assign n_10788 = ~n_10786 & ~n_10787;
assign n_10789 = ~n_10785 &  n_10788;
assign n_10790 = ~n_10784 &  n_10789;
assign n_10791 = ~n_10783 &  n_10790;
assign n_10792 =  x_2689 & ~n_10791;
assign n_10793 = ~x_2689 &  n_10791;
assign n_10794 = ~n_10792 & ~n_10793;
assign n_10795 =  x_2688 &  n_10482;
assign n_10796 =  x_3837 &  n_10472;
assign n_10797 =  x_3613 &  n_10474;
assign n_10798 =  x_4781 &  n_10479;
assign n_10799 =  x_1936 &  n_10476;
assign n_10800 = ~n_10798 & ~n_10799;
assign n_10801 = ~n_10797 &  n_10800;
assign n_10802 = ~n_10796 &  n_10801;
assign n_10803 = ~n_10795 &  n_10802;
assign n_10804 =  x_2688 & ~n_10803;
assign n_10805 = ~x_2688 &  n_10803;
assign n_10806 = ~n_10804 & ~n_10805;
assign n_10807 =  x_2687 &  n_10482;
assign n_10808 =  x_3836 &  n_10472;
assign n_10809 =  x_3612 &  n_10474;
assign n_10810 =  x_4780 &  n_10479;
assign n_10811 =  x_1935 &  n_10476;
assign n_10812 = ~n_10810 & ~n_10811;
assign n_10813 = ~n_10809 &  n_10812;
assign n_10814 = ~n_10808 &  n_10813;
assign n_10815 = ~n_10807 &  n_10814;
assign n_10816 =  x_2687 & ~n_10815;
assign n_10817 = ~x_2687 &  n_10815;
assign n_10818 = ~n_10816 & ~n_10817;
assign n_10819 =  x_2686 &  n_10482;
assign n_10820 =  x_3835 &  n_10472;
assign n_10821 =  x_3611 &  n_10474;
assign n_10822 =  x_4779 &  n_10479;
assign n_10823 =  x_1934 &  n_10476;
assign n_10824 = ~n_10822 & ~n_10823;
assign n_10825 = ~n_10821 &  n_10824;
assign n_10826 = ~n_10820 &  n_10825;
assign n_10827 = ~n_10819 &  n_10826;
assign n_10828 =  x_2686 & ~n_10827;
assign n_10829 = ~x_2686 &  n_10827;
assign n_10830 = ~n_10828 & ~n_10829;
assign n_10831 =  x_2685 &  n_10482;
assign n_10832 =  x_3834 &  n_10472;
assign n_10833 =  x_3610 &  n_10474;
assign n_10834 =  x_4778 &  n_10479;
assign n_10835 =  x_1933 &  n_10476;
assign n_10836 = ~n_10834 & ~n_10835;
assign n_10837 = ~n_10833 &  n_10836;
assign n_10838 = ~n_10832 &  n_10837;
assign n_10839 = ~n_10831 &  n_10838;
assign n_10840 =  x_2685 & ~n_10839;
assign n_10841 = ~x_2685 &  n_10839;
assign n_10842 = ~n_10840 & ~n_10841;
assign n_10843 =  x_2684 &  n_10482;
assign n_10844 =  x_3833 &  n_10472;
assign n_10845 =  x_3609 &  n_10474;
assign n_10846 =  x_4777 &  n_10479;
assign n_10847 =  x_1932 &  n_10476;
assign n_10848 = ~n_10846 & ~n_10847;
assign n_10849 = ~n_10845 &  n_10848;
assign n_10850 = ~n_10844 &  n_10849;
assign n_10851 = ~n_10843 &  n_10850;
assign n_10852 =  x_2684 & ~n_10851;
assign n_10853 = ~x_2684 &  n_10851;
assign n_10854 = ~n_10852 & ~n_10853;
assign n_10855 =  x_2683 &  n_10482;
assign n_10856 =  x_3832 &  n_10472;
assign n_10857 =  x_3608 &  n_10474;
assign n_10858 =  x_4776 &  n_10479;
assign n_10859 =  x_1931 &  n_10476;
assign n_10860 = ~n_10858 & ~n_10859;
assign n_10861 = ~n_10857 &  n_10860;
assign n_10862 = ~n_10856 &  n_10861;
assign n_10863 = ~n_10855 &  n_10862;
assign n_10864 =  x_2683 & ~n_10863;
assign n_10865 = ~x_2683 &  n_10863;
assign n_10866 = ~n_10864 & ~n_10865;
assign n_10867 =  n_765 &  n_1041;
assign n_10868 =  x_40 &  n_152;
assign n_10869 =  n_10867 &  n_10868;
assign n_10870 = ~x_43 &  n_10869;
assign n_10871 =  x_43 &  n_3630;
assign n_10872 = ~x_40 &  n_1038;
assign n_10873 =  n_10872 &  n_10867;
assign n_10874 =  n_554 &  n_1305;
assign n_10875 =  n_1306 &  n_10874;
assign n_10876 = ~n_10873 & ~n_10875;
assign n_10877 = ~n_10871 &  n_10876;
assign n_10878 = ~n_10870 &  n_10877;
assign n_10879 =  x_2682 &  n_10878;
assign n_10880 =  x_2026 &  x_3831;
assign n_10881 = ~x_2026 & ~x_3831;
assign n_10882 = ~n_10880 & ~n_10881;
assign n_10883 =  n_10870 &  n_10882;
assign n_10884 =  x_2250 &  x_3767;
assign n_10885 = ~x_2250 & ~x_3767;
assign n_10886 = ~n_10884 & ~n_10885;
assign n_10887 =  n_10871 &  n_10886;
assign n_10888 =  x_4839 &  n_10875;
assign n_10889 =  x_1514 &  x_4200;
assign n_10890 = ~x_1514 & ~x_4200;
assign n_10891 = ~n_10889 & ~n_10890;
assign n_10892 =  n_10873 &  n_10891;
assign n_10893 = ~n_10888 & ~n_10892;
assign n_10894 = ~n_10887 &  n_10893;
assign n_10895 = ~n_10883 &  n_10894;
assign n_10896 = ~n_10879 &  n_10895;
assign n_10897 =  x_2682 & ~n_10896;
assign n_10898 = ~x_2682 &  n_10896;
assign n_10899 = ~n_10897 & ~n_10898;
assign n_10900 =  x_2681 &  n_10878;
assign n_10901 =  x_4838 &  n_10875;
assign n_10902 = ~x_1513 & ~x_1514;
assign n_10903 =  x_1513 &  x_1514;
assign n_10904 = ~n_10902 & ~n_10903;
assign n_10905 =  x_4199 &  n_10904;
assign n_10906 = ~x_4199 & ~n_10904;
assign n_10907 = ~n_10905 & ~n_10906;
assign n_10908 =  n_10889 &  n_10907;
assign n_10909 = ~n_10889 & ~n_10907;
assign n_10910 =  n_10873 & ~n_10909;
assign n_10911 = ~n_10908 &  n_10910;
assign n_10912 = ~n_10901 & ~n_10911;
assign n_10913 = ~x_2025 & ~x_2026;
assign n_10914 =  x_2025 &  x_2026;
assign n_10915 = ~n_10913 & ~n_10914;
assign n_10916 =  x_3830 &  n_10915;
assign n_10917 = ~x_3830 & ~n_10915;
assign n_10918 = ~n_10916 & ~n_10917;
assign n_10919 =  n_10880 &  n_10918;
assign n_10920 = ~n_10880 & ~n_10918;
assign n_10921 =  n_10870 & ~n_10920;
assign n_10922 = ~n_10919 &  n_10921;
assign n_10923 = ~x_3766 & ~x_3767;
assign n_10924 =  x_3766 &  x_3767;
assign n_10925 = ~n_10923 & ~n_10924;
assign n_10926 =  x_2249 &  n_10925;
assign n_10927 = ~x_2249 & ~n_10925;
assign n_10928 = ~n_10926 & ~n_10927;
assign n_10929 = ~n_10884 & ~n_10928;
assign n_10930 =  n_10884 &  n_10928;
assign n_10931 =  n_10871 & ~n_10930;
assign n_10932 = ~n_10929 &  n_10931;
assign n_10933 = ~n_10922 & ~n_10932;
assign n_10934 =  n_10912 &  n_10933;
assign n_10935 = ~n_10900 &  n_10934;
assign n_10936 =  x_2681 & ~n_10935;
assign n_10937 = ~x_2681 &  n_10935;
assign n_10938 = ~n_10936 & ~n_10937;
assign n_10939 = ~x_1512 &  n_10902;
assign n_10940 =  x_1512 & ~n_10902;
assign n_10941 = ~n_10939 & ~n_10940;
assign n_10942 =  x_1513 & ~x_4199;
assign n_10943 =  n_10889 & ~n_10942;
assign n_10944 = ~n_10943 & ~n_10905;
assign n_10945 =  n_10941 & ~n_10944;
assign n_10946 = ~n_10941 &  n_10944;
assign n_10947 = ~n_10945 & ~n_10946;
assign n_10948 = ~x_4198 & ~n_10947;
assign n_10949 =  x_4198 & ~n_10946;
assign n_10950 = ~n_10945 &  n_10949;
assign n_10951 =  n_10873 & ~n_10950;
assign n_10952 = ~n_10948 &  n_10951;
assign n_10953 =  x_2680 &  n_10878;
assign n_10954 =  x_4837 &  n_10875;
assign n_10955 = ~n_10953 & ~n_10954;
assign n_10956 = ~n_10952 &  n_10955;
assign n_10957 = ~x_2024 &  n_10913;
assign n_10958 =  x_2024 & ~n_10913;
assign n_10959 = ~n_10957 & ~n_10958;
assign n_10960 =  x_2025 & ~x_3830;
assign n_10961 =  n_10880 & ~n_10960;
assign n_10962 = ~n_10961 & ~n_10916;
assign n_10963 =  n_10959 & ~n_10962;
assign n_10964 = ~n_10959 &  n_10962;
assign n_10965 = ~n_10963 & ~n_10964;
assign n_10966 = ~x_3829 & ~n_10965;
assign n_10967 =  x_3829 & ~n_10964;
assign n_10968 = ~n_10963 &  n_10967;
assign n_10969 =  n_10870 & ~n_10968;
assign n_10970 = ~n_10966 &  n_10969;
assign n_10971 = ~x_3765 &  n_10923;
assign n_10972 =  x_3765 & ~n_10923;
assign n_10973 = ~n_10971 & ~n_10972;
assign n_10974 = ~x_2249 &  x_3766;
assign n_10975 =  n_10884 & ~n_10974;
assign n_10976 = ~n_10975 & ~n_10926;
assign n_10977 =  n_10973 & ~n_10976;
assign n_10978 = ~n_10973 &  n_10976;
assign n_10979 = ~n_10977 & ~n_10978;
assign n_10980 =  x_2248 &  n_10979;
assign n_10981 = ~x_2248 & ~n_10979;
assign n_10982 =  n_10871 & ~n_10981;
assign n_10983 = ~n_10980 &  n_10982;
assign n_10984 = ~n_10970 & ~n_10983;
assign n_10985 =  n_10956 &  n_10984;
assign n_10986 =  x_2680 & ~n_10985;
assign n_10987 = ~x_2680 &  n_10985;
assign n_10988 = ~n_10986 & ~n_10987;
assign n_10989 = ~x_2023 &  n_10957;
assign n_10990 =  x_2023 & ~n_10957;
assign n_10991 = ~n_10989 & ~n_10990;
assign n_10992 = ~n_10963 & ~n_10967;
assign n_10993 =  n_10991 & ~n_10992;
assign n_10994 = ~n_10991 &  n_10992;
assign n_10995 = ~n_10993 & ~n_10994;
assign n_10996 = ~x_3828 & ~n_10995;
assign n_10997 =  x_3828 & ~n_10994;
assign n_10998 = ~n_10993 &  n_10997;
assign n_10999 =  n_10870 & ~n_10998;
assign n_11000 = ~n_10996 &  n_10999;
assign n_11001 =  x_2679 &  n_10878;
assign n_11002 =  x_4836 &  n_10875;
assign n_11003 = ~n_11001 & ~n_11002;
assign n_11004 = ~n_11000 &  n_11003;
assign n_11005 = ~x_1511 &  n_10939;
assign n_11006 =  x_1511 & ~n_10939;
assign n_11007 = ~n_11005 & ~n_11006;
assign n_11008 = ~n_10945 & ~n_10949;
assign n_11009 =  n_11007 & ~n_11008;
assign n_11010 = ~n_11007 &  n_11008;
assign n_11011 = ~n_11009 & ~n_11010;
assign n_11012 = ~x_4197 & ~n_11011;
assign n_11013 =  x_4197 & ~n_11010;
assign n_11014 = ~n_11009 &  n_11013;
assign n_11015 =  n_10873 & ~n_11014;
assign n_11016 = ~n_11012 &  n_11015;
assign n_11017 = ~x_3764 &  n_10971;
assign n_11018 =  x_3764 & ~n_10971;
assign n_11019 = ~n_11017 & ~n_11018;
assign n_11020 =  x_2248 & ~n_10978;
assign n_11021 = ~n_10977 & ~n_11020;
assign n_11022 =  n_11019 & ~n_11021;
assign n_11023 = ~n_11019 &  n_11021;
assign n_11024 = ~n_11022 & ~n_11023;
assign n_11025 = ~x_2247 & ~n_11024;
assign n_11026 =  x_2247 & ~n_11023;
assign n_11027 = ~n_11022 &  n_11026;
assign n_11028 =  n_10871 & ~n_11027;
assign n_11029 = ~n_11025 &  n_11028;
assign n_11030 = ~n_11016 & ~n_11029;
assign n_11031 =  n_11004 &  n_11030;
assign n_11032 =  x_2679 & ~n_11031;
assign n_11033 = ~x_2679 &  n_11031;
assign n_11034 = ~n_11032 & ~n_11033;
assign n_11035 = ~x_3763 &  n_11017;
assign n_11036 =  x_3763 & ~n_11017;
assign n_11037 = ~n_11035 & ~n_11036;
assign n_11038 = ~n_11022 & ~n_11026;
assign n_11039 =  n_11037 & ~n_11038;
assign n_11040 = ~n_11037 &  n_11038;
assign n_11041 = ~n_11039 & ~n_11040;
assign n_11042 = ~x_2246 & ~n_11041;
assign n_11043 =  x_2246 & ~n_11040;
assign n_11044 = ~n_11039 &  n_11043;
assign n_11045 =  n_10871 & ~n_11044;
assign n_11046 = ~n_11042 &  n_11045;
assign n_11047 =  x_2678 &  n_10878;
assign n_11048 =  x_4835 &  n_10875;
assign n_11049 = ~n_11047 & ~n_11048;
assign n_11050 = ~n_11046 &  n_11049;
assign n_11051 = ~x_1510 &  n_11005;
assign n_11052 =  x_1510 & ~n_11005;
assign n_11053 = ~n_11051 & ~n_11052;
assign n_11054 = ~n_11009 & ~n_11013;
assign n_11055 =  n_11053 & ~n_11054;
assign n_11056 = ~n_11053 &  n_11054;
assign n_11057 = ~n_11055 & ~n_11056;
assign n_11058 = ~x_4196 & ~n_11057;
assign n_11059 =  x_4196 & ~n_11056;
assign n_11060 = ~n_11055 &  n_11059;
assign n_11061 =  n_10873 & ~n_11060;
assign n_11062 = ~n_11058 &  n_11061;
assign n_11063 = ~x_2022 &  n_10989;
assign n_11064 =  x_2022 & ~n_10989;
assign n_11065 = ~n_11063 & ~n_11064;
assign n_11066 = ~n_10993 & ~n_10997;
assign n_11067 =  n_11065 & ~n_11066;
assign n_11068 = ~n_11065 &  n_11066;
assign n_11069 = ~n_11067 & ~n_11068;
assign n_11070 = ~x_3827 & ~n_11069;
assign n_11071 =  x_3827 & ~n_11068;
assign n_11072 = ~n_11067 &  n_11071;
assign n_11073 =  n_10870 & ~n_11072;
assign n_11074 = ~n_11070 &  n_11073;
assign n_11075 = ~n_11062 & ~n_11074;
assign n_11076 =  n_11050 &  n_11075;
assign n_11077 =  x_2678 & ~n_11076;
assign n_11078 = ~x_2678 &  n_11076;
assign n_11079 = ~n_11077 & ~n_11078;
assign n_11080 = ~x_3762 &  n_11035;
assign n_11081 =  x_3762 & ~n_11035;
assign n_11082 = ~n_11080 & ~n_11081;
assign n_11083 = ~n_11039 & ~n_11043;
assign n_11084 =  n_11082 & ~n_11083;
assign n_11085 = ~n_11082 &  n_11083;
assign n_11086 = ~n_11084 & ~n_11085;
assign n_11087 = ~x_2245 & ~n_11086;
assign n_11088 =  x_2245 & ~n_11085;
assign n_11089 = ~n_11084 &  n_11088;
assign n_11090 =  n_10871 & ~n_11089;
assign n_11091 = ~n_11087 &  n_11090;
assign n_11092 =  x_2677 &  n_10878;
assign n_11093 =  x_4834 &  n_10875;
assign n_11094 = ~n_11092 & ~n_11093;
assign n_11095 = ~n_11091 &  n_11094;
assign n_11096 = ~x_1509 &  n_11051;
assign n_11097 =  x_1509 & ~n_11051;
assign n_11098 = ~n_11096 & ~n_11097;
assign n_11099 = ~n_11055 & ~n_11059;
assign n_11100 =  n_11098 & ~n_11099;
assign n_11101 = ~n_11098 &  n_11099;
assign n_11102 = ~n_11100 & ~n_11101;
assign n_11103 = ~x_4195 & ~n_11102;
assign n_11104 =  x_4195 & ~n_11101;
assign n_11105 = ~n_11100 &  n_11104;
assign n_11106 =  n_10873 & ~n_11105;
assign n_11107 = ~n_11103 &  n_11106;
assign n_11108 = ~x_2021 &  n_11063;
assign n_11109 =  x_2021 & ~n_11063;
assign n_11110 = ~n_11108 & ~n_11109;
assign n_11111 = ~n_11067 & ~n_11071;
assign n_11112 =  n_11110 & ~n_11111;
assign n_11113 = ~n_11110 &  n_11111;
assign n_11114 = ~n_11112 & ~n_11113;
assign n_11115 = ~x_3826 & ~n_11114;
assign n_11116 =  x_3826 & ~n_11113;
assign n_11117 = ~n_11112 &  n_11116;
assign n_11118 =  n_10870 & ~n_11117;
assign n_11119 = ~n_11115 &  n_11118;
assign n_11120 = ~n_11107 & ~n_11119;
assign n_11121 =  n_11095 &  n_11120;
assign n_11122 =  x_2677 & ~n_11121;
assign n_11123 = ~x_2677 &  n_11121;
assign n_11124 = ~n_11122 & ~n_11123;
assign n_11125 = ~x_3761 &  n_11080;
assign n_11126 =  x_3761 & ~n_11080;
assign n_11127 = ~n_11125 & ~n_11126;
assign n_11128 = ~n_11084 & ~n_11088;
assign n_11129 =  n_11127 & ~n_11128;
assign n_11130 = ~n_11127 &  n_11128;
assign n_11131 = ~n_11129 & ~n_11130;
assign n_11132 = ~x_2244 & ~n_11131;
assign n_11133 =  x_2244 & ~n_11130;
assign n_11134 = ~n_11129 &  n_11133;
assign n_11135 =  n_10871 & ~n_11134;
assign n_11136 = ~n_11132 &  n_11135;
assign n_11137 =  x_2676 &  n_10878;
assign n_11138 =  x_4833 &  n_10875;
assign n_11139 = ~n_11137 & ~n_11138;
assign n_11140 = ~n_11136 &  n_11139;
assign n_11141 = ~x_1508 &  n_11096;
assign n_11142 =  x_1508 & ~n_11096;
assign n_11143 = ~n_11141 & ~n_11142;
assign n_11144 = ~n_11100 & ~n_11104;
assign n_11145 =  n_11143 & ~n_11144;
assign n_11146 = ~n_11143 &  n_11144;
assign n_11147 = ~n_11145 & ~n_11146;
assign n_11148 = ~x_4194 & ~n_11147;
assign n_11149 =  x_4194 & ~n_11146;
assign n_11150 = ~n_11145 &  n_11149;
assign n_11151 =  n_10873 & ~n_11150;
assign n_11152 = ~n_11148 &  n_11151;
assign n_11153 = ~x_2020 &  n_11108;
assign n_11154 =  x_2020 & ~n_11108;
assign n_11155 = ~n_11153 & ~n_11154;
assign n_11156 = ~n_11112 & ~n_11116;
assign n_11157 =  n_11155 & ~n_11156;
assign n_11158 = ~n_11155 &  n_11156;
assign n_11159 = ~n_11157 & ~n_11158;
assign n_11160 = ~x_3825 & ~n_11159;
assign n_11161 =  x_3825 & ~n_11158;
assign n_11162 = ~n_11157 &  n_11161;
assign n_11163 =  n_10870 & ~n_11162;
assign n_11164 = ~n_11160 &  n_11163;
assign n_11165 = ~n_11152 & ~n_11164;
assign n_11166 =  n_11140 &  n_11165;
assign n_11167 =  x_2676 & ~n_11166;
assign n_11168 = ~x_2676 &  n_11166;
assign n_11169 = ~n_11167 & ~n_11168;
assign n_11170 = ~x_3760 &  n_11125;
assign n_11171 =  x_3760 & ~n_11125;
assign n_11172 = ~n_11170 & ~n_11171;
assign n_11173 = ~n_11129 & ~n_11133;
assign n_11174 =  n_11172 & ~n_11173;
assign n_11175 = ~n_11172 &  n_11173;
assign n_11176 = ~n_11174 & ~n_11175;
assign n_11177 = ~x_2243 & ~n_11176;
assign n_11178 =  x_2243 & ~n_11175;
assign n_11179 = ~n_11174 &  n_11178;
assign n_11180 =  n_10871 & ~n_11179;
assign n_11181 = ~n_11177 &  n_11180;
assign n_11182 =  x_2675 &  n_10878;
assign n_11183 =  x_4832 &  n_10875;
assign n_11184 = ~n_11182 & ~n_11183;
assign n_11185 = ~n_11181 &  n_11184;
assign n_11186 = ~x_1507 &  n_11141;
assign n_11187 =  x_1507 & ~n_11141;
assign n_11188 = ~n_11186 & ~n_11187;
assign n_11189 = ~n_11145 & ~n_11149;
assign n_11190 =  n_11188 & ~n_11189;
assign n_11191 = ~n_11188 &  n_11189;
assign n_11192 = ~n_11190 & ~n_11191;
assign n_11193 = ~x_4193 & ~n_11192;
assign n_11194 =  x_4193 & ~n_11191;
assign n_11195 = ~n_11190 &  n_11194;
assign n_11196 =  n_10873 & ~n_11195;
assign n_11197 = ~n_11193 &  n_11196;
assign n_11198 = ~x_2019 &  n_11153;
assign n_11199 =  x_2019 & ~n_11153;
assign n_11200 = ~n_11198 & ~n_11199;
assign n_11201 = ~n_11157 & ~n_11161;
assign n_11202 =  n_11200 & ~n_11201;
assign n_11203 = ~n_11200 &  n_11201;
assign n_11204 = ~n_11202 & ~n_11203;
assign n_11205 = ~x_3824 & ~n_11204;
assign n_11206 =  x_3824 & ~n_11203;
assign n_11207 = ~n_11202 &  n_11206;
assign n_11208 =  n_10870 & ~n_11207;
assign n_11209 = ~n_11205 &  n_11208;
assign n_11210 = ~n_11197 & ~n_11209;
assign n_11211 =  n_11185 &  n_11210;
assign n_11212 =  x_2675 & ~n_11211;
assign n_11213 = ~x_2675 &  n_11211;
assign n_11214 = ~n_11212 & ~n_11213;
assign n_11215 = ~x_3759 &  n_11170;
assign n_11216 =  x_3759 & ~n_11170;
assign n_11217 = ~n_11215 & ~n_11216;
assign n_11218 = ~n_11174 & ~n_11178;
assign n_11219 =  n_11217 & ~n_11218;
assign n_11220 = ~n_11217 &  n_11218;
assign n_11221 = ~n_11219 & ~n_11220;
assign n_11222 = ~x_2242 & ~n_11221;
assign n_11223 =  x_2242 & ~n_11220;
assign n_11224 = ~n_11219 &  n_11223;
assign n_11225 =  n_10871 & ~n_11224;
assign n_11226 = ~n_11222 &  n_11225;
assign n_11227 =  x_2674 &  n_10878;
assign n_11228 =  x_4831 &  n_10875;
assign n_11229 = ~n_11227 & ~n_11228;
assign n_11230 = ~n_11226 &  n_11229;
assign n_11231 = ~x_1506 &  n_11186;
assign n_11232 =  x_1506 & ~n_11186;
assign n_11233 = ~n_11231 & ~n_11232;
assign n_11234 = ~n_11190 & ~n_11194;
assign n_11235 =  n_11233 & ~n_11234;
assign n_11236 = ~n_11233 &  n_11234;
assign n_11237 = ~n_11235 & ~n_11236;
assign n_11238 = ~x_4192 & ~n_11237;
assign n_11239 =  x_4192 & ~n_11236;
assign n_11240 = ~n_11235 &  n_11239;
assign n_11241 =  n_10873 & ~n_11240;
assign n_11242 = ~n_11238 &  n_11241;
assign n_11243 = ~x_2018 &  n_11198;
assign n_11244 =  x_2018 & ~n_11198;
assign n_11245 = ~n_11243 & ~n_11244;
assign n_11246 = ~n_11202 & ~n_11206;
assign n_11247 =  n_11245 & ~n_11246;
assign n_11248 = ~n_11245 &  n_11246;
assign n_11249 = ~n_11247 & ~n_11248;
assign n_11250 = ~x_3823 & ~n_11249;
assign n_11251 =  x_3823 & ~n_11248;
assign n_11252 = ~n_11247 &  n_11251;
assign n_11253 =  n_10870 & ~n_11252;
assign n_11254 = ~n_11250 &  n_11253;
assign n_11255 = ~n_11242 & ~n_11254;
assign n_11256 =  n_11230 &  n_11255;
assign n_11257 =  x_2674 & ~n_11256;
assign n_11258 = ~x_2674 &  n_11256;
assign n_11259 = ~n_11257 & ~n_11258;
assign n_11260 = ~x_3758 &  n_11215;
assign n_11261 =  x_3758 & ~n_11215;
assign n_11262 = ~n_11260 & ~n_11261;
assign n_11263 = ~n_11219 & ~n_11223;
assign n_11264 =  n_11262 & ~n_11263;
assign n_11265 = ~n_11262 &  n_11263;
assign n_11266 = ~n_11264 & ~n_11265;
assign n_11267 = ~x_2241 & ~n_11266;
assign n_11268 =  x_2241 & ~n_11265;
assign n_11269 = ~n_11264 &  n_11268;
assign n_11270 =  n_10871 & ~n_11269;
assign n_11271 = ~n_11267 &  n_11270;
assign n_11272 =  x_2673 &  n_10878;
assign n_11273 =  x_4830 &  n_10875;
assign n_11274 = ~n_11272 & ~n_11273;
assign n_11275 = ~n_11271 &  n_11274;
assign n_11276 = ~x_1505 &  n_11231;
assign n_11277 =  x_1505 & ~n_11231;
assign n_11278 = ~n_11276 & ~n_11277;
assign n_11279 = ~n_11235 & ~n_11239;
assign n_11280 =  n_11278 & ~n_11279;
assign n_11281 = ~n_11278 &  n_11279;
assign n_11282 = ~n_11280 & ~n_11281;
assign n_11283 = ~x_4191 & ~n_11282;
assign n_11284 =  x_4191 & ~n_11281;
assign n_11285 = ~n_11280 &  n_11284;
assign n_11286 =  n_10873 & ~n_11285;
assign n_11287 = ~n_11283 &  n_11286;
assign n_11288 = ~x_2017 &  n_11243;
assign n_11289 =  x_2017 & ~n_11243;
assign n_11290 = ~n_11288 & ~n_11289;
assign n_11291 = ~n_11247 & ~n_11251;
assign n_11292 =  n_11290 & ~n_11291;
assign n_11293 = ~n_11290 &  n_11291;
assign n_11294 = ~n_11292 & ~n_11293;
assign n_11295 = ~x_3822 & ~n_11294;
assign n_11296 =  x_3822 & ~n_11293;
assign n_11297 = ~n_11292 &  n_11296;
assign n_11298 =  n_10870 & ~n_11297;
assign n_11299 = ~n_11295 &  n_11298;
assign n_11300 = ~n_11287 & ~n_11299;
assign n_11301 =  n_11275 &  n_11300;
assign n_11302 =  x_2673 & ~n_11301;
assign n_11303 = ~x_2673 &  n_11301;
assign n_11304 = ~n_11302 & ~n_11303;
assign n_11305 = ~x_3757 &  n_11260;
assign n_11306 =  x_3757 & ~n_11260;
assign n_11307 = ~n_11305 & ~n_11306;
assign n_11308 = ~n_11264 & ~n_11268;
assign n_11309 =  n_11307 & ~n_11308;
assign n_11310 = ~n_11307 &  n_11308;
assign n_11311 = ~n_11309 & ~n_11310;
assign n_11312 = ~x_2240 & ~n_11311;
assign n_11313 =  x_2240 & ~n_11310;
assign n_11314 = ~n_11309 &  n_11313;
assign n_11315 =  n_10871 & ~n_11314;
assign n_11316 = ~n_11312 &  n_11315;
assign n_11317 =  x_2672 &  n_10878;
assign n_11318 =  x_4829 &  n_10875;
assign n_11319 = ~n_11317 & ~n_11318;
assign n_11320 = ~n_11316 &  n_11319;
assign n_11321 = ~x_1504 &  n_11276;
assign n_11322 =  x_1504 & ~n_11276;
assign n_11323 = ~n_11321 & ~n_11322;
assign n_11324 = ~n_11280 & ~n_11284;
assign n_11325 =  n_11323 & ~n_11324;
assign n_11326 = ~n_11323 &  n_11324;
assign n_11327 = ~n_11325 & ~n_11326;
assign n_11328 = ~x_4190 & ~n_11327;
assign n_11329 =  x_4190 & ~n_11326;
assign n_11330 = ~n_11325 &  n_11329;
assign n_11331 =  n_10873 & ~n_11330;
assign n_11332 = ~n_11328 &  n_11331;
assign n_11333 = ~x_2016 &  n_11288;
assign n_11334 =  x_2016 & ~n_11288;
assign n_11335 = ~n_11333 & ~n_11334;
assign n_11336 = ~n_11292 & ~n_11296;
assign n_11337 =  n_11335 & ~n_11336;
assign n_11338 = ~n_11335 &  n_11336;
assign n_11339 = ~n_11337 & ~n_11338;
assign n_11340 = ~x_3821 & ~n_11339;
assign n_11341 =  x_3821 & ~n_11338;
assign n_11342 = ~n_11337 &  n_11341;
assign n_11343 =  n_10870 & ~n_11342;
assign n_11344 = ~n_11340 &  n_11343;
assign n_11345 = ~n_11332 & ~n_11344;
assign n_11346 =  n_11320 &  n_11345;
assign n_11347 =  x_2672 & ~n_11346;
assign n_11348 = ~x_2672 &  n_11346;
assign n_11349 = ~n_11347 & ~n_11348;
assign n_11350 = ~x_3756 &  n_11305;
assign n_11351 =  x_3756 & ~n_11305;
assign n_11352 = ~n_11350 & ~n_11351;
assign n_11353 = ~n_11309 & ~n_11313;
assign n_11354 =  n_11352 & ~n_11353;
assign n_11355 = ~n_11352 &  n_11353;
assign n_11356 = ~n_11354 & ~n_11355;
assign n_11357 = ~x_2239 & ~n_11356;
assign n_11358 =  x_2239 & ~n_11355;
assign n_11359 = ~n_11354 &  n_11358;
assign n_11360 =  n_10871 & ~n_11359;
assign n_11361 = ~n_11357 &  n_11360;
assign n_11362 =  x_2671 &  n_10878;
assign n_11363 =  x_4828 &  n_10875;
assign n_11364 = ~n_11362 & ~n_11363;
assign n_11365 = ~n_11361 &  n_11364;
assign n_11366 = ~x_1503 &  n_11321;
assign n_11367 =  x_1503 & ~n_11321;
assign n_11368 = ~n_11366 & ~n_11367;
assign n_11369 = ~n_11325 & ~n_11329;
assign n_11370 =  n_11368 & ~n_11369;
assign n_11371 = ~n_11368 &  n_11369;
assign n_11372 = ~n_11370 & ~n_11371;
assign n_11373 = ~x_4189 & ~n_11372;
assign n_11374 =  x_4189 & ~n_11371;
assign n_11375 = ~n_11370 &  n_11374;
assign n_11376 =  n_10873 & ~n_11375;
assign n_11377 = ~n_11373 &  n_11376;
assign n_11378 = ~x_2015 &  n_11333;
assign n_11379 =  x_2015 & ~n_11333;
assign n_11380 = ~n_11378 & ~n_11379;
assign n_11381 = ~n_11337 & ~n_11341;
assign n_11382 =  n_11380 & ~n_11381;
assign n_11383 = ~n_11380 &  n_11381;
assign n_11384 = ~n_11382 & ~n_11383;
assign n_11385 = ~x_3820 & ~n_11384;
assign n_11386 =  x_3820 & ~n_11383;
assign n_11387 = ~n_11382 &  n_11386;
assign n_11388 =  n_10870 & ~n_11387;
assign n_11389 = ~n_11385 &  n_11388;
assign n_11390 = ~n_11377 & ~n_11389;
assign n_11391 =  n_11365 &  n_11390;
assign n_11392 =  x_2671 & ~n_11391;
assign n_11393 = ~x_2671 &  n_11391;
assign n_11394 = ~n_11392 & ~n_11393;
assign n_11395 = ~x_3755 &  n_11350;
assign n_11396 =  x_3755 & ~n_11350;
assign n_11397 = ~n_11395 & ~n_11396;
assign n_11398 = ~n_11354 & ~n_11358;
assign n_11399 =  n_11397 & ~n_11398;
assign n_11400 = ~n_11397 &  n_11398;
assign n_11401 = ~n_11399 & ~n_11400;
assign n_11402 = ~x_2238 & ~n_11401;
assign n_11403 =  x_2238 & ~n_11400;
assign n_11404 = ~n_11399 &  n_11403;
assign n_11405 =  n_10871 & ~n_11404;
assign n_11406 = ~n_11402 &  n_11405;
assign n_11407 =  x_2670 &  n_10878;
assign n_11408 =  x_4827 &  n_10875;
assign n_11409 = ~n_11407 & ~n_11408;
assign n_11410 = ~n_11406 &  n_11409;
assign n_11411 = ~x_1502 &  n_11366;
assign n_11412 =  x_1502 & ~n_11366;
assign n_11413 = ~n_11411 & ~n_11412;
assign n_11414 = ~n_11370 & ~n_11374;
assign n_11415 =  n_11413 & ~n_11414;
assign n_11416 = ~n_11413 &  n_11414;
assign n_11417 = ~n_11415 & ~n_11416;
assign n_11418 = ~x_4188 & ~n_11417;
assign n_11419 =  x_4188 & ~n_11416;
assign n_11420 = ~n_11415 &  n_11419;
assign n_11421 =  n_10873 & ~n_11420;
assign n_11422 = ~n_11418 &  n_11421;
assign n_11423 = ~x_2014 &  n_11378;
assign n_11424 =  x_2014 & ~n_11378;
assign n_11425 = ~n_11423 & ~n_11424;
assign n_11426 = ~n_11382 & ~n_11386;
assign n_11427 =  n_11425 & ~n_11426;
assign n_11428 = ~n_11425 &  n_11426;
assign n_11429 = ~n_11427 & ~n_11428;
assign n_11430 = ~x_3819 & ~n_11429;
assign n_11431 =  x_3819 & ~n_11428;
assign n_11432 = ~n_11427 &  n_11431;
assign n_11433 =  n_10870 & ~n_11432;
assign n_11434 = ~n_11430 &  n_11433;
assign n_11435 = ~n_11422 & ~n_11434;
assign n_11436 =  n_11410 &  n_11435;
assign n_11437 =  x_2670 & ~n_11436;
assign n_11438 = ~x_2670 &  n_11436;
assign n_11439 = ~n_11437 & ~n_11438;
assign n_11440 = ~x_3754 &  n_11395;
assign n_11441 =  x_3754 & ~n_11395;
assign n_11442 = ~n_11440 & ~n_11441;
assign n_11443 = ~n_11399 & ~n_11403;
assign n_11444 =  n_11442 & ~n_11443;
assign n_11445 = ~n_11442 &  n_11443;
assign n_11446 = ~n_11444 & ~n_11445;
assign n_11447 = ~x_2237 & ~n_11446;
assign n_11448 =  x_2237 & ~n_11445;
assign n_11449 = ~n_11444 &  n_11448;
assign n_11450 =  n_10871 & ~n_11449;
assign n_11451 = ~n_11447 &  n_11450;
assign n_11452 =  x_2669 &  n_10878;
assign n_11453 =  x_4826 &  n_10875;
assign n_11454 = ~n_11452 & ~n_11453;
assign n_11455 = ~n_11451 &  n_11454;
assign n_11456 = ~x_1501 &  n_11411;
assign n_11457 =  x_1501 & ~n_11411;
assign n_11458 = ~n_11456 & ~n_11457;
assign n_11459 = ~n_11415 & ~n_11419;
assign n_11460 =  n_11458 & ~n_11459;
assign n_11461 = ~n_11458 &  n_11459;
assign n_11462 = ~n_11460 & ~n_11461;
assign n_11463 = ~x_4187 & ~n_11462;
assign n_11464 =  x_4187 & ~n_11461;
assign n_11465 = ~n_11460 &  n_11464;
assign n_11466 =  n_10873 & ~n_11465;
assign n_11467 = ~n_11463 &  n_11466;
assign n_11468 = ~x_2013 &  n_11423;
assign n_11469 =  x_2013 & ~n_11423;
assign n_11470 = ~n_11468 & ~n_11469;
assign n_11471 = ~n_11427 & ~n_11431;
assign n_11472 =  n_11470 & ~n_11471;
assign n_11473 = ~n_11470 &  n_11471;
assign n_11474 = ~n_11472 & ~n_11473;
assign n_11475 = ~x_3818 & ~n_11474;
assign n_11476 =  x_3818 & ~n_11473;
assign n_11477 = ~n_11472 &  n_11476;
assign n_11478 =  n_10870 & ~n_11477;
assign n_11479 = ~n_11475 &  n_11478;
assign n_11480 = ~n_11467 & ~n_11479;
assign n_11481 =  n_11455 &  n_11480;
assign n_11482 =  x_2669 & ~n_11481;
assign n_11483 = ~x_2669 &  n_11481;
assign n_11484 = ~n_11482 & ~n_11483;
assign n_11485 = ~x_3753 &  n_11440;
assign n_11486 =  x_3753 & ~n_11440;
assign n_11487 = ~n_11485 & ~n_11486;
assign n_11488 = ~n_11444 & ~n_11448;
assign n_11489 =  n_11487 & ~n_11488;
assign n_11490 = ~n_11487 &  n_11488;
assign n_11491 = ~n_11489 & ~n_11490;
assign n_11492 = ~x_2236 & ~n_11491;
assign n_11493 =  x_2236 & ~n_11490;
assign n_11494 = ~n_11489 &  n_11493;
assign n_11495 =  n_10871 & ~n_11494;
assign n_11496 = ~n_11492 &  n_11495;
assign n_11497 =  x_2668 &  n_10878;
assign n_11498 =  x_4825 &  n_10875;
assign n_11499 = ~n_11497 & ~n_11498;
assign n_11500 = ~n_11496 &  n_11499;
assign n_11501 = ~x_1500 &  n_11456;
assign n_11502 =  x_1500 & ~n_11456;
assign n_11503 = ~n_11501 & ~n_11502;
assign n_11504 = ~n_11460 & ~n_11464;
assign n_11505 =  n_11503 & ~n_11504;
assign n_11506 = ~n_11503 &  n_11504;
assign n_11507 = ~n_11505 & ~n_11506;
assign n_11508 = ~x_4186 & ~n_11507;
assign n_11509 =  x_4186 & ~n_11506;
assign n_11510 = ~n_11505 &  n_11509;
assign n_11511 =  n_10873 & ~n_11510;
assign n_11512 = ~n_11508 &  n_11511;
assign n_11513 = ~x_2012 &  n_11468;
assign n_11514 =  x_2012 & ~n_11468;
assign n_11515 = ~n_11513 & ~n_11514;
assign n_11516 = ~n_11472 & ~n_11476;
assign n_11517 =  n_11515 & ~n_11516;
assign n_11518 = ~n_11515 &  n_11516;
assign n_11519 = ~n_11517 & ~n_11518;
assign n_11520 = ~x_3817 & ~n_11519;
assign n_11521 =  x_3817 & ~n_11518;
assign n_11522 = ~n_11517 &  n_11521;
assign n_11523 =  n_10870 & ~n_11522;
assign n_11524 = ~n_11520 &  n_11523;
assign n_11525 = ~n_11512 & ~n_11524;
assign n_11526 =  n_11500 &  n_11525;
assign n_11527 =  x_2668 & ~n_11526;
assign n_11528 = ~x_2668 &  n_11526;
assign n_11529 = ~n_11527 & ~n_11528;
assign n_11530 = ~x_3752 &  n_11485;
assign n_11531 =  x_3752 & ~n_11485;
assign n_11532 = ~n_11530 & ~n_11531;
assign n_11533 = ~n_11489 & ~n_11493;
assign n_11534 =  n_11532 & ~n_11533;
assign n_11535 = ~n_11532 &  n_11533;
assign n_11536 = ~n_11534 & ~n_11535;
assign n_11537 = ~x_2235 & ~n_11536;
assign n_11538 =  x_2235 & ~n_11535;
assign n_11539 = ~n_11534 &  n_11538;
assign n_11540 =  n_10871 & ~n_11539;
assign n_11541 = ~n_11537 &  n_11540;
assign n_11542 =  x_2667 &  n_10878;
assign n_11543 =  x_4824 &  n_10875;
assign n_11544 = ~n_11542 & ~n_11543;
assign n_11545 = ~n_11541 &  n_11544;
assign n_11546 = ~x_1499 &  n_11501;
assign n_11547 =  x_1499 & ~n_11501;
assign n_11548 = ~n_11546 & ~n_11547;
assign n_11549 = ~n_11505 & ~n_11509;
assign n_11550 =  n_11548 & ~n_11549;
assign n_11551 = ~n_11548 &  n_11549;
assign n_11552 = ~n_11550 & ~n_11551;
assign n_11553 = ~x_4185 & ~n_11552;
assign n_11554 =  x_4185 & ~n_11551;
assign n_11555 = ~n_11550 &  n_11554;
assign n_11556 =  n_10873 & ~n_11555;
assign n_11557 = ~n_11553 &  n_11556;
assign n_11558 = ~x_2011 &  n_11513;
assign n_11559 =  x_2011 & ~n_11513;
assign n_11560 = ~n_11558 & ~n_11559;
assign n_11561 = ~n_11517 & ~n_11521;
assign n_11562 =  n_11560 & ~n_11561;
assign n_11563 = ~n_11560 &  n_11561;
assign n_11564 = ~n_11562 & ~n_11563;
assign n_11565 = ~x_3816 & ~n_11564;
assign n_11566 =  x_3816 & ~n_11563;
assign n_11567 = ~n_11562 &  n_11566;
assign n_11568 =  n_10870 & ~n_11567;
assign n_11569 = ~n_11565 &  n_11568;
assign n_11570 = ~n_11557 & ~n_11569;
assign n_11571 =  n_11545 &  n_11570;
assign n_11572 =  x_2667 & ~n_11571;
assign n_11573 = ~x_2667 &  n_11571;
assign n_11574 = ~n_11572 & ~n_11573;
assign n_11575 = ~x_3751 &  n_11530;
assign n_11576 =  x_3751 & ~n_11530;
assign n_11577 = ~n_11575 & ~n_11576;
assign n_11578 = ~n_11534 & ~n_11538;
assign n_11579 =  n_11577 & ~n_11578;
assign n_11580 = ~n_11577 &  n_11578;
assign n_11581 = ~n_11579 & ~n_11580;
assign n_11582 = ~x_2234 & ~n_11581;
assign n_11583 =  x_2234 & ~n_11580;
assign n_11584 = ~n_11579 &  n_11583;
assign n_11585 =  n_10871 & ~n_11584;
assign n_11586 = ~n_11582 &  n_11585;
assign n_11587 =  x_2666 &  n_10878;
assign n_11588 =  x_4823 &  n_10875;
assign n_11589 = ~n_11587 & ~n_11588;
assign n_11590 = ~n_11586 &  n_11589;
assign n_11591 = ~x_1498 &  n_11546;
assign n_11592 =  x_1498 & ~n_11546;
assign n_11593 = ~n_11591 & ~n_11592;
assign n_11594 = ~n_11550 & ~n_11554;
assign n_11595 =  n_11593 & ~n_11594;
assign n_11596 = ~n_11593 &  n_11594;
assign n_11597 = ~n_11595 & ~n_11596;
assign n_11598 = ~x_4184 & ~n_11597;
assign n_11599 =  x_4184 & ~n_11596;
assign n_11600 = ~n_11595 &  n_11599;
assign n_11601 =  n_10873 & ~n_11600;
assign n_11602 = ~n_11598 &  n_11601;
assign n_11603 = ~x_2010 &  n_11558;
assign n_11604 =  x_2010 & ~n_11558;
assign n_11605 = ~n_11603 & ~n_11604;
assign n_11606 = ~n_11562 & ~n_11566;
assign n_11607 =  n_11605 & ~n_11606;
assign n_11608 = ~n_11605 &  n_11606;
assign n_11609 = ~n_11607 & ~n_11608;
assign n_11610 = ~x_3815 & ~n_11609;
assign n_11611 =  x_3815 & ~n_11608;
assign n_11612 = ~n_11607 &  n_11611;
assign n_11613 =  n_10870 & ~n_11612;
assign n_11614 = ~n_11610 &  n_11613;
assign n_11615 = ~n_11602 & ~n_11614;
assign n_11616 =  n_11590 &  n_11615;
assign n_11617 =  x_2666 & ~n_11616;
assign n_11618 = ~x_2666 &  n_11616;
assign n_11619 = ~n_11617 & ~n_11618;
assign n_11620 = ~x_3750 &  n_11575;
assign n_11621 =  x_3750 & ~n_11575;
assign n_11622 = ~n_11620 & ~n_11621;
assign n_11623 = ~n_11579 & ~n_11583;
assign n_11624 =  n_11622 & ~n_11623;
assign n_11625 = ~n_11622 &  n_11623;
assign n_11626 = ~n_11624 & ~n_11625;
assign n_11627 = ~x_2233 & ~n_11626;
assign n_11628 =  x_2233 & ~n_11625;
assign n_11629 = ~n_11624 &  n_11628;
assign n_11630 =  n_10871 & ~n_11629;
assign n_11631 = ~n_11627 &  n_11630;
assign n_11632 =  x_2665 &  n_10878;
assign n_11633 =  x_4822 &  n_10875;
assign n_11634 = ~n_11632 & ~n_11633;
assign n_11635 = ~n_11631 &  n_11634;
assign n_11636 = ~x_1497 &  n_11591;
assign n_11637 =  x_1497 & ~n_11591;
assign n_11638 = ~n_11636 & ~n_11637;
assign n_11639 = ~n_11595 & ~n_11599;
assign n_11640 =  n_11638 & ~n_11639;
assign n_11641 = ~n_11638 &  n_11639;
assign n_11642 = ~n_11640 & ~n_11641;
assign n_11643 = ~x_4183 & ~n_11642;
assign n_11644 =  x_4183 & ~n_11641;
assign n_11645 = ~n_11640 &  n_11644;
assign n_11646 =  n_10873 & ~n_11645;
assign n_11647 = ~n_11643 &  n_11646;
assign n_11648 = ~x_2009 &  n_11603;
assign n_11649 =  x_2009 & ~n_11603;
assign n_11650 = ~n_11648 & ~n_11649;
assign n_11651 = ~n_11607 & ~n_11611;
assign n_11652 =  n_11650 & ~n_11651;
assign n_11653 = ~n_11650 &  n_11651;
assign n_11654 = ~n_11652 & ~n_11653;
assign n_11655 = ~x_3814 & ~n_11654;
assign n_11656 =  x_3814 & ~n_11653;
assign n_11657 = ~n_11652 &  n_11656;
assign n_11658 =  n_10870 & ~n_11657;
assign n_11659 = ~n_11655 &  n_11658;
assign n_11660 = ~n_11647 & ~n_11659;
assign n_11661 =  n_11635 &  n_11660;
assign n_11662 =  x_2665 & ~n_11661;
assign n_11663 = ~x_2665 &  n_11661;
assign n_11664 = ~n_11662 & ~n_11663;
assign n_11665 = ~x_3749 &  n_11620;
assign n_11666 =  x_3749 & ~n_11620;
assign n_11667 = ~n_11665 & ~n_11666;
assign n_11668 = ~n_11624 & ~n_11628;
assign n_11669 =  n_11667 & ~n_11668;
assign n_11670 = ~n_11667 &  n_11668;
assign n_11671 = ~n_11669 & ~n_11670;
assign n_11672 = ~x_2232 & ~n_11671;
assign n_11673 =  x_2232 & ~n_11670;
assign n_11674 = ~n_11669 &  n_11673;
assign n_11675 =  n_10871 & ~n_11674;
assign n_11676 = ~n_11672 &  n_11675;
assign n_11677 =  x_2664 &  n_10878;
assign n_11678 =  x_4821 &  n_10875;
assign n_11679 = ~n_11677 & ~n_11678;
assign n_11680 = ~n_11676 &  n_11679;
assign n_11681 = ~x_1496 &  n_11636;
assign n_11682 =  x_1496 & ~n_11636;
assign n_11683 = ~n_11681 & ~n_11682;
assign n_11684 = ~n_11640 & ~n_11644;
assign n_11685 =  n_11683 & ~n_11684;
assign n_11686 = ~n_11683 &  n_11684;
assign n_11687 = ~n_11685 & ~n_11686;
assign n_11688 = ~x_4182 & ~n_11687;
assign n_11689 =  x_4182 & ~n_11686;
assign n_11690 = ~n_11685 &  n_11689;
assign n_11691 =  n_10873 & ~n_11690;
assign n_11692 = ~n_11688 &  n_11691;
assign n_11693 = ~x_2008 &  n_11648;
assign n_11694 =  x_2008 & ~n_11648;
assign n_11695 = ~n_11693 & ~n_11694;
assign n_11696 = ~n_11652 & ~n_11656;
assign n_11697 =  n_11695 & ~n_11696;
assign n_11698 = ~n_11695 &  n_11696;
assign n_11699 = ~n_11697 & ~n_11698;
assign n_11700 = ~x_3813 & ~n_11699;
assign n_11701 =  x_3813 & ~n_11698;
assign n_11702 = ~n_11697 &  n_11701;
assign n_11703 =  n_10870 & ~n_11702;
assign n_11704 = ~n_11700 &  n_11703;
assign n_11705 = ~n_11692 & ~n_11704;
assign n_11706 =  n_11680 &  n_11705;
assign n_11707 =  x_2664 & ~n_11706;
assign n_11708 = ~x_2664 &  n_11706;
assign n_11709 = ~n_11707 & ~n_11708;
assign n_11710 = ~x_3748 &  n_11665;
assign n_11711 =  x_3748 & ~n_11665;
assign n_11712 = ~n_11710 & ~n_11711;
assign n_11713 = ~n_11669 & ~n_11673;
assign n_11714 =  n_11712 & ~n_11713;
assign n_11715 = ~n_11712 &  n_11713;
assign n_11716 = ~n_11714 & ~n_11715;
assign n_11717 = ~x_2231 & ~n_11716;
assign n_11718 =  x_2231 & ~n_11715;
assign n_11719 = ~n_11714 &  n_11718;
assign n_11720 =  n_10871 & ~n_11719;
assign n_11721 = ~n_11717 &  n_11720;
assign n_11722 =  x_2663 &  n_10878;
assign n_11723 =  x_4820 &  n_10875;
assign n_11724 = ~n_11722 & ~n_11723;
assign n_11725 = ~n_11721 &  n_11724;
assign n_11726 = ~x_1495 &  n_11681;
assign n_11727 =  x_1495 & ~n_11681;
assign n_11728 = ~n_11726 & ~n_11727;
assign n_11729 = ~n_11685 & ~n_11689;
assign n_11730 =  n_11728 & ~n_11729;
assign n_11731 = ~n_11728 &  n_11729;
assign n_11732 = ~n_11730 & ~n_11731;
assign n_11733 = ~x_4181 & ~n_11732;
assign n_11734 =  x_4181 & ~n_11731;
assign n_11735 = ~n_11730 &  n_11734;
assign n_11736 =  n_10873 & ~n_11735;
assign n_11737 = ~n_11733 &  n_11736;
assign n_11738 = ~x_2007 &  n_11693;
assign n_11739 =  x_2007 & ~n_11693;
assign n_11740 = ~n_11738 & ~n_11739;
assign n_11741 = ~n_11697 & ~n_11701;
assign n_11742 =  n_11740 & ~n_11741;
assign n_11743 = ~n_11740 &  n_11741;
assign n_11744 = ~n_11742 & ~n_11743;
assign n_11745 = ~x_3812 & ~n_11744;
assign n_11746 =  x_3812 & ~n_11743;
assign n_11747 = ~n_11742 &  n_11746;
assign n_11748 =  n_10870 & ~n_11747;
assign n_11749 = ~n_11745 &  n_11748;
assign n_11750 = ~n_11737 & ~n_11749;
assign n_11751 =  n_11725 &  n_11750;
assign n_11752 =  x_2663 & ~n_11751;
assign n_11753 = ~x_2663 &  n_11751;
assign n_11754 = ~n_11752 & ~n_11753;
assign n_11755 = ~x_3747 &  n_11710;
assign n_11756 =  x_3747 & ~n_11710;
assign n_11757 = ~n_11755 & ~n_11756;
assign n_11758 = ~n_11714 & ~n_11718;
assign n_11759 =  n_11757 & ~n_11758;
assign n_11760 = ~n_11757 &  n_11758;
assign n_11761 = ~n_11759 & ~n_11760;
assign n_11762 = ~x_2230 & ~n_11761;
assign n_11763 =  x_2230 & ~n_11760;
assign n_11764 = ~n_11759 &  n_11763;
assign n_11765 =  n_10871 & ~n_11764;
assign n_11766 = ~n_11762 &  n_11765;
assign n_11767 =  x_2662 &  n_10878;
assign n_11768 =  x_4819 &  n_10875;
assign n_11769 = ~n_11767 & ~n_11768;
assign n_11770 = ~n_11766 &  n_11769;
assign n_11771 = ~x_1494 &  n_11726;
assign n_11772 =  x_1494 & ~n_11726;
assign n_11773 = ~n_11771 & ~n_11772;
assign n_11774 = ~n_11730 & ~n_11734;
assign n_11775 =  n_11773 & ~n_11774;
assign n_11776 = ~n_11773 &  n_11774;
assign n_11777 = ~n_11775 & ~n_11776;
assign n_11778 = ~x_4180 & ~n_11777;
assign n_11779 =  x_4180 & ~n_11776;
assign n_11780 = ~n_11775 &  n_11779;
assign n_11781 =  n_10873 & ~n_11780;
assign n_11782 = ~n_11778 &  n_11781;
assign n_11783 = ~x_2006 &  n_11738;
assign n_11784 =  x_2006 & ~n_11738;
assign n_11785 = ~n_11783 & ~n_11784;
assign n_11786 = ~n_11742 & ~n_11746;
assign n_11787 =  n_11785 & ~n_11786;
assign n_11788 = ~n_11785 &  n_11786;
assign n_11789 = ~n_11787 & ~n_11788;
assign n_11790 = ~x_3811 & ~n_11789;
assign n_11791 =  x_3811 & ~n_11788;
assign n_11792 = ~n_11787 &  n_11791;
assign n_11793 =  n_10870 & ~n_11792;
assign n_11794 = ~n_11790 &  n_11793;
assign n_11795 = ~n_11782 & ~n_11794;
assign n_11796 =  n_11770 &  n_11795;
assign n_11797 =  x_2662 & ~n_11796;
assign n_11798 = ~x_2662 &  n_11796;
assign n_11799 = ~n_11797 & ~n_11798;
assign n_11800 = ~x_3746 &  n_11755;
assign n_11801 =  x_3746 & ~n_11755;
assign n_11802 = ~n_11800 & ~n_11801;
assign n_11803 = ~n_11759 & ~n_11763;
assign n_11804 =  n_11802 & ~n_11803;
assign n_11805 = ~n_11802 &  n_11803;
assign n_11806 = ~n_11804 & ~n_11805;
assign n_11807 = ~x_2229 & ~n_11806;
assign n_11808 =  x_2229 & ~n_11805;
assign n_11809 = ~n_11804 &  n_11808;
assign n_11810 =  n_10871 & ~n_11809;
assign n_11811 = ~n_11807 &  n_11810;
assign n_11812 =  x_2661 &  n_10878;
assign n_11813 =  x_4818 &  n_10875;
assign n_11814 = ~n_11812 & ~n_11813;
assign n_11815 = ~n_11811 &  n_11814;
assign n_11816 = ~x_1493 &  n_11771;
assign n_11817 =  x_1493 & ~n_11771;
assign n_11818 = ~n_11816 & ~n_11817;
assign n_11819 = ~n_11775 & ~n_11779;
assign n_11820 =  n_11818 & ~n_11819;
assign n_11821 = ~n_11818 &  n_11819;
assign n_11822 = ~n_11820 & ~n_11821;
assign n_11823 = ~x_4179 & ~n_11822;
assign n_11824 =  x_4179 & ~n_11821;
assign n_11825 = ~n_11820 &  n_11824;
assign n_11826 =  n_10873 & ~n_11825;
assign n_11827 = ~n_11823 &  n_11826;
assign n_11828 = ~x_2005 &  n_11783;
assign n_11829 =  x_2005 & ~n_11783;
assign n_11830 = ~n_11828 & ~n_11829;
assign n_11831 = ~n_11787 & ~n_11791;
assign n_11832 =  n_11830 & ~n_11831;
assign n_11833 = ~n_11830 &  n_11831;
assign n_11834 = ~n_11832 & ~n_11833;
assign n_11835 = ~x_3810 & ~n_11834;
assign n_11836 =  x_3810 & ~n_11833;
assign n_11837 = ~n_11832 &  n_11836;
assign n_11838 =  n_10870 & ~n_11837;
assign n_11839 = ~n_11835 &  n_11838;
assign n_11840 = ~n_11827 & ~n_11839;
assign n_11841 =  n_11815 &  n_11840;
assign n_11842 =  x_2661 & ~n_11841;
assign n_11843 = ~x_2661 &  n_11841;
assign n_11844 = ~n_11842 & ~n_11843;
assign n_11845 = ~x_3745 &  n_11800;
assign n_11846 =  x_3745 & ~n_11800;
assign n_11847 = ~n_11845 & ~n_11846;
assign n_11848 = ~n_11804 & ~n_11808;
assign n_11849 =  n_11847 & ~n_11848;
assign n_11850 = ~n_11847 &  n_11848;
assign n_11851 = ~n_11849 & ~n_11850;
assign n_11852 = ~x_2228 & ~n_11851;
assign n_11853 =  x_2228 & ~n_11850;
assign n_11854 = ~n_11849 &  n_11853;
assign n_11855 =  n_10871 & ~n_11854;
assign n_11856 = ~n_11852 &  n_11855;
assign n_11857 =  x_2660 &  n_10878;
assign n_11858 =  x_4817 &  n_10875;
assign n_11859 = ~n_11857 & ~n_11858;
assign n_11860 = ~n_11856 &  n_11859;
assign n_11861 = ~x_1492 &  n_11816;
assign n_11862 =  x_1492 & ~n_11816;
assign n_11863 = ~n_11861 & ~n_11862;
assign n_11864 = ~n_11820 & ~n_11824;
assign n_11865 =  n_11863 & ~n_11864;
assign n_11866 = ~n_11863 &  n_11864;
assign n_11867 = ~n_11865 & ~n_11866;
assign n_11868 = ~x_4178 & ~n_11867;
assign n_11869 =  x_4178 & ~n_11866;
assign n_11870 = ~n_11865 &  n_11869;
assign n_11871 =  n_10873 & ~n_11870;
assign n_11872 = ~n_11868 &  n_11871;
assign n_11873 = ~x_2004 &  n_11828;
assign n_11874 =  x_2004 & ~n_11828;
assign n_11875 = ~n_11873 & ~n_11874;
assign n_11876 = ~n_11832 & ~n_11836;
assign n_11877 =  n_11875 & ~n_11876;
assign n_11878 = ~n_11875 &  n_11876;
assign n_11879 = ~n_11877 & ~n_11878;
assign n_11880 = ~x_3809 & ~n_11879;
assign n_11881 =  x_3809 & ~n_11878;
assign n_11882 = ~n_11877 &  n_11881;
assign n_11883 =  n_10870 & ~n_11882;
assign n_11884 = ~n_11880 &  n_11883;
assign n_11885 = ~n_11872 & ~n_11884;
assign n_11886 =  n_11860 &  n_11885;
assign n_11887 =  x_2660 & ~n_11886;
assign n_11888 = ~x_2660 &  n_11886;
assign n_11889 = ~n_11887 & ~n_11888;
assign n_11890 = ~x_3744 &  n_11845;
assign n_11891 =  x_3744 & ~n_11845;
assign n_11892 = ~n_11890 & ~n_11891;
assign n_11893 = ~n_11849 & ~n_11853;
assign n_11894 =  n_11892 & ~n_11893;
assign n_11895 = ~n_11892 &  n_11893;
assign n_11896 = ~n_11894 & ~n_11895;
assign n_11897 = ~x_2227 & ~n_11896;
assign n_11898 =  x_2227 & ~n_11895;
assign n_11899 = ~n_11894 &  n_11898;
assign n_11900 =  n_10871 & ~n_11899;
assign n_11901 = ~n_11897 &  n_11900;
assign n_11902 =  x_2659 &  n_10878;
assign n_11903 =  x_4816 &  n_10875;
assign n_11904 = ~n_11902 & ~n_11903;
assign n_11905 = ~n_11901 &  n_11904;
assign n_11906 = ~x_1491 &  n_11861;
assign n_11907 =  x_1491 & ~n_11861;
assign n_11908 = ~n_11906 & ~n_11907;
assign n_11909 = ~n_11865 & ~n_11869;
assign n_11910 =  n_11908 & ~n_11909;
assign n_11911 = ~n_11908 &  n_11909;
assign n_11912 = ~n_11910 & ~n_11911;
assign n_11913 = ~x_4177 & ~n_11912;
assign n_11914 =  x_4177 & ~n_11911;
assign n_11915 = ~n_11910 &  n_11914;
assign n_11916 =  n_10873 & ~n_11915;
assign n_11917 = ~n_11913 &  n_11916;
assign n_11918 = ~x_2003 &  n_11873;
assign n_11919 =  x_2003 & ~n_11873;
assign n_11920 = ~n_11918 & ~n_11919;
assign n_11921 = ~n_11877 & ~n_11881;
assign n_11922 =  n_11920 & ~n_11921;
assign n_11923 = ~n_11920 &  n_11921;
assign n_11924 = ~n_11922 & ~n_11923;
assign n_11925 = ~x_3808 & ~n_11924;
assign n_11926 =  x_3808 & ~n_11923;
assign n_11927 = ~n_11922 &  n_11926;
assign n_11928 =  n_10870 & ~n_11927;
assign n_11929 = ~n_11925 &  n_11928;
assign n_11930 = ~n_11917 & ~n_11929;
assign n_11931 =  n_11905 &  n_11930;
assign n_11932 =  x_2659 & ~n_11931;
assign n_11933 = ~x_2659 &  n_11931;
assign n_11934 = ~n_11932 & ~n_11933;
assign n_11935 = ~x_3743 &  n_11890;
assign n_11936 =  x_3743 & ~n_11890;
assign n_11937 = ~n_11935 & ~n_11936;
assign n_11938 = ~n_11894 & ~n_11898;
assign n_11939 =  n_11937 & ~n_11938;
assign n_11940 = ~n_11937 &  n_11938;
assign n_11941 = ~n_11939 & ~n_11940;
assign n_11942 = ~x_2226 & ~n_11941;
assign n_11943 =  x_2226 & ~n_11940;
assign n_11944 = ~n_11939 &  n_11943;
assign n_11945 =  n_10871 & ~n_11944;
assign n_11946 = ~n_11942 &  n_11945;
assign n_11947 =  x_2658 &  n_10878;
assign n_11948 =  x_4815 &  n_10875;
assign n_11949 = ~n_11947 & ~n_11948;
assign n_11950 = ~n_11946 &  n_11949;
assign n_11951 = ~x_1490 &  n_11906;
assign n_11952 =  x_1490 & ~n_11906;
assign n_11953 = ~n_11951 & ~n_11952;
assign n_11954 = ~n_11910 & ~n_11914;
assign n_11955 =  n_11953 & ~n_11954;
assign n_11956 = ~n_11953 &  n_11954;
assign n_11957 = ~n_11955 & ~n_11956;
assign n_11958 = ~x_4176 & ~n_11957;
assign n_11959 =  x_4176 & ~n_11956;
assign n_11960 = ~n_11955 &  n_11959;
assign n_11961 =  n_10873 & ~n_11960;
assign n_11962 = ~n_11958 &  n_11961;
assign n_11963 = ~x_2002 &  n_11918;
assign n_11964 =  x_2002 & ~n_11918;
assign n_11965 = ~n_11963 & ~n_11964;
assign n_11966 = ~n_11922 & ~n_11926;
assign n_11967 =  n_11965 & ~n_11966;
assign n_11968 = ~n_11965 &  n_11966;
assign n_11969 = ~n_11967 & ~n_11968;
assign n_11970 = ~x_3807 & ~n_11969;
assign n_11971 =  x_3807 & ~n_11968;
assign n_11972 = ~n_11967 &  n_11971;
assign n_11973 =  n_10870 & ~n_11972;
assign n_11974 = ~n_11970 &  n_11973;
assign n_11975 = ~n_11962 & ~n_11974;
assign n_11976 =  n_11950 &  n_11975;
assign n_11977 =  x_2658 & ~n_11976;
assign n_11978 = ~x_2658 &  n_11976;
assign n_11979 = ~n_11977 & ~n_11978;
assign n_11980 = ~x_3742 &  n_11935;
assign n_11981 =  x_3742 & ~n_11935;
assign n_11982 = ~n_11980 & ~n_11981;
assign n_11983 = ~n_11939 & ~n_11943;
assign n_11984 =  n_11982 & ~n_11983;
assign n_11985 = ~n_11982 &  n_11983;
assign n_11986 = ~n_11984 & ~n_11985;
assign n_11987 = ~x_2225 & ~n_11986;
assign n_11988 =  x_2225 & ~n_11985;
assign n_11989 = ~n_11984 &  n_11988;
assign n_11990 =  n_10871 & ~n_11989;
assign n_11991 = ~n_11987 &  n_11990;
assign n_11992 =  x_2657 &  n_10878;
assign n_11993 =  x_4814 &  n_10875;
assign n_11994 = ~n_11992 & ~n_11993;
assign n_11995 = ~n_11991 &  n_11994;
assign n_11996 = ~x_1489 &  n_11951;
assign n_11997 =  x_1489 & ~n_11951;
assign n_11998 = ~n_11996 & ~n_11997;
assign n_11999 = ~n_11955 & ~n_11959;
assign n_12000 =  n_11998 & ~n_11999;
assign n_12001 = ~n_11998 &  n_11999;
assign n_12002 = ~n_12000 & ~n_12001;
assign n_12003 = ~x_4175 & ~n_12002;
assign n_12004 =  x_4175 & ~n_12001;
assign n_12005 = ~n_12000 &  n_12004;
assign n_12006 =  n_10873 & ~n_12005;
assign n_12007 = ~n_12003 &  n_12006;
assign n_12008 = ~x_2001 &  n_11963;
assign n_12009 =  x_2001 & ~n_11963;
assign n_12010 = ~n_12008 & ~n_12009;
assign n_12011 = ~n_11967 & ~n_11971;
assign n_12012 =  n_12010 & ~n_12011;
assign n_12013 = ~n_12010 &  n_12011;
assign n_12014 = ~n_12012 & ~n_12013;
assign n_12015 = ~x_3806 & ~n_12014;
assign n_12016 =  x_3806 & ~n_12013;
assign n_12017 = ~n_12012 &  n_12016;
assign n_12018 =  n_10870 & ~n_12017;
assign n_12019 = ~n_12015 &  n_12018;
assign n_12020 = ~n_12007 & ~n_12019;
assign n_12021 =  n_11995 &  n_12020;
assign n_12022 =  x_2657 & ~n_12021;
assign n_12023 = ~x_2657 &  n_12021;
assign n_12024 = ~n_12022 & ~n_12023;
assign n_12025 = ~x_3741 &  n_11980;
assign n_12026 =  x_3741 & ~n_11980;
assign n_12027 = ~n_12025 & ~n_12026;
assign n_12028 = ~n_11984 & ~n_11988;
assign n_12029 =  n_12027 & ~n_12028;
assign n_12030 = ~n_12027 &  n_12028;
assign n_12031 = ~n_12029 & ~n_12030;
assign n_12032 = ~x_2224 & ~n_12031;
assign n_12033 =  x_2224 & ~n_12030;
assign n_12034 = ~n_12029 &  n_12033;
assign n_12035 =  n_10871 & ~n_12034;
assign n_12036 = ~n_12032 &  n_12035;
assign n_12037 =  x_2656 &  n_10878;
assign n_12038 =  x_4813 &  n_10875;
assign n_12039 = ~n_12037 & ~n_12038;
assign n_12040 = ~n_12036 &  n_12039;
assign n_12041 = ~x_1488 &  n_11996;
assign n_12042 =  x_1488 & ~n_11996;
assign n_12043 = ~n_12041 & ~n_12042;
assign n_12044 = ~n_12000 & ~n_12004;
assign n_12045 =  n_12043 & ~n_12044;
assign n_12046 = ~n_12043 &  n_12044;
assign n_12047 = ~n_12045 & ~n_12046;
assign n_12048 = ~x_4174 & ~n_12047;
assign n_12049 =  x_4174 & ~n_12046;
assign n_12050 = ~n_12045 &  n_12049;
assign n_12051 =  n_10873 & ~n_12050;
assign n_12052 = ~n_12048 &  n_12051;
assign n_12053 = ~x_2000 &  n_12008;
assign n_12054 =  x_2000 & ~n_12008;
assign n_12055 = ~n_12053 & ~n_12054;
assign n_12056 = ~n_12012 & ~n_12016;
assign n_12057 =  n_12055 & ~n_12056;
assign n_12058 = ~n_12055 &  n_12056;
assign n_12059 = ~n_12057 & ~n_12058;
assign n_12060 = ~x_3805 & ~n_12059;
assign n_12061 =  x_3805 & ~n_12058;
assign n_12062 = ~n_12057 &  n_12061;
assign n_12063 =  n_10870 & ~n_12062;
assign n_12064 = ~n_12060 &  n_12063;
assign n_12065 = ~n_12052 & ~n_12064;
assign n_12066 =  n_12040 &  n_12065;
assign n_12067 =  x_2656 & ~n_12066;
assign n_12068 = ~x_2656 &  n_12066;
assign n_12069 = ~n_12067 & ~n_12068;
assign n_12070 = ~x_3740 &  n_12025;
assign n_12071 =  x_3740 & ~n_12025;
assign n_12072 = ~n_12070 & ~n_12071;
assign n_12073 = ~n_12029 & ~n_12033;
assign n_12074 =  n_12072 & ~n_12073;
assign n_12075 = ~n_12072 &  n_12073;
assign n_12076 = ~n_12074 & ~n_12075;
assign n_12077 = ~x_2223 & ~n_12076;
assign n_12078 =  x_2223 & ~n_12075;
assign n_12079 = ~n_12074 &  n_12078;
assign n_12080 =  n_10871 & ~n_12079;
assign n_12081 = ~n_12077 &  n_12080;
assign n_12082 =  x_2655 &  n_10878;
assign n_12083 =  x_4812 &  n_10875;
assign n_12084 = ~n_12082 & ~n_12083;
assign n_12085 = ~n_12081 &  n_12084;
assign n_12086 = ~x_1487 &  n_12041;
assign n_12087 =  x_1487 & ~n_12041;
assign n_12088 = ~n_12086 & ~n_12087;
assign n_12089 = ~n_12045 & ~n_12049;
assign n_12090 =  n_12088 & ~n_12089;
assign n_12091 = ~n_12088 &  n_12089;
assign n_12092 = ~n_12090 & ~n_12091;
assign n_12093 = ~x_4173 & ~n_12092;
assign n_12094 =  x_4173 & ~n_12091;
assign n_12095 = ~n_12090 &  n_12094;
assign n_12096 =  n_10873 & ~n_12095;
assign n_12097 = ~n_12093 &  n_12096;
assign n_12098 = ~x_1999 &  n_12053;
assign n_12099 =  x_1999 & ~n_12053;
assign n_12100 = ~n_12098 & ~n_12099;
assign n_12101 = ~n_12057 & ~n_12061;
assign n_12102 =  n_12100 & ~n_12101;
assign n_12103 = ~n_12100 &  n_12101;
assign n_12104 = ~n_12102 & ~n_12103;
assign n_12105 = ~x_3804 & ~n_12104;
assign n_12106 =  x_3804 & ~n_12103;
assign n_12107 = ~n_12102 &  n_12106;
assign n_12108 =  n_10870 & ~n_12107;
assign n_12109 = ~n_12105 &  n_12108;
assign n_12110 = ~n_12097 & ~n_12109;
assign n_12111 =  n_12085 &  n_12110;
assign n_12112 =  x_2655 & ~n_12111;
assign n_12113 = ~x_2655 &  n_12111;
assign n_12114 = ~n_12112 & ~n_12113;
assign n_12115 = ~x_3739 &  n_12070;
assign n_12116 =  x_3739 & ~n_12070;
assign n_12117 = ~n_12115 & ~n_12116;
assign n_12118 = ~n_12074 & ~n_12078;
assign n_12119 =  n_12117 & ~n_12118;
assign n_12120 = ~n_12117 &  n_12118;
assign n_12121 = ~n_12119 & ~n_12120;
assign n_12122 = ~x_2222 & ~n_12121;
assign n_12123 =  x_2222 & ~n_12120;
assign n_12124 = ~n_12119 &  n_12123;
assign n_12125 =  n_10871 & ~n_12124;
assign n_12126 = ~n_12122 &  n_12125;
assign n_12127 =  x_2654 &  n_10878;
assign n_12128 =  x_4811 &  n_10875;
assign n_12129 = ~n_12127 & ~n_12128;
assign n_12130 = ~n_12126 &  n_12129;
assign n_12131 = ~x_1486 &  n_12086;
assign n_12132 =  x_1486 & ~n_12086;
assign n_12133 = ~n_12131 & ~n_12132;
assign n_12134 = ~n_12090 & ~n_12094;
assign n_12135 =  n_12133 & ~n_12134;
assign n_12136 = ~n_12133 &  n_12134;
assign n_12137 = ~n_12135 & ~n_12136;
assign n_12138 = ~x_4172 & ~n_12137;
assign n_12139 =  x_4172 & ~n_12136;
assign n_12140 = ~n_12135 &  n_12139;
assign n_12141 =  n_10873 & ~n_12140;
assign n_12142 = ~n_12138 &  n_12141;
assign n_12143 = ~x_1998 &  n_12098;
assign n_12144 =  x_1998 & ~n_12098;
assign n_12145 = ~n_12143 & ~n_12144;
assign n_12146 = ~n_12102 & ~n_12106;
assign n_12147 =  n_12145 & ~n_12146;
assign n_12148 = ~n_12145 &  n_12146;
assign n_12149 = ~n_12147 & ~n_12148;
assign n_12150 = ~x_3803 & ~n_12149;
assign n_12151 =  x_3803 & ~n_12148;
assign n_12152 = ~n_12147 &  n_12151;
assign n_12153 =  n_10870 & ~n_12152;
assign n_12154 = ~n_12150 &  n_12153;
assign n_12155 = ~n_12142 & ~n_12154;
assign n_12156 =  n_12130 &  n_12155;
assign n_12157 =  x_2654 & ~n_12156;
assign n_12158 = ~x_2654 &  n_12156;
assign n_12159 = ~n_12157 & ~n_12158;
assign n_12160 = ~x_3738 &  n_12115;
assign n_12161 =  x_3738 & ~n_12115;
assign n_12162 = ~n_12160 & ~n_12161;
assign n_12163 = ~n_12119 & ~n_12123;
assign n_12164 =  n_12162 & ~n_12163;
assign n_12165 = ~n_12162 &  n_12163;
assign n_12166 = ~n_12164 & ~n_12165;
assign n_12167 = ~x_2221 & ~n_12166;
assign n_12168 =  x_2221 & ~n_12165;
assign n_12169 = ~n_12164 &  n_12168;
assign n_12170 =  n_10871 & ~n_12169;
assign n_12171 = ~n_12167 &  n_12170;
assign n_12172 =  x_2653 &  n_10878;
assign n_12173 =  x_4810 &  n_10875;
assign n_12174 = ~n_12172 & ~n_12173;
assign n_12175 = ~n_12171 &  n_12174;
assign n_12176 = ~x_1485 &  n_12131;
assign n_12177 =  x_1485 & ~n_12131;
assign n_12178 = ~n_12176 & ~n_12177;
assign n_12179 = ~n_12135 & ~n_12139;
assign n_12180 =  n_12178 & ~n_12179;
assign n_12181 = ~n_12178 &  n_12179;
assign n_12182 = ~n_12180 & ~n_12181;
assign n_12183 = ~x_4171 & ~n_12182;
assign n_12184 =  x_4171 & ~n_12181;
assign n_12185 = ~n_12180 &  n_12184;
assign n_12186 =  n_10873 & ~n_12185;
assign n_12187 = ~n_12183 &  n_12186;
assign n_12188 = ~x_1997 &  n_12143;
assign n_12189 =  x_1997 & ~n_12143;
assign n_12190 = ~n_12188 & ~n_12189;
assign n_12191 = ~n_12147 & ~n_12151;
assign n_12192 =  n_12190 & ~n_12191;
assign n_12193 = ~n_12190 &  n_12191;
assign n_12194 = ~n_12192 & ~n_12193;
assign n_12195 = ~x_3802 & ~n_12194;
assign n_12196 =  x_3802 & ~n_12193;
assign n_12197 = ~n_12192 &  n_12196;
assign n_12198 =  n_10870 & ~n_12197;
assign n_12199 = ~n_12195 &  n_12198;
assign n_12200 = ~n_12187 & ~n_12199;
assign n_12201 =  n_12175 &  n_12200;
assign n_12202 =  x_2653 & ~n_12201;
assign n_12203 = ~x_2653 &  n_12201;
assign n_12204 = ~n_12202 & ~n_12203;
assign n_12205 = ~x_3737 &  n_12160;
assign n_12206 =  x_3737 & ~n_12160;
assign n_12207 = ~n_12205 & ~n_12206;
assign n_12208 = ~n_12164 & ~n_12168;
assign n_12209 =  n_12207 & ~n_12208;
assign n_12210 = ~n_12207 &  n_12208;
assign n_12211 = ~n_12209 & ~n_12210;
assign n_12212 = ~x_2220 & ~n_12211;
assign n_12213 =  x_2220 & ~n_12210;
assign n_12214 = ~n_12209 &  n_12213;
assign n_12215 =  n_10871 & ~n_12214;
assign n_12216 = ~n_12212 &  n_12215;
assign n_12217 =  x_2652 &  n_10878;
assign n_12218 =  x_4809 &  n_10875;
assign n_12219 = ~n_12217 & ~n_12218;
assign n_12220 = ~n_12216 &  n_12219;
assign n_12221 = ~x_1484 &  n_12176;
assign n_12222 =  x_1484 & ~n_12176;
assign n_12223 = ~n_12221 & ~n_12222;
assign n_12224 = ~n_12180 & ~n_12184;
assign n_12225 =  n_12223 & ~n_12224;
assign n_12226 = ~n_12223 &  n_12224;
assign n_12227 = ~n_12225 & ~n_12226;
assign n_12228 = ~x_4170 & ~n_12227;
assign n_12229 =  x_4170 & ~n_12226;
assign n_12230 = ~n_12225 &  n_12229;
assign n_12231 =  n_10873 & ~n_12230;
assign n_12232 = ~n_12228 &  n_12231;
assign n_12233 = ~x_1996 &  n_12188;
assign n_12234 =  x_1996 & ~n_12188;
assign n_12235 = ~n_12233 & ~n_12234;
assign n_12236 = ~n_12192 & ~n_12196;
assign n_12237 =  n_12235 & ~n_12236;
assign n_12238 = ~n_12235 &  n_12236;
assign n_12239 = ~n_12237 & ~n_12238;
assign n_12240 = ~x_3801 & ~n_12239;
assign n_12241 =  x_3801 & ~n_12238;
assign n_12242 = ~n_12237 &  n_12241;
assign n_12243 =  n_10870 & ~n_12242;
assign n_12244 = ~n_12240 &  n_12243;
assign n_12245 = ~n_12232 & ~n_12244;
assign n_12246 =  n_12220 &  n_12245;
assign n_12247 =  x_2652 & ~n_12246;
assign n_12248 = ~x_2652 &  n_12246;
assign n_12249 = ~n_12247 & ~n_12248;
assign n_12250 = ~n_12237 & ~n_12241;
assign n_12251 =  x_1995 & ~x_3800;
assign n_12252 = ~x_1995 &  x_3800;
assign n_12253 = ~n_12251 & ~n_12252;
assign n_12254 =  n_12233 &  n_12253;
assign n_12255 = ~n_12233 & ~n_12253;
assign n_12256 = ~n_12254 & ~n_12255;
assign n_12257 =  n_12250 & ~n_12256;
assign n_12258 = ~n_12250 &  n_12256;
assign n_12259 =  n_10870 & ~n_12258;
assign n_12260 = ~n_12257 &  n_12259;
assign n_12261 =  x_4808 &  n_10875;
assign n_12262 =  x_2651 &  n_10878;
assign n_12263 = ~n_12261 & ~n_12262;
assign n_12264 = ~n_12260 &  n_12263;
assign n_12265 = ~n_12209 & ~n_12213;
assign n_12266 =  x_2219 & ~x_3736;
assign n_12267 = ~x_2219 &  x_3736;
assign n_12268 = ~n_12266 & ~n_12267;
assign n_12269 =  n_12205 &  n_12268;
assign n_12270 = ~n_12205 & ~n_12268;
assign n_12271 = ~n_12269 & ~n_12270;
assign n_12272 =  n_12265 & ~n_12271;
assign n_12273 = ~n_12265 &  n_12271;
assign n_12274 =  n_10871 & ~n_12273;
assign n_12275 = ~n_12272 &  n_12274;
assign n_12276 = ~n_12225 & ~n_12229;
assign n_12277 =  x_1483 & ~x_4169;
assign n_12278 = ~x_1483 &  x_4169;
assign n_12279 = ~n_12277 & ~n_12278;
assign n_12280 =  n_12221 &  n_12279;
assign n_12281 = ~n_12221 & ~n_12279;
assign n_12282 = ~n_12280 & ~n_12281;
assign n_12283 =  n_12276 & ~n_12282;
assign n_12284 = ~n_12276 &  n_12282;
assign n_12285 =  n_10873 & ~n_12284;
assign n_12286 = ~n_12283 &  n_12285;
assign n_12287 = ~n_12275 & ~n_12286;
assign n_12288 =  n_12264 &  n_12287;
assign n_12289 =  x_2651 & ~n_12288;
assign n_12290 = ~x_2651 &  n_12288;
assign n_12291 = ~n_12289 & ~n_12290;
assign n_12292 =  n_6 &  n_356;
assign n_12293 =  n_554 &  n_12292;
assign n_12294 = ~x_1603 &  x_1604;
assign n_12295 =  x_1605 &  n_12294;
assign n_12296 = ~x_1599 &  x_1600;
assign n_12297 = ~x_1601 &  x_1602;
assign n_12298 =  n_12296 &  n_12297;
assign n_12299 = ~x_1595 & ~x_1596;
assign n_12300 = ~x_1597 & ~x_1598;
assign n_12301 =  n_12299 &  n_12300;
assign n_12302 =  n_12298 &  n_12301;
assign n_12303 =  n_12295 &  n_12302;
assign n_12304 = ~x_1583 & ~x_1584;
assign n_12305 = ~x_1585 & ~x_1586;
assign n_12306 =  n_12304 &  n_12305;
assign n_12307 = ~x_1579 & ~x_1580;
assign n_12308 = ~x_1581 & ~x_1582;
assign n_12309 =  n_12307 &  n_12308;
assign n_12310 =  n_12306 &  n_12309;
assign n_12311 = ~x_1591 & ~x_1592;
assign n_12312 = ~x_1593 & ~x_1594;
assign n_12313 =  n_12311 &  n_12312;
assign n_12314 = ~x_1587 & ~x_1588;
assign n_12315 = ~x_1589 & ~x_1590;
assign n_12316 =  n_12314 &  n_12315;
assign n_12317 =  n_12313 &  n_12316;
assign n_12318 =  n_12310 &  n_12317;
assign n_12319 =  n_12303 &  n_12318;
assign n_12320 = ~x_1606 &  x_1607;
assign n_12321 =  x_1608 &  x_1609;
assign n_12322 =  n_12320 &  n_12321;
assign n_12323 =  n_12319 &  n_12322;
assign n_12324 =  x_1610 &  n_12323;
assign n_12325 =  x_1606 & ~x_1607;
assign n_12326 = ~x_1608 &  n_12325;
assign n_12327 =  n_12319 &  n_12326;
assign n_12328 =  x_1609 &  n_12327;
assign n_12329 = ~x_1610 &  n_12328;
assign n_12330 = ~x_1609 &  n_12327;
assign n_12331 =  x_1610 &  n_12330;
assign n_12332 = ~x_1610 &  n_12330;
assign n_12333 =  i_32 & ~n_12332;
assign n_12334 =  x_3064 &  n_12332;
assign n_12335 = ~n_12333 & ~n_12334;
assign n_12336 = ~n_12331 & ~n_12335;
assign n_12337 =  x_3032 &  n_12331;
assign n_12338 = ~n_12336 & ~n_12337;
assign n_12339 = ~n_12329 & ~n_12338;
assign n_12340 =  x_2906 &  n_12329;
assign n_12341 = ~n_12339 & ~n_12340;
assign n_12342 = ~n_12324 & ~n_12341;
assign n_12343 =  x_2842 &  n_12324;
assign n_12344 = ~n_12342 & ~n_12343;
assign n_12345 =  n_12293 & ~n_12344;
assign n_12346 =  x_2650 & ~n_12293;
assign n_12347 = ~n_12345 & ~n_12346;
assign n_12348 =  x_2650 & ~n_12347;
assign n_12349 = ~x_2650 &  n_12347;
assign n_12350 = ~n_12348 & ~n_12349;
assign n_12351 =  i_31 & ~n_12332;
assign n_12352 =  x_3063 &  n_12332;
assign n_12353 = ~n_12351 & ~n_12352;
assign n_12354 = ~n_12331 & ~n_12353;
assign n_12355 =  x_3031 &  n_12331;
assign n_12356 = ~n_12354 & ~n_12355;
assign n_12357 = ~n_12329 & ~n_12356;
assign n_12358 =  x_2905 &  n_12329;
assign n_12359 = ~n_12357 & ~n_12358;
assign n_12360 = ~n_12324 & ~n_12359;
assign n_12361 =  x_2841 &  n_12324;
assign n_12362 = ~n_12360 & ~n_12361;
assign n_12363 =  n_12293 & ~n_12362;
assign n_12364 =  x_2649 & ~n_12293;
assign n_12365 = ~n_12363 & ~n_12364;
assign n_12366 =  x_2649 & ~n_12365;
assign n_12367 = ~x_2649 &  n_12365;
assign n_12368 = ~n_12366 & ~n_12367;
assign n_12369 =  i_30 & ~n_12332;
assign n_12370 =  x_3062 &  n_12332;
assign n_12371 = ~n_12369 & ~n_12370;
assign n_12372 = ~n_12331 & ~n_12371;
assign n_12373 =  x_3030 &  n_12331;
assign n_12374 = ~n_12372 & ~n_12373;
assign n_12375 = ~n_12329 & ~n_12374;
assign n_12376 =  x_2904 &  n_12329;
assign n_12377 = ~n_12375 & ~n_12376;
assign n_12378 = ~n_12324 & ~n_12377;
assign n_12379 =  x_2840 &  n_12324;
assign n_12380 = ~n_12378 & ~n_12379;
assign n_12381 =  n_12293 & ~n_12380;
assign n_12382 =  x_2648 & ~n_12293;
assign n_12383 = ~n_12381 & ~n_12382;
assign n_12384 =  x_2648 & ~n_12383;
assign n_12385 = ~x_2648 &  n_12383;
assign n_12386 = ~n_12384 & ~n_12385;
assign n_12387 =  i_29 & ~n_12332;
assign n_12388 =  x_3061 &  n_12332;
assign n_12389 = ~n_12387 & ~n_12388;
assign n_12390 = ~n_12331 & ~n_12389;
assign n_12391 =  x_3029 &  n_12331;
assign n_12392 = ~n_12390 & ~n_12391;
assign n_12393 = ~n_12329 & ~n_12392;
assign n_12394 =  x_2903 &  n_12329;
assign n_12395 = ~n_12393 & ~n_12394;
assign n_12396 = ~n_12324 & ~n_12395;
assign n_12397 =  x_2839 &  n_12324;
assign n_12398 = ~n_12396 & ~n_12397;
assign n_12399 =  n_12293 & ~n_12398;
assign n_12400 =  x_2647 & ~n_12293;
assign n_12401 = ~n_12399 & ~n_12400;
assign n_12402 =  x_2647 & ~n_12401;
assign n_12403 = ~x_2647 &  n_12401;
assign n_12404 = ~n_12402 & ~n_12403;
assign n_12405 =  i_28 & ~n_12332;
assign n_12406 =  x_3060 &  n_12332;
assign n_12407 = ~n_12405 & ~n_12406;
assign n_12408 = ~n_12331 & ~n_12407;
assign n_12409 =  x_3028 &  n_12331;
assign n_12410 = ~n_12408 & ~n_12409;
assign n_12411 = ~n_12329 & ~n_12410;
assign n_12412 =  x_2902 &  n_12329;
assign n_12413 = ~n_12411 & ~n_12412;
assign n_12414 = ~n_12324 & ~n_12413;
assign n_12415 =  x_2838 &  n_12324;
assign n_12416 = ~n_12414 & ~n_12415;
assign n_12417 =  n_12293 & ~n_12416;
assign n_12418 =  x_2646 & ~n_12293;
assign n_12419 = ~n_12417 & ~n_12418;
assign n_12420 =  x_2646 & ~n_12419;
assign n_12421 = ~x_2646 &  n_12419;
assign n_12422 = ~n_12420 & ~n_12421;
assign n_12423 =  i_27 & ~n_12332;
assign n_12424 =  x_3059 &  n_12332;
assign n_12425 = ~n_12423 & ~n_12424;
assign n_12426 = ~n_12331 & ~n_12425;
assign n_12427 =  x_3027 &  n_12331;
assign n_12428 = ~n_12426 & ~n_12427;
assign n_12429 = ~n_12329 & ~n_12428;
assign n_12430 =  x_2901 &  n_12329;
assign n_12431 = ~n_12429 & ~n_12430;
assign n_12432 = ~n_12324 & ~n_12431;
assign n_12433 =  x_2837 &  n_12324;
assign n_12434 = ~n_12432 & ~n_12433;
assign n_12435 =  n_12293 & ~n_12434;
assign n_12436 =  x_2645 & ~n_12293;
assign n_12437 = ~n_12435 & ~n_12436;
assign n_12438 =  x_2645 & ~n_12437;
assign n_12439 = ~x_2645 &  n_12437;
assign n_12440 = ~n_12438 & ~n_12439;
assign n_12441 =  i_26 & ~n_12332;
assign n_12442 =  x_3058 &  n_12332;
assign n_12443 = ~n_12441 & ~n_12442;
assign n_12444 = ~n_12331 & ~n_12443;
assign n_12445 =  x_3026 &  n_12331;
assign n_12446 = ~n_12444 & ~n_12445;
assign n_12447 = ~n_12329 & ~n_12446;
assign n_12448 =  x_2900 &  n_12329;
assign n_12449 = ~n_12447 & ~n_12448;
assign n_12450 = ~n_12324 & ~n_12449;
assign n_12451 =  x_2836 &  n_12324;
assign n_12452 = ~n_12450 & ~n_12451;
assign n_12453 =  n_12293 & ~n_12452;
assign n_12454 =  x_2644 & ~n_12293;
assign n_12455 = ~n_12453 & ~n_12454;
assign n_12456 =  x_2644 & ~n_12455;
assign n_12457 = ~x_2644 &  n_12455;
assign n_12458 = ~n_12456 & ~n_12457;
assign n_12459 =  i_25 & ~n_12332;
assign n_12460 =  x_3057 &  n_12332;
assign n_12461 = ~n_12459 & ~n_12460;
assign n_12462 = ~n_12331 & ~n_12461;
assign n_12463 =  x_3025 &  n_12331;
assign n_12464 = ~n_12462 & ~n_12463;
assign n_12465 = ~n_12329 & ~n_12464;
assign n_12466 =  x_2899 &  n_12329;
assign n_12467 = ~n_12465 & ~n_12466;
assign n_12468 = ~n_12324 & ~n_12467;
assign n_12469 =  x_2835 &  n_12324;
assign n_12470 = ~n_12468 & ~n_12469;
assign n_12471 =  n_12293 & ~n_12470;
assign n_12472 =  x_2643 & ~n_12293;
assign n_12473 = ~n_12471 & ~n_12472;
assign n_12474 =  x_2643 & ~n_12473;
assign n_12475 = ~x_2643 &  n_12473;
assign n_12476 = ~n_12474 & ~n_12475;
assign n_12477 =  i_24 & ~n_12332;
assign n_12478 =  x_3056 &  n_12332;
assign n_12479 = ~n_12477 & ~n_12478;
assign n_12480 = ~n_12331 & ~n_12479;
assign n_12481 =  x_3024 &  n_12331;
assign n_12482 = ~n_12480 & ~n_12481;
assign n_12483 = ~n_12329 & ~n_12482;
assign n_12484 =  x_2898 &  n_12329;
assign n_12485 = ~n_12483 & ~n_12484;
assign n_12486 = ~n_12324 & ~n_12485;
assign n_12487 =  x_2834 &  n_12324;
assign n_12488 = ~n_12486 & ~n_12487;
assign n_12489 =  n_12293 & ~n_12488;
assign n_12490 =  x_2642 & ~n_12293;
assign n_12491 = ~n_12489 & ~n_12490;
assign n_12492 =  x_2642 & ~n_12491;
assign n_12493 = ~x_2642 &  n_12491;
assign n_12494 = ~n_12492 & ~n_12493;
assign n_12495 =  i_23 & ~n_12332;
assign n_12496 =  x_3055 &  n_12332;
assign n_12497 = ~n_12495 & ~n_12496;
assign n_12498 = ~n_12331 & ~n_12497;
assign n_12499 =  x_3023 &  n_12331;
assign n_12500 = ~n_12498 & ~n_12499;
assign n_12501 = ~n_12329 & ~n_12500;
assign n_12502 =  x_2897 &  n_12329;
assign n_12503 = ~n_12501 & ~n_12502;
assign n_12504 = ~n_12324 & ~n_12503;
assign n_12505 =  x_2833 &  n_12324;
assign n_12506 = ~n_12504 & ~n_12505;
assign n_12507 =  n_12293 & ~n_12506;
assign n_12508 =  x_2641 & ~n_12293;
assign n_12509 = ~n_12507 & ~n_12508;
assign n_12510 =  x_2641 & ~n_12509;
assign n_12511 = ~x_2641 &  n_12509;
assign n_12512 = ~n_12510 & ~n_12511;
assign n_12513 =  i_22 & ~n_12332;
assign n_12514 =  x_3054 &  n_12332;
assign n_12515 = ~n_12513 & ~n_12514;
assign n_12516 = ~n_12331 & ~n_12515;
assign n_12517 =  x_3022 &  n_12331;
assign n_12518 = ~n_12516 & ~n_12517;
assign n_12519 = ~n_12329 & ~n_12518;
assign n_12520 =  x_2896 &  n_12329;
assign n_12521 = ~n_12519 & ~n_12520;
assign n_12522 = ~n_12324 & ~n_12521;
assign n_12523 =  x_2832 &  n_12324;
assign n_12524 = ~n_12522 & ~n_12523;
assign n_12525 =  n_12293 & ~n_12524;
assign n_12526 =  x_2640 & ~n_12293;
assign n_12527 = ~n_12525 & ~n_12526;
assign n_12528 =  x_2640 & ~n_12527;
assign n_12529 = ~x_2640 &  n_12527;
assign n_12530 = ~n_12528 & ~n_12529;
assign n_12531 =  i_21 & ~n_12332;
assign n_12532 =  x_3053 &  n_12332;
assign n_12533 = ~n_12531 & ~n_12532;
assign n_12534 = ~n_12331 & ~n_12533;
assign n_12535 =  x_3021 &  n_12331;
assign n_12536 = ~n_12534 & ~n_12535;
assign n_12537 = ~n_12329 & ~n_12536;
assign n_12538 =  x_2895 &  n_12329;
assign n_12539 = ~n_12537 & ~n_12538;
assign n_12540 = ~n_12324 & ~n_12539;
assign n_12541 =  x_2831 &  n_12324;
assign n_12542 = ~n_12540 & ~n_12541;
assign n_12543 =  n_12293 & ~n_12542;
assign n_12544 =  x_2639 & ~n_12293;
assign n_12545 = ~n_12543 & ~n_12544;
assign n_12546 =  x_2639 & ~n_12545;
assign n_12547 = ~x_2639 &  n_12545;
assign n_12548 = ~n_12546 & ~n_12547;
assign n_12549 =  i_20 & ~n_12332;
assign n_12550 =  x_3052 &  n_12332;
assign n_12551 = ~n_12549 & ~n_12550;
assign n_12552 = ~n_12331 & ~n_12551;
assign n_12553 =  x_3020 &  n_12331;
assign n_12554 = ~n_12552 & ~n_12553;
assign n_12555 = ~n_12329 & ~n_12554;
assign n_12556 =  x_2894 &  n_12329;
assign n_12557 = ~n_12555 & ~n_12556;
assign n_12558 = ~n_12324 & ~n_12557;
assign n_12559 =  x_2830 &  n_12324;
assign n_12560 = ~n_12558 & ~n_12559;
assign n_12561 =  n_12293 & ~n_12560;
assign n_12562 =  x_2638 & ~n_12293;
assign n_12563 = ~n_12561 & ~n_12562;
assign n_12564 =  x_2638 & ~n_12563;
assign n_12565 = ~x_2638 &  n_12563;
assign n_12566 = ~n_12564 & ~n_12565;
assign n_12567 =  i_19 & ~n_12332;
assign n_12568 =  x_3051 &  n_12332;
assign n_12569 = ~n_12567 & ~n_12568;
assign n_12570 = ~n_12331 & ~n_12569;
assign n_12571 =  x_3019 &  n_12331;
assign n_12572 = ~n_12570 & ~n_12571;
assign n_12573 = ~n_12329 & ~n_12572;
assign n_12574 =  x_2893 &  n_12329;
assign n_12575 = ~n_12573 & ~n_12574;
assign n_12576 = ~n_12324 & ~n_12575;
assign n_12577 =  x_2829 &  n_12324;
assign n_12578 = ~n_12576 & ~n_12577;
assign n_12579 =  n_12293 & ~n_12578;
assign n_12580 =  x_2637 & ~n_12293;
assign n_12581 = ~n_12579 & ~n_12580;
assign n_12582 =  x_2637 & ~n_12581;
assign n_12583 = ~x_2637 &  n_12581;
assign n_12584 = ~n_12582 & ~n_12583;
assign n_12585 =  i_18 & ~n_12332;
assign n_12586 =  x_3050 &  n_12332;
assign n_12587 = ~n_12585 & ~n_12586;
assign n_12588 = ~n_12331 & ~n_12587;
assign n_12589 =  x_3018 &  n_12331;
assign n_12590 = ~n_12588 & ~n_12589;
assign n_12591 = ~n_12329 & ~n_12590;
assign n_12592 =  x_2892 &  n_12329;
assign n_12593 = ~n_12591 & ~n_12592;
assign n_12594 = ~n_12324 & ~n_12593;
assign n_12595 =  x_2828 &  n_12324;
assign n_12596 = ~n_12594 & ~n_12595;
assign n_12597 =  n_12293 & ~n_12596;
assign n_12598 =  x_2636 & ~n_12293;
assign n_12599 = ~n_12597 & ~n_12598;
assign n_12600 =  x_2636 & ~n_12599;
assign n_12601 = ~x_2636 &  n_12599;
assign n_12602 = ~n_12600 & ~n_12601;
assign n_12603 =  i_17 & ~n_12332;
assign n_12604 =  x_3049 &  n_12332;
assign n_12605 = ~n_12603 & ~n_12604;
assign n_12606 = ~n_12331 & ~n_12605;
assign n_12607 =  x_3017 &  n_12331;
assign n_12608 = ~n_12606 & ~n_12607;
assign n_12609 = ~n_12329 & ~n_12608;
assign n_12610 =  x_2891 &  n_12329;
assign n_12611 = ~n_12609 & ~n_12610;
assign n_12612 = ~n_12324 & ~n_12611;
assign n_12613 =  x_2827 &  n_12324;
assign n_12614 = ~n_12612 & ~n_12613;
assign n_12615 =  n_12293 & ~n_12614;
assign n_12616 =  x_2635 & ~n_12293;
assign n_12617 = ~n_12615 & ~n_12616;
assign n_12618 =  x_2635 & ~n_12617;
assign n_12619 = ~x_2635 &  n_12617;
assign n_12620 = ~n_12618 & ~n_12619;
assign n_12621 =  i_16 & ~n_12332;
assign n_12622 =  x_3048 &  n_12332;
assign n_12623 = ~n_12621 & ~n_12622;
assign n_12624 = ~n_12331 & ~n_12623;
assign n_12625 =  x_3016 &  n_12331;
assign n_12626 = ~n_12624 & ~n_12625;
assign n_12627 = ~n_12329 & ~n_12626;
assign n_12628 =  x_2890 &  n_12329;
assign n_12629 = ~n_12627 & ~n_12628;
assign n_12630 = ~n_12324 & ~n_12629;
assign n_12631 =  x_2826 &  n_12324;
assign n_12632 = ~n_12630 & ~n_12631;
assign n_12633 =  n_12293 & ~n_12632;
assign n_12634 =  x_2634 & ~n_12293;
assign n_12635 = ~n_12633 & ~n_12634;
assign n_12636 =  x_2634 & ~n_12635;
assign n_12637 = ~x_2634 &  n_12635;
assign n_12638 = ~n_12636 & ~n_12637;
assign n_12639 =  i_15 & ~n_12332;
assign n_12640 =  x_3047 &  n_12332;
assign n_12641 = ~n_12639 & ~n_12640;
assign n_12642 = ~n_12331 & ~n_12641;
assign n_12643 =  x_3015 &  n_12331;
assign n_12644 = ~n_12642 & ~n_12643;
assign n_12645 = ~n_12329 & ~n_12644;
assign n_12646 =  x_2889 &  n_12329;
assign n_12647 = ~n_12645 & ~n_12646;
assign n_12648 = ~n_12324 & ~n_12647;
assign n_12649 =  x_2825 &  n_12324;
assign n_12650 = ~n_12648 & ~n_12649;
assign n_12651 =  n_12293 & ~n_12650;
assign n_12652 =  x_2633 & ~n_12293;
assign n_12653 = ~n_12651 & ~n_12652;
assign n_12654 =  x_2633 & ~n_12653;
assign n_12655 = ~x_2633 &  n_12653;
assign n_12656 = ~n_12654 & ~n_12655;
assign n_12657 =  i_14 & ~n_12332;
assign n_12658 =  x_3046 &  n_12332;
assign n_12659 = ~n_12657 & ~n_12658;
assign n_12660 = ~n_12331 & ~n_12659;
assign n_12661 =  x_3014 &  n_12331;
assign n_12662 = ~n_12660 & ~n_12661;
assign n_12663 = ~n_12329 & ~n_12662;
assign n_12664 =  x_2888 &  n_12329;
assign n_12665 = ~n_12663 & ~n_12664;
assign n_12666 = ~n_12324 & ~n_12665;
assign n_12667 =  x_2824 &  n_12324;
assign n_12668 = ~n_12666 & ~n_12667;
assign n_12669 =  n_12293 & ~n_12668;
assign n_12670 =  x_2632 & ~n_12293;
assign n_12671 = ~n_12669 & ~n_12670;
assign n_12672 =  x_2632 & ~n_12671;
assign n_12673 = ~x_2632 &  n_12671;
assign n_12674 = ~n_12672 & ~n_12673;
assign n_12675 =  i_13 & ~n_12332;
assign n_12676 =  x_3045 &  n_12332;
assign n_12677 = ~n_12675 & ~n_12676;
assign n_12678 = ~n_12331 & ~n_12677;
assign n_12679 =  x_3013 &  n_12331;
assign n_12680 = ~n_12678 & ~n_12679;
assign n_12681 = ~n_12329 & ~n_12680;
assign n_12682 =  x_2887 &  n_12329;
assign n_12683 = ~n_12681 & ~n_12682;
assign n_12684 = ~n_12324 & ~n_12683;
assign n_12685 =  x_2823 &  n_12324;
assign n_12686 = ~n_12684 & ~n_12685;
assign n_12687 =  n_12293 & ~n_12686;
assign n_12688 =  x_2631 & ~n_12293;
assign n_12689 = ~n_12687 & ~n_12688;
assign n_12690 =  x_2631 & ~n_12689;
assign n_12691 = ~x_2631 &  n_12689;
assign n_12692 = ~n_12690 & ~n_12691;
assign n_12693 =  i_12 & ~n_12332;
assign n_12694 =  x_3044 &  n_12332;
assign n_12695 = ~n_12693 & ~n_12694;
assign n_12696 = ~n_12331 & ~n_12695;
assign n_12697 =  x_3012 &  n_12331;
assign n_12698 = ~n_12696 & ~n_12697;
assign n_12699 = ~n_12329 & ~n_12698;
assign n_12700 =  x_2886 &  n_12329;
assign n_12701 = ~n_12699 & ~n_12700;
assign n_12702 = ~n_12324 & ~n_12701;
assign n_12703 =  x_2822 &  n_12324;
assign n_12704 = ~n_12702 & ~n_12703;
assign n_12705 =  n_12293 & ~n_12704;
assign n_12706 =  x_2630 & ~n_12293;
assign n_12707 = ~n_12705 & ~n_12706;
assign n_12708 =  x_2630 & ~n_12707;
assign n_12709 = ~x_2630 &  n_12707;
assign n_12710 = ~n_12708 & ~n_12709;
assign n_12711 =  i_11 & ~n_12332;
assign n_12712 =  x_3043 &  n_12332;
assign n_12713 = ~n_12711 & ~n_12712;
assign n_12714 = ~n_12331 & ~n_12713;
assign n_12715 =  x_3011 &  n_12331;
assign n_12716 = ~n_12714 & ~n_12715;
assign n_12717 = ~n_12329 & ~n_12716;
assign n_12718 =  x_2885 &  n_12329;
assign n_12719 = ~n_12717 & ~n_12718;
assign n_12720 = ~n_12324 & ~n_12719;
assign n_12721 =  x_2821 &  n_12324;
assign n_12722 = ~n_12720 & ~n_12721;
assign n_12723 =  n_12293 & ~n_12722;
assign n_12724 =  x_2629 & ~n_12293;
assign n_12725 = ~n_12723 & ~n_12724;
assign n_12726 =  x_2629 & ~n_12725;
assign n_12727 = ~x_2629 &  n_12725;
assign n_12728 = ~n_12726 & ~n_12727;
assign n_12729 =  i_10 & ~n_12332;
assign n_12730 =  x_3042 &  n_12332;
assign n_12731 = ~n_12729 & ~n_12730;
assign n_12732 = ~n_12331 & ~n_12731;
assign n_12733 =  x_3010 &  n_12331;
assign n_12734 = ~n_12732 & ~n_12733;
assign n_12735 = ~n_12329 & ~n_12734;
assign n_12736 =  x_2884 &  n_12329;
assign n_12737 = ~n_12735 & ~n_12736;
assign n_12738 = ~n_12324 & ~n_12737;
assign n_12739 =  x_2820 &  n_12324;
assign n_12740 = ~n_12738 & ~n_12739;
assign n_12741 =  n_12293 & ~n_12740;
assign n_12742 =  x_2628 & ~n_12293;
assign n_12743 = ~n_12741 & ~n_12742;
assign n_12744 =  x_2628 & ~n_12743;
assign n_12745 = ~x_2628 &  n_12743;
assign n_12746 = ~n_12744 & ~n_12745;
assign n_12747 =  i_9 & ~n_12332;
assign n_12748 =  x_3041 &  n_12332;
assign n_12749 = ~n_12747 & ~n_12748;
assign n_12750 = ~n_12331 & ~n_12749;
assign n_12751 =  x_3009 &  n_12331;
assign n_12752 = ~n_12750 & ~n_12751;
assign n_12753 = ~n_12329 & ~n_12752;
assign n_12754 =  x_2883 &  n_12329;
assign n_12755 = ~n_12753 & ~n_12754;
assign n_12756 = ~n_12324 & ~n_12755;
assign n_12757 =  x_2819 &  n_12324;
assign n_12758 = ~n_12756 & ~n_12757;
assign n_12759 =  n_12293 & ~n_12758;
assign n_12760 =  x_2627 & ~n_12293;
assign n_12761 = ~n_12759 & ~n_12760;
assign n_12762 =  x_2627 & ~n_12761;
assign n_12763 = ~x_2627 &  n_12761;
assign n_12764 = ~n_12762 & ~n_12763;
assign n_12765 =  i_8 & ~n_12332;
assign n_12766 =  x_3040 &  n_12332;
assign n_12767 = ~n_12765 & ~n_12766;
assign n_12768 = ~n_12331 & ~n_12767;
assign n_12769 =  x_3008 &  n_12331;
assign n_12770 = ~n_12768 & ~n_12769;
assign n_12771 = ~n_12329 & ~n_12770;
assign n_12772 =  x_2882 &  n_12329;
assign n_12773 = ~n_12771 & ~n_12772;
assign n_12774 = ~n_12324 & ~n_12773;
assign n_12775 =  x_2818 &  n_12324;
assign n_12776 = ~n_12774 & ~n_12775;
assign n_12777 =  n_12293 & ~n_12776;
assign n_12778 =  x_2626 & ~n_12293;
assign n_12779 = ~n_12777 & ~n_12778;
assign n_12780 =  x_2626 & ~n_12779;
assign n_12781 = ~x_2626 &  n_12779;
assign n_12782 = ~n_12780 & ~n_12781;
assign n_12783 =  i_7 & ~n_12332;
assign n_12784 =  x_3039 &  n_12332;
assign n_12785 = ~n_12783 & ~n_12784;
assign n_12786 = ~n_12331 & ~n_12785;
assign n_12787 =  x_3007 &  n_12331;
assign n_12788 = ~n_12786 & ~n_12787;
assign n_12789 = ~n_12329 & ~n_12788;
assign n_12790 =  x_2881 &  n_12329;
assign n_12791 = ~n_12789 & ~n_12790;
assign n_12792 = ~n_12324 & ~n_12791;
assign n_12793 =  x_2817 &  n_12324;
assign n_12794 = ~n_12792 & ~n_12793;
assign n_12795 =  n_12293 & ~n_12794;
assign n_12796 =  x_2625 & ~n_12293;
assign n_12797 = ~n_12795 & ~n_12796;
assign n_12798 =  x_2625 & ~n_12797;
assign n_12799 = ~x_2625 &  n_12797;
assign n_12800 = ~n_12798 & ~n_12799;
assign n_12801 =  i_6 & ~n_12332;
assign n_12802 =  x_3038 &  n_12332;
assign n_12803 = ~n_12801 & ~n_12802;
assign n_12804 = ~n_12331 & ~n_12803;
assign n_12805 =  x_3006 &  n_12331;
assign n_12806 = ~n_12804 & ~n_12805;
assign n_12807 = ~n_12329 & ~n_12806;
assign n_12808 =  x_2880 &  n_12329;
assign n_12809 = ~n_12807 & ~n_12808;
assign n_12810 = ~n_12324 & ~n_12809;
assign n_12811 =  x_2816 &  n_12324;
assign n_12812 = ~n_12810 & ~n_12811;
assign n_12813 =  n_12293 & ~n_12812;
assign n_12814 =  x_2624 & ~n_12293;
assign n_12815 = ~n_12813 & ~n_12814;
assign n_12816 =  x_2624 & ~n_12815;
assign n_12817 = ~x_2624 &  n_12815;
assign n_12818 = ~n_12816 & ~n_12817;
assign n_12819 =  i_5 & ~n_12332;
assign n_12820 =  x_3037 &  n_12332;
assign n_12821 = ~n_12819 & ~n_12820;
assign n_12822 = ~n_12331 & ~n_12821;
assign n_12823 =  x_3005 &  n_12331;
assign n_12824 = ~n_12822 & ~n_12823;
assign n_12825 = ~n_12329 & ~n_12824;
assign n_12826 =  x_2879 &  n_12329;
assign n_12827 = ~n_12825 & ~n_12826;
assign n_12828 = ~n_12324 & ~n_12827;
assign n_12829 =  x_2815 &  n_12324;
assign n_12830 = ~n_12828 & ~n_12829;
assign n_12831 =  n_12293 & ~n_12830;
assign n_12832 =  x_2623 & ~n_12293;
assign n_12833 = ~n_12831 & ~n_12832;
assign n_12834 =  x_2623 & ~n_12833;
assign n_12835 = ~x_2623 &  n_12833;
assign n_12836 = ~n_12834 & ~n_12835;
assign n_12837 =  i_4 & ~n_12332;
assign n_12838 =  x_3036 &  n_12332;
assign n_12839 = ~n_12837 & ~n_12838;
assign n_12840 = ~n_12331 & ~n_12839;
assign n_12841 =  x_3004 &  n_12331;
assign n_12842 = ~n_12840 & ~n_12841;
assign n_12843 = ~n_12329 & ~n_12842;
assign n_12844 =  x_2878 &  n_12329;
assign n_12845 = ~n_12843 & ~n_12844;
assign n_12846 = ~n_12324 & ~n_12845;
assign n_12847 =  x_2814 &  n_12324;
assign n_12848 = ~n_12846 & ~n_12847;
assign n_12849 =  n_12293 & ~n_12848;
assign n_12850 =  x_2622 & ~n_12293;
assign n_12851 = ~n_12849 & ~n_12850;
assign n_12852 =  x_2622 & ~n_12851;
assign n_12853 = ~x_2622 &  n_12851;
assign n_12854 = ~n_12852 & ~n_12853;
assign n_12855 =  i_3 & ~n_12332;
assign n_12856 =  x_3035 &  n_12332;
assign n_12857 = ~n_12855 & ~n_12856;
assign n_12858 = ~n_12331 & ~n_12857;
assign n_12859 =  x_3003 &  n_12331;
assign n_12860 = ~n_12858 & ~n_12859;
assign n_12861 = ~n_12329 & ~n_12860;
assign n_12862 =  x_2877 &  n_12329;
assign n_12863 = ~n_12861 & ~n_12862;
assign n_12864 = ~n_12324 & ~n_12863;
assign n_12865 =  x_2813 &  n_12324;
assign n_12866 = ~n_12864 & ~n_12865;
assign n_12867 =  n_12293 & ~n_12866;
assign n_12868 =  x_2621 & ~n_12293;
assign n_12869 = ~n_12867 & ~n_12868;
assign n_12870 =  x_2621 & ~n_12869;
assign n_12871 = ~x_2621 &  n_12869;
assign n_12872 = ~n_12870 & ~n_12871;
assign n_12873 =  i_2 & ~n_12332;
assign n_12874 =  x_3034 &  n_12332;
assign n_12875 = ~n_12873 & ~n_12874;
assign n_12876 = ~n_12331 & ~n_12875;
assign n_12877 =  x_3002 &  n_12331;
assign n_12878 = ~n_12876 & ~n_12877;
assign n_12879 = ~n_12329 & ~n_12878;
assign n_12880 =  x_2876 &  n_12329;
assign n_12881 = ~n_12879 & ~n_12880;
assign n_12882 = ~n_12324 & ~n_12881;
assign n_12883 =  x_2812 &  n_12324;
assign n_12884 = ~n_12882 & ~n_12883;
assign n_12885 =  n_12293 & ~n_12884;
assign n_12886 =  x_2620 & ~n_12293;
assign n_12887 = ~n_12885 & ~n_12886;
assign n_12888 =  x_2620 & ~n_12887;
assign n_12889 = ~x_2620 &  n_12887;
assign n_12890 = ~n_12888 & ~n_12889;
assign n_12891 =  i_1 & ~n_12332;
assign n_12892 =  x_3033 &  n_12332;
assign n_12893 = ~n_12891 & ~n_12892;
assign n_12894 = ~n_12331 & ~n_12893;
assign n_12895 =  x_3001 &  n_12331;
assign n_12896 = ~n_12894 & ~n_12895;
assign n_12897 = ~n_12329 & ~n_12896;
assign n_12898 =  x_2875 &  n_12329;
assign n_12899 = ~n_12897 & ~n_12898;
assign n_12900 = ~n_12324 & ~n_12899;
assign n_12901 =  x_2811 &  n_12324;
assign n_12902 = ~n_12900 & ~n_12901;
assign n_12903 =  n_12293 & ~n_12902;
assign n_12904 =  x_2619 & ~n_12293;
assign n_12905 = ~n_12903 & ~n_12904;
assign n_12906 =  x_2619 & ~n_12905;
assign n_12907 = ~x_2619 &  n_12905;
assign n_12908 = ~n_12906 & ~n_12907;
assign n_12909 =  n_2095 &  n_10478;
assign n_12910 = ~x_43 &  n_5983;
assign n_12911 = ~n_12909 & ~n_12910;
assign n_12912 =  i_32 & ~n_12911;
assign n_12913 =  x_2618 &  n_12911;
assign n_12914 = ~n_12912 & ~n_12913;
assign n_12915 =  x_2618 & ~n_12914;
assign n_12916 = ~x_2618 &  n_12914;
assign n_12917 = ~n_12915 & ~n_12916;
assign n_12918 =  i_31 & ~n_12911;
assign n_12919 =  x_2617 &  n_12911;
assign n_12920 = ~n_12918 & ~n_12919;
assign n_12921 =  x_2617 & ~n_12920;
assign n_12922 = ~x_2617 &  n_12920;
assign n_12923 = ~n_12921 & ~n_12922;
assign n_12924 =  i_30 & ~n_12911;
assign n_12925 =  x_2616 &  n_12911;
assign n_12926 = ~n_12924 & ~n_12925;
assign n_12927 =  x_2616 & ~n_12926;
assign n_12928 = ~x_2616 &  n_12926;
assign n_12929 = ~n_12927 & ~n_12928;
assign n_12930 =  i_29 & ~n_12911;
assign n_12931 =  x_2615 &  n_12911;
assign n_12932 = ~n_12930 & ~n_12931;
assign n_12933 =  x_2615 & ~n_12932;
assign n_12934 = ~x_2615 &  n_12932;
assign n_12935 = ~n_12933 & ~n_12934;
assign n_12936 =  i_28 & ~n_12911;
assign n_12937 =  x_2614 &  n_12911;
assign n_12938 = ~n_12936 & ~n_12937;
assign n_12939 =  x_2614 & ~n_12938;
assign n_12940 = ~x_2614 &  n_12938;
assign n_12941 = ~n_12939 & ~n_12940;
assign n_12942 =  i_27 & ~n_12911;
assign n_12943 =  x_2613 &  n_12911;
assign n_12944 = ~n_12942 & ~n_12943;
assign n_12945 =  x_2613 & ~n_12944;
assign n_12946 = ~x_2613 &  n_12944;
assign n_12947 = ~n_12945 & ~n_12946;
assign n_12948 =  i_26 & ~n_12911;
assign n_12949 =  x_2612 &  n_12911;
assign n_12950 = ~n_12948 & ~n_12949;
assign n_12951 =  x_2612 & ~n_12950;
assign n_12952 = ~x_2612 &  n_12950;
assign n_12953 = ~n_12951 & ~n_12952;
assign n_12954 =  i_25 & ~n_12911;
assign n_12955 =  x_2611 &  n_12911;
assign n_12956 = ~n_12954 & ~n_12955;
assign n_12957 =  x_2611 & ~n_12956;
assign n_12958 = ~x_2611 &  n_12956;
assign n_12959 = ~n_12957 & ~n_12958;
assign n_12960 =  i_24 & ~n_12911;
assign n_12961 =  x_2610 &  n_12911;
assign n_12962 = ~n_12960 & ~n_12961;
assign n_12963 =  x_2610 & ~n_12962;
assign n_12964 = ~x_2610 &  n_12962;
assign n_12965 = ~n_12963 & ~n_12964;
assign n_12966 =  i_23 & ~n_12911;
assign n_12967 =  x_2609 &  n_12911;
assign n_12968 = ~n_12966 & ~n_12967;
assign n_12969 =  x_2609 & ~n_12968;
assign n_12970 = ~x_2609 &  n_12968;
assign n_12971 = ~n_12969 & ~n_12970;
assign n_12972 =  i_22 & ~n_12911;
assign n_12973 =  x_2608 &  n_12911;
assign n_12974 = ~n_12972 & ~n_12973;
assign n_12975 =  x_2608 & ~n_12974;
assign n_12976 = ~x_2608 &  n_12974;
assign n_12977 = ~n_12975 & ~n_12976;
assign n_12978 =  i_21 & ~n_12911;
assign n_12979 =  x_2607 &  n_12911;
assign n_12980 = ~n_12978 & ~n_12979;
assign n_12981 =  x_2607 & ~n_12980;
assign n_12982 = ~x_2607 &  n_12980;
assign n_12983 = ~n_12981 & ~n_12982;
assign n_12984 =  i_20 & ~n_12911;
assign n_12985 =  x_2606 &  n_12911;
assign n_12986 = ~n_12984 & ~n_12985;
assign n_12987 =  x_2606 & ~n_12986;
assign n_12988 = ~x_2606 &  n_12986;
assign n_12989 = ~n_12987 & ~n_12988;
assign n_12990 =  i_19 & ~n_12911;
assign n_12991 =  x_2605 &  n_12911;
assign n_12992 = ~n_12990 & ~n_12991;
assign n_12993 =  x_2605 & ~n_12992;
assign n_12994 = ~x_2605 &  n_12992;
assign n_12995 = ~n_12993 & ~n_12994;
assign n_12996 =  i_18 & ~n_12911;
assign n_12997 =  x_2604 &  n_12911;
assign n_12998 = ~n_12996 & ~n_12997;
assign n_12999 =  x_2604 & ~n_12998;
assign n_13000 = ~x_2604 &  n_12998;
assign n_13001 = ~n_12999 & ~n_13000;
assign n_13002 =  i_17 & ~n_12911;
assign n_13003 =  x_2603 &  n_12911;
assign n_13004 = ~n_13002 & ~n_13003;
assign n_13005 =  x_2603 & ~n_13004;
assign n_13006 = ~x_2603 &  n_13004;
assign n_13007 = ~n_13005 & ~n_13006;
assign n_13008 =  i_16 & ~n_12911;
assign n_13009 =  x_2602 &  n_12911;
assign n_13010 = ~n_13008 & ~n_13009;
assign n_13011 =  x_2602 & ~n_13010;
assign n_13012 = ~x_2602 &  n_13010;
assign n_13013 = ~n_13011 & ~n_13012;
assign n_13014 =  i_15 & ~n_12911;
assign n_13015 =  x_2601 &  n_12911;
assign n_13016 = ~n_13014 & ~n_13015;
assign n_13017 =  x_2601 & ~n_13016;
assign n_13018 = ~x_2601 &  n_13016;
assign n_13019 = ~n_13017 & ~n_13018;
assign n_13020 =  i_14 & ~n_12911;
assign n_13021 =  x_2600 &  n_12911;
assign n_13022 = ~n_13020 & ~n_13021;
assign n_13023 =  x_2600 & ~n_13022;
assign n_13024 = ~x_2600 &  n_13022;
assign n_13025 = ~n_13023 & ~n_13024;
assign n_13026 =  i_13 & ~n_12911;
assign n_13027 =  x_2599 &  n_12911;
assign n_13028 = ~n_13026 & ~n_13027;
assign n_13029 =  x_2599 & ~n_13028;
assign n_13030 = ~x_2599 &  n_13028;
assign n_13031 = ~n_13029 & ~n_13030;
assign n_13032 =  i_12 & ~n_12911;
assign n_13033 =  x_2598 &  n_12911;
assign n_13034 = ~n_13032 & ~n_13033;
assign n_13035 =  x_2598 & ~n_13034;
assign n_13036 = ~x_2598 &  n_13034;
assign n_13037 = ~n_13035 & ~n_13036;
assign n_13038 =  i_11 & ~n_12911;
assign n_13039 =  x_2597 &  n_12911;
assign n_13040 = ~n_13038 & ~n_13039;
assign n_13041 =  x_2597 & ~n_13040;
assign n_13042 = ~x_2597 &  n_13040;
assign n_13043 = ~n_13041 & ~n_13042;
assign n_13044 =  i_10 & ~n_12911;
assign n_13045 =  x_2596 &  n_12911;
assign n_13046 = ~n_13044 & ~n_13045;
assign n_13047 =  x_2596 & ~n_13046;
assign n_13048 = ~x_2596 &  n_13046;
assign n_13049 = ~n_13047 & ~n_13048;
assign n_13050 =  i_9 & ~n_12911;
assign n_13051 =  x_2595 &  n_12911;
assign n_13052 = ~n_13050 & ~n_13051;
assign n_13053 =  x_2595 & ~n_13052;
assign n_13054 = ~x_2595 &  n_13052;
assign n_13055 = ~n_13053 & ~n_13054;
assign n_13056 =  i_8 & ~n_12911;
assign n_13057 =  x_2594 &  n_12911;
assign n_13058 = ~n_13056 & ~n_13057;
assign n_13059 =  x_2594 & ~n_13058;
assign n_13060 = ~x_2594 &  n_13058;
assign n_13061 = ~n_13059 & ~n_13060;
assign n_13062 =  i_7 & ~n_12911;
assign n_13063 =  x_2593 &  n_12911;
assign n_13064 = ~n_13062 & ~n_13063;
assign n_13065 =  x_2593 & ~n_13064;
assign n_13066 = ~x_2593 &  n_13064;
assign n_13067 = ~n_13065 & ~n_13066;
assign n_13068 =  i_6 & ~n_12911;
assign n_13069 =  x_2592 &  n_12911;
assign n_13070 = ~n_13068 & ~n_13069;
assign n_13071 =  x_2592 & ~n_13070;
assign n_13072 = ~x_2592 &  n_13070;
assign n_13073 = ~n_13071 & ~n_13072;
assign n_13074 =  i_5 & ~n_12911;
assign n_13075 =  x_2591 &  n_12911;
assign n_13076 = ~n_13074 & ~n_13075;
assign n_13077 =  x_2591 & ~n_13076;
assign n_13078 = ~x_2591 &  n_13076;
assign n_13079 = ~n_13077 & ~n_13078;
assign n_13080 =  i_4 & ~n_12911;
assign n_13081 =  x_2590 &  n_12911;
assign n_13082 = ~n_13080 & ~n_13081;
assign n_13083 =  x_2590 & ~n_13082;
assign n_13084 = ~x_2590 &  n_13082;
assign n_13085 = ~n_13083 & ~n_13084;
assign n_13086 =  i_3 & ~n_12911;
assign n_13087 =  x_2589 &  n_12911;
assign n_13088 = ~n_13086 & ~n_13087;
assign n_13089 =  x_2589 & ~n_13088;
assign n_13090 = ~x_2589 &  n_13088;
assign n_13091 = ~n_13089 & ~n_13090;
assign n_13092 =  i_2 & ~n_12911;
assign n_13093 =  x_2588 &  n_12911;
assign n_13094 = ~n_13092 & ~n_13093;
assign n_13095 =  x_2588 & ~n_13094;
assign n_13096 = ~x_2588 &  n_13094;
assign n_13097 = ~n_13095 & ~n_13096;
assign n_13098 =  i_1 & ~n_12911;
assign n_13099 =  x_2587 &  n_12911;
assign n_13100 = ~n_13098 & ~n_13099;
assign n_13101 =  x_2587 & ~n_13100;
assign n_13102 = ~x_2587 &  n_13100;
assign n_13103 = ~n_13101 & ~n_13102;
assign n_13104 =  n_561 &  n_5654;
assign n_13105 =  n_13104 &  n_3619;
assign n_13106 = ~x_4768 &  x_4769;
assign n_13107 =  x_4770 &  n_13106;
assign n_13108 = ~x_4764 &  x_4765;
assign n_13109 = ~x_4766 &  x_4767;
assign n_13110 =  n_13108 &  n_13109;
assign n_13111 = ~x_4760 & ~x_4761;
assign n_13112 = ~x_4762 & ~x_4763;
assign n_13113 =  n_13111 &  n_13112;
assign n_13114 =  n_13110 &  n_13113;
assign n_13115 =  n_13107 &  n_13114;
assign n_13116 = ~x_4748 & ~x_4749;
assign n_13117 = ~x_4750 & ~x_4751;
assign n_13118 =  n_13116 &  n_13117;
assign n_13119 = ~x_4744 & ~x_4745;
assign n_13120 = ~x_4746 & ~x_4747;
assign n_13121 =  n_13119 &  n_13120;
assign n_13122 =  n_13118 &  n_13121;
assign n_13123 = ~x_4756 & ~x_4757;
assign n_13124 = ~x_4758 & ~x_4759;
assign n_13125 =  n_13123 &  n_13124;
assign n_13126 = ~x_4752 & ~x_4753;
assign n_13127 = ~x_4754 & ~x_4755;
assign n_13128 =  n_13126 &  n_13127;
assign n_13129 =  n_13125 &  n_13128;
assign n_13130 =  n_13122 &  n_13129;
assign n_13131 =  n_13115 &  n_13130;
assign n_13132 = ~x_4771 &  x_4772;
assign n_13133 =  x_4773 &  x_4774;
assign n_13134 =  n_13132 &  n_13133;
assign n_13135 =  n_13131 &  n_13134;
assign n_13136 =  x_4775 &  n_13135;
assign n_13137 =  x_4771 & ~x_4772;
assign n_13138 = ~x_4773 &  n_13137;
assign n_13139 =  n_13131 &  n_13138;
assign n_13140 =  x_4774 &  n_13139;
assign n_13141 = ~x_4775 &  n_13140;
assign n_13142 = ~x_4774 &  n_13139;
assign n_13143 =  x_4775 &  n_13142;
assign n_13144 = ~x_3032 &  n_13143;
assign n_13145 = ~x_4775 &  n_13142;
assign n_13146 = ~x_3064 &  n_13145;
assign n_13147 = ~i_32 & ~n_13142;
assign n_13148 = ~n_13146 & ~n_13147;
assign n_13149 = ~n_13144 &  n_13148;
assign n_13150 = ~n_13141 & ~n_13149;
assign n_13151 = ~x_2906 &  n_13141;
assign n_13152 = ~n_13150 & ~n_13151;
assign n_13153 = ~n_13136 & ~n_13152;
assign n_13154 = ~x_2842 &  n_13136;
assign n_13155 = ~n_13153 & ~n_13154;
assign n_13156 =  n_13105 & ~n_13155;
assign n_13157 = ~x_2586 & ~n_13105;
assign n_13158 = ~n_13156 & ~n_13157;
assign n_13159 =  x_2586 &  n_13158;
assign n_13160 = ~x_2586 & ~n_13158;
assign n_13161 = ~n_13159 & ~n_13160;
assign n_13162 = ~x_3031 &  n_13143;
assign n_13163 = ~x_3063 &  n_13145;
assign n_13164 = ~i_31 & ~n_13142;
assign n_13165 = ~n_13163 & ~n_13164;
assign n_13166 = ~n_13162 &  n_13165;
assign n_13167 = ~n_13141 & ~n_13166;
assign n_13168 = ~x_2905 &  n_13141;
assign n_13169 = ~n_13167 & ~n_13168;
assign n_13170 = ~n_13136 & ~n_13169;
assign n_13171 = ~x_2841 &  n_13136;
assign n_13172 = ~n_13170 & ~n_13171;
assign n_13173 =  n_13105 & ~n_13172;
assign n_13174 = ~x_2585 & ~n_13105;
assign n_13175 = ~n_13173 & ~n_13174;
assign n_13176 =  x_2585 &  n_13175;
assign n_13177 = ~x_2585 & ~n_13175;
assign n_13178 = ~n_13176 & ~n_13177;
assign n_13179 = ~x_3030 &  n_13143;
assign n_13180 = ~x_3062 &  n_13145;
assign n_13181 = ~i_30 & ~n_13142;
assign n_13182 = ~n_13180 & ~n_13181;
assign n_13183 = ~n_13179 &  n_13182;
assign n_13184 = ~n_13141 & ~n_13183;
assign n_13185 = ~x_2904 &  n_13141;
assign n_13186 = ~n_13184 & ~n_13185;
assign n_13187 = ~n_13136 & ~n_13186;
assign n_13188 = ~x_2840 &  n_13136;
assign n_13189 = ~n_13187 & ~n_13188;
assign n_13190 =  n_13105 & ~n_13189;
assign n_13191 = ~x_2584 & ~n_13105;
assign n_13192 = ~n_13190 & ~n_13191;
assign n_13193 =  x_2584 &  n_13192;
assign n_13194 = ~x_2584 & ~n_13192;
assign n_13195 = ~n_13193 & ~n_13194;
assign n_13196 = ~x_3029 &  n_13143;
assign n_13197 = ~x_3061 &  n_13145;
assign n_13198 = ~i_29 & ~n_13142;
assign n_13199 = ~n_13197 & ~n_13198;
assign n_13200 = ~n_13196 &  n_13199;
assign n_13201 = ~n_13141 & ~n_13200;
assign n_13202 = ~x_2903 &  n_13141;
assign n_13203 = ~n_13201 & ~n_13202;
assign n_13204 = ~n_13136 & ~n_13203;
assign n_13205 = ~x_2839 &  n_13136;
assign n_13206 = ~n_13204 & ~n_13205;
assign n_13207 =  n_13105 & ~n_13206;
assign n_13208 = ~x_2583 & ~n_13105;
assign n_13209 = ~n_13207 & ~n_13208;
assign n_13210 =  x_2583 &  n_13209;
assign n_13211 = ~x_2583 & ~n_13209;
assign n_13212 = ~n_13210 & ~n_13211;
assign n_13213 = ~x_3028 &  n_13143;
assign n_13214 = ~x_3060 &  n_13145;
assign n_13215 = ~i_28 & ~n_13142;
assign n_13216 = ~n_13214 & ~n_13215;
assign n_13217 = ~n_13213 &  n_13216;
assign n_13218 = ~n_13141 & ~n_13217;
assign n_13219 = ~x_2902 &  n_13141;
assign n_13220 = ~n_13218 & ~n_13219;
assign n_13221 = ~n_13136 & ~n_13220;
assign n_13222 = ~x_2838 &  n_13136;
assign n_13223 = ~n_13221 & ~n_13222;
assign n_13224 =  n_13105 & ~n_13223;
assign n_13225 = ~x_2582 & ~n_13105;
assign n_13226 = ~n_13224 & ~n_13225;
assign n_13227 =  x_2582 &  n_13226;
assign n_13228 = ~x_2582 & ~n_13226;
assign n_13229 = ~n_13227 & ~n_13228;
assign n_13230 =  n_2290 &  n_3615;
assign n_13231 =  n_13104 &  n_13230;
assign n_13232 =  x_1331 & ~n_13231;
assign n_13233 =  i_9 &  n_13231;
assign n_13234 = ~n_13232 & ~n_13233;
assign n_13235 =  x_1331 & ~n_13234;
assign n_13236 = ~x_1331 &  n_13234;
assign n_13237 = ~n_13235 & ~n_13236;
assign n_13238 =  x_1330 & ~n_13231;
assign n_13239 =  i_8 &  n_13231;
assign n_13240 = ~n_13238 & ~n_13239;
assign n_13241 =  x_1330 & ~n_13240;
assign n_13242 = ~x_1330 &  n_13240;
assign n_13243 = ~n_13241 & ~n_13242;
assign n_13244 =  x_1329 & ~n_13231;
assign n_13245 =  i_7 &  n_13231;
assign n_13246 = ~n_13244 & ~n_13245;
assign n_13247 =  x_1329 & ~n_13246;
assign n_13248 = ~x_1329 &  n_13246;
assign n_13249 = ~n_13247 & ~n_13248;
assign n_13250 =  x_1328 & ~n_13231;
assign n_13251 =  i_6 &  n_13231;
assign n_13252 = ~n_13250 & ~n_13251;
assign n_13253 =  x_1328 & ~n_13252;
assign n_13254 = ~x_1328 &  n_13252;
assign n_13255 = ~n_13253 & ~n_13254;
assign n_13256 =  x_1327 & ~n_13231;
assign n_13257 =  i_5 &  n_13231;
assign n_13258 = ~n_13256 & ~n_13257;
assign n_13259 =  x_1327 & ~n_13258;
assign n_13260 = ~x_1327 &  n_13258;
assign n_13261 = ~n_13259 & ~n_13260;
assign n_13262 =  x_1326 & ~n_13231;
assign n_13263 =  i_4 &  n_13231;
assign n_13264 = ~n_13262 & ~n_13263;
assign n_13265 =  x_1326 & ~n_13264;
assign n_13266 = ~x_1326 &  n_13264;
assign n_13267 = ~n_13265 & ~n_13266;
assign n_13268 =  x_1325 & ~n_13231;
assign n_13269 =  i_3 &  n_13231;
assign n_13270 = ~n_13268 & ~n_13269;
assign n_13271 =  x_1325 & ~n_13270;
assign n_13272 = ~x_1325 &  n_13270;
assign n_13273 = ~n_13271 & ~n_13272;
assign n_13274 =  x_1324 & ~n_13231;
assign n_13275 =  i_2 &  n_13231;
assign n_13276 = ~n_13274 & ~n_13275;
assign n_13277 =  x_1324 & ~n_13276;
assign n_13278 = ~x_1324 &  n_13276;
assign n_13279 = ~n_13277 & ~n_13278;
assign n_13280 =  x_1323 & ~n_13231;
assign n_13281 =  i_1 &  n_13231;
assign n_13282 = ~n_13280 & ~n_13281;
assign n_13283 =  x_1323 & ~n_13282;
assign n_13284 = ~x_1323 &  n_13282;
assign n_13285 = ~n_13283 & ~n_13284;
assign n_13286 =  n_555 &  n_13230;
assign n_13287 =  x_1322 & ~n_13286;
assign n_13288 =  i_32 &  n_13286;
assign n_13289 = ~n_13287 & ~n_13288;
assign n_13290 =  x_1322 & ~n_13289;
assign n_13291 = ~x_1322 &  n_13289;
assign n_13292 = ~n_13290 & ~n_13291;
assign n_13293 =  x_1321 & ~n_13286;
assign n_13294 =  i_31 &  n_13286;
assign n_13295 = ~n_13293 & ~n_13294;
assign n_13296 =  x_1321 & ~n_13295;
assign n_13297 = ~x_1321 &  n_13295;
assign n_13298 = ~n_13296 & ~n_13297;
assign n_13299 =  x_1320 & ~n_13286;
assign n_13300 =  i_30 &  n_13286;
assign n_13301 = ~n_13299 & ~n_13300;
assign n_13302 =  x_1320 & ~n_13301;
assign n_13303 = ~x_1320 &  n_13301;
assign n_13304 = ~n_13302 & ~n_13303;
assign n_13305 =  x_1319 & ~n_13286;
assign n_13306 =  i_29 &  n_13286;
assign n_13307 = ~n_13305 & ~n_13306;
assign n_13308 =  x_1319 & ~n_13307;
assign n_13309 = ~x_1319 &  n_13307;
assign n_13310 = ~n_13308 & ~n_13309;
assign n_13311 =  x_1318 & ~n_13286;
assign n_13312 =  i_28 &  n_13286;
assign n_13313 = ~n_13311 & ~n_13312;
assign n_13314 =  x_1318 & ~n_13313;
assign n_13315 = ~x_1318 &  n_13313;
assign n_13316 = ~n_13314 & ~n_13315;
assign n_13317 =  x_1317 & ~n_13286;
assign n_13318 =  i_27 &  n_13286;
assign n_13319 = ~n_13317 & ~n_13318;
assign n_13320 =  x_1317 & ~n_13319;
assign n_13321 = ~x_1317 &  n_13319;
assign n_13322 = ~n_13320 & ~n_13321;
assign n_13323 =  x_1316 & ~n_13286;
assign n_13324 =  i_26 &  n_13286;
assign n_13325 = ~n_13323 & ~n_13324;
assign n_13326 =  x_1316 & ~n_13325;
assign n_13327 = ~x_1316 &  n_13325;
assign n_13328 = ~n_13326 & ~n_13327;
assign n_13329 =  x_1315 & ~n_13286;
assign n_13330 =  i_25 &  n_13286;
assign n_13331 = ~n_13329 & ~n_13330;
assign n_13332 =  x_1315 & ~n_13331;
assign n_13333 = ~x_1315 &  n_13331;
assign n_13334 = ~n_13332 & ~n_13333;
assign n_13335 =  x_1314 & ~n_13286;
assign n_13336 =  i_24 &  n_13286;
assign n_13337 = ~n_13335 & ~n_13336;
assign n_13338 =  x_1314 & ~n_13337;
assign n_13339 = ~x_1314 &  n_13337;
assign n_13340 = ~n_13338 & ~n_13339;
assign n_13341 =  x_1313 & ~n_13286;
assign n_13342 =  i_23 &  n_13286;
assign n_13343 = ~n_13341 & ~n_13342;
assign n_13344 =  x_1313 & ~n_13343;
assign n_13345 = ~x_1313 &  n_13343;
assign n_13346 = ~n_13344 & ~n_13345;
assign n_13347 =  x_1312 & ~n_13286;
assign n_13348 =  i_22 &  n_13286;
assign n_13349 = ~n_13347 & ~n_13348;
assign n_13350 =  x_1312 & ~n_13349;
assign n_13351 = ~x_1312 &  n_13349;
assign n_13352 = ~n_13350 & ~n_13351;
assign n_13353 =  x_1311 & ~n_13286;
assign n_13354 =  i_21 &  n_13286;
assign n_13355 = ~n_13353 & ~n_13354;
assign n_13356 =  x_1311 & ~n_13355;
assign n_13357 = ~x_1311 &  n_13355;
assign n_13358 = ~n_13356 & ~n_13357;
assign n_13359 =  x_1310 & ~n_13286;
assign n_13360 =  i_20 &  n_13286;
assign n_13361 = ~n_13359 & ~n_13360;
assign n_13362 =  x_1310 & ~n_13361;
assign n_13363 = ~x_1310 &  n_13361;
assign n_13364 = ~n_13362 & ~n_13363;
assign n_13365 =  x_1309 & ~n_13286;
assign n_13366 =  i_19 &  n_13286;
assign n_13367 = ~n_13365 & ~n_13366;
assign n_13368 =  x_1309 & ~n_13367;
assign n_13369 = ~x_1309 &  n_13367;
assign n_13370 = ~n_13368 & ~n_13369;
assign n_13371 =  x_1308 & ~n_13286;
assign n_13372 =  i_18 &  n_13286;
assign n_13373 = ~n_13371 & ~n_13372;
assign n_13374 =  x_1308 & ~n_13373;
assign n_13375 = ~x_1308 &  n_13373;
assign n_13376 = ~n_13374 & ~n_13375;
assign n_13377 =  x_1307 & ~n_13286;
assign n_13378 =  i_17 &  n_13286;
assign n_13379 = ~n_13377 & ~n_13378;
assign n_13380 =  x_1307 & ~n_13379;
assign n_13381 = ~x_1307 &  n_13379;
assign n_13382 = ~n_13380 & ~n_13381;
assign n_13383 =  x_1306 & ~n_13286;
assign n_13384 =  i_16 &  n_13286;
assign n_13385 = ~n_13383 & ~n_13384;
assign n_13386 =  x_1306 & ~n_13385;
assign n_13387 = ~x_1306 &  n_13385;
assign n_13388 = ~n_13386 & ~n_13387;
assign n_13389 =  x_1305 & ~n_13286;
assign n_13390 =  i_15 &  n_13286;
assign n_13391 = ~n_13389 & ~n_13390;
assign n_13392 =  x_1305 & ~n_13391;
assign n_13393 = ~x_1305 &  n_13391;
assign n_13394 = ~n_13392 & ~n_13393;
assign n_13395 =  x_1304 & ~n_13286;
assign n_13396 =  i_14 &  n_13286;
assign n_13397 = ~n_13395 & ~n_13396;
assign n_13398 =  x_1304 & ~n_13397;
assign n_13399 = ~x_1304 &  n_13397;
assign n_13400 = ~n_13398 & ~n_13399;
assign n_13401 =  x_1303 & ~n_13286;
assign n_13402 =  i_13 &  n_13286;
assign n_13403 = ~n_13401 & ~n_13402;
assign n_13404 =  x_1303 & ~n_13403;
assign n_13405 = ~x_1303 &  n_13403;
assign n_13406 = ~n_13404 & ~n_13405;
assign n_13407 =  x_1302 & ~n_13286;
assign n_13408 =  i_12 &  n_13286;
assign n_13409 = ~n_13407 & ~n_13408;
assign n_13410 =  x_1302 & ~n_13409;
assign n_13411 = ~x_1302 &  n_13409;
assign n_13412 = ~n_13410 & ~n_13411;
assign n_13413 =  x_1301 & ~n_13286;
assign n_13414 =  i_11 &  n_13286;
assign n_13415 = ~n_13413 & ~n_13414;
assign n_13416 =  x_1301 & ~n_13415;
assign n_13417 = ~x_1301 &  n_13415;
assign n_13418 = ~n_13416 & ~n_13417;
assign n_13419 =  x_1300 & ~n_13286;
assign n_13420 =  i_10 &  n_13286;
assign n_13421 = ~n_13419 & ~n_13420;
assign n_13422 =  x_1300 & ~n_13421;
assign n_13423 = ~x_1300 &  n_13421;
assign n_13424 = ~n_13422 & ~n_13423;
assign n_13425 =  x_1299 & ~n_13286;
assign n_13426 =  i_9 &  n_13286;
assign n_13427 = ~n_13425 & ~n_13426;
assign n_13428 =  x_1299 & ~n_13427;
assign n_13429 = ~x_1299 &  n_13427;
assign n_13430 = ~n_13428 & ~n_13429;
assign n_13431 =  x_1298 & ~n_13286;
assign n_13432 =  i_8 &  n_13286;
assign n_13433 = ~n_13431 & ~n_13432;
assign n_13434 =  x_1298 & ~n_13433;
assign n_13435 = ~x_1298 &  n_13433;
assign n_13436 = ~n_13434 & ~n_13435;
assign n_13437 =  x_1297 & ~n_13286;
assign n_13438 =  i_7 &  n_13286;
assign n_13439 = ~n_13437 & ~n_13438;
assign n_13440 =  x_1297 & ~n_13439;
assign n_13441 = ~x_1297 &  n_13439;
assign n_13442 = ~n_13440 & ~n_13441;
assign n_13443 =  x_1296 & ~n_13286;
assign n_13444 =  i_6 &  n_13286;
assign n_13445 = ~n_13443 & ~n_13444;
assign n_13446 =  x_1296 & ~n_13445;
assign n_13447 = ~x_1296 &  n_13445;
assign n_13448 = ~n_13446 & ~n_13447;
assign n_13449 =  x_1295 & ~n_13286;
assign n_13450 =  i_5 &  n_13286;
assign n_13451 = ~n_13449 & ~n_13450;
assign n_13452 =  x_1295 & ~n_13451;
assign n_13453 = ~x_1295 &  n_13451;
assign n_13454 = ~n_13452 & ~n_13453;
assign n_13455 =  x_1294 & ~n_13286;
assign n_13456 =  i_4 &  n_13286;
assign n_13457 = ~n_13455 & ~n_13456;
assign n_13458 =  x_1294 & ~n_13457;
assign n_13459 = ~x_1294 &  n_13457;
assign n_13460 = ~n_13458 & ~n_13459;
assign n_13461 =  x_1293 & ~n_13286;
assign n_13462 =  i_3 &  n_13286;
assign n_13463 = ~n_13461 & ~n_13462;
assign n_13464 =  x_1293 & ~n_13463;
assign n_13465 = ~x_1293 &  n_13463;
assign n_13466 = ~n_13464 & ~n_13465;
assign n_13467 =  x_1292 & ~n_13286;
assign n_13468 =  i_2 &  n_13286;
assign n_13469 = ~n_13467 & ~n_13468;
assign n_13470 =  x_1292 & ~n_13469;
assign n_13471 = ~x_1292 &  n_13469;
assign n_13472 = ~n_13470 & ~n_13471;
assign n_13473 =  x_1291 & ~n_13286;
assign n_13474 =  i_1 &  n_13286;
assign n_13475 = ~n_13473 & ~n_13474;
assign n_13476 =  x_1291 & ~n_13475;
assign n_13477 = ~x_1291 &  n_13475;
assign n_13478 = ~n_13476 & ~n_13477;
assign n_13479 =  n_6525 &  n_13230;
assign n_13480 =  x_1290 & ~n_13479;
assign n_13481 =  i_32 &  n_13479;
assign n_13482 = ~n_13480 & ~n_13481;
assign n_13483 =  x_1290 & ~n_13482;
assign n_13484 = ~x_1290 &  n_13482;
assign n_13485 = ~n_13483 & ~n_13484;
assign n_13486 =  x_1289 & ~n_13479;
assign n_13487 =  i_31 &  n_13479;
assign n_13488 = ~n_13486 & ~n_13487;
assign n_13489 =  x_1289 & ~n_13488;
assign n_13490 = ~x_1289 &  n_13488;
assign n_13491 = ~n_13489 & ~n_13490;
assign n_13492 =  x_1288 & ~n_13479;
assign n_13493 =  i_30 &  n_13479;
assign n_13494 = ~n_13492 & ~n_13493;
assign n_13495 =  x_1288 & ~n_13494;
assign n_13496 = ~x_1288 &  n_13494;
assign n_13497 = ~n_13495 & ~n_13496;
assign n_13498 =  x_1287 & ~n_13479;
assign n_13499 =  i_29 &  n_13479;
assign n_13500 = ~n_13498 & ~n_13499;
assign n_13501 =  x_1287 & ~n_13500;
assign n_13502 = ~x_1287 &  n_13500;
assign n_13503 = ~n_13501 & ~n_13502;
assign n_13504 =  x_1286 & ~n_13479;
assign n_13505 =  i_28 &  n_13479;
assign n_13506 = ~n_13504 & ~n_13505;
assign n_13507 =  x_1286 & ~n_13506;
assign n_13508 = ~x_1286 &  n_13506;
assign n_13509 = ~n_13507 & ~n_13508;
assign n_13510 =  x_1285 & ~n_13479;
assign n_13511 =  i_27 &  n_13479;
assign n_13512 = ~n_13510 & ~n_13511;
assign n_13513 =  x_1285 & ~n_13512;
assign n_13514 = ~x_1285 &  n_13512;
assign n_13515 = ~n_13513 & ~n_13514;
assign n_13516 =  x_1284 & ~n_13479;
assign n_13517 =  i_26 &  n_13479;
assign n_13518 = ~n_13516 & ~n_13517;
assign n_13519 =  x_1284 & ~n_13518;
assign n_13520 = ~x_1284 &  n_13518;
assign n_13521 = ~n_13519 & ~n_13520;
assign n_13522 =  x_1283 & ~n_13479;
assign n_13523 =  i_25 &  n_13479;
assign n_13524 = ~n_13522 & ~n_13523;
assign n_13525 =  x_1283 & ~n_13524;
assign n_13526 = ~x_1283 &  n_13524;
assign n_13527 = ~n_13525 & ~n_13526;
assign n_13528 =  x_1282 & ~n_13479;
assign n_13529 =  i_24 &  n_13479;
assign n_13530 = ~n_13528 & ~n_13529;
assign n_13531 =  x_1282 & ~n_13530;
assign n_13532 = ~x_1282 &  n_13530;
assign n_13533 = ~n_13531 & ~n_13532;
assign n_13534 =  x_1281 & ~n_13479;
assign n_13535 =  i_23 &  n_13479;
assign n_13536 = ~n_13534 & ~n_13535;
assign n_13537 =  x_1281 & ~n_13536;
assign n_13538 = ~x_1281 &  n_13536;
assign n_13539 = ~n_13537 & ~n_13538;
assign n_13540 =  x_1280 & ~n_13479;
assign n_13541 =  i_22 &  n_13479;
assign n_13542 = ~n_13540 & ~n_13541;
assign n_13543 =  x_1280 & ~n_13542;
assign n_13544 = ~x_1280 &  n_13542;
assign n_13545 = ~n_13543 & ~n_13544;
assign n_13546 =  x_1279 & ~n_13479;
assign n_13547 =  i_21 &  n_13479;
assign n_13548 = ~n_13546 & ~n_13547;
assign n_13549 =  x_1279 & ~n_13548;
assign n_13550 = ~x_1279 &  n_13548;
assign n_13551 = ~n_13549 & ~n_13550;
assign n_13552 =  x_1278 & ~n_13479;
assign n_13553 =  i_20 &  n_13479;
assign n_13554 = ~n_13552 & ~n_13553;
assign n_13555 =  x_1278 & ~n_13554;
assign n_13556 = ~x_1278 &  n_13554;
assign n_13557 = ~n_13555 & ~n_13556;
assign n_13558 =  x_1277 & ~n_13479;
assign n_13559 =  i_19 &  n_13479;
assign n_13560 = ~n_13558 & ~n_13559;
assign n_13561 =  x_1277 & ~n_13560;
assign n_13562 = ~x_1277 &  n_13560;
assign n_13563 = ~n_13561 & ~n_13562;
assign n_13564 =  x_1276 & ~n_13479;
assign n_13565 =  i_18 &  n_13479;
assign n_13566 = ~n_13564 & ~n_13565;
assign n_13567 =  x_1276 & ~n_13566;
assign n_13568 = ~x_1276 &  n_13566;
assign n_13569 = ~n_13567 & ~n_13568;
assign n_13570 =  x_1275 & ~n_13479;
assign n_13571 =  i_17 &  n_13479;
assign n_13572 = ~n_13570 & ~n_13571;
assign n_13573 =  x_1275 & ~n_13572;
assign n_13574 = ~x_1275 &  n_13572;
assign n_13575 = ~n_13573 & ~n_13574;
assign n_13576 =  x_1274 & ~n_13479;
assign n_13577 =  i_16 &  n_13479;
assign n_13578 = ~n_13576 & ~n_13577;
assign n_13579 =  x_1274 & ~n_13578;
assign n_13580 = ~x_1274 &  n_13578;
assign n_13581 = ~n_13579 & ~n_13580;
assign n_13582 =  x_1273 & ~n_13479;
assign n_13583 =  i_15 &  n_13479;
assign n_13584 = ~n_13582 & ~n_13583;
assign n_13585 =  x_1273 & ~n_13584;
assign n_13586 = ~x_1273 &  n_13584;
assign n_13587 = ~n_13585 & ~n_13586;
assign n_13588 =  x_1272 & ~n_13479;
assign n_13589 =  i_14 &  n_13479;
assign n_13590 = ~n_13588 & ~n_13589;
assign n_13591 =  x_1272 & ~n_13590;
assign n_13592 = ~x_1272 &  n_13590;
assign n_13593 = ~n_13591 & ~n_13592;
assign n_13594 =  x_1271 & ~n_13479;
assign n_13595 =  i_13 &  n_13479;
assign n_13596 = ~n_13594 & ~n_13595;
assign n_13597 =  x_1271 & ~n_13596;
assign n_13598 = ~x_1271 &  n_13596;
assign n_13599 = ~n_13597 & ~n_13598;
assign n_13600 =  x_1270 & ~n_13479;
assign n_13601 =  i_12 &  n_13479;
assign n_13602 = ~n_13600 & ~n_13601;
assign n_13603 =  x_1270 & ~n_13602;
assign n_13604 = ~x_1270 &  n_13602;
assign n_13605 = ~n_13603 & ~n_13604;
assign n_13606 =  x_1269 & ~n_13479;
assign n_13607 =  i_11 &  n_13479;
assign n_13608 = ~n_13606 & ~n_13607;
assign n_13609 =  x_1269 & ~n_13608;
assign n_13610 = ~x_1269 &  n_13608;
assign n_13611 = ~n_13609 & ~n_13610;
assign n_13612 =  x_1268 & ~n_13479;
assign n_13613 =  i_10 &  n_13479;
assign n_13614 = ~n_13612 & ~n_13613;
assign n_13615 =  x_1268 & ~n_13614;
assign n_13616 = ~x_1268 &  n_13614;
assign n_13617 = ~n_13615 & ~n_13616;
assign n_13618 =  x_1267 & ~n_13479;
assign n_13619 =  i_9 &  n_13479;
assign n_13620 = ~n_13618 & ~n_13619;
assign n_13621 =  x_1267 & ~n_13620;
assign n_13622 = ~x_1267 &  n_13620;
assign n_13623 = ~n_13621 & ~n_13622;
assign n_13624 =  x_1266 & ~n_13479;
assign n_13625 =  i_8 &  n_13479;
assign n_13626 = ~n_13624 & ~n_13625;
assign n_13627 =  x_1266 & ~n_13626;
assign n_13628 = ~x_1266 &  n_13626;
assign n_13629 = ~n_13627 & ~n_13628;
assign n_13630 =  x_1265 & ~n_13479;
assign n_13631 =  i_7 &  n_13479;
assign n_13632 = ~n_13630 & ~n_13631;
assign n_13633 =  x_1265 & ~n_13632;
assign n_13634 = ~x_1265 &  n_13632;
assign n_13635 = ~n_13633 & ~n_13634;
assign n_13636 =  x_1264 & ~n_13479;
assign n_13637 =  i_6 &  n_13479;
assign n_13638 = ~n_13636 & ~n_13637;
assign n_13639 =  x_1264 & ~n_13638;
assign n_13640 = ~x_1264 &  n_13638;
assign n_13641 = ~n_13639 & ~n_13640;
assign n_13642 =  x_1263 & ~n_13479;
assign n_13643 =  i_5 &  n_13479;
assign n_13644 = ~n_13642 & ~n_13643;
assign n_13645 =  x_1263 & ~n_13644;
assign n_13646 = ~x_1263 &  n_13644;
assign n_13647 = ~n_13645 & ~n_13646;
assign n_13648 =  x_1262 & ~n_13479;
assign n_13649 =  i_4 &  n_13479;
assign n_13650 = ~n_13648 & ~n_13649;
assign n_13651 =  x_1262 & ~n_13650;
assign n_13652 = ~x_1262 &  n_13650;
assign n_13653 = ~n_13651 & ~n_13652;
assign n_13654 =  x_1261 & ~n_13479;
assign n_13655 =  i_3 &  n_13479;
assign n_13656 = ~n_13654 & ~n_13655;
assign n_13657 =  x_1261 & ~n_13656;
assign n_13658 = ~x_1261 &  n_13656;
assign n_13659 = ~n_13657 & ~n_13658;
assign n_13660 =  x_1260 & ~n_13479;
assign n_13661 =  i_2 &  n_13479;
assign n_13662 = ~n_13660 & ~n_13661;
assign n_13663 =  x_1260 & ~n_13662;
assign n_13664 = ~x_1260 &  n_13662;
assign n_13665 = ~n_13663 & ~n_13664;
assign n_13666 =  x_1259 & ~n_13479;
assign n_13667 =  i_1 &  n_13479;
assign n_13668 = ~n_13666 & ~n_13667;
assign n_13669 =  x_1259 & ~n_13668;
assign n_13670 = ~x_1259 &  n_13668;
assign n_13671 = ~n_13669 & ~n_13670;
assign n_13672 =  n_2 &  n_5651;
assign n_13673 =  n_3615 &  n_13672;
assign n_13674 =  x_1258 & ~n_13673;
assign n_13675 =  i_32 &  n_13673;
assign n_13676 = ~n_13674 & ~n_13675;
assign n_13677 =  x_1258 & ~n_13676;
assign n_13678 = ~x_1258 &  n_13676;
assign n_13679 = ~n_13677 & ~n_13678;
assign n_13680 =  x_1257 & ~n_13673;
assign n_13681 =  i_31 &  n_13673;
assign n_13682 = ~n_13680 & ~n_13681;
assign n_13683 =  x_1257 & ~n_13682;
assign n_13684 = ~x_1257 &  n_13682;
assign n_13685 = ~n_13683 & ~n_13684;
assign n_13686 =  x_1256 & ~n_13673;
assign n_13687 =  i_30 &  n_13673;
assign n_13688 = ~n_13686 & ~n_13687;
assign n_13689 =  x_1256 & ~n_13688;
assign n_13690 = ~x_1256 &  n_13688;
assign n_13691 = ~n_13689 & ~n_13690;
assign n_13692 =  x_1255 & ~n_13673;
assign n_13693 =  i_29 &  n_13673;
assign n_13694 = ~n_13692 & ~n_13693;
assign n_13695 =  x_1255 & ~n_13694;
assign n_13696 = ~x_1255 &  n_13694;
assign n_13697 = ~n_13695 & ~n_13696;
assign n_13698 =  x_1254 & ~n_13673;
assign n_13699 =  i_28 &  n_13673;
assign n_13700 = ~n_13698 & ~n_13699;
assign n_13701 =  x_1254 & ~n_13700;
assign n_13702 = ~x_1254 &  n_13700;
assign n_13703 = ~n_13701 & ~n_13702;
assign n_13704 =  x_1253 & ~n_13673;
assign n_13705 =  i_27 &  n_13673;
assign n_13706 = ~n_13704 & ~n_13705;
assign n_13707 =  x_1253 & ~n_13706;
assign n_13708 = ~x_1253 &  n_13706;
assign n_13709 = ~n_13707 & ~n_13708;
assign n_13710 =  x_1252 & ~n_13673;
assign n_13711 =  i_26 &  n_13673;
assign n_13712 = ~n_13710 & ~n_13711;
assign n_13713 =  x_1252 & ~n_13712;
assign n_13714 = ~x_1252 &  n_13712;
assign n_13715 = ~n_13713 & ~n_13714;
assign n_13716 =  x_1251 & ~n_13673;
assign n_13717 =  i_25 &  n_13673;
assign n_13718 = ~n_13716 & ~n_13717;
assign n_13719 =  x_1251 & ~n_13718;
assign n_13720 = ~x_1251 &  n_13718;
assign n_13721 = ~n_13719 & ~n_13720;
assign n_13722 =  x_1250 & ~n_13673;
assign n_13723 =  i_24 &  n_13673;
assign n_13724 = ~n_13722 & ~n_13723;
assign n_13725 =  x_1250 & ~n_13724;
assign n_13726 = ~x_1250 &  n_13724;
assign n_13727 = ~n_13725 & ~n_13726;
assign n_13728 =  x_1249 & ~n_13673;
assign n_13729 =  i_23 &  n_13673;
assign n_13730 = ~n_13728 & ~n_13729;
assign n_13731 =  x_1249 & ~n_13730;
assign n_13732 = ~x_1249 &  n_13730;
assign n_13733 = ~n_13731 & ~n_13732;
assign n_13734 =  x_1248 & ~n_13673;
assign n_13735 =  i_22 &  n_13673;
assign n_13736 = ~n_13734 & ~n_13735;
assign n_13737 =  x_1248 & ~n_13736;
assign n_13738 = ~x_1248 &  n_13736;
assign n_13739 = ~n_13737 & ~n_13738;
assign n_13740 =  x_1247 & ~n_13673;
assign n_13741 =  i_21 &  n_13673;
assign n_13742 = ~n_13740 & ~n_13741;
assign n_13743 =  x_1247 & ~n_13742;
assign n_13744 = ~x_1247 &  n_13742;
assign n_13745 = ~n_13743 & ~n_13744;
assign n_13746 =  x_1246 & ~n_13673;
assign n_13747 =  i_20 &  n_13673;
assign n_13748 = ~n_13746 & ~n_13747;
assign n_13749 =  x_1246 & ~n_13748;
assign n_13750 = ~x_1246 &  n_13748;
assign n_13751 = ~n_13749 & ~n_13750;
assign n_13752 =  x_1245 & ~n_13673;
assign n_13753 =  i_19 &  n_13673;
assign n_13754 = ~n_13752 & ~n_13753;
assign n_13755 =  x_1245 & ~n_13754;
assign n_13756 = ~x_1245 &  n_13754;
assign n_13757 = ~n_13755 & ~n_13756;
assign n_13758 =  x_1244 & ~n_13673;
assign n_13759 =  i_18 &  n_13673;
assign n_13760 = ~n_13758 & ~n_13759;
assign n_13761 =  x_1244 & ~n_13760;
assign n_13762 = ~x_1244 &  n_13760;
assign n_13763 = ~n_13761 & ~n_13762;
assign n_13764 =  x_1243 & ~n_13673;
assign n_13765 =  i_17 &  n_13673;
assign n_13766 = ~n_13764 & ~n_13765;
assign n_13767 =  x_1243 & ~n_13766;
assign n_13768 = ~x_1243 &  n_13766;
assign n_13769 = ~n_13767 & ~n_13768;
assign n_13770 =  x_1242 & ~n_13673;
assign n_13771 =  i_16 &  n_13673;
assign n_13772 = ~n_13770 & ~n_13771;
assign n_13773 =  x_1242 & ~n_13772;
assign n_13774 = ~x_1242 &  n_13772;
assign n_13775 = ~n_13773 & ~n_13774;
assign n_13776 =  x_1241 & ~n_13673;
assign n_13777 =  i_15 &  n_13673;
assign n_13778 = ~n_13776 & ~n_13777;
assign n_13779 =  x_1241 & ~n_13778;
assign n_13780 = ~x_1241 &  n_13778;
assign n_13781 = ~n_13779 & ~n_13780;
assign n_13782 =  x_1240 & ~n_13673;
assign n_13783 =  i_14 &  n_13673;
assign n_13784 = ~n_13782 & ~n_13783;
assign n_13785 =  x_1240 & ~n_13784;
assign n_13786 = ~x_1240 &  n_13784;
assign n_13787 = ~n_13785 & ~n_13786;
assign n_13788 =  x_1239 & ~n_13673;
assign n_13789 =  i_13 &  n_13673;
assign n_13790 = ~n_13788 & ~n_13789;
assign n_13791 =  x_1239 & ~n_13790;
assign n_13792 = ~x_1239 &  n_13790;
assign n_13793 = ~n_13791 & ~n_13792;
assign n_13794 =  x_1238 & ~n_13673;
assign n_13795 =  i_12 &  n_13673;
assign n_13796 = ~n_13794 & ~n_13795;
assign n_13797 =  x_1238 & ~n_13796;
assign n_13798 = ~x_1238 &  n_13796;
assign n_13799 = ~n_13797 & ~n_13798;
assign n_13800 =  x_1237 & ~n_13673;
assign n_13801 =  i_11 &  n_13673;
assign n_13802 = ~n_13800 & ~n_13801;
assign n_13803 =  x_1237 & ~n_13802;
assign n_13804 = ~x_1237 &  n_13802;
assign n_13805 = ~n_13803 & ~n_13804;
assign n_13806 =  x_1236 & ~n_13673;
assign n_13807 =  i_10 &  n_13673;
assign n_13808 = ~n_13806 & ~n_13807;
assign n_13809 =  x_1236 & ~n_13808;
assign n_13810 = ~x_1236 &  n_13808;
assign n_13811 = ~n_13809 & ~n_13810;
assign n_13812 =  x_1235 & ~n_13673;
assign n_13813 =  i_9 &  n_13673;
assign n_13814 = ~n_13812 & ~n_13813;
assign n_13815 =  x_1235 & ~n_13814;
assign n_13816 = ~x_1235 &  n_13814;
assign n_13817 = ~n_13815 & ~n_13816;
assign n_13818 =  x_1234 & ~n_13673;
assign n_13819 =  i_8 &  n_13673;
assign n_13820 = ~n_13818 & ~n_13819;
assign n_13821 =  x_1234 & ~n_13820;
assign n_13822 = ~x_1234 &  n_13820;
assign n_13823 = ~n_13821 & ~n_13822;
assign n_13824 =  x_1233 & ~n_13673;
assign n_13825 =  i_7 &  n_13673;
assign n_13826 = ~n_13824 & ~n_13825;
assign n_13827 =  x_1233 & ~n_13826;
assign n_13828 = ~x_1233 &  n_13826;
assign n_13829 = ~n_13827 & ~n_13828;
assign n_13830 =  x_1232 & ~n_13673;
assign n_13831 =  i_6 &  n_13673;
assign n_13832 = ~n_13830 & ~n_13831;
assign n_13833 =  x_1232 & ~n_13832;
assign n_13834 = ~x_1232 &  n_13832;
assign n_13835 = ~n_13833 & ~n_13834;
assign n_13836 =  x_1231 & ~n_13673;
assign n_13837 =  i_5 &  n_13673;
assign n_13838 = ~n_13836 & ~n_13837;
assign n_13839 =  x_1231 & ~n_13838;
assign n_13840 = ~x_1231 &  n_13838;
assign n_13841 = ~n_13839 & ~n_13840;
assign n_13842 =  x_1230 & ~n_13673;
assign n_13843 =  i_4 &  n_13673;
assign n_13844 = ~n_13842 & ~n_13843;
assign n_13845 =  x_1230 & ~n_13844;
assign n_13846 = ~x_1230 &  n_13844;
assign n_13847 = ~n_13845 & ~n_13846;
assign n_13848 =  x_1229 & ~n_13673;
assign n_13849 =  i_3 &  n_13673;
assign n_13850 = ~n_13848 & ~n_13849;
assign n_13851 =  x_1229 & ~n_13850;
assign n_13852 = ~x_1229 &  n_13850;
assign n_13853 = ~n_13851 & ~n_13852;
assign n_13854 =  x_1228 & ~n_13673;
assign n_13855 =  i_2 &  n_13673;
assign n_13856 = ~n_13854 & ~n_13855;
assign n_13857 =  x_1228 & ~n_13856;
assign n_13858 = ~x_1228 &  n_13856;
assign n_13859 = ~n_13857 & ~n_13858;
assign n_13860 =  x_1227 & ~n_13673;
assign n_13861 =  i_1 &  n_13673;
assign n_13862 = ~n_13860 & ~n_13861;
assign n_13863 =  x_1227 & ~n_13862;
assign n_13864 = ~x_1227 &  n_13862;
assign n_13865 = ~n_13863 & ~n_13864;
assign n_13866 =  x_38 &  n_1175;
assign n_13867 =  n_2486 &  n_13866;
assign n_13868 =  n_2291 &  n_10872;
assign n_13869 = ~n_13867 & ~n_13868;
assign n_13870 =  n_1174 &  n_2;
assign n_13871 =  n_13870 &  n_8354;
assign n_13872 =  n_3141 &  n_6181;
assign n_13873 =  n_13872 &  n_8361;
assign n_13874 = ~n_13871 & ~n_13873;
assign n_13875 =  n_13869 &  n_13874;
assign n_13876 =  x_1226 &  n_13875;
assign n_13877 =  x_4072 &  n_13873;
assign n_13878 =  x_523 &  n_13871;
assign n_13879 = ~n_13877 & ~n_13878;
assign n_13880 =  x_1898 &  n_13867;
assign n_13881 =  x_3543 &  n_13868;
assign n_13882 = ~n_13880 & ~n_13881;
assign n_13883 =  n_13879 &  n_13882;
assign n_13884 = ~n_13876 &  n_13883;
assign n_13885 =  x_1226 & ~n_13884;
assign n_13886 = ~x_1226 &  n_13884;
assign n_13887 = ~n_13885 & ~n_13886;
assign n_13888 =  x_1225 &  n_13875;
assign n_13889 =  x_4071 &  n_13873;
assign n_13890 =  x_522 &  n_13871;
assign n_13891 = ~n_13889 & ~n_13890;
assign n_13892 =  x_1897 &  n_13867;
assign n_13893 =  x_3542 &  n_13868;
assign n_13894 = ~n_13892 & ~n_13893;
assign n_13895 =  n_13891 &  n_13894;
assign n_13896 = ~n_13888 &  n_13895;
assign n_13897 =  x_1225 & ~n_13896;
assign n_13898 = ~x_1225 &  n_13896;
assign n_13899 = ~n_13897 & ~n_13898;
assign n_13900 =  x_1224 &  n_13875;
assign n_13901 =  x_4070 &  n_13873;
assign n_13902 =  x_521 &  n_13871;
assign n_13903 = ~n_13901 & ~n_13902;
assign n_13904 =  x_1896 &  n_13867;
assign n_13905 =  x_3541 &  n_13868;
assign n_13906 = ~n_13904 & ~n_13905;
assign n_13907 =  n_13903 &  n_13906;
assign n_13908 = ~n_13900 &  n_13907;
assign n_13909 =  x_1224 & ~n_13908;
assign n_13910 = ~x_1224 &  n_13908;
assign n_13911 = ~n_13909 & ~n_13910;
assign n_13912 =  x_1223 &  n_13875;
assign n_13913 =  x_4069 &  n_13873;
assign n_13914 =  x_520 &  n_13871;
assign n_13915 = ~n_13913 & ~n_13914;
assign n_13916 =  x_1895 &  n_13867;
assign n_13917 =  x_3540 &  n_13868;
assign n_13918 = ~n_13916 & ~n_13917;
assign n_13919 =  n_13915 &  n_13918;
assign n_13920 = ~n_13912 &  n_13919;
assign n_13921 =  x_1223 & ~n_13920;
assign n_13922 = ~x_1223 &  n_13920;
assign n_13923 = ~n_13921 & ~n_13922;
assign n_13924 =  x_1222 &  n_13875;
assign n_13925 =  x_4068 &  n_13873;
assign n_13926 =  x_519 &  n_13871;
assign n_13927 = ~n_13925 & ~n_13926;
assign n_13928 =  x_1894 &  n_13867;
assign n_13929 =  x_3539 &  n_13868;
assign n_13930 = ~n_13928 & ~n_13929;
assign n_13931 =  n_13927 &  n_13930;
assign n_13932 = ~n_13924 &  n_13931;
assign n_13933 =  x_1222 & ~n_13932;
assign n_13934 = ~x_1222 &  n_13932;
assign n_13935 = ~n_13933 & ~n_13934;
assign n_13936 =  x_1221 &  n_13875;
assign n_13937 =  x_4067 &  n_13873;
assign n_13938 =  x_518 &  n_13871;
assign n_13939 = ~n_13937 & ~n_13938;
assign n_13940 =  x_1893 &  n_13867;
assign n_13941 =  x_3538 &  n_13868;
assign n_13942 = ~n_13940 & ~n_13941;
assign n_13943 =  n_13939 &  n_13942;
assign n_13944 = ~n_13936 &  n_13943;
assign n_13945 =  x_1221 & ~n_13944;
assign n_13946 = ~x_1221 &  n_13944;
assign n_13947 = ~n_13945 & ~n_13946;
assign n_13948 =  x_1220 &  n_13875;
assign n_13949 =  x_4066 &  n_13873;
assign n_13950 =  x_517 &  n_13871;
assign n_13951 = ~n_13949 & ~n_13950;
assign n_13952 =  x_1892 &  n_13867;
assign n_13953 =  x_3537 &  n_13868;
assign n_13954 = ~n_13952 & ~n_13953;
assign n_13955 =  n_13951 &  n_13954;
assign n_13956 = ~n_13948 &  n_13955;
assign n_13957 =  x_1220 & ~n_13956;
assign n_13958 = ~x_1220 &  n_13956;
assign n_13959 = ~n_13957 & ~n_13958;
assign n_13960 =  x_1219 &  n_13875;
assign n_13961 =  x_4065 &  n_13873;
assign n_13962 =  x_516 &  n_13871;
assign n_13963 = ~n_13961 & ~n_13962;
assign n_13964 =  x_1891 &  n_13867;
assign n_13965 =  x_3536 &  n_13868;
assign n_13966 = ~n_13964 & ~n_13965;
assign n_13967 =  n_13963 &  n_13966;
assign n_13968 = ~n_13960 &  n_13967;
assign n_13969 =  x_1219 & ~n_13968;
assign n_13970 = ~x_1219 &  n_13968;
assign n_13971 = ~n_13969 & ~n_13970;
assign n_13972 =  x_1218 &  n_13875;
assign n_13973 =  x_4064 &  n_13873;
assign n_13974 =  x_515 &  n_13871;
assign n_13975 = ~n_13973 & ~n_13974;
assign n_13976 =  x_1890 &  n_13867;
assign n_13977 =  x_3535 &  n_13868;
assign n_13978 = ~n_13976 & ~n_13977;
assign n_13979 =  n_13975 &  n_13978;
assign n_13980 = ~n_13972 &  n_13979;
assign n_13981 =  x_1218 & ~n_13980;
assign n_13982 = ~x_1218 &  n_13980;
assign n_13983 = ~n_13981 & ~n_13982;
assign n_13984 =  x_1217 &  n_13875;
assign n_13985 =  x_4063 &  n_13873;
assign n_13986 =  x_514 &  n_13871;
assign n_13987 = ~n_13985 & ~n_13986;
assign n_13988 =  x_1889 &  n_13867;
assign n_13989 =  x_3534 &  n_13868;
assign n_13990 = ~n_13988 & ~n_13989;
assign n_13991 =  n_13987 &  n_13990;
assign n_13992 = ~n_13984 &  n_13991;
assign n_13993 =  x_1217 & ~n_13992;
assign n_13994 = ~x_1217 &  n_13992;
assign n_13995 = ~n_13993 & ~n_13994;
assign n_13996 =  x_1216 &  n_13875;
assign n_13997 =  x_4062 &  n_13873;
assign n_13998 =  x_513 &  n_13871;
assign n_13999 = ~n_13997 & ~n_13998;
assign n_14000 =  x_1888 &  n_13867;
assign n_14001 =  x_3533 &  n_13868;
assign n_14002 = ~n_14000 & ~n_14001;
assign n_14003 =  n_13999 &  n_14002;
assign n_14004 = ~n_13996 &  n_14003;
assign n_14005 =  x_1216 & ~n_14004;
assign n_14006 = ~x_1216 &  n_14004;
assign n_14007 = ~n_14005 & ~n_14006;
assign n_14008 =  x_1215 &  n_13875;
assign n_14009 =  x_4061 &  n_13873;
assign n_14010 =  x_512 &  n_13871;
assign n_14011 = ~n_14009 & ~n_14010;
assign n_14012 =  x_1887 &  n_13867;
assign n_14013 =  x_3532 &  n_13868;
assign n_14014 = ~n_14012 & ~n_14013;
assign n_14015 =  n_14011 &  n_14014;
assign n_14016 = ~n_14008 &  n_14015;
assign n_14017 =  x_1215 & ~n_14016;
assign n_14018 = ~x_1215 &  n_14016;
assign n_14019 = ~n_14017 & ~n_14018;
assign n_14020 =  x_1214 &  n_13875;
assign n_14021 =  x_4060 &  n_13873;
assign n_14022 =  x_511 &  n_13871;
assign n_14023 = ~n_14021 & ~n_14022;
assign n_14024 =  x_1886 &  n_13867;
assign n_14025 =  x_3531 &  n_13868;
assign n_14026 = ~n_14024 & ~n_14025;
assign n_14027 =  n_14023 &  n_14026;
assign n_14028 = ~n_14020 &  n_14027;
assign n_14029 =  x_1214 & ~n_14028;
assign n_14030 = ~x_1214 &  n_14028;
assign n_14031 = ~n_14029 & ~n_14030;
assign n_14032 =  x_1213 &  n_13875;
assign n_14033 =  x_4059 &  n_13873;
assign n_14034 =  x_510 &  n_13871;
assign n_14035 = ~n_14033 & ~n_14034;
assign n_14036 =  x_1885 &  n_13867;
assign n_14037 =  x_3530 &  n_13868;
assign n_14038 = ~n_14036 & ~n_14037;
assign n_14039 =  n_14035 &  n_14038;
assign n_14040 = ~n_14032 &  n_14039;
assign n_14041 =  x_1213 & ~n_14040;
assign n_14042 = ~x_1213 &  n_14040;
assign n_14043 = ~n_14041 & ~n_14042;
assign n_14044 =  x_1212 &  n_13875;
assign n_14045 =  x_4058 &  n_13873;
assign n_14046 =  x_509 &  n_13871;
assign n_14047 = ~n_14045 & ~n_14046;
assign n_14048 =  x_1884 &  n_13867;
assign n_14049 =  x_3529 &  n_13868;
assign n_14050 = ~n_14048 & ~n_14049;
assign n_14051 =  n_14047 &  n_14050;
assign n_14052 = ~n_14044 &  n_14051;
assign n_14053 =  x_1212 & ~n_14052;
assign n_14054 = ~x_1212 &  n_14052;
assign n_14055 = ~n_14053 & ~n_14054;
assign n_14056 =  x_1211 &  n_13875;
assign n_14057 =  x_4057 &  n_13873;
assign n_14058 =  x_508 &  n_13871;
assign n_14059 = ~n_14057 & ~n_14058;
assign n_14060 =  x_1883 &  n_13867;
assign n_14061 =  x_3528 &  n_13868;
assign n_14062 = ~n_14060 & ~n_14061;
assign n_14063 =  n_14059 &  n_14062;
assign n_14064 = ~n_14056 &  n_14063;
assign n_14065 =  x_1211 & ~n_14064;
assign n_14066 = ~x_1211 &  n_14064;
assign n_14067 = ~n_14065 & ~n_14066;
assign n_14068 =  x_1210 &  n_13875;
assign n_14069 =  x_4056 &  n_13873;
assign n_14070 =  x_507 &  n_13871;
assign n_14071 = ~n_14069 & ~n_14070;
assign n_14072 =  x_1882 &  n_13867;
assign n_14073 =  x_3527 &  n_13868;
assign n_14074 = ~n_14072 & ~n_14073;
assign n_14075 =  n_14071 &  n_14074;
assign n_14076 = ~n_14068 &  n_14075;
assign n_14077 =  x_1210 & ~n_14076;
assign n_14078 = ~x_1210 &  n_14076;
assign n_14079 = ~n_14077 & ~n_14078;
assign n_14080 =  x_1209 &  n_13875;
assign n_14081 =  x_4055 &  n_13873;
assign n_14082 =  x_506 &  n_13871;
assign n_14083 = ~n_14081 & ~n_14082;
assign n_14084 =  x_1881 &  n_13867;
assign n_14085 =  x_3526 &  n_13868;
assign n_14086 = ~n_14084 & ~n_14085;
assign n_14087 =  n_14083 &  n_14086;
assign n_14088 = ~n_14080 &  n_14087;
assign n_14089 =  x_1209 & ~n_14088;
assign n_14090 = ~x_1209 &  n_14088;
assign n_14091 = ~n_14089 & ~n_14090;
assign n_14092 =  x_1208 &  n_13875;
assign n_14093 =  x_4054 &  n_13873;
assign n_14094 =  x_505 &  n_13871;
assign n_14095 = ~n_14093 & ~n_14094;
assign n_14096 =  x_1880 &  n_13867;
assign n_14097 =  x_3525 &  n_13868;
assign n_14098 = ~n_14096 & ~n_14097;
assign n_14099 =  n_14095 &  n_14098;
assign n_14100 = ~n_14092 &  n_14099;
assign n_14101 =  x_1208 & ~n_14100;
assign n_14102 = ~x_1208 &  n_14100;
assign n_14103 = ~n_14101 & ~n_14102;
assign n_14104 =  x_1207 &  n_13875;
assign n_14105 =  x_4053 &  n_13873;
assign n_14106 =  x_504 &  n_13871;
assign n_14107 = ~n_14105 & ~n_14106;
assign n_14108 =  x_1879 &  n_13867;
assign n_14109 =  x_3524 &  n_13868;
assign n_14110 = ~n_14108 & ~n_14109;
assign n_14111 =  n_14107 &  n_14110;
assign n_14112 = ~n_14104 &  n_14111;
assign n_14113 =  x_1207 & ~n_14112;
assign n_14114 = ~x_1207 &  n_14112;
assign n_14115 = ~n_14113 & ~n_14114;
assign n_14116 =  x_1206 &  n_13875;
assign n_14117 =  x_4052 &  n_13873;
assign n_14118 =  x_503 &  n_13871;
assign n_14119 = ~n_14117 & ~n_14118;
assign n_14120 =  x_1878 &  n_13867;
assign n_14121 =  x_3523 &  n_13868;
assign n_14122 = ~n_14120 & ~n_14121;
assign n_14123 =  n_14119 &  n_14122;
assign n_14124 = ~n_14116 &  n_14123;
assign n_14125 =  x_1206 & ~n_14124;
assign n_14126 = ~x_1206 &  n_14124;
assign n_14127 = ~n_14125 & ~n_14126;
assign n_14128 =  x_1205 &  n_13875;
assign n_14129 =  x_4051 &  n_13873;
assign n_14130 =  x_502 &  n_13871;
assign n_14131 = ~n_14129 & ~n_14130;
assign n_14132 =  x_1877 &  n_13867;
assign n_14133 =  x_3522 &  n_13868;
assign n_14134 = ~n_14132 & ~n_14133;
assign n_14135 =  n_14131 &  n_14134;
assign n_14136 = ~n_14128 &  n_14135;
assign n_14137 =  x_1205 & ~n_14136;
assign n_14138 = ~x_1205 &  n_14136;
assign n_14139 = ~n_14137 & ~n_14138;
assign n_14140 =  x_1204 &  n_13875;
assign n_14141 =  x_4050 &  n_13873;
assign n_14142 =  x_501 &  n_13871;
assign n_14143 = ~n_14141 & ~n_14142;
assign n_14144 =  x_1876 &  n_13867;
assign n_14145 =  x_3521 &  n_13868;
assign n_14146 = ~n_14144 & ~n_14145;
assign n_14147 =  n_14143 &  n_14146;
assign n_14148 = ~n_14140 &  n_14147;
assign n_14149 =  x_1204 & ~n_14148;
assign n_14150 = ~x_1204 &  n_14148;
assign n_14151 = ~n_14149 & ~n_14150;
assign n_14152 =  x_1203 &  n_13875;
assign n_14153 =  x_4049 &  n_13873;
assign n_14154 =  x_500 &  n_13871;
assign n_14155 = ~n_14153 & ~n_14154;
assign n_14156 =  x_1875 &  n_13867;
assign n_14157 =  x_3520 &  n_13868;
assign n_14158 = ~n_14156 & ~n_14157;
assign n_14159 =  n_14155 &  n_14158;
assign n_14160 = ~n_14152 &  n_14159;
assign n_14161 =  x_1203 & ~n_14160;
assign n_14162 = ~x_1203 &  n_14160;
assign n_14163 = ~n_14161 & ~n_14162;
assign n_14164 =  x_1202 &  n_13875;
assign n_14165 =  x_4048 &  n_13873;
assign n_14166 =  x_499 &  n_13871;
assign n_14167 = ~n_14165 & ~n_14166;
assign n_14168 =  x_1874 &  n_13867;
assign n_14169 =  x_3519 &  n_13868;
assign n_14170 = ~n_14168 & ~n_14169;
assign n_14171 =  n_14167 &  n_14170;
assign n_14172 = ~n_14164 &  n_14171;
assign n_14173 =  x_1202 & ~n_14172;
assign n_14174 = ~x_1202 &  n_14172;
assign n_14175 = ~n_14173 & ~n_14174;
assign n_14176 =  x_1201 &  n_13875;
assign n_14177 =  x_4047 &  n_13873;
assign n_14178 =  x_498 &  n_13871;
assign n_14179 = ~n_14177 & ~n_14178;
assign n_14180 =  x_1873 &  n_13867;
assign n_14181 =  x_3518 &  n_13868;
assign n_14182 = ~n_14180 & ~n_14181;
assign n_14183 =  n_14179 &  n_14182;
assign n_14184 = ~n_14176 &  n_14183;
assign n_14185 =  x_1201 & ~n_14184;
assign n_14186 = ~x_1201 &  n_14184;
assign n_14187 = ~n_14185 & ~n_14186;
assign n_14188 =  x_1200 &  n_13875;
assign n_14189 =  x_4046 &  n_13873;
assign n_14190 =  x_497 &  n_13871;
assign n_14191 = ~n_14189 & ~n_14190;
assign n_14192 =  x_1872 &  n_13867;
assign n_14193 =  x_3517 &  n_13868;
assign n_14194 = ~n_14192 & ~n_14193;
assign n_14195 =  n_14191 &  n_14194;
assign n_14196 = ~n_14188 &  n_14195;
assign n_14197 =  x_1200 & ~n_14196;
assign n_14198 = ~x_1200 &  n_14196;
assign n_14199 = ~n_14197 & ~n_14198;
assign n_14200 =  x_1199 &  n_13875;
assign n_14201 =  x_4045 &  n_13873;
assign n_14202 =  x_496 &  n_13871;
assign n_14203 = ~n_14201 & ~n_14202;
assign n_14204 =  x_1871 &  n_13867;
assign n_14205 =  x_3516 &  n_13868;
assign n_14206 = ~n_14204 & ~n_14205;
assign n_14207 =  n_14203 &  n_14206;
assign n_14208 = ~n_14200 &  n_14207;
assign n_14209 =  x_1199 & ~n_14208;
assign n_14210 = ~x_1199 &  n_14208;
assign n_14211 = ~n_14209 & ~n_14210;
assign n_14212 =  x_1198 &  n_13875;
assign n_14213 =  x_4044 &  n_13873;
assign n_14214 =  x_495 &  n_13871;
assign n_14215 = ~n_14213 & ~n_14214;
assign n_14216 =  x_1870 &  n_13867;
assign n_14217 =  x_3515 &  n_13868;
assign n_14218 = ~n_14216 & ~n_14217;
assign n_14219 =  n_14215 &  n_14218;
assign n_14220 = ~n_14212 &  n_14219;
assign n_14221 =  x_1198 & ~n_14220;
assign n_14222 = ~x_1198 &  n_14220;
assign n_14223 = ~n_14221 & ~n_14222;
assign n_14224 =  x_1197 &  n_13875;
assign n_14225 =  x_4043 &  n_13873;
assign n_14226 =  x_494 &  n_13871;
assign n_14227 = ~n_14225 & ~n_14226;
assign n_14228 =  x_1869 &  n_13867;
assign n_14229 =  x_3514 &  n_13868;
assign n_14230 = ~n_14228 & ~n_14229;
assign n_14231 =  n_14227 &  n_14230;
assign n_14232 = ~n_14224 &  n_14231;
assign n_14233 =  x_1197 & ~n_14232;
assign n_14234 = ~x_1197 &  n_14232;
assign n_14235 = ~n_14233 & ~n_14234;
assign n_14236 =  x_1196 &  n_13875;
assign n_14237 =  x_4042 &  n_13873;
assign n_14238 =  x_493 &  n_13871;
assign n_14239 = ~n_14237 & ~n_14238;
assign n_14240 =  x_1868 &  n_13867;
assign n_14241 =  x_3513 &  n_13868;
assign n_14242 = ~n_14240 & ~n_14241;
assign n_14243 =  n_14239 &  n_14242;
assign n_14244 = ~n_14236 &  n_14243;
assign n_14245 =  x_1196 & ~n_14244;
assign n_14246 = ~x_1196 &  n_14244;
assign n_14247 = ~n_14245 & ~n_14246;
assign n_14248 =  x_1195 &  n_13875;
assign n_14249 =  x_4041 &  n_13873;
assign n_14250 =  x_492 &  n_13871;
assign n_14251 = ~n_14249 & ~n_14250;
assign n_14252 =  x_1867 &  n_13867;
assign n_14253 =  x_3512 &  n_13868;
assign n_14254 = ~n_14252 & ~n_14253;
assign n_14255 =  n_14251 &  n_14254;
assign n_14256 = ~n_14248 &  n_14255;
assign n_14257 =  x_1195 & ~n_14256;
assign n_14258 = ~x_1195 &  n_14256;
assign n_14259 = ~n_14257 & ~n_14258;
assign n_14260 =  n_6378 &  n_2486;
assign n_14261 =  n_2682 &  n_8354;
assign n_14262 = ~n_14260 & ~n_14261;
assign n_14263 =  n_349 &  n_8352;
assign n_14264 =  x_38 &  n_14263;
assign n_14265 =  n_2486 &  n_14264;
assign n_14266 =  n_3341 &  n_5648;
assign n_14267 =  n_2486 &  n_14266;
assign n_14268 = ~x_43 &  n_14267;
assign n_14269 = ~n_14265 & ~n_14268;
assign n_14270 =  n_14262 &  n_14269;
assign n_14271 =  x_1194 &  n_14270;
assign n_14272 =  x_3976 &  n_14268;
assign n_14273 =  x_1866 &  n_14261;
assign n_14274 = ~n_14272 & ~n_14273;
assign n_14275 =  x_3511 &  n_14265;
assign n_14276 =  x_363 &  n_14260;
assign n_14277 = ~n_14275 & ~n_14276;
assign n_14278 =  n_14274 &  n_14277;
assign n_14279 = ~n_14271 &  n_14278;
assign n_14280 =  x_1194 & ~n_14279;
assign n_14281 = ~x_1194 &  n_14279;
assign n_14282 = ~n_14280 & ~n_14281;
assign n_14283 =  x_1193 &  n_14270;
assign n_14284 =  x_3975 &  n_14268;
assign n_14285 =  x_1865 &  n_14261;
assign n_14286 = ~n_14284 & ~n_14285;
assign n_14287 =  x_3510 &  n_14265;
assign n_14288 =  x_362 &  n_14260;
assign n_14289 = ~n_14287 & ~n_14288;
assign n_14290 =  n_14286 &  n_14289;
assign n_14291 = ~n_14283 &  n_14290;
assign n_14292 =  x_1193 & ~n_14291;
assign n_14293 = ~x_1193 &  n_14291;
assign n_14294 = ~n_14292 & ~n_14293;
assign n_14295 =  x_1192 &  n_14270;
assign n_14296 =  x_3974 &  n_14268;
assign n_14297 =  x_1864 &  n_14261;
assign n_14298 = ~n_14296 & ~n_14297;
assign n_14299 =  x_3509 &  n_14265;
assign n_14300 =  x_361 &  n_14260;
assign n_14301 = ~n_14299 & ~n_14300;
assign n_14302 =  n_14298 &  n_14301;
assign n_14303 = ~n_14295 &  n_14302;
assign n_14304 =  x_1192 & ~n_14303;
assign n_14305 = ~x_1192 &  n_14303;
assign n_14306 = ~n_14304 & ~n_14305;
assign n_14307 =  x_1191 &  n_14270;
assign n_14308 =  x_3973 &  n_14268;
assign n_14309 =  x_1863 &  n_14261;
assign n_14310 = ~n_14308 & ~n_14309;
assign n_14311 =  x_3508 &  n_14265;
assign n_14312 =  x_360 &  n_14260;
assign n_14313 = ~n_14311 & ~n_14312;
assign n_14314 =  n_14310 &  n_14313;
assign n_14315 = ~n_14307 &  n_14314;
assign n_14316 =  x_1191 & ~n_14315;
assign n_14317 = ~x_1191 &  n_14315;
assign n_14318 = ~n_14316 & ~n_14317;
assign n_14319 =  x_1190 &  n_14270;
assign n_14320 =  x_3972 &  n_14268;
assign n_14321 =  x_1862 &  n_14261;
assign n_14322 = ~n_14320 & ~n_14321;
assign n_14323 =  x_3507 &  n_14265;
assign n_14324 =  x_359 &  n_14260;
assign n_14325 = ~n_14323 & ~n_14324;
assign n_14326 =  n_14322 &  n_14325;
assign n_14327 = ~n_14319 &  n_14326;
assign n_14328 =  x_1190 & ~n_14327;
assign n_14329 = ~x_1190 &  n_14327;
assign n_14330 = ~n_14328 & ~n_14329;
assign n_14331 =  x_1189 &  n_14270;
assign n_14332 =  x_3971 &  n_14268;
assign n_14333 =  x_1861 &  n_14261;
assign n_14334 = ~n_14332 & ~n_14333;
assign n_14335 =  x_3506 &  n_14265;
assign n_14336 =  x_358 &  n_14260;
assign n_14337 = ~n_14335 & ~n_14336;
assign n_14338 =  n_14334 &  n_14337;
assign n_14339 = ~n_14331 &  n_14338;
assign n_14340 =  x_1189 & ~n_14339;
assign n_14341 = ~x_1189 &  n_14339;
assign n_14342 = ~n_14340 & ~n_14341;
assign n_14343 =  x_1188 &  n_14270;
assign n_14344 =  x_3970 &  n_14268;
assign n_14345 =  x_1860 &  n_14261;
assign n_14346 = ~n_14344 & ~n_14345;
assign n_14347 =  x_3505 &  n_14265;
assign n_14348 =  x_357 &  n_14260;
assign n_14349 = ~n_14347 & ~n_14348;
assign n_14350 =  n_14346 &  n_14349;
assign n_14351 = ~n_14343 &  n_14350;
assign n_14352 =  x_1188 & ~n_14351;
assign n_14353 = ~x_1188 &  n_14351;
assign n_14354 = ~n_14352 & ~n_14353;
assign n_14355 =  x_1187 &  n_14270;
assign n_14356 =  x_3969 &  n_14268;
assign n_14357 =  x_1859 &  n_14261;
assign n_14358 = ~n_14356 & ~n_14357;
assign n_14359 =  x_3504 &  n_14265;
assign n_14360 =  x_356 &  n_14260;
assign n_14361 = ~n_14359 & ~n_14360;
assign n_14362 =  n_14358 &  n_14361;
assign n_14363 = ~n_14355 &  n_14362;
assign n_14364 =  x_1187 & ~n_14363;
assign n_14365 = ~x_1187 &  n_14363;
assign n_14366 = ~n_14364 & ~n_14365;
assign n_14367 =  x_1186 &  n_14270;
assign n_14368 =  x_3968 &  n_14268;
assign n_14369 =  x_1858 &  n_14261;
assign n_14370 = ~n_14368 & ~n_14369;
assign n_14371 =  x_3503 &  n_14265;
assign n_14372 =  x_355 &  n_14260;
assign n_14373 = ~n_14371 & ~n_14372;
assign n_14374 =  n_14370 &  n_14373;
assign n_14375 = ~n_14367 &  n_14374;
assign n_14376 =  x_1186 & ~n_14375;
assign n_14377 = ~x_1186 &  n_14375;
assign n_14378 = ~n_14376 & ~n_14377;
assign n_14379 =  x_1185 &  n_14270;
assign n_14380 =  x_3967 &  n_14268;
assign n_14381 =  x_1857 &  n_14261;
assign n_14382 = ~n_14380 & ~n_14381;
assign n_14383 =  x_3502 &  n_14265;
assign n_14384 =  x_354 &  n_14260;
assign n_14385 = ~n_14383 & ~n_14384;
assign n_14386 =  n_14382 &  n_14385;
assign n_14387 = ~n_14379 &  n_14386;
assign n_14388 =  x_1185 & ~n_14387;
assign n_14389 = ~x_1185 &  n_14387;
assign n_14390 = ~n_14388 & ~n_14389;
assign n_14391 =  x_1184 &  n_14270;
assign n_14392 =  x_3966 &  n_14268;
assign n_14393 =  x_1856 &  n_14261;
assign n_14394 = ~n_14392 & ~n_14393;
assign n_14395 =  x_3501 &  n_14265;
assign n_14396 =  x_353 &  n_14260;
assign n_14397 = ~n_14395 & ~n_14396;
assign n_14398 =  n_14394 &  n_14397;
assign n_14399 = ~n_14391 &  n_14398;
assign n_14400 =  x_1184 & ~n_14399;
assign n_14401 = ~x_1184 &  n_14399;
assign n_14402 = ~n_14400 & ~n_14401;
assign n_14403 =  x_1183 &  n_14270;
assign n_14404 =  x_3965 &  n_14268;
assign n_14405 =  x_1855 &  n_14261;
assign n_14406 = ~n_14404 & ~n_14405;
assign n_14407 =  x_3500 &  n_14265;
assign n_14408 =  x_352 &  n_14260;
assign n_14409 = ~n_14407 & ~n_14408;
assign n_14410 =  n_14406 &  n_14409;
assign n_14411 = ~n_14403 &  n_14410;
assign n_14412 =  x_1183 & ~n_14411;
assign n_14413 = ~x_1183 &  n_14411;
assign n_14414 = ~n_14412 & ~n_14413;
assign n_14415 =  x_1182 &  n_14270;
assign n_14416 =  x_3964 &  n_14268;
assign n_14417 =  x_1854 &  n_14261;
assign n_14418 = ~n_14416 & ~n_14417;
assign n_14419 =  x_3499 &  n_14265;
assign n_14420 =  x_351 &  n_14260;
assign n_14421 = ~n_14419 & ~n_14420;
assign n_14422 =  n_14418 &  n_14421;
assign n_14423 = ~n_14415 &  n_14422;
assign n_14424 =  x_1182 & ~n_14423;
assign n_14425 = ~x_1182 &  n_14423;
assign n_14426 = ~n_14424 & ~n_14425;
assign n_14427 =  x_1181 &  n_14270;
assign n_14428 =  x_3963 &  n_14268;
assign n_14429 =  x_1853 &  n_14261;
assign n_14430 = ~n_14428 & ~n_14429;
assign n_14431 =  x_3498 &  n_14265;
assign n_14432 =  x_350 &  n_14260;
assign n_14433 = ~n_14431 & ~n_14432;
assign n_14434 =  n_14430 &  n_14433;
assign n_14435 = ~n_14427 &  n_14434;
assign n_14436 =  x_1181 & ~n_14435;
assign n_14437 = ~x_1181 &  n_14435;
assign n_14438 = ~n_14436 & ~n_14437;
assign n_14439 =  x_1180 &  n_14270;
assign n_14440 =  x_3962 &  n_14268;
assign n_14441 =  x_1852 &  n_14261;
assign n_14442 = ~n_14440 & ~n_14441;
assign n_14443 =  x_3497 &  n_14265;
assign n_14444 =  x_349 &  n_14260;
assign n_14445 = ~n_14443 & ~n_14444;
assign n_14446 =  n_14442 &  n_14445;
assign n_14447 = ~n_14439 &  n_14446;
assign n_14448 =  x_1180 & ~n_14447;
assign n_14449 = ~x_1180 &  n_14447;
assign n_14450 = ~n_14448 & ~n_14449;
assign n_14451 =  x_1179 &  n_14270;
assign n_14452 =  x_3961 &  n_14268;
assign n_14453 =  x_1851 &  n_14261;
assign n_14454 = ~n_14452 & ~n_14453;
assign n_14455 =  x_3496 &  n_14265;
assign n_14456 =  x_348 &  n_14260;
assign n_14457 = ~n_14455 & ~n_14456;
assign n_14458 =  n_14454 &  n_14457;
assign n_14459 = ~n_14451 &  n_14458;
assign n_14460 =  x_1179 & ~n_14459;
assign n_14461 = ~x_1179 &  n_14459;
assign n_14462 = ~n_14460 & ~n_14461;
assign n_14463 =  x_1178 &  n_14270;
assign n_14464 =  x_3960 &  n_14268;
assign n_14465 =  x_1850 &  n_14261;
assign n_14466 = ~n_14464 & ~n_14465;
assign n_14467 =  x_3495 &  n_14265;
assign n_14468 =  x_347 &  n_14260;
assign n_14469 = ~n_14467 & ~n_14468;
assign n_14470 =  n_14466 &  n_14469;
assign n_14471 = ~n_14463 &  n_14470;
assign n_14472 =  x_1178 & ~n_14471;
assign n_14473 = ~x_1178 &  n_14471;
assign n_14474 = ~n_14472 & ~n_14473;
assign n_14475 =  x_1177 &  n_14270;
assign n_14476 =  x_3959 &  n_14268;
assign n_14477 =  x_1849 &  n_14261;
assign n_14478 = ~n_14476 & ~n_14477;
assign n_14479 =  x_3494 &  n_14265;
assign n_14480 =  x_346 &  n_14260;
assign n_14481 = ~n_14479 & ~n_14480;
assign n_14482 =  n_14478 &  n_14481;
assign n_14483 = ~n_14475 &  n_14482;
assign n_14484 =  x_1177 & ~n_14483;
assign n_14485 = ~x_1177 &  n_14483;
assign n_14486 = ~n_14484 & ~n_14485;
assign n_14487 =  x_1176 &  n_14270;
assign n_14488 =  x_3958 &  n_14268;
assign n_14489 =  x_1848 &  n_14261;
assign n_14490 = ~n_14488 & ~n_14489;
assign n_14491 =  x_3493 &  n_14265;
assign n_14492 =  x_345 &  n_14260;
assign n_14493 = ~n_14491 & ~n_14492;
assign n_14494 =  n_14490 &  n_14493;
assign n_14495 = ~n_14487 &  n_14494;
assign n_14496 =  x_1176 & ~n_14495;
assign n_14497 = ~x_1176 &  n_14495;
assign n_14498 = ~n_14496 & ~n_14497;
assign n_14499 =  x_1175 &  n_14270;
assign n_14500 =  x_3957 &  n_14268;
assign n_14501 =  x_1847 &  n_14261;
assign n_14502 = ~n_14500 & ~n_14501;
assign n_14503 =  x_3492 &  n_14265;
assign n_14504 =  x_344 &  n_14260;
assign n_14505 = ~n_14503 & ~n_14504;
assign n_14506 =  n_14502 &  n_14505;
assign n_14507 = ~n_14499 &  n_14506;
assign n_14508 =  x_1175 & ~n_14507;
assign n_14509 = ~x_1175 &  n_14507;
assign n_14510 = ~n_14508 & ~n_14509;
assign n_14511 =  x_1174 &  n_14270;
assign n_14512 =  x_3956 &  n_14268;
assign n_14513 =  x_1846 &  n_14261;
assign n_14514 = ~n_14512 & ~n_14513;
assign n_14515 =  x_3491 &  n_14265;
assign n_14516 =  x_343 &  n_14260;
assign n_14517 = ~n_14515 & ~n_14516;
assign n_14518 =  n_14514 &  n_14517;
assign n_14519 = ~n_14511 &  n_14518;
assign n_14520 =  x_1174 & ~n_14519;
assign n_14521 = ~x_1174 &  n_14519;
assign n_14522 = ~n_14520 & ~n_14521;
assign n_14523 =  x_1173 &  n_14270;
assign n_14524 =  x_3955 &  n_14268;
assign n_14525 =  x_1845 &  n_14261;
assign n_14526 = ~n_14524 & ~n_14525;
assign n_14527 =  x_3490 &  n_14265;
assign n_14528 =  x_342 &  n_14260;
assign n_14529 = ~n_14527 & ~n_14528;
assign n_14530 =  n_14526 &  n_14529;
assign n_14531 = ~n_14523 &  n_14530;
assign n_14532 =  x_1173 & ~n_14531;
assign n_14533 = ~x_1173 &  n_14531;
assign n_14534 = ~n_14532 & ~n_14533;
assign n_14535 =  x_1172 &  n_14270;
assign n_14536 =  x_3954 &  n_14268;
assign n_14537 =  x_1844 &  n_14261;
assign n_14538 = ~n_14536 & ~n_14537;
assign n_14539 =  x_3489 &  n_14265;
assign n_14540 =  x_341 &  n_14260;
assign n_14541 = ~n_14539 & ~n_14540;
assign n_14542 =  n_14538 &  n_14541;
assign n_14543 = ~n_14535 &  n_14542;
assign n_14544 =  x_1172 & ~n_14543;
assign n_14545 = ~x_1172 &  n_14543;
assign n_14546 = ~n_14544 & ~n_14545;
assign n_14547 =  x_1171 &  n_14270;
assign n_14548 =  x_3953 &  n_14268;
assign n_14549 =  x_1843 &  n_14261;
assign n_14550 = ~n_14548 & ~n_14549;
assign n_14551 =  x_3488 &  n_14265;
assign n_14552 =  x_340 &  n_14260;
assign n_14553 = ~n_14551 & ~n_14552;
assign n_14554 =  n_14550 &  n_14553;
assign n_14555 = ~n_14547 &  n_14554;
assign n_14556 =  x_1171 & ~n_14555;
assign n_14557 = ~x_1171 &  n_14555;
assign n_14558 = ~n_14556 & ~n_14557;
assign n_14559 =  x_1170 &  n_14270;
assign n_14560 =  x_3952 &  n_14268;
assign n_14561 =  x_1842 &  n_14261;
assign n_14562 = ~n_14560 & ~n_14561;
assign n_14563 =  x_3487 &  n_14265;
assign n_14564 =  x_339 &  n_14260;
assign n_14565 = ~n_14563 & ~n_14564;
assign n_14566 =  n_14562 &  n_14565;
assign n_14567 = ~n_14559 &  n_14566;
assign n_14568 =  x_1170 & ~n_14567;
assign n_14569 = ~x_1170 &  n_14567;
assign n_14570 = ~n_14568 & ~n_14569;
assign n_14571 =  x_1169 &  n_14270;
assign n_14572 =  x_3951 &  n_14268;
assign n_14573 =  x_1841 &  n_14261;
assign n_14574 = ~n_14572 & ~n_14573;
assign n_14575 =  x_3486 &  n_14265;
assign n_14576 =  x_338 &  n_14260;
assign n_14577 = ~n_14575 & ~n_14576;
assign n_14578 =  n_14574 &  n_14577;
assign n_14579 = ~n_14571 &  n_14578;
assign n_14580 =  x_1169 & ~n_14579;
assign n_14581 = ~x_1169 &  n_14579;
assign n_14582 = ~n_14580 & ~n_14581;
assign n_14583 =  x_1168 &  n_14270;
assign n_14584 =  x_3950 &  n_14268;
assign n_14585 =  x_1840 &  n_14261;
assign n_14586 = ~n_14584 & ~n_14585;
assign n_14587 =  x_3485 &  n_14265;
assign n_14588 =  x_337 &  n_14260;
assign n_14589 = ~n_14587 & ~n_14588;
assign n_14590 =  n_14586 &  n_14589;
assign n_14591 = ~n_14583 &  n_14590;
assign n_14592 =  x_1168 & ~n_14591;
assign n_14593 = ~x_1168 &  n_14591;
assign n_14594 = ~n_14592 & ~n_14593;
assign n_14595 =  x_1167 &  n_14270;
assign n_14596 =  x_3949 &  n_14268;
assign n_14597 =  x_1839 &  n_14261;
assign n_14598 = ~n_14596 & ~n_14597;
assign n_14599 =  x_3484 &  n_14265;
assign n_14600 =  x_336 &  n_14260;
assign n_14601 = ~n_14599 & ~n_14600;
assign n_14602 =  n_14598 &  n_14601;
assign n_14603 = ~n_14595 &  n_14602;
assign n_14604 =  x_1167 & ~n_14603;
assign n_14605 = ~x_1167 &  n_14603;
assign n_14606 = ~n_14604 & ~n_14605;
assign n_14607 =  x_1166 &  n_14270;
assign n_14608 =  x_3948 &  n_14268;
assign n_14609 =  x_1838 &  n_14261;
assign n_14610 = ~n_14608 & ~n_14609;
assign n_14611 =  x_3483 &  n_14265;
assign n_14612 =  x_335 &  n_14260;
assign n_14613 = ~n_14611 & ~n_14612;
assign n_14614 =  n_14610 &  n_14613;
assign n_14615 = ~n_14607 &  n_14614;
assign n_14616 =  x_1166 & ~n_14615;
assign n_14617 = ~x_1166 &  n_14615;
assign n_14618 = ~n_14616 & ~n_14617;
assign n_14619 =  x_1165 &  n_14270;
assign n_14620 =  x_3947 &  n_14268;
assign n_14621 =  x_1837 &  n_14261;
assign n_14622 = ~n_14620 & ~n_14621;
assign n_14623 =  x_3482 &  n_14265;
assign n_14624 =  x_334 &  n_14260;
assign n_14625 = ~n_14623 & ~n_14624;
assign n_14626 =  n_14622 &  n_14625;
assign n_14627 = ~n_14619 &  n_14626;
assign n_14628 =  x_1165 & ~n_14627;
assign n_14629 = ~x_1165 &  n_14627;
assign n_14630 = ~n_14628 & ~n_14629;
assign n_14631 =  x_1164 &  n_14270;
assign n_14632 =  x_3946 &  n_14268;
assign n_14633 =  x_1836 &  n_14261;
assign n_14634 = ~n_14632 & ~n_14633;
assign n_14635 =  x_3481 &  n_14265;
assign n_14636 =  x_333 &  n_14260;
assign n_14637 = ~n_14635 & ~n_14636;
assign n_14638 =  n_14634 &  n_14637;
assign n_14639 = ~n_14631 &  n_14638;
assign n_14640 =  x_1164 & ~n_14639;
assign n_14641 = ~x_1164 &  n_14639;
assign n_14642 = ~n_14640 & ~n_14641;
assign n_14643 =  x_1163 &  n_14270;
assign n_14644 =  x_3945 &  n_14268;
assign n_14645 =  x_1835 &  n_14261;
assign n_14646 = ~n_14644 & ~n_14645;
assign n_14647 =  x_3480 &  n_14265;
assign n_14648 =  x_332 &  n_14260;
assign n_14649 = ~n_14647 & ~n_14648;
assign n_14650 =  n_14646 &  n_14649;
assign n_14651 = ~n_14643 &  n_14650;
assign n_14652 =  x_1163 & ~n_14651;
assign n_14653 = ~x_1163 &  n_14651;
assign n_14654 = ~n_14652 & ~n_14653;
assign n_14655 =  n_759 &  n_4290;
assign n_14656 =  n_1038 &  n_14655;
assign n_14657 =  x_1162 & ~n_14656;
assign n_14658 =  x_1162 &  n_14657;
assign n_14659 = ~x_1162 & ~n_14657;
assign n_14660 = ~n_14658 & ~n_14659;
assign n_14661 =  x_1161 & ~n_14656;
assign n_14662 =  x_1161 &  n_14661;
assign n_14663 = ~x_1161 & ~n_14661;
assign n_14664 = ~n_14662 & ~n_14663;
assign n_14665 =  x_1160 & ~n_14656;
assign n_14666 =  x_1160 &  n_14665;
assign n_14667 = ~x_1160 & ~n_14665;
assign n_14668 = ~n_14666 & ~n_14667;
assign n_14669 =  x_1159 & ~n_14656;
assign n_14670 =  x_1159 &  n_14669;
assign n_14671 = ~x_1159 & ~n_14669;
assign n_14672 = ~n_14670 & ~n_14671;
assign n_14673 =  x_1158 & ~n_14656;
assign n_14674 =  x_1158 &  n_14673;
assign n_14675 = ~x_1158 & ~n_14673;
assign n_14676 = ~n_14674 & ~n_14675;
assign n_14677 =  x_1157 & ~n_14656;
assign n_14678 =  x_1157 &  n_14677;
assign n_14679 = ~x_1157 & ~n_14677;
assign n_14680 = ~n_14678 & ~n_14679;
assign n_14681 =  x_1156 & ~n_14656;
assign n_14682 =  x_1156 &  n_14681;
assign n_14683 = ~x_1156 & ~n_14681;
assign n_14684 = ~n_14682 & ~n_14683;
assign n_14685 =  x_1155 & ~n_14656;
assign n_14686 =  x_1155 &  n_14685;
assign n_14687 = ~x_1155 & ~n_14685;
assign n_14688 = ~n_14686 & ~n_14687;
assign n_14689 =  x_1154 & ~n_14656;
assign n_14690 =  x_1154 &  n_14689;
assign n_14691 = ~x_1154 & ~n_14689;
assign n_14692 = ~n_14690 & ~n_14691;
assign n_14693 =  x_1153 & ~n_14656;
assign n_14694 =  x_1153 &  n_14693;
assign n_14695 = ~x_1153 & ~n_14693;
assign n_14696 = ~n_14694 & ~n_14695;
assign n_14697 =  x_1152 & ~n_14656;
assign n_14698 =  x_1152 &  n_14697;
assign n_14699 = ~x_1152 & ~n_14697;
assign n_14700 = ~n_14698 & ~n_14699;
assign n_14701 =  x_1151 & ~n_14656;
assign n_14702 =  x_1151 &  n_14701;
assign n_14703 = ~x_1151 & ~n_14701;
assign n_14704 = ~n_14702 & ~n_14703;
assign n_14705 =  x_1150 & ~n_14656;
assign n_14706 =  x_1150 &  n_14705;
assign n_14707 = ~x_1150 & ~n_14705;
assign n_14708 = ~n_14706 & ~n_14707;
assign n_14709 =  x_1149 & ~n_14656;
assign n_14710 =  x_1149 &  n_14709;
assign n_14711 = ~x_1149 & ~n_14709;
assign n_14712 = ~n_14710 & ~n_14711;
assign n_14713 =  x_1148 & ~n_14656;
assign n_14714 =  x_1148 &  n_14713;
assign n_14715 = ~x_1148 & ~n_14713;
assign n_14716 = ~n_14714 & ~n_14715;
assign n_14717 =  x_1147 & ~n_14656;
assign n_14718 =  x_1147 &  n_14717;
assign n_14719 = ~x_1147 & ~n_14717;
assign n_14720 = ~n_14718 & ~n_14719;
assign n_14721 =  x_1146 & ~n_14656;
assign n_14722 =  x_1146 &  n_14721;
assign n_14723 = ~x_1146 & ~n_14721;
assign n_14724 = ~n_14722 & ~n_14723;
assign n_14725 =  x_1145 & ~n_14656;
assign n_14726 =  x_1145 &  n_14725;
assign n_14727 = ~x_1145 & ~n_14725;
assign n_14728 = ~n_14726 & ~n_14727;
assign n_14729 =  x_1144 & ~n_14656;
assign n_14730 =  x_1144 &  n_14729;
assign n_14731 = ~x_1144 & ~n_14729;
assign n_14732 = ~n_14730 & ~n_14731;
assign n_14733 =  x_1143 & ~n_14656;
assign n_14734 =  x_1143 &  n_14733;
assign n_14735 = ~x_1143 & ~n_14733;
assign n_14736 = ~n_14734 & ~n_14735;
assign n_14737 =  x_1142 & ~n_14656;
assign n_14738 =  x_1142 &  n_14737;
assign n_14739 = ~x_1142 & ~n_14737;
assign n_14740 = ~n_14738 & ~n_14739;
assign n_14741 =  x_1141 & ~n_14656;
assign n_14742 =  x_1141 &  n_14741;
assign n_14743 = ~x_1141 & ~n_14741;
assign n_14744 = ~n_14742 & ~n_14743;
assign n_14745 =  x_1140 & ~n_14656;
assign n_14746 =  x_1140 &  n_14745;
assign n_14747 = ~x_1140 & ~n_14745;
assign n_14748 = ~n_14746 & ~n_14747;
assign n_14749 =  x_1139 & ~n_14656;
assign n_14750 =  x_1139 &  n_14749;
assign n_14751 = ~x_1139 & ~n_14749;
assign n_14752 = ~n_14750 & ~n_14751;
assign n_14753 =  x_1138 & ~n_14656;
assign n_14754 =  x_1138 &  n_14753;
assign n_14755 = ~x_1138 & ~n_14753;
assign n_14756 = ~n_14754 & ~n_14755;
assign n_14757 =  x_1137 & ~n_14656;
assign n_14758 =  x_1137 &  n_14757;
assign n_14759 = ~x_1137 & ~n_14757;
assign n_14760 = ~n_14758 & ~n_14759;
assign n_14761 =  x_1136 & ~n_14656;
assign n_14762 =  x_1136 &  n_14761;
assign n_14763 = ~x_1136 & ~n_14761;
assign n_14764 = ~n_14762 & ~n_14763;
assign n_14765 =  x_1135 & ~n_14656;
assign n_14766 =  x_1135 &  n_14765;
assign n_14767 = ~x_1135 & ~n_14765;
assign n_14768 = ~n_14766 & ~n_14767;
assign n_14769 =  x_1134 & ~n_14656;
assign n_14770 =  x_1134 &  n_14769;
assign n_14771 = ~x_1134 & ~n_14769;
assign n_14772 = ~n_14770 & ~n_14771;
assign n_14773 =  x_1133 & ~n_14656;
assign n_14774 =  x_1133 &  n_14773;
assign n_14775 = ~x_1133 & ~n_14773;
assign n_14776 = ~n_14774 & ~n_14775;
assign n_14777 =  x_1132 & ~n_14656;
assign n_14778 =  x_1132 &  n_14777;
assign n_14779 = ~x_1132 & ~n_14777;
assign n_14780 = ~n_14778 & ~n_14779;
assign n_14781 =  x_1131 & ~n_14656;
assign n_14782 =  x_1131 &  n_14781;
assign n_14783 = ~x_1131 & ~n_14781;
assign n_14784 = ~n_14782 & ~n_14783;
assign n_14785 =  x_39 &  n_356;
assign n_14786 =  n_9689 &  n_14785;
assign n_14787 =  x_43 &  n_14786;
assign n_14788 = ~x_1610 &  n_12323;
assign n_14789 =  x_1610 &  n_12328;
assign n_14790 =  i_32 & ~n_12331;
assign n_14791 =  x_3064 &  n_12331;
assign n_14792 = ~n_14790 & ~n_14791;
assign n_14793 = ~n_12329 & ~n_14792;
assign n_14794 =  x_3032 &  n_12329;
assign n_14795 = ~n_14793 & ~n_14794;
assign n_14796 = ~n_14789 & ~n_14795;
assign n_14797 =  x_2906 &  n_14789;
assign n_14798 = ~n_14796 & ~n_14797;
assign n_14799 = ~n_14788 & ~n_14798;
assign n_14800 =  x_2842 &  n_14788;
assign n_14801 = ~n_14799 & ~n_14800;
assign n_14802 =  n_14787 & ~n_14801;
assign n_14803 =  x_1130 & ~n_14787;
assign n_14804 = ~n_14802 & ~n_14803;
assign n_14805 =  x_1130 & ~n_14804;
assign n_14806 = ~x_1130 &  n_14804;
assign n_14807 = ~n_14805 & ~n_14806;
assign n_14808 =  i_31 & ~n_12331;
assign n_14809 =  x_3063 &  n_12331;
assign n_14810 = ~n_14808 & ~n_14809;
assign n_14811 = ~n_12329 & ~n_14810;
assign n_14812 =  x_3031 &  n_12329;
assign n_14813 = ~n_14811 & ~n_14812;
assign n_14814 = ~n_14789 & ~n_14813;
assign n_14815 =  x_2905 &  n_14789;
assign n_14816 = ~n_14814 & ~n_14815;
assign n_14817 = ~n_14788 & ~n_14816;
assign n_14818 =  x_2841 &  n_14788;
assign n_14819 = ~n_14817 & ~n_14818;
assign n_14820 =  n_14787 & ~n_14819;
assign n_14821 =  x_1129 & ~n_14787;
assign n_14822 = ~n_14820 & ~n_14821;
assign n_14823 =  x_1129 & ~n_14822;
assign n_14824 = ~x_1129 &  n_14822;
assign n_14825 = ~n_14823 & ~n_14824;
assign n_14826 =  i_30 & ~n_12331;
assign n_14827 =  x_3062 &  n_12331;
assign n_14828 = ~n_14826 & ~n_14827;
assign n_14829 = ~n_12329 & ~n_14828;
assign n_14830 =  x_3030 &  n_12329;
assign n_14831 = ~n_14829 & ~n_14830;
assign n_14832 = ~n_14789 & ~n_14831;
assign n_14833 =  x_2904 &  n_14789;
assign n_14834 = ~n_14832 & ~n_14833;
assign n_14835 = ~n_14788 & ~n_14834;
assign n_14836 =  x_2840 &  n_14788;
assign n_14837 = ~n_14835 & ~n_14836;
assign n_14838 =  n_14787 & ~n_14837;
assign n_14839 =  x_1128 & ~n_14787;
assign n_14840 = ~n_14838 & ~n_14839;
assign n_14841 =  x_1128 & ~n_14840;
assign n_14842 = ~x_1128 &  n_14840;
assign n_14843 = ~n_14841 & ~n_14842;
assign n_14844 =  i_29 & ~n_12331;
assign n_14845 =  x_3061 &  n_12331;
assign n_14846 = ~n_14844 & ~n_14845;
assign n_14847 = ~n_12329 & ~n_14846;
assign n_14848 =  x_3029 &  n_12329;
assign n_14849 = ~n_14847 & ~n_14848;
assign n_14850 = ~n_14789 & ~n_14849;
assign n_14851 =  x_2903 &  n_14789;
assign n_14852 = ~n_14850 & ~n_14851;
assign n_14853 = ~n_14788 & ~n_14852;
assign n_14854 =  x_2839 &  n_14788;
assign n_14855 = ~n_14853 & ~n_14854;
assign n_14856 =  n_14787 & ~n_14855;
assign n_14857 =  x_1127 & ~n_14787;
assign n_14858 = ~n_14856 & ~n_14857;
assign n_14859 =  x_1127 & ~n_14858;
assign n_14860 = ~x_1127 &  n_14858;
assign n_14861 = ~n_14859 & ~n_14860;
assign n_14862 =  i_28 & ~n_12331;
assign n_14863 =  x_3060 &  n_12331;
assign n_14864 = ~n_14862 & ~n_14863;
assign n_14865 = ~n_12329 & ~n_14864;
assign n_14866 =  x_3028 &  n_12329;
assign n_14867 = ~n_14865 & ~n_14866;
assign n_14868 = ~n_14789 & ~n_14867;
assign n_14869 =  x_2902 &  n_14789;
assign n_14870 = ~n_14868 & ~n_14869;
assign n_14871 = ~n_14788 & ~n_14870;
assign n_14872 =  x_2838 &  n_14788;
assign n_14873 = ~n_14871 & ~n_14872;
assign n_14874 =  n_14787 & ~n_14873;
assign n_14875 =  x_1126 & ~n_14787;
assign n_14876 = ~n_14874 & ~n_14875;
assign n_14877 =  x_1126 & ~n_14876;
assign n_14878 = ~x_1126 &  n_14876;
assign n_14879 = ~n_14877 & ~n_14878;
assign n_14880 =  i_27 & ~n_12331;
assign n_14881 =  x_3059 &  n_12331;
assign n_14882 = ~n_14880 & ~n_14881;
assign n_14883 = ~n_12329 & ~n_14882;
assign n_14884 =  x_3027 &  n_12329;
assign n_14885 = ~n_14883 & ~n_14884;
assign n_14886 = ~n_14789 & ~n_14885;
assign n_14887 =  x_2901 &  n_14789;
assign n_14888 = ~n_14886 & ~n_14887;
assign n_14889 = ~n_14788 & ~n_14888;
assign n_14890 =  x_2837 &  n_14788;
assign n_14891 = ~n_14889 & ~n_14890;
assign n_14892 =  n_14787 & ~n_14891;
assign n_14893 =  x_1125 & ~n_14787;
assign n_14894 = ~n_14892 & ~n_14893;
assign n_14895 =  x_1125 & ~n_14894;
assign n_14896 = ~x_1125 &  n_14894;
assign n_14897 = ~n_14895 & ~n_14896;
assign n_14898 =  i_26 & ~n_12331;
assign n_14899 =  x_3058 &  n_12331;
assign n_14900 = ~n_14898 & ~n_14899;
assign n_14901 = ~n_12329 & ~n_14900;
assign n_14902 =  x_3026 &  n_12329;
assign n_14903 = ~n_14901 & ~n_14902;
assign n_14904 = ~n_14789 & ~n_14903;
assign n_14905 =  x_2900 &  n_14789;
assign n_14906 = ~n_14904 & ~n_14905;
assign n_14907 = ~n_14788 & ~n_14906;
assign n_14908 =  x_2836 &  n_14788;
assign n_14909 = ~n_14907 & ~n_14908;
assign n_14910 =  n_14787 & ~n_14909;
assign n_14911 =  x_1124 & ~n_14787;
assign n_14912 = ~n_14910 & ~n_14911;
assign n_14913 =  x_1124 & ~n_14912;
assign n_14914 = ~x_1124 &  n_14912;
assign n_14915 = ~n_14913 & ~n_14914;
assign n_14916 =  i_25 & ~n_12331;
assign n_14917 =  x_3057 &  n_12331;
assign n_14918 = ~n_14916 & ~n_14917;
assign n_14919 = ~n_12329 & ~n_14918;
assign n_14920 =  x_3025 &  n_12329;
assign n_14921 = ~n_14919 & ~n_14920;
assign n_14922 = ~n_14789 & ~n_14921;
assign n_14923 =  x_2899 &  n_14789;
assign n_14924 = ~n_14922 & ~n_14923;
assign n_14925 = ~n_14788 & ~n_14924;
assign n_14926 =  x_2835 &  n_14788;
assign n_14927 = ~n_14925 & ~n_14926;
assign n_14928 =  n_14787 & ~n_14927;
assign n_14929 =  x_1123 & ~n_14787;
assign n_14930 = ~n_14928 & ~n_14929;
assign n_14931 =  x_1123 & ~n_14930;
assign n_14932 = ~x_1123 &  n_14930;
assign n_14933 = ~n_14931 & ~n_14932;
assign n_14934 =  i_24 & ~n_12331;
assign n_14935 =  x_3056 &  n_12331;
assign n_14936 = ~n_14934 & ~n_14935;
assign n_14937 = ~n_12329 & ~n_14936;
assign n_14938 =  x_3024 &  n_12329;
assign n_14939 = ~n_14937 & ~n_14938;
assign n_14940 = ~n_14789 & ~n_14939;
assign n_14941 =  x_2898 &  n_14789;
assign n_14942 = ~n_14940 & ~n_14941;
assign n_14943 = ~n_14788 & ~n_14942;
assign n_14944 =  x_2834 &  n_14788;
assign n_14945 = ~n_14943 & ~n_14944;
assign n_14946 =  n_14787 & ~n_14945;
assign n_14947 =  x_1122 & ~n_14787;
assign n_14948 = ~n_14946 & ~n_14947;
assign n_14949 =  x_1122 & ~n_14948;
assign n_14950 = ~x_1122 &  n_14948;
assign n_14951 = ~n_14949 & ~n_14950;
assign n_14952 =  i_23 & ~n_12331;
assign n_14953 =  x_3055 &  n_12331;
assign n_14954 = ~n_14952 & ~n_14953;
assign n_14955 = ~n_12329 & ~n_14954;
assign n_14956 =  x_3023 &  n_12329;
assign n_14957 = ~n_14955 & ~n_14956;
assign n_14958 = ~n_14789 & ~n_14957;
assign n_14959 =  x_2897 &  n_14789;
assign n_14960 = ~n_14958 & ~n_14959;
assign n_14961 = ~n_14788 & ~n_14960;
assign n_14962 =  x_2833 &  n_14788;
assign n_14963 = ~n_14961 & ~n_14962;
assign n_14964 =  n_14787 & ~n_14963;
assign n_14965 =  x_1121 & ~n_14787;
assign n_14966 = ~n_14964 & ~n_14965;
assign n_14967 =  x_1121 & ~n_14966;
assign n_14968 = ~x_1121 &  n_14966;
assign n_14969 = ~n_14967 & ~n_14968;
assign n_14970 =  i_22 & ~n_12331;
assign n_14971 =  x_3054 &  n_12331;
assign n_14972 = ~n_14970 & ~n_14971;
assign n_14973 = ~n_12329 & ~n_14972;
assign n_14974 =  x_3022 &  n_12329;
assign n_14975 = ~n_14973 & ~n_14974;
assign n_14976 = ~n_14789 & ~n_14975;
assign n_14977 =  x_2896 &  n_14789;
assign n_14978 = ~n_14976 & ~n_14977;
assign n_14979 = ~n_14788 & ~n_14978;
assign n_14980 =  x_2832 &  n_14788;
assign n_14981 = ~n_14979 & ~n_14980;
assign n_14982 =  n_14787 & ~n_14981;
assign n_14983 =  x_1120 & ~n_14787;
assign n_14984 = ~n_14982 & ~n_14983;
assign n_14985 =  x_1120 & ~n_14984;
assign n_14986 = ~x_1120 &  n_14984;
assign n_14987 = ~n_14985 & ~n_14986;
assign n_14988 =  i_21 & ~n_12331;
assign n_14989 =  x_3053 &  n_12331;
assign n_14990 = ~n_14988 & ~n_14989;
assign n_14991 = ~n_12329 & ~n_14990;
assign n_14992 =  x_3021 &  n_12329;
assign n_14993 = ~n_14991 & ~n_14992;
assign n_14994 = ~n_14789 & ~n_14993;
assign n_14995 =  x_2895 &  n_14789;
assign n_14996 = ~n_14994 & ~n_14995;
assign n_14997 = ~n_14788 & ~n_14996;
assign n_14998 =  x_2831 &  n_14788;
assign n_14999 = ~n_14997 & ~n_14998;
assign n_15000 =  n_14787 & ~n_14999;
assign n_15001 =  x_1119 & ~n_14787;
assign n_15002 = ~n_15000 & ~n_15001;
assign n_15003 =  x_1119 & ~n_15002;
assign n_15004 = ~x_1119 &  n_15002;
assign n_15005 = ~n_15003 & ~n_15004;
assign n_15006 =  i_20 & ~n_12331;
assign n_15007 =  x_3052 &  n_12331;
assign n_15008 = ~n_15006 & ~n_15007;
assign n_15009 = ~n_12329 & ~n_15008;
assign n_15010 =  x_3020 &  n_12329;
assign n_15011 = ~n_15009 & ~n_15010;
assign n_15012 = ~n_14789 & ~n_15011;
assign n_15013 =  x_2894 &  n_14789;
assign n_15014 = ~n_15012 & ~n_15013;
assign n_15015 = ~n_14788 & ~n_15014;
assign n_15016 =  x_2830 &  n_14788;
assign n_15017 = ~n_15015 & ~n_15016;
assign n_15018 =  n_14787 & ~n_15017;
assign n_15019 =  x_1118 & ~n_14787;
assign n_15020 = ~n_15018 & ~n_15019;
assign n_15021 =  x_1118 & ~n_15020;
assign n_15022 = ~x_1118 &  n_15020;
assign n_15023 = ~n_15021 & ~n_15022;
assign n_15024 =  i_19 & ~n_12331;
assign n_15025 =  x_3051 &  n_12331;
assign n_15026 = ~n_15024 & ~n_15025;
assign n_15027 = ~n_12329 & ~n_15026;
assign n_15028 =  x_3019 &  n_12329;
assign n_15029 = ~n_15027 & ~n_15028;
assign n_15030 = ~n_14789 & ~n_15029;
assign n_15031 =  x_2893 &  n_14789;
assign n_15032 = ~n_15030 & ~n_15031;
assign n_15033 = ~n_14788 & ~n_15032;
assign n_15034 =  x_2829 &  n_14788;
assign n_15035 = ~n_15033 & ~n_15034;
assign n_15036 =  n_14787 & ~n_15035;
assign n_15037 =  x_1117 & ~n_14787;
assign n_15038 = ~n_15036 & ~n_15037;
assign n_15039 =  x_1117 & ~n_15038;
assign n_15040 = ~x_1117 &  n_15038;
assign n_15041 = ~n_15039 & ~n_15040;
assign n_15042 =  i_18 & ~n_12331;
assign n_15043 =  x_3050 &  n_12331;
assign n_15044 = ~n_15042 & ~n_15043;
assign n_15045 = ~n_12329 & ~n_15044;
assign n_15046 =  x_3018 &  n_12329;
assign n_15047 = ~n_15045 & ~n_15046;
assign n_15048 = ~n_14789 & ~n_15047;
assign n_15049 =  x_2892 &  n_14789;
assign n_15050 = ~n_15048 & ~n_15049;
assign n_15051 = ~n_14788 & ~n_15050;
assign n_15052 =  x_2828 &  n_14788;
assign n_15053 = ~n_15051 & ~n_15052;
assign n_15054 =  n_14787 & ~n_15053;
assign n_15055 =  x_1116 & ~n_14787;
assign n_15056 = ~n_15054 & ~n_15055;
assign n_15057 =  x_1116 & ~n_15056;
assign n_15058 = ~x_1116 &  n_15056;
assign n_15059 = ~n_15057 & ~n_15058;
assign n_15060 =  i_17 & ~n_12331;
assign n_15061 =  x_3049 &  n_12331;
assign n_15062 = ~n_15060 & ~n_15061;
assign n_15063 = ~n_12329 & ~n_15062;
assign n_15064 =  x_3017 &  n_12329;
assign n_15065 = ~n_15063 & ~n_15064;
assign n_15066 = ~n_14789 & ~n_15065;
assign n_15067 =  x_2891 &  n_14789;
assign n_15068 = ~n_15066 & ~n_15067;
assign n_15069 = ~n_14788 & ~n_15068;
assign n_15070 =  x_2827 &  n_14788;
assign n_15071 = ~n_15069 & ~n_15070;
assign n_15072 =  n_14787 & ~n_15071;
assign n_15073 =  x_1115 & ~n_14787;
assign n_15074 = ~n_15072 & ~n_15073;
assign n_15075 =  x_1115 & ~n_15074;
assign n_15076 = ~x_1115 &  n_15074;
assign n_15077 = ~n_15075 & ~n_15076;
assign n_15078 =  i_16 & ~n_12331;
assign n_15079 =  x_3048 &  n_12331;
assign n_15080 = ~n_15078 & ~n_15079;
assign n_15081 = ~n_12329 & ~n_15080;
assign n_15082 =  x_3016 &  n_12329;
assign n_15083 = ~n_15081 & ~n_15082;
assign n_15084 = ~n_14789 & ~n_15083;
assign n_15085 =  x_2890 &  n_14789;
assign n_15086 = ~n_15084 & ~n_15085;
assign n_15087 = ~n_14788 & ~n_15086;
assign n_15088 =  x_2826 &  n_14788;
assign n_15089 = ~n_15087 & ~n_15088;
assign n_15090 =  n_14787 & ~n_15089;
assign n_15091 =  x_1114 & ~n_14787;
assign n_15092 = ~n_15090 & ~n_15091;
assign n_15093 =  x_1114 & ~n_15092;
assign n_15094 = ~x_1114 &  n_15092;
assign n_15095 = ~n_15093 & ~n_15094;
assign n_15096 =  i_15 & ~n_12331;
assign n_15097 =  x_3047 &  n_12331;
assign n_15098 = ~n_15096 & ~n_15097;
assign n_15099 = ~n_12329 & ~n_15098;
assign n_15100 =  x_3015 &  n_12329;
assign n_15101 = ~n_15099 & ~n_15100;
assign n_15102 = ~n_14789 & ~n_15101;
assign n_15103 =  x_2889 &  n_14789;
assign n_15104 = ~n_15102 & ~n_15103;
assign n_15105 = ~n_14788 & ~n_15104;
assign n_15106 =  x_2825 &  n_14788;
assign n_15107 = ~n_15105 & ~n_15106;
assign n_15108 =  n_14787 & ~n_15107;
assign n_15109 =  x_1113 & ~n_14787;
assign n_15110 = ~n_15108 & ~n_15109;
assign n_15111 =  x_1113 & ~n_15110;
assign n_15112 = ~x_1113 &  n_15110;
assign n_15113 = ~n_15111 & ~n_15112;
assign n_15114 =  i_14 & ~n_12331;
assign n_15115 =  x_3046 &  n_12331;
assign n_15116 = ~n_15114 & ~n_15115;
assign n_15117 = ~n_12329 & ~n_15116;
assign n_15118 =  x_3014 &  n_12329;
assign n_15119 = ~n_15117 & ~n_15118;
assign n_15120 = ~n_14789 & ~n_15119;
assign n_15121 =  x_2888 &  n_14789;
assign n_15122 = ~n_15120 & ~n_15121;
assign n_15123 = ~n_14788 & ~n_15122;
assign n_15124 =  x_2824 &  n_14788;
assign n_15125 = ~n_15123 & ~n_15124;
assign n_15126 =  n_14787 & ~n_15125;
assign n_15127 =  x_1112 & ~n_14787;
assign n_15128 = ~n_15126 & ~n_15127;
assign n_15129 =  x_1112 & ~n_15128;
assign n_15130 = ~x_1112 &  n_15128;
assign n_15131 = ~n_15129 & ~n_15130;
assign n_15132 =  i_13 & ~n_12331;
assign n_15133 =  x_3045 &  n_12331;
assign n_15134 = ~n_15132 & ~n_15133;
assign n_15135 = ~n_12329 & ~n_15134;
assign n_15136 =  x_3013 &  n_12329;
assign n_15137 = ~n_15135 & ~n_15136;
assign n_15138 = ~n_14789 & ~n_15137;
assign n_15139 =  x_2887 &  n_14789;
assign n_15140 = ~n_15138 & ~n_15139;
assign n_15141 = ~n_14788 & ~n_15140;
assign n_15142 =  x_2823 &  n_14788;
assign n_15143 = ~n_15141 & ~n_15142;
assign n_15144 =  n_14787 & ~n_15143;
assign n_15145 =  x_1111 & ~n_14787;
assign n_15146 = ~n_15144 & ~n_15145;
assign n_15147 =  x_1111 & ~n_15146;
assign n_15148 = ~x_1111 &  n_15146;
assign n_15149 = ~n_15147 & ~n_15148;
assign n_15150 =  i_12 & ~n_12331;
assign n_15151 =  x_3044 &  n_12331;
assign n_15152 = ~n_15150 & ~n_15151;
assign n_15153 = ~n_12329 & ~n_15152;
assign n_15154 =  x_3012 &  n_12329;
assign n_15155 = ~n_15153 & ~n_15154;
assign n_15156 = ~n_14789 & ~n_15155;
assign n_15157 =  x_2886 &  n_14789;
assign n_15158 = ~n_15156 & ~n_15157;
assign n_15159 = ~n_14788 & ~n_15158;
assign n_15160 =  x_2822 &  n_14788;
assign n_15161 = ~n_15159 & ~n_15160;
assign n_15162 =  n_14787 & ~n_15161;
assign n_15163 =  x_1110 & ~n_14787;
assign n_15164 = ~n_15162 & ~n_15163;
assign n_15165 =  x_1110 & ~n_15164;
assign n_15166 = ~x_1110 &  n_15164;
assign n_15167 = ~n_15165 & ~n_15166;
assign n_15168 =  i_11 & ~n_12331;
assign n_15169 =  x_3043 &  n_12331;
assign n_15170 = ~n_15168 & ~n_15169;
assign n_15171 = ~n_12329 & ~n_15170;
assign n_15172 =  x_3011 &  n_12329;
assign n_15173 = ~n_15171 & ~n_15172;
assign n_15174 = ~n_14789 & ~n_15173;
assign n_15175 =  x_2885 &  n_14789;
assign n_15176 = ~n_15174 & ~n_15175;
assign n_15177 = ~n_14788 & ~n_15176;
assign n_15178 =  x_2821 &  n_14788;
assign n_15179 = ~n_15177 & ~n_15178;
assign n_15180 =  n_14787 & ~n_15179;
assign n_15181 =  x_1109 & ~n_14787;
assign n_15182 = ~n_15180 & ~n_15181;
assign n_15183 =  x_1109 & ~n_15182;
assign n_15184 = ~x_1109 &  n_15182;
assign n_15185 = ~n_15183 & ~n_15184;
assign n_15186 =  i_10 & ~n_12331;
assign n_15187 =  x_3042 &  n_12331;
assign n_15188 = ~n_15186 & ~n_15187;
assign n_15189 = ~n_12329 & ~n_15188;
assign n_15190 =  x_3010 &  n_12329;
assign n_15191 = ~n_15189 & ~n_15190;
assign n_15192 = ~n_14789 & ~n_15191;
assign n_15193 =  x_2884 &  n_14789;
assign n_15194 = ~n_15192 & ~n_15193;
assign n_15195 = ~n_14788 & ~n_15194;
assign n_15196 =  x_2820 &  n_14788;
assign n_15197 = ~n_15195 & ~n_15196;
assign n_15198 =  n_14787 & ~n_15197;
assign n_15199 =  x_1108 & ~n_14787;
assign n_15200 = ~n_15198 & ~n_15199;
assign n_15201 =  x_1108 & ~n_15200;
assign n_15202 = ~x_1108 &  n_15200;
assign n_15203 = ~n_15201 & ~n_15202;
assign n_15204 =  i_9 & ~n_12331;
assign n_15205 =  x_3041 &  n_12331;
assign n_15206 = ~n_15204 & ~n_15205;
assign n_15207 = ~n_12329 & ~n_15206;
assign n_15208 =  x_3009 &  n_12329;
assign n_15209 = ~n_15207 & ~n_15208;
assign n_15210 = ~n_14789 & ~n_15209;
assign n_15211 =  x_2883 &  n_14789;
assign n_15212 = ~n_15210 & ~n_15211;
assign n_15213 = ~n_14788 & ~n_15212;
assign n_15214 =  x_2819 &  n_14788;
assign n_15215 = ~n_15213 & ~n_15214;
assign n_15216 =  n_14787 & ~n_15215;
assign n_15217 =  x_1107 & ~n_14787;
assign n_15218 = ~n_15216 & ~n_15217;
assign n_15219 =  x_1107 & ~n_15218;
assign n_15220 = ~x_1107 &  n_15218;
assign n_15221 = ~n_15219 & ~n_15220;
assign n_15222 =  i_8 & ~n_12331;
assign n_15223 =  x_3040 &  n_12331;
assign n_15224 = ~n_15222 & ~n_15223;
assign n_15225 = ~n_12329 & ~n_15224;
assign n_15226 =  x_3008 &  n_12329;
assign n_15227 = ~n_15225 & ~n_15226;
assign n_15228 = ~n_14789 & ~n_15227;
assign n_15229 =  x_2882 &  n_14789;
assign n_15230 = ~n_15228 & ~n_15229;
assign n_15231 = ~n_14788 & ~n_15230;
assign n_15232 =  x_2818 &  n_14788;
assign n_15233 = ~n_15231 & ~n_15232;
assign n_15234 =  n_14787 & ~n_15233;
assign n_15235 =  x_1106 & ~n_14787;
assign n_15236 = ~n_15234 & ~n_15235;
assign n_15237 =  x_1106 & ~n_15236;
assign n_15238 = ~x_1106 &  n_15236;
assign n_15239 = ~n_15237 & ~n_15238;
assign n_15240 =  i_7 & ~n_12331;
assign n_15241 =  x_3039 &  n_12331;
assign n_15242 = ~n_15240 & ~n_15241;
assign n_15243 = ~n_12329 & ~n_15242;
assign n_15244 =  x_3007 &  n_12329;
assign n_15245 = ~n_15243 & ~n_15244;
assign n_15246 = ~n_14789 & ~n_15245;
assign n_15247 =  x_2881 &  n_14789;
assign n_15248 = ~n_15246 & ~n_15247;
assign n_15249 = ~n_14788 & ~n_15248;
assign n_15250 =  x_2817 &  n_14788;
assign n_15251 = ~n_15249 & ~n_15250;
assign n_15252 =  n_14787 & ~n_15251;
assign n_15253 =  x_1105 & ~n_14787;
assign n_15254 = ~n_15252 & ~n_15253;
assign n_15255 =  x_1105 & ~n_15254;
assign n_15256 = ~x_1105 &  n_15254;
assign n_15257 = ~n_15255 & ~n_15256;
assign n_15258 =  i_6 & ~n_12331;
assign n_15259 =  x_3038 &  n_12331;
assign n_15260 = ~n_15258 & ~n_15259;
assign n_15261 = ~n_12329 & ~n_15260;
assign n_15262 =  x_3006 &  n_12329;
assign n_15263 = ~n_15261 & ~n_15262;
assign n_15264 = ~n_14789 & ~n_15263;
assign n_15265 =  x_2880 &  n_14789;
assign n_15266 = ~n_15264 & ~n_15265;
assign n_15267 = ~n_14788 & ~n_15266;
assign n_15268 =  x_2816 &  n_14788;
assign n_15269 = ~n_15267 & ~n_15268;
assign n_15270 =  n_14787 & ~n_15269;
assign n_15271 =  x_1104 & ~n_14787;
assign n_15272 = ~n_15270 & ~n_15271;
assign n_15273 =  x_1104 & ~n_15272;
assign n_15274 = ~x_1104 &  n_15272;
assign n_15275 = ~n_15273 & ~n_15274;
assign n_15276 =  i_5 & ~n_12331;
assign n_15277 =  x_3037 &  n_12331;
assign n_15278 = ~n_15276 & ~n_15277;
assign n_15279 = ~n_12329 & ~n_15278;
assign n_15280 =  x_3005 &  n_12329;
assign n_15281 = ~n_15279 & ~n_15280;
assign n_15282 = ~n_14789 & ~n_15281;
assign n_15283 =  x_2879 &  n_14789;
assign n_15284 = ~n_15282 & ~n_15283;
assign n_15285 = ~n_14788 & ~n_15284;
assign n_15286 =  x_2815 &  n_14788;
assign n_15287 = ~n_15285 & ~n_15286;
assign n_15288 =  n_14787 & ~n_15287;
assign n_15289 =  x_1103 & ~n_14787;
assign n_15290 = ~n_15288 & ~n_15289;
assign n_15291 =  x_1103 & ~n_15290;
assign n_15292 = ~x_1103 &  n_15290;
assign n_15293 = ~n_15291 & ~n_15292;
assign n_15294 =  i_4 & ~n_12331;
assign n_15295 =  x_3036 &  n_12331;
assign n_15296 = ~n_15294 & ~n_15295;
assign n_15297 = ~n_12329 & ~n_15296;
assign n_15298 =  x_3004 &  n_12329;
assign n_15299 = ~n_15297 & ~n_15298;
assign n_15300 = ~n_14789 & ~n_15299;
assign n_15301 =  x_2878 &  n_14789;
assign n_15302 = ~n_15300 & ~n_15301;
assign n_15303 = ~n_14788 & ~n_15302;
assign n_15304 =  x_2814 &  n_14788;
assign n_15305 = ~n_15303 & ~n_15304;
assign n_15306 =  n_14787 & ~n_15305;
assign n_15307 =  x_1102 & ~n_14787;
assign n_15308 = ~n_15306 & ~n_15307;
assign n_15309 =  x_1102 & ~n_15308;
assign n_15310 = ~x_1102 &  n_15308;
assign n_15311 = ~n_15309 & ~n_15310;
assign n_15312 =  i_3 & ~n_12331;
assign n_15313 =  x_3035 &  n_12331;
assign n_15314 = ~n_15312 & ~n_15313;
assign n_15315 = ~n_12329 & ~n_15314;
assign n_15316 =  x_3003 &  n_12329;
assign n_15317 = ~n_15315 & ~n_15316;
assign n_15318 = ~n_14789 & ~n_15317;
assign n_15319 =  x_2877 &  n_14789;
assign n_15320 = ~n_15318 & ~n_15319;
assign n_15321 = ~n_14788 & ~n_15320;
assign n_15322 =  x_2813 &  n_14788;
assign n_15323 = ~n_15321 & ~n_15322;
assign n_15324 =  n_14787 & ~n_15323;
assign n_15325 =  x_1101 & ~n_14787;
assign n_15326 = ~n_15324 & ~n_15325;
assign n_15327 =  x_1101 & ~n_15326;
assign n_15328 = ~x_1101 &  n_15326;
assign n_15329 = ~n_15327 & ~n_15328;
assign n_15330 =  i_2 & ~n_12331;
assign n_15331 =  x_3034 &  n_12331;
assign n_15332 = ~n_15330 & ~n_15331;
assign n_15333 = ~n_12329 & ~n_15332;
assign n_15334 =  x_3002 &  n_12329;
assign n_15335 = ~n_15333 & ~n_15334;
assign n_15336 = ~n_14789 & ~n_15335;
assign n_15337 =  x_2876 &  n_14789;
assign n_15338 = ~n_15336 & ~n_15337;
assign n_15339 = ~n_14788 & ~n_15338;
assign n_15340 =  x_2812 &  n_14788;
assign n_15341 = ~n_15339 & ~n_15340;
assign n_15342 =  n_14787 & ~n_15341;
assign n_15343 =  x_1100 & ~n_14787;
assign n_15344 = ~n_15342 & ~n_15343;
assign n_15345 =  x_1100 & ~n_15344;
assign n_15346 = ~x_1100 &  n_15344;
assign n_15347 = ~n_15345 & ~n_15346;
assign n_15348 =  i_1 & ~n_12331;
assign n_15349 =  x_3033 &  n_12331;
assign n_15350 = ~n_15348 & ~n_15349;
assign n_15351 = ~n_12329 & ~n_15350;
assign n_15352 =  x_3001 &  n_12329;
assign n_15353 = ~n_15351 & ~n_15352;
assign n_15354 = ~n_14789 & ~n_15353;
assign n_15355 =  x_2875 &  n_14789;
assign n_15356 = ~n_15354 & ~n_15355;
assign n_15357 = ~n_14788 & ~n_15356;
assign n_15358 =  x_2811 &  n_14788;
assign n_15359 = ~n_15357 & ~n_15358;
assign n_15360 =  n_14787 & ~n_15359;
assign n_15361 =  x_1099 & ~n_14787;
assign n_15362 = ~n_15360 & ~n_15361;
assign n_15363 =  x_1099 & ~n_15362;
assign n_15364 = ~x_1099 &  n_15362;
assign n_15365 = ~n_15363 & ~n_15364;
assign n_15366 =  x_40 &  n_5645;
assign n_15367 =  n_15366 &  n_3619;
assign n_15368 =  x_1098 & ~n_15367;
assign n_15369 = ~x_3064 &  n_13143;
assign n_15370 = ~i_32 & ~n_13143;
assign n_15371 = ~n_13140 & ~n_15370;
assign n_15372 = ~n_15369 &  n_15371;
assign n_15373 =  x_4775 &  n_13140;
assign n_15374 =  x_2906 &  n_15373;
assign n_15375 = ~x_4775 &  n_13135;
assign n_15376 =  x_3032 &  n_13141;
assign n_15377 = ~n_15375 & ~n_15376;
assign n_15378 = ~n_15374 &  n_15377;
assign n_15379 = ~n_15372 &  n_15378;
assign n_15380 = ~x_2842 &  n_15375;
assign n_15381 =  n_15367 & ~n_15380;
assign n_15382 = ~n_15379 &  n_15381;
assign n_15383 = ~n_15368 & ~n_15382;
assign n_15384 =  x_1098 & ~n_15383;
assign n_15385 = ~x_1098 &  n_15383;
assign n_15386 = ~n_15384 & ~n_15385;
assign n_15387 =  x_1097 & ~n_15367;
assign n_15388 = ~x_3063 &  n_13143;
assign n_15389 = ~i_31 & ~n_13143;
assign n_15390 = ~n_13140 & ~n_15389;
assign n_15391 = ~n_15388 &  n_15390;
assign n_15392 =  x_2905 &  n_15373;
assign n_15393 =  x_3031 &  n_13141;
assign n_15394 = ~n_15375 & ~n_15393;
assign n_15395 = ~n_15392 &  n_15394;
assign n_15396 = ~n_15391 &  n_15395;
assign n_15397 = ~x_2841 &  n_15375;
assign n_15398 =  n_15367 & ~n_15397;
assign n_15399 = ~n_15396 &  n_15398;
assign n_15400 = ~n_15387 & ~n_15399;
assign n_15401 =  x_1097 & ~n_15400;
assign n_15402 = ~x_1097 &  n_15400;
assign n_15403 = ~n_15401 & ~n_15402;
assign n_15404 =  x_1096 & ~n_15367;
assign n_15405 = ~x_3062 &  n_13143;
assign n_15406 = ~i_30 & ~n_13143;
assign n_15407 = ~n_13140 & ~n_15406;
assign n_15408 = ~n_15405 &  n_15407;
assign n_15409 =  x_2904 &  n_15373;
assign n_15410 =  x_3030 &  n_13141;
assign n_15411 = ~n_15375 & ~n_15410;
assign n_15412 = ~n_15409 &  n_15411;
assign n_15413 = ~n_15408 &  n_15412;
assign n_15414 = ~x_2840 &  n_15375;
assign n_15415 =  n_15367 & ~n_15414;
assign n_15416 = ~n_15413 &  n_15415;
assign n_15417 = ~n_15404 & ~n_15416;
assign n_15418 =  x_1096 & ~n_15417;
assign n_15419 = ~x_1096 &  n_15417;
assign n_15420 = ~n_15418 & ~n_15419;
assign n_15421 =  x_1095 & ~n_15367;
assign n_15422 = ~x_3061 &  n_13143;
assign n_15423 = ~i_29 & ~n_13143;
assign n_15424 = ~n_13140 & ~n_15423;
assign n_15425 = ~n_15422 &  n_15424;
assign n_15426 =  x_2903 &  n_15373;
assign n_15427 =  x_3029 &  n_13141;
assign n_15428 = ~n_15375 & ~n_15427;
assign n_15429 = ~n_15426 &  n_15428;
assign n_15430 = ~n_15425 &  n_15429;
assign n_15431 = ~x_2839 &  n_15375;
assign n_15432 =  n_15367 & ~n_15431;
assign n_15433 = ~n_15430 &  n_15432;
assign n_15434 = ~n_15421 & ~n_15433;
assign n_15435 =  x_1095 & ~n_15434;
assign n_15436 = ~x_1095 &  n_15434;
assign n_15437 = ~n_15435 & ~n_15436;
assign n_15438 =  x_1094 & ~n_15367;
assign n_15439 = ~x_3060 &  n_13143;
assign n_15440 = ~i_28 & ~n_13143;
assign n_15441 = ~n_13140 & ~n_15440;
assign n_15442 = ~n_15439 &  n_15441;
assign n_15443 =  x_2902 &  n_15373;
assign n_15444 =  x_3028 &  n_13141;
assign n_15445 = ~n_15375 & ~n_15444;
assign n_15446 = ~n_15443 &  n_15445;
assign n_15447 = ~n_15442 &  n_15446;
assign n_15448 = ~x_2838 &  n_15375;
assign n_15449 =  n_15367 & ~n_15448;
assign n_15450 = ~n_15447 &  n_15449;
assign n_15451 = ~n_15438 & ~n_15450;
assign n_15452 =  x_1094 & ~n_15451;
assign n_15453 = ~x_1094 &  n_15451;
assign n_15454 = ~n_15452 & ~n_15453;
assign n_15455 =  x_1093 & ~n_15367;
assign n_15456 = ~x_3059 &  n_13143;
assign n_15457 = ~i_27 & ~n_13143;
assign n_15458 = ~n_13140 & ~n_15457;
assign n_15459 = ~n_15456 &  n_15458;
assign n_15460 =  x_2901 &  n_15373;
assign n_15461 =  x_3027 &  n_13141;
assign n_15462 = ~n_15375 & ~n_15461;
assign n_15463 = ~n_15460 &  n_15462;
assign n_15464 = ~n_15459 &  n_15463;
assign n_15465 = ~x_2837 &  n_15375;
assign n_15466 =  n_15367 & ~n_15465;
assign n_15467 = ~n_15464 &  n_15466;
assign n_15468 = ~n_15455 & ~n_15467;
assign n_15469 =  x_1093 & ~n_15468;
assign n_15470 = ~x_1093 &  n_15468;
assign n_15471 = ~n_15469 & ~n_15470;
assign n_15472 =  x_1092 & ~n_15367;
assign n_15473 = ~x_3058 &  n_13143;
assign n_15474 = ~i_26 & ~n_13143;
assign n_15475 = ~n_13140 & ~n_15474;
assign n_15476 = ~n_15473 &  n_15475;
assign n_15477 =  x_2900 &  n_15373;
assign n_15478 =  x_3026 &  n_13141;
assign n_15479 = ~n_15375 & ~n_15478;
assign n_15480 = ~n_15477 &  n_15479;
assign n_15481 = ~n_15476 &  n_15480;
assign n_15482 = ~x_2836 &  n_15375;
assign n_15483 =  n_15367 & ~n_15482;
assign n_15484 = ~n_15481 &  n_15483;
assign n_15485 = ~n_15472 & ~n_15484;
assign n_15486 =  x_1092 & ~n_15485;
assign n_15487 = ~x_1092 &  n_15485;
assign n_15488 = ~n_15486 & ~n_15487;
assign n_15489 =  x_1091 & ~n_15367;
assign n_15490 = ~x_3057 &  n_13143;
assign n_15491 = ~i_25 & ~n_13143;
assign n_15492 = ~n_13140 & ~n_15491;
assign n_15493 = ~n_15490 &  n_15492;
assign n_15494 =  x_2899 &  n_15373;
assign n_15495 =  x_3025 &  n_13141;
assign n_15496 = ~n_15375 & ~n_15495;
assign n_15497 = ~n_15494 &  n_15496;
assign n_15498 = ~n_15493 &  n_15497;
assign n_15499 = ~x_2835 &  n_15375;
assign n_15500 =  n_15367 & ~n_15499;
assign n_15501 = ~n_15498 &  n_15500;
assign n_15502 = ~n_15489 & ~n_15501;
assign n_15503 =  x_1091 & ~n_15502;
assign n_15504 = ~x_1091 &  n_15502;
assign n_15505 = ~n_15503 & ~n_15504;
assign n_15506 =  x_1090 & ~n_15367;
assign n_15507 = ~x_3056 &  n_13143;
assign n_15508 = ~i_24 & ~n_13143;
assign n_15509 = ~n_13140 & ~n_15508;
assign n_15510 = ~n_15507 &  n_15509;
assign n_15511 =  x_2898 &  n_15373;
assign n_15512 =  x_3024 &  n_13141;
assign n_15513 = ~n_15375 & ~n_15512;
assign n_15514 = ~n_15511 &  n_15513;
assign n_15515 = ~n_15510 &  n_15514;
assign n_15516 = ~x_2834 &  n_15375;
assign n_15517 =  n_15367 & ~n_15516;
assign n_15518 = ~n_15515 &  n_15517;
assign n_15519 = ~n_15506 & ~n_15518;
assign n_15520 =  x_1090 & ~n_15519;
assign n_15521 = ~x_1090 &  n_15519;
assign n_15522 = ~n_15520 & ~n_15521;
assign n_15523 =  x_1089 & ~n_15367;
assign n_15524 = ~x_3055 &  n_13143;
assign n_15525 = ~i_23 & ~n_13143;
assign n_15526 = ~n_13140 & ~n_15525;
assign n_15527 = ~n_15524 &  n_15526;
assign n_15528 =  x_2897 &  n_15373;
assign n_15529 =  x_3023 &  n_13141;
assign n_15530 = ~n_15375 & ~n_15529;
assign n_15531 = ~n_15528 &  n_15530;
assign n_15532 = ~n_15527 &  n_15531;
assign n_15533 = ~x_2833 &  n_15375;
assign n_15534 =  n_15367 & ~n_15533;
assign n_15535 = ~n_15532 &  n_15534;
assign n_15536 = ~n_15523 & ~n_15535;
assign n_15537 =  x_1089 & ~n_15536;
assign n_15538 = ~x_1089 &  n_15536;
assign n_15539 = ~n_15537 & ~n_15538;
assign n_15540 =  x_1088 & ~n_15367;
assign n_15541 = ~x_3054 &  n_13143;
assign n_15542 = ~i_22 & ~n_13143;
assign n_15543 = ~n_13140 & ~n_15542;
assign n_15544 = ~n_15541 &  n_15543;
assign n_15545 =  x_2896 &  n_15373;
assign n_15546 =  x_3022 &  n_13141;
assign n_15547 = ~n_15375 & ~n_15546;
assign n_15548 = ~n_15545 &  n_15547;
assign n_15549 = ~n_15544 &  n_15548;
assign n_15550 = ~x_2832 &  n_15375;
assign n_15551 =  n_15367 & ~n_15550;
assign n_15552 = ~n_15549 &  n_15551;
assign n_15553 = ~n_15540 & ~n_15552;
assign n_15554 =  x_1088 & ~n_15553;
assign n_15555 = ~x_1088 &  n_15553;
assign n_15556 = ~n_15554 & ~n_15555;
assign n_15557 =  x_1087 & ~n_15367;
assign n_15558 = ~x_3053 &  n_13143;
assign n_15559 = ~i_21 & ~n_13143;
assign n_15560 = ~n_13140 & ~n_15559;
assign n_15561 = ~n_15558 &  n_15560;
assign n_15562 =  x_2895 &  n_15373;
assign n_15563 =  x_3021 &  n_13141;
assign n_15564 = ~n_15375 & ~n_15563;
assign n_15565 = ~n_15562 &  n_15564;
assign n_15566 = ~n_15561 &  n_15565;
assign n_15567 = ~x_2831 &  n_15375;
assign n_15568 =  n_15367 & ~n_15567;
assign n_15569 = ~n_15566 &  n_15568;
assign n_15570 = ~n_15557 & ~n_15569;
assign n_15571 =  x_1087 & ~n_15570;
assign n_15572 = ~x_1087 &  n_15570;
assign n_15573 = ~n_15571 & ~n_15572;
assign n_15574 =  x_1086 & ~n_15367;
assign n_15575 = ~x_3052 &  n_13143;
assign n_15576 = ~i_20 & ~n_13143;
assign n_15577 = ~n_13140 & ~n_15576;
assign n_15578 = ~n_15575 &  n_15577;
assign n_15579 =  x_2894 &  n_15373;
assign n_15580 =  x_3020 &  n_13141;
assign n_15581 = ~n_15375 & ~n_15580;
assign n_15582 = ~n_15579 &  n_15581;
assign n_15583 = ~n_15578 &  n_15582;
assign n_15584 = ~x_2830 &  n_15375;
assign n_15585 =  n_15367 & ~n_15584;
assign n_15586 = ~n_15583 &  n_15585;
assign n_15587 = ~n_15574 & ~n_15586;
assign n_15588 =  x_1086 & ~n_15587;
assign n_15589 = ~x_1086 &  n_15587;
assign n_15590 = ~n_15588 & ~n_15589;
assign n_15591 =  x_1085 & ~n_15367;
assign n_15592 = ~x_3051 &  n_13143;
assign n_15593 = ~i_19 & ~n_13143;
assign n_15594 = ~n_13140 & ~n_15593;
assign n_15595 = ~n_15592 &  n_15594;
assign n_15596 =  x_2893 &  n_15373;
assign n_15597 =  x_3019 &  n_13141;
assign n_15598 = ~n_15375 & ~n_15597;
assign n_15599 = ~n_15596 &  n_15598;
assign n_15600 = ~n_15595 &  n_15599;
assign n_15601 = ~x_2829 &  n_15375;
assign n_15602 =  n_15367 & ~n_15601;
assign n_15603 = ~n_15600 &  n_15602;
assign n_15604 = ~n_15591 & ~n_15603;
assign n_15605 =  x_1085 & ~n_15604;
assign n_15606 = ~x_1085 &  n_15604;
assign n_15607 = ~n_15605 & ~n_15606;
assign n_15608 =  x_1084 & ~n_15367;
assign n_15609 = ~x_3050 &  n_13143;
assign n_15610 = ~i_18 & ~n_13143;
assign n_15611 = ~n_13140 & ~n_15610;
assign n_15612 = ~n_15609 &  n_15611;
assign n_15613 =  x_2892 &  n_15373;
assign n_15614 =  x_3018 &  n_13141;
assign n_15615 = ~n_15375 & ~n_15614;
assign n_15616 = ~n_15613 &  n_15615;
assign n_15617 = ~n_15612 &  n_15616;
assign n_15618 = ~x_2828 &  n_15375;
assign n_15619 =  n_15367 & ~n_15618;
assign n_15620 = ~n_15617 &  n_15619;
assign n_15621 = ~n_15608 & ~n_15620;
assign n_15622 =  x_1084 & ~n_15621;
assign n_15623 = ~x_1084 &  n_15621;
assign n_15624 = ~n_15622 & ~n_15623;
assign n_15625 =  x_1083 & ~n_15367;
assign n_15626 = ~x_3049 &  n_13143;
assign n_15627 = ~i_17 & ~n_13143;
assign n_15628 = ~n_13140 & ~n_15627;
assign n_15629 = ~n_15626 &  n_15628;
assign n_15630 =  x_2891 &  n_15373;
assign n_15631 =  x_3017 &  n_13141;
assign n_15632 = ~n_15375 & ~n_15631;
assign n_15633 = ~n_15630 &  n_15632;
assign n_15634 = ~n_15629 &  n_15633;
assign n_15635 = ~x_2827 &  n_15375;
assign n_15636 =  n_15367 & ~n_15635;
assign n_15637 = ~n_15634 &  n_15636;
assign n_15638 = ~n_15625 & ~n_15637;
assign n_15639 =  x_1083 & ~n_15638;
assign n_15640 = ~x_1083 &  n_15638;
assign n_15641 = ~n_15639 & ~n_15640;
assign n_15642 =  x_1082 & ~n_15367;
assign n_15643 = ~x_3048 &  n_13143;
assign n_15644 = ~i_16 & ~n_13143;
assign n_15645 = ~n_13140 & ~n_15644;
assign n_15646 = ~n_15643 &  n_15645;
assign n_15647 =  x_2890 &  n_15373;
assign n_15648 =  x_3016 &  n_13141;
assign n_15649 = ~n_15375 & ~n_15648;
assign n_15650 = ~n_15647 &  n_15649;
assign n_15651 = ~n_15646 &  n_15650;
assign n_15652 = ~x_2826 &  n_15375;
assign n_15653 =  n_15367 & ~n_15652;
assign n_15654 = ~n_15651 &  n_15653;
assign n_15655 = ~n_15642 & ~n_15654;
assign n_15656 =  x_1082 & ~n_15655;
assign n_15657 = ~x_1082 &  n_15655;
assign n_15658 = ~n_15656 & ~n_15657;
assign n_15659 =  x_1081 & ~n_15367;
assign n_15660 = ~x_3047 &  n_13143;
assign n_15661 = ~i_15 & ~n_13143;
assign n_15662 = ~n_13140 & ~n_15661;
assign n_15663 = ~n_15660 &  n_15662;
assign n_15664 =  x_2889 &  n_15373;
assign n_15665 =  x_3015 &  n_13141;
assign n_15666 = ~n_15375 & ~n_15665;
assign n_15667 = ~n_15664 &  n_15666;
assign n_15668 = ~n_15663 &  n_15667;
assign n_15669 = ~x_2825 &  n_15375;
assign n_15670 =  n_15367 & ~n_15669;
assign n_15671 = ~n_15668 &  n_15670;
assign n_15672 = ~n_15659 & ~n_15671;
assign n_15673 =  x_1081 & ~n_15672;
assign n_15674 = ~x_1081 &  n_15672;
assign n_15675 = ~n_15673 & ~n_15674;
assign n_15676 =  x_1080 & ~n_15367;
assign n_15677 = ~x_3046 &  n_13143;
assign n_15678 = ~i_14 & ~n_13143;
assign n_15679 = ~n_13140 & ~n_15678;
assign n_15680 = ~n_15677 &  n_15679;
assign n_15681 =  x_2888 &  n_15373;
assign n_15682 =  x_3014 &  n_13141;
assign n_15683 = ~n_15375 & ~n_15682;
assign n_15684 = ~n_15681 &  n_15683;
assign n_15685 = ~n_15680 &  n_15684;
assign n_15686 = ~x_2824 &  n_15375;
assign n_15687 =  n_15367 & ~n_15686;
assign n_15688 = ~n_15685 &  n_15687;
assign n_15689 = ~n_15676 & ~n_15688;
assign n_15690 =  x_1080 & ~n_15689;
assign n_15691 = ~x_1080 &  n_15689;
assign n_15692 = ~n_15690 & ~n_15691;
assign n_15693 =  x_1079 & ~n_15367;
assign n_15694 = ~x_3045 &  n_13143;
assign n_15695 = ~i_13 & ~n_13143;
assign n_15696 = ~n_13140 & ~n_15695;
assign n_15697 = ~n_15694 &  n_15696;
assign n_15698 =  x_2887 &  n_15373;
assign n_15699 =  x_3013 &  n_13141;
assign n_15700 = ~n_15375 & ~n_15699;
assign n_15701 = ~n_15698 &  n_15700;
assign n_15702 = ~n_15697 &  n_15701;
assign n_15703 = ~x_2823 &  n_15375;
assign n_15704 =  n_15367 & ~n_15703;
assign n_15705 = ~n_15702 &  n_15704;
assign n_15706 = ~n_15693 & ~n_15705;
assign n_15707 =  x_1079 & ~n_15706;
assign n_15708 = ~x_1079 &  n_15706;
assign n_15709 = ~n_15707 & ~n_15708;
assign n_15710 =  x_1078 & ~n_15367;
assign n_15711 = ~x_3044 &  n_13143;
assign n_15712 = ~i_12 & ~n_13143;
assign n_15713 = ~n_13140 & ~n_15712;
assign n_15714 = ~n_15711 &  n_15713;
assign n_15715 =  x_2886 &  n_15373;
assign n_15716 =  x_3012 &  n_13141;
assign n_15717 = ~n_15375 & ~n_15716;
assign n_15718 = ~n_15715 &  n_15717;
assign n_15719 = ~n_15714 &  n_15718;
assign n_15720 = ~x_2822 &  n_15375;
assign n_15721 =  n_15367 & ~n_15720;
assign n_15722 = ~n_15719 &  n_15721;
assign n_15723 = ~n_15710 & ~n_15722;
assign n_15724 =  x_1078 & ~n_15723;
assign n_15725 = ~x_1078 &  n_15723;
assign n_15726 = ~n_15724 & ~n_15725;
assign n_15727 =  x_1077 & ~n_15367;
assign n_15728 = ~x_3043 &  n_13143;
assign n_15729 = ~i_11 & ~n_13143;
assign n_15730 = ~n_13140 & ~n_15729;
assign n_15731 = ~n_15728 &  n_15730;
assign n_15732 =  x_2885 &  n_15373;
assign n_15733 =  x_3011 &  n_13141;
assign n_15734 = ~n_15375 & ~n_15733;
assign n_15735 = ~n_15732 &  n_15734;
assign n_15736 = ~n_15731 &  n_15735;
assign n_15737 = ~x_2821 &  n_15375;
assign n_15738 =  n_15367 & ~n_15737;
assign n_15739 = ~n_15736 &  n_15738;
assign n_15740 = ~n_15727 & ~n_15739;
assign n_15741 =  x_1077 & ~n_15740;
assign n_15742 = ~x_1077 &  n_15740;
assign n_15743 = ~n_15741 & ~n_15742;
assign n_15744 =  x_1076 & ~n_15367;
assign n_15745 = ~x_3042 &  n_13143;
assign n_15746 = ~i_10 & ~n_13143;
assign n_15747 = ~n_13140 & ~n_15746;
assign n_15748 = ~n_15745 &  n_15747;
assign n_15749 =  x_2884 &  n_15373;
assign n_15750 =  x_3010 &  n_13141;
assign n_15751 = ~n_15375 & ~n_15750;
assign n_15752 = ~n_15749 &  n_15751;
assign n_15753 = ~n_15748 &  n_15752;
assign n_15754 = ~x_2820 &  n_15375;
assign n_15755 =  n_15367 & ~n_15754;
assign n_15756 = ~n_15753 &  n_15755;
assign n_15757 = ~n_15744 & ~n_15756;
assign n_15758 =  x_1076 & ~n_15757;
assign n_15759 = ~x_1076 &  n_15757;
assign n_15760 = ~n_15758 & ~n_15759;
assign n_15761 =  x_1075 & ~n_15367;
assign n_15762 = ~x_3041 &  n_13143;
assign n_15763 = ~i_9 & ~n_13143;
assign n_15764 = ~n_13140 & ~n_15763;
assign n_15765 = ~n_15762 &  n_15764;
assign n_15766 =  x_2883 &  n_15373;
assign n_15767 =  x_3009 &  n_13141;
assign n_15768 = ~n_15375 & ~n_15767;
assign n_15769 = ~n_15766 &  n_15768;
assign n_15770 = ~n_15765 &  n_15769;
assign n_15771 = ~x_2819 &  n_15375;
assign n_15772 =  n_15367 & ~n_15771;
assign n_15773 = ~n_15770 &  n_15772;
assign n_15774 = ~n_15761 & ~n_15773;
assign n_15775 =  x_1075 & ~n_15774;
assign n_15776 = ~x_1075 &  n_15774;
assign n_15777 = ~n_15775 & ~n_15776;
assign n_15778 =  x_1074 & ~n_15367;
assign n_15779 = ~x_3040 &  n_13143;
assign n_15780 = ~i_8 & ~n_13143;
assign n_15781 = ~n_13140 & ~n_15780;
assign n_15782 = ~n_15779 &  n_15781;
assign n_15783 =  x_2882 &  n_15373;
assign n_15784 =  x_3008 &  n_13141;
assign n_15785 = ~n_15375 & ~n_15784;
assign n_15786 = ~n_15783 &  n_15785;
assign n_15787 = ~n_15782 &  n_15786;
assign n_15788 = ~x_2818 &  n_15375;
assign n_15789 =  n_15367 & ~n_15788;
assign n_15790 = ~n_15787 &  n_15789;
assign n_15791 = ~n_15778 & ~n_15790;
assign n_15792 =  x_1074 & ~n_15791;
assign n_15793 = ~x_1074 &  n_15791;
assign n_15794 = ~n_15792 & ~n_15793;
assign n_15795 =  x_1073 & ~n_15367;
assign n_15796 = ~x_3039 &  n_13143;
assign n_15797 = ~i_7 & ~n_13143;
assign n_15798 = ~n_13140 & ~n_15797;
assign n_15799 = ~n_15796 &  n_15798;
assign n_15800 =  x_2881 &  n_15373;
assign n_15801 =  x_3007 &  n_13141;
assign n_15802 = ~n_15375 & ~n_15801;
assign n_15803 = ~n_15800 &  n_15802;
assign n_15804 = ~n_15799 &  n_15803;
assign n_15805 = ~x_2817 &  n_15375;
assign n_15806 =  n_15367 & ~n_15805;
assign n_15807 = ~n_15804 &  n_15806;
assign n_15808 = ~n_15795 & ~n_15807;
assign n_15809 =  x_1073 & ~n_15808;
assign n_15810 = ~x_1073 &  n_15808;
assign n_15811 = ~n_15809 & ~n_15810;
assign n_15812 =  x_1072 & ~n_15367;
assign n_15813 = ~x_3038 &  n_13143;
assign n_15814 = ~i_6 & ~n_13143;
assign n_15815 = ~n_13140 & ~n_15814;
assign n_15816 = ~n_15813 &  n_15815;
assign n_15817 =  x_2880 &  n_15373;
assign n_15818 =  x_3006 &  n_13141;
assign n_15819 = ~n_15375 & ~n_15818;
assign n_15820 = ~n_15817 &  n_15819;
assign n_15821 = ~n_15816 &  n_15820;
assign n_15822 = ~x_2816 &  n_15375;
assign n_15823 =  n_15367 & ~n_15822;
assign n_15824 = ~n_15821 &  n_15823;
assign n_15825 = ~n_15812 & ~n_15824;
assign n_15826 =  x_1072 & ~n_15825;
assign n_15827 = ~x_1072 &  n_15825;
assign n_15828 = ~n_15826 & ~n_15827;
assign n_15829 =  x_1071 & ~n_15367;
assign n_15830 = ~x_3037 &  n_13143;
assign n_15831 = ~i_5 & ~n_13143;
assign n_15832 = ~n_13140 & ~n_15831;
assign n_15833 = ~n_15830 &  n_15832;
assign n_15834 =  x_2879 &  n_15373;
assign n_15835 =  x_3005 &  n_13141;
assign n_15836 = ~n_15375 & ~n_15835;
assign n_15837 = ~n_15834 &  n_15836;
assign n_15838 = ~n_15833 &  n_15837;
assign n_15839 = ~x_2815 &  n_15375;
assign n_15840 =  n_15367 & ~n_15839;
assign n_15841 = ~n_15838 &  n_15840;
assign n_15842 = ~n_15829 & ~n_15841;
assign n_15843 =  x_1071 & ~n_15842;
assign n_15844 = ~x_1071 &  n_15842;
assign n_15845 = ~n_15843 & ~n_15844;
assign n_15846 =  x_1070 & ~n_15367;
assign n_15847 = ~x_3036 &  n_13143;
assign n_15848 = ~i_4 & ~n_13143;
assign n_15849 = ~n_13140 & ~n_15848;
assign n_15850 = ~n_15847 &  n_15849;
assign n_15851 =  x_2878 &  n_15373;
assign n_15852 =  x_3004 &  n_13141;
assign n_15853 = ~n_15375 & ~n_15852;
assign n_15854 = ~n_15851 &  n_15853;
assign n_15855 = ~n_15850 &  n_15854;
assign n_15856 = ~x_2814 &  n_15375;
assign n_15857 =  n_15367 & ~n_15856;
assign n_15858 = ~n_15855 &  n_15857;
assign n_15859 = ~n_15846 & ~n_15858;
assign n_15860 =  x_1070 & ~n_15859;
assign n_15861 = ~x_1070 &  n_15859;
assign n_15862 = ~n_15860 & ~n_15861;
assign n_15863 =  x_1069 & ~n_15367;
assign n_15864 = ~x_3035 &  n_13143;
assign n_15865 = ~i_3 & ~n_13143;
assign n_15866 = ~n_13140 & ~n_15865;
assign n_15867 = ~n_15864 &  n_15866;
assign n_15868 =  x_2877 &  n_15373;
assign n_15869 =  x_3003 &  n_13141;
assign n_15870 = ~n_15375 & ~n_15869;
assign n_15871 = ~n_15868 &  n_15870;
assign n_15872 = ~n_15867 &  n_15871;
assign n_15873 = ~x_2813 &  n_15375;
assign n_15874 =  n_15367 & ~n_15873;
assign n_15875 = ~n_15872 &  n_15874;
assign n_15876 = ~n_15863 & ~n_15875;
assign n_15877 =  x_1069 & ~n_15876;
assign n_15878 = ~x_1069 &  n_15876;
assign n_15879 = ~n_15877 & ~n_15878;
assign n_15880 =  x_1068 & ~n_15367;
assign n_15881 = ~x_3034 &  n_13143;
assign n_15882 = ~i_2 & ~n_13143;
assign n_15883 = ~n_13140 & ~n_15882;
assign n_15884 = ~n_15881 &  n_15883;
assign n_15885 =  x_2876 &  n_15373;
assign n_15886 =  x_3002 &  n_13141;
assign n_15887 = ~n_15375 & ~n_15886;
assign n_15888 = ~n_15885 &  n_15887;
assign n_15889 = ~n_15884 &  n_15888;
assign n_15890 = ~x_2812 &  n_15375;
assign n_15891 =  n_15367 & ~n_15890;
assign n_15892 = ~n_15889 &  n_15891;
assign n_15893 = ~n_15880 & ~n_15892;
assign n_15894 =  x_1068 & ~n_15893;
assign n_15895 = ~x_1068 &  n_15893;
assign n_15896 = ~n_15894 & ~n_15895;
assign n_15897 =  x_1067 & ~n_15367;
assign n_15898 =  x_3033 &  n_13143;
assign n_15899 =  i_1 & ~n_13143;
assign n_15900 = ~n_15375 & ~n_13140;
assign n_15901 = ~n_15899 &  n_15900;
assign n_15902 = ~n_15898 &  n_15901;
assign n_15903 = ~x_2875 &  x_4775;
assign n_15904 = ~x_3001 & ~x_4775;
assign n_15905 = ~n_13135 &  n_15904;
assign n_15906 = ~n_15903 & ~n_15905;
assign n_15907 =  n_13140 & ~n_15906;
assign n_15908 = ~x_2811 &  n_15375;
assign n_15909 =  n_15367 & ~n_15908;
assign n_15910 = ~n_15907 &  n_15909;
assign n_15911 = ~n_15902 &  n_15910;
assign n_15912 = ~n_15897 & ~n_15911;
assign n_15913 =  x_1067 & ~n_15912;
assign n_15914 = ~x_1067 &  n_15912;
assign n_15915 = ~n_15913 & ~n_15914;
assign n_15916 =  n_759 &  n_767;
assign n_15917 = ~x_36 &  n_15916;
assign n_15918 =  n_1897 &  n_15917;
assign n_15919 =  n_2 &  n_15918;
assign n_15920 =  x_1066 & ~n_15919;
assign n_15921 =  x_4455 &  n_15919;
assign n_15922 = ~n_15920 & ~n_15921;
assign n_15923 =  x_1066 & ~n_15922;
assign n_15924 = ~x_1066 &  n_15922;
assign n_15925 = ~n_15923 & ~n_15924;
assign n_15926 =  x_1065 & ~n_15919;
assign n_15927 =  x_4454 &  n_15919;
assign n_15928 = ~n_15926 & ~n_15927;
assign n_15929 =  x_1065 & ~n_15928;
assign n_15930 = ~x_1065 &  n_15928;
assign n_15931 = ~n_15929 & ~n_15930;
assign n_15932 =  x_1064 & ~n_15919;
assign n_15933 =  x_4453 &  n_15919;
assign n_15934 = ~n_15932 & ~n_15933;
assign n_15935 =  x_1064 & ~n_15934;
assign n_15936 = ~x_1064 &  n_15934;
assign n_15937 = ~n_15935 & ~n_15936;
assign n_15938 =  x_1063 & ~n_15919;
assign n_15939 =  x_4452 &  n_15919;
assign n_15940 = ~n_15938 & ~n_15939;
assign n_15941 =  x_1063 & ~n_15940;
assign n_15942 = ~x_1063 &  n_15940;
assign n_15943 = ~n_15941 & ~n_15942;
assign n_15944 =  x_1062 & ~n_15919;
assign n_15945 =  x_4451 &  n_15919;
assign n_15946 = ~n_15944 & ~n_15945;
assign n_15947 =  x_1062 & ~n_15946;
assign n_15948 = ~x_1062 &  n_15946;
assign n_15949 = ~n_15947 & ~n_15948;
assign n_15950 =  x_1061 & ~n_15919;
assign n_15951 =  x_4450 &  n_15919;
assign n_15952 = ~n_15950 & ~n_15951;
assign n_15953 =  x_1061 & ~n_15952;
assign n_15954 = ~x_1061 &  n_15952;
assign n_15955 = ~n_15953 & ~n_15954;
assign n_15956 =  x_1060 & ~n_15919;
assign n_15957 =  x_4449 &  n_15919;
assign n_15958 = ~n_15956 & ~n_15957;
assign n_15959 =  x_1060 & ~n_15958;
assign n_15960 = ~x_1060 &  n_15958;
assign n_15961 = ~n_15959 & ~n_15960;
assign n_15962 =  x_1059 & ~n_15919;
assign n_15963 =  x_4448 &  n_15919;
assign n_15964 = ~n_15962 & ~n_15963;
assign n_15965 =  x_1059 & ~n_15964;
assign n_15966 = ~x_1059 &  n_15964;
assign n_15967 = ~n_15965 & ~n_15966;
assign n_15968 =  x_1058 & ~n_15919;
assign n_15969 =  x_4447 &  n_15919;
assign n_15970 = ~n_15968 & ~n_15969;
assign n_15971 =  x_1058 & ~n_15970;
assign n_15972 = ~x_1058 &  n_15970;
assign n_15973 = ~n_15971 & ~n_15972;
assign n_15974 =  x_1057 & ~n_15919;
assign n_15975 =  x_4446 &  n_15919;
assign n_15976 = ~n_15974 & ~n_15975;
assign n_15977 =  x_1057 & ~n_15976;
assign n_15978 = ~x_1057 &  n_15976;
assign n_15979 = ~n_15977 & ~n_15978;
assign n_15980 =  x_1056 & ~n_15919;
assign n_15981 =  x_4445 &  n_15919;
assign n_15982 = ~n_15980 & ~n_15981;
assign n_15983 =  x_1056 & ~n_15982;
assign n_15984 = ~x_1056 &  n_15982;
assign n_15985 = ~n_15983 & ~n_15984;
assign n_15986 =  x_1055 & ~n_15919;
assign n_15987 =  x_4444 &  n_15919;
assign n_15988 = ~n_15986 & ~n_15987;
assign n_15989 =  x_1055 & ~n_15988;
assign n_15990 = ~x_1055 &  n_15988;
assign n_15991 = ~n_15989 & ~n_15990;
assign n_15992 =  x_1054 & ~n_15919;
assign n_15993 =  x_4443 &  n_15919;
assign n_15994 = ~n_15992 & ~n_15993;
assign n_15995 =  x_1054 & ~n_15994;
assign n_15996 = ~x_1054 &  n_15994;
assign n_15997 = ~n_15995 & ~n_15996;
assign n_15998 =  x_1053 & ~n_15919;
assign n_15999 =  x_4442 &  n_15919;
assign n_16000 = ~n_15998 & ~n_15999;
assign n_16001 =  x_1053 & ~n_16000;
assign n_16002 = ~x_1053 &  n_16000;
assign n_16003 = ~n_16001 & ~n_16002;
assign n_16004 =  x_1052 & ~n_15919;
assign n_16005 =  x_4441 &  n_15919;
assign n_16006 = ~n_16004 & ~n_16005;
assign n_16007 =  x_1052 & ~n_16006;
assign n_16008 = ~x_1052 &  n_16006;
assign n_16009 = ~n_16007 & ~n_16008;
assign n_16010 =  x_1051 & ~n_15919;
assign n_16011 =  x_4440 &  n_15919;
assign n_16012 = ~n_16010 & ~n_16011;
assign n_16013 =  x_1051 & ~n_16012;
assign n_16014 = ~x_1051 &  n_16012;
assign n_16015 = ~n_16013 & ~n_16014;
assign n_16016 =  x_1050 & ~n_15919;
assign n_16017 =  x_4439 &  n_15919;
assign n_16018 = ~n_16016 & ~n_16017;
assign n_16019 =  x_1050 & ~n_16018;
assign n_16020 = ~x_1050 &  n_16018;
assign n_16021 = ~n_16019 & ~n_16020;
assign n_16022 =  x_1049 & ~n_15919;
assign n_16023 =  x_4438 &  n_15919;
assign n_16024 = ~n_16022 & ~n_16023;
assign n_16025 =  x_1049 & ~n_16024;
assign n_16026 = ~x_1049 &  n_16024;
assign n_16027 = ~n_16025 & ~n_16026;
assign n_16028 =  x_1048 & ~n_15919;
assign n_16029 =  x_4437 &  n_15919;
assign n_16030 = ~n_16028 & ~n_16029;
assign n_16031 =  x_1048 & ~n_16030;
assign n_16032 = ~x_1048 &  n_16030;
assign n_16033 = ~n_16031 & ~n_16032;
assign n_16034 =  x_1047 & ~n_15919;
assign n_16035 =  x_4436 &  n_15919;
assign n_16036 = ~n_16034 & ~n_16035;
assign n_16037 =  x_1047 & ~n_16036;
assign n_16038 = ~x_1047 &  n_16036;
assign n_16039 = ~n_16037 & ~n_16038;
assign n_16040 =  x_1046 & ~n_15919;
assign n_16041 =  x_4435 &  n_15919;
assign n_16042 = ~n_16040 & ~n_16041;
assign n_16043 =  x_1046 & ~n_16042;
assign n_16044 = ~x_1046 &  n_16042;
assign n_16045 = ~n_16043 & ~n_16044;
assign n_16046 =  x_1045 & ~n_15919;
assign n_16047 =  x_4434 &  n_15919;
assign n_16048 = ~n_16046 & ~n_16047;
assign n_16049 =  x_1045 & ~n_16048;
assign n_16050 = ~x_1045 &  n_16048;
assign n_16051 = ~n_16049 & ~n_16050;
assign n_16052 =  x_1044 & ~n_15919;
assign n_16053 =  x_4433 &  n_15919;
assign n_16054 = ~n_16052 & ~n_16053;
assign n_16055 =  x_1044 & ~n_16054;
assign n_16056 = ~x_1044 &  n_16054;
assign n_16057 = ~n_16055 & ~n_16056;
assign n_16058 =  x_1043 & ~n_15919;
assign n_16059 =  x_4432 &  n_15919;
assign n_16060 = ~n_16058 & ~n_16059;
assign n_16061 =  x_1043 & ~n_16060;
assign n_16062 = ~x_1043 &  n_16060;
assign n_16063 = ~n_16061 & ~n_16062;
assign n_16064 =  x_1042 & ~n_15919;
assign n_16065 =  x_4431 &  n_15919;
assign n_16066 = ~n_16064 & ~n_16065;
assign n_16067 =  x_1042 & ~n_16066;
assign n_16068 = ~x_1042 &  n_16066;
assign n_16069 = ~n_16067 & ~n_16068;
assign n_16070 =  x_1041 & ~n_15919;
assign n_16071 =  x_4430 &  n_15919;
assign n_16072 = ~n_16070 & ~n_16071;
assign n_16073 =  x_1041 & ~n_16072;
assign n_16074 = ~x_1041 &  n_16072;
assign n_16075 = ~n_16073 & ~n_16074;
assign n_16076 =  x_1040 & ~n_15919;
assign n_16077 =  x_4429 &  n_15919;
assign n_16078 = ~n_16076 & ~n_16077;
assign n_16079 =  x_1040 & ~n_16078;
assign n_16080 = ~x_1040 &  n_16078;
assign n_16081 = ~n_16079 & ~n_16080;
assign n_16082 =  x_1039 & ~n_15919;
assign n_16083 =  x_4428 &  n_15919;
assign n_16084 = ~n_16082 & ~n_16083;
assign n_16085 =  x_1039 & ~n_16084;
assign n_16086 = ~x_1039 &  n_16084;
assign n_16087 = ~n_16085 & ~n_16086;
assign n_16088 =  x_1038 & ~n_15919;
assign n_16089 =  x_4427 &  n_15919;
assign n_16090 = ~n_16088 & ~n_16089;
assign n_16091 =  x_1038 & ~n_16090;
assign n_16092 = ~x_1038 &  n_16090;
assign n_16093 = ~n_16091 & ~n_16092;
assign n_16094 =  x_1037 & ~n_15919;
assign n_16095 =  x_4426 &  n_15919;
assign n_16096 = ~n_16094 & ~n_16095;
assign n_16097 =  x_1037 & ~n_16096;
assign n_16098 = ~x_1037 &  n_16096;
assign n_16099 = ~n_16097 & ~n_16098;
assign n_16100 =  x_1036 & ~n_15919;
assign n_16101 =  x_4425 &  n_15919;
assign n_16102 = ~n_16100 & ~n_16101;
assign n_16103 =  x_1036 & ~n_16102;
assign n_16104 = ~x_1036 &  n_16102;
assign n_16105 = ~n_16103 & ~n_16104;
assign n_16106 =  x_1035 & ~n_15919;
assign n_16107 =  x_1035 &  n_16106;
assign n_16108 = ~x_1035 & ~n_16106;
assign n_16109 = ~n_16107 & ~n_16108;
assign n_16110 =  n_152 &  n_15918;
assign n_16111 =  x_43 &  n_16110;
assign n_16112 =  x_1034 & ~n_16111;
assign n_16113 =  x_3223 &  n_16111;
assign n_16114 = ~n_16112 & ~n_16113;
assign n_16115 =  x_1034 & ~n_16114;
assign n_16116 = ~x_1034 &  n_16114;
assign n_16117 = ~n_16115 & ~n_16116;
assign n_16118 =  x_1033 & ~n_16111;
assign n_16119 =  x_3222 &  n_16111;
assign n_16120 = ~n_16118 & ~n_16119;
assign n_16121 =  x_1033 & ~n_16120;
assign n_16122 = ~x_1033 &  n_16120;
assign n_16123 = ~n_16121 & ~n_16122;
assign n_16124 =  x_1032 & ~n_16111;
assign n_16125 =  x_3221 &  n_16111;
assign n_16126 = ~n_16124 & ~n_16125;
assign n_16127 =  x_1032 & ~n_16126;
assign n_16128 = ~x_1032 &  n_16126;
assign n_16129 = ~n_16127 & ~n_16128;
assign n_16130 =  x_1031 & ~n_16111;
assign n_16131 =  x_3220 &  n_16111;
assign n_16132 = ~n_16130 & ~n_16131;
assign n_16133 =  x_1031 & ~n_16132;
assign n_16134 = ~x_1031 &  n_16132;
assign n_16135 = ~n_16133 & ~n_16134;
assign n_16136 =  x_1030 & ~n_16111;
assign n_16137 =  x_3219 &  n_16111;
assign n_16138 = ~n_16136 & ~n_16137;
assign n_16139 =  x_1030 & ~n_16138;
assign n_16140 = ~x_1030 &  n_16138;
assign n_16141 = ~n_16139 & ~n_16140;
assign n_16142 =  x_1029 & ~n_16111;
assign n_16143 =  x_3218 &  n_16111;
assign n_16144 = ~n_16142 & ~n_16143;
assign n_16145 =  x_1029 & ~n_16144;
assign n_16146 = ~x_1029 &  n_16144;
assign n_16147 = ~n_16145 & ~n_16146;
assign n_16148 =  x_1028 & ~n_16111;
assign n_16149 =  x_3217 &  n_16111;
assign n_16150 = ~n_16148 & ~n_16149;
assign n_16151 =  x_1028 & ~n_16150;
assign n_16152 = ~x_1028 &  n_16150;
assign n_16153 = ~n_16151 & ~n_16152;
assign n_16154 =  x_1027 & ~n_16111;
assign n_16155 =  x_3216 &  n_16111;
assign n_16156 = ~n_16154 & ~n_16155;
assign n_16157 =  x_1027 & ~n_16156;
assign n_16158 = ~x_1027 &  n_16156;
assign n_16159 = ~n_16157 & ~n_16158;
assign n_16160 =  x_1026 & ~n_16111;
assign n_16161 =  x_3215 &  n_16111;
assign n_16162 = ~n_16160 & ~n_16161;
assign n_16163 =  x_1026 & ~n_16162;
assign n_16164 = ~x_1026 &  n_16162;
assign n_16165 = ~n_16163 & ~n_16164;
assign n_16166 =  x_1025 & ~n_16111;
assign n_16167 =  x_3214 &  n_16111;
assign n_16168 = ~n_16166 & ~n_16167;
assign n_16169 =  x_1025 & ~n_16168;
assign n_16170 = ~x_1025 &  n_16168;
assign n_16171 = ~n_16169 & ~n_16170;
assign n_16172 =  x_1024 & ~n_16111;
assign n_16173 =  x_3213 &  n_16111;
assign n_16174 = ~n_16172 & ~n_16173;
assign n_16175 =  x_1024 & ~n_16174;
assign n_16176 = ~x_1024 &  n_16174;
assign n_16177 = ~n_16175 & ~n_16176;
assign n_16178 =  x_1023 & ~n_16111;
assign n_16179 =  x_3212 &  n_16111;
assign n_16180 = ~n_16178 & ~n_16179;
assign n_16181 =  x_1023 & ~n_16180;
assign n_16182 = ~x_1023 &  n_16180;
assign n_16183 = ~n_16181 & ~n_16182;
assign n_16184 =  x_1022 & ~n_16111;
assign n_16185 =  x_3211 &  n_16111;
assign n_16186 = ~n_16184 & ~n_16185;
assign n_16187 =  x_1022 & ~n_16186;
assign n_16188 = ~x_1022 &  n_16186;
assign n_16189 = ~n_16187 & ~n_16188;
assign n_16190 =  x_1021 & ~n_16111;
assign n_16191 =  x_3210 &  n_16111;
assign n_16192 = ~n_16190 & ~n_16191;
assign n_16193 =  x_1021 & ~n_16192;
assign n_16194 = ~x_1021 &  n_16192;
assign n_16195 = ~n_16193 & ~n_16194;
assign n_16196 =  x_1020 & ~n_16111;
assign n_16197 =  x_3209 &  n_16111;
assign n_16198 = ~n_16196 & ~n_16197;
assign n_16199 =  x_1020 & ~n_16198;
assign n_16200 = ~x_1020 &  n_16198;
assign n_16201 = ~n_16199 & ~n_16200;
assign n_16202 =  x_1019 & ~n_16111;
assign n_16203 =  x_3208 &  n_16111;
assign n_16204 = ~n_16202 & ~n_16203;
assign n_16205 =  x_1019 & ~n_16204;
assign n_16206 = ~x_1019 &  n_16204;
assign n_16207 = ~n_16205 & ~n_16206;
assign n_16208 =  x_1018 & ~n_16111;
assign n_16209 =  x_3207 &  n_16111;
assign n_16210 = ~n_16208 & ~n_16209;
assign n_16211 =  x_1018 & ~n_16210;
assign n_16212 = ~x_1018 &  n_16210;
assign n_16213 = ~n_16211 & ~n_16212;
assign n_16214 =  x_1017 & ~n_16111;
assign n_16215 =  x_3206 &  n_16111;
assign n_16216 = ~n_16214 & ~n_16215;
assign n_16217 =  x_1017 & ~n_16216;
assign n_16218 = ~x_1017 &  n_16216;
assign n_16219 = ~n_16217 & ~n_16218;
assign n_16220 =  x_1016 & ~n_16111;
assign n_16221 =  x_3205 &  n_16111;
assign n_16222 = ~n_16220 & ~n_16221;
assign n_16223 =  x_1016 & ~n_16222;
assign n_16224 = ~x_1016 &  n_16222;
assign n_16225 = ~n_16223 & ~n_16224;
assign n_16226 =  x_1015 & ~n_16111;
assign n_16227 =  x_3204 &  n_16111;
assign n_16228 = ~n_16226 & ~n_16227;
assign n_16229 =  x_1015 & ~n_16228;
assign n_16230 = ~x_1015 &  n_16228;
assign n_16231 = ~n_16229 & ~n_16230;
assign n_16232 =  x_1014 & ~n_16111;
assign n_16233 =  x_3203 &  n_16111;
assign n_16234 = ~n_16232 & ~n_16233;
assign n_16235 =  x_1014 & ~n_16234;
assign n_16236 = ~x_1014 &  n_16234;
assign n_16237 = ~n_16235 & ~n_16236;
assign n_16238 =  x_1013 & ~n_16111;
assign n_16239 =  x_3202 &  n_16111;
assign n_16240 = ~n_16238 & ~n_16239;
assign n_16241 =  x_1013 & ~n_16240;
assign n_16242 = ~x_1013 &  n_16240;
assign n_16243 = ~n_16241 & ~n_16242;
assign n_16244 =  x_1012 & ~n_16111;
assign n_16245 =  x_3201 &  n_16111;
assign n_16246 = ~n_16244 & ~n_16245;
assign n_16247 =  x_1012 & ~n_16246;
assign n_16248 = ~x_1012 &  n_16246;
assign n_16249 = ~n_16247 & ~n_16248;
assign n_16250 =  x_1011 & ~n_16111;
assign n_16251 =  x_3200 &  n_16111;
assign n_16252 = ~n_16250 & ~n_16251;
assign n_16253 =  x_1011 & ~n_16252;
assign n_16254 = ~x_1011 &  n_16252;
assign n_16255 = ~n_16253 & ~n_16254;
assign n_16256 =  x_1010 & ~n_16111;
assign n_16257 =  x_3199 &  n_16111;
assign n_16258 = ~n_16256 & ~n_16257;
assign n_16259 =  x_1010 & ~n_16258;
assign n_16260 = ~x_1010 &  n_16258;
assign n_16261 = ~n_16259 & ~n_16260;
assign n_16262 =  x_1009 & ~n_16111;
assign n_16263 =  x_3198 &  n_16111;
assign n_16264 = ~n_16262 & ~n_16263;
assign n_16265 =  x_1009 & ~n_16264;
assign n_16266 = ~x_1009 &  n_16264;
assign n_16267 = ~n_16265 & ~n_16266;
assign n_16268 =  x_1008 & ~n_16111;
assign n_16269 =  x_3197 &  n_16111;
assign n_16270 = ~n_16268 & ~n_16269;
assign n_16271 =  x_1008 & ~n_16270;
assign n_16272 = ~x_1008 &  n_16270;
assign n_16273 = ~n_16271 & ~n_16272;
assign n_16274 =  x_1007 & ~n_16111;
assign n_16275 =  x_3196 &  n_16111;
assign n_16276 = ~n_16274 & ~n_16275;
assign n_16277 =  x_1007 & ~n_16276;
assign n_16278 = ~x_1007 &  n_16276;
assign n_16279 = ~n_16277 & ~n_16278;
assign n_16280 =  x_1006 & ~n_16111;
assign n_16281 =  x_3195 &  n_16111;
assign n_16282 = ~n_16280 & ~n_16281;
assign n_16283 =  x_1006 & ~n_16282;
assign n_16284 = ~x_1006 &  n_16282;
assign n_16285 = ~n_16283 & ~n_16284;
assign n_16286 =  x_1005 & ~n_16111;
assign n_16287 =  x_3194 &  n_16111;
assign n_16288 = ~n_16286 & ~n_16287;
assign n_16289 =  x_1005 & ~n_16288;
assign n_16290 = ~x_1005 &  n_16288;
assign n_16291 = ~n_16289 & ~n_16290;
assign n_16292 =  x_1004 & ~n_16111;
assign n_16293 =  x_3193 &  n_16111;
assign n_16294 = ~n_16292 & ~n_16293;
assign n_16295 =  x_1004 & ~n_16294;
assign n_16296 = ~x_1004 &  n_16294;
assign n_16297 = ~n_16295 & ~n_16296;
assign n_16298 =  x_1003 & ~n_16111;
assign n_16299 =  x_1003 &  n_16298;
assign n_16300 = ~x_1003 & ~n_16298;
assign n_16301 = ~n_16299 & ~n_16300;
assign n_16302 =  n_6525 &  n_6182;
assign n_16303 =  x_1002 & ~n_16302;
assign n_16304 =  i_32 &  n_16302;
assign n_16305 = ~n_16303 & ~n_16304;
assign n_16306 =  x_1002 & ~n_16305;
assign n_16307 = ~x_1002 &  n_16305;
assign n_16308 = ~n_16306 & ~n_16307;
assign n_16309 =  x_1001 & ~n_16302;
assign n_16310 =  i_31 &  n_16302;
assign n_16311 = ~n_16309 & ~n_16310;
assign n_16312 =  x_1001 & ~n_16311;
assign n_16313 = ~x_1001 &  n_16311;
assign n_16314 = ~n_16312 & ~n_16313;
assign n_16315 =  x_1000 & ~n_16302;
assign n_16316 =  i_30 &  n_16302;
assign n_16317 = ~n_16315 & ~n_16316;
assign n_16318 =  x_1000 & ~n_16317;
assign n_16319 = ~x_1000 &  n_16317;
assign n_16320 = ~n_16318 & ~n_16319;
assign n_16321 =  x_999 & ~n_16302;
assign n_16322 =  i_29 &  n_16302;
assign n_16323 = ~n_16321 & ~n_16322;
assign n_16324 =  x_999 & ~n_16323;
assign n_16325 = ~x_999 &  n_16323;
assign n_16326 = ~n_16324 & ~n_16325;
assign n_16327 =  x_998 & ~n_16302;
assign n_16328 =  i_28 &  n_16302;
assign n_16329 = ~n_16327 & ~n_16328;
assign n_16330 =  x_998 & ~n_16329;
assign n_16331 = ~x_998 &  n_16329;
assign n_16332 = ~n_16330 & ~n_16331;
assign n_16333 =  x_997 & ~n_16302;
assign n_16334 =  i_27 &  n_16302;
assign n_16335 = ~n_16333 & ~n_16334;
assign n_16336 =  x_997 & ~n_16335;
assign n_16337 = ~x_997 &  n_16335;
assign n_16338 = ~n_16336 & ~n_16337;
assign n_16339 =  x_996 & ~n_16302;
assign n_16340 =  i_26 &  n_16302;
assign n_16341 = ~n_16339 & ~n_16340;
assign n_16342 =  x_996 & ~n_16341;
assign n_16343 = ~x_996 &  n_16341;
assign n_16344 = ~n_16342 & ~n_16343;
assign n_16345 =  x_995 & ~n_16302;
assign n_16346 =  i_25 &  n_16302;
assign n_16347 = ~n_16345 & ~n_16346;
assign n_16348 =  x_995 & ~n_16347;
assign n_16349 = ~x_995 &  n_16347;
assign n_16350 = ~n_16348 & ~n_16349;
assign n_16351 =  x_994 & ~n_16302;
assign n_16352 =  i_24 &  n_16302;
assign n_16353 = ~n_16351 & ~n_16352;
assign n_16354 =  x_994 & ~n_16353;
assign n_16355 = ~x_994 &  n_16353;
assign n_16356 = ~n_16354 & ~n_16355;
assign n_16357 =  x_993 & ~n_16302;
assign n_16358 =  i_23 &  n_16302;
assign n_16359 = ~n_16357 & ~n_16358;
assign n_16360 =  x_993 & ~n_16359;
assign n_16361 = ~x_993 &  n_16359;
assign n_16362 = ~n_16360 & ~n_16361;
assign n_16363 =  x_992 & ~n_16302;
assign n_16364 =  i_22 &  n_16302;
assign n_16365 = ~n_16363 & ~n_16364;
assign n_16366 =  x_992 & ~n_16365;
assign n_16367 = ~x_992 &  n_16365;
assign n_16368 = ~n_16366 & ~n_16367;
assign n_16369 =  x_991 & ~n_16302;
assign n_16370 =  i_21 &  n_16302;
assign n_16371 = ~n_16369 & ~n_16370;
assign n_16372 =  x_991 & ~n_16371;
assign n_16373 = ~x_991 &  n_16371;
assign n_16374 = ~n_16372 & ~n_16373;
assign n_16375 =  x_990 & ~n_16302;
assign n_16376 =  i_20 &  n_16302;
assign n_16377 = ~n_16375 & ~n_16376;
assign n_16378 =  x_990 & ~n_16377;
assign n_16379 = ~x_990 &  n_16377;
assign n_16380 = ~n_16378 & ~n_16379;
assign n_16381 =  x_989 & ~n_16302;
assign n_16382 =  i_19 &  n_16302;
assign n_16383 = ~n_16381 & ~n_16382;
assign n_16384 =  x_989 & ~n_16383;
assign n_16385 = ~x_989 &  n_16383;
assign n_16386 = ~n_16384 & ~n_16385;
assign n_16387 =  x_988 & ~n_16302;
assign n_16388 =  i_18 &  n_16302;
assign n_16389 = ~n_16387 & ~n_16388;
assign n_16390 =  x_988 & ~n_16389;
assign n_16391 = ~x_988 &  n_16389;
assign n_16392 = ~n_16390 & ~n_16391;
assign n_16393 =  x_987 & ~n_16302;
assign n_16394 =  i_17 &  n_16302;
assign n_16395 = ~n_16393 & ~n_16394;
assign n_16396 =  x_987 & ~n_16395;
assign n_16397 = ~x_987 &  n_16395;
assign n_16398 = ~n_16396 & ~n_16397;
assign n_16399 =  x_986 & ~n_16302;
assign n_16400 =  i_16 &  n_16302;
assign n_16401 = ~n_16399 & ~n_16400;
assign n_16402 =  x_986 & ~n_16401;
assign n_16403 = ~x_986 &  n_16401;
assign n_16404 = ~n_16402 & ~n_16403;
assign n_16405 =  x_985 & ~n_16302;
assign n_16406 =  i_15 &  n_16302;
assign n_16407 = ~n_16405 & ~n_16406;
assign n_16408 =  x_985 & ~n_16407;
assign n_16409 = ~x_985 &  n_16407;
assign n_16410 = ~n_16408 & ~n_16409;
assign n_16411 =  x_984 & ~n_16302;
assign n_16412 =  i_14 &  n_16302;
assign n_16413 = ~n_16411 & ~n_16412;
assign n_16414 =  x_984 & ~n_16413;
assign n_16415 = ~x_984 &  n_16413;
assign n_16416 = ~n_16414 & ~n_16415;
assign n_16417 =  x_983 & ~n_16302;
assign n_16418 =  i_13 &  n_16302;
assign n_16419 = ~n_16417 & ~n_16418;
assign n_16420 =  x_983 & ~n_16419;
assign n_16421 = ~x_983 &  n_16419;
assign n_16422 = ~n_16420 & ~n_16421;
assign n_16423 =  x_982 & ~n_16302;
assign n_16424 =  i_12 &  n_16302;
assign n_16425 = ~n_16423 & ~n_16424;
assign n_16426 =  x_982 & ~n_16425;
assign n_16427 = ~x_982 &  n_16425;
assign n_16428 = ~n_16426 & ~n_16427;
assign n_16429 =  x_981 & ~n_16302;
assign n_16430 =  i_11 &  n_16302;
assign n_16431 = ~n_16429 & ~n_16430;
assign n_16432 =  x_981 & ~n_16431;
assign n_16433 = ~x_981 &  n_16431;
assign n_16434 = ~n_16432 & ~n_16433;
assign n_16435 =  x_980 & ~n_16302;
assign n_16436 =  i_10 &  n_16302;
assign n_16437 = ~n_16435 & ~n_16436;
assign n_16438 =  x_980 & ~n_16437;
assign n_16439 = ~x_980 &  n_16437;
assign n_16440 = ~n_16438 & ~n_16439;
assign n_16441 =  x_979 & ~n_16302;
assign n_16442 =  i_9 &  n_16302;
assign n_16443 = ~n_16441 & ~n_16442;
assign n_16444 =  x_979 & ~n_16443;
assign n_16445 = ~x_979 &  n_16443;
assign n_16446 = ~n_16444 & ~n_16445;
assign n_16447 =  x_978 & ~n_16302;
assign n_16448 =  i_8 &  n_16302;
assign n_16449 = ~n_16447 & ~n_16448;
assign n_16450 =  x_978 & ~n_16449;
assign n_16451 = ~x_978 &  n_16449;
assign n_16452 = ~n_16450 & ~n_16451;
assign n_16453 =  x_977 & ~n_16302;
assign n_16454 =  i_7 &  n_16302;
assign n_16455 = ~n_16453 & ~n_16454;
assign n_16456 =  x_977 & ~n_16455;
assign n_16457 = ~x_977 &  n_16455;
assign n_16458 = ~n_16456 & ~n_16457;
assign n_16459 =  x_976 & ~n_16302;
assign n_16460 =  i_6 &  n_16302;
assign n_16461 = ~n_16459 & ~n_16460;
assign n_16462 =  x_976 & ~n_16461;
assign n_16463 = ~x_976 &  n_16461;
assign n_16464 = ~n_16462 & ~n_16463;
assign n_16465 =  x_975 & ~n_16302;
assign n_16466 =  i_5 &  n_16302;
assign n_16467 = ~n_16465 & ~n_16466;
assign n_16468 =  x_975 & ~n_16467;
assign n_16469 = ~x_975 &  n_16467;
assign n_16470 = ~n_16468 & ~n_16469;
assign n_16471 =  x_974 & ~n_16302;
assign n_16472 =  i_4 &  n_16302;
assign n_16473 = ~n_16471 & ~n_16472;
assign n_16474 =  x_974 & ~n_16473;
assign n_16475 = ~x_974 &  n_16473;
assign n_16476 = ~n_16474 & ~n_16475;
assign n_16477 =  x_973 & ~n_16302;
assign n_16478 =  i_3 &  n_16302;
assign n_16479 = ~n_16477 & ~n_16478;
assign n_16480 =  x_973 & ~n_16479;
assign n_16481 = ~x_973 &  n_16479;
assign n_16482 = ~n_16480 & ~n_16481;
assign n_16483 =  x_972 & ~n_16302;
assign n_16484 =  i_2 &  n_16302;
assign n_16485 = ~n_16483 & ~n_16484;
assign n_16486 =  x_972 & ~n_16485;
assign n_16487 = ~x_972 &  n_16485;
assign n_16488 = ~n_16486 & ~n_16487;
assign n_16489 =  x_971 & ~n_16302;
assign n_16490 =  i_1 &  n_16302;
assign n_16491 = ~n_16489 & ~n_16490;
assign n_16492 =  x_971 & ~n_16491;
assign n_16493 = ~x_971 &  n_16491;
assign n_16494 = ~n_16492 & ~n_16493;
assign n_16495 =  n_151 &  n_15366;
assign n_16496 =  n_6379 &  n_16495;
assign n_16497 =  x_970 & ~n_16496;
assign n_16498 =  i_32 &  n_16496;
assign n_16499 = ~n_16497 & ~n_16498;
assign n_16500 =  x_970 & ~n_16499;
assign n_16501 = ~x_970 &  n_16499;
assign n_16502 = ~n_16500 & ~n_16501;
assign n_16503 =  x_969 & ~n_16496;
assign n_16504 =  i_31 &  n_16496;
assign n_16505 = ~n_16503 & ~n_16504;
assign n_16506 =  x_969 & ~n_16505;
assign n_16507 = ~x_969 &  n_16505;
assign n_16508 = ~n_16506 & ~n_16507;
assign n_16509 =  x_968 & ~n_16496;
assign n_16510 =  i_30 &  n_16496;
assign n_16511 = ~n_16509 & ~n_16510;
assign n_16512 =  x_968 & ~n_16511;
assign n_16513 = ~x_968 &  n_16511;
assign n_16514 = ~n_16512 & ~n_16513;
assign n_16515 =  x_967 & ~n_16496;
assign n_16516 =  i_29 &  n_16496;
assign n_16517 = ~n_16515 & ~n_16516;
assign n_16518 =  x_967 & ~n_16517;
assign n_16519 = ~x_967 &  n_16517;
assign n_16520 = ~n_16518 & ~n_16519;
assign n_16521 =  x_966 & ~n_16496;
assign n_16522 =  i_28 &  n_16496;
assign n_16523 = ~n_16521 & ~n_16522;
assign n_16524 =  x_966 & ~n_16523;
assign n_16525 = ~x_966 &  n_16523;
assign n_16526 = ~n_16524 & ~n_16525;
assign n_16527 =  x_965 & ~n_16496;
assign n_16528 =  i_27 &  n_16496;
assign n_16529 = ~n_16527 & ~n_16528;
assign n_16530 =  x_965 & ~n_16529;
assign n_16531 = ~x_965 &  n_16529;
assign n_16532 = ~n_16530 & ~n_16531;
assign n_16533 =  x_964 & ~n_16496;
assign n_16534 =  i_26 &  n_16496;
assign n_16535 = ~n_16533 & ~n_16534;
assign n_16536 =  x_964 & ~n_16535;
assign n_16537 = ~x_964 &  n_16535;
assign n_16538 = ~n_16536 & ~n_16537;
assign n_16539 =  x_963 & ~n_16496;
assign n_16540 =  i_25 &  n_16496;
assign n_16541 = ~n_16539 & ~n_16540;
assign n_16542 =  x_963 & ~n_16541;
assign n_16543 = ~x_963 &  n_16541;
assign n_16544 = ~n_16542 & ~n_16543;
assign n_16545 =  x_962 & ~n_16496;
assign n_16546 =  i_24 &  n_16496;
assign n_16547 = ~n_16545 & ~n_16546;
assign n_16548 =  x_962 & ~n_16547;
assign n_16549 = ~x_962 &  n_16547;
assign n_16550 = ~n_16548 & ~n_16549;
assign n_16551 =  x_961 & ~n_16496;
assign n_16552 =  i_23 &  n_16496;
assign n_16553 = ~n_16551 & ~n_16552;
assign n_16554 =  x_961 & ~n_16553;
assign n_16555 = ~x_961 &  n_16553;
assign n_16556 = ~n_16554 & ~n_16555;
assign n_16557 =  x_960 & ~n_16496;
assign n_16558 =  i_22 &  n_16496;
assign n_16559 = ~n_16557 & ~n_16558;
assign n_16560 =  x_960 & ~n_16559;
assign n_16561 = ~x_960 &  n_16559;
assign n_16562 = ~n_16560 & ~n_16561;
assign n_16563 =  x_959 & ~n_16496;
assign n_16564 =  i_21 &  n_16496;
assign n_16565 = ~n_16563 & ~n_16564;
assign n_16566 =  x_959 & ~n_16565;
assign n_16567 = ~x_959 &  n_16565;
assign n_16568 = ~n_16566 & ~n_16567;
assign n_16569 =  x_958 & ~n_16496;
assign n_16570 =  i_20 &  n_16496;
assign n_16571 = ~n_16569 & ~n_16570;
assign n_16572 =  x_958 & ~n_16571;
assign n_16573 = ~x_958 &  n_16571;
assign n_16574 = ~n_16572 & ~n_16573;
assign n_16575 =  x_957 & ~n_16496;
assign n_16576 =  i_19 &  n_16496;
assign n_16577 = ~n_16575 & ~n_16576;
assign n_16578 =  x_957 & ~n_16577;
assign n_16579 = ~x_957 &  n_16577;
assign n_16580 = ~n_16578 & ~n_16579;
assign n_16581 =  x_956 & ~n_16496;
assign n_16582 =  i_18 &  n_16496;
assign n_16583 = ~n_16581 & ~n_16582;
assign n_16584 =  x_956 & ~n_16583;
assign n_16585 = ~x_956 &  n_16583;
assign n_16586 = ~n_16584 & ~n_16585;
assign n_16587 =  x_955 & ~n_16496;
assign n_16588 =  i_17 &  n_16496;
assign n_16589 = ~n_16587 & ~n_16588;
assign n_16590 =  x_955 & ~n_16589;
assign n_16591 = ~x_955 &  n_16589;
assign n_16592 = ~n_16590 & ~n_16591;
assign n_16593 =  x_954 & ~n_16496;
assign n_16594 =  i_16 &  n_16496;
assign n_16595 = ~n_16593 & ~n_16594;
assign n_16596 =  x_954 & ~n_16595;
assign n_16597 = ~x_954 &  n_16595;
assign n_16598 = ~n_16596 & ~n_16597;
assign n_16599 =  x_953 & ~n_16496;
assign n_16600 =  i_15 &  n_16496;
assign n_16601 = ~n_16599 & ~n_16600;
assign n_16602 =  x_953 & ~n_16601;
assign n_16603 = ~x_953 &  n_16601;
assign n_16604 = ~n_16602 & ~n_16603;
assign n_16605 =  x_952 & ~n_16496;
assign n_16606 =  i_14 &  n_16496;
assign n_16607 = ~n_16605 & ~n_16606;
assign n_16608 =  x_952 & ~n_16607;
assign n_16609 = ~x_952 &  n_16607;
assign n_16610 = ~n_16608 & ~n_16609;
assign n_16611 =  x_951 & ~n_16496;
assign n_16612 =  i_13 &  n_16496;
assign n_16613 = ~n_16611 & ~n_16612;
assign n_16614 =  x_951 & ~n_16613;
assign n_16615 = ~x_951 &  n_16613;
assign n_16616 = ~n_16614 & ~n_16615;
assign n_16617 =  x_950 & ~n_16496;
assign n_16618 =  i_12 &  n_16496;
assign n_16619 = ~n_16617 & ~n_16618;
assign n_16620 =  x_950 & ~n_16619;
assign n_16621 = ~x_950 &  n_16619;
assign n_16622 = ~n_16620 & ~n_16621;
assign n_16623 =  x_949 & ~n_16496;
assign n_16624 =  i_11 &  n_16496;
assign n_16625 = ~n_16623 & ~n_16624;
assign n_16626 =  x_949 & ~n_16625;
assign n_16627 = ~x_949 &  n_16625;
assign n_16628 = ~n_16626 & ~n_16627;
assign n_16629 =  x_948 & ~n_16496;
assign n_16630 =  i_10 &  n_16496;
assign n_16631 = ~n_16629 & ~n_16630;
assign n_16632 =  x_948 & ~n_16631;
assign n_16633 = ~x_948 &  n_16631;
assign n_16634 = ~n_16632 & ~n_16633;
assign n_16635 =  x_947 & ~n_16496;
assign n_16636 =  i_9 &  n_16496;
assign n_16637 = ~n_16635 & ~n_16636;
assign n_16638 =  x_947 & ~n_16637;
assign n_16639 = ~x_947 &  n_16637;
assign n_16640 = ~n_16638 & ~n_16639;
assign n_16641 =  x_946 & ~n_16496;
assign n_16642 =  i_8 &  n_16496;
assign n_16643 = ~n_16641 & ~n_16642;
assign n_16644 =  x_946 & ~n_16643;
assign n_16645 = ~x_946 &  n_16643;
assign n_16646 = ~n_16644 & ~n_16645;
assign n_16647 =  x_945 & ~n_16496;
assign n_16648 =  i_7 &  n_16496;
assign n_16649 = ~n_16647 & ~n_16648;
assign n_16650 =  x_945 & ~n_16649;
assign n_16651 = ~x_945 &  n_16649;
assign n_16652 = ~n_16650 & ~n_16651;
assign n_16653 =  x_944 & ~n_16496;
assign n_16654 =  i_6 &  n_16496;
assign n_16655 = ~n_16653 & ~n_16654;
assign n_16656 =  x_944 & ~n_16655;
assign n_16657 = ~x_944 &  n_16655;
assign n_16658 = ~n_16656 & ~n_16657;
assign n_16659 =  x_943 & ~n_16496;
assign n_16660 =  i_5 &  n_16496;
assign n_16661 = ~n_16659 & ~n_16660;
assign n_16662 =  x_943 & ~n_16661;
assign n_16663 = ~x_943 &  n_16661;
assign n_16664 = ~n_16662 & ~n_16663;
assign n_16665 =  x_942 & ~n_16496;
assign n_16666 =  i_4 &  n_16496;
assign n_16667 = ~n_16665 & ~n_16666;
assign n_16668 =  x_942 & ~n_16667;
assign n_16669 = ~x_942 &  n_16667;
assign n_16670 = ~n_16668 & ~n_16669;
assign n_16671 =  x_941 & ~n_16496;
assign n_16672 =  i_3 &  n_16496;
assign n_16673 = ~n_16671 & ~n_16672;
assign n_16674 =  x_941 & ~n_16673;
assign n_16675 = ~x_941 &  n_16673;
assign n_16676 = ~n_16674 & ~n_16675;
assign n_16677 =  x_940 & ~n_16496;
assign n_16678 =  i_2 &  n_16496;
assign n_16679 = ~n_16677 & ~n_16678;
assign n_16680 =  x_940 & ~n_16679;
assign n_16681 = ~x_940 &  n_16679;
assign n_16682 = ~n_16680 & ~n_16681;
assign n_16683 =  x_939 & ~n_16496;
assign n_16684 =  i_1 &  n_16496;
assign n_16685 = ~n_16683 & ~n_16684;
assign n_16686 =  x_939 & ~n_16685;
assign n_16687 = ~x_939 &  n_16685;
assign n_16688 = ~n_16686 & ~n_16687;
assign n_16689 =  n_1895 &  n_2487;
assign n_16690 =  x_938 & ~n_16689;
assign n_16691 =  i_32 &  n_16689;
assign n_16692 = ~n_16690 & ~n_16691;
assign n_16693 =  x_938 & ~n_16692;
assign n_16694 = ~x_938 &  n_16692;
assign n_16695 = ~n_16693 & ~n_16694;
assign n_16696 =  x_937 & ~n_16689;
assign n_16697 =  i_31 &  n_16689;
assign n_16698 = ~n_16696 & ~n_16697;
assign n_16699 =  x_937 & ~n_16698;
assign n_16700 = ~x_937 &  n_16698;
assign n_16701 = ~n_16699 & ~n_16700;
assign n_16702 =  x_936 & ~n_16689;
assign n_16703 =  i_30 &  n_16689;
assign n_16704 = ~n_16702 & ~n_16703;
assign n_16705 =  x_936 & ~n_16704;
assign n_16706 = ~x_936 &  n_16704;
assign n_16707 = ~n_16705 & ~n_16706;
assign n_16708 =  x_935 & ~n_16689;
assign n_16709 =  i_29 &  n_16689;
assign n_16710 = ~n_16708 & ~n_16709;
assign n_16711 =  x_935 & ~n_16710;
assign n_16712 = ~x_935 &  n_16710;
assign n_16713 = ~n_16711 & ~n_16712;
assign n_16714 =  x_934 & ~n_16689;
assign n_16715 =  i_28 &  n_16689;
assign n_16716 = ~n_16714 & ~n_16715;
assign n_16717 =  x_934 & ~n_16716;
assign n_16718 = ~x_934 &  n_16716;
assign n_16719 = ~n_16717 & ~n_16718;
assign n_16720 =  x_933 & ~n_16689;
assign n_16721 =  i_27 &  n_16689;
assign n_16722 = ~n_16720 & ~n_16721;
assign n_16723 =  x_933 & ~n_16722;
assign n_16724 = ~x_933 &  n_16722;
assign n_16725 = ~n_16723 & ~n_16724;
assign n_16726 =  x_932 & ~n_16689;
assign n_16727 =  i_26 &  n_16689;
assign n_16728 = ~n_16726 & ~n_16727;
assign n_16729 =  x_932 & ~n_16728;
assign n_16730 = ~x_932 &  n_16728;
assign n_16731 = ~n_16729 & ~n_16730;
assign n_16732 =  x_931 & ~n_16689;
assign n_16733 =  i_25 &  n_16689;
assign n_16734 = ~n_16732 & ~n_16733;
assign n_16735 =  x_931 & ~n_16734;
assign n_16736 = ~x_931 &  n_16734;
assign n_16737 = ~n_16735 & ~n_16736;
assign n_16738 =  x_930 & ~n_16689;
assign n_16739 =  i_24 &  n_16689;
assign n_16740 = ~n_16738 & ~n_16739;
assign n_16741 =  x_930 & ~n_16740;
assign n_16742 = ~x_930 &  n_16740;
assign n_16743 = ~n_16741 & ~n_16742;
assign n_16744 =  x_929 & ~n_16689;
assign n_16745 =  i_23 &  n_16689;
assign n_16746 = ~n_16744 & ~n_16745;
assign n_16747 =  x_929 & ~n_16746;
assign n_16748 = ~x_929 &  n_16746;
assign n_16749 = ~n_16747 & ~n_16748;
assign n_16750 =  x_928 & ~n_16689;
assign n_16751 =  i_22 &  n_16689;
assign n_16752 = ~n_16750 & ~n_16751;
assign n_16753 =  x_928 & ~n_16752;
assign n_16754 = ~x_928 &  n_16752;
assign n_16755 = ~n_16753 & ~n_16754;
assign n_16756 =  x_927 & ~n_16689;
assign n_16757 =  i_21 &  n_16689;
assign n_16758 = ~n_16756 & ~n_16757;
assign n_16759 =  x_927 & ~n_16758;
assign n_16760 = ~x_927 &  n_16758;
assign n_16761 = ~n_16759 & ~n_16760;
assign n_16762 =  x_926 & ~n_16689;
assign n_16763 =  i_20 &  n_16689;
assign n_16764 = ~n_16762 & ~n_16763;
assign n_16765 =  x_926 & ~n_16764;
assign n_16766 = ~x_926 &  n_16764;
assign n_16767 = ~n_16765 & ~n_16766;
assign n_16768 =  x_925 & ~n_16689;
assign n_16769 =  i_19 &  n_16689;
assign n_16770 = ~n_16768 & ~n_16769;
assign n_16771 =  x_925 & ~n_16770;
assign n_16772 = ~x_925 &  n_16770;
assign n_16773 = ~n_16771 & ~n_16772;
assign n_16774 =  x_924 & ~n_16689;
assign n_16775 =  i_18 &  n_16689;
assign n_16776 = ~n_16774 & ~n_16775;
assign n_16777 =  x_924 & ~n_16776;
assign n_16778 = ~x_924 &  n_16776;
assign n_16779 = ~n_16777 & ~n_16778;
assign n_16780 =  x_923 & ~n_16689;
assign n_16781 =  i_17 &  n_16689;
assign n_16782 = ~n_16780 & ~n_16781;
assign n_16783 =  x_923 & ~n_16782;
assign n_16784 = ~x_923 &  n_16782;
assign n_16785 = ~n_16783 & ~n_16784;
assign n_16786 =  x_922 & ~n_16689;
assign n_16787 =  i_16 &  n_16689;
assign n_16788 = ~n_16786 & ~n_16787;
assign n_16789 =  x_922 & ~n_16788;
assign n_16790 = ~x_922 &  n_16788;
assign n_16791 = ~n_16789 & ~n_16790;
assign n_16792 =  x_921 & ~n_16689;
assign n_16793 =  i_15 &  n_16689;
assign n_16794 = ~n_16792 & ~n_16793;
assign n_16795 =  x_921 & ~n_16794;
assign n_16796 = ~x_921 &  n_16794;
assign n_16797 = ~n_16795 & ~n_16796;
assign n_16798 =  x_920 & ~n_16689;
assign n_16799 =  i_14 &  n_16689;
assign n_16800 = ~n_16798 & ~n_16799;
assign n_16801 =  x_920 & ~n_16800;
assign n_16802 = ~x_920 &  n_16800;
assign n_16803 = ~n_16801 & ~n_16802;
assign n_16804 =  x_919 & ~n_16689;
assign n_16805 =  i_13 &  n_16689;
assign n_16806 = ~n_16804 & ~n_16805;
assign n_16807 =  x_919 & ~n_16806;
assign n_16808 = ~x_919 &  n_16806;
assign n_16809 = ~n_16807 & ~n_16808;
assign n_16810 =  x_918 & ~n_16689;
assign n_16811 =  i_12 &  n_16689;
assign n_16812 = ~n_16810 & ~n_16811;
assign n_16813 =  x_918 & ~n_16812;
assign n_16814 = ~x_918 &  n_16812;
assign n_16815 = ~n_16813 & ~n_16814;
assign n_16816 =  x_917 & ~n_16689;
assign n_16817 =  i_11 &  n_16689;
assign n_16818 = ~n_16816 & ~n_16817;
assign n_16819 =  x_917 & ~n_16818;
assign n_16820 = ~x_917 &  n_16818;
assign n_16821 = ~n_16819 & ~n_16820;
assign n_16822 =  x_916 & ~n_16689;
assign n_16823 =  i_10 &  n_16689;
assign n_16824 = ~n_16822 & ~n_16823;
assign n_16825 =  x_916 & ~n_16824;
assign n_16826 = ~x_916 &  n_16824;
assign n_16827 = ~n_16825 & ~n_16826;
assign n_16828 =  x_915 & ~n_16689;
assign n_16829 =  i_9 &  n_16689;
assign n_16830 = ~n_16828 & ~n_16829;
assign n_16831 =  x_915 & ~n_16830;
assign n_16832 = ~x_915 &  n_16830;
assign n_16833 = ~n_16831 & ~n_16832;
assign n_16834 =  x_914 & ~n_16689;
assign n_16835 =  i_8 &  n_16689;
assign n_16836 = ~n_16834 & ~n_16835;
assign n_16837 =  x_914 & ~n_16836;
assign n_16838 = ~x_914 &  n_16836;
assign n_16839 = ~n_16837 & ~n_16838;
assign n_16840 =  x_913 & ~n_16689;
assign n_16841 =  i_7 &  n_16689;
assign n_16842 = ~n_16840 & ~n_16841;
assign n_16843 =  x_913 & ~n_16842;
assign n_16844 = ~x_913 &  n_16842;
assign n_16845 = ~n_16843 & ~n_16844;
assign n_16846 =  x_912 & ~n_16689;
assign n_16847 =  i_6 &  n_16689;
assign n_16848 = ~n_16846 & ~n_16847;
assign n_16849 =  x_912 & ~n_16848;
assign n_16850 = ~x_912 &  n_16848;
assign n_16851 = ~n_16849 & ~n_16850;
assign n_16852 =  x_911 & ~n_16689;
assign n_16853 =  i_5 &  n_16689;
assign n_16854 = ~n_16852 & ~n_16853;
assign n_16855 =  x_911 & ~n_16854;
assign n_16856 = ~x_911 &  n_16854;
assign n_16857 = ~n_16855 & ~n_16856;
assign n_16858 =  x_910 & ~n_16689;
assign n_16859 =  i_4 &  n_16689;
assign n_16860 = ~n_16858 & ~n_16859;
assign n_16861 =  x_910 & ~n_16860;
assign n_16862 = ~x_910 &  n_16860;
assign n_16863 = ~n_16861 & ~n_16862;
assign n_16864 =  x_909 & ~n_16689;
assign n_16865 =  i_3 &  n_16689;
assign n_16866 = ~n_16864 & ~n_16865;
assign n_16867 =  x_909 & ~n_16866;
assign n_16868 = ~x_909 &  n_16866;
assign n_16869 = ~n_16867 & ~n_16868;
assign n_16870 =  x_908 & ~n_16689;
assign n_16871 =  i_2 &  n_16689;
assign n_16872 = ~n_16870 & ~n_16871;
assign n_16873 =  x_908 & ~n_16872;
assign n_16874 = ~x_908 &  n_16872;
assign n_16875 = ~n_16873 & ~n_16874;
assign n_16876 =  x_907 & ~n_16689;
assign n_16877 =  i_1 &  n_16689;
assign n_16878 = ~n_16876 & ~n_16877;
assign n_16879 =  x_907 & ~n_16878;
assign n_16880 = ~x_907 &  n_16878;
assign n_16881 = ~n_16879 & ~n_16880;
assign n_16882 =  n_154 &  n_560;
assign n_16883 =  x_2969 &  n_16882;
assign n_16884 = ~n_9300 & ~n_16882;
assign n_16885 =  x_906 &  n_16884;
assign n_16886 = ~n_16883 & ~n_16885;
assign n_16887 =  x_906 & ~n_16886;
assign n_16888 = ~x_906 &  n_16886;
assign n_16889 = ~n_16887 & ~n_16888;
assign n_16890 =  x_2968 &  n_16882;
assign n_16891 =  x_905 &  n_16884;
assign n_16892 = ~n_16890 & ~n_16891;
assign n_16893 =  x_905 & ~n_16892;
assign n_16894 = ~x_905 &  n_16892;
assign n_16895 = ~n_16893 & ~n_16894;
assign n_16896 =  x_2967 &  n_16882;
assign n_16897 =  x_904 &  n_16884;
assign n_16898 = ~n_16896 & ~n_16897;
assign n_16899 =  x_904 & ~n_16898;
assign n_16900 = ~x_904 &  n_16898;
assign n_16901 = ~n_16899 & ~n_16900;
assign n_16902 =  x_2966 &  n_16882;
assign n_16903 =  x_903 &  n_16884;
assign n_16904 = ~n_16902 & ~n_16903;
assign n_16905 =  x_903 & ~n_16904;
assign n_16906 = ~x_903 &  n_16904;
assign n_16907 = ~n_16905 & ~n_16906;
assign n_16908 =  x_2965 &  n_16882;
assign n_16909 =  x_902 &  n_16884;
assign n_16910 = ~n_16908 & ~n_16909;
assign n_16911 =  x_902 & ~n_16910;
assign n_16912 = ~x_902 &  n_16910;
assign n_16913 = ~n_16911 & ~n_16912;
assign n_16914 =  x_2964 &  n_16882;
assign n_16915 =  x_901 &  n_16884;
assign n_16916 = ~n_16914 & ~n_16915;
assign n_16917 =  x_901 & ~n_16916;
assign n_16918 = ~x_901 &  n_16916;
assign n_16919 = ~n_16917 & ~n_16918;
assign n_16920 =  x_2963 &  n_16882;
assign n_16921 =  x_900 &  n_16884;
assign n_16922 = ~n_16920 & ~n_16921;
assign n_16923 =  x_900 & ~n_16922;
assign n_16924 = ~x_900 &  n_16922;
assign n_16925 = ~n_16923 & ~n_16924;
assign n_16926 =  x_2962 &  n_16882;
assign n_16927 =  x_899 &  n_16884;
assign n_16928 = ~n_16926 & ~n_16927;
assign n_16929 =  x_899 & ~n_16928;
assign n_16930 = ~x_899 &  n_16928;
assign n_16931 = ~n_16929 & ~n_16930;
assign n_16932 =  x_2961 &  n_16882;
assign n_16933 =  x_898 &  n_16884;
assign n_16934 = ~n_16932 & ~n_16933;
assign n_16935 =  x_898 & ~n_16934;
assign n_16936 = ~x_898 &  n_16934;
assign n_16937 = ~n_16935 & ~n_16936;
assign n_16938 =  x_2960 &  n_16882;
assign n_16939 =  x_897 &  n_16884;
assign n_16940 = ~n_16938 & ~n_16939;
assign n_16941 =  x_897 & ~n_16940;
assign n_16942 = ~x_897 &  n_16940;
assign n_16943 = ~n_16941 & ~n_16942;
assign n_16944 =  x_2959 &  n_16882;
assign n_16945 =  x_896 &  n_16884;
assign n_16946 = ~n_16944 & ~n_16945;
assign n_16947 =  x_896 & ~n_16946;
assign n_16948 = ~x_896 &  n_16946;
assign n_16949 = ~n_16947 & ~n_16948;
assign n_16950 =  x_2958 &  n_16882;
assign n_16951 =  x_895 &  n_16884;
assign n_16952 = ~n_16950 & ~n_16951;
assign n_16953 =  x_895 & ~n_16952;
assign n_16954 = ~x_895 &  n_16952;
assign n_16955 = ~n_16953 & ~n_16954;
assign n_16956 =  x_2957 &  n_16882;
assign n_16957 =  x_894 &  n_16884;
assign n_16958 = ~n_16956 & ~n_16957;
assign n_16959 =  x_894 & ~n_16958;
assign n_16960 = ~x_894 &  n_16958;
assign n_16961 = ~n_16959 & ~n_16960;
assign n_16962 =  x_2956 &  n_16882;
assign n_16963 =  x_893 &  n_16884;
assign n_16964 = ~n_16962 & ~n_16963;
assign n_16965 =  x_893 & ~n_16964;
assign n_16966 = ~x_893 &  n_16964;
assign n_16967 = ~n_16965 & ~n_16966;
assign n_16968 =  x_2955 &  n_16882;
assign n_16969 =  x_892 &  n_16884;
assign n_16970 = ~n_16968 & ~n_16969;
assign n_16971 =  x_892 & ~n_16970;
assign n_16972 = ~x_892 &  n_16970;
assign n_16973 = ~n_16971 & ~n_16972;
assign n_16974 =  x_2954 &  n_16882;
assign n_16975 =  x_891 &  n_16884;
assign n_16976 = ~n_16974 & ~n_16975;
assign n_16977 =  x_891 & ~n_16976;
assign n_16978 = ~x_891 &  n_16976;
assign n_16979 = ~n_16977 & ~n_16978;
assign n_16980 =  x_2953 &  n_16882;
assign n_16981 =  x_890 &  n_16884;
assign n_16982 = ~n_16980 & ~n_16981;
assign n_16983 =  x_890 & ~n_16982;
assign n_16984 = ~x_890 &  n_16982;
assign n_16985 = ~n_16983 & ~n_16984;
assign n_16986 =  x_2952 &  n_16882;
assign n_16987 =  x_889 &  n_16884;
assign n_16988 = ~n_16986 & ~n_16987;
assign n_16989 =  x_889 & ~n_16988;
assign n_16990 = ~x_889 &  n_16988;
assign n_16991 = ~n_16989 & ~n_16990;
assign n_16992 =  x_2951 &  n_16882;
assign n_16993 =  x_888 &  n_16884;
assign n_16994 = ~n_16992 & ~n_16993;
assign n_16995 =  x_888 & ~n_16994;
assign n_16996 = ~x_888 &  n_16994;
assign n_16997 = ~n_16995 & ~n_16996;
assign n_16998 =  x_2950 &  n_16882;
assign n_16999 =  x_887 &  n_16884;
assign n_17000 = ~n_16998 & ~n_16999;
assign n_17001 =  x_887 & ~n_17000;
assign n_17002 = ~x_887 &  n_17000;
assign n_17003 = ~n_17001 & ~n_17002;
assign n_17004 =  x_2949 &  n_16882;
assign n_17005 =  x_886 &  n_16884;
assign n_17006 = ~n_17004 & ~n_17005;
assign n_17007 =  x_886 & ~n_17006;
assign n_17008 = ~x_886 &  n_17006;
assign n_17009 = ~n_17007 & ~n_17008;
assign n_17010 =  x_2948 &  n_16882;
assign n_17011 =  x_885 &  n_16884;
assign n_17012 = ~n_17010 & ~n_17011;
assign n_17013 =  x_885 & ~n_17012;
assign n_17014 = ~x_885 &  n_17012;
assign n_17015 = ~n_17013 & ~n_17014;
assign n_17016 =  x_2947 &  n_16882;
assign n_17017 =  x_884 &  n_16884;
assign n_17018 = ~n_17016 & ~n_17017;
assign n_17019 =  x_884 & ~n_17018;
assign n_17020 = ~x_884 &  n_17018;
assign n_17021 = ~n_17019 & ~n_17020;
assign n_17022 =  x_2946 &  n_16882;
assign n_17023 =  x_883 &  n_16884;
assign n_17024 = ~n_17022 & ~n_17023;
assign n_17025 =  x_883 & ~n_17024;
assign n_17026 = ~x_883 &  n_17024;
assign n_17027 = ~n_17025 & ~n_17026;
assign n_17028 =  x_2945 &  n_16882;
assign n_17029 =  x_882 &  n_16884;
assign n_17030 = ~n_17028 & ~n_17029;
assign n_17031 =  x_882 & ~n_17030;
assign n_17032 = ~x_882 &  n_17030;
assign n_17033 = ~n_17031 & ~n_17032;
assign n_17034 =  x_2944 &  n_16882;
assign n_17035 =  x_881 &  n_16884;
assign n_17036 = ~n_17034 & ~n_17035;
assign n_17037 =  x_881 & ~n_17036;
assign n_17038 = ~x_881 &  n_17036;
assign n_17039 = ~n_17037 & ~n_17038;
assign n_17040 =  x_2943 &  n_16882;
assign n_17041 =  x_880 &  n_16884;
assign n_17042 = ~n_17040 & ~n_17041;
assign n_17043 =  x_880 & ~n_17042;
assign n_17044 = ~x_880 &  n_17042;
assign n_17045 = ~n_17043 & ~n_17044;
assign n_17046 =  x_2942 &  n_16882;
assign n_17047 =  x_879 &  n_16884;
assign n_17048 = ~n_17046 & ~n_17047;
assign n_17049 =  x_879 & ~n_17048;
assign n_17050 = ~x_879 &  n_17048;
assign n_17051 = ~n_17049 & ~n_17050;
assign n_17052 =  x_2941 &  n_16882;
assign n_17053 =  x_878 &  n_16884;
assign n_17054 = ~n_17052 & ~n_17053;
assign n_17055 =  x_878 & ~n_17054;
assign n_17056 = ~x_878 &  n_17054;
assign n_17057 = ~n_17055 & ~n_17056;
assign n_17058 =  x_2940 &  n_16882;
assign n_17059 =  x_877 &  n_16884;
assign n_17060 = ~n_17058 & ~n_17059;
assign n_17061 =  x_877 & ~n_17060;
assign n_17062 = ~x_877 &  n_17060;
assign n_17063 = ~n_17061 & ~n_17062;
assign n_17064 =  x_2939 &  n_16882;
assign n_17065 =  x_876 &  n_16884;
assign n_17066 = ~n_17064 & ~n_17065;
assign n_17067 =  x_876 & ~n_17066;
assign n_17068 = ~x_876 &  n_17066;
assign n_17069 = ~n_17067 & ~n_17068;
assign n_17070 =  x_2938 &  n_16882;
assign n_17071 =  x_875 &  n_16884;
assign n_17072 = ~n_17070 & ~n_17071;
assign n_17073 =  x_875 & ~n_17072;
assign n_17074 = ~x_875 &  n_17072;
assign n_17075 = ~n_17073 & ~n_17074;
assign n_17076 =  n_349 &  n_8347;
assign n_17077 =  n_3628 &  n_17076;
assign n_17078 =  x_843 & ~n_17077;
assign n_17079 =  x_843 &  n_17078;
assign n_17080 = ~x_843 & ~n_17078;
assign n_17081 = ~n_17079 & ~n_17080;
assign n_17082 =  x_842 & ~n_17077;
assign n_17083 =  x_842 &  n_17082;
assign n_17084 = ~x_842 & ~n_17082;
assign n_17085 = ~n_17083 & ~n_17084;
assign n_17086 =  x_841 & ~n_17077;
assign n_17087 =  x_841 &  n_17086;
assign n_17088 = ~x_841 & ~n_17086;
assign n_17089 = ~n_17087 & ~n_17088;
assign n_17090 =  x_840 & ~n_17077;
assign n_17091 =  x_840 &  n_17090;
assign n_17092 = ~x_840 & ~n_17090;
assign n_17093 = ~n_17091 & ~n_17092;
assign n_17094 =  x_839 & ~n_17077;
assign n_17095 =  x_839 &  n_17094;
assign n_17096 = ~x_839 & ~n_17094;
assign n_17097 = ~n_17095 & ~n_17096;
assign n_17098 =  x_838 & ~n_17077;
assign n_17099 =  x_838 &  n_17098;
assign n_17100 = ~x_838 & ~n_17098;
assign n_17101 = ~n_17099 & ~n_17100;
assign n_17102 =  x_837 & ~n_17077;
assign n_17103 =  x_837 &  n_17102;
assign n_17104 = ~x_837 & ~n_17102;
assign n_17105 = ~n_17103 & ~n_17104;
assign n_17106 =  x_836 & ~n_17077;
assign n_17107 =  x_836 &  n_17106;
assign n_17108 = ~x_836 & ~n_17106;
assign n_17109 = ~n_17107 & ~n_17108;
assign n_17110 =  x_835 & ~n_17077;
assign n_17111 =  x_835 &  n_17110;
assign n_17112 = ~x_835 & ~n_17110;
assign n_17113 = ~n_17111 & ~n_17112;
assign n_17114 =  x_834 & ~n_17077;
assign n_17115 =  x_834 &  n_17114;
assign n_17116 = ~x_834 & ~n_17114;
assign n_17117 = ~n_17115 & ~n_17116;
assign n_17118 =  x_833 & ~n_17077;
assign n_17119 =  x_833 &  n_17118;
assign n_17120 = ~x_833 & ~n_17118;
assign n_17121 = ~n_17119 & ~n_17120;
assign n_17122 =  x_832 & ~n_17077;
assign n_17123 =  x_832 &  n_17122;
assign n_17124 = ~x_832 & ~n_17122;
assign n_17125 = ~n_17123 & ~n_17124;
assign n_17126 =  x_831 & ~n_17077;
assign n_17127 =  x_831 &  n_17126;
assign n_17128 = ~x_831 & ~n_17126;
assign n_17129 = ~n_17127 & ~n_17128;
assign n_17130 =  x_830 & ~n_17077;
assign n_17131 =  x_830 &  n_17130;
assign n_17132 = ~x_830 & ~n_17130;
assign n_17133 = ~n_17131 & ~n_17132;
assign n_17134 =  x_829 & ~n_17077;
assign n_17135 =  x_829 &  n_17134;
assign n_17136 = ~x_829 & ~n_17134;
assign n_17137 = ~n_17135 & ~n_17136;
assign n_17138 =  x_828 & ~n_17077;
assign n_17139 =  x_828 &  n_17138;
assign n_17140 = ~x_828 & ~n_17138;
assign n_17141 = ~n_17139 & ~n_17140;
assign n_17142 =  x_827 & ~n_17077;
assign n_17143 =  x_827 &  n_17142;
assign n_17144 = ~x_827 & ~n_17142;
assign n_17145 = ~n_17143 & ~n_17144;
assign n_17146 =  x_826 & ~n_17077;
assign n_17147 =  x_826 &  n_17146;
assign n_17148 = ~x_826 & ~n_17146;
assign n_17149 = ~n_17147 & ~n_17148;
assign n_17150 =  x_825 & ~n_17077;
assign n_17151 =  x_825 &  n_17150;
assign n_17152 = ~x_825 & ~n_17150;
assign n_17153 = ~n_17151 & ~n_17152;
assign n_17154 =  x_824 & ~n_17077;
assign n_17155 =  x_824 &  n_17154;
assign n_17156 = ~x_824 & ~n_17154;
assign n_17157 = ~n_17155 & ~n_17156;
assign n_17158 =  x_823 & ~n_17077;
assign n_17159 =  x_823 &  n_17158;
assign n_17160 = ~x_823 & ~n_17158;
assign n_17161 = ~n_17159 & ~n_17160;
assign n_17162 =  x_822 & ~n_17077;
assign n_17163 =  x_822 &  n_17162;
assign n_17164 = ~x_822 & ~n_17162;
assign n_17165 = ~n_17163 & ~n_17164;
assign n_17166 =  x_821 & ~n_17077;
assign n_17167 =  x_821 &  n_17166;
assign n_17168 = ~x_821 & ~n_17166;
assign n_17169 = ~n_17167 & ~n_17168;
assign n_17170 =  x_820 & ~n_17077;
assign n_17171 =  x_820 &  n_17170;
assign n_17172 = ~x_820 & ~n_17170;
assign n_17173 = ~n_17171 & ~n_17172;
assign n_17174 =  x_819 & ~n_17077;
assign n_17175 =  x_819 &  n_17174;
assign n_17176 = ~x_819 & ~n_17174;
assign n_17177 = ~n_17175 & ~n_17176;
assign n_17178 =  x_818 & ~n_17077;
assign n_17179 =  x_818 &  n_17178;
assign n_17180 = ~x_818 & ~n_17178;
assign n_17181 = ~n_17179 & ~n_17180;
assign n_17182 =  x_817 & ~n_17077;
assign n_17183 =  x_817 &  n_17182;
assign n_17184 = ~x_817 & ~n_17182;
assign n_17185 = ~n_17183 & ~n_17184;
assign n_17186 =  x_816 & ~n_17077;
assign n_17187 =  x_816 &  n_17186;
assign n_17188 = ~x_816 & ~n_17186;
assign n_17189 = ~n_17187 & ~n_17188;
assign n_17190 =  x_815 & ~n_17077;
assign n_17191 =  x_815 &  n_17190;
assign n_17192 = ~x_815 & ~n_17190;
assign n_17193 = ~n_17191 & ~n_17192;
assign n_17194 =  x_814 & ~n_17077;
assign n_17195 =  x_814 &  n_17194;
assign n_17196 = ~x_814 & ~n_17194;
assign n_17197 = ~n_17195 & ~n_17196;
assign n_17198 =  x_813 & ~n_17077;
assign n_17199 =  x_813 &  n_17198;
assign n_17200 = ~x_813 & ~n_17198;
assign n_17201 = ~n_17199 & ~n_17200;
assign n_17202 =  x_812 & ~n_17077;
assign n_17203 =  x_812 &  n_17202;
assign n_17204 = ~x_812 & ~n_17202;
assign n_17205 = ~n_17203 & ~n_17204;
assign n_17206 = ~x_3248 &  x_3249;
assign n_17207 =  x_3250 &  n_17206;
assign n_17208 = ~x_3244 &  x_3245;
assign n_17209 = ~x_3246 &  x_3247;
assign n_17210 =  n_17208 &  n_17209;
assign n_17211 = ~x_3240 & ~x_3241;
assign n_17212 = ~x_3242 & ~x_3243;
assign n_17213 =  n_17211 &  n_17212;
assign n_17214 =  n_17210 &  n_17213;
assign n_17215 =  n_17207 &  n_17214;
assign n_17216 = ~x_3228 & ~x_3229;
assign n_17217 = ~x_3230 & ~x_3231;
assign n_17218 =  n_17216 &  n_17217;
assign n_17219 = ~x_3224 & ~x_3225;
assign n_17220 = ~x_3226 & ~x_3227;
assign n_17221 =  n_17219 &  n_17220;
assign n_17222 =  n_17218 &  n_17221;
assign n_17223 = ~x_3236 & ~x_3237;
assign n_17224 = ~x_3238 & ~x_3239;
assign n_17225 =  n_17223 &  n_17224;
assign n_17226 = ~x_3232 & ~x_3233;
assign n_17227 = ~x_3234 & ~x_3235;
assign n_17228 =  n_17226 &  n_17227;
assign n_17229 =  n_17225 &  n_17228;
assign n_17230 =  n_17222 &  n_17229;
assign n_17231 =  n_17215 &  n_17230;
assign n_17232 =  x_3251 & ~x_3252;
assign n_17233 = ~x_3253 & ~x_3254;
assign n_17234 =  n_17232 &  n_17233;
assign n_17235 =  n_17231 &  n_17234;
assign n_17236 = ~x_2842 & ~x_3255;
assign n_17237 = ~x_2906 &  x_3255;
assign n_17238 = ~n_17236 & ~n_17237;
assign n_17239 =  n_17235 &  n_17238;
assign n_17240 = ~x_3251 &  n_8081;
assign n_17241 =  n_17231 &  n_17240;
assign n_17242 = ~x_3064 &  n_17241;
assign n_17243 = ~i_32 & ~n_17241;
assign n_17244 = ~n_17235 & ~n_17243;
assign n_17245 = ~n_17242 &  n_17244;
assign n_17246 = ~n_17239 & ~n_17245;
assign n_17247 =  n_8055 & ~n_17246;
assign n_17248 =  x_2842 &  n_761;
assign n_17249 =  x_811 & ~n_8051;
assign n_17250 = ~n_17248 & ~n_17249;
assign n_17251 = ~n_17247 &  n_17250;
assign n_17252 =  x_811 & ~n_17251;
assign n_17253 = ~x_811 &  n_17251;
assign n_17254 = ~n_17252 & ~n_17253;
assign n_17255 = ~x_2841 & ~x_3255;
assign n_17256 = ~x_2905 &  x_3255;
assign n_17257 = ~n_17255 & ~n_17256;
assign n_17258 =  n_17235 &  n_17257;
assign n_17259 = ~x_3063 &  n_17241;
assign n_17260 = ~i_31 & ~n_17241;
assign n_17261 = ~n_17235 & ~n_17260;
assign n_17262 = ~n_17259 &  n_17261;
assign n_17263 = ~n_17258 & ~n_17262;
assign n_17264 =  n_8055 & ~n_17263;
assign n_17265 =  x_2841 &  n_761;
assign n_17266 =  x_810 & ~n_8051;
assign n_17267 = ~n_17265 & ~n_17266;
assign n_17268 = ~n_17264 &  n_17267;
assign n_17269 =  x_810 & ~n_17268;
assign n_17270 = ~x_810 &  n_17268;
assign n_17271 = ~n_17269 & ~n_17270;
assign n_17272 = ~x_2840 & ~x_3255;
assign n_17273 = ~x_2904 &  x_3255;
assign n_17274 = ~n_17272 & ~n_17273;
assign n_17275 =  n_17235 &  n_17274;
assign n_17276 = ~x_3062 &  n_17241;
assign n_17277 = ~i_30 & ~n_17241;
assign n_17278 = ~n_17235 & ~n_17277;
assign n_17279 = ~n_17276 &  n_17278;
assign n_17280 = ~n_17275 & ~n_17279;
assign n_17281 =  n_8055 & ~n_17280;
assign n_17282 =  x_2840 &  n_761;
assign n_17283 =  x_809 & ~n_8051;
assign n_17284 = ~n_17282 & ~n_17283;
assign n_17285 = ~n_17281 &  n_17284;
assign n_17286 =  x_809 & ~n_17285;
assign n_17287 = ~x_809 &  n_17285;
assign n_17288 = ~n_17286 & ~n_17287;
assign n_17289 = ~x_2839 & ~x_3255;
assign n_17290 = ~x_2903 &  x_3255;
assign n_17291 = ~n_17289 & ~n_17290;
assign n_17292 =  n_17235 &  n_17291;
assign n_17293 = ~x_3061 &  n_17241;
assign n_17294 = ~i_29 & ~n_17241;
assign n_17295 = ~n_17235 & ~n_17294;
assign n_17296 = ~n_17293 &  n_17295;
assign n_17297 = ~n_17292 & ~n_17296;
assign n_17298 =  n_8055 & ~n_17297;
assign n_17299 =  x_2839 &  n_761;
assign n_17300 =  x_808 & ~n_8051;
assign n_17301 = ~n_17299 & ~n_17300;
assign n_17302 = ~n_17298 &  n_17301;
assign n_17303 =  x_808 & ~n_17302;
assign n_17304 = ~x_808 &  n_17302;
assign n_17305 = ~n_17303 & ~n_17304;
assign n_17306 = ~x_2838 & ~x_3255;
assign n_17307 = ~x_2902 &  x_3255;
assign n_17308 = ~n_17306 & ~n_17307;
assign n_17309 =  n_17235 &  n_17308;
assign n_17310 = ~x_3060 &  n_17241;
assign n_17311 = ~i_28 & ~n_17241;
assign n_17312 = ~n_17235 & ~n_17311;
assign n_17313 = ~n_17310 &  n_17312;
assign n_17314 = ~n_17309 & ~n_17313;
assign n_17315 =  n_8055 & ~n_17314;
assign n_17316 =  x_2838 &  n_761;
assign n_17317 =  x_807 & ~n_8051;
assign n_17318 = ~n_17316 & ~n_17317;
assign n_17319 = ~n_17315 &  n_17318;
assign n_17320 =  x_807 & ~n_17319;
assign n_17321 = ~x_807 &  n_17319;
assign n_17322 = ~n_17320 & ~n_17321;
assign n_17323 = ~x_2837 & ~x_3255;
assign n_17324 = ~x_2901 &  x_3255;
assign n_17325 = ~n_17323 & ~n_17324;
assign n_17326 =  n_17235 &  n_17325;
assign n_17327 = ~x_3059 &  n_17241;
assign n_17328 = ~i_27 & ~n_17241;
assign n_17329 = ~n_17235 & ~n_17328;
assign n_17330 = ~n_17327 &  n_17329;
assign n_17331 = ~n_17326 & ~n_17330;
assign n_17332 =  n_8055 & ~n_17331;
assign n_17333 =  x_2837 &  n_761;
assign n_17334 =  x_806 & ~n_8051;
assign n_17335 = ~n_17333 & ~n_17334;
assign n_17336 = ~n_17332 &  n_17335;
assign n_17337 =  x_806 & ~n_17336;
assign n_17338 = ~x_806 &  n_17336;
assign n_17339 = ~n_17337 & ~n_17338;
assign n_17340 = ~x_2836 & ~x_3255;
assign n_17341 = ~x_2900 &  x_3255;
assign n_17342 = ~n_17340 & ~n_17341;
assign n_17343 =  n_17235 &  n_17342;
assign n_17344 = ~x_3058 &  n_17241;
assign n_17345 = ~i_26 & ~n_17241;
assign n_17346 = ~n_17235 & ~n_17345;
assign n_17347 = ~n_17344 &  n_17346;
assign n_17348 = ~n_17343 & ~n_17347;
assign n_17349 =  n_8055 & ~n_17348;
assign n_17350 =  x_2836 &  n_761;
assign n_17351 =  x_805 & ~n_8051;
assign n_17352 = ~n_17350 & ~n_17351;
assign n_17353 = ~n_17349 &  n_17352;
assign n_17354 =  x_805 & ~n_17353;
assign n_17355 = ~x_805 &  n_17353;
assign n_17356 = ~n_17354 & ~n_17355;
assign n_17357 = ~x_2835 & ~x_3255;
assign n_17358 = ~x_2899 &  x_3255;
assign n_17359 = ~n_17357 & ~n_17358;
assign n_17360 =  n_17235 &  n_17359;
assign n_17361 = ~x_3057 &  n_17241;
assign n_17362 = ~i_25 & ~n_17241;
assign n_17363 = ~n_17235 & ~n_17362;
assign n_17364 = ~n_17361 &  n_17363;
assign n_17365 = ~n_17360 & ~n_17364;
assign n_17366 =  n_8055 & ~n_17365;
assign n_17367 =  x_2835 &  n_761;
assign n_17368 =  x_804 & ~n_8051;
assign n_17369 = ~n_17367 & ~n_17368;
assign n_17370 = ~n_17366 &  n_17369;
assign n_17371 =  x_804 & ~n_17370;
assign n_17372 = ~x_804 &  n_17370;
assign n_17373 = ~n_17371 & ~n_17372;
assign n_17374 = ~x_2834 & ~x_3255;
assign n_17375 = ~x_2898 &  x_3255;
assign n_17376 = ~n_17374 & ~n_17375;
assign n_17377 =  n_17235 &  n_17376;
assign n_17378 = ~x_3056 &  n_17241;
assign n_17379 = ~i_24 & ~n_17241;
assign n_17380 = ~n_17235 & ~n_17379;
assign n_17381 = ~n_17378 &  n_17380;
assign n_17382 = ~n_17377 & ~n_17381;
assign n_17383 =  n_8055 & ~n_17382;
assign n_17384 =  x_2834 &  n_761;
assign n_17385 =  x_803 & ~n_8051;
assign n_17386 = ~n_17384 & ~n_17385;
assign n_17387 = ~n_17383 &  n_17386;
assign n_17388 =  x_803 & ~n_17387;
assign n_17389 = ~x_803 &  n_17387;
assign n_17390 = ~n_17388 & ~n_17389;
assign n_17391 = ~x_2833 & ~x_3255;
assign n_17392 = ~x_2897 &  x_3255;
assign n_17393 = ~n_17391 & ~n_17392;
assign n_17394 =  n_17235 &  n_17393;
assign n_17395 = ~x_3055 &  n_17241;
assign n_17396 = ~i_23 & ~n_17241;
assign n_17397 = ~n_17235 & ~n_17396;
assign n_17398 = ~n_17395 &  n_17397;
assign n_17399 = ~n_17394 & ~n_17398;
assign n_17400 =  n_8055 & ~n_17399;
assign n_17401 =  x_2833 &  n_761;
assign n_17402 =  x_802 & ~n_8051;
assign n_17403 = ~n_17401 & ~n_17402;
assign n_17404 = ~n_17400 &  n_17403;
assign n_17405 =  x_802 & ~n_17404;
assign n_17406 = ~x_802 &  n_17404;
assign n_17407 = ~n_17405 & ~n_17406;
assign n_17408 = ~x_2832 & ~x_3255;
assign n_17409 = ~x_2896 &  x_3255;
assign n_17410 = ~n_17408 & ~n_17409;
assign n_17411 =  n_17235 &  n_17410;
assign n_17412 = ~x_3054 &  n_17241;
assign n_17413 = ~i_22 & ~n_17241;
assign n_17414 = ~n_17235 & ~n_17413;
assign n_17415 = ~n_17412 &  n_17414;
assign n_17416 = ~n_17411 & ~n_17415;
assign n_17417 =  n_8055 & ~n_17416;
assign n_17418 =  x_2832 &  n_761;
assign n_17419 =  x_801 & ~n_8051;
assign n_17420 = ~n_17418 & ~n_17419;
assign n_17421 = ~n_17417 &  n_17420;
assign n_17422 =  x_801 & ~n_17421;
assign n_17423 = ~x_801 &  n_17421;
assign n_17424 = ~n_17422 & ~n_17423;
assign n_17425 = ~x_2831 & ~x_3255;
assign n_17426 = ~x_2895 &  x_3255;
assign n_17427 = ~n_17425 & ~n_17426;
assign n_17428 =  n_17235 &  n_17427;
assign n_17429 = ~x_3053 &  n_17241;
assign n_17430 = ~i_21 & ~n_17241;
assign n_17431 = ~n_17235 & ~n_17430;
assign n_17432 = ~n_17429 &  n_17431;
assign n_17433 = ~n_17428 & ~n_17432;
assign n_17434 =  n_8055 & ~n_17433;
assign n_17435 =  x_2831 &  n_761;
assign n_17436 =  x_800 & ~n_8051;
assign n_17437 = ~n_17435 & ~n_17436;
assign n_17438 = ~n_17434 &  n_17437;
assign n_17439 =  x_800 & ~n_17438;
assign n_17440 = ~x_800 &  n_17438;
assign n_17441 = ~n_17439 & ~n_17440;
assign n_17442 = ~x_2830 & ~x_3255;
assign n_17443 = ~x_2894 &  x_3255;
assign n_17444 = ~n_17442 & ~n_17443;
assign n_17445 =  n_17235 &  n_17444;
assign n_17446 = ~x_3052 &  n_17241;
assign n_17447 = ~i_20 & ~n_17241;
assign n_17448 = ~n_17235 & ~n_17447;
assign n_17449 = ~n_17446 &  n_17448;
assign n_17450 = ~n_17445 & ~n_17449;
assign n_17451 =  n_8055 & ~n_17450;
assign n_17452 =  x_2830 &  n_761;
assign n_17453 =  x_799 & ~n_8051;
assign n_17454 = ~n_17452 & ~n_17453;
assign n_17455 = ~n_17451 &  n_17454;
assign n_17456 =  x_799 & ~n_17455;
assign n_17457 = ~x_799 &  n_17455;
assign n_17458 = ~n_17456 & ~n_17457;
assign n_17459 = ~x_2829 & ~x_3255;
assign n_17460 = ~x_2893 &  x_3255;
assign n_17461 = ~n_17459 & ~n_17460;
assign n_17462 =  n_17235 &  n_17461;
assign n_17463 = ~x_3051 &  n_17241;
assign n_17464 = ~i_19 & ~n_17241;
assign n_17465 = ~n_17235 & ~n_17464;
assign n_17466 = ~n_17463 &  n_17465;
assign n_17467 = ~n_17462 & ~n_17466;
assign n_17468 =  n_8055 & ~n_17467;
assign n_17469 =  x_2829 &  n_761;
assign n_17470 =  x_798 & ~n_8051;
assign n_17471 = ~n_17469 & ~n_17470;
assign n_17472 = ~n_17468 &  n_17471;
assign n_17473 =  x_798 & ~n_17472;
assign n_17474 = ~x_798 &  n_17472;
assign n_17475 = ~n_17473 & ~n_17474;
assign n_17476 = ~x_2828 & ~x_3255;
assign n_17477 = ~x_2892 &  x_3255;
assign n_17478 = ~n_17476 & ~n_17477;
assign n_17479 =  n_17235 &  n_17478;
assign n_17480 = ~x_3050 &  n_17241;
assign n_17481 = ~i_18 & ~n_17241;
assign n_17482 = ~n_17235 & ~n_17481;
assign n_17483 = ~n_17480 &  n_17482;
assign n_17484 = ~n_17479 & ~n_17483;
assign n_17485 =  n_8055 & ~n_17484;
assign n_17486 =  x_2828 &  n_761;
assign n_17487 =  x_797 & ~n_8051;
assign n_17488 = ~n_17486 & ~n_17487;
assign n_17489 = ~n_17485 &  n_17488;
assign n_17490 =  x_797 & ~n_17489;
assign n_17491 = ~x_797 &  n_17489;
assign n_17492 = ~n_17490 & ~n_17491;
assign n_17493 = ~x_2827 & ~x_3255;
assign n_17494 = ~x_2891 &  x_3255;
assign n_17495 = ~n_17493 & ~n_17494;
assign n_17496 =  n_17235 &  n_17495;
assign n_17497 = ~x_3049 &  n_17241;
assign n_17498 = ~i_17 & ~n_17241;
assign n_17499 = ~n_17235 & ~n_17498;
assign n_17500 = ~n_17497 &  n_17499;
assign n_17501 = ~n_17496 & ~n_17500;
assign n_17502 =  n_8055 & ~n_17501;
assign n_17503 =  x_2827 &  n_761;
assign n_17504 =  x_796 & ~n_8051;
assign n_17505 = ~n_17503 & ~n_17504;
assign n_17506 = ~n_17502 &  n_17505;
assign n_17507 =  x_796 & ~n_17506;
assign n_17508 = ~x_796 &  n_17506;
assign n_17509 = ~n_17507 & ~n_17508;
assign n_17510 = ~x_2826 & ~x_3255;
assign n_17511 = ~x_2890 &  x_3255;
assign n_17512 = ~n_17510 & ~n_17511;
assign n_17513 =  n_17235 &  n_17512;
assign n_17514 = ~x_3048 &  n_17241;
assign n_17515 = ~i_16 & ~n_17241;
assign n_17516 = ~n_17235 & ~n_17515;
assign n_17517 = ~n_17514 &  n_17516;
assign n_17518 = ~n_17513 & ~n_17517;
assign n_17519 =  n_8055 & ~n_17518;
assign n_17520 =  x_2826 &  n_761;
assign n_17521 =  x_795 & ~n_8051;
assign n_17522 = ~n_17520 & ~n_17521;
assign n_17523 = ~n_17519 &  n_17522;
assign n_17524 =  x_795 & ~n_17523;
assign n_17525 = ~x_795 &  n_17523;
assign n_17526 = ~n_17524 & ~n_17525;
assign n_17527 = ~x_2825 & ~x_3255;
assign n_17528 = ~x_2889 &  x_3255;
assign n_17529 = ~n_17527 & ~n_17528;
assign n_17530 =  n_17235 &  n_17529;
assign n_17531 = ~x_3047 &  n_17241;
assign n_17532 = ~i_15 & ~n_17241;
assign n_17533 = ~n_17235 & ~n_17532;
assign n_17534 = ~n_17531 &  n_17533;
assign n_17535 = ~n_17530 & ~n_17534;
assign n_17536 =  n_8055 & ~n_17535;
assign n_17537 =  x_2825 &  n_761;
assign n_17538 =  x_794 & ~n_8051;
assign n_17539 = ~n_17537 & ~n_17538;
assign n_17540 = ~n_17536 &  n_17539;
assign n_17541 =  x_794 & ~n_17540;
assign n_17542 = ~x_794 &  n_17540;
assign n_17543 = ~n_17541 & ~n_17542;
assign n_17544 = ~x_2824 & ~x_3255;
assign n_17545 = ~x_2888 &  x_3255;
assign n_17546 = ~n_17544 & ~n_17545;
assign n_17547 =  n_17235 &  n_17546;
assign n_17548 = ~x_3046 &  n_17241;
assign n_17549 = ~i_14 & ~n_17241;
assign n_17550 = ~n_17235 & ~n_17549;
assign n_17551 = ~n_17548 &  n_17550;
assign n_17552 = ~n_17547 & ~n_17551;
assign n_17553 =  n_8055 & ~n_17552;
assign n_17554 =  x_2824 &  n_761;
assign n_17555 =  x_793 & ~n_8051;
assign n_17556 = ~n_17554 & ~n_17555;
assign n_17557 = ~n_17553 &  n_17556;
assign n_17558 =  x_793 & ~n_17557;
assign n_17559 = ~x_793 &  n_17557;
assign n_17560 = ~n_17558 & ~n_17559;
assign n_17561 = ~x_2823 & ~x_3255;
assign n_17562 = ~x_2887 &  x_3255;
assign n_17563 = ~n_17561 & ~n_17562;
assign n_17564 =  n_17235 &  n_17563;
assign n_17565 = ~x_3045 &  n_17241;
assign n_17566 = ~i_13 & ~n_17241;
assign n_17567 = ~n_17235 & ~n_17566;
assign n_17568 = ~n_17565 &  n_17567;
assign n_17569 = ~n_17564 & ~n_17568;
assign n_17570 =  n_8055 & ~n_17569;
assign n_17571 =  x_2823 &  n_761;
assign n_17572 =  x_792 & ~n_8051;
assign n_17573 = ~n_17571 & ~n_17572;
assign n_17574 = ~n_17570 &  n_17573;
assign n_17575 =  x_792 & ~n_17574;
assign n_17576 = ~x_792 &  n_17574;
assign n_17577 = ~n_17575 & ~n_17576;
assign n_17578 = ~x_2822 & ~x_3255;
assign n_17579 = ~x_2886 &  x_3255;
assign n_17580 = ~n_17578 & ~n_17579;
assign n_17581 =  n_17235 &  n_17580;
assign n_17582 = ~x_3044 &  n_17241;
assign n_17583 = ~i_12 & ~n_17241;
assign n_17584 = ~n_17235 & ~n_17583;
assign n_17585 = ~n_17582 &  n_17584;
assign n_17586 = ~n_17581 & ~n_17585;
assign n_17587 =  n_8055 & ~n_17586;
assign n_17588 =  x_2822 &  n_761;
assign n_17589 =  x_791 & ~n_8051;
assign n_17590 = ~n_17588 & ~n_17589;
assign n_17591 = ~n_17587 &  n_17590;
assign n_17592 =  x_791 & ~n_17591;
assign n_17593 = ~x_791 &  n_17591;
assign n_17594 = ~n_17592 & ~n_17593;
assign n_17595 = ~x_2821 & ~x_3255;
assign n_17596 = ~x_2885 &  x_3255;
assign n_17597 = ~n_17595 & ~n_17596;
assign n_17598 =  n_17235 &  n_17597;
assign n_17599 = ~x_3043 &  n_17241;
assign n_17600 = ~i_11 & ~n_17241;
assign n_17601 = ~n_17235 & ~n_17600;
assign n_17602 = ~n_17599 &  n_17601;
assign n_17603 = ~n_17598 & ~n_17602;
assign n_17604 =  n_8055 & ~n_17603;
assign n_17605 =  x_2821 &  n_761;
assign n_17606 =  x_790 & ~n_8051;
assign n_17607 = ~n_17605 & ~n_17606;
assign n_17608 = ~n_17604 &  n_17607;
assign n_17609 =  x_790 & ~n_17608;
assign n_17610 = ~x_790 &  n_17608;
assign n_17611 = ~n_17609 & ~n_17610;
assign n_17612 = ~x_2820 & ~x_3255;
assign n_17613 = ~x_2884 &  x_3255;
assign n_17614 = ~n_17612 & ~n_17613;
assign n_17615 =  n_17235 &  n_17614;
assign n_17616 = ~x_3042 &  n_17241;
assign n_17617 = ~i_10 & ~n_17241;
assign n_17618 = ~n_17235 & ~n_17617;
assign n_17619 = ~n_17616 &  n_17618;
assign n_17620 = ~n_17615 & ~n_17619;
assign n_17621 =  n_8055 & ~n_17620;
assign n_17622 =  x_2820 &  n_761;
assign n_17623 =  x_789 & ~n_8051;
assign n_17624 = ~n_17622 & ~n_17623;
assign n_17625 = ~n_17621 &  n_17624;
assign n_17626 =  x_789 & ~n_17625;
assign n_17627 = ~x_789 &  n_17625;
assign n_17628 = ~n_17626 & ~n_17627;
assign n_17629 = ~x_2819 & ~x_3255;
assign n_17630 = ~x_2883 &  x_3255;
assign n_17631 = ~n_17629 & ~n_17630;
assign n_17632 =  n_17235 &  n_17631;
assign n_17633 = ~x_3041 &  n_17241;
assign n_17634 = ~i_9 & ~n_17241;
assign n_17635 = ~n_17235 & ~n_17634;
assign n_17636 = ~n_17633 &  n_17635;
assign n_17637 = ~n_17632 & ~n_17636;
assign n_17638 =  n_8055 & ~n_17637;
assign n_17639 =  x_2819 &  n_761;
assign n_17640 =  x_788 & ~n_8051;
assign n_17641 = ~n_17639 & ~n_17640;
assign n_17642 = ~n_17638 &  n_17641;
assign n_17643 =  x_788 & ~n_17642;
assign n_17644 = ~x_788 &  n_17642;
assign n_17645 = ~n_17643 & ~n_17644;
assign n_17646 = ~x_2818 & ~x_3255;
assign n_17647 = ~x_2882 &  x_3255;
assign n_17648 = ~n_17646 & ~n_17647;
assign n_17649 =  n_17235 &  n_17648;
assign n_17650 = ~x_3040 &  n_17241;
assign n_17651 = ~i_8 & ~n_17241;
assign n_17652 = ~n_17235 & ~n_17651;
assign n_17653 = ~n_17650 &  n_17652;
assign n_17654 = ~n_17649 & ~n_17653;
assign n_17655 =  n_8055 & ~n_17654;
assign n_17656 =  x_2818 &  n_761;
assign n_17657 =  x_787 & ~n_8051;
assign n_17658 = ~n_17656 & ~n_17657;
assign n_17659 = ~n_17655 &  n_17658;
assign n_17660 =  x_787 & ~n_17659;
assign n_17661 = ~x_787 &  n_17659;
assign n_17662 = ~n_17660 & ~n_17661;
assign n_17663 = ~x_2817 & ~x_3255;
assign n_17664 = ~x_2881 &  x_3255;
assign n_17665 = ~n_17663 & ~n_17664;
assign n_17666 =  n_17235 &  n_17665;
assign n_17667 = ~x_3039 &  n_17241;
assign n_17668 = ~i_7 & ~n_17241;
assign n_17669 = ~n_17235 & ~n_17668;
assign n_17670 = ~n_17667 &  n_17669;
assign n_17671 = ~n_17666 & ~n_17670;
assign n_17672 =  n_8055 & ~n_17671;
assign n_17673 =  x_2817 &  n_761;
assign n_17674 =  x_786 & ~n_8051;
assign n_17675 = ~n_17673 & ~n_17674;
assign n_17676 = ~n_17672 &  n_17675;
assign n_17677 =  x_786 & ~n_17676;
assign n_17678 = ~x_786 &  n_17676;
assign n_17679 = ~n_17677 & ~n_17678;
assign n_17680 = ~x_2816 & ~x_3255;
assign n_17681 = ~x_2880 &  x_3255;
assign n_17682 = ~n_17680 & ~n_17681;
assign n_17683 =  n_17235 &  n_17682;
assign n_17684 = ~x_3038 &  n_17241;
assign n_17685 = ~i_6 & ~n_17241;
assign n_17686 = ~n_17235 & ~n_17685;
assign n_17687 = ~n_17684 &  n_17686;
assign n_17688 = ~n_17683 & ~n_17687;
assign n_17689 =  n_8055 & ~n_17688;
assign n_17690 =  x_2816 &  n_761;
assign n_17691 =  x_785 & ~n_8051;
assign n_17692 = ~n_17690 & ~n_17691;
assign n_17693 = ~n_17689 &  n_17692;
assign n_17694 =  x_785 & ~n_17693;
assign n_17695 = ~x_785 &  n_17693;
assign n_17696 = ~n_17694 & ~n_17695;
assign n_17697 = ~x_2815 & ~x_3255;
assign n_17698 = ~x_2879 &  x_3255;
assign n_17699 = ~n_17697 & ~n_17698;
assign n_17700 =  n_17235 &  n_17699;
assign n_17701 = ~x_3037 &  n_17241;
assign n_17702 = ~i_5 & ~n_17241;
assign n_17703 = ~n_17235 & ~n_17702;
assign n_17704 = ~n_17701 &  n_17703;
assign n_17705 = ~n_17700 & ~n_17704;
assign n_17706 =  n_8055 & ~n_17705;
assign n_17707 =  x_2815 &  n_761;
assign n_17708 =  x_784 & ~n_8051;
assign n_17709 = ~n_17707 & ~n_17708;
assign n_17710 = ~n_17706 &  n_17709;
assign n_17711 =  x_784 & ~n_17710;
assign n_17712 = ~x_784 &  n_17710;
assign n_17713 = ~n_17711 & ~n_17712;
assign n_17714 = ~x_2814 & ~x_3255;
assign n_17715 = ~x_2878 &  x_3255;
assign n_17716 = ~n_17714 & ~n_17715;
assign n_17717 =  n_17235 &  n_17716;
assign n_17718 = ~x_3036 &  n_17241;
assign n_17719 = ~i_4 & ~n_17241;
assign n_17720 = ~n_17235 & ~n_17719;
assign n_17721 = ~n_17718 &  n_17720;
assign n_17722 = ~n_17717 & ~n_17721;
assign n_17723 =  n_8055 & ~n_17722;
assign n_17724 =  x_2814 &  n_761;
assign n_17725 =  x_783 & ~n_8051;
assign n_17726 = ~n_17724 & ~n_17725;
assign n_17727 = ~n_17723 &  n_17726;
assign n_17728 =  x_783 & ~n_17727;
assign n_17729 = ~x_783 &  n_17727;
assign n_17730 = ~n_17728 & ~n_17729;
assign n_17731 = ~x_2813 & ~x_3255;
assign n_17732 = ~x_2877 &  x_3255;
assign n_17733 = ~n_17731 & ~n_17732;
assign n_17734 =  n_17235 &  n_17733;
assign n_17735 = ~x_3035 &  n_17241;
assign n_17736 = ~i_3 & ~n_17241;
assign n_17737 = ~n_17235 & ~n_17736;
assign n_17738 = ~n_17735 &  n_17737;
assign n_17739 = ~n_17734 & ~n_17738;
assign n_17740 =  n_8055 & ~n_17739;
assign n_17741 =  x_2813 &  n_761;
assign n_17742 =  x_782 & ~n_8051;
assign n_17743 = ~n_17741 & ~n_17742;
assign n_17744 = ~n_17740 &  n_17743;
assign n_17745 =  x_782 & ~n_17744;
assign n_17746 = ~x_782 &  n_17744;
assign n_17747 = ~n_17745 & ~n_17746;
assign n_17748 = ~x_2812 & ~x_3255;
assign n_17749 = ~x_2876 &  x_3255;
assign n_17750 = ~n_17748 & ~n_17749;
assign n_17751 =  n_17235 &  n_17750;
assign n_17752 = ~x_3034 &  n_17241;
assign n_17753 = ~i_2 & ~n_17241;
assign n_17754 = ~n_17235 & ~n_17753;
assign n_17755 = ~n_17752 &  n_17754;
assign n_17756 = ~n_17751 & ~n_17755;
assign n_17757 =  n_8055 & ~n_17756;
assign n_17758 =  x_2812 &  n_761;
assign n_17759 =  x_781 & ~n_8051;
assign n_17760 = ~n_17758 & ~n_17759;
assign n_17761 = ~n_17757 &  n_17760;
assign n_17762 =  x_781 & ~n_17761;
assign n_17763 = ~x_781 &  n_17761;
assign n_17764 = ~n_17762 & ~n_17763;
assign n_17765 = ~x_2811 & ~x_3255;
assign n_17766 = ~x_2875 &  x_3255;
assign n_17767 = ~n_17765 & ~n_17766;
assign n_17768 =  n_17235 &  n_17767;
assign n_17769 = ~x_3033 &  n_17241;
assign n_17770 = ~i_1 & ~n_17241;
assign n_17771 = ~n_17235 & ~n_17770;
assign n_17772 = ~n_17769 &  n_17771;
assign n_17773 = ~n_17768 & ~n_17772;
assign n_17774 =  n_8055 & ~n_17773;
assign n_17775 =  x_2811 &  n_761;
assign n_17776 =  x_780 & ~n_8051;
assign n_17777 = ~n_17775 & ~n_17776;
assign n_17778 = ~n_17774 &  n_17777;
assign n_17779 =  x_780 & ~n_17778;
assign n_17780 = ~x_780 &  n_17778;
assign n_17781 = ~n_17779 & ~n_17780;
assign n_17782 =  x_37 &  n_765;
assign n_17783 = ~x_38 &  n_17782;
assign n_17784 =  x_39 &  n_17783;
assign n_17785 = ~x_42 &  n_561;
assign n_17786 =  n_17784 &  n_17785;
assign n_17787 = ~x_43 &  n_17786;
assign n_17788 =  x_779 & ~n_17787;
assign n_17789 =  i_32 &  n_17787;
assign n_17790 = ~n_17788 & ~n_17789;
assign n_17791 =  x_779 & ~n_17790;
assign n_17792 = ~x_779 &  n_17790;
assign n_17793 = ~n_17791 & ~n_17792;
assign n_17794 =  x_778 & ~n_17787;
assign n_17795 =  i_31 &  n_17787;
assign n_17796 = ~n_17794 & ~n_17795;
assign n_17797 =  x_778 & ~n_17796;
assign n_17798 = ~x_778 &  n_17796;
assign n_17799 = ~n_17797 & ~n_17798;
assign n_17800 =  x_777 & ~n_17787;
assign n_17801 =  i_30 &  n_17787;
assign n_17802 = ~n_17800 & ~n_17801;
assign n_17803 =  x_777 & ~n_17802;
assign n_17804 = ~x_777 &  n_17802;
assign n_17805 = ~n_17803 & ~n_17804;
assign n_17806 =  x_776 & ~n_17787;
assign n_17807 =  i_29 &  n_17787;
assign n_17808 = ~n_17806 & ~n_17807;
assign n_17809 =  x_776 & ~n_17808;
assign n_17810 = ~x_776 &  n_17808;
assign n_17811 = ~n_17809 & ~n_17810;
assign n_17812 =  x_775 & ~n_17787;
assign n_17813 =  i_28 &  n_17787;
assign n_17814 = ~n_17812 & ~n_17813;
assign n_17815 =  x_775 & ~n_17814;
assign n_17816 = ~x_775 &  n_17814;
assign n_17817 = ~n_17815 & ~n_17816;
assign n_17818 =  x_774 & ~n_17787;
assign n_17819 =  i_27 &  n_17787;
assign n_17820 = ~n_17818 & ~n_17819;
assign n_17821 =  x_774 & ~n_17820;
assign n_17822 = ~x_774 &  n_17820;
assign n_17823 = ~n_17821 & ~n_17822;
assign n_17824 =  x_773 & ~n_17787;
assign n_17825 =  i_26 &  n_17787;
assign n_17826 = ~n_17824 & ~n_17825;
assign n_17827 =  x_773 & ~n_17826;
assign n_17828 = ~x_773 &  n_17826;
assign n_17829 = ~n_17827 & ~n_17828;
assign n_17830 =  x_772 & ~n_17787;
assign n_17831 =  i_25 &  n_17787;
assign n_17832 = ~n_17830 & ~n_17831;
assign n_17833 =  x_772 & ~n_17832;
assign n_17834 = ~x_772 &  n_17832;
assign n_17835 = ~n_17833 & ~n_17834;
assign n_17836 =  x_771 & ~n_17787;
assign n_17837 =  i_24 &  n_17787;
assign n_17838 = ~n_17836 & ~n_17837;
assign n_17839 =  x_771 & ~n_17838;
assign n_17840 = ~x_771 &  n_17838;
assign n_17841 = ~n_17839 & ~n_17840;
assign n_17842 =  x_770 & ~n_17787;
assign n_17843 =  i_23 &  n_17787;
assign n_17844 = ~n_17842 & ~n_17843;
assign n_17845 =  x_770 & ~n_17844;
assign n_17846 = ~x_770 &  n_17844;
assign n_17847 = ~n_17845 & ~n_17846;
assign n_17848 =  x_769 & ~n_17787;
assign n_17849 =  i_22 &  n_17787;
assign n_17850 = ~n_17848 & ~n_17849;
assign n_17851 =  x_769 & ~n_17850;
assign n_17852 = ~x_769 &  n_17850;
assign n_17853 = ~n_17851 & ~n_17852;
assign n_17854 =  x_768 & ~n_17787;
assign n_17855 =  i_21 &  n_17787;
assign n_17856 = ~n_17854 & ~n_17855;
assign n_17857 =  x_768 & ~n_17856;
assign n_17858 = ~x_768 &  n_17856;
assign n_17859 = ~n_17857 & ~n_17858;
assign n_17860 =  x_767 & ~n_17787;
assign n_17861 =  i_20 &  n_17787;
assign n_17862 = ~n_17860 & ~n_17861;
assign n_17863 =  x_767 & ~n_17862;
assign n_17864 = ~x_767 &  n_17862;
assign n_17865 = ~n_17863 & ~n_17864;
assign n_17866 =  x_766 & ~n_17787;
assign n_17867 =  i_19 &  n_17787;
assign n_17868 = ~n_17866 & ~n_17867;
assign n_17869 =  x_766 & ~n_17868;
assign n_17870 = ~x_766 &  n_17868;
assign n_17871 = ~n_17869 & ~n_17870;
assign n_17872 =  x_765 & ~n_17787;
assign n_17873 =  i_18 &  n_17787;
assign n_17874 = ~n_17872 & ~n_17873;
assign n_17875 =  x_765 & ~n_17874;
assign n_17876 = ~x_765 &  n_17874;
assign n_17877 = ~n_17875 & ~n_17876;
assign n_17878 =  x_764 & ~n_17787;
assign n_17879 =  i_17 &  n_17787;
assign n_17880 = ~n_17878 & ~n_17879;
assign n_17881 =  x_764 & ~n_17880;
assign n_17882 = ~x_764 &  n_17880;
assign n_17883 = ~n_17881 & ~n_17882;
assign n_17884 =  x_763 & ~n_17787;
assign n_17885 =  i_16 &  n_17787;
assign n_17886 = ~n_17884 & ~n_17885;
assign n_17887 =  x_763 & ~n_17886;
assign n_17888 = ~x_763 &  n_17886;
assign n_17889 = ~n_17887 & ~n_17888;
assign n_17890 =  x_762 & ~n_17787;
assign n_17891 =  i_15 &  n_17787;
assign n_17892 = ~n_17890 & ~n_17891;
assign n_17893 =  x_762 & ~n_17892;
assign n_17894 = ~x_762 &  n_17892;
assign n_17895 = ~n_17893 & ~n_17894;
assign n_17896 =  x_761 & ~n_17787;
assign n_17897 =  i_14 &  n_17787;
assign n_17898 = ~n_17896 & ~n_17897;
assign n_17899 =  x_761 & ~n_17898;
assign n_17900 = ~x_761 &  n_17898;
assign n_17901 = ~n_17899 & ~n_17900;
assign n_17902 =  x_760 & ~n_17787;
assign n_17903 =  i_13 &  n_17787;
assign n_17904 = ~n_17902 & ~n_17903;
assign n_17905 =  x_760 & ~n_17904;
assign n_17906 = ~x_760 &  n_17904;
assign n_17907 = ~n_17905 & ~n_17906;
assign n_17908 =  x_759 & ~n_17787;
assign n_17909 =  i_12 &  n_17787;
assign n_17910 = ~n_17908 & ~n_17909;
assign n_17911 =  x_759 & ~n_17910;
assign n_17912 = ~x_759 &  n_17910;
assign n_17913 = ~n_17911 & ~n_17912;
assign n_17914 =  x_758 & ~n_17787;
assign n_17915 =  i_11 &  n_17787;
assign n_17916 = ~n_17914 & ~n_17915;
assign n_17917 =  x_758 & ~n_17916;
assign n_17918 = ~x_758 &  n_17916;
assign n_17919 = ~n_17917 & ~n_17918;
assign n_17920 =  x_757 & ~n_17787;
assign n_17921 =  i_10 &  n_17787;
assign n_17922 = ~n_17920 & ~n_17921;
assign n_17923 =  x_757 & ~n_17922;
assign n_17924 = ~x_757 &  n_17922;
assign n_17925 = ~n_17923 & ~n_17924;
assign n_17926 =  x_756 & ~n_17787;
assign n_17927 =  i_9 &  n_17787;
assign n_17928 = ~n_17926 & ~n_17927;
assign n_17929 =  x_756 & ~n_17928;
assign n_17930 = ~x_756 &  n_17928;
assign n_17931 = ~n_17929 & ~n_17930;
assign n_17932 =  x_755 & ~n_17787;
assign n_17933 =  i_8 &  n_17787;
assign n_17934 = ~n_17932 & ~n_17933;
assign n_17935 =  x_755 & ~n_17934;
assign n_17936 = ~x_755 &  n_17934;
assign n_17937 = ~n_17935 & ~n_17936;
assign n_17938 =  x_754 & ~n_17787;
assign n_17939 =  i_7 &  n_17787;
assign n_17940 = ~n_17938 & ~n_17939;
assign n_17941 =  x_754 & ~n_17940;
assign n_17942 = ~x_754 &  n_17940;
assign n_17943 = ~n_17941 & ~n_17942;
assign n_17944 =  x_753 & ~n_17787;
assign n_17945 =  i_6 &  n_17787;
assign n_17946 = ~n_17944 & ~n_17945;
assign n_17947 =  x_753 & ~n_17946;
assign n_17948 = ~x_753 &  n_17946;
assign n_17949 = ~n_17947 & ~n_17948;
assign n_17950 =  x_752 & ~n_17787;
assign n_17951 =  i_5 &  n_17787;
assign n_17952 = ~n_17950 & ~n_17951;
assign n_17953 =  x_752 & ~n_17952;
assign n_17954 = ~x_752 &  n_17952;
assign n_17955 = ~n_17953 & ~n_17954;
assign n_17956 =  x_751 & ~n_17787;
assign n_17957 =  i_4 &  n_17787;
assign n_17958 = ~n_17956 & ~n_17957;
assign n_17959 =  x_751 & ~n_17958;
assign n_17960 = ~x_751 &  n_17958;
assign n_17961 = ~n_17959 & ~n_17960;
assign n_17962 =  x_750 & ~n_17787;
assign n_17963 =  i_3 &  n_17787;
assign n_17964 = ~n_17962 & ~n_17963;
assign n_17965 =  x_750 & ~n_17964;
assign n_17966 = ~x_750 &  n_17964;
assign n_17967 = ~n_17965 & ~n_17966;
assign n_17968 =  x_749 & ~n_17787;
assign n_17969 =  i_2 &  n_17787;
assign n_17970 = ~n_17968 & ~n_17969;
assign n_17971 =  x_749 & ~n_17970;
assign n_17972 = ~x_749 &  n_17970;
assign n_17973 = ~n_17971 & ~n_17972;
assign n_17974 =  x_748 & ~n_17787;
assign n_17975 =  i_1 &  n_17787;
assign n_17976 = ~n_17974 & ~n_17975;
assign n_17977 =  x_748 & ~n_17976;
assign n_17978 = ~x_748 &  n_17976;
assign n_17979 = ~n_17977 & ~n_17978;
assign n_17980 =  n_15366 &  n_2096;
assign n_17981 =  x_747 & ~n_17980;
assign n_17982 =  x_747 &  n_17981;
assign n_17983 = ~x_747 & ~n_17981;
assign n_17984 = ~n_17982 & ~n_17983;
assign n_17985 =  x_746 & ~n_17980;
assign n_17986 =  x_746 &  n_17985;
assign n_17987 = ~x_746 & ~n_17985;
assign n_17988 = ~n_17986 & ~n_17987;
assign n_17989 =  x_745 & ~n_17980;
assign n_17990 =  x_745 &  n_17989;
assign n_17991 = ~x_745 & ~n_17989;
assign n_17992 = ~n_17990 & ~n_17991;
assign n_17993 =  x_744 & ~n_17980;
assign n_17994 =  x_744 &  n_17993;
assign n_17995 = ~x_744 & ~n_17993;
assign n_17996 = ~n_17994 & ~n_17995;
assign n_17997 =  x_743 & ~n_17980;
assign n_17998 =  x_743 &  n_17997;
assign n_17999 = ~x_743 & ~n_17997;
assign n_18000 = ~n_17998 & ~n_17999;
assign n_18001 =  x_742 & ~n_17980;
assign n_18002 =  x_742 &  n_18001;
assign n_18003 = ~x_742 & ~n_18001;
assign n_18004 = ~n_18002 & ~n_18003;
assign n_18005 =  x_741 & ~n_17980;
assign n_18006 =  x_741 &  n_18005;
assign n_18007 = ~x_741 & ~n_18005;
assign n_18008 = ~n_18006 & ~n_18007;
assign n_18009 =  x_740 & ~n_17980;
assign n_18010 =  x_740 &  n_18009;
assign n_18011 = ~x_740 & ~n_18009;
assign n_18012 = ~n_18010 & ~n_18011;
assign n_18013 =  x_739 & ~n_17980;
assign n_18014 =  x_739 &  n_18013;
assign n_18015 = ~x_739 & ~n_18013;
assign n_18016 = ~n_18014 & ~n_18015;
assign n_18017 =  x_738 & ~n_17980;
assign n_18018 =  x_738 &  n_18017;
assign n_18019 = ~x_738 & ~n_18017;
assign n_18020 = ~n_18018 & ~n_18019;
assign n_18021 =  x_737 & ~n_17980;
assign n_18022 =  x_737 &  n_18021;
assign n_18023 = ~x_737 & ~n_18021;
assign n_18024 = ~n_18022 & ~n_18023;
assign n_18025 =  x_736 & ~n_17980;
assign n_18026 =  x_736 &  n_18025;
assign n_18027 = ~x_736 & ~n_18025;
assign n_18028 = ~n_18026 & ~n_18027;
assign n_18029 =  x_735 & ~n_17980;
assign n_18030 =  x_735 &  n_18029;
assign n_18031 = ~x_735 & ~n_18029;
assign n_18032 = ~n_18030 & ~n_18031;
assign n_18033 =  x_734 & ~n_17980;
assign n_18034 =  x_734 &  n_18033;
assign n_18035 = ~x_734 & ~n_18033;
assign n_18036 = ~n_18034 & ~n_18035;
assign n_18037 =  x_733 & ~n_17980;
assign n_18038 =  x_733 &  n_18037;
assign n_18039 = ~x_733 & ~n_18037;
assign n_18040 = ~n_18038 & ~n_18039;
assign n_18041 =  x_732 & ~n_17980;
assign n_18042 =  x_732 &  n_18041;
assign n_18043 = ~x_732 & ~n_18041;
assign n_18044 = ~n_18042 & ~n_18043;
assign n_18045 =  x_731 & ~n_17980;
assign n_18046 =  x_731 &  n_18045;
assign n_18047 = ~x_731 & ~n_18045;
assign n_18048 = ~n_18046 & ~n_18047;
assign n_18049 =  x_730 & ~n_17980;
assign n_18050 =  x_730 &  n_18049;
assign n_18051 = ~x_730 & ~n_18049;
assign n_18052 = ~n_18050 & ~n_18051;
assign n_18053 =  x_729 & ~n_17980;
assign n_18054 =  x_729 &  n_18053;
assign n_18055 = ~x_729 & ~n_18053;
assign n_18056 = ~n_18054 & ~n_18055;
assign n_18057 =  x_728 & ~n_17980;
assign n_18058 =  x_728 &  n_18057;
assign n_18059 = ~x_728 & ~n_18057;
assign n_18060 = ~n_18058 & ~n_18059;
assign n_18061 =  x_727 & ~n_17980;
assign n_18062 =  x_727 &  n_18061;
assign n_18063 = ~x_727 & ~n_18061;
assign n_18064 = ~n_18062 & ~n_18063;
assign n_18065 =  x_726 & ~n_17980;
assign n_18066 =  x_726 &  n_18065;
assign n_18067 = ~x_726 & ~n_18065;
assign n_18068 = ~n_18066 & ~n_18067;
assign n_18069 =  x_725 & ~n_17980;
assign n_18070 =  x_725 &  n_18069;
assign n_18071 = ~x_725 & ~n_18069;
assign n_18072 = ~n_18070 & ~n_18071;
assign n_18073 =  x_724 & ~n_17980;
assign n_18074 =  x_724 &  n_18073;
assign n_18075 = ~x_724 & ~n_18073;
assign n_18076 = ~n_18074 & ~n_18075;
assign n_18077 =  x_723 & ~n_17980;
assign n_18078 =  x_723 &  n_18077;
assign n_18079 = ~x_723 & ~n_18077;
assign n_18080 = ~n_18078 & ~n_18079;
assign n_18081 =  x_722 & ~n_17980;
assign n_18082 =  x_722 &  n_18081;
assign n_18083 = ~x_722 & ~n_18081;
assign n_18084 = ~n_18082 & ~n_18083;
assign n_18085 =  x_721 & ~n_17980;
assign n_18086 =  x_721 &  n_18085;
assign n_18087 = ~x_721 & ~n_18085;
assign n_18088 = ~n_18086 & ~n_18087;
assign n_18089 =  x_720 & ~n_17980;
assign n_18090 =  x_720 &  n_18089;
assign n_18091 = ~x_720 & ~n_18089;
assign n_18092 = ~n_18090 & ~n_18091;
assign n_18093 =  x_719 & ~n_17980;
assign n_18094 =  x_719 &  n_18093;
assign n_18095 = ~x_719 & ~n_18093;
assign n_18096 = ~n_18094 & ~n_18095;
assign n_18097 =  x_718 & ~n_17980;
assign n_18098 =  x_718 &  n_18097;
assign n_18099 = ~x_718 & ~n_18097;
assign n_18100 = ~n_18098 & ~n_18099;
assign n_18101 =  x_717 & ~n_17980;
assign n_18102 =  x_717 &  n_18101;
assign n_18103 = ~x_717 & ~n_18101;
assign n_18104 = ~n_18102 & ~n_18103;
assign n_18105 =  x_716 & ~n_17980;
assign n_18106 =  x_716 &  n_18105;
assign n_18107 = ~x_716 & ~n_18105;
assign n_18108 = ~n_18106 & ~n_18107;
assign n_18109 =  n_4290 &  n_3625;
assign n_18110 =  x_715 & ~n_18109;
assign n_18111 =  i_32 &  n_18109;
assign n_18112 = ~n_18110 & ~n_18111;
assign n_18113 =  x_715 & ~n_18112;
assign n_18114 = ~x_715 &  n_18112;
assign n_18115 = ~n_18113 & ~n_18114;
assign n_18116 =  x_714 & ~n_18109;
assign n_18117 =  i_31 &  n_18109;
assign n_18118 = ~n_18116 & ~n_18117;
assign n_18119 =  x_714 & ~n_18118;
assign n_18120 = ~x_714 &  n_18118;
assign n_18121 = ~n_18119 & ~n_18120;
assign n_18122 =  x_713 & ~n_18109;
assign n_18123 =  i_30 &  n_18109;
assign n_18124 = ~n_18122 & ~n_18123;
assign n_18125 =  x_713 & ~n_18124;
assign n_18126 = ~x_713 &  n_18124;
assign n_18127 = ~n_18125 & ~n_18126;
assign n_18128 =  x_712 & ~n_18109;
assign n_18129 =  i_29 &  n_18109;
assign n_18130 = ~n_18128 & ~n_18129;
assign n_18131 =  x_712 & ~n_18130;
assign n_18132 = ~x_712 &  n_18130;
assign n_18133 = ~n_18131 & ~n_18132;
assign n_18134 =  x_711 & ~n_18109;
assign n_18135 =  i_28 &  n_18109;
assign n_18136 = ~n_18134 & ~n_18135;
assign n_18137 =  x_711 & ~n_18136;
assign n_18138 = ~x_711 &  n_18136;
assign n_18139 = ~n_18137 & ~n_18138;
assign n_18140 =  x_710 & ~n_18109;
assign n_18141 =  i_27 &  n_18109;
assign n_18142 = ~n_18140 & ~n_18141;
assign n_18143 =  x_710 & ~n_18142;
assign n_18144 = ~x_710 &  n_18142;
assign n_18145 = ~n_18143 & ~n_18144;
assign n_18146 =  x_709 & ~n_18109;
assign n_18147 =  i_26 &  n_18109;
assign n_18148 = ~n_18146 & ~n_18147;
assign n_18149 =  x_709 & ~n_18148;
assign n_18150 = ~x_709 &  n_18148;
assign n_18151 = ~n_18149 & ~n_18150;
assign n_18152 =  x_708 & ~n_18109;
assign n_18153 =  i_25 &  n_18109;
assign n_18154 = ~n_18152 & ~n_18153;
assign n_18155 =  x_708 & ~n_18154;
assign n_18156 = ~x_708 &  n_18154;
assign n_18157 = ~n_18155 & ~n_18156;
assign n_18158 =  x_707 & ~n_18109;
assign n_18159 =  i_24 &  n_18109;
assign n_18160 = ~n_18158 & ~n_18159;
assign n_18161 =  x_707 & ~n_18160;
assign n_18162 = ~x_707 &  n_18160;
assign n_18163 = ~n_18161 & ~n_18162;
assign n_18164 =  x_706 & ~n_18109;
assign n_18165 =  i_23 &  n_18109;
assign n_18166 = ~n_18164 & ~n_18165;
assign n_18167 =  x_706 & ~n_18166;
assign n_18168 = ~x_706 &  n_18166;
assign n_18169 = ~n_18167 & ~n_18168;
assign n_18170 =  x_705 & ~n_18109;
assign n_18171 =  i_22 &  n_18109;
assign n_18172 = ~n_18170 & ~n_18171;
assign n_18173 =  x_705 & ~n_18172;
assign n_18174 = ~x_705 &  n_18172;
assign n_18175 = ~n_18173 & ~n_18174;
assign n_18176 =  x_704 & ~n_18109;
assign n_18177 =  i_21 &  n_18109;
assign n_18178 = ~n_18176 & ~n_18177;
assign n_18179 =  x_704 & ~n_18178;
assign n_18180 = ~x_704 &  n_18178;
assign n_18181 = ~n_18179 & ~n_18180;
assign n_18182 =  x_703 & ~n_18109;
assign n_18183 =  i_20 &  n_18109;
assign n_18184 = ~n_18182 & ~n_18183;
assign n_18185 =  x_703 & ~n_18184;
assign n_18186 = ~x_703 &  n_18184;
assign n_18187 = ~n_18185 & ~n_18186;
assign n_18188 =  x_702 & ~n_18109;
assign n_18189 =  i_19 &  n_18109;
assign n_18190 = ~n_18188 & ~n_18189;
assign n_18191 =  x_702 & ~n_18190;
assign n_18192 = ~x_702 &  n_18190;
assign n_18193 = ~n_18191 & ~n_18192;
assign n_18194 =  x_701 & ~n_18109;
assign n_18195 =  i_18 &  n_18109;
assign n_18196 = ~n_18194 & ~n_18195;
assign n_18197 =  x_701 & ~n_18196;
assign n_18198 = ~x_701 &  n_18196;
assign n_18199 = ~n_18197 & ~n_18198;
assign n_18200 =  x_700 & ~n_18109;
assign n_18201 =  i_17 &  n_18109;
assign n_18202 = ~n_18200 & ~n_18201;
assign n_18203 =  x_700 & ~n_18202;
assign n_18204 = ~x_700 &  n_18202;
assign n_18205 = ~n_18203 & ~n_18204;
assign n_18206 =  x_699 & ~n_18109;
assign n_18207 =  i_16 &  n_18109;
assign n_18208 = ~n_18206 & ~n_18207;
assign n_18209 =  x_699 & ~n_18208;
assign n_18210 = ~x_699 &  n_18208;
assign n_18211 = ~n_18209 & ~n_18210;
assign n_18212 =  x_698 & ~n_18109;
assign n_18213 =  i_15 &  n_18109;
assign n_18214 = ~n_18212 & ~n_18213;
assign n_18215 =  x_698 & ~n_18214;
assign n_18216 = ~x_698 &  n_18214;
assign n_18217 = ~n_18215 & ~n_18216;
assign n_18218 =  x_697 & ~n_18109;
assign n_18219 =  i_14 &  n_18109;
assign n_18220 = ~n_18218 & ~n_18219;
assign n_18221 =  x_697 & ~n_18220;
assign n_18222 = ~x_697 &  n_18220;
assign n_18223 = ~n_18221 & ~n_18222;
assign n_18224 =  x_696 & ~n_18109;
assign n_18225 =  i_13 &  n_18109;
assign n_18226 = ~n_18224 & ~n_18225;
assign n_18227 =  x_696 & ~n_18226;
assign n_18228 = ~x_696 &  n_18226;
assign n_18229 = ~n_18227 & ~n_18228;
assign n_18230 =  x_695 & ~n_18109;
assign n_18231 =  i_12 &  n_18109;
assign n_18232 = ~n_18230 & ~n_18231;
assign n_18233 =  x_695 & ~n_18232;
assign n_18234 = ~x_695 &  n_18232;
assign n_18235 = ~n_18233 & ~n_18234;
assign n_18236 =  x_694 & ~n_18109;
assign n_18237 =  i_11 &  n_18109;
assign n_18238 = ~n_18236 & ~n_18237;
assign n_18239 =  x_694 & ~n_18238;
assign n_18240 = ~x_694 &  n_18238;
assign n_18241 = ~n_18239 & ~n_18240;
assign n_18242 =  x_693 & ~n_18109;
assign n_18243 =  i_10 &  n_18109;
assign n_18244 = ~n_18242 & ~n_18243;
assign n_18245 =  x_693 & ~n_18244;
assign n_18246 = ~x_693 &  n_18244;
assign n_18247 = ~n_18245 & ~n_18246;
assign n_18248 =  x_692 & ~n_18109;
assign n_18249 =  i_9 &  n_18109;
assign n_18250 = ~n_18248 & ~n_18249;
assign n_18251 =  x_692 & ~n_18250;
assign n_18252 = ~x_692 &  n_18250;
assign n_18253 = ~n_18251 & ~n_18252;
assign n_18254 =  x_691 & ~n_18109;
assign n_18255 =  i_8 &  n_18109;
assign n_18256 = ~n_18254 & ~n_18255;
assign n_18257 =  x_691 & ~n_18256;
assign n_18258 = ~x_691 &  n_18256;
assign n_18259 = ~n_18257 & ~n_18258;
assign n_18260 =  x_690 & ~n_18109;
assign n_18261 =  i_7 &  n_18109;
assign n_18262 = ~n_18260 & ~n_18261;
assign n_18263 =  x_690 & ~n_18262;
assign n_18264 = ~x_690 &  n_18262;
assign n_18265 = ~n_18263 & ~n_18264;
assign n_18266 =  x_689 & ~n_18109;
assign n_18267 =  i_6 &  n_18109;
assign n_18268 = ~n_18266 & ~n_18267;
assign n_18269 =  x_689 & ~n_18268;
assign n_18270 = ~x_689 &  n_18268;
assign n_18271 = ~n_18269 & ~n_18270;
assign n_18272 =  x_688 & ~n_18109;
assign n_18273 =  i_5 &  n_18109;
assign n_18274 = ~n_18272 & ~n_18273;
assign n_18275 =  x_688 & ~n_18274;
assign n_18276 = ~x_688 &  n_18274;
assign n_18277 = ~n_18275 & ~n_18276;
assign n_18278 =  x_687 & ~n_18109;
assign n_18279 =  i_4 &  n_18109;
assign n_18280 = ~n_18278 & ~n_18279;
assign n_18281 =  x_687 & ~n_18280;
assign n_18282 = ~x_687 &  n_18280;
assign n_18283 = ~n_18281 & ~n_18282;
assign n_18284 =  x_686 & ~n_18109;
assign n_18285 =  i_3 &  n_18109;
assign n_18286 = ~n_18284 & ~n_18285;
assign n_18287 =  x_686 & ~n_18286;
assign n_18288 = ~x_686 &  n_18286;
assign n_18289 = ~n_18287 & ~n_18288;
assign n_18290 =  x_685 & ~n_18109;
assign n_18291 =  i_2 &  n_18109;
assign n_18292 = ~n_18290 & ~n_18291;
assign n_18293 =  x_685 & ~n_18292;
assign n_18294 = ~x_685 &  n_18292;
assign n_18295 = ~n_18293 & ~n_18294;
assign n_18296 =  x_684 & ~n_18109;
assign n_18297 =  i_1 &  n_18109;
assign n_18298 = ~n_18296 & ~n_18297;
assign n_18299 =  x_684 & ~n_18298;
assign n_18300 = ~x_684 &  n_18298;
assign n_18301 = ~n_18299 & ~n_18300;
assign n_18302 =  x_43 &  n_17786;
assign n_18303 =  x_683 & ~n_18302;
assign n_18304 =  i_32 &  n_18302;
assign n_18305 = ~n_18303 & ~n_18304;
assign n_18306 =  x_683 & ~n_18305;
assign n_18307 = ~x_683 &  n_18305;
assign n_18308 = ~n_18306 & ~n_18307;
assign n_18309 =  x_682 & ~n_18302;
assign n_18310 =  i_31 &  n_18302;
assign n_18311 = ~n_18309 & ~n_18310;
assign n_18312 =  x_682 & ~n_18311;
assign n_18313 = ~x_682 &  n_18311;
assign n_18314 = ~n_18312 & ~n_18313;
assign n_18315 =  x_681 & ~n_18302;
assign n_18316 =  i_30 &  n_18302;
assign n_18317 = ~n_18315 & ~n_18316;
assign n_18318 =  x_681 & ~n_18317;
assign n_18319 = ~x_681 &  n_18317;
assign n_18320 = ~n_18318 & ~n_18319;
assign n_18321 =  x_680 & ~n_18302;
assign n_18322 =  i_29 &  n_18302;
assign n_18323 = ~n_18321 & ~n_18322;
assign n_18324 =  x_680 & ~n_18323;
assign n_18325 = ~x_680 &  n_18323;
assign n_18326 = ~n_18324 & ~n_18325;
assign n_18327 =  x_679 & ~n_18302;
assign n_18328 =  i_28 &  n_18302;
assign n_18329 = ~n_18327 & ~n_18328;
assign n_18330 =  x_679 & ~n_18329;
assign n_18331 = ~x_679 &  n_18329;
assign n_18332 = ~n_18330 & ~n_18331;
assign n_18333 =  x_678 & ~n_18302;
assign n_18334 =  i_27 &  n_18302;
assign n_18335 = ~n_18333 & ~n_18334;
assign n_18336 =  x_678 & ~n_18335;
assign n_18337 = ~x_678 &  n_18335;
assign n_18338 = ~n_18336 & ~n_18337;
assign n_18339 =  x_677 & ~n_18302;
assign n_18340 =  i_26 &  n_18302;
assign n_18341 = ~n_18339 & ~n_18340;
assign n_18342 =  x_677 & ~n_18341;
assign n_18343 = ~x_677 &  n_18341;
assign n_18344 = ~n_18342 & ~n_18343;
assign n_18345 =  x_676 & ~n_18302;
assign n_18346 =  i_25 &  n_18302;
assign n_18347 = ~n_18345 & ~n_18346;
assign n_18348 =  x_676 & ~n_18347;
assign n_18349 = ~x_676 &  n_18347;
assign n_18350 = ~n_18348 & ~n_18349;
assign n_18351 =  x_675 & ~n_18302;
assign n_18352 =  i_24 &  n_18302;
assign n_18353 = ~n_18351 & ~n_18352;
assign n_18354 =  x_675 & ~n_18353;
assign n_18355 = ~x_675 &  n_18353;
assign n_18356 = ~n_18354 & ~n_18355;
assign n_18357 =  x_674 & ~n_18302;
assign n_18358 =  i_23 &  n_18302;
assign n_18359 = ~n_18357 & ~n_18358;
assign n_18360 =  x_674 & ~n_18359;
assign n_18361 = ~x_674 &  n_18359;
assign n_18362 = ~n_18360 & ~n_18361;
assign n_18363 =  x_673 & ~n_18302;
assign n_18364 =  i_22 &  n_18302;
assign n_18365 = ~n_18363 & ~n_18364;
assign n_18366 =  x_673 & ~n_18365;
assign n_18367 = ~x_673 &  n_18365;
assign n_18368 = ~n_18366 & ~n_18367;
assign n_18369 =  x_672 & ~n_18302;
assign n_18370 =  i_21 &  n_18302;
assign n_18371 = ~n_18369 & ~n_18370;
assign n_18372 =  x_672 & ~n_18371;
assign n_18373 = ~x_672 &  n_18371;
assign n_18374 = ~n_18372 & ~n_18373;
assign n_18375 =  x_671 & ~n_18302;
assign n_18376 =  i_20 &  n_18302;
assign n_18377 = ~n_18375 & ~n_18376;
assign n_18378 =  x_671 & ~n_18377;
assign n_18379 = ~x_671 &  n_18377;
assign n_18380 = ~n_18378 & ~n_18379;
assign n_18381 =  x_670 & ~n_18302;
assign n_18382 =  i_19 &  n_18302;
assign n_18383 = ~n_18381 & ~n_18382;
assign n_18384 =  x_670 & ~n_18383;
assign n_18385 = ~x_670 &  n_18383;
assign n_18386 = ~n_18384 & ~n_18385;
assign n_18387 =  x_669 & ~n_18302;
assign n_18388 =  i_18 &  n_18302;
assign n_18389 = ~n_18387 & ~n_18388;
assign n_18390 =  x_669 & ~n_18389;
assign n_18391 = ~x_669 &  n_18389;
assign n_18392 = ~n_18390 & ~n_18391;
assign n_18393 =  x_668 & ~n_18302;
assign n_18394 =  i_17 &  n_18302;
assign n_18395 = ~n_18393 & ~n_18394;
assign n_18396 =  x_668 & ~n_18395;
assign n_18397 = ~x_668 &  n_18395;
assign n_18398 = ~n_18396 & ~n_18397;
assign n_18399 =  x_667 & ~n_18302;
assign n_18400 =  i_16 &  n_18302;
assign n_18401 = ~n_18399 & ~n_18400;
assign n_18402 =  x_667 & ~n_18401;
assign n_18403 = ~x_667 &  n_18401;
assign n_18404 = ~n_18402 & ~n_18403;
assign n_18405 =  x_666 & ~n_18302;
assign n_18406 =  i_15 &  n_18302;
assign n_18407 = ~n_18405 & ~n_18406;
assign n_18408 =  x_666 & ~n_18407;
assign n_18409 = ~x_666 &  n_18407;
assign n_18410 = ~n_18408 & ~n_18409;
assign n_18411 =  x_665 & ~n_18302;
assign n_18412 =  i_14 &  n_18302;
assign n_18413 = ~n_18411 & ~n_18412;
assign n_18414 =  x_665 & ~n_18413;
assign n_18415 = ~x_665 &  n_18413;
assign n_18416 = ~n_18414 & ~n_18415;
assign n_18417 =  x_664 & ~n_18302;
assign n_18418 =  i_13 &  n_18302;
assign n_18419 = ~n_18417 & ~n_18418;
assign n_18420 =  x_664 & ~n_18419;
assign n_18421 = ~x_664 &  n_18419;
assign n_18422 = ~n_18420 & ~n_18421;
assign n_18423 =  x_663 & ~n_18302;
assign n_18424 =  i_12 &  n_18302;
assign n_18425 = ~n_18423 & ~n_18424;
assign n_18426 =  x_663 & ~n_18425;
assign n_18427 = ~x_663 &  n_18425;
assign n_18428 = ~n_18426 & ~n_18427;
assign n_18429 =  x_662 & ~n_18302;
assign n_18430 =  i_11 &  n_18302;
assign n_18431 = ~n_18429 & ~n_18430;
assign n_18432 =  x_662 & ~n_18431;
assign n_18433 = ~x_662 &  n_18431;
assign n_18434 = ~n_18432 & ~n_18433;
assign n_18435 =  x_661 & ~n_18302;
assign n_18436 =  i_10 &  n_18302;
assign n_18437 = ~n_18435 & ~n_18436;
assign n_18438 =  x_661 & ~n_18437;
assign n_18439 = ~x_661 &  n_18437;
assign n_18440 = ~n_18438 & ~n_18439;
assign n_18441 =  x_660 & ~n_18302;
assign n_18442 =  i_9 &  n_18302;
assign n_18443 = ~n_18441 & ~n_18442;
assign n_18444 =  x_660 & ~n_18443;
assign n_18445 = ~x_660 &  n_18443;
assign n_18446 = ~n_18444 & ~n_18445;
assign n_18447 =  x_659 & ~n_18302;
assign n_18448 =  i_8 &  n_18302;
assign n_18449 = ~n_18447 & ~n_18448;
assign n_18450 =  x_659 & ~n_18449;
assign n_18451 = ~x_659 &  n_18449;
assign n_18452 = ~n_18450 & ~n_18451;
assign n_18453 =  x_658 & ~n_18302;
assign n_18454 =  i_7 &  n_18302;
assign n_18455 = ~n_18453 & ~n_18454;
assign n_18456 =  x_658 & ~n_18455;
assign n_18457 = ~x_658 &  n_18455;
assign n_18458 = ~n_18456 & ~n_18457;
assign n_18459 =  x_657 & ~n_18302;
assign n_18460 =  i_6 &  n_18302;
assign n_18461 = ~n_18459 & ~n_18460;
assign n_18462 =  x_657 & ~n_18461;
assign n_18463 = ~x_657 &  n_18461;
assign n_18464 = ~n_18462 & ~n_18463;
assign n_18465 =  x_656 & ~n_18302;
assign n_18466 =  i_5 &  n_18302;
assign n_18467 = ~n_18465 & ~n_18466;
assign n_18468 =  x_656 & ~n_18467;
assign n_18469 = ~x_656 &  n_18467;
assign n_18470 = ~n_18468 & ~n_18469;
assign n_18471 =  x_655 & ~n_18302;
assign n_18472 =  i_4 &  n_18302;
assign n_18473 = ~n_18471 & ~n_18472;
assign n_18474 =  x_655 & ~n_18473;
assign n_18475 = ~x_655 &  n_18473;
assign n_18476 = ~n_18474 & ~n_18475;
assign n_18477 =  x_654 & ~n_18302;
assign n_18478 =  i_3 &  n_18302;
assign n_18479 = ~n_18477 & ~n_18478;
assign n_18480 =  x_654 & ~n_18479;
assign n_18481 = ~x_654 &  n_18479;
assign n_18482 = ~n_18480 & ~n_18481;
assign n_18483 =  x_653 & ~n_18302;
assign n_18484 =  i_2 &  n_18302;
assign n_18485 = ~n_18483 & ~n_18484;
assign n_18486 =  x_653 & ~n_18485;
assign n_18487 = ~x_653 &  n_18485;
assign n_18488 = ~n_18486 & ~n_18487;
assign n_18489 =  x_652 & ~n_18302;
assign n_18490 =  i_1 &  n_18302;
assign n_18491 = ~n_18489 & ~n_18490;
assign n_18492 =  x_652 & ~n_18491;
assign n_18493 = ~x_652 &  n_18491;
assign n_18494 = ~n_18492 & ~n_18493;
assign n_18495 =  n_2 &  n_1043;
assign n_18496 =  x_651 & ~n_18495;
assign n_18497 =  x_651 &  n_18496;
assign n_18498 = ~x_651 & ~n_18496;
assign n_18499 = ~n_18497 & ~n_18498;
assign n_18500 =  x_650 & ~n_18495;
assign n_18501 =  x_650 &  n_18500;
assign n_18502 = ~x_650 & ~n_18500;
assign n_18503 = ~n_18501 & ~n_18502;
assign n_18504 =  x_649 & ~n_18495;
assign n_18505 =  x_649 &  n_18504;
assign n_18506 = ~x_649 & ~n_18504;
assign n_18507 = ~n_18505 & ~n_18506;
assign n_18508 =  x_648 & ~n_18495;
assign n_18509 =  x_648 &  n_18508;
assign n_18510 = ~x_648 & ~n_18508;
assign n_18511 = ~n_18509 & ~n_18510;
assign n_18512 =  x_647 & ~n_18495;
assign n_18513 =  x_647 &  n_18512;
assign n_18514 = ~x_647 & ~n_18512;
assign n_18515 = ~n_18513 & ~n_18514;
assign n_18516 =  x_646 & ~n_18495;
assign n_18517 =  x_646 &  n_18516;
assign n_18518 = ~x_646 & ~n_18516;
assign n_18519 = ~n_18517 & ~n_18518;
assign n_18520 =  x_645 & ~n_18495;
assign n_18521 =  x_645 &  n_18520;
assign n_18522 = ~x_645 & ~n_18520;
assign n_18523 = ~n_18521 & ~n_18522;
assign n_18524 =  x_644 & ~n_18495;
assign n_18525 =  x_644 &  n_18524;
assign n_18526 = ~x_644 & ~n_18524;
assign n_18527 = ~n_18525 & ~n_18526;
assign n_18528 =  x_643 & ~n_18495;
assign n_18529 =  x_643 &  n_18528;
assign n_18530 = ~x_643 & ~n_18528;
assign n_18531 = ~n_18529 & ~n_18530;
assign n_18532 =  x_642 & ~n_18495;
assign n_18533 =  x_642 &  n_18532;
assign n_18534 = ~x_642 & ~n_18532;
assign n_18535 = ~n_18533 & ~n_18534;
assign n_18536 =  x_641 & ~n_18495;
assign n_18537 =  x_641 &  n_18536;
assign n_18538 = ~x_641 & ~n_18536;
assign n_18539 = ~n_18537 & ~n_18538;
assign n_18540 =  x_640 & ~n_18495;
assign n_18541 =  x_640 &  n_18540;
assign n_18542 = ~x_640 & ~n_18540;
assign n_18543 = ~n_18541 & ~n_18542;
assign n_18544 =  x_639 & ~n_18495;
assign n_18545 =  x_639 &  n_18544;
assign n_18546 = ~x_639 & ~n_18544;
assign n_18547 = ~n_18545 & ~n_18546;
assign n_18548 =  x_638 & ~n_18495;
assign n_18549 =  x_638 &  n_18548;
assign n_18550 = ~x_638 & ~n_18548;
assign n_18551 = ~n_18549 & ~n_18550;
assign n_18552 =  x_637 & ~n_18495;
assign n_18553 =  x_637 &  n_18552;
assign n_18554 = ~x_637 & ~n_18552;
assign n_18555 = ~n_18553 & ~n_18554;
assign n_18556 =  x_636 & ~n_18495;
assign n_18557 =  x_636 &  n_18556;
assign n_18558 = ~x_636 & ~n_18556;
assign n_18559 = ~n_18557 & ~n_18558;
assign n_18560 =  x_635 & ~n_18495;
assign n_18561 =  x_635 &  n_18560;
assign n_18562 = ~x_635 & ~n_18560;
assign n_18563 = ~n_18561 & ~n_18562;
assign n_18564 =  x_634 & ~n_18495;
assign n_18565 =  x_634 &  n_18564;
assign n_18566 = ~x_634 & ~n_18564;
assign n_18567 = ~n_18565 & ~n_18566;
assign n_18568 =  x_633 & ~n_18495;
assign n_18569 =  x_633 &  n_18568;
assign n_18570 = ~x_633 & ~n_18568;
assign n_18571 = ~n_18569 & ~n_18570;
assign n_18572 =  x_632 & ~n_18495;
assign n_18573 =  x_632 &  n_18572;
assign n_18574 = ~x_632 & ~n_18572;
assign n_18575 = ~n_18573 & ~n_18574;
assign n_18576 =  x_631 & ~n_18495;
assign n_18577 =  x_631 &  n_18576;
assign n_18578 = ~x_631 & ~n_18576;
assign n_18579 = ~n_18577 & ~n_18578;
assign n_18580 =  x_630 & ~n_18495;
assign n_18581 =  x_630 &  n_18580;
assign n_18582 = ~x_630 & ~n_18580;
assign n_18583 = ~n_18581 & ~n_18582;
assign n_18584 =  x_629 & ~n_18495;
assign n_18585 =  x_629 &  n_18584;
assign n_18586 = ~x_629 & ~n_18584;
assign n_18587 = ~n_18585 & ~n_18586;
assign n_18588 =  x_628 & ~n_18495;
assign n_18589 =  x_628 &  n_18588;
assign n_18590 = ~x_628 & ~n_18588;
assign n_18591 = ~n_18589 & ~n_18590;
assign n_18592 =  x_627 & ~n_18495;
assign n_18593 =  x_627 &  n_18592;
assign n_18594 = ~x_627 & ~n_18592;
assign n_18595 = ~n_18593 & ~n_18594;
assign n_18596 =  x_626 & ~n_18495;
assign n_18597 =  x_626 &  n_18596;
assign n_18598 = ~x_626 & ~n_18596;
assign n_18599 = ~n_18597 & ~n_18598;
assign n_18600 =  x_625 & ~n_18495;
assign n_18601 =  x_625 &  n_18600;
assign n_18602 = ~x_625 & ~n_18600;
assign n_18603 = ~n_18601 & ~n_18602;
assign n_18604 =  x_624 & ~n_18495;
assign n_18605 =  x_624 &  n_18604;
assign n_18606 = ~x_624 & ~n_18604;
assign n_18607 = ~n_18605 & ~n_18606;
assign n_18608 =  x_623 & ~n_18495;
assign n_18609 =  x_623 &  n_18608;
assign n_18610 = ~x_623 & ~n_18608;
assign n_18611 = ~n_18609 & ~n_18610;
assign n_18612 =  x_622 & ~n_18495;
assign n_18613 =  x_622 &  n_18612;
assign n_18614 = ~x_622 & ~n_18612;
assign n_18615 = ~n_18613 & ~n_18614;
assign n_18616 =  x_621 & ~n_18495;
assign n_18617 =  x_621 &  n_18616;
assign n_18618 = ~x_621 & ~n_18616;
assign n_18619 = ~n_18617 & ~n_18618;
assign n_18620 =  x_620 & ~n_18495;
assign n_18621 =  x_620 &  n_18620;
assign n_18622 = ~x_620 & ~n_18620;
assign n_18623 = ~n_18621 & ~n_18622;
assign n_18624 =  n_1896 &  n_13104;
assign n_18625 =  n_552 &  n_18624;
assign n_18626 =  x_619 & ~n_18625;
assign n_18627 =  x_619 &  n_18626;
assign n_18628 = ~x_619 & ~n_18626;
assign n_18629 = ~n_18627 & ~n_18628;
assign n_18630 =  x_618 & ~n_18625;
assign n_18631 =  x_618 &  n_18630;
assign n_18632 = ~x_618 & ~n_18630;
assign n_18633 = ~n_18631 & ~n_18632;
assign n_18634 =  x_617 & ~n_18625;
assign n_18635 =  x_617 &  n_18634;
assign n_18636 = ~x_617 & ~n_18634;
assign n_18637 = ~n_18635 & ~n_18636;
assign n_18638 =  x_616 & ~n_18625;
assign n_18639 =  x_616 &  n_18638;
assign n_18640 = ~x_616 & ~n_18638;
assign n_18641 = ~n_18639 & ~n_18640;
assign n_18642 =  x_615 & ~n_18625;
assign n_18643 =  x_615 &  n_18642;
assign n_18644 = ~x_615 & ~n_18642;
assign n_18645 = ~n_18643 & ~n_18644;
assign n_18646 =  x_614 & ~n_18625;
assign n_18647 =  x_614 &  n_18646;
assign n_18648 = ~x_614 & ~n_18646;
assign n_18649 = ~n_18647 & ~n_18648;
assign n_18650 =  x_613 & ~n_18625;
assign n_18651 =  x_613 &  n_18650;
assign n_18652 = ~x_613 & ~n_18650;
assign n_18653 = ~n_18651 & ~n_18652;
assign n_18654 =  x_612 & ~n_18625;
assign n_18655 =  x_612 &  n_18654;
assign n_18656 = ~x_612 & ~n_18654;
assign n_18657 = ~n_18655 & ~n_18656;
assign n_18658 =  x_611 & ~n_18625;
assign n_18659 =  x_611 &  n_18658;
assign n_18660 = ~x_611 & ~n_18658;
assign n_18661 = ~n_18659 & ~n_18660;
assign n_18662 =  x_610 & ~n_18625;
assign n_18663 =  x_610 &  n_18662;
assign n_18664 = ~x_610 & ~n_18662;
assign n_18665 = ~n_18663 & ~n_18664;
assign n_18666 =  x_609 & ~n_18625;
assign n_18667 =  x_609 &  n_18666;
assign n_18668 = ~x_609 & ~n_18666;
assign n_18669 = ~n_18667 & ~n_18668;
assign n_18670 =  x_608 & ~n_18625;
assign n_18671 =  x_608 &  n_18670;
assign n_18672 = ~x_608 & ~n_18670;
assign n_18673 = ~n_18671 & ~n_18672;
assign n_18674 =  x_607 & ~n_18625;
assign n_18675 =  x_607 &  n_18674;
assign n_18676 = ~x_607 & ~n_18674;
assign n_18677 = ~n_18675 & ~n_18676;
assign n_18678 =  x_606 & ~n_18625;
assign n_18679 =  x_606 &  n_18678;
assign n_18680 = ~x_606 & ~n_18678;
assign n_18681 = ~n_18679 & ~n_18680;
assign n_18682 =  x_605 & ~n_18625;
assign n_18683 =  x_605 &  n_18682;
assign n_18684 = ~x_605 & ~n_18682;
assign n_18685 = ~n_18683 & ~n_18684;
assign n_18686 =  x_604 & ~n_18625;
assign n_18687 =  x_604 &  n_18686;
assign n_18688 = ~x_604 & ~n_18686;
assign n_18689 = ~n_18687 & ~n_18688;
assign n_18690 =  x_603 & ~n_18625;
assign n_18691 =  x_603 &  n_18690;
assign n_18692 = ~x_603 & ~n_18690;
assign n_18693 = ~n_18691 & ~n_18692;
assign n_18694 =  x_602 & ~n_18625;
assign n_18695 =  x_602 &  n_18694;
assign n_18696 = ~x_602 & ~n_18694;
assign n_18697 = ~n_18695 & ~n_18696;
assign n_18698 =  x_601 & ~n_18625;
assign n_18699 =  x_601 &  n_18698;
assign n_18700 = ~x_601 & ~n_18698;
assign n_18701 = ~n_18699 & ~n_18700;
assign n_18702 =  x_600 & ~n_18625;
assign n_18703 =  x_600 &  n_18702;
assign n_18704 = ~x_600 & ~n_18702;
assign n_18705 = ~n_18703 & ~n_18704;
assign n_18706 =  x_599 & ~n_18625;
assign n_18707 =  x_599 &  n_18706;
assign n_18708 = ~x_599 & ~n_18706;
assign n_18709 = ~n_18707 & ~n_18708;
assign n_18710 =  x_598 & ~n_18625;
assign n_18711 =  x_598 &  n_18710;
assign n_18712 = ~x_598 & ~n_18710;
assign n_18713 = ~n_18711 & ~n_18712;
assign n_18714 =  x_597 & ~n_18625;
assign n_18715 =  x_597 &  n_18714;
assign n_18716 = ~x_597 & ~n_18714;
assign n_18717 = ~n_18715 & ~n_18716;
assign n_18718 =  x_596 & ~n_18625;
assign n_18719 =  x_596 &  n_18718;
assign n_18720 = ~x_596 & ~n_18718;
assign n_18721 = ~n_18719 & ~n_18720;
assign n_18722 =  x_595 & ~n_18625;
assign n_18723 =  x_595 &  n_18722;
assign n_18724 = ~x_595 & ~n_18722;
assign n_18725 = ~n_18723 & ~n_18724;
assign n_18726 =  x_594 & ~n_18625;
assign n_18727 =  x_594 &  n_18726;
assign n_18728 = ~x_594 & ~n_18726;
assign n_18729 = ~n_18727 & ~n_18728;
assign n_18730 =  x_593 & ~n_18625;
assign n_18731 =  x_593 &  n_18730;
assign n_18732 = ~x_593 & ~n_18730;
assign n_18733 = ~n_18731 & ~n_18732;
assign n_18734 =  x_592 & ~n_18625;
assign n_18735 =  x_592 &  n_18734;
assign n_18736 = ~x_592 & ~n_18734;
assign n_18737 = ~n_18735 & ~n_18736;
assign n_18738 =  x_591 & ~n_18625;
assign n_18739 =  x_591 &  n_18738;
assign n_18740 = ~x_591 & ~n_18738;
assign n_18741 = ~n_18739 & ~n_18740;
assign n_18742 =  x_590 & ~n_18625;
assign n_18743 =  x_590 &  n_18742;
assign n_18744 = ~x_590 & ~n_18742;
assign n_18745 = ~n_18743 & ~n_18744;
assign n_18746 =  x_589 & ~n_18625;
assign n_18747 =  x_589 &  n_18746;
assign n_18748 = ~x_589 & ~n_18746;
assign n_18749 = ~n_18747 & ~n_18748;
assign n_18750 =  x_588 & ~n_18625;
assign n_18751 =  x_588 &  n_18750;
assign n_18752 = ~x_588 & ~n_18750;
assign n_18753 = ~n_18751 & ~n_18752;
assign n_18754 =  x_587 & ~n_7274;
assign n_18755 = ~n_18754 & ~n_7275;
assign n_18756 =  x_587 & ~n_18755;
assign n_18757 = ~x_587 &  n_18755;
assign n_18758 = ~n_18756 & ~n_18757;
assign n_18759 =  x_586 & ~n_7274;
assign n_18760 = ~n_18759 & ~n_7281;
assign n_18761 =  x_586 & ~n_18760;
assign n_18762 = ~x_586 &  n_18760;
assign n_18763 = ~n_18761 & ~n_18762;
assign n_18764 =  x_585 & ~n_7274;
assign n_18765 = ~n_18764 & ~n_7287;
assign n_18766 =  x_585 & ~n_18765;
assign n_18767 = ~x_585 &  n_18765;
assign n_18768 = ~n_18766 & ~n_18767;
assign n_18769 =  x_584 & ~n_7274;
assign n_18770 = ~n_18769 & ~n_7293;
assign n_18771 =  x_584 & ~n_18770;
assign n_18772 = ~x_584 &  n_18770;
assign n_18773 = ~n_18771 & ~n_18772;
assign n_18774 =  x_583 & ~n_7274;
assign n_18775 = ~n_18774 & ~n_7299;
assign n_18776 =  x_583 & ~n_18775;
assign n_18777 = ~x_583 &  n_18775;
assign n_18778 = ~n_18776 & ~n_18777;
assign n_18779 =  x_582 & ~n_7274;
assign n_18780 = ~n_18779 & ~n_7305;
assign n_18781 =  x_582 & ~n_18780;
assign n_18782 = ~x_582 &  n_18780;
assign n_18783 = ~n_18781 & ~n_18782;
assign n_18784 =  x_581 & ~n_7274;
assign n_18785 = ~n_18784 & ~n_7311;
assign n_18786 =  x_581 & ~n_18785;
assign n_18787 = ~x_581 &  n_18785;
assign n_18788 = ~n_18786 & ~n_18787;
assign n_18789 =  x_580 & ~n_7274;
assign n_18790 = ~n_18789 & ~n_7317;
assign n_18791 =  x_580 & ~n_18790;
assign n_18792 = ~x_580 &  n_18790;
assign n_18793 = ~n_18791 & ~n_18792;
assign n_18794 =  x_579 & ~n_7274;
assign n_18795 = ~n_18794 & ~n_7323;
assign n_18796 =  x_579 & ~n_18795;
assign n_18797 = ~x_579 &  n_18795;
assign n_18798 = ~n_18796 & ~n_18797;
assign n_18799 =  x_578 & ~n_7274;
assign n_18800 = ~n_18799 & ~n_7329;
assign n_18801 =  x_578 & ~n_18800;
assign n_18802 = ~x_578 &  n_18800;
assign n_18803 = ~n_18801 & ~n_18802;
assign n_18804 =  x_577 & ~n_7274;
assign n_18805 = ~n_18804 & ~n_7335;
assign n_18806 =  x_577 & ~n_18805;
assign n_18807 = ~x_577 &  n_18805;
assign n_18808 = ~n_18806 & ~n_18807;
assign n_18809 =  x_576 & ~n_7274;
assign n_18810 = ~n_18809 & ~n_7341;
assign n_18811 =  x_576 & ~n_18810;
assign n_18812 = ~x_576 &  n_18810;
assign n_18813 = ~n_18811 & ~n_18812;
assign n_18814 =  x_575 & ~n_7274;
assign n_18815 = ~n_18814 & ~n_7347;
assign n_18816 =  x_575 & ~n_18815;
assign n_18817 = ~x_575 &  n_18815;
assign n_18818 = ~n_18816 & ~n_18817;
assign n_18819 =  x_574 & ~n_7274;
assign n_18820 = ~n_18819 & ~n_7353;
assign n_18821 =  x_574 & ~n_18820;
assign n_18822 = ~x_574 &  n_18820;
assign n_18823 = ~n_18821 & ~n_18822;
assign n_18824 =  x_573 & ~n_7274;
assign n_18825 = ~n_18824 & ~n_7359;
assign n_18826 =  x_573 & ~n_18825;
assign n_18827 = ~x_573 &  n_18825;
assign n_18828 = ~n_18826 & ~n_18827;
assign n_18829 =  x_572 & ~n_7274;
assign n_18830 = ~n_18829 & ~n_7365;
assign n_18831 =  x_572 & ~n_18830;
assign n_18832 = ~x_572 &  n_18830;
assign n_18833 = ~n_18831 & ~n_18832;
assign n_18834 =  x_571 & ~n_7274;
assign n_18835 = ~n_18834 & ~n_7371;
assign n_18836 =  x_571 & ~n_18835;
assign n_18837 = ~x_571 &  n_18835;
assign n_18838 = ~n_18836 & ~n_18837;
assign n_18839 =  x_570 & ~n_7274;
assign n_18840 = ~n_18839 & ~n_7377;
assign n_18841 =  x_570 & ~n_18840;
assign n_18842 = ~x_570 &  n_18840;
assign n_18843 = ~n_18841 & ~n_18842;
assign n_18844 =  x_569 & ~n_7274;
assign n_18845 = ~n_18844 & ~n_7383;
assign n_18846 =  x_569 & ~n_18845;
assign n_18847 = ~x_569 &  n_18845;
assign n_18848 = ~n_18846 & ~n_18847;
assign n_18849 =  x_568 & ~n_7274;
assign n_18850 = ~n_18849 & ~n_7389;
assign n_18851 =  x_568 & ~n_18850;
assign n_18852 = ~x_568 &  n_18850;
assign n_18853 = ~n_18851 & ~n_18852;
assign n_18854 =  x_567 & ~n_7274;
assign n_18855 = ~n_18854 & ~n_7395;
assign n_18856 =  x_567 & ~n_18855;
assign n_18857 = ~x_567 &  n_18855;
assign n_18858 = ~n_18856 & ~n_18857;
assign n_18859 =  x_566 & ~n_7274;
assign n_18860 = ~n_18859 & ~n_7401;
assign n_18861 =  x_566 & ~n_18860;
assign n_18862 = ~x_566 &  n_18860;
assign n_18863 = ~n_18861 & ~n_18862;
assign n_18864 =  x_565 & ~n_7274;
assign n_18865 = ~n_18864 & ~n_7407;
assign n_18866 =  x_565 & ~n_18865;
assign n_18867 = ~x_565 &  n_18865;
assign n_18868 = ~n_18866 & ~n_18867;
assign n_18869 =  x_564 & ~n_7274;
assign n_18870 = ~n_18869 & ~n_7413;
assign n_18871 =  x_564 & ~n_18870;
assign n_18872 = ~x_564 &  n_18870;
assign n_18873 = ~n_18871 & ~n_18872;
assign n_18874 =  x_563 & ~n_7274;
assign n_18875 = ~n_18874 & ~n_7419;
assign n_18876 =  x_563 & ~n_18875;
assign n_18877 = ~x_563 &  n_18875;
assign n_18878 = ~n_18876 & ~n_18877;
assign n_18879 =  x_562 & ~n_7274;
assign n_18880 = ~n_18879 & ~n_7425;
assign n_18881 =  x_562 & ~n_18880;
assign n_18882 = ~x_562 &  n_18880;
assign n_18883 = ~n_18881 & ~n_18882;
assign n_18884 =  x_561 & ~n_7274;
assign n_18885 = ~n_18884 & ~n_7431;
assign n_18886 =  x_561 & ~n_18885;
assign n_18887 = ~x_561 &  n_18885;
assign n_18888 = ~n_18886 & ~n_18887;
assign n_18889 =  x_560 & ~n_7274;
assign n_18890 = ~n_18889 & ~n_7437;
assign n_18891 =  x_560 & ~n_18890;
assign n_18892 = ~x_560 &  n_18890;
assign n_18893 = ~n_18891 & ~n_18892;
assign n_18894 =  x_559 & ~n_7274;
assign n_18895 = ~n_18894 & ~n_7443;
assign n_18896 =  x_559 & ~n_18895;
assign n_18897 = ~x_559 &  n_18895;
assign n_18898 = ~n_18896 & ~n_18897;
assign n_18899 =  x_558 & ~n_7274;
assign n_18900 = ~n_18899 & ~n_7449;
assign n_18901 =  x_558 & ~n_18900;
assign n_18902 = ~x_558 &  n_18900;
assign n_18903 = ~n_18901 & ~n_18902;
assign n_18904 =  x_557 & ~n_7274;
assign n_18905 = ~n_18904 & ~n_7455;
assign n_18906 =  x_557 & ~n_18905;
assign n_18907 = ~x_557 &  n_18905;
assign n_18908 = ~n_18906 & ~n_18907;
assign n_18909 =  x_556 & ~n_7274;
assign n_18910 = ~n_18909 & ~n_7461;
assign n_18911 =  x_556 & ~n_18910;
assign n_18912 = ~x_556 &  n_18910;
assign n_18913 = ~n_18911 & ~n_18912;
assign n_18914 =  n_2095 &  n_1896;
assign n_18915 =  n_8344 &  n_18914;
assign n_18916 =  x_555 & ~n_18915;
assign n_18917 =  i_32 &  n_18915;
assign n_18918 = ~n_18916 & ~n_18917;
assign n_18919 =  x_555 & ~n_18918;
assign n_18920 = ~x_555 &  n_18918;
assign n_18921 = ~n_18919 & ~n_18920;
assign n_18922 =  x_554 & ~n_18915;
assign n_18923 =  i_31 &  n_18915;
assign n_18924 = ~n_18922 & ~n_18923;
assign n_18925 =  x_554 & ~n_18924;
assign n_18926 = ~x_554 &  n_18924;
assign n_18927 = ~n_18925 & ~n_18926;
assign n_18928 =  x_553 & ~n_18915;
assign n_18929 =  i_30 &  n_18915;
assign n_18930 = ~n_18928 & ~n_18929;
assign n_18931 =  x_553 & ~n_18930;
assign n_18932 = ~x_553 &  n_18930;
assign n_18933 = ~n_18931 & ~n_18932;
assign n_18934 =  x_552 & ~n_18915;
assign n_18935 =  i_29 &  n_18915;
assign n_18936 = ~n_18934 & ~n_18935;
assign n_18937 =  x_552 & ~n_18936;
assign n_18938 = ~x_552 &  n_18936;
assign n_18939 = ~n_18937 & ~n_18938;
assign n_18940 =  x_551 & ~n_18915;
assign n_18941 =  i_28 &  n_18915;
assign n_18942 = ~n_18940 & ~n_18941;
assign n_18943 =  x_551 & ~n_18942;
assign n_18944 = ~x_551 &  n_18942;
assign n_18945 = ~n_18943 & ~n_18944;
assign n_18946 =  x_550 & ~n_18915;
assign n_18947 =  i_27 &  n_18915;
assign n_18948 = ~n_18946 & ~n_18947;
assign n_18949 =  x_550 & ~n_18948;
assign n_18950 = ~x_550 &  n_18948;
assign n_18951 = ~n_18949 & ~n_18950;
assign n_18952 =  x_549 & ~n_18915;
assign n_18953 =  i_26 &  n_18915;
assign n_18954 = ~n_18952 & ~n_18953;
assign n_18955 =  x_549 & ~n_18954;
assign n_18956 = ~x_549 &  n_18954;
assign n_18957 = ~n_18955 & ~n_18956;
assign n_18958 =  x_548 & ~n_18915;
assign n_18959 =  i_25 &  n_18915;
assign n_18960 = ~n_18958 & ~n_18959;
assign n_18961 =  x_548 & ~n_18960;
assign n_18962 = ~x_548 &  n_18960;
assign n_18963 = ~n_18961 & ~n_18962;
assign n_18964 =  x_547 & ~n_18915;
assign n_18965 =  i_24 &  n_18915;
assign n_18966 = ~n_18964 & ~n_18965;
assign n_18967 =  x_547 & ~n_18966;
assign n_18968 = ~x_547 &  n_18966;
assign n_18969 = ~n_18967 & ~n_18968;
assign n_18970 =  x_546 & ~n_18915;
assign n_18971 =  i_23 &  n_18915;
assign n_18972 = ~n_18970 & ~n_18971;
assign n_18973 =  x_546 & ~n_18972;
assign n_18974 = ~x_546 &  n_18972;
assign n_18975 = ~n_18973 & ~n_18974;
assign n_18976 =  x_545 & ~n_18915;
assign n_18977 =  i_22 &  n_18915;
assign n_18978 = ~n_18976 & ~n_18977;
assign n_18979 =  x_545 & ~n_18978;
assign n_18980 = ~x_545 &  n_18978;
assign n_18981 = ~n_18979 & ~n_18980;
assign n_18982 =  x_544 & ~n_18915;
assign n_18983 =  i_21 &  n_18915;
assign n_18984 = ~n_18982 & ~n_18983;
assign n_18985 =  x_544 & ~n_18984;
assign n_18986 = ~x_544 &  n_18984;
assign n_18987 = ~n_18985 & ~n_18986;
assign n_18988 =  x_543 & ~n_18915;
assign n_18989 =  i_20 &  n_18915;
assign n_18990 = ~n_18988 & ~n_18989;
assign n_18991 =  x_543 & ~n_18990;
assign n_18992 = ~x_543 &  n_18990;
assign n_18993 = ~n_18991 & ~n_18992;
assign n_18994 =  x_542 & ~n_18915;
assign n_18995 =  i_19 &  n_18915;
assign n_18996 = ~n_18994 & ~n_18995;
assign n_18997 =  x_542 & ~n_18996;
assign n_18998 = ~x_542 &  n_18996;
assign n_18999 = ~n_18997 & ~n_18998;
assign n_19000 =  x_541 & ~n_18915;
assign n_19001 =  i_18 &  n_18915;
assign n_19002 = ~n_19000 & ~n_19001;
assign n_19003 =  x_541 & ~n_19002;
assign n_19004 = ~x_541 &  n_19002;
assign n_19005 = ~n_19003 & ~n_19004;
assign n_19006 =  x_540 & ~n_18915;
assign n_19007 =  i_17 &  n_18915;
assign n_19008 = ~n_19006 & ~n_19007;
assign n_19009 =  x_540 & ~n_19008;
assign n_19010 = ~x_540 &  n_19008;
assign n_19011 = ~n_19009 & ~n_19010;
assign n_19012 =  x_539 & ~n_18915;
assign n_19013 =  i_16 &  n_18915;
assign n_19014 = ~n_19012 & ~n_19013;
assign n_19015 =  x_539 & ~n_19014;
assign n_19016 = ~x_539 &  n_19014;
assign n_19017 = ~n_19015 & ~n_19016;
assign n_19018 =  x_538 & ~n_18915;
assign n_19019 =  i_15 &  n_18915;
assign n_19020 = ~n_19018 & ~n_19019;
assign n_19021 =  x_538 & ~n_19020;
assign n_19022 = ~x_538 &  n_19020;
assign n_19023 = ~n_19021 & ~n_19022;
assign n_19024 =  x_537 & ~n_18915;
assign n_19025 =  i_14 &  n_18915;
assign n_19026 = ~n_19024 & ~n_19025;
assign n_19027 =  x_537 & ~n_19026;
assign n_19028 = ~x_537 &  n_19026;
assign n_19029 = ~n_19027 & ~n_19028;
assign n_19030 =  x_536 & ~n_18915;
assign n_19031 =  i_13 &  n_18915;
assign n_19032 = ~n_19030 & ~n_19031;
assign n_19033 =  x_536 & ~n_19032;
assign n_19034 = ~x_536 &  n_19032;
assign n_19035 = ~n_19033 & ~n_19034;
assign n_19036 =  x_535 & ~n_18915;
assign n_19037 =  i_12 &  n_18915;
assign n_19038 = ~n_19036 & ~n_19037;
assign n_19039 =  x_535 & ~n_19038;
assign n_19040 = ~x_535 &  n_19038;
assign n_19041 = ~n_19039 & ~n_19040;
assign n_19042 =  x_534 & ~n_18915;
assign n_19043 =  i_11 &  n_18915;
assign n_19044 = ~n_19042 & ~n_19043;
assign n_19045 =  x_534 & ~n_19044;
assign n_19046 = ~x_534 &  n_19044;
assign n_19047 = ~n_19045 & ~n_19046;
assign n_19048 =  x_533 & ~n_18915;
assign n_19049 =  i_10 &  n_18915;
assign n_19050 = ~n_19048 & ~n_19049;
assign n_19051 =  x_533 & ~n_19050;
assign n_19052 = ~x_533 &  n_19050;
assign n_19053 = ~n_19051 & ~n_19052;
assign n_19054 =  x_532 & ~n_18915;
assign n_19055 =  i_9 &  n_18915;
assign n_19056 = ~n_19054 & ~n_19055;
assign n_19057 =  x_532 & ~n_19056;
assign n_19058 = ~x_532 &  n_19056;
assign n_19059 = ~n_19057 & ~n_19058;
assign n_19060 =  x_531 & ~n_18915;
assign n_19061 =  i_8 &  n_18915;
assign n_19062 = ~n_19060 & ~n_19061;
assign n_19063 =  x_531 & ~n_19062;
assign n_19064 = ~x_531 &  n_19062;
assign n_19065 = ~n_19063 & ~n_19064;
assign n_19066 =  x_530 & ~n_18915;
assign n_19067 =  i_7 &  n_18915;
assign n_19068 = ~n_19066 & ~n_19067;
assign n_19069 =  x_530 & ~n_19068;
assign n_19070 = ~x_530 &  n_19068;
assign n_19071 = ~n_19069 & ~n_19070;
assign n_19072 =  x_529 & ~n_18915;
assign n_19073 =  i_6 &  n_18915;
assign n_19074 = ~n_19072 & ~n_19073;
assign n_19075 =  x_529 & ~n_19074;
assign n_19076 = ~x_529 &  n_19074;
assign n_19077 = ~n_19075 & ~n_19076;
assign n_19078 =  x_528 & ~n_18915;
assign n_19079 =  i_5 &  n_18915;
assign n_19080 = ~n_19078 & ~n_19079;
assign n_19081 =  x_528 & ~n_19080;
assign n_19082 = ~x_528 &  n_19080;
assign n_19083 = ~n_19081 & ~n_19082;
assign n_19084 =  x_527 & ~n_18915;
assign n_19085 =  i_4 &  n_18915;
assign n_19086 = ~n_19084 & ~n_19085;
assign n_19087 =  x_527 & ~n_19086;
assign n_19088 = ~x_527 &  n_19086;
assign n_19089 = ~n_19087 & ~n_19088;
assign n_19090 =  x_526 & ~n_18915;
assign n_19091 =  i_3 &  n_18915;
assign n_19092 = ~n_19090 & ~n_19091;
assign n_19093 =  x_526 & ~n_19092;
assign n_19094 = ~x_526 &  n_19092;
assign n_19095 = ~n_19093 & ~n_19094;
assign n_19096 =  x_525 & ~n_18915;
assign n_19097 =  i_2 &  n_18915;
assign n_19098 = ~n_19096 & ~n_19097;
assign n_19099 =  x_525 & ~n_19098;
assign n_19100 = ~x_525 &  n_19098;
assign n_19101 = ~n_19099 & ~n_19100;
assign n_19102 =  x_524 & ~n_18915;
assign n_19103 =  i_1 &  n_18915;
assign n_19104 = ~n_19102 & ~n_19103;
assign n_19105 =  x_524 & ~n_19104;
assign n_19106 = ~x_524 &  n_19104;
assign n_19107 = ~n_19105 & ~n_19106;
assign n_19108 =  n_555 &  n_13872;
assign n_19109 =  x_523 & ~n_19108;
assign n_19110 =  i_32 &  n_19108;
assign n_19111 = ~n_19109 & ~n_19110;
assign n_19112 =  x_523 & ~n_19111;
assign n_19113 = ~x_523 &  n_19111;
assign n_19114 = ~n_19112 & ~n_19113;
assign n_19115 =  x_522 & ~n_19108;
assign n_19116 =  i_31 &  n_19108;
assign n_19117 = ~n_19115 & ~n_19116;
assign n_19118 =  x_522 & ~n_19117;
assign n_19119 = ~x_522 &  n_19117;
assign n_19120 = ~n_19118 & ~n_19119;
assign n_19121 =  x_521 & ~n_19108;
assign n_19122 =  i_30 &  n_19108;
assign n_19123 = ~n_19121 & ~n_19122;
assign n_19124 =  x_521 & ~n_19123;
assign n_19125 = ~x_521 &  n_19123;
assign n_19126 = ~n_19124 & ~n_19125;
assign n_19127 =  x_520 & ~n_19108;
assign n_19128 =  i_29 &  n_19108;
assign n_19129 = ~n_19127 & ~n_19128;
assign n_19130 =  x_520 & ~n_19129;
assign n_19131 = ~x_520 &  n_19129;
assign n_19132 = ~n_19130 & ~n_19131;
assign n_19133 =  x_519 & ~n_19108;
assign n_19134 =  i_28 &  n_19108;
assign n_19135 = ~n_19133 & ~n_19134;
assign n_19136 =  x_519 & ~n_19135;
assign n_19137 = ~x_519 &  n_19135;
assign n_19138 = ~n_19136 & ~n_19137;
assign n_19139 =  x_518 & ~n_19108;
assign n_19140 =  i_27 &  n_19108;
assign n_19141 = ~n_19139 & ~n_19140;
assign n_19142 =  x_518 & ~n_19141;
assign n_19143 = ~x_518 &  n_19141;
assign n_19144 = ~n_19142 & ~n_19143;
assign n_19145 =  x_517 & ~n_19108;
assign n_19146 =  i_26 &  n_19108;
assign n_19147 = ~n_19145 & ~n_19146;
assign n_19148 =  x_517 & ~n_19147;
assign n_19149 = ~x_517 &  n_19147;
assign n_19150 = ~n_19148 & ~n_19149;
assign n_19151 =  x_516 & ~n_19108;
assign n_19152 =  i_25 &  n_19108;
assign n_19153 = ~n_19151 & ~n_19152;
assign n_19154 =  x_516 & ~n_19153;
assign n_19155 = ~x_516 &  n_19153;
assign n_19156 = ~n_19154 & ~n_19155;
assign n_19157 =  x_515 & ~n_19108;
assign n_19158 =  i_24 &  n_19108;
assign n_19159 = ~n_19157 & ~n_19158;
assign n_19160 =  x_515 & ~n_19159;
assign n_19161 = ~x_515 &  n_19159;
assign n_19162 = ~n_19160 & ~n_19161;
assign n_19163 =  x_514 & ~n_19108;
assign n_19164 =  i_23 &  n_19108;
assign n_19165 = ~n_19163 & ~n_19164;
assign n_19166 =  x_514 & ~n_19165;
assign n_19167 = ~x_514 &  n_19165;
assign n_19168 = ~n_19166 & ~n_19167;
assign n_19169 =  x_513 & ~n_19108;
assign n_19170 =  i_22 &  n_19108;
assign n_19171 = ~n_19169 & ~n_19170;
assign n_19172 =  x_513 & ~n_19171;
assign n_19173 = ~x_513 &  n_19171;
assign n_19174 = ~n_19172 & ~n_19173;
assign n_19175 =  x_512 & ~n_19108;
assign n_19176 =  i_21 &  n_19108;
assign n_19177 = ~n_19175 & ~n_19176;
assign n_19178 =  x_512 & ~n_19177;
assign n_19179 = ~x_512 &  n_19177;
assign n_19180 = ~n_19178 & ~n_19179;
assign n_19181 =  x_511 & ~n_19108;
assign n_19182 =  i_20 &  n_19108;
assign n_19183 = ~n_19181 & ~n_19182;
assign n_19184 =  x_511 & ~n_19183;
assign n_19185 = ~x_511 &  n_19183;
assign n_19186 = ~n_19184 & ~n_19185;
assign n_19187 =  x_510 & ~n_19108;
assign n_19188 =  i_19 &  n_19108;
assign n_19189 = ~n_19187 & ~n_19188;
assign n_19190 =  x_510 & ~n_19189;
assign n_19191 = ~x_510 &  n_19189;
assign n_19192 = ~n_19190 & ~n_19191;
assign n_19193 =  x_509 & ~n_19108;
assign n_19194 =  i_18 &  n_19108;
assign n_19195 = ~n_19193 & ~n_19194;
assign n_19196 =  x_509 & ~n_19195;
assign n_19197 = ~x_509 &  n_19195;
assign n_19198 = ~n_19196 & ~n_19197;
assign n_19199 =  x_508 & ~n_19108;
assign n_19200 =  i_17 &  n_19108;
assign n_19201 = ~n_19199 & ~n_19200;
assign n_19202 =  x_508 & ~n_19201;
assign n_19203 = ~x_508 &  n_19201;
assign n_19204 = ~n_19202 & ~n_19203;
assign n_19205 =  x_507 & ~n_19108;
assign n_19206 =  i_16 &  n_19108;
assign n_19207 = ~n_19205 & ~n_19206;
assign n_19208 =  x_507 & ~n_19207;
assign n_19209 = ~x_507 &  n_19207;
assign n_19210 = ~n_19208 & ~n_19209;
assign n_19211 =  x_506 & ~n_19108;
assign n_19212 =  i_15 &  n_19108;
assign n_19213 = ~n_19211 & ~n_19212;
assign n_19214 =  x_506 & ~n_19213;
assign n_19215 = ~x_506 &  n_19213;
assign n_19216 = ~n_19214 & ~n_19215;
assign n_19217 =  x_505 & ~n_19108;
assign n_19218 =  i_14 &  n_19108;
assign n_19219 = ~n_19217 & ~n_19218;
assign n_19220 =  x_505 & ~n_19219;
assign n_19221 = ~x_505 &  n_19219;
assign n_19222 = ~n_19220 & ~n_19221;
assign n_19223 =  x_504 & ~n_19108;
assign n_19224 =  i_13 &  n_19108;
assign n_19225 = ~n_19223 & ~n_19224;
assign n_19226 =  x_504 & ~n_19225;
assign n_19227 = ~x_504 &  n_19225;
assign n_19228 = ~n_19226 & ~n_19227;
assign n_19229 =  x_503 & ~n_19108;
assign n_19230 =  i_12 &  n_19108;
assign n_19231 = ~n_19229 & ~n_19230;
assign n_19232 =  x_503 & ~n_19231;
assign n_19233 = ~x_503 &  n_19231;
assign n_19234 = ~n_19232 & ~n_19233;
assign n_19235 =  x_502 & ~n_19108;
assign n_19236 =  i_11 &  n_19108;
assign n_19237 = ~n_19235 & ~n_19236;
assign n_19238 =  x_502 & ~n_19237;
assign n_19239 = ~x_502 &  n_19237;
assign n_19240 = ~n_19238 & ~n_19239;
assign n_19241 =  x_501 & ~n_19108;
assign n_19242 =  i_10 &  n_19108;
assign n_19243 = ~n_19241 & ~n_19242;
assign n_19244 =  x_501 & ~n_19243;
assign n_19245 = ~x_501 &  n_19243;
assign n_19246 = ~n_19244 & ~n_19245;
assign n_19247 =  x_500 & ~n_19108;
assign n_19248 =  i_9 &  n_19108;
assign n_19249 = ~n_19247 & ~n_19248;
assign n_19250 =  x_500 & ~n_19249;
assign n_19251 = ~x_500 &  n_19249;
assign n_19252 = ~n_19250 & ~n_19251;
assign n_19253 =  x_499 & ~n_19108;
assign n_19254 =  i_8 &  n_19108;
assign n_19255 = ~n_19253 & ~n_19254;
assign n_19256 =  x_499 & ~n_19255;
assign n_19257 = ~x_499 &  n_19255;
assign n_19258 = ~n_19256 & ~n_19257;
assign n_19259 =  x_498 & ~n_19108;
assign n_19260 =  i_7 &  n_19108;
assign n_19261 = ~n_19259 & ~n_19260;
assign n_19262 =  x_498 & ~n_19261;
assign n_19263 = ~x_498 &  n_19261;
assign n_19264 = ~n_19262 & ~n_19263;
assign n_19265 =  x_497 & ~n_19108;
assign n_19266 =  i_6 &  n_19108;
assign n_19267 = ~n_19265 & ~n_19266;
assign n_19268 =  x_497 & ~n_19267;
assign n_19269 = ~x_497 &  n_19267;
assign n_19270 = ~n_19268 & ~n_19269;
assign n_19271 =  x_496 & ~n_19108;
assign n_19272 =  i_5 &  n_19108;
assign n_19273 = ~n_19271 & ~n_19272;
assign n_19274 =  x_496 & ~n_19273;
assign n_19275 = ~x_496 &  n_19273;
assign n_19276 = ~n_19274 & ~n_19275;
assign n_19277 =  x_495 & ~n_19108;
assign n_19278 =  i_4 &  n_19108;
assign n_19279 = ~n_19277 & ~n_19278;
assign n_19280 =  x_495 & ~n_19279;
assign n_19281 = ~x_495 &  n_19279;
assign n_19282 = ~n_19280 & ~n_19281;
assign n_19283 =  x_494 & ~n_19108;
assign n_19284 =  i_3 &  n_19108;
assign n_19285 = ~n_19283 & ~n_19284;
assign n_19286 =  x_494 & ~n_19285;
assign n_19287 = ~x_494 &  n_19285;
assign n_19288 = ~n_19286 & ~n_19287;
assign n_19289 =  x_493 & ~n_19108;
assign n_19290 =  i_2 &  n_19108;
assign n_19291 = ~n_19289 & ~n_19290;
assign n_19292 =  x_493 & ~n_19291;
assign n_19293 = ~x_493 &  n_19291;
assign n_19294 = ~n_19292 & ~n_19293;
assign n_19295 =  x_492 & ~n_19108;
assign n_19296 =  i_1 &  n_19108;
assign n_19297 = ~n_19295 & ~n_19296;
assign n_19298 =  x_492 & ~n_19297;
assign n_19299 = ~x_492 &  n_19297;
assign n_19300 = ~n_19298 & ~n_19299;
assign n_19301 =  x_491 & ~n_1701;
assign n_19302 =  x_2058 &  n_1701;
assign n_19303 = ~n_19301 & ~n_19302;
assign n_19304 =  x_491 & ~n_19303;
assign n_19305 = ~x_491 &  n_19303;
assign n_19306 = ~n_19304 & ~n_19305;
assign n_19307 =  x_490 & ~n_1701;
assign n_19308 =  x_2057 &  n_1701;
assign n_19309 = ~n_19307 & ~n_19308;
assign n_19310 =  x_490 & ~n_19309;
assign n_19311 = ~x_490 &  n_19309;
assign n_19312 = ~n_19310 & ~n_19311;
assign n_19313 =  x_489 & ~n_1701;
assign n_19314 =  x_2056 &  n_1701;
assign n_19315 = ~n_19313 & ~n_19314;
assign n_19316 =  x_489 & ~n_19315;
assign n_19317 = ~x_489 &  n_19315;
assign n_19318 = ~n_19316 & ~n_19317;
assign n_19319 =  x_488 & ~n_1701;
assign n_19320 =  x_2055 &  n_1701;
assign n_19321 = ~n_19319 & ~n_19320;
assign n_19322 =  x_488 & ~n_19321;
assign n_19323 = ~x_488 &  n_19321;
assign n_19324 = ~n_19322 & ~n_19323;
assign n_19325 =  x_487 & ~n_1701;
assign n_19326 =  x_2054 &  n_1701;
assign n_19327 = ~n_19325 & ~n_19326;
assign n_19328 =  x_487 & ~n_19327;
assign n_19329 = ~x_487 &  n_19327;
assign n_19330 = ~n_19328 & ~n_19329;
assign n_19331 =  x_486 & ~n_1701;
assign n_19332 =  x_2053 &  n_1701;
assign n_19333 = ~n_19331 & ~n_19332;
assign n_19334 =  x_486 & ~n_19333;
assign n_19335 = ~x_486 &  n_19333;
assign n_19336 = ~n_19334 & ~n_19335;
assign n_19337 =  x_485 & ~n_1701;
assign n_19338 =  x_2052 &  n_1701;
assign n_19339 = ~n_19337 & ~n_19338;
assign n_19340 =  x_485 & ~n_19339;
assign n_19341 = ~x_485 &  n_19339;
assign n_19342 = ~n_19340 & ~n_19341;
assign n_19343 =  x_484 & ~n_1701;
assign n_19344 =  x_2051 &  n_1701;
assign n_19345 = ~n_19343 & ~n_19344;
assign n_19346 =  x_484 & ~n_19345;
assign n_19347 = ~x_484 &  n_19345;
assign n_19348 = ~n_19346 & ~n_19347;
assign n_19349 =  x_483 & ~n_1701;
assign n_19350 =  x_2050 &  n_1701;
assign n_19351 = ~n_19349 & ~n_19350;
assign n_19352 =  x_483 & ~n_19351;
assign n_19353 = ~x_483 &  n_19351;
assign n_19354 = ~n_19352 & ~n_19353;
assign n_19355 =  x_482 & ~n_1701;
assign n_19356 =  x_2049 &  n_1701;
assign n_19357 = ~n_19355 & ~n_19356;
assign n_19358 =  x_482 & ~n_19357;
assign n_19359 = ~x_482 &  n_19357;
assign n_19360 = ~n_19358 & ~n_19359;
assign n_19361 =  x_481 & ~n_1701;
assign n_19362 =  x_2048 &  n_1701;
assign n_19363 = ~n_19361 & ~n_19362;
assign n_19364 =  x_481 & ~n_19363;
assign n_19365 = ~x_481 &  n_19363;
assign n_19366 = ~n_19364 & ~n_19365;
assign n_19367 =  x_480 & ~n_1701;
assign n_19368 =  x_2047 &  n_1701;
assign n_19369 = ~n_19367 & ~n_19368;
assign n_19370 =  x_480 & ~n_19369;
assign n_19371 = ~x_480 &  n_19369;
assign n_19372 = ~n_19370 & ~n_19371;
assign n_19373 =  x_479 & ~n_1701;
assign n_19374 =  x_2046 &  n_1701;
assign n_19375 = ~n_19373 & ~n_19374;
assign n_19376 =  x_479 & ~n_19375;
assign n_19377 = ~x_479 &  n_19375;
assign n_19378 = ~n_19376 & ~n_19377;
assign n_19379 =  x_478 & ~n_1701;
assign n_19380 =  x_2045 &  n_1701;
assign n_19381 = ~n_19379 & ~n_19380;
assign n_19382 =  x_478 & ~n_19381;
assign n_19383 = ~x_478 &  n_19381;
assign n_19384 = ~n_19382 & ~n_19383;
assign n_19385 =  x_477 & ~n_1701;
assign n_19386 =  x_2044 &  n_1701;
assign n_19387 = ~n_19385 & ~n_19386;
assign n_19388 =  x_477 & ~n_19387;
assign n_19389 = ~x_477 &  n_19387;
assign n_19390 = ~n_19388 & ~n_19389;
assign n_19391 =  x_476 & ~n_1701;
assign n_19392 =  x_2043 &  n_1701;
assign n_19393 = ~n_19391 & ~n_19392;
assign n_19394 =  x_476 & ~n_19393;
assign n_19395 = ~x_476 &  n_19393;
assign n_19396 = ~n_19394 & ~n_19395;
assign n_19397 =  x_475 & ~n_1701;
assign n_19398 =  x_2042 &  n_1701;
assign n_19399 = ~n_19397 & ~n_19398;
assign n_19400 =  x_475 & ~n_19399;
assign n_19401 = ~x_475 &  n_19399;
assign n_19402 = ~n_19400 & ~n_19401;
assign n_19403 =  x_474 & ~n_1701;
assign n_19404 =  x_2041 &  n_1701;
assign n_19405 = ~n_19403 & ~n_19404;
assign n_19406 =  x_474 & ~n_19405;
assign n_19407 = ~x_474 &  n_19405;
assign n_19408 = ~n_19406 & ~n_19407;
assign n_19409 =  x_473 & ~n_1701;
assign n_19410 =  x_2040 &  n_1701;
assign n_19411 = ~n_19409 & ~n_19410;
assign n_19412 =  x_473 & ~n_19411;
assign n_19413 = ~x_473 &  n_19411;
assign n_19414 = ~n_19412 & ~n_19413;
assign n_19415 =  x_472 & ~n_1701;
assign n_19416 =  x_2039 &  n_1701;
assign n_19417 = ~n_19415 & ~n_19416;
assign n_19418 =  x_472 & ~n_19417;
assign n_19419 = ~x_472 &  n_19417;
assign n_19420 = ~n_19418 & ~n_19419;
assign n_19421 =  x_471 & ~n_1701;
assign n_19422 =  x_2038 &  n_1701;
assign n_19423 = ~n_19421 & ~n_19422;
assign n_19424 =  x_471 & ~n_19423;
assign n_19425 = ~x_471 &  n_19423;
assign n_19426 = ~n_19424 & ~n_19425;
assign n_19427 =  x_470 & ~n_1701;
assign n_19428 =  x_2037 &  n_1701;
assign n_19429 = ~n_19427 & ~n_19428;
assign n_19430 =  x_470 & ~n_19429;
assign n_19431 = ~x_470 &  n_19429;
assign n_19432 = ~n_19430 & ~n_19431;
assign n_19433 =  x_469 & ~n_1701;
assign n_19434 =  x_2036 &  n_1701;
assign n_19435 = ~n_19433 & ~n_19434;
assign n_19436 =  x_469 & ~n_19435;
assign n_19437 = ~x_469 &  n_19435;
assign n_19438 = ~n_19436 & ~n_19437;
assign n_19439 =  x_468 & ~n_1701;
assign n_19440 =  x_2035 &  n_1701;
assign n_19441 = ~n_19439 & ~n_19440;
assign n_19442 =  x_468 & ~n_19441;
assign n_19443 = ~x_468 &  n_19441;
assign n_19444 = ~n_19442 & ~n_19443;
assign n_19445 =  x_467 & ~n_1701;
assign n_19446 =  x_2034 &  n_1701;
assign n_19447 = ~n_19445 & ~n_19446;
assign n_19448 =  x_467 & ~n_19447;
assign n_19449 = ~x_467 &  n_19447;
assign n_19450 = ~n_19448 & ~n_19449;
assign n_19451 =  x_466 & ~n_1701;
assign n_19452 =  x_2033 &  n_1701;
assign n_19453 = ~n_19451 & ~n_19452;
assign n_19454 =  x_466 & ~n_19453;
assign n_19455 = ~x_466 &  n_19453;
assign n_19456 = ~n_19454 & ~n_19455;
assign n_19457 =  x_465 & ~n_1701;
assign n_19458 =  x_2032 &  n_1701;
assign n_19459 = ~n_19457 & ~n_19458;
assign n_19460 =  x_465 & ~n_19459;
assign n_19461 = ~x_465 &  n_19459;
assign n_19462 = ~n_19460 & ~n_19461;
assign n_19463 =  x_464 & ~n_1701;
assign n_19464 =  x_2031 &  n_1701;
assign n_19465 = ~n_19463 & ~n_19464;
assign n_19466 =  x_464 & ~n_19465;
assign n_19467 = ~x_464 &  n_19465;
assign n_19468 = ~n_19466 & ~n_19467;
assign n_19469 =  x_463 & ~n_1701;
assign n_19470 =  x_2030 &  n_1701;
assign n_19471 = ~n_19469 & ~n_19470;
assign n_19472 =  x_463 & ~n_19471;
assign n_19473 = ~x_463 &  n_19471;
assign n_19474 = ~n_19472 & ~n_19473;
assign n_19475 =  x_462 & ~n_1701;
assign n_19476 =  x_2029 &  n_1701;
assign n_19477 = ~n_19475 & ~n_19476;
assign n_19478 =  x_462 & ~n_19477;
assign n_19479 = ~x_462 &  n_19477;
assign n_19480 = ~n_19478 & ~n_19479;
assign n_19481 =  x_461 & ~n_1701;
assign n_19482 =  x_2028 &  n_1701;
assign n_19483 = ~n_19481 & ~n_19482;
assign n_19484 =  x_461 & ~n_19483;
assign n_19485 = ~x_461 &  n_19483;
assign n_19486 = ~n_19484 & ~n_19485;
assign n_19487 =  x_460 & ~n_1701;
assign n_19488 =  x_2027 &  n_1701;
assign n_19489 = ~n_19487 & ~n_19488;
assign n_19490 =  x_460 & ~n_19489;
assign n_19491 = ~x_460 &  n_19489;
assign n_19492 = ~n_19490 & ~n_19491;
assign n_19493 =  n_556 &  n_1899;
assign n_19494 =  n_2094 &  n_19493;
assign n_19495 =  x_1034 &  n_19494;
assign n_19496 =  n_1037 &  n_770;
assign n_19497 =  n_8359 &  n_556;
assign n_19498 =  n_555 &  n_19497;
assign n_19499 = ~n_19496 & ~n_19498;
assign n_19500 =  n_10872 &  n_8360;
assign n_19501 = ~n_19494 & ~n_19500;
assign n_19502 =  n_19499 &  n_19501;
assign n_19503 =  x_459 &  n_19502;
assign n_19504 = ~n_19495 & ~n_19503;
assign n_19505 =  x_459 & ~n_19504;
assign n_19506 = ~x_459 &  n_19504;
assign n_19507 = ~n_19505 & ~n_19506;
assign n_19508 =  x_1033 &  n_19494;
assign n_19509 =  x_458 &  n_19502;
assign n_19510 = ~n_19508 & ~n_19509;
assign n_19511 =  x_458 & ~n_19510;
assign n_19512 = ~x_458 &  n_19510;
assign n_19513 = ~n_19511 & ~n_19512;
assign n_19514 =  x_1032 &  n_19494;
assign n_19515 =  x_457 &  n_19502;
assign n_19516 = ~n_19514 & ~n_19515;
assign n_19517 =  x_457 & ~n_19516;
assign n_19518 = ~x_457 &  n_19516;
assign n_19519 = ~n_19517 & ~n_19518;
assign n_19520 =  x_1031 &  n_19494;
assign n_19521 =  x_456 &  n_19502;
assign n_19522 = ~n_19520 & ~n_19521;
assign n_19523 =  x_456 & ~n_19522;
assign n_19524 = ~x_456 &  n_19522;
assign n_19525 = ~n_19523 & ~n_19524;
assign n_19526 =  x_1030 &  n_19494;
assign n_19527 =  x_455 &  n_19502;
assign n_19528 = ~n_19526 & ~n_19527;
assign n_19529 =  x_455 & ~n_19528;
assign n_19530 = ~x_455 &  n_19528;
assign n_19531 = ~n_19529 & ~n_19530;
assign n_19532 =  x_1029 &  n_19494;
assign n_19533 =  x_454 &  n_19502;
assign n_19534 = ~n_19532 & ~n_19533;
assign n_19535 =  x_454 & ~n_19534;
assign n_19536 = ~x_454 &  n_19534;
assign n_19537 = ~n_19535 & ~n_19536;
assign n_19538 =  x_1028 &  n_19494;
assign n_19539 =  x_453 &  n_19502;
assign n_19540 = ~n_19538 & ~n_19539;
assign n_19541 =  x_453 & ~n_19540;
assign n_19542 = ~x_453 &  n_19540;
assign n_19543 = ~n_19541 & ~n_19542;
assign n_19544 =  x_1027 &  n_19494;
assign n_19545 =  x_452 &  n_19502;
assign n_19546 = ~n_19544 & ~n_19545;
assign n_19547 =  x_452 & ~n_19546;
assign n_19548 = ~x_452 &  n_19546;
assign n_19549 = ~n_19547 & ~n_19548;
assign n_19550 =  x_1026 &  n_19494;
assign n_19551 =  x_451 &  n_19502;
assign n_19552 = ~n_19550 & ~n_19551;
assign n_19553 =  x_451 & ~n_19552;
assign n_19554 = ~x_451 &  n_19552;
assign n_19555 = ~n_19553 & ~n_19554;
assign n_19556 =  x_1025 &  n_19494;
assign n_19557 =  x_450 &  n_19502;
assign n_19558 = ~n_19556 & ~n_19557;
assign n_19559 =  x_450 & ~n_19558;
assign n_19560 = ~x_450 &  n_19558;
assign n_19561 = ~n_19559 & ~n_19560;
assign n_19562 =  x_1024 &  n_19494;
assign n_19563 =  x_449 &  n_19502;
assign n_19564 = ~n_19562 & ~n_19563;
assign n_19565 =  x_449 & ~n_19564;
assign n_19566 = ~x_449 &  n_19564;
assign n_19567 = ~n_19565 & ~n_19566;
assign n_19568 =  x_1023 &  n_19494;
assign n_19569 =  x_448 &  n_19502;
assign n_19570 = ~n_19568 & ~n_19569;
assign n_19571 =  x_448 & ~n_19570;
assign n_19572 = ~x_448 &  n_19570;
assign n_19573 = ~n_19571 & ~n_19572;
assign n_19574 =  x_1022 &  n_19494;
assign n_19575 =  x_447 &  n_19502;
assign n_19576 = ~n_19574 & ~n_19575;
assign n_19577 =  x_447 & ~n_19576;
assign n_19578 = ~x_447 &  n_19576;
assign n_19579 = ~n_19577 & ~n_19578;
assign n_19580 =  x_1021 &  n_19494;
assign n_19581 =  x_446 &  n_19502;
assign n_19582 = ~n_19580 & ~n_19581;
assign n_19583 =  x_446 & ~n_19582;
assign n_19584 = ~x_446 &  n_19582;
assign n_19585 = ~n_19583 & ~n_19584;
assign n_19586 =  x_1020 &  n_19494;
assign n_19587 =  x_445 &  n_19502;
assign n_19588 = ~n_19586 & ~n_19587;
assign n_19589 =  x_445 & ~n_19588;
assign n_19590 = ~x_445 &  n_19588;
assign n_19591 = ~n_19589 & ~n_19590;
assign n_19592 =  x_1019 &  n_19494;
assign n_19593 =  x_444 &  n_19502;
assign n_19594 = ~n_19592 & ~n_19593;
assign n_19595 =  x_444 & ~n_19594;
assign n_19596 = ~x_444 &  n_19594;
assign n_19597 = ~n_19595 & ~n_19596;
assign n_19598 =  x_1018 &  n_19494;
assign n_19599 =  x_443 &  n_19502;
assign n_19600 = ~n_19598 & ~n_19599;
assign n_19601 =  x_443 & ~n_19600;
assign n_19602 = ~x_443 &  n_19600;
assign n_19603 = ~n_19601 & ~n_19602;
assign n_19604 =  x_1017 &  n_19494;
assign n_19605 =  x_442 &  n_19502;
assign n_19606 = ~n_19604 & ~n_19605;
assign n_19607 =  x_442 & ~n_19606;
assign n_19608 = ~x_442 &  n_19606;
assign n_19609 = ~n_19607 & ~n_19608;
assign n_19610 =  x_1016 &  n_19494;
assign n_19611 =  x_441 &  n_19502;
assign n_19612 = ~n_19610 & ~n_19611;
assign n_19613 =  x_441 & ~n_19612;
assign n_19614 = ~x_441 &  n_19612;
assign n_19615 = ~n_19613 & ~n_19614;
assign n_19616 =  x_1015 &  n_19494;
assign n_19617 =  x_440 &  n_19502;
assign n_19618 = ~n_19616 & ~n_19617;
assign n_19619 =  x_440 & ~n_19618;
assign n_19620 = ~x_440 &  n_19618;
assign n_19621 = ~n_19619 & ~n_19620;
assign n_19622 =  x_1014 &  n_19494;
assign n_19623 =  x_439 &  n_19502;
assign n_19624 = ~n_19622 & ~n_19623;
assign n_19625 =  x_439 & ~n_19624;
assign n_19626 = ~x_439 &  n_19624;
assign n_19627 = ~n_19625 & ~n_19626;
assign n_19628 =  x_1013 &  n_19494;
assign n_19629 =  x_438 &  n_19502;
assign n_19630 = ~n_19628 & ~n_19629;
assign n_19631 =  x_438 & ~n_19630;
assign n_19632 = ~x_438 &  n_19630;
assign n_19633 = ~n_19631 & ~n_19632;
assign n_19634 =  x_1012 &  n_19494;
assign n_19635 =  x_437 &  n_19502;
assign n_19636 = ~n_19634 & ~n_19635;
assign n_19637 =  x_437 & ~n_19636;
assign n_19638 = ~x_437 &  n_19636;
assign n_19639 = ~n_19637 & ~n_19638;
assign n_19640 =  x_1011 &  n_19494;
assign n_19641 =  x_436 &  n_19502;
assign n_19642 = ~n_19640 & ~n_19641;
assign n_19643 =  x_436 & ~n_19642;
assign n_19644 = ~x_436 &  n_19642;
assign n_19645 = ~n_19643 & ~n_19644;
assign n_19646 =  x_1010 &  n_19494;
assign n_19647 =  x_435 &  n_19502;
assign n_19648 = ~n_19646 & ~n_19647;
assign n_19649 =  x_435 & ~n_19648;
assign n_19650 = ~x_435 &  n_19648;
assign n_19651 = ~n_19649 & ~n_19650;
assign n_19652 =  x_1009 &  n_19494;
assign n_19653 =  x_434 &  n_19502;
assign n_19654 = ~n_19652 & ~n_19653;
assign n_19655 =  x_434 & ~n_19654;
assign n_19656 = ~x_434 &  n_19654;
assign n_19657 = ~n_19655 & ~n_19656;
assign n_19658 =  x_1008 &  n_19494;
assign n_19659 =  x_433 &  n_19502;
assign n_19660 = ~n_19658 & ~n_19659;
assign n_19661 =  x_433 & ~n_19660;
assign n_19662 = ~x_433 &  n_19660;
assign n_19663 = ~n_19661 & ~n_19662;
assign n_19664 =  x_1007 &  n_19494;
assign n_19665 =  x_432 &  n_19502;
assign n_19666 = ~n_19664 & ~n_19665;
assign n_19667 =  x_432 & ~n_19666;
assign n_19668 = ~x_432 &  n_19666;
assign n_19669 = ~n_19667 & ~n_19668;
assign n_19670 =  x_1006 &  n_19494;
assign n_19671 =  x_431 &  n_19502;
assign n_19672 = ~n_19670 & ~n_19671;
assign n_19673 =  x_431 & ~n_19672;
assign n_19674 = ~x_431 &  n_19672;
assign n_19675 = ~n_19673 & ~n_19674;
assign n_19676 =  x_1005 &  n_19494;
assign n_19677 =  x_430 &  n_19502;
assign n_19678 = ~n_19676 & ~n_19677;
assign n_19679 =  x_430 & ~n_19678;
assign n_19680 = ~x_430 &  n_19678;
assign n_19681 = ~n_19679 & ~n_19680;
assign n_19682 =  x_1004 &  n_19494;
assign n_19683 =  x_429 &  n_19502;
assign n_19684 = ~n_19682 & ~n_19683;
assign n_19685 =  x_429 & ~n_19684;
assign n_19686 = ~x_429 &  n_19684;
assign n_19687 = ~n_19685 & ~n_19686;
assign n_19688 =  x_1003 &  n_19494;
assign n_19689 =  x_428 &  n_19502;
assign n_19690 = ~n_19688 & ~n_19689;
assign n_19691 =  x_428 & ~n_19690;
assign n_19692 = ~x_428 &  n_19690;
assign n_19693 = ~n_19691 & ~n_19692;
assign n_19694 =  n_8361 &  n_1900;
assign n_19695 =  x_427 & ~n_19694;
assign n_19696 =  x_2458 &  n_19694;
assign n_19697 = ~n_19695 & ~n_19696;
assign n_19698 =  x_427 & ~n_19697;
assign n_19699 = ~x_427 &  n_19697;
assign n_19700 = ~n_19698 & ~n_19699;
assign n_19701 =  x_426 & ~n_19694;
assign n_19702 =  x_2457 &  n_19694;
assign n_19703 = ~n_19701 & ~n_19702;
assign n_19704 =  x_426 & ~n_19703;
assign n_19705 = ~x_426 &  n_19703;
assign n_19706 = ~n_19704 & ~n_19705;
assign n_19707 =  x_425 & ~n_19694;
assign n_19708 =  x_2456 &  n_19694;
assign n_19709 = ~n_19707 & ~n_19708;
assign n_19710 =  x_425 & ~n_19709;
assign n_19711 = ~x_425 &  n_19709;
assign n_19712 = ~n_19710 & ~n_19711;
assign n_19713 =  x_424 & ~n_19694;
assign n_19714 =  x_2455 &  n_19694;
assign n_19715 = ~n_19713 & ~n_19714;
assign n_19716 =  x_424 & ~n_19715;
assign n_19717 = ~x_424 &  n_19715;
assign n_19718 = ~n_19716 & ~n_19717;
assign n_19719 =  x_423 & ~n_19694;
assign n_19720 =  x_2454 &  n_19694;
assign n_19721 = ~n_19719 & ~n_19720;
assign n_19722 =  x_423 & ~n_19721;
assign n_19723 = ~x_423 &  n_19721;
assign n_19724 = ~n_19722 & ~n_19723;
assign n_19725 =  x_422 & ~n_19694;
assign n_19726 =  x_2453 &  n_19694;
assign n_19727 = ~n_19725 & ~n_19726;
assign n_19728 =  x_422 & ~n_19727;
assign n_19729 = ~x_422 &  n_19727;
assign n_19730 = ~n_19728 & ~n_19729;
assign n_19731 =  x_421 & ~n_19694;
assign n_19732 =  x_2452 &  n_19694;
assign n_19733 = ~n_19731 & ~n_19732;
assign n_19734 =  x_421 & ~n_19733;
assign n_19735 = ~x_421 &  n_19733;
assign n_19736 = ~n_19734 & ~n_19735;
assign n_19737 =  x_420 & ~n_19694;
assign n_19738 =  x_2451 &  n_19694;
assign n_19739 = ~n_19737 & ~n_19738;
assign n_19740 =  x_420 & ~n_19739;
assign n_19741 = ~x_420 &  n_19739;
assign n_19742 = ~n_19740 & ~n_19741;
assign n_19743 =  x_419 & ~n_19694;
assign n_19744 =  x_2450 &  n_19694;
assign n_19745 = ~n_19743 & ~n_19744;
assign n_19746 =  x_419 & ~n_19745;
assign n_19747 = ~x_419 &  n_19745;
assign n_19748 = ~n_19746 & ~n_19747;
assign n_19749 =  x_418 & ~n_19694;
assign n_19750 =  x_2449 &  n_19694;
assign n_19751 = ~n_19749 & ~n_19750;
assign n_19752 =  x_418 & ~n_19751;
assign n_19753 = ~x_418 &  n_19751;
assign n_19754 = ~n_19752 & ~n_19753;
assign n_19755 =  x_417 & ~n_19694;
assign n_19756 =  x_2448 &  n_19694;
assign n_19757 = ~n_19755 & ~n_19756;
assign n_19758 =  x_417 & ~n_19757;
assign n_19759 = ~x_417 &  n_19757;
assign n_19760 = ~n_19758 & ~n_19759;
assign n_19761 =  x_416 & ~n_19694;
assign n_19762 =  x_2447 &  n_19694;
assign n_19763 = ~n_19761 & ~n_19762;
assign n_19764 =  x_416 & ~n_19763;
assign n_19765 = ~x_416 &  n_19763;
assign n_19766 = ~n_19764 & ~n_19765;
assign n_19767 =  x_415 & ~n_19694;
assign n_19768 =  x_2446 &  n_19694;
assign n_19769 = ~n_19767 & ~n_19768;
assign n_19770 =  x_415 & ~n_19769;
assign n_19771 = ~x_415 &  n_19769;
assign n_19772 = ~n_19770 & ~n_19771;
assign n_19773 =  x_414 & ~n_19694;
assign n_19774 =  x_2445 &  n_19694;
assign n_19775 = ~n_19773 & ~n_19774;
assign n_19776 =  x_414 & ~n_19775;
assign n_19777 = ~x_414 &  n_19775;
assign n_19778 = ~n_19776 & ~n_19777;
assign n_19779 =  x_413 & ~n_19694;
assign n_19780 =  x_2444 &  n_19694;
assign n_19781 = ~n_19779 & ~n_19780;
assign n_19782 =  x_413 & ~n_19781;
assign n_19783 = ~x_413 &  n_19781;
assign n_19784 = ~n_19782 & ~n_19783;
assign n_19785 =  x_412 & ~n_19694;
assign n_19786 =  x_2443 &  n_19694;
assign n_19787 = ~n_19785 & ~n_19786;
assign n_19788 =  x_412 & ~n_19787;
assign n_19789 = ~x_412 &  n_19787;
assign n_19790 = ~n_19788 & ~n_19789;
assign n_19791 =  x_411 & ~n_19694;
assign n_19792 =  x_2442 &  n_19694;
assign n_19793 = ~n_19791 & ~n_19792;
assign n_19794 =  x_411 & ~n_19793;
assign n_19795 = ~x_411 &  n_19793;
assign n_19796 = ~n_19794 & ~n_19795;
assign n_19797 =  x_410 & ~n_19694;
assign n_19798 =  x_2441 &  n_19694;
assign n_19799 = ~n_19797 & ~n_19798;
assign n_19800 =  x_410 & ~n_19799;
assign n_19801 = ~x_410 &  n_19799;
assign n_19802 = ~n_19800 & ~n_19801;
assign n_19803 =  x_409 & ~n_19694;
assign n_19804 =  x_2440 &  n_19694;
assign n_19805 = ~n_19803 & ~n_19804;
assign n_19806 =  x_409 & ~n_19805;
assign n_19807 = ~x_409 &  n_19805;
assign n_19808 = ~n_19806 & ~n_19807;
assign n_19809 =  x_408 & ~n_19694;
assign n_19810 =  x_2439 &  n_19694;
assign n_19811 = ~n_19809 & ~n_19810;
assign n_19812 =  x_408 & ~n_19811;
assign n_19813 = ~x_408 &  n_19811;
assign n_19814 = ~n_19812 & ~n_19813;
assign n_19815 =  x_407 & ~n_19694;
assign n_19816 =  x_2438 &  n_19694;
assign n_19817 = ~n_19815 & ~n_19816;
assign n_19818 =  x_407 & ~n_19817;
assign n_19819 = ~x_407 &  n_19817;
assign n_19820 = ~n_19818 & ~n_19819;
assign n_19821 =  x_406 & ~n_19694;
assign n_19822 =  x_2437 &  n_19694;
assign n_19823 = ~n_19821 & ~n_19822;
assign n_19824 =  x_406 & ~n_19823;
assign n_19825 = ~x_406 &  n_19823;
assign n_19826 = ~n_19824 & ~n_19825;
assign n_19827 =  x_405 & ~n_19694;
assign n_19828 =  x_2436 &  n_19694;
assign n_19829 = ~n_19827 & ~n_19828;
assign n_19830 =  x_405 & ~n_19829;
assign n_19831 = ~x_405 &  n_19829;
assign n_19832 = ~n_19830 & ~n_19831;
assign n_19833 =  x_404 & ~n_19694;
assign n_19834 =  x_2435 &  n_19694;
assign n_19835 = ~n_19833 & ~n_19834;
assign n_19836 =  x_404 & ~n_19835;
assign n_19837 = ~x_404 &  n_19835;
assign n_19838 = ~n_19836 & ~n_19837;
assign n_19839 =  x_403 & ~n_19694;
assign n_19840 =  x_2434 &  n_19694;
assign n_19841 = ~n_19839 & ~n_19840;
assign n_19842 =  x_403 & ~n_19841;
assign n_19843 = ~x_403 &  n_19841;
assign n_19844 = ~n_19842 & ~n_19843;
assign n_19845 =  x_402 & ~n_19694;
assign n_19846 =  x_2433 &  n_19694;
assign n_19847 = ~n_19845 & ~n_19846;
assign n_19848 =  x_402 & ~n_19847;
assign n_19849 = ~x_402 &  n_19847;
assign n_19850 = ~n_19848 & ~n_19849;
assign n_19851 =  x_401 & ~n_19694;
assign n_19852 =  x_2432 &  n_19694;
assign n_19853 = ~n_19851 & ~n_19852;
assign n_19854 =  x_401 & ~n_19853;
assign n_19855 = ~x_401 &  n_19853;
assign n_19856 = ~n_19854 & ~n_19855;
assign n_19857 =  x_400 & ~n_19694;
assign n_19858 =  x_2431 &  n_19694;
assign n_19859 = ~n_19857 & ~n_19858;
assign n_19860 =  x_400 & ~n_19859;
assign n_19861 = ~x_400 &  n_19859;
assign n_19862 = ~n_19860 & ~n_19861;
assign n_19863 =  x_399 & ~n_19694;
assign n_19864 =  x_2430 &  n_19694;
assign n_19865 = ~n_19863 & ~n_19864;
assign n_19866 =  x_399 & ~n_19865;
assign n_19867 = ~x_399 &  n_19865;
assign n_19868 = ~n_19866 & ~n_19867;
assign n_19869 =  x_398 & ~n_19694;
assign n_19870 =  x_2429 &  n_19694;
assign n_19871 = ~n_19869 & ~n_19870;
assign n_19872 =  x_398 & ~n_19871;
assign n_19873 = ~x_398 &  n_19871;
assign n_19874 = ~n_19872 & ~n_19873;
assign n_19875 =  x_397 & ~n_19694;
assign n_19876 =  x_2428 &  n_19694;
assign n_19877 = ~n_19875 & ~n_19876;
assign n_19878 =  x_397 & ~n_19877;
assign n_19879 = ~x_397 &  n_19877;
assign n_19880 = ~n_19878 & ~n_19879;
assign n_19881 =  x_396 & ~n_19694;
assign n_19882 =  x_396 &  n_19881;
assign n_19883 = ~x_396 & ~n_19881;
assign n_19884 = ~n_19882 & ~n_19883;
assign n_19885 =  x_2186 &  n_16882;
assign n_19886 =  x_395 &  n_16884;
assign n_19887 = ~n_19885 & ~n_19886;
assign n_19888 =  x_395 & ~n_19887;
assign n_19889 = ~x_395 &  n_19887;
assign n_19890 = ~n_19888 & ~n_19889;
assign n_19891 =  x_2185 &  n_16882;
assign n_19892 =  x_394 &  n_16884;
assign n_19893 = ~n_19891 & ~n_19892;
assign n_19894 =  x_394 & ~n_19893;
assign n_19895 = ~x_394 &  n_19893;
assign n_19896 = ~n_19894 & ~n_19895;
assign n_19897 =  x_2184 &  n_16882;
assign n_19898 =  x_393 &  n_16884;
assign n_19899 = ~n_19897 & ~n_19898;
assign n_19900 =  x_393 & ~n_19899;
assign n_19901 = ~x_393 &  n_19899;
assign n_19902 = ~n_19900 & ~n_19901;
assign n_19903 =  x_2183 &  n_16882;
assign n_19904 =  x_392 &  n_16884;
assign n_19905 = ~n_19903 & ~n_19904;
assign n_19906 =  x_392 & ~n_19905;
assign n_19907 = ~x_392 &  n_19905;
assign n_19908 = ~n_19906 & ~n_19907;
assign n_19909 =  x_2182 &  n_16882;
assign n_19910 =  x_391 &  n_16884;
assign n_19911 = ~n_19909 & ~n_19910;
assign n_19912 =  x_391 & ~n_19911;
assign n_19913 = ~x_391 &  n_19911;
assign n_19914 = ~n_19912 & ~n_19913;
assign n_19915 =  x_2181 &  n_16882;
assign n_19916 =  x_390 &  n_16884;
assign n_19917 = ~n_19915 & ~n_19916;
assign n_19918 =  x_390 & ~n_19917;
assign n_19919 = ~x_390 &  n_19917;
assign n_19920 = ~n_19918 & ~n_19919;
assign n_19921 =  x_2180 &  n_16882;
assign n_19922 =  x_389 &  n_16884;
assign n_19923 = ~n_19921 & ~n_19922;
assign n_19924 =  x_389 & ~n_19923;
assign n_19925 = ~x_389 &  n_19923;
assign n_19926 = ~n_19924 & ~n_19925;
assign n_19927 =  x_2179 &  n_16882;
assign n_19928 =  x_388 &  n_16884;
assign n_19929 = ~n_19927 & ~n_19928;
assign n_19930 =  x_388 & ~n_19929;
assign n_19931 = ~x_388 &  n_19929;
assign n_19932 = ~n_19930 & ~n_19931;
assign n_19933 =  x_2178 &  n_16882;
assign n_19934 =  x_387 &  n_16884;
assign n_19935 = ~n_19933 & ~n_19934;
assign n_19936 =  x_387 & ~n_19935;
assign n_19937 = ~x_387 &  n_19935;
assign n_19938 = ~n_19936 & ~n_19937;
assign n_19939 =  x_2177 &  n_16882;
assign n_19940 =  x_386 &  n_16884;
assign n_19941 = ~n_19939 & ~n_19940;
assign n_19942 =  x_386 & ~n_19941;
assign n_19943 = ~x_386 &  n_19941;
assign n_19944 = ~n_19942 & ~n_19943;
assign n_19945 =  x_2176 &  n_16882;
assign n_19946 =  x_385 &  n_16884;
assign n_19947 = ~n_19945 & ~n_19946;
assign n_19948 =  x_385 & ~n_19947;
assign n_19949 = ~x_385 &  n_19947;
assign n_19950 = ~n_19948 & ~n_19949;
assign n_19951 =  x_2175 &  n_16882;
assign n_19952 =  x_384 &  n_16884;
assign n_19953 = ~n_19951 & ~n_19952;
assign n_19954 =  x_384 & ~n_19953;
assign n_19955 = ~x_384 &  n_19953;
assign n_19956 = ~n_19954 & ~n_19955;
assign n_19957 =  x_2174 &  n_16882;
assign n_19958 =  x_383 &  n_16884;
assign n_19959 = ~n_19957 & ~n_19958;
assign n_19960 =  x_383 & ~n_19959;
assign n_19961 = ~x_383 &  n_19959;
assign n_19962 = ~n_19960 & ~n_19961;
assign n_19963 =  x_2173 &  n_16882;
assign n_19964 =  x_382 &  n_16884;
assign n_19965 = ~n_19963 & ~n_19964;
assign n_19966 =  x_382 & ~n_19965;
assign n_19967 = ~x_382 &  n_19965;
assign n_19968 = ~n_19966 & ~n_19967;
assign n_19969 =  x_2172 &  n_16882;
assign n_19970 =  x_381 &  n_16884;
assign n_19971 = ~n_19969 & ~n_19970;
assign n_19972 =  x_381 & ~n_19971;
assign n_19973 = ~x_381 &  n_19971;
assign n_19974 = ~n_19972 & ~n_19973;
assign n_19975 =  x_2171 &  n_16882;
assign n_19976 =  x_380 &  n_16884;
assign n_19977 = ~n_19975 & ~n_19976;
assign n_19978 =  x_380 & ~n_19977;
assign n_19979 = ~x_380 &  n_19977;
assign n_19980 = ~n_19978 & ~n_19979;
assign n_19981 =  x_2170 &  n_16882;
assign n_19982 =  x_379 &  n_16884;
assign n_19983 = ~n_19981 & ~n_19982;
assign n_19984 =  x_379 & ~n_19983;
assign n_19985 = ~x_379 &  n_19983;
assign n_19986 = ~n_19984 & ~n_19985;
assign n_19987 =  x_2169 &  n_16882;
assign n_19988 =  x_378 &  n_16884;
assign n_19989 = ~n_19987 & ~n_19988;
assign n_19990 =  x_378 & ~n_19989;
assign n_19991 = ~x_378 &  n_19989;
assign n_19992 = ~n_19990 & ~n_19991;
assign n_19993 =  x_2168 &  n_16882;
assign n_19994 =  x_377 &  n_16884;
assign n_19995 = ~n_19993 & ~n_19994;
assign n_19996 =  x_377 & ~n_19995;
assign n_19997 = ~x_377 &  n_19995;
assign n_19998 = ~n_19996 & ~n_19997;
assign n_19999 =  x_2167 &  n_16882;
assign n_20000 =  x_376 &  n_16884;
assign n_20001 = ~n_19999 & ~n_20000;
assign n_20002 =  x_376 & ~n_20001;
assign n_20003 = ~x_376 &  n_20001;
assign n_20004 = ~n_20002 & ~n_20003;
assign n_20005 =  x_2166 &  n_16882;
assign n_20006 =  x_375 &  n_16884;
assign n_20007 = ~n_20005 & ~n_20006;
assign n_20008 =  x_375 & ~n_20007;
assign n_20009 = ~x_375 &  n_20007;
assign n_20010 = ~n_20008 & ~n_20009;
assign n_20011 =  x_2165 &  n_16882;
assign n_20012 =  x_374 &  n_16884;
assign n_20013 = ~n_20011 & ~n_20012;
assign n_20014 =  x_374 & ~n_20013;
assign n_20015 = ~x_374 &  n_20013;
assign n_20016 = ~n_20014 & ~n_20015;
assign n_20017 =  x_2164 &  n_16882;
assign n_20018 =  x_373 &  n_16884;
assign n_20019 = ~n_20017 & ~n_20018;
assign n_20020 =  x_373 & ~n_20019;
assign n_20021 = ~x_373 &  n_20019;
assign n_20022 = ~n_20020 & ~n_20021;
assign n_20023 =  x_2163 &  n_16882;
assign n_20024 =  x_372 &  n_16884;
assign n_20025 = ~n_20023 & ~n_20024;
assign n_20026 =  x_372 & ~n_20025;
assign n_20027 = ~x_372 &  n_20025;
assign n_20028 = ~n_20026 & ~n_20027;
assign n_20029 =  x_2162 &  n_16882;
assign n_20030 =  x_371 &  n_16884;
assign n_20031 = ~n_20029 & ~n_20030;
assign n_20032 =  x_371 & ~n_20031;
assign n_20033 = ~x_371 &  n_20031;
assign n_20034 = ~n_20032 & ~n_20033;
assign n_20035 =  x_2161 &  n_16882;
assign n_20036 =  x_370 &  n_16884;
assign n_20037 = ~n_20035 & ~n_20036;
assign n_20038 =  x_370 & ~n_20037;
assign n_20039 = ~x_370 &  n_20037;
assign n_20040 = ~n_20038 & ~n_20039;
assign n_20041 =  x_2160 &  n_16882;
assign n_20042 =  x_369 &  n_16884;
assign n_20043 = ~n_20041 & ~n_20042;
assign n_20044 =  x_369 & ~n_20043;
assign n_20045 = ~x_369 &  n_20043;
assign n_20046 = ~n_20044 & ~n_20045;
assign n_20047 =  x_2159 &  n_16882;
assign n_20048 =  x_368 &  n_16884;
assign n_20049 = ~n_20047 & ~n_20048;
assign n_20050 =  x_368 & ~n_20049;
assign n_20051 = ~x_368 &  n_20049;
assign n_20052 = ~n_20050 & ~n_20051;
assign n_20053 =  x_2158 &  n_16882;
assign n_20054 =  x_367 &  n_16884;
assign n_20055 = ~n_20053 & ~n_20054;
assign n_20056 =  x_367 & ~n_20055;
assign n_20057 = ~x_367 &  n_20055;
assign n_20058 = ~n_20056 & ~n_20057;
assign n_20059 =  x_2157 &  n_16882;
assign n_20060 =  x_366 &  n_16884;
assign n_20061 = ~n_20059 & ~n_20060;
assign n_20062 =  x_366 & ~n_20061;
assign n_20063 = ~x_366 &  n_20061;
assign n_20064 = ~n_20062 & ~n_20063;
assign n_20065 =  x_2156 &  n_16882;
assign n_20066 =  x_365 &  n_16884;
assign n_20067 = ~n_20065 & ~n_20066;
assign n_20068 =  x_365 & ~n_20067;
assign n_20069 = ~x_365 &  n_20067;
assign n_20070 = ~n_20068 & ~n_20069;
assign n_20071 =  x_2155 &  n_16882;
assign n_20072 =  x_364 &  n_16884;
assign n_20073 = ~n_20071 & ~n_20072;
assign n_20074 =  x_364 & ~n_20073;
assign n_20075 = ~x_364 &  n_20073;
assign n_20076 = ~n_20074 & ~n_20075;
assign n_20077 =  n_5651 &  n_2486;
assign n_20078 =  n_5645 &  n_20077;
assign n_20079 =  x_363 & ~n_20078;
assign n_20080 =  x_363 &  n_20079;
assign n_20081 = ~x_363 & ~n_20079;
assign n_20082 = ~n_20080 & ~n_20081;
assign n_20083 =  x_362 & ~n_20078;
assign n_20084 =  x_362 &  n_20083;
assign n_20085 = ~x_362 & ~n_20083;
assign n_20086 = ~n_20084 & ~n_20085;
assign n_20087 =  x_361 & ~n_20078;
assign n_20088 =  x_361 &  n_20087;
assign n_20089 = ~x_361 & ~n_20087;
assign n_20090 = ~n_20088 & ~n_20089;
assign n_20091 =  x_360 & ~n_20078;
assign n_20092 =  x_360 &  n_20091;
assign n_20093 = ~x_360 & ~n_20091;
assign n_20094 = ~n_20092 & ~n_20093;
assign n_20095 =  x_359 & ~n_20078;
assign n_20096 =  x_359 &  n_20095;
assign n_20097 = ~x_359 & ~n_20095;
assign n_20098 = ~n_20096 & ~n_20097;
assign n_20099 =  x_358 & ~n_20078;
assign n_20100 =  x_358 &  n_20099;
assign n_20101 = ~x_358 & ~n_20099;
assign n_20102 = ~n_20100 & ~n_20101;
assign n_20103 =  x_357 & ~n_20078;
assign n_20104 =  x_357 &  n_20103;
assign n_20105 = ~x_357 & ~n_20103;
assign n_20106 = ~n_20104 & ~n_20105;
assign n_20107 =  x_356 & ~n_20078;
assign n_20108 =  x_356 &  n_20107;
assign n_20109 = ~x_356 & ~n_20107;
assign n_20110 = ~n_20108 & ~n_20109;
assign n_20111 =  x_355 & ~n_20078;
assign n_20112 =  x_355 &  n_20111;
assign n_20113 = ~x_355 & ~n_20111;
assign n_20114 = ~n_20112 & ~n_20113;
assign n_20115 =  x_354 & ~n_20078;
assign n_20116 =  x_354 &  n_20115;
assign n_20117 = ~x_354 & ~n_20115;
assign n_20118 = ~n_20116 & ~n_20117;
assign n_20119 =  x_353 & ~n_20078;
assign n_20120 =  x_353 &  n_20119;
assign n_20121 = ~x_353 & ~n_20119;
assign n_20122 = ~n_20120 & ~n_20121;
assign n_20123 =  x_352 & ~n_20078;
assign n_20124 =  x_352 &  n_20123;
assign n_20125 = ~x_352 & ~n_20123;
assign n_20126 = ~n_20124 & ~n_20125;
assign n_20127 =  x_351 & ~n_20078;
assign n_20128 =  x_351 &  n_20127;
assign n_20129 = ~x_351 & ~n_20127;
assign n_20130 = ~n_20128 & ~n_20129;
assign n_20131 =  x_350 & ~n_20078;
assign n_20132 =  x_350 &  n_20131;
assign n_20133 = ~x_350 & ~n_20131;
assign n_20134 = ~n_20132 & ~n_20133;
assign n_20135 =  x_349 & ~n_20078;
assign n_20136 =  x_349 &  n_20135;
assign n_20137 = ~x_349 & ~n_20135;
assign n_20138 = ~n_20136 & ~n_20137;
assign n_20139 =  x_348 & ~n_20078;
assign n_20140 =  x_348 &  n_20139;
assign n_20141 = ~x_348 & ~n_20139;
assign n_20142 = ~n_20140 & ~n_20141;
assign n_20143 =  x_347 & ~n_20078;
assign n_20144 =  x_347 &  n_20143;
assign n_20145 = ~x_347 & ~n_20143;
assign n_20146 = ~n_20144 & ~n_20145;
assign n_20147 =  x_346 & ~n_20078;
assign n_20148 =  x_346 &  n_20147;
assign n_20149 = ~x_346 & ~n_20147;
assign n_20150 = ~n_20148 & ~n_20149;
assign n_20151 =  x_345 & ~n_20078;
assign n_20152 =  x_345 &  n_20151;
assign n_20153 = ~x_345 & ~n_20151;
assign n_20154 = ~n_20152 & ~n_20153;
assign n_20155 =  x_344 & ~n_20078;
assign n_20156 =  x_344 &  n_20155;
assign n_20157 = ~x_344 & ~n_20155;
assign n_20158 = ~n_20156 & ~n_20157;
assign n_20159 =  x_343 & ~n_20078;
assign n_20160 =  x_343 &  n_20159;
assign n_20161 = ~x_343 & ~n_20159;
assign n_20162 = ~n_20160 & ~n_20161;
assign n_20163 =  x_342 & ~n_20078;
assign n_20164 =  x_342 &  n_20163;
assign n_20165 = ~x_342 & ~n_20163;
assign n_20166 = ~n_20164 & ~n_20165;
assign n_20167 =  x_341 & ~n_20078;
assign n_20168 =  x_341 &  n_20167;
assign n_20169 = ~x_341 & ~n_20167;
assign n_20170 = ~n_20168 & ~n_20169;
assign n_20171 =  x_340 & ~n_20078;
assign n_20172 =  x_340 &  n_20171;
assign n_20173 = ~x_340 & ~n_20171;
assign n_20174 = ~n_20172 & ~n_20173;
assign n_20175 =  x_339 & ~n_20078;
assign n_20176 =  x_339 &  n_20175;
assign n_20177 = ~x_339 & ~n_20175;
assign n_20178 = ~n_20176 & ~n_20177;
assign n_20179 =  x_338 & ~n_20078;
assign n_20180 =  x_338 &  n_20179;
assign n_20181 = ~x_338 & ~n_20179;
assign n_20182 = ~n_20180 & ~n_20181;
assign n_20183 =  x_337 & ~n_20078;
assign n_20184 =  x_337 &  n_20183;
assign n_20185 = ~x_337 & ~n_20183;
assign n_20186 = ~n_20184 & ~n_20185;
assign n_20187 =  x_336 & ~n_20078;
assign n_20188 =  x_336 &  n_20187;
assign n_20189 = ~x_336 & ~n_20187;
assign n_20190 = ~n_20188 & ~n_20189;
assign n_20191 =  x_335 & ~n_20078;
assign n_20192 =  x_335 &  n_20191;
assign n_20193 = ~x_335 & ~n_20191;
assign n_20194 = ~n_20192 & ~n_20193;
assign n_20195 =  x_334 & ~n_20078;
assign n_20196 =  x_334 &  n_20195;
assign n_20197 = ~x_334 & ~n_20195;
assign n_20198 = ~n_20196 & ~n_20197;
assign n_20199 =  x_333 & ~n_20078;
assign n_20200 =  x_333 &  n_20199;
assign n_20201 = ~x_333 & ~n_20199;
assign n_20202 = ~n_20200 & ~n_20201;
assign n_20203 =  x_332 & ~n_20078;
assign n_20204 =  x_332 &  n_20203;
assign n_20205 = ~x_332 & ~n_20203;
assign n_20206 = ~n_20204 & ~n_20205;
assign n_20207 =  n_2290 &  n_7467;
assign n_20208 =  n_150 &  n_20207;
assign n_20209 =  x_331 & ~n_20208;
assign n_20210 =  i_32 &  n_20208;
assign n_20211 = ~n_20209 & ~n_20210;
assign n_20212 =  x_331 & ~n_20211;
assign n_20213 = ~x_331 &  n_20211;
assign n_20214 = ~n_20212 & ~n_20213;
assign n_20215 =  x_330 & ~n_20208;
assign n_20216 =  i_31 &  n_20208;
assign n_20217 = ~n_20215 & ~n_20216;
assign n_20218 =  x_330 & ~n_20217;
assign n_20219 = ~x_330 &  n_20217;
assign n_20220 = ~n_20218 & ~n_20219;
assign n_20221 =  x_329 & ~n_20208;
assign n_20222 =  i_30 &  n_20208;
assign n_20223 = ~n_20221 & ~n_20222;
assign n_20224 =  x_329 & ~n_20223;
assign n_20225 = ~x_329 &  n_20223;
assign n_20226 = ~n_20224 & ~n_20225;
assign n_20227 =  x_328 & ~n_20208;
assign n_20228 =  i_29 &  n_20208;
assign n_20229 = ~n_20227 & ~n_20228;
assign n_20230 =  x_328 & ~n_20229;
assign n_20231 = ~x_328 &  n_20229;
assign n_20232 = ~n_20230 & ~n_20231;
assign n_20233 =  x_327 & ~n_20208;
assign n_20234 =  i_28 &  n_20208;
assign n_20235 = ~n_20233 & ~n_20234;
assign n_20236 =  x_327 & ~n_20235;
assign n_20237 = ~x_327 &  n_20235;
assign n_20238 = ~n_20236 & ~n_20237;
assign n_20239 =  x_326 & ~n_20208;
assign n_20240 =  i_27 &  n_20208;
assign n_20241 = ~n_20239 & ~n_20240;
assign n_20242 =  x_326 & ~n_20241;
assign n_20243 = ~x_326 &  n_20241;
assign n_20244 = ~n_20242 & ~n_20243;
assign n_20245 =  x_325 & ~n_20208;
assign n_20246 =  i_26 &  n_20208;
assign n_20247 = ~n_20245 & ~n_20246;
assign n_20248 =  x_325 & ~n_20247;
assign n_20249 = ~x_325 &  n_20247;
assign n_20250 = ~n_20248 & ~n_20249;
assign n_20251 =  x_324 & ~n_20208;
assign n_20252 =  i_25 &  n_20208;
assign n_20253 = ~n_20251 & ~n_20252;
assign n_20254 =  x_324 & ~n_20253;
assign n_20255 = ~x_324 &  n_20253;
assign n_20256 = ~n_20254 & ~n_20255;
assign n_20257 =  x_323 & ~n_20208;
assign n_20258 =  i_24 &  n_20208;
assign n_20259 = ~n_20257 & ~n_20258;
assign n_20260 =  x_323 & ~n_20259;
assign n_20261 = ~x_323 &  n_20259;
assign n_20262 = ~n_20260 & ~n_20261;
assign n_20263 =  x_322 & ~n_20208;
assign n_20264 =  i_23 &  n_20208;
assign n_20265 = ~n_20263 & ~n_20264;
assign n_20266 =  x_322 & ~n_20265;
assign n_20267 = ~x_322 &  n_20265;
assign n_20268 = ~n_20266 & ~n_20267;
assign n_20269 =  x_321 & ~n_20208;
assign n_20270 =  i_22 &  n_20208;
assign n_20271 = ~n_20269 & ~n_20270;
assign n_20272 =  x_321 & ~n_20271;
assign n_20273 = ~x_321 &  n_20271;
assign n_20274 = ~n_20272 & ~n_20273;
assign n_20275 =  x_320 & ~n_20208;
assign n_20276 =  i_21 &  n_20208;
assign n_20277 = ~n_20275 & ~n_20276;
assign n_20278 =  x_320 & ~n_20277;
assign n_20279 = ~x_320 &  n_20277;
assign n_20280 = ~n_20278 & ~n_20279;
assign n_20281 =  x_319 & ~n_20208;
assign n_20282 =  i_20 &  n_20208;
assign n_20283 = ~n_20281 & ~n_20282;
assign n_20284 =  x_319 & ~n_20283;
assign n_20285 = ~x_319 &  n_20283;
assign n_20286 = ~n_20284 & ~n_20285;
assign n_20287 =  x_318 & ~n_20208;
assign n_20288 =  i_19 &  n_20208;
assign n_20289 = ~n_20287 & ~n_20288;
assign n_20290 =  x_318 & ~n_20289;
assign n_20291 = ~x_318 &  n_20289;
assign n_20292 = ~n_20290 & ~n_20291;
assign n_20293 =  x_317 & ~n_20208;
assign n_20294 =  i_18 &  n_20208;
assign n_20295 = ~n_20293 & ~n_20294;
assign n_20296 =  x_317 & ~n_20295;
assign n_20297 = ~x_317 &  n_20295;
assign n_20298 = ~n_20296 & ~n_20297;
assign n_20299 =  x_316 & ~n_20208;
assign n_20300 =  i_17 &  n_20208;
assign n_20301 = ~n_20299 & ~n_20300;
assign n_20302 =  x_316 & ~n_20301;
assign n_20303 = ~x_316 &  n_20301;
assign n_20304 = ~n_20302 & ~n_20303;
assign n_20305 =  x_315 & ~n_20208;
assign n_20306 =  i_16 &  n_20208;
assign n_20307 = ~n_20305 & ~n_20306;
assign n_20308 =  x_315 & ~n_20307;
assign n_20309 = ~x_315 &  n_20307;
assign n_20310 = ~n_20308 & ~n_20309;
assign n_20311 =  x_314 & ~n_20208;
assign n_20312 =  i_15 &  n_20208;
assign n_20313 = ~n_20311 & ~n_20312;
assign n_20314 =  x_314 & ~n_20313;
assign n_20315 = ~x_314 &  n_20313;
assign n_20316 = ~n_20314 & ~n_20315;
assign n_20317 =  x_313 & ~n_20208;
assign n_20318 =  i_14 &  n_20208;
assign n_20319 = ~n_20317 & ~n_20318;
assign n_20320 =  x_313 & ~n_20319;
assign n_20321 = ~x_313 &  n_20319;
assign n_20322 = ~n_20320 & ~n_20321;
assign n_20323 =  x_312 & ~n_20208;
assign n_20324 =  i_13 &  n_20208;
assign n_20325 = ~n_20323 & ~n_20324;
assign n_20326 =  x_312 & ~n_20325;
assign n_20327 = ~x_312 &  n_20325;
assign n_20328 = ~n_20326 & ~n_20327;
assign n_20329 =  x_311 & ~n_20208;
assign n_20330 =  i_12 &  n_20208;
assign n_20331 = ~n_20329 & ~n_20330;
assign n_20332 =  x_311 & ~n_20331;
assign n_20333 = ~x_311 &  n_20331;
assign n_20334 = ~n_20332 & ~n_20333;
assign n_20335 =  x_310 & ~n_20208;
assign n_20336 =  i_11 &  n_20208;
assign n_20337 = ~n_20335 & ~n_20336;
assign n_20338 =  x_310 & ~n_20337;
assign n_20339 = ~x_310 &  n_20337;
assign n_20340 = ~n_20338 & ~n_20339;
assign n_20341 =  x_309 & ~n_20208;
assign n_20342 =  i_10 &  n_20208;
assign n_20343 = ~n_20341 & ~n_20342;
assign n_20344 =  x_309 & ~n_20343;
assign n_20345 = ~x_309 &  n_20343;
assign n_20346 = ~n_20344 & ~n_20345;
assign n_20347 =  x_308 & ~n_20208;
assign n_20348 =  i_9 &  n_20208;
assign n_20349 = ~n_20347 & ~n_20348;
assign n_20350 =  x_308 & ~n_20349;
assign n_20351 = ~x_308 &  n_20349;
assign n_20352 = ~n_20350 & ~n_20351;
assign n_20353 =  x_307 & ~n_20208;
assign n_20354 =  i_8 &  n_20208;
assign n_20355 = ~n_20353 & ~n_20354;
assign n_20356 =  x_307 & ~n_20355;
assign n_20357 = ~x_307 &  n_20355;
assign n_20358 = ~n_20356 & ~n_20357;
assign n_20359 =  x_306 & ~n_20208;
assign n_20360 =  i_7 &  n_20208;
assign n_20361 = ~n_20359 & ~n_20360;
assign n_20362 =  x_306 & ~n_20361;
assign n_20363 = ~x_306 &  n_20361;
assign n_20364 = ~n_20362 & ~n_20363;
assign n_20365 =  x_305 & ~n_20208;
assign n_20366 =  i_6 &  n_20208;
assign n_20367 = ~n_20365 & ~n_20366;
assign n_20368 =  x_305 & ~n_20367;
assign n_20369 = ~x_305 &  n_20367;
assign n_20370 = ~n_20368 & ~n_20369;
assign n_20371 =  x_304 & ~n_20208;
assign n_20372 =  i_5 &  n_20208;
assign n_20373 = ~n_20371 & ~n_20372;
assign n_20374 =  x_304 & ~n_20373;
assign n_20375 = ~x_304 &  n_20373;
assign n_20376 = ~n_20374 & ~n_20375;
assign n_20377 =  x_303 & ~n_20208;
assign n_20378 =  i_4 &  n_20208;
assign n_20379 = ~n_20377 & ~n_20378;
assign n_20380 =  x_303 & ~n_20379;
assign n_20381 = ~x_303 &  n_20379;
assign n_20382 = ~n_20380 & ~n_20381;
assign n_20383 =  x_302 & ~n_20208;
assign n_20384 =  i_3 &  n_20208;
assign n_20385 = ~n_20383 & ~n_20384;
assign n_20386 =  x_302 & ~n_20385;
assign n_20387 = ~x_302 &  n_20385;
assign n_20388 = ~n_20386 & ~n_20387;
assign n_20389 =  x_301 & ~n_20208;
assign n_20390 =  i_2 &  n_20208;
assign n_20391 = ~n_20389 & ~n_20390;
assign n_20392 =  x_301 & ~n_20391;
assign n_20393 = ~x_301 &  n_20391;
assign n_20394 = ~n_20392 & ~n_20393;
assign n_20395 =  x_300 & ~n_20208;
assign n_20396 =  i_1 &  n_20208;
assign n_20397 = ~n_20395 & ~n_20396;
assign n_20398 =  x_300 & ~n_20397;
assign n_20399 = ~x_300 &  n_20397;
assign n_20400 = ~n_20398 & ~n_20399;
assign n_20401 = ~x_40 &  n_2290;
assign n_20402 =  n_150 &  n_20401;
assign n_20403 =  n_554 &  n_20402;
assign n_20404 =  x_299 & ~n_20403;
assign n_20405 =  i_32 &  n_20403;
assign n_20406 = ~n_20404 & ~n_20405;
assign n_20407 =  x_299 & ~n_20406;
assign n_20408 = ~x_299 &  n_20406;
assign n_20409 = ~n_20407 & ~n_20408;
assign n_20410 =  x_298 & ~n_20403;
assign n_20411 =  i_31 &  n_20403;
assign n_20412 = ~n_20410 & ~n_20411;
assign n_20413 =  x_298 & ~n_20412;
assign n_20414 = ~x_298 &  n_20412;
assign n_20415 = ~n_20413 & ~n_20414;
assign n_20416 =  x_297 & ~n_20403;
assign n_20417 =  i_30 &  n_20403;
assign n_20418 = ~n_20416 & ~n_20417;
assign n_20419 =  x_297 & ~n_20418;
assign n_20420 = ~x_297 &  n_20418;
assign n_20421 = ~n_20419 & ~n_20420;
assign n_20422 =  x_296 & ~n_20403;
assign n_20423 =  i_29 &  n_20403;
assign n_20424 = ~n_20422 & ~n_20423;
assign n_20425 =  x_296 & ~n_20424;
assign n_20426 = ~x_296 &  n_20424;
assign n_20427 = ~n_20425 & ~n_20426;
assign n_20428 =  x_295 & ~n_20403;
assign n_20429 =  i_28 &  n_20403;
assign n_20430 = ~n_20428 & ~n_20429;
assign n_20431 =  x_295 & ~n_20430;
assign n_20432 = ~x_295 &  n_20430;
assign n_20433 = ~n_20431 & ~n_20432;
assign n_20434 =  x_294 & ~n_20403;
assign n_20435 =  i_27 &  n_20403;
assign n_20436 = ~n_20434 & ~n_20435;
assign n_20437 =  x_294 & ~n_20436;
assign n_20438 = ~x_294 &  n_20436;
assign n_20439 = ~n_20437 & ~n_20438;
assign n_20440 =  x_293 & ~n_20403;
assign n_20441 =  i_26 &  n_20403;
assign n_20442 = ~n_20440 & ~n_20441;
assign n_20443 =  x_293 & ~n_20442;
assign n_20444 = ~x_293 &  n_20442;
assign n_20445 = ~n_20443 & ~n_20444;
assign n_20446 =  x_292 & ~n_20403;
assign n_20447 =  i_25 &  n_20403;
assign n_20448 = ~n_20446 & ~n_20447;
assign n_20449 =  x_292 & ~n_20448;
assign n_20450 = ~x_292 &  n_20448;
assign n_20451 = ~n_20449 & ~n_20450;
assign n_20452 =  x_291 & ~n_20403;
assign n_20453 =  i_24 &  n_20403;
assign n_20454 = ~n_20452 & ~n_20453;
assign n_20455 =  x_291 & ~n_20454;
assign n_20456 = ~x_291 &  n_20454;
assign n_20457 = ~n_20455 & ~n_20456;
assign n_20458 =  x_290 & ~n_20403;
assign n_20459 =  i_23 &  n_20403;
assign n_20460 = ~n_20458 & ~n_20459;
assign n_20461 =  x_290 & ~n_20460;
assign n_20462 = ~x_290 &  n_20460;
assign n_20463 = ~n_20461 & ~n_20462;
assign n_20464 =  x_289 & ~n_20403;
assign n_20465 =  i_22 &  n_20403;
assign n_20466 = ~n_20464 & ~n_20465;
assign n_20467 =  x_289 & ~n_20466;
assign n_20468 = ~x_289 &  n_20466;
assign n_20469 = ~n_20467 & ~n_20468;
assign n_20470 =  x_288 & ~n_20403;
assign n_20471 =  i_21 &  n_20403;
assign n_20472 = ~n_20470 & ~n_20471;
assign n_20473 =  x_288 & ~n_20472;
assign n_20474 = ~x_288 &  n_20472;
assign n_20475 = ~n_20473 & ~n_20474;
assign n_20476 =  x_287 & ~n_20403;
assign n_20477 =  i_20 &  n_20403;
assign n_20478 = ~n_20476 & ~n_20477;
assign n_20479 =  x_287 & ~n_20478;
assign n_20480 = ~x_287 &  n_20478;
assign n_20481 = ~n_20479 & ~n_20480;
assign n_20482 =  x_286 & ~n_20403;
assign n_20483 =  i_19 &  n_20403;
assign n_20484 = ~n_20482 & ~n_20483;
assign n_20485 =  x_286 & ~n_20484;
assign n_20486 = ~x_286 &  n_20484;
assign n_20487 = ~n_20485 & ~n_20486;
assign n_20488 =  x_285 & ~n_20403;
assign n_20489 =  i_18 &  n_20403;
assign n_20490 = ~n_20488 & ~n_20489;
assign n_20491 =  x_285 & ~n_20490;
assign n_20492 = ~x_285 &  n_20490;
assign n_20493 = ~n_20491 & ~n_20492;
assign n_20494 =  x_284 & ~n_20403;
assign n_20495 =  i_17 &  n_20403;
assign n_20496 = ~n_20494 & ~n_20495;
assign n_20497 =  x_284 & ~n_20496;
assign n_20498 = ~x_284 &  n_20496;
assign n_20499 = ~n_20497 & ~n_20498;
assign n_20500 =  x_283 & ~n_20403;
assign n_20501 =  i_16 &  n_20403;
assign n_20502 = ~n_20500 & ~n_20501;
assign n_20503 =  x_283 & ~n_20502;
assign n_20504 = ~x_283 &  n_20502;
assign n_20505 = ~n_20503 & ~n_20504;
assign n_20506 =  x_282 & ~n_20403;
assign n_20507 =  i_15 &  n_20403;
assign n_20508 = ~n_20506 & ~n_20507;
assign n_20509 =  x_282 & ~n_20508;
assign n_20510 = ~x_282 &  n_20508;
assign n_20511 = ~n_20509 & ~n_20510;
assign n_20512 =  x_281 & ~n_20403;
assign n_20513 =  i_14 &  n_20403;
assign n_20514 = ~n_20512 & ~n_20513;
assign n_20515 =  x_281 & ~n_20514;
assign n_20516 = ~x_281 &  n_20514;
assign n_20517 = ~n_20515 & ~n_20516;
assign n_20518 =  x_280 & ~n_20403;
assign n_20519 =  i_13 &  n_20403;
assign n_20520 = ~n_20518 & ~n_20519;
assign n_20521 =  x_280 & ~n_20520;
assign n_20522 = ~x_280 &  n_20520;
assign n_20523 = ~n_20521 & ~n_20522;
assign n_20524 =  x_279 & ~n_20403;
assign n_20525 =  i_12 &  n_20403;
assign n_20526 = ~n_20524 & ~n_20525;
assign n_20527 =  x_279 & ~n_20526;
assign n_20528 = ~x_279 &  n_20526;
assign n_20529 = ~n_20527 & ~n_20528;
assign n_20530 =  x_278 & ~n_20403;
assign n_20531 =  i_11 &  n_20403;
assign n_20532 = ~n_20530 & ~n_20531;
assign n_20533 =  x_278 & ~n_20532;
assign n_20534 = ~x_278 &  n_20532;
assign n_20535 = ~n_20533 & ~n_20534;
assign n_20536 =  x_277 & ~n_20403;
assign n_20537 =  i_10 &  n_20403;
assign n_20538 = ~n_20536 & ~n_20537;
assign n_20539 =  x_277 & ~n_20538;
assign n_20540 = ~x_277 &  n_20538;
assign n_20541 = ~n_20539 & ~n_20540;
assign n_20542 =  x_276 & ~n_20403;
assign n_20543 =  i_9 &  n_20403;
assign n_20544 = ~n_20542 & ~n_20543;
assign n_20545 =  x_276 & ~n_20544;
assign n_20546 = ~x_276 &  n_20544;
assign n_20547 = ~n_20545 & ~n_20546;
assign n_20548 =  x_275 & ~n_20403;
assign n_20549 =  i_8 &  n_20403;
assign n_20550 = ~n_20548 & ~n_20549;
assign n_20551 =  x_275 & ~n_20550;
assign n_20552 = ~x_275 &  n_20550;
assign n_20553 = ~n_20551 & ~n_20552;
assign n_20554 =  x_274 & ~n_20403;
assign n_20555 =  i_7 &  n_20403;
assign n_20556 = ~n_20554 & ~n_20555;
assign n_20557 =  x_274 & ~n_20556;
assign n_20558 = ~x_274 &  n_20556;
assign n_20559 = ~n_20557 & ~n_20558;
assign n_20560 =  x_273 & ~n_20403;
assign n_20561 =  i_6 &  n_20403;
assign n_20562 = ~n_20560 & ~n_20561;
assign n_20563 =  x_273 & ~n_20562;
assign n_20564 = ~x_273 &  n_20562;
assign n_20565 = ~n_20563 & ~n_20564;
assign n_20566 =  x_272 & ~n_20403;
assign n_20567 =  i_5 &  n_20403;
assign n_20568 = ~n_20566 & ~n_20567;
assign n_20569 =  x_272 & ~n_20568;
assign n_20570 = ~x_272 &  n_20568;
assign n_20571 = ~n_20569 & ~n_20570;
assign n_20572 =  x_271 & ~n_20403;
assign n_20573 =  i_4 &  n_20403;
assign n_20574 = ~n_20572 & ~n_20573;
assign n_20575 =  x_271 & ~n_20574;
assign n_20576 = ~x_271 &  n_20574;
assign n_20577 = ~n_20575 & ~n_20576;
assign n_20578 =  x_270 & ~n_20403;
assign n_20579 =  i_3 &  n_20403;
assign n_20580 = ~n_20578 & ~n_20579;
assign n_20581 =  x_270 & ~n_20580;
assign n_20582 = ~x_270 &  n_20580;
assign n_20583 = ~n_20581 & ~n_20582;
assign n_20584 =  x_269 & ~n_20403;
assign n_20585 =  i_2 &  n_20403;
assign n_20586 = ~n_20584 & ~n_20585;
assign n_20587 =  x_269 & ~n_20586;
assign n_20588 = ~x_269 &  n_20586;
assign n_20589 = ~n_20587 & ~n_20588;
assign n_20590 =  x_268 & ~n_20403;
assign n_20591 =  i_1 &  n_20403;
assign n_20592 = ~n_20590 & ~n_20591;
assign n_20593 =  x_268 & ~n_20592;
assign n_20594 = ~x_268 &  n_20592;
assign n_20595 = ~n_20593 & ~n_20594;
assign n_20596 =  n_151 &  n_552;
assign n_20597 =  n_8365 &  n_20596;
assign n_20598 =  x_267 & ~n_20597;
assign n_20599 =  i_32 &  n_20597;
assign n_20600 = ~n_20598 & ~n_20599;
assign n_20601 =  x_267 & ~n_20600;
assign n_20602 = ~x_267 &  n_20600;
assign n_20603 = ~n_20601 & ~n_20602;
assign n_20604 =  x_266 & ~n_20597;
assign n_20605 =  i_31 &  n_20597;
assign n_20606 = ~n_20604 & ~n_20605;
assign n_20607 =  x_266 & ~n_20606;
assign n_20608 = ~x_266 &  n_20606;
assign n_20609 = ~n_20607 & ~n_20608;
assign n_20610 =  x_265 & ~n_20597;
assign n_20611 =  i_30 &  n_20597;
assign n_20612 = ~n_20610 & ~n_20611;
assign n_20613 =  x_265 & ~n_20612;
assign n_20614 = ~x_265 &  n_20612;
assign n_20615 = ~n_20613 & ~n_20614;
assign n_20616 =  x_264 & ~n_20597;
assign n_20617 =  i_29 &  n_20597;
assign n_20618 = ~n_20616 & ~n_20617;
assign n_20619 =  x_264 & ~n_20618;
assign n_20620 = ~x_264 &  n_20618;
assign n_20621 = ~n_20619 & ~n_20620;
assign n_20622 =  x_263 & ~n_20597;
assign n_20623 =  i_28 &  n_20597;
assign n_20624 = ~n_20622 & ~n_20623;
assign n_20625 =  x_263 & ~n_20624;
assign n_20626 = ~x_263 &  n_20624;
assign n_20627 = ~n_20625 & ~n_20626;
assign n_20628 =  x_262 & ~n_20597;
assign n_20629 =  i_27 &  n_20597;
assign n_20630 = ~n_20628 & ~n_20629;
assign n_20631 =  x_262 & ~n_20630;
assign n_20632 = ~x_262 &  n_20630;
assign n_20633 = ~n_20631 & ~n_20632;
assign n_20634 =  x_261 & ~n_20597;
assign n_20635 =  i_26 &  n_20597;
assign n_20636 = ~n_20634 & ~n_20635;
assign n_20637 =  x_261 & ~n_20636;
assign n_20638 = ~x_261 &  n_20636;
assign n_20639 = ~n_20637 & ~n_20638;
assign n_20640 =  x_260 & ~n_20597;
assign n_20641 =  i_25 &  n_20597;
assign n_20642 = ~n_20640 & ~n_20641;
assign n_20643 =  x_260 & ~n_20642;
assign n_20644 = ~x_260 &  n_20642;
assign n_20645 = ~n_20643 & ~n_20644;
assign n_20646 =  x_259 & ~n_20597;
assign n_20647 =  i_24 &  n_20597;
assign n_20648 = ~n_20646 & ~n_20647;
assign n_20649 =  x_259 & ~n_20648;
assign n_20650 = ~x_259 &  n_20648;
assign n_20651 = ~n_20649 & ~n_20650;
assign n_20652 =  x_258 & ~n_20597;
assign n_20653 =  i_23 &  n_20597;
assign n_20654 = ~n_20652 & ~n_20653;
assign n_20655 =  x_258 & ~n_20654;
assign n_20656 = ~x_258 &  n_20654;
assign n_20657 = ~n_20655 & ~n_20656;
assign n_20658 =  x_257 & ~n_20597;
assign n_20659 =  i_22 &  n_20597;
assign n_20660 = ~n_20658 & ~n_20659;
assign n_20661 =  x_257 & ~n_20660;
assign n_20662 = ~x_257 &  n_20660;
assign n_20663 = ~n_20661 & ~n_20662;
assign n_20664 =  x_256 & ~n_20597;
assign n_20665 =  i_21 &  n_20597;
assign n_20666 = ~n_20664 & ~n_20665;
assign n_20667 =  x_256 & ~n_20666;
assign n_20668 = ~x_256 &  n_20666;
assign n_20669 = ~n_20667 & ~n_20668;
assign n_20670 =  x_255 & ~n_20597;
assign n_20671 =  i_20 &  n_20597;
assign n_20672 = ~n_20670 & ~n_20671;
assign n_20673 =  x_255 & ~n_20672;
assign n_20674 = ~x_255 &  n_20672;
assign n_20675 = ~n_20673 & ~n_20674;
assign n_20676 =  x_254 & ~n_20597;
assign n_20677 =  i_19 &  n_20597;
assign n_20678 = ~n_20676 & ~n_20677;
assign n_20679 =  x_254 & ~n_20678;
assign n_20680 = ~x_254 &  n_20678;
assign n_20681 = ~n_20679 & ~n_20680;
assign n_20682 =  x_253 & ~n_20597;
assign n_20683 =  i_18 &  n_20597;
assign n_20684 = ~n_20682 & ~n_20683;
assign n_20685 =  x_253 & ~n_20684;
assign n_20686 = ~x_253 &  n_20684;
assign n_20687 = ~n_20685 & ~n_20686;
assign n_20688 =  x_252 & ~n_20597;
assign n_20689 =  i_17 &  n_20597;
assign n_20690 = ~n_20688 & ~n_20689;
assign n_20691 =  x_252 & ~n_20690;
assign n_20692 = ~x_252 &  n_20690;
assign n_20693 = ~n_20691 & ~n_20692;
assign n_20694 =  x_251 & ~n_20597;
assign n_20695 =  i_16 &  n_20597;
assign n_20696 = ~n_20694 & ~n_20695;
assign n_20697 =  x_251 & ~n_20696;
assign n_20698 = ~x_251 &  n_20696;
assign n_20699 = ~n_20697 & ~n_20698;
assign n_20700 =  x_250 & ~n_20597;
assign n_20701 =  i_15 &  n_20597;
assign n_20702 = ~n_20700 & ~n_20701;
assign n_20703 =  x_250 & ~n_20702;
assign n_20704 = ~x_250 &  n_20702;
assign n_20705 = ~n_20703 & ~n_20704;
assign n_20706 =  x_249 & ~n_20597;
assign n_20707 =  i_14 &  n_20597;
assign n_20708 = ~n_20706 & ~n_20707;
assign n_20709 =  x_249 & ~n_20708;
assign n_20710 = ~x_249 &  n_20708;
assign n_20711 = ~n_20709 & ~n_20710;
assign n_20712 =  x_248 & ~n_20597;
assign n_20713 =  i_13 &  n_20597;
assign n_20714 = ~n_20712 & ~n_20713;
assign n_20715 =  x_248 & ~n_20714;
assign n_20716 = ~x_248 &  n_20714;
assign n_20717 = ~n_20715 & ~n_20716;
assign n_20718 =  x_247 & ~n_20597;
assign n_20719 =  i_12 &  n_20597;
assign n_20720 = ~n_20718 & ~n_20719;
assign n_20721 =  x_247 & ~n_20720;
assign n_20722 = ~x_247 &  n_20720;
assign n_20723 = ~n_20721 & ~n_20722;
assign n_20724 =  x_246 & ~n_20597;
assign n_20725 =  i_11 &  n_20597;
assign n_20726 = ~n_20724 & ~n_20725;
assign n_20727 =  x_246 & ~n_20726;
assign n_20728 = ~x_246 &  n_20726;
assign n_20729 = ~n_20727 & ~n_20728;
assign n_20730 =  x_245 & ~n_20597;
assign n_20731 =  i_10 &  n_20597;
assign n_20732 = ~n_20730 & ~n_20731;
assign n_20733 =  x_245 & ~n_20732;
assign n_20734 = ~x_245 &  n_20732;
assign n_20735 = ~n_20733 & ~n_20734;
assign n_20736 =  x_244 & ~n_20597;
assign n_20737 =  i_9 &  n_20597;
assign n_20738 = ~n_20736 & ~n_20737;
assign n_20739 =  x_244 & ~n_20738;
assign n_20740 = ~x_244 &  n_20738;
assign n_20741 = ~n_20739 & ~n_20740;
assign n_20742 =  x_243 & ~n_20597;
assign n_20743 =  i_8 &  n_20597;
assign n_20744 = ~n_20742 & ~n_20743;
assign n_20745 =  x_243 & ~n_20744;
assign n_20746 = ~x_243 &  n_20744;
assign n_20747 = ~n_20745 & ~n_20746;
assign n_20748 =  x_242 & ~n_20597;
assign n_20749 =  i_7 &  n_20597;
assign n_20750 = ~n_20748 & ~n_20749;
assign n_20751 =  x_242 & ~n_20750;
assign n_20752 = ~x_242 &  n_20750;
assign n_20753 = ~n_20751 & ~n_20752;
assign n_20754 =  x_241 & ~n_20597;
assign n_20755 =  i_6 &  n_20597;
assign n_20756 = ~n_20754 & ~n_20755;
assign n_20757 =  x_241 & ~n_20756;
assign n_20758 = ~x_241 &  n_20756;
assign n_20759 = ~n_20757 & ~n_20758;
assign n_20760 =  x_240 & ~n_20597;
assign n_20761 =  i_5 &  n_20597;
assign n_20762 = ~n_20760 & ~n_20761;
assign n_20763 =  x_240 & ~n_20762;
assign n_20764 = ~x_240 &  n_20762;
assign n_20765 = ~n_20763 & ~n_20764;
assign n_20766 =  x_239 & ~n_20597;
assign n_20767 =  i_4 &  n_20597;
assign n_20768 = ~n_20766 & ~n_20767;
assign n_20769 =  x_239 & ~n_20768;
assign n_20770 = ~x_239 &  n_20768;
assign n_20771 = ~n_20769 & ~n_20770;
assign n_20772 =  x_238 & ~n_20597;
assign n_20773 =  i_3 &  n_20597;
assign n_20774 = ~n_20772 & ~n_20773;
assign n_20775 =  x_238 & ~n_20774;
assign n_20776 = ~x_238 &  n_20774;
assign n_20777 = ~n_20775 & ~n_20776;
assign n_20778 =  x_237 & ~n_20597;
assign n_20779 =  i_2 &  n_20597;
assign n_20780 = ~n_20778 & ~n_20779;
assign n_20781 =  x_237 & ~n_20780;
assign n_20782 = ~x_237 &  n_20780;
assign n_20783 = ~n_20781 & ~n_20782;
assign n_20784 =  x_236 & ~n_20597;
assign n_20785 =  i_1 &  n_20597;
assign n_20786 = ~n_20784 & ~n_20785;
assign n_20787 =  x_236 & ~n_20786;
assign n_20788 = ~x_236 &  n_20786;
assign n_20789 = ~n_20787 & ~n_20788;
assign n_20790 =  n_151 &  n_9884;
assign n_20791 =  n_20790 &  n_3615;
assign n_20792 =  x_235 & ~n_20791;
assign n_20793 =  i_32 &  n_20791;
assign n_20794 = ~n_20792 & ~n_20793;
assign n_20795 =  x_235 & ~n_20794;
assign n_20796 = ~x_235 &  n_20794;
assign n_20797 = ~n_20795 & ~n_20796;
assign n_20798 =  x_234 & ~n_20791;
assign n_20799 =  i_31 &  n_20791;
assign n_20800 = ~n_20798 & ~n_20799;
assign n_20801 =  x_234 & ~n_20800;
assign n_20802 = ~x_234 &  n_20800;
assign n_20803 = ~n_20801 & ~n_20802;
assign n_20804 =  x_233 & ~n_20791;
assign n_20805 =  i_30 &  n_20791;
assign n_20806 = ~n_20804 & ~n_20805;
assign n_20807 =  x_233 & ~n_20806;
assign n_20808 = ~x_233 &  n_20806;
assign n_20809 = ~n_20807 & ~n_20808;
assign n_20810 =  x_232 & ~n_20791;
assign n_20811 =  i_29 &  n_20791;
assign n_20812 = ~n_20810 & ~n_20811;
assign n_20813 =  x_232 & ~n_20812;
assign n_20814 = ~x_232 &  n_20812;
assign n_20815 = ~n_20813 & ~n_20814;
assign n_20816 =  x_231 & ~n_20791;
assign n_20817 =  i_28 &  n_20791;
assign n_20818 = ~n_20816 & ~n_20817;
assign n_20819 =  x_231 & ~n_20818;
assign n_20820 = ~x_231 &  n_20818;
assign n_20821 = ~n_20819 & ~n_20820;
assign n_20822 =  x_230 & ~n_20791;
assign n_20823 =  i_27 &  n_20791;
assign n_20824 = ~n_20822 & ~n_20823;
assign n_20825 =  x_230 & ~n_20824;
assign n_20826 = ~x_230 &  n_20824;
assign n_20827 = ~n_20825 & ~n_20826;
assign n_20828 =  x_229 & ~n_20791;
assign n_20829 =  i_26 &  n_20791;
assign n_20830 = ~n_20828 & ~n_20829;
assign n_20831 =  x_229 & ~n_20830;
assign n_20832 = ~x_229 &  n_20830;
assign n_20833 = ~n_20831 & ~n_20832;
assign n_20834 =  x_228 & ~n_20791;
assign n_20835 =  i_25 &  n_20791;
assign n_20836 = ~n_20834 & ~n_20835;
assign n_20837 =  x_228 & ~n_20836;
assign n_20838 = ~x_228 &  n_20836;
assign n_20839 = ~n_20837 & ~n_20838;
assign n_20840 =  x_227 & ~n_20791;
assign n_20841 =  i_24 &  n_20791;
assign n_20842 = ~n_20840 & ~n_20841;
assign n_20843 =  x_227 & ~n_20842;
assign n_20844 = ~x_227 &  n_20842;
assign n_20845 = ~n_20843 & ~n_20844;
assign n_20846 =  x_226 & ~n_20791;
assign n_20847 =  i_23 &  n_20791;
assign n_20848 = ~n_20846 & ~n_20847;
assign n_20849 =  x_226 & ~n_20848;
assign n_20850 = ~x_226 &  n_20848;
assign n_20851 = ~n_20849 & ~n_20850;
assign n_20852 =  x_225 & ~n_20791;
assign n_20853 =  i_22 &  n_20791;
assign n_20854 = ~n_20852 & ~n_20853;
assign n_20855 =  x_225 & ~n_20854;
assign n_20856 = ~x_225 &  n_20854;
assign n_20857 = ~n_20855 & ~n_20856;
assign n_20858 =  x_224 & ~n_20791;
assign n_20859 =  i_21 &  n_20791;
assign n_20860 = ~n_20858 & ~n_20859;
assign n_20861 =  x_224 & ~n_20860;
assign n_20862 = ~x_224 &  n_20860;
assign n_20863 = ~n_20861 & ~n_20862;
assign n_20864 =  x_223 & ~n_20791;
assign n_20865 =  i_20 &  n_20791;
assign n_20866 = ~n_20864 & ~n_20865;
assign n_20867 =  x_223 & ~n_20866;
assign n_20868 = ~x_223 &  n_20866;
assign n_20869 = ~n_20867 & ~n_20868;
assign n_20870 =  x_222 & ~n_20791;
assign n_20871 =  i_19 &  n_20791;
assign n_20872 = ~n_20870 & ~n_20871;
assign n_20873 =  x_222 & ~n_20872;
assign n_20874 = ~x_222 &  n_20872;
assign n_20875 = ~n_20873 & ~n_20874;
assign n_20876 =  x_221 & ~n_20791;
assign n_20877 =  i_18 &  n_20791;
assign n_20878 = ~n_20876 & ~n_20877;
assign n_20879 =  x_221 & ~n_20878;
assign n_20880 = ~x_221 &  n_20878;
assign n_20881 = ~n_20879 & ~n_20880;
assign n_20882 =  x_220 & ~n_20791;
assign n_20883 =  i_17 &  n_20791;
assign n_20884 = ~n_20882 & ~n_20883;
assign n_20885 =  x_220 & ~n_20884;
assign n_20886 = ~x_220 &  n_20884;
assign n_20887 = ~n_20885 & ~n_20886;
assign n_20888 =  x_219 & ~n_20791;
assign n_20889 =  i_16 &  n_20791;
assign n_20890 = ~n_20888 & ~n_20889;
assign n_20891 =  x_219 & ~n_20890;
assign n_20892 = ~x_219 &  n_20890;
assign n_20893 = ~n_20891 & ~n_20892;
assign n_20894 =  x_218 & ~n_20791;
assign n_20895 =  i_15 &  n_20791;
assign n_20896 = ~n_20894 & ~n_20895;
assign n_20897 =  x_218 & ~n_20896;
assign n_20898 = ~x_218 &  n_20896;
assign n_20899 = ~n_20897 & ~n_20898;
assign n_20900 =  x_217 & ~n_20791;
assign n_20901 =  i_14 &  n_20791;
assign n_20902 = ~n_20900 & ~n_20901;
assign n_20903 =  x_217 & ~n_20902;
assign n_20904 = ~x_217 &  n_20902;
assign n_20905 = ~n_20903 & ~n_20904;
assign n_20906 =  x_216 & ~n_20791;
assign n_20907 =  i_13 &  n_20791;
assign n_20908 = ~n_20906 & ~n_20907;
assign n_20909 =  x_216 & ~n_20908;
assign n_20910 = ~x_216 &  n_20908;
assign n_20911 = ~n_20909 & ~n_20910;
assign n_20912 =  x_215 & ~n_20791;
assign n_20913 =  i_12 &  n_20791;
assign n_20914 = ~n_20912 & ~n_20913;
assign n_20915 =  x_215 & ~n_20914;
assign n_20916 = ~x_215 &  n_20914;
assign n_20917 = ~n_20915 & ~n_20916;
assign n_20918 =  x_214 & ~n_20791;
assign n_20919 =  i_11 &  n_20791;
assign n_20920 = ~n_20918 & ~n_20919;
assign n_20921 =  x_214 & ~n_20920;
assign n_20922 = ~x_214 &  n_20920;
assign n_20923 = ~n_20921 & ~n_20922;
assign n_20924 =  x_213 & ~n_20791;
assign n_20925 =  i_10 &  n_20791;
assign n_20926 = ~n_20924 & ~n_20925;
assign n_20927 =  x_213 & ~n_20926;
assign n_20928 = ~x_213 &  n_20926;
assign n_20929 = ~n_20927 & ~n_20928;
assign n_20930 =  x_212 & ~n_20791;
assign n_20931 =  i_9 &  n_20791;
assign n_20932 = ~n_20930 & ~n_20931;
assign n_20933 =  x_212 & ~n_20932;
assign n_20934 = ~x_212 &  n_20932;
assign n_20935 = ~n_20933 & ~n_20934;
assign n_20936 =  x_211 & ~n_20791;
assign n_20937 =  i_8 &  n_20791;
assign n_20938 = ~n_20936 & ~n_20937;
assign n_20939 =  x_211 & ~n_20938;
assign n_20940 = ~x_211 &  n_20938;
assign n_20941 = ~n_20939 & ~n_20940;
assign n_20942 =  x_210 & ~n_20791;
assign n_20943 =  i_7 &  n_20791;
assign n_20944 = ~n_20942 & ~n_20943;
assign n_20945 =  x_210 & ~n_20944;
assign n_20946 = ~x_210 &  n_20944;
assign n_20947 = ~n_20945 & ~n_20946;
assign n_20948 =  x_209 & ~n_20791;
assign n_20949 =  i_6 &  n_20791;
assign n_20950 = ~n_20948 & ~n_20949;
assign n_20951 =  x_209 & ~n_20950;
assign n_20952 = ~x_209 &  n_20950;
assign n_20953 = ~n_20951 & ~n_20952;
assign n_20954 =  x_208 & ~n_20791;
assign n_20955 =  i_5 &  n_20791;
assign n_20956 = ~n_20954 & ~n_20955;
assign n_20957 =  x_208 & ~n_20956;
assign n_20958 = ~x_208 &  n_20956;
assign n_20959 = ~n_20957 & ~n_20958;
assign n_20960 =  x_207 & ~n_20791;
assign n_20961 =  i_4 &  n_20791;
assign n_20962 = ~n_20960 & ~n_20961;
assign n_20963 =  x_207 & ~n_20962;
assign n_20964 = ~x_207 &  n_20962;
assign n_20965 = ~n_20963 & ~n_20964;
assign n_20966 =  x_206 & ~n_20791;
assign n_20967 =  i_3 &  n_20791;
assign n_20968 = ~n_20966 & ~n_20967;
assign n_20969 =  x_206 & ~n_20968;
assign n_20970 = ~x_206 &  n_20968;
assign n_20971 = ~n_20969 & ~n_20970;
assign n_20972 =  x_205 & ~n_20791;
assign n_20973 =  i_2 &  n_20791;
assign n_20974 = ~n_20972 & ~n_20973;
assign n_20975 =  x_205 & ~n_20974;
assign n_20976 = ~x_205 &  n_20974;
assign n_20977 = ~n_20975 & ~n_20976;
assign n_20978 =  x_204 & ~n_20791;
assign n_20979 =  i_1 &  n_20791;
assign n_20980 = ~n_20978 & ~n_20979;
assign n_20981 =  x_204 & ~n_20980;
assign n_20982 = ~x_204 &  n_20980;
assign n_20983 = ~n_20981 & ~n_20982;
assign n_20984 =  n_553 &  n_1699;
assign n_20985 =  x_43 &  n_20984;
assign n_20986 =  x_203 & ~n_20985;
assign n_20987 =  x_491 &  n_20985;
assign n_20988 = ~n_20986 & ~n_20987;
assign n_20989 =  x_203 & ~n_20988;
assign n_20990 = ~x_203 &  n_20988;
assign n_20991 = ~n_20989 & ~n_20990;
assign n_20992 =  x_202 & ~n_20985;
assign n_20993 =  x_490 &  n_20985;
assign n_20994 = ~n_20992 & ~n_20993;
assign n_20995 =  x_202 & ~n_20994;
assign n_20996 = ~x_202 &  n_20994;
assign n_20997 = ~n_20995 & ~n_20996;
assign n_20998 =  x_201 & ~n_20985;
assign n_20999 =  x_489 &  n_20985;
assign n_21000 = ~n_20998 & ~n_20999;
assign n_21001 =  x_201 & ~n_21000;
assign n_21002 = ~x_201 &  n_21000;
assign n_21003 = ~n_21001 & ~n_21002;
assign n_21004 =  x_200 & ~n_20985;
assign n_21005 =  x_488 &  n_20985;
assign n_21006 = ~n_21004 & ~n_21005;
assign n_21007 =  x_200 & ~n_21006;
assign n_21008 = ~x_200 &  n_21006;
assign n_21009 = ~n_21007 & ~n_21008;
assign n_21010 =  x_199 & ~n_20985;
assign n_21011 =  x_487 &  n_20985;
assign n_21012 = ~n_21010 & ~n_21011;
assign n_21013 =  x_199 & ~n_21012;
assign n_21014 = ~x_199 &  n_21012;
assign n_21015 = ~n_21013 & ~n_21014;
assign n_21016 =  x_198 & ~n_20985;
assign n_21017 =  x_486 &  n_20985;
assign n_21018 = ~n_21016 & ~n_21017;
assign n_21019 =  x_198 & ~n_21018;
assign n_21020 = ~x_198 &  n_21018;
assign n_21021 = ~n_21019 & ~n_21020;
assign n_21022 =  x_197 & ~n_20985;
assign n_21023 =  x_485 &  n_20985;
assign n_21024 = ~n_21022 & ~n_21023;
assign n_21025 =  x_197 & ~n_21024;
assign n_21026 = ~x_197 &  n_21024;
assign n_21027 = ~n_21025 & ~n_21026;
assign n_21028 =  x_196 & ~n_20985;
assign n_21029 =  x_484 &  n_20985;
assign n_21030 = ~n_21028 & ~n_21029;
assign n_21031 =  x_196 & ~n_21030;
assign n_21032 = ~x_196 &  n_21030;
assign n_21033 = ~n_21031 & ~n_21032;
assign n_21034 =  x_195 & ~n_20985;
assign n_21035 =  x_483 &  n_20985;
assign n_21036 = ~n_21034 & ~n_21035;
assign n_21037 =  x_195 & ~n_21036;
assign n_21038 = ~x_195 &  n_21036;
assign n_21039 = ~n_21037 & ~n_21038;
assign n_21040 =  x_194 & ~n_20985;
assign n_21041 =  x_482 &  n_20985;
assign n_21042 = ~n_21040 & ~n_21041;
assign n_21043 =  x_194 & ~n_21042;
assign n_21044 = ~x_194 &  n_21042;
assign n_21045 = ~n_21043 & ~n_21044;
assign n_21046 =  x_193 & ~n_20985;
assign n_21047 =  x_481 &  n_20985;
assign n_21048 = ~n_21046 & ~n_21047;
assign n_21049 =  x_193 & ~n_21048;
assign n_21050 = ~x_193 &  n_21048;
assign n_21051 = ~n_21049 & ~n_21050;
assign n_21052 =  x_192 & ~n_20985;
assign n_21053 =  x_480 &  n_20985;
assign n_21054 = ~n_21052 & ~n_21053;
assign n_21055 =  x_192 & ~n_21054;
assign n_21056 = ~x_192 &  n_21054;
assign n_21057 = ~n_21055 & ~n_21056;
assign n_21058 =  x_191 & ~n_20985;
assign n_21059 =  x_479 &  n_20985;
assign n_21060 = ~n_21058 & ~n_21059;
assign n_21061 =  x_191 & ~n_21060;
assign n_21062 = ~x_191 &  n_21060;
assign n_21063 = ~n_21061 & ~n_21062;
assign n_21064 =  x_190 & ~n_20985;
assign n_21065 =  x_478 &  n_20985;
assign n_21066 = ~n_21064 & ~n_21065;
assign n_21067 =  x_190 & ~n_21066;
assign n_21068 = ~x_190 &  n_21066;
assign n_21069 = ~n_21067 & ~n_21068;
assign n_21070 =  x_189 & ~n_20985;
assign n_21071 =  x_477 &  n_20985;
assign n_21072 = ~n_21070 & ~n_21071;
assign n_21073 =  x_189 & ~n_21072;
assign n_21074 = ~x_189 &  n_21072;
assign n_21075 = ~n_21073 & ~n_21074;
assign n_21076 =  x_188 & ~n_20985;
assign n_21077 =  x_476 &  n_20985;
assign n_21078 = ~n_21076 & ~n_21077;
assign n_21079 =  x_188 & ~n_21078;
assign n_21080 = ~x_188 &  n_21078;
assign n_21081 = ~n_21079 & ~n_21080;
assign n_21082 =  x_187 & ~n_20985;
assign n_21083 =  x_475 &  n_20985;
assign n_21084 = ~n_21082 & ~n_21083;
assign n_21085 =  x_187 & ~n_21084;
assign n_21086 = ~x_187 &  n_21084;
assign n_21087 = ~n_21085 & ~n_21086;
assign n_21088 =  x_186 & ~n_20985;
assign n_21089 =  x_474 &  n_20985;
assign n_21090 = ~n_21088 & ~n_21089;
assign n_21091 =  x_186 & ~n_21090;
assign n_21092 = ~x_186 &  n_21090;
assign n_21093 = ~n_21091 & ~n_21092;
assign n_21094 =  x_185 & ~n_20985;
assign n_21095 =  x_473 &  n_20985;
assign n_21096 = ~n_21094 & ~n_21095;
assign n_21097 =  x_185 & ~n_21096;
assign n_21098 = ~x_185 &  n_21096;
assign n_21099 = ~n_21097 & ~n_21098;
assign n_21100 =  x_184 & ~n_20985;
assign n_21101 =  x_472 &  n_20985;
assign n_21102 = ~n_21100 & ~n_21101;
assign n_21103 =  x_184 & ~n_21102;
assign n_21104 = ~x_184 &  n_21102;
assign n_21105 = ~n_21103 & ~n_21104;
assign n_21106 =  x_183 & ~n_20985;
assign n_21107 =  x_471 &  n_20985;
assign n_21108 = ~n_21106 & ~n_21107;
assign n_21109 =  x_183 & ~n_21108;
assign n_21110 = ~x_183 &  n_21108;
assign n_21111 = ~n_21109 & ~n_21110;
assign n_21112 =  x_182 & ~n_20985;
assign n_21113 =  x_470 &  n_20985;
assign n_21114 = ~n_21112 & ~n_21113;
assign n_21115 =  x_182 & ~n_21114;
assign n_21116 = ~x_182 &  n_21114;
assign n_21117 = ~n_21115 & ~n_21116;
assign n_21118 =  x_181 & ~n_20985;
assign n_21119 =  x_469 &  n_20985;
assign n_21120 = ~n_21118 & ~n_21119;
assign n_21121 =  x_181 & ~n_21120;
assign n_21122 = ~x_181 &  n_21120;
assign n_21123 = ~n_21121 & ~n_21122;
assign n_21124 =  x_180 & ~n_20985;
assign n_21125 =  x_468 &  n_20985;
assign n_21126 = ~n_21124 & ~n_21125;
assign n_21127 =  x_180 & ~n_21126;
assign n_21128 = ~x_180 &  n_21126;
assign n_21129 = ~n_21127 & ~n_21128;
assign n_21130 =  x_179 & ~n_20985;
assign n_21131 =  x_467 &  n_20985;
assign n_21132 = ~n_21130 & ~n_21131;
assign n_21133 =  x_179 & ~n_21132;
assign n_21134 = ~x_179 &  n_21132;
assign n_21135 = ~n_21133 & ~n_21134;
assign n_21136 =  x_178 & ~n_20985;
assign n_21137 =  x_466 &  n_20985;
assign n_21138 = ~n_21136 & ~n_21137;
assign n_21139 =  x_178 & ~n_21138;
assign n_21140 = ~x_178 &  n_21138;
assign n_21141 = ~n_21139 & ~n_21140;
assign n_21142 =  x_177 & ~n_20985;
assign n_21143 =  x_465 &  n_20985;
assign n_21144 = ~n_21142 & ~n_21143;
assign n_21145 =  x_177 & ~n_21144;
assign n_21146 = ~x_177 &  n_21144;
assign n_21147 = ~n_21145 & ~n_21146;
assign n_21148 =  x_176 & ~n_20985;
assign n_21149 =  x_464 &  n_20985;
assign n_21150 = ~n_21148 & ~n_21149;
assign n_21151 =  x_176 & ~n_21150;
assign n_21152 = ~x_176 &  n_21150;
assign n_21153 = ~n_21151 & ~n_21152;
assign n_21154 =  x_175 & ~n_20985;
assign n_21155 =  x_463 &  n_20985;
assign n_21156 = ~n_21154 & ~n_21155;
assign n_21157 =  x_175 & ~n_21156;
assign n_21158 = ~x_175 &  n_21156;
assign n_21159 = ~n_21157 & ~n_21158;
assign n_21160 =  x_174 & ~n_20985;
assign n_21161 =  x_462 &  n_20985;
assign n_21162 = ~n_21160 & ~n_21161;
assign n_21163 =  x_174 & ~n_21162;
assign n_21164 = ~x_174 &  n_21162;
assign n_21165 = ~n_21163 & ~n_21164;
assign n_21166 =  x_173 & ~n_20985;
assign n_21167 =  x_461 &  n_20985;
assign n_21168 = ~n_21166 & ~n_21167;
assign n_21169 =  x_173 & ~n_21168;
assign n_21170 = ~x_173 &  n_21168;
assign n_21171 = ~n_21169 & ~n_21170;
assign n_21172 =  x_172 & ~n_20985;
assign n_21173 =  x_460 &  n_20985;
assign n_21174 = ~n_21172 & ~n_21173;
assign n_21175 =  x_172 & ~n_21174;
assign n_21176 = ~x_172 &  n_21174;
assign n_21177 = ~n_21175 & ~n_21176;
assign n_21178 =  n_14 &  n_13866;
assign n_21179 =  x_171 & ~n_21178;
assign n_21180 =  i_32 &  n_21178;
assign n_21181 = ~n_21179 & ~n_21180;
assign n_21182 =  x_171 & ~n_21181;
assign n_21183 = ~x_171 &  n_21181;
assign n_21184 = ~n_21182 & ~n_21183;
assign n_21185 =  x_170 & ~n_21178;
assign n_21186 =  i_31 &  n_21178;
assign n_21187 = ~n_21185 & ~n_21186;
assign n_21188 =  x_170 & ~n_21187;
assign n_21189 = ~x_170 &  n_21187;
assign n_21190 = ~n_21188 & ~n_21189;
assign n_21191 =  x_169 & ~n_21178;
assign n_21192 =  i_30 &  n_21178;
assign n_21193 = ~n_21191 & ~n_21192;
assign n_21194 =  x_169 & ~n_21193;
assign n_21195 = ~x_169 &  n_21193;
assign n_21196 = ~n_21194 & ~n_21195;
assign n_21197 =  x_168 & ~n_21178;
assign n_21198 =  i_29 &  n_21178;
assign n_21199 = ~n_21197 & ~n_21198;
assign n_21200 =  x_168 & ~n_21199;
assign n_21201 = ~x_168 &  n_21199;
assign n_21202 = ~n_21200 & ~n_21201;
assign n_21203 =  x_167 & ~n_21178;
assign n_21204 =  i_28 &  n_21178;
assign n_21205 = ~n_21203 & ~n_21204;
assign n_21206 =  x_167 & ~n_21205;
assign n_21207 = ~x_167 &  n_21205;
assign n_21208 = ~n_21206 & ~n_21207;
assign n_21209 =  x_166 & ~n_21178;
assign n_21210 =  i_27 &  n_21178;
assign n_21211 = ~n_21209 & ~n_21210;
assign n_21212 =  x_166 & ~n_21211;
assign n_21213 = ~x_166 &  n_21211;
assign n_21214 = ~n_21212 & ~n_21213;
assign n_21215 =  x_165 & ~n_21178;
assign n_21216 =  i_26 &  n_21178;
assign n_21217 = ~n_21215 & ~n_21216;
assign n_21218 =  x_165 & ~n_21217;
assign n_21219 = ~x_165 &  n_21217;
assign n_21220 = ~n_21218 & ~n_21219;
assign n_21221 =  x_164 & ~n_21178;
assign n_21222 =  i_25 &  n_21178;
assign n_21223 = ~n_21221 & ~n_21222;
assign n_21224 =  x_164 & ~n_21223;
assign n_21225 = ~x_164 &  n_21223;
assign n_21226 = ~n_21224 & ~n_21225;
assign n_21227 =  x_163 & ~n_21178;
assign n_21228 =  i_24 &  n_21178;
assign n_21229 = ~n_21227 & ~n_21228;
assign n_21230 =  x_163 & ~n_21229;
assign n_21231 = ~x_163 &  n_21229;
assign n_21232 = ~n_21230 & ~n_21231;
assign n_21233 =  x_162 & ~n_21178;
assign n_21234 =  i_23 &  n_21178;
assign n_21235 = ~n_21233 & ~n_21234;
assign n_21236 =  x_162 & ~n_21235;
assign n_21237 = ~x_162 &  n_21235;
assign n_21238 = ~n_21236 & ~n_21237;
assign n_21239 =  x_161 & ~n_21178;
assign n_21240 =  i_22 &  n_21178;
assign n_21241 = ~n_21239 & ~n_21240;
assign n_21242 =  x_161 & ~n_21241;
assign n_21243 = ~x_161 &  n_21241;
assign n_21244 = ~n_21242 & ~n_21243;
assign n_21245 =  x_160 & ~n_21178;
assign n_21246 =  i_21 &  n_21178;
assign n_21247 = ~n_21245 & ~n_21246;
assign n_21248 =  x_160 & ~n_21247;
assign n_21249 = ~x_160 &  n_21247;
assign n_21250 = ~n_21248 & ~n_21249;
assign n_21251 =  x_159 & ~n_21178;
assign n_21252 =  i_20 &  n_21178;
assign n_21253 = ~n_21251 & ~n_21252;
assign n_21254 =  x_159 & ~n_21253;
assign n_21255 = ~x_159 &  n_21253;
assign n_21256 = ~n_21254 & ~n_21255;
assign n_21257 =  x_158 & ~n_21178;
assign n_21258 =  i_19 &  n_21178;
assign n_21259 = ~n_21257 & ~n_21258;
assign n_21260 =  x_158 & ~n_21259;
assign n_21261 = ~x_158 &  n_21259;
assign n_21262 = ~n_21260 & ~n_21261;
assign n_21263 =  x_157 & ~n_21178;
assign n_21264 =  i_18 &  n_21178;
assign n_21265 = ~n_21263 & ~n_21264;
assign n_21266 =  x_157 & ~n_21265;
assign n_21267 = ~x_157 &  n_21265;
assign n_21268 = ~n_21266 & ~n_21267;
assign n_21269 =  x_156 & ~n_21178;
assign n_21270 =  i_17 &  n_21178;
assign n_21271 = ~n_21269 & ~n_21270;
assign n_21272 =  x_156 & ~n_21271;
assign n_21273 = ~x_156 &  n_21271;
assign n_21274 = ~n_21272 & ~n_21273;
assign n_21275 =  x_155 & ~n_21178;
assign n_21276 =  i_16 &  n_21178;
assign n_21277 = ~n_21275 & ~n_21276;
assign n_21278 =  x_155 & ~n_21277;
assign n_21279 = ~x_155 &  n_21277;
assign n_21280 = ~n_21278 & ~n_21279;
assign n_21281 =  x_154 & ~n_21178;
assign n_21282 =  i_15 &  n_21178;
assign n_21283 = ~n_21281 & ~n_21282;
assign n_21284 =  x_154 & ~n_21283;
assign n_21285 = ~x_154 &  n_21283;
assign n_21286 = ~n_21284 & ~n_21285;
assign n_21287 =  x_153 & ~n_21178;
assign n_21288 =  i_14 &  n_21178;
assign n_21289 = ~n_21287 & ~n_21288;
assign n_21290 =  x_153 & ~n_21289;
assign n_21291 = ~x_153 &  n_21289;
assign n_21292 = ~n_21290 & ~n_21291;
assign n_21293 =  x_152 & ~n_21178;
assign n_21294 =  i_13 &  n_21178;
assign n_21295 = ~n_21293 & ~n_21294;
assign n_21296 =  x_152 & ~n_21295;
assign n_21297 = ~x_152 &  n_21295;
assign n_21298 = ~n_21296 & ~n_21297;
assign n_21299 =  x_151 & ~n_21178;
assign n_21300 =  i_12 &  n_21178;
assign n_21301 = ~n_21299 & ~n_21300;
assign n_21302 =  x_151 & ~n_21301;
assign n_21303 = ~x_151 &  n_21301;
assign n_21304 = ~n_21302 & ~n_21303;
assign n_21305 =  x_150 & ~n_21178;
assign n_21306 =  i_11 &  n_21178;
assign n_21307 = ~n_21305 & ~n_21306;
assign n_21308 =  x_150 & ~n_21307;
assign n_21309 = ~x_150 &  n_21307;
assign n_21310 = ~n_21308 & ~n_21309;
assign n_21311 =  x_149 & ~n_21178;
assign n_21312 =  i_10 &  n_21178;
assign n_21313 = ~n_21311 & ~n_21312;
assign n_21314 =  x_149 & ~n_21313;
assign n_21315 = ~x_149 &  n_21313;
assign n_21316 = ~n_21314 & ~n_21315;
assign n_21317 =  x_148 & ~n_21178;
assign n_21318 =  i_9 &  n_21178;
assign n_21319 = ~n_21317 & ~n_21318;
assign n_21320 =  x_148 & ~n_21319;
assign n_21321 = ~x_148 &  n_21319;
assign n_21322 = ~n_21320 & ~n_21321;
assign n_21323 =  x_147 & ~n_21178;
assign n_21324 =  i_8 &  n_21178;
assign n_21325 = ~n_21323 & ~n_21324;
assign n_21326 =  x_147 & ~n_21325;
assign n_21327 = ~x_147 &  n_21325;
assign n_21328 = ~n_21326 & ~n_21327;
assign n_21329 =  x_146 & ~n_21178;
assign n_21330 =  i_7 &  n_21178;
assign n_21331 = ~n_21329 & ~n_21330;
assign n_21332 =  x_146 & ~n_21331;
assign n_21333 = ~x_146 &  n_21331;
assign n_21334 = ~n_21332 & ~n_21333;
assign n_21335 =  x_145 & ~n_21178;
assign n_21336 =  i_6 &  n_21178;
assign n_21337 = ~n_21335 & ~n_21336;
assign n_21338 =  x_145 & ~n_21337;
assign n_21339 = ~x_145 &  n_21337;
assign n_21340 = ~n_21338 & ~n_21339;
assign n_21341 =  x_144 & ~n_21178;
assign n_21342 =  i_5 &  n_21178;
assign n_21343 = ~n_21341 & ~n_21342;
assign n_21344 =  x_144 & ~n_21343;
assign n_21345 = ~x_144 &  n_21343;
assign n_21346 = ~n_21344 & ~n_21345;
assign n_21347 =  x_143 & ~n_21178;
assign n_21348 =  i_4 &  n_21178;
assign n_21349 = ~n_21347 & ~n_21348;
assign n_21350 =  x_143 & ~n_21349;
assign n_21351 = ~x_143 &  n_21349;
assign n_21352 = ~n_21350 & ~n_21351;
assign n_21353 =  x_142 & ~n_21178;
assign n_21354 =  i_3 &  n_21178;
assign n_21355 = ~n_21353 & ~n_21354;
assign n_21356 =  x_142 & ~n_21355;
assign n_21357 = ~x_142 &  n_21355;
assign n_21358 = ~n_21356 & ~n_21357;
assign n_21359 =  x_141 & ~n_21178;
assign n_21360 =  i_2 &  n_21178;
assign n_21361 = ~n_21359 & ~n_21360;
assign n_21362 =  x_141 & ~n_21361;
assign n_21363 = ~x_141 &  n_21361;
assign n_21364 = ~n_21362 & ~n_21363;
assign n_21365 =  x_140 & ~n_21178;
assign n_21366 =  i_1 &  n_21178;
assign n_21367 = ~n_21365 & ~n_21366;
assign n_21368 =  x_140 & ~n_21367;
assign n_21369 = ~x_140 &  n_21367;
assign n_21370 = ~n_21368 & ~n_21369;
assign n_21371 =  n_6378 &  n_3615;
assign n_21372 =  x_139 & ~n_21371;
assign n_21373 =  i_32 &  n_21371;
assign n_21374 = ~n_21372 & ~n_21373;
assign n_21375 =  x_139 & ~n_21374;
assign n_21376 = ~x_139 &  n_21374;
assign n_21377 = ~n_21375 & ~n_21376;
assign n_21378 =  x_138 & ~n_21371;
assign n_21379 =  i_31 &  n_21371;
assign n_21380 = ~n_21378 & ~n_21379;
assign n_21381 =  x_138 & ~n_21380;
assign n_21382 = ~x_138 &  n_21380;
assign n_21383 = ~n_21381 & ~n_21382;
assign n_21384 =  x_137 & ~n_21371;
assign n_21385 =  i_30 &  n_21371;
assign n_21386 = ~n_21384 & ~n_21385;
assign n_21387 =  x_137 & ~n_21386;
assign n_21388 = ~x_137 &  n_21386;
assign n_21389 = ~n_21387 & ~n_21388;
assign n_21390 =  x_136 & ~n_21371;
assign n_21391 =  i_29 &  n_21371;
assign n_21392 = ~n_21390 & ~n_21391;
assign n_21393 =  x_136 & ~n_21392;
assign n_21394 = ~x_136 &  n_21392;
assign n_21395 = ~n_21393 & ~n_21394;
assign n_21396 =  x_135 & ~n_21371;
assign n_21397 =  i_28 &  n_21371;
assign n_21398 = ~n_21396 & ~n_21397;
assign n_21399 =  x_135 & ~n_21398;
assign n_21400 = ~x_135 &  n_21398;
assign n_21401 = ~n_21399 & ~n_21400;
assign n_21402 =  x_134 & ~n_21371;
assign n_21403 =  i_27 &  n_21371;
assign n_21404 = ~n_21402 & ~n_21403;
assign n_21405 =  x_134 & ~n_21404;
assign n_21406 = ~x_134 &  n_21404;
assign n_21407 = ~n_21405 & ~n_21406;
assign n_21408 =  x_133 & ~n_21371;
assign n_21409 =  i_26 &  n_21371;
assign n_21410 = ~n_21408 & ~n_21409;
assign n_21411 =  x_133 & ~n_21410;
assign n_21412 = ~x_133 &  n_21410;
assign n_21413 = ~n_21411 & ~n_21412;
assign n_21414 =  x_132 & ~n_21371;
assign n_21415 =  i_25 &  n_21371;
assign n_21416 = ~n_21414 & ~n_21415;
assign n_21417 =  x_132 & ~n_21416;
assign n_21418 = ~x_132 &  n_21416;
assign n_21419 = ~n_21417 & ~n_21418;
assign n_21420 =  x_131 & ~n_21371;
assign n_21421 =  i_24 &  n_21371;
assign n_21422 = ~n_21420 & ~n_21421;
assign n_21423 =  x_131 & ~n_21422;
assign n_21424 = ~x_131 &  n_21422;
assign n_21425 = ~n_21423 & ~n_21424;
assign n_21426 =  x_130 & ~n_21371;
assign n_21427 =  i_23 &  n_21371;
assign n_21428 = ~n_21426 & ~n_21427;
assign n_21429 =  x_130 & ~n_21428;
assign n_21430 = ~x_130 &  n_21428;
assign n_21431 = ~n_21429 & ~n_21430;
assign n_21432 =  x_129 & ~n_21371;
assign n_21433 =  i_22 &  n_21371;
assign n_21434 = ~n_21432 & ~n_21433;
assign n_21435 =  x_129 & ~n_21434;
assign n_21436 = ~x_129 &  n_21434;
assign n_21437 = ~n_21435 & ~n_21436;
assign n_21438 =  x_128 & ~n_21371;
assign n_21439 =  i_21 &  n_21371;
assign n_21440 = ~n_21438 & ~n_21439;
assign n_21441 =  x_128 & ~n_21440;
assign n_21442 = ~x_128 &  n_21440;
assign n_21443 = ~n_21441 & ~n_21442;
assign n_21444 =  x_127 & ~n_21371;
assign n_21445 =  i_20 &  n_21371;
assign n_21446 = ~n_21444 & ~n_21445;
assign n_21447 =  x_127 & ~n_21446;
assign n_21448 = ~x_127 &  n_21446;
assign n_21449 = ~n_21447 & ~n_21448;
assign n_21450 =  x_126 & ~n_21371;
assign n_21451 =  i_19 &  n_21371;
assign n_21452 = ~n_21450 & ~n_21451;
assign n_21453 =  x_126 & ~n_21452;
assign n_21454 = ~x_126 &  n_21452;
assign n_21455 = ~n_21453 & ~n_21454;
assign n_21456 =  x_125 & ~n_21371;
assign n_21457 =  i_18 &  n_21371;
assign n_21458 = ~n_21456 & ~n_21457;
assign n_21459 =  x_125 & ~n_21458;
assign n_21460 = ~x_125 &  n_21458;
assign n_21461 = ~n_21459 & ~n_21460;
assign n_21462 =  x_124 & ~n_21371;
assign n_21463 =  i_17 &  n_21371;
assign n_21464 = ~n_21462 & ~n_21463;
assign n_21465 =  x_124 & ~n_21464;
assign n_21466 = ~x_124 &  n_21464;
assign n_21467 = ~n_21465 & ~n_21466;
assign n_21468 =  x_123 & ~n_21371;
assign n_21469 =  i_16 &  n_21371;
assign n_21470 = ~n_21468 & ~n_21469;
assign n_21471 =  x_123 & ~n_21470;
assign n_21472 = ~x_123 &  n_21470;
assign n_21473 = ~n_21471 & ~n_21472;
assign n_21474 =  x_122 & ~n_21371;
assign n_21475 =  i_15 &  n_21371;
assign n_21476 = ~n_21474 & ~n_21475;
assign n_21477 =  x_122 & ~n_21476;
assign n_21478 = ~x_122 &  n_21476;
assign n_21479 = ~n_21477 & ~n_21478;
assign n_21480 =  x_121 & ~n_21371;
assign n_21481 =  i_14 &  n_21371;
assign n_21482 = ~n_21480 & ~n_21481;
assign n_21483 =  x_121 & ~n_21482;
assign n_21484 = ~x_121 &  n_21482;
assign n_21485 = ~n_21483 & ~n_21484;
assign n_21486 =  x_120 & ~n_21371;
assign n_21487 =  i_13 &  n_21371;
assign n_21488 = ~n_21486 & ~n_21487;
assign n_21489 =  x_120 & ~n_21488;
assign n_21490 = ~x_120 &  n_21488;
assign n_21491 = ~n_21489 & ~n_21490;
assign n_21492 =  x_119 & ~n_21371;
assign n_21493 =  i_12 &  n_21371;
assign n_21494 = ~n_21492 & ~n_21493;
assign n_21495 =  x_119 & ~n_21494;
assign n_21496 = ~x_119 &  n_21494;
assign n_21497 = ~n_21495 & ~n_21496;
assign n_21498 =  x_118 & ~n_21371;
assign n_21499 =  i_11 &  n_21371;
assign n_21500 = ~n_21498 & ~n_21499;
assign n_21501 =  x_118 & ~n_21500;
assign n_21502 = ~x_118 &  n_21500;
assign n_21503 = ~n_21501 & ~n_21502;
assign n_21504 =  x_117 & ~n_21371;
assign n_21505 =  i_10 &  n_21371;
assign n_21506 = ~n_21504 & ~n_21505;
assign n_21507 =  x_117 & ~n_21506;
assign n_21508 = ~x_117 &  n_21506;
assign n_21509 = ~n_21507 & ~n_21508;
assign n_21510 =  x_116 & ~n_21371;
assign n_21511 =  i_9 &  n_21371;
assign n_21512 = ~n_21510 & ~n_21511;
assign n_21513 =  x_116 & ~n_21512;
assign n_21514 = ~x_116 &  n_21512;
assign n_21515 = ~n_21513 & ~n_21514;
assign n_21516 =  x_115 & ~n_21371;
assign n_21517 =  i_8 &  n_21371;
assign n_21518 = ~n_21516 & ~n_21517;
assign n_21519 =  x_115 & ~n_21518;
assign n_21520 = ~x_115 &  n_21518;
assign n_21521 = ~n_21519 & ~n_21520;
assign n_21522 =  x_114 & ~n_21371;
assign n_21523 =  i_7 &  n_21371;
assign n_21524 = ~n_21522 & ~n_21523;
assign n_21525 =  x_114 & ~n_21524;
assign n_21526 = ~x_114 &  n_21524;
assign n_21527 = ~n_21525 & ~n_21526;
assign n_21528 =  x_113 & ~n_21371;
assign n_21529 =  i_6 &  n_21371;
assign n_21530 = ~n_21528 & ~n_21529;
assign n_21531 =  x_113 & ~n_21530;
assign n_21532 = ~x_113 &  n_21530;
assign n_21533 = ~n_21531 & ~n_21532;
assign n_21534 =  x_112 & ~n_21371;
assign n_21535 =  i_5 &  n_21371;
assign n_21536 = ~n_21534 & ~n_21535;
assign n_21537 =  x_112 & ~n_21536;
assign n_21538 = ~x_112 &  n_21536;
assign n_21539 = ~n_21537 & ~n_21538;
assign n_21540 =  x_111 & ~n_21371;
assign n_21541 =  i_4 &  n_21371;
assign n_21542 = ~n_21540 & ~n_21541;
assign n_21543 =  x_111 & ~n_21542;
assign n_21544 = ~x_111 &  n_21542;
assign n_21545 = ~n_21543 & ~n_21544;
assign n_21546 =  x_110 & ~n_21371;
assign n_21547 =  i_3 &  n_21371;
assign n_21548 = ~n_21546 & ~n_21547;
assign n_21549 =  x_110 & ~n_21548;
assign n_21550 = ~x_110 &  n_21548;
assign n_21551 = ~n_21549 & ~n_21550;
assign n_21552 =  x_109 & ~n_21371;
assign n_21553 =  i_2 &  n_21371;
assign n_21554 = ~n_21552 & ~n_21553;
assign n_21555 =  x_109 & ~n_21554;
assign n_21556 = ~x_109 &  n_21554;
assign n_21557 = ~n_21555 & ~n_21556;
assign n_21558 =  x_108 & ~n_21371;
assign n_21559 =  i_1 &  n_21371;
assign n_21560 = ~n_21558 & ~n_21559;
assign n_21561 =  x_108 & ~n_21560;
assign n_21562 = ~x_108 &  n_21560;
assign n_21563 = ~n_21561 & ~n_21562;
assign n_21564 =  n_1174 &  n_153;
assign n_21565 =  n_21564 &  n_7079;
assign n_21566 =  x_107 & ~n_21565;
assign n_21567 =  i_32 &  n_21565;
assign n_21568 = ~n_21566 & ~n_21567;
assign n_21569 =  x_107 & ~n_21568;
assign n_21570 = ~x_107 &  n_21568;
assign n_21571 = ~n_21569 & ~n_21570;
assign n_21572 =  x_106 & ~n_21565;
assign n_21573 =  i_31 &  n_21565;
assign n_21574 = ~n_21572 & ~n_21573;
assign n_21575 =  x_106 & ~n_21574;
assign n_21576 = ~x_106 &  n_21574;
assign n_21577 = ~n_21575 & ~n_21576;
assign n_21578 =  x_105 & ~n_21565;
assign n_21579 =  i_30 &  n_21565;
assign n_21580 = ~n_21578 & ~n_21579;
assign n_21581 =  x_105 & ~n_21580;
assign n_21582 = ~x_105 &  n_21580;
assign n_21583 = ~n_21581 & ~n_21582;
assign n_21584 =  x_104 & ~n_21565;
assign n_21585 =  i_29 &  n_21565;
assign n_21586 = ~n_21584 & ~n_21585;
assign n_21587 =  x_104 & ~n_21586;
assign n_21588 = ~x_104 &  n_21586;
assign n_21589 = ~n_21587 & ~n_21588;
assign n_21590 =  x_103 & ~n_21565;
assign n_21591 =  i_28 &  n_21565;
assign n_21592 = ~n_21590 & ~n_21591;
assign n_21593 =  x_103 & ~n_21592;
assign n_21594 = ~x_103 &  n_21592;
assign n_21595 = ~n_21593 & ~n_21594;
assign n_21596 =  x_102 & ~n_21565;
assign n_21597 =  i_27 &  n_21565;
assign n_21598 = ~n_21596 & ~n_21597;
assign n_21599 =  x_102 & ~n_21598;
assign n_21600 = ~x_102 &  n_21598;
assign n_21601 = ~n_21599 & ~n_21600;
assign n_21602 =  x_101 & ~n_21565;
assign n_21603 =  i_26 &  n_21565;
assign n_21604 = ~n_21602 & ~n_21603;
assign n_21605 =  x_101 & ~n_21604;
assign n_21606 = ~x_101 &  n_21604;
assign n_21607 = ~n_21605 & ~n_21606;
assign n_21608 =  x_100 & ~n_21565;
assign n_21609 =  i_25 &  n_21565;
assign n_21610 = ~n_21608 & ~n_21609;
assign n_21611 =  x_100 & ~n_21610;
assign n_21612 = ~x_100 &  n_21610;
assign n_21613 = ~n_21611 & ~n_21612;
assign n_21614 =  x_99 & ~n_21565;
assign n_21615 =  i_24 &  n_21565;
assign n_21616 = ~n_21614 & ~n_21615;
assign n_21617 =  x_99 & ~n_21616;
assign n_21618 = ~x_99 &  n_21616;
assign n_21619 = ~n_21617 & ~n_21618;
assign n_21620 =  x_98 & ~n_21565;
assign n_21621 =  i_23 &  n_21565;
assign n_21622 = ~n_21620 & ~n_21621;
assign n_21623 =  x_98 & ~n_21622;
assign n_21624 = ~x_98 &  n_21622;
assign n_21625 = ~n_21623 & ~n_21624;
assign n_21626 =  x_97 & ~n_21565;
assign n_21627 =  i_22 &  n_21565;
assign n_21628 = ~n_21626 & ~n_21627;
assign n_21629 =  x_97 & ~n_21628;
assign n_21630 = ~x_97 &  n_21628;
assign n_21631 = ~n_21629 & ~n_21630;
assign n_21632 =  x_96 & ~n_21565;
assign n_21633 =  i_21 &  n_21565;
assign n_21634 = ~n_21632 & ~n_21633;
assign n_21635 =  x_96 & ~n_21634;
assign n_21636 = ~x_96 &  n_21634;
assign n_21637 = ~n_21635 & ~n_21636;
assign n_21638 =  x_95 & ~n_21565;
assign n_21639 =  i_20 &  n_21565;
assign n_21640 = ~n_21638 & ~n_21639;
assign n_21641 =  x_95 & ~n_21640;
assign n_21642 = ~x_95 &  n_21640;
assign n_21643 = ~n_21641 & ~n_21642;
assign n_21644 =  x_94 & ~n_21565;
assign n_21645 =  i_19 &  n_21565;
assign n_21646 = ~n_21644 & ~n_21645;
assign n_21647 =  x_94 & ~n_21646;
assign n_21648 = ~x_94 &  n_21646;
assign n_21649 = ~n_21647 & ~n_21648;
assign n_21650 =  x_93 & ~n_21565;
assign n_21651 =  i_18 &  n_21565;
assign n_21652 = ~n_21650 & ~n_21651;
assign n_21653 =  x_93 & ~n_21652;
assign n_21654 = ~x_93 &  n_21652;
assign n_21655 = ~n_21653 & ~n_21654;
assign n_21656 =  x_92 & ~n_21565;
assign n_21657 =  i_17 &  n_21565;
assign n_21658 = ~n_21656 & ~n_21657;
assign n_21659 =  x_92 & ~n_21658;
assign n_21660 = ~x_92 &  n_21658;
assign n_21661 = ~n_21659 & ~n_21660;
assign n_21662 =  x_91 & ~n_21565;
assign n_21663 =  i_16 &  n_21565;
assign n_21664 = ~n_21662 & ~n_21663;
assign n_21665 =  x_91 & ~n_21664;
assign n_21666 = ~x_91 &  n_21664;
assign n_21667 = ~n_21665 & ~n_21666;
assign n_21668 =  x_90 & ~n_21565;
assign n_21669 =  i_15 &  n_21565;
assign n_21670 = ~n_21668 & ~n_21669;
assign n_21671 =  x_90 & ~n_21670;
assign n_21672 = ~x_90 &  n_21670;
assign n_21673 = ~n_21671 & ~n_21672;
assign n_21674 =  x_89 & ~n_21565;
assign n_21675 =  i_14 &  n_21565;
assign n_21676 = ~n_21674 & ~n_21675;
assign n_21677 =  x_89 & ~n_21676;
assign n_21678 = ~x_89 &  n_21676;
assign n_21679 = ~n_21677 & ~n_21678;
assign n_21680 =  x_88 & ~n_21565;
assign n_21681 =  i_13 &  n_21565;
assign n_21682 = ~n_21680 & ~n_21681;
assign n_21683 =  x_88 & ~n_21682;
assign n_21684 = ~x_88 &  n_21682;
assign n_21685 = ~n_21683 & ~n_21684;
assign n_21686 =  x_87 & ~n_21565;
assign n_21687 =  i_12 &  n_21565;
assign n_21688 = ~n_21686 & ~n_21687;
assign n_21689 =  x_87 & ~n_21688;
assign n_21690 = ~x_87 &  n_21688;
assign n_21691 = ~n_21689 & ~n_21690;
assign n_21692 =  x_86 & ~n_21565;
assign n_21693 =  i_11 &  n_21565;
assign n_21694 = ~n_21692 & ~n_21693;
assign n_21695 =  x_86 & ~n_21694;
assign n_21696 = ~x_86 &  n_21694;
assign n_21697 = ~n_21695 & ~n_21696;
assign n_21698 =  x_85 & ~n_21565;
assign n_21699 =  i_10 &  n_21565;
assign n_21700 = ~n_21698 & ~n_21699;
assign n_21701 =  x_85 & ~n_21700;
assign n_21702 = ~x_85 &  n_21700;
assign n_21703 = ~n_21701 & ~n_21702;
assign n_21704 =  x_84 & ~n_21565;
assign n_21705 =  i_9 &  n_21565;
assign n_21706 = ~n_21704 & ~n_21705;
assign n_21707 =  x_84 & ~n_21706;
assign n_21708 = ~x_84 &  n_21706;
assign n_21709 = ~n_21707 & ~n_21708;
assign n_21710 =  x_83 & ~n_21565;
assign n_21711 =  i_8 &  n_21565;
assign n_21712 = ~n_21710 & ~n_21711;
assign n_21713 =  x_83 & ~n_21712;
assign n_21714 = ~x_83 &  n_21712;
assign n_21715 = ~n_21713 & ~n_21714;
assign n_21716 =  x_82 & ~n_21565;
assign n_21717 =  i_7 &  n_21565;
assign n_21718 = ~n_21716 & ~n_21717;
assign n_21719 =  x_82 & ~n_21718;
assign n_21720 = ~x_82 &  n_21718;
assign n_21721 = ~n_21719 & ~n_21720;
assign n_21722 =  x_81 & ~n_21565;
assign n_21723 =  i_6 &  n_21565;
assign n_21724 = ~n_21722 & ~n_21723;
assign n_21725 =  x_81 & ~n_21724;
assign n_21726 = ~x_81 &  n_21724;
assign n_21727 = ~n_21725 & ~n_21726;
assign n_21728 =  x_80 & ~n_21565;
assign n_21729 =  i_5 &  n_21565;
assign n_21730 = ~n_21728 & ~n_21729;
assign n_21731 =  x_80 & ~n_21730;
assign n_21732 = ~x_80 &  n_21730;
assign n_21733 = ~n_21731 & ~n_21732;
assign n_21734 =  x_79 & ~n_21565;
assign n_21735 =  i_4 &  n_21565;
assign n_21736 = ~n_21734 & ~n_21735;
assign n_21737 =  x_79 & ~n_21736;
assign n_21738 = ~x_79 &  n_21736;
assign n_21739 = ~n_21737 & ~n_21738;
assign n_21740 =  x_78 & ~n_21565;
assign n_21741 =  i_3 &  n_21565;
assign n_21742 = ~n_21740 & ~n_21741;
assign n_21743 =  x_78 & ~n_21742;
assign n_21744 = ~x_78 &  n_21742;
assign n_21745 = ~n_21743 & ~n_21744;
assign n_21746 =  x_77 & ~n_21565;
assign n_21747 =  i_2 &  n_21565;
assign n_21748 = ~n_21746 & ~n_21747;
assign n_21749 =  x_77 & ~n_21748;
assign n_21750 = ~x_77 &  n_21748;
assign n_21751 = ~n_21749 & ~n_21750;
assign n_21752 =  x_76 & ~n_21565;
assign n_21753 =  i_1 &  n_21565;
assign n_21754 = ~n_21752 & ~n_21753;
assign n_21755 =  x_76 & ~n_21754;
assign n_21756 = ~x_76 &  n_21754;
assign n_21757 = ~n_21755 & ~n_21756;
assign n_21758 = ~x_38 &  n_1175;
assign n_21759 =  n_14 &  n_21758;
assign n_21760 =  x_75 & ~n_21759;
assign n_21761 =  i_32 &  n_21759;
assign n_21762 = ~n_21760 & ~n_21761;
assign n_21763 =  x_75 & ~n_21762;
assign n_21764 = ~x_75 &  n_21762;
assign n_21765 = ~n_21763 & ~n_21764;
assign n_21766 =  x_74 & ~n_21759;
assign n_21767 =  i_31 &  n_21759;
assign n_21768 = ~n_21766 & ~n_21767;
assign n_21769 =  x_74 & ~n_21768;
assign n_21770 = ~x_74 &  n_21768;
assign n_21771 = ~n_21769 & ~n_21770;
assign n_21772 =  x_73 & ~n_21759;
assign n_21773 =  i_30 &  n_21759;
assign n_21774 = ~n_21772 & ~n_21773;
assign n_21775 =  x_73 & ~n_21774;
assign n_21776 = ~x_73 &  n_21774;
assign n_21777 = ~n_21775 & ~n_21776;
assign n_21778 =  x_72 & ~n_21759;
assign n_21779 =  i_29 &  n_21759;
assign n_21780 = ~n_21778 & ~n_21779;
assign n_21781 =  x_72 & ~n_21780;
assign n_21782 = ~x_72 &  n_21780;
assign n_21783 = ~n_21781 & ~n_21782;
assign n_21784 =  x_71 & ~n_21759;
assign n_21785 =  i_28 &  n_21759;
assign n_21786 = ~n_21784 & ~n_21785;
assign n_21787 =  x_71 & ~n_21786;
assign n_21788 = ~x_71 &  n_21786;
assign n_21789 = ~n_21787 & ~n_21788;
assign n_21790 =  x_70 & ~n_21759;
assign n_21791 =  i_27 &  n_21759;
assign n_21792 = ~n_21790 & ~n_21791;
assign n_21793 =  x_70 & ~n_21792;
assign n_21794 = ~x_70 &  n_21792;
assign n_21795 = ~n_21793 & ~n_21794;
assign n_21796 =  x_69 & ~n_21759;
assign n_21797 =  i_26 &  n_21759;
assign n_21798 = ~n_21796 & ~n_21797;
assign n_21799 =  x_69 & ~n_21798;
assign n_21800 = ~x_69 &  n_21798;
assign n_21801 = ~n_21799 & ~n_21800;
assign n_21802 =  x_68 & ~n_21759;
assign n_21803 =  i_25 &  n_21759;
assign n_21804 = ~n_21802 & ~n_21803;
assign n_21805 =  x_68 & ~n_21804;
assign n_21806 = ~x_68 &  n_21804;
assign n_21807 = ~n_21805 & ~n_21806;
assign n_21808 =  x_67 & ~n_21759;
assign n_21809 =  i_24 &  n_21759;
assign n_21810 = ~n_21808 & ~n_21809;
assign n_21811 =  x_67 & ~n_21810;
assign n_21812 = ~x_67 &  n_21810;
assign n_21813 = ~n_21811 & ~n_21812;
assign n_21814 =  x_66 & ~n_21759;
assign n_21815 =  i_23 &  n_21759;
assign n_21816 = ~n_21814 & ~n_21815;
assign n_21817 =  x_66 & ~n_21816;
assign n_21818 = ~x_66 &  n_21816;
assign n_21819 = ~n_21817 & ~n_21818;
assign n_21820 =  x_65 & ~n_21759;
assign n_21821 =  i_22 &  n_21759;
assign n_21822 = ~n_21820 & ~n_21821;
assign n_21823 =  x_65 & ~n_21822;
assign n_21824 = ~x_65 &  n_21822;
assign n_21825 = ~n_21823 & ~n_21824;
assign n_21826 =  x_64 & ~n_21759;
assign n_21827 =  i_21 &  n_21759;
assign n_21828 = ~n_21826 & ~n_21827;
assign n_21829 =  x_64 & ~n_21828;
assign n_21830 = ~x_64 &  n_21828;
assign n_21831 = ~n_21829 & ~n_21830;
assign n_21832 =  x_63 & ~n_21759;
assign n_21833 =  i_20 &  n_21759;
assign n_21834 = ~n_21832 & ~n_21833;
assign n_21835 =  x_63 & ~n_21834;
assign n_21836 = ~x_63 &  n_21834;
assign n_21837 = ~n_21835 & ~n_21836;
assign n_21838 =  x_62 & ~n_21759;
assign n_21839 =  i_19 &  n_21759;
assign n_21840 = ~n_21838 & ~n_21839;
assign n_21841 =  x_62 & ~n_21840;
assign n_21842 = ~x_62 &  n_21840;
assign n_21843 = ~n_21841 & ~n_21842;
assign n_21844 =  x_61 & ~n_21759;
assign n_21845 =  i_18 &  n_21759;
assign n_21846 = ~n_21844 & ~n_21845;
assign n_21847 =  x_61 & ~n_21846;
assign n_21848 = ~x_61 &  n_21846;
assign n_21849 = ~n_21847 & ~n_21848;
assign n_21850 =  x_60 & ~n_21759;
assign n_21851 =  i_17 &  n_21759;
assign n_21852 = ~n_21850 & ~n_21851;
assign n_21853 =  x_60 & ~n_21852;
assign n_21854 = ~x_60 &  n_21852;
assign n_21855 = ~n_21853 & ~n_21854;
assign n_21856 =  x_59 & ~n_21759;
assign n_21857 =  i_16 &  n_21759;
assign n_21858 = ~n_21856 & ~n_21857;
assign n_21859 =  x_59 & ~n_21858;
assign n_21860 = ~x_59 &  n_21858;
assign n_21861 = ~n_21859 & ~n_21860;
assign n_21862 =  x_58 & ~n_21759;
assign n_21863 =  i_15 &  n_21759;
assign n_21864 = ~n_21862 & ~n_21863;
assign n_21865 =  x_58 & ~n_21864;
assign n_21866 = ~x_58 &  n_21864;
assign n_21867 = ~n_21865 & ~n_21866;
assign n_21868 =  x_57 & ~n_21759;
assign n_21869 =  i_14 &  n_21759;
assign n_21870 = ~n_21868 & ~n_21869;
assign n_21871 =  x_57 & ~n_21870;
assign n_21872 = ~x_57 &  n_21870;
assign n_21873 = ~n_21871 & ~n_21872;
assign n_21874 =  x_56 & ~n_21759;
assign n_21875 =  i_13 &  n_21759;
assign n_21876 = ~n_21874 & ~n_21875;
assign n_21877 =  x_56 & ~n_21876;
assign n_21878 = ~x_56 &  n_21876;
assign n_21879 = ~n_21877 & ~n_21878;
assign n_21880 =  x_55 & ~n_21759;
assign n_21881 =  i_12 &  n_21759;
assign n_21882 = ~n_21880 & ~n_21881;
assign n_21883 =  x_55 & ~n_21882;
assign n_21884 = ~x_55 &  n_21882;
assign n_21885 = ~n_21883 & ~n_21884;
assign n_21886 =  x_54 & ~n_21759;
assign n_21887 =  i_11 &  n_21759;
assign n_21888 = ~n_21886 & ~n_21887;
assign n_21889 =  x_54 & ~n_21888;
assign n_21890 = ~x_54 &  n_21888;
assign n_21891 = ~n_21889 & ~n_21890;
assign n_21892 =  x_53 & ~n_21759;
assign n_21893 =  i_10 &  n_21759;
assign n_21894 = ~n_21892 & ~n_21893;
assign n_21895 =  x_53 & ~n_21894;
assign n_21896 = ~x_53 &  n_21894;
assign n_21897 = ~n_21895 & ~n_21896;
assign n_21898 =  x_52 & ~n_21759;
assign n_21899 =  i_9 &  n_21759;
assign n_21900 = ~n_21898 & ~n_21899;
assign n_21901 =  x_52 & ~n_21900;
assign n_21902 = ~x_52 &  n_21900;
assign n_21903 = ~n_21901 & ~n_21902;
assign n_21904 =  x_51 & ~n_21759;
assign n_21905 =  i_8 &  n_21759;
assign n_21906 = ~n_21904 & ~n_21905;
assign n_21907 =  x_51 & ~n_21906;
assign n_21908 = ~x_51 &  n_21906;
assign n_21909 = ~n_21907 & ~n_21908;
assign n_21910 =  x_50 & ~n_21759;
assign n_21911 =  i_7 &  n_21759;
assign n_21912 = ~n_21910 & ~n_21911;
assign n_21913 =  x_50 & ~n_21912;
assign n_21914 = ~x_50 &  n_21912;
assign n_21915 = ~n_21913 & ~n_21914;
assign n_21916 =  x_49 & ~n_21759;
assign n_21917 =  i_6 &  n_21759;
assign n_21918 = ~n_21916 & ~n_21917;
assign n_21919 =  x_49 & ~n_21918;
assign n_21920 = ~x_49 &  n_21918;
assign n_21921 = ~n_21919 & ~n_21920;
assign n_21922 =  x_48 & ~n_21759;
assign n_21923 =  i_5 &  n_21759;
assign n_21924 = ~n_21922 & ~n_21923;
assign n_21925 =  x_48 & ~n_21924;
assign n_21926 = ~x_48 &  n_21924;
assign n_21927 = ~n_21925 & ~n_21926;
assign n_21928 =  x_47 & ~n_21759;
assign n_21929 =  i_4 &  n_21759;
assign n_21930 = ~n_21928 & ~n_21929;
assign n_21931 =  x_47 & ~n_21930;
assign n_21932 = ~x_47 &  n_21930;
assign n_21933 = ~n_21931 & ~n_21932;
assign n_21934 =  x_46 & ~n_21759;
assign n_21935 =  i_3 &  n_21759;
assign n_21936 = ~n_21934 & ~n_21935;
assign n_21937 =  x_46 & ~n_21936;
assign n_21938 = ~x_46 &  n_21936;
assign n_21939 = ~n_21937 & ~n_21938;
assign n_21940 =  x_45 & ~n_21759;
assign n_21941 =  i_2 &  n_21759;
assign n_21942 = ~n_21940 & ~n_21941;
assign n_21943 =  x_45 & ~n_21942;
assign n_21944 = ~x_45 &  n_21942;
assign n_21945 = ~n_21943 & ~n_21944;
assign n_21946 =  x_44 & ~n_21759;
assign n_21947 =  i_1 &  n_21759;
assign n_21948 = ~n_21946 & ~n_21947;
assign n_21949 =  x_44 & ~n_21948;
assign n_21950 = ~x_44 &  n_21948;
assign n_21951 = ~n_21949 & ~n_21950;
assign n_21952 =  x_33 &  n_3;
assign n_21953 =  x_36 &  n_21952;
assign n_21954 =  n_6 &  n_756;
assign n_21955 =  n_21953 &  n_21954;
assign n_21956 =  n_21955 &  n_5645;
assign n_21957 = ~x_364 &  x_1579;
assign n_21958 =  x_364 & ~x_1579;
assign n_21959 =  x_365 & ~x_1580;
assign n_21960 = ~x_365 &  x_1580;
assign n_21961 =  x_366 & ~x_1581;
assign n_21962 = ~x_366 &  x_1581;
assign n_21963 =  x_367 & ~x_1582;
assign n_21964 = ~x_367 &  x_1582;
assign n_21965 =  x_368 & ~x_1583;
assign n_21966 = ~x_368 &  x_1583;
assign n_21967 =  x_369 & ~x_1584;
assign n_21968 = ~x_369 &  x_1584;
assign n_21969 =  x_370 & ~x_1585;
assign n_21970 = ~x_370 &  x_1585;
assign n_21971 =  x_371 & ~x_1586;
assign n_21972 = ~x_371 &  x_1586;
assign n_21973 =  x_372 & ~x_1587;
assign n_21974 = ~x_372 &  x_1587;
assign n_21975 =  x_373 & ~x_1588;
assign n_21976 = ~x_373 &  x_1588;
assign n_21977 =  x_374 & ~x_1589;
assign n_21978 = ~x_374 &  x_1589;
assign n_21979 =  x_375 & ~x_1590;
assign n_21980 = ~x_375 &  x_1590;
assign n_21981 =  x_376 & ~x_1591;
assign n_21982 = ~x_376 &  x_1591;
assign n_21983 =  x_377 & ~x_1592;
assign n_21984 = ~x_377 &  x_1592;
assign n_21985 =  x_378 & ~x_1593;
assign n_21986 = ~x_378 &  x_1593;
assign n_21987 =  x_379 & ~x_1594;
assign n_21988 = ~x_379 &  x_1594;
assign n_21989 =  x_380 & ~x_1595;
assign n_21990 = ~x_380 &  x_1595;
assign n_21991 =  x_381 & ~x_1596;
assign n_21992 = ~x_381 &  x_1596;
assign n_21993 =  x_382 & ~x_1597;
assign n_21994 = ~x_382 &  x_1597;
assign n_21995 =  x_383 & ~x_1598;
assign n_21996 = ~x_383 &  x_1598;
assign n_21997 =  x_384 & ~x_1599;
assign n_21998 = ~x_384 &  x_1599;
assign n_21999 =  x_385 & ~x_1600;
assign n_22000 = ~x_385 &  x_1600;
assign n_22001 =  x_386 & ~x_1601;
assign n_22002 = ~x_386 &  x_1601;
assign n_22003 =  x_387 & ~x_1602;
assign n_22004 = ~x_387 &  x_1602;
assign n_22005 =  x_388 & ~x_1603;
assign n_22006 = ~x_388 &  x_1603;
assign n_22007 =  x_389 & ~x_1604;
assign n_22008 = ~x_389 &  x_1604;
assign n_22009 =  x_390 & ~x_1605;
assign n_22010 = ~x_390 &  x_1605;
assign n_22011 =  x_391 & ~x_1606;
assign n_22012 = ~x_391 &  x_1606;
assign n_22013 =  x_392 & ~x_1607;
assign n_22014 = ~x_392 &  x_1607;
assign n_22015 =  x_394 & ~x_1609;
assign n_22016 = ~x_394 &  x_1609;
assign n_22017 =  x_395 & ~x_1610;
assign n_22018 = ~n_22016 &  n_22017;
assign n_22019 = ~n_22015 & ~n_22018;
assign n_22020 =  x_1608 &  n_22019;
assign n_22021 =  x_393 & ~n_22020;
assign n_22022 = ~x_1608 & ~n_22019;
assign n_22023 = ~n_22021 & ~n_22022;
assign n_22024 = ~n_22014 & ~n_22023;
assign n_22025 = ~n_22013 & ~n_22024;
assign n_22026 = ~n_22012 & ~n_22025;
assign n_22027 = ~n_22011 & ~n_22026;
assign n_22028 = ~n_22010 & ~n_22027;
assign n_22029 = ~n_22009 & ~n_22028;
assign n_22030 = ~n_22008 & ~n_22029;
assign n_22031 = ~n_22007 & ~n_22030;
assign n_22032 = ~n_22006 & ~n_22031;
assign n_22033 = ~n_22005 & ~n_22032;
assign n_22034 = ~n_22004 & ~n_22033;
assign n_22035 = ~n_22003 & ~n_22034;
assign n_22036 = ~n_22002 & ~n_22035;
assign n_22037 = ~n_22001 & ~n_22036;
assign n_22038 = ~n_22000 & ~n_22037;
assign n_22039 = ~n_21999 & ~n_22038;
assign n_22040 = ~n_21998 & ~n_22039;
assign n_22041 = ~n_21997 & ~n_22040;
assign n_22042 = ~n_21996 & ~n_22041;
assign n_22043 = ~n_21995 & ~n_22042;
assign n_22044 = ~n_21994 & ~n_22043;
assign n_22045 = ~n_21993 & ~n_22044;
assign n_22046 = ~n_21992 & ~n_22045;
assign n_22047 = ~n_21991 & ~n_22046;
assign n_22048 = ~n_21990 & ~n_22047;
assign n_22049 = ~n_21989 & ~n_22048;
assign n_22050 = ~n_21988 & ~n_22049;
assign n_22051 = ~n_21987 & ~n_22050;
assign n_22052 = ~n_21986 & ~n_22051;
assign n_22053 = ~n_21985 & ~n_22052;
assign n_22054 = ~n_21984 & ~n_22053;
assign n_22055 = ~n_21983 & ~n_22054;
assign n_22056 = ~n_21982 & ~n_22055;
assign n_22057 = ~n_21981 & ~n_22056;
assign n_22058 = ~n_21980 & ~n_22057;
assign n_22059 = ~n_21979 & ~n_22058;
assign n_22060 = ~n_21978 & ~n_22059;
assign n_22061 = ~n_21977 & ~n_22060;
assign n_22062 = ~n_21976 & ~n_22061;
assign n_22063 = ~n_21975 & ~n_22062;
assign n_22064 = ~n_21974 & ~n_22063;
assign n_22065 = ~n_21973 & ~n_22064;
assign n_22066 = ~n_21972 & ~n_22065;
assign n_22067 = ~n_21971 & ~n_22066;
assign n_22068 = ~n_21970 & ~n_22067;
assign n_22069 = ~n_21969 & ~n_22068;
assign n_22070 = ~n_21968 & ~n_22069;
assign n_22071 = ~n_21967 & ~n_22070;
assign n_22072 = ~n_21966 & ~n_22071;
assign n_22073 = ~n_21965 & ~n_22072;
assign n_22074 = ~n_21964 & ~n_22073;
assign n_22075 = ~n_21963 & ~n_22074;
assign n_22076 = ~n_21962 & ~n_22075;
assign n_22077 = ~n_21961 & ~n_22076;
assign n_22078 = ~n_21960 & ~n_22077;
assign n_22079 = ~n_21959 & ~n_22078;
assign n_22080 = ~n_21958 & ~n_22079;
assign n_22081 = ~n_21957 & ~n_22080;
assign n_22082 =  n_21956 & ~n_22081;
assign n_22083 =  n_21955 &  n_758;
assign n_22084 = ~x_875 &  x_1579;
assign n_22085 =  x_875 & ~x_1579;
assign n_22086 =  x_876 & ~x_1580;
assign n_22087 = ~x_876 &  x_1580;
assign n_22088 =  x_877 & ~x_1581;
assign n_22089 = ~x_877 &  x_1581;
assign n_22090 =  x_878 & ~x_1582;
assign n_22091 = ~x_878 &  x_1582;
assign n_22092 =  x_879 & ~x_1583;
assign n_22093 = ~x_879 &  x_1583;
assign n_22094 =  x_880 & ~x_1584;
assign n_22095 = ~x_880 &  x_1584;
assign n_22096 =  x_881 & ~x_1585;
assign n_22097 = ~x_881 &  x_1585;
assign n_22098 =  x_882 & ~x_1586;
assign n_22099 = ~x_882 &  x_1586;
assign n_22100 =  x_883 & ~x_1587;
assign n_22101 = ~x_883 &  x_1587;
assign n_22102 =  x_884 & ~x_1588;
assign n_22103 = ~x_884 &  x_1588;
assign n_22104 =  x_885 & ~x_1589;
assign n_22105 = ~x_885 &  x_1589;
assign n_22106 =  x_886 & ~x_1590;
assign n_22107 = ~x_886 &  x_1590;
assign n_22108 =  x_887 & ~x_1591;
assign n_22109 = ~x_887 &  x_1591;
assign n_22110 =  x_888 & ~x_1592;
assign n_22111 = ~x_888 &  x_1592;
assign n_22112 =  x_889 & ~x_1593;
assign n_22113 = ~x_889 &  x_1593;
assign n_22114 =  x_890 & ~x_1594;
assign n_22115 = ~x_890 &  x_1594;
assign n_22116 =  x_891 & ~x_1595;
assign n_22117 = ~x_891 &  x_1595;
assign n_22118 =  x_892 & ~x_1596;
assign n_22119 = ~x_892 &  x_1596;
assign n_22120 =  x_893 & ~x_1597;
assign n_22121 = ~x_893 &  x_1597;
assign n_22122 =  x_894 & ~x_1598;
assign n_22123 = ~x_894 &  x_1598;
assign n_22124 =  x_895 & ~x_1599;
assign n_22125 = ~x_895 &  x_1599;
assign n_22126 =  x_896 & ~x_1600;
assign n_22127 = ~x_896 &  x_1600;
assign n_22128 =  x_897 & ~x_1601;
assign n_22129 = ~x_897 &  x_1601;
assign n_22130 =  x_898 & ~x_1602;
assign n_22131 = ~x_898 &  x_1602;
assign n_22132 =  x_899 & ~x_1603;
assign n_22133 = ~x_899 &  x_1603;
assign n_22134 =  x_900 & ~x_1604;
assign n_22135 = ~x_900 &  x_1604;
assign n_22136 =  x_901 & ~x_1605;
assign n_22137 = ~x_901 &  x_1605;
assign n_22138 =  x_902 & ~x_1606;
assign n_22139 = ~x_902 &  x_1606;
assign n_22140 =  x_903 & ~x_1607;
assign n_22141 = ~x_903 &  x_1607;
assign n_22142 =  x_905 & ~x_1609;
assign n_22143 = ~x_905 &  x_1609;
assign n_22144 =  x_906 & ~x_1610;
assign n_22145 = ~n_22143 &  n_22144;
assign n_22146 = ~n_22142 & ~n_22145;
assign n_22147 =  x_1608 &  n_22146;
assign n_22148 =  x_904 & ~n_22147;
assign n_22149 = ~x_1608 & ~n_22146;
assign n_22150 = ~n_22148 & ~n_22149;
assign n_22151 = ~n_22141 & ~n_22150;
assign n_22152 = ~n_22140 & ~n_22151;
assign n_22153 = ~n_22139 & ~n_22152;
assign n_22154 = ~n_22138 & ~n_22153;
assign n_22155 = ~n_22137 & ~n_22154;
assign n_22156 = ~n_22136 & ~n_22155;
assign n_22157 = ~n_22135 & ~n_22156;
assign n_22158 = ~n_22134 & ~n_22157;
assign n_22159 = ~n_22133 & ~n_22158;
assign n_22160 = ~n_22132 & ~n_22159;
assign n_22161 = ~n_22131 & ~n_22160;
assign n_22162 = ~n_22130 & ~n_22161;
assign n_22163 = ~n_22129 & ~n_22162;
assign n_22164 = ~n_22128 & ~n_22163;
assign n_22165 = ~n_22127 & ~n_22164;
assign n_22166 = ~n_22126 & ~n_22165;
assign n_22167 = ~n_22125 & ~n_22166;
assign n_22168 = ~n_22124 & ~n_22167;
assign n_22169 = ~n_22123 & ~n_22168;
assign n_22170 = ~n_22122 & ~n_22169;
assign n_22171 = ~n_22121 & ~n_22170;
assign n_22172 = ~n_22120 & ~n_22171;
assign n_22173 = ~n_22119 & ~n_22172;
assign n_22174 = ~n_22118 & ~n_22173;
assign n_22175 = ~n_22117 & ~n_22174;
assign n_22176 = ~n_22116 & ~n_22175;
assign n_22177 = ~n_22115 & ~n_22176;
assign n_22178 = ~n_22114 & ~n_22177;
assign n_22179 = ~n_22113 & ~n_22178;
assign n_22180 = ~n_22112 & ~n_22179;
assign n_22181 = ~n_22111 & ~n_22180;
assign n_22182 = ~n_22110 & ~n_22181;
assign n_22183 = ~n_22109 & ~n_22182;
assign n_22184 = ~n_22108 & ~n_22183;
assign n_22185 = ~n_22107 & ~n_22184;
assign n_22186 = ~n_22106 & ~n_22185;
assign n_22187 = ~n_22105 & ~n_22186;
assign n_22188 = ~n_22104 & ~n_22187;
assign n_22189 = ~n_22103 & ~n_22188;
assign n_22190 = ~n_22102 & ~n_22189;
assign n_22191 = ~n_22101 & ~n_22190;
assign n_22192 = ~n_22100 & ~n_22191;
assign n_22193 = ~n_22099 & ~n_22192;
assign n_22194 = ~n_22098 & ~n_22193;
assign n_22195 = ~n_22097 & ~n_22194;
assign n_22196 = ~n_22096 & ~n_22195;
assign n_22197 = ~n_22095 & ~n_22196;
assign n_22198 = ~n_22094 & ~n_22197;
assign n_22199 = ~n_22093 & ~n_22198;
assign n_22200 = ~n_22092 & ~n_22199;
assign n_22201 = ~n_22091 & ~n_22200;
assign n_22202 = ~n_22090 & ~n_22201;
assign n_22203 = ~n_22089 & ~n_22202;
assign n_22204 = ~n_22088 & ~n_22203;
assign n_22205 = ~n_22087 & ~n_22204;
assign n_22206 = ~n_22086 & ~n_22205;
assign n_22207 = ~n_22085 & ~n_22206;
assign n_22208 = ~n_22084 & ~n_22207;
assign n_22209 =  n_22083 &  n_22208;
assign n_22210 =  n_1038 &  n_9;
assign n_22211 = ~x_1707 &  x_3913;
assign n_22212 =  x_1707 & ~x_3913;
assign n_22213 =  x_1708 & ~x_3914;
assign n_22214 = ~x_1708 &  x_3914;
assign n_22215 =  x_1709 & ~x_3915;
assign n_22216 = ~x_1709 &  x_3915;
assign n_22217 =  x_1710 & ~x_3916;
assign n_22218 = ~x_1710 &  x_3916;
assign n_22219 =  x_1711 & ~x_3917;
assign n_22220 =  x_1712 & ~x_3918;
assign n_22221 = ~x_1713 &  x_3919;
assign n_22222 =  x_1713 & ~x_3919;
assign n_22223 = ~x_1714 &  x_3920;
assign n_22224 =  x_1714 & ~x_3920;
assign n_22225 = ~x_1715 &  x_3921;
assign n_22226 =  x_1715 & ~x_3921;
assign n_22227 = ~x_1716 &  x_3922;
assign n_22228 =  x_1716 & ~x_3922;
assign n_22229 = ~x_1717 &  x_3923;
assign n_22230 =  x_1717 & ~x_3923;
assign n_22231 = ~x_1718 &  x_3924;
assign n_22232 =  x_1718 & ~x_3924;
assign n_22233 = ~x_1719 &  x_3925;
assign n_22234 =  x_1719 & ~x_3925;
assign n_22235 = ~x_1720 &  x_3926;
assign n_22236 =  x_1720 & ~x_3926;
assign n_22237 = ~x_1721 &  x_3927;
assign n_22238 =  x_1721 & ~x_3927;
assign n_22239 = ~x_1722 &  x_3928;
assign n_22240 =  x_1722 & ~x_3928;
assign n_22241 = ~x_1723 &  x_3929;
assign n_22242 =  x_1723 & ~x_3929;
assign n_22243 = ~x_1724 &  x_3930;
assign n_22244 =  x_1724 & ~x_3930;
assign n_22245 = ~x_1725 &  x_3931;
assign n_22246 =  x_1725 & ~x_3931;
assign n_22247 = ~x_1726 &  x_3932;
assign n_22248 =  x_1726 & ~x_3932;
assign n_22249 = ~x_1727 &  x_3933;
assign n_22250 =  x_1727 & ~x_3933;
assign n_22251 = ~x_1728 &  x_3934;
assign n_22252 =  x_1728 & ~x_3934;
assign n_22253 = ~x_1729 &  x_3935;
assign n_22254 =  x_1729 & ~x_3935;
assign n_22255 = ~x_1730 &  x_3936;
assign n_22256 =  x_1730 & ~x_3936;
assign n_22257 = ~x_1731 &  x_3937;
assign n_22258 =  x_1731 & ~x_3937;
assign n_22259 = ~x_1732 &  x_3938;
assign n_22260 =  x_1732 & ~x_3938;
assign n_22261 = ~x_1733 &  x_3939;
assign n_22262 =  x_1733 & ~x_3939;
assign n_22263 = ~x_1734 &  x_3940;
assign n_22264 =  x_1734 & ~x_3940;
assign n_22265 = ~x_1735 &  x_3941;
assign n_22266 =  x_1735 & ~x_3941;
assign n_22267 = ~x_1737 &  x_3943;
assign n_22268 =  x_1738 & ~x_3944;
assign n_22269 = ~n_22267 &  n_22268;
assign n_22270 =  x_1737 & ~x_3943;
assign n_22271 =  x_1736 & ~x_3942;
assign n_22272 = ~n_22270 & ~n_22271;
assign n_22273 = ~n_22269 &  n_22272;
assign n_22274 = ~x_1736 &  x_3942;
assign n_22275 = ~n_22273 & ~n_22274;
assign n_22276 = ~n_22266 & ~n_22275;
assign n_22277 = ~n_22265 & ~n_22276;
assign n_22278 = ~n_22264 & ~n_22277;
assign n_22279 = ~n_22263 & ~n_22278;
assign n_22280 = ~n_22262 & ~n_22279;
assign n_22281 = ~n_22261 & ~n_22280;
assign n_22282 = ~n_22260 & ~n_22281;
assign n_22283 = ~n_22259 & ~n_22282;
assign n_22284 = ~n_22258 & ~n_22283;
assign n_22285 = ~n_22257 & ~n_22284;
assign n_22286 = ~n_22256 & ~n_22285;
assign n_22287 = ~n_22255 & ~n_22286;
assign n_22288 = ~n_22254 & ~n_22287;
assign n_22289 = ~n_22253 & ~n_22288;
assign n_22290 = ~n_22252 & ~n_22289;
assign n_22291 = ~n_22251 & ~n_22290;
assign n_22292 = ~n_22250 & ~n_22291;
assign n_22293 = ~n_22249 & ~n_22292;
assign n_22294 = ~n_22248 & ~n_22293;
assign n_22295 = ~n_22247 & ~n_22294;
assign n_22296 = ~n_22246 & ~n_22295;
assign n_22297 = ~n_22245 & ~n_22296;
assign n_22298 = ~n_22244 & ~n_22297;
assign n_22299 = ~n_22243 & ~n_22298;
assign n_22300 = ~n_22242 & ~n_22299;
assign n_22301 = ~n_22241 & ~n_22300;
assign n_22302 = ~n_22240 & ~n_22301;
assign n_22303 = ~n_22239 & ~n_22302;
assign n_22304 = ~n_22238 & ~n_22303;
assign n_22305 = ~n_22237 & ~n_22304;
assign n_22306 = ~n_22236 & ~n_22305;
assign n_22307 = ~n_22235 & ~n_22306;
assign n_22308 = ~n_22234 & ~n_22307;
assign n_22309 = ~n_22233 & ~n_22308;
assign n_22310 = ~n_22232 & ~n_22309;
assign n_22311 = ~n_22231 & ~n_22310;
assign n_22312 = ~n_22230 & ~n_22311;
assign n_22313 = ~n_22229 & ~n_22312;
assign n_22314 = ~n_22228 & ~n_22313;
assign n_22315 = ~n_22227 & ~n_22314;
assign n_22316 = ~n_22226 & ~n_22315;
assign n_22317 = ~n_22225 & ~n_22316;
assign n_22318 = ~n_22224 & ~n_22317;
assign n_22319 = ~n_22223 & ~n_22318;
assign n_22320 = ~n_22222 & ~n_22319;
assign n_22321 = ~n_22221 & ~n_22320;
assign n_22322 = ~n_22220 & ~n_22321;
assign n_22323 = ~x_1712 &  x_3918;
assign n_22324 = ~x_1711 &  x_3917;
assign n_22325 = ~n_22323 & ~n_22324;
assign n_22326 = ~n_22322 &  n_22325;
assign n_22327 = ~n_22219 & ~n_22326;
assign n_22328 = ~n_22218 & ~n_22327;
assign n_22329 = ~n_22217 & ~n_22328;
assign n_22330 = ~n_22216 & ~n_22329;
assign n_22331 = ~n_22215 & ~n_22330;
assign n_22332 = ~n_22214 & ~n_22331;
assign n_22333 = ~n_22213 & ~n_22332;
assign n_22334 = ~n_22212 & ~n_22333;
assign n_22335 = ~n_22211 & ~n_22334;
assign n_22336 =  n_22210 & ~n_22335;
assign n_22337 =  n_8344 &  n_3616;
assign n_22338 = ~x_1675 &  x_2315;
assign n_22339 =  x_1675 & ~x_2315;
assign n_22340 =  x_1676 & ~x_2316;
assign n_22341 = ~x_1676 &  x_2316;
assign n_22342 =  x_1677 & ~x_2317;
assign n_22343 = ~x_1677 &  x_2317;
assign n_22344 =  x_1678 & ~x_2318;
assign n_22345 = ~x_1678 &  x_2318;
assign n_22346 =  x_1679 & ~x_2319;
assign n_22347 =  x_1680 & ~x_2320;
assign n_22348 = ~x_1681 &  x_2321;
assign n_22349 =  x_1681 & ~x_2321;
assign n_22350 = ~x_1682 &  x_2322;
assign n_22351 =  x_1682 & ~x_2322;
assign n_22352 = ~x_1683 &  x_2323;
assign n_22353 =  x_1683 & ~x_2323;
assign n_22354 = ~x_1684 &  x_2324;
assign n_22355 =  x_1684 & ~x_2324;
assign n_22356 = ~x_1685 &  x_2325;
assign n_22357 =  x_1685 & ~x_2325;
assign n_22358 = ~x_1686 &  x_2326;
assign n_22359 =  x_1686 & ~x_2326;
assign n_22360 = ~x_1687 &  x_2327;
assign n_22361 =  x_1687 & ~x_2327;
assign n_22362 = ~x_1688 &  x_2328;
assign n_22363 =  x_1688 & ~x_2328;
assign n_22364 = ~x_1689 &  x_2329;
assign n_22365 =  x_1689 & ~x_2329;
assign n_22366 = ~x_1690 &  x_2330;
assign n_22367 =  x_1690 & ~x_2330;
assign n_22368 = ~x_1691 &  x_2331;
assign n_22369 =  x_1691 & ~x_2331;
assign n_22370 = ~x_1692 &  x_2332;
assign n_22371 =  x_1692 & ~x_2332;
assign n_22372 = ~x_1693 &  x_2333;
assign n_22373 =  x_1693 & ~x_2333;
assign n_22374 = ~x_1694 &  x_2334;
assign n_22375 =  x_1694 & ~x_2334;
assign n_22376 = ~x_1695 &  x_2335;
assign n_22377 =  x_1695 & ~x_2335;
assign n_22378 = ~x_1696 &  x_2336;
assign n_22379 =  x_1696 & ~x_2336;
assign n_22380 = ~x_1697 &  x_2337;
assign n_22381 =  x_1697 & ~x_2337;
assign n_22382 = ~x_1698 &  x_2338;
assign n_22383 =  x_1698 & ~x_2338;
assign n_22384 = ~x_1699 &  x_2339;
assign n_22385 =  x_1699 & ~x_2339;
assign n_22386 = ~x_1700 &  x_2340;
assign n_22387 =  x_1700 & ~x_2340;
assign n_22388 = ~x_1701 &  x_2341;
assign n_22389 =  x_1701 & ~x_2341;
assign n_22390 = ~x_1702 &  x_2342;
assign n_22391 =  x_1702 & ~x_2342;
assign n_22392 = ~x_1703 &  x_2343;
assign n_22393 =  x_1703 & ~x_2343;
assign n_22394 = ~x_1705 &  x_2345;
assign n_22395 =  x_1706 & ~x_2346;
assign n_22396 = ~n_22394 &  n_22395;
assign n_22397 =  x_1705 & ~x_2345;
assign n_22398 =  x_1704 & ~x_2344;
assign n_22399 = ~n_22397 & ~n_22398;
assign n_22400 = ~n_22396 &  n_22399;
assign n_22401 = ~x_1704 &  x_2344;
assign n_22402 = ~n_22400 & ~n_22401;
assign n_22403 = ~n_22393 & ~n_22402;
assign n_22404 = ~n_22392 & ~n_22403;
assign n_22405 = ~n_22391 & ~n_22404;
assign n_22406 = ~n_22390 & ~n_22405;
assign n_22407 = ~n_22389 & ~n_22406;
assign n_22408 = ~n_22388 & ~n_22407;
assign n_22409 = ~n_22387 & ~n_22408;
assign n_22410 = ~n_22386 & ~n_22409;
assign n_22411 = ~n_22385 & ~n_22410;
assign n_22412 = ~n_22384 & ~n_22411;
assign n_22413 = ~n_22383 & ~n_22412;
assign n_22414 = ~n_22382 & ~n_22413;
assign n_22415 = ~n_22381 & ~n_22414;
assign n_22416 = ~n_22380 & ~n_22415;
assign n_22417 = ~n_22379 & ~n_22416;
assign n_22418 = ~n_22378 & ~n_22417;
assign n_22419 = ~n_22377 & ~n_22418;
assign n_22420 = ~n_22376 & ~n_22419;
assign n_22421 = ~n_22375 & ~n_22420;
assign n_22422 = ~n_22374 & ~n_22421;
assign n_22423 = ~n_22373 & ~n_22422;
assign n_22424 = ~n_22372 & ~n_22423;
assign n_22425 = ~n_22371 & ~n_22424;
assign n_22426 = ~n_22370 & ~n_22425;
assign n_22427 = ~n_22369 & ~n_22426;
assign n_22428 = ~n_22368 & ~n_22427;
assign n_22429 = ~n_22367 & ~n_22428;
assign n_22430 = ~n_22366 & ~n_22429;
assign n_22431 = ~n_22365 & ~n_22430;
assign n_22432 = ~n_22364 & ~n_22431;
assign n_22433 = ~n_22363 & ~n_22432;
assign n_22434 = ~n_22362 & ~n_22433;
assign n_22435 = ~n_22361 & ~n_22434;
assign n_22436 = ~n_22360 & ~n_22435;
assign n_22437 = ~n_22359 & ~n_22436;
assign n_22438 = ~n_22358 & ~n_22437;
assign n_22439 = ~n_22357 & ~n_22438;
assign n_22440 = ~n_22356 & ~n_22439;
assign n_22441 = ~n_22355 & ~n_22440;
assign n_22442 = ~n_22354 & ~n_22441;
assign n_22443 = ~n_22353 & ~n_22442;
assign n_22444 = ~n_22352 & ~n_22443;
assign n_22445 = ~n_22351 & ~n_22444;
assign n_22446 = ~n_22350 & ~n_22445;
assign n_22447 = ~n_22349 & ~n_22446;
assign n_22448 = ~n_22348 & ~n_22447;
assign n_22449 = ~n_22347 & ~n_22448;
assign n_22450 = ~x_1680 &  x_2320;
assign n_22451 = ~x_1679 &  x_2319;
assign n_22452 = ~n_22450 & ~n_22451;
assign n_22453 = ~n_22449 &  n_22452;
assign n_22454 = ~n_22346 & ~n_22453;
assign n_22455 = ~n_22345 & ~n_22454;
assign n_22456 = ~n_22344 & ~n_22455;
assign n_22457 = ~n_22343 & ~n_22456;
assign n_22458 = ~n_22342 & ~n_22457;
assign n_22459 = ~n_22341 & ~n_22458;
assign n_22460 = ~n_22340 & ~n_22459;
assign n_22461 = ~n_22339 & ~n_22460;
assign n_22462 = ~n_22338 & ~n_22461;
assign n_22463 =  n_22337 & ~n_22462;
assign n_22464 = ~n_22336 & ~n_22463;
assign n_22465 =  n_153 &  n_3346;
assign n_22466 = ~x_2587 &  x_4265;
assign n_22467 =  x_2587 & ~x_4265;
assign n_22468 =  x_2588 & ~x_4266;
assign n_22469 = ~x_2588 &  x_4266;
assign n_22470 =  x_2589 & ~x_4267;
assign n_22471 = ~x_2589 &  x_4267;
assign n_22472 =  x_2590 & ~x_4268;
assign n_22473 = ~x_2590 &  x_4268;
assign n_22474 =  x_2591 & ~x_4269;
assign n_22475 =  x_2592 & ~x_4270;
assign n_22476 = ~x_2593 &  x_4271;
assign n_22477 =  x_2593 & ~x_4271;
assign n_22478 = ~x_2594 &  x_4272;
assign n_22479 =  x_2594 & ~x_4272;
assign n_22480 = ~x_2595 &  x_4273;
assign n_22481 =  x_2595 & ~x_4273;
assign n_22482 = ~x_2596 &  x_4274;
assign n_22483 =  x_2596 & ~x_4274;
assign n_22484 = ~x_2597 &  x_4275;
assign n_22485 =  x_2597 & ~x_4275;
assign n_22486 = ~x_2598 &  x_4276;
assign n_22487 =  x_2598 & ~x_4276;
assign n_22488 = ~x_2599 &  x_4277;
assign n_22489 =  x_2599 & ~x_4277;
assign n_22490 = ~x_2600 &  x_4278;
assign n_22491 =  x_2600 & ~x_4278;
assign n_22492 = ~x_2601 &  x_4279;
assign n_22493 =  x_2601 & ~x_4279;
assign n_22494 = ~x_2602 &  x_4280;
assign n_22495 =  x_2602 & ~x_4280;
assign n_22496 = ~x_2603 &  x_4281;
assign n_22497 =  x_2603 & ~x_4281;
assign n_22498 = ~x_2604 &  x_4282;
assign n_22499 =  x_2604 & ~x_4282;
assign n_22500 = ~x_2605 &  x_4283;
assign n_22501 =  x_2605 & ~x_4283;
assign n_22502 = ~x_2606 &  x_4284;
assign n_22503 =  x_2606 & ~x_4284;
assign n_22504 = ~x_2607 &  x_4285;
assign n_22505 =  x_2607 & ~x_4285;
assign n_22506 = ~x_2608 &  x_4286;
assign n_22507 =  x_2608 & ~x_4286;
assign n_22508 = ~x_2609 &  x_4287;
assign n_22509 =  x_2609 & ~x_4287;
assign n_22510 = ~x_2610 &  x_4288;
assign n_22511 =  x_2610 & ~x_4288;
assign n_22512 = ~x_2611 &  x_4289;
assign n_22513 =  x_2611 & ~x_4289;
assign n_22514 = ~x_2612 &  x_4290;
assign n_22515 =  x_2612 & ~x_4290;
assign n_22516 = ~x_2613 &  x_4291;
assign n_22517 =  x_2613 & ~x_4291;
assign n_22518 = ~x_2614 &  x_4292;
assign n_22519 =  x_2614 & ~x_4292;
assign n_22520 = ~x_2615 &  x_4293;
assign n_22521 =  x_2615 & ~x_4293;
assign n_22522 = ~x_2617 &  x_4295;
assign n_22523 =  x_2618 & ~x_4296;
assign n_22524 = ~n_22522 &  n_22523;
assign n_22525 =  x_2617 & ~x_4295;
assign n_22526 =  x_2616 & ~x_4294;
assign n_22527 = ~n_22525 & ~n_22526;
assign n_22528 = ~n_22524 &  n_22527;
assign n_22529 = ~x_2616 &  x_4294;
assign n_22530 = ~n_22528 & ~n_22529;
assign n_22531 = ~n_22521 & ~n_22530;
assign n_22532 = ~n_22520 & ~n_22531;
assign n_22533 = ~n_22519 & ~n_22532;
assign n_22534 = ~n_22518 & ~n_22533;
assign n_22535 = ~n_22517 & ~n_22534;
assign n_22536 = ~n_22516 & ~n_22535;
assign n_22537 = ~n_22515 & ~n_22536;
assign n_22538 = ~n_22514 & ~n_22537;
assign n_22539 = ~n_22513 & ~n_22538;
assign n_22540 = ~n_22512 & ~n_22539;
assign n_22541 = ~n_22511 & ~n_22540;
assign n_22542 = ~n_22510 & ~n_22541;
assign n_22543 = ~n_22509 & ~n_22542;
assign n_22544 = ~n_22508 & ~n_22543;
assign n_22545 = ~n_22507 & ~n_22544;
assign n_22546 = ~n_22506 & ~n_22545;
assign n_22547 = ~n_22505 & ~n_22546;
assign n_22548 = ~n_22504 & ~n_22547;
assign n_22549 = ~n_22503 & ~n_22548;
assign n_22550 = ~n_22502 & ~n_22549;
assign n_22551 = ~n_22501 & ~n_22550;
assign n_22552 = ~n_22500 & ~n_22551;
assign n_22553 = ~n_22499 & ~n_22552;
assign n_22554 = ~n_22498 & ~n_22553;
assign n_22555 = ~n_22497 & ~n_22554;
assign n_22556 = ~n_22496 & ~n_22555;
assign n_22557 = ~n_22495 & ~n_22556;
assign n_22558 = ~n_22494 & ~n_22557;
assign n_22559 = ~n_22493 & ~n_22558;
assign n_22560 = ~n_22492 & ~n_22559;
assign n_22561 = ~n_22491 & ~n_22560;
assign n_22562 = ~n_22490 & ~n_22561;
assign n_22563 = ~n_22489 & ~n_22562;
assign n_22564 = ~n_22488 & ~n_22563;
assign n_22565 = ~n_22487 & ~n_22564;
assign n_22566 = ~n_22486 & ~n_22565;
assign n_22567 = ~n_22485 & ~n_22566;
assign n_22568 = ~n_22484 & ~n_22567;
assign n_22569 = ~n_22483 & ~n_22568;
assign n_22570 = ~n_22482 & ~n_22569;
assign n_22571 = ~n_22481 & ~n_22570;
assign n_22572 = ~n_22480 & ~n_22571;
assign n_22573 = ~n_22479 & ~n_22572;
assign n_22574 = ~n_22478 & ~n_22573;
assign n_22575 = ~n_22477 & ~n_22574;
assign n_22576 = ~n_22476 & ~n_22575;
assign n_22577 = ~n_22475 & ~n_22576;
assign n_22578 = ~x_2592 &  x_4270;
assign n_22579 = ~x_2591 &  x_4269;
assign n_22580 = ~n_22578 & ~n_22579;
assign n_22581 = ~n_22577 &  n_22580;
assign n_22582 = ~n_22474 & ~n_22581;
assign n_22583 = ~n_22473 & ~n_22582;
assign n_22584 = ~n_22472 & ~n_22583;
assign n_22585 = ~n_22471 & ~n_22584;
assign n_22586 = ~n_22470 & ~n_22585;
assign n_22587 = ~n_22469 & ~n_22586;
assign n_22588 = ~n_22468 & ~n_22587;
assign n_22589 = ~n_22467 & ~n_22588;
assign n_22590 = ~n_22466 & ~n_22589;
assign n_22591 =  n_22465 & ~n_22590;
assign n_22592 =  x_560 & ~x_3356;
assign n_22593 = ~x_561 &  x_3357;
assign n_22594 =  x_561 & ~x_3357;
assign n_22595 = ~x_562 &  x_3358;
assign n_22596 =  x_562 & ~x_3358;
assign n_22597 = ~x_563 &  x_3359;
assign n_22598 =  x_563 & ~x_3359;
assign n_22599 = ~x_564 &  x_3360;
assign n_22600 =  x_564 & ~x_3360;
assign n_22601 = ~x_565 &  x_3361;
assign n_22602 =  x_565 & ~x_3361;
assign n_22603 = ~x_566 &  x_3362;
assign n_22604 =  x_566 & ~x_3362;
assign n_22605 = ~x_567 &  x_3363;
assign n_22606 =  x_567 & ~x_3363;
assign n_22607 = ~x_568 &  x_3364;
assign n_22608 =  x_568 & ~x_3364;
assign n_22609 = ~x_569 &  x_3365;
assign n_22610 =  x_569 & ~x_3365;
assign n_22611 = ~x_570 &  x_3366;
assign n_22612 =  x_570 & ~x_3366;
assign n_22613 = ~x_571 &  x_3367;
assign n_22614 =  x_571 & ~x_3367;
assign n_22615 = ~x_572 &  x_3368;
assign n_22616 =  x_572 & ~x_3368;
assign n_22617 = ~x_573 &  x_3369;
assign n_22618 =  x_573 & ~x_3369;
assign n_22619 = ~x_574 &  x_3370;
assign n_22620 =  x_574 & ~x_3370;
assign n_22621 = ~x_575 &  x_3371;
assign n_22622 =  x_575 & ~x_3371;
assign n_22623 = ~x_576 &  x_3372;
assign n_22624 =  x_576 & ~x_3372;
assign n_22625 = ~x_577 &  x_3373;
assign n_22626 =  x_577 & ~x_3373;
assign n_22627 = ~x_578 &  x_3374;
assign n_22628 =  x_578 & ~x_3374;
assign n_22629 = ~x_579 &  x_3375;
assign n_22630 =  x_579 & ~x_3375;
assign n_22631 = ~x_580 &  x_3376;
assign n_22632 =  x_580 & ~x_3376;
assign n_22633 = ~x_581 &  x_3377;
assign n_22634 =  x_581 & ~x_3377;
assign n_22635 = ~x_582 &  x_3378;
assign n_22636 =  x_582 & ~x_3378;
assign n_22637 = ~x_583 &  x_3379;
assign n_22638 =  x_583 & ~x_3379;
assign n_22639 = ~x_584 &  x_3380;
assign n_22640 =  x_584 & ~x_3380;
assign n_22641 = ~x_586 &  x_3382;
assign n_22642 =  x_586 & ~x_3382;
assign n_22643 = ~x_587 &  x_3383;
assign n_22644 = ~n_22642 &  n_22643;
assign n_22645 = ~n_22641 & ~n_22644;
assign n_22646 =  x_585 &  n_22645;
assign n_22647 =  x_3381 & ~n_22646;
assign n_22648 = ~x_585 & ~n_22645;
assign n_22649 = ~n_22647 & ~n_22648;
assign n_22650 = ~n_22640 & ~n_22649;
assign n_22651 = ~n_22639 & ~n_22650;
assign n_22652 = ~n_22638 & ~n_22651;
assign n_22653 = ~n_22637 & ~n_22652;
assign n_22654 = ~n_22636 & ~n_22653;
assign n_22655 = ~n_22635 & ~n_22654;
assign n_22656 = ~n_22634 & ~n_22655;
assign n_22657 = ~n_22633 & ~n_22656;
assign n_22658 = ~n_22632 & ~n_22657;
assign n_22659 = ~n_22631 & ~n_22658;
assign n_22660 = ~n_22630 & ~n_22659;
assign n_22661 = ~n_22629 & ~n_22660;
assign n_22662 = ~n_22628 & ~n_22661;
assign n_22663 = ~n_22627 & ~n_22662;
assign n_22664 = ~n_22626 & ~n_22663;
assign n_22665 = ~n_22625 & ~n_22664;
assign n_22666 = ~n_22624 & ~n_22665;
assign n_22667 = ~n_22623 & ~n_22666;
assign n_22668 = ~n_22622 & ~n_22667;
assign n_22669 = ~n_22621 & ~n_22668;
assign n_22670 = ~n_22620 & ~n_22669;
assign n_22671 = ~n_22619 & ~n_22670;
assign n_22672 = ~n_22618 & ~n_22671;
assign n_22673 = ~n_22617 & ~n_22672;
assign n_22674 = ~n_22616 & ~n_22673;
assign n_22675 = ~n_22615 & ~n_22674;
assign n_22676 = ~n_22614 & ~n_22675;
assign n_22677 = ~n_22613 & ~n_22676;
assign n_22678 = ~n_22612 & ~n_22677;
assign n_22679 = ~n_22611 & ~n_22678;
assign n_22680 = ~n_22610 & ~n_22679;
assign n_22681 = ~n_22609 & ~n_22680;
assign n_22682 = ~n_22608 & ~n_22681;
assign n_22683 = ~n_22607 & ~n_22682;
assign n_22684 = ~n_22606 & ~n_22683;
assign n_22685 = ~n_22605 & ~n_22684;
assign n_22686 = ~n_22604 & ~n_22685;
assign n_22687 = ~n_22603 & ~n_22686;
assign n_22688 = ~n_22602 & ~n_22687;
assign n_22689 = ~n_22601 & ~n_22688;
assign n_22690 = ~n_22600 & ~n_22689;
assign n_22691 = ~n_22599 & ~n_22690;
assign n_22692 = ~n_22598 & ~n_22691;
assign n_22693 = ~n_22597 & ~n_22692;
assign n_22694 = ~n_22596 & ~n_22693;
assign n_22695 = ~n_22595 & ~n_22694;
assign n_22696 = ~n_22594 & ~n_22695;
assign n_22697 = ~n_22593 & ~n_22696;
assign n_22698 = ~n_22592 & ~n_22697;
assign n_22699 = ~x_560 &  x_3356;
assign n_22700 = ~x_559 &  x_3355;
assign n_22701 = ~n_22699 & ~n_22700;
assign n_22702 = ~n_22698 &  n_22701;
assign n_22703 =  x_558 & ~x_3354;
assign n_22704 =  x_559 & ~x_3355;
assign n_22705 = ~n_22703 & ~n_22704;
assign n_22706 = ~n_22702 &  n_22705;
assign n_22707 = ~x_558 &  x_3354;
assign n_22708 = ~x_557 &  x_3353;
assign n_22709 = ~n_22707 & ~n_22708;
assign n_22710 = ~n_22706 &  n_22709;
assign n_22711 =  x_557 & ~x_3353;
assign n_22712 = ~x_556 &  x_3352;
assign n_22713 = ~n_22711 & ~n_22712;
assign n_22714 = ~n_22710 &  n_22713;
assign n_22715 = ~x_36 &  n_21952;
assign n_22716 =  n_22715 &  n_3142;
assign n_22717 =  n_758 &  n_22716;
assign n_22718 =  x_556 & ~x_3352;
assign n_22719 =  n_22717 & ~n_22718;
assign n_22720 = ~n_22714 &  n_22719;
assign n_22721 =  n_555 &  n_17784;
assign n_22722 =  x_778 &  x_779;
assign n_22723 =  x_777 &  n_22722;
assign n_22724 =  x_776 &  n_22723;
assign n_22725 =  x_775 &  n_22724;
assign n_22726 =  x_774 &  n_22725;
assign n_22727 =  x_773 &  n_22726;
assign n_22728 =  x_772 &  n_22727;
assign n_22729 =  x_771 &  n_22728;
assign n_22730 =  x_770 &  n_22729;
assign n_22731 =  x_769 &  n_22730;
assign n_22732 =  x_768 &  n_22731;
assign n_22733 =  x_767 &  n_22732;
assign n_22734 =  x_766 &  n_22733;
assign n_22735 =  x_765 &  n_22734;
assign n_22736 =  x_764 &  n_22735;
assign n_22737 =  x_763 &  n_22736;
assign n_22738 =  x_762 &  n_22737;
assign n_22739 =  x_761 &  n_22738;
assign n_22740 =  x_760 &  n_22739;
assign n_22741 =  x_759 &  n_22740;
assign n_22742 =  x_758 &  n_22741;
assign n_22743 =  x_757 &  n_22742;
assign n_22744 =  x_756 &  n_22743;
assign n_22745 =  x_755 &  n_22744;
assign n_22746 =  x_754 &  n_22745;
assign n_22747 =  x_753 &  n_22746;
assign n_22748 =  x_752 &  n_22747;
assign n_22749 =  x_751 &  n_22748;
assign n_22750 =  x_750 &  n_22749;
assign n_22751 =  x_749 &  n_22750;
assign n_22752 = ~x_749 & ~n_22750;
assign n_22753 = ~n_22751 & ~n_22752;
assign n_22754 = ~x_653 &  n_22753;
assign n_22755 = ~x_750 & ~n_22749;
assign n_22756 = ~n_22750 & ~n_22755;
assign n_22757 =  x_654 & ~n_22756;
assign n_22758 = ~x_751 & ~n_22748;
assign n_22759 = ~n_22749 & ~n_22758;
assign n_22760 =  x_655 & ~n_22759;
assign n_22761 = ~x_752 & ~n_22747;
assign n_22762 = ~n_22748 & ~n_22761;
assign n_22763 = ~x_656 &  n_22762;
assign n_22764 =  x_656 & ~n_22762;
assign n_22765 = ~x_753 & ~n_22746;
assign n_22766 = ~n_22747 & ~n_22765;
assign n_22767 = ~x_657 &  n_22766;
assign n_22768 =  x_657 & ~n_22766;
assign n_22769 = ~x_754 & ~n_22745;
assign n_22770 = ~n_22746 & ~n_22769;
assign n_22771 = ~x_658 &  n_22770;
assign n_22772 =  x_658 & ~n_22770;
assign n_22773 = ~x_755 & ~n_22744;
assign n_22774 = ~n_22745 & ~n_22773;
assign n_22775 = ~x_659 &  n_22774;
assign n_22776 =  x_659 & ~n_22774;
assign n_22777 = ~x_756 & ~n_22743;
assign n_22778 = ~n_22744 & ~n_22777;
assign n_22779 = ~x_660 &  n_22778;
assign n_22780 =  x_660 & ~n_22778;
assign n_22781 = ~x_757 & ~n_22742;
assign n_22782 = ~n_22743 & ~n_22781;
assign n_22783 = ~x_661 &  n_22782;
assign n_22784 =  x_661 & ~n_22782;
assign n_22785 = ~x_758 & ~n_22741;
assign n_22786 = ~n_22742 & ~n_22785;
assign n_22787 = ~x_662 &  n_22786;
assign n_22788 =  x_662 & ~n_22786;
assign n_22789 = ~x_759 & ~n_22740;
assign n_22790 = ~n_22741 & ~n_22789;
assign n_22791 = ~x_663 &  n_22790;
assign n_22792 =  x_663 & ~n_22790;
assign n_22793 = ~x_760 & ~n_22739;
assign n_22794 = ~n_22740 & ~n_22793;
assign n_22795 = ~x_664 &  n_22794;
assign n_22796 =  x_664 & ~n_22794;
assign n_22797 = ~x_761 & ~n_22738;
assign n_22798 = ~n_22739 & ~n_22797;
assign n_22799 = ~x_665 &  n_22798;
assign n_22800 =  x_665 & ~n_22798;
assign n_22801 = ~x_762 & ~n_22737;
assign n_22802 = ~n_22738 & ~n_22801;
assign n_22803 = ~x_666 &  n_22802;
assign n_22804 =  x_666 & ~n_22802;
assign n_22805 = ~x_763 & ~n_22736;
assign n_22806 = ~n_22737 & ~n_22805;
assign n_22807 = ~x_667 &  n_22806;
assign n_22808 =  x_667 & ~n_22806;
assign n_22809 = ~x_764 & ~n_22735;
assign n_22810 = ~n_22736 & ~n_22809;
assign n_22811 = ~x_668 &  n_22810;
assign n_22812 =  x_668 & ~n_22810;
assign n_22813 = ~x_765 & ~n_22734;
assign n_22814 = ~n_22735 & ~n_22813;
assign n_22815 = ~x_669 &  n_22814;
assign n_22816 =  x_669 & ~n_22814;
assign n_22817 = ~x_766 & ~n_22733;
assign n_22818 = ~n_22734 & ~n_22817;
assign n_22819 = ~x_670 &  n_22818;
assign n_22820 =  x_670 & ~n_22818;
assign n_22821 = ~x_767 & ~n_22732;
assign n_22822 = ~n_22733 & ~n_22821;
assign n_22823 = ~x_671 &  n_22822;
assign n_22824 =  x_671 & ~n_22822;
assign n_22825 = ~x_768 & ~n_22731;
assign n_22826 = ~n_22732 & ~n_22825;
assign n_22827 = ~x_672 &  n_22826;
assign n_22828 =  x_672 & ~n_22826;
assign n_22829 = ~x_769 & ~n_22730;
assign n_22830 = ~n_22731 & ~n_22829;
assign n_22831 = ~x_673 &  n_22830;
assign n_22832 =  x_673 & ~n_22830;
assign n_22833 = ~x_770 & ~n_22729;
assign n_22834 = ~n_22730 & ~n_22833;
assign n_22835 = ~x_674 &  n_22834;
assign n_22836 = ~x_771 & ~n_22728;
assign n_22837 = ~n_22729 & ~n_22836;
assign n_22838 = ~x_675 &  n_22837;
assign n_22839 = ~x_772 & ~n_22727;
assign n_22840 = ~n_22728 & ~n_22839;
assign n_22841 =  x_676 & ~n_22840;
assign n_22842 = ~x_774 & ~n_22725;
assign n_22843 = ~n_22726 & ~n_22842;
assign n_22844 = ~x_678 &  n_22843;
assign n_22845 = ~x_775 & ~n_22724;
assign n_22846 = ~n_22725 & ~n_22845;
assign n_22847 =  x_679 & ~n_22846;
assign n_22848 = ~x_776 & ~n_22723;
assign n_22849 = ~n_22724 & ~n_22848;
assign n_22850 =  x_680 & ~n_22849;
assign n_22851 = ~x_777 & ~n_22722;
assign n_22852 = ~n_22723 & ~n_22851;
assign n_22853 = ~x_681 &  n_22852;
assign n_22854 =  x_681 & ~n_22852;
assign n_22855 =  x_682 & ~x_778;
assign n_22856 = ~n_22722 & ~n_22855;
assign n_22857 =  x_682 &  x_778;
assign n_22858 = ~x_683 &  x_779;
assign n_22859 = ~n_22857 &  n_22858;
assign n_22860 = ~n_22856 & ~n_22859;
assign n_22861 = ~n_22854 & ~n_22860;
assign n_22862 = ~n_22853 & ~n_22861;
assign n_22863 = ~n_22850 & ~n_22862;
assign n_22864 = ~x_680 &  n_22849;
assign n_22865 = ~x_679 &  n_22846;
assign n_22866 = ~n_22864 & ~n_22865;
assign n_22867 = ~n_22863 &  n_22866;
assign n_22868 = ~n_22847 & ~n_22867;
assign n_22869 = ~n_22844 & ~n_22868;
assign n_22870 =  x_678 & ~n_22843;
assign n_22871 = ~x_773 & ~n_22726;
assign n_22872 = ~n_22727 & ~n_22871;
assign n_22873 =  x_677 & ~n_22872;
assign n_22874 = ~n_22870 & ~n_22873;
assign n_22875 = ~n_22869 &  n_22874;
assign n_22876 = ~x_677 &  n_22872;
assign n_22877 = ~x_676 &  n_22840;
assign n_22878 = ~n_22876 & ~n_22877;
assign n_22879 = ~n_22875 &  n_22878;
assign n_22880 = ~n_22841 & ~n_22879;
assign n_22881 = ~n_22838 & ~n_22880;
assign n_22882 =  x_675 & ~n_22837;
assign n_22883 =  x_674 & ~n_22834;
assign n_22884 = ~n_22882 & ~n_22883;
assign n_22885 = ~n_22881 &  n_22884;
assign n_22886 = ~n_22835 & ~n_22885;
assign n_22887 = ~n_22832 & ~n_22886;
assign n_22888 = ~n_22831 & ~n_22887;
assign n_22889 = ~n_22828 & ~n_22888;
assign n_22890 = ~n_22827 & ~n_22889;
assign n_22891 = ~n_22824 & ~n_22890;
assign n_22892 = ~n_22823 & ~n_22891;
assign n_22893 = ~n_22820 & ~n_22892;
assign n_22894 = ~n_22819 & ~n_22893;
assign n_22895 = ~n_22816 & ~n_22894;
assign n_22896 = ~n_22815 & ~n_22895;
assign n_22897 = ~n_22812 & ~n_22896;
assign n_22898 = ~n_22811 & ~n_22897;
assign n_22899 = ~n_22808 & ~n_22898;
assign n_22900 = ~n_22807 & ~n_22899;
assign n_22901 = ~n_22804 & ~n_22900;
assign n_22902 = ~n_22803 & ~n_22901;
assign n_22903 = ~n_22800 & ~n_22902;
assign n_22904 = ~n_22799 & ~n_22903;
assign n_22905 = ~n_22796 & ~n_22904;
assign n_22906 = ~n_22795 & ~n_22905;
assign n_22907 = ~n_22792 & ~n_22906;
assign n_22908 = ~n_22791 & ~n_22907;
assign n_22909 = ~n_22788 & ~n_22908;
assign n_22910 = ~n_22787 & ~n_22909;
assign n_22911 = ~n_22784 & ~n_22910;
assign n_22912 = ~n_22783 & ~n_22911;
assign n_22913 = ~n_22780 & ~n_22912;
assign n_22914 = ~n_22779 & ~n_22913;
assign n_22915 = ~n_22776 & ~n_22914;
assign n_22916 = ~n_22775 & ~n_22915;
assign n_22917 = ~n_22772 & ~n_22916;
assign n_22918 = ~n_22771 & ~n_22917;
assign n_22919 = ~n_22768 & ~n_22918;
assign n_22920 = ~n_22767 & ~n_22919;
assign n_22921 = ~n_22764 & ~n_22920;
assign n_22922 = ~n_22763 & ~n_22921;
assign n_22923 = ~n_22760 & ~n_22922;
assign n_22924 = ~x_655 &  n_22759;
assign n_22925 = ~x_654 &  n_22756;
assign n_22926 = ~n_22924 & ~n_22925;
assign n_22927 = ~n_22923 &  n_22926;
assign n_22928 = ~n_22757 & ~n_22927;
assign n_22929 = ~n_22754 & ~n_22928;
assign n_22930 =  x_653 & ~n_22753;
assign n_22931 =  x_748 & ~n_22751;
assign n_22932 = ~x_652 &  n_22931;
assign n_22933 = ~n_22930 & ~n_22932;
assign n_22934 = ~n_22929 &  n_22933;
assign n_22935 =  x_652 & ~n_22931;
assign n_22936 = ~x_748 &  n_22751;
assign n_22937 = ~n_22935 & ~n_22936;
assign n_22938 = ~n_22934 &  n_22937;
assign n_22939 =  n_22721 & ~n_22938;
assign n_22940 =  n_2 &  n_5648;
assign n_22941 = ~x_1726 & ~x_1727;
assign n_22942 = ~x_1728 & ~x_1729;
assign n_22943 =  n_22941 &  n_22942;
assign n_22944 = ~x_1722 & ~x_1723;
assign n_22945 = ~x_1724 & ~x_1725;
assign n_22946 =  n_22944 &  n_22945;
assign n_22947 =  n_22943 &  n_22946;
assign n_22948 = ~x_1734 & ~x_1735;
assign n_22949 = ~x_1736 &  n_22948;
assign n_22950 = ~x_1730 & ~x_1731;
assign n_22951 = ~x_1732 & ~x_1733;
assign n_22952 =  n_22950 &  n_22951;
assign n_22953 =  n_22949 &  n_22952;
assign n_22954 =  n_22947 &  n_22953;
assign n_22955 = ~x_1708 & ~x_1709;
assign n_22956 = ~x_1710 & ~x_1711;
assign n_22957 = ~x_1712 & ~x_1713;
assign n_22958 =  n_22956 &  n_22957;
assign n_22959 =  n_22955 &  n_22958;
assign n_22960 = ~x_1718 & ~x_1719;
assign n_22961 = ~x_1720 & ~x_1721;
assign n_22962 =  n_22960 &  n_22961;
assign n_22963 = ~x_1714 & ~x_1715;
assign n_22964 = ~x_1716 & ~x_1717;
assign n_22965 =  n_22963 &  n_22964;
assign n_22966 =  n_22962 &  n_22965;
assign n_22967 =  n_22959 &  n_22966;
assign n_22968 =  n_22954 &  n_22967;
assign n_22969 = ~x_1737 &  n_22968;
assign n_22970 = ~x_1738 &  n_22969;
assign n_22971 = ~x_1707 & ~n_22970;
assign n_22972 =  n_150 &  n_22971;
assign n_22973 =  n_22940 &  n_22972;
assign n_22974 = ~x_4284 & ~x_4285;
assign n_22975 = ~x_4286 & ~x_4287;
assign n_22976 =  n_22974 &  n_22975;
assign n_22977 = ~x_4280 & ~x_4281;
assign n_22978 = ~x_4282 & ~x_4283;
assign n_22979 =  n_22977 &  n_22978;
assign n_22980 =  n_22976 &  n_22979;
assign n_22981 = ~x_4292 & ~x_4293;
assign n_22982 = ~x_4294 &  n_22981;
assign n_22983 = ~x_4288 & ~x_4289;
assign n_22984 = ~x_4290 & ~x_4291;
assign n_22985 =  n_22983 &  n_22984;
assign n_22986 =  n_22982 &  n_22985;
assign n_22987 =  n_22980 &  n_22986;
assign n_22988 = ~x_4266 & ~x_4267;
assign n_22989 = ~x_4268 & ~x_4269;
assign n_22990 = ~x_4270 & ~x_4271;
assign n_22991 =  n_22989 &  n_22990;
assign n_22992 =  n_22988 &  n_22991;
assign n_22993 = ~x_4276 & ~x_4277;
assign n_22994 = ~x_4278 & ~x_4279;
assign n_22995 =  n_22993 &  n_22994;
assign n_22996 = ~x_4272 & ~x_4273;
assign n_22997 = ~x_4274 & ~x_4275;
assign n_22998 =  n_22996 &  n_22997;
assign n_22999 =  n_22995 &  n_22998;
assign n_23000 =  n_22992 &  n_22999;
assign n_23001 =  n_22987 &  n_23000;
assign n_23002 = ~x_4295 &  n_23001;
assign n_23003 = ~x_4296 &  n_23002;
assign n_23004 = ~x_4265 & ~n_23003;
assign n_23005 =  n_12 &  n_556;
assign n_23006 =  n_11 &  n_23005;
assign n_23007 =  n_23006 &  n_2486;
assign n_23008 =  n_23004 &  n_23007;
assign n_23009 =  x_33 &  x_34;
assign n_23010 =  x_1771 &  n_23009;
assign n_23011 =  n_149 &  n_23010;
assign n_23012 =  n_12 &  n_1896;
assign n_23013 =  n_11 &  n_23012;
assign n_23014 =  n_23011 &  n_23013;
assign n_23015 = ~n_23008 & ~n_23014;
assign n_23016 = ~n_22973 &  n_23015;
assign n_23017 = ~x_3932 & ~x_3933;
assign n_23018 = ~x_3934 & ~x_3935;
assign n_23019 =  n_23017 &  n_23018;
assign n_23020 = ~x_3928 & ~x_3929;
assign n_23021 = ~x_3930 & ~x_3931;
assign n_23022 =  n_23020 &  n_23021;
assign n_23023 =  n_23019 &  n_23022;
assign n_23024 = ~x_3940 & ~x_3941;
assign n_23025 = ~x_3942 &  n_23024;
assign n_23026 = ~x_3936 & ~x_3937;
assign n_23027 = ~x_3938 & ~x_3939;
assign n_23028 =  n_23026 &  n_23027;
assign n_23029 =  n_23025 &  n_23028;
assign n_23030 =  n_23023 &  n_23029;
assign n_23031 = ~x_3914 & ~x_3915;
assign n_23032 = ~x_3916 & ~x_3917;
assign n_23033 = ~x_3918 & ~x_3919;
assign n_23034 =  n_23032 &  n_23033;
assign n_23035 =  n_23031 &  n_23034;
assign n_23036 = ~x_3924 & ~x_3925;
assign n_23037 = ~x_3926 & ~x_3927;
assign n_23038 =  n_23036 &  n_23037;
assign n_23039 = ~x_3920 & ~x_3921;
assign n_23040 = ~x_3922 & ~x_3923;
assign n_23041 =  n_23039 &  n_23040;
assign n_23042 =  n_23038 &  n_23041;
assign n_23043 =  n_23035 &  n_23042;
assign n_23044 =  n_23030 &  n_23043;
assign n_23045 =  x_3943 &  x_3944;
assign n_23046 =  n_23044 & ~n_23045;
assign n_23047 = ~x_3913 & ~n_23046;
assign n_23048 =  n_15366 &  n_6182;
assign n_23049 = ~n_23047 &  n_23048;
assign n_23050 =  x_38 &  n_2683;
assign n_23051 =  x_3416 &  n_21952;
assign n_23052 =  n_23050 &  n_23051;
assign n_23053 =  n_23052 &  n_7855;
assign n_23054 = ~n_23049 & ~n_23053;
assign n_23055 =  x_1737 &  x_1738;
assign n_23056 =  n_22968 & ~n_23055;
assign n_23057 = ~x_1707 & ~n_23056;
assign n_23058 =  n_4089 &  n_4290;
assign n_23059 = ~n_23057 &  n_23058;
assign n_23060 = ~x_1707 & ~n_22969;
assign n_23061 =  n_1173 &  n_21564;
assign n_23062 = ~n_23060 &  n_23061;
assign n_23063 = ~n_23059 & ~n_23062;
assign n_23064 =  n_23054 &  n_23063;
assign n_23065 =  n_2879 &  n_5656;
assign n_23066 =  n_1040 &  n_23065;
assign n_23067 =  n_2879 &  n_14263;
assign n_23068 = ~x_2606 & ~x_2607;
assign n_23069 = ~x_2608 & ~x_2609;
assign n_23070 =  n_23068 &  n_23069;
assign n_23071 = ~x_2602 & ~x_2603;
assign n_23072 = ~x_2604 & ~x_2605;
assign n_23073 =  n_23071 &  n_23072;
assign n_23074 =  n_23070 &  n_23073;
assign n_23075 = ~x_2614 & ~x_2615;
assign n_23076 = ~x_2616 &  n_23075;
assign n_23077 = ~x_2610 & ~x_2611;
assign n_23078 = ~x_2612 & ~x_2613;
assign n_23079 =  n_23077 &  n_23078;
assign n_23080 =  n_23076 &  n_23079;
assign n_23081 =  n_23074 &  n_23080;
assign n_23082 = ~x_2588 & ~x_2589;
assign n_23083 = ~x_2590 & ~x_2591;
assign n_23084 = ~x_2592 & ~x_2593;
assign n_23085 =  n_23083 &  n_23084;
assign n_23086 =  n_23082 &  n_23085;
assign n_23087 = ~x_2598 & ~x_2599;
assign n_23088 = ~x_2600 & ~x_2601;
assign n_23089 =  n_23087 &  n_23088;
assign n_23090 = ~x_2594 & ~x_2595;
assign n_23091 = ~x_2596 & ~x_2597;
assign n_23092 =  n_23090 &  n_23091;
assign n_23093 =  n_23089 &  n_23092;
assign n_23094 =  n_23086 &  n_23093;
assign n_23095 =  n_23081 &  n_23094;
assign n_23096 =  x_2617 &  x_2618;
assign n_23097 =  n_23095 & ~n_23096;
assign n_23098 = ~x_2587 & ~n_23097;
assign n_23099 =  n_1040 &  n_23098;
assign n_23100 =  n_23067 &  n_23099;
assign n_23101 = ~n_23066 & ~n_23100;
assign n_23102 =  n_23064 &  n_23101;
assign n_23103 =  n_23016 &  n_23102;
assign n_23104 = ~x_3692 & ~x_3693;
assign n_23105 = ~x_3694 & ~x_3695;
assign n_23106 =  n_23104 &  n_23105;
assign n_23107 = ~x_3688 & ~x_3689;
assign n_23108 = ~x_3690 & ~x_3691;
assign n_23109 =  n_23107 &  n_23108;
assign n_23110 =  n_23106 &  n_23109;
assign n_23111 = ~x_3700 & ~x_3701;
assign n_23112 = ~x_3702 & ~x_3703;
assign n_23113 =  n_23111 &  n_23112;
assign n_23114 = ~x_3696 & ~x_3697;
assign n_23115 = ~x_3698 & ~x_3699;
assign n_23116 =  n_23114 &  n_23115;
assign n_23117 =  n_23113 &  n_23116;
assign n_23118 =  n_23110 &  n_23117;
assign n_23119 = ~x_3676 & ~x_3677;
assign n_23120 = ~x_3678 & ~x_3679;
assign n_23121 =  n_23119 &  n_23120;
assign n_23122 = ~x_3672 & ~x_3673;
assign n_23123 = ~x_3674 & ~x_3675;
assign n_23124 =  n_23122 &  n_23123;
assign n_23125 =  n_23121 &  n_23124;
assign n_23126 = ~x_3684 & ~x_3685;
assign n_23127 = ~x_3686 & ~x_3687;
assign n_23128 =  n_23126 &  n_23127;
assign n_23129 = ~x_3680 & ~x_3681;
assign n_23130 = ~x_3682 & ~x_3683;
assign n_23131 =  n_23129 &  n_23130;
assign n_23132 =  n_23128 &  n_23131;
assign n_23133 =  n_23125 &  n_23132;
assign n_23134 =  n_23118 &  n_23133;
assign n_23135 = ~x_39 &  n_15366;
assign n_23136 =  n_23135 &  n_1698;
assign n_23137 = ~n_23134 &  n_23136;
assign n_23138 =  n_2290 &  n_351;
assign n_23139 =  n_552 &  n_23138;
assign n_23140 =  n_8054 &  n_10276;
assign n_23141 = ~n_23139 & ~n_23140;
assign n_23142 = ~n_23137 &  n_23141;
assign n_23143 = ~x_1535 & ~x_1536;
assign n_23144 = ~x_1537 & ~x_1538;
assign n_23145 =  n_23143 &  n_23144;
assign n_23146 = ~x_1531 & ~x_1532;
assign n_23147 = ~x_1533 & ~x_1534;
assign n_23148 =  n_23146 &  n_23147;
assign n_23149 =  n_23145 &  n_23148;
assign n_23150 = ~x_1543 & ~x_1544;
assign n_23151 = ~x_1545 & ~x_1546;
assign n_23152 =  n_23150 &  n_23151;
assign n_23153 = ~x_1539 & ~x_1540;
assign n_23154 = ~x_1541 & ~x_1542;
assign n_23155 =  n_23153 &  n_23154;
assign n_23156 =  n_23152 &  n_23155;
assign n_23157 =  n_23149 &  n_23156;
assign n_23158 = ~x_1519 & ~x_1520;
assign n_23159 = ~x_1521 & ~x_1522;
assign n_23160 =  n_23158 &  n_23159;
assign n_23161 = ~x_1515 & ~x_1516;
assign n_23162 = ~x_1517 & ~x_1518;
assign n_23163 =  n_23161 &  n_23162;
assign n_23164 =  n_23160 &  n_23163;
assign n_23165 = ~x_1527 & ~x_1528;
assign n_23166 = ~x_1529 & ~x_1530;
assign n_23167 =  n_23165 &  n_23166;
assign n_23168 = ~x_1523 & ~x_1524;
assign n_23169 = ~x_1525 & ~x_1526;
assign n_23170 =  n_23168 &  n_23169;
assign n_23171 =  n_23167 &  n_23170;
assign n_23172 =  n_23164 &  n_23171;
assign n_23173 =  n_23157 &  n_23172;
assign n_23174 =  x_43 &  n_3341;
assign n_23175 =  n_5648 &  n_3615;
assign n_23176 =  n_23174 &  n_23175;
assign n_23177 =  n_23173 &  n_23176;
assign n_23178 =  n_5648 &  n_3143;
assign n_23179 =  n_23178 &  n_3615;
assign n_23180 = ~x_1471 & ~x_1472;
assign n_23181 = ~x_1473 & ~x_1474;
assign n_23182 =  n_23180 &  n_23181;
assign n_23183 = ~x_1467 & ~x_1468;
assign n_23184 = ~x_1469 & ~x_1470;
assign n_23185 =  n_23183 &  n_23184;
assign n_23186 =  n_23182 &  n_23185;
assign n_23187 = ~x_1479 & ~x_1480;
assign n_23188 = ~x_1481 & ~x_1482;
assign n_23189 =  n_23187 &  n_23188;
assign n_23190 = ~x_1475 & ~x_1476;
assign n_23191 = ~x_1477 & ~x_1478;
assign n_23192 =  n_23190 &  n_23191;
assign n_23193 =  n_23189 &  n_23192;
assign n_23194 =  n_23186 &  n_23193;
assign n_23195 = ~x_1455 & ~x_1456;
assign n_23196 = ~x_1457 & ~x_1458;
assign n_23197 =  n_23195 &  n_23196;
assign n_23198 = ~x_1451 & ~x_1452;
assign n_23199 = ~x_1453 & ~x_1454;
assign n_23200 =  n_23198 &  n_23199;
assign n_23201 =  n_23197 &  n_23200;
assign n_23202 = ~x_1463 & ~x_1464;
assign n_23203 = ~x_1465 & ~x_1466;
assign n_23204 =  n_23202 &  n_23203;
assign n_23205 = ~x_1459 & ~x_1460;
assign n_23206 = ~x_1461 & ~x_1462;
assign n_23207 =  n_23205 &  n_23206;
assign n_23208 =  n_23204 &  n_23207;
assign n_23209 =  n_23201 &  n_23208;
assign n_23210 =  n_23194 &  n_23209;
assign n_23211 =  n_23179 &  n_23210;
assign n_23212 = ~n_23177 & ~n_23211;
assign n_23213 =  n_23142 &  n_23212;
assign n_23214 = ~x_3564 & ~x_3565;
assign n_23215 = ~x_3566 & ~x_3567;
assign n_23216 =  n_23214 &  n_23215;
assign n_23217 = ~x_3560 & ~x_3561;
assign n_23218 = ~x_3562 & ~x_3563;
assign n_23219 =  n_23217 &  n_23218;
assign n_23220 =  n_23216 &  n_23219;
assign n_23221 = ~x_3572 & ~x_3573;
assign n_23222 = ~x_3574 & ~x_3575;
assign n_23223 =  n_23221 &  n_23222;
assign n_23224 = ~x_3568 & ~x_3569;
assign n_23225 = ~x_3570 & ~x_3571;
assign n_23226 =  n_23224 &  n_23225;
assign n_23227 =  n_23223 &  n_23226;
assign n_23228 =  n_23220 &  n_23227;
assign n_23229 = ~x_3548 & ~x_3549;
assign n_23230 = ~x_3550 & ~x_3551;
assign n_23231 =  n_23229 &  n_23230;
assign n_23232 = ~x_3544 & ~x_3545;
assign n_23233 = ~x_3546 & ~x_3547;
assign n_23234 =  n_23232 &  n_23233;
assign n_23235 =  n_23231 &  n_23234;
assign n_23236 = ~x_3556 & ~x_3557;
assign n_23237 = ~x_3558 & ~x_3559;
assign n_23238 =  n_23236 &  n_23237;
assign n_23239 = ~x_3552 & ~x_3553;
assign n_23240 = ~x_3554 & ~x_3555;
assign n_23241 =  n_23239 &  n_23240;
assign n_23242 =  n_23238 &  n_23241;
assign n_23243 =  n_23235 &  n_23242;
assign n_23244 =  n_23228 &  n_23243;
assign n_23245 =  n_6379 &  n_10475;
assign n_23246 =  n_23244 &  n_23245;
assign n_23247 =  n_19497 &  n_10872;
assign n_23248 = ~n_23247 & ~n_20984;
assign n_23249 = ~n_23246 &  n_23248;
assign n_23250 =  n_23213 &  n_23249;
assign n_23251 =  n_21758 &  n_3615;
assign n_23252 =  n_1038 &  n_1174;
assign n_23253 = ~x_38 &  n_23252;
assign n_23254 =  n_23253 &  n_3615;
assign n_23255 =  n_5645 &  n_23175;
assign n_23256 = ~n_23254 & ~n_23255;
assign n_23257 = ~n_23251 &  n_23256;
assign n_23258 = ~n_9885 &  n_23257;
assign n_23259 =  n_23067 &  n_1040;
assign n_23260 = ~n_23098 &  n_23259;
assign n_23261 =  n_23258 & ~n_23260;
assign n_23262 =  n_23250 &  n_23261;
assign n_23263 = ~x_1694 & ~x_1695;
assign n_23264 = ~x_1696 & ~x_1697;
assign n_23265 =  n_23263 &  n_23264;
assign n_23266 = ~x_1690 & ~x_1691;
assign n_23267 = ~x_1692 & ~x_1693;
assign n_23268 =  n_23266 &  n_23267;
assign n_23269 =  n_23265 &  n_23268;
assign n_23270 = ~x_1702 & ~x_1703;
assign n_23271 = ~x_1704 &  n_23270;
assign n_23272 = ~x_1698 & ~x_1699;
assign n_23273 = ~x_1700 & ~x_1701;
assign n_23274 =  n_23272 &  n_23273;
assign n_23275 =  n_23271 &  n_23274;
assign n_23276 =  n_23269 &  n_23275;
assign n_23277 = ~x_1676 & ~x_1677;
assign n_23278 = ~x_1678 & ~x_1679;
assign n_23279 = ~x_1680 & ~x_1681;
assign n_23280 =  n_23278 &  n_23279;
assign n_23281 =  n_23277 &  n_23280;
assign n_23282 = ~x_1686 & ~x_1687;
assign n_23283 = ~x_1688 & ~x_1689;
assign n_23284 =  n_23282 &  n_23283;
assign n_23285 = ~x_1682 & ~x_1683;
assign n_23286 = ~x_1684 & ~x_1685;
assign n_23287 =  n_23285 &  n_23286;
assign n_23288 =  n_23284 &  n_23287;
assign n_23289 =  n_23281 &  n_23288;
assign n_23290 =  n_23276 &  n_23289;
assign n_23291 = ~x_1705 &  n_23290;
assign n_23292 = ~x_1675 & ~n_23291;
assign n_23293 =  n_16495 &  n_1502;
assign n_23294 =  n_23292 &  n_23293;
assign n_23295 = ~x_2334 & ~x_2335;
assign n_23296 = ~x_2336 & ~x_2337;
assign n_23297 =  n_23295 &  n_23296;
assign n_23298 = ~x_2330 & ~x_2331;
assign n_23299 = ~x_2332 & ~x_2333;
assign n_23300 =  n_23298 &  n_23299;
assign n_23301 =  n_23297 &  n_23300;
assign n_23302 = ~x_2342 & ~x_2343;
assign n_23303 = ~x_2344 &  n_23302;
assign n_23304 = ~x_2338 & ~x_2339;
assign n_23305 = ~x_2340 & ~x_2341;
assign n_23306 =  n_23304 &  n_23305;
assign n_23307 =  n_23303 &  n_23306;
assign n_23308 =  n_23301 &  n_23307;
assign n_23309 = ~x_2316 & ~x_2317;
assign n_23310 = ~x_2318 & ~x_2319;
assign n_23311 = ~x_2320 & ~x_2321;
assign n_23312 =  n_23310 &  n_23311;
assign n_23313 =  n_23309 &  n_23312;
assign n_23314 = ~x_2326 & ~x_2327;
assign n_23315 = ~x_2328 & ~x_2329;
assign n_23316 =  n_23314 &  n_23315;
assign n_23317 = ~x_2322 & ~x_2323;
assign n_23318 = ~x_2324 & ~x_2325;
assign n_23319 =  n_23317 &  n_23318;
assign n_23320 =  n_23316 &  n_23319;
assign n_23321 =  n_23313 &  n_23320;
assign n_23322 =  n_23308 &  n_23321;
assign n_23323 =  x_2345 &  x_2346;
assign n_23324 =  n_23322 & ~n_23323;
assign n_23325 = ~x_2315 & ~n_23324;
assign n_23326 =  n_557 &  n_355;
assign n_23327 =  n_23325 &  n_23326;
assign n_23328 = ~n_23294 & ~n_23327;
assign n_23329 =  x_40 &  n_23174;
assign n_23330 =  n_17784 &  n_23329;
assign n_23331 =  n_19493 &  n_7467;
assign n_23332 = ~n_23330 & ~n_23331;
assign n_23333 =  n_10478 &  n_3615;
assign n_23334 = ~x_1247 & ~x_1248;
assign n_23335 = ~x_1249 & ~x_1250;
assign n_23336 =  n_23334 &  n_23335;
assign n_23337 = ~x_1243 & ~x_1244;
assign n_23338 = ~x_1245 & ~x_1246;
assign n_23339 =  n_23337 &  n_23338;
assign n_23340 =  n_23336 &  n_23339;
assign n_23341 = ~x_1255 & ~x_1256;
assign n_23342 = ~x_1257 & ~x_1258;
assign n_23343 =  n_23341 &  n_23342;
assign n_23344 = ~x_1251 & ~x_1252;
assign n_23345 = ~x_1253 & ~x_1254;
assign n_23346 =  n_23344 &  n_23345;
assign n_23347 =  n_23343 &  n_23346;
assign n_23348 =  n_23340 &  n_23347;
assign n_23349 = ~x_1231 & ~x_1232;
assign n_23350 = ~x_1233 & ~x_1234;
assign n_23351 =  n_23349 &  n_23350;
assign n_23352 = ~x_1227 & ~x_1228;
assign n_23353 = ~x_1229 & ~x_1230;
assign n_23354 =  n_23352 &  n_23353;
assign n_23355 =  n_23351 &  n_23354;
assign n_23356 = ~x_1239 & ~x_1240;
assign n_23357 = ~x_1241 & ~x_1242;
assign n_23358 =  n_23356 &  n_23357;
assign n_23359 = ~x_1235 & ~x_1236;
assign n_23360 = ~x_1237 & ~x_1238;
assign n_23361 =  n_23359 &  n_23360;
assign n_23362 =  n_23358 &  n_23361;
assign n_23363 =  n_23355 &  n_23362;
assign n_23364 =  n_23348 &  n_23363;
assign n_23365 =  n_23333 & ~n_23364;
assign n_23366 = ~n_23173 &  n_23176;
assign n_23367 = ~n_23365 & ~n_23366;
assign n_23368 =  n_23332 &  n_23367;
assign n_23369 =  n_6525 &  n_357;
assign n_23370 = ~n_23369 & ~n_1701;
assign n_23371 =  n_23368 &  n_23370;
assign n_23372 =  n_23328 &  n_23371;
assign n_23373 =  n_23262 &  n_23372;
assign n_23374 = ~x_38 &  n_4285;
assign n_23375 =  n_349 &  n_23374;
assign n_23376 = ~n_23375 & ~n_23013;
assign n_23377 =  n_17782 & ~n_23376;
assign n_23378 =  n_552 &  n_5652;
assign n_23379 = ~n_23377 & ~n_23378;
assign n_23380 = ~n_16882 &  n_23379;
assign n_23381 =  n_1039 &  n_353;
assign n_23382 =  x_37 &  n_23381;
assign n_23383 =  n_561 &  n_556;
assign n_23384 =  n_23382 &  n_23383;
assign n_23385 = ~x_43 & ~x_1771;
assign n_23386 =  n_23384 &  n_23385;
assign n_23387 = ~x_42 &  n_23386;
assign n_23388 =  n_554 &  n_3141;
assign n_23389 =  n_23388 &  n_3628;
assign n_23390 = ~x_4636 & ~x_4637;
assign n_23391 = ~x_4638 & ~x_4639;
assign n_23392 =  n_23390 &  n_23391;
assign n_23393 = ~x_4632 & ~x_4633;
assign n_23394 = ~x_4634 & ~x_4635;
assign n_23395 =  n_23393 &  n_23394;
assign n_23396 =  n_23392 &  n_23395;
assign n_23397 = ~x_4644 & ~x_4645;
assign n_23398 = ~x_4646 & ~x_4647;
assign n_23399 =  n_23397 &  n_23398;
assign n_23400 = ~x_4640 & ~x_4641;
assign n_23401 = ~x_4642 & ~x_4643;
assign n_23402 =  n_23400 &  n_23401;
assign n_23403 =  n_23399 &  n_23402;
assign n_23404 =  n_23396 &  n_23403;
assign n_23405 = ~x_4620 & ~x_4621;
assign n_23406 = ~x_4622 & ~x_4623;
assign n_23407 =  n_23405 &  n_23406;
assign n_23408 = ~x_4616 & ~x_4617;
assign n_23409 = ~x_4618 & ~x_4619;
assign n_23410 =  n_23408 &  n_23409;
assign n_23411 =  n_23407 &  n_23410;
assign n_23412 = ~x_4628 & ~x_4629;
assign n_23413 = ~x_4630 & ~x_4631;
assign n_23414 =  n_23412 &  n_23413;
assign n_23415 = ~x_4624 & ~x_4625;
assign n_23416 = ~x_4626 & ~x_4627;
assign n_23417 =  n_23415 &  n_23416;
assign n_23418 =  n_23414 &  n_23417;
assign n_23419 =  n_23411 &  n_23418;
assign n_23420 =  n_23404 &  n_23419;
assign n_23421 =  n_23389 &  n_23420;
assign n_23422 =  n_11 &  n_8347;
assign n_23423 =  n_6882 &  n_23422;
assign n_23424 = ~x_4668 & ~x_4669;
assign n_23425 = ~x_4670 & ~x_4671;
assign n_23426 =  n_23424 &  n_23425;
assign n_23427 = ~x_4664 & ~x_4665;
assign n_23428 = ~x_4666 & ~x_4667;
assign n_23429 =  n_23427 &  n_23428;
assign n_23430 =  n_23426 &  n_23429;
assign n_23431 = ~x_4676 & ~x_4677;
assign n_23432 = ~x_4678 & ~x_4679;
assign n_23433 =  n_23431 &  n_23432;
assign n_23434 = ~x_4672 & ~x_4673;
assign n_23435 = ~x_4674 & ~x_4675;
assign n_23436 =  n_23434 &  n_23435;
assign n_23437 =  n_23433 &  n_23436;
assign n_23438 =  n_23430 &  n_23437;
assign n_23439 = ~x_4652 & ~x_4653;
assign n_23440 = ~x_4654 & ~x_4655;
assign n_23441 =  n_23439 &  n_23440;
assign n_23442 = ~x_4648 & ~x_4649;
assign n_23443 = ~x_4650 & ~x_4651;
assign n_23444 =  n_23442 &  n_23443;
assign n_23445 =  n_23441 &  n_23444;
assign n_23446 = ~x_4660 & ~x_4661;
assign n_23447 = ~x_4662 & ~x_4663;
assign n_23448 =  n_23446 &  n_23447;
assign n_23449 = ~x_4656 & ~x_4657;
assign n_23450 = ~x_4658 & ~x_4659;
assign n_23451 =  n_23449 &  n_23450;
assign n_23452 =  n_23448 &  n_23451;
assign n_23453 =  n_23445 &  n_23452;
assign n_23454 =  n_23438 &  n_23453;
assign n_23455 =  n_23423 & ~n_23454;
assign n_23456 = ~n_23421 & ~n_23455;
assign n_23457 = ~n_23387 &  n_23456;
assign n_23458 =  n_23380 &  n_23457;
assign n_23459 = ~x_35 &  n_23009;
assign n_23460 = ~x_36 &  n_23459;
assign n_23461 =  n_349 &  n_23460;
assign n_23462 =  n_2879 &  n_4285;
assign n_23463 =  n_23461 &  n_23462;
assign n_23464 = ~x_1547 &  n_23463;
assign n_23465 =  n_12 &  n_768;
assign n_23466 =  x_3416 &  n_23381;
assign n_23467 =  n_23465 &  n_23466;
assign n_23468 =  n_11 &  n_23467;
assign n_23469 =  n_23253 &  n_1502;
assign n_23470 = ~n_23468 & ~n_23469;
assign n_23471 = ~n_10472 &  n_23470;
assign n_23472 = ~n_23464 &  n_23471;
assign n_23473 =  n_150 &  n_21758;
assign n_23474 =  n_23060 &  n_23473;
assign n_23475 =  n_23472 & ~n_23474;
assign n_23476 =  n_23458 &  n_23475;
assign n_23477 =  n_760 &  n_15;
assign n_23478 = ~x_64 & ~x_65;
assign n_23479 = ~x_66 & ~x_67;
assign n_23480 =  n_23478 &  n_23479;
assign n_23481 = ~x_60 & ~x_61;
assign n_23482 = ~x_62 & ~x_63;
assign n_23483 =  n_23481 &  n_23482;
assign n_23484 =  n_23480 &  n_23483;
assign n_23485 = ~x_72 & ~x_73;
assign n_23486 = ~x_74 & ~x_75;
assign n_23487 =  n_23485 &  n_23486;
assign n_23488 = ~x_68 & ~x_69;
assign n_23489 = ~x_70 & ~x_71;
assign n_23490 =  n_23488 &  n_23489;
assign n_23491 =  n_23487 &  n_23490;
assign n_23492 =  n_23484 &  n_23491;
assign n_23493 = ~x_48 & ~x_49;
assign n_23494 = ~x_50 & ~x_51;
assign n_23495 =  n_23493 &  n_23494;
assign n_23496 = ~x_44 & ~x_45;
assign n_23497 = ~x_46 & ~x_47;
assign n_23498 =  n_23496 &  n_23497;
assign n_23499 =  n_23495 &  n_23498;
assign n_23500 = ~x_56 & ~x_57;
assign n_23501 = ~x_58 & ~x_59;
assign n_23502 =  n_23500 &  n_23501;
assign n_23503 = ~x_52 & ~x_53;
assign n_23504 = ~x_54 & ~x_55;
assign n_23505 =  n_23503 &  n_23504;
assign n_23506 =  n_23502 &  n_23505;
assign n_23507 =  n_23499 &  n_23506;
assign n_23508 =  n_23492 &  n_23507;
assign n_23509 =  n_23477 &  n_23508;
assign n_23510 = ~x_96 & ~x_97;
assign n_23511 = ~x_98 & ~x_99;
assign n_23512 =  n_23510 &  n_23511;
assign n_23513 = ~x_92 & ~x_93;
assign n_23514 = ~x_94 & ~x_95;
assign n_23515 =  n_23513 &  n_23514;
assign n_23516 =  n_23512 &  n_23515;
assign n_23517 = ~x_104 & ~x_105;
assign n_23518 = ~x_106 & ~x_107;
assign n_23519 =  n_23517 &  n_23518;
assign n_23520 = ~x_100 & ~x_101;
assign n_23521 = ~x_102 & ~x_103;
assign n_23522 =  n_23520 &  n_23521;
assign n_23523 =  n_23519 &  n_23522;
assign n_23524 =  n_23516 &  n_23523;
assign n_23525 = ~x_80 & ~x_81;
assign n_23526 = ~x_82 & ~x_83;
assign n_23527 =  n_23525 &  n_23526;
assign n_23528 = ~x_76 & ~x_77;
assign n_23529 = ~x_78 & ~x_79;
assign n_23530 =  n_23528 &  n_23529;
assign n_23531 =  n_23527 &  n_23530;
assign n_23532 = ~x_88 & ~x_89;
assign n_23533 = ~x_90 & ~x_91;
assign n_23534 =  n_23532 &  n_23533;
assign n_23535 = ~x_84 & ~x_85;
assign n_23536 = ~x_86 & ~x_87;
assign n_23537 =  n_23535 &  n_23536;
assign n_23538 =  n_23534 &  n_23537;
assign n_23539 =  n_23531 &  n_23538;
assign n_23540 =  n_23524 &  n_23539;
assign n_23541 =  n_23252 &  n_7079;
assign n_23542 =  n_23540 &  n_23541;
assign n_23543 = ~n_23509 & ~n_23542;
assign n_23544 =  n_23253 &  n_8359;
assign n_23545 =  n_8359 &  n_10475;
assign n_23546 = ~n_23544 & ~n_23545;
assign n_23547 =  n_23543 &  n_23546;
assign n_23548 =  n_765 &  n_767;
assign n_23549 =  n_1174 &  n_3143;
assign n_23550 =  n_23548 &  n_23549;
assign n_23551 = ~n_23550 & ~n_14787;
assign n_23552 =  n_23547 &  n_23551;
assign n_23553 = ~x_38 &  n_8352;
assign n_23554 =  n_1037 &  n_23553;
assign n_23555 =  n_23554 &  n_1502;
assign n_23556 = ~x_1675 & ~n_23290;
assign n_23557 =  n_23555 & ~n_23556;
assign n_23558 =  n_13870 &  n_15;
assign n_23559 = ~n_23558 & ~n_10870;
assign n_23560 = ~n_23557 &  n_23559;
assign n_23561 =  n_2 &  n_5646;
assign n_23562 = ~x_4317 & ~x_4318;
assign n_23563 = ~x_4319 & ~x_4320;
assign n_23564 =  n_23562 &  n_23563;
assign n_23565 = ~x_4313 & ~x_4314;
assign n_23566 = ~x_4315 & ~x_4316;
assign n_23567 =  n_23565 &  n_23566;
assign n_23568 =  n_23564 &  n_23567;
assign n_23569 = ~x_4325 & ~x_4326;
assign n_23570 = ~x_4327 & ~x_4328;
assign n_23571 =  n_23569 &  n_23570;
assign n_23572 = ~x_4321 & ~x_4322;
assign n_23573 = ~x_4323 & ~x_4324;
assign n_23574 =  n_23572 &  n_23573;
assign n_23575 =  n_23571 &  n_23574;
assign n_23576 =  n_23568 &  n_23575;
assign n_23577 = ~x_4301 & ~x_4302;
assign n_23578 = ~x_4303 & ~x_4304;
assign n_23579 =  n_23577 &  n_23578;
assign n_23580 = ~x_4297 & ~x_4298;
assign n_23581 = ~x_4299 & ~x_4300;
assign n_23582 =  n_23580 &  n_23581;
assign n_23583 =  n_23579 &  n_23582;
assign n_23584 = ~x_4309 & ~x_4310;
assign n_23585 = ~x_4311 & ~x_4312;
assign n_23586 =  n_23584 &  n_23585;
assign n_23587 = ~x_4305 & ~x_4306;
assign n_23588 = ~x_4307 & ~x_4308;
assign n_23589 =  n_23587 &  n_23588;
assign n_23590 =  n_23586 &  n_23589;
assign n_23591 =  n_23583 &  n_23590;
assign n_23592 =  n_23576 &  n_23591;
assign n_23593 =  n_23561 &  n_23592;
assign n_23594 =  n_1041 &  n_9690;
assign n_23595 =  n_4288 &  n_23594;
assign n_23596 =  x_37 &  n_22715;
assign n_23597 =  x_3416 &  n_23596;
assign n_23598 =  n_20790 &  n_23597;
assign n_23599 = ~n_23595 & ~n_23598;
assign n_23600 = ~n_23593 &  n_23599;
assign n_23601 =  n_23560 &  n_23600;
assign n_23602 =  n_23552 &  n_23601;
assign n_23603 =  n_23476 &  n_23602;
assign n_23604 =  n_23373 &  n_23603;
assign n_23605 =  n_23103 &  n_23604;
assign n_23606 = ~x_39 &  n_2879;
assign n_23607 =  n_1040 &  n_23606;
assign n_23608 =  n_8344 &  n_23607;
assign n_23609 = ~x_2617 &  n_23095;
assign n_23610 = ~x_2587 & ~n_23609;
assign n_23611 =  n_23608 & ~n_23610;
assign n_23612 = ~x_1771 &  n_23009;
assign n_23613 =  n_149 &  n_23612;
assign n_23614 = ~x_43 &  n_23012;
assign n_23615 =  n_23613 &  n_23614;
assign n_23616 = ~x_42 &  n_23615;
assign n_23617 =  n_10872 &  n_23606;
assign n_23618 = ~x_3913 & ~n_23044;
assign n_23619 =  n_5 & ~n_23618;
assign n_23620 =  n_23617 &  n_23619;
assign n_23621 = ~n_23616 & ~n_23620;
assign n_23622 = ~n_23611 &  n_23621;
assign n_23623 =  n_23011 &  n_13866;
assign n_23624 =  n_1040 &  n_3144;
assign n_23625 =  n_23624 &  n_23610;
assign n_23626 = ~n_23623 & ~n_23625;
assign n_23627 = ~n_23004 &  n_23007;
assign n_23628 = ~x_3943 &  n_23044;
assign n_23629 = ~x_3944 &  n_23628;
assign n_23630 = ~x_3913 & ~n_23629;
assign n_23631 =  n_6379 &  n_13672;
assign n_23632 =  n_23630 &  n_23631;
assign n_23633 = ~n_23627 & ~n_23632;
assign n_23634 =  n_23626 &  n_23633;
assign n_23635 =  n_23622 &  n_23634;
assign n_23636 =  n_349 &  n_23005;
assign n_23637 = ~x_1706 &  n_23291;
assign n_23638 = ~x_1675 & ~n_23637;
assign n_23639 =  n_1502 & ~n_23638;
assign n_23640 =  n_23636 &  n_23639;
assign n_23641 =  n_2683 &  n_23553;
assign n_23642 =  n_23051 &  n_23641;
assign n_23643 =  n_11 &  n_23642;
assign n_23644 = ~x_3596 & ~x_3597;
assign n_23645 = ~x_3598 & ~x_3599;
assign n_23646 =  n_23644 &  n_23645;
assign n_23647 = ~x_3592 & ~x_3593;
assign n_23648 = ~x_3594 & ~x_3595;
assign n_23649 =  n_23647 &  n_23648;
assign n_23650 =  n_23646 &  n_23649;
assign n_23651 = ~x_3604 & ~x_3605;
assign n_23652 = ~x_3606 & ~x_3607;
assign n_23653 =  n_23651 &  n_23652;
assign n_23654 = ~x_3600 & ~x_3601;
assign n_23655 = ~x_3602 & ~x_3603;
assign n_23656 =  n_23654 &  n_23655;
assign n_23657 =  n_23653 &  n_23656;
assign n_23658 =  n_23650 &  n_23657;
assign n_23659 = ~x_3580 & ~x_3581;
assign n_23660 = ~x_3582 & ~x_3583;
assign n_23661 =  n_23659 &  n_23660;
assign n_23662 = ~x_3576 & ~x_3577;
assign n_23663 = ~x_3578 & ~x_3579;
assign n_23664 =  n_23662 &  n_23663;
assign n_23665 =  n_23661 &  n_23664;
assign n_23666 = ~x_3588 & ~x_3589;
assign n_23667 = ~x_3590 & ~x_3591;
assign n_23668 =  n_23666 &  n_23667;
assign n_23669 = ~x_3584 & ~x_3585;
assign n_23670 = ~x_3586 & ~x_3587;
assign n_23671 =  n_23669 &  n_23670;
assign n_23672 =  n_23668 &  n_23671;
assign n_23673 =  n_23665 &  n_23672;
assign n_23674 =  n_23658 &  n_23673;
assign n_23675 =  n_6182 &  n_23674;
assign n_23676 =  n_10872 &  n_23675;
assign n_23677 = ~n_23643 & ~n_23676;
assign n_23678 = ~x_4265 & ~n_23002;
assign n_23679 =  n_13872 &  n_23329;
assign n_23680 = ~n_23678 &  n_23679;
assign n_23681 =  n_7 &  n_23459;
assign n_23682 =  n_23252 &  n_23681;
assign n_23683 =  n_561 &  n_1896;
assign n_23684 =  n_1037 &  n_23683;
assign n_23685 =  n_23459 &  n_2485;
assign n_23686 =  n_23684 &  n_23685;
assign n_23687 =  n_21953 &  n_6181;
assign n_23688 =  n_10872 &  n_23687;
assign n_23689 = ~n_23686 & ~n_23688;
assign n_23690 = ~n_23682 &  n_23689;
assign n_23691 =  n_766 &  n_556;
assign n_23692 =  n_349 &  n_23691;
assign n_23693 =  n_23692 &  n_23613;
assign n_23694 =  n_758 &  n_3629;
assign n_23695 = ~x_2671 & ~x_2672;
assign n_23696 = ~x_2673 & ~x_2674;
assign n_23697 =  n_23695 &  n_23696;
assign n_23698 = ~x_2667 & ~x_2668;
assign n_23699 = ~x_2669 & ~x_2670;
assign n_23700 =  n_23698 &  n_23699;
assign n_23701 =  n_23697 &  n_23700;
assign n_23702 = ~x_2679 & ~x_2680;
assign n_23703 = ~x_2681 & ~x_2682;
assign n_23704 =  n_23702 &  n_23703;
assign n_23705 = ~x_2675 & ~x_2676;
assign n_23706 = ~x_2677 & ~x_2678;
assign n_23707 =  n_23705 &  n_23706;
assign n_23708 =  n_23704 &  n_23707;
assign n_23709 =  n_23701 &  n_23708;
assign n_23710 = ~x_2655 & ~x_2656;
assign n_23711 = ~x_2657 & ~x_2658;
assign n_23712 =  n_23710 &  n_23711;
assign n_23713 = ~x_2651 & ~x_2652;
assign n_23714 = ~x_2653 & ~x_2654;
assign n_23715 =  n_23713 &  n_23714;
assign n_23716 =  n_23712 &  n_23715;
assign n_23717 = ~x_2663 & ~x_2664;
assign n_23718 = ~x_2665 & ~x_2666;
assign n_23719 =  n_23717 &  n_23718;
assign n_23720 = ~x_2659 & ~x_2660;
assign n_23721 = ~x_2661 & ~x_2662;
assign n_23722 =  n_23720 &  n_23721;
assign n_23723 =  n_23719 &  n_23722;
assign n_23724 =  n_23716 &  n_23723;
assign n_23725 =  n_23709 &  n_23724;
assign n_23726 =  n_23694 & ~n_23725;
assign n_23727 = ~n_23693 & ~n_23726;
assign n_23728 =  n_23690 &  n_23727;
assign n_23729 = ~n_23680 &  n_23728;
assign n_23730 =  n_23677 &  n_23729;
assign n_23731 = ~n_23640 &  n_23730;
assign n_23732 =  n_555 &  n_5982;
assign n_23733 = ~x_4540 & ~x_4541;
assign n_23734 = ~x_4542 & ~x_4543;
assign n_23735 =  n_23733 &  n_23734;
assign n_23736 = ~x_4536 & ~x_4537;
assign n_23737 = ~x_4538 & ~x_4539;
assign n_23738 =  n_23736 &  n_23737;
assign n_23739 =  n_23735 &  n_23738;
assign n_23740 = ~x_4548 & ~x_4549;
assign n_23741 = ~x_4550 & ~x_4551;
assign n_23742 =  n_23740 &  n_23741;
assign n_23743 = ~x_4544 & ~x_4545;
assign n_23744 = ~x_4546 & ~x_4547;
assign n_23745 =  n_23743 &  n_23744;
assign n_23746 =  n_23742 &  n_23745;
assign n_23747 =  n_23739 &  n_23746;
assign n_23748 = ~x_4524 & ~x_4525;
assign n_23749 = ~x_4526 & ~x_4527;
assign n_23750 =  n_23748 &  n_23749;
assign n_23751 = ~x_4520 & ~x_4521;
assign n_23752 = ~x_4522 & ~x_4523;
assign n_23753 =  n_23751 &  n_23752;
assign n_23754 =  n_23750 &  n_23753;
assign n_23755 = ~x_4532 & ~x_4533;
assign n_23756 = ~x_4534 & ~x_4535;
assign n_23757 =  n_23755 &  n_23756;
assign n_23758 = ~x_4528 & ~x_4529;
assign n_23759 = ~x_4530 & ~x_4531;
assign n_23760 =  n_23758 &  n_23759;
assign n_23761 =  n_23757 &  n_23760;
assign n_23762 =  n_23754 &  n_23761;
assign n_23763 =  n_23747 &  n_23762;
assign n_23764 =  n_23732 &  n_23763;
assign n_23765 =  n_8359 &  n_21758;
assign n_23766 =  n_6181 &  n_9690;
assign n_23767 =  n_764 &  n_147;
assign n_23768 =  n_23766 &  n_23767;
assign n_23769 = ~n_23765 & ~n_23768;
assign n_23770 = ~n_23764 &  n_23769;
assign n_23771 =  n_7078 &  n_356;
assign n_23772 = ~x_2799 & ~x_2800;
assign n_23773 = ~x_2801 & ~x_2802;
assign n_23774 =  n_23772 &  n_23773;
assign n_23775 = ~x_2795 & ~x_2796;
assign n_23776 = ~x_2797 & ~x_2798;
assign n_23777 =  n_23775 &  n_23776;
assign n_23778 =  n_23774 &  n_23777;
assign n_23779 = ~x_2807 & ~x_2808;
assign n_23780 = ~x_2809 & ~x_2810;
assign n_23781 =  n_23779 &  n_23780;
assign n_23782 = ~x_2803 & ~x_2804;
assign n_23783 = ~x_2805 & ~x_2806;
assign n_23784 =  n_23782 &  n_23783;
assign n_23785 =  n_23781 &  n_23784;
assign n_23786 =  n_23778 &  n_23785;
assign n_23787 = ~x_2783 & ~x_2784;
assign n_23788 = ~x_2785 & ~x_2786;
assign n_23789 =  n_23787 &  n_23788;
assign n_23790 = ~x_2779 & ~x_2780;
assign n_23791 = ~x_2781 & ~x_2782;
assign n_23792 =  n_23790 &  n_23791;
assign n_23793 =  n_23789 &  n_23792;
assign n_23794 = ~x_2791 & ~x_2792;
assign n_23795 = ~x_2793 & ~x_2794;
assign n_23796 =  n_23794 &  n_23795;
assign n_23797 = ~x_2787 & ~x_2788;
assign n_23798 = ~x_2789 & ~x_2790;
assign n_23799 =  n_23797 &  n_23798;
assign n_23800 =  n_23796 &  n_23799;
assign n_23801 =  n_23793 &  n_23800;
assign n_23802 =  n_23786 &  n_23801;
assign n_23803 =  n_23771 & ~n_23802;
assign n_23804 =  n_351 &  n_3619;
assign n_23805 = ~n_23134 &  n_23804;
assign n_23806 = ~n_23803 & ~n_23805;
assign n_23807 =  n_23770 &  n_23806;
assign n_23808 =  n_10867 & ~n_23725;
assign n_23809 =  n_23329 &  n_23808;
assign n_23810 = ~n_13868 & ~n_13105;
assign n_23811 = ~n_14268 &  n_23810;
assign n_23812 =  n_9884 &  n_18914;
assign n_23813 =  n_5652 &  n_355;
assign n_23814 = ~n_23812 & ~n_23813;
assign n_23815 =  n_2290 &  n_12;
assign n_23816 =  n_1898 &  n_23459;
assign n_23817 =  n_5654 &  n_23816;
assign n_23818 =  n_23815 &  n_23817;
assign n_23819 = ~x_39 &  n_756;
assign n_23820 =  n_23819 &  n_23460;
assign n_23821 =  n_10872 &  n_23820;
assign n_23822 = ~n_23818 & ~n_23821;
assign n_23823 =  n_23814 &  n_23822;
assign n_23824 =  n_23811 &  n_23823;
assign n_23825 = ~n_23809 &  n_23824;
assign n_23826 =  n_23807 &  n_23825;
assign n_23827 =  n_5 &  n_23618;
assign n_23828 =  n_23827 &  n_23617;
assign n_23829 = ~x_38 &  n_8818;
assign n_23830 =  n_150 &  n_23829;
assign n_23831 = ~n_23828 & ~n_23830;
assign n_23832 = ~x_1707 & ~n_22968;
assign n_23833 = ~n_23828 &  n_23832;
assign n_23834 = ~n_23831 & ~n_23833;
assign n_23835 =  n_23826 & ~n_23834;
assign n_23836 =  n_23731 &  n_23835;
assign n_23837 =  n_23635 &  n_23836;
assign n_23838 =  n_23605 &  n_23837;
assign n_23839 =  n_2094 &  n_8360;
assign n_23840 =  x_38 &  n_23816;
assign n_23841 =  n_23840 &  n_8818;
assign n_23842 = ~n_23839 & ~n_23841;
assign n_23843 =  n_23009 &  n_1501;
assign n_23844 =  n_1896 &  n_23843;
assign n_23845 =  n_23844 &  n_8365;
assign n_23846 = ~n_20208 & ~n_23845;
assign n_23847 =  n_23842 &  n_23846;
assign n_23848 =  n_23381 &  n_768;
assign n_23849 =  n_13104 &  n_23848;
assign n_23850 = ~n_23849 & ~n_5650;
assign n_23851 =  n_2 &  n_20402;
assign n_23852 = ~n_18109 & ~n_23851;
assign n_23853 =  n_23850 &  n_23852;
assign n_23854 =  n_23847 &  n_23853;
assign n_23855 =  n_1037 &  n_4283;
assign n_23856 = ~x_43 &  n_16110;
assign n_23857 = ~n_23855 & ~n_23856;
assign n_23858 =  n_23857 & ~n_7662;
assign n_23859 =  n_23854 &  n_23858;
assign n_23860 = ~x_2379 & ~x_2380;
assign n_23861 = ~x_2381 & ~x_2382;
assign n_23862 = ~x_2383 & ~x_2384;
assign n_23863 =  n_23861 &  n_23862;
assign n_23864 =  n_23860 &  n_23863;
assign n_23865 = ~x_2389 & ~x_2390;
assign n_23866 = ~x_2391 & ~x_2392;
assign n_23867 =  n_23865 &  n_23866;
assign n_23868 = ~x_2385 & ~x_2386;
assign n_23869 = ~x_2387 & ~x_2388;
assign n_23870 =  n_23868 &  n_23869;
assign n_23871 =  n_23867 &  n_23870;
assign n_23872 =  n_23864 &  n_23871;
assign n_23873 = ~x_2393 &  n_23872;
assign n_23874 =  x_2394 &  n_23873;
assign n_23875 = ~x_43 &  x_2395;
assign n_23876 =  x_42 &  n_12;
assign n_23877 =  n_1896 &  n_552;
assign n_23878 =  n_23876 &  n_23877;
assign n_23879 =  n_23875 &  n_23878;
assign n_23880 =  n_23874 &  n_23879;
assign n_23881 =  n_23050 &  n_23459;
assign n_23882 =  n_8353 &  n_23881;
assign n_23883 =  n_2683 &  n_23459;
assign n_23884 =  n_151 &  n_23329;
assign n_23885 =  n_23883 &  n_23884;
assign n_23886 = ~n_23882 & ~n_23885;
assign n_23887 =  n_23460 &  n_23766;
assign n_23888 = ~x_36 & ~x_37;
assign n_23889 =  n_23459 &  n_23888;
assign n_23890 =  n_10478 &  n_23889;
assign n_23891 = ~n_23887 & ~n_23890;
assign n_23892 =  n_23886 &  n_23891;
assign n_23893 = ~n_23880 &  n_23892;
assign n_23894 =  n_5654 &  n_4283;
assign n_23895 =  n_4289 &  n_22940;
assign n_23896 = ~n_23894 & ~n_23895;
assign n_23897 =  n_23375 &  n_2486;
assign n_23898 =  n_13104 &  n_19493;
assign n_23899 = ~n_23897 & ~n_23898;
assign n_23900 =  n_8344 &  n_23820;
assign n_23901 =  n_8353 &  n_23840;
assign n_23902 = ~n_23900 & ~n_23901;
assign n_23903 =  n_23899 &  n_23902;
assign n_23904 =  n_23896 &  n_23903;
assign n_23905 =  n_23893 &  n_23904;
assign n_23906 =  n_23859 &  n_23905;
assign n_23907 =  n_3622 & ~n_18302;
assign n_23908 = ~x_3788 & ~x_3789;
assign n_23909 = ~x_3790 & ~x_3791;
assign n_23910 =  n_23908 &  n_23909;
assign n_23911 = ~x_3784 & ~x_3785;
assign n_23912 = ~x_3786 & ~x_3787;
assign n_23913 =  n_23911 &  n_23912;
assign n_23914 =  n_23910 &  n_23913;
assign n_23915 = ~x_3796 & ~x_3797;
assign n_23916 = ~x_3798 & ~x_3799;
assign n_23917 =  n_23915 &  n_23916;
assign n_23918 = ~x_3792 & ~x_3793;
assign n_23919 = ~x_3794 & ~x_3795;
assign n_23920 =  n_23918 &  n_23919;
assign n_23921 =  n_23917 &  n_23920;
assign n_23922 =  n_23914 &  n_23921;
assign n_23923 = ~x_3772 & ~x_3773;
assign n_23924 = ~x_3774 & ~x_3775;
assign n_23925 =  n_23923 &  n_23924;
assign n_23926 = ~x_3768 & ~x_3769;
assign n_23927 = ~x_3770 & ~x_3771;
assign n_23928 =  n_23926 &  n_23927;
assign n_23929 =  n_23925 &  n_23928;
assign n_23930 = ~x_3780 & ~x_3781;
assign n_23931 = ~x_3782 & ~x_3783;
assign n_23932 =  n_23930 &  n_23931;
assign n_23933 = ~x_3776 & ~x_3777;
assign n_23934 = ~x_3778 & ~x_3779;
assign n_23935 =  n_23933 &  n_23934;
assign n_23936 =  n_23932 &  n_23935;
assign n_23937 =  n_23929 &  n_23936;
assign n_23938 =  n_23922 &  n_23937;
assign n_23939 =  n_9690 &  n_357;
assign n_23940 =  n_23938 &  n_23939;
assign n_23941 =  n_6379 &  n_6877;
assign n_23942 =  n_21953 &  n_23819;
assign n_23943 =  n_10872 &  n_23942;
assign n_23944 = ~n_23941 & ~n_23943;
assign n_23945 =  n_2290 &  n_6379;
assign n_23946 =  n_555 &  n_23945;
assign n_23947 = ~n_23946 & ~n_21178;
assign n_23948 =  n_23944 &  n_23947;
assign n_23949 = ~n_23940 &  n_23948;
assign n_23950 =  n_23907 &  n_23949;
assign n_23951 =  n_23174 &  n_3346;
assign n_23952 = ~x_4508 & ~x_4509;
assign n_23953 = ~x_4510 & ~x_4511;
assign n_23954 =  n_23952 &  n_23953;
assign n_23955 = ~x_4504 & ~x_4505;
assign n_23956 = ~x_4506 & ~x_4507;
assign n_23957 =  n_23955 &  n_23956;
assign n_23958 =  n_23954 &  n_23957;
assign n_23959 = ~x_4516 & ~x_4517;
assign n_23960 = ~x_4518 & ~x_4519;
assign n_23961 =  n_23959 &  n_23960;
assign n_23962 = ~x_4512 & ~x_4513;
assign n_23963 = ~x_4514 & ~x_4515;
assign n_23964 =  n_23962 &  n_23963;
assign n_23965 =  n_23961 &  n_23964;
assign n_23966 =  n_23958 &  n_23965;
assign n_23967 = ~x_4492 & ~x_4493;
assign n_23968 = ~x_4494 & ~x_4495;
assign n_23969 =  n_23967 &  n_23968;
assign n_23970 = ~x_4488 & ~x_4489;
assign n_23971 = ~x_4490 & ~x_4491;
assign n_23972 =  n_23970 &  n_23971;
assign n_23973 =  n_23969 &  n_23972;
assign n_23974 = ~x_4500 & ~x_4501;
assign n_23975 = ~x_4502 & ~x_4503;
assign n_23976 =  n_23974 &  n_23975;
assign n_23977 = ~x_4496 & ~x_4497;
assign n_23978 = ~x_4498 & ~x_4499;
assign n_23979 =  n_23977 &  n_23978;
assign n_23980 =  n_23976 &  n_23979;
assign n_23981 =  n_23973 &  n_23980;
assign n_23982 =  n_23966 &  n_23981;
assign n_23983 =  n_23951 &  n_23982;
assign n_23984 =  n_10867 &  n_23725;
assign n_23985 =  n_23329 &  n_23984;
assign n_23986 = ~n_23983 & ~n_23985;
assign n_23987 =  n_21952 &  n_2485;
assign n_23988 =  n_10478 &  n_23987;
assign n_23989 =  x_41 &  n_1174;
assign n_23990 = ~x_38 &  n_23989;
assign n_23991 =  n_23990 &  n_23843;
assign n_23992 =  n_1037 &  n_23991;
assign n_23993 =  n_1037 &  n_23012;
assign n_23994 =  n_23843 &  n_23993;
assign n_23995 = ~n_23992 & ~n_23994;
assign n_23996 = ~n_23988 &  n_23995;
assign n_23997 =  n_154 &  n_1900;
assign n_23998 = ~n_3145 & ~n_23997;
assign n_23999 = ~n_5983 &  n_23998;
assign n_24000 =  n_23996 &  n_23999;
assign n_24001 =  n_23986 &  n_24000;
assign n_24002 =  n_23950 &  n_24001;
assign n_24003 =  n_23906 &  n_24002;
assign n_24004 =  n_23329 &  n_3619;
assign n_24005 =  n_154 &  n_3619;
assign n_24006 = ~n_24004 & ~n_24005;
assign n_24007 =  n_17783 &  n_2682;
assign n_24008 =  n_765 &  n_6181;
assign n_24009 =  n_6180 &  n_24008;
assign n_24010 =  x_43 &  n_24009;
assign n_24011 = ~n_24007 & ~n_24010;
assign n_24012 =  n_24006 &  n_24011;
assign n_24013 = ~x_3416 &  n_21952;
assign n_24014 =  n_2485 &  n_24013;
assign n_24015 =  n_2094 &  n_556;
assign n_24016 =  n_24014 &  n_24015;
assign n_24017 =  n_5 &  n_768;
assign n_24018 =  n_350 &  n_24017;
assign n_24019 =  x_42 &  n_24018;
assign n_24020 = ~n_24016 & ~n_24019;
assign n_24021 =  n_15366 &  n_3616;
assign n_24022 =  n_8344 &  n_3619;
assign n_24023 = ~n_24021 & ~n_24022;
assign n_24024 =  n_24020 &  n_24023;
assign n_24025 =  n_24012 &  n_24024;
assign n_24026 =  n_4289 &  n_6377;
assign n_24027 =  n_1037 &  n_24026;
assign n_24028 =  n_769 &  n_354;
assign n_24029 =  n_5654 &  n_24028;
assign n_24030 = ~n_24027 & ~n_24029;
assign n_24031 =  n_1037 &  n_8348;
assign n_24032 = ~n_21564 & ~n_6525;
assign n_24033 =  n_757 & ~n_24032;
assign n_24034 = ~n_24031 & ~n_24033;
assign n_24035 =  n_24030 &  n_24034;
assign n_24036 =  n_2094 &  n_3619;
assign n_24037 =  n_552 &  n_23683;
assign n_24038 =  x_42 &  n_24037;
assign n_24039 = ~n_24036 & ~n_24038;
assign n_24040 = ~x_3416 &  n_23381;
assign n_24041 =  n_24040 &  n_23465;
assign n_24042 =  n_349 &  n_24041;
assign n_24043 =  n_756 &  n_23381;
assign n_24044 =  n_1305 &  n_24043;
assign n_24045 =  n_152 &  n_24044;
assign n_24046 = ~n_24042 & ~n_24045;
assign n_24047 =  n_24039 &  n_24046;
assign n_24048 =  n_24035 &  n_24047;
assign n_24049 =  n_24025 &  n_24048;
assign n_24050 =  n_2290 &  n_2684;
assign n_24051 =  n_10872 &  n_24050;
assign n_24052 = ~n_20403 & ~n_24051;
assign n_24053 = ~n_4291 & ~n_21759;
assign n_24054 =  n_24052 &  n_24053;
assign n_24055 = ~x_38 &  n_23685;
assign n_24056 =  n_3625 &  n_24055;
assign n_24057 =  n_23005 &  n_23817;
assign n_24058 = ~n_24056 & ~n_24057;
assign n_24059 =  x_38 &  n_23889;
assign n_24060 =  n_5656 &  n_24059;
assign n_24061 = ~n_24060 & ~n_2488;
assign n_24062 =  n_24058 &  n_24061;
assign n_24063 =  n_24054 &  n_24062;
assign n_24064 =  n_24013 &  n_23888;
assign n_24065 =  n_23692 &  n_24064;
assign n_24066 = ~n_19496 & ~n_24065;
assign n_24067 =  x_3448 &  n_23816;
assign n_24068 =  n_20207 &  n_24067;
assign n_24069 =  n_2485 &  n_23051;
assign n_24070 =  n_16495 &  n_24069;
assign n_24071 = ~n_24068 & ~n_24070;
assign n_24072 =  n_24066 &  n_24071;
assign n_24073 =  n_5651 &  n_14;
assign n_24074 =  n_152 &  n_24073;
assign n_24075 = ~n_6380 & ~n_24074;
assign n_24076 = ~x_43 &  n_3633;
assign n_24077 =  n_21955 &  n_153;
assign n_24078 = ~n_24076 & ~n_24077;
assign n_24079 =  n_24075 &  n_24078;
assign n_24080 =  n_24072 &  n_24079;
assign n_24081 =  n_24063 &  n_24080;
assign n_24082 =  n_24049 &  n_24081;
assign n_24083 = ~x_2143 & ~x_2144;
assign n_24084 = ~x_2145 & ~x_2146;
assign n_24085 =  n_24083 &  n_24084;
assign n_24086 = ~x_2139 & ~x_2140;
assign n_24087 = ~x_2141 & ~x_2142;
assign n_24088 =  n_24086 &  n_24087;
assign n_24089 =  n_24085 &  n_24088;
assign n_24090 = ~x_2151 & ~x_2152;
assign n_24091 = ~x_2153 & ~x_2154;
assign n_24092 =  n_24090 &  n_24091;
assign n_24093 = ~x_2147 & ~x_2148;
assign n_24094 = ~x_2149 & ~x_2150;
assign n_24095 =  n_24093 &  n_24094;
assign n_24096 =  n_24092 &  n_24095;
assign n_24097 =  n_24089 &  n_24096;
assign n_24098 = ~x_2127 & ~x_2128;
assign n_24099 = ~x_2129 & ~x_2130;
assign n_24100 =  n_24098 &  n_24099;
assign n_24101 = ~x_2123 & ~x_2124;
assign n_24102 = ~x_2125 & ~x_2126;
assign n_24103 =  n_24101 &  n_24102;
assign n_24104 =  n_24100 &  n_24103;
assign n_24105 = ~x_2135 & ~x_2136;
assign n_24106 = ~x_2137 & ~x_2138;
assign n_24107 =  n_24105 &  n_24106;
assign n_24108 = ~x_2131 & ~x_2132;
assign n_24109 = ~x_2133 & ~x_2134;
assign n_24110 =  n_24108 &  n_24109;
assign n_24111 =  n_24107 &  n_24110;
assign n_24112 =  n_24104 &  n_24111;
assign n_24113 =  n_24097 &  n_24112;
assign n_24114 =  n_18914 &  n_24113;
assign n_24115 =  n_24114 &  n_8365;
assign n_24116 = ~x_40 &  n_1042;
assign n_24117 =  n_554 &  n_24116;
assign n_24118 = ~n_24115 & ~n_24117;
assign n_24119 =  n_1896 &  n_350;
assign n_24120 =  n_8359 &  n_24119;
assign n_24121 =  n_1037 &  n_24120;
assign n_24122 =  n_23548 &  n_2682;
assign n_24123 = ~n_24121 & ~n_24122;
assign n_24124 =  n_23884 &  n_23987;
assign n_24125 =  n_14263 &  n_1173;
assign n_24126 = ~n_24124 & ~n_24125;
assign n_24127 =  n_24123 &  n_24126;
assign n_24128 = ~x_4572 & ~x_4573;
assign n_24129 = ~x_4574 & ~x_4575;
assign n_24130 =  n_24128 &  n_24129;
assign n_24131 = ~x_4568 & ~x_4569;
assign n_24132 = ~x_4570 & ~x_4571;
assign n_24133 =  n_24131 &  n_24132;
assign n_24134 =  n_24130 &  n_24133;
assign n_24135 = ~x_4580 & ~x_4581;
assign n_24136 = ~x_4582 & ~x_4583;
assign n_24137 =  n_24135 &  n_24136;
assign n_24138 = ~x_4576 & ~x_4577;
assign n_24139 = ~x_4578 & ~x_4579;
assign n_24140 =  n_24138 &  n_24139;
assign n_24141 =  n_24137 &  n_24140;
assign n_24142 =  n_24134 &  n_24141;
assign n_24143 = ~x_4556 & ~x_4557;
assign n_24144 = ~x_4558 & ~x_4559;
assign n_24145 =  n_24143 &  n_24144;
assign n_24146 = ~x_4552 & ~x_4553;
assign n_24147 = ~x_4554 & ~x_4555;
assign n_24148 =  n_24146 &  n_24147;
assign n_24149 =  n_24145 &  n_24148;
assign n_24150 = ~x_4564 & ~x_4565;
assign n_24151 = ~x_4566 & ~x_4567;
assign n_24152 =  n_24150 &  n_24151;
assign n_24153 = ~x_4560 & ~x_4561;
assign n_24154 = ~x_4562 & ~x_4563;
assign n_24155 =  n_24153 &  n_24154;
assign n_24156 =  n_24152 &  n_24155;
assign n_24157 =  n_24149 &  n_24156;
assign n_24158 =  n_24142 &  n_24157;
assign n_24159 =  n_17782 &  n_10477;
assign n_24160 =  n_349 &  n_24159;
assign n_24161 = ~n_24158 &  n_24160;
assign n_24162 = ~x_1791 & ~x_1792;
assign n_24163 = ~x_1793 & ~x_1794;
assign n_24164 =  n_24162 &  n_24163;
assign n_24165 = ~x_1787 & ~x_1788;
assign n_24166 = ~x_1789 & ~x_1790;
assign n_24167 =  n_24165 &  n_24166;
assign n_24168 =  n_24164 &  n_24167;
assign n_24169 = ~x_1799 & ~x_1800;
assign n_24170 = ~x_1801 & ~x_1802;
assign n_24171 =  n_24169 &  n_24170;
assign n_24172 = ~x_1795 & ~x_1796;
assign n_24173 = ~x_1797 & ~x_1798;
assign n_24174 =  n_24172 &  n_24173;
assign n_24175 =  n_24171 &  n_24174;
assign n_24176 =  n_24168 &  n_24175;
assign n_24177 = ~x_1775 & ~x_1776;
assign n_24178 = ~x_1777 & ~x_1778;
assign n_24179 =  n_24177 &  n_24178;
assign n_24180 = ~x_1771 & ~x_1772;
assign n_24181 = ~x_1773 & ~x_1774;
assign n_24182 =  n_24180 &  n_24181;
assign n_24183 =  n_24179 &  n_24182;
assign n_24184 = ~x_1783 & ~x_1784;
assign n_24185 = ~x_1785 & ~x_1786;
assign n_24186 =  n_24184 &  n_24185;
assign n_24187 = ~x_1779 & ~x_1780;
assign n_24188 = ~x_1781 & ~x_1782;
assign n_24189 =  n_24187 &  n_24188;
assign n_24190 =  n_24186 &  n_24189;
assign n_24191 =  n_24183 &  n_24190;
assign n_24192 =  n_24176 &  n_24191;
assign n_24193 =  n_1305 &  n_767;
assign n_24194 =  n_17076 &  n_24193;
assign n_24195 =  n_24192 &  n_24194;
assign n_24196 = ~n_24161 & ~n_24195;
assign n_24197 =  n_24127 &  n_24196;
assign n_24198 =  n_24118 &  n_24197;
assign n_24199 =  n_554 &  n_5984;
assign n_24200 =  n_3141 &  n_5654;
assign n_24201 =  n_23465 &  n_24200;
assign n_24202 = ~n_13867 & ~n_24201;
assign n_24203 = ~n_24199 &  n_24202;
assign n_24204 =  n_5654 &  n_24018;
assign n_24205 =  n_6180 &  n_13230;
assign n_24206 =  n_8344 &  n_1900;
assign n_24207 = ~n_24205 & ~n_24206;
assign n_24208 = ~n_24204 &  n_24207;
assign n_24209 =  n_24203 &  n_24208;
assign n_24210 =  n_150 &  n_16495;
assign n_24211 =  x_1771 &  n_23384;
assign n_24212 =  n_11 &  n_24211;
assign n_24213 = ~n_24210 & ~n_24212;
assign n_24214 =  n_1 &  n_1043;
assign n_24215 =  n_24213 & ~n_24214;
assign n_24216 =  n_24209 &  n_24215;
assign n_24217 =  n_24198 &  n_24216;
assign n_24218 =  n_24082 &  n_24217;
assign n_24219 =  n_24003 &  n_24218;
assign n_24220 =  n_349 &  n_4283;
assign n_24221 =  n_6378 &  n_150;
assign n_24222 =  n_554 &  n_10078;
assign n_24223 =  n_1040 &  n_24222;
assign n_24224 = ~n_24221 & ~n_24223;
assign n_24225 = ~n_24220 &  n_24224;
assign n_24226 =  n_24043 &  n_13870;
assign n_24227 =  n_2094 &  n_19497;
assign n_24228 = ~n_24226 & ~n_24227;
assign n_24229 =  n_23388 &  n_15916;
assign n_24230 =  n_17782 &  n_22940;
assign n_24231 =  n_11 &  n_24120;
assign n_24232 = ~n_24230 & ~n_24231;
assign n_24233 = ~n_24229 &  n_24232;
assign n_24234 =  n_24228 &  n_24233;
assign n_24235 =  n_24225 &  n_24234;
assign n_24236 = ~x_3997 & ~x_3998;
assign n_24237 = ~x_3999 & ~x_4000;
assign n_24238 =  n_24236 &  n_24237;
assign n_24239 = ~x_3993 & ~x_3994;
assign n_24240 = ~x_3995 & ~x_3996;
assign n_24241 =  n_24239 &  n_24240;
assign n_24242 =  n_24238 &  n_24241;
assign n_24243 = ~x_4005 & ~x_4006;
assign n_24244 = ~x_4007 & ~x_4008;
assign n_24245 =  n_24243 &  n_24244;
assign n_24246 = ~x_4001 & ~x_4002;
assign n_24247 = ~x_4003 & ~x_4004;
assign n_24248 =  n_24246 &  n_24247;
assign n_24249 =  n_24245 &  n_24248;
assign n_24250 =  n_24242 &  n_24249;
assign n_24251 = ~x_3981 & ~x_3982;
assign n_24252 = ~x_3983 & ~x_3984;
assign n_24253 =  n_24251 &  n_24252;
assign n_24254 = ~x_3977 & ~x_3978;
assign n_24255 = ~x_3979 & ~x_3980;
assign n_24256 =  n_24254 &  n_24255;
assign n_24257 =  n_24253 &  n_24256;
assign n_24258 = ~x_3989 & ~x_3990;
assign n_24259 = ~x_3991 & ~x_3992;
assign n_24260 =  n_24258 &  n_24259;
assign n_24261 = ~x_3985 & ~x_3986;
assign n_24262 = ~x_3987 & ~x_3988;
assign n_24263 =  n_24261 &  n_24262;
assign n_24264 =  n_24260 &  n_24263;
assign n_24265 =  n_24257 &  n_24264;
assign n_24266 =  n_24250 &  n_24265;
assign n_24267 =  n_1899 &  n_23006;
assign n_24268 =  n_24266 &  n_24267;
assign n_24269 =  n_758 &  n_4288;
assign n_24270 =  n_6882 &  n_24269;
assign n_24271 = ~x_288 & ~x_289;
assign n_24272 = ~x_290 & ~x_291;
assign n_24273 =  n_24271 &  n_24272;
assign n_24274 = ~x_284 & ~x_285;
assign n_24275 = ~x_286 & ~x_287;
assign n_24276 =  n_24274 &  n_24275;
assign n_24277 =  n_24273 &  n_24276;
assign n_24278 = ~x_296 & ~x_297;
assign n_24279 = ~x_298 & ~x_299;
assign n_24280 =  n_24278 &  n_24279;
assign n_24281 = ~x_292 & ~x_293;
assign n_24282 = ~x_294 & ~x_295;
assign n_24283 =  n_24281 &  n_24282;
assign n_24284 =  n_24280 &  n_24283;
assign n_24285 =  n_24277 &  n_24284;
assign n_24286 = ~x_272 & ~x_273;
assign n_24287 = ~x_274 & ~x_275;
assign n_24288 =  n_24286 &  n_24287;
assign n_24289 = ~x_268 & ~x_269;
assign n_24290 = ~x_270 & ~x_271;
assign n_24291 =  n_24289 &  n_24290;
assign n_24292 =  n_24288 &  n_24291;
assign n_24293 = ~x_280 & ~x_281;
assign n_24294 = ~x_282 & ~x_283;
assign n_24295 =  n_24293 &  n_24294;
assign n_24296 = ~x_276 & ~x_277;
assign n_24297 = ~x_278 & ~x_279;
assign n_24298 =  n_24296 &  n_24297;
assign n_24299 =  n_24295 &  n_24298;
assign n_24300 =  n_24292 &  n_24299;
assign n_24301 =  n_24285 &  n_24300;
assign n_24302 =  n_24270 & ~n_24301;
assign n_24303 = ~n_24268 & ~n_24302;
assign n_24304 =  n_1899 &  n_23636;
assign n_24305 =  n_24303 & ~n_24304;
assign n_24306 =  n_7 &  n_23381;
assign n_24307 =  n_24306 &  n_3339;
assign n_24308 = ~n_24307 & ~n_1176;
assign n_24309 =  n_21952 &  n_23050;
assign n_24310 = ~x_39 &  n_10872;
assign n_24311 =  n_24309 &  n_24310;
assign n_24312 =  n_24308 & ~n_24311;
assign n_24313 =  n_20790 &  n_6379;
assign n_24314 =  n_22715 &  n_7;
assign n_24315 =  n_24314 &  n_8353;
assign n_24316 = ~n_24313 & ~n_24315;
assign n_24317 =  n_23596 &  n_10478;
assign n_24318 = ~x_38 &  n_23883;
assign n_24319 =  n_24310 &  n_24318;
assign n_24320 = ~n_24317 & ~n_24319;
assign n_24321 =  n_24316 &  n_24320;
assign n_24322 =  n_24312 &  n_24321;
assign n_24323 =  n_24305 &  n_24322;
assign n_24324 =  n_24235 &  n_24323;
assign n_24325 = ~x_3660 & ~x_3661;
assign n_24326 = ~x_3662 & ~x_3663;
assign n_24327 =  n_24325 &  n_24326;
assign n_24328 = ~x_3656 & ~x_3657;
assign n_24329 = ~x_3658 & ~x_3659;
assign n_24330 =  n_24328 &  n_24329;
assign n_24331 =  n_24327 &  n_24330;
assign n_24332 = ~x_3668 & ~x_3669;
assign n_24333 = ~x_3670 & ~x_3671;
assign n_24334 =  n_24332 &  n_24333;
assign n_24335 = ~x_3664 & ~x_3665;
assign n_24336 = ~x_3666 & ~x_3667;
assign n_24337 =  n_24335 &  n_24336;
assign n_24338 =  n_24334 &  n_24337;
assign n_24339 =  n_24331 &  n_24338;
assign n_24340 = ~x_3644 & ~x_3645;
assign n_24341 = ~x_3646 & ~x_3647;
assign n_24342 =  n_24340 &  n_24341;
assign n_24343 = ~x_3640 & ~x_3641;
assign n_24344 = ~x_3642 & ~x_3643;
assign n_24345 =  n_24343 &  n_24344;
assign n_24346 =  n_24342 &  n_24345;
assign n_24347 = ~x_3652 & ~x_3653;
assign n_24348 = ~x_3654 & ~x_3655;
assign n_24349 =  n_24347 &  n_24348;
assign n_24350 = ~x_3648 & ~x_3649;
assign n_24351 = ~x_3650 & ~x_3651;
assign n_24352 =  n_24350 &  n_24351;
assign n_24353 =  n_24349 &  n_24352;
assign n_24354 =  n_24346 &  n_24353;
assign n_24355 =  n_24339 &  n_24354;
assign n_24356 =  n_1305 &  n_4290;
assign n_24357 =  n_1038 &  n_24356;
assign n_24358 = ~n_24355 &  n_24357;
assign n_24359 =  n_5 &  n_23067;
assign n_24360 = ~x_1439 & ~x_1440;
assign n_24361 = ~x_1441 & ~x_1442;
assign n_24362 =  n_24360 &  n_24361;
assign n_24363 = ~x_1435 & ~x_1436;
assign n_24364 = ~x_1437 & ~x_1438;
assign n_24365 =  n_24363 &  n_24364;
assign n_24366 =  n_24362 &  n_24365;
assign n_24367 = ~x_1447 & ~x_1448;
assign n_24368 = ~x_1449 & ~x_1450;
assign n_24369 =  n_24367 &  n_24368;
assign n_24370 = ~x_1443 & ~x_1444;
assign n_24371 = ~x_1445 & ~x_1446;
assign n_24372 =  n_24370 &  n_24371;
assign n_24373 =  n_24369 &  n_24372;
assign n_24374 =  n_24366 &  n_24373;
assign n_24375 = ~x_1423 & ~x_1424;
assign n_24376 = ~x_1425 & ~x_1426;
assign n_24377 =  n_24375 &  n_24376;
assign n_24378 = ~x_1419 & ~x_1420;
assign n_24379 = ~x_1421 & ~x_1422;
assign n_24380 =  n_24378 &  n_24379;
assign n_24381 =  n_24377 &  n_24380;
assign n_24382 = ~x_1431 & ~x_1432;
assign n_24383 = ~x_1433 & ~x_1434;
assign n_24384 =  n_24382 &  n_24383;
assign n_24385 = ~x_1427 & ~x_1428;
assign n_24386 = ~x_1429 & ~x_1430;
assign n_24387 =  n_24385 &  n_24386;
assign n_24388 =  n_24384 &  n_24387;
assign n_24389 =  n_24381 &  n_24388;
assign n_24390 =  n_24374 &  n_24389;
assign n_24391 =  n_24359 & ~n_24390;
assign n_24392 = ~n_24358 & ~n_24391;
assign n_24393 = ~x_1215 & ~x_1216;
assign n_24394 = ~x_1217 & ~x_1218;
assign n_24395 =  n_24393 &  n_24394;
assign n_24396 = ~x_1211 & ~x_1212;
assign n_24397 = ~x_1213 & ~x_1214;
assign n_24398 =  n_24396 &  n_24397;
assign n_24399 =  n_24395 &  n_24398;
assign n_24400 = ~x_1223 & ~x_1224;
assign n_24401 = ~x_1225 & ~x_1226;
assign n_24402 =  n_24400 &  n_24401;
assign n_24403 = ~x_1219 & ~x_1220;
assign n_24404 = ~x_1221 & ~x_1222;
assign n_24405 =  n_24403 &  n_24404;
assign n_24406 =  n_24402 &  n_24405;
assign n_24407 =  n_24399 &  n_24406;
assign n_24408 = ~x_1199 & ~x_1200;
assign n_24409 = ~x_1201 & ~x_1202;
assign n_24410 =  n_24408 &  n_24409;
assign n_24411 = ~x_1195 & ~x_1196;
assign n_24412 = ~x_1197 & ~x_1198;
assign n_24413 =  n_24411 &  n_24412;
assign n_24414 =  n_24410 &  n_24413;
assign n_24415 = ~x_1207 & ~x_1208;
assign n_24416 = ~x_1209 & ~x_1210;
assign n_24417 =  n_24415 &  n_24416;
assign n_24418 = ~x_1203 & ~x_1204;
assign n_24419 = ~x_1205 & ~x_1206;
assign n_24420 =  n_24418 &  n_24419;
assign n_24421 =  n_24417 &  n_24420;
assign n_24422 =  n_24414 &  n_24421;
assign n_24423 =  n_24407 &  n_24422;
assign n_24424 =  n_13872 & ~n_24423;
assign n_24425 =  n_2094 &  n_24424;
assign n_24426 = ~x_2587 & ~n_23095;
assign n_24427 =  n_2095 &  n_6378;
assign n_24428 = ~n_24426 &  n_24427;
assign n_24429 = ~n_24425 & ~n_24428;
assign n_24430 =  n_24392 &  n_24429;
assign n_24431 =  n_1895 &  n_24017;
assign n_24432 = ~n_23630 &  n_24431;
assign n_24433 =  n_24430 & ~n_24432;
assign n_24434 =  n_24324 &  n_24433;
assign n_24435 =  n_14263 &  n_8053;
assign n_24436 = ~x_448 & ~x_449;
assign n_24437 = ~x_450 & ~x_451;
assign n_24438 =  n_24436 &  n_24437;
assign n_24439 = ~x_444 & ~x_445;
assign n_24440 = ~x_446 & ~x_447;
assign n_24441 =  n_24439 &  n_24440;
assign n_24442 =  n_24438 &  n_24441;
assign n_24443 = ~x_456 & ~x_457;
assign n_24444 = ~x_458 & ~x_459;
assign n_24445 =  n_24443 &  n_24444;
assign n_24446 = ~x_452 & ~x_453;
assign n_24447 = ~x_454 & ~x_455;
assign n_24448 =  n_24446 &  n_24447;
assign n_24449 =  n_24445 &  n_24448;
assign n_24450 =  n_24442 &  n_24449;
assign n_24451 = ~x_432 & ~x_433;
assign n_24452 = ~x_434 & ~x_435;
assign n_24453 =  n_24451 &  n_24452;
assign n_24454 = ~x_428 & ~x_429;
assign n_24455 = ~x_430 & ~x_431;
assign n_24456 =  n_24454 &  n_24455;
assign n_24457 =  n_24453 &  n_24456;
assign n_24458 = ~x_440 & ~x_441;
assign n_24459 = ~x_442 & ~x_443;
assign n_24460 =  n_24458 &  n_24459;
assign n_24461 = ~x_436 & ~x_437;
assign n_24462 = ~x_438 & ~x_439;
assign n_24463 =  n_24461 &  n_24462;
assign n_24464 =  n_24460 &  n_24463;
assign n_24465 =  n_24457 &  n_24464;
assign n_24466 =  n_24450 &  n_24465;
assign n_24467 =  n_24435 & ~n_24466;
assign n_24468 =  n_3339 &  n_8053;
assign n_24469 = ~x_2111 & ~x_2112;
assign n_24470 = ~x_2113 & ~x_2114;
assign n_24471 =  n_24469 &  n_24470;
assign n_24472 = ~x_2107 & ~x_2108;
assign n_24473 = ~x_2109 & ~x_2110;
assign n_24474 =  n_24472 &  n_24473;
assign n_24475 =  n_24471 &  n_24474;
assign n_24476 = ~x_2119 & ~x_2120;
assign n_24477 = ~x_2121 &  x_2122;
assign n_24478 =  n_24476 &  n_24477;
assign n_24479 = ~x_2115 & ~x_2116;
assign n_24480 = ~x_2117 & ~x_2118;
assign n_24481 =  n_24479 &  n_24480;
assign n_24482 =  n_24478 &  n_24481;
assign n_24483 =  n_24475 &  n_24482;
assign n_24484 = ~x_2095 & ~x_2096;
assign n_24485 = ~x_2097 & ~x_2098;
assign n_24486 =  n_24484 &  n_24485;
assign n_24487 = ~x_2091 & ~x_2092;
assign n_24488 = ~x_2093 & ~x_2094;
assign n_24489 =  n_24487 &  n_24488;
assign n_24490 =  n_24486 &  n_24489;
assign n_24491 = ~x_2103 & ~x_2104;
assign n_24492 = ~x_2105 & ~x_2106;
assign n_24493 =  n_24491 &  n_24492;
assign n_24494 = ~x_2099 & ~x_2100;
assign n_24495 = ~x_2101 & ~x_2102;
assign n_24496 =  n_24494 &  n_24495;
assign n_24497 =  n_24493 &  n_24496;
assign n_24498 =  n_24490 &  n_24497;
assign n_24499 =  n_24483 &  n_24498;
assign n_24500 =  n_24468 &  n_24499;
assign n_24501 = ~n_24467 & ~n_24500;
assign n_24502 =  x_38 &  n_2095;
assign n_24503 =  n_3623 &  n_24502;
assign n_24504 =  n_1042 &  n_8365;
assign n_24505 = ~n_24503 & ~n_24504;
assign n_24506 =  n_24501 &  n_24505;
assign n_24507 =  x_2393 &  n_23872;
assign n_24508 = ~x_43 & ~x_2395;
assign n_24509 =  x_2394 &  n_24508;
assign n_24510 =  n_4088 &  n_24509;
assign n_24511 =  n_8053 &  n_24510;
assign n_24512 =  n_24507 &  n_24511;
assign n_24513 =  n_153 &  n_3617;
assign n_24514 = ~n_24512 & ~n_24513;
assign n_24515 =  n_24013 &  n_23641;
assign n_24516 = ~x_43 &  n_24515;
assign n_24517 = ~x_42 &  n_24516;
assign n_24518 =  n_24514 & ~n_24517;
assign n_24519 =  n_24506 &  n_24518;
assign n_24520 =  n_23596 &  n_23684;
assign n_24521 =  n_23329 &  n_2096;
assign n_24522 = ~n_24520 & ~n_24521;
assign n_24523 =  n_1 &  n_12292;
assign n_24524 =  n_24522 & ~n_24523;
assign n_24525 =  n_9884 &  n_23808;
assign n_24526 =  n_24524 & ~n_24525;
assign n_24527 =  n_8344 &  n_23848;
assign n_24528 = ~n_24527 & ~n_14656;
assign n_24529 =  n_22940 &  n_23987;
assign n_24530 =  n_24318 &  n_3625;
assign n_24531 = ~n_24529 & ~n_24530;
assign n_24532 =  n_23329 &  n_24008;
assign n_24533 = ~x_608 & ~x_609;
assign n_24534 = ~x_610 & ~x_611;
assign n_24535 =  n_24533 &  n_24534;
assign n_24536 = ~x_604 & ~x_605;
assign n_24537 = ~x_606 & ~x_607;
assign n_24538 =  n_24536 &  n_24537;
assign n_24539 =  n_24535 &  n_24538;
assign n_24540 = ~x_616 & ~x_617;
assign n_24541 = ~x_618 & ~x_619;
assign n_24542 =  n_24540 &  n_24541;
assign n_24543 = ~x_612 & ~x_613;
assign n_24544 = ~x_614 & ~x_615;
assign n_24545 =  n_24543 &  n_24544;
assign n_24546 =  n_24542 &  n_24545;
assign n_24547 =  n_24539 &  n_24546;
assign n_24548 = ~x_592 & ~x_593;
assign n_24549 = ~x_594 & ~x_595;
assign n_24550 =  n_24548 &  n_24549;
assign n_24551 = ~x_588 & ~x_589;
assign n_24552 = ~x_590 & ~x_591;
assign n_24553 =  n_24551 &  n_24552;
assign n_24554 =  n_24550 &  n_24553;
assign n_24555 = ~x_600 & ~x_601;
assign n_24556 = ~x_602 & ~x_603;
assign n_24557 =  n_24555 &  n_24556;
assign n_24558 = ~x_596 & ~x_597;
assign n_24559 = ~x_598 & ~x_599;
assign n_24560 =  n_24558 &  n_24559;
assign n_24561 =  n_24557 &  n_24560;
assign n_24562 =  n_24554 &  n_24561;
assign n_24563 =  n_24547 &  n_24562;
assign n_24564 =  n_24532 & ~n_24563;
assign n_24565 =  n_24531 & ~n_24564;
assign n_24566 =  n_24528 &  n_24565;
assign n_24567 =  n_24526 &  n_24566;
assign n_24568 =  n_24519 &  n_24567;
assign n_24569 =  x_42 &  n_561;
assign n_24570 =  n_2290 &  n_14;
assign n_24571 =  n_24569 &  n_24570;
assign n_24572 =  x_43 &  n_24571;
assign n_24573 =  n_1038 &  n_762;
assign n_24574 = ~n_24572 & ~n_24573;
assign n_24575 =  n_21954 &  n_551;
assign n_24576 = ~n_6883 & ~n_24575;
assign n_24577 =  n_1 & ~n_24576;
assign n_24578 = ~n_6881 & ~n_24577;
assign n_24579 =  x_43 & ~n_24578;
assign n_24580 =  n_24574 & ~n_24579;
assign n_24581 =  n_10078 &  n_354;
assign n_24582 =  n_5645 &  n_24581;
assign n_24583 =  n_24582 & ~n_23556;
assign n_24584 = ~x_33 &  n_3;
assign n_24585 =  n_2683 &  n_1896;
assign n_24586 =  n_24584 &  n_24585;
assign n_24587 =  n_7467 &  n_24586;
assign n_24588 =  n_24587 & ~n_23832;
assign n_24589 = ~n_24583 & ~n_24588;
assign n_24590 =  n_24580 &  n_24589;
assign n_24591 =  n_3141 &  n_23594;
assign n_24592 =  n_23252 &  n_8354;
assign n_24593 = ~n_24591 & ~n_24592;
assign n_24594 = ~n_6527 &  n_24593;
assign n_24595 =  n_18624 &  n_1502;
assign n_24596 = ~x_2703 & ~x_2704;
assign n_24597 = ~x_2705 & ~x_2706;
assign n_24598 =  n_24596 &  n_24597;
assign n_24599 = ~x_2699 & ~x_2700;
assign n_24600 = ~x_2701 & ~x_2702;
assign n_24601 =  n_24599 &  n_24600;
assign n_24602 =  n_24598 &  n_24601;
assign n_24603 = ~x_2711 & ~x_2712;
assign n_24604 = ~x_2713 & ~x_2714;
assign n_24605 =  n_24603 &  n_24604;
assign n_24606 = ~x_2707 & ~x_2708;
assign n_24607 = ~x_2709 & ~x_2710;
assign n_24608 =  n_24606 &  n_24607;
assign n_24609 =  n_24605 &  n_24608;
assign n_24610 =  n_24602 &  n_24609;
assign n_24611 = ~x_2687 & ~x_2688;
assign n_24612 = ~x_2689 & ~x_2690;
assign n_24613 =  n_24611 &  n_24612;
assign n_24614 = ~x_2683 & ~x_2684;
assign n_24615 = ~x_2685 & ~x_2686;
assign n_24616 =  n_24614 &  n_24615;
assign n_24617 =  n_24613 &  n_24616;
assign n_24618 = ~x_2695 & ~x_2696;
assign n_24619 = ~x_2697 & ~x_2698;
assign n_24620 =  n_24618 &  n_24619;
assign n_24621 = ~x_2691 & ~x_2692;
assign n_24622 = ~x_2693 & ~x_2694;
assign n_24623 =  n_24621 &  n_24622;
assign n_24624 =  n_24620 &  n_24623;
assign n_24625 =  n_24617 &  n_24624;
assign n_24626 =  n_24610 &  n_24625;
assign n_24627 =  n_24595 &  n_24626;
assign n_24628 =  n_756 &  n_22715;
assign n_24629 =  n_23252 &  n_24628;
assign n_24630 =  n_554 &  n_5651;
assign n_24631 =  n_23843 &  n_24630;
assign n_24632 =  x_1771 &  n_24631;
assign n_24633 = ~n_24629 & ~n_24632;
assign n_24634 = ~n_24627 &  n_24633;
assign n_24635 =  n_24594 &  n_24634;
assign n_24636 = ~x_2767 & ~x_2768;
assign n_24637 = ~x_2769 & ~x_2770;
assign n_24638 =  n_24636 &  n_24637;
assign n_24639 = ~x_2763 & ~x_2764;
assign n_24640 = ~x_2765 & ~x_2766;
assign n_24641 =  n_24639 &  n_24640;
assign n_24642 =  n_24638 &  n_24641;
assign n_24643 = ~x_2775 & ~x_2776;
assign n_24644 = ~x_2777 & ~x_2778;
assign n_24645 =  n_24643 &  n_24644;
assign n_24646 = ~x_2771 & ~x_2772;
assign n_24647 = ~x_2773 & ~x_2774;
assign n_24648 =  n_24646 &  n_24647;
assign n_24649 =  n_24645 &  n_24648;
assign n_24650 =  n_24642 &  n_24649;
assign n_24651 = ~x_2751 & ~x_2752;
assign n_24652 = ~x_2753 & ~x_2754;
assign n_24653 =  n_24651 &  n_24652;
assign n_24654 = ~x_2747 & ~x_2748;
assign n_24655 = ~x_2749 & ~x_2750;
assign n_24656 =  n_24654 &  n_24655;
assign n_24657 =  n_24653 &  n_24656;
assign n_24658 = ~x_2759 & ~x_2760;
assign n_24659 = ~x_2761 & ~x_2762;
assign n_24660 =  n_24658 &  n_24659;
assign n_24661 = ~x_2755 & ~x_2756;
assign n_24662 = ~x_2757 & ~x_2758;
assign n_24663 =  n_24661 &  n_24662;
assign n_24664 =  n_24660 &  n_24663;
assign n_24665 =  n_24657 &  n_24664;
assign n_24666 =  n_24650 &  n_24665;
assign n_24667 =  n_8353 & ~n_24666;
assign n_24668 =  n_10276 &  n_24667;
assign n_24669 = ~x_43 &  n_24064;
assign n_24670 =  n_23815 &  n_24669;
assign n_24671 = ~x_42 &  n_24670;
assign n_24672 = ~n_24668 & ~n_24671;
assign n_24673 =  n_24635 &  n_24672;
assign n_24674 =  n_24590 &  n_24673;
assign n_24675 =  n_24568 &  n_24674;
assign n_24676 =  n_24434 &  n_24675;
assign n_24677 =  n_24219 &  n_24676;
assign n_24678 = ~x_4265 & ~n_23001;
assign n_24679 =  n_3141 &  n_24678;
assign n_24680 =  n_153 &  n_2880;
assign n_24681 =  n_24679 &  n_24680;
assign n_24682 =  n_24043 &  n_8054;
assign n_24683 = ~n_15919 & ~n_24682;
assign n_24684 =  n_151 &  n_23843;
assign n_24685 =  n_23329 &  n_24684;
assign n_24686 =  n_10478 &  n_23685;
assign n_24687 =  n_23993 &  n_23889;
assign n_24688 = ~n_24686 & ~n_24687;
assign n_24689 =  n_23816 &  n_23829;
assign n_24690 =  n_24688 & ~n_24689;
assign n_24691 = ~n_24685 &  n_24690;
assign n_24692 =  n_24683 &  n_24691;
assign n_24693 = ~n_24681 &  n_24692;
assign n_24694 =  n_3143 &  n_3346;
assign n_24695 = ~n_8819 & ~n_24694;
assign n_24696 =  n_13872 &  n_6180;
assign n_24697 =  n_24695 & ~n_24696;
assign n_24698 =  n_23057 &  n_23058;
assign n_24699 =  n_24697 & ~n_24698;
assign n_24700 =  n_24693 &  n_24699;
assign n_24701 =  n_22716 &  n_23174;
assign n_24702 = ~n_24701 & ~n_1044;
assign n_24703 =  n_24222 &  n_551;
assign n_24704 = ~x_2735 & ~x_2736;
assign n_24705 = ~x_2737 & ~x_2738;
assign n_24706 =  n_24704 &  n_24705;
assign n_24707 = ~x_2731 & ~x_2732;
assign n_24708 = ~x_2733 & ~x_2734;
assign n_24709 =  n_24707 &  n_24708;
assign n_24710 =  n_24706 &  n_24709;
assign n_24711 = ~x_2743 & ~x_2744;
assign n_24712 = ~x_2745 & ~x_2746;
assign n_24713 =  n_24711 &  n_24712;
assign n_24714 = ~x_2739 & ~x_2740;
assign n_24715 = ~x_2741 & ~x_2742;
assign n_24716 =  n_24714 &  n_24715;
assign n_24717 =  n_24713 &  n_24716;
assign n_24718 =  n_24710 &  n_24717;
assign n_24719 = ~x_2719 & ~x_2720;
assign n_24720 = ~x_2721 & ~x_2722;
assign n_24721 =  n_24719 &  n_24720;
assign n_24722 = ~x_2715 & ~x_2716;
assign n_24723 = ~x_2717 & ~x_2718;
assign n_24724 =  n_24722 &  n_24723;
assign n_24725 =  n_24721 &  n_24724;
assign n_24726 = ~x_2727 & ~x_2728;
assign n_24727 = ~x_2729 & ~x_2730;
assign n_24728 =  n_24726 &  n_24727;
assign n_24729 = ~x_2723 & ~x_2724;
assign n_24730 = ~x_2725 & ~x_2726;
assign n_24731 =  n_24729 &  n_24730;
assign n_24732 =  n_24728 &  n_24731;
assign n_24733 =  n_24725 &  n_24732;
assign n_24734 =  n_24718 &  n_24733;
assign n_24735 =  n_24703 &  n_24734;
assign n_24736 =  x_43 &  n_24575;
assign n_24737 = ~n_2881 & ~n_24736;
assign n_24738 = ~n_2 & ~n_24737;
assign n_24739 =  n_24119 &  n_23883;
assign n_24740 = ~x_43 & ~x_3416;
assign n_24741 =  n_24739 &  n_24740;
assign n_24742 = ~x_42 &  n_24741;
assign n_24743 = ~n_24738 & ~n_24742;
assign n_24744 = ~n_24735 &  n_24743;
assign n_24745 =  n_24702 &  n_24744;
assign n_24746 =  n_561 &  n_2290;
assign n_24747 = ~x_1771 &  n_21952;
assign n_24748 =  n_2683 &  n_24747;
assign n_24749 =  n_24746 &  n_24748;
assign n_24750 =  n_349 &  n_24749;
assign n_24751 =  n_24424 &  n_154;
assign n_24752 = ~n_24750 & ~n_24751;
assign n_24753 = ~x_37 &  n_14264;
assign n_24754 =  n_23827 &  n_24753;
assign n_24755 =  n_24752 & ~n_24754;
assign n_24756 =  n_24745 &  n_24755;
assign n_24757 =  n_24700 &  n_24756;
assign n_24758 =  n_1173 &  n_13870;
assign n_24759 =  x_39 &  n_24309;
assign n_24760 =  n_10872 &  n_24759;
assign n_24761 = ~n_24758 & ~n_24760;
assign n_24762 =  n_153 &  n_1307;
assign n_24763 =  n_1502 &  n_13672;
assign n_24764 =  n_1038 &  n_3629;
assign n_24765 = ~n_24763 & ~n_24764;
assign n_24766 = ~n_24762 &  n_24765;
assign n_24767 = ~n_6878 &  n_24766;
assign n_24768 =  n_24761 &  n_24767;
assign n_24769 = ~x_41 &  n_3628;
assign n_24770 =  n_1037 &  n_24769;
assign n_24771 = ~x_2315 & ~n_23322;
assign n_24772 =  n_354 &  n_24771;
assign n_24773 =  n_24770 &  n_24772;
assign n_24774 =  n_24768 & ~n_24773;
assign n_24775 =  n_556 &  n_6525;
assign n_24776 =  n_24775 &  n_1502;
assign n_24777 = ~n_23292 &  n_24776;
assign n_24778 =  n_2486 &  n_23178;
assign n_24779 =  n_23678 &  n_24778;
assign n_24780 = ~n_24777 & ~n_24779;
assign n_24781 =  n_24774 &  n_24780;
assign n_24782 =  n_23878 &  n_24508;
assign n_24783 =  n_23874 &  n_24782;
assign n_24784 =  n_10872 &  n_19493;
assign n_24785 = ~n_24783 & ~n_24784;
assign n_24786 =  n_13872 &  n_24423;
assign n_24787 =  n_154 &  n_24786;
assign n_24788 =  n_353 &  n_23010;
assign n_24789 = ~x_37 &  n_24788;
assign n_24790 =  n_13866 &  n_24789;
assign n_24791 = ~n_24787 & ~n_24790;
assign n_24792 =  n_24785 &  n_24791;
assign n_24793 = ~n_156 & ~n_16689;
assign n_24794 = ~n_4284 &  n_24793;
assign n_24795 = ~n_1895 & ~n_10872;
assign n_24796 =  n_6182 & ~n_24795;
assign n_24797 = ~n_23674 &  n_24796;
assign n_24798 = ~n_24797 & ~n_16111;
assign n_24799 =  n_24794 &  n_24798;
assign n_24800 =  n_3141 & ~n_24678;
assign n_24801 =  n_24680 &  n_24800;
assign n_24802 =  n_24799 & ~n_24801;
assign n_24803 =  n_24792 &  n_24802;
assign n_24804 =  n_24781 &  n_24803;
assign n_24805 =  n_24757 &  n_24804;
assign n_24806 =  n_4288 &  n_767;
assign n_24807 =  n_5656 &  n_24806;
assign n_24808 = ~x_3404 & ~x_3405;
assign n_24809 = ~x_3406 & ~x_3407;
assign n_24810 =  n_24808 &  n_24809;
assign n_24811 = ~x_3400 & ~x_3401;
assign n_24812 = ~x_3402 & ~x_3403;
assign n_24813 =  n_24811 &  n_24812;
assign n_24814 =  n_24810 &  n_24813;
assign n_24815 = ~x_3412 & ~x_3413;
assign n_24816 = ~x_3414 & ~x_3415;
assign n_24817 =  n_24815 &  n_24816;
assign n_24818 = ~x_3408 & ~x_3409;
assign n_24819 = ~x_3410 & ~x_3411;
assign n_24820 =  n_24818 &  n_24819;
assign n_24821 =  n_24817 &  n_24820;
assign n_24822 =  n_24814 &  n_24821;
assign n_24823 = ~x_3388 & ~x_3389;
assign n_24824 = ~x_3390 & ~x_3391;
assign n_24825 =  n_24823 &  n_24824;
assign n_24826 = ~x_3384 & ~x_3385;
assign n_24827 = ~x_3386 & ~x_3387;
assign n_24828 =  n_24826 &  n_24827;
assign n_24829 =  n_24825 &  n_24828;
assign n_24830 = ~x_3396 & ~x_3397;
assign n_24831 = ~x_3398 & ~x_3399;
assign n_24832 =  n_24830 &  n_24831;
assign n_24833 = ~x_3392 & ~x_3393;
assign n_24834 = ~x_3394 & ~x_3395;
assign n_24835 =  n_24833 &  n_24834;
assign n_24836 =  n_24832 &  n_24835;
assign n_24837 =  n_24829 &  n_24836;
assign n_24838 =  n_24822 &  n_24837;
assign n_24839 =  n_24807 & ~n_24838;
assign n_24840 =  n_5645 &  n_7273;
assign n_24841 = ~x_576 & ~x_577;
assign n_24842 = ~x_578 & ~x_579;
assign n_24843 =  n_24841 &  n_24842;
assign n_24844 = ~x_572 & ~x_573;
assign n_24845 = ~x_574 & ~x_575;
assign n_24846 =  n_24844 &  n_24845;
assign n_24847 =  n_24843 &  n_24846;
assign n_24848 = ~x_584 & ~x_585;
assign n_24849 = ~x_586 & ~x_587;
assign n_24850 =  n_24848 &  n_24849;
assign n_24851 = ~x_580 & ~x_581;
assign n_24852 = ~x_582 & ~x_583;
assign n_24853 =  n_24851 &  n_24852;
assign n_24854 =  n_24850 &  n_24853;
assign n_24855 =  n_24847 &  n_24854;
assign n_24856 = ~x_560 & ~x_561;
assign n_24857 = ~x_562 & ~x_563;
assign n_24858 =  n_24856 &  n_24857;
assign n_24859 = ~x_556 & ~x_557;
assign n_24860 = ~x_558 & ~x_559;
assign n_24861 =  n_24859 &  n_24860;
assign n_24862 =  n_24858 &  n_24861;
assign n_24863 = ~x_568 & ~x_569;
assign n_24864 = ~x_570 & ~x_571;
assign n_24865 =  n_24863 &  n_24864;
assign n_24866 = ~x_564 & ~x_565;
assign n_24867 = ~x_566 & ~x_567;
assign n_24868 =  n_24866 &  n_24867;
assign n_24869 =  n_24865 &  n_24868;
assign n_24870 =  n_24862 &  n_24869;
assign n_24871 =  n_24855 &  n_24870;
assign n_24872 =  n_24840 & ~n_24871;
assign n_24873 = ~n_24839 & ~n_24872;
assign n_24874 =  n_9884 &  n_19497;
assign n_24875 = ~n_9300 & ~n_24874;
assign n_24876 = ~x_3900 & ~x_3901;
assign n_24877 = ~x_3902 & ~x_3903;
assign n_24878 =  n_24876 &  n_24877;
assign n_24879 = ~x_3896 & ~x_3897;
assign n_24880 = ~x_3898 & ~x_3899;
assign n_24881 =  n_24879 &  n_24880;
assign n_24882 =  n_24878 &  n_24881;
assign n_24883 = ~x_3908 & ~x_3909;
assign n_24884 = ~x_3910 &  n_24883;
assign n_24885 = ~x_3904 & ~x_3905;
assign n_24886 = ~x_3906 & ~x_3907;
assign n_24887 =  n_24885 &  n_24886;
assign n_24888 =  n_24884 &  n_24887;
assign n_24889 =  n_24882 &  n_24888;
assign n_24890 = ~x_3911 &  x_3912;
assign n_24891 =  n_13104 &  n_24890;
assign n_24892 =  n_24889 &  n_24891;
assign n_24893 =  n_24570 &  n_24892;
assign n_24894 =  n_24875 & ~n_24893;
assign n_24895 =  n_24873 &  n_24894;
assign n_24896 = ~x_428 &  n_1039;
assign n_24897 = ~x_43 &  n_24896;
assign n_24898 =  n_353 &  n_24769;
assign n_24899 =  n_24897 &  n_24898;
assign n_24900 = ~x_42 &  n_24899;
assign n_24901 =  n_22940 &  n_552;
assign n_24902 = ~n_24901 & ~n_3634;
assign n_24903 =  n_4088 &  n_757;
assign n_24904 = ~n_24903 & ~n_18625;
assign n_24905 =  n_24902 &  n_24904;
assign n_24906 = ~n_24900 &  n_24905;
assign n_24907 =  n_23382 &  n_24775;
assign n_24908 = ~n_24907 & ~n_2292;
assign n_24909 =  n_561 &  n_23819;
assign n_24910 =  n_11 &  n_24909;
assign n_24911 =  n_24788 &  n_24910;
assign n_24912 =  n_24908 & ~n_24911;
assign n_24913 =  n_24906 &  n_24912;
assign n_24914 =  n_24895 &  n_24913;
assign n_24915 =  n_23382 &  n_20401;
assign n_24916 =  n_23174 &  n_24915;
assign n_24917 =  x_38 &  n_23252;
assign n_24918 =  n_22715 &  n_24917;
assign n_24919 = ~n_24916 & ~n_24918;
assign n_24920 =  n_24359 &  n_24390;
assign n_24921 =  n_24919 & ~n_24920;
assign n_24922 =  n_2291 &  n_17785;
assign n_24923 =  x_43 &  n_24922;
assign n_24924 =  n_23050 &  n_24013;
assign n_24925 =  n_3338 &  n_24924;
assign n_24926 =  n_349 &  n_24925;
assign n_24927 = ~n_24923 & ~n_24926;
assign n_24928 =  n_24921 &  n_24927;
assign n_24929 =  n_23816 &  n_23884;
assign n_24930 =  n_23843 &  n_5652;
assign n_24931 = ~n_24929 & ~n_24930;
assign n_24932 =  n_1895 &  n_19493;
assign n_24933 =  n_24684 &  n_6525;
assign n_24934 = ~n_24932 & ~n_24933;
assign n_24935 =  n_24931 &  n_24934;
assign n_24936 =  n_12 &  n_23942;
assign n_24937 =  n_1037 &  n_24936;
assign n_24938 =  n_22715 &  n_24909;
assign n_24939 =  n_1037 &  n_24938;
assign n_24940 =  n_23883 &  n_23554;
assign n_24941 = ~n_24939 & ~n_24940;
assign n_24942 = ~n_24937 &  n_24941;
assign n_24943 =  n_24935 &  n_24942;
assign n_24944 =  n_24928 &  n_24943;
assign n_24945 =  n_24914 &  n_24944;
assign n_24946 =  n_6379 &  n_23884;
assign n_24947 =  n_23942 &  n_23329;
assign n_24948 = ~n_24946 & ~n_24947;
assign n_24949 =  x_39 &  n_15366;
assign n_24950 =  n_23548 &  n_24949;
assign n_24951 =  n_24318 &  n_3623;
assign n_24952 = ~n_24950 & ~n_24951;
assign n_24953 =  n_24948 &  n_24952;
assign n_24954 =  n_6378 &  n_8359;
assign n_24955 =  x_1771 &  n_21952;
assign n_24956 =  n_2683 &  n_24955;
assign n_24957 =  n_24956 &  n_23006;
assign n_24958 = ~n_24954 & ~n_24957;
assign n_24959 =  n_2682 &  n_24628;
assign n_24960 =  n_24747 &  n_15917;
assign n_24961 =  n_24960 &  n_3143;
assign n_24962 = ~n_24959 & ~n_24961;
assign n_24963 =  n_24958 &  n_24962;
assign n_24964 =  n_24953 &  n_24963;
assign n_24965 =  n_6378 &  n_23596;
assign n_24966 = ~n_2097 & ~n_24965;
assign n_24967 =  n_758 &  n_5651;
assign n_24968 =  n_353 &  n_23612;
assign n_24969 =  x_37 &  n_24968;
assign n_24970 =  n_24967 &  n_24969;
assign n_24971 =  x_3384 &  n_23816;
assign n_24972 =  n_24971 &  n_13866;
assign n_24973 = ~n_24970 & ~n_24972;
assign n_24974 =  n_24966 &  n_24973;
assign n_24975 =  x_39 &  n_756;
assign n_24976 =  n_764 &  n_24975;
assign n_24977 =  n_23612 &  n_24976;
assign n_24978 =  n_351 &  n_24977;
assign n_24979 =  n_24306 &  n_4285;
assign n_24980 =  n_1037 &  n_24979;
assign n_24981 = ~n_24978 & ~n_24980;
assign n_24982 =  n_23596 &  n_23993;
assign n_24983 = ~n_24982 & ~n_18915;
assign n_24984 =  n_24981 &  n_24983;
assign n_24985 =  n_24974 &  n_24984;
assign n_24986 =  n_24964 &  n_24985;
assign n_24987 =  n_23816 &  n_13672;
assign n_24988 = ~n_24987 & ~n_3624;
assign n_24989 =  n_8344 &  n_24017;
assign n_24990 =  n_5654 &  n_23005;
assign n_24991 =  n_6379 &  n_24990;
assign n_24992 = ~n_24989 & ~n_24991;
assign n_24993 =  n_24988 &  n_24992;
assign n_24994 =  n_154 &  n_10867;
assign n_24995 = ~n_24994 & ~n_3630;
assign n_24996 =  n_1038 &  n_6883;
assign n_24997 = ~n_24996 & ~n_16302;
assign n_24998 =  n_24995 &  n_24997;
assign n_24999 =  n_24993 &  n_24998;
assign n_25000 =  n_20790 &  n_552;
assign n_25001 = ~n_25000 & ~n_10277;
assign n_25002 = ~x_42 &  n_2681;
assign n_25003 =  n_10276 &  n_25002;
assign n_25004 =  n_153 &  n_7273;
assign n_25005 = ~n_25003 & ~n_25004;
assign n_25006 =  n_25001 &  n_25005;
assign n_25007 =  n_14 &  n_13672;
assign n_25008 =  n_23006 &  n_3615;
assign n_25009 = ~n_25007 & ~n_25008;
assign n_25010 =  n_23382 &  n_24990;
assign n_25011 =  n_23548 &  n_21564;
assign n_25012 = ~n_25010 & ~n_25011;
assign n_25013 =  n_25009 &  n_25012;
assign n_25014 =  n_25006 &  n_25013;
assign n_25015 =  n_24999 &  n_25014;
assign n_25016 =  n_24748 &  n_23636;
assign n_25017 =  n_10478 &  n_552;
assign n_25018 =  n_24569 &  n_23607;
assign n_25019 = ~n_25017 & ~n_25018;
assign n_25020 = ~n_25016 &  n_25019;
assign n_25021 =  n_13104 &  n_24759;
assign n_25022 = ~n_25021 & ~n_1901;
assign n_25023 =  n_25020 &  n_25022;
assign n_25024 =  n_4289 &  n_6378;
assign n_25025 =  n_7467 &  n_10867;
assign n_25026 = ~n_25024 & ~n_25025;
assign n_25027 =  n_554 &  n_9;
assign n_25028 =  n_23174 &  n_6883;
assign n_25029 = ~n_25027 & ~n_25028;
assign n_25030 =  n_25026 &  n_25029;
assign n_25031 =  n_153 &  n_15916;
assign n_25032 =  n_765 &  n_25031;
assign n_25033 =  n_150 &  n_23993;
assign n_25034 = ~n_25032 & ~n_25033;
assign n_25035 =  n_23848 &  n_9690;
assign n_25036 =  n_24309 &  n_3623;
assign n_25037 = ~n_25035 & ~n_25036;
assign n_25038 =  n_25034 &  n_25037;
assign n_25039 =  n_25030 &  n_25038;
assign n_25040 =  n_25023 &  n_25039;
assign n_25041 =  n_25015 &  n_25040;
assign n_25042 =  n_24986 &  n_25041;
assign n_25043 =  n_24945 &  n_25042;
assign n_25044 =  n_8359 &  n_1896;
assign n_25045 =  n_5981 &  n_25044;
assign n_25046 =  x_43 &  n_25045;
assign n_25047 =  n_3615 &  n_24990;
assign n_25048 = ~x_1407 & ~x_1408;
assign n_25049 = ~x_1409 & ~x_1410;
assign n_25050 =  n_25048 &  n_25049;
assign n_25051 = ~x_1403 & ~x_1404;
assign n_25052 = ~x_1405 & ~x_1406;
assign n_25053 =  n_25051 &  n_25052;
assign n_25054 =  n_25050 &  n_25053;
assign n_25055 = ~x_1415 & ~x_1416;
assign n_25056 = ~x_1417 & ~x_1418;
assign n_25057 =  n_25055 &  n_25056;
assign n_25058 = ~x_1411 & ~x_1412;
assign n_25059 = ~x_1413 & ~x_1414;
assign n_25060 =  n_25058 &  n_25059;
assign n_25061 =  n_25057 &  n_25060;
assign n_25062 =  n_25054 &  n_25061;
assign n_25063 = ~x_1391 & ~x_1392;
assign n_25064 = ~x_1393 & ~x_1394;
assign n_25065 =  n_25063 &  n_25064;
assign n_25066 = ~x_1387 & ~x_1388;
assign n_25067 = ~x_1389 & ~x_1390;
assign n_25068 =  n_25066 &  n_25067;
assign n_25069 =  n_25065 &  n_25068;
assign n_25070 = ~x_1399 & ~x_1400;
assign n_25071 = ~x_1401 & ~x_1402;
assign n_25072 =  n_25070 &  n_25071;
assign n_25073 = ~x_1395 & ~x_1396;
assign n_25074 = ~x_1397 & ~x_1398;
assign n_25075 =  n_25073 &  n_25074;
assign n_25076 =  n_25072 &  n_25075;
assign n_25077 =  n_25069 &  n_25076;
assign n_25078 =  n_25062 &  n_25077;
assign n_25079 =  n_25047 &  n_25078;
assign n_25080 = ~n_25046 & ~n_25079;
assign n_25081 =  n_4290 &  n_4285;
assign n_25082 =  n_1037 &  n_25081;
assign n_25083 =  n_18624 &  n_2684;
assign n_25084 =  n_154 &  n_23942;
assign n_25085 = ~n_25083 & ~n_25084;
assign n_25086 = ~n_25082 &  n_25085;
assign n_25087 =  n_25080 &  n_25086;
assign n_25088 =  n_8361 &  n_23877;
assign n_25089 =  n_351 &  n_20596;
assign n_25090 = ~n_25088 & ~n_25089;
assign n_25091 =  x_41 &  n_8;
assign n_25092 = ~x_43 &  n_24040;
assign n_25093 =  n_25091 &  n_25092;
assign n_25094 = ~x_42 &  n_25093;
assign n_25095 =  n_25090 & ~n_25094;
assign n_25096 =  n_1037 &  n_4285;
assign n_25097 =  n_24043 &  n_25096;
assign n_25098 =  n_1037 &  n_23384;
assign n_25099 = ~n_25097 & ~n_25098;
assign n_25100 =  n_6378 &  n_23889;
assign n_25101 = ~n_25100 & ~n_9691;
assign n_25102 =  n_25099 &  n_25101;
assign n_25103 =  n_25095 &  n_25102;
assign n_25104 =  n_25087 &  n_25103;
assign n_25105 =  n_24909 &  n_23461;
assign n_25106 = ~x_3416 &  n_25105;
assign n_25107 =  n_768 &  n_23460;
assign n_25108 = ~x_1771 &  n_25107;
assign n_25109 = ~n_1895 & ~n_8361;
assign n_25110 =  n_25108 & ~n_25109;
assign n_25111 = ~n_25106 & ~n_25110;
assign n_25112 = ~n_1305 & ~n_23989;
assign n_25113 =  n_1037 & ~n_25112;
assign n_25114 = ~n_6876 & ~n_25113;
assign n_25115 =  n_757 & ~n_25114;
assign n_25116 =  n_350 &  n_24050;
assign n_25117 =  x_43 &  n_25116;
assign n_25118 = ~n_25115 & ~n_25117;
assign n_25119 =  n_25111 &  n_25118;
assign n_25120 = ~x_2271 & ~x_2272;
assign n_25121 = ~x_2273 & ~x_2274;
assign n_25122 =  n_25120 &  n_25121;
assign n_25123 = ~x_2267 & ~x_2268;
assign n_25124 = ~x_2269 & ~x_2270;
assign n_25125 =  n_25123 &  n_25124;
assign n_25126 =  n_25122 &  n_25125;
assign n_25127 = ~x_2279 & ~x_2280;
assign n_25128 = ~x_2281 & ~x_2282;
assign n_25129 =  n_25127 &  n_25128;
assign n_25130 = ~x_2275 & ~x_2276;
assign n_25131 = ~x_2277 & ~x_2278;
assign n_25132 =  n_25130 &  n_25131;
assign n_25133 =  n_25129 &  n_25132;
assign n_25134 =  n_25126 &  n_25133;
assign n_25135 = ~x_2255 & ~x_2256;
assign n_25136 = ~x_2257 & ~x_2258;
assign n_25137 =  n_25135 &  n_25136;
assign n_25138 = ~x_2251 & ~x_2252;
assign n_25139 = ~x_2253 & ~x_2254;
assign n_25140 =  n_25138 &  n_25139;
assign n_25141 =  n_25137 &  n_25140;
assign n_25142 = ~x_2263 & ~x_2264;
assign n_25143 = ~x_2265 & ~x_2266;
assign n_25144 =  n_25142 &  n_25143;
assign n_25145 = ~x_2259 & ~x_2260;
assign n_25146 = ~x_2261 & ~x_2262;
assign n_25147 =  n_25145 &  n_25146;
assign n_25148 =  n_25144 &  n_25147;
assign n_25149 =  n_25141 &  n_25148;
assign n_25150 =  n_25134 &  n_25149;
assign n_25151 =  n_15366 &  n_23607;
assign n_25152 = ~n_25150 &  n_25151;
assign n_25153 =  n_1174 &  n_757;
assign n_25154 =  n_23174 &  n_25153;
assign n_25155 = ~n_7274 & ~n_25154;
assign n_25156 = ~n_25152 &  n_25155;
assign n_25157 =  n_2094 &  n_24684;
assign n_25158 = ~x_1771 &  n_25157;
assign n_25159 = ~x_37 &  n_24968;
assign n_25160 =  n_349 &  n_25159;
assign n_25161 =  n_23374 &  n_25160;
assign n_25162 = ~n_25158 & ~n_25161;
assign n_25163 =  n_25156 &  n_25162;
assign n_25164 =  n_25119 &  n_25163;
assign n_25165 =  n_25104 &  n_25164;
assign n_25166 =  n_7079 &  n_23135;
assign n_25167 =  n_23174 &  n_20077;
assign n_25168 = ~n_25166 & ~n_25167;
assign n_25169 =  n_5654 &  n_8348;
assign n_25170 =  n_8361 &  n_24017;
assign n_25171 = ~n_25169 & ~n_25170;
assign n_25172 =  n_25168 &  n_25171;
assign n_25173 =  n_23460 &  n_24770;
assign n_25174 = ~n_17077 & ~n_25173;
assign n_25175 =  n_10872 &  n_6526;
assign n_25176 = ~x_1183 & ~x_1184;
assign n_25177 = ~x_1185 & ~x_1186;
assign n_25178 =  n_25176 &  n_25177;
assign n_25179 = ~x_1179 & ~x_1180;
assign n_25180 = ~x_1181 & ~x_1182;
assign n_25181 =  n_25179 &  n_25180;
assign n_25182 =  n_25178 &  n_25181;
assign n_25183 = ~x_1191 & ~x_1192;
assign n_25184 = ~x_1193 & ~x_1194;
assign n_25185 =  n_25183 &  n_25184;
assign n_25186 = ~x_1187 & ~x_1188;
assign n_25187 = ~x_1189 & ~x_1190;
assign n_25188 =  n_25186 &  n_25187;
assign n_25189 =  n_25185 &  n_25188;
assign n_25190 =  n_25182 &  n_25189;
assign n_25191 = ~x_1167 & ~x_1168;
assign n_25192 = ~x_1169 & ~x_1170;
assign n_25193 =  n_25191 &  n_25192;
assign n_25194 = ~x_1163 & ~x_1164;
assign n_25195 = ~x_1165 & ~x_1166;
assign n_25196 =  n_25194 &  n_25195;
assign n_25197 =  n_25193 &  n_25196;
assign n_25198 = ~x_1175 & ~x_1176;
assign n_25199 = ~x_1177 & ~x_1178;
assign n_25200 =  n_25198 &  n_25199;
assign n_25201 = ~x_1171 & ~x_1172;
assign n_25202 = ~x_1173 & ~x_1174;
assign n_25203 =  n_25201 &  n_25202;
assign n_25204 =  n_25200 &  n_25203;
assign n_25205 =  n_25197 &  n_25204;
assign n_25206 =  n_25190 &  n_25205;
assign n_25207 =  n_25175 &  n_25206;
assign n_25208 =  n_25174 & ~n_25207;
assign n_25209 =  n_25172 &  n_25208;
assign n_25210 =  n_1895 &  n_1042;
assign n_25211 = ~n_25150 &  n_25210;
assign n_25212 = ~x_3416 &  n_23843;
assign n_25213 =  n_23614 &  n_25212;
assign n_25214 = ~x_42 &  n_25213;
assign n_25215 = ~n_25211 & ~n_25214;
assign n_25216 =  x_43 &  n_3343;
assign n_25217 = ~x_428 &  n_561;
assign n_25218 =  n_23844 &  n_25217;
assign n_25219 =  n_349 &  n_25218;
assign n_25220 = ~n_25216 & ~n_25219;
assign n_25221 =  n_25215 &  n_25220;
assign n_25222 =  n_25209 &  n_25221;
assign n_25223 =  x_428 &  n_1039;
assign n_25224 =  n_25223 &  n_24898;
assign n_25225 =  n_11 &  n_25224;
assign n_25226 =  n_10872 &  n_23844;
assign n_25227 =  n_21955 &  n_23174;
assign n_25228 = ~n_25226 & ~n_25227;
assign n_25229 = ~n_25225 &  n_25228;
assign n_25230 =  n_6525 &  n_10470;
assign n_25231 =  n_17785 &  n_10867;
assign n_25232 =  x_43 &  n_25231;
assign n_25233 = ~n_25230 & ~n_25232;
assign n_25234 =  n_25233 & ~n_9429;
assign n_25235 =  n_25229 &  n_25234;
assign n_25236 =  n_4088 &  n_15;
assign n_25237 =  n_10078 &  n_3632;
assign n_25238 = ~n_25236 & ~n_25237;
assign n_25239 =  n_22940 &  n_2486;
assign n_25240 =  n_25239 &  n_25206;
assign n_25241 =  n_25238 & ~n_25240;
assign n_25242 = ~x_41 &  n_21954;
assign n_25243 =  x_1547 &  n_11;
assign n_25244 =  n_23460 &  n_25243;
assign n_25245 =  n_25242 &  n_25244;
assign n_25246 =  x_1547 &  n_23987;
assign n_25247 =  n_24630 &  n_25246;
assign n_25248 = ~n_25245 & ~n_25247;
assign n_25249 =  n_760 &  n_24502;
assign n_25250 =  n_6377 &  n_23987;
assign n_25251 =  n_1037 &  n_25250;
assign n_25252 = ~n_25249 & ~n_25251;
assign n_25253 =  n_25248 &  n_25252;
assign n_25254 =  n_25241 &  n_25253;
assign n_25255 =  n_25235 &  n_25254;
assign n_25256 =  n_25222 &  n_25255;
assign n_25257 =  n_25165 &  n_25256;
assign n_25258 =  n_25043 &  n_25257;
assign n_25259 =  n_24805 &  n_25258;
assign n_25260 =  n_24677 &  n_25259;
assign n_25261 =  n_1502 &  n_24626;
assign n_25262 =  n_5652 &  n_25261;
assign n_25263 =  n_1502 &  n_23638;
assign n_25264 =  n_23636 &  n_25263;
assign n_25265 = ~n_25262 & ~n_25264;
assign n_25266 = ~x_3913 & ~n_23628;
assign n_25267 =  n_6379 &  n_25266;
assign n_25268 =  n_24630 &  n_25267;
assign n_25269 =  n_23047 &  n_23048;
assign n_25270 = ~n_25268 & ~n_25269;
assign n_25271 =  n_1042 &  n_15366;
assign n_25272 = ~x_2618 &  n_23609;
assign n_25273 = ~x_2587 & ~n_25272;
assign n_25274 =  n_25271 &  n_25273;
assign n_25275 =  x_42 &  x_3416;
assign n_25276 = ~x_43 &  n_23991;
assign n_25277 =  n_25275 &  n_25276;
assign n_25278 =  x_428 &  n_23683;
assign n_25279 =  n_23843 &  n_25278;
assign n_25280 =  n_11 &  n_25279;
assign n_25281 =  n_6525 &  n_23844;
assign n_25282 = ~n_25280 & ~n_25281;
assign n_25283 = ~n_25277 &  n_25282;
assign n_25284 = ~n_25274 &  n_25283;
assign n_25285 =  n_25270 &  n_25284;
assign n_25286 =  n_25265 &  n_25285;
assign n_25287 =  x_1771 &  n_25107;
assign n_25288 =  n_7467 &  n_25287;
assign n_25289 =  n_3143 &  n_3342;
assign n_25290 = ~n_24426 &  n_25289;
assign n_25291 = ~n_25288 & ~n_25290;
assign n_25292 =  n_2 &  n_24581;
assign n_25293 =  n_2682 &  n_356;
assign n_25294 = ~n_24771 &  n_25293;
assign n_25295 = ~n_25292 & ~n_25294;
assign n_25296 =  n_7078 &  n_1503;
assign n_25297 = ~x_2416 & ~x_2417;
assign n_25298 = ~x_2418 & ~x_2419;
assign n_25299 =  n_25297 &  n_25298;
assign n_25300 = ~x_2412 & ~x_2413;
assign n_25301 = ~x_2414 & ~x_2415;
assign n_25302 =  n_25300 &  n_25301;
assign n_25303 =  n_25299 &  n_25302;
assign n_25304 = ~x_2424 & ~x_2425;
assign n_25305 = ~x_2426 & ~x_2427;
assign n_25306 =  n_25304 &  n_25305;
assign n_25307 = ~x_2420 & ~x_2421;
assign n_25308 = ~x_2422 & ~x_2423;
assign n_25309 =  n_25307 &  n_25308;
assign n_25310 =  n_25306 &  n_25309;
assign n_25311 =  n_25303 &  n_25310;
assign n_25312 = ~x_2400 & ~x_2401;
assign n_25313 = ~x_2402 & ~x_2403;
assign n_25314 =  n_25312 &  n_25313;
assign n_25315 = ~x_2396 & ~x_2397;
assign n_25316 = ~x_2398 & ~x_2399;
assign n_25317 =  n_25315 &  n_25316;
assign n_25318 =  n_25314 &  n_25317;
assign n_25319 = ~x_2408 & ~x_2409;
assign n_25320 = ~x_2410 & ~x_2411;
assign n_25321 =  n_25319 &  n_25320;
assign n_25322 = ~x_2404 & ~x_2405;
assign n_25323 = ~x_2406 & ~x_2407;
assign n_25324 =  n_25322 &  n_25323;
assign n_25325 =  n_25321 &  n_25324;
assign n_25326 =  n_25318 &  n_25325;
assign n_25327 =  n_25311 &  n_25326;
assign n_25328 =  n_25296 & ~n_25327;
assign n_25329 =  x_3416 &  n_12;
assign n_25330 =  n_23844 &  n_25329;
assign n_25331 =  n_11 &  n_25330;
assign n_25332 =  n_23691 &  n_25160;
assign n_25333 = ~n_25331 & ~n_25332;
assign n_25334 = ~n_25328 &  n_25333;
assign n_25335 =  n_25295 &  n_25334;
assign n_25336 =  n_25291 &  n_25335;
assign n_25337 =  n_24355 &  n_24357;
assign n_25338 =  n_24158 &  n_24160;
assign n_25339 =  n_153 &  n_24915;
assign n_25340 = ~n_25338 & ~n_25339;
assign n_25341 = ~n_25337 &  n_25340;
assign n_25342 = ~x_4137 &  n_23381;
assign n_25343 =  n_769 &  n_25342;
assign n_25344 =  n_349 &  n_25343;
assign n_25345 =  n_11 &  n_24979;
assign n_25346 =  x_1771 &  n_25345;
assign n_25347 = ~n_25344 & ~n_25346;
assign n_25348 =  n_10872 &  n_13230;
assign n_25349 = ~x_1343 & ~x_1344;
assign n_25350 = ~x_1345 & ~x_1346;
assign n_25351 =  n_25349 &  n_25350;
assign n_25352 = ~x_1339 & ~x_1340;
assign n_25353 = ~x_1341 & ~x_1342;
assign n_25354 =  n_25352 &  n_25353;
assign n_25355 =  n_25351 &  n_25354;
assign n_25356 = ~x_1351 & ~x_1352;
assign n_25357 = ~x_1353 & ~x_1354;
assign n_25358 =  n_25356 &  n_25357;
assign n_25359 = ~x_1347 & ~x_1348;
assign n_25360 = ~x_1349 & ~x_1350;
assign n_25361 =  n_25359 &  n_25360;
assign n_25362 =  n_25358 &  n_25361;
assign n_25363 =  n_25355 &  n_25362;
assign n_25364 = ~x_1327 & ~x_1328;
assign n_25365 = ~x_1329 & ~x_1330;
assign n_25366 =  n_25364 &  n_25365;
assign n_25367 = ~x_1323 & ~x_1324;
assign n_25368 = ~x_1325 & ~x_1326;
assign n_25369 =  n_25367 &  n_25368;
assign n_25370 =  n_25366 &  n_25369;
assign n_25371 = ~x_1335 & ~x_1336;
assign n_25372 = ~x_1337 & ~x_1338;
assign n_25373 =  n_25371 &  n_25372;
assign n_25374 = ~x_1331 & ~x_1332;
assign n_25375 = ~x_1333 & ~x_1334;
assign n_25376 =  n_25374 &  n_25375;
assign n_25377 =  n_25373 &  n_25376;
assign n_25378 =  n_25370 &  n_25377;
assign n_25379 =  n_25363 &  n_25378;
assign n_25380 =  n_25348 & ~n_25379;
assign n_25381 = ~x_43 &  n_24909;
assign n_25382 =  n_24968 &  n_25381;
assign n_25383 = ~x_42 &  n_25382;
assign n_25384 = ~n_25380 & ~n_25383;
assign n_25385 =  n_25347 &  n_25384;
assign n_25386 =  n_25341 &  n_25385;
assign n_25387 =  n_8361 &  n_23945;
assign n_25388 = ~x_160 & ~x_161;
assign n_25389 = ~x_162 & ~x_163;
assign n_25390 =  n_25388 &  n_25389;
assign n_25391 = ~x_156 & ~x_157;
assign n_25392 = ~x_158 & ~x_159;
assign n_25393 =  n_25391 &  n_25392;
assign n_25394 =  n_25390 &  n_25393;
assign n_25395 = ~x_168 & ~x_169;
assign n_25396 = ~x_170 & ~x_171;
assign n_25397 =  n_25395 &  n_25396;
assign n_25398 = ~x_164 & ~x_165;
assign n_25399 = ~x_166 & ~x_167;
assign n_25400 =  n_25398 &  n_25399;
assign n_25401 =  n_25397 &  n_25400;
assign n_25402 =  n_25394 &  n_25401;
assign n_25403 = ~x_144 & ~x_145;
assign n_25404 = ~x_146 & ~x_147;
assign n_25405 =  n_25403 &  n_25404;
assign n_25406 = ~x_140 & ~x_141;
assign n_25407 = ~x_142 & ~x_143;
assign n_25408 =  n_25406 &  n_25407;
assign n_25409 =  n_25405 &  n_25408;
assign n_25410 = ~x_152 & ~x_153;
assign n_25411 = ~x_154 & ~x_155;
assign n_25412 =  n_25410 &  n_25411;
assign n_25413 = ~x_148 & ~x_149;
assign n_25414 = ~x_150 & ~x_151;
assign n_25415 =  n_25413 &  n_25414;
assign n_25416 =  n_25412 &  n_25415;
assign n_25417 =  n_25409 &  n_25416;
assign n_25418 =  n_25402 &  n_25417;
assign n_25419 =  n_25387 &  n_25418;
assign n_25420 = ~x_2367 & ~x_2368;
assign n_25421 = ~x_2369 & ~x_2370;
assign n_25422 =  n_25420 &  n_25421;
assign n_25423 = ~x_2363 & ~x_2364;
assign n_25424 = ~x_2365 & ~x_2366;
assign n_25425 =  n_25423 &  n_25424;
assign n_25426 =  n_25422 &  n_25425;
assign n_25427 = ~x_2375 & ~x_2376;
assign n_25428 = ~x_2377 & ~x_2378;
assign n_25429 =  n_25427 &  n_25428;
assign n_25430 = ~x_2371 & ~x_2372;
assign n_25431 = ~x_2373 & ~x_2374;
assign n_25432 =  n_25430 &  n_25431;
assign n_25433 =  n_25429 &  n_25432;
assign n_25434 =  n_25426 &  n_25433;
assign n_25435 = ~x_2351 & ~x_2352;
assign n_25436 = ~x_2353 & ~x_2354;
assign n_25437 =  n_25435 &  n_25436;
assign n_25438 = ~x_2347 & ~x_2348;
assign n_25439 = ~x_2349 & ~x_2350;
assign n_25440 =  n_25438 &  n_25439;
assign n_25441 =  n_25437 &  n_25440;
assign n_25442 = ~x_2359 & ~x_2360;
assign n_25443 = ~x_2361 & ~x_2362;
assign n_25444 =  n_25442 &  n_25443;
assign n_25445 = ~x_2355 & ~x_2356;
assign n_25446 = ~x_2357 & ~x_2358;
assign n_25447 =  n_25445 &  n_25446;
assign n_25448 =  n_25444 &  n_25447;
assign n_25449 =  n_25441 &  n_25448;
assign n_25450 =  n_25434 &  n_25449;
assign n_25451 =  n_1895 &  n_3616;
assign n_25452 =  n_25450 &  n_25451;
assign n_25453 = ~n_25419 & ~n_25452;
assign n_25454 = ~n_23540 &  n_23541;
assign n_25455 =  n_153 &  n_9;
assign n_25456 = ~x_5052 & ~x_5053;
assign n_25457 = ~x_5054 & ~x_5055;
assign n_25458 =  n_25456 &  n_25457;
assign n_25459 = ~x_5048 & ~x_5049;
assign n_25460 = ~x_5050 & ~x_5051;
assign n_25461 =  n_25459 &  n_25460;
assign n_25462 =  n_25458 &  n_25461;
assign n_25463 = ~x_5060 & ~x_5061;
assign n_25464 = ~x_5062 & ~x_5063;
assign n_25465 =  n_25463 &  n_25464;
assign n_25466 = ~x_5056 & ~x_5057;
assign n_25467 = ~x_5058 & ~x_5059;
assign n_25468 =  n_25466 &  n_25467;
assign n_25469 =  n_25465 &  n_25468;
assign n_25470 =  n_25462 &  n_25469;
assign n_25471 = ~x_5036 & ~x_5037;
assign n_25472 = ~x_5038 & ~x_5039;
assign n_25473 =  n_25471 &  n_25472;
assign n_25474 = ~x_5032 & ~x_5033;
assign n_25475 = ~x_5034 & ~x_5035;
assign n_25476 =  n_25474 &  n_25475;
assign n_25477 =  n_25473 &  n_25476;
assign n_25478 = ~x_5044 & ~x_5045;
assign n_25479 = ~x_5046 & ~x_5047;
assign n_25480 =  n_25478 &  n_25479;
assign n_25481 = ~x_5040 & ~x_5041;
assign n_25482 = ~x_5042 & ~x_5043;
assign n_25483 =  n_25481 &  n_25482;
assign n_25484 =  n_25480 &  n_25483;
assign n_25485 =  n_25477 &  n_25484;
assign n_25486 =  n_25470 &  n_25485;
assign n_25487 =  n_25455 &  n_25486;
assign n_25488 = ~n_25454 & ~n_25487;
assign n_25489 =  n_25453 &  n_25488;
assign n_25490 =  n_21953 &  n_8345;
assign n_25491 =  n_23816 &  n_23993;
assign n_25492 = ~n_25490 & ~n_25491;
assign n_25493 =  x_4137 &  n_1039;
assign n_25494 =  n_353 &  n_25493;
assign n_25495 =  n_769 &  n_25494;
assign n_25496 =  n_11 &  n_25495;
assign n_25497 = ~n_4292 & ~n_25496;
assign n_25498 =  n_25492 &  n_25497;
assign n_25499 = ~x_43 &  n_5655;
assign n_25500 =  n_24924 &  n_25499;
assign n_25501 = ~x_42 &  n_25500;
assign n_25502 =  n_2291 &  n_8361;
assign n_25503 =  n_14264 &  n_24064;
assign n_25504 = ~n_25502 & ~n_25503;
assign n_25505 = ~n_25501 &  n_25504;
assign n_25506 =  n_25498 &  n_25505;
assign n_25507 =  n_25489 &  n_25506;
assign n_25508 =  n_25386 &  n_25507;
assign n_25509 =  n_25336 &  n_25508;
assign n_25510 =  n_23459 &  n_23641;
assign n_25511 = ~x_1547 &  n_25510;
assign n_25512 = ~x_588 &  n_24936;
assign n_25513 = ~n_25511 & ~n_25512;
assign n_25514 =  x_36 &  n_2879;
assign n_25515 =  n_13 &  n_25514;
assign n_25516 =  n_24747 &  n_25515;
assign n_25517 = ~x_3416 &  n_23460;
assign n_25518 =  n_25517 &  n_24769;
assign n_25519 = ~n_25516 & ~n_25518;
assign n_25520 = ~x_3416 &  n_23596;
assign n_25521 = ~n_10477 & ~n_23691;
assign n_25522 =  n_25520 & ~n_25521;
assign n_25523 =  n_25519 & ~n_25522;
assign n_25524 =  n_25513 &  n_25523;
assign n_25525 =  n_1501 &  n_23990;
assign n_25526 =  n_25525 &  n_24896;
assign n_25527 = ~x_3416 &  n_23991;
assign n_25528 = ~x_3448 &  n_23816;
assign n_25529 = ~x_38 &  n_10274;
assign n_25530 =  n_25528 &  n_25529;
assign n_25531 = ~n_25527 & ~n_25530;
assign n_25532 = ~n_25526 &  n_25531;
assign n_25533 =  n_24014 &  n_23374;
assign n_25534 = ~x_3384 &  n_23989;
assign n_25535 =  n_23840 &  n_25534;
assign n_25536 = ~n_25533 & ~n_25535;
assign n_25537 = ~x_4137 &  n_24938;
assign n_25538 = ~x_1771 &  n_24979;
assign n_25539 = ~n_25537 & ~n_25538;
assign n_25540 =  n_25536 &  n_25539;
assign n_25541 =  n_24119 &  n_25528;
assign n_25542 =  n_23613 &  n_23815;
assign n_25543 = ~n_25541 & ~n_25542;
assign n_25544 = ~x_1547 &  n_25250;
assign n_25545 = ~x_1547 &  n_23460;
assign n_25546 =  n_25545 &  n_25242;
assign n_25547 = ~n_25544 & ~n_25546;
assign n_25548 =  n_25543 &  n_25547;
assign n_25549 =  n_25540 &  n_25548;
assign n_25550 =  n_25532 &  n_25549;
assign n_25551 =  n_25524 &  n_25550;
assign n_25552 =  n_349 & ~n_25551;
assign n_25553 =  n_25509 & ~n_25552;
assign n_25554 =  n_25286 &  n_25553;
assign n_25555 =  n_24679 &  n_24222;
assign n_25556 =  n_24306 &  n_21564;
assign n_25557 = ~n_25555 & ~n_25556;
assign n_25558 =  n_3143 &  n_14655;
assign n_25559 = ~x_4349 & ~x_4350;
assign n_25560 = ~x_4351 & ~x_4352;
assign n_25561 =  n_25559 &  n_25560;
assign n_25562 = ~x_4345 & ~x_4346;
assign n_25563 = ~x_4347 & ~x_4348;
assign n_25564 =  n_25562 &  n_25563;
assign n_25565 =  n_25561 &  n_25564;
assign n_25566 = ~x_4357 & ~x_4358;
assign n_25567 = ~x_4359 & ~x_4360;
assign n_25568 =  n_25566 &  n_25567;
assign n_25569 = ~x_4353 & ~x_4354;
assign n_25570 = ~x_4355 & ~x_4356;
assign n_25571 =  n_25569 &  n_25570;
assign n_25572 =  n_25568 &  n_25571;
assign n_25573 =  n_25565 &  n_25572;
assign n_25574 = ~x_4333 & ~x_4334;
assign n_25575 = ~x_4335 & ~x_4336;
assign n_25576 =  n_25574 &  n_25575;
assign n_25577 = ~x_4329 & ~x_4330;
assign n_25578 = ~x_4331 & ~x_4332;
assign n_25579 =  n_25577 &  n_25578;
assign n_25580 =  n_25576 &  n_25579;
assign n_25581 = ~x_4341 & ~x_4342;
assign n_25582 = ~x_4343 & ~x_4344;
assign n_25583 =  n_25581 &  n_25582;
assign n_25584 = ~x_4337 & ~x_4338;
assign n_25585 = ~x_4339 & ~x_4340;
assign n_25586 =  n_25584 &  n_25585;
assign n_25587 =  n_25583 &  n_25586;
assign n_25588 =  n_25580 &  n_25587;
assign n_25589 =  n_25573 &  n_25588;
assign n_25590 =  n_25558 & ~n_25589;
assign n_25591 =  n_2880 &  n_10080;
assign n_25592 = ~x_4157 & ~x_4158;
assign n_25593 = ~x_4159 & ~x_4160;
assign n_25594 =  n_25592 &  n_25593;
assign n_25595 = ~x_4153 & ~x_4154;
assign n_25596 = ~x_4155 & ~x_4156;
assign n_25597 =  n_25595 &  n_25596;
assign n_25598 =  n_25594 &  n_25597;
assign n_25599 = ~x_4165 & ~x_4166;
assign n_25600 = ~x_4167 & ~x_4168;
assign n_25601 =  n_25599 &  n_25600;
assign n_25602 = ~x_4161 & ~x_4162;
assign n_25603 = ~x_4163 & ~x_4164;
assign n_25604 =  n_25602 &  n_25603;
assign n_25605 =  n_25601 &  n_25604;
assign n_25606 =  n_25598 &  n_25605;
assign n_25607 = ~x_4141 & ~x_4142;
assign n_25608 = ~x_4143 & ~x_4144;
assign n_25609 =  n_25607 &  n_25608;
assign n_25610 = ~x_4137 & ~x_4138;
assign n_25611 = ~x_4139 & ~x_4140;
assign n_25612 =  n_25610 &  n_25611;
assign n_25613 =  n_25609 &  n_25612;
assign n_25614 = ~x_4149 & ~x_4150;
assign n_25615 = ~x_4151 & ~x_4152;
assign n_25616 =  n_25614 &  n_25615;
assign n_25617 = ~x_4145 & ~x_4146;
assign n_25618 = ~x_4147 & ~x_4148;
assign n_25619 =  n_25617 &  n_25618;
assign n_25620 =  n_25616 &  n_25619;
assign n_25621 =  n_25613 &  n_25620;
assign n_25622 =  n_25606 &  n_25621;
assign n_25623 =  n_25591 &  n_25622;
assign n_25624 =  n_24468 & ~n_24499;
assign n_25625 =  n_13104 &  n_23844;
assign n_25626 =  n_155 &  n_23987;
assign n_25627 = ~n_25625 & ~n_25626;
assign n_25628 = ~n_25624 &  n_25627;
assign n_25629 = ~n_25623 &  n_25628;
assign n_25630 = ~n_25590 &  n_25629;
assign n_25631 =  n_25557 &  n_25630;
assign n_25632 =  n_1038 &  n_24116;
assign n_25633 =  n_758 &  n_24960;
assign n_25634 =  n_24955 &  n_15917;
assign n_25635 =  n_5645 &  n_25634;
assign n_25636 = ~n_25633 & ~n_25635;
assign n_25637 =  n_23596 &  n_18624;
assign n_25638 =  x_43 &  n_10473;
assign n_25639 = ~n_25637 & ~n_25638;
assign n_25640 =  n_25636 &  n_25639;
assign n_25641 =  n_3341 &  n_24073;
assign n_25642 =  x_43 &  n_25641;
assign n_25643 =  n_9884 &  n_2291;
assign n_25644 = ~n_24423 &  n_25643;
assign n_25645 = ~n_25642 & ~n_25644;
assign n_25646 =  n_25640 &  n_25645;
assign n_25647 = ~n_25632 &  n_25646;
assign n_25648 =  n_18914 &  n_9690;
assign n_25649 =  n_24113 &  n_25648;
assign n_25650 =  n_23884 &  n_2486;
assign n_25651 =  n_9690 &  n_6182;
assign n_25652 =  n_5981 &  n_6182;
assign n_25653 = ~x_43 &  n_25652;
assign n_25654 = ~n_25651 & ~n_25653;
assign n_25655 = ~n_25650 &  n_25654;
assign n_25656 = ~n_25649 &  n_25655;
assign n_25657 =  n_3339 &  n_8354;
assign n_25658 = ~x_42 &  n_6379;
assign n_25659 =  n_6377 &  n_25658;
assign n_25660 = ~x_43 &  n_25659;
assign n_25661 = ~n_25657 & ~n_25660;
assign n_25662 =  n_23683 &  n_24969;
assign n_25663 = ~x_43 &  n_25662;
assign n_25664 = ~x_42 &  n_25663;
assign n_25665 =  n_25661 & ~n_25664;
assign n_25666 =  n_25656 &  n_25665;
assign n_25667 =  n_25647 &  n_25666;
assign n_25668 =  n_25631 &  n_25667;
assign n_25669 =  n_23135 &  n_1503;
assign n_25670 = ~n_3626 & ~n_25669;
assign n_25671 = ~x_39 &  n_1503;
assign n_25672 =  n_9884 &  n_25671;
assign n_25673 = ~n_25672 & ~n_17787;
assign n_25674 =  n_25670 &  n_25673;
assign n_25675 =  n_14785 &  n_23938;
assign n_25676 =  n_154 &  n_25675;
assign n_25677 = ~n_23325 &  n_23326;
assign n_25678 = ~n_25676 & ~n_25677;
assign n_25679 =  n_25674 &  n_25678;
assign n_25680 = ~x_2345 &  n_23322;
assign n_25681 = ~x_2346 &  n_25680;
assign n_25682 = ~x_2315 & ~n_25681;
assign n_25683 =  n_14264 &  n_355;
assign n_25684 =  n_25682 &  n_25683;
assign n_25685 =  n_25271 & ~n_25273;
assign n_25686 = ~n_25684 & ~n_25685;
assign n_25687 =  n_25679 &  n_25686;
assign n_25688 =  n_25668 &  n_25687;
assign n_25689 =  n_150 & ~n_22971;
assign n_25690 =  n_24015 &  n_25689;
assign n_25691 =  n_6379 & ~n_25266;
assign n_25692 =  n_556 &  n_13104;
assign n_25693 =  n_25691 &  n_25692;
assign n_25694 = ~n_25690 & ~n_25693;
assign n_25695 = ~n_25682 &  n_25683;
assign n_25696 = ~x_2315 & ~n_25680;
assign n_25697 =  n_5645 &  n_12292;
assign n_25698 =  n_25696 &  n_25697;
assign n_25699 = ~n_25695 & ~n_25698;
assign n_25700 =  n_8365 &  n_3619;
assign n_25701 = ~n_25696 &  n_25700;
assign n_25702 =  n_25699 & ~n_25701;
assign n_25703 =  n_25694 &  n_25702;
assign n_25704 =  n_25688 &  n_25703;
assign n_25705 =  n_25554 &  n_25704;
assign n_25706 =  n_25260 &  n_25705;
assign n_25707 =  n_23838 &  n_25706;
assign n_25708 = ~n_22939 &  n_25707;
assign n_25709 = ~n_22720 &  n_25708;
assign n_25710 = ~n_22591 &  n_25709;
assign n_25711 =  n_22464 &  n_25710;
assign n_25712 = ~n_22209 &  n_25711;
assign n_25713 = ~n_22082 &  n_25712;
assign n_25714 =  x_43 &  n_25713;
assign n_25715 = ~x_43 & ~n_25713;
assign n_25716 = ~n_25714 & ~n_25715;
assign n_25717 = ~n_22717 & ~n_22209;
assign n_25718 =  n_5652 &  n_3615;
assign n_25719 = ~x_108 &  x_204;
assign n_25720 =  x_108 & ~x_204;
assign n_25721 =  x_109 & ~x_205;
assign n_25722 = ~x_109 &  x_205;
assign n_25723 =  x_110 & ~x_206;
assign n_25724 = ~x_110 &  x_206;
assign n_25725 =  x_111 & ~x_207;
assign n_25726 = ~x_111 &  x_207;
assign n_25727 =  x_112 & ~x_208;
assign n_25728 = ~x_112 &  x_208;
assign n_25729 =  x_113 & ~x_209;
assign n_25730 = ~x_113 &  x_209;
assign n_25731 =  x_114 & ~x_210;
assign n_25732 = ~x_114 &  x_210;
assign n_25733 =  x_115 & ~x_211;
assign n_25734 = ~x_115 &  x_211;
assign n_25735 =  x_116 & ~x_212;
assign n_25736 = ~x_116 &  x_212;
assign n_25737 =  x_117 & ~x_213;
assign n_25738 = ~x_117 &  x_213;
assign n_25739 =  x_118 & ~x_214;
assign n_25740 = ~x_118 &  x_214;
assign n_25741 =  x_119 & ~x_215;
assign n_25742 = ~x_119 &  x_215;
assign n_25743 =  x_120 & ~x_216;
assign n_25744 = ~x_120 &  x_216;
assign n_25745 =  x_121 & ~x_217;
assign n_25746 = ~x_121 &  x_217;
assign n_25747 =  x_122 & ~x_218;
assign n_25748 = ~x_122 &  x_218;
assign n_25749 =  x_123 & ~x_219;
assign n_25750 = ~x_123 &  x_219;
assign n_25751 =  x_124 & ~x_220;
assign n_25752 = ~x_124 &  x_220;
assign n_25753 =  x_125 & ~x_221;
assign n_25754 = ~x_125 &  x_221;
assign n_25755 =  x_126 & ~x_222;
assign n_25756 = ~x_126 &  x_222;
assign n_25757 =  x_127 & ~x_223;
assign n_25758 = ~x_127 &  x_223;
assign n_25759 =  x_128 & ~x_224;
assign n_25760 = ~x_128 &  x_224;
assign n_25761 =  x_129 & ~x_225;
assign n_25762 = ~x_129 &  x_225;
assign n_25763 =  x_130 & ~x_226;
assign n_25764 = ~x_130 &  x_226;
assign n_25765 =  x_131 & ~x_227;
assign n_25766 = ~x_131 &  x_227;
assign n_25767 =  x_132 & ~x_228;
assign n_25768 = ~x_132 &  x_228;
assign n_25769 =  x_133 & ~x_229;
assign n_25770 = ~x_133 &  x_229;
assign n_25771 =  x_134 & ~x_230;
assign n_25772 = ~x_134 &  x_230;
assign n_25773 =  x_135 & ~x_231;
assign n_25774 = ~x_135 &  x_231;
assign n_25775 =  x_136 & ~x_232;
assign n_25776 = ~x_136 &  x_232;
assign n_25777 =  x_138 & ~x_234;
assign n_25778 = ~x_138 &  x_234;
assign n_25779 =  x_139 & ~x_235;
assign n_25780 = ~n_25778 &  n_25779;
assign n_25781 = ~n_25777 & ~n_25780;
assign n_25782 =  x_233 &  n_25781;
assign n_25783 =  x_137 & ~n_25782;
assign n_25784 = ~x_233 & ~n_25781;
assign n_25785 = ~n_25783 & ~n_25784;
assign n_25786 = ~n_25776 & ~n_25785;
assign n_25787 = ~n_25775 & ~n_25786;
assign n_25788 = ~n_25774 & ~n_25787;
assign n_25789 = ~n_25773 & ~n_25788;
assign n_25790 = ~n_25772 & ~n_25789;
assign n_25791 = ~n_25771 & ~n_25790;
assign n_25792 = ~n_25770 & ~n_25791;
assign n_25793 = ~n_25769 & ~n_25792;
assign n_25794 = ~n_25768 & ~n_25793;
assign n_25795 = ~n_25767 & ~n_25794;
assign n_25796 = ~n_25766 & ~n_25795;
assign n_25797 = ~n_25765 & ~n_25796;
assign n_25798 = ~n_25764 & ~n_25797;
assign n_25799 = ~n_25763 & ~n_25798;
assign n_25800 = ~n_25762 & ~n_25799;
assign n_25801 = ~n_25761 & ~n_25800;
assign n_25802 = ~n_25760 & ~n_25801;
assign n_25803 = ~n_25759 & ~n_25802;
assign n_25804 = ~n_25758 & ~n_25803;
assign n_25805 = ~n_25757 & ~n_25804;
assign n_25806 = ~n_25756 & ~n_25805;
assign n_25807 = ~n_25755 & ~n_25806;
assign n_25808 = ~n_25754 & ~n_25807;
assign n_25809 = ~n_25753 & ~n_25808;
assign n_25810 = ~n_25752 & ~n_25809;
assign n_25811 = ~n_25751 & ~n_25810;
assign n_25812 = ~n_25750 & ~n_25811;
assign n_25813 = ~n_25749 & ~n_25812;
assign n_25814 = ~n_25748 & ~n_25813;
assign n_25815 = ~n_25747 & ~n_25814;
assign n_25816 = ~n_25746 & ~n_25815;
assign n_25817 = ~n_25745 & ~n_25816;
assign n_25818 = ~n_25744 & ~n_25817;
assign n_25819 = ~n_25743 & ~n_25818;
assign n_25820 = ~n_25742 & ~n_25819;
assign n_25821 = ~n_25741 & ~n_25820;
assign n_25822 = ~n_25740 & ~n_25821;
assign n_25823 = ~n_25739 & ~n_25822;
assign n_25824 = ~n_25738 & ~n_25823;
assign n_25825 = ~n_25737 & ~n_25824;
assign n_25826 = ~n_25736 & ~n_25825;
assign n_25827 = ~n_25735 & ~n_25826;
assign n_25828 = ~n_25734 & ~n_25827;
assign n_25829 = ~n_25733 & ~n_25828;
assign n_25830 = ~n_25732 & ~n_25829;
assign n_25831 = ~n_25731 & ~n_25830;
assign n_25832 = ~n_25730 & ~n_25831;
assign n_25833 = ~n_25729 & ~n_25832;
assign n_25834 = ~n_25728 & ~n_25833;
assign n_25835 = ~n_25727 & ~n_25834;
assign n_25836 = ~n_25726 & ~n_25835;
assign n_25837 = ~n_25725 & ~n_25836;
assign n_25838 = ~n_25724 & ~n_25837;
assign n_25839 = ~n_25723 & ~n_25838;
assign n_25840 = ~n_25722 & ~n_25839;
assign n_25841 = ~n_25721 & ~n_25840;
assign n_25842 = ~n_25720 & ~n_25841;
assign n_25843 = ~n_25719 & ~n_25842;
assign n_25844 =  n_25718 &  n_25843;
assign n_25845 =  n_22083 & ~n_22208;
assign n_25846 =  n_22465 &  n_22590;
assign n_25847 =  n_23178 &  n_25261;
assign n_25848 =  n_23292 &  n_24776;
assign n_25849 = ~n_25847 & ~n_25848;
assign n_25850 =  n_23624 & ~n_23610;
assign n_25851 =  n_24753 &  n_23619;
assign n_25852 = ~n_25851 & ~n_23985;
assign n_25853 = ~n_25850 &  n_25852;
assign n_25854 =  n_25849 &  n_25853;
assign n_25855 =  n_25265 &  n_25854;
assign n_25856 =  n_5651 &  n_3143;
assign n_25857 =  n_23987 &  n_25856;
assign n_25858 = ~n_25226 & ~n_25857;
assign n_25859 = ~n_2292 & ~n_24689;
assign n_25860 =  n_25858 &  n_25859;
assign n_25861 = ~n_12910 &  n_25860;
assign n_25862 =  n_25558 &  n_25589;
assign n_25863 =  n_23840 &  n_23549;
assign n_25864 =  n_6877 &  n_2684;
assign n_25865 =  n_24628 &  n_3623;
assign n_25866 = ~n_25864 & ~n_25865;
assign n_25867 = ~n_25863 &  n_25866;
assign n_25868 = ~n_23940 &  n_25867;
assign n_25869 = ~n_25862 &  n_25868;
assign n_25870 =  n_25861 &  n_25869;
assign n_25871 =  n_1895 &  n_23675;
assign n_25872 = ~n_25871 & ~n_24070;
assign n_25873 =  n_6379 &  n_23375;
assign n_25874 =  n_25873 &  n_23244;
assign n_25875 =  n_25872 & ~n_25874;
assign n_25876 =  n_1895 &  n_14785;
assign n_25877 = ~n_25876 & ~n_24036;
assign n_25878 =  n_758 &  n_12292;
assign n_25879 = ~n_23813 & ~n_25878;
assign n_25880 =  n_25877 &  n_25879;
assign n_25881 =  n_25875 &  n_25880;
assign n_25882 =  n_2095 &  n_23253;
assign n_25883 =  n_25882 & ~n_25273;
assign n_25884 = ~n_25047 &  n_24501;
assign n_25885 = ~n_25883 &  n_25884;
assign n_25886 =  n_25881 &  n_25885;
assign n_25887 =  n_25870 &  n_25886;
assign n_25888 =  n_25855 &  n_25887;
assign n_25889 =  n_23635 &  n_25888;
assign n_25890 =  n_349 &  n_24739;
assign n_25891 = ~n_25890 & ~n_24939;
assign n_25892 =  n_23596 &  n_23692;
assign n_25893 = ~n_24311 & ~n_25892;
assign n_25894 =  n_25891 &  n_25893;
assign n_25895 =  x_1547 &  n_2879;
assign n_25896 =  n_23460 &  n_25895;
assign n_25897 =  n_8054 &  n_25896;
assign n_25898 = ~n_24947 & ~n_25897;
assign n_25899 =  n_349 &  n_24909;
assign n_25900 =  n_24788 &  n_25899;
assign n_25901 = ~n_24121 & ~n_25900;
assign n_25902 =  n_25898 &  n_25901;
assign n_25903 =  n_25894 &  n_25902;
assign n_25904 =  n_6525 &  n_23687;
assign n_25905 =  n_5654 &  n_23991;
assign n_25906 = ~n_25904 & ~n_25905;
assign n_25907 =  n_5656 &  n_8354;
assign n_25908 = ~n_24051 & ~n_25907;
assign n_25909 =  n_25906 &  n_25908;
assign n_25910 =  x_37 &  n_24788;
assign n_25911 =  n_20790 &  n_25910;
assign n_25912 = ~n_25036 & ~n_5657;
assign n_25913 = ~n_25911 &  n_25912;
assign n_25914 = ~n_19694 & ~n_25175;
assign n_25915 =  n_25913 &  n_25914;
assign n_25916 =  n_25909 &  n_25915;
assign n_25917 =  n_25903 &  n_25916;
assign n_25918 =  n_23843 &  n_23178;
assign n_25919 = ~n_24307 & ~n_25918;
assign n_25920 = ~n_25016 &  n_25919;
assign n_25921 =  n_1895 &  n_2290;
assign n_25922 =  n_23816 &  n_25921;
assign n_25923 =  n_349 &  n_23384;
assign n_25924 = ~n_25922 & ~n_25923;
assign n_25925 =  n_25920 &  n_25924;
assign n_25926 = ~n_24532 & ~n_25028;
assign n_25927 =  n_24967 &  n_14;
assign n_25928 = ~n_23550 & ~n_25927;
assign n_25929 =  n_25926 &  n_25928;
assign n_25930 = ~n_3145 & ~n_24778;
assign n_25931 =  n_7078 &  n_1306;
assign n_25932 = ~n_10476 & ~n_25931;
assign n_25933 =  n_25930 &  n_25932;
assign n_25934 =  n_25929 &  n_25933;
assign n_25935 =  n_25925 &  n_25934;
assign n_25936 =  n_23942 &  n_8361;
assign n_25937 =  n_21954 &  n_23422;
assign n_25938 = ~n_25936 & ~n_25937;
assign n_25939 =  n_349 &  n_25495;
assign n_25940 =  n_758 &  n_25634;
assign n_25941 = ~n_25939 & ~n_25940;
assign n_25942 =  n_25938 &  n_25941;
assign n_25943 =  n_23816 &  n_14264;
assign n_25944 = ~n_25943 & ~n_23247;
assign n_25945 = ~n_25105 & ~n_24959;
assign n_25946 =  n_25944 &  n_25945;
assign n_25947 =  n_25942 &  n_25946;
assign n_25948 =  n_25935 &  n_25947;
assign n_25949 =  n_25917 &  n_25948;
assign n_25950 = ~n_1037 & ~n_349;
assign n_25951 = ~n_25950 &  n_24026;
assign n_25952 = ~n_1038 & ~n_3143;
assign n_25953 = ~n_25952 &  n_25153;
assign n_25954 = ~n_25951 & ~n_25953;
assign n_25955 =  n_1895 &  n_25107;
assign n_25956 =  n_17782 &  n_23554;
assign n_25957 = ~n_25955 & ~n_25956;
assign n_25958 =  n_25954 &  n_25957;
assign n_25959 = ~n_23254 & ~n_24004;
assign n_25960 = ~n_8055 &  n_23141;
assign n_25961 =  n_25959 &  n_25960;
assign n_25962 =  n_25958 &  n_25961;
assign n_25963 =  n_351 &  n_24684;
assign n_25964 = ~n_13873 & ~n_25963;
assign n_25965 = ~n_25950 &  n_24018;
assign n_25966 = ~n_25965 & ~n_1308;
assign n_25967 =  n_25964 &  n_25966;
assign n_25968 =  n_24909 &  n_10079;
assign n_25969 =  n_10872 &  n_23607;
assign n_25970 = ~n_25968 & ~n_25969;
assign n_25971 =  n_6882 &  n_551;
assign n_25972 =  n_1 &  n_25971;
assign n_25973 = ~x_43 &  n_25972;
assign n_25974 =  n_25970 & ~n_25973;
assign n_25975 =  n_3623 &  n_1503;
assign n_25976 = ~n_24042 & ~n_25975;
assign n_25977 =  n_25974 &  n_25976;
assign n_25978 =  n_25967 &  n_25977;
assign n_25979 =  n_25962 &  n_25978;
assign n_25980 =  n_8054 &  n_15;
assign n_25981 = ~n_23053 & ~n_25980;
assign n_25982 =  n_24015 &  n_24069;
assign n_25983 = ~n_7080 & ~n_25982;
assign n_25984 =  n_25981 &  n_25983;
assign n_25985 =  n_8361 &  n_6526;
assign n_25986 =  n_23883 &  n_6877;
assign n_25987 = ~n_25985 & ~n_25986;
assign n_25988 =  n_8354 &  n_23549;
assign n_25989 = ~n_25247 & ~n_25988;
assign n_25990 =  n_25987 &  n_25989;
assign n_25991 =  n_25984 &  n_25990;
assign n_25992 = ~n_25625 & ~n_21565;
assign n_25993 =  n_2879 &  n_3625;
assign n_25994 =  n_354 &  n_25993;
assign n_25995 = ~n_13479 & ~n_25994;
assign n_25996 =  n_25992 &  n_25995;
assign n_25997 = ~x_43 &  n_6884;
assign n_25998 =  n_1895 &  n_23945;
assign n_25999 = ~n_25997 & ~n_25998;
assign n_26000 =  n_24066 &  n_25999;
assign n_26001 =  n_25996 &  n_26000;
assign n_26002 =  n_25991 &  n_26001;
assign n_26003 =  n_25979 &  n_26002;
assign n_26004 =  n_25949 &  n_26003;
assign n_26005 =  n_23051 &  n_23888;
assign n_26006 =  n_11 &  n_26005;
assign n_26007 =  n_23815 &  n_26006;
assign n_26008 =  n_1899 &  n_23990;
assign n_26009 =  n_5654 &  n_26008;
assign n_26010 =  n_23462 &  n_25244;
assign n_26011 = ~n_26009 & ~n_26010;
assign n_26012 = ~n_26007 &  n_26011;
assign n_26013 =  n_6378 &  n_2684;
assign n_26014 =  n_23816 &  n_155;
assign n_26015 = ~n_26013 & ~n_26014;
assign n_26016 =  n_23850 &  n_26015;
assign n_26017 =  n_26012 &  n_26016;
assign n_26018 = ~n_24192 &  n_24194;
assign n_26019 = ~n_26018 & ~n_25219;
assign n_26020 =  n_150 &  n_25856;
assign n_26021 =  n_24314 &  n_6876;
assign n_26022 = ~n_26020 & ~n_26021;
assign n_26023 =  n_349 &  n_4286;
assign n_26024 =  n_26022 & ~n_26023;
assign n_26025 =  n_26019 &  n_26024;
assign n_26026 =  n_26017 &  n_26025;
assign n_26027 =  n_24628 &  n_7078;
assign n_26028 = ~n_26027 & ~n_25157;
assign n_26029 =  n_26028 &  n_24593;
assign n_26030 =  n_24956 &  n_23636;
assign n_26031 = ~n_26030 & ~n_24016;
assign n_26032 =  n_9884 &  n_13230;
assign n_26033 = ~x_1375 & ~x_1376;
assign n_26034 = ~x_1377 & ~x_1378;
assign n_26035 =  n_26033 &  n_26034;
assign n_26036 = ~x_1371 & ~x_1372;
assign n_26037 = ~x_1373 & ~x_1374;
assign n_26038 =  n_26036 &  n_26037;
assign n_26039 =  n_26035 &  n_26038;
assign n_26040 = ~x_1383 & ~x_1384;
assign n_26041 = ~x_1385 & ~x_1386;
assign n_26042 =  n_26040 &  n_26041;
assign n_26043 = ~x_1379 & ~x_1380;
assign n_26044 = ~x_1381 & ~x_1382;
assign n_26045 =  n_26043 &  n_26044;
assign n_26046 =  n_26042 &  n_26045;
assign n_26047 =  n_26039 &  n_26046;
assign n_26048 = ~x_1359 & ~x_1360;
assign n_26049 = ~x_1361 & ~x_1362;
assign n_26050 =  n_26048 &  n_26049;
assign n_26051 = ~x_1355 & ~x_1356;
assign n_26052 = ~x_1357 & ~x_1358;
assign n_26053 =  n_26051 &  n_26052;
assign n_26054 =  n_26050 &  n_26053;
assign n_26055 = ~x_1367 & ~x_1368;
assign n_26056 = ~x_1369 & ~x_1370;
assign n_26057 =  n_26055 &  n_26056;
assign n_26058 = ~x_1363 & ~x_1364;
assign n_26059 = ~x_1365 & ~x_1366;
assign n_26060 =  n_26058 &  n_26059;
assign n_26061 =  n_26057 &  n_26060;
assign n_26062 =  n_26054 &  n_26061;
assign n_26063 =  n_26047 &  n_26062;
assign n_26064 =  n_26032 &  n_26063;
assign n_26065 =  n_26031 & ~n_26064;
assign n_26066 =  n_26029 &  n_26065;
assign n_26067 =  n_5654 &  n_24119;
assign n_26068 =  n_23596 &  n_26067;
assign n_26069 = ~n_2488 & ~n_26068;
assign n_26070 =  n_557 &  n_24069;
assign n_26071 =  n_2880 &  n_24269;
assign n_26072 = ~n_26070 & ~n_26071;
assign n_26073 =  n_26069 &  n_26072;
assign n_26074 =  n_23389 & ~n_23420;
assign n_26075 = ~n_3349 & ~n_26074;
assign n_26076 =  n_26073 &  n_26075;
assign n_26077 =  n_26066 &  n_26076;
assign n_26078 =  n_26026 &  n_26077;
assign n_26079 =  n_349 &  n_26005;
assign n_26080 =  n_26079 &  n_23815;
assign n_26081 =  n_23011 &  n_23815;
assign n_26082 = ~n_26081 & ~n_25542;
assign n_26083 =  n_349 & ~n_26082;
assign n_26084 = ~n_26080 & ~n_26083;
assign n_26085 =  n_24955 &  n_25515;
assign n_26086 =  n_349 &  n_26085;
assign n_26087 =  n_349 &  n_25516;
assign n_26088 = ~n_26086 & ~n_26087;
assign n_26089 =  n_26088 & ~n_24893;
assign n_26090 =  n_26084 &  n_26089;
assign n_26091 =  n_349 &  n_25510;
assign n_26092 =  n_23174 &  n_24575;
assign n_26093 = ~n_25952 &  n_25971;
assign n_26094 = ~n_26092 & ~n_26093;
assign n_26095 =  n_757 &  n_8054;
assign n_26096 = ~n_25952 &  n_24575;
assign n_26097 = ~n_26095 & ~n_26096;
assign n_26098 =  n_26094 &  n_26097;
assign n_26099 = ~n_26091 &  n_26098;
assign n_26100 =  n_2095 &  n_155;
assign n_26101 = ~n_23900 & ~n_26100;
assign n_26102 =  n_23883 &  n_23375;
assign n_26103 =  n_26101 & ~n_26102;
assign n_26104 =  n_26099 &  n_26103;
assign n_26105 =  n_26090 &  n_26104;
assign n_26106 =  x_3416 &  n_23460;
assign n_26107 =  n_24769 &  n_26106;
assign n_26108 =  n_349 &  n_26107;
assign n_26109 =  n_2 &  n_20401;
assign n_26110 =  n_8359 &  n_26109;
assign n_26111 = ~n_25251 & ~n_26110;
assign n_26112 = ~n_26108 &  n_26111;
assign n_26113 =  n_3338 &  n_23052;
assign n_26114 =  n_349 &  n_26113;
assign n_26115 =  n_24320 & ~n_26114;
assign n_26116 =  n_26112 &  n_26115;
assign n_26117 = ~n_25150 &  n_23066;
assign n_26118 =  n_4089 &  n_24043;
assign n_26119 =  n_19497 &  n_6525;
assign n_26120 = ~n_26118 & ~n_26119;
assign n_26121 = ~n_26117 &  n_26120;
assign n_26122 =  n_153 &  n_10078;
assign n_26123 = ~n_23067 & ~n_26122;
assign n_26124 =  n_1040 & ~n_26123;
assign n_26125 = ~n_24937 & ~n_26124;
assign n_26126 =  n_26121 &  n_26125;
assign n_26127 =  n_26116 &  n_26126;
assign n_26128 =  n_26105 &  n_26127;
assign n_26129 =  n_26078 &  n_26128;
assign n_26130 =  n_26004 &  n_26129;
assign n_26131 =  n_7078 &  n_1698;
assign n_26132 = ~n_358 & ~n_26131;
assign n_26133 =  n_23820 &  n_6525;
assign n_26134 = ~n_26133 & ~n_25626;
assign n_26135 =  n_23883 &  n_155;
assign n_26136 = ~n_26135 & ~n_24057;
assign n_26137 =  n_26134 &  n_26136;
assign n_26138 =  n_26132 &  n_26137;
assign n_26139 =  n_24426 &  n_25289;
assign n_26140 =  n_24119 &  n_26006;
assign n_26141 =  n_2486 &  n_21758;
assign n_26142 =  n_26141 & ~n_25206;
assign n_26143 = ~n_26140 & ~n_26142;
assign n_26144 = ~n_26139 &  n_26143;
assign n_26145 =  n_26138 &  n_26144;
assign n_26146 =  n_25223 &  n_25525;
assign n_26147 =  n_11 &  n_26146;
assign n_26148 = ~n_25225 & ~n_26147;
assign n_26149 =  n_3143 &  n_1307;
assign n_26150 = ~n_26149 & ~n_24996;
assign n_26151 = ~n_1505 &  n_26150;
assign n_26152 =  n_26148 &  n_26151;
assign n_26153 = ~x_2394 &  n_24507;
assign n_26154 =  n_24782 &  n_26153;
assign n_26155 = ~x_43 &  n_24074;
assign n_26156 = ~x_43 &  n_25231;
assign n_26157 = ~n_10870 & ~n_26156;
assign n_26158 = ~n_26155 &  n_26157;
assign n_26159 = ~n_26154 &  n_26158;
assign n_26160 =  n_26152 &  n_26159;
assign n_26161 =  n_26145 &  n_26160;
assign n_26162 =  n_349 &  n_26146;
assign n_26163 =  n_25525 &  n_24897;
assign n_26164 = ~x_42 &  n_26163;
assign n_26165 = ~n_26162 & ~n_26164;
assign n_26166 =  n_6378 &  n_23685;
assign n_26167 = ~n_26166 & ~n_24685;
assign n_26168 =  n_5652 &  n_2684;
assign n_26169 =  n_26167 & ~n_26168;
assign n_26170 =  n_26165 &  n_26169;
assign n_26171 =  n_758 &  n_20402;
assign n_26172 = ~n_26171 & ~n_25082;
assign n_26173 =  n_22940 &  n_3615;
assign n_26174 =  n_6525 &  n_14785;
assign n_26175 = ~n_26173 & ~n_26174;
assign n_26176 =  n_26172 &  n_26175;
assign n_26177 =  n_26170 &  n_26176;
assign n_26178 =  n_3144 &  n_354;
assign n_26179 = ~n_24771 &  n_26178;
assign n_26180 =  n_23595 &  n_25589;
assign n_26181 = ~n_23841 & ~n_24520;
assign n_26182 = ~n_26180 &  n_26181;
assign n_26183 = ~n_26179 &  n_26182;
assign n_26184 =  n_26005 &  n_14264;
assign n_26185 =  n_23011 &  n_23012;
assign n_26186 = ~n_24120 & ~n_26185;
assign n_26187 =  n_349 & ~n_26186;
assign n_26188 = ~n_26184 & ~n_26187;
assign n_26189 =  n_1042 &  n_6180;
assign n_26190 = ~x_43 &  n_26189;
assign n_26191 =  n_26188 & ~n_26190;
assign n_26192 =  n_26183 &  n_26191;
assign n_26193 =  n_26177 &  n_26192;
assign n_26194 =  n_26161 &  n_26193;
assign n_26195 =  n_24746 &  n_24956;
assign n_26196 =  n_349 &  n_26195;
assign n_26197 = ~n_25211 & ~n_26196;
assign n_26198 =  n_7078 &  n_23052;
assign n_26199 = ~n_24926 & ~n_26198;
assign n_26200 =  n_26197 &  n_26199;
assign n_26201 =  n_349 &  n_25330;
assign n_26202 = ~n_26201 & ~n_25214;
assign n_26203 = ~n_24425 &  n_26202;
assign n_26204 =  n_26200 &  n_26203;
assign n_26205 =  n_3143 &  n_25634;
assign n_26206 = ~n_26205 & ~n_24961;
assign n_26207 =  n_24688 &  n_26206;
assign n_26208 =  n_26207 & ~n_23880;
assign n_26209 =  n_24306 &  n_2682;
assign n_26210 =  n_2095 &  n_24967;
assign n_26211 = ~n_26209 & ~n_26210;
assign n_26212 =  n_23692 &  n_23011;
assign n_26213 = ~n_23693 & ~n_26212;
assign n_26214 =  n_26211 &  n_26213;
assign n_26215 =  n_8353 &  n_24306;
assign n_26216 = ~n_25556 & ~n_26215;
assign n_26217 =  n_153 &  n_24044;
assign n_26218 =  n_26216 & ~n_26217;
assign n_26219 =  n_26214 &  n_26218;
assign n_26220 =  n_26219 &  n_23892;
assign n_26221 =  n_26208 &  n_26220;
assign n_26222 =  n_26204 &  n_26221;
assign n_26223 = ~n_23676 &  n_23996;
assign n_26224 =  n_16495 &  n_24789;
assign n_26225 =  n_25239 & ~n_25206;
assign n_26226 = ~n_26224 & ~n_26225;
assign n_26227 = ~n_16689 & ~n_3347;
assign n_26228 =  n_26226 &  n_26227;
assign n_26229 =  n_26223 &  n_26228;
assign n_26230 =  n_24695 & ~n_24783;
assign n_26231 =  n_2094 &  n_24786;
assign n_26232 =  n_3345 & ~n_26231;
assign n_26233 =  n_26230 &  n_26232;
assign n_26234 =  n_26229 &  n_26233;
assign n_26235 =  n_26222 &  n_26234;
assign n_26236 =  n_26194 &  n_26235;
assign n_26237 =  n_26130 &  n_26236;
assign n_26238 = ~n_25173 & ~n_25098;
assign n_26239 = ~n_13868 &  n_26238;
assign n_26240 = ~x_43 &  n_24922;
assign n_26241 = ~n_23901 & ~n_24982;
assign n_26242 = ~n_2097 & ~n_23943;
assign n_26243 =  n_26241 &  n_26242;
assign n_26244 = ~n_26240 &  n_26243;
assign n_26245 =  n_26239 &  n_26244;
assign n_26246 =  n_18914 & ~n_24113;
assign n_26247 =  n_26246 &  n_8365;
assign n_26248 =  n_23942 &  n_6525;
assign n_26249 = ~n_26248 & ~n_18915;
assign n_26250 = ~n_23818 &  n_26249;
assign n_26251 = ~n_26247 &  n_26250;
assign n_26252 =  n_26251 & ~n_23680;
assign n_26253 =  n_26245 &  n_26252;
assign n_26254 =  n_23694 &  n_23725;
assign n_26255 = ~n_24195 & ~n_24632;
assign n_26256 = ~n_26254 &  n_26255;
assign n_26257 =  n_23691 &  n_26079;
assign n_26258 =  n_555 &  n_26246;
assign n_26259 = ~n_26257 & ~n_26258;
assign n_26260 =  n_26256 &  n_26259;
assign n_26261 =  n_24356 &  n_23174;
assign n_26262 =  n_554 &  n_24356;
assign n_26263 = ~n_26261 & ~n_26262;
assign n_26264 =  n_150 &  n_6876;
assign n_26265 =  n_26263 & ~n_26264;
assign n_26266 =  n_26265 &  n_23472;
assign n_26267 =  n_26260 &  n_26266;
assign n_26268 =  n_26253 &  n_26267;
assign n_26269 =  n_8359 &  n_24630;
assign n_26270 = ~n_14265 & ~n_26269;
assign n_26271 = ~n_25088 & ~n_25010;
assign n_26272 =  n_26270 &  n_26271;
assign n_26273 = ~n_25685 &  n_26272;
assign n_26274 = ~n_22973 &  n_26273;
assign n_26275 =  n_26268 &  n_26274;
assign n_26276 = ~x_43 &  n_24577;
assign n_26277 = ~n_25152 & ~n_26276;
assign n_26278 =  n_23423 &  n_23454;
assign n_26279 =  n_23134 &  n_23804;
assign n_26280 = ~n_26278 & ~n_26279;
assign n_26281 =  n_26277 &  n_26280;
assign n_26282 = ~n_10081 & ~n_10277;
assign n_26283 =  n_23816 &  n_18624;
assign n_26284 = ~n_26283 & ~n_24933;
assign n_26285 =  n_26282 &  n_26284;
assign n_26286 =  n_8348 & ~n_25950;
assign n_26287 = ~n_24918 & ~n_26286;
assign n_26288 = ~n_23803 &  n_26287;
assign n_26289 =  n_26285 &  n_26288;
assign n_26290 =  n_26281 &  n_26289;
assign n_26291 =  n_349 &  n_25081;
assign n_26292 = ~n_25950 &  n_25116;
assign n_26293 = ~n_25950 &  n_763;
assign n_26294 = ~n_26292 & ~n_26293;
assign n_26295 = ~n_26291 &  n_26294;
assign n_26296 =  n_349 &  n_25533;
assign n_26297 =  n_25155 & ~n_26296;
assign n_26298 =  n_1173 &  n_760;
assign n_26299 =  n_26298 &  n_23592;
assign n_26300 = ~x_42 &  n_24028;
assign n_26301 = ~x_43 &  n_26300;
assign n_26302 = ~n_26299 & ~n_26301;
assign n_26303 =  n_26297 &  n_26302;
assign n_26304 =  n_26295 &  n_26303;
assign n_26305 =  n_26290 &  n_26304;
assign n_26306 =  n_23375 &  n_24069;
assign n_26307 = ~n_24916 & ~n_26306;
assign n_26308 = ~n_13673 & ~n_21371;
assign n_26309 =  n_26307 &  n_26308;
assign n_26310 = ~n_24527 & ~n_24124;
assign n_26311 =  n_758 &  n_20077;
assign n_26312 = ~n_24682 & ~n_26311;
assign n_26313 =  n_26310 &  n_26312;
assign n_26314 =  n_26309 &  n_26313;
assign n_26315 =  n_24910 &  n_26106;
assign n_26316 = ~n_24989 & ~n_6184;
assign n_26317 = ~n_26315 &  n_26316;
assign n_26318 =  n_8361 &  n_13230;
assign n_26319 = ~n_13231 & ~n_26318;
assign n_26320 =  n_26319 & ~n_23365;
assign n_26321 =  n_26317 &  n_26320;
assign n_26322 =  n_26314 &  n_26321;
assign n_26323 = ~n_24113 &  n_25648;
assign n_26324 = ~n_23176 & ~n_23179;
assign n_26325 = ~n_26323 &  n_26324;
assign n_26326 =  n_24435 &  n_24466;
assign n_26327 = ~n_25624 & ~n_26326;
assign n_26328 =  n_26325 &  n_26327;
assign n_26329 = ~n_16882 & ~n_25000;
assign n_26330 =  n_24306 &  n_760;
assign n_26331 = ~n_24315 & ~n_26330;
assign n_26332 =  n_26329 &  n_26331;
assign n_26333 =  n_11 &  n_24159;
assign n_26334 =  n_26333 &  n_24563;
assign n_26335 =  n_349 &  n_24979;
assign n_26336 =  n_23461 &  n_25242;
assign n_26337 = ~n_26335 & ~n_26336;
assign n_26338 = ~n_26334 &  n_26337;
assign n_26339 =  n_26332 &  n_26338;
assign n_26340 =  n_26328 &  n_26339;
assign n_26341 =  n_26322 &  n_26340;
assign n_26342 =  n_26305 &  n_26341;
assign n_26343 =  n_5654 &  n_24938;
assign n_26344 = ~n_26343 & ~n_7662;
assign n_26345 =  n_4288 &  n_24680;
assign n_26346 =  n_24531 & ~n_26345;
assign n_26347 = ~n_13871 &  n_26346;
assign n_26348 =  n_26344 &  n_26347;
assign n_26349 =  n_25696 &  n_25700;
assign n_26350 =  n_760 &  n_23840;
assign n_26351 =  n_25910 &  n_23683;
assign n_26352 =  n_349 &  n_26351;
assign n_26353 =  n_9884 &  n_25287;
assign n_26354 = ~n_26352 & ~n_26353;
assign n_26355 = ~n_26350 &  n_26354;
assign n_26356 = ~n_26349 &  n_26355;
assign n_26357 =  n_26348 &  n_26356;
assign n_26358 =  n_349 &  n_25224;
assign n_26359 =  n_349 &  n_25279;
assign n_26360 = ~n_26358 & ~n_26359;
assign n_26361 = ~n_24900 &  n_26360;
assign n_26362 = ~n_25227 & ~n_25035;
assign n_26363 =  n_23596 &  n_24967;
assign n_26364 = ~n_23821 & ~n_26363;
assign n_26365 = ~n_24760 &  n_26364;
assign n_26366 =  n_26362 &  n_26365;
assign n_26367 =  n_26361 &  n_26366;
assign n_26368 =  n_13104 &  n_24017;
assign n_26369 = ~n_26368 & ~n_14260;
assign n_26370 =  n_23857 &  n_26369;
assign n_26371 =  n_25910 &  n_24967;
assign n_26372 = ~n_26371 & ~n_24970;
assign n_26373 =  n_25510 &  n_25243;
assign n_26374 = ~n_26373 & ~n_24972;
assign n_26375 =  n_26372 &  n_26374;
assign n_26376 =  n_26370 &  n_26375;
assign n_26377 =  n_26367 &  n_26376;
assign n_26378 =  n_26357 &  n_26377;
assign n_26379 =  n_26342 &  n_26378;
assign n_26380 =  n_26275 &  n_26379;
assign n_26381 =  n_26237 &  n_26380;
assign n_26382 =  n_6378 &  n_25263;
assign n_26383 = ~n_23555 & ~n_24773;
assign n_26384 = ~n_26382 &  n_26383;
assign n_26385 = ~n_25518 & ~n_24037;
assign n_26386 = ~x_42 & ~n_26385;
assign n_26387 = ~n_25003 & ~n_26386;
assign n_26388 = ~x_43 & ~n_26387;
assign n_26389 = ~n_26388 &  n_25666;
assign n_26390 =  n_25647 &  n_26389;
assign n_26391 =  n_26384 &  n_26390;
assign n_26392 =  n_25509 &  n_26391;
assign n_26393 =  n_25692 &  n_25267;
assign n_26394 =  n_1038 &  n_20077;
assign n_26395 = ~n_23004 &  n_26394;
assign n_26396 = ~n_26393 & ~n_26395;
assign n_26397 =  n_6876 &  n_356;
assign n_26398 =  n_25682 &  n_26397;
assign n_26399 = ~n_26398 & ~n_25684;
assign n_26400 =  n_26396 &  n_26399;
assign n_26401 =  n_1900 &  n_23876;
assign n_26402 =  n_2880 &  n_3632;
assign n_26403 = ~n_26401 & ~n_26402;
assign n_26404 =  x_43 & ~n_26403;
assign n_26405 = ~n_6881 & ~n_25236;
assign n_26406 =  x_43 & ~n_26405;
assign n_26407 = ~n_26404 & ~n_26406;
assign n_26408 =  n_24574 &  n_26407;
assign n_26409 =  n_764 &  n_25493;
assign n_26410 =  n_24910 &  n_26409;
assign n_26411 =  n_552 &  n_25692;
assign n_26412 =  n_24310 &  n_8053;
assign n_26413 = ~n_26411 & ~n_26412;
assign n_26414 = ~n_26410 &  n_26413;
assign n_26415 =  n_23690 &  n_26414;
assign n_26416 =  n_23769 & ~n_25011;
assign n_26417 = ~n_24671 &  n_26416;
assign n_26418 =  n_26415 &  n_26417;
assign n_26419 =  n_26408 &  n_26418;
assign n_26420 =  n_26195 &  n_11;
assign n_26421 =  n_24752 & ~n_26420;
assign n_26422 =  n_26421 &  n_23831;
assign n_26423 =  n_26419 &  n_26422;
assign n_26424 =  n_26400 &  n_26423;
assign n_26425 =  n_23060 &  n_23061;
assign n_26426 =  n_6379 &  n_155;
assign n_26427 = ~n_26425 & ~n_26426;
assign n_26428 =  n_2094 &  n_25675;
assign n_26429 =  n_23134 &  n_24022;
assign n_26430 =  n_25150 &  n_25210;
assign n_26431 =  n_23692 &  n_24789;
assign n_26432 = ~n_26430 & ~n_26431;
assign n_26433 = ~n_26429 &  n_26432;
assign n_26434 = ~n_26428 &  n_26433;
assign n_26435 =  n_26427 &  n_26434;
assign n_26436 =  n_24806 &  n_23135;
assign n_26437 = ~n_24930 & ~n_26436;
assign n_26438 = ~n_24929 & ~n_23378;
assign n_26439 = ~x_43 &  n_24009;
assign n_26440 = ~n_20597 & ~n_26439;
assign n_26441 =  n_26438 &  n_26440;
assign n_26442 =  n_26437 &  n_26441;
assign n_26443 = ~n_17787 &  n_26442;
assign n_26444 =  n_23174 &  n_25971;
assign n_26445 = ~n_24629 & ~n_26444;
assign n_26446 =  n_351 &  n_18914;
assign n_26447 = ~n_24940 & ~n_26446;
assign n_26448 =  n_26445 &  n_26447;
assign n_26449 =  n_4089 &  n_24306;
assign n_26450 = ~n_24980 & ~n_26449;
assign n_26451 =  n_349 &  n_23642;
assign n_26452 =  n_26450 & ~n_26451;
assign n_26453 =  n_26448 &  n_26452;
assign n_26454 = ~n_24517 &  n_26453;
assign n_26455 =  n_26443 &  n_26454;
assign n_26456 =  n_26435 &  n_26455;
assign n_26457 = ~n_14787 & ~n_20985;
assign n_26458 =  n_24746 &  n_25658;
assign n_26459 =  x_43 &  n_26458;
assign n_26460 = ~n_26459 & ~n_24007;
assign n_26461 = ~n_23377 &  n_26460;
assign n_26462 =  n_26457 &  n_26461;
assign n_26463 =  x_3911 &  n_20401;
assign n_26464 =  n_14 &  n_26463;
assign n_26465 =  n_24889 &  n_26464;
assign n_26466 = ~x_3912 &  n_153;
assign n_26467 =  n_26465 &  n_26466;
assign n_26468 =  x_42 &  n_26008;
assign n_26469 =  x_43 &  n_26468;
assign n_26470 = ~n_26467 & ~n_26469;
assign n_26471 =  n_349 &  n_23467;
assign n_26472 =  n_25091 &  n_23466;
assign n_26473 = ~x_43 &  n_26472;
assign n_26474 = ~x_42 &  n_26473;
assign n_26475 = ~n_26471 & ~n_26474;
assign n_26476 = ~n_25094 &  n_26475;
assign n_26477 =  n_26470 &  n_26476;
assign n_26478 =  n_26462 &  n_26477;
assign n_26479 =  n_23477 & ~n_23508;
assign n_26480 = ~n_23542 & ~n_26479;
assign n_26481 =  n_24314 &  n_3625;
assign n_26482 = ~n_23509 & ~n_26481;
assign n_26483 =  n_25455 & ~n_25486;
assign n_26484 =  n_23010 &  n_24976;
assign n_26485 =  n_15366 &  n_26484;
assign n_26486 =  n_554 &  n_25634;
assign n_26487 = ~n_26485 & ~n_26486;
assign n_26488 = ~n_26483 &  n_26487;
assign n_26489 =  n_26482 &  n_26488;
assign n_26490 =  n_26480 &  n_26489;
assign n_26491 = ~x_43 &  n_24214;
assign n_26492 = ~n_24701 & ~n_26491;
assign n_26493 =  n_26490 &  n_26492;
assign n_26494 =  n_26478 &  n_26493;
assign n_26495 =  n_26456 &  n_26494;
assign n_26496 =  n_26424 &  n_26495;
assign n_26497 =  n_26392 &  n_26496;
assign n_26498 =  n_26381 &  n_26497;
assign n_26499 =  n_25889 &  n_26498;
assign n_26500 = ~n_25846 &  n_26499;
assign n_26501 =  n_22464 &  n_26500;
assign n_26502 = ~n_25845 &  n_26501;
assign n_26503 = ~n_25844 &  n_26502;
assign n_26504 =  n_25717 &  n_26503;
assign n_26505 =  x_42 & ~n_26504;
assign n_26506 = ~x_42 &  n_26504;
assign n_26507 = ~n_26505 & ~n_26506;
assign n_26508 =  n_4089 &  n_24314;
assign n_26509 =  x_556 & ~x_3097;
assign n_26510 = ~x_556 &  x_3097;
assign n_26511 = ~x_557 &  x_3098;
assign n_26512 =  x_557 & ~x_3098;
assign n_26513 = ~x_558 &  x_3099;
assign n_26514 =  x_558 & ~x_3099;
assign n_26515 = ~x_559 &  x_3100;
assign n_26516 =  x_559 & ~x_3100;
assign n_26517 = ~x_560 &  x_3101;
assign n_26518 =  x_560 & ~x_3101;
assign n_26519 = ~x_561 &  x_3102;
assign n_26520 =  x_561 & ~x_3102;
assign n_26521 = ~x_562 &  x_3103;
assign n_26522 =  x_562 & ~x_3103;
assign n_26523 = ~x_563 &  x_3104;
assign n_26524 =  x_563 & ~x_3104;
assign n_26525 = ~x_564 &  x_3105;
assign n_26526 =  x_564 & ~x_3105;
assign n_26527 = ~x_565 &  x_3106;
assign n_26528 =  x_565 & ~x_3106;
assign n_26529 = ~x_566 &  x_3107;
assign n_26530 =  x_566 & ~x_3107;
assign n_26531 = ~x_567 &  x_3108;
assign n_26532 =  x_567 & ~x_3108;
assign n_26533 = ~x_568 &  x_3109;
assign n_26534 =  x_568 & ~x_3109;
assign n_26535 = ~x_569 &  x_3110;
assign n_26536 =  x_569 & ~x_3110;
assign n_26537 = ~x_570 &  x_3111;
assign n_26538 =  x_570 & ~x_3111;
assign n_26539 = ~x_571 &  x_3112;
assign n_26540 =  x_571 & ~x_3112;
assign n_26541 = ~x_572 &  x_3113;
assign n_26542 =  x_572 & ~x_3113;
assign n_26543 = ~x_573 &  x_3114;
assign n_26544 =  x_573 & ~x_3114;
assign n_26545 = ~x_574 &  x_3115;
assign n_26546 =  x_574 & ~x_3115;
assign n_26547 = ~x_575 &  x_3116;
assign n_26548 =  x_575 & ~x_3116;
assign n_26549 = ~x_576 &  x_3117;
assign n_26550 =  x_576 & ~x_3117;
assign n_26551 = ~x_577 &  x_3118;
assign n_26552 =  x_577 & ~x_3118;
assign n_26553 = ~x_578 &  x_3119;
assign n_26554 =  x_578 & ~x_3119;
assign n_26555 = ~x_579 &  x_3120;
assign n_26556 =  x_579 & ~x_3120;
assign n_26557 = ~x_580 &  x_3121;
assign n_26558 =  x_580 & ~x_3121;
assign n_26559 = ~x_581 &  x_3122;
assign n_26560 =  x_581 & ~x_3122;
assign n_26561 = ~x_582 &  x_3123;
assign n_26562 =  x_582 & ~x_3123;
assign n_26563 = ~x_583 &  x_3124;
assign n_26564 =  x_583 & ~x_3124;
assign n_26565 = ~x_584 &  x_3125;
assign n_26566 =  x_584 & ~x_3125;
assign n_26567 = ~x_586 &  x_3127;
assign n_26568 =  x_586 & ~x_3127;
assign n_26569 = ~x_587 &  x_3128;
assign n_26570 = ~n_26568 &  n_26569;
assign n_26571 = ~n_26567 & ~n_26570;
assign n_26572 =  x_585 &  n_26571;
assign n_26573 =  x_3126 & ~n_26572;
assign n_26574 = ~x_585 & ~n_26571;
assign n_26575 = ~n_26573 & ~n_26574;
assign n_26576 = ~n_26566 & ~n_26575;
assign n_26577 = ~n_26565 & ~n_26576;
assign n_26578 = ~n_26564 & ~n_26577;
assign n_26579 = ~n_26563 & ~n_26578;
assign n_26580 = ~n_26562 & ~n_26579;
assign n_26581 = ~n_26561 & ~n_26580;
assign n_26582 = ~n_26560 & ~n_26581;
assign n_26583 = ~n_26559 & ~n_26582;
assign n_26584 = ~n_26558 & ~n_26583;
assign n_26585 = ~n_26557 & ~n_26584;
assign n_26586 = ~n_26556 & ~n_26585;
assign n_26587 = ~n_26555 & ~n_26586;
assign n_26588 = ~n_26554 & ~n_26587;
assign n_26589 = ~n_26553 & ~n_26588;
assign n_26590 = ~n_26552 & ~n_26589;
assign n_26591 = ~n_26551 & ~n_26590;
assign n_26592 = ~n_26550 & ~n_26591;
assign n_26593 = ~n_26549 & ~n_26592;
assign n_26594 = ~n_26548 & ~n_26593;
assign n_26595 = ~n_26547 & ~n_26594;
assign n_26596 = ~n_26546 & ~n_26595;
assign n_26597 = ~n_26545 & ~n_26596;
assign n_26598 = ~n_26544 & ~n_26597;
assign n_26599 = ~n_26543 & ~n_26598;
assign n_26600 = ~n_26542 & ~n_26599;
assign n_26601 = ~n_26541 & ~n_26600;
assign n_26602 = ~n_26540 & ~n_26601;
assign n_26603 = ~n_26539 & ~n_26602;
assign n_26604 = ~n_26538 & ~n_26603;
assign n_26605 = ~n_26537 & ~n_26604;
assign n_26606 = ~n_26536 & ~n_26605;
assign n_26607 = ~n_26535 & ~n_26606;
assign n_26608 = ~n_26534 & ~n_26607;
assign n_26609 = ~n_26533 & ~n_26608;
assign n_26610 = ~n_26532 & ~n_26609;
assign n_26611 = ~n_26531 & ~n_26610;
assign n_26612 = ~n_26530 & ~n_26611;
assign n_26613 = ~n_26529 & ~n_26612;
assign n_26614 = ~n_26528 & ~n_26613;
assign n_26615 = ~n_26527 & ~n_26614;
assign n_26616 = ~n_26526 & ~n_26615;
assign n_26617 = ~n_26525 & ~n_26616;
assign n_26618 = ~n_26524 & ~n_26617;
assign n_26619 = ~n_26523 & ~n_26618;
assign n_26620 = ~n_26522 & ~n_26619;
assign n_26621 = ~n_26521 & ~n_26620;
assign n_26622 = ~n_26520 & ~n_26621;
assign n_26623 = ~n_26519 & ~n_26622;
assign n_26624 = ~n_26518 & ~n_26623;
assign n_26625 = ~n_26517 & ~n_26624;
assign n_26626 = ~n_26516 & ~n_26625;
assign n_26627 = ~n_26515 & ~n_26626;
assign n_26628 = ~n_26514 & ~n_26627;
assign n_26629 = ~n_26513 & ~n_26628;
assign n_26630 = ~n_26512 & ~n_26629;
assign n_26631 = ~n_26511 & ~n_26630;
assign n_26632 = ~n_26510 & ~n_26631;
assign n_26633 = ~n_26509 & ~n_26632;
assign n_26634 =  n_26508 &  n_26633;
assign n_26635 = ~n_26634 & ~n_22465;
assign n_26636 = ~n_22082 &  n_26635;
assign n_26637 =  n_26508 & ~n_26633;
assign n_26638 =  n_21956 &  n_22081;
assign n_26639 =  n_22337 &  n_22462;
assign n_26640 =  n_554 &  n_1897;
assign n_26641 =  n_15917 &  n_26640;
assign n_26642 = ~x_1567 & ~x_1568;
assign n_26643 = ~x_1569 & ~x_1570;
assign n_26644 =  n_26642 &  n_26643;
assign n_26645 = ~x_1563 & ~x_1564;
assign n_26646 = ~x_1565 & ~x_1566;
assign n_26647 =  n_26645 &  n_26646;
assign n_26648 =  n_26644 &  n_26647;
assign n_26649 = ~x_1575 & ~x_1576;
assign n_26650 = ~x_1577 & ~x_1578;
assign n_26651 =  n_26649 &  n_26650;
assign n_26652 = ~x_1571 & ~x_1572;
assign n_26653 = ~x_1573 & ~x_1574;
assign n_26654 =  n_26652 &  n_26653;
assign n_26655 =  n_26651 &  n_26654;
assign n_26656 =  n_26648 &  n_26655;
assign n_26657 = ~x_1551 & ~x_1552;
assign n_26658 = ~x_1553 & ~x_1554;
assign n_26659 =  n_26657 &  n_26658;
assign n_26660 = ~x_1547 & ~x_1548;
assign n_26661 = ~x_1549 & ~x_1550;
assign n_26662 =  n_26660 &  n_26661;
assign n_26663 =  n_26659 &  n_26662;
assign n_26664 = ~x_1559 & ~x_1560;
assign n_26665 = ~x_1561 & ~x_1562;
assign n_26666 =  n_26664 &  n_26665;
assign n_26667 = ~x_1555 & ~x_1556;
assign n_26668 = ~x_1557 & ~x_1558;
assign n_26669 =  n_26667 &  n_26668;
assign n_26670 =  n_26666 &  n_26669;
assign n_26671 =  n_26663 &  n_26670;
assign n_26672 =  n_26656 &  n_26671;
assign n_26673 =  n_26641 & ~n_26672;
assign n_26674 =  n_2684 &  n_23829;
assign n_26675 =  n_26674 & ~n_26672;
assign n_26676 =  n_24785 & ~n_26675;
assign n_26677 = ~n_26673 &  n_26676;
assign n_26678 =  n_26122 &  n_23099;
assign n_26679 = ~n_24582 & ~n_26179;
assign n_26680 = ~n_26678 &  n_26679;
assign n_26681 =  n_26677 &  n_26680;
assign n_26682 = ~n_23060 &  n_23473;
assign n_26683 =  n_24270 &  n_24301;
assign n_26684 =  n_23333 &  n_23364;
assign n_26685 = ~n_26683 & ~n_26684;
assign n_26686 = ~n_26064 &  n_26685;
assign n_26687 = ~n_25337 &  n_26686;
assign n_26688 = ~n_26682 &  n_26687;
assign n_26689 =  n_26688 &  n_23730;
assign n_26690 =  n_26681 &  n_26689;
assign n_26691 =  n_9884 &  n_10867;
assign n_26692 = ~n_25847 & ~n_26691;
assign n_26693 = ~n_25262 &  n_26692;
assign n_26694 = ~n_24777 & ~n_23294;
assign n_26695 =  n_26693 &  n_26694;
assign n_26696 =  x_1705 &  x_1706;
assign n_26697 =  n_23290 & ~n_26696;
assign n_26698 = ~x_1675 & ~n_26697;
assign n_26699 = ~n_26698 &  n_25025;
assign n_26700 =  n_26005 &  n_13866;
assign n_26701 = ~n_26699 & ~n_26700;
assign n_26702 = ~n_23620 &  n_26701;
assign n_26703 =  n_26695 &  n_26702;
assign n_26704 = ~n_24513 & ~n_26300;
assign n_26705 = ~n_26674 & ~n_26641;
assign n_26706 = ~n_26705 &  n_26672;
assign n_26707 = ~n_26706 & ~n_26139;
assign n_26708 =  n_26704 &  n_26707;
assign n_26709 =  n_23329 &  n_357;
assign n_26710 =  n_1175 &  n_23548;
assign n_26711 = ~n_7080 & ~n_26710;
assign n_26712 =  n_23840 &  n_6876;
assign n_26713 = ~n_26013 & ~n_26712;
assign n_26714 =  n_26711 &  n_26713;
assign n_26715 = ~n_26709 &  n_26714;
assign n_26716 =  n_23258 &  n_26715;
assign n_26717 =  n_26708 &  n_26716;
assign n_26718 = ~n_23134 &  n_24022;
assign n_26719 =  n_23329 &  n_14785;
assign n_26720 =  n_23325 &  n_26719;
assign n_26721 = ~n_26718 & ~n_26720;
assign n_26722 =  n_26721 &  n_25678;
assign n_26723 =  n_26717 &  n_26722;
assign n_26724 =  n_26703 &  n_26723;
assign n_26725 =  n_26690 &  n_26724;
assign n_26726 = ~n_26428 &  n_25702;
assign n_26727 =  n_25870 & ~n_23834;
assign n_26728 =  n_23826 &  n_26727;
assign n_26729 =  n_26726 &  n_26728;
assign n_26730 =  n_26725 &  n_26729;
assign n_26731 =  n_25171 & ~n_4284;
assign n_26732 =  n_23329 &  n_23877;
assign n_26733 = ~n_24077 & ~n_26732;
assign n_26734 =  n_26733 &  n_25252;
assign n_26735 =  n_26731 &  n_26734;
assign n_26736 = ~n_26373 & ~n_25207;
assign n_26737 = ~n_24051 & ~n_25986;
assign n_26738 = ~n_25277 &  n_26737;
assign n_26739 =  n_26736 &  n_26738;
assign n_26740 =  n_26735 &  n_26739;
assign n_26741 = ~n_24311 & ~n_24068;
assign n_26742 = ~n_26481 & ~n_19496;
assign n_26743 =  n_26741 &  n_26742;
assign n_26744 = ~x_2863 & ~x_2864;
assign n_26745 = ~x_2865 & ~x_2866;
assign n_26746 =  n_26744 &  n_26745;
assign n_26747 = ~x_2859 & ~x_2860;
assign n_26748 = ~x_2861 & ~x_2862;
assign n_26749 =  n_26747 &  n_26748;
assign n_26750 =  n_26746 &  n_26749;
assign n_26751 = ~x_2871 & ~x_2872;
assign n_26752 = ~x_2873 & ~x_2874;
assign n_26753 =  n_26751 &  n_26752;
assign n_26754 = ~x_2867 & ~x_2868;
assign n_26755 = ~x_2869 & ~x_2870;
assign n_26756 =  n_26754 &  n_26755;
assign n_26757 =  n_26753 &  n_26756;
assign n_26758 =  n_26750 &  n_26757;
assign n_26759 = ~x_2847 & ~x_2848;
assign n_26760 = ~x_2849 & ~x_2850;
assign n_26761 =  n_26759 &  n_26760;
assign n_26762 = ~x_2843 & ~x_2844;
assign n_26763 = ~x_2845 & ~x_2846;
assign n_26764 =  n_26762 &  n_26763;
assign n_26765 =  n_26761 &  n_26764;
assign n_26766 = ~x_2855 & ~x_2856;
assign n_26767 = ~x_2857 & ~x_2858;
assign n_26768 =  n_26766 &  n_26767;
assign n_26769 = ~x_2851 & ~x_2852;
assign n_26770 = ~x_2853 & ~x_2854;
assign n_26771 =  n_26769 &  n_26770;
assign n_26772 =  n_26768 &  n_26771;
assign n_26773 =  n_26765 &  n_26772;
assign n_26774 =  n_26758 &  n_26773;
assign n_26775 =  n_24304 & ~n_26774;
assign n_26776 = ~n_26775 & ~n_1700;
assign n_26777 =  n_26743 &  n_26776;
assign n_26778 =  n_25873 & ~n_23244;
assign n_26779 = ~n_26778 &  n_26437;
assign n_26780 = ~x_3436 & ~x_3437;
assign n_26781 = ~x_3438 & ~x_3439;
assign n_26782 =  n_26780 &  n_26781;
assign n_26783 = ~x_3432 & ~x_3433;
assign n_26784 = ~x_3434 & ~x_3435;
assign n_26785 =  n_26783 &  n_26784;
assign n_26786 =  n_26782 &  n_26785;
assign n_26787 = ~x_3444 & ~x_3445;
assign n_26788 = ~x_3446 & ~x_3447;
assign n_26789 =  n_26787 &  n_26788;
assign n_26790 = ~x_3440 & ~x_3441;
assign n_26791 = ~x_3442 & ~x_3443;
assign n_26792 =  n_26790 &  n_26791;
assign n_26793 =  n_26789 &  n_26792;
assign n_26794 =  n_26786 &  n_26793;
assign n_26795 = ~x_3420 & ~x_3421;
assign n_26796 = ~x_3422 & ~x_3423;
assign n_26797 =  n_26795 &  n_26796;
assign n_26798 = ~x_3416 & ~x_3417;
assign n_26799 = ~x_3418 & ~x_3419;
assign n_26800 =  n_26798 &  n_26799;
assign n_26801 =  n_26797 &  n_26800;
assign n_26802 = ~x_3428 & ~x_3429;
assign n_26803 = ~x_3430 & ~x_3431;
assign n_26804 =  n_26802 &  n_26803;
assign n_26805 = ~x_3424 & ~x_3425;
assign n_26806 = ~x_3426 & ~x_3427;
assign n_26807 =  n_26805 &  n_26806;
assign n_26808 =  n_26804 &  n_26807;
assign n_26809 =  n_26801 &  n_26808;
assign n_26810 =  n_26794 &  n_26809;
assign n_26811 =  n_554 &  n_24073;
assign n_26812 = ~n_26810 &  n_26811;
assign n_26813 = ~n_26147 & ~n_26812;
assign n_26814 =  n_26779 &  n_26813;
assign n_26815 =  n_26777 &  n_26814;
assign n_26816 =  n_26740 &  n_26815;
assign n_26817 =  n_11 &  n_25541;
assign n_26818 = ~n_26817 & ~n_25271;
assign n_26819 = ~n_23841 & ~n_12909;
assign n_26820 =  n_24875 &  n_26819;
assign n_26821 =  n_26818 &  n_26820;
assign n_26822 =  n_20790 &  n_25520;
assign n_26823 =  n_24306 &  n_8818;
assign n_26824 =  n_5645 &  n_3629;
assign n_26825 = ~x_41 & ~n_11;
assign n_26826 = ~n_554 & ~n_26825;
assign n_26827 =  n_24575 &  n_26826;
assign n_26828 = ~n_26824 & ~n_26827;
assign n_26829 = ~n_26823 &  n_26828;
assign n_26830 = ~n_26822 &  n_26829;
assign n_26831 = ~n_8364 & ~n_24520;
assign n_26832 = ~n_25167 & ~n_8358;
assign n_26833 =  n_26831 &  n_26832;
assign n_26834 =  n_26830 &  n_26833;
assign n_26835 =  n_26821 &  n_26834;
assign n_26836 =  n_16495 &  n_25159;
assign n_26837 = ~n_26212 & ~n_26836;
assign n_26838 =  n_26837 &  n_26011;
assign n_26839 =  n_20790 &  n_24969;
assign n_26840 =  n_25912 & ~n_26839;
assign n_26841 = ~n_25216 &  n_26840;
assign n_26842 =  n_26838 &  n_26841;
assign n_26843 =  x_42 &  n_24741;
assign n_26844 =  n_24308 & ~n_26843;
assign n_26845 =  n_9884 &  n_25108;
assign n_26846 = ~n_26162 & ~n_26845;
assign n_26847 =  n_26844 &  n_26846;
assign n_26848 =  n_26842 &  n_26847;
assign n_26849 =  n_26835 &  n_26848;
assign n_26850 =  n_26816 &  n_26849;
assign n_26851 =  n_11 &  n_25533;
assign n_26852 = ~n_26851 &  n_26284;
assign n_26853 = ~x_43 &  n_25641;
assign n_26854 =  n_26287 & ~n_26853;
assign n_26855 =  n_26852 &  n_26854;
assign n_26856 = ~n_24572 &  n_25085;
assign n_26857 =  n_23179 & ~n_23210;
assign n_26858 = ~n_25328 & ~n_26857;
assign n_26859 =  n_26856 &  n_26858;
assign n_26860 =  n_26855 &  n_26859;
assign n_26861 =  n_24119 &  n_24669;
assign n_26862 =  x_42 &  n_26861;
assign n_26863 = ~n_26862 & ~n_25900;
assign n_26864 =  n_24752 &  n_26863;
assign n_26865 =  n_26860 &  n_26864;
assign n_26866 =  n_23942 &  n_13104;
assign n_26867 = ~n_25232 & ~n_26866;
assign n_26868 =  n_26867 & ~n_26180;
assign n_26869 =  n_23771 &  n_23802;
assign n_26870 = ~n_26869 & ~n_25094;
assign n_26871 =  n_26868 &  n_26870;
assign n_26872 = ~n_24005 & ~n_15367;
assign n_26873 = ~n_3145 & ~n_2686;
assign n_26874 =  n_26872 &  n_26873;
assign n_26875 = ~n_26209 & ~n_23247;
assign n_26876 = ~n_26014 & ~n_2488;
assign n_26877 =  n_26875 &  n_26876;
assign n_26878 =  n_26874 &  n_26877;
assign n_26879 =  n_26871 &  n_26878;
assign n_26880 = ~n_26100 & ~n_2097;
assign n_26881 = ~n_24500 &  n_26880;
assign n_26882 = ~n_26071 & ~n_25980;
assign n_26883 =  n_26298 & ~n_23592;
assign n_26884 =  n_26882 & ~n_26883;
assign n_26885 =  n_26881 &  n_26884;
assign n_26886 = ~n_24229 & ~n_25035;
assign n_26887 = ~n_24762 & ~n_23550;
assign n_26888 =  n_26886 &  n_26887;
assign n_26889 =  n_9884 &  n_24017;
assign n_26890 = ~n_26889 & ~n_26156;
assign n_26891 = ~x_4700 & ~x_4701;
assign n_26892 = ~x_4702 & ~x_4703;
assign n_26893 =  n_26891 &  n_26892;
assign n_26894 = ~x_4696 & ~x_4697;
assign n_26895 = ~x_4698 & ~x_4699;
assign n_26896 =  n_26894 &  n_26895;
assign n_26897 =  n_26893 &  n_26896;
assign n_26898 = ~x_4708 & ~x_4709;
assign n_26899 = ~x_4710 & ~x_4711;
assign n_26900 =  n_26898 &  n_26899;
assign n_26901 = ~x_4704 & ~x_4705;
assign n_26902 = ~x_4706 & ~x_4707;
assign n_26903 =  n_26901 &  n_26902;
assign n_26904 =  n_26900 &  n_26903;
assign n_26905 =  n_26897 &  n_26904;
assign n_26906 = ~x_4684 & ~x_4685;
assign n_26907 = ~x_4686 & ~x_4687;
assign n_26908 =  n_26906 &  n_26907;
assign n_26909 = ~x_4680 & ~x_4681;
assign n_26910 = ~x_4682 & ~x_4683;
assign n_26911 =  n_26909 &  n_26910;
assign n_26912 =  n_26908 &  n_26911;
assign n_26913 = ~x_4692 & ~x_4693;
assign n_26914 = ~x_4694 & ~x_4695;
assign n_26915 =  n_26913 &  n_26914;
assign n_26916 = ~x_4688 & ~x_4689;
assign n_26917 = ~x_4690 & ~x_4691;
assign n_26918 =  n_26916 &  n_26917;
assign n_26919 =  n_26915 &  n_26918;
assign n_26920 =  n_26912 &  n_26919;
assign n_26921 =  n_26905 &  n_26920;
assign n_26922 =  n_25937 &  n_26921;
assign n_26923 =  n_26890 & ~n_26922;
assign n_26924 =  n_26888 &  n_26923;
assign n_26925 =  n_26885 &  n_26924;
assign n_26926 =  n_26879 &  n_26925;
assign n_26927 =  n_26865 &  n_26926;
assign n_26928 =  n_26850 &  n_26927;
assign n_26929 =  x_3416 &  n_24739;
assign n_26930 = ~n_26472 & ~n_26929;
assign n_26931 =  n_11 & ~n_26930;
assign n_26932 =  n_13870 &  n_24306;
assign n_26933 = ~n_26932 & ~n_5647;
assign n_26934 = ~n_26931 &  n_26933;
assign n_26935 =  n_15366 &  n_24050;
assign n_26936 = ~n_20078 & ~n_26935;
assign n_26937 =  n_24593 &  n_26936;
assign n_26938 =  x_43 &  n_24074;
assign n_26939 = ~n_10479 & ~n_26938;
assign n_26940 =  n_26937 &  n_26939;
assign n_26941 =  n_26934 &  n_26940;
assign n_26942 =  n_24807 &  n_24838;
assign n_26943 = ~n_26942 & ~n_25419;
assign n_26944 = ~n_26359 & ~n_25219;
assign n_26945 =  n_26943 &  n_26944;
assign n_26946 = ~x_43 &  n_23462;
assign n_26947 =  n_25545 &  n_26946;
assign n_26948 =  x_42 &  n_26947;
assign n_26949 = ~n_24221 & ~n_24319;
assign n_26950 = ~n_26948 &  n_26949;
assign n_26951 =  n_24695 &  n_26950;
assign n_26952 =  n_26945 &  n_26951;
assign n_26953 =  n_26941 &  n_26952;
assign n_26954 =  n_8357 &  n_26354;
assign n_26955 = ~n_1901 & ~n_25011;
assign n_26956 = ~n_25098 & ~n_19500;
assign n_26957 =  n_26955 &  n_26956;
assign n_26958 = ~n_26166 & ~n_24893;
assign n_26959 =  n_26957 &  n_26958;
assign n_26960 =  n_26954 &  n_26959;
assign n_26961 = ~n_26257 & ~n_24065;
assign n_26962 =  n_2682 &  n_7079;
assign n_26963 =  x_588 &  n_11;
assign n_26964 =  n_24936 &  n_26963;
assign n_26965 = ~n_26962 & ~n_26964;
assign n_26966 =  n_26961 &  n_26965;
assign n_26967 =  n_24119 &  n_24067;
assign n_26968 = ~n_25330 & ~n_26967;
assign n_26969 =  n_11 & ~n_26968;
assign n_26970 = ~n_14656 & ~n_24760;
assign n_26971 = ~n_26969 &  n_26970;
assign n_26972 =  n_26966 &  n_26971;
assign n_26973 =  n_26960 &  n_26972;
assign n_26974 =  n_26953 &  n_26973;
assign n_26975 =  n_23329 &  n_2487;
assign n_26976 = ~n_23845 & ~n_26975;
assign n_26977 = ~n_25100 & ~n_25905;
assign n_26978 =  n_26976 &  n_26977;
assign n_26979 = ~n_24231 & ~n_24922;
assign n_26980 =  n_24977 &  n_15366;
assign n_26981 = ~n_26980 & ~n_23943;
assign n_26982 =  n_26979 &  n_26981;
assign n_26983 =  n_26978 &  n_26982;
assign n_26984 = ~n_23053 & ~n_10871;
assign n_26985 = ~n_6878 & ~n_25669;
assign n_26986 =  n_26984 &  n_26985;
assign n_26987 = ~n_14260 & ~n_25245;
assign n_26988 = ~n_25988 & ~n_26171;
assign n_26989 =  n_26987 &  n_26988;
assign n_26990 =  n_26986 &  n_26989;
assign n_26991 =  n_26983 &  n_26990;
assign n_26992 =  n_15366 &  n_10867;
assign n_26993 = ~n_26345 & ~n_26992;
assign n_26994 =  n_6876 &  n_23881;
assign n_26995 = ~n_26368 & ~n_26994;
assign n_26996 =  n_26993 &  n_26995;
assign n_26997 = ~n_25017 & ~n_25151;
assign n_26998 = ~n_24313 & ~n_26020;
assign n_26999 =  n_26997 &  n_26998;
assign n_27000 =  n_26996 &  n_26999;
assign n_27001 =  n_758 &  n_9;
assign n_27002 = ~n_27001 & ~n_20791;
assign n_27003 =  n_6883 & ~n_25952;
assign n_27004 = ~n_25008 & ~n_27003;
assign n_27005 =  n_27002 &  n_27004;
assign n_27006 = ~n_25024 & ~n_25931;
assign n_27007 =  n_13870 &  n_24309;
assign n_27008 = ~n_10 & ~n_27007;
assign n_27009 =  n_27006 &  n_27008;
assign n_27010 =  n_27005 &  n_27009;
assign n_27011 =  n_27000 &  n_27010;
assign n_27012 =  n_11 &  n_25542;
assign n_27013 = ~n_24951 & ~n_27012;
assign n_27014 = ~n_23066 & ~n_17980;
assign n_27015 =  n_27013 &  n_27014;
assign n_27016 =  n_23329 &  n_18914;
assign n_27017 = ~n_27016 & ~n_25105;
assign n_27018 = ~n_25157 & ~n_24961;
assign n_27019 =  n_27017 &  n_27018;
assign n_27020 =  n_27015 &  n_27019;
assign n_27021 =  n_27011 &  n_27020;
assign n_27022 =  n_26991 &  n_27021;
assign n_27023 =  n_9884 &  n_1900;
assign n_27024 = ~n_24573 & ~n_27023;
assign n_27025 =  n_25970 &  n_27024;
assign n_27026 = ~x_43 &  n_6881;
assign n_27027 = ~n_25955 & ~n_27026;
assign n_27028 = ~x_42 &  n_24037;
assign n_27029 = ~n_25638 & ~n_27028;
assign n_27030 =  n_27027 &  n_27029;
assign n_27031 =  n_27025 &  n_27030;
assign n_27032 =  x_42 &  n_24899;
assign n_27033 = ~n_27032 & ~n_25345;
assign n_27034 = ~n_25632 &  n_27033;
assign n_27035 =  n_27031 &  n_27034;
assign n_27036 = ~n_21565 & ~n_23136;
assign n_27037 = ~n_13231 & ~n_21371;
assign n_27038 =  n_27036 &  n_27037;
assign n_27039 = ~n_23541 & ~n_16496;
assign n_27040 =  n_22715 &  n_25993;
assign n_27041 = ~n_24016 & ~n_27040;
assign n_27042 =  n_27039 &  n_27041;
assign n_27043 =  n_27038 &  n_27042;
assign n_27044 =  n_1307 & ~n_25952;
assign n_27045 =  n_24314 &  n_5656;
assign n_27046 = ~n_27044 & ~n_27045;
assign n_27047 =  n_152 &  n_5649;
assign n_27048 = ~n_24682 & ~n_25651;
assign n_27049 = ~n_27047 &  n_27048;
assign n_27050 =  n_27046 &  n_27049;
assign n_27051 = ~n_8362 & ~n_19498;
assign n_27052 =  n_23006 &  n_552;
assign n_27053 = ~n_27052 & ~n_10277;
assign n_27054 = ~n_19494 &  n_27053;
assign n_27055 =  n_27051 &  n_27054;
assign n_27056 =  n_27050 &  n_27055;
assign n_27057 =  n_27043 &  n_27056;
assign n_27058 =  n_27035 &  n_27057;
assign n_27059 =  n_27022 &  n_27058;
assign n_27060 =  n_26974 &  n_27059;
assign n_27061 =  n_26928 &  n_27060;
assign n_27062 = ~n_24041 &  n_25519;
assign n_27063 =  n_11 & ~n_27062;
assign n_27064 =  n_26265 & ~n_27063;
assign n_27065 =  x_4295 &  x_4296;
assign n_27066 =  n_23001 & ~n_27065;
assign n_27067 = ~x_4265 & ~n_27066;
assign n_27068 =  n_25502 & ~n_27067;
assign n_27069 = ~n_27068 &  n_23380;
assign n_27070 =  n_27064 &  n_27069;
assign n_27071 = ~n_23469 & ~n_24994;
assign n_27072 =  n_1037 &  n_16;
assign n_27073 = ~n_10870 & ~n_27072;
assign n_27074 =  n_27071 &  n_27073;
assign n_27075 =  n_5645 &  n_762;
assign n_27076 = ~n_27075 & ~n_25649;
assign n_27077 = ~n_1044 &  n_27076;
assign n_27078 =  n_27074 &  n_27077;
assign n_27079 =  n_2682 &  n_1306;
assign n_27080 =  n_27079 &  n_26698;
assign n_27081 = ~n_27080 &  n_23457;
assign n_27082 =  n_27078 &  n_27081;
assign n_27083 =  n_27070 &  n_27082;
assign n_27084 =  n_23613 &  n_23013;
assign n_27085 = ~n_23627 & ~n_27084;
assign n_27086 =  n_22940 &  n_25689;
assign n_27087 =  n_27085 & ~n_27086;
assign n_27088 =  n_27083 &  n_27087;
assign n_27089 = ~n_24987 & ~n_25625;
assign n_27090 = ~n_24230 & ~n_24939;
assign n_27091 = ~n_14261 &  n_27090;
assign n_27092 =  n_27089 &  n_27091;
assign n_27093 =  n_27092 &  n_25673;
assign n_27094 =  n_26032 & ~n_26063;
assign n_27095 = ~n_26459 & ~n_26155;
assign n_27096 = ~n_27094 &  n_27095;
assign n_27097 = ~n_26485 & ~n_23983;
assign n_27098 =  n_27096 &  n_27097;
assign n_27099 =  n_27093 &  n_27098;
assign n_27100 = ~n_26114 & ~n_25501;
assign n_27101 =  n_26199 &  n_27100;
assign n_27102 =  n_27067 &  n_25907;
assign n_27103 =  n_27101 & ~n_27102;
assign n_27104 =  n_25387 & ~n_25418;
assign n_27105 = ~n_23509 & ~n_25455;
assign n_27106 = ~n_27104 &  n_27105;
assign n_27107 = ~n_24801 &  n_27106;
assign n_27108 =  n_27103 &  n_27107;
assign n_27109 =  n_27099 &  n_27108;
assign n_27110 = ~n_26231 & ~n_25290;
assign n_27111 =  x_42 &  n_25213;
assign n_27112 = ~n_25892 &  n_26216;
assign n_27113 = ~n_26431 &  n_27112;
assign n_27114 = ~n_27111 &  n_27113;
assign n_27115 =  n_27110 &  n_27114;
assign n_27116 =  n_11 &  n_25546;
assign n_27117 = ~n_25918 & ~n_27116;
assign n_27118 = ~n_26474 &  n_27117;
assign n_27119 = ~n_24787 & ~n_25951;
assign n_27120 =  n_27118 &  n_27119;
assign n_27121 =  n_27115 &  n_27120;
assign n_27122 =  n_8344 &  n_6182;
assign n_27123 = ~n_27122 & ~n_6380;
assign n_27124 = ~x_43 &  n_24019;
assign n_27125 = ~n_25998 & ~n_27124;
assign n_27126 =  n_27123 &  n_27125;
assign n_27127 =  n_26457 &  n_27126;
assign n_27128 =  n_23879 &  n_26153;
assign n_27129 = ~n_25871 & ~n_27128;
assign n_27130 = ~n_25982 & ~n_25332;
assign n_27131 =  n_26810 &  n_26811;
assign n_27132 = ~n_24266 &  n_24267;
assign n_27133 = ~n_27131 & ~n_27132;
assign n_27134 =  n_27130 &  n_27133;
assign n_27135 =  n_27129 &  n_27134;
assign n_27136 =  n_27127 &  n_27135;
assign n_27137 =  n_27121 &  n_27136;
assign n_27138 =  n_27109 &  n_27137;
assign n_27139 =  n_27088 &  n_27138;
assign n_27140 =  n_27061 &  n_27139;
assign n_27141 =  n_24043 &  n_8353;
assign n_27142 = ~n_25911 & ~n_27141;
assign n_27143 = ~n_25643 & ~n_23544;
assign n_27144 =  n_27142 &  n_27143;
assign n_27145 = ~n_26430 &  n_27144;
assign n_27146 =  n_26197 &  n_27145;
assign n_27147 = ~n_24681 & ~n_25555;
assign n_27148 =  n_27146 &  n_27147;
assign n_27149 =  n_24430 &  n_27148;
assign n_27150 =  n_23253 &  n_6379;
assign n_27151 = ~n_23047 &  n_27150;
assign n_27152 =  n_23006 &  n_355;
assign n_27153 =  n_23555 &  n_23556;
assign n_27154 = ~n_27152 & ~n_27153;
assign n_27155 = ~n_27151 &  n_27154;
assign n_27156 = ~n_23640 &  n_27155;
assign n_27157 =  n_27149 &  n_27156;
assign n_27158 =  n_11 &  n_26113;
assign n_27159 = ~n_27158 & ~n_26393;
assign n_27160 =  n_24630 &  n_25691;
assign n_27161 = ~n_27160 & ~n_25269;
assign n_27162 =  n_27159 &  n_27161;
assign n_27163 = ~n_18302 &  n_26427;
assign n_27164 = ~n_26382 &  n_27163;
assign n_27165 =  n_27162 &  n_27164;
assign n_27166 =  n_27157 &  n_27165;
assign n_27167 =  n_25661 &  n_24634;
assign n_27168 = ~n_24668 &  n_27167;
assign n_27169 =  x_42 &  n_24516;
assign n_27170 =  n_26414 & ~n_27169;
assign n_27171 =  x_42 &  n_24670;
assign n_27172 = ~n_25664 & ~n_27171;
assign n_27173 =  n_27170 &  n_27172;
assign n_27174 =  n_27168 &  n_27173;
assign n_27175 = ~x_43 &  n_25511;
assign n_27176 =  x_42 &  n_27175;
assign n_27177 = ~n_25939 & ~n_25344;
assign n_27178 =  n_27177 & ~n_26027;
assign n_27179 = ~n_27176 &  n_27178;
assign n_27180 =  n_1173 &  n_24310;
assign n_27181 = ~n_23057 &  n_27180;
assign n_27182 = ~n_27181 & ~n_24698;
assign n_27183 =  n_27179 &  n_27182;
assign n_27184 =  n_27174 &  n_27183;
assign n_27185 = ~n_23244 &  n_23245;
assign n_27186 = ~n_27185 & ~n_24021;
assign n_27187 =  n_26470 &  n_27186;
assign n_27188 =  n_25921 &  n_1502;
assign n_27189 = ~x_2511 & ~x_2512;
assign n_27190 = ~x_2513 & ~x_2514;
assign n_27191 =  n_27189 &  n_27190;
assign n_27192 = ~x_2507 & ~x_2508;
assign n_27193 = ~x_2509 & ~x_2510;
assign n_27194 =  n_27192 &  n_27193;
assign n_27195 =  n_27191 &  n_27194;
assign n_27196 = ~x_2519 & ~x_2520;
assign n_27197 = ~x_2521 & ~x_2522;
assign n_27198 =  n_27196 &  n_27197;
assign n_27199 = ~x_2515 & ~x_2516;
assign n_27200 = ~x_2517 & ~x_2518;
assign n_27201 =  n_27199 &  n_27200;
assign n_27202 =  n_27198 &  n_27201;
assign n_27203 =  n_27195 &  n_27202;
assign n_27204 = ~x_2495 & ~x_2496;
assign n_27205 = ~x_2497 & ~x_2498;
assign n_27206 =  n_27204 &  n_27205;
assign n_27207 = ~x_2491 & ~x_2492;
assign n_27208 = ~x_2493 & ~x_2494;
assign n_27209 =  n_27207 &  n_27208;
assign n_27210 =  n_27206 &  n_27209;
assign n_27211 = ~x_2503 & ~x_2504;
assign n_27212 = ~x_2505 & ~x_2506;
assign n_27213 =  n_27211 &  n_27212;
assign n_27214 = ~x_2499 & ~x_2500;
assign n_27215 = ~x_2501 & ~x_2502;
assign n_27216 =  n_27214 &  n_27215;
assign n_27217 =  n_27213 &  n_27216;
assign n_27218 =  n_27210 &  n_27217;
assign n_27219 =  n_27203 &  n_27218;
assign n_27220 =  n_27188 &  n_27219;
assign n_27221 = ~n_24512 & ~n_27220;
assign n_27222 = ~n_24949 & ~n_21564;
assign n_27223 =  n_757 & ~n_27222;
assign n_27224 = ~n_27223 & ~n_25953;
assign n_27225 =  n_27221 &  n_27224;
assign n_27226 =  n_27187 &  n_27225;
assign n_27227 = ~n_23608 & ~n_23887;
assign n_27228 = ~n_23997 & ~n_16689;
assign n_27229 =  n_27227 &  n_27228;
assign n_27230 =  n_5645 &  n_24960;
assign n_27231 = ~n_24839 & ~n_27230;
assign n_27232 =  n_27229 &  n_27231;
assign n_27233 = ~x_3181 & ~x_3182;
assign n_27234 = ~x_3183 & ~x_3184;
assign n_27235 =  n_27233 &  n_27234;
assign n_27236 = ~x_3177 & ~x_3178;
assign n_27237 = ~x_3179 & ~x_3180;
assign n_27238 =  n_27236 &  n_27237;
assign n_27239 =  n_27235 &  n_27238;
assign n_27240 = ~x_3189 & ~x_3190;
assign n_27241 = ~x_3191 & ~x_3192;
assign n_27242 =  n_27240 &  n_27241;
assign n_27243 = ~x_3185 & ~x_3186;
assign n_27244 = ~x_3187 & ~x_3188;
assign n_27245 =  n_27243 &  n_27244;
assign n_27246 =  n_27242 &  n_27245;
assign n_27247 =  n_27239 &  n_27246;
assign n_27248 = ~x_3165 & ~x_3166;
assign n_27249 = ~x_3167 & ~x_3168;
assign n_27250 =  n_27248 &  n_27249;
assign n_27251 = ~x_3161 & ~x_3162;
assign n_27252 = ~x_3163 & ~x_3164;
assign n_27253 =  n_27251 &  n_27252;
assign n_27254 =  n_27250 &  n_27253;
assign n_27255 = ~x_3173 & ~x_3174;
assign n_27256 = ~x_3175 & ~x_3176;
assign n_27257 =  n_27255 &  n_27256;
assign n_27258 = ~x_3169 & ~x_3170;
assign n_27259 = ~x_3171 & ~x_3172;
assign n_27260 =  n_27258 &  n_27259;
assign n_27261 =  n_27257 &  n_27260;
assign n_27262 =  n_27254 &  n_27261;
assign n_27263 =  n_27247 &  n_27262;
assign n_27264 =  n_24954 &  n_27263;
assign n_27265 = ~n_26205 & ~n_27264;
assign n_27266 =  n_23561 & ~n_23592;
assign n_27267 =  n_27265 & ~n_27266;
assign n_27268 =  n_27232 &  n_27267;
assign n_27269 =  n_27226 &  n_27268;
assign n_27270 = ~n_25922 & ~n_26164;
assign n_27271 = ~n_6876 & ~n_23135;
assign n_27272 =  n_757 & ~n_27271;
assign n_27273 =  x_41 &  x_43;
assign n_27274 =  n_2881 &  n_27273;
assign n_27275 = ~n_27274 & ~n_26093;
assign n_27276 = ~n_27272 &  n_27275;
assign n_27277 =  n_27270 &  n_27276;
assign n_27278 = ~x_41 &  n_8049;
assign n_27279 =  x_42 &  n_27278;
assign n_27280 =  n_25384 & ~n_27279;
assign n_27281 =  n_27277 &  n_27280;
assign n_27282 = ~x_43 &  n_23005;
assign n_27283 =  n_24748 &  n_27282;
assign n_27284 =  x_42 &  n_27283;
assign n_27285 = ~n_27284 & ~n_26269;
assign n_27286 =  n_25877 &  n_27285;
assign n_27287 =  n_26333 & ~n_24563;
assign n_27288 = ~n_24210 & ~n_23992;
assign n_27289 = ~n_27287 &  n_27288;
assign n_27290 =  n_21954 &  n_24269;
assign n_27291 = ~x_320 & ~x_321;
assign n_27292 = ~x_322 & ~x_323;
assign n_27293 =  n_27291 &  n_27292;
assign n_27294 = ~x_316 & ~x_317;
assign n_27295 = ~x_318 & ~x_319;
assign n_27296 =  n_27294 &  n_27295;
assign n_27297 =  n_27293 &  n_27296;
assign n_27298 = ~x_328 & ~x_329;
assign n_27299 = ~x_330 & ~x_331;
assign n_27300 =  n_27298 &  n_27299;
assign n_27301 = ~x_324 & ~x_325;
assign n_27302 = ~x_326 & ~x_327;
assign n_27303 =  n_27301 &  n_27302;
assign n_27304 =  n_27300 &  n_27303;
assign n_27305 =  n_27297 &  n_27304;
assign n_27306 = ~x_304 & ~x_305;
assign n_27307 = ~x_306 & ~x_307;
assign n_27308 =  n_27306 &  n_27307;
assign n_27309 = ~x_300 & ~x_301;
assign n_27310 = ~x_302 & ~x_303;
assign n_27311 =  n_27309 &  n_27310;
assign n_27312 =  n_27308 &  n_27311;
assign n_27313 = ~x_312 & ~x_313;
assign n_27314 = ~x_314 & ~x_315;
assign n_27315 =  n_27313 &  n_27314;
assign n_27316 = ~x_308 & ~x_309;
assign n_27317 = ~x_310 & ~x_311;
assign n_27318 =  n_27316 &  n_27317;
assign n_27319 =  n_27315 &  n_27318;
assign n_27320 =  n_27312 &  n_27319;
assign n_27321 =  n_27305 &  n_27320;
assign n_27322 =  n_27290 & ~n_27321;
assign n_27323 = ~n_24201 & ~n_8366;
assign n_27324 = ~n_27322 &  n_27323;
assign n_27325 =  n_27289 &  n_27324;
assign n_27326 =  n_27286 &  n_27325;
assign n_27327 =  n_27281 &  n_27326;
assign n_27328 =  n_27269 &  n_27327;
assign n_27329 =  n_27184 &  n_27328;
assign n_27330 =  n_349 &  n_24211;
assign n_27331 = ~x_43 &  n_25512;
assign n_27332 =  x_42 &  n_27331;
assign n_27333 = ~n_27330 & ~n_27332;
assign n_27334 = ~n_24911 & ~n_23260;
assign n_27335 =  n_27333 &  n_27334;
assign n_27336 =  n_23951 & ~n_23982;
assign n_27337 = ~n_4287 & ~n_4090;
assign n_27338 =  n_11 &  n_25081;
assign n_27339 = ~n_16110 & ~n_27338;
assign n_27340 =  n_27337 &  n_27339;
assign n_27341 = ~n_27336 &  n_27340;
assign n_27342 =  n_27341 &  n_23626;
assign n_27343 =  n_27335 &  n_27342;
assign n_27344 =  n_23678 &  n_23679;
assign n_27345 = ~n_27344 & ~n_24779;
assign n_27346 = ~n_23008 &  n_27345;
assign n_27347 = ~n_23630 &  n_23631;
assign n_27348 = ~n_27347 & ~n_26398;
assign n_27349 =  n_27346 &  n_27348;
assign n_27350 =  n_27343 &  n_27349;
assign n_27351 =  n_27329 &  n_27350;
assign n_27352 =  n_27166 &  n_27351;
assign n_27353 =  n_27140 &  n_27352;
assign n_27354 =  n_26730 &  n_27353;
assign n_27355 = ~n_22336 &  n_27354;
assign n_27356 = ~n_26639 &  n_27355;
assign n_27357 = ~n_26638 &  n_27356;
assign n_27358 = ~n_26637 &  n_27357;
assign n_27359 =  n_26636 &  n_27358;
assign n_27360 =  x_41 & ~n_27359;
assign n_27361 = ~x_41 &  n_27359;
assign n_27362 = ~n_27360 & ~n_27361;
assign n_27363 =  n_22210 &  n_22335;
assign n_27364 = ~x_1262 &  x_1294;
assign n_27365 =  x_1263 & ~x_1295;
assign n_27366 = ~x_1263 &  x_1295;
assign n_27367 =  x_1264 & ~x_1296;
assign n_27368 = ~x_1264 &  x_1296;
assign n_27369 =  x_1265 & ~x_1297;
assign n_27370 = ~x_1265 &  x_1297;
assign n_27371 =  x_1266 & ~x_1298;
assign n_27372 = ~x_1266 &  x_1298;
assign n_27373 =  x_1267 & ~x_1299;
assign n_27374 = ~x_1267 &  x_1299;
assign n_27375 =  x_1268 & ~x_1300;
assign n_27376 = ~x_1268 &  x_1300;
assign n_27377 =  x_1269 & ~x_1301;
assign n_27378 = ~x_1269 &  x_1301;
assign n_27379 =  x_1270 & ~x_1302;
assign n_27380 = ~x_1270 &  x_1302;
assign n_27381 =  x_1271 & ~x_1303;
assign n_27382 = ~x_1271 &  x_1303;
assign n_27383 =  x_1272 & ~x_1304;
assign n_27384 = ~x_1272 &  x_1304;
assign n_27385 =  x_1273 & ~x_1305;
assign n_27386 = ~x_1273 &  x_1305;
assign n_27387 =  x_1274 & ~x_1306;
assign n_27388 = ~x_1274 &  x_1306;
assign n_27389 =  x_1275 & ~x_1307;
assign n_27390 = ~x_1275 &  x_1307;
assign n_27391 =  x_1276 & ~x_1308;
assign n_27392 = ~x_1276 &  x_1308;
assign n_27393 =  x_1277 & ~x_1309;
assign n_27394 = ~x_1277 &  x_1309;
assign n_27395 =  x_1278 & ~x_1310;
assign n_27396 = ~x_1278 &  x_1310;
assign n_27397 =  x_1279 & ~x_1311;
assign n_27398 = ~x_1279 &  x_1311;
assign n_27399 =  x_1280 & ~x_1312;
assign n_27400 = ~x_1280 &  x_1312;
assign n_27401 =  x_1281 & ~x_1313;
assign n_27402 = ~x_1281 &  x_1313;
assign n_27403 =  x_1282 & ~x_1314;
assign n_27404 = ~x_1282 &  x_1314;
assign n_27405 =  x_1283 & ~x_1315;
assign n_27406 = ~x_1283 &  x_1315;
assign n_27407 =  x_1284 & ~x_1316;
assign n_27408 = ~x_1284 &  x_1316;
assign n_27409 =  x_1285 & ~x_1317;
assign n_27410 = ~x_1285 &  x_1317;
assign n_27411 =  x_1286 & ~x_1318;
assign n_27412 = ~x_1286 &  x_1318;
assign n_27413 =  x_1287 & ~x_1319;
assign n_27414 = ~x_1287 &  x_1319;
assign n_27415 =  x_1289 & ~x_1321;
assign n_27416 = ~x_1289 &  x_1321;
assign n_27417 =  x_1290 & ~x_1322;
assign n_27418 = ~n_27416 &  n_27417;
assign n_27419 = ~n_27415 & ~n_27418;
assign n_27420 =  x_1320 &  n_27419;
assign n_27421 =  x_1288 & ~n_27420;
assign n_27422 = ~x_1320 & ~n_27419;
assign n_27423 = ~n_27421 & ~n_27422;
assign n_27424 = ~n_27414 & ~n_27423;
assign n_27425 = ~n_27413 & ~n_27424;
assign n_27426 = ~n_27412 & ~n_27425;
assign n_27427 = ~n_27411 & ~n_27426;
assign n_27428 = ~n_27410 & ~n_27427;
assign n_27429 = ~n_27409 & ~n_27428;
assign n_27430 = ~n_27408 & ~n_27429;
assign n_27431 = ~n_27407 & ~n_27430;
assign n_27432 = ~n_27406 & ~n_27431;
assign n_27433 = ~n_27405 & ~n_27432;
assign n_27434 = ~n_27404 & ~n_27433;
assign n_27435 = ~n_27403 & ~n_27434;
assign n_27436 = ~n_27402 & ~n_27435;
assign n_27437 = ~n_27401 & ~n_27436;
assign n_27438 = ~n_27400 & ~n_27437;
assign n_27439 = ~n_27399 & ~n_27438;
assign n_27440 = ~n_27398 & ~n_27439;
assign n_27441 = ~n_27397 & ~n_27440;
assign n_27442 = ~n_27396 & ~n_27441;
assign n_27443 = ~n_27395 & ~n_27442;
assign n_27444 = ~n_27394 & ~n_27443;
assign n_27445 = ~n_27393 & ~n_27444;
assign n_27446 = ~n_27392 & ~n_27445;
assign n_27447 = ~n_27391 & ~n_27446;
assign n_27448 = ~n_27390 & ~n_27447;
assign n_27449 = ~n_27389 & ~n_27448;
assign n_27450 = ~n_27388 & ~n_27449;
assign n_27451 = ~n_27387 & ~n_27450;
assign n_27452 = ~n_27386 & ~n_27451;
assign n_27453 = ~n_27385 & ~n_27452;
assign n_27454 = ~n_27384 & ~n_27453;
assign n_27455 = ~n_27383 & ~n_27454;
assign n_27456 = ~n_27382 & ~n_27455;
assign n_27457 = ~n_27381 & ~n_27456;
assign n_27458 = ~n_27380 & ~n_27457;
assign n_27459 = ~n_27379 & ~n_27458;
assign n_27460 = ~n_27378 & ~n_27459;
assign n_27461 = ~n_27377 & ~n_27460;
assign n_27462 = ~n_27376 & ~n_27461;
assign n_27463 = ~n_27375 & ~n_27462;
assign n_27464 = ~n_27374 & ~n_27463;
assign n_27465 = ~n_27373 & ~n_27464;
assign n_27466 = ~n_27372 & ~n_27465;
assign n_27467 = ~n_27371 & ~n_27466;
assign n_27468 = ~n_27370 & ~n_27467;
assign n_27469 = ~n_27369 & ~n_27468;
assign n_27470 = ~n_27368 & ~n_27469;
assign n_27471 = ~n_27367 & ~n_27470;
assign n_27472 = ~n_27366 & ~n_27471;
assign n_27473 = ~n_27365 & ~n_27472;
assign n_27474 = ~n_27364 & ~n_27473;
assign n_27475 =  x_1262 & ~x_1294;
assign n_27476 =  x_1261 & ~x_1293;
assign n_27477 = ~n_27475 & ~n_27476;
assign n_27478 = ~n_27474 &  n_27477;
assign n_27479 = ~x_1260 &  x_1292;
assign n_27480 = ~x_1261 &  x_1293;
assign n_27481 = ~n_27479 & ~n_27480;
assign n_27482 = ~n_27478 &  n_27481;
assign n_27483 =  x_1260 & ~x_1292;
assign n_27484 = ~x_1259 &  x_1291;
assign n_27485 = ~n_27483 & ~n_27484;
assign n_27486 = ~n_27482 &  n_27485;
assign n_27487 =  n_23554 &  n_3615;
assign n_27488 =  x_1259 & ~x_1291;
assign n_27489 =  n_27487 & ~n_27488;
assign n_27490 = ~n_27486 &  n_27489;
assign n_27491 =  n_22721 &  n_22938;
assign n_27492 =  n_6378 &  n_23639;
assign n_27493 =  n_1502 & ~n_24626;
assign n_27494 =  n_5652 &  n_27493;
assign n_27495 = ~n_26014 & ~n_25292;
assign n_27496 = ~n_24065 &  n_27495;
assign n_27497 = ~n_27494 &  n_27496;
assign n_27498 =  n_26676 &  n_27497;
assign n_27499 = ~n_27492 &  n_27498;
assign n_27500 =  n_26680 &  n_27499;
assign n_27501 =  n_24015 &  n_22972;
assign n_27502 =  n_23057 &  n_27180;
assign n_27503 = ~n_26425 & ~n_27502;
assign n_27504 = ~n_27086 &  n_27503;
assign n_27505 = ~n_27501 &  n_27504;
assign n_27506 = ~x_2543 & ~x_2544;
assign n_27507 = ~x_2545 & ~x_2546;
assign n_27508 =  n_27506 &  n_27507;
assign n_27509 = ~x_2539 & ~x_2540;
assign n_27510 = ~x_2541 & ~x_2542;
assign n_27511 =  n_27509 &  n_27510;
assign n_27512 =  n_27508 &  n_27511;
assign n_27513 = ~x_2551 & ~x_2552;
assign n_27514 = ~x_2553 & ~x_2554;
assign n_27515 =  n_27513 &  n_27514;
assign n_27516 = ~x_2547 & ~x_2548;
assign n_27517 = ~x_2549 & ~x_2550;
assign n_27518 =  n_27516 &  n_27517;
assign n_27519 =  n_27515 &  n_27518;
assign n_27520 =  n_27512 &  n_27519;
assign n_27521 = ~x_2527 & ~x_2528;
assign n_27522 = ~x_2529 & ~x_2530;
assign n_27523 =  n_27521 &  n_27522;
assign n_27524 = ~x_2523 & ~x_2524;
assign n_27525 = ~x_2525 & ~x_2526;
assign n_27526 =  n_27524 &  n_27525;
assign n_27527 =  n_27523 &  n_27526;
assign n_27528 = ~x_2535 & ~x_2536;
assign n_27529 = ~x_2537 & ~x_2538;
assign n_27530 =  n_27528 &  n_27529;
assign n_27531 = ~x_2531 & ~x_2532;
assign n_27532 = ~x_2533 & ~x_2534;
assign n_27533 =  n_27531 &  n_27532;
assign n_27534 =  n_27530 &  n_27533;
assign n_27535 =  n_27527 &  n_27534;
assign n_27536 =  n_27520 &  n_27535;
assign n_27537 =  n_24949 & ~n_27536;
assign n_27538 = ~x_1663 & ~x_1664;
assign n_27539 = ~x_1665 & ~x_1666;
assign n_27540 =  n_27538 &  n_27539;
assign n_27541 = ~x_1659 & ~x_1660;
assign n_27542 = ~x_1661 & ~x_1662;
assign n_27543 =  n_27541 &  n_27542;
assign n_27544 =  n_27540 &  n_27543;
assign n_27545 = ~x_1671 & ~x_1672;
assign n_27546 = ~x_1673 & ~x_1674;
assign n_27547 =  n_27545 &  n_27546;
assign n_27548 = ~x_1667 & ~x_1668;
assign n_27549 = ~x_1669 & ~x_1670;
assign n_27550 =  n_27548 &  n_27549;
assign n_27551 =  n_27547 &  n_27550;
assign n_27552 =  n_27544 &  n_27551;
assign n_27553 = ~x_1647 & ~x_1648;
assign n_27554 = ~x_1649 & ~x_1650;
assign n_27555 =  n_27553 &  n_27554;
assign n_27556 = ~x_1643 & ~x_1644;
assign n_27557 = ~x_1645 & ~x_1646;
assign n_27558 =  n_27556 &  n_27557;
assign n_27559 =  n_27555 &  n_27558;
assign n_27560 = ~x_1655 & ~x_1656;
assign n_27561 = ~x_1657 & ~x_1658;
assign n_27562 =  n_27560 &  n_27561;
assign n_27563 = ~x_1651 & ~x_1652;
assign n_27564 = ~x_1653 & ~x_1654;
assign n_27565 =  n_27563 &  n_27564;
assign n_27566 =  n_27562 &  n_27565;
assign n_27567 =  n_27559 &  n_27566;
assign n_27568 =  n_27552 &  n_27567;
assign n_27569 =  n_4089 & ~n_27568;
assign n_27570 = ~n_27537 & ~n_27569;
assign n_27571 = ~n_24667 &  n_27570;
assign n_27572 =  n_10276 & ~n_27571;
assign n_27573 =  n_24840 &  n_24871;
assign n_27574 = ~n_26007 & ~n_27573;
assign n_27575 = ~n_27266 &  n_27574;
assign n_27576 = ~n_27572 &  n_27575;
assign n_27577 =  n_27576 &  n_25270;
assign n_27578 =  n_26688 &  n_27577;
assign n_27579 =  n_27505 &  n_27578;
assign n_27580 =  n_27500 &  n_27579;
assign n_27581 =  n_555 &  n_24114;
assign n_27582 =  n_11 &  n_25544;
assign n_27583 = ~n_27581 & ~n_27582;
assign n_27584 =  n_24968 &  n_24910;
assign n_27585 = ~x_42 &  n_25081;
assign n_27586 = ~n_27585 &  n_26282;
assign n_27587 = ~n_27584 &  n_27586;
assign n_27588 =  n_27583 &  n_27587;
assign n_27589 =  n_13104 &  n_23820;
assign n_27590 = ~n_27589 & ~n_18495;
assign n_27591 =  n_27590 & ~n_26491;
assign n_27592 =  n_27588 &  n_27591;
assign n_27593 =  x_42 &  n_25093;
assign n_27594 = ~n_27593 & ~n_26469;
assign n_27595 =  n_11 &  n_24026;
assign n_27596 = ~n_26932 & ~n_27595;
assign n_27597 =  n_27596 & ~n_12293;
assign n_27598 =  n_27594 &  n_27597;
assign n_27599 =  n_26270 & ~n_24564;
assign n_27600 = ~n_24972 & ~n_26010;
assign n_27601 = ~n_24689 & ~n_25035;
assign n_27602 =  n_27600 &  n_27601;
assign n_27603 =  n_27599 &  n_27602;
assign n_27604 =  n_27598 &  n_27603;
assign n_27605 =  n_26882 & ~n_25079;
assign n_27606 =  n_25937 & ~n_26921;
assign n_27607 = ~n_27606 & ~n_26326;
assign n_27608 =  n_27605 &  n_27607;
assign n_27609 = ~n_16882 & ~n_558;
assign n_27610 =  n_27609 & ~n_26883;
assign n_27611 =  n_24595 & ~n_24626;
assign n_27612 = ~n_24570 & ~n_20596;
assign n_27613 =  n_555 & ~n_27612;
assign n_27614 = ~n_27611 & ~n_27613;
assign n_27615 =  n_27610 &  n_27614;
assign n_27616 =  n_27608 &  n_27615;
assign n_27617 =  n_27604 &  n_27616;
assign n_27618 =  n_27592 &  n_27617;
assign n_27619 =  n_351 &  n_26484;
assign n_27620 = ~x_927 & ~x_928;
assign n_27621 = ~x_929 & ~x_930;
assign n_27622 =  n_27620 &  n_27621;
assign n_27623 = ~x_923 & ~x_924;
assign n_27624 = ~x_925 & ~x_926;
assign n_27625 =  n_27623 &  n_27624;
assign n_27626 =  n_27622 &  n_27625;
assign n_27627 = ~x_935 & ~x_936;
assign n_27628 = ~x_937 & ~x_938;
assign n_27629 =  n_27627 &  n_27628;
assign n_27630 = ~x_931 & ~x_932;
assign n_27631 = ~x_933 & ~x_934;
assign n_27632 =  n_27630 &  n_27631;
assign n_27633 =  n_27629 &  n_27632;
assign n_27634 =  n_27626 &  n_27633;
assign n_27635 = ~x_911 & ~x_912;
assign n_27636 = ~x_913 & ~x_914;
assign n_27637 =  n_27635 &  n_27636;
assign n_27638 = ~x_907 & ~x_908;
assign n_27639 = ~x_909 & ~x_910;
assign n_27640 =  n_27638 &  n_27639;
assign n_27641 =  n_27637 &  n_27640;
assign n_27642 = ~x_919 & ~x_920;
assign n_27643 = ~x_921 & ~x_922;
assign n_27644 =  n_27642 &  n_27643;
assign n_27645 = ~x_915 & ~x_916;
assign n_27646 = ~x_917 & ~x_918;
assign n_27647 =  n_27645 &  n_27646;
assign n_27648 =  n_27644 &  n_27647;
assign n_27649 =  n_27641 &  n_27648;
assign n_27650 =  n_27634 &  n_27649;
assign n_27651 =  n_24199 &  n_27650;
assign n_27652 = ~n_27619 & ~n_27651;
assign n_27653 = ~n_27067 &  n_25907;
assign n_27654 =  n_27652 & ~n_27653;
assign n_27655 =  x_43 &  n_5983;
assign n_27656 = ~n_26931 & ~n_27655;
assign n_27657 = ~n_26074 & ~n_27336;
assign n_27658 =  n_27656 &  n_27657;
assign n_27659 =  n_27654 &  n_27658;
assign n_27660 = ~n_26184 & ~n_25151;
assign n_27661 = ~n_25503 &  n_27660;
assign n_27662 =  n_24934 &  n_26120;
assign n_27663 =  n_27661 &  n_27662;
assign n_27664 = ~n_24681 &  n_27663;
assign n_27665 =  n_554 &  n_24960;
assign n_27666 = ~n_26162 & ~n_27665;
assign n_27667 =  n_11 &  n_25537;
assign n_27668 = ~n_24978 & ~n_26980;
assign n_27669 = ~n_27667 &  n_27668;
assign n_27670 =  n_27666 &  n_27669;
assign n_27671 =  n_27670 & ~n_27181;
assign n_27672 =  n_27664 &  n_27671;
assign n_27673 =  n_27659 &  n_27672;
assign n_27674 =  n_27618 &  n_27673;
assign n_27675 = ~n_24951 & ~n_24124;
assign n_27676 = ~n_23841 & ~n_23992;
assign n_27677 =  n_27675 &  n_27676;
assign n_27678 = ~n_26100 & ~n_2292;
assign n_27679 =  n_25517 &  n_24910;
assign n_27680 = ~n_27679 & ~n_26286;
assign n_27681 =  n_27678 &  n_27680;
assign n_27682 =  n_27677 &  n_27681;
assign n_27683 = ~n_23818 & ~n_26009;
assign n_27684 =  n_27228 &  n_27683;
assign n_27685 = ~n_1176 & ~n_24685;
assign n_27686 = ~n_24315 & ~n_23901;
assign n_27687 =  n_27685 &  n_27686;
assign n_27688 =  n_27684 &  n_27687;
assign n_27689 =  n_27682 &  n_27688;
assign n_27690 = ~n_25718 & ~n_16302;
assign n_27691 =  n_554 &  n_551;
assign n_27692 =  n_3628 &  n_27691;
assign n_27693 = ~n_27003 & ~n_27692;
assign n_27694 =  n_27690 &  n_27693;
assign n_27695 =  n_23685 &  n_26067;
assign n_27696 = ~n_27695 & ~n_25239;
assign n_27697 =  n_27696 &  n_26993;
assign n_27698 =  n_27694 &  n_27697;
assign n_27699 =  n_11 &  n_24749;
assign n_27700 = ~n_23140 & ~n_25004;
assign n_27701 = ~n_25972 &  n_27700;
assign n_27702 = ~n_27699 &  n_27701;
assign n_27703 =  n_27698 &  n_27702;
assign n_27704 = ~n_25021 & ~n_26306;
assign n_27705 = ~n_24957 & ~n_24201;
assign n_27706 =  n_27704 &  n_27705;
assign n_27707 = ~n_24221 & ~n_23882;
assign n_27708 = ~n_24226 & ~n_26368;
assign n_27709 =  n_27707 &  n_27708;
assign n_27710 = ~n_24120 & ~n_25918;
assign n_27711 = ~n_23331 &  n_27710;
assign n_27712 =  n_27709 &  n_27711;
assign n_27713 =  n_27706 &  n_27712;
assign n_27714 =  n_27703 &  n_27713;
assign n_27715 =  n_27689 &  n_27714;
assign n_27716 = ~n_23259 & ~n_26439;
assign n_27717 =  n_27048 & ~n_25955;
assign n_27718 =  n_27716 &  n_27717;
assign n_27719 = ~n_27141 & ~n_23545;
assign n_27720 = ~n_23804 &  n_27719;
assign n_27721 =  n_23329 &  n_560;
assign n_27722 = ~n_25683 & ~n_27721;
assign n_27723 =  n_27720 &  n_27722;
assign n_27724 =  n_27718 &  n_27723;
assign n_27725 =  n_554 &  n_762;
assign n_27726 = ~n_10474 &  n_3635;
assign n_27727 = ~n_27725 &  n_27726;
assign n_27728 =  n_23422 &  n_3628;
assign n_27729 = ~n_27728 & ~n_25863;
assign n_27730 =  n_4089 &  n_15;
assign n_27731 = ~n_25956 & ~n_27730;
assign n_27732 =  n_27729 &  n_27731;
assign n_27733 =  n_27727 &  n_27732;
assign n_27734 =  n_27724 &  n_27733;
assign n_27735 = ~n_25116 & ~n_26135;
assign n_27736 = ~n_24530 & ~n_4291;
assign n_27737 =  n_27735 &  n_27736;
assign n_27738 = ~n_25905 & ~n_23830;
assign n_27739 = ~n_26394 & ~n_3348;
assign n_27740 =  n_27738 &  n_27739;
assign n_27741 =  n_27737 &  n_27740;
assign n_27742 = ~n_23946 & ~n_25084;
assign n_27743 = ~n_3631 & ~n_13286;
assign n_27744 =  n_27742 &  n_27743;
assign n_27745 = ~n_156 & ~n_7856;
assign n_27746 = ~n_5650 & ~n_23293;
assign n_27747 =  n_27745 &  n_27746;
assign n_27748 =  n_27744 &  n_27747;
assign n_27749 =  n_27741 &  n_27748;
assign n_27750 =  n_27734 &  n_27749;
assign n_27751 =  n_27715 &  n_27750;
assign n_27752 =  n_27071 &  n_25670;
assign n_27753 = ~n_555 & ~n_6525;
assign n_27754 =  n_25671 & ~n_27753;
assign n_27755 = ~n_27754 & ~n_25454;
assign n_27756 =  n_27752 &  n_27755;
assign n_27757 =  n_24304 &  n_26774;
assign n_27758 = ~n_9300 & ~n_24947;
assign n_27759 = ~n_27757 &  n_27758;
assign n_27760 =  n_25282 & ~n_26147;
assign n_27761 =  n_27759 &  n_27760;
assign n_27762 =  n_27756 &  n_27761;
assign n_27763 =  n_24954 & ~n_27263;
assign n_27764 =  n_23256 & ~n_27763;
assign n_27765 = ~n_23897 & ~n_24946;
assign n_27766 =  n_27765 & ~n_26673;
assign n_27767 =  n_27764 &  n_27766;
assign n_27768 = ~n_23643 & ~n_27124;
assign n_27769 = ~n_26718 & ~n_23369;
assign n_27770 =  n_27768 &  n_27769;
assign n_27771 =  n_27767 &  n_27770;
assign n_27772 =  n_27762 &  n_27771;
assign n_27773 =  x_42 &  n_23386;
assign n_27774 = ~n_26947 & ~n_25897;
assign n_27775 = ~n_27773 &  n_27774;
assign n_27776 = ~n_25637 & ~n_17980;
assign n_27777 = ~n_24220 &  n_27776;
assign n_27778 =  n_27775 &  n_27777;
assign n_27779 = ~n_27016 & ~n_23941;
assign n_27780 =  n_27779 & ~n_26091;
assign n_27781 =  n_23883 &  n_23692;
assign n_27782 = ~n_27781 & ~n_23421;
assign n_27783 =  n_27780 &  n_27782;
assign n_27784 =  n_27778 &  n_27783;
assign n_27785 = ~n_3344 & ~n_4287;
assign n_27786 = ~n_26994 & ~n_20403;
assign n_27787 =  n_25168 &  n_27786;
assign n_27788 =  n_27785 &  n_27787;
assign n_27789 = ~x_256 & ~x_257;
assign n_27790 = ~x_258 & ~x_259;
assign n_27791 =  n_27789 &  n_27790;
assign n_27792 = ~x_252 & ~x_253;
assign n_27793 = ~x_254 & ~x_255;
assign n_27794 =  n_27792 &  n_27793;
assign n_27795 =  n_27791 &  n_27794;
assign n_27796 = ~x_264 & ~x_265;
assign n_27797 = ~x_266 & ~x_267;
assign n_27798 =  n_27796 &  n_27797;
assign n_27799 = ~x_260 & ~x_261;
assign n_27800 = ~x_262 & ~x_263;
assign n_27801 =  n_27799 &  n_27800;
assign n_27802 =  n_27798 &  n_27801;
assign n_27803 =  n_27795 &  n_27802;
assign n_27804 = ~x_240 & ~x_241;
assign n_27805 = ~x_242 & ~x_243;
assign n_27806 =  n_27804 &  n_27805;
assign n_27807 = ~x_236 & ~x_237;
assign n_27808 = ~x_238 & ~x_239;
assign n_27809 =  n_27807 &  n_27808;
assign n_27810 =  n_27806 &  n_27809;
assign n_27811 = ~x_248 & ~x_249;
assign n_27812 = ~x_250 & ~x_251;
assign n_27813 =  n_27811 &  n_27812;
assign n_27814 = ~x_244 & ~x_245;
assign n_27815 = ~x_246 & ~x_247;
assign n_27816 =  n_27814 &  n_27815;
assign n_27817 =  n_27813 &  n_27816;
assign n_27818 =  n_27810 &  n_27817;
assign n_27819 =  n_27803 &  n_27818;
assign n_27820 =  n_25017 &  n_27819;
assign n_27821 = ~n_25211 & ~n_27820;
assign n_27822 = ~n_24391 & ~n_22465;
assign n_27823 =  n_27821 &  n_27822;
assign n_27824 =  n_27788 &  n_27823;
assign n_27825 =  n_27784 &  n_27824;
assign n_27826 =  n_27772 &  n_27825;
assign n_27827 =  n_27751 &  n_27826;
assign n_27828 =  n_27674 &  n_27827;
assign n_27829 = ~n_27344 & ~n_26224;
assign n_27830 =  n_27829 & ~n_24778;
assign n_27831 = ~n_27278 & ~n_24038;
assign n_27832 = ~n_1037 & ~n_27831;
assign n_27833 =  n_23560 & ~n_23611;
assign n_27834 = ~n_27832 &  n_27833;
assign n_27835 =  n_27830 &  n_27834;
assign n_27836 =  n_11 &  n_25538;
assign n_27837 =  n_27177 & ~n_27836;
assign n_27838 = ~n_11 &  n_24018;
assign n_27839 =  n_349 &  n_13;
assign n_27840 =  n_24043 &  n_27839;
assign n_27841 = ~n_27840 & ~n_26168;
assign n_27842 = ~n_27838 &  n_27841;
assign n_27843 = ~n_25998 &  n_27842;
assign n_27844 = ~n_23137 &  n_27843;
assign n_27845 =  n_27837 &  n_27844;
assign n_27846 = ~n_27176 &  n_27845;
assign n_27847 = ~n_22973 &  n_27846;
assign n_27848 =  n_27835 &  n_27847;
assign n_27849 = ~n_24004 &  n_26872;
assign n_27850 = ~n_25876 &  n_27849;
assign n_27851 =  n_23732 & ~n_23763;
assign n_27852 =  n_24569 &  n_24050;
assign n_27853 = ~x_43 &  n_27852;
assign n_27854 = ~n_27853 & ~n_25864;
assign n_27855 = ~n_27851 &  n_27854;
assign n_27856 =  n_27850 &  n_27855;
assign n_27857 = ~x_43 &  n_20984;
assign n_27858 = ~n_358 & ~n_27857;
assign n_27859 = ~n_25701 &  n_27858;
assign n_27860 =  n_27856 &  n_27859;
assign n_27861 =  n_23178 &  n_27493;
assign n_27862 = ~n_23985 & ~n_27861;
assign n_27863 = ~n_23059 &  n_27862;
assign n_27864 = ~n_26720 & ~n_23327;
assign n_27865 =  n_27863 &  n_27864;
assign n_27866 =  n_27860 &  n_27865;
assign n_27867 = ~n_24839 & ~n_25635;
assign n_27868 =  n_27867 & ~n_24631;
assign n_27869 =  n_27079 & ~n_26698;
assign n_27870 =  n_27868 & ~n_27869;
assign n_27871 =  n_23600 &  n_27077;
assign n_27872 =  n_27870 &  n_27871;
assign n_27873 =  n_11 &  n_25218;
assign n_27874 =  n_23065 &  n_23460;
assign n_27875 = ~n_13871 & ~n_25027;
assign n_27876 = ~n_27874 &  n_27875;
assign n_27877 = ~n_27873 &  n_27876;
assign n_27878 = ~n_26343 & ~n_26023;
assign n_27879 = ~n_7661 &  n_27878;
assign n_27880 =  n_27877 &  n_27879;
assign n_27881 =  n_11 &  n_26107;
assign n_27882 = ~n_27881 & ~n_25487;
assign n_27883 =  n_27882 &  n_27221;
assign n_27884 =  x_3912 &  n_153;
assign n_27885 =  n_26465 &  n_27884;
assign n_27886 = ~n_27885 & ~n_27044;
assign n_27887 = ~n_24314 & ~n_23681;
assign n_27888 =  n_23252 & ~n_27887;
assign n_27889 = ~n_27888 &  n_26887;
assign n_27890 =  n_27886 &  n_27889;
assign n_27891 =  n_27883 &  n_27890;
assign n_27892 =  n_27880 &  n_27891;
assign n_27893 =  n_27872 &  n_27892;
assign n_27894 =  n_27866 &  n_27893;
assign n_27895 =  n_27848 &  n_27894;
assign n_27896 =  n_27828 &  n_27895;
assign n_27897 = ~n_23062 & ~n_25690;
assign n_27898 =  n_555 &  n_357;
assign n_27899 = ~n_26398 & ~n_27898;
assign n_27900 =  n_23134 &  n_23136;
assign n_27901 = ~n_27900 & ~n_23940;
assign n_27902 = ~n_24021 & ~n_13479;
assign n_27903 =  n_27901 &  n_27902;
assign n_27904 =  n_27899 &  n_27903;
assign n_27905 =  n_25875 &  n_25630;
assign n_27906 =  n_26454 &  n_27905;
assign n_27907 =  n_27904 &  n_27906;
assign n_27908 =  n_27897 &  n_27907;
assign n_27909 =  n_24014 &  n_557;
assign n_27910 = ~n_26215 & ~n_27909;
assign n_27911 =  n_6379 &  n_557;
assign n_27912 = ~n_27911 & ~n_26700;
assign n_27913 =  n_27910 &  n_27912;
assign n_27914 = ~n_26812 & ~n_27040;
assign n_27915 =  n_27913 &  n_27914;
assign n_27916 = ~n_26300 & ~n_26709;
assign n_27917 = ~n_14787 &  n_27916;
assign n_27918 =  n_27915 &  n_27917;
assign n_27919 = ~n_26426 & ~n_26142;
assign n_27920 =  n_27919 & ~n_26969;
assign n_27921 = ~x_42 &  n_8352;
assign n_27922 =  n_7079 &  n_27921;
assign n_27923 = ~n_27922 & ~n_25028;
assign n_27924 = ~n_6878 &  n_27923;
assign n_27925 = ~n_26154 &  n_27924;
assign n_27926 =  n_27920 &  n_27925;
assign n_27927 =  n_27918 &  n_27926;
assign n_27928 =  n_26324 & ~n_24901;
assign n_27929 =  n_27928 &  n_23543;
assign n_27930 = ~n_24515 & ~n_25662;
assign n_27931 =  n_11 & ~n_27930;
assign n_27932 = ~n_27931 &  n_27270;
assign n_27933 =  n_27929 &  n_27932;
assign n_27934 =  n_25296 &  n_25327;
assign n_27935 = ~n_24929 & ~n_26436;
assign n_27936 = ~n_27934 &  n_27935;
assign n_27937 =  x_37 &  n_24918;
assign n_27938 = ~n_26335 & ~n_27937;
assign n_27939 =  n_27936 &  n_27938;
assign n_27940 = ~n_24077 & ~n_26964;
assign n_27941 = ~n_23885 & ~n_23887;
assign n_27942 = ~n_10471 &  n_27941;
assign n_27943 =  n_27940 &  n_27942;
assign n_27944 =  n_27939 &  n_27943;
assign n_27945 =  n_27933 &  n_27944;
assign n_27946 =  n_27927 &  n_27945;
assign n_27947 = ~n_24965 & ~n_5653;
assign n_27948 =  n_27947 & ~n_26264;
assign n_27949 =  n_24303 &  n_27948;
assign n_27950 = ~n_26117 & ~n_26257;
assign n_27951 =  n_27950 & ~n_26862;
assign n_27952 =  n_27949 &  n_27951;
assign n_27953 = ~n_26817 & ~n_25943;
assign n_27954 =  x_42 &  n_25500;
assign n_27955 =  n_555 &  n_25044;
assign n_27956 = ~n_1901 & ~n_27955;
assign n_27957 = ~n_27954 &  n_27956;
assign n_27958 =  n_27953 &  n_27957;
assign n_27959 = ~n_26102 & ~n_25271;
assign n_27960 =  n_11 &  n_24925;
assign n_27961 = ~n_27960 & ~n_24911;
assign n_27962 =  n_27959 &  n_27961;
assign n_27963 =  n_27958 &  n_27962;
assign n_27964 =  n_27952 &  n_27963;
assign n_27965 =  n_11 &  n_26351;
assign n_27966 =  n_25175 & ~n_25206;
assign n_27967 = ~n_27965 & ~n_27966;
assign n_27968 =  n_27967 & ~n_24787;
assign n_27969 = ~n_3347 & ~n_12910;
assign n_27970 = ~n_26975 & ~n_25653;
assign n_27971 = ~n_16496 &  n_27970;
assign n_27972 =  n_27969 &  n_27971;
assign n_27973 =  n_27968 &  n_27972;
assign n_27974 = ~x_43 &  n_25533;
assign n_27975 = ~n_27974 & ~n_25892;
assign n_27976 =  x_3416 &  n_25890;
assign n_27977 = ~n_24741 & ~n_27976;
assign n_27978 =  n_27975 &  n_27977;
assign n_27979 =  n_24695 &  n_26263;
assign n_27980 =  n_27978 &  n_27979;
assign n_27981 =  n_27973 &  n_27980;
assign n_27982 =  n_27964 &  n_27981;
assign n_27983 =  n_27946 &  n_27982;
assign n_27984 =  n_3144 &  n_24772;
assign n_27985 =  n_11 &  n_26081;
assign n_27986 = ~n_26430 & ~n_27985;
assign n_27987 = ~n_27984 &  n_27986;
assign n_27988 =  n_25678 &  n_27987;
assign n_27989 = ~n_23693 & ~n_23623;
assign n_27990 =  n_25153 &  n_26825;
assign n_27991 =  n_21954 &  n_27691;
assign n_27992 = ~n_27990 & ~n_27991;
assign n_27993 =  n_26837 &  n_27992;
assign n_27994 =  n_27989 &  n_27993;
assign n_27995 =  n_27224 &  n_27994;
assign n_27996 =  n_25849 &  n_27995;
assign n_27997 =  n_27988 &  n_27996;
assign n_27998 =  n_24222 &  n_24800;
assign n_27999 = ~n_27998 & ~n_24801;
assign n_28000 =  n_27276 &  n_26172;
assign n_28001 =  n_26175 &  n_24594;
assign n_28002 =  n_28000 &  n_28001;
assign n_28003 =  n_27999 &  n_28002;
assign n_28004 =  n_3622 &  n_26742;
assign n_28005 = ~n_26712 & ~n_26866;
assign n_28006 =  n_28004 &  n_28005;
assign n_28007 = ~n_25988 & ~n_14267;
assign n_28008 =  n_28007 & ~n_19108;
assign n_28009 = ~n_21565 & ~n_10873;
assign n_28010 =  n_24630 &  n_1502;
assign n_28011 = ~n_3624 & ~n_28010;
assign n_28012 = ~n_26485 &  n_28011;
assign n_28013 = ~n_26942 &  n_28012;
assign n_28014 =  n_28009 &  n_28013;
assign n_28015 =  n_28008 &  n_28014;
assign n_28016 =  n_28006 &  n_28015;
assign n_28017 =  n_28003 &  n_28016;
assign n_28018 =  n_27997 &  n_28017;
assign n_28019 =  n_27983 &  n_28018;
assign n_28020 =  n_27908 &  n_28019;
assign n_28021 =  n_27896 &  n_28020;
assign n_28022 =  n_27580 &  n_28021;
assign n_28023 = ~n_27491 &  n_28022;
assign n_28024 = ~n_27490 &  n_28023;
assign n_28025 = ~n_27363 &  n_28024;
assign n_28026 = ~n_22082 &  n_28025;
assign n_28027 =  x_40 & ~n_28026;
assign n_28028 = ~x_40 &  n_28026;
assign n_28029 = ~n_28027 & ~n_28028;
assign n_28030 = ~n_26638 & ~n_22465;
assign n_28031 = ~n_22209 &  n_28030;
assign n_28032 =  n_25718 & ~n_25843;
assign n_28033 = ~n_22210 & ~n_27487;
assign n_28034 = ~n_22337 &  n_28033;
assign n_28035 = ~n_28032 &  n_28034;
assign n_28036 = ~n_27998 & ~n_3347;
assign n_28037 =  n_26259 &  n_28036;
assign n_28038 =  n_28037 &  n_25885;
assign n_28039 =  n_25881 &  n_28038;
assign n_28040 =  n_27159 &  n_25699;
assign n_28041 =  n_25528 &  n_20207;
assign n_28042 = ~n_28041 &  n_24934;
assign n_28043 =  n_26372 &  n_28042;
assign n_28044 = ~n_23386 & ~n_27330;
assign n_28045 = ~x_43 &  n_25544;
assign n_28046 =  n_25856 &  n_25246;
assign n_28047 = ~n_28045 & ~n_28046;
assign n_28048 = ~x_43 &  n_25535;
assign n_28049 = ~x_42 &  n_28048;
assign n_28050 =  n_28047 & ~n_28049;
assign n_28051 =  n_28044 &  n_28050;
assign n_28052 =  n_28043 &  n_28051;
assign n_28053 =  n_23004 &  n_26394;
assign n_28054 = ~n_25240 & ~n_28053;
assign n_28055 =  n_28052 &  n_28054;
assign n_28056 =  n_28040 &  n_28055;
assign n_28057 =  n_28039 &  n_28056;
assign n_28058 =  n_25855 &  n_28057;
assign n_28059 = ~n_23988 & ~n_24954;
assign n_28060 =  n_6378 &  n_23987;
assign n_28061 = ~n_28060 & ~n_25093;
assign n_28062 =  n_28059 &  n_28061;
assign n_28063 = ~n_24212 & ~n_27960;
assign n_28064 =  n_28062 &  n_28063;
assign n_28065 = ~n_25231 & ~n_10479;
assign n_28066 = ~n_28010 & ~n_25010;
assign n_28067 =  n_28065 &  n_28066;
assign n_28068 = ~n_12909 & ~n_26992;
assign n_28069 = ~n_25455 & ~n_27122;
assign n_28070 =  n_28068 &  n_28069;
assign n_28071 =  n_28067 &  n_28070;
assign n_28072 =  n_552 &  n_24630;
assign n_28073 = ~n_28072 & ~n_26827;
assign n_28074 =  n_13672 &  n_355;
assign n_28075 = ~n_28074 & ~n_26092;
assign n_28076 =  n_28073 &  n_28075;
assign n_28077 = ~n_27052 & ~n_26411;
assign n_28078 =  n_554 &  n_25971;
assign n_28079 = ~n_23140 & ~n_28078;
assign n_28080 =  n_28077 &  n_28079;
assign n_28081 =  n_28076 &  n_28080;
assign n_28082 =  n_28071 &  n_28081;
assign n_28083 =  n_28064 &  n_28082;
assign n_28084 = ~n_22721 &  n_24228;
assign n_28085 = ~n_24694 &  n_27947;
assign n_28086 =  n_28084 &  n_28085;
assign n_28087 = ~n_25937 & ~n_23423;
assign n_28088 =  n_28087 & ~n_26102;
assign n_28089 =  n_11 &  n_26085;
assign n_28090 = ~n_27985 & ~n_28089;
assign n_28091 =  n_8350 &  n_28090;
assign n_28092 =  n_28088 &  n_28091;
assign n_28093 =  n_28086 &  n_28092;
assign n_28094 =  n_28083 &  n_28093;
assign n_28095 = ~n_24592 & ~n_3340;
assign n_28096 = ~n_26486 & ~n_24074;
assign n_28097 =  n_28095 &  n_28096;
assign n_28098 = ~n_25289 & ~n_24060;
assign n_28099 = ~n_26068 & ~n_26070;
assign n_28100 =  n_28098 &  n_28099;
assign n_28101 =  n_28097 &  n_28100;
assign n_28102 = ~n_24703 & ~n_10875;
assign n_28103 = ~n_23804 &  n_28102;
assign n_28104 = ~n_24010 & ~n_27047;
assign n_28105 =  n_28103 &  n_28104;
assign n_28106 =  n_11 &  n_770;
assign n_28107 = ~n_28106 & ~n_24065;
assign n_28108 = ~n_24005 & ~n_24021;
assign n_28109 =  n_28107 &  n_28108;
assign n_28110 =  n_28105 &  n_28109;
assign n_28111 =  n_28101 &  n_28110;
assign n_28112 =  n_11 &  n_25343;
assign n_28113 = ~n_24946 & ~n_28112;
assign n_28114 = ~n_23839 & ~n_24980;
assign n_28115 =  n_28113 &  n_28114;
assign n_28116 = ~n_24907 & ~n_27840;
assign n_28117 = ~n_26210 & ~n_23890;
assign n_28118 =  n_28116 &  n_28117;
assign n_28119 = ~x_43 &  n_25516;
assign n_28120 =  n_23692 &  n_24971;
assign n_28121 = ~n_28119 & ~n_28120;
assign n_28122 =  n_28118 &  n_28121;
assign n_28123 =  n_28115 &  n_28122;
assign n_28124 =  n_24224 & ~n_23818;
assign n_28125 = ~n_25904 & ~n_3343;
assign n_28126 =  n_28124 &  n_28125;
assign n_28127 = ~n_24427 & ~n_25251;
assign n_28128 = ~n_25227 & ~n_26363;
assign n_28129 =  n_28127 &  n_28128;
assign n_28130 =  n_28126 &  n_28129;
assign n_28131 =  n_28123 &  n_28130;
assign n_28132 =  n_28111 &  n_28131;
assign n_28133 =  n_28094 &  n_28132;
assign n_28134 = ~n_6183 & ~n_26866;
assign n_28135 = ~n_8364 & ~n_24686;
assign n_28136 =  n_28134 &  n_28135;
assign n_28137 =  n_27290 &  n_27321;
assign n_28138 = ~n_28137 & ~n_26180;
assign n_28139 =  n_28136 &  n_28138;
assign n_28140 = ~n_27836 &  n_23256;
assign n_28141 = ~n_25027 & ~n_25641;
assign n_28142 =  n_28141 &  n_26312;
assign n_28143 =  n_28140 &  n_28142;
assign n_28144 =  n_28139 &  n_28143;
assign n_28145 = ~n_26323 & ~n_25624;
assign n_28146 =  n_27596 &  n_27609;
assign n_28147 =  n_28145 &  n_28146;
assign n_28148 =  n_7467 &  n_25108;
assign n_28149 = ~n_28148 &  n_26337;
assign n_28150 = ~n_27278 & ~n_12293;
assign n_28151 =  n_28149 &  n_28150;
assign n_28152 =  n_28147 &  n_28151;
assign n_28153 =  n_28144 &  n_28152;
assign n_28154 =  n_6379 &  n_23829;
assign n_28155 = ~n_28154 & ~n_27911;
assign n_28156 =  n_28155 &  n_24761;
assign n_28157 = ~n_14260 & ~n_13871;
assign n_28158 = ~n_25338 &  n_28157;
assign n_28159 =  n_28156 &  n_28158;
assign n_28160 =  n_23846 & ~n_27132;
assign n_28161 = ~n_4287 & ~n_23598;
assign n_28162 =  n_28160 &  n_28161;
assign n_28163 =  n_28159 &  n_28162;
assign n_28164 = ~n_25651 & ~n_25652;
assign n_28165 = ~n_16496 &  n_28164;
assign n_28166 = ~n_24307 & ~n_25927;
assign n_28167 = ~n_25098 &  n_28166;
assign n_28168 =  n_28165 &  n_28167;
assign n_28169 = ~n_24313 & ~n_24124;
assign n_28170 =  n_28169 & ~n_23365;
assign n_28171 =  n_28168 &  n_28170;
assign n_28172 = ~n_1176 & ~n_24317;
assign n_28173 =  n_28172 &  n_28009;
assign n_28174 = ~n_23558 & ~n_25659;
assign n_28175 =  n_554 &  n_6883;
assign n_28176 = ~n_28175 & ~n_26173;
assign n_28177 = ~n_25007 & ~n_20791;
assign n_28178 =  n_28176 &  n_28177;
assign n_28179 =  n_28174 &  n_28178;
assign n_28180 =  n_28173 &  n_28179;
assign n_28181 =  n_28171 &  n_28180;
assign n_28182 =  n_28163 &  n_28181;
assign n_28183 =  n_28153 &  n_28182;
assign n_28184 =  n_28133 &  n_28183;
assign n_28185 = ~n_23137 & ~n_25865;
assign n_28186 =  n_28185 &  n_27130;
assign n_28187 = ~n_24696 & ~n_25004;
assign n_28188 =  n_13872 &  n_24569;
assign n_28189 = ~n_28188 & ~n_27045;
assign n_28190 =  n_28187 &  n_28189;
assign n_28191 =  n_9884 &  n_23984;
assign n_28192 =  n_28190 & ~n_28191;
assign n_28193 =  n_28186 &  n_28192;
assign n_28194 = ~n_1038 & ~n_152;
assign n_28195 =  n_24581 & ~n_28194;
assign n_28196 =  n_26308 & ~n_28195;
assign n_28197 = ~n_26706 &  n_28196;
assign n_28198 = ~n_25911 & ~n_26839;
assign n_28199 =  n_26875 &  n_28198;
assign n_28200 =  n_8363 & ~n_24564;
assign n_28201 =  n_28199 &  n_28200;
assign n_28202 =  n_28197 &  n_28201;
assign n_28203 =  n_28193 &  n_28202;
assign n_28204 =  n_26165 &  n_27928;
assign n_28205 =  n_27285 &  n_24514;
assign n_28206 =  n_28204 &  n_28205;
assign n_28207 = ~n_4283 & ~n_26473;
assign n_28208 =  x_42 & ~n_28207;
assign n_28209 =  n_27942 & ~n_28208;
assign n_28210 =  n_24505 & ~n_26190;
assign n_28211 =  n_28209 &  n_28210;
assign n_28212 =  n_28206 &  n_28211;
assign n_28213 =  n_28203 &  n_28212;
assign n_28214 =  n_27776 & ~n_8351;
assign n_28215 =  n_28214 & ~n_26247;
assign n_28216 = ~n_9691 & ~n_24057;
assign n_28217 =  n_28216 &  n_26015;
assign n_28218 =  n_7467 &  n_6526;
assign n_28219 = ~n_28218 & ~n_3349;
assign n_28220 =  n_28217 &  n_28219;
assign n_28221 =  n_28215 &  n_28220;
assign n_28222 = ~n_24629 & ~n_25157;
assign n_28223 = ~n_27885 &  n_28222;
assign n_28224 =  x_41 &  n_2882;
assign n_28225 = ~n_9 & ~n_24575;
assign n_28226 =  n_1 & ~n_28225;
assign n_28227 = ~n_28226 & ~n_13105;
assign n_28228 = ~n_28224 &  n_28227;
assign n_28229 =  n_28223 &  n_28228;
assign n_28230 = ~n_25632 & ~n_1044;
assign n_28231 =  n_28229 &  n_28230;
assign n_28232 =  n_28221 &  n_28231;
assign n_28233 = ~n_23688 & ~n_27007;
assign n_28234 = ~n_24918 & ~n_25626;
assign n_28235 =  n_28233 &  n_28234;
assign n_28236 = ~n_24926 & ~n_26114;
assign n_28237 =  n_28235 &  n_28236;
assign n_28238 = ~n_26154 & ~n_25676;
assign n_28239 =  n_28237 &  n_28238;
assign n_28240 =  n_28007 & ~n_25024;
assign n_28241 =  n_28240 & ~n_27336;
assign n_28242 = ~n_26262 & ~n_24529;
assign n_28243 = ~n_23676 &  n_28242;
assign n_28244 =  n_28241 &  n_28243;
assign n_28245 =  n_28239 &  n_28244;
assign n_28246 =  n_28232 &  n_28245;
assign n_28247 =  n_28213 &  n_28246;
assign n_28248 =  n_28184 &  n_28247;
assign n_28249 = ~n_26491 & ~n_8355;
assign n_28250 =  n_27590 &  n_28249;
assign n_28251 = ~x_42 &  n_1504;
assign n_28252 = ~n_2882 & ~n_28251;
assign n_28253 = ~x_41 & ~n_28252;
assign n_28254 = ~n_28253 &  n_27868;
assign n_28255 =  n_27074 &  n_23547;
assign n_28256 =  n_28254 &  n_28255;
assign n_28257 =  n_28250 &  n_28256;
assign n_28258 = ~n_27501 &  n_23015;
assign n_28259 =  n_28257 &  n_28258;
assign n_28260 = ~n_26231 & ~n_25288;
assign n_28261 =  n_28260 & ~n_24779;
assign n_28262 =  n_25248 & ~n_26812;
assign n_28263 = ~n_25454 &  n_28262;
assign n_28264 = ~n_26306 & ~n_26822;
assign n_28265 = ~n_27974 &  n_28264;
assign n_28266 =  n_28263 &  n_28265;
assign n_28267 =  n_28261 &  n_28266;
assign n_28268 = ~n_24893 &  n_27774;
assign n_28269 =  n_24196 &  n_28268;
assign n_28270 =  n_27188 & ~n_27219;
assign n_28271 =  n_25591 & ~n_25622;
assign n_28272 = ~n_28270 & ~n_28271;
assign n_28273 =  n_25348 &  n_25379;
assign n_28274 = ~n_28273 &  n_26880;
assign n_28275 =  n_28272 &  n_28274;
assign n_28276 =  n_28269 &  n_28275;
assign n_28277 = ~n_20078 & ~n_6881;
assign n_28278 = ~n_24591 &  n_28277;
assign n_28279 =  n_23896 &  n_28278;
assign n_28280 =  n_28279 &  n_24785;
assign n_28281 =  n_28276 &  n_28280;
assign n_28282 =  n_28267 &  n_28281;
assign n_28283 =  n_3341 &  n_3620;
assign n_28284 = ~n_23326 & ~n_7274;
assign n_28285 = ~n_25700 &  n_28284;
assign n_28286 = ~n_28283 &  n_28285;
assign n_28287 =  n_28286 &  n_27118;
assign n_28288 =  n_27119 &  n_23551;
assign n_28289 =  n_28287 &  n_28288;
assign n_28290 = ~n_26135 & ~n_25100;
assign n_28291 = ~n_25892 &  n_28290;
assign n_28292 = ~n_27909 & ~n_25016;
assign n_28293 =  n_28292 &  n_26031;
assign n_28294 =  n_28291 &  n_28293;
assign n_28295 =  n_28294 & ~n_23294;
assign n_28296 =  n_24753 &  n_354;
assign n_28297 =  n_8818 &  n_1698;
assign n_28298 = ~n_25008 & ~n_28297;
assign n_28299 = ~n_28296 &  n_28298;
assign n_28300 =  n_356 &  n_10874;
assign n_28301 = ~n_27152 & ~n_28300;
assign n_28302 = ~n_26174 &  n_28301;
assign n_28303 =  n_28299 &  n_28302;
assign n_28304 =  n_1040 &  n_26122;
assign n_28305 = ~n_23098 &  n_28304;
assign n_28306 =  n_28303 & ~n_28305;
assign n_28307 =  n_28295 &  n_28306;
assign n_28308 =  n_28289 &  n_28307;
assign n_28309 =  n_28282 &  n_28308;
assign n_28310 =  n_28259 &  n_28309;
assign n_28311 =  n_28248 &  n_28310;
assign n_28312 =  n_23630 &  n_24431;
assign n_28313 = ~n_24587 & ~n_23632;
assign n_28314 = ~n_28312 &  n_28313;
assign n_28315 =  n_28314 &  n_27164;
assign n_28316 =  n_25285 &  n_28315;
assign n_28317 = ~n_24358 & ~n_26775;
assign n_28318 = ~n_24391 & ~n_26086;
assign n_28319 =  n_28317 &  n_28318;
assign n_28320 =  n_27829 &  n_28319;
assign n_28321 = ~n_26467 & ~n_25496;
assign n_28322 = ~n_26942 & ~n_26964;
assign n_28323 = ~n_26410 &  n_28322;
assign n_28324 =  n_28321 &  n_28323;
assign n_28325 =  n_26721 &  n_28324;
assign n_28326 =  n_28320 &  n_28325;
assign n_28327 = ~n_23330 & ~n_25032;
assign n_28328 =  n_24875 & ~n_25490;
assign n_28329 =  n_23899 &  n_28328;
assign n_28330 =  n_28327 &  n_28329;
assign n_28331 =  n_26169 &  n_27324;
assign n_28332 =  n_27289 &  n_28331;
assign n_28333 =  n_28330 &  n_28332;
assign n_28334 = ~n_23682 &  n_26022;
assign n_28335 = ~n_25950 &  n_25081;
assign n_28336 = ~n_26023 & ~n_28335;
assign n_28337 =  n_26011 &  n_28336;
assign n_28338 =  n_28334 &  n_28337;
assign n_28339 =  n_27668 &  n_27652;
assign n_28340 =  n_28338 &  n_28339;
assign n_28341 =  n_28333 &  n_28340;
assign n_28342 =  n_28326 &  n_28341;
assign n_28343 = ~n_22973 & ~n_26140;
assign n_28344 =  n_27995 &  n_26434;
assign n_28345 =  n_26443 &  n_28344;
assign n_28346 =  n_28343 &  n_28345;
assign n_28347 =  n_28342 &  n_28346;
assign n_28348 =  n_28316 &  n_28347;
assign n_28349 =  n_28311 &  n_28348;
assign n_28350 =  n_28058 &  n_28349;
assign n_28351 = ~n_25845 &  n_28350;
assign n_28352 = ~n_26637 &  n_28351;
assign n_28353 =  n_28035 &  n_28352;
assign n_28354 =  n_28031 &  n_28353;
assign n_28355 =  x_39 & ~n_28354;
assign n_28356 = ~x_39 &  n_28354;
assign n_28357 = ~n_28355 & ~n_28356;
assign n_28358 =  n_27576 & ~n_25264;
assign n_28359 =  n_28037 &  n_28358;
assign n_28360 =  n_27505 &  n_28359;
assign n_28361 =  n_27500 &  n_28360;
assign n_28362 = ~n_24521 & ~n_25632;
assign n_28363 = ~n_26334 & ~n_25331;
assign n_28364 = ~x_43 &  n_26468;
assign n_28365 = ~n_28364 &  n_26890;
assign n_28366 =  n_28363 &  n_28365;
assign n_28367 =  n_28362 &  n_28366;
assign n_28368 =  n_24392 &  n_27590;
assign n_28369 =  n_28367 &  n_28368;
assign n_28370 =  n_25090 &  n_26329;
assign n_28371 = ~n_26869 &  n_25099;
assign n_28372 =  n_28370 &  n_28371;
assign n_28373 = ~n_26411 & ~n_558;
assign n_28374 = ~n_25346 &  n_28373;
assign n_28375 =  n_26867 &  n_27989;
assign n_28376 =  n_28374 &  n_28375;
assign n_28377 =  n_28372 &  n_28376;
assign n_28378 =  n_26886 & ~n_27593;
assign n_28379 = ~n_25046 & ~n_26922;
assign n_28380 =  n_28378 &  n_28379;
assign n_28381 =  x_42 &  n_26163;
assign n_28382 = ~n_28137 & ~n_28381;
assign n_28383 =  n_25101 &  n_26331;
assign n_28384 =  n_28382 &  n_28383;
assign n_28385 =  n_28380 &  n_28384;
assign n_28386 =  n_28377 &  n_28385;
assign n_28387 =  n_28369 &  n_28386;
assign n_28388 = ~n_27344 & ~n_25851;
assign n_28389 = ~n_23676 & ~n_26778;
assign n_28390 = ~n_25175 & ~n_25907;
assign n_28391 = ~n_26133 &  n_28390;
assign n_28392 = ~n_27965 &  n_28391;
assign n_28393 =  n_28389 &  n_28392;
assign n_28394 =  n_28388 &  n_28393;
assign n_28395 = ~n_26352 & ~n_25663;
assign n_28396 = ~n_26845 &  n_28395;
assign n_28397 =  n_26251 &  n_28396;
assign n_28398 = ~n_27181 &  n_24791;
assign n_28399 =  n_28397 &  n_28398;
assign n_28400 =  n_28394 &  n_28399;
assign n_28401 =  n_28387 &  n_28400;
assign n_28402 = ~n_25988 & ~n_14261;
assign n_28403 = ~n_6527 & ~n_25236;
assign n_28404 =  n_28402 &  n_28403;
assign n_28405 = ~n_23468 & ~n_2686;
assign n_28406 = ~n_25905 & ~n_26068;
assign n_28407 =  n_28405 &  n_28406;
assign n_28408 =  n_28404 &  n_28407;
assign n_28409 = ~n_22337 & ~n_26131;
assign n_28410 =  n_17785 &  n_3619;
assign n_28411 = ~n_23251 & ~n_28410;
assign n_28412 =  n_28409 &  n_28411;
assign n_28413 = ~n_10473 & ~n_10;
assign n_28414 = ~n_27911 &  n_28413;
assign n_28415 = ~n_25339 & ~n_25625;
assign n_28416 =  n_28414 &  n_28415;
assign n_28417 =  n_28412 &  n_28416;
assign n_28418 =  n_28408 &  n_28417;
assign n_28419 =  n_25212 &  n_21758;
assign n_28420 = ~n_26205 & ~n_28419;
assign n_28421 = ~n_24121 & ~n_23887;
assign n_28422 =  n_28420 &  n_28421;
assign n_28423 = ~x_43 &  n_24041;
assign n_28424 = ~n_28423 & ~n_25648;
assign n_28425 = ~n_24210 & ~n_28112;
assign n_28426 =  n_28424 &  n_28425;
assign n_28427 =  n_28422 &  n_28426;
assign n_28428 = ~n_22717 & ~n_24965;
assign n_28429 = ~n_24591 & ~n_26021;
assign n_28430 =  n_28428 &  n_28429;
assign n_28431 = ~n_28089 & ~n_24760;
assign n_28432 = ~n_26508 & ~n_4283;
assign n_28433 =  n_28431 &  n_28432;
assign n_28434 =  n_28430 &  n_28433;
assign n_28435 =  n_28427 &  n_28434;
assign n_28436 =  n_28418 &  n_28435;
assign n_28437 = ~n_27581 & ~n_24115;
assign n_28438 = ~n_26401 & ~n_19694;
assign n_28439 =  n_28438 & ~n_25216;
assign n_28440 =  n_24312 &  n_28439;
assign n_28441 =  n_28437 &  n_28440;
assign n_28442 = ~n_10081 &  n_25492;
assign n_28443 =  n_554 &  n_25153;
assign n_28444 =  x_42 &  n_770;
assign n_28445 = ~n_28443 & ~n_28444;
assign n_28446 =  n_28442 &  n_28445;
assign n_28447 = ~n_24005 & ~n_19500;
assign n_28448 =  n_27053 &  n_28102;
assign n_28449 =  n_28447 &  n_28448;
assign n_28450 =  n_28446 &  n_28449;
assign n_28451 = ~n_24957 & ~n_27284;
assign n_28452 =  n_28292 & ~n_26350;
assign n_28453 =  n_28451 &  n_28452;
assign n_28454 =  n_28450 &  n_28453;
assign n_28455 =  n_28441 &  n_28454;
assign n_28456 =  n_28436 &  n_28455;
assign n_28457 = ~n_23558 & ~n_27838;
assign n_28458 =  n_28457 & ~n_26225;
assign n_28459 =  n_26031 & ~n_26315;
assign n_28460 =  n_28458 &  n_28459;
assign n_28461 = ~n_24592 & ~n_25985;
assign n_28462 =  n_26241 &  n_28461;
assign n_28463 = ~n_10476 & ~n_26992;
assign n_28464 = ~n_21759 &  n_28463;
assign n_28465 =  n_25168 &  n_28464;
assign n_28466 =  n_28462 &  n_28465;
assign n_28467 =  n_28460 &  n_28466;
assign n_28468 = ~n_27721 & ~n_8055;
assign n_28469 = ~n_26673 &  n_28468;
assign n_28470 = ~n_24468 & ~n_24435;
assign n_28471 = ~n_24874 & ~n_27955;
assign n_28472 =  n_28470 &  n_28471;
assign n_28473 =  n_28469 &  n_28472;
assign n_28474 = ~n_27900 & ~n_26718;
assign n_28475 =  n_23689 & ~n_27851;
assign n_28476 =  n_28474 &  n_28475;
assign n_28477 =  n_28473 &  n_28476;
assign n_28478 =  n_28467 &  n_28477;
assign n_28479 = ~n_23849 & ~n_24009;
assign n_28480 = ~n_24595 & ~n_25652;
assign n_28481 =  n_28479 &  n_28480;
assign n_28482 = ~n_26209 & ~n_26212;
assign n_28483 = ~n_24313 & ~n_5657;
assign n_28484 =  n_28482 &  n_28483;
assign n_28485 =  n_28481 &  n_28484;
assign n_28486 = ~n_27152 & ~n_25047;
assign n_28487 = ~n_28195 & ~n_25003;
assign n_28488 =  n_28486 &  n_28487;
assign n_28489 = ~n_27079 & ~n_10869;
assign n_28490 = ~n_24587 & ~n_10873;
assign n_28491 =  n_28489 &  n_28490;
assign n_28492 =  n_28488 &  n_28491;
assign n_28493 =  n_28485 &  n_28492;
assign n_28494 = ~n_25226 & ~n_25882;
assign n_28495 =  n_18914 &  n_5981;
assign n_28496 = ~n_27016 & ~n_28495;
assign n_28497 =  n_28494 &  n_28496;
assign n_28498 =  n_24043 &  n_10275;
assign n_28499 = ~n_25033 & ~n_28498;
assign n_28500 = ~n_23994 & ~n_23882;
assign n_28501 =  n_28499 &  n_28500;
assign n_28502 = ~n_28060 & ~n_23545;
assign n_28503 = ~n_24687 & ~n_23615;
assign n_28504 =  n_28502 &  n_28503;
assign n_28505 =  n_28501 &  n_28504;
assign n_28506 =  n_28497 &  n_28505;
assign n_28507 =  n_28493 &  n_28506;
assign n_28508 =  n_24232 & ~n_26189;
assign n_28509 = ~n_26420 & ~n_24302;
assign n_28510 =  n_28508 &  n_28509;
assign n_28511 = ~n_17077 & ~n_23812;
assign n_28512 = ~n_25021 & ~n_23624;
assign n_28513 =  n_28511 &  n_28512;
assign n_28514 = ~n_24872 & ~n_24195;
assign n_28515 =  n_28513 &  n_28514;
assign n_28516 =  n_28510 &  n_28515;
assign n_28517 =  n_28507 &  n_28516;
assign n_28518 =  n_28478 &  n_28517;
assign n_28519 =  n_28456 &  n_28518;
assign n_28520 =  n_28401 &  n_28519;
assign n_28521 = ~n_23678 &  n_24778;
assign n_28522 =  n_26141 &  n_25206;
assign n_28523 = ~n_28521 & ~n_28522;
assign n_28524 =  n_27862 &  n_28523;
assign n_28525 =  n_27110 &  n_27883;
assign n_28526 =  n_23250 &  n_28525;
assign n_28527 =  n_28524 &  n_28526;
assign n_28528 =  n_14785 & ~n_23938;
assign n_28529 =  n_154 &  n_28528;
assign n_28530 = ~n_28529 & ~n_23804;
assign n_28531 =  n_27953 & ~n_28120;
assign n_28532 = ~x_2394 &  n_23875;
assign n_28533 =  n_4088 &  n_28532;
assign n_28534 =  n_8053 &  n_28533;
assign n_28535 =  n_23873 &  n_28534;
assign n_28536 = ~n_27820 & ~n_28535;
assign n_28537 =  n_28536 & ~n_19494;
assign n_28538 =  n_28531 &  n_28537;
assign n_28539 =  n_28530 &  n_28538;
assign n_28540 = ~n_23008 & ~n_26395;
assign n_28541 =  n_28539 &  n_28540;
assign n_28542 =  n_28527 &  n_28541;
assign n_28543 = ~x_43 &  n_14786;
assign n_28544 = ~n_15919 & ~n_25651;
assign n_28545 = ~n_28543 &  n_28544;
assign n_28546 =  n_8053 &  n_24949;
assign n_28547 = ~n_24037 & ~n_19498;
assign n_28548 = ~n_28546 &  n_28547;
assign n_28549 = ~n_9429 &  n_28548;
assign n_28550 =  n_28545 &  n_28549;
assign n_28551 = ~n_27665 & ~n_24961;
assign n_28552 =  n_25248 &  n_28551;
assign n_28553 =  n_27600 &  n_28552;
assign n_28554 = ~n_25940 & ~n_25633;
assign n_28555 =  n_28554 &  n_27231;
assign n_28556 =  n_28553 &  n_28555;
assign n_28557 =  n_28550 &  n_28556;
assign n_28558 = ~n_26217 & ~n_24201;
assign n_28559 = ~n_14265 &  n_28558;
assign n_28560 =  n_26450 &  n_28559;
assign n_28561 = ~n_27960 & ~n_26198;
assign n_28562 = ~n_25500 &  n_28561;
assign n_28563 =  n_28560 &  n_28562;
assign n_28564 = ~n_27122 & ~n_27124;
assign n_28565 = ~n_23455 & ~n_27763;
assign n_28566 =  n_28564 &  n_28565;
assign n_28567 = ~x_4604 & ~x_4605;
assign n_28568 = ~x_4606 & ~x_4607;
assign n_28569 =  n_28567 &  n_28568;
assign n_28570 = ~x_4600 & ~x_4601;
assign n_28571 = ~x_4602 & ~x_4603;
assign n_28572 =  n_28570 &  n_28571;
assign n_28573 =  n_28569 &  n_28572;
assign n_28574 = ~x_4612 & ~x_4613;
assign n_28575 = ~x_4614 & ~x_4615;
assign n_28576 =  n_28574 &  n_28575;
assign n_28577 = ~x_4608 & ~x_4609;
assign n_28578 = ~x_4610 & ~x_4611;
assign n_28579 =  n_28577 &  n_28578;
assign n_28580 =  n_28576 &  n_28579;
assign n_28581 =  n_28573 &  n_28580;
assign n_28582 = ~x_4588 & ~x_4589;
assign n_28583 = ~x_4590 & ~x_4591;
assign n_28584 =  n_28582 &  n_28583;
assign n_28585 = ~x_4584 & ~x_4585;
assign n_28586 = ~x_4586 & ~x_4587;
assign n_28587 =  n_28585 &  n_28586;
assign n_28588 =  n_28584 &  n_28587;
assign n_28589 = ~x_4596 & ~x_4597;
assign n_28590 = ~x_4598 & ~x_4599;
assign n_28591 =  n_28589 &  n_28590;
assign n_28592 = ~x_4592 & ~x_4593;
assign n_28593 = ~x_4594 & ~x_4595;
assign n_28594 =  n_28592 &  n_28593;
assign n_28595 =  n_28591 &  n_28594;
assign n_28596 =  n_28588 &  n_28595;
assign n_28597 =  n_28581 &  n_28596;
assign n_28598 =  n_25083 & ~n_28597;
assign n_28599 = ~n_24056 & ~n_27695;
assign n_28600 = ~n_26018 &  n_28599;
assign n_28601 = ~n_28598 &  n_28600;
assign n_28602 =  n_28566 &  n_28601;
assign n_28603 =  n_28563 &  n_28602;
assign n_28604 =  n_28557 &  n_28603;
assign n_28605 =  n_27129 &  n_27877;
assign n_28606 =  n_27890 &  n_27114;
assign n_28607 =  n_28605 &  n_28606;
assign n_28608 = ~n_28305 &  n_28286;
assign n_28609 =  n_27134 &  n_27879;
assign n_28610 =  n_28608 &  n_28609;
assign n_28611 =  n_28607 &  n_28610;
assign n_28612 =  n_28604 &  n_28611;
assign n_28613 =  n_28542 &  n_28612;
assign n_28614 =  n_28520 &  n_28613;
assign n_28615 =  n_26477 &  n_26492;
assign n_28616 =  n_26490 &  n_28615;
assign n_28617 = ~n_25695 & ~n_25274;
assign n_28618 =  n_27341 &  n_27987;
assign n_28619 =  n_28617 &  n_28618;
assign n_28620 =  n_28616 &  n_28619;
assign n_28621 =  n_27161 & ~n_27150;
assign n_28622 = ~n_25682 &  n_26397;
assign n_28623 = ~n_25696 &  n_25697;
assign n_28624 = ~n_28623 & ~n_25684;
assign n_28625 = ~n_28622 &  n_28624;
assign n_28626 =  n_28621 &  n_28625;
assign n_28627 =  n_28620 &  n_28626;
assign n_28628 = ~n_23593 &  n_27938;
assign n_28629 =  n_28190 &  n_24528;
assign n_28630 =  n_28628 &  n_28629;
assign n_28631 =  n_26143 &  n_27186;
assign n_28632 =  n_26182 & ~n_28191;
assign n_28633 =  n_28631 &  n_28632;
assign n_28634 =  n_28630 &  n_28633;
assign n_28635 =  n_26202 &  n_26944;
assign n_28636 =  n_27977 &  n_28635;
assign n_28637 =  n_24565 &  n_26188;
assign n_28638 =  n_27940 &  n_28637;
assign n_28639 =  n_28636 &  n_28638;
assign n_28640 =  n_28634 &  n_28639;
assign n_28641 = ~n_23598 & ~n_23473;
assign n_28642 =  n_1175 &  n_1503;
assign n_28643 = ~n_25931 & ~n_22210;
assign n_28644 = ~n_28642 &  n_28643;
assign n_28645 = ~n_27072 &  n_28644;
assign n_28646 =  n_28641 &  n_28645;
assign n_28647 = ~n_27001 & ~n_24991;
assign n_28648 =  n_26316 &  n_28647;
assign n_28649 =  n_26148 &  n_28648;
assign n_28650 =  n_28646 &  n_28649;
assign n_28651 = ~n_26298 & ~n_22465;
assign n_28652 =  n_24695 &  n_28651;
assign n_28653 =  n_3345 &  n_28219;
assign n_28654 =  n_28652 &  n_28653;
assign n_28655 =  n_28650 &  n_28654;
assign n_28656 =  n_26704 & ~n_26139;
assign n_28657 =  n_28044 & ~n_28049;
assign n_28658 =  n_28656 &  n_28657;
assign n_28659 = ~n_23938 &  n_23939;
assign n_28660 = ~n_28659 &  n_28299;
assign n_28661 =  n_27837 & ~n_1701;
assign n_28662 =  n_28660 &  n_28661;
assign n_28663 =  n_28658 &  n_28662;
assign n_28664 =  n_28655 &  n_28663;
assign n_28665 =  n_28640 &  n_28664;
assign n_28666 = ~n_26393 & ~n_28312;
assign n_28667 = ~n_23325 &  n_26719;
assign n_28668 =  n_2094 &  n_28528;
assign n_28669 = ~n_28668 & ~n_26429;
assign n_28670 = ~n_28667 &  n_28669;
assign n_28671 = ~n_27347 &  n_28670;
assign n_28672 =  n_28666 &  n_28671;
assign n_28673 =  n_24199 & ~n_27650;
assign n_28674 =  n_1894 &  n_25108;
assign n_28675 =  n_1895 &  n_25287;
assign n_28676 = ~n_28674 & ~n_28675;
assign n_28677 = ~n_1044 &  n_28676;
assign n_28678 = ~n_28673 &  n_28677;
assign n_28679 = ~n_23292 &  n_23293;
assign n_28680 = ~n_25848 & ~n_28679;
assign n_28681 =  n_28678 &  n_28680;
assign n_28682 = ~n_25555 & ~n_24754;
assign n_28683 = ~n_26861 &  n_28236;
assign n_28684 =  n_23999 &  n_28683;
assign n_28685 =  n_28682 &  n_28684;
assign n_28686 =  n_28681 &  n_28685;
assign n_28687 =  n_28672 &  n_28686;
assign n_28688 =  n_28665 &  n_28687;
assign n_28689 =  n_28627 &  n_28688;
assign n_28690 =  n_28614 &  n_28689;
assign n_28691 =  n_28361 &  n_28690;
assign n_28692 = ~n_22082 &  n_28691;
assign n_28693 =  x_38 & ~n_28692;
assign n_28694 = ~x_38 &  n_28692;
assign n_28695 = ~n_28693 & ~n_28694;
assign n_28696 =  n_28625 & ~n_26349;
assign n_28697 =  n_26726 &  n_28696;
assign n_28698 =  n_28670 & ~n_23327;
assign n_28699 =  n_26722 &  n_28698;
assign n_28700 =  n_28699 &  n_27156;
assign n_28701 =  n_27162 &  n_27897;
assign n_28702 =  n_28700 &  n_28701;
assign n_28703 =  n_26462 &  n_27334;
assign n_28704 =  n_25557 &  n_28703;
assign n_28705 = ~n_25268 & ~n_28312;
assign n_28706 =  n_23370 & ~n_25994;
assign n_28707 =  n_28706 &  n_28324;
assign n_28708 =  n_28705 &  n_28707;
assign n_28709 =  n_28704 &  n_28708;
assign n_28710 =  n_28260 &  n_24791;
assign n_28711 = ~n_27653 & ~n_25207;
assign n_28712 = ~n_5654 &  n_24026;
assign n_28713 = ~n_28712 &  n_26072;
assign n_28714 = ~n_27102 &  n_28713;
assign n_28715 =  n_28711 &  n_28714;
assign n_28716 =  n_28710 &  n_28715;
assign n_28717 =  n_26226 &  n_27345;
assign n_28718 =  n_26702 &  n_28717;
assign n_28719 =  n_28716 &  n_28718;
assign n_28720 =  n_28709 &  n_28719;
assign n_28721 =  n_28702 &  n_28720;
assign n_28722 =  n_28697 &  n_28721;
assign n_28723 =  n_28054 &  n_28539;
assign n_28724 =  n_28052 &  n_28723;
assign n_28725 =  n_26677 &  n_23101;
assign n_28726 =  n_26273 &  n_28540;
assign n_28727 =  n_28725 &  n_28726;
assign n_28728 = ~n_26363 & ~n_24512;
assign n_28729 = ~n_26064 &  n_28728;
assign n_28730 =  n_25340 &  n_28729;
assign n_28731 =  n_28265 &  n_28730;
assign n_28732 =  n_26698 &  n_25025;
assign n_28733 = ~n_23014 & ~n_23809;
assign n_28734 = ~n_24801 &  n_28733;
assign n_28735 = ~n_28732 &  n_28734;
assign n_28736 =  n_28731 &  n_28735;
assign n_28737 =  n_553 &  n_12292;
assign n_28738 = ~n_25873 & ~n_28410;
assign n_28739 = ~n_23246 &  n_28738;
assign n_28740 = ~n_28737 &  n_28739;
assign n_28741 =  n_25872 &  n_28740;
assign n_28742 =  n_23677 &  n_27850;
assign n_28743 =  n_28741 &  n_28742;
assign n_28744 =  n_28743 &  n_27899;
assign n_28745 =  n_28736 &  n_28744;
assign n_28746 =  n_28727 &  n_28745;
assign n_28747 =  n_28724 &  n_28746;
assign n_28748 =  n_17783 &  n_27921;
assign n_28749 = ~n_28106 & ~n_28748;
assign n_28750 = ~n_27838 & ~n_27040;
assign n_28751 =  n_28749 &  n_28750;
assign n_28752 = ~n_23463 & ~n_23053;
assign n_28753 = ~n_26333 & ~n_24077;
assign n_28754 =  n_28752 &  n_28753;
assign n_28755 =  n_28751 &  n_28754;
assign n_28756 = ~n_349 &  n_26008;
assign n_28757 = ~n_20597 & ~n_28756;
assign n_28758 =  n_9689 &  n_6526;
assign n_28759 = ~n_28758 & ~n_25591;
assign n_28760 =  n_28757 &  n_28759;
assign n_28761 = ~n_28297 & ~n_28300;
assign n_28762 = ~n_23771 & ~n_26131;
assign n_28763 =  n_28761 &  n_28762;
assign n_28764 =  n_28760 &  n_28763;
assign n_28765 =  n_28755 &  n_28764;
assign n_28766 = ~n_23423 & ~n_25166;
assign n_28767 = ~n_25939 & ~n_24916;
assign n_28768 =  n_28766 &  n_28767;
assign n_28769 = ~n_25167 & ~n_27909;
assign n_28770 = ~n_25922 & ~n_24899;
assign n_28771 =  n_28769 &  n_28770;
assign n_28772 =  n_28768 &  n_28771;
assign n_28773 = ~n_24696 & ~n_18109;
assign n_28774 = ~n_24592 & ~n_23058;
assign n_28775 =  n_28773 &  n_28774;
assign n_28776 =  n_23613 &  n_13866;
assign n_28777 = ~n_28776 & ~n_25045;
assign n_28778 = ~n_24231 & ~n_20078;
assign n_28779 =  n_28777 &  n_28778;
assign n_28780 =  n_28775 &  n_28779;
assign n_28781 =  n_28772 &  n_28780;
assign n_28782 =  n_28765 &  n_28781;
assign n_28783 = ~n_27132 & ~n_26683;
assign n_28784 =  n_28783 &  n_27967;
assign n_28785 = ~n_4291 & ~n_25558;
assign n_28786 =  n_26346 &  n_28785;
assign n_28787 =  n_28784 &  n_28786;
assign n_28788 = ~n_24946 & ~n_26286;
assign n_28789 = ~n_24758 &  n_28788;
assign n_28790 =  n_1173 &  n_6876;
assign n_28791 = ~n_9884 & ~n_24569;
assign n_28792 = ~n_5981 &  n_28791;
assign n_28793 =  n_20596 & ~n_28792;
assign n_28794 = ~n_28790 & ~n_28793;
assign n_28795 = ~n_8366 & ~n_16882;
assign n_28796 =  n_28794 &  n_28795;
assign n_28797 =  n_28789 &  n_28796;
assign n_28798 = ~n_24951 &  n_26088;
assign n_28799 =  n_25159 &  n_13866;
assign n_28800 = ~n_25663 & ~n_28799;
assign n_28801 =  n_28798 &  n_28800;
assign n_28802 =  n_28797 &  n_28801;
assign n_28803 =  n_28787 &  n_28802;
assign n_28804 =  n_28782 &  n_28803;
assign n_28805 = ~n_27104 & ~n_26684;
assign n_28806 = ~n_17786 & ~n_26174;
assign n_28807 =  n_28805 &  n_28806;
assign n_28808 =  n_28216 & ~n_26948;
assign n_28809 = ~n_25905 & ~n_24060;
assign n_28810 = ~n_24009 & ~n_21178;
assign n_28811 =  n_28809 &  n_28810;
assign n_28812 =  n_28808 &  n_28811;
assign n_28813 =  n_28807 &  n_28812;
assign n_28814 = ~n_27937 &  n_23769;
assign n_28815 =  n_28468 &  n_28470;
assign n_28816 =  n_28814 &  n_28815;
assign n_28817 = ~n_24223 & ~n_24229;
assign n_28818 =  n_28817 &  n_26134;
assign n_28819 =  n_25083 &  n_28597;
assign n_28820 = ~n_9885 & ~n_28819;
assign n_28821 =  n_28818 &  n_28820;
assign n_28822 =  n_28816 &  n_28821;
assign n_28823 =  n_28813 &  n_28822;
assign n_28824 = ~n_26471 & ~n_28423;
assign n_28825 =  n_24017 &  n_23876;
assign n_28826 = ~n_27692 & ~n_28825;
assign n_28827 = ~n_26824 &  n_28826;
assign n_28828 =  n_28824 &  n_28827;
assign n_28829 =  x_42 &  n_28119;
assign n_28830 = ~n_28829 & ~n_27885;
assign n_28831 =  n_28828 &  n_28830;
assign n_28832 = ~n_25033 & ~n_25036;
assign n_28833 = ~n_23895 & ~n_6881;
assign n_28834 =  n_28832 &  n_28833;
assign n_28835 =  n_23987 &  n_24015;
assign n_28836 = ~n_28835 & ~n_25018;
assign n_28837 = ~n_23988 & ~n_25151;
assign n_28838 =  n_28836 &  n_28837;
assign n_28839 =  n_28834 &  n_28838;
assign n_28840 = ~n_23631 & ~n_27007;
assign n_28841 = ~n_23139 & ~n_27052;
assign n_28842 =  n_28840 &  n_28841;
assign n_28843 = ~n_26368 & ~n_3630;
assign n_28844 = ~n_3341 & ~n_152;
assign n_28845 = ~n_28844 &  n_2881;
assign n_28846 = ~n_28845 & ~n_3633;
assign n_28847 =  n_28843 &  n_28846;
assign n_28848 =  n_28842 &  n_28847;
assign n_28849 =  n_28839 &  n_28848;
assign n_28850 =  n_28831 &  n_28849;
assign n_28851 = ~n_26845 & ~n_28335;
assign n_28852 =  n_13866 &  n_23597;
assign n_28853 =  n_23842 & ~n_28852;
assign n_28854 =  n_28851 &  n_28853;
assign n_28855 =  n_1042 &  n_7467;
assign n_28856 = ~n_28855 &  n_24123;
assign n_28857 = ~n_25211 &  n_26241;
assign n_28858 =  n_28856 &  n_28857;
assign n_28859 =  n_28854 &  n_28858;
assign n_28860 =  n_28850 &  n_28859;
assign n_28861 =  n_28823 &  n_28860;
assign n_28862 =  n_28804 &  n_28861;
assign n_28863 = ~n_26171 & ~n_7856;
assign n_28864 = ~n_25980 & ~n_14261;
assign n_28865 =  n_28863 &  n_28864;
assign n_28866 = ~n_28188 & ~n_4292;
assign n_28867 = ~n_27338 &  n_28866;
assign n_28868 =  n_28865 &  n_28867;
assign n_28869 =  n_28240 &  n_28868;
assign n_28870 =  n_25347 &  n_27936;
assign n_28871 =  n_28185 &  n_28870;
assign n_28872 =  n_28869 &  n_28871;
assign n_28873 =  n_28438 & ~n_16302;
assign n_28874 = ~n_25660 &  n_28873;
assign n_28875 =  n_27971 &  n_28874;
assign n_28876 =  n_28523 &  n_28875;
assign n_28877 =  n_28872 &  n_28876;
assign n_28878 = ~n_25294 &  n_8357;
assign n_28879 =  n_26957 &  n_24524;
assign n_28880 =  n_28878 &  n_28879;
assign n_28881 = ~n_16110 &  n_28157;
assign n_28882 =  n_28291 &  n_28881;
assign n_28883 =  n_1894 &  n_556;
assign n_28884 =  n_24064 &  n_28883;
assign n_28885 =  x_42 &  n_28884;
assign n_28886 = ~n_26402 & ~n_23550;
assign n_28887 = ~n_28885 &  n_28886;
assign n_28888 = ~n_26074 & ~n_23764;
assign n_28889 =  n_28887 &  n_28888;
assign n_28890 =  n_28882 &  n_28889;
assign n_28891 =  n_28880 &  n_28890;
assign n_28892 =  n_28199 & ~n_24525;
assign n_28893 =  n_23830 &  n_23832;
assign n_28894 = ~n_28893 &  n_27265;
assign n_28895 =  n_28892 &  n_28894;
assign n_28896 =  n_28200 &  n_26958;
assign n_28897 =  n_27229 &  n_27916;
assign n_28898 =  n_28896 &  n_28897;
assign n_28899 =  n_28895 &  n_28898;
assign n_28900 =  n_28891 &  n_28899;
assign n_28901 =  n_28877 &  n_28900;
assign n_28902 =  n_28862 &  n_28901;
assign n_28903 =  n_28545 &  n_27126;
assign n_28904 =  n_23047 &  n_27150;
assign n_28905 = ~n_28904 &  n_26256;
assign n_28906 =  n_28903 &  n_28905;
assign n_28907 = ~n_26358 & ~n_28112;
assign n_28908 = ~n_25450 &  n_25451;
assign n_28909 =  n_23689 & ~n_28908;
assign n_28910 =  n_28907 &  n_28909;
assign n_28911 =  n_28910 &  n_28549;
assign n_28912 =  n_27097 &  n_26355;
assign n_28913 =  n_28911 &  n_28912;
assign n_28914 =  n_28906 &  n_28913;
assign n_28915 = ~x_43 &  n_25518;
assign n_28916 = ~n_28915 & ~n_24920;
assign n_28917 = ~n_26108 &  n_28916;
assign n_28918 =  n_24426 &  n_24427;
assign n_28919 = ~n_26283 & ~n_25491;
assign n_28920 =  n_26111 &  n_28919;
assign n_28921 = ~n_28918 &  n_28920;
assign n_28922 =  n_28676 &  n_28921;
assign n_28923 =  n_28917 &  n_28922;
assign n_28924 =  n_28555 &  n_27858;
assign n_28925 =  n_28553 &  n_28924;
assign n_28926 =  n_28923 &  n_28925;
assign n_28927 =  n_28914 &  n_28926;
assign n_28928 = ~n_24056 & ~n_25904;
assign n_28929 = ~n_25337 &  n_28928;
assign n_28930 =  n_5654 &  n_24936;
assign n_28931 = ~n_28930 & ~n_27695;
assign n_28932 = ~n_27131 &  n_28931;
assign n_28933 =  n_28929 &  n_28932;
assign n_28934 = ~n_25985 & ~n_25084;
assign n_28935 = ~n_27874 & ~n_6527;
assign n_28936 =  n_28934 &  n_28935;
assign n_28937 = ~n_23946 &  n_28936;
assign n_28938 =  n_25282 &  n_26148;
assign n_28939 =  n_28937 &  n_28938;
assign n_28940 =  n_28933 &  n_28939;
assign n_28941 =  n_26310 &  n_28134;
assign n_28942 =  n_28373 &  n_26876;
assign n_28943 =  n_28941 &  n_28942;
assign n_28944 =  n_28471 &  n_27601;
assign n_28945 =  n_26312 &  n_3627;
assign n_28946 =  n_28944 &  n_28945;
assign n_28947 =  n_28943 &  n_28946;
assign n_28948 =  n_26263 &  n_25174;
assign n_28949 =  n_23595 & ~n_25589;
assign n_28950 = ~n_28949 & ~n_23726;
assign n_28951 =  n_28135 &  n_28950;
assign n_28952 =  n_28948 &  n_28951;
assign n_28953 =  n_28947 &  n_28952;
assign n_28954 =  n_28940 &  n_28953;
assign n_28955 = ~n_24777 &  n_28317;
assign n_28956 = ~n_28659 & ~n_27185;
assign n_28957 =  n_28956 &  n_27901;
assign n_28958 =  n_28955 &  n_28957;
assign n_28959 = ~n_27881 &  n_28172;
assign n_28960 = ~n_26315 &  n_28959;
assign n_28961 = ~n_26154 & ~n_27128;
assign n_28962 =  n_28960 &  n_28961;
assign n_28963 =  n_27919 &  n_28155;
assign n_28964 =  n_28963 &  n_28004;
assign n_28965 =  n_28962 &  n_28964;
assign n_28966 =  n_28958 &  n_28965;
assign n_28967 =  n_28954 &  n_28966;
assign n_28968 =  n_28927 &  n_28967;
assign n_28969 =  n_28902 &  n_28968;
assign n_28970 =  n_28747 &  n_28969;
assign n_28971 =  n_28722 &  n_28970;
assign n_28972 = ~n_27491 &  n_28971;
assign n_28973 = ~n_22082 &  n_28972;
assign n_28974 = ~n_25844 &  n_28973;
assign n_28975 =  x_37 & ~n_28974;
assign n_28976 = ~x_37 &  n_28974;
assign n_28977 = ~n_28975 & ~n_28976;
assign n_28978 = ~n_26196 & ~n_24750;
assign n_28979 =  n_25252 &  n_28978;
assign n_28980 = ~n_28218 & ~n_3348;
assign n_28981 = ~n_25657 &  n_28980;
assign n_28982 =  n_26937 &  n_28981;
assign n_28983 =  n_28979 &  n_28982;
assign n_28984 =  n_24697 &  n_28983;
assign n_28985 =  n_28984 &  n_27846;
assign n_28986 =  n_26717 &  n_28743;
assign n_28987 =  n_28985 &  n_28986;
assign n_28988 =  n_28910 &  n_27855;
assign n_28989 =  n_27096 &  n_28530;
assign n_28990 =  n_28988 &  n_28989;
assign n_28991 =  n_28956 &  n_28560;
assign n_28992 =  n_28562 &  n_28566;
assign n_28993 =  n_28991 &  n_28992;
assign n_28994 =  n_28990 &  n_28993;
assign n_28995 =  n_25295 &  n_25291;
assign n_28996 =  n_28601 &  n_28995;
assign n_28997 =  n_27830 &  n_28996;
assign n_28998 =  n_28994 &  n_28997;
assign n_28999 =  n_24532 &  n_24563;
assign n_29000 =  n_27765 & ~n_28999;
assign n_29001 = ~n_28819 &  n_29000;
assign n_29002 =  n_26873 &  n_28141;
assign n_29003 =  n_26307 & ~n_23177;
assign n_29004 =  n_29002 &  n_29003;
assign n_29005 =  n_29001 &  n_29004;
assign n_29006 = ~n_26451 & ~n_24516;
assign n_29007 = ~n_26352 &  n_29006;
assign n_29008 = ~n_23880 & ~n_26371;
assign n_29009 =  n_29007 &  n_29008;
assign n_29010 =  n_29005 &  n_29009;
assign n_29011 = ~n_26483 &  n_28174;
assign n_29012 =  n_28178 & ~n_24523;
assign n_29013 =  n_29011 &  n_29012;
assign n_29014 = ~n_26315 &  n_28157;
assign n_29015 =  n_27089 &  n_26319;
assign n_29016 =  n_29014 &  n_29015;
assign n_29017 =  n_29013 &  n_29016;
assign n_29018 =  n_28817 &  n_26487;
assign n_29019 =  n_29018 &  n_28168;
assign n_29020 = ~n_20984 & ~n_14786;
assign n_29021 = ~n_26426 & ~n_28154;
assign n_29022 =  n_28169 &  n_29021;
assign n_29023 =  n_29020 &  n_29022;
assign n_29024 =  n_29019 &  n_29023;
assign n_29025 =  n_29017 &  n_29024;
assign n_29026 =  n_29010 &  n_29025;
assign n_29027 = ~n_26969 &  n_26741;
assign n_29028 =  n_29027 & ~n_23620;
assign n_29029 =  n_28303 &  n_23368;
assign n_29030 =  n_29028 &  n_29029;
assign n_29031 =  n_24305 &  n_24791;
assign n_29032 = ~n_27102 & ~n_25851;
assign n_29033 =  n_29031 &  n_29032;
assign n_29034 =  n_29030 &  n_29033;
assign n_29035 =  n_29026 &  n_29034;
assign n_29036 =  n_28998 &  n_29035;
assign n_29037 =  n_28987 &  n_29036;
assign n_29038 = ~n_26394 &  n_27999;
assign n_29039 =  n_23015 &  n_29038;
assign n_29040 =  n_29039 &  n_28699;
assign n_29041 =  n_27904 &  n_29040;
assign n_29042 =  n_27719 & ~n_23771;
assign n_29043 =  n_1175 &  n_8053;
assign n_29044 = ~n_25348 & ~n_29043;
assign n_29045 =  n_29042 &  n_29044;
assign n_29046 = ~n_21565 & ~n_13286;
assign n_29047 =  n_25159 &  n_28883;
assign n_29048 =  n_8365 &  n_13230;
assign n_29049 = ~n_29047 & ~n_29048;
assign n_29050 =  n_29046 &  n_29049;
assign n_29051 =  n_29045 &  n_29050;
assign n_29052 = ~x_43 &  n_10477;
assign n_29053 =  n_24969 &  n_29052;
assign n_29054 = ~n_29053 & ~n_25169;
assign n_29055 = ~n_24947 &  n_29054;
assign n_29056 = ~n_26091 & ~n_26335;
assign n_29057 =  n_29055 &  n_29056;
assign n_29058 =  n_29051 &  n_29057;
assign n_29059 = ~n_24319 & ~n_3343;
assign n_29060 = ~n_5983 & ~n_14261;
assign n_29061 =  n_29059 &  n_29060;
assign n_29062 = ~n_25936 & ~n_25382;
assign n_29063 = ~n_23386 & ~n_26086;
assign n_29064 =  n_29062 &  n_29063;
assign n_29065 =  n_29061 &  n_29064;
assign n_29066 = ~n_26732 & ~n_26962;
assign n_29067 = ~n_23541 & ~n_24503;
assign n_29068 =  n_29066 &  n_29067;
assign n_29069 = ~n_24571 & ~n_21759;
assign n_29070 = ~n_23477 & ~n_25236;
assign n_29071 =  n_29069 &  n_29070;
assign n_29072 =  n_29068 &  n_29071;
assign n_29073 =  n_29065 &  n_29072;
assign n_29074 =  n_29058 &  n_29073;
assign n_29075 =  n_27967 & ~n_26231;
assign n_29076 =  n_28936 &  n_26227;
assign n_29077 =  n_29075 &  n_29076;
assign n_29078 = ~n_23839 & ~n_24937;
assign n_29079 = ~n_24950 & ~n_25097;
assign n_29080 = ~n_25890 &  n_29079;
assign n_29081 =  n_29078 &  n_29080;
assign n_29082 = ~n_26102 & ~n_26431;
assign n_29083 = ~n_24358 &  n_29082;
assign n_29084 =  n_29081 &  n_29083;
assign n_29085 =  n_29077 &  n_29084;
assign n_29086 =  n_29074 &  n_29085;
assign n_29087 =  n_28809 &  n_26069;
assign n_29088 = ~n_26311 & ~n_26975;
assign n_29089 = ~n_26373 &  n_29088;
assign n_29090 =  n_29087 &  n_29089;
assign n_29091 =  n_24228 & ~n_26474;
assign n_29092 = ~n_27974 & ~n_27820;
assign n_29093 =  n_29091 &  n_29092;
assign n_29094 =  n_29090 &  n_29093;
assign n_29095 = ~n_27104 & ~n_27072;
assign n_29096 =  n_26031 & ~n_26938;
assign n_29097 =  n_29095 &  n_29096;
assign n_29098 = ~n_24940 & ~n_25900;
assign n_29099 =  n_29098 &  n_26737;
assign n_29100 = ~n_25239 & ~n_26141;
assign n_29101 =  n_29100 & ~n_23951;
assign n_29102 =  n_29099 &  n_29101;
assign n_29103 =  n_29097 &  n_29102;
assign n_29104 =  n_29094 &  n_29103;
assign n_29105 =  n_23252 &  n_23881;
assign n_29106 = ~n_26178 & ~n_29105;
assign n_29107 = ~n_27003 &  n_29106;
assign n_29108 = ~n_27007 & ~n_25047;
assign n_29109 = ~n_23179 & ~n_24582;
assign n_29110 =  n_29108 &  n_29109;
assign n_29111 =  n_29107 &  n_29110;
assign n_29112 =  n_28824 & ~n_25663;
assign n_29113 =  n_29111 &  n_29112;
assign n_29114 = ~n_24899 & ~n_27283;
assign n_29115 = ~n_28119 & ~n_24210;
assign n_29116 =  n_29114 &  n_29115;
assign n_29117 = ~n_25032 & ~n_25490;
assign n_29118 = ~n_24122 & ~n_10;
assign n_29119 =  n_29117 &  n_29118;
assign n_29120 = ~n_23988 & ~n_24686;
assign n_29121 = ~n_25093 &  n_29120;
assign n_29122 =  n_29119 &  n_29121;
assign n_29123 =  n_29116 &  n_29122;
assign n_29124 =  n_29113 &  n_29123;
assign n_29125 = ~n_26330 & ~n_28498;
assign n_29126 = ~n_27075 &  n_29125;
assign n_29127 =  n_29126 &  n_23886;
assign n_29128 = ~n_26843 &  n_26362;
assign n_29129 =  n_29127 &  n_29128;
assign n_29130 =  n_13866 &  n_25520;
assign n_29131 = ~n_29130 & ~n_24161;
assign n_29132 = ~n_25033 & ~n_24527;
assign n_29133 = ~n_26836 &  n_29132;
assign n_29134 =  n_29133 &  n_26120;
assign n_29135 =  n_29131 &  n_29134;
assign n_29136 =  n_29129 &  n_29135;
assign n_29137 =  n_29124 &  n_29136;
assign n_29138 =  n_29104 &  n_29137;
assign n_29139 =  n_29086 &  n_29138;
assign n_29140 =  n_28711 &  n_28706;
assign n_29141 =  n_27333 &  n_29140;
assign n_29142 =  x_42 &  n_28048;
assign n_29143 = ~n_29142 &  n_26132;
assign n_29144 =  n_27924 &  n_27882;
assign n_29145 =  n_29143 &  n_29144;
assign n_29146 = ~n_27699 & ~n_25982;
assign n_29147 =  n_28047 &  n_29146;
assign n_29148 =  n_28008 &  n_28236;
assign n_29149 =  n_29147 &  n_29148;
assign n_29150 =  n_29145 &  n_29149;
assign n_29151 =  n_28888 &  n_26970;
assign n_29152 =  n_23948 &  n_29151;
assign n_29153 =  n_27913 &  n_26137;
assign n_29154 =  n_28196 &  n_27914;
assign n_29155 =  n_29153 &  n_29154;
assign n_29156 =  n_29152 &  n_29155;
assign n_29157 =  n_29150 &  n_29156;
assign n_29158 =  n_29141 &  n_29157;
assign n_29159 =  n_29139 &  n_29158;
assign n_29160 =  n_29041 &  n_29159;
assign n_29161 = ~n_11 &  n_25116;
assign n_29162 = ~n_26889 & ~n_29161;
assign n_29163 =  n_28648 &  n_29162;
assign n_29164 = ~n_25268 &  n_29163;
assign n_29165 = ~n_27347 &  n_29164;
assign n_29166 =  n_27159 &  n_29165;
assign n_29167 =  n_28621 &  n_28314;
assign n_29168 =  n_29166 &  n_29167;
assign n_29169 =  n_29168 &  n_28697;
assign n_29170 =  n_29160 &  n_29169;
assign n_29171 =  n_29037 &  n_29170;
assign n_29172 = ~n_22939 &  n_29171;
assign n_29173 = ~n_25845 &  n_29172;
assign n_29174 =  n_28035 &  n_29173;
assign n_29175 =  n_28031 &  n_29174;
assign n_29176 =  x_36 & ~n_29175;
assign n_29177 = ~x_36 &  n_29175;
assign n_29178 = ~n_29176 & ~n_29177;
assign n_29179 = ~n_26638 &  n_25717;
assign n_29180 = ~n_27998 & ~n_25851;
assign n_29181 =  n_27106 &  n_28937;
assign n_29182 =  n_29180 &  n_29181;
assign n_29183 =  n_25233 & ~n_27754;
assign n_29184 = ~n_23643 &  n_29183;
assign n_29185 =  n_27758 &  n_28457;
assign n_29186 =  n_26028 &  n_27071;
assign n_29187 =  n_29185 &  n_29186;
assign n_29188 =  n_29184 &  n_29187;
assign n_29189 = ~n_29130 & ~n_24670;
assign n_29190 = ~n_26080 &  n_29189;
assign n_29191 = ~n_26468 & ~n_26018;
assign n_29192 = ~n_26467 &  n_29191;
assign n_29193 =  n_29190 &  n_29192;
assign n_29194 =  n_29188 &  n_29193;
assign n_29195 =  n_29182 &  n_29194;
assign n_29196 =  n_28963 &  n_29027;
assign n_29197 =  n_25872 &  n_28294;
assign n_29198 =  n_29196 &  n_29197;
assign n_29199 =  n_28389 &  n_24768;
assign n_29200 =  n_28938 &  n_28263;
assign n_29201 =  n_29199 &  n_29200;
assign n_29202 =  n_29198 &  n_29201;
assign n_29203 =  n_29195 &  n_29202;
assign n_29204 = ~n_24701 & ~n_24946;
assign n_29205 = ~n_28419 & ~n_26184;
assign n_29206 =  n_29204 &  n_29205;
assign n_29207 = ~n_25490 & ~n_25083;
assign n_29208 = ~n_25500 &  n_29207;
assign n_29209 = ~n_28119 & ~n_24629;
assign n_29210 =  n_29208 &  n_29209;
assign n_29211 =  n_29206 &  n_29210;
assign n_29212 = ~x_1771 &  n_24631;
assign n_29213 = ~n_29212 & ~n_27852;
assign n_29214 = ~n_25986 & ~n_26311;
assign n_29215 =  n_29213 &  n_29214;
assign n_29216 = ~n_24950 & ~n_24685;
assign n_29217 = ~n_24982 & ~n_3343;
assign n_29218 =  n_29216 &  n_29217;
assign n_29219 =  n_29215 &  n_29218;
assign n_29220 =  n_29211 &  n_29219;
assign n_29221 =  x_588 &  n_25936;
assign n_29222 = ~n_29221 &  n_28554;
assign n_29223 = ~n_26201 & ~n_27284;
assign n_29224 =  n_29222 &  n_29223;
assign n_29225 = ~n_23245 & ~n_28845;
assign n_29226 = ~n_24595 & ~n_28175;
assign n_29227 =  n_29225 &  n_29226;
assign n_29228 =  n_3341 &  n_3629;
assign n_29229 = ~n_29228 & ~n_25651;
assign n_29230 =  n_8361 &  n_10867;
assign n_29231 = ~n_25027 & ~n_29230;
assign n_29232 =  n_29229 &  n_29231;
assign n_29233 =  n_29227 &  n_29232;
assign n_29234 =  n_25017 & ~n_27819;
assign n_29235 = ~n_24532 & ~n_23694;
assign n_29236 = ~n_27079 &  n_29235;
assign n_29237 = ~n_29234 &  n_29236;
assign n_29238 =  n_29233 &  n_29237;
assign n_29239 =  n_29224 &  n_29238;
assign n_29240 =  n_29220 &  n_29239;
assign n_29241 = ~n_24959 & ~n_14656;
assign n_29242 =  n_29006 &  n_29241;
assign n_29243 = ~n_24872 & ~n_27230;
assign n_29244 =  n_28327 &  n_29243;
assign n_29245 =  n_29242 &  n_29244;
assign n_29246 = ~n_14265 & ~n_28106;
assign n_29247 = ~n_3631 & ~n_24076;
assign n_29248 =  n_29246 &  n_29247;
assign n_29249 = ~n_25296 & ~n_26333;
assign n_29250 = ~n_24571 & ~n_27188;
assign n_29251 =  n_29249 &  n_29250;
assign n_29252 =  n_29248 &  n_29251;
assign n_29253 =  n_28413 & ~n_27040;
assign n_29254 =  n_1 &  n_24073;
assign n_29255 = ~n_29254 & ~n_25997;
assign n_29256 =  n_29253 &  n_29255;
assign n_29257 = ~n_25641 & ~n_10871;
assign n_29258 = ~n_24503 & ~n_28748;
assign n_29259 =  n_29257 &  n_29258;
assign n_29260 =  n_29256 &  n_29259;
assign n_29261 =  n_29252 &  n_29260;
assign n_29262 =  n_29245 &  n_29261;
assign n_29263 =  n_29240 &  n_29262;
assign n_29264 = ~n_25874 &  n_28599;
assign n_29265 =  n_29264 &  n_25241;
assign n_29266 =  n_28464 &  n_28810;
assign n_29267 =  n_27123 & ~n_25452;
assign n_29268 =  n_29266 &  n_29267;
assign n_29269 =  n_29265 &  n_29268;
assign n_29270 =  n_26437 & ~n_10472;
assign n_29271 =  n_24522 & ~n_26459;
assign n_29272 =  n_29270 &  n_29271;
assign n_29273 =  n_27923 &  n_26733;
assign n_29274 = ~n_26684 &  n_25228;
assign n_29275 =  n_29273 &  n_29274;
assign n_29276 =  n_29272 &  n_29275;
assign n_29277 =  n_29269 &  n_29276;
assign n_29278 =  n_24316 & ~n_24937;
assign n_29279 = ~n_22721 &  n_26011;
assign n_29280 =  n_29278 &  n_29279;
assign n_29281 =  n_26206 & ~n_24161;
assign n_29282 = ~n_25213 & ~n_25918;
assign n_29283 =  n_29282 &  n_24126;
assign n_29284 =  n_29281 &  n_29283;
assign n_29285 =  n_29280 &  n_29284;
assign n_29286 = ~n_23544 & ~n_23732;
assign n_29287 =  n_29286 & ~n_27873;
assign n_29288 =  n_23944 &  n_26711;
assign n_29289 =  n_29287 &  n_29288;
assign n_29290 =  n_24683 & ~n_26373;
assign n_29291 = ~n_2686 & ~n_25864;
assign n_29292 =  n_29291 & ~n_27132;
assign n_29293 =  n_29290 &  n_29292;
assign n_29294 =  n_29289 &  n_29293;
assign n_29295 =  n_29285 &  n_29294;
assign n_29296 =  n_29277 &  n_29295;
assign n_29297 =  n_29263 &  n_29296;
assign n_29298 =  n_29203 &  n_29297;
assign n_29299 =  n_28524 & ~n_27492;
assign n_29300 =  n_28731 &  n_26695;
assign n_29301 =  n_29299 &  n_29300;
assign n_29302 = ~n_25289 &  n_26705;
assign n_29303 =  n_29302 &  n_29087;
assign n_29304 =  n_28217 &  n_29303;
assign n_29305 =  n_24785 &  n_29304;
assign n_29306 =  n_27092 &  n_28392;
assign n_29307 =  n_28962 &  n_29306;
assign n_29308 =  n_29305 &  n_29307;
assign n_29309 =  n_28735 &  n_28984;
assign n_29310 =  n_29308 &  n_29309;
assign n_29311 =  n_29301 &  n_29310;
assign n_29312 =  n_29298 &  n_29311;
assign n_29313 =  n_28682 &  n_28006;
assign n_29314 =  n_28015 &  n_28319;
assign n_29315 =  n_29313 &  n_29314;
assign n_29316 =  n_26384 &  n_29315;
assign n_29317 =  n_28718 &  n_29316;
assign n_29318 =  n_28881 &  n_26158;
assign n_29319 =  n_28887 &  n_29318;
assign n_29320 = ~n_18302 &  n_28235;
assign n_29321 =  n_27125 &  n_26480;
assign n_29322 =  n_29320 &  n_29321;
assign n_29323 =  n_29319 &  n_29322;
assign n_29324 = ~n_26163 & ~n_27619;
assign n_29325 =  n_27670 &  n_29324;
assign n_29326 =  n_29325 &  n_28710;
assign n_29327 =  n_29323 &  n_29326;
assign n_29328 =  n_28242 &  n_26939;
assign n_29329 =  n_28561 &  n_23996;
assign n_29330 =  n_29328 &  n_29329;
assign n_29331 =  n_24225 &  n_26944;
assign n_29332 = ~n_27651 &  n_28645;
assign n_29333 =  n_29331 &  n_29332;
assign n_29334 =  n_29330 &  n_29333;
assign n_29335 =  n_28047 &  n_26961;
assign n_29336 =  n_26151 & ~n_27494;
assign n_29337 =  n_29335 &  n_29336;
assign n_29338 = ~n_27331 &  n_26965;
assign n_29339 =  n_26227 &  n_29146;
assign n_29340 =  n_29338 &  n_29339;
assign n_29341 =  n_29337 &  n_29340;
assign n_29342 =  n_29334 &  n_29341;
assign n_29343 =  n_29327 &  n_29342;
assign n_29344 =  n_28680 &  n_25674;
assign n_29345 =  n_28875 &  n_28684;
assign n_29346 =  n_29344 &  n_29345;
assign n_29347 = ~n_26486 & ~n_23983;
assign n_29348 =  n_27657 &  n_29347;
assign n_29349 = ~n_23008 &  n_29348;
assign n_29350 = ~n_26394 &  n_29349;
assign n_29351 =  n_29346 &  n_29350;
assign n_29352 =  n_29343 &  n_29351;
assign n_29353 =  n_29317 &  n_29352;
assign n_29354 =  n_29168 &  n_29353;
assign n_29355 =  n_29312 &  n_29354;
assign n_29356 = ~n_25845 &  n_29355;
assign n_29357 = ~n_25844 &  n_29356;
assign n_29358 =  n_29179 &  n_29357;
assign n_29359 =  n_26636 &  n_29358;
assign n_29360 =  x_35 & ~n_29359;
assign n_29361 = ~x_35 &  n_29359;
assign n_29362 = ~n_29360 & ~n_29361;
assign n_29363 =  n_28917 &  n_28396;
assign n_29364 =  n_29192 &  n_28279;
assign n_29365 =  n_29363 &  n_29364;
assign n_29366 = ~n_27116 & ~n_26336;
assign n_29367 = ~n_28048 &  n_29366;
assign n_29368 = ~n_24754 &  n_29367;
assign n_29369 = ~n_26083 & ~n_27012;
assign n_29370 = ~n_24117 &  n_29369;
assign n_29371 =  n_23995 &  n_23892;
assign n_29372 =  n_29370 &  n_29371;
assign n_29373 =  n_29368 &  n_29372;
assign n_29374 =  n_29365 &  n_29373;
assign n_29375 =  n_28929 &  n_26370;
assign n_29376 =  n_26344 &  n_28932;
assign n_29377 =  n_29375 &  n_29376;
assign n_29378 =  n_24692 &  n_24697;
assign n_29379 =  n_26375 &  n_28948;
assign n_29380 =  n_29378 &  n_29379;
assign n_29381 =  n_29377 &  n_29380;
assign n_29382 =  n_29374 &  n_29381;
assign n_29383 =  n_8354 &  n_27921;
assign n_29384 = ~n_29383 & ~n_25116;
assign n_29385 = ~n_23463 & ~n_26485;
assign n_29386 =  n_29384 &  n_29385;
assign n_29387 = ~n_26436 & ~n_29212;
assign n_29388 = ~n_23468 & ~n_23595;
assign n_29389 =  n_29387 &  n_29388;
assign n_29390 =  n_29386 &  n_29389;
assign n_29391 =  n_24931 & ~n_23686;
assign n_29392 =  n_29391 & ~n_27175;
assign n_29393 =  n_29390 &  n_29392;
assign n_29394 = ~n_23615 & ~n_25491;
assign n_29395 = ~n_24230 & ~n_7468;
assign n_29396 =  n_29394 &  n_29395;
assign n_29397 = ~n_1901 & ~n_26350;
assign n_29398 =  n_29396 &  n_29397;
assign n_29399 = ~n_23331 & ~n_25226;
assign n_29400 = ~n_3145 & ~n_25083;
assign n_29401 = ~n_27290 &  n_29400;
assign n_29402 =  n_29399 &  n_29401;
assign n_29403 =  n_29398 &  n_29402;
assign n_29404 = ~n_28041 & ~n_23821;
assign n_29405 = ~n_24229 & ~n_23997;
assign n_29406 =  n_29404 &  n_29405;
assign n_29407 = ~n_25157 & ~n_24201;
assign n_29408 = ~n_25382 & ~n_24932;
assign n_29409 =  n_29407 &  n_29408;
assign n_29410 =  n_29406 &  n_29409;
assign n_29411 =  n_29403 &  n_29410;
assign n_29412 =  n_29393 &  n_29411;
assign n_29413 =  n_23903 &  n_29082;
assign n_29414 =  n_29413 &  n_23854;
assign n_29415 =  n_26943 &  n_28439;
assign n_29416 =  n_27949 &  n_29415;
assign n_29417 =  n_29414 &  n_29416;
assign n_29418 =  n_29412 &  n_29417;
assign n_29419 =  n_29286 & ~n_27111;
assign n_29420 =  n_25172 &  n_29419;
assign n_29421 =  n_28290 &  n_27786;
assign n_29422 =  n_28461 & ~n_25277;
assign n_29423 =  n_29421 &  n_29422;
assign n_29424 =  n_29420 &  n_29423;
assign n_29425 =  n_25248 & ~n_27757;
assign n_29426 =  n_29100 &  n_29425;
assign n_29427 =  n_28531 &  n_29426;
assign n_29428 =  n_29424 &  n_29427;
assign n_29429 =  n_26840 & ~n_26007;
assign n_29430 = ~n_23561 & ~n_28852;
assign n_29431 =  n_29429 &  n_29430;
assign n_29432 =  n_349 &  n_26185;
assign n_29433 = ~n_29432 & ~n_25922;
assign n_29434 = ~n_25105 & ~n_27679;
assign n_29435 =  n_29433 &  n_29434;
assign n_29436 = ~n_24839 &  n_26837;
assign n_29437 =  n_29435 &  n_29436;
assign n_29438 =  n_29431 &  n_29437;
assign n_29439 = ~n_23613 & ~n_25159;
assign n_29440 =  n_28883 & ~n_29439;
assign n_29441 = ~n_29440 &  n_29098;
assign n_29442 =  n_26737 & ~n_27873;
assign n_29443 =  n_29441 &  n_29442;
assign n_29444 = ~n_25275 &  n_25276;
assign n_29445 = ~n_27853 & ~n_29444;
assign n_29446 =  n_29088 &  n_29291;
assign n_29447 =  n_29445 &  n_29446;
assign n_29448 =  n_29443 &  n_29447;
assign n_29449 =  n_29438 &  n_29448;
assign n_29450 =  n_29428 &  n_29449;
assign n_29451 =  n_29418 &  n_29450;
assign n_29452 =  n_29382 &  n_29451;
assign n_29453 =  n_27656 &  n_26347;
assign n_29454 =  n_24799 &  n_29453;
assign n_29455 =  n_29305 &  n_29454;
assign n_29456 =  n_27830 &  n_23064;
assign n_29457 =  n_29455 &  n_29456;
assign n_29458 =  n_27505 &  n_29457;
assign n_29459 =  n_29452 &  n_29458;
assign n_29460 =  n_29039 &  n_25694;
assign n_29461 =  n_28343 &  n_29460;
assign n_29462 =  n_28338 &  n_27182;
assign n_29463 =  n_28339 & ~n_24432;
assign n_29464 =  n_29462 &  n_29463;
assign n_29465 =  n_26933 &  n_3345;
assign n_29466 =  n_27969 &  n_27337;
assign n_29467 =  n_29465 &  n_29466;
assign n_29468 =  n_26950 &  n_28651;
assign n_29469 =  n_28784 &  n_29468;
assign n_29470 =  n_29467 &  n_29469;
assign n_29471 =  n_28219 &  n_28641;
assign n_29472 =  x_1547 &  n_26091;
assign n_29473 =  n_28785 & ~n_29472;
assign n_29474 =  n_29471 &  n_29473;
assign n_29475 =  n_28636 &  n_29474;
assign n_29476 =  n_29470 &  n_29475;
assign n_29477 =  n_29464 &  n_29476;
assign n_29478 =  n_23831 &  n_28869;
assign n_29479 =  n_29348 &  n_28678;
assign n_29480 =  n_29478 &  n_29479;
assign n_29481 =  n_28716 &  n_29480;
assign n_29482 =  n_29477 &  n_29481;
assign n_29483 =  n_29461 &  n_29482;
assign n_29484 =  n_29459 &  n_29483;
assign n_29485 =  x_34 & ~n_29484;
assign n_29486 = ~x_34 &  n_29484;
assign n_29487 = ~n_29485 & ~n_29486;
assign n_29488 =  n_24235 &  n_26421;
assign n_29489 =  n_24323 &  n_29325;
assign n_29490 =  n_29488 &  n_29489;
assign n_29491 =  n_29078 &  n_28536;
assign n_29492 =  n_27975 &  n_29491;
assign n_29493 =  n_29391 &  n_29080;
assign n_29494 =  n_27950 &  n_26219;
assign n_29495 =  n_29493 &  n_29494;
assign n_29496 =  n_29492 &  n_29495;
assign n_29497 =  n_27179 &  n_28330;
assign n_29498 =  n_29496 &  n_29497;
assign n_29499 =  n_29490 &  n_29498;
assign n_29500 =  n_27149 &  n_29499;
assign n_29501 =  n_29282 &  n_29133;
assign n_29502 =  n_29126 &  n_26819;
assign n_29503 =  n_29501 &  n_29502;
assign n_29504 =  n_25150 &  n_23066;
assign n_29505 = ~n_27773 & ~n_29504;
assign n_29506 =  n_29222 &  n_29505;
assign n_29507 =  n_29503 &  n_29506;
assign n_29508 =  n_24919 &  n_26167;
assign n_29509 = ~n_26124 &  n_26450;
assign n_29510 =  n_29508 &  n_29509;
assign n_29511 = ~n_26843 &  n_8350;
assign n_29512 =  n_24941 &  n_28090;
assign n_29513 =  n_29511 &  n_29512;
assign n_29514 =  n_29510 &  n_29513;
assign n_29515 =  n_29507 &  n_29514;
assign n_29516 =  n_29433 &  n_26101;
assign n_29517 =  n_28059 &  n_24908;
assign n_29518 =  n_29516 &  n_29517;
assign n_29519 =  n_28061 & ~n_29234;
assign n_29520 = ~n_26201 &  n_26831;
assign n_29521 =  n_29519 &  n_29520;
assign n_29522 =  n_29518 &  n_29521;
assign n_29523 =  n_28824 & ~n_27781;
assign n_29524 =  n_28087 & ~n_28829;
assign n_29525 =  n_29523 &  n_29524;
assign n_29526 =  n_27779 & ~n_23421;
assign n_29527 =  n_29434 &  n_28511;
assign n_29528 =  n_29526 &  n_29527;
assign n_29529 =  n_29525 &  n_29528;
assign n_29530 =  n_29522 &  n_29529;
assign n_29531 =  n_29515 &  n_29530;
assign n_29532 =  n_28362 &  n_24702;
assign n_29533 =  n_29007 & ~n_24754;
assign n_29534 =  n_29532 &  n_29533;
assign n_29535 = ~n_26474 & ~n_28855;
assign n_29536 = ~n_26189 & ~n_24923;
assign n_29537 =  n_29535 &  n_29536;
assign n_29538 =  n_26361 &  n_29537;
assign n_29539 =  n_28531 &  n_27583;
assign n_29540 =  n_29538 &  n_29539;
assign n_29541 =  n_29534 &  n_29540;
assign n_29542 =  n_29531 &  n_29541;
assign n_29543 =  n_27867 &  n_27959;
assign n_29544 = ~n_26258 &  n_28789;
assign n_29545 =  n_29543 &  n_29544;
assign n_29546 =  n_29241 &  n_24213;
assign n_29547 =  n_28223 &  n_26207;
assign n_29548 =  n_29546 &  n_29547;
assign n_29549 =  n_29545 &  n_29548;
assign n_29550 = ~n_24115 &  n_28798;
assign n_29551 =  n_28214 &  n_24127;
assign n_29552 =  n_29550 &  n_29551;
assign n_29553 =  n_28800 &  n_27033;
assign n_29554 =  n_29243 &  n_29055;
assign n_29555 =  n_29553 &  n_29554;
assign n_29556 =  n_29552 &  n_29555;
assign n_29557 =  n_29549 &  n_29556;
assign n_29558 = ~n_25648 & ~n_25166;
assign n_29559 = ~n_28884 & ~n_25382;
assign n_29560 =  n_29558 &  n_29559;
assign n_29561 =  n_9884 &  n_25107;
assign n_29562 = ~n_29561 & ~n_28495;
assign n_29563 = ~n_23688 & ~n_23247;
assign n_29564 =  n_29562 &  n_29563;
assign n_29565 =  n_29560 &  n_29564;
assign n_29566 = ~n_28419 & ~n_23623;
assign n_29567 =  n_29566 &  n_28777;
assign n_29568 = ~n_555 & ~n_6180;
assign n_29569 =  n_8360 & ~n_29568;
assign n_29570 = ~n_29569 & ~n_23616;
assign n_29571 = ~n_25249 & ~n_28112;
assign n_29572 =  n_29570 &  n_29571;
assign n_29573 =  n_29567 &  n_29572;
assign n_29574 =  n_29565 &  n_29573;
assign n_29575 = ~n_27699 &  n_29399;
assign n_29576 =  n_26832 &  n_28512;
assign n_29577 =  n_29575 &  n_29576;
assign n_29578 =  n_28836 & ~n_25882;
assign n_29579 = ~n_25923 & ~n_24689;
assign n_29580 =  n_29578 &  n_29579;
assign n_29581 = ~n_23608 & ~n_27840;
assign n_29582 = ~n_26168 & ~n_25857;
assign n_29583 =  n_29581 &  n_29582;
assign n_29584 = ~n_23682 & ~n_24631;
assign n_29585 = ~n_23545 & ~n_25170;
assign n_29586 =  n_29584 &  n_29585;
assign n_29587 =  n_29583 &  n_29586;
assign n_29588 =  n_29580 &  n_29587;
assign n_29589 =  n_29577 &  n_29588;
assign n_29590 =  n_29574 &  n_29589;
assign n_29591 =  n_27957 &  n_28451;
assign n_29592 =  n_24203 &  n_27961;
assign n_29593 =  n_29591 &  n_29592;
assign n_29594 = ~n_25502 & ~n_28041;
assign n_29595 = ~n_26030 &  n_29594;
assign n_29596 =  n_28452 &  n_29595;
assign n_29597 =  n_28264 &  n_29056;
assign n_29598 =  n_29596 &  n_29597;
assign n_29599 =  n_29593 &  n_29598;
assign n_29600 =  n_29590 &  n_29599;
assign n_29601 =  n_29557 &  n_29600;
assign n_29602 =  n_29542 &  n_29601;
assign n_29603 =  n_27085 &  n_28923;
assign n_29604 =  n_26253 &  n_29603;
assign n_29605 = ~n_25512 & ~n_25218;
assign n_29606 = ~x_43 & ~n_29605;
assign n_29607 = ~n_29606 &  n_27663;
assign n_29608 =  n_26863 &  n_29008;
assign n_29609 =  n_29607 &  n_29608;
assign n_29610 =  n_29367 &  n_29190;
assign n_29611 =  n_29370 &  n_28269;
assign n_29612 =  n_29610 &  n_29611;
assign n_29613 =  n_29609 &  n_29612;
assign n_29614 =  n_29371 &  n_26366;
assign n_29615 =  n_27101 &  n_29614;
assign n_29616 =  n_28250 &  n_29615;
assign n_29617 =  n_29613 &  n_29616;
assign n_29618 =  n_29604 &  n_29617;
assign n_29619 =  n_29602 &  n_29618;
assign n_29620 =  n_29500 &  n_29619;
assign n_29621 = ~n_22939 &  n_29620;
assign n_29622 = ~n_25845 &  n_29621;
assign n_29623 = ~n_26634 &  n_29622;
assign n_29624 =  n_29179 &  n_29623;
assign n_29625 =  x_33 & ~n_29624;
assign n_29626 = ~x_33 &  n_29624;
assign n_29627 = ~n_29625 & ~n_29626;
assign n_29628 = ~x_3027 &  n_13143;
assign n_29629 = ~x_3059 &  n_13145;
assign n_29630 = ~i_27 & ~n_13142;
assign n_29631 = ~n_29629 & ~n_29630;
assign n_29632 = ~n_29628 &  n_29631;
assign n_29633 = ~n_13141 & ~n_29632;
assign n_29634 = ~x_2901 &  n_13141;
assign n_29635 = ~n_29633 & ~n_29634;
assign n_29636 = ~n_13136 & ~n_29635;
assign n_29637 = ~x_2837 &  n_13136;
assign n_29638 = ~n_29636 & ~n_29637;
assign n_29639 =  n_13105 & ~n_29638;
assign n_29640 = ~x_2581 & ~n_13105;
assign n_29641 = ~n_29639 & ~n_29640;
assign n_29642 =  x_2581 &  n_29641;
assign n_29643 = ~x_2581 & ~n_29641;
assign n_29644 = ~n_29642 & ~n_29643;
assign n_29645 = ~x_3026 &  n_13143;
assign n_29646 = ~x_3058 &  n_13145;
assign n_29647 = ~i_26 & ~n_13142;
assign n_29648 = ~n_29646 & ~n_29647;
assign n_29649 = ~n_29645 &  n_29648;
assign n_29650 = ~n_13141 & ~n_29649;
assign n_29651 = ~x_2900 &  n_13141;
assign n_29652 = ~n_29650 & ~n_29651;
assign n_29653 = ~n_13136 & ~n_29652;
assign n_29654 = ~x_2836 &  n_13136;
assign n_29655 = ~n_29653 & ~n_29654;
assign n_29656 =  n_13105 & ~n_29655;
assign n_29657 = ~x_2580 & ~n_13105;
assign n_29658 = ~n_29656 & ~n_29657;
assign n_29659 =  x_2580 &  n_29658;
assign n_29660 = ~x_2580 & ~n_29658;
assign n_29661 = ~n_29659 & ~n_29660;
assign n_29662 = ~x_3025 &  n_13143;
assign n_29663 = ~x_3057 &  n_13145;
assign n_29664 = ~i_25 & ~n_13142;
assign n_29665 = ~n_29663 & ~n_29664;
assign n_29666 = ~n_29662 &  n_29665;
assign n_29667 = ~n_13141 & ~n_29666;
assign n_29668 = ~x_2899 &  n_13141;
assign n_29669 = ~n_29667 & ~n_29668;
assign n_29670 = ~n_13136 & ~n_29669;
assign n_29671 = ~x_2835 &  n_13136;
assign n_29672 = ~n_29670 & ~n_29671;
assign n_29673 =  n_13105 & ~n_29672;
assign n_29674 = ~x_2579 & ~n_13105;
assign n_29675 = ~n_29673 & ~n_29674;
assign n_29676 =  x_2579 &  n_29675;
assign n_29677 = ~x_2579 & ~n_29675;
assign n_29678 = ~n_29676 & ~n_29677;
assign n_29679 = ~x_3024 &  n_13143;
assign n_29680 = ~x_3056 &  n_13145;
assign n_29681 = ~i_24 & ~n_13142;
assign n_29682 = ~n_29680 & ~n_29681;
assign n_29683 = ~n_29679 &  n_29682;
assign n_29684 = ~n_13141 & ~n_29683;
assign n_29685 = ~x_2898 &  n_13141;
assign n_29686 = ~n_29684 & ~n_29685;
assign n_29687 = ~n_13136 & ~n_29686;
assign n_29688 = ~x_2834 &  n_13136;
assign n_29689 = ~n_29687 & ~n_29688;
assign n_29690 =  n_13105 & ~n_29689;
assign n_29691 = ~x_2578 & ~n_13105;
assign n_29692 = ~n_29690 & ~n_29691;
assign n_29693 =  x_2578 &  n_29692;
assign n_29694 = ~x_2578 & ~n_29692;
assign n_29695 = ~n_29693 & ~n_29694;
assign n_29696 = ~x_3023 &  n_13143;
assign n_29697 = ~x_3055 &  n_13145;
assign n_29698 = ~i_23 & ~n_13142;
assign n_29699 = ~n_29697 & ~n_29698;
assign n_29700 = ~n_29696 &  n_29699;
assign n_29701 = ~n_13141 & ~n_29700;
assign n_29702 = ~x_2897 &  n_13141;
assign n_29703 = ~n_29701 & ~n_29702;
assign n_29704 = ~n_13136 & ~n_29703;
assign n_29705 = ~x_2833 &  n_13136;
assign n_29706 = ~n_29704 & ~n_29705;
assign n_29707 =  n_13105 & ~n_29706;
assign n_29708 = ~x_2577 & ~n_13105;
assign n_29709 = ~n_29707 & ~n_29708;
assign n_29710 =  x_2577 &  n_29709;
assign n_29711 = ~x_2577 & ~n_29709;
assign n_29712 = ~n_29710 & ~n_29711;
assign n_29713 = ~x_3022 &  n_13143;
assign n_29714 = ~x_3054 &  n_13145;
assign n_29715 = ~i_22 & ~n_13142;
assign n_29716 = ~n_29714 & ~n_29715;
assign n_29717 = ~n_29713 &  n_29716;
assign n_29718 = ~n_13141 & ~n_29717;
assign n_29719 = ~x_2896 &  n_13141;
assign n_29720 = ~n_29718 & ~n_29719;
assign n_29721 = ~n_13136 & ~n_29720;
assign n_29722 = ~x_2832 &  n_13136;
assign n_29723 = ~n_29721 & ~n_29722;
assign n_29724 =  n_13105 & ~n_29723;
assign n_29725 = ~x_2576 & ~n_13105;
assign n_29726 = ~n_29724 & ~n_29725;
assign n_29727 =  x_2576 &  n_29726;
assign n_29728 = ~x_2576 & ~n_29726;
assign n_29729 = ~n_29727 & ~n_29728;
assign n_29730 = ~x_3021 &  n_13143;
assign n_29731 = ~x_3053 &  n_13145;
assign n_29732 = ~i_21 & ~n_13142;
assign n_29733 = ~n_29731 & ~n_29732;
assign n_29734 = ~n_29730 &  n_29733;
assign n_29735 = ~n_13141 & ~n_29734;
assign n_29736 = ~x_2895 &  n_13141;
assign n_29737 = ~n_29735 & ~n_29736;
assign n_29738 = ~n_13136 & ~n_29737;
assign n_29739 = ~x_2831 &  n_13136;
assign n_29740 = ~n_29738 & ~n_29739;
assign n_29741 =  n_13105 & ~n_29740;
assign n_29742 = ~x_2575 & ~n_13105;
assign n_29743 = ~n_29741 & ~n_29742;
assign n_29744 =  x_2575 &  n_29743;
assign n_29745 = ~x_2575 & ~n_29743;
assign n_29746 = ~n_29744 & ~n_29745;
assign n_29747 = ~x_3020 &  n_13143;
assign n_29748 = ~x_3052 &  n_13145;
assign n_29749 = ~i_20 & ~n_13142;
assign n_29750 = ~n_29748 & ~n_29749;
assign n_29751 = ~n_29747 &  n_29750;
assign n_29752 = ~n_13141 & ~n_29751;
assign n_29753 = ~x_2894 &  n_13141;
assign n_29754 = ~n_29752 & ~n_29753;
assign n_29755 = ~n_13136 & ~n_29754;
assign n_29756 = ~x_2830 &  n_13136;
assign n_29757 = ~n_29755 & ~n_29756;
assign n_29758 =  n_13105 & ~n_29757;
assign n_29759 = ~x_2574 & ~n_13105;
assign n_29760 = ~n_29758 & ~n_29759;
assign n_29761 =  x_2574 &  n_29760;
assign n_29762 = ~x_2574 & ~n_29760;
assign n_29763 = ~n_29761 & ~n_29762;
assign n_29764 = ~x_3019 &  n_13143;
assign n_29765 = ~x_3051 &  n_13145;
assign n_29766 = ~i_19 & ~n_13142;
assign n_29767 = ~n_29765 & ~n_29766;
assign n_29768 = ~n_29764 &  n_29767;
assign n_29769 = ~n_13141 & ~n_29768;
assign n_29770 = ~x_2893 &  n_13141;
assign n_29771 = ~n_29769 & ~n_29770;
assign n_29772 = ~n_13136 & ~n_29771;
assign n_29773 = ~x_2829 &  n_13136;
assign n_29774 = ~n_29772 & ~n_29773;
assign n_29775 =  n_13105 & ~n_29774;
assign n_29776 = ~x_2573 & ~n_13105;
assign n_29777 = ~n_29775 & ~n_29776;
assign n_29778 =  x_2573 &  n_29777;
assign n_29779 = ~x_2573 & ~n_29777;
assign n_29780 = ~n_29778 & ~n_29779;
assign n_29781 = ~x_3018 &  n_13143;
assign n_29782 = ~x_3050 &  n_13145;
assign n_29783 = ~i_18 & ~n_13142;
assign n_29784 = ~n_29782 & ~n_29783;
assign n_29785 = ~n_29781 &  n_29784;
assign n_29786 = ~n_13141 & ~n_29785;
assign n_29787 = ~x_2892 &  n_13141;
assign n_29788 = ~n_29786 & ~n_29787;
assign n_29789 = ~n_13136 & ~n_29788;
assign n_29790 = ~x_2828 &  n_13136;
assign n_29791 = ~n_29789 & ~n_29790;
assign n_29792 =  n_13105 & ~n_29791;
assign n_29793 = ~x_2572 & ~n_13105;
assign n_29794 = ~n_29792 & ~n_29793;
assign n_29795 =  x_2572 &  n_29794;
assign n_29796 = ~x_2572 & ~n_29794;
assign n_29797 = ~n_29795 & ~n_29796;
assign n_29798 = ~x_3017 &  n_13143;
assign n_29799 = ~x_3049 &  n_13145;
assign n_29800 = ~i_17 & ~n_13142;
assign n_29801 = ~n_29799 & ~n_29800;
assign n_29802 = ~n_29798 &  n_29801;
assign n_29803 = ~n_13141 & ~n_29802;
assign n_29804 = ~x_2891 &  n_13141;
assign n_29805 = ~n_29803 & ~n_29804;
assign n_29806 = ~n_13136 & ~n_29805;
assign n_29807 = ~x_2827 &  n_13136;
assign n_29808 = ~n_29806 & ~n_29807;
assign n_29809 =  n_13105 & ~n_29808;
assign n_29810 = ~x_2571 & ~n_13105;
assign n_29811 = ~n_29809 & ~n_29810;
assign n_29812 =  x_2571 &  n_29811;
assign n_29813 = ~x_2571 & ~n_29811;
assign n_29814 = ~n_29812 & ~n_29813;
assign n_29815 = ~x_3016 &  n_13143;
assign n_29816 = ~x_3048 &  n_13145;
assign n_29817 = ~i_16 & ~n_13142;
assign n_29818 = ~n_29816 & ~n_29817;
assign n_29819 = ~n_29815 &  n_29818;
assign n_29820 = ~n_13141 & ~n_29819;
assign n_29821 = ~x_2890 &  n_13141;
assign n_29822 = ~n_29820 & ~n_29821;
assign n_29823 = ~n_13136 & ~n_29822;
assign n_29824 = ~x_2826 &  n_13136;
assign n_29825 = ~n_29823 & ~n_29824;
assign n_29826 =  n_13105 & ~n_29825;
assign n_29827 = ~x_2570 & ~n_13105;
assign n_29828 = ~n_29826 & ~n_29827;
assign n_29829 =  x_2570 &  n_29828;
assign n_29830 = ~x_2570 & ~n_29828;
assign n_29831 = ~n_29829 & ~n_29830;
assign n_29832 = ~x_3015 &  n_13143;
assign n_29833 = ~x_3047 &  n_13145;
assign n_29834 = ~i_15 & ~n_13142;
assign n_29835 = ~n_29833 & ~n_29834;
assign n_29836 = ~n_29832 &  n_29835;
assign n_29837 = ~n_13141 & ~n_29836;
assign n_29838 = ~x_2889 &  n_13141;
assign n_29839 = ~n_29837 & ~n_29838;
assign n_29840 = ~n_13136 & ~n_29839;
assign n_29841 = ~x_2825 &  n_13136;
assign n_29842 = ~n_29840 & ~n_29841;
assign n_29843 =  n_13105 & ~n_29842;
assign n_29844 = ~x_2569 & ~n_13105;
assign n_29845 = ~n_29843 & ~n_29844;
assign n_29846 =  x_2569 &  n_29845;
assign n_29847 = ~x_2569 & ~n_29845;
assign n_29848 = ~n_29846 & ~n_29847;
assign n_29849 = ~x_3014 &  n_13143;
assign n_29850 = ~x_3046 &  n_13145;
assign n_29851 = ~i_14 & ~n_13142;
assign n_29852 = ~n_29850 & ~n_29851;
assign n_29853 = ~n_29849 &  n_29852;
assign n_29854 = ~n_13141 & ~n_29853;
assign n_29855 = ~x_2888 &  n_13141;
assign n_29856 = ~n_29854 & ~n_29855;
assign n_29857 = ~n_13136 & ~n_29856;
assign n_29858 = ~x_2824 &  n_13136;
assign n_29859 = ~n_29857 & ~n_29858;
assign n_29860 =  n_13105 & ~n_29859;
assign n_29861 = ~x_2568 & ~n_13105;
assign n_29862 = ~n_29860 & ~n_29861;
assign n_29863 =  x_2568 &  n_29862;
assign n_29864 = ~x_2568 & ~n_29862;
assign n_29865 = ~n_29863 & ~n_29864;
assign n_29866 = ~x_3013 &  n_13143;
assign n_29867 = ~x_3045 &  n_13145;
assign n_29868 = ~i_13 & ~n_13142;
assign n_29869 = ~n_29867 & ~n_29868;
assign n_29870 = ~n_29866 &  n_29869;
assign n_29871 = ~n_13141 & ~n_29870;
assign n_29872 = ~x_2887 &  n_13141;
assign n_29873 = ~n_29871 & ~n_29872;
assign n_29874 = ~n_13136 & ~n_29873;
assign n_29875 = ~x_2823 &  n_13136;
assign n_29876 = ~n_29874 & ~n_29875;
assign n_29877 =  n_13105 & ~n_29876;
assign n_29878 = ~x_2567 & ~n_13105;
assign n_29879 = ~n_29877 & ~n_29878;
assign n_29880 =  x_2567 &  n_29879;
assign n_29881 = ~x_2567 & ~n_29879;
assign n_29882 = ~n_29880 & ~n_29881;
assign n_29883 = ~x_3012 &  n_13143;
assign n_29884 = ~x_3044 &  n_13145;
assign n_29885 = ~i_12 & ~n_13142;
assign n_29886 = ~n_29884 & ~n_29885;
assign n_29887 = ~n_29883 &  n_29886;
assign n_29888 = ~n_13141 & ~n_29887;
assign n_29889 = ~x_2886 &  n_13141;
assign n_29890 = ~n_29888 & ~n_29889;
assign n_29891 = ~n_13136 & ~n_29890;
assign n_29892 = ~x_2822 &  n_13136;
assign n_29893 = ~n_29891 & ~n_29892;
assign n_29894 =  n_13105 & ~n_29893;
assign n_29895 = ~x_2566 & ~n_13105;
assign n_29896 = ~n_29894 & ~n_29895;
assign n_29897 =  x_2566 &  n_29896;
assign n_29898 = ~x_2566 & ~n_29896;
assign n_29899 = ~n_29897 & ~n_29898;
assign n_29900 = ~x_3011 &  n_13143;
assign n_29901 = ~x_3043 &  n_13145;
assign n_29902 = ~i_11 & ~n_13142;
assign n_29903 = ~n_29901 & ~n_29902;
assign n_29904 = ~n_29900 &  n_29903;
assign n_29905 = ~n_13141 & ~n_29904;
assign n_29906 = ~x_2885 &  n_13141;
assign n_29907 = ~n_29905 & ~n_29906;
assign n_29908 = ~n_13136 & ~n_29907;
assign n_29909 = ~x_2821 &  n_13136;
assign n_29910 = ~n_29908 & ~n_29909;
assign n_29911 =  n_13105 & ~n_29910;
assign n_29912 = ~x_2565 & ~n_13105;
assign n_29913 = ~n_29911 & ~n_29912;
assign n_29914 =  x_2565 &  n_29913;
assign n_29915 = ~x_2565 & ~n_29913;
assign n_29916 = ~n_29914 & ~n_29915;
assign n_29917 = ~x_3010 &  n_13143;
assign n_29918 = ~x_3042 &  n_13145;
assign n_29919 = ~i_10 & ~n_13142;
assign n_29920 = ~n_29918 & ~n_29919;
assign n_29921 = ~n_29917 &  n_29920;
assign n_29922 = ~n_13141 & ~n_29921;
assign n_29923 = ~x_2884 &  n_13141;
assign n_29924 = ~n_29922 & ~n_29923;
assign n_29925 = ~n_13136 & ~n_29924;
assign n_29926 = ~x_2820 &  n_13136;
assign n_29927 = ~n_29925 & ~n_29926;
assign n_29928 =  n_13105 & ~n_29927;
assign n_29929 = ~x_2564 & ~n_13105;
assign n_29930 = ~n_29928 & ~n_29929;
assign n_29931 =  x_2564 &  n_29930;
assign n_29932 = ~x_2564 & ~n_29930;
assign n_29933 = ~n_29931 & ~n_29932;
assign n_29934 = ~x_3009 &  n_13143;
assign n_29935 = ~x_3041 &  n_13145;
assign n_29936 = ~i_9 & ~n_13142;
assign n_29937 = ~n_29935 & ~n_29936;
assign n_29938 = ~n_29934 &  n_29937;
assign n_29939 = ~n_13141 & ~n_29938;
assign n_29940 = ~x_2883 &  n_13141;
assign n_29941 = ~n_29939 & ~n_29940;
assign n_29942 = ~n_13136 & ~n_29941;
assign n_29943 = ~x_2819 &  n_13136;
assign n_29944 = ~n_29942 & ~n_29943;
assign n_29945 =  n_13105 & ~n_29944;
assign n_29946 = ~x_2563 & ~n_13105;
assign n_29947 = ~n_29945 & ~n_29946;
assign n_29948 =  x_2563 &  n_29947;
assign n_29949 = ~x_2563 & ~n_29947;
assign n_29950 = ~n_29948 & ~n_29949;
assign n_29951 = ~x_3008 &  n_13143;
assign n_29952 = ~x_3040 &  n_13145;
assign n_29953 = ~i_8 & ~n_13142;
assign n_29954 = ~n_29952 & ~n_29953;
assign n_29955 = ~n_29951 &  n_29954;
assign n_29956 = ~n_13141 & ~n_29955;
assign n_29957 = ~x_2882 &  n_13141;
assign n_29958 = ~n_29956 & ~n_29957;
assign n_29959 = ~n_13136 & ~n_29958;
assign n_29960 = ~x_2818 &  n_13136;
assign n_29961 = ~n_29959 & ~n_29960;
assign n_29962 =  n_13105 & ~n_29961;
assign n_29963 = ~x_2562 & ~n_13105;
assign n_29964 = ~n_29962 & ~n_29963;
assign n_29965 =  x_2562 &  n_29964;
assign n_29966 = ~x_2562 & ~n_29964;
assign n_29967 = ~n_29965 & ~n_29966;
assign n_29968 = ~x_3007 &  n_13143;
assign n_29969 = ~x_3039 &  n_13145;
assign n_29970 = ~i_7 & ~n_13142;
assign n_29971 = ~n_29969 & ~n_29970;
assign n_29972 = ~n_29968 &  n_29971;
assign n_29973 = ~n_13141 & ~n_29972;
assign n_29974 = ~x_2881 &  n_13141;
assign n_29975 = ~n_29973 & ~n_29974;
assign n_29976 = ~n_13136 & ~n_29975;
assign n_29977 = ~x_2817 &  n_13136;
assign n_29978 = ~n_29976 & ~n_29977;
assign n_29979 =  n_13105 & ~n_29978;
assign n_29980 = ~x_2561 & ~n_13105;
assign n_29981 = ~n_29979 & ~n_29980;
assign n_29982 =  x_2561 &  n_29981;
assign n_29983 = ~x_2561 & ~n_29981;
assign n_29984 = ~n_29982 & ~n_29983;
assign n_29985 = ~x_3006 &  n_13143;
assign n_29986 = ~x_3038 &  n_13145;
assign n_29987 = ~i_6 & ~n_13142;
assign n_29988 = ~n_29986 & ~n_29987;
assign n_29989 = ~n_29985 &  n_29988;
assign n_29990 = ~n_13141 & ~n_29989;
assign n_29991 = ~x_2880 &  n_13141;
assign n_29992 = ~n_29990 & ~n_29991;
assign n_29993 = ~n_13136 & ~n_29992;
assign n_29994 = ~x_2816 &  n_13136;
assign n_29995 = ~n_29993 & ~n_29994;
assign n_29996 =  n_13105 & ~n_29995;
assign n_29997 = ~x_2560 & ~n_13105;
assign n_29998 = ~n_29996 & ~n_29997;
assign n_29999 =  x_2560 &  n_29998;
assign n_30000 = ~x_2560 & ~n_29998;
assign n_30001 = ~n_29999 & ~n_30000;
assign n_30002 = ~x_3005 &  n_13143;
assign n_30003 = ~x_3037 &  n_13145;
assign n_30004 = ~i_5 & ~n_13142;
assign n_30005 = ~n_30003 & ~n_30004;
assign n_30006 = ~n_30002 &  n_30005;
assign n_30007 = ~n_13141 & ~n_30006;
assign n_30008 = ~x_2879 &  n_13141;
assign n_30009 = ~n_30007 & ~n_30008;
assign n_30010 = ~n_13136 & ~n_30009;
assign n_30011 = ~x_2815 &  n_13136;
assign n_30012 = ~n_30010 & ~n_30011;
assign n_30013 =  n_13105 & ~n_30012;
assign n_30014 = ~x_2559 & ~n_13105;
assign n_30015 = ~n_30013 & ~n_30014;
assign n_30016 =  x_2559 &  n_30015;
assign n_30017 = ~x_2559 & ~n_30015;
assign n_30018 = ~n_30016 & ~n_30017;
assign n_30019 = ~x_3004 &  n_13143;
assign n_30020 = ~x_3036 &  n_13145;
assign n_30021 = ~i_4 & ~n_13142;
assign n_30022 = ~n_30020 & ~n_30021;
assign n_30023 = ~n_30019 &  n_30022;
assign n_30024 = ~n_13141 & ~n_30023;
assign n_30025 = ~x_2878 &  n_13141;
assign n_30026 = ~n_30024 & ~n_30025;
assign n_30027 = ~n_13136 & ~n_30026;
assign n_30028 = ~x_2814 &  n_13136;
assign n_30029 = ~n_30027 & ~n_30028;
assign n_30030 =  n_13105 & ~n_30029;
assign n_30031 = ~x_2558 & ~n_13105;
assign n_30032 = ~n_30030 & ~n_30031;
assign n_30033 =  x_2558 &  n_30032;
assign n_30034 = ~x_2558 & ~n_30032;
assign n_30035 = ~n_30033 & ~n_30034;
assign n_30036 = ~x_3003 &  n_13143;
assign n_30037 = ~x_3035 &  n_13145;
assign n_30038 = ~i_3 & ~n_13142;
assign n_30039 = ~n_30037 & ~n_30038;
assign n_30040 = ~n_30036 &  n_30039;
assign n_30041 = ~n_13141 & ~n_30040;
assign n_30042 = ~x_2877 &  n_13141;
assign n_30043 = ~n_30041 & ~n_30042;
assign n_30044 = ~n_13136 & ~n_30043;
assign n_30045 = ~x_2813 &  n_13136;
assign n_30046 = ~n_30044 & ~n_30045;
assign n_30047 =  n_13105 & ~n_30046;
assign n_30048 = ~x_2557 & ~n_13105;
assign n_30049 = ~n_30047 & ~n_30048;
assign n_30050 =  x_2557 &  n_30049;
assign n_30051 = ~x_2557 & ~n_30049;
assign n_30052 = ~n_30050 & ~n_30051;
assign n_30053 = ~x_3002 &  n_13143;
assign n_30054 = ~x_3034 &  n_13145;
assign n_30055 = ~i_2 & ~n_13142;
assign n_30056 = ~n_30054 & ~n_30055;
assign n_30057 = ~n_30053 &  n_30056;
assign n_30058 = ~n_13141 & ~n_30057;
assign n_30059 = ~x_2876 &  n_13141;
assign n_30060 = ~n_30058 & ~n_30059;
assign n_30061 = ~n_13136 & ~n_30060;
assign n_30062 = ~x_2812 &  n_13136;
assign n_30063 = ~n_30061 & ~n_30062;
assign n_30064 =  n_13105 & ~n_30063;
assign n_30065 = ~x_2556 & ~n_13105;
assign n_30066 = ~n_30064 & ~n_30065;
assign n_30067 =  x_2556 &  n_30066;
assign n_30068 = ~x_2556 & ~n_30066;
assign n_30069 = ~n_30067 & ~n_30068;
assign n_30070 = ~i_1 & ~n_13145;
assign n_30071 = ~x_3033 &  n_13145;
assign n_30072 = ~n_30070 & ~n_30071;
assign n_30073 = ~n_13143 & ~n_30072;
assign n_30074 = ~x_3001 &  n_13143;
assign n_30075 = ~n_30073 & ~n_30074;
assign n_30076 = ~n_13141 & ~n_30075;
assign n_30077 = ~x_2875 &  n_13141;
assign n_30078 = ~n_30076 & ~n_30077;
assign n_30079 = ~n_13136 & ~n_30078;
assign n_30080 = ~x_2811 &  n_13136;
assign n_30081 = ~n_30079 & ~n_30080;
assign n_30082 =  n_13105 & ~n_30081;
assign n_30083 = ~x_2555 & ~n_13105;
assign n_30084 = ~n_30082 & ~n_30083;
assign n_30085 =  x_2555 &  n_30084;
assign n_30086 = ~x_2555 & ~n_30084;
assign n_30087 = ~n_30085 & ~n_30086;
assign n_30088 =  x_2554 & ~n_23140;
assign n_30089 =  i_32 &  n_23140;
assign n_30090 = ~n_30088 & ~n_30089;
assign n_30091 =  x_2554 & ~n_30090;
assign n_30092 = ~x_2554 &  n_30090;
assign n_30093 = ~n_30091 & ~n_30092;
assign n_30094 =  x_2553 & ~n_23140;
assign n_30095 =  i_31 &  n_23140;
assign n_30096 = ~n_30094 & ~n_30095;
assign n_30097 =  x_2553 & ~n_30096;
assign n_30098 = ~x_2553 &  n_30096;
assign n_30099 = ~n_30097 & ~n_30098;
assign n_30100 =  x_2552 & ~n_23140;
assign n_30101 =  i_30 &  n_23140;
assign n_30102 = ~n_30100 & ~n_30101;
assign n_30103 =  x_2552 & ~n_30102;
assign n_30104 = ~x_2552 &  n_30102;
assign n_30105 = ~n_30103 & ~n_30104;
assign n_30106 =  x_2551 & ~n_23140;
assign n_30107 =  i_29 &  n_23140;
assign n_30108 = ~n_30106 & ~n_30107;
assign n_30109 =  x_2551 & ~n_30108;
assign n_30110 = ~x_2551 &  n_30108;
assign n_30111 = ~n_30109 & ~n_30110;
assign n_30112 =  x_2550 & ~n_23140;
assign n_30113 =  i_28 &  n_23140;
assign n_30114 = ~n_30112 & ~n_30113;
assign n_30115 =  x_2550 & ~n_30114;
assign n_30116 = ~x_2550 &  n_30114;
assign n_30117 = ~n_30115 & ~n_30116;
assign n_30118 =  x_2549 & ~n_23140;
assign n_30119 =  i_27 &  n_23140;
assign n_30120 = ~n_30118 & ~n_30119;
assign n_30121 =  x_2549 & ~n_30120;
assign n_30122 = ~x_2549 &  n_30120;
assign n_30123 = ~n_30121 & ~n_30122;
assign n_30124 =  x_2548 & ~n_23140;
assign n_30125 =  i_26 &  n_23140;
assign n_30126 = ~n_30124 & ~n_30125;
assign n_30127 =  x_2548 & ~n_30126;
assign n_30128 = ~x_2548 &  n_30126;
assign n_30129 = ~n_30127 & ~n_30128;
assign n_30130 =  x_2547 & ~n_23140;
assign n_30131 =  i_25 &  n_23140;
assign n_30132 = ~n_30130 & ~n_30131;
assign n_30133 =  x_2547 & ~n_30132;
assign n_30134 = ~x_2547 &  n_30132;
assign n_30135 = ~n_30133 & ~n_30134;
assign n_30136 =  x_2546 & ~n_23140;
assign n_30137 =  i_24 &  n_23140;
assign n_30138 = ~n_30136 & ~n_30137;
assign n_30139 =  x_2546 & ~n_30138;
assign n_30140 = ~x_2546 &  n_30138;
assign n_30141 = ~n_30139 & ~n_30140;
assign n_30142 =  x_2545 & ~n_23140;
assign n_30143 =  i_23 &  n_23140;
assign n_30144 = ~n_30142 & ~n_30143;
assign n_30145 =  x_2545 & ~n_30144;
assign n_30146 = ~x_2545 &  n_30144;
assign n_30147 = ~n_30145 & ~n_30146;
assign n_30148 =  x_2544 & ~n_23140;
assign n_30149 =  i_22 &  n_23140;
assign n_30150 = ~n_30148 & ~n_30149;
assign n_30151 =  x_2544 & ~n_30150;
assign n_30152 = ~x_2544 &  n_30150;
assign n_30153 = ~n_30151 & ~n_30152;
assign n_30154 =  x_2543 & ~n_23140;
assign n_30155 =  i_21 &  n_23140;
assign n_30156 = ~n_30154 & ~n_30155;
assign n_30157 =  x_2543 & ~n_30156;
assign n_30158 = ~x_2543 &  n_30156;
assign n_30159 = ~n_30157 & ~n_30158;
assign n_30160 =  x_2542 & ~n_23140;
assign n_30161 =  i_20 &  n_23140;
assign n_30162 = ~n_30160 & ~n_30161;
assign n_30163 =  x_2542 & ~n_30162;
assign n_30164 = ~x_2542 &  n_30162;
assign n_30165 = ~n_30163 & ~n_30164;
assign n_30166 =  x_2541 & ~n_23140;
assign n_30167 =  i_19 &  n_23140;
assign n_30168 = ~n_30166 & ~n_30167;
assign n_30169 =  x_2541 & ~n_30168;
assign n_30170 = ~x_2541 &  n_30168;
assign n_30171 = ~n_30169 & ~n_30170;
assign n_30172 =  x_2540 & ~n_23140;
assign n_30173 =  i_18 &  n_23140;
assign n_30174 = ~n_30172 & ~n_30173;
assign n_30175 =  x_2540 & ~n_30174;
assign n_30176 = ~x_2540 &  n_30174;
assign n_30177 = ~n_30175 & ~n_30176;
assign n_30178 =  x_2539 & ~n_23140;
assign n_30179 =  i_17 &  n_23140;
assign n_30180 = ~n_30178 & ~n_30179;
assign n_30181 =  x_2539 & ~n_30180;
assign n_30182 = ~x_2539 &  n_30180;
assign n_30183 = ~n_30181 & ~n_30182;
assign n_30184 =  x_2538 & ~n_23140;
assign n_30185 =  i_16 &  n_23140;
assign n_30186 = ~n_30184 & ~n_30185;
assign n_30187 =  x_2538 & ~n_30186;
assign n_30188 = ~x_2538 &  n_30186;
assign n_30189 = ~n_30187 & ~n_30188;
assign n_30190 =  x_2537 & ~n_23140;
assign n_30191 =  i_15 &  n_23140;
assign n_30192 = ~n_30190 & ~n_30191;
assign n_30193 =  x_2537 & ~n_30192;
assign n_30194 = ~x_2537 &  n_30192;
assign n_30195 = ~n_30193 & ~n_30194;
assign n_30196 =  x_2536 & ~n_23140;
assign n_30197 =  i_14 &  n_23140;
assign n_30198 = ~n_30196 & ~n_30197;
assign n_30199 =  x_2536 & ~n_30198;
assign n_30200 = ~x_2536 &  n_30198;
assign n_30201 = ~n_30199 & ~n_30200;
assign n_30202 =  x_2535 & ~n_23140;
assign n_30203 =  i_13 &  n_23140;
assign n_30204 = ~n_30202 & ~n_30203;
assign n_30205 =  x_2535 & ~n_30204;
assign n_30206 = ~x_2535 &  n_30204;
assign n_30207 = ~n_30205 & ~n_30206;
assign n_30208 =  x_2534 & ~n_23140;
assign n_30209 =  i_12 &  n_23140;
assign n_30210 = ~n_30208 & ~n_30209;
assign n_30211 =  x_2534 & ~n_30210;
assign n_30212 = ~x_2534 &  n_30210;
assign n_30213 = ~n_30211 & ~n_30212;
assign n_30214 =  x_2533 & ~n_23140;
assign n_30215 =  i_11 &  n_23140;
assign n_30216 = ~n_30214 & ~n_30215;
assign n_30217 =  x_2533 & ~n_30216;
assign n_30218 = ~x_2533 &  n_30216;
assign n_30219 = ~n_30217 & ~n_30218;
assign n_30220 =  x_2532 & ~n_23140;
assign n_30221 =  i_10 &  n_23140;
assign n_30222 = ~n_30220 & ~n_30221;
assign n_30223 =  x_2532 & ~n_30222;
assign n_30224 = ~x_2532 &  n_30222;
assign n_30225 = ~n_30223 & ~n_30224;
assign n_30226 =  x_2531 & ~n_23140;
assign n_30227 =  i_9 &  n_23140;
assign n_30228 = ~n_30226 & ~n_30227;
assign n_30229 =  x_2531 & ~n_30228;
assign n_30230 = ~x_2531 &  n_30228;
assign n_30231 = ~n_30229 & ~n_30230;
assign n_30232 =  x_2530 & ~n_23140;
assign n_30233 =  i_8 &  n_23140;
assign n_30234 = ~n_30232 & ~n_30233;
assign n_30235 =  x_2530 & ~n_30234;
assign n_30236 = ~x_2530 &  n_30234;
assign n_30237 = ~n_30235 & ~n_30236;
assign n_30238 =  x_2529 & ~n_23140;
assign n_30239 =  i_7 &  n_23140;
assign n_30240 = ~n_30238 & ~n_30239;
assign n_30241 =  x_2529 & ~n_30240;
assign n_30242 = ~x_2529 &  n_30240;
assign n_30243 = ~n_30241 & ~n_30242;
assign n_30244 =  x_2528 & ~n_23140;
assign n_30245 =  i_6 &  n_23140;
assign n_30246 = ~n_30244 & ~n_30245;
assign n_30247 =  x_2528 & ~n_30246;
assign n_30248 = ~x_2528 &  n_30246;
assign n_30249 = ~n_30247 & ~n_30248;
assign n_30250 =  x_2527 & ~n_23140;
assign n_30251 =  i_5 &  n_23140;
assign n_30252 = ~n_30250 & ~n_30251;
assign n_30253 =  x_2527 & ~n_30252;
assign n_30254 = ~x_2527 &  n_30252;
assign n_30255 = ~n_30253 & ~n_30254;
assign n_30256 =  x_2526 & ~n_23140;
assign n_30257 =  i_4 &  n_23140;
assign n_30258 = ~n_30256 & ~n_30257;
assign n_30259 =  x_2526 & ~n_30258;
assign n_30260 = ~x_2526 &  n_30258;
assign n_30261 = ~n_30259 & ~n_30260;
assign n_30262 =  x_2525 & ~n_23140;
assign n_30263 =  i_3 &  n_23140;
assign n_30264 = ~n_30262 & ~n_30263;
assign n_30265 =  x_2525 & ~n_30264;
assign n_30266 = ~x_2525 &  n_30264;
assign n_30267 = ~n_30265 & ~n_30266;
assign n_30268 =  x_2524 & ~n_23140;
assign n_30269 =  i_2 &  n_23140;
assign n_30270 = ~n_30268 & ~n_30269;
assign n_30271 =  x_2524 & ~n_30270;
assign n_30272 = ~x_2524 &  n_30270;
assign n_30273 = ~n_30271 & ~n_30272;
assign n_30274 =  x_2523 & ~n_23140;
assign n_30275 =  i_1 &  n_23140;
assign n_30276 = ~n_30274 & ~n_30275;
assign n_30277 =  x_2523 & ~n_30276;
assign n_30278 = ~x_2523 &  n_30276;
assign n_30279 = ~n_30277 & ~n_30278;
assign n_30280 =  x_2522 & ~n_25669;
assign n_30281 =  i_32 &  n_25669;
assign n_30282 = ~n_30280 & ~n_30281;
assign n_30283 =  x_2522 & ~n_30282;
assign n_30284 = ~x_2522 &  n_30282;
assign n_30285 = ~n_30283 & ~n_30284;
assign n_30286 =  x_2521 & ~n_25669;
assign n_30287 =  i_31 &  n_25669;
assign n_30288 = ~n_30286 & ~n_30287;
assign n_30289 =  x_2521 & ~n_30288;
assign n_30290 = ~x_2521 &  n_30288;
assign n_30291 = ~n_30289 & ~n_30290;
assign n_30292 =  x_2520 & ~n_25669;
assign n_30293 =  i_30 &  n_25669;
assign n_30294 = ~n_30292 & ~n_30293;
assign n_30295 =  x_2520 & ~n_30294;
assign n_30296 = ~x_2520 &  n_30294;
assign n_30297 = ~n_30295 & ~n_30296;
assign n_30298 =  x_2519 & ~n_25669;
assign n_30299 =  i_29 &  n_25669;
assign n_30300 = ~n_30298 & ~n_30299;
assign n_30301 =  x_2519 & ~n_30300;
assign n_30302 = ~x_2519 &  n_30300;
assign n_30303 = ~n_30301 & ~n_30302;
assign n_30304 =  x_2518 & ~n_25669;
assign n_30305 =  i_28 &  n_25669;
assign n_30306 = ~n_30304 & ~n_30305;
assign n_30307 =  x_2518 & ~n_30306;
assign n_30308 = ~x_2518 &  n_30306;
assign n_30309 = ~n_30307 & ~n_30308;
assign n_30310 =  x_2517 & ~n_25669;
assign n_30311 =  i_27 &  n_25669;
assign n_30312 = ~n_30310 & ~n_30311;
assign n_30313 =  x_2517 & ~n_30312;
assign n_30314 = ~x_2517 &  n_30312;
assign n_30315 = ~n_30313 & ~n_30314;
assign n_30316 =  x_2516 & ~n_25669;
assign n_30317 =  i_26 &  n_25669;
assign n_30318 = ~n_30316 & ~n_30317;
assign n_30319 =  x_2516 & ~n_30318;
assign n_30320 = ~x_2516 &  n_30318;
assign n_30321 = ~n_30319 & ~n_30320;
assign n_30322 =  x_2515 & ~n_25669;
assign n_30323 =  i_25 &  n_25669;
assign n_30324 = ~n_30322 & ~n_30323;
assign n_30325 =  x_2515 & ~n_30324;
assign n_30326 = ~x_2515 &  n_30324;
assign n_30327 = ~n_30325 & ~n_30326;
assign n_30328 =  x_2514 & ~n_25669;
assign n_30329 =  i_24 &  n_25669;
assign n_30330 = ~n_30328 & ~n_30329;
assign n_30331 =  x_2514 & ~n_30330;
assign n_30332 = ~x_2514 &  n_30330;
assign n_30333 = ~n_30331 & ~n_30332;
assign n_30334 =  x_2513 & ~n_25669;
assign n_30335 =  i_23 &  n_25669;
assign n_30336 = ~n_30334 & ~n_30335;
assign n_30337 =  x_2513 & ~n_30336;
assign n_30338 = ~x_2513 &  n_30336;
assign n_30339 = ~n_30337 & ~n_30338;
assign n_30340 =  x_2512 & ~n_25669;
assign n_30341 =  i_22 &  n_25669;
assign n_30342 = ~n_30340 & ~n_30341;
assign n_30343 =  x_2512 & ~n_30342;
assign n_30344 = ~x_2512 &  n_30342;
assign n_30345 = ~n_30343 & ~n_30344;
assign n_30346 =  x_2511 & ~n_25669;
assign n_30347 =  i_21 &  n_25669;
assign n_30348 = ~n_30346 & ~n_30347;
assign n_30349 =  x_2511 & ~n_30348;
assign n_30350 = ~x_2511 &  n_30348;
assign n_30351 = ~n_30349 & ~n_30350;
assign n_30352 =  x_2510 & ~n_25669;
assign n_30353 =  i_20 &  n_25669;
assign n_30354 = ~n_30352 & ~n_30353;
assign n_30355 =  x_2510 & ~n_30354;
assign n_30356 = ~x_2510 &  n_30354;
assign n_30357 = ~n_30355 & ~n_30356;
assign n_30358 =  x_2509 & ~n_25669;
assign n_30359 =  i_19 &  n_25669;
assign n_30360 = ~n_30358 & ~n_30359;
assign n_30361 =  x_2509 & ~n_30360;
assign n_30362 = ~x_2509 &  n_30360;
assign n_30363 = ~n_30361 & ~n_30362;
assign n_30364 =  x_2508 & ~n_25669;
assign n_30365 =  i_18 &  n_25669;
assign n_30366 = ~n_30364 & ~n_30365;
assign n_30367 =  x_2508 & ~n_30366;
assign n_30368 = ~x_2508 &  n_30366;
assign n_30369 = ~n_30367 & ~n_30368;
assign n_30370 =  x_2507 & ~n_25669;
assign n_30371 =  i_17 &  n_25669;
assign n_30372 = ~n_30370 & ~n_30371;
assign n_30373 =  x_2507 & ~n_30372;
assign n_30374 = ~x_2507 &  n_30372;
assign n_30375 = ~n_30373 & ~n_30374;
assign n_30376 =  x_2506 & ~n_25669;
assign n_30377 =  i_16 &  n_25669;
assign n_30378 = ~n_30376 & ~n_30377;
assign n_30379 =  x_2506 & ~n_30378;
assign n_30380 = ~x_2506 &  n_30378;
assign n_30381 = ~n_30379 & ~n_30380;
assign n_30382 =  x_2505 & ~n_25669;
assign n_30383 =  i_15 &  n_25669;
assign n_30384 = ~n_30382 & ~n_30383;
assign n_30385 =  x_2505 & ~n_30384;
assign n_30386 = ~x_2505 &  n_30384;
assign n_30387 = ~n_30385 & ~n_30386;
assign n_30388 =  x_2504 & ~n_25669;
assign n_30389 =  i_14 &  n_25669;
assign n_30390 = ~n_30388 & ~n_30389;
assign n_30391 =  x_2504 & ~n_30390;
assign n_30392 = ~x_2504 &  n_30390;
assign n_30393 = ~n_30391 & ~n_30392;
assign n_30394 =  x_2503 & ~n_25669;
assign n_30395 =  i_13 &  n_25669;
assign n_30396 = ~n_30394 & ~n_30395;
assign n_30397 =  x_2503 & ~n_30396;
assign n_30398 = ~x_2503 &  n_30396;
assign n_30399 = ~n_30397 & ~n_30398;
assign n_30400 =  x_2502 & ~n_25669;
assign n_30401 =  i_12 &  n_25669;
assign n_30402 = ~n_30400 & ~n_30401;
assign n_30403 =  x_2502 & ~n_30402;
assign n_30404 = ~x_2502 &  n_30402;
assign n_30405 = ~n_30403 & ~n_30404;
assign n_30406 =  x_2501 & ~n_25669;
assign n_30407 =  i_11 &  n_25669;
assign n_30408 = ~n_30406 & ~n_30407;
assign n_30409 =  x_2501 & ~n_30408;
assign n_30410 = ~x_2501 &  n_30408;
assign n_30411 = ~n_30409 & ~n_30410;
assign n_30412 =  x_2500 & ~n_25669;
assign n_30413 =  i_10 &  n_25669;
assign n_30414 = ~n_30412 & ~n_30413;
assign n_30415 =  x_2500 & ~n_30414;
assign n_30416 = ~x_2500 &  n_30414;
assign n_30417 = ~n_30415 & ~n_30416;
assign n_30418 =  x_2499 & ~n_25669;
assign n_30419 =  i_9 &  n_25669;
assign n_30420 = ~n_30418 & ~n_30419;
assign n_30421 =  x_2499 & ~n_30420;
assign n_30422 = ~x_2499 &  n_30420;
assign n_30423 = ~n_30421 & ~n_30422;
assign n_30424 =  x_2498 & ~n_25669;
assign n_30425 =  i_8 &  n_25669;
assign n_30426 = ~n_30424 & ~n_30425;
assign n_30427 =  x_2498 & ~n_30426;
assign n_30428 = ~x_2498 &  n_30426;
assign n_30429 = ~n_30427 & ~n_30428;
assign n_30430 =  x_2497 & ~n_25669;
assign n_30431 =  i_7 &  n_25669;
assign n_30432 = ~n_30430 & ~n_30431;
assign n_30433 =  x_2497 & ~n_30432;
assign n_30434 = ~x_2497 &  n_30432;
assign n_30435 = ~n_30433 & ~n_30434;
assign n_30436 =  x_2496 & ~n_25669;
assign n_30437 =  i_6 &  n_25669;
assign n_30438 = ~n_30436 & ~n_30437;
assign n_30439 =  x_2496 & ~n_30438;
assign n_30440 = ~x_2496 &  n_30438;
assign n_30441 = ~n_30439 & ~n_30440;
assign n_30442 =  x_2495 & ~n_25669;
assign n_30443 =  i_5 &  n_25669;
assign n_30444 = ~n_30442 & ~n_30443;
assign n_30445 =  x_2495 & ~n_30444;
assign n_30446 = ~x_2495 &  n_30444;
assign n_30447 = ~n_30445 & ~n_30446;
assign n_30448 =  x_2494 & ~n_25669;
assign n_30449 =  i_4 &  n_25669;
assign n_30450 = ~n_30448 & ~n_30449;
assign n_30451 =  x_2494 & ~n_30450;
assign n_30452 = ~x_2494 &  n_30450;
assign n_30453 = ~n_30451 & ~n_30452;
assign n_30454 =  x_2493 & ~n_25669;
assign n_30455 =  i_3 &  n_25669;
assign n_30456 = ~n_30454 & ~n_30455;
assign n_30457 =  x_2493 & ~n_30456;
assign n_30458 = ~x_2493 &  n_30456;
assign n_30459 = ~n_30457 & ~n_30458;
assign n_30460 =  x_2492 & ~n_25669;
assign n_30461 =  i_2 &  n_25669;
assign n_30462 = ~n_30460 & ~n_30461;
assign n_30463 =  x_2492 & ~n_30462;
assign n_30464 = ~x_2492 &  n_30462;
assign n_30465 = ~n_30463 & ~n_30464;
assign n_30466 =  x_2491 & ~n_25669;
assign n_30467 =  i_1 &  n_25669;
assign n_30468 = ~n_30466 & ~n_30467;
assign n_30469 =  x_2491 & ~n_30468;
assign n_30470 = ~x_2491 &  n_30468;
assign n_30471 = ~n_30469 & ~n_30470;
assign n_30472 =  x_2490 & ~n_24989;
assign n_30473 =  i_32 &  n_24989;
assign n_30474 = ~n_30472 & ~n_30473;
assign n_30475 =  x_2490 & ~n_30474;
assign n_30476 = ~x_2490 &  n_30474;
assign n_30477 = ~n_30475 & ~n_30476;
assign n_30478 =  x_2489 & ~n_24989;
assign n_30479 =  i_31 &  n_24989;
assign n_30480 = ~n_30478 & ~n_30479;
assign n_30481 =  x_2489 & ~n_30480;
assign n_30482 = ~x_2489 &  n_30480;
assign n_30483 = ~n_30481 & ~n_30482;
assign n_30484 =  x_2488 & ~n_24989;
assign n_30485 =  i_30 &  n_24989;
assign n_30486 = ~n_30484 & ~n_30485;
assign n_30487 =  x_2488 & ~n_30486;
assign n_30488 = ~x_2488 &  n_30486;
assign n_30489 = ~n_30487 & ~n_30488;
assign n_30490 =  x_2487 & ~n_24989;
assign n_30491 =  i_29 &  n_24989;
assign n_30492 = ~n_30490 & ~n_30491;
assign n_30493 =  x_2487 & ~n_30492;
assign n_30494 = ~x_2487 &  n_30492;
assign n_30495 = ~n_30493 & ~n_30494;
assign n_30496 =  x_2486 & ~n_24989;
assign n_30497 =  i_28 &  n_24989;
assign n_30498 = ~n_30496 & ~n_30497;
assign n_30499 =  x_2486 & ~n_30498;
assign n_30500 = ~x_2486 &  n_30498;
assign n_30501 = ~n_30499 & ~n_30500;
assign n_30502 =  x_2485 & ~n_24989;
assign n_30503 =  i_27 &  n_24989;
assign n_30504 = ~n_30502 & ~n_30503;
assign n_30505 =  x_2485 & ~n_30504;
assign n_30506 = ~x_2485 &  n_30504;
assign n_30507 = ~n_30505 & ~n_30506;
assign n_30508 =  x_2484 & ~n_24989;
assign n_30509 =  i_26 &  n_24989;
assign n_30510 = ~n_30508 & ~n_30509;
assign n_30511 =  x_2484 & ~n_30510;
assign n_30512 = ~x_2484 &  n_30510;
assign n_30513 = ~n_30511 & ~n_30512;
assign n_30514 =  x_2483 & ~n_24989;
assign n_30515 =  i_25 &  n_24989;
assign n_30516 = ~n_30514 & ~n_30515;
assign n_30517 =  x_2483 & ~n_30516;
assign n_30518 = ~x_2483 &  n_30516;
assign n_30519 = ~n_30517 & ~n_30518;
assign n_30520 =  x_2482 & ~n_24989;
assign n_30521 =  i_24 &  n_24989;
assign n_30522 = ~n_30520 & ~n_30521;
assign n_30523 =  x_2482 & ~n_30522;
assign n_30524 = ~x_2482 &  n_30522;
assign n_30525 = ~n_30523 & ~n_30524;
assign n_30526 =  x_2481 & ~n_24989;
assign n_30527 =  i_23 &  n_24989;
assign n_30528 = ~n_30526 & ~n_30527;
assign n_30529 =  x_2481 & ~n_30528;
assign n_30530 = ~x_2481 &  n_30528;
assign n_30531 = ~n_30529 & ~n_30530;
assign n_30532 =  x_2480 & ~n_24989;
assign n_30533 =  i_22 &  n_24989;
assign n_30534 = ~n_30532 & ~n_30533;
assign n_30535 =  x_2480 & ~n_30534;
assign n_30536 = ~x_2480 &  n_30534;
assign n_30537 = ~n_30535 & ~n_30536;
assign n_30538 =  x_2479 & ~n_24989;
assign n_30539 =  i_21 &  n_24989;
assign n_30540 = ~n_30538 & ~n_30539;
assign n_30541 =  x_2479 & ~n_30540;
assign n_30542 = ~x_2479 &  n_30540;
assign n_30543 = ~n_30541 & ~n_30542;
assign n_30544 =  x_2478 & ~n_24989;
assign n_30545 =  i_20 &  n_24989;
assign n_30546 = ~n_30544 & ~n_30545;
assign n_30547 =  x_2478 & ~n_30546;
assign n_30548 = ~x_2478 &  n_30546;
assign n_30549 = ~n_30547 & ~n_30548;
assign n_30550 =  x_2477 & ~n_24989;
assign n_30551 =  i_19 &  n_24989;
assign n_30552 = ~n_30550 & ~n_30551;
assign n_30553 =  x_2477 & ~n_30552;
assign n_30554 = ~x_2477 &  n_30552;
assign n_30555 = ~n_30553 & ~n_30554;
assign n_30556 =  x_2476 & ~n_24989;
assign n_30557 =  i_18 &  n_24989;
assign n_30558 = ~n_30556 & ~n_30557;
assign n_30559 =  x_2476 & ~n_30558;
assign n_30560 = ~x_2476 &  n_30558;
assign n_30561 = ~n_30559 & ~n_30560;
assign n_30562 =  x_2475 & ~n_24989;
assign n_30563 =  i_17 &  n_24989;
assign n_30564 = ~n_30562 & ~n_30563;
assign n_30565 =  x_2475 & ~n_30564;
assign n_30566 = ~x_2475 &  n_30564;
assign n_30567 = ~n_30565 & ~n_30566;
assign n_30568 =  x_2474 & ~n_24989;
assign n_30569 =  i_16 &  n_24989;
assign n_30570 = ~n_30568 & ~n_30569;
assign n_30571 =  x_2474 & ~n_30570;
assign n_30572 = ~x_2474 &  n_30570;
assign n_30573 = ~n_30571 & ~n_30572;
assign n_30574 =  x_2473 & ~n_24989;
assign n_30575 =  i_15 &  n_24989;
assign n_30576 = ~n_30574 & ~n_30575;
assign n_30577 =  x_2473 & ~n_30576;
assign n_30578 = ~x_2473 &  n_30576;
assign n_30579 = ~n_30577 & ~n_30578;
assign n_30580 =  x_2472 & ~n_24989;
assign n_30581 =  i_14 &  n_24989;
assign n_30582 = ~n_30580 & ~n_30581;
assign n_30583 =  x_2472 & ~n_30582;
assign n_30584 = ~x_2472 &  n_30582;
assign n_30585 = ~n_30583 & ~n_30584;
assign n_30586 =  x_2471 & ~n_24989;
assign n_30587 =  i_13 &  n_24989;
assign n_30588 = ~n_30586 & ~n_30587;
assign n_30589 =  x_2471 & ~n_30588;
assign n_30590 = ~x_2471 &  n_30588;
assign n_30591 = ~n_30589 & ~n_30590;
assign n_30592 =  x_2470 & ~n_24989;
assign n_30593 =  i_12 &  n_24989;
assign n_30594 = ~n_30592 & ~n_30593;
assign n_30595 =  x_2470 & ~n_30594;
assign n_30596 = ~x_2470 &  n_30594;
assign n_30597 = ~n_30595 & ~n_30596;
assign n_30598 =  x_2469 & ~n_24989;
assign n_30599 =  i_11 &  n_24989;
assign n_30600 = ~n_30598 & ~n_30599;
assign n_30601 =  x_2469 & ~n_30600;
assign n_30602 = ~x_2469 &  n_30600;
assign n_30603 = ~n_30601 & ~n_30602;
assign n_30604 =  x_2468 & ~n_24989;
assign n_30605 =  i_10 &  n_24989;
assign n_30606 = ~n_30604 & ~n_30605;
assign n_30607 =  x_2468 & ~n_30606;
assign n_30608 = ~x_2468 &  n_30606;
assign n_30609 = ~n_30607 & ~n_30608;
assign n_30610 =  x_2467 & ~n_24989;
assign n_30611 =  i_9 &  n_24989;
assign n_30612 = ~n_30610 & ~n_30611;
assign n_30613 =  x_2467 & ~n_30612;
assign n_30614 = ~x_2467 &  n_30612;
assign n_30615 = ~n_30613 & ~n_30614;
assign n_30616 =  x_2466 & ~n_24989;
assign n_30617 =  i_8 &  n_24989;
assign n_30618 = ~n_30616 & ~n_30617;
assign n_30619 =  x_2466 & ~n_30618;
assign n_30620 = ~x_2466 &  n_30618;
assign n_30621 = ~n_30619 & ~n_30620;
assign n_30622 =  x_2465 & ~n_24989;
assign n_30623 =  i_7 &  n_24989;
assign n_30624 = ~n_30622 & ~n_30623;
assign n_30625 =  x_2465 & ~n_30624;
assign n_30626 = ~x_2465 &  n_30624;
assign n_30627 = ~n_30625 & ~n_30626;
assign n_30628 =  x_2464 & ~n_24989;
assign n_30629 =  i_6 &  n_24989;
assign n_30630 = ~n_30628 & ~n_30629;
assign n_30631 =  x_2464 & ~n_30630;
assign n_30632 = ~x_2464 &  n_30630;
assign n_30633 = ~n_30631 & ~n_30632;
assign n_30634 =  x_2463 & ~n_24989;
assign n_30635 =  i_5 &  n_24989;
assign n_30636 = ~n_30634 & ~n_30635;
assign n_30637 =  x_2463 & ~n_30636;
assign n_30638 = ~x_2463 &  n_30636;
assign n_30639 = ~n_30637 & ~n_30638;
assign n_30640 =  x_2462 & ~n_24989;
assign n_30641 =  i_4 &  n_24989;
assign n_30642 = ~n_30640 & ~n_30641;
assign n_30643 =  x_2462 & ~n_30642;
assign n_30644 = ~x_2462 &  n_30642;
assign n_30645 = ~n_30643 & ~n_30644;
assign n_30646 =  x_2461 & ~n_24989;
assign n_30647 =  i_3 &  n_24989;
assign n_30648 = ~n_30646 & ~n_30647;
assign n_30649 =  x_2461 & ~n_30648;
assign n_30650 = ~x_2461 &  n_30648;
assign n_30651 = ~n_30649 & ~n_30650;
assign n_30652 =  x_2460 & ~n_24989;
assign n_30653 =  i_2 &  n_24989;
assign n_30654 = ~n_30652 & ~n_30653;
assign n_30655 =  x_2460 & ~n_30654;
assign n_30656 = ~x_2460 &  n_30654;
assign n_30657 = ~n_30655 & ~n_30656;
assign n_30658 =  x_2459 & ~n_24989;
assign n_30659 =  i_1 &  n_24989;
assign n_30660 = ~n_30658 & ~n_30659;
assign n_30661 =  x_2459 & ~n_30660;
assign n_30662 = ~x_2459 &  n_30660;
assign n_30663 = ~n_30661 & ~n_30662;
assign n_30664 =  x_2427 & ~n_25672;
assign n_30665 =  i_32 &  n_25672;
assign n_30666 = ~n_30664 & ~n_30665;
assign n_30667 =  x_2427 & ~n_30666;
assign n_30668 = ~x_2427 &  n_30666;
assign n_30669 = ~n_30667 & ~n_30668;
assign n_30670 =  x_2426 & ~n_25672;
assign n_30671 =  i_31 &  n_25672;
assign n_30672 = ~n_30670 & ~n_30671;
assign n_30673 =  x_2426 & ~n_30672;
assign n_30674 = ~x_2426 &  n_30672;
assign n_30675 = ~n_30673 & ~n_30674;
assign n_30676 =  x_2425 & ~n_25672;
assign n_30677 =  i_30 &  n_25672;
assign n_30678 = ~n_30676 & ~n_30677;
assign n_30679 =  x_2425 & ~n_30678;
assign n_30680 = ~x_2425 &  n_30678;
assign n_30681 = ~n_30679 & ~n_30680;
assign n_30682 =  x_2424 & ~n_25672;
assign n_30683 =  i_29 &  n_25672;
assign n_30684 = ~n_30682 & ~n_30683;
assign n_30685 =  x_2424 & ~n_30684;
assign n_30686 = ~x_2424 &  n_30684;
assign n_30687 = ~n_30685 & ~n_30686;
assign n_30688 =  x_2423 & ~n_25672;
assign n_30689 =  i_28 &  n_25672;
assign n_30690 = ~n_30688 & ~n_30689;
assign n_30691 =  x_2423 & ~n_30690;
assign n_30692 = ~x_2423 &  n_30690;
assign n_30693 = ~n_30691 & ~n_30692;
assign n_30694 =  x_2422 & ~n_25672;
assign n_30695 =  i_27 &  n_25672;
assign n_30696 = ~n_30694 & ~n_30695;
assign n_30697 =  x_2422 & ~n_30696;
assign n_30698 = ~x_2422 &  n_30696;
assign n_30699 = ~n_30697 & ~n_30698;
assign n_30700 =  x_2421 & ~n_25672;
assign n_30701 =  i_26 &  n_25672;
assign n_30702 = ~n_30700 & ~n_30701;
assign n_30703 =  x_2421 & ~n_30702;
assign n_30704 = ~x_2421 &  n_30702;
assign n_30705 = ~n_30703 & ~n_30704;
assign n_30706 =  x_2420 & ~n_25672;
assign n_30707 =  i_25 &  n_25672;
assign n_30708 = ~n_30706 & ~n_30707;
assign n_30709 =  x_2420 & ~n_30708;
assign n_30710 = ~x_2420 &  n_30708;
assign n_30711 = ~n_30709 & ~n_30710;
assign n_30712 =  x_2419 & ~n_25672;
assign n_30713 =  i_24 &  n_25672;
assign n_30714 = ~n_30712 & ~n_30713;
assign n_30715 =  x_2419 & ~n_30714;
assign n_30716 = ~x_2419 &  n_30714;
assign n_30717 = ~n_30715 & ~n_30716;
assign n_30718 =  x_2418 & ~n_25672;
assign n_30719 =  i_23 &  n_25672;
assign n_30720 = ~n_30718 & ~n_30719;
assign n_30721 =  x_2418 & ~n_30720;
assign n_30722 = ~x_2418 &  n_30720;
assign n_30723 = ~n_30721 & ~n_30722;
assign n_30724 =  x_2417 & ~n_25672;
assign n_30725 =  i_22 &  n_25672;
assign n_30726 = ~n_30724 & ~n_30725;
assign n_30727 =  x_2417 & ~n_30726;
assign n_30728 = ~x_2417 &  n_30726;
assign n_30729 = ~n_30727 & ~n_30728;
assign n_30730 =  x_2416 & ~n_25672;
assign n_30731 =  i_21 &  n_25672;
assign n_30732 = ~n_30730 & ~n_30731;
assign n_30733 =  x_2416 & ~n_30732;
assign n_30734 = ~x_2416 &  n_30732;
assign n_30735 = ~n_30733 & ~n_30734;
assign n_30736 =  x_2415 & ~n_25672;
assign n_30737 =  i_20 &  n_25672;
assign n_30738 = ~n_30736 & ~n_30737;
assign n_30739 =  x_2415 & ~n_30738;
assign n_30740 = ~x_2415 &  n_30738;
assign n_30741 = ~n_30739 & ~n_30740;
assign n_30742 =  x_2414 & ~n_25672;
assign n_30743 =  i_19 &  n_25672;
assign n_30744 = ~n_30742 & ~n_30743;
assign n_30745 =  x_2414 & ~n_30744;
assign n_30746 = ~x_2414 &  n_30744;
assign n_30747 = ~n_30745 & ~n_30746;
assign n_30748 =  x_2413 & ~n_25672;
assign n_30749 =  i_18 &  n_25672;
assign n_30750 = ~n_30748 & ~n_30749;
assign n_30751 =  x_2413 & ~n_30750;
assign n_30752 = ~x_2413 &  n_30750;
assign n_30753 = ~n_30751 & ~n_30752;
assign n_30754 =  x_2412 & ~n_25672;
assign n_30755 =  i_17 &  n_25672;
assign n_30756 = ~n_30754 & ~n_30755;
assign n_30757 =  x_2412 & ~n_30756;
assign n_30758 = ~x_2412 &  n_30756;
assign n_30759 = ~n_30757 & ~n_30758;
assign n_30760 =  x_2411 & ~n_25672;
assign n_30761 =  i_16 &  n_25672;
assign n_30762 = ~n_30760 & ~n_30761;
assign n_30763 =  x_2411 & ~n_30762;
assign n_30764 = ~x_2411 &  n_30762;
assign n_30765 = ~n_30763 & ~n_30764;
assign n_30766 =  x_2410 & ~n_25672;
assign n_30767 =  i_15 &  n_25672;
assign n_30768 = ~n_30766 & ~n_30767;
assign n_30769 =  x_2410 & ~n_30768;
assign n_30770 = ~x_2410 &  n_30768;
assign n_30771 = ~n_30769 & ~n_30770;
assign n_30772 =  x_2409 & ~n_25672;
assign n_30773 =  i_14 &  n_25672;
assign n_30774 = ~n_30772 & ~n_30773;
assign n_30775 =  x_2409 & ~n_30774;
assign n_30776 = ~x_2409 &  n_30774;
assign n_30777 = ~n_30775 & ~n_30776;
assign n_30778 =  x_2408 & ~n_25672;
assign n_30779 =  i_13 &  n_25672;
assign n_30780 = ~n_30778 & ~n_30779;
assign n_30781 =  x_2408 & ~n_30780;
assign n_30782 = ~x_2408 &  n_30780;
assign n_30783 = ~n_30781 & ~n_30782;
assign n_30784 =  x_2407 & ~n_25672;
assign n_30785 =  i_12 &  n_25672;
assign n_30786 = ~n_30784 & ~n_30785;
assign n_30787 =  x_2407 & ~n_30786;
assign n_30788 = ~x_2407 &  n_30786;
assign n_30789 = ~n_30787 & ~n_30788;
assign n_30790 =  x_2406 & ~n_25672;
assign n_30791 =  i_11 &  n_25672;
assign n_30792 = ~n_30790 & ~n_30791;
assign n_30793 =  x_2406 & ~n_30792;
assign n_30794 = ~x_2406 &  n_30792;
assign n_30795 = ~n_30793 & ~n_30794;
assign n_30796 =  x_2405 & ~n_25672;
assign n_30797 =  i_10 &  n_25672;
assign n_30798 = ~n_30796 & ~n_30797;
assign n_30799 =  x_2405 & ~n_30798;
assign n_30800 = ~x_2405 &  n_30798;
assign n_30801 = ~n_30799 & ~n_30800;
assign n_30802 =  x_2404 & ~n_25672;
assign n_30803 =  i_9 &  n_25672;
assign n_30804 = ~n_30802 & ~n_30803;
assign n_30805 =  x_2404 & ~n_30804;
assign n_30806 = ~x_2404 &  n_30804;
assign n_30807 = ~n_30805 & ~n_30806;
assign n_30808 =  x_2403 & ~n_25672;
assign n_30809 =  i_8 &  n_25672;
assign n_30810 = ~n_30808 & ~n_30809;
assign n_30811 =  x_2403 & ~n_30810;
assign n_30812 = ~x_2403 &  n_30810;
assign n_30813 = ~n_30811 & ~n_30812;
assign n_30814 =  x_2402 & ~n_25672;
assign n_30815 =  i_7 &  n_25672;
assign n_30816 = ~n_30814 & ~n_30815;
assign n_30817 =  x_2402 & ~n_30816;
assign n_30818 = ~x_2402 &  n_30816;
assign n_30819 = ~n_30817 & ~n_30818;
assign n_30820 =  x_2401 & ~n_25672;
assign n_30821 =  i_6 &  n_25672;
assign n_30822 = ~n_30820 & ~n_30821;
assign n_30823 =  x_2401 & ~n_30822;
assign n_30824 = ~x_2401 &  n_30822;
assign n_30825 = ~n_30823 & ~n_30824;
assign n_30826 =  x_2400 & ~n_25672;
assign n_30827 =  i_5 &  n_25672;
assign n_30828 = ~n_30826 & ~n_30827;
assign n_30829 =  x_2400 & ~n_30828;
assign n_30830 = ~x_2400 &  n_30828;
assign n_30831 = ~n_30829 & ~n_30830;
assign n_30832 =  x_2399 & ~n_25672;
assign n_30833 =  i_4 &  n_25672;
assign n_30834 = ~n_30832 & ~n_30833;
assign n_30835 =  x_2399 & ~n_30834;
assign n_30836 = ~x_2399 &  n_30834;
assign n_30837 = ~n_30835 & ~n_30836;
assign n_30838 =  x_2398 & ~n_25672;
assign n_30839 =  i_3 &  n_25672;
assign n_30840 = ~n_30838 & ~n_30839;
assign n_30841 =  x_2398 & ~n_30840;
assign n_30842 = ~x_2398 &  n_30840;
assign n_30843 = ~n_30841 & ~n_30842;
assign n_30844 =  x_2397 & ~n_25672;
assign n_30845 =  i_2 &  n_25672;
assign n_30846 = ~n_30844 & ~n_30845;
assign n_30847 =  x_2397 & ~n_30846;
assign n_30848 = ~x_2397 &  n_30846;
assign n_30849 = ~n_30847 & ~n_30848;
assign n_30850 =  x_2396 & ~n_25672;
assign n_30851 =  i_1 &  n_25672;
assign n_30852 = ~n_30850 & ~n_30851;
assign n_30853 =  x_2396 & ~n_30852;
assign n_30854 = ~x_2396 &  n_30852;
assign n_30855 = ~n_30853 & ~n_30854;
assign n_30856 = ~n_23544 & ~n_24122;
assign n_30857 = ~n_24950 & ~n_24932;
assign n_30858 = ~n_24230 &  n_30856;
assign n_30859 =  n_30857 &  n_30858;
assign n_30860 =  x_2395 &  n_30859;
assign n_30861 =  n_30856 & ~n_30860;
assign n_30862 =  x_2395 & ~n_30861;
assign n_30863 = ~x_2395 &  n_30861;
assign n_30864 = ~n_30862 & ~n_30863;
assign n_30865 =  x_2394 &  n_30858;
assign n_30866 =  n_30857 & ~n_30865;
assign n_30867 =  x_2394 & ~n_30866;
assign n_30868 = ~x_2394 &  n_30866;
assign n_30869 = ~n_30867 & ~n_30868;
assign n_30870 =  x_2393 &  n_30859;
assign n_30871 = ~n_24230 & ~n_24122;
assign n_30872 = ~n_24950 &  n_30871;
assign n_30873 = ~n_30870 &  n_30872;
assign n_30874 =  x_2393 & ~n_30873;
assign n_30875 = ~x_2393 &  n_30873;
assign n_30876 = ~n_30874 & ~n_30875;
assign n_30877 =  x_2392 &  n_30859;
assign n_30878 =  x_2392 &  n_30877;
assign n_30879 = ~x_2392 & ~n_30877;
assign n_30880 = ~n_30878 & ~n_30879;
assign n_30881 =  x_2391 &  n_30859;
assign n_30882 =  x_2391 &  n_30881;
assign n_30883 = ~x_2391 & ~n_30881;
assign n_30884 = ~n_30882 & ~n_30883;
assign n_30885 =  x_2390 &  n_30859;
assign n_30886 =  x_2390 &  n_30885;
assign n_30887 = ~x_2390 & ~n_30885;
assign n_30888 = ~n_30886 & ~n_30887;
assign n_30889 =  x_2389 &  n_30859;
assign n_30890 =  x_2389 &  n_30889;
assign n_30891 = ~x_2389 & ~n_30889;
assign n_30892 = ~n_30890 & ~n_30891;
assign n_30893 =  x_2388 &  n_30859;
assign n_30894 =  x_2388 &  n_30893;
assign n_30895 = ~x_2388 & ~n_30893;
assign n_30896 = ~n_30894 & ~n_30895;
assign n_30897 =  x_2387 &  n_30859;
assign n_30898 =  x_2387 &  n_30897;
assign n_30899 = ~x_2387 & ~n_30897;
assign n_30900 = ~n_30898 & ~n_30899;
assign n_30901 =  x_2386 &  n_30859;
assign n_30902 =  x_2386 &  n_30901;
assign n_30903 = ~x_2386 & ~n_30901;
assign n_30904 = ~n_30902 & ~n_30903;
assign n_30905 =  x_2385 &  n_30859;
assign n_30906 =  x_2385 &  n_30905;
assign n_30907 = ~x_2385 & ~n_30905;
assign n_30908 = ~n_30906 & ~n_30907;
assign n_30909 =  x_2384 &  n_30859;
assign n_30910 =  x_2384 &  n_30909;
assign n_30911 = ~x_2384 & ~n_30909;
assign n_30912 = ~n_30910 & ~n_30911;
assign n_30913 =  x_2383 &  n_30859;
assign n_30914 =  x_2383 &  n_30913;
assign n_30915 = ~x_2383 & ~n_30913;
assign n_30916 = ~n_30914 & ~n_30915;
assign n_30917 =  x_2382 &  n_30859;
assign n_30918 =  x_2382 &  n_30917;
assign n_30919 = ~x_2382 & ~n_30917;
assign n_30920 = ~n_30918 & ~n_30919;
assign n_30921 =  x_2381 &  n_30859;
assign n_30922 =  x_2381 &  n_30921;
assign n_30923 = ~x_2381 & ~n_30921;
assign n_30924 = ~n_30922 & ~n_30923;
assign n_30925 =  x_2380 &  n_30859;
assign n_30926 =  x_2380 &  n_30925;
assign n_30927 = ~x_2380 & ~n_30925;
assign n_30928 = ~n_30926 & ~n_30927;
assign n_30929 =  x_2379 &  n_30859;
assign n_30930 =  x_2379 &  n_30929;
assign n_30931 = ~x_2379 & ~n_30929;
assign n_30932 = ~n_30930 & ~n_30931;
assign n_30933 =  x_2378 & ~n_24021;
assign n_30934 =  i_32 &  n_24021;
assign n_30935 = ~n_30933 & ~n_30934;
assign n_30936 =  x_2378 & ~n_30935;
assign n_30937 = ~x_2378 &  n_30935;
assign n_30938 = ~n_30936 & ~n_30937;
assign n_30939 =  x_2377 & ~n_24021;
assign n_30940 =  i_31 &  n_24021;
assign n_30941 = ~n_30939 & ~n_30940;
assign n_30942 =  x_2377 & ~n_30941;
assign n_30943 = ~x_2377 &  n_30941;
assign n_30944 = ~n_30942 & ~n_30943;
assign n_30945 =  x_2376 & ~n_24021;
assign n_30946 =  i_30 &  n_24021;
assign n_30947 = ~n_30945 & ~n_30946;
assign n_30948 =  x_2376 & ~n_30947;
assign n_30949 = ~x_2376 &  n_30947;
assign n_30950 = ~n_30948 & ~n_30949;
assign n_30951 =  x_2375 & ~n_24021;
assign n_30952 =  i_29 &  n_24021;
assign n_30953 = ~n_30951 & ~n_30952;
assign n_30954 =  x_2375 & ~n_30953;
assign n_30955 = ~x_2375 &  n_30953;
assign n_30956 = ~n_30954 & ~n_30955;
assign n_30957 =  x_2374 & ~n_24021;
assign n_30958 =  i_28 &  n_24021;
assign n_30959 = ~n_30957 & ~n_30958;
assign n_30960 =  x_2374 & ~n_30959;
assign n_30961 = ~x_2374 &  n_30959;
assign n_30962 = ~n_30960 & ~n_30961;
assign n_30963 =  x_2373 & ~n_24021;
assign n_30964 =  i_27 &  n_24021;
assign n_30965 = ~n_30963 & ~n_30964;
assign n_30966 =  x_2373 & ~n_30965;
assign n_30967 = ~x_2373 &  n_30965;
assign n_30968 = ~n_30966 & ~n_30967;
assign n_30969 =  x_2372 & ~n_24021;
assign n_30970 =  i_26 &  n_24021;
assign n_30971 = ~n_30969 & ~n_30970;
assign n_30972 =  x_2372 & ~n_30971;
assign n_30973 = ~x_2372 &  n_30971;
assign n_30974 = ~n_30972 & ~n_30973;
assign n_30975 =  x_2371 & ~n_24021;
assign n_30976 =  i_25 &  n_24021;
assign n_30977 = ~n_30975 & ~n_30976;
assign n_30978 =  x_2371 & ~n_30977;
assign n_30979 = ~x_2371 &  n_30977;
assign n_30980 = ~n_30978 & ~n_30979;
assign n_30981 =  x_2370 & ~n_24021;
assign n_30982 =  i_24 &  n_24021;
assign n_30983 = ~n_30981 & ~n_30982;
assign n_30984 =  x_2370 & ~n_30983;
assign n_30985 = ~x_2370 &  n_30983;
assign n_30986 = ~n_30984 & ~n_30985;
assign n_30987 =  x_2369 & ~n_24021;
assign n_30988 =  i_23 &  n_24021;
assign n_30989 = ~n_30987 & ~n_30988;
assign n_30990 =  x_2369 & ~n_30989;
assign n_30991 = ~x_2369 &  n_30989;
assign n_30992 = ~n_30990 & ~n_30991;
assign n_30993 =  x_2368 & ~n_24021;
assign n_30994 =  i_22 &  n_24021;
assign n_30995 = ~n_30993 & ~n_30994;
assign n_30996 =  x_2368 & ~n_30995;
assign n_30997 = ~x_2368 &  n_30995;
assign n_30998 = ~n_30996 & ~n_30997;
assign n_30999 =  x_2367 & ~n_24021;
assign n_31000 =  i_21 &  n_24021;
assign n_31001 = ~n_30999 & ~n_31000;
assign n_31002 =  x_2367 & ~n_31001;
assign n_31003 = ~x_2367 &  n_31001;
assign n_31004 = ~n_31002 & ~n_31003;
assign n_31005 =  x_2366 & ~n_24021;
assign n_31006 =  i_20 &  n_24021;
assign n_31007 = ~n_31005 & ~n_31006;
assign n_31008 =  x_2366 & ~n_31007;
assign n_31009 = ~x_2366 &  n_31007;
assign n_31010 = ~n_31008 & ~n_31009;
assign n_31011 =  x_2365 & ~n_24021;
assign n_31012 =  i_19 &  n_24021;
assign n_31013 = ~n_31011 & ~n_31012;
assign n_31014 =  x_2365 & ~n_31013;
assign n_31015 = ~x_2365 &  n_31013;
assign n_31016 = ~n_31014 & ~n_31015;
assign n_31017 =  x_2364 & ~n_24021;
assign n_31018 =  i_18 &  n_24021;
assign n_31019 = ~n_31017 & ~n_31018;
assign n_31020 =  x_2364 & ~n_31019;
assign n_31021 = ~x_2364 &  n_31019;
assign n_31022 = ~n_31020 & ~n_31021;
assign n_31023 =  x_2363 & ~n_24021;
assign n_31024 =  i_17 &  n_24021;
assign n_31025 = ~n_31023 & ~n_31024;
assign n_31026 =  x_2363 & ~n_31025;
assign n_31027 = ~x_2363 &  n_31025;
assign n_31028 = ~n_31026 & ~n_31027;
assign n_31029 =  x_2362 & ~n_24021;
assign n_31030 =  i_16 &  n_24021;
assign n_31031 = ~n_31029 & ~n_31030;
assign n_31032 =  x_2362 & ~n_31031;
assign n_31033 = ~x_2362 &  n_31031;
assign n_31034 = ~n_31032 & ~n_31033;
assign n_31035 =  x_2361 & ~n_24021;
assign n_31036 =  i_15 &  n_24021;
assign n_31037 = ~n_31035 & ~n_31036;
assign n_31038 =  x_2361 & ~n_31037;
assign n_31039 = ~x_2361 &  n_31037;
assign n_31040 = ~n_31038 & ~n_31039;
assign n_31041 =  x_2360 & ~n_24021;
assign n_31042 =  i_14 &  n_24021;
assign n_31043 = ~n_31041 & ~n_31042;
assign n_31044 =  x_2360 & ~n_31043;
assign n_31045 = ~x_2360 &  n_31043;
assign n_31046 = ~n_31044 & ~n_31045;
assign n_31047 =  x_2359 & ~n_24021;
assign n_31048 =  i_13 &  n_24021;
assign n_31049 = ~n_31047 & ~n_31048;
assign n_31050 =  x_2359 & ~n_31049;
assign n_31051 = ~x_2359 &  n_31049;
assign n_31052 = ~n_31050 & ~n_31051;
assign n_31053 =  x_2358 & ~n_24021;
assign n_31054 =  i_12 &  n_24021;
assign n_31055 = ~n_31053 & ~n_31054;
assign n_31056 =  x_2358 & ~n_31055;
assign n_31057 = ~x_2358 &  n_31055;
assign n_31058 = ~n_31056 & ~n_31057;
assign n_31059 =  x_2357 & ~n_24021;
assign n_31060 =  i_11 &  n_24021;
assign n_31061 = ~n_31059 & ~n_31060;
assign n_31062 =  x_2357 & ~n_31061;
assign n_31063 = ~x_2357 &  n_31061;
assign n_31064 = ~n_31062 & ~n_31063;
assign n_31065 =  x_2356 & ~n_24021;
assign n_31066 =  i_10 &  n_24021;
assign n_31067 = ~n_31065 & ~n_31066;
assign n_31068 =  x_2356 & ~n_31067;
assign n_31069 = ~x_2356 &  n_31067;
assign n_31070 = ~n_31068 & ~n_31069;
assign n_31071 =  x_2355 & ~n_24021;
assign n_31072 =  i_9 &  n_24021;
assign n_31073 = ~n_31071 & ~n_31072;
assign n_31074 =  x_2355 & ~n_31073;
assign n_31075 = ~x_2355 &  n_31073;
assign n_31076 = ~n_31074 & ~n_31075;
assign n_31077 =  x_2354 & ~n_24021;
assign n_31078 =  i_8 &  n_24021;
assign n_31079 = ~n_31077 & ~n_31078;
assign n_31080 =  x_2354 & ~n_31079;
assign n_31081 = ~x_2354 &  n_31079;
assign n_31082 = ~n_31080 & ~n_31081;
assign n_31083 =  x_2353 & ~n_24021;
assign n_31084 =  i_7 &  n_24021;
assign n_31085 = ~n_31083 & ~n_31084;
assign n_31086 =  x_2353 & ~n_31085;
assign n_31087 = ~x_2353 &  n_31085;
assign n_31088 = ~n_31086 & ~n_31087;
assign n_31089 =  x_2352 & ~n_24021;
assign n_31090 =  i_6 &  n_24021;
assign n_31091 = ~n_31089 & ~n_31090;
assign n_31092 =  x_2352 & ~n_31091;
assign n_31093 = ~x_2352 &  n_31091;
assign n_31094 = ~n_31092 & ~n_31093;
assign n_31095 =  x_2351 & ~n_24021;
assign n_31096 =  i_5 &  n_24021;
assign n_31097 = ~n_31095 & ~n_31096;
assign n_31098 =  x_2351 & ~n_31097;
assign n_31099 = ~x_2351 &  n_31097;
assign n_31100 = ~n_31098 & ~n_31099;
assign n_31101 =  x_2350 & ~n_24021;
assign n_31102 =  i_4 &  n_24021;
assign n_31103 = ~n_31101 & ~n_31102;
assign n_31104 =  x_2350 & ~n_31103;
assign n_31105 = ~x_2350 &  n_31103;
assign n_31106 = ~n_31104 & ~n_31105;
assign n_31107 =  x_2349 & ~n_24021;
assign n_31108 =  i_3 &  n_24021;
assign n_31109 = ~n_31107 & ~n_31108;
assign n_31110 =  x_2349 & ~n_31109;
assign n_31111 = ~x_2349 &  n_31109;
assign n_31112 = ~n_31110 & ~n_31111;
assign n_31113 =  x_2348 & ~n_24021;
assign n_31114 =  i_2 &  n_24021;
assign n_31115 = ~n_31113 & ~n_31114;
assign n_31116 =  x_2348 & ~n_31115;
assign n_31117 = ~x_2348 &  n_31115;
assign n_31118 = ~n_31116 & ~n_31117;
assign n_31119 =  x_2347 & ~n_24021;
assign n_31120 =  i_1 &  n_24021;
assign n_31121 = ~n_31119 & ~n_31120;
assign n_31122 =  x_2347 & ~n_31121;
assign n_31123 = ~x_2347 &  n_31121;
assign n_31124 = ~n_31122 & ~n_31123;
assign n_31125 =  n_553 &  n_23175;
assign n_31126 =  n_6180 &  n_357;
assign n_31127 = ~n_31125 & ~n_31126;
assign n_31128 =  x_43 & ~n_31127;
assign n_31129 =  x_2346 & ~n_31128;
assign n_31130 =  i_32 &  n_31128;
assign n_31131 = ~n_31129 & ~n_31130;
assign n_31132 =  x_2346 & ~n_31131;
assign n_31133 = ~x_2346 &  n_31131;
assign n_31134 = ~n_31132 & ~n_31133;
assign n_31135 =  x_2345 & ~n_31128;
assign n_31136 =  i_31 &  n_31128;
assign n_31137 = ~n_31135 & ~n_31136;
assign n_31138 =  x_2345 & ~n_31137;
assign n_31139 = ~x_2345 &  n_31137;
assign n_31140 = ~n_31138 & ~n_31139;
assign n_31141 =  x_2344 & ~n_31128;
assign n_31142 =  i_30 &  n_31128;
assign n_31143 = ~n_31141 & ~n_31142;
assign n_31144 =  x_2344 & ~n_31143;
assign n_31145 = ~x_2344 &  n_31143;
assign n_31146 = ~n_31144 & ~n_31145;
assign n_31147 =  x_2343 & ~n_31128;
assign n_31148 =  i_29 &  n_31128;
assign n_31149 = ~n_31147 & ~n_31148;
assign n_31150 =  x_2343 & ~n_31149;
assign n_31151 = ~x_2343 &  n_31149;
assign n_31152 = ~n_31150 & ~n_31151;
assign n_31153 =  x_2342 & ~n_31128;
assign n_31154 =  i_28 &  n_31128;
assign n_31155 = ~n_31153 & ~n_31154;
assign n_31156 =  x_2342 & ~n_31155;
assign n_31157 = ~x_2342 &  n_31155;
assign n_31158 = ~n_31156 & ~n_31157;
assign n_31159 =  x_2341 & ~n_31128;
assign n_31160 =  i_27 &  n_31128;
assign n_31161 = ~n_31159 & ~n_31160;
assign n_31162 =  x_2341 & ~n_31161;
assign n_31163 = ~x_2341 &  n_31161;
assign n_31164 = ~n_31162 & ~n_31163;
assign n_31165 =  x_2340 & ~n_31128;
assign n_31166 =  i_26 &  n_31128;
assign n_31167 = ~n_31165 & ~n_31166;
assign n_31168 =  x_2340 & ~n_31167;
assign n_31169 = ~x_2340 &  n_31167;
assign n_31170 = ~n_31168 & ~n_31169;
assign n_31171 =  x_2339 & ~n_31128;
assign n_31172 =  i_25 &  n_31128;
assign n_31173 = ~n_31171 & ~n_31172;
assign n_31174 =  x_2339 & ~n_31173;
assign n_31175 = ~x_2339 &  n_31173;
assign n_31176 = ~n_31174 & ~n_31175;
assign n_31177 =  x_2338 & ~n_31128;
assign n_31178 =  i_24 &  n_31128;
assign n_31179 = ~n_31177 & ~n_31178;
assign n_31180 =  x_2338 & ~n_31179;
assign n_31181 = ~x_2338 &  n_31179;
assign n_31182 = ~n_31180 & ~n_31181;
assign n_31183 =  x_2337 & ~n_31128;
assign n_31184 =  i_23 &  n_31128;
assign n_31185 = ~n_31183 & ~n_31184;
assign n_31186 =  x_2337 & ~n_31185;
assign n_31187 = ~x_2337 &  n_31185;
assign n_31188 = ~n_31186 & ~n_31187;
assign n_31189 =  x_2336 & ~n_31128;
assign n_31190 =  i_22 &  n_31128;
assign n_31191 = ~n_31189 & ~n_31190;
assign n_31192 =  x_2336 & ~n_31191;
assign n_31193 = ~x_2336 &  n_31191;
assign n_31194 = ~n_31192 & ~n_31193;
assign n_31195 =  x_2335 & ~n_31128;
assign n_31196 =  i_21 &  n_31128;
assign n_31197 = ~n_31195 & ~n_31196;
assign n_31198 =  x_2335 & ~n_31197;
assign n_31199 = ~x_2335 &  n_31197;
assign n_31200 = ~n_31198 & ~n_31199;
assign n_31201 =  x_2334 & ~n_31128;
assign n_31202 =  i_20 &  n_31128;
assign n_31203 = ~n_31201 & ~n_31202;
assign n_31204 =  x_2334 & ~n_31203;
assign n_31205 = ~x_2334 &  n_31203;
assign n_31206 = ~n_31204 & ~n_31205;
assign n_31207 =  x_2333 & ~n_31128;
assign n_31208 =  i_19 &  n_31128;
assign n_31209 = ~n_31207 & ~n_31208;
assign n_31210 =  x_2333 & ~n_31209;
assign n_31211 = ~x_2333 &  n_31209;
assign n_31212 = ~n_31210 & ~n_31211;
assign n_31213 =  x_2332 & ~n_31128;
assign n_31214 =  i_18 &  n_31128;
assign n_31215 = ~n_31213 & ~n_31214;
assign n_31216 =  x_2332 & ~n_31215;
assign n_31217 = ~x_2332 &  n_31215;
assign n_31218 = ~n_31216 & ~n_31217;
assign n_31219 =  x_2331 & ~n_31128;
assign n_31220 =  i_17 &  n_31128;
assign n_31221 = ~n_31219 & ~n_31220;
assign n_31222 =  x_2331 & ~n_31221;
assign n_31223 = ~x_2331 &  n_31221;
assign n_31224 = ~n_31222 & ~n_31223;
assign n_31225 =  x_2330 & ~n_31128;
assign n_31226 =  i_16 &  n_31128;
assign n_31227 = ~n_31225 & ~n_31226;
assign n_31228 =  x_2330 & ~n_31227;
assign n_31229 = ~x_2330 &  n_31227;
assign n_31230 = ~n_31228 & ~n_31229;
assign n_31231 =  x_2329 & ~n_31128;
assign n_31232 =  i_15 &  n_31128;
assign n_31233 = ~n_31231 & ~n_31232;
assign n_31234 =  x_2329 & ~n_31233;
assign n_31235 = ~x_2329 &  n_31233;
assign n_31236 = ~n_31234 & ~n_31235;
assign n_31237 =  x_2328 & ~n_31128;
assign n_31238 =  i_14 &  n_31128;
assign n_31239 = ~n_31237 & ~n_31238;
assign n_31240 =  x_2328 & ~n_31239;
assign n_31241 = ~x_2328 &  n_31239;
assign n_31242 = ~n_31240 & ~n_31241;
assign n_31243 =  x_2327 & ~n_31128;
assign n_31244 =  i_13 &  n_31128;
assign n_31245 = ~n_31243 & ~n_31244;
assign n_31246 =  x_2327 & ~n_31245;
assign n_31247 = ~x_2327 &  n_31245;
assign n_31248 = ~n_31246 & ~n_31247;
assign n_31249 =  x_2326 & ~n_31128;
assign n_31250 =  i_12 &  n_31128;
assign n_31251 = ~n_31249 & ~n_31250;
assign n_31252 =  x_2326 & ~n_31251;
assign n_31253 = ~x_2326 &  n_31251;
assign n_31254 = ~n_31252 & ~n_31253;
assign n_31255 =  x_2325 & ~n_31128;
assign n_31256 =  i_11 &  n_31128;
assign n_31257 = ~n_31255 & ~n_31256;
assign n_31258 =  x_2325 & ~n_31257;
assign n_31259 = ~x_2325 &  n_31257;
assign n_31260 = ~n_31258 & ~n_31259;
assign n_31261 =  x_2324 & ~n_31128;
assign n_31262 =  i_10 &  n_31128;
assign n_31263 = ~n_31261 & ~n_31262;
assign n_31264 =  x_2324 & ~n_31263;
assign n_31265 = ~x_2324 &  n_31263;
assign n_31266 = ~n_31264 & ~n_31265;
assign n_31267 =  x_2323 & ~n_31128;
assign n_31268 =  i_9 &  n_31128;
assign n_31269 = ~n_31267 & ~n_31268;
assign n_31270 =  x_2323 & ~n_31269;
assign n_31271 = ~x_2323 &  n_31269;
assign n_31272 = ~n_31270 & ~n_31271;
assign n_31273 =  x_2322 & ~n_31128;
assign n_31274 =  i_8 &  n_31128;
assign n_31275 = ~n_31273 & ~n_31274;
assign n_31276 =  x_2322 & ~n_31275;
assign n_31277 = ~x_2322 &  n_31275;
assign n_31278 = ~n_31276 & ~n_31277;
assign n_31279 =  x_2321 & ~n_31128;
assign n_31280 =  i_7 &  n_31128;
assign n_31281 = ~n_31279 & ~n_31280;
assign n_31282 =  x_2321 & ~n_31281;
assign n_31283 = ~x_2321 &  n_31281;
assign n_31284 = ~n_31282 & ~n_31283;
assign n_31285 =  x_2320 & ~n_31128;
assign n_31286 =  i_6 &  n_31128;
assign n_31287 = ~n_31285 & ~n_31286;
assign n_31288 =  x_2320 & ~n_31287;
assign n_31289 = ~x_2320 &  n_31287;
assign n_31290 = ~n_31288 & ~n_31289;
assign n_31291 =  x_2319 & ~n_31128;
assign n_31292 =  i_5 &  n_31128;
assign n_31293 = ~n_31291 & ~n_31292;
assign n_31294 =  x_2319 & ~n_31293;
assign n_31295 = ~x_2319 &  n_31293;
assign n_31296 = ~n_31294 & ~n_31295;
assign n_31297 =  x_2318 & ~n_31128;
assign n_31298 =  i_4 &  n_31128;
assign n_31299 = ~n_31297 & ~n_31298;
assign n_31300 =  x_2318 & ~n_31299;
assign n_31301 = ~x_2318 &  n_31299;
assign n_31302 = ~n_31300 & ~n_31301;
assign n_31303 =  x_2317 & ~n_31128;
assign n_31304 =  i_3 &  n_31128;
assign n_31305 = ~n_31303 & ~n_31304;
assign n_31306 =  x_2317 & ~n_31305;
assign n_31307 = ~x_2317 &  n_31305;
assign n_31308 = ~n_31306 & ~n_31307;
assign n_31309 =  x_2316 & ~n_31128;
assign n_31310 =  i_2 &  n_31128;
assign n_31311 = ~n_31309 & ~n_31310;
assign n_31312 =  x_2316 & ~n_31311;
assign n_31313 = ~x_2316 &  n_31311;
assign n_31314 = ~n_31312 & ~n_31313;
assign n_31315 =  x_2315 & ~n_31128;
assign n_31316 =  i_1 &  n_31128;
assign n_31317 = ~n_31315 & ~n_31316;
assign n_31318 =  x_2315 & ~n_31317;
assign n_31319 = ~x_2315 &  n_31317;
assign n_31320 = ~n_31318 & ~n_31319;
assign n_31321 =  x_2314 & ~n_1901;
assign n_31322 =  x_1066 &  n_1901;
assign n_31323 = ~n_31321 & ~n_31322;
assign n_31324 =  x_2314 & ~n_31323;
assign n_31325 = ~x_2314 &  n_31323;
assign n_31326 = ~n_31324 & ~n_31325;
assign n_31327 =  x_2313 & ~n_1901;
assign n_31328 =  x_1065 &  n_1901;
assign n_31329 = ~n_31327 & ~n_31328;
assign n_31330 =  x_2313 & ~n_31329;
assign n_31331 = ~x_2313 &  n_31329;
assign n_31332 = ~n_31330 & ~n_31331;
assign n_31333 =  x_2312 & ~n_1901;
assign n_31334 =  x_1064 &  n_1901;
assign n_31335 = ~n_31333 & ~n_31334;
assign n_31336 =  x_2312 & ~n_31335;
assign n_31337 = ~x_2312 &  n_31335;
assign n_31338 = ~n_31336 & ~n_31337;
assign n_31339 =  x_2311 & ~n_1901;
assign n_31340 =  x_1063 &  n_1901;
assign n_31341 = ~n_31339 & ~n_31340;
assign n_31342 =  x_2311 & ~n_31341;
assign n_31343 = ~x_2311 &  n_31341;
assign n_31344 = ~n_31342 & ~n_31343;
assign n_31345 =  x_2310 & ~n_1901;
assign n_31346 =  x_1062 &  n_1901;
assign n_31347 = ~n_31345 & ~n_31346;
assign n_31348 =  x_2310 & ~n_31347;
assign n_31349 = ~x_2310 &  n_31347;
assign n_31350 = ~n_31348 & ~n_31349;
assign n_31351 =  x_2309 & ~n_1901;
assign n_31352 =  x_1061 &  n_1901;
assign n_31353 = ~n_31351 & ~n_31352;
assign n_31354 =  x_2309 & ~n_31353;
assign n_31355 = ~x_2309 &  n_31353;
assign n_31356 = ~n_31354 & ~n_31355;
assign n_31357 =  x_2308 & ~n_1901;
assign n_31358 =  x_1060 &  n_1901;
assign n_31359 = ~n_31357 & ~n_31358;
assign n_31360 =  x_2308 & ~n_31359;
assign n_31361 = ~x_2308 &  n_31359;
assign n_31362 = ~n_31360 & ~n_31361;
assign n_31363 =  x_2307 & ~n_1901;
assign n_31364 =  x_1059 &  n_1901;
assign n_31365 = ~n_31363 & ~n_31364;
assign n_31366 =  x_2307 & ~n_31365;
assign n_31367 = ~x_2307 &  n_31365;
assign n_31368 = ~n_31366 & ~n_31367;
assign n_31369 =  x_2306 & ~n_1901;
assign n_31370 =  x_1058 &  n_1901;
assign n_31371 = ~n_31369 & ~n_31370;
assign n_31372 =  x_2306 & ~n_31371;
assign n_31373 = ~x_2306 &  n_31371;
assign n_31374 = ~n_31372 & ~n_31373;
assign n_31375 =  x_2305 & ~n_1901;
assign n_31376 =  x_1057 &  n_1901;
assign n_31377 = ~n_31375 & ~n_31376;
assign n_31378 =  x_2305 & ~n_31377;
assign n_31379 = ~x_2305 &  n_31377;
assign n_31380 = ~n_31378 & ~n_31379;
assign n_31381 =  x_2304 & ~n_1901;
assign n_31382 =  x_1056 &  n_1901;
assign n_31383 = ~n_31381 & ~n_31382;
assign n_31384 =  x_2304 & ~n_31383;
assign n_31385 = ~x_2304 &  n_31383;
assign n_31386 = ~n_31384 & ~n_31385;
assign n_31387 =  x_2303 & ~n_1901;
assign n_31388 =  x_1055 &  n_1901;
assign n_31389 = ~n_31387 & ~n_31388;
assign n_31390 =  x_2303 & ~n_31389;
assign n_31391 = ~x_2303 &  n_31389;
assign n_31392 = ~n_31390 & ~n_31391;
assign n_31393 =  x_2302 & ~n_1901;
assign n_31394 =  x_1054 &  n_1901;
assign n_31395 = ~n_31393 & ~n_31394;
assign n_31396 =  x_2302 & ~n_31395;
assign n_31397 = ~x_2302 &  n_31395;
assign n_31398 = ~n_31396 & ~n_31397;
assign n_31399 =  x_2301 & ~n_1901;
assign n_31400 =  x_1053 &  n_1901;
assign n_31401 = ~n_31399 & ~n_31400;
assign n_31402 =  x_2301 & ~n_31401;
assign n_31403 = ~x_2301 &  n_31401;
assign n_31404 = ~n_31402 & ~n_31403;
assign n_31405 =  x_2300 & ~n_1901;
assign n_31406 =  x_1052 &  n_1901;
assign n_31407 = ~n_31405 & ~n_31406;
assign n_31408 =  x_2300 & ~n_31407;
assign n_31409 = ~x_2300 &  n_31407;
assign n_31410 = ~n_31408 & ~n_31409;
assign n_31411 =  x_2299 & ~n_1901;
assign n_31412 =  x_1051 &  n_1901;
assign n_31413 = ~n_31411 & ~n_31412;
assign n_31414 =  x_2299 & ~n_31413;
assign n_31415 = ~x_2299 &  n_31413;
assign n_31416 = ~n_31414 & ~n_31415;
assign n_31417 =  x_2298 & ~n_1901;
assign n_31418 =  x_1050 &  n_1901;
assign n_31419 = ~n_31417 & ~n_31418;
assign n_31420 =  x_2298 & ~n_31419;
assign n_31421 = ~x_2298 &  n_31419;
assign n_31422 = ~n_31420 & ~n_31421;
assign n_31423 =  x_2297 & ~n_1901;
assign n_31424 =  x_1049 &  n_1901;
assign n_31425 = ~n_31423 & ~n_31424;
assign n_31426 =  x_2297 & ~n_31425;
assign n_31427 = ~x_2297 &  n_31425;
assign n_31428 = ~n_31426 & ~n_31427;
assign n_31429 =  x_2296 & ~n_1901;
assign n_31430 =  x_1048 &  n_1901;
assign n_31431 = ~n_31429 & ~n_31430;
assign n_31432 =  x_2296 & ~n_31431;
assign n_31433 = ~x_2296 &  n_31431;
assign n_31434 = ~n_31432 & ~n_31433;
assign n_31435 =  x_2295 & ~n_1901;
assign n_31436 =  x_1047 &  n_1901;
assign n_31437 = ~n_31435 & ~n_31436;
assign n_31438 =  x_2295 & ~n_31437;
assign n_31439 = ~x_2295 &  n_31437;
assign n_31440 = ~n_31438 & ~n_31439;
assign n_31441 =  x_2294 & ~n_1901;
assign n_31442 =  x_1046 &  n_1901;
assign n_31443 = ~n_31441 & ~n_31442;
assign n_31444 =  x_2294 & ~n_31443;
assign n_31445 = ~x_2294 &  n_31443;
assign n_31446 = ~n_31444 & ~n_31445;
assign n_31447 =  x_2293 & ~n_1901;
assign n_31448 =  x_1045 &  n_1901;
assign n_31449 = ~n_31447 & ~n_31448;
assign n_31450 =  x_2293 & ~n_31449;
assign n_31451 = ~x_2293 &  n_31449;
assign n_31452 = ~n_31450 & ~n_31451;
assign n_31453 =  x_2292 & ~n_1901;
assign n_31454 =  x_1044 &  n_1901;
assign n_31455 = ~n_31453 & ~n_31454;
assign n_31456 =  x_2292 & ~n_31455;
assign n_31457 = ~x_2292 &  n_31455;
assign n_31458 = ~n_31456 & ~n_31457;
assign n_31459 =  x_2291 & ~n_1901;
assign n_31460 =  x_1043 &  n_1901;
assign n_31461 = ~n_31459 & ~n_31460;
assign n_31462 =  x_2291 & ~n_31461;
assign n_31463 = ~x_2291 &  n_31461;
assign n_31464 = ~n_31462 & ~n_31463;
assign n_31465 =  x_2290 & ~n_1901;
assign n_31466 =  x_1042 &  n_1901;
assign n_31467 = ~n_31465 & ~n_31466;
assign n_31468 =  x_2290 & ~n_31467;
assign n_31469 = ~x_2290 &  n_31467;
assign n_31470 = ~n_31468 & ~n_31469;
assign n_31471 =  x_2289 & ~n_1901;
assign n_31472 =  x_1041 &  n_1901;
assign n_31473 = ~n_31471 & ~n_31472;
assign n_31474 =  x_2289 & ~n_31473;
assign n_31475 = ~x_2289 &  n_31473;
assign n_31476 = ~n_31474 & ~n_31475;
assign n_31477 =  x_2288 & ~n_1901;
assign n_31478 =  x_1040 &  n_1901;
assign n_31479 = ~n_31477 & ~n_31478;
assign n_31480 =  x_2288 & ~n_31479;
assign n_31481 = ~x_2288 &  n_31479;
assign n_31482 = ~n_31480 & ~n_31481;
assign n_31483 =  x_2287 & ~n_1901;
assign n_31484 =  x_1039 &  n_1901;
assign n_31485 = ~n_31483 & ~n_31484;
assign n_31486 =  x_2287 & ~n_31485;
assign n_31487 = ~x_2287 &  n_31485;
assign n_31488 = ~n_31486 & ~n_31487;
assign n_31489 =  x_2286 & ~n_1901;
assign n_31490 =  x_1038 &  n_1901;
assign n_31491 = ~n_31489 & ~n_31490;
assign n_31492 =  x_2286 & ~n_31491;
assign n_31493 = ~x_2286 &  n_31491;
assign n_31494 = ~n_31492 & ~n_31493;
assign n_31495 =  x_2285 & ~n_1901;
assign n_31496 =  x_1037 &  n_1901;
assign n_31497 = ~n_31495 & ~n_31496;
assign n_31498 =  x_2285 & ~n_31497;
assign n_31499 = ~x_2285 &  n_31497;
assign n_31500 = ~n_31498 & ~n_31499;
assign n_31501 =  x_2284 & ~n_1901;
assign n_31502 =  x_1036 &  n_1901;
assign n_31503 = ~n_31501 & ~n_31502;
assign n_31504 =  x_2284 & ~n_31503;
assign n_31505 = ~x_2284 &  n_31503;
assign n_31506 = ~n_31504 & ~n_31505;
assign n_31507 =  x_2283 & ~n_1901;
assign n_31508 =  x_1035 &  n_1901;
assign n_31509 = ~n_31507 & ~n_31508;
assign n_31510 =  x_2283 & ~n_31509;
assign n_31511 = ~x_2283 &  n_31509;
assign n_31512 = ~n_31510 & ~n_31511;
assign n_31513 = ~n_26110 & ~n_27728;
assign n_31514 = ~n_24031 &  n_31513;
assign n_31515 = ~n_26491 &  n_31514;
assign n_31516 =  x_2282 &  n_31515;
assign n_31517 =  x_651 &  n_26491;
assign n_31518 =  x_1994 &  x_2218;
assign n_31519 = ~x_1994 & ~x_2218;
assign n_31520 = ~n_31518 & ~n_31519;
assign n_31521 =  n_24031 &  n_31520;
assign n_31522 =  x_843 &  x_3735;
assign n_31523 = ~x_843 & ~x_3735;
assign n_31524 = ~n_31522 & ~n_31523;
assign n_31525 =  n_27728 &  n_31524;
assign n_31526 =  x_4104 &  x_4903;
assign n_31527 = ~x_4104 & ~x_4903;
assign n_31528 = ~n_31526 & ~n_31527;
assign n_31529 =  n_26110 &  n_31528;
assign n_31530 = ~n_31525 & ~n_31529;
assign n_31531 = ~n_31521 &  n_31530;
assign n_31532 = ~n_31517 &  n_31531;
assign n_31533 = ~n_31516 &  n_31532;
assign n_31534 =  x_2282 & ~n_31533;
assign n_31535 = ~x_2282 &  n_31533;
assign n_31536 = ~n_31534 & ~n_31535;
assign n_31537 =  x_2281 &  n_31515;
assign n_31538 =  x_650 &  n_26491;
assign n_31539 = ~x_4103 & ~x_4104;
assign n_31540 =  x_4103 &  x_4104;
assign n_31541 = ~n_31539 & ~n_31540;
assign n_31542 =  x_4902 &  n_31541;
assign n_31543 = ~x_4902 & ~n_31541;
assign n_31544 = ~n_31542 & ~n_31543;
assign n_31545 =  n_31526 &  n_31544;
assign n_31546 = ~n_31526 & ~n_31544;
assign n_31547 =  n_26110 & ~n_31546;
assign n_31548 = ~n_31545 &  n_31547;
assign n_31549 = ~x_1993 & ~x_1994;
assign n_31550 =  x_1993 &  x_1994;
assign n_31551 = ~n_31549 & ~n_31550;
assign n_31552 =  x_2217 &  n_31551;
assign n_31553 = ~x_2217 & ~n_31551;
assign n_31554 = ~n_31552 & ~n_31553;
assign n_31555 = ~n_31518 & ~n_31554;
assign n_31556 =  n_31518 &  n_31554;
assign n_31557 =  n_24031 & ~n_31556;
assign n_31558 = ~n_31555 &  n_31557;
assign n_31559 = ~x_3734 & ~x_3735;
assign n_31560 =  x_3734 &  x_3735;
assign n_31561 = ~n_31559 & ~n_31560;
assign n_31562 =  x_842 &  n_31561;
assign n_31563 = ~x_842 & ~n_31561;
assign n_31564 = ~n_31562 & ~n_31563;
assign n_31565 = ~n_31522 & ~n_31564;
assign n_31566 =  n_31522 &  n_31564;
assign n_31567 =  n_27728 & ~n_31566;
assign n_31568 = ~n_31565 &  n_31567;
assign n_31569 = ~n_31558 & ~n_31568;
assign n_31570 = ~n_31548 &  n_31569;
assign n_31571 = ~n_31538 &  n_31570;
assign n_31572 = ~n_31537 &  n_31571;
assign n_31573 =  x_2281 & ~n_31572;
assign n_31574 = ~x_2281 &  n_31572;
assign n_31575 = ~n_31573 & ~n_31574;
assign n_31576 =  x_2280 &  n_31515;
assign n_31577 =  x_649 &  n_26491;
assign n_31578 = ~x_4102 &  n_31539;
assign n_31579 =  x_4102 & ~n_31539;
assign n_31580 = ~n_31578 & ~n_31579;
assign n_31581 =  x_4103 & ~x_4902;
assign n_31582 =  n_31526 & ~n_31581;
assign n_31583 = ~n_31582 & ~n_31542;
assign n_31584 =  n_31580 & ~n_31583;
assign n_31585 = ~n_31580 &  n_31583;
assign n_31586 = ~n_31584 & ~n_31585;
assign n_31587 = ~x_4901 & ~n_31586;
assign n_31588 =  x_4901 & ~n_31585;
assign n_31589 = ~n_31584 &  n_31588;
assign n_31590 =  n_26110 & ~n_31589;
assign n_31591 = ~n_31587 &  n_31590;
assign n_31592 = ~n_31577 & ~n_31591;
assign n_31593 = ~x_3733 &  n_31559;
assign n_31594 =  x_3733 & ~n_31559;
assign n_31595 = ~n_31593 & ~n_31594;
assign n_31596 = ~x_842 &  x_3734;
assign n_31597 =  n_31522 & ~n_31596;
assign n_31598 = ~n_31597 & ~n_31562;
assign n_31599 =  n_31595 & ~n_31598;
assign n_31600 = ~n_31595 &  n_31598;
assign n_31601 = ~n_31599 & ~n_31600;
assign n_31602 = ~x_841 & ~n_31601;
assign n_31603 =  x_841 & ~n_31600;
assign n_31604 = ~n_31599 &  n_31603;
assign n_31605 =  n_27728 & ~n_31604;
assign n_31606 = ~n_31602 &  n_31605;
assign n_31607 = ~x_1992 &  n_31549;
assign n_31608 =  x_1992 & ~n_31549;
assign n_31609 = ~n_31607 & ~n_31608;
assign n_31610 =  x_1993 & ~x_2217;
assign n_31611 =  n_31518 & ~n_31610;
assign n_31612 = ~n_31611 & ~n_31552;
assign n_31613 =  n_31609 & ~n_31612;
assign n_31614 = ~n_31609 &  n_31612;
assign n_31615 = ~n_31613 & ~n_31614;
assign n_31616 = ~x_2216 & ~n_31615;
assign n_31617 =  x_2216 & ~n_31614;
assign n_31618 = ~n_31613 &  n_31617;
assign n_31619 =  n_24031 & ~n_31618;
assign n_31620 = ~n_31616 &  n_31619;
assign n_31621 = ~n_31606 & ~n_31620;
assign n_31622 =  n_31592 &  n_31621;
assign n_31623 = ~n_31576 &  n_31622;
assign n_31624 =  x_2280 & ~n_31623;
assign n_31625 = ~x_2280 &  n_31623;
assign n_31626 = ~n_31624 & ~n_31625;
assign n_31627 = ~x_1991 &  n_31607;
assign n_31628 =  x_1991 & ~n_31607;
assign n_31629 = ~n_31627 & ~n_31628;
assign n_31630 = ~n_31613 & ~n_31617;
assign n_31631 =  n_31629 & ~n_31630;
assign n_31632 = ~n_31629 &  n_31630;
assign n_31633 = ~n_31631 & ~n_31632;
assign n_31634 = ~x_2215 & ~n_31633;
assign n_31635 =  x_2215 & ~n_31632;
assign n_31636 = ~n_31631 &  n_31635;
assign n_31637 =  n_24031 & ~n_31636;
assign n_31638 = ~n_31634 &  n_31637;
assign n_31639 =  x_2279 &  n_31515;
assign n_31640 =  x_648 &  n_26491;
assign n_31641 = ~n_31639 & ~n_31640;
assign n_31642 = ~n_31638 &  n_31641;
assign n_31643 = ~x_4101 &  n_31578;
assign n_31644 =  x_4101 & ~n_31578;
assign n_31645 = ~n_31643 & ~n_31644;
assign n_31646 = ~n_31584 & ~n_31588;
assign n_31647 =  n_31645 & ~n_31646;
assign n_31648 = ~n_31645 &  n_31646;
assign n_31649 = ~n_31647 & ~n_31648;
assign n_31650 = ~x_4900 & ~n_31649;
assign n_31651 =  x_4900 & ~n_31648;
assign n_31652 = ~n_31647 &  n_31651;
assign n_31653 =  n_26110 & ~n_31652;
assign n_31654 = ~n_31650 &  n_31653;
assign n_31655 = ~x_3732 &  n_31593;
assign n_31656 =  x_3732 & ~n_31593;
assign n_31657 = ~n_31655 & ~n_31656;
assign n_31658 = ~n_31599 & ~n_31603;
assign n_31659 =  n_31657 & ~n_31658;
assign n_31660 = ~n_31657 &  n_31658;
assign n_31661 = ~n_31659 & ~n_31660;
assign n_31662 = ~x_840 & ~n_31661;
assign n_31663 =  x_840 & ~n_31660;
assign n_31664 = ~n_31659 &  n_31663;
assign n_31665 =  n_27728 & ~n_31664;
assign n_31666 = ~n_31662 &  n_31665;
assign n_31667 = ~n_31654 & ~n_31666;
assign n_31668 =  n_31642 &  n_31667;
assign n_31669 =  x_2279 & ~n_31668;
assign n_31670 = ~x_2279 &  n_31668;
assign n_31671 = ~n_31669 & ~n_31670;
assign n_31672 = ~x_1990 &  n_31627;
assign n_31673 =  x_1990 & ~n_31627;
assign n_31674 = ~n_31672 & ~n_31673;
assign n_31675 = ~n_31631 & ~n_31635;
assign n_31676 =  n_31674 & ~n_31675;
assign n_31677 = ~n_31674 &  n_31675;
assign n_31678 = ~n_31676 & ~n_31677;
assign n_31679 = ~x_2214 & ~n_31678;
assign n_31680 =  x_2214 & ~n_31677;
assign n_31681 = ~n_31676 &  n_31680;
assign n_31682 =  n_24031 & ~n_31681;
assign n_31683 = ~n_31679 &  n_31682;
assign n_31684 =  x_2278 &  n_31515;
assign n_31685 =  x_647 &  n_26491;
assign n_31686 = ~n_31684 & ~n_31685;
assign n_31687 = ~n_31683 &  n_31686;
assign n_31688 = ~x_4100 &  n_31643;
assign n_31689 =  x_4100 & ~n_31643;
assign n_31690 = ~n_31688 & ~n_31689;
assign n_31691 = ~n_31647 & ~n_31651;
assign n_31692 =  n_31690 & ~n_31691;
assign n_31693 = ~n_31690 &  n_31691;
assign n_31694 = ~n_31692 & ~n_31693;
assign n_31695 = ~x_4899 & ~n_31694;
assign n_31696 =  x_4899 & ~n_31693;
assign n_31697 = ~n_31692 &  n_31696;
assign n_31698 =  n_26110 & ~n_31697;
assign n_31699 = ~n_31695 &  n_31698;
assign n_31700 = ~x_3731 &  n_31655;
assign n_31701 =  x_3731 & ~n_31655;
assign n_31702 = ~n_31700 & ~n_31701;
assign n_31703 = ~n_31659 & ~n_31663;
assign n_31704 =  n_31702 & ~n_31703;
assign n_31705 = ~n_31702 &  n_31703;
assign n_31706 = ~n_31704 & ~n_31705;
assign n_31707 = ~x_839 & ~n_31706;
assign n_31708 =  x_839 & ~n_31705;
assign n_31709 = ~n_31704 &  n_31708;
assign n_31710 =  n_27728 & ~n_31709;
assign n_31711 = ~n_31707 &  n_31710;
assign n_31712 = ~n_31699 & ~n_31711;
assign n_31713 =  n_31687 &  n_31712;
assign n_31714 =  x_2278 & ~n_31713;
assign n_31715 = ~x_2278 &  n_31713;
assign n_31716 = ~n_31714 & ~n_31715;
assign n_31717 = ~x_1989 &  n_31672;
assign n_31718 =  x_1989 & ~n_31672;
assign n_31719 = ~n_31717 & ~n_31718;
assign n_31720 = ~n_31676 & ~n_31680;
assign n_31721 =  n_31719 & ~n_31720;
assign n_31722 = ~n_31719 &  n_31720;
assign n_31723 = ~n_31721 & ~n_31722;
assign n_31724 = ~x_2213 & ~n_31723;
assign n_31725 =  x_2213 & ~n_31722;
assign n_31726 = ~n_31721 &  n_31725;
assign n_31727 =  n_24031 & ~n_31726;
assign n_31728 = ~n_31724 &  n_31727;
assign n_31729 =  x_2277 &  n_31515;
assign n_31730 =  x_646 &  n_26491;
assign n_31731 = ~n_31729 & ~n_31730;
assign n_31732 = ~n_31728 &  n_31731;
assign n_31733 = ~x_4099 &  n_31688;
assign n_31734 =  x_4099 & ~n_31688;
assign n_31735 = ~n_31733 & ~n_31734;
assign n_31736 = ~n_31692 & ~n_31696;
assign n_31737 =  n_31735 & ~n_31736;
assign n_31738 = ~n_31735 &  n_31736;
assign n_31739 = ~n_31737 & ~n_31738;
assign n_31740 = ~x_4898 & ~n_31739;
assign n_31741 =  x_4898 & ~n_31738;
assign n_31742 = ~n_31737 &  n_31741;
assign n_31743 =  n_26110 & ~n_31742;
assign n_31744 = ~n_31740 &  n_31743;
assign n_31745 = ~x_3730 &  n_31700;
assign n_31746 =  x_3730 & ~n_31700;
assign n_31747 = ~n_31745 & ~n_31746;
assign n_31748 = ~n_31704 & ~n_31708;
assign n_31749 =  n_31747 & ~n_31748;
assign n_31750 = ~n_31747 &  n_31748;
assign n_31751 = ~n_31749 & ~n_31750;
assign n_31752 = ~x_838 & ~n_31751;
assign n_31753 =  x_838 & ~n_31750;
assign n_31754 = ~n_31749 &  n_31753;
assign n_31755 =  n_27728 & ~n_31754;
assign n_31756 = ~n_31752 &  n_31755;
assign n_31757 = ~n_31744 & ~n_31756;
assign n_31758 =  n_31732 &  n_31757;
assign n_31759 =  x_2277 & ~n_31758;
assign n_31760 = ~x_2277 &  n_31758;
assign n_31761 = ~n_31759 & ~n_31760;
assign n_31762 = ~x_1988 &  n_31717;
assign n_31763 =  x_1988 & ~n_31717;
assign n_31764 = ~n_31762 & ~n_31763;
assign n_31765 = ~n_31721 & ~n_31725;
assign n_31766 =  n_31764 & ~n_31765;
assign n_31767 = ~n_31764 &  n_31765;
assign n_31768 = ~n_31766 & ~n_31767;
assign n_31769 = ~x_2212 & ~n_31768;
assign n_31770 =  x_2212 & ~n_31767;
assign n_31771 = ~n_31766 &  n_31770;
assign n_31772 =  n_24031 & ~n_31771;
assign n_31773 = ~n_31769 &  n_31772;
assign n_31774 =  x_2276 &  n_31515;
assign n_31775 =  x_645 &  n_26491;
assign n_31776 = ~n_31774 & ~n_31775;
assign n_31777 = ~n_31773 &  n_31776;
assign n_31778 = ~x_4098 &  n_31733;
assign n_31779 =  x_4098 & ~n_31733;
assign n_31780 = ~n_31778 & ~n_31779;
assign n_31781 = ~n_31737 & ~n_31741;
assign n_31782 =  n_31780 & ~n_31781;
assign n_31783 = ~n_31780 &  n_31781;
assign n_31784 = ~n_31782 & ~n_31783;
assign n_31785 = ~x_4897 & ~n_31784;
assign n_31786 =  x_4897 & ~n_31783;
assign n_31787 = ~n_31782 &  n_31786;
assign n_31788 =  n_26110 & ~n_31787;
assign n_31789 = ~n_31785 &  n_31788;
assign n_31790 = ~x_3729 &  n_31745;
assign n_31791 =  x_3729 & ~n_31745;
assign n_31792 = ~n_31790 & ~n_31791;
assign n_31793 = ~n_31749 & ~n_31753;
assign n_31794 =  n_31792 & ~n_31793;
assign n_31795 = ~n_31792 &  n_31793;
assign n_31796 = ~n_31794 & ~n_31795;
assign n_31797 = ~x_837 & ~n_31796;
assign n_31798 =  x_837 & ~n_31795;
assign n_31799 = ~n_31794 &  n_31798;
assign n_31800 =  n_27728 & ~n_31799;
assign n_31801 = ~n_31797 &  n_31800;
assign n_31802 = ~n_31789 & ~n_31801;
assign n_31803 =  n_31777 &  n_31802;
assign n_31804 =  x_2276 & ~n_31803;
assign n_31805 = ~x_2276 &  n_31803;
assign n_31806 = ~n_31804 & ~n_31805;
assign n_31807 = ~x_1987 &  n_31762;
assign n_31808 =  x_1987 & ~n_31762;
assign n_31809 = ~n_31807 & ~n_31808;
assign n_31810 = ~n_31766 & ~n_31770;
assign n_31811 =  n_31809 & ~n_31810;
assign n_31812 = ~n_31809 &  n_31810;
assign n_31813 = ~n_31811 & ~n_31812;
assign n_31814 = ~x_2211 & ~n_31813;
assign n_31815 =  x_2211 & ~n_31812;
assign n_31816 = ~n_31811 &  n_31815;
assign n_31817 =  n_24031 & ~n_31816;
assign n_31818 = ~n_31814 &  n_31817;
assign n_31819 =  x_2275 &  n_31515;
assign n_31820 =  x_644 &  n_26491;
assign n_31821 = ~n_31819 & ~n_31820;
assign n_31822 = ~n_31818 &  n_31821;
assign n_31823 = ~x_4097 &  n_31778;
assign n_31824 =  x_4097 & ~n_31778;
assign n_31825 = ~n_31823 & ~n_31824;
assign n_31826 = ~n_31782 & ~n_31786;
assign n_31827 =  n_31825 & ~n_31826;
assign n_31828 = ~n_31825 &  n_31826;
assign n_31829 = ~n_31827 & ~n_31828;
assign n_31830 = ~x_4896 & ~n_31829;
assign n_31831 =  x_4896 & ~n_31828;
assign n_31832 = ~n_31827 &  n_31831;
assign n_31833 =  n_26110 & ~n_31832;
assign n_31834 = ~n_31830 &  n_31833;
assign n_31835 = ~x_3728 &  n_31790;
assign n_31836 =  x_3728 & ~n_31790;
assign n_31837 = ~n_31835 & ~n_31836;
assign n_31838 = ~n_31794 & ~n_31798;
assign n_31839 =  n_31837 & ~n_31838;
assign n_31840 = ~n_31837 &  n_31838;
assign n_31841 = ~n_31839 & ~n_31840;
assign n_31842 = ~x_836 & ~n_31841;
assign n_31843 =  x_836 & ~n_31840;
assign n_31844 = ~n_31839 &  n_31843;
assign n_31845 =  n_27728 & ~n_31844;
assign n_31846 = ~n_31842 &  n_31845;
assign n_31847 = ~n_31834 & ~n_31846;
assign n_31848 =  n_31822 &  n_31847;
assign n_31849 =  x_2275 & ~n_31848;
assign n_31850 = ~x_2275 &  n_31848;
assign n_31851 = ~n_31849 & ~n_31850;
assign n_31852 = ~x_1986 &  n_31807;
assign n_31853 =  x_1986 & ~n_31807;
assign n_31854 = ~n_31852 & ~n_31853;
assign n_31855 = ~n_31811 & ~n_31815;
assign n_31856 =  n_31854 & ~n_31855;
assign n_31857 = ~n_31854 &  n_31855;
assign n_31858 = ~n_31856 & ~n_31857;
assign n_31859 = ~x_2210 & ~n_31858;
assign n_31860 =  x_2210 & ~n_31857;
assign n_31861 = ~n_31856 &  n_31860;
assign n_31862 =  n_24031 & ~n_31861;
assign n_31863 = ~n_31859 &  n_31862;
assign n_31864 =  x_2274 &  n_31515;
assign n_31865 =  x_643 &  n_26491;
assign n_31866 = ~n_31864 & ~n_31865;
assign n_31867 = ~n_31863 &  n_31866;
assign n_31868 = ~x_4096 &  n_31823;
assign n_31869 =  x_4096 & ~n_31823;
assign n_31870 = ~n_31868 & ~n_31869;
assign n_31871 = ~n_31827 & ~n_31831;
assign n_31872 =  n_31870 & ~n_31871;
assign n_31873 = ~n_31870 &  n_31871;
assign n_31874 = ~n_31872 & ~n_31873;
assign n_31875 = ~x_4895 & ~n_31874;
assign n_31876 =  x_4895 & ~n_31873;
assign n_31877 = ~n_31872 &  n_31876;
assign n_31878 =  n_26110 & ~n_31877;
assign n_31879 = ~n_31875 &  n_31878;
assign n_31880 = ~x_3727 &  n_31835;
assign n_31881 =  x_3727 & ~n_31835;
assign n_31882 = ~n_31880 & ~n_31881;
assign n_31883 = ~n_31839 & ~n_31843;
assign n_31884 =  n_31882 & ~n_31883;
assign n_31885 = ~n_31882 &  n_31883;
assign n_31886 = ~n_31884 & ~n_31885;
assign n_31887 = ~x_835 & ~n_31886;
assign n_31888 =  x_835 & ~n_31885;
assign n_31889 = ~n_31884 &  n_31888;
assign n_31890 =  n_27728 & ~n_31889;
assign n_31891 = ~n_31887 &  n_31890;
assign n_31892 = ~n_31879 & ~n_31891;
assign n_31893 =  n_31867 &  n_31892;
assign n_31894 =  x_2274 & ~n_31893;
assign n_31895 = ~x_2274 &  n_31893;
assign n_31896 = ~n_31894 & ~n_31895;
assign n_31897 = ~x_1985 &  n_31852;
assign n_31898 =  x_1985 & ~n_31852;
assign n_31899 = ~n_31897 & ~n_31898;
assign n_31900 = ~n_31856 & ~n_31860;
assign n_31901 =  n_31899 & ~n_31900;
assign n_31902 = ~n_31899 &  n_31900;
assign n_31903 = ~n_31901 & ~n_31902;
assign n_31904 = ~x_2209 & ~n_31903;
assign n_31905 =  x_2209 & ~n_31902;
assign n_31906 = ~n_31901 &  n_31905;
assign n_31907 =  n_24031 & ~n_31906;
assign n_31908 = ~n_31904 &  n_31907;
assign n_31909 =  x_2273 &  n_31515;
assign n_31910 =  x_642 &  n_26491;
assign n_31911 = ~n_31909 & ~n_31910;
assign n_31912 = ~n_31908 &  n_31911;
assign n_31913 = ~x_4095 &  n_31868;
assign n_31914 =  x_4095 & ~n_31868;
assign n_31915 = ~n_31913 & ~n_31914;
assign n_31916 = ~n_31872 & ~n_31876;
assign n_31917 =  n_31915 & ~n_31916;
assign n_31918 = ~n_31915 &  n_31916;
assign n_31919 = ~n_31917 & ~n_31918;
assign n_31920 = ~x_4894 & ~n_31919;
assign n_31921 =  x_4894 & ~n_31918;
assign n_31922 = ~n_31917 &  n_31921;
assign n_31923 =  n_26110 & ~n_31922;
assign n_31924 = ~n_31920 &  n_31923;
assign n_31925 = ~x_3726 &  n_31880;
assign n_31926 =  x_3726 & ~n_31880;
assign n_31927 = ~n_31925 & ~n_31926;
assign n_31928 = ~n_31884 & ~n_31888;
assign n_31929 =  n_31927 & ~n_31928;
assign n_31930 = ~n_31927 &  n_31928;
assign n_31931 = ~n_31929 & ~n_31930;
assign n_31932 = ~x_834 & ~n_31931;
assign n_31933 =  x_834 & ~n_31930;
assign n_31934 = ~n_31929 &  n_31933;
assign n_31935 =  n_27728 & ~n_31934;
assign n_31936 = ~n_31932 &  n_31935;
assign n_31937 = ~n_31924 & ~n_31936;
assign n_31938 =  n_31912 &  n_31937;
assign n_31939 =  x_2273 & ~n_31938;
assign n_31940 = ~x_2273 &  n_31938;
assign n_31941 = ~n_31939 & ~n_31940;
assign n_31942 = ~x_1984 &  n_31897;
assign n_31943 =  x_1984 & ~n_31897;
assign n_31944 = ~n_31942 & ~n_31943;
assign n_31945 = ~n_31901 & ~n_31905;
assign n_31946 =  n_31944 & ~n_31945;
assign n_31947 = ~n_31944 &  n_31945;
assign n_31948 = ~n_31946 & ~n_31947;
assign n_31949 = ~x_2208 & ~n_31948;
assign n_31950 =  x_2208 & ~n_31947;
assign n_31951 = ~n_31946 &  n_31950;
assign n_31952 =  n_24031 & ~n_31951;
assign n_31953 = ~n_31949 &  n_31952;
assign n_31954 =  x_2272 &  n_31515;
assign n_31955 =  x_641 &  n_26491;
assign n_31956 = ~n_31954 & ~n_31955;
assign n_31957 = ~n_31953 &  n_31956;
assign n_31958 = ~x_4094 &  n_31913;
assign n_31959 =  x_4094 & ~n_31913;
assign n_31960 = ~n_31958 & ~n_31959;
assign n_31961 = ~n_31917 & ~n_31921;
assign n_31962 =  n_31960 & ~n_31961;
assign n_31963 = ~n_31960 &  n_31961;
assign n_31964 = ~n_31962 & ~n_31963;
assign n_31965 = ~x_4893 & ~n_31964;
assign n_31966 =  x_4893 & ~n_31963;
assign n_31967 = ~n_31962 &  n_31966;
assign n_31968 =  n_26110 & ~n_31967;
assign n_31969 = ~n_31965 &  n_31968;
assign n_31970 = ~x_3725 &  n_31925;
assign n_31971 =  x_3725 & ~n_31925;
assign n_31972 = ~n_31970 & ~n_31971;
assign n_31973 = ~n_31929 & ~n_31933;
assign n_31974 =  n_31972 & ~n_31973;
assign n_31975 = ~n_31972 &  n_31973;
assign n_31976 = ~n_31974 & ~n_31975;
assign n_31977 = ~x_833 & ~n_31976;
assign n_31978 =  x_833 & ~n_31975;
assign n_31979 = ~n_31974 &  n_31978;
assign n_31980 =  n_27728 & ~n_31979;
assign n_31981 = ~n_31977 &  n_31980;
assign n_31982 = ~n_31969 & ~n_31981;
assign n_31983 =  n_31957 &  n_31982;
assign n_31984 =  x_2272 & ~n_31983;
assign n_31985 = ~x_2272 &  n_31983;
assign n_31986 = ~n_31984 & ~n_31985;
assign n_31987 = ~x_1983 &  n_31942;
assign n_31988 =  x_1983 & ~n_31942;
assign n_31989 = ~n_31987 & ~n_31988;
assign n_31990 = ~n_31946 & ~n_31950;
assign n_31991 =  n_31989 & ~n_31990;
assign n_31992 = ~n_31989 &  n_31990;
assign n_31993 = ~n_31991 & ~n_31992;
assign n_31994 = ~x_2207 & ~n_31993;
assign n_31995 =  x_2207 & ~n_31992;
assign n_31996 = ~n_31991 &  n_31995;
assign n_31997 =  n_24031 & ~n_31996;
assign n_31998 = ~n_31994 &  n_31997;
assign n_31999 =  x_2271 &  n_31515;
assign n_32000 =  x_640 &  n_26491;
assign n_32001 = ~n_31999 & ~n_32000;
assign n_32002 = ~n_31998 &  n_32001;
assign n_32003 = ~x_4093 &  n_31958;
assign n_32004 =  x_4093 & ~n_31958;
assign n_32005 = ~n_32003 & ~n_32004;
assign n_32006 = ~n_31962 & ~n_31966;
assign n_32007 =  n_32005 & ~n_32006;
assign n_32008 = ~n_32005 &  n_32006;
assign n_32009 = ~n_32007 & ~n_32008;
assign n_32010 = ~x_4892 & ~n_32009;
assign n_32011 =  x_4892 & ~n_32008;
assign n_32012 = ~n_32007 &  n_32011;
assign n_32013 =  n_26110 & ~n_32012;
assign n_32014 = ~n_32010 &  n_32013;
assign n_32015 = ~x_3724 &  n_31970;
assign n_32016 =  x_3724 & ~n_31970;
assign n_32017 = ~n_32015 & ~n_32016;
assign n_32018 = ~n_31974 & ~n_31978;
assign n_32019 =  n_32017 & ~n_32018;
assign n_32020 = ~n_32017 &  n_32018;
assign n_32021 = ~n_32019 & ~n_32020;
assign n_32022 = ~x_832 & ~n_32021;
assign n_32023 =  x_832 & ~n_32020;
assign n_32024 = ~n_32019 &  n_32023;
assign n_32025 =  n_27728 & ~n_32024;
assign n_32026 = ~n_32022 &  n_32025;
assign n_32027 = ~n_32014 & ~n_32026;
assign n_32028 =  n_32002 &  n_32027;
assign n_32029 =  x_2271 & ~n_32028;
assign n_32030 = ~x_2271 &  n_32028;
assign n_32031 = ~n_32029 & ~n_32030;
assign n_32032 = ~x_1982 &  n_31987;
assign n_32033 =  x_1982 & ~n_31987;
assign n_32034 = ~n_32032 & ~n_32033;
assign n_32035 = ~n_31991 & ~n_31995;
assign n_32036 =  n_32034 & ~n_32035;
assign n_32037 = ~n_32034 &  n_32035;
assign n_32038 = ~n_32036 & ~n_32037;
assign n_32039 = ~x_2206 & ~n_32038;
assign n_32040 =  x_2206 & ~n_32037;
assign n_32041 = ~n_32036 &  n_32040;
assign n_32042 =  n_24031 & ~n_32041;
assign n_32043 = ~n_32039 &  n_32042;
assign n_32044 =  x_2270 &  n_31515;
assign n_32045 =  x_639 &  n_26491;
assign n_32046 = ~n_32044 & ~n_32045;
assign n_32047 = ~n_32043 &  n_32046;
assign n_32048 = ~x_4092 &  n_32003;
assign n_32049 =  x_4092 & ~n_32003;
assign n_32050 = ~n_32048 & ~n_32049;
assign n_32051 = ~n_32007 & ~n_32011;
assign n_32052 =  n_32050 & ~n_32051;
assign n_32053 = ~n_32050 &  n_32051;
assign n_32054 = ~n_32052 & ~n_32053;
assign n_32055 = ~x_4891 & ~n_32054;
assign n_32056 =  x_4891 & ~n_32053;
assign n_32057 = ~n_32052 &  n_32056;
assign n_32058 =  n_26110 & ~n_32057;
assign n_32059 = ~n_32055 &  n_32058;
assign n_32060 = ~x_3723 &  n_32015;
assign n_32061 =  x_3723 & ~n_32015;
assign n_32062 = ~n_32060 & ~n_32061;
assign n_32063 = ~n_32019 & ~n_32023;
assign n_32064 =  n_32062 & ~n_32063;
assign n_32065 = ~n_32062 &  n_32063;
assign n_32066 = ~n_32064 & ~n_32065;
assign n_32067 = ~x_831 & ~n_32066;
assign n_32068 =  x_831 & ~n_32065;
assign n_32069 = ~n_32064 &  n_32068;
assign n_32070 =  n_27728 & ~n_32069;
assign n_32071 = ~n_32067 &  n_32070;
assign n_32072 = ~n_32059 & ~n_32071;
assign n_32073 =  n_32047 &  n_32072;
assign n_32074 =  x_2270 & ~n_32073;
assign n_32075 = ~x_2270 &  n_32073;
assign n_32076 = ~n_32074 & ~n_32075;
assign n_32077 = ~x_1981 &  n_32032;
assign n_32078 =  x_1981 & ~n_32032;
assign n_32079 = ~n_32077 & ~n_32078;
assign n_32080 = ~n_32036 & ~n_32040;
assign n_32081 =  n_32079 & ~n_32080;
assign n_32082 = ~n_32079 &  n_32080;
assign n_32083 = ~n_32081 & ~n_32082;
assign n_32084 = ~x_2205 & ~n_32083;
assign n_32085 =  x_2205 & ~n_32082;
assign n_32086 = ~n_32081 &  n_32085;
assign n_32087 =  n_24031 & ~n_32086;
assign n_32088 = ~n_32084 &  n_32087;
assign n_32089 =  x_2269 &  n_31515;
assign n_32090 =  x_638 &  n_26491;
assign n_32091 = ~n_32089 & ~n_32090;
assign n_32092 = ~n_32088 &  n_32091;
assign n_32093 = ~x_4091 &  n_32048;
assign n_32094 =  x_4091 & ~n_32048;
assign n_32095 = ~n_32093 & ~n_32094;
assign n_32096 = ~n_32052 & ~n_32056;
assign n_32097 =  n_32095 & ~n_32096;
assign n_32098 = ~n_32095 &  n_32096;
assign n_32099 = ~n_32097 & ~n_32098;
assign n_32100 = ~x_4890 & ~n_32099;
assign n_32101 =  x_4890 & ~n_32098;
assign n_32102 = ~n_32097 &  n_32101;
assign n_32103 =  n_26110 & ~n_32102;
assign n_32104 = ~n_32100 &  n_32103;
assign n_32105 = ~x_3722 &  n_32060;
assign n_32106 =  x_3722 & ~n_32060;
assign n_32107 = ~n_32105 & ~n_32106;
assign n_32108 = ~n_32064 & ~n_32068;
assign n_32109 =  n_32107 & ~n_32108;
assign n_32110 = ~n_32107 &  n_32108;
assign n_32111 = ~n_32109 & ~n_32110;
assign n_32112 = ~x_830 & ~n_32111;
assign n_32113 =  x_830 & ~n_32110;
assign n_32114 = ~n_32109 &  n_32113;
assign n_32115 =  n_27728 & ~n_32114;
assign n_32116 = ~n_32112 &  n_32115;
assign n_32117 = ~n_32104 & ~n_32116;
assign n_32118 =  n_32092 &  n_32117;
assign n_32119 =  x_2269 & ~n_32118;
assign n_32120 = ~x_2269 &  n_32118;
assign n_32121 = ~n_32119 & ~n_32120;
assign n_32122 = ~x_1980 &  n_32077;
assign n_32123 =  x_1980 & ~n_32077;
assign n_32124 = ~n_32122 & ~n_32123;
assign n_32125 = ~n_32081 & ~n_32085;
assign n_32126 =  n_32124 & ~n_32125;
assign n_32127 = ~n_32124 &  n_32125;
assign n_32128 = ~n_32126 & ~n_32127;
assign n_32129 = ~x_2204 & ~n_32128;
assign n_32130 =  x_2204 & ~n_32127;
assign n_32131 = ~n_32126 &  n_32130;
assign n_32132 =  n_24031 & ~n_32131;
assign n_32133 = ~n_32129 &  n_32132;
assign n_32134 =  x_2268 &  n_31515;
assign n_32135 =  x_637 &  n_26491;
assign n_32136 = ~n_32134 & ~n_32135;
assign n_32137 = ~n_32133 &  n_32136;
assign n_32138 = ~x_4090 &  n_32093;
assign n_32139 =  x_4090 & ~n_32093;
assign n_32140 = ~n_32138 & ~n_32139;
assign n_32141 = ~n_32097 & ~n_32101;
assign n_32142 =  n_32140 & ~n_32141;
assign n_32143 = ~n_32140 &  n_32141;
assign n_32144 = ~n_32142 & ~n_32143;
assign n_32145 = ~x_4889 & ~n_32144;
assign n_32146 =  x_4889 & ~n_32143;
assign n_32147 = ~n_32142 &  n_32146;
assign n_32148 =  n_26110 & ~n_32147;
assign n_32149 = ~n_32145 &  n_32148;
assign n_32150 = ~x_3721 &  n_32105;
assign n_32151 =  x_3721 & ~n_32105;
assign n_32152 = ~n_32150 & ~n_32151;
assign n_32153 = ~n_32109 & ~n_32113;
assign n_32154 =  n_32152 & ~n_32153;
assign n_32155 = ~n_32152 &  n_32153;
assign n_32156 = ~n_32154 & ~n_32155;
assign n_32157 = ~x_829 & ~n_32156;
assign n_32158 =  x_829 & ~n_32155;
assign n_32159 = ~n_32154 &  n_32158;
assign n_32160 =  n_27728 & ~n_32159;
assign n_32161 = ~n_32157 &  n_32160;
assign n_32162 = ~n_32149 & ~n_32161;
assign n_32163 =  n_32137 &  n_32162;
assign n_32164 =  x_2268 & ~n_32163;
assign n_32165 = ~x_2268 &  n_32163;
assign n_32166 = ~n_32164 & ~n_32165;
assign n_32167 = ~x_1979 &  n_32122;
assign n_32168 =  x_1979 & ~n_32122;
assign n_32169 = ~n_32167 & ~n_32168;
assign n_32170 = ~n_32126 & ~n_32130;
assign n_32171 =  n_32169 & ~n_32170;
assign n_32172 = ~n_32169 &  n_32170;
assign n_32173 = ~n_32171 & ~n_32172;
assign n_32174 = ~x_2203 & ~n_32173;
assign n_32175 =  x_2203 & ~n_32172;
assign n_32176 = ~n_32171 &  n_32175;
assign n_32177 =  n_24031 & ~n_32176;
assign n_32178 = ~n_32174 &  n_32177;
assign n_32179 =  x_2267 &  n_31515;
assign n_32180 =  x_636 &  n_26491;
assign n_32181 = ~n_32179 & ~n_32180;
assign n_32182 = ~n_32178 &  n_32181;
assign n_32183 = ~x_4089 &  n_32138;
assign n_32184 =  x_4089 & ~n_32138;
assign n_32185 = ~n_32183 & ~n_32184;
assign n_32186 = ~n_32142 & ~n_32146;
assign n_32187 =  n_32185 & ~n_32186;
assign n_32188 = ~n_32185 &  n_32186;
assign n_32189 = ~n_32187 & ~n_32188;
assign n_32190 = ~x_4888 & ~n_32189;
assign n_32191 =  x_4888 & ~n_32188;
assign n_32192 = ~n_32187 &  n_32191;
assign n_32193 =  n_26110 & ~n_32192;
assign n_32194 = ~n_32190 &  n_32193;
assign n_32195 = ~x_3720 &  n_32150;
assign n_32196 =  x_3720 & ~n_32150;
assign n_32197 = ~n_32195 & ~n_32196;
assign n_32198 = ~n_32154 & ~n_32158;
assign n_32199 =  n_32197 & ~n_32198;
assign n_32200 = ~n_32197 &  n_32198;
assign n_32201 = ~n_32199 & ~n_32200;
assign n_32202 = ~x_828 & ~n_32201;
assign n_32203 =  x_828 & ~n_32200;
assign n_32204 = ~n_32199 &  n_32203;
assign n_32205 =  n_27728 & ~n_32204;
assign n_32206 = ~n_32202 &  n_32205;
assign n_32207 = ~n_32194 & ~n_32206;
assign n_32208 =  n_32182 &  n_32207;
assign n_32209 =  x_2267 & ~n_32208;
assign n_32210 = ~x_2267 &  n_32208;
assign n_32211 = ~n_32209 & ~n_32210;
assign n_32212 = ~x_1978 &  n_32167;
assign n_32213 =  x_1978 & ~n_32167;
assign n_32214 = ~n_32212 & ~n_32213;
assign n_32215 = ~n_32171 & ~n_32175;
assign n_32216 =  n_32214 & ~n_32215;
assign n_32217 = ~n_32214 &  n_32215;
assign n_32218 = ~n_32216 & ~n_32217;
assign n_32219 = ~x_2202 & ~n_32218;
assign n_32220 =  x_2202 & ~n_32217;
assign n_32221 = ~n_32216 &  n_32220;
assign n_32222 =  n_24031 & ~n_32221;
assign n_32223 = ~n_32219 &  n_32222;
assign n_32224 =  x_2266 &  n_31515;
assign n_32225 =  x_635 &  n_26491;
assign n_32226 = ~n_32224 & ~n_32225;
assign n_32227 = ~n_32223 &  n_32226;
assign n_32228 = ~x_4088 &  n_32183;
assign n_32229 =  x_4088 & ~n_32183;
assign n_32230 = ~n_32228 & ~n_32229;
assign n_32231 = ~n_32187 & ~n_32191;
assign n_32232 =  n_32230 & ~n_32231;
assign n_32233 = ~n_32230 &  n_32231;
assign n_32234 = ~n_32232 & ~n_32233;
assign n_32235 = ~x_4887 & ~n_32234;
assign n_32236 =  x_4887 & ~n_32233;
assign n_32237 = ~n_32232 &  n_32236;
assign n_32238 =  n_26110 & ~n_32237;
assign n_32239 = ~n_32235 &  n_32238;
assign n_32240 = ~x_3719 &  n_32195;
assign n_32241 =  x_3719 & ~n_32195;
assign n_32242 = ~n_32240 & ~n_32241;
assign n_32243 = ~n_32199 & ~n_32203;
assign n_32244 =  n_32242 & ~n_32243;
assign n_32245 = ~n_32242 &  n_32243;
assign n_32246 = ~n_32244 & ~n_32245;
assign n_32247 = ~x_827 & ~n_32246;
assign n_32248 =  x_827 & ~n_32245;
assign n_32249 = ~n_32244 &  n_32248;
assign n_32250 =  n_27728 & ~n_32249;
assign n_32251 = ~n_32247 &  n_32250;
assign n_32252 = ~n_32239 & ~n_32251;
assign n_32253 =  n_32227 &  n_32252;
assign n_32254 =  x_2266 & ~n_32253;
assign n_32255 = ~x_2266 &  n_32253;
assign n_32256 = ~n_32254 & ~n_32255;
assign n_32257 = ~x_1977 &  n_32212;
assign n_32258 =  x_1977 & ~n_32212;
assign n_32259 = ~n_32257 & ~n_32258;
assign n_32260 = ~n_32216 & ~n_32220;
assign n_32261 =  n_32259 & ~n_32260;
assign n_32262 = ~n_32259 &  n_32260;
assign n_32263 = ~n_32261 & ~n_32262;
assign n_32264 = ~x_2201 & ~n_32263;
assign n_32265 =  x_2201 & ~n_32262;
assign n_32266 = ~n_32261 &  n_32265;
assign n_32267 =  n_24031 & ~n_32266;
assign n_32268 = ~n_32264 &  n_32267;
assign n_32269 =  x_2265 &  n_31515;
assign n_32270 =  x_634 &  n_26491;
assign n_32271 = ~n_32269 & ~n_32270;
assign n_32272 = ~n_32268 &  n_32271;
assign n_32273 = ~x_4087 &  n_32228;
assign n_32274 =  x_4087 & ~n_32228;
assign n_32275 = ~n_32273 & ~n_32274;
assign n_32276 = ~n_32232 & ~n_32236;
assign n_32277 =  n_32275 & ~n_32276;
assign n_32278 = ~n_32275 &  n_32276;
assign n_32279 = ~n_32277 & ~n_32278;
assign n_32280 = ~x_4886 & ~n_32279;
assign n_32281 =  x_4886 & ~n_32278;
assign n_32282 = ~n_32277 &  n_32281;
assign n_32283 =  n_26110 & ~n_32282;
assign n_32284 = ~n_32280 &  n_32283;
assign n_32285 = ~x_3718 &  n_32240;
assign n_32286 =  x_3718 & ~n_32240;
assign n_32287 = ~n_32285 & ~n_32286;
assign n_32288 = ~n_32244 & ~n_32248;
assign n_32289 =  n_32287 & ~n_32288;
assign n_32290 = ~n_32287 &  n_32288;
assign n_32291 = ~n_32289 & ~n_32290;
assign n_32292 = ~x_826 & ~n_32291;
assign n_32293 =  x_826 & ~n_32290;
assign n_32294 = ~n_32289 &  n_32293;
assign n_32295 =  n_27728 & ~n_32294;
assign n_32296 = ~n_32292 &  n_32295;
assign n_32297 = ~n_32284 & ~n_32296;
assign n_32298 =  n_32272 &  n_32297;
assign n_32299 =  x_2265 & ~n_32298;
assign n_32300 = ~x_2265 &  n_32298;
assign n_32301 = ~n_32299 & ~n_32300;
assign n_32302 = ~x_1976 &  n_32257;
assign n_32303 =  x_1976 & ~n_32257;
assign n_32304 = ~n_32302 & ~n_32303;
assign n_32305 = ~n_32261 & ~n_32265;
assign n_32306 =  n_32304 & ~n_32305;
assign n_32307 = ~n_32304 &  n_32305;
assign n_32308 = ~n_32306 & ~n_32307;
assign n_32309 = ~x_2200 & ~n_32308;
assign n_32310 =  x_2200 & ~n_32307;
assign n_32311 = ~n_32306 &  n_32310;
assign n_32312 =  n_24031 & ~n_32311;
assign n_32313 = ~n_32309 &  n_32312;
assign n_32314 =  x_2264 &  n_31515;
assign n_32315 =  x_633 &  n_26491;
assign n_32316 = ~n_32314 & ~n_32315;
assign n_32317 = ~n_32313 &  n_32316;
assign n_32318 = ~x_4086 &  n_32273;
assign n_32319 =  x_4086 & ~n_32273;
assign n_32320 = ~n_32318 & ~n_32319;
assign n_32321 = ~n_32277 & ~n_32281;
assign n_32322 =  n_32320 & ~n_32321;
assign n_32323 = ~n_32320 &  n_32321;
assign n_32324 = ~n_32322 & ~n_32323;
assign n_32325 = ~x_4885 & ~n_32324;
assign n_32326 =  x_4885 & ~n_32323;
assign n_32327 = ~n_32322 &  n_32326;
assign n_32328 =  n_26110 & ~n_32327;
assign n_32329 = ~n_32325 &  n_32328;
assign n_32330 = ~x_3717 &  n_32285;
assign n_32331 =  x_3717 & ~n_32285;
assign n_32332 = ~n_32330 & ~n_32331;
assign n_32333 = ~n_32289 & ~n_32293;
assign n_32334 =  n_32332 & ~n_32333;
assign n_32335 = ~n_32332 &  n_32333;
assign n_32336 = ~n_32334 & ~n_32335;
assign n_32337 = ~x_825 & ~n_32336;
assign n_32338 =  x_825 & ~n_32335;
assign n_32339 = ~n_32334 &  n_32338;
assign n_32340 =  n_27728 & ~n_32339;
assign n_32341 = ~n_32337 &  n_32340;
assign n_32342 = ~n_32329 & ~n_32341;
assign n_32343 =  n_32317 &  n_32342;
assign n_32344 =  x_2264 & ~n_32343;
assign n_32345 = ~x_2264 &  n_32343;
assign n_32346 = ~n_32344 & ~n_32345;
assign n_32347 = ~x_1975 &  n_32302;
assign n_32348 =  x_1975 & ~n_32302;
assign n_32349 = ~n_32347 & ~n_32348;
assign n_32350 = ~n_32306 & ~n_32310;
assign n_32351 =  n_32349 & ~n_32350;
assign n_32352 = ~n_32349 &  n_32350;
assign n_32353 = ~n_32351 & ~n_32352;
assign n_32354 = ~x_2199 & ~n_32353;
assign n_32355 =  x_2199 & ~n_32352;
assign n_32356 = ~n_32351 &  n_32355;
assign n_32357 =  n_24031 & ~n_32356;
assign n_32358 = ~n_32354 &  n_32357;
assign n_32359 =  x_2263 &  n_31515;
assign n_32360 =  x_632 &  n_26491;
assign n_32361 = ~n_32359 & ~n_32360;
assign n_32362 = ~n_32358 &  n_32361;
assign n_32363 = ~x_4085 &  n_32318;
assign n_32364 =  x_4085 & ~n_32318;
assign n_32365 = ~n_32363 & ~n_32364;
assign n_32366 = ~n_32322 & ~n_32326;
assign n_32367 =  n_32365 & ~n_32366;
assign n_32368 = ~n_32365 &  n_32366;
assign n_32369 = ~n_32367 & ~n_32368;
assign n_32370 = ~x_4884 & ~n_32369;
assign n_32371 =  x_4884 & ~n_32368;
assign n_32372 = ~n_32367 &  n_32371;
assign n_32373 =  n_26110 & ~n_32372;
assign n_32374 = ~n_32370 &  n_32373;
assign n_32375 = ~x_3716 &  n_32330;
assign n_32376 =  x_3716 & ~n_32330;
assign n_32377 = ~n_32375 & ~n_32376;
assign n_32378 = ~n_32334 & ~n_32338;
assign n_32379 =  n_32377 & ~n_32378;
assign n_32380 = ~n_32377 &  n_32378;
assign n_32381 = ~n_32379 & ~n_32380;
assign n_32382 = ~x_824 & ~n_32381;
assign n_32383 =  x_824 & ~n_32380;
assign n_32384 = ~n_32379 &  n_32383;
assign n_32385 =  n_27728 & ~n_32384;
assign n_32386 = ~n_32382 &  n_32385;
assign n_32387 = ~n_32374 & ~n_32386;
assign n_32388 =  n_32362 &  n_32387;
assign n_32389 =  x_2263 & ~n_32388;
assign n_32390 = ~x_2263 &  n_32388;
assign n_32391 = ~n_32389 & ~n_32390;
assign n_32392 = ~x_1974 &  n_32347;
assign n_32393 =  x_1974 & ~n_32347;
assign n_32394 = ~n_32392 & ~n_32393;
assign n_32395 = ~n_32351 & ~n_32355;
assign n_32396 =  n_32394 & ~n_32395;
assign n_32397 = ~n_32394 &  n_32395;
assign n_32398 = ~n_32396 & ~n_32397;
assign n_32399 = ~x_2198 & ~n_32398;
assign n_32400 =  x_2198 & ~n_32397;
assign n_32401 = ~n_32396 &  n_32400;
assign n_32402 =  n_24031 & ~n_32401;
assign n_32403 = ~n_32399 &  n_32402;
assign n_32404 =  x_2262 &  n_31515;
assign n_32405 =  x_631 &  n_26491;
assign n_32406 = ~n_32404 & ~n_32405;
assign n_32407 = ~n_32403 &  n_32406;
assign n_32408 = ~x_4084 &  n_32363;
assign n_32409 =  x_4084 & ~n_32363;
assign n_32410 = ~n_32408 & ~n_32409;
assign n_32411 = ~n_32367 & ~n_32371;
assign n_32412 =  n_32410 & ~n_32411;
assign n_32413 = ~n_32410 &  n_32411;
assign n_32414 = ~n_32412 & ~n_32413;
assign n_32415 = ~x_4883 & ~n_32414;
assign n_32416 =  x_4883 & ~n_32413;
assign n_32417 = ~n_32412 &  n_32416;
assign n_32418 =  n_26110 & ~n_32417;
assign n_32419 = ~n_32415 &  n_32418;
assign n_32420 = ~x_3715 &  n_32375;
assign n_32421 =  x_3715 & ~n_32375;
assign n_32422 = ~n_32420 & ~n_32421;
assign n_32423 = ~n_32379 & ~n_32383;
assign n_32424 =  n_32422 & ~n_32423;
assign n_32425 = ~n_32422 &  n_32423;
assign n_32426 = ~n_32424 & ~n_32425;
assign n_32427 = ~x_823 & ~n_32426;
assign n_32428 =  x_823 & ~n_32425;
assign n_32429 = ~n_32424 &  n_32428;
assign n_32430 =  n_27728 & ~n_32429;
assign n_32431 = ~n_32427 &  n_32430;
assign n_32432 = ~n_32419 & ~n_32431;
assign n_32433 =  n_32407 &  n_32432;
assign n_32434 =  x_2262 & ~n_32433;
assign n_32435 = ~x_2262 &  n_32433;
assign n_32436 = ~n_32434 & ~n_32435;
assign n_32437 = ~x_1973 &  n_32392;
assign n_32438 =  x_1973 & ~n_32392;
assign n_32439 = ~n_32437 & ~n_32438;
assign n_32440 = ~n_32396 & ~n_32400;
assign n_32441 =  n_32439 & ~n_32440;
assign n_32442 = ~n_32439 &  n_32440;
assign n_32443 = ~n_32441 & ~n_32442;
assign n_32444 = ~x_2197 & ~n_32443;
assign n_32445 =  x_2197 & ~n_32442;
assign n_32446 = ~n_32441 &  n_32445;
assign n_32447 =  n_24031 & ~n_32446;
assign n_32448 = ~n_32444 &  n_32447;
assign n_32449 =  x_2261 &  n_31515;
assign n_32450 =  x_630 &  n_26491;
assign n_32451 = ~n_32449 & ~n_32450;
assign n_32452 = ~n_32448 &  n_32451;
assign n_32453 = ~x_4083 &  n_32408;
assign n_32454 =  x_4083 & ~n_32408;
assign n_32455 = ~n_32453 & ~n_32454;
assign n_32456 = ~n_32412 & ~n_32416;
assign n_32457 =  n_32455 & ~n_32456;
assign n_32458 = ~n_32455 &  n_32456;
assign n_32459 = ~n_32457 & ~n_32458;
assign n_32460 = ~x_4882 & ~n_32459;
assign n_32461 =  x_4882 & ~n_32458;
assign n_32462 = ~n_32457 &  n_32461;
assign n_32463 =  n_26110 & ~n_32462;
assign n_32464 = ~n_32460 &  n_32463;
assign n_32465 = ~x_3714 &  n_32420;
assign n_32466 =  x_3714 & ~n_32420;
assign n_32467 = ~n_32465 & ~n_32466;
assign n_32468 = ~n_32424 & ~n_32428;
assign n_32469 =  n_32467 & ~n_32468;
assign n_32470 = ~n_32467 &  n_32468;
assign n_32471 = ~n_32469 & ~n_32470;
assign n_32472 = ~x_822 & ~n_32471;
assign n_32473 =  x_822 & ~n_32470;
assign n_32474 = ~n_32469 &  n_32473;
assign n_32475 =  n_27728 & ~n_32474;
assign n_32476 = ~n_32472 &  n_32475;
assign n_32477 = ~n_32464 & ~n_32476;
assign n_32478 =  n_32452 &  n_32477;
assign n_32479 =  x_2261 & ~n_32478;
assign n_32480 = ~x_2261 &  n_32478;
assign n_32481 = ~n_32479 & ~n_32480;
assign n_32482 = ~x_1972 &  n_32437;
assign n_32483 =  x_1972 & ~n_32437;
assign n_32484 = ~n_32482 & ~n_32483;
assign n_32485 = ~n_32441 & ~n_32445;
assign n_32486 =  n_32484 & ~n_32485;
assign n_32487 = ~n_32484 &  n_32485;
assign n_32488 = ~n_32486 & ~n_32487;
assign n_32489 = ~x_2196 & ~n_32488;
assign n_32490 =  x_2196 & ~n_32487;
assign n_32491 = ~n_32486 &  n_32490;
assign n_32492 =  n_24031 & ~n_32491;
assign n_32493 = ~n_32489 &  n_32492;
assign n_32494 =  x_2260 &  n_31515;
assign n_32495 =  x_629 &  n_26491;
assign n_32496 = ~n_32494 & ~n_32495;
assign n_32497 = ~n_32493 &  n_32496;
assign n_32498 = ~x_4082 &  n_32453;
assign n_32499 =  x_4082 & ~n_32453;
assign n_32500 = ~n_32498 & ~n_32499;
assign n_32501 = ~n_32457 & ~n_32461;
assign n_32502 =  n_32500 & ~n_32501;
assign n_32503 = ~n_32500 &  n_32501;
assign n_32504 = ~n_32502 & ~n_32503;
assign n_32505 = ~x_4881 & ~n_32504;
assign n_32506 =  x_4881 & ~n_32503;
assign n_32507 = ~n_32502 &  n_32506;
assign n_32508 =  n_26110 & ~n_32507;
assign n_32509 = ~n_32505 &  n_32508;
assign n_32510 = ~x_3713 &  n_32465;
assign n_32511 =  x_3713 & ~n_32465;
assign n_32512 = ~n_32510 & ~n_32511;
assign n_32513 = ~n_32469 & ~n_32473;
assign n_32514 =  n_32512 & ~n_32513;
assign n_32515 = ~n_32512 &  n_32513;
assign n_32516 = ~n_32514 & ~n_32515;
assign n_32517 = ~x_821 & ~n_32516;
assign n_32518 =  x_821 & ~n_32515;
assign n_32519 = ~n_32514 &  n_32518;
assign n_32520 =  n_27728 & ~n_32519;
assign n_32521 = ~n_32517 &  n_32520;
assign n_32522 = ~n_32509 & ~n_32521;
assign n_32523 =  n_32497 &  n_32522;
assign n_32524 =  x_2260 & ~n_32523;
assign n_32525 = ~x_2260 &  n_32523;
assign n_32526 = ~n_32524 & ~n_32525;
assign n_32527 = ~x_1971 &  n_32482;
assign n_32528 =  x_1971 & ~n_32482;
assign n_32529 = ~n_32527 & ~n_32528;
assign n_32530 = ~n_32486 & ~n_32490;
assign n_32531 =  n_32529 & ~n_32530;
assign n_32532 = ~n_32529 &  n_32530;
assign n_32533 = ~n_32531 & ~n_32532;
assign n_32534 = ~x_2195 & ~n_32533;
assign n_32535 =  x_2195 & ~n_32532;
assign n_32536 = ~n_32531 &  n_32535;
assign n_32537 =  n_24031 & ~n_32536;
assign n_32538 = ~n_32534 &  n_32537;
assign n_32539 =  x_2259 &  n_31515;
assign n_32540 =  x_628 &  n_26491;
assign n_32541 = ~n_32539 & ~n_32540;
assign n_32542 = ~n_32538 &  n_32541;
assign n_32543 = ~x_4081 &  n_32498;
assign n_32544 =  x_4081 & ~n_32498;
assign n_32545 = ~n_32543 & ~n_32544;
assign n_32546 = ~n_32502 & ~n_32506;
assign n_32547 =  n_32545 & ~n_32546;
assign n_32548 = ~n_32545 &  n_32546;
assign n_32549 = ~n_32547 & ~n_32548;
assign n_32550 = ~x_4880 & ~n_32549;
assign n_32551 =  x_4880 & ~n_32548;
assign n_32552 = ~n_32547 &  n_32551;
assign n_32553 =  n_26110 & ~n_32552;
assign n_32554 = ~n_32550 &  n_32553;
assign n_32555 = ~x_3712 &  n_32510;
assign n_32556 =  x_3712 & ~n_32510;
assign n_32557 = ~n_32555 & ~n_32556;
assign n_32558 = ~n_32514 & ~n_32518;
assign n_32559 =  n_32557 & ~n_32558;
assign n_32560 = ~n_32557 &  n_32558;
assign n_32561 = ~n_32559 & ~n_32560;
assign n_32562 = ~x_820 & ~n_32561;
assign n_32563 =  x_820 & ~n_32560;
assign n_32564 = ~n_32559 &  n_32563;
assign n_32565 =  n_27728 & ~n_32564;
assign n_32566 = ~n_32562 &  n_32565;
assign n_32567 = ~n_32554 & ~n_32566;
assign n_32568 =  n_32542 &  n_32567;
assign n_32569 =  x_2259 & ~n_32568;
assign n_32570 = ~x_2259 &  n_32568;
assign n_32571 = ~n_32569 & ~n_32570;
assign n_32572 = ~x_1970 &  n_32527;
assign n_32573 =  x_1970 & ~n_32527;
assign n_32574 = ~n_32572 & ~n_32573;
assign n_32575 = ~n_32531 & ~n_32535;
assign n_32576 =  n_32574 & ~n_32575;
assign n_32577 = ~n_32574 &  n_32575;
assign n_32578 = ~n_32576 & ~n_32577;
assign n_32579 = ~x_2194 & ~n_32578;
assign n_32580 =  x_2194 & ~n_32577;
assign n_32581 = ~n_32576 &  n_32580;
assign n_32582 =  n_24031 & ~n_32581;
assign n_32583 = ~n_32579 &  n_32582;
assign n_32584 =  x_2258 &  n_31515;
assign n_32585 =  x_627 &  n_26491;
assign n_32586 = ~n_32584 & ~n_32585;
assign n_32587 = ~n_32583 &  n_32586;
assign n_32588 = ~x_4080 &  n_32543;
assign n_32589 =  x_4080 & ~n_32543;
assign n_32590 = ~n_32588 & ~n_32589;
assign n_32591 = ~n_32547 & ~n_32551;
assign n_32592 =  n_32590 & ~n_32591;
assign n_32593 = ~n_32590 &  n_32591;
assign n_32594 = ~n_32592 & ~n_32593;
assign n_32595 = ~x_4879 & ~n_32594;
assign n_32596 =  x_4879 & ~n_32593;
assign n_32597 = ~n_32592 &  n_32596;
assign n_32598 =  n_26110 & ~n_32597;
assign n_32599 = ~n_32595 &  n_32598;
assign n_32600 = ~x_3711 &  n_32555;
assign n_32601 =  x_3711 & ~n_32555;
assign n_32602 = ~n_32600 & ~n_32601;
assign n_32603 = ~n_32559 & ~n_32563;
assign n_32604 =  n_32602 & ~n_32603;
assign n_32605 = ~n_32602 &  n_32603;
assign n_32606 = ~n_32604 & ~n_32605;
assign n_32607 = ~x_819 & ~n_32606;
assign n_32608 =  x_819 & ~n_32605;
assign n_32609 = ~n_32604 &  n_32608;
assign n_32610 =  n_27728 & ~n_32609;
assign n_32611 = ~n_32607 &  n_32610;
assign n_32612 = ~n_32599 & ~n_32611;
assign n_32613 =  n_32587 &  n_32612;
assign n_32614 =  x_2258 & ~n_32613;
assign n_32615 = ~x_2258 &  n_32613;
assign n_32616 = ~n_32614 & ~n_32615;
assign n_32617 = ~x_1969 &  n_32572;
assign n_32618 =  x_1969 & ~n_32572;
assign n_32619 = ~n_32617 & ~n_32618;
assign n_32620 = ~n_32576 & ~n_32580;
assign n_32621 =  n_32619 & ~n_32620;
assign n_32622 = ~n_32619 &  n_32620;
assign n_32623 = ~n_32621 & ~n_32622;
assign n_32624 = ~x_2193 & ~n_32623;
assign n_32625 =  x_2193 & ~n_32622;
assign n_32626 = ~n_32621 &  n_32625;
assign n_32627 =  n_24031 & ~n_32626;
assign n_32628 = ~n_32624 &  n_32627;
assign n_32629 =  x_2257 &  n_31515;
assign n_32630 =  x_626 &  n_26491;
assign n_32631 = ~n_32629 & ~n_32630;
assign n_32632 = ~n_32628 &  n_32631;
assign n_32633 = ~x_4079 &  n_32588;
assign n_32634 =  x_4079 & ~n_32588;
assign n_32635 = ~n_32633 & ~n_32634;
assign n_32636 = ~n_32592 & ~n_32596;
assign n_32637 =  n_32635 & ~n_32636;
assign n_32638 = ~n_32635 &  n_32636;
assign n_32639 = ~n_32637 & ~n_32638;
assign n_32640 = ~x_4878 & ~n_32639;
assign n_32641 =  x_4878 & ~n_32638;
assign n_32642 = ~n_32637 &  n_32641;
assign n_32643 =  n_26110 & ~n_32642;
assign n_32644 = ~n_32640 &  n_32643;
assign n_32645 = ~x_3710 &  n_32600;
assign n_32646 =  x_3710 & ~n_32600;
assign n_32647 = ~n_32645 & ~n_32646;
assign n_32648 = ~n_32604 & ~n_32608;
assign n_32649 =  n_32647 & ~n_32648;
assign n_32650 = ~n_32647 &  n_32648;
assign n_32651 = ~n_32649 & ~n_32650;
assign n_32652 = ~x_818 & ~n_32651;
assign n_32653 =  x_818 & ~n_32650;
assign n_32654 = ~n_32649 &  n_32653;
assign n_32655 =  n_27728 & ~n_32654;
assign n_32656 = ~n_32652 &  n_32655;
assign n_32657 = ~n_32644 & ~n_32656;
assign n_32658 =  n_32632 &  n_32657;
assign n_32659 =  x_2257 & ~n_32658;
assign n_32660 = ~x_2257 &  n_32658;
assign n_32661 = ~n_32659 & ~n_32660;
assign n_32662 = ~x_1968 &  n_32617;
assign n_32663 =  x_1968 & ~n_32617;
assign n_32664 = ~n_32662 & ~n_32663;
assign n_32665 = ~n_32621 & ~n_32625;
assign n_32666 =  n_32664 & ~n_32665;
assign n_32667 = ~n_32664 &  n_32665;
assign n_32668 = ~n_32666 & ~n_32667;
assign n_32669 = ~x_2192 & ~n_32668;
assign n_32670 =  x_2192 & ~n_32667;
assign n_32671 = ~n_32666 &  n_32670;
assign n_32672 =  n_24031 & ~n_32671;
assign n_32673 = ~n_32669 &  n_32672;
assign n_32674 =  x_2256 &  n_31515;
assign n_32675 =  x_625 &  n_26491;
assign n_32676 = ~n_32674 & ~n_32675;
assign n_32677 = ~n_32673 &  n_32676;
assign n_32678 = ~x_4078 &  n_32633;
assign n_32679 =  x_4078 & ~n_32633;
assign n_32680 = ~n_32678 & ~n_32679;
assign n_32681 = ~n_32637 & ~n_32641;
assign n_32682 =  n_32680 & ~n_32681;
assign n_32683 = ~n_32680 &  n_32681;
assign n_32684 = ~n_32682 & ~n_32683;
assign n_32685 = ~x_4877 & ~n_32684;
assign n_32686 =  x_4877 & ~n_32683;
assign n_32687 = ~n_32682 &  n_32686;
assign n_32688 =  n_26110 & ~n_32687;
assign n_32689 = ~n_32685 &  n_32688;
assign n_32690 = ~x_3709 &  n_32645;
assign n_32691 =  x_3709 & ~n_32645;
assign n_32692 = ~n_32690 & ~n_32691;
assign n_32693 = ~n_32649 & ~n_32653;
assign n_32694 =  n_32692 & ~n_32693;
assign n_32695 = ~n_32692 &  n_32693;
assign n_32696 = ~n_32694 & ~n_32695;
assign n_32697 = ~x_817 & ~n_32696;
assign n_32698 =  x_817 & ~n_32695;
assign n_32699 = ~n_32694 &  n_32698;
assign n_32700 =  n_27728 & ~n_32699;
assign n_32701 = ~n_32697 &  n_32700;
assign n_32702 = ~n_32689 & ~n_32701;
assign n_32703 =  n_32677 &  n_32702;
assign n_32704 =  x_2256 & ~n_32703;
assign n_32705 = ~x_2256 &  n_32703;
assign n_32706 = ~n_32704 & ~n_32705;
assign n_32707 = ~x_1967 &  n_32662;
assign n_32708 =  x_1967 & ~n_32662;
assign n_32709 = ~n_32707 & ~n_32708;
assign n_32710 = ~n_32666 & ~n_32670;
assign n_32711 =  n_32709 & ~n_32710;
assign n_32712 = ~n_32709 &  n_32710;
assign n_32713 = ~n_32711 & ~n_32712;
assign n_32714 = ~x_2191 & ~n_32713;
assign n_32715 =  x_2191 & ~n_32712;
assign n_32716 = ~n_32711 &  n_32715;
assign n_32717 =  n_24031 & ~n_32716;
assign n_32718 = ~n_32714 &  n_32717;
assign n_32719 =  x_2255 &  n_31515;
assign n_32720 =  x_624 &  n_26491;
assign n_32721 = ~n_32719 & ~n_32720;
assign n_32722 = ~n_32718 &  n_32721;
assign n_32723 = ~x_4077 &  n_32678;
assign n_32724 =  x_4077 & ~n_32678;
assign n_32725 = ~n_32723 & ~n_32724;
assign n_32726 = ~n_32682 & ~n_32686;
assign n_32727 =  n_32725 & ~n_32726;
assign n_32728 = ~n_32725 &  n_32726;
assign n_32729 = ~n_32727 & ~n_32728;
assign n_32730 = ~x_4876 & ~n_32729;
assign n_32731 =  x_4876 & ~n_32728;
assign n_32732 = ~n_32727 &  n_32731;
assign n_32733 =  n_26110 & ~n_32732;
assign n_32734 = ~n_32730 &  n_32733;
assign n_32735 = ~x_3708 &  n_32690;
assign n_32736 =  x_3708 & ~n_32690;
assign n_32737 = ~n_32735 & ~n_32736;
assign n_32738 = ~n_32694 & ~n_32698;
assign n_32739 =  n_32737 & ~n_32738;
assign n_32740 = ~n_32737 &  n_32738;
assign n_32741 = ~n_32739 & ~n_32740;
assign n_32742 = ~x_816 & ~n_32741;
assign n_32743 =  x_816 & ~n_32740;
assign n_32744 = ~n_32739 &  n_32743;
assign n_32745 =  n_27728 & ~n_32744;
assign n_32746 = ~n_32742 &  n_32745;
assign n_32747 = ~n_32734 & ~n_32746;
assign n_32748 =  n_32722 &  n_32747;
assign n_32749 =  x_2255 & ~n_32748;
assign n_32750 = ~x_2255 &  n_32748;
assign n_32751 = ~n_32749 & ~n_32750;
assign n_32752 = ~x_1966 &  n_32707;
assign n_32753 =  x_1966 & ~n_32707;
assign n_32754 = ~n_32752 & ~n_32753;
assign n_32755 = ~n_32711 & ~n_32715;
assign n_32756 =  n_32754 & ~n_32755;
assign n_32757 = ~n_32754 &  n_32755;
assign n_32758 = ~n_32756 & ~n_32757;
assign n_32759 = ~x_2190 & ~n_32758;
assign n_32760 =  x_2190 & ~n_32757;
assign n_32761 = ~n_32756 &  n_32760;
assign n_32762 =  n_24031 & ~n_32761;
assign n_32763 = ~n_32759 &  n_32762;
assign n_32764 =  x_2254 &  n_31515;
assign n_32765 =  x_623 &  n_26491;
assign n_32766 = ~n_32764 & ~n_32765;
assign n_32767 = ~n_32763 &  n_32766;
assign n_32768 = ~x_4076 &  n_32723;
assign n_32769 =  x_4076 & ~n_32723;
assign n_32770 = ~n_32768 & ~n_32769;
assign n_32771 = ~n_32727 & ~n_32731;
assign n_32772 =  n_32770 & ~n_32771;
assign n_32773 = ~n_32770 &  n_32771;
assign n_32774 = ~n_32772 & ~n_32773;
assign n_32775 = ~x_4875 & ~n_32774;
assign n_32776 =  x_4875 & ~n_32773;
assign n_32777 = ~n_32772 &  n_32776;
assign n_32778 =  n_26110 & ~n_32777;
assign n_32779 = ~n_32775 &  n_32778;
assign n_32780 = ~x_3707 &  n_32735;
assign n_32781 =  x_3707 & ~n_32735;
assign n_32782 = ~n_32780 & ~n_32781;
assign n_32783 = ~n_32739 & ~n_32743;
assign n_32784 =  n_32782 & ~n_32783;
assign n_32785 = ~n_32782 &  n_32783;
assign n_32786 = ~n_32784 & ~n_32785;
assign n_32787 = ~x_815 & ~n_32786;
assign n_32788 =  x_815 & ~n_32785;
assign n_32789 = ~n_32784 &  n_32788;
assign n_32790 =  n_27728 & ~n_32789;
assign n_32791 = ~n_32787 &  n_32790;
assign n_32792 = ~n_32779 & ~n_32791;
assign n_32793 =  n_32767 &  n_32792;
assign n_32794 =  x_2254 & ~n_32793;
assign n_32795 = ~x_2254 &  n_32793;
assign n_32796 = ~n_32794 & ~n_32795;
assign n_32797 = ~x_1965 &  n_32752;
assign n_32798 =  x_1965 & ~n_32752;
assign n_32799 = ~n_32797 & ~n_32798;
assign n_32800 = ~n_32756 & ~n_32760;
assign n_32801 =  n_32799 & ~n_32800;
assign n_32802 = ~n_32799 &  n_32800;
assign n_32803 = ~n_32801 & ~n_32802;
assign n_32804 = ~x_2189 & ~n_32803;
assign n_32805 =  x_2189 & ~n_32802;
assign n_32806 = ~n_32801 &  n_32805;
assign n_32807 =  n_24031 & ~n_32806;
assign n_32808 = ~n_32804 &  n_32807;
assign n_32809 =  x_2253 &  n_31515;
assign n_32810 =  x_622 &  n_26491;
assign n_32811 = ~n_32809 & ~n_32810;
assign n_32812 = ~n_32808 &  n_32811;
assign n_32813 = ~x_4075 &  n_32768;
assign n_32814 =  x_4075 & ~n_32768;
assign n_32815 = ~n_32813 & ~n_32814;
assign n_32816 = ~n_32772 & ~n_32776;
assign n_32817 =  n_32815 & ~n_32816;
assign n_32818 = ~n_32815 &  n_32816;
assign n_32819 = ~n_32817 & ~n_32818;
assign n_32820 = ~x_4874 & ~n_32819;
assign n_32821 =  x_4874 & ~n_32818;
assign n_32822 = ~n_32817 &  n_32821;
assign n_32823 =  n_26110 & ~n_32822;
assign n_32824 = ~n_32820 &  n_32823;
assign n_32825 = ~x_3706 &  n_32780;
assign n_32826 =  x_3706 & ~n_32780;
assign n_32827 = ~n_32825 & ~n_32826;
assign n_32828 = ~n_32784 & ~n_32788;
assign n_32829 =  n_32827 & ~n_32828;
assign n_32830 = ~n_32827 &  n_32828;
assign n_32831 = ~n_32829 & ~n_32830;
assign n_32832 = ~x_814 & ~n_32831;
assign n_32833 =  x_814 & ~n_32830;
assign n_32834 = ~n_32829 &  n_32833;
assign n_32835 =  n_27728 & ~n_32834;
assign n_32836 = ~n_32832 &  n_32835;
assign n_32837 = ~n_32824 & ~n_32836;
assign n_32838 =  n_32812 &  n_32837;
assign n_32839 =  x_2253 & ~n_32838;
assign n_32840 = ~x_2253 &  n_32838;
assign n_32841 = ~n_32839 & ~n_32840;
assign n_32842 = ~x_1964 &  n_32797;
assign n_32843 =  x_1964 & ~n_32797;
assign n_32844 = ~n_32842 & ~n_32843;
assign n_32845 = ~n_32801 & ~n_32805;
assign n_32846 =  n_32844 & ~n_32845;
assign n_32847 = ~n_32844 &  n_32845;
assign n_32848 = ~n_32846 & ~n_32847;
assign n_32849 = ~x_2188 & ~n_32848;
assign n_32850 =  x_2188 & ~n_32847;
assign n_32851 = ~n_32846 &  n_32850;
assign n_32852 =  n_24031 & ~n_32851;
assign n_32853 = ~n_32849 &  n_32852;
assign n_32854 =  x_2252 &  n_31515;
assign n_32855 =  x_621 &  n_26491;
assign n_32856 = ~n_32854 & ~n_32855;
assign n_32857 = ~n_32853 &  n_32856;
assign n_32858 = ~x_4074 &  n_32813;
assign n_32859 =  x_4074 & ~n_32813;
assign n_32860 = ~n_32858 & ~n_32859;
assign n_32861 = ~n_32817 & ~n_32821;
assign n_32862 =  n_32860 & ~n_32861;
assign n_32863 = ~n_32860 &  n_32861;
assign n_32864 = ~n_32862 & ~n_32863;
assign n_32865 = ~x_4873 & ~n_32864;
assign n_32866 =  x_4873 & ~n_32863;
assign n_32867 = ~n_32862 &  n_32866;
assign n_32868 =  n_26110 & ~n_32867;
assign n_32869 = ~n_32865 &  n_32868;
assign n_32870 = ~x_3705 &  n_32825;
assign n_32871 =  x_3705 & ~n_32825;
assign n_32872 = ~n_32870 & ~n_32871;
assign n_32873 = ~n_32829 & ~n_32833;
assign n_32874 =  n_32872 & ~n_32873;
assign n_32875 = ~n_32872 &  n_32873;
assign n_32876 = ~n_32874 & ~n_32875;
assign n_32877 = ~x_813 & ~n_32876;
assign n_32878 =  x_813 & ~n_32875;
assign n_32879 = ~n_32874 &  n_32878;
assign n_32880 =  n_27728 & ~n_32879;
assign n_32881 = ~n_32877 &  n_32880;
assign n_32882 = ~n_32869 & ~n_32881;
assign n_32883 =  n_32857 &  n_32882;
assign n_32884 =  x_2252 & ~n_32883;
assign n_32885 = ~x_2252 &  n_32883;
assign n_32886 = ~n_32884 & ~n_32885;
assign n_32887 = ~n_32846 & ~n_32850;
assign n_32888 =  x_1963 & ~x_2187;
assign n_32889 = ~x_1963 &  x_2187;
assign n_32890 = ~n_32888 & ~n_32889;
assign n_32891 =  n_32842 &  n_32890;
assign n_32892 = ~n_32842 & ~n_32890;
assign n_32893 = ~n_32891 & ~n_32892;
assign n_32894 =  n_32887 & ~n_32893;
assign n_32895 = ~n_32887 &  n_32893;
assign n_32896 =  n_24031 & ~n_32895;
assign n_32897 = ~n_32894 &  n_32896;
assign n_32898 =  x_620 &  n_26491;
assign n_32899 =  x_2251 &  n_31515;
assign n_32900 = ~n_32898 & ~n_32899;
assign n_32901 = ~n_32897 &  n_32900;
assign n_32902 = ~n_32874 & ~n_32878;
assign n_32903 =  x_812 & ~x_3704;
assign n_32904 = ~x_812 &  x_3704;
assign n_32905 = ~n_32903 & ~n_32904;
assign n_32906 =  n_32870 &  n_32905;
assign n_32907 = ~n_32870 & ~n_32905;
assign n_32908 = ~n_32906 & ~n_32907;
assign n_32909 =  n_32902 & ~n_32908;
assign n_32910 = ~n_32902 &  n_32908;
assign n_32911 =  n_27728 & ~n_32910;
assign n_32912 = ~n_32909 &  n_32911;
assign n_32913 = ~n_32862 & ~n_32866;
assign n_32914 =  x_4073 & ~x_4872;
assign n_32915 = ~x_4073 &  x_4872;
assign n_32916 = ~n_32914 & ~n_32915;
assign n_32917 =  n_32858 &  n_32916;
assign n_32918 = ~n_32858 & ~n_32916;
assign n_32919 = ~n_32917 & ~n_32918;
assign n_32920 = ~n_32913 &  n_32919;
assign n_32921 =  n_32913 & ~n_32919;
assign n_32922 =  n_26110 & ~n_32921;
assign n_32923 = ~n_32920 &  n_32922;
assign n_32924 = ~n_32912 & ~n_32923;
assign n_32925 =  n_32901 &  n_32924;
assign n_32926 =  x_2251 & ~n_32925;
assign n_32927 = ~x_2251 &  n_32925;
assign n_32928 = ~n_32926 & ~n_32927;
assign n_32929 =  x_2250 & ~n_24007;
assign n_32930 =  x_2250 &  n_32929;
assign n_32931 = ~x_2250 & ~n_32929;
assign n_32932 = ~n_32930 & ~n_32931;
assign n_32933 =  x_2249 & ~n_24007;
assign n_32934 =  x_2249 &  n_32933;
assign n_32935 = ~x_2249 & ~n_32933;
assign n_32936 = ~n_32934 & ~n_32935;
assign n_32937 =  x_2248 & ~n_24007;
assign n_32938 =  x_2248 &  n_32937;
assign n_32939 = ~x_2248 & ~n_32937;
assign n_32940 = ~n_32938 & ~n_32939;
assign n_32941 =  x_2247 & ~n_24007;
assign n_32942 =  x_2247 &  n_32941;
assign n_32943 = ~x_2247 & ~n_32941;
assign n_32944 = ~n_32942 & ~n_32943;
assign n_32945 =  x_2246 & ~n_24007;
assign n_32946 =  x_2246 &  n_32945;
assign n_32947 = ~x_2246 & ~n_32945;
assign n_32948 = ~n_32946 & ~n_32947;
assign n_32949 =  x_2245 & ~n_24007;
assign n_32950 =  x_2245 &  n_32949;
assign n_32951 = ~x_2245 & ~n_32949;
assign n_32952 = ~n_32950 & ~n_32951;
assign n_32953 =  x_2244 & ~n_24007;
assign n_32954 =  x_2244 &  n_32953;
assign n_32955 = ~x_2244 & ~n_32953;
assign n_32956 = ~n_32954 & ~n_32955;
assign n_32957 =  x_2243 & ~n_24007;
assign n_32958 =  x_2243 &  n_32957;
assign n_32959 = ~x_2243 & ~n_32957;
assign n_32960 = ~n_32958 & ~n_32959;
assign n_32961 =  x_2242 & ~n_24007;
assign n_32962 =  x_2242 &  n_32961;
assign n_32963 = ~x_2242 & ~n_32961;
assign n_32964 = ~n_32962 & ~n_32963;
assign n_32965 =  x_2241 & ~n_24007;
assign n_32966 =  x_2241 &  n_32965;
assign n_32967 = ~x_2241 & ~n_32965;
assign n_32968 = ~n_32966 & ~n_32967;
assign n_32969 =  x_2240 & ~n_24007;
assign n_32970 =  x_2240 &  n_32969;
assign n_32971 = ~x_2240 & ~n_32969;
assign n_32972 = ~n_32970 & ~n_32971;
assign n_32973 =  x_2239 & ~n_24007;
assign n_32974 =  x_2239 &  n_32973;
assign n_32975 = ~x_2239 & ~n_32973;
assign n_32976 = ~n_32974 & ~n_32975;
assign n_32977 =  x_2238 & ~n_24007;
assign n_32978 =  x_2238 &  n_32977;
assign n_32979 = ~x_2238 & ~n_32977;
assign n_32980 = ~n_32978 & ~n_32979;
assign n_32981 =  x_2237 & ~n_24007;
assign n_32982 =  x_2237 &  n_32981;
assign n_32983 = ~x_2237 & ~n_32981;
assign n_32984 = ~n_32982 & ~n_32983;
assign n_32985 =  x_2236 & ~n_24007;
assign n_32986 =  x_2236 &  n_32985;
assign n_32987 = ~x_2236 & ~n_32985;
assign n_32988 = ~n_32986 & ~n_32987;
assign n_32989 =  x_2235 & ~n_24007;
assign n_32990 =  x_2235 &  n_32989;
assign n_32991 = ~x_2235 & ~n_32989;
assign n_32992 = ~n_32990 & ~n_32991;
assign n_32993 =  x_2234 & ~n_24007;
assign n_32994 =  x_2234 &  n_32993;
assign n_32995 = ~x_2234 & ~n_32993;
assign n_32996 = ~n_32994 & ~n_32995;
assign n_32997 =  x_2233 & ~n_24007;
assign n_32998 =  x_2233 &  n_32997;
assign n_32999 = ~x_2233 & ~n_32997;
assign n_33000 = ~n_32998 & ~n_32999;
assign n_33001 =  x_2232 & ~n_24007;
assign n_33002 =  x_2232 &  n_33001;
assign n_33003 = ~x_2232 & ~n_33001;
assign n_33004 = ~n_33002 & ~n_33003;
assign n_33005 =  x_2231 & ~n_24007;
assign n_33006 =  x_2231 &  n_33005;
assign n_33007 = ~x_2231 & ~n_33005;
assign n_33008 = ~n_33006 & ~n_33007;
assign n_33009 =  x_2230 & ~n_24007;
assign n_33010 =  x_2230 &  n_33009;
assign n_33011 = ~x_2230 & ~n_33009;
assign n_33012 = ~n_33010 & ~n_33011;
assign n_33013 =  x_2229 & ~n_24007;
assign n_33014 =  x_2229 &  n_33013;
assign n_33015 = ~x_2229 & ~n_33013;
assign n_33016 = ~n_33014 & ~n_33015;
assign n_33017 =  x_2228 & ~n_24007;
assign n_33018 =  x_2228 &  n_33017;
assign n_33019 = ~x_2228 & ~n_33017;
assign n_33020 = ~n_33018 & ~n_33019;
assign n_33021 =  x_2227 & ~n_24007;
assign n_33022 =  x_2227 &  n_33021;
assign n_33023 = ~x_2227 & ~n_33021;
assign n_33024 = ~n_33022 & ~n_33023;
assign n_33025 =  x_2226 & ~n_24007;
assign n_33026 =  x_2226 &  n_33025;
assign n_33027 = ~x_2226 & ~n_33025;
assign n_33028 = ~n_33026 & ~n_33027;
assign n_33029 =  x_2225 & ~n_24007;
assign n_33030 =  x_2225 &  n_33029;
assign n_33031 = ~x_2225 & ~n_33029;
assign n_33032 = ~n_33030 & ~n_33031;
assign n_33033 =  x_2224 & ~n_24007;
assign n_33034 =  x_2224 &  n_33033;
assign n_33035 = ~x_2224 & ~n_33033;
assign n_33036 = ~n_33034 & ~n_33035;
assign n_33037 =  x_2223 & ~n_24007;
assign n_33038 =  x_2223 &  n_33037;
assign n_33039 = ~x_2223 & ~n_33037;
assign n_33040 = ~n_33038 & ~n_33039;
assign n_33041 =  x_2222 & ~n_24007;
assign n_33042 =  x_2222 &  n_33041;
assign n_33043 = ~x_2222 & ~n_33041;
assign n_33044 = ~n_33042 & ~n_33043;
assign n_33045 =  x_2221 & ~n_24007;
assign n_33046 =  x_2221 &  n_33045;
assign n_33047 = ~x_2221 & ~n_33045;
assign n_33048 = ~n_33046 & ~n_33047;
assign n_33049 =  x_2220 & ~n_24007;
assign n_33050 =  x_2220 &  n_33049;
assign n_33051 = ~x_2220 & ~n_33049;
assign n_33052 = ~n_33050 & ~n_33051;
assign n_33053 =  x_2219 & ~n_24007;
assign n_33054 =  x_2219 &  n_33053;
assign n_33055 = ~x_2219 & ~n_33053;
assign n_33056 = ~n_33054 & ~n_33055;
assign n_33057 =  x_2218 & ~n_25169;
assign n_33058 =  x_2218 &  n_33057;
assign n_33059 = ~x_2218 & ~n_33057;
assign n_33060 = ~n_33058 & ~n_33059;
assign n_33061 =  x_2217 & ~n_25169;
assign n_33062 =  x_2217 &  n_33061;
assign n_33063 = ~x_2217 & ~n_33061;
assign n_33064 = ~n_33062 & ~n_33063;
assign n_33065 =  x_2216 & ~n_25169;
assign n_33066 =  x_2216 &  n_33065;
assign n_33067 = ~x_2216 & ~n_33065;
assign n_33068 = ~n_33066 & ~n_33067;
assign n_33069 =  x_2215 & ~n_25169;
assign n_33070 =  x_2215 &  n_33069;
assign n_33071 = ~x_2215 & ~n_33069;
assign n_33072 = ~n_33070 & ~n_33071;
assign n_33073 =  x_2214 & ~n_25169;
assign n_33074 =  x_2214 &  n_33073;
assign n_33075 = ~x_2214 & ~n_33073;
assign n_33076 = ~n_33074 & ~n_33075;
assign n_33077 =  x_2213 & ~n_25169;
assign n_33078 =  x_2213 &  n_33077;
assign n_33079 = ~x_2213 & ~n_33077;
assign n_33080 = ~n_33078 & ~n_33079;
assign n_33081 =  x_2212 & ~n_25169;
assign n_33082 =  x_2212 &  n_33081;
assign n_33083 = ~x_2212 & ~n_33081;
assign n_33084 = ~n_33082 & ~n_33083;
assign n_33085 =  x_2211 & ~n_25169;
assign n_33086 =  x_2211 &  n_33085;
assign n_33087 = ~x_2211 & ~n_33085;
assign n_33088 = ~n_33086 & ~n_33087;
assign n_33089 =  x_2210 & ~n_25169;
assign n_33090 =  x_2210 &  n_33089;
assign n_33091 = ~x_2210 & ~n_33089;
assign n_33092 = ~n_33090 & ~n_33091;
assign n_33093 =  x_2209 & ~n_25169;
assign n_33094 =  x_2209 &  n_33093;
assign n_33095 = ~x_2209 & ~n_33093;
assign n_33096 = ~n_33094 & ~n_33095;
assign n_33097 =  x_2208 & ~n_25169;
assign n_33098 =  x_2208 &  n_33097;
assign n_33099 = ~x_2208 & ~n_33097;
assign n_33100 = ~n_33098 & ~n_33099;
assign n_33101 =  x_2207 & ~n_25169;
assign n_33102 =  x_2207 &  n_33101;
assign n_33103 = ~x_2207 & ~n_33101;
assign n_33104 = ~n_33102 & ~n_33103;
assign n_33105 =  x_2206 & ~n_25169;
assign n_33106 =  x_2206 &  n_33105;
assign n_33107 = ~x_2206 & ~n_33105;
assign n_33108 = ~n_33106 & ~n_33107;
assign n_33109 =  x_2205 & ~n_25169;
assign n_33110 =  x_2205 &  n_33109;
assign n_33111 = ~x_2205 & ~n_33109;
assign n_33112 = ~n_33110 & ~n_33111;
assign n_33113 =  x_2204 & ~n_25169;
assign n_33114 =  x_2204 &  n_33113;
assign n_33115 = ~x_2204 & ~n_33113;
assign n_33116 = ~n_33114 & ~n_33115;
assign n_33117 =  x_2203 & ~n_25169;
assign n_33118 =  x_2203 &  n_33117;
assign n_33119 = ~x_2203 & ~n_33117;
assign n_33120 = ~n_33118 & ~n_33119;
assign n_33121 =  x_2202 & ~n_25169;
assign n_33122 =  x_2202 &  n_33121;
assign n_33123 = ~x_2202 & ~n_33121;
assign n_33124 = ~n_33122 & ~n_33123;
assign n_33125 =  x_2201 & ~n_25169;
assign n_33126 =  x_2201 &  n_33125;
assign n_33127 = ~x_2201 & ~n_33125;
assign n_33128 = ~n_33126 & ~n_33127;
assign n_33129 =  x_2200 & ~n_25169;
assign n_33130 =  x_2200 &  n_33129;
assign n_33131 = ~x_2200 & ~n_33129;
assign n_33132 = ~n_33130 & ~n_33131;
assign n_33133 =  x_2199 & ~n_25169;
assign n_33134 =  x_2199 &  n_33133;
assign n_33135 = ~x_2199 & ~n_33133;
assign n_33136 = ~n_33134 & ~n_33135;
assign n_33137 =  x_2198 & ~n_25169;
assign n_33138 =  x_2198 &  n_33137;
assign n_33139 = ~x_2198 & ~n_33137;
assign n_33140 = ~n_33138 & ~n_33139;
assign n_33141 =  x_2197 & ~n_25169;
assign n_33142 =  x_2197 &  n_33141;
assign n_33143 = ~x_2197 & ~n_33141;
assign n_33144 = ~n_33142 & ~n_33143;
assign n_33145 =  x_2196 & ~n_25169;
assign n_33146 =  x_2196 &  n_33145;
assign n_33147 = ~x_2196 & ~n_33145;
assign n_33148 = ~n_33146 & ~n_33147;
assign n_33149 =  x_2195 & ~n_25169;
assign n_33150 =  x_2195 &  n_33149;
assign n_33151 = ~x_2195 & ~n_33149;
assign n_33152 = ~n_33150 & ~n_33151;
assign n_33153 =  x_2194 & ~n_25169;
assign n_33154 =  x_2194 &  n_33153;
assign n_33155 = ~x_2194 & ~n_33153;
assign n_33156 = ~n_33154 & ~n_33155;
assign n_33157 =  x_2193 & ~n_25169;
assign n_33158 =  x_2193 &  n_33157;
assign n_33159 = ~x_2193 & ~n_33157;
assign n_33160 = ~n_33158 & ~n_33159;
assign n_33161 =  x_2192 & ~n_25169;
assign n_33162 =  x_2192 &  n_33161;
assign n_33163 = ~x_2192 & ~n_33161;
assign n_33164 = ~n_33162 & ~n_33163;
assign n_33165 =  x_2191 & ~n_25169;
assign n_33166 =  x_2191 &  n_33165;
assign n_33167 = ~x_2191 & ~n_33165;
assign n_33168 = ~n_33166 & ~n_33167;
assign n_33169 =  x_2190 & ~n_25169;
assign n_33170 =  x_2190 &  n_33169;
assign n_33171 = ~x_2190 & ~n_33169;
assign n_33172 = ~n_33170 & ~n_33171;
assign n_33173 =  x_2189 & ~n_25169;
assign n_33174 =  x_2189 &  n_33173;
assign n_33175 = ~x_2189 & ~n_33173;
assign n_33176 = ~n_33174 & ~n_33175;
assign n_33177 =  x_2188 & ~n_25169;
assign n_33178 =  x_2188 &  n_33177;
assign n_33179 = ~x_2188 & ~n_33177;
assign n_33180 = ~n_33178 & ~n_33179;
assign n_33181 =  x_2187 & ~n_25169;
assign n_33182 =  x_2187 &  n_33181;
assign n_33183 = ~x_2187 & ~n_33181;
assign n_33184 = ~n_33182 & ~n_33183;
assign n_33185 = ~n_27721 &  n_9430;
assign n_33186 = ~n_33185 & ~n_9428;
assign n_33187 =  x_2186 & ~n_33186;
assign n_33188 =  x_3255 &  n_27721;
assign n_33189 =  x_4935 &  n_558;
assign n_33190 = ~n_33188 & ~n_33189;
assign n_33191 = ~n_33187 &  n_33190;
assign n_33192 =  x_2186 & ~n_33191;
assign n_33193 = ~x_2186 &  n_33191;
assign n_33194 = ~n_33192 & ~n_33193;
assign n_33195 =  x_2185 & ~n_33186;
assign n_33196 =  x_3254 &  n_27721;
assign n_33197 =  x_4934 &  n_558;
assign n_33198 = ~n_33196 & ~n_33197;
assign n_33199 = ~n_33195 &  n_33198;
assign n_33200 =  x_2185 & ~n_33199;
assign n_33201 = ~x_2185 &  n_33199;
assign n_33202 = ~n_33200 & ~n_33201;
assign n_33203 =  x_2184 & ~n_33186;
assign n_33204 =  x_3253 &  n_27721;
assign n_33205 =  x_4933 &  n_558;
assign n_33206 = ~n_33204 & ~n_33205;
assign n_33207 = ~n_33203 &  n_33206;
assign n_33208 =  x_2184 & ~n_33207;
assign n_33209 = ~x_2184 &  n_33207;
assign n_33210 = ~n_33208 & ~n_33209;
assign n_33211 =  x_2183 & ~n_33186;
assign n_33212 =  x_3252 &  n_27721;
assign n_33213 =  x_4932 &  n_558;
assign n_33214 = ~n_33212 & ~n_33213;
assign n_33215 = ~n_33211 &  n_33214;
assign n_33216 =  x_2183 & ~n_33215;
assign n_33217 = ~x_2183 &  n_33215;
assign n_33218 = ~n_33216 & ~n_33217;
assign n_33219 =  x_2182 & ~n_33186;
assign n_33220 =  x_3251 &  n_27721;
assign n_33221 =  x_4931 &  n_558;
assign n_33222 = ~n_33220 & ~n_33221;
assign n_33223 = ~n_33219 &  n_33222;
assign n_33224 =  x_2182 & ~n_33223;
assign n_33225 = ~x_2182 &  n_33223;
assign n_33226 = ~n_33224 & ~n_33225;
assign n_33227 =  x_2181 & ~n_33186;
assign n_33228 =  x_3250 &  n_27721;
assign n_33229 =  x_4930 &  n_558;
assign n_33230 = ~n_33228 & ~n_33229;
assign n_33231 = ~n_33227 &  n_33230;
assign n_33232 =  x_2181 & ~n_33231;
assign n_33233 = ~x_2181 &  n_33231;
assign n_33234 = ~n_33232 & ~n_33233;
assign n_33235 =  x_2180 & ~n_33186;
assign n_33236 =  x_3249 &  n_27721;
assign n_33237 =  x_4929 &  n_558;
assign n_33238 = ~n_33236 & ~n_33237;
assign n_33239 = ~n_33235 &  n_33238;
assign n_33240 =  x_2180 & ~n_33239;
assign n_33241 = ~x_2180 &  n_33239;
assign n_33242 = ~n_33240 & ~n_33241;
assign n_33243 =  x_2179 & ~n_33186;
assign n_33244 =  x_3248 &  n_27721;
assign n_33245 =  x_4928 &  n_558;
assign n_33246 = ~n_33244 & ~n_33245;
assign n_33247 = ~n_33243 &  n_33246;
assign n_33248 =  x_2179 & ~n_33247;
assign n_33249 = ~x_2179 &  n_33247;
assign n_33250 = ~n_33248 & ~n_33249;
assign n_33251 =  x_2178 & ~n_33186;
assign n_33252 =  x_3247 &  n_27721;
assign n_33253 =  x_4927 &  n_558;
assign n_33254 = ~n_33252 & ~n_33253;
assign n_33255 = ~n_33251 &  n_33254;
assign n_33256 =  x_2178 & ~n_33255;
assign n_33257 = ~x_2178 &  n_33255;
assign n_33258 = ~n_33256 & ~n_33257;
assign n_33259 =  x_2177 & ~n_33186;
assign n_33260 =  x_3246 &  n_27721;
assign n_33261 =  x_4926 &  n_558;
assign n_33262 = ~n_33260 & ~n_33261;
assign n_33263 = ~n_33259 &  n_33262;
assign n_33264 =  x_2177 & ~n_33263;
assign n_33265 = ~x_2177 &  n_33263;
assign n_33266 = ~n_33264 & ~n_33265;
assign n_33267 =  x_2176 & ~n_33186;
assign n_33268 =  x_3245 &  n_27721;
assign n_33269 =  x_4925 &  n_558;
assign n_33270 = ~n_33268 & ~n_33269;
assign n_33271 = ~n_33267 &  n_33270;
assign n_33272 =  x_2176 & ~n_33271;
assign n_33273 = ~x_2176 &  n_33271;
assign n_33274 = ~n_33272 & ~n_33273;
assign n_33275 =  x_2175 & ~n_33186;
assign n_33276 =  x_3244 &  n_27721;
assign n_33277 =  x_4924 &  n_558;
assign n_33278 = ~n_33276 & ~n_33277;
assign n_33279 = ~n_33275 &  n_33278;
assign n_33280 =  x_2175 & ~n_33279;
assign n_33281 = ~x_2175 &  n_33279;
assign n_33282 = ~n_33280 & ~n_33281;
assign n_33283 =  x_2174 & ~n_33186;
assign n_33284 =  x_3243 &  n_27721;
assign n_33285 =  x_4923 &  n_558;
assign n_33286 = ~n_33284 & ~n_33285;
assign n_33287 = ~n_33283 &  n_33286;
assign n_33288 =  x_2174 & ~n_33287;
assign n_33289 = ~x_2174 &  n_33287;
assign n_33290 = ~n_33288 & ~n_33289;
assign n_33291 =  x_2173 & ~n_33186;
assign n_33292 =  x_3242 &  n_27721;
assign n_33293 =  x_4922 &  n_558;
assign n_33294 = ~n_33292 & ~n_33293;
assign n_33295 = ~n_33291 &  n_33294;
assign n_33296 =  x_2173 & ~n_33295;
assign n_33297 = ~x_2173 &  n_33295;
assign n_33298 = ~n_33296 & ~n_33297;
assign n_33299 =  x_2172 & ~n_33186;
assign n_33300 =  x_3241 &  n_27721;
assign n_33301 =  x_4921 &  n_558;
assign n_33302 = ~n_33300 & ~n_33301;
assign n_33303 = ~n_33299 &  n_33302;
assign n_33304 =  x_2172 & ~n_33303;
assign n_33305 = ~x_2172 &  n_33303;
assign n_33306 = ~n_33304 & ~n_33305;
assign n_33307 =  x_2171 & ~n_33186;
assign n_33308 =  x_3240 &  n_27721;
assign n_33309 =  x_4920 &  n_558;
assign n_33310 = ~n_33308 & ~n_33309;
assign n_33311 = ~n_33307 &  n_33310;
assign n_33312 =  x_2171 & ~n_33311;
assign n_33313 = ~x_2171 &  n_33311;
assign n_33314 = ~n_33312 & ~n_33313;
assign n_33315 =  x_2170 & ~n_33186;
assign n_33316 =  x_3239 &  n_27721;
assign n_33317 =  x_4919 &  n_558;
assign n_33318 = ~n_33316 & ~n_33317;
assign n_33319 = ~n_33315 &  n_33318;
assign n_33320 =  x_2170 & ~n_33319;
assign n_33321 = ~x_2170 &  n_33319;
assign n_33322 = ~n_33320 & ~n_33321;
assign n_33323 =  x_2169 & ~n_33186;
assign n_33324 =  x_3238 &  n_27721;
assign n_33325 =  x_4918 &  n_558;
assign n_33326 = ~n_33324 & ~n_33325;
assign n_33327 = ~n_33323 &  n_33326;
assign n_33328 =  x_2169 & ~n_33327;
assign n_33329 = ~x_2169 &  n_33327;
assign n_33330 = ~n_33328 & ~n_33329;
assign n_33331 =  x_2168 & ~n_33186;
assign n_33332 =  x_3237 &  n_27721;
assign n_33333 =  x_4917 &  n_558;
assign n_33334 = ~n_33332 & ~n_33333;
assign n_33335 = ~n_33331 &  n_33334;
assign n_33336 =  x_2168 & ~n_33335;
assign n_33337 = ~x_2168 &  n_33335;
assign n_33338 = ~n_33336 & ~n_33337;
assign n_33339 =  x_2167 & ~n_33186;
assign n_33340 =  x_3236 &  n_27721;
assign n_33341 =  x_4916 &  n_558;
assign n_33342 = ~n_33340 & ~n_33341;
assign n_33343 = ~n_33339 &  n_33342;
assign n_33344 =  x_2167 & ~n_33343;
assign n_33345 = ~x_2167 &  n_33343;
assign n_33346 = ~n_33344 & ~n_33345;
assign n_33347 =  x_2166 & ~n_33186;
assign n_33348 =  x_3235 &  n_27721;
assign n_33349 =  x_4915 &  n_558;
assign n_33350 = ~n_33348 & ~n_33349;
assign n_33351 = ~n_33347 &  n_33350;
assign n_33352 =  x_2166 & ~n_33351;
assign n_33353 = ~x_2166 &  n_33351;
assign n_33354 = ~n_33352 & ~n_33353;
assign n_33355 =  x_2165 & ~n_33186;
assign n_33356 =  x_3234 &  n_27721;
assign n_33357 =  x_4914 &  n_558;
assign n_33358 = ~n_33356 & ~n_33357;
assign n_33359 = ~n_33355 &  n_33358;
assign n_33360 =  x_2165 & ~n_33359;
assign n_33361 = ~x_2165 &  n_33359;
assign n_33362 = ~n_33360 & ~n_33361;
assign n_33363 =  x_2164 & ~n_33186;
assign n_33364 =  x_3233 &  n_27721;
assign n_33365 =  x_4913 &  n_558;
assign n_33366 = ~n_33364 & ~n_33365;
assign n_33367 = ~n_33363 &  n_33366;
assign n_33368 =  x_2164 & ~n_33367;
assign n_33369 = ~x_2164 &  n_33367;
assign n_33370 = ~n_33368 & ~n_33369;
assign n_33371 =  x_2163 & ~n_33186;
assign n_33372 =  x_3232 &  n_27721;
assign n_33373 =  x_4912 &  n_558;
assign n_33374 = ~n_33372 & ~n_33373;
assign n_33375 = ~n_33371 &  n_33374;
assign n_33376 =  x_2163 & ~n_33375;
assign n_33377 = ~x_2163 &  n_33375;
assign n_33378 = ~n_33376 & ~n_33377;
assign n_33379 =  x_2162 & ~n_33186;
assign n_33380 =  x_3231 &  n_27721;
assign n_33381 =  x_4911 &  n_558;
assign n_33382 = ~n_33380 & ~n_33381;
assign n_33383 = ~n_33379 &  n_33382;
assign n_33384 =  x_2162 & ~n_33383;
assign n_33385 = ~x_2162 &  n_33383;
assign n_33386 = ~n_33384 & ~n_33385;
assign n_33387 =  x_2161 & ~n_33186;
assign n_33388 =  x_3230 &  n_27721;
assign n_33389 =  x_4910 &  n_558;
assign n_33390 = ~n_33388 & ~n_33389;
assign n_33391 = ~n_33387 &  n_33390;
assign n_33392 =  x_2161 & ~n_33391;
assign n_33393 = ~x_2161 &  n_33391;
assign n_33394 = ~n_33392 & ~n_33393;
assign n_33395 =  x_2160 & ~n_33186;
assign n_33396 =  x_3229 &  n_27721;
assign n_33397 =  x_4909 &  n_558;
assign n_33398 = ~n_33396 & ~n_33397;
assign n_33399 = ~n_33395 &  n_33398;
assign n_33400 =  x_2160 & ~n_33399;
assign n_33401 = ~x_2160 &  n_33399;
assign n_33402 = ~n_33400 & ~n_33401;
assign n_33403 =  x_2159 & ~n_33186;
assign n_33404 =  x_3228 &  n_27721;
assign n_33405 =  x_4908 &  n_558;
assign n_33406 = ~n_33404 & ~n_33405;
assign n_33407 = ~n_33403 &  n_33406;
assign n_33408 =  x_2159 & ~n_33407;
assign n_33409 = ~x_2159 &  n_33407;
assign n_33410 = ~n_33408 & ~n_33409;
assign n_33411 =  x_2158 & ~n_33186;
assign n_33412 =  x_3227 &  n_27721;
assign n_33413 =  x_4907 &  n_558;
assign n_33414 = ~n_33412 & ~n_33413;
assign n_33415 = ~n_33411 &  n_33414;
assign n_33416 =  x_2158 & ~n_33415;
assign n_33417 = ~x_2158 &  n_33415;
assign n_33418 = ~n_33416 & ~n_33417;
assign n_33419 =  x_2157 & ~n_33186;
assign n_33420 =  x_3226 &  n_27721;
assign n_33421 =  x_4906 &  n_558;
assign n_33422 = ~n_33420 & ~n_33421;
assign n_33423 = ~n_33419 &  n_33422;
assign n_33424 =  x_2157 & ~n_33423;
assign n_33425 = ~x_2157 &  n_33423;
assign n_33426 = ~n_33424 & ~n_33425;
assign n_33427 =  x_2156 & ~n_33186;
assign n_33428 =  x_3225 &  n_27721;
assign n_33429 =  x_4905 &  n_558;
assign n_33430 = ~n_33428 & ~n_33429;
assign n_33431 = ~n_33427 &  n_33430;
assign n_33432 =  x_2156 & ~n_33431;
assign n_33433 = ~x_2156 &  n_33431;
assign n_33434 = ~n_33432 & ~n_33433;
assign n_33435 =  x_2155 & ~n_33186;
assign n_33436 =  x_4904 &  n_558;
assign n_33437 =  x_3224 &  n_27721;
assign n_33438 = ~n_33436 & ~n_33437;
assign n_33439 = ~n_33435 &  n_33438;
assign n_33440 =  x_2155 & ~n_33439;
assign n_33441 = ~x_2155 &  n_33439;
assign n_33442 = ~n_33440 & ~n_33441;
assign n_33443 = ~n_26100 & ~n_27016;
assign n_33444 = ~n_23812 &  n_33443;
assign n_33445 = ~n_26190 &  n_33444;
assign n_33446 =  x_2154 &  n_33445;
assign n_33447 =  x_2090 &  n_26190;
assign n_33448 =  x_555 &  n_23812;
assign n_33449 =  x_747 &  n_26100;
assign n_33450 =  x_1930 &  n_27016;
assign n_33451 = ~n_33449 & ~n_33450;
assign n_33452 = ~n_33448 &  n_33451;
assign n_33453 = ~n_33447 &  n_33452;
assign n_33454 = ~n_33446 &  n_33453;
assign n_33455 =  x_2154 & ~n_33454;
assign n_33456 = ~x_2154 &  n_33454;
assign n_33457 = ~n_33455 & ~n_33456;
assign n_33458 =  x_2153 &  n_33445;
assign n_33459 =  x_2089 &  n_26190;
assign n_33460 =  x_554 &  n_23812;
assign n_33461 =  x_746 &  n_26100;
assign n_33462 =  x_1929 &  n_27016;
assign n_33463 = ~n_33461 & ~n_33462;
assign n_33464 = ~n_33460 &  n_33463;
assign n_33465 = ~n_33459 &  n_33464;
assign n_33466 = ~n_33458 &  n_33465;
assign n_33467 =  x_2153 & ~n_33466;
assign n_33468 = ~x_2153 &  n_33466;
assign n_33469 = ~n_33467 & ~n_33468;
assign n_33470 =  x_2152 &  n_33445;
assign n_33471 =  x_2088 &  n_26190;
assign n_33472 =  x_553 &  n_23812;
assign n_33473 =  x_745 &  n_26100;
assign n_33474 =  x_1928 &  n_27016;
assign n_33475 = ~n_33473 & ~n_33474;
assign n_33476 = ~n_33472 &  n_33475;
assign n_33477 = ~n_33471 &  n_33476;
assign n_33478 = ~n_33470 &  n_33477;
assign n_33479 =  x_2152 & ~n_33478;
assign n_33480 = ~x_2152 &  n_33478;
assign n_33481 = ~n_33479 & ~n_33480;
assign n_33482 =  x_2151 &  n_33445;
assign n_33483 =  x_2087 &  n_26190;
assign n_33484 =  x_552 &  n_23812;
assign n_33485 =  x_744 &  n_26100;
assign n_33486 =  x_1927 &  n_27016;
assign n_33487 = ~n_33485 & ~n_33486;
assign n_33488 = ~n_33484 &  n_33487;
assign n_33489 = ~n_33483 &  n_33488;
assign n_33490 = ~n_33482 &  n_33489;
assign n_33491 =  x_2151 & ~n_33490;
assign n_33492 = ~x_2151 &  n_33490;
assign n_33493 = ~n_33491 & ~n_33492;
assign n_33494 =  x_2150 &  n_33445;
assign n_33495 =  x_2086 &  n_26190;
assign n_33496 =  x_551 &  n_23812;
assign n_33497 =  x_743 &  n_26100;
assign n_33498 =  x_1926 &  n_27016;
assign n_33499 = ~n_33497 & ~n_33498;
assign n_33500 = ~n_33496 &  n_33499;
assign n_33501 = ~n_33495 &  n_33500;
assign n_33502 = ~n_33494 &  n_33501;
assign n_33503 =  x_2150 & ~n_33502;
assign n_33504 = ~x_2150 &  n_33502;
assign n_33505 = ~n_33503 & ~n_33504;
assign n_33506 =  x_2149 &  n_33445;
assign n_33507 =  x_2085 &  n_26190;
assign n_33508 =  x_550 &  n_23812;
assign n_33509 =  x_742 &  n_26100;
assign n_33510 =  x_1925 &  n_27016;
assign n_33511 = ~n_33509 & ~n_33510;
assign n_33512 = ~n_33508 &  n_33511;
assign n_33513 = ~n_33507 &  n_33512;
assign n_33514 = ~n_33506 &  n_33513;
assign n_33515 =  x_2149 & ~n_33514;
assign n_33516 = ~x_2149 &  n_33514;
assign n_33517 = ~n_33515 & ~n_33516;
assign n_33518 =  x_2148 &  n_33445;
assign n_33519 =  x_2084 &  n_26190;
assign n_33520 =  x_549 &  n_23812;
assign n_33521 =  x_741 &  n_26100;
assign n_33522 =  x_1924 &  n_27016;
assign n_33523 = ~n_33521 & ~n_33522;
assign n_33524 = ~n_33520 &  n_33523;
assign n_33525 = ~n_33519 &  n_33524;
assign n_33526 = ~n_33518 &  n_33525;
assign n_33527 =  x_2148 & ~n_33526;
assign n_33528 = ~x_2148 &  n_33526;
assign n_33529 = ~n_33527 & ~n_33528;
assign n_33530 =  x_2147 &  n_33445;
assign n_33531 =  x_2083 &  n_26190;
assign n_33532 =  x_548 &  n_23812;
assign n_33533 =  x_740 &  n_26100;
assign n_33534 =  x_1923 &  n_27016;
assign n_33535 = ~n_33533 & ~n_33534;
assign n_33536 = ~n_33532 &  n_33535;
assign n_33537 = ~n_33531 &  n_33536;
assign n_33538 = ~n_33530 &  n_33537;
assign n_33539 =  x_2147 & ~n_33538;
assign n_33540 = ~x_2147 &  n_33538;
assign n_33541 = ~n_33539 & ~n_33540;
assign n_33542 =  x_2146 &  n_33445;
assign n_33543 =  x_2082 &  n_26190;
assign n_33544 =  x_547 &  n_23812;
assign n_33545 =  x_739 &  n_26100;
assign n_33546 =  x_1922 &  n_27016;
assign n_33547 = ~n_33545 & ~n_33546;
assign n_33548 = ~n_33544 &  n_33547;
assign n_33549 = ~n_33543 &  n_33548;
assign n_33550 = ~n_33542 &  n_33549;
assign n_33551 =  x_2146 & ~n_33550;
assign n_33552 = ~x_2146 &  n_33550;
assign n_33553 = ~n_33551 & ~n_33552;
assign n_33554 =  x_2145 &  n_33445;
assign n_33555 =  x_2081 &  n_26190;
assign n_33556 =  x_546 &  n_23812;
assign n_33557 =  x_738 &  n_26100;
assign n_33558 =  x_1921 &  n_27016;
assign n_33559 = ~n_33557 & ~n_33558;
assign n_33560 = ~n_33556 &  n_33559;
assign n_33561 = ~n_33555 &  n_33560;
assign n_33562 = ~n_33554 &  n_33561;
assign n_33563 =  x_2145 & ~n_33562;
assign n_33564 = ~x_2145 &  n_33562;
assign n_33565 = ~n_33563 & ~n_33564;
assign n_33566 =  x_2144 &  n_33445;
assign n_33567 =  x_2080 &  n_26190;
assign n_33568 =  x_545 &  n_23812;
assign n_33569 =  x_737 &  n_26100;
assign n_33570 =  x_1920 &  n_27016;
assign n_33571 = ~n_33569 & ~n_33570;
assign n_33572 = ~n_33568 &  n_33571;
assign n_33573 = ~n_33567 &  n_33572;
assign n_33574 = ~n_33566 &  n_33573;
assign n_33575 =  x_2144 & ~n_33574;
assign n_33576 = ~x_2144 &  n_33574;
assign n_33577 = ~n_33575 & ~n_33576;
assign n_33578 =  x_2143 &  n_33445;
assign n_33579 =  x_2079 &  n_26190;
assign n_33580 =  x_544 &  n_23812;
assign n_33581 =  x_736 &  n_26100;
assign n_33582 =  x_1919 &  n_27016;
assign n_33583 = ~n_33581 & ~n_33582;
assign n_33584 = ~n_33580 &  n_33583;
assign n_33585 = ~n_33579 &  n_33584;
assign n_33586 = ~n_33578 &  n_33585;
assign n_33587 =  x_2143 & ~n_33586;
assign n_33588 = ~x_2143 &  n_33586;
assign n_33589 = ~n_33587 & ~n_33588;
assign n_33590 =  x_2142 &  n_33445;
assign n_33591 =  x_2078 &  n_26190;
assign n_33592 =  x_543 &  n_23812;
assign n_33593 =  x_735 &  n_26100;
assign n_33594 =  x_1918 &  n_27016;
assign n_33595 = ~n_33593 & ~n_33594;
assign n_33596 = ~n_33592 &  n_33595;
assign n_33597 = ~n_33591 &  n_33596;
assign n_33598 = ~n_33590 &  n_33597;
assign n_33599 =  x_2142 & ~n_33598;
assign n_33600 = ~x_2142 &  n_33598;
assign n_33601 = ~n_33599 & ~n_33600;
assign n_33602 =  x_2141 &  n_33445;
assign n_33603 =  x_2077 &  n_26190;
assign n_33604 =  x_542 &  n_23812;
assign n_33605 =  x_734 &  n_26100;
assign n_33606 =  x_1917 &  n_27016;
assign n_33607 = ~n_33605 & ~n_33606;
assign n_33608 = ~n_33604 &  n_33607;
assign n_33609 = ~n_33603 &  n_33608;
assign n_33610 = ~n_33602 &  n_33609;
assign n_33611 =  x_2141 & ~n_33610;
assign n_33612 = ~x_2141 &  n_33610;
assign n_33613 = ~n_33611 & ~n_33612;
assign n_33614 =  x_2140 &  n_33445;
assign n_33615 =  x_2076 &  n_26190;
assign n_33616 =  x_541 &  n_23812;
assign n_33617 =  x_733 &  n_26100;
assign n_33618 =  x_1916 &  n_27016;
assign n_33619 = ~n_33617 & ~n_33618;
assign n_33620 = ~n_33616 &  n_33619;
assign n_33621 = ~n_33615 &  n_33620;
assign n_33622 = ~n_33614 &  n_33621;
assign n_33623 =  x_2140 & ~n_33622;
assign n_33624 = ~x_2140 &  n_33622;
assign n_33625 = ~n_33623 & ~n_33624;
assign n_33626 =  x_2139 &  n_33445;
assign n_33627 =  x_2075 &  n_26190;
assign n_33628 =  x_540 &  n_23812;
assign n_33629 =  x_732 &  n_26100;
assign n_33630 =  x_1915 &  n_27016;
assign n_33631 = ~n_33629 & ~n_33630;
assign n_33632 = ~n_33628 &  n_33631;
assign n_33633 = ~n_33627 &  n_33632;
assign n_33634 = ~n_33626 &  n_33633;
assign n_33635 =  x_2139 & ~n_33634;
assign n_33636 = ~x_2139 &  n_33634;
assign n_33637 = ~n_33635 & ~n_33636;
assign n_33638 =  x_2138 &  n_33445;
assign n_33639 =  x_2074 &  n_26190;
assign n_33640 =  x_539 &  n_23812;
assign n_33641 =  x_731 &  n_26100;
assign n_33642 =  x_1914 &  n_27016;
assign n_33643 = ~n_33641 & ~n_33642;
assign n_33644 = ~n_33640 &  n_33643;
assign n_33645 = ~n_33639 &  n_33644;
assign n_33646 = ~n_33638 &  n_33645;
assign n_33647 =  x_2138 & ~n_33646;
assign n_33648 = ~x_2138 &  n_33646;
assign n_33649 = ~n_33647 & ~n_33648;
assign n_33650 =  x_2137 &  n_33445;
assign n_33651 =  x_2073 &  n_26190;
assign n_33652 =  x_538 &  n_23812;
assign n_33653 =  x_730 &  n_26100;
assign n_33654 =  x_1913 &  n_27016;
assign n_33655 = ~n_33653 & ~n_33654;
assign n_33656 = ~n_33652 &  n_33655;
assign n_33657 = ~n_33651 &  n_33656;
assign n_33658 = ~n_33650 &  n_33657;
assign n_33659 =  x_2137 & ~n_33658;
assign n_33660 = ~x_2137 &  n_33658;
assign n_33661 = ~n_33659 & ~n_33660;
assign n_33662 =  x_2136 &  n_33445;
assign n_33663 =  x_2072 &  n_26190;
assign n_33664 =  x_537 &  n_23812;
assign n_33665 =  x_729 &  n_26100;
assign n_33666 =  x_1912 &  n_27016;
assign n_33667 = ~n_33665 & ~n_33666;
assign n_33668 = ~n_33664 &  n_33667;
assign n_33669 = ~n_33663 &  n_33668;
assign n_33670 = ~n_33662 &  n_33669;
assign n_33671 =  x_2136 & ~n_33670;
assign n_33672 = ~x_2136 &  n_33670;
assign n_33673 = ~n_33671 & ~n_33672;
assign n_33674 =  x_2135 &  n_33445;
assign n_33675 =  x_2071 &  n_26190;
assign n_33676 =  x_536 &  n_23812;
assign n_33677 =  x_728 &  n_26100;
assign n_33678 =  x_1911 &  n_27016;
assign n_33679 = ~n_33677 & ~n_33678;
assign n_33680 = ~n_33676 &  n_33679;
assign n_33681 = ~n_33675 &  n_33680;
assign n_33682 = ~n_33674 &  n_33681;
assign n_33683 =  x_2135 & ~n_33682;
assign n_33684 = ~x_2135 &  n_33682;
assign n_33685 = ~n_33683 & ~n_33684;
assign n_33686 =  x_2134 &  n_33445;
assign n_33687 =  x_2070 &  n_26190;
assign n_33688 =  x_535 &  n_23812;
assign n_33689 =  x_727 &  n_26100;
assign n_33690 =  x_1910 &  n_27016;
assign n_33691 = ~n_33689 & ~n_33690;
assign n_33692 = ~n_33688 &  n_33691;
assign n_33693 = ~n_33687 &  n_33692;
assign n_33694 = ~n_33686 &  n_33693;
assign n_33695 =  x_2134 & ~n_33694;
assign n_33696 = ~x_2134 &  n_33694;
assign n_33697 = ~n_33695 & ~n_33696;
assign n_33698 =  x_2133 &  n_33445;
assign n_33699 =  x_2069 &  n_26190;
assign n_33700 =  x_534 &  n_23812;
assign n_33701 =  x_726 &  n_26100;
assign n_33702 =  x_1909 &  n_27016;
assign n_33703 = ~n_33701 & ~n_33702;
assign n_33704 = ~n_33700 &  n_33703;
assign n_33705 = ~n_33699 &  n_33704;
assign n_33706 = ~n_33698 &  n_33705;
assign n_33707 =  x_2133 & ~n_33706;
assign n_33708 = ~x_2133 &  n_33706;
assign n_33709 = ~n_33707 & ~n_33708;
assign n_33710 =  x_2132 &  n_33445;
assign n_33711 =  x_2068 &  n_26190;
assign n_33712 =  x_533 &  n_23812;
assign n_33713 =  x_725 &  n_26100;
assign n_33714 =  x_1908 &  n_27016;
assign n_33715 = ~n_33713 & ~n_33714;
assign n_33716 = ~n_33712 &  n_33715;
assign n_33717 = ~n_33711 &  n_33716;
assign n_33718 = ~n_33710 &  n_33717;
assign n_33719 =  x_2132 & ~n_33718;
assign n_33720 = ~x_2132 &  n_33718;
assign n_33721 = ~n_33719 & ~n_33720;
assign n_33722 =  x_2131 &  n_33445;
assign n_33723 =  x_2067 &  n_26190;
assign n_33724 =  x_532 &  n_23812;
assign n_33725 =  x_724 &  n_26100;
assign n_33726 =  x_1907 &  n_27016;
assign n_33727 = ~n_33725 & ~n_33726;
assign n_33728 = ~n_33724 &  n_33727;
assign n_33729 = ~n_33723 &  n_33728;
assign n_33730 = ~n_33722 &  n_33729;
assign n_33731 =  x_2131 & ~n_33730;
assign n_33732 = ~x_2131 &  n_33730;
assign n_33733 = ~n_33731 & ~n_33732;
assign n_33734 =  x_2130 &  n_33445;
assign n_33735 =  x_2066 &  n_26190;
assign n_33736 =  x_531 &  n_23812;
assign n_33737 =  x_723 &  n_26100;
assign n_33738 =  x_1906 &  n_27016;
assign n_33739 = ~n_33737 & ~n_33738;
assign n_33740 = ~n_33736 &  n_33739;
assign n_33741 = ~n_33735 &  n_33740;
assign n_33742 = ~n_33734 &  n_33741;
assign n_33743 =  x_2130 & ~n_33742;
assign n_33744 = ~x_2130 &  n_33742;
assign n_33745 = ~n_33743 & ~n_33744;
assign n_33746 =  x_2129 &  n_33445;
assign n_33747 =  x_2065 &  n_26190;
assign n_33748 =  x_530 &  n_23812;
assign n_33749 =  x_722 &  n_26100;
assign n_33750 =  x_1905 &  n_27016;
assign n_33751 = ~n_33749 & ~n_33750;
assign n_33752 = ~n_33748 &  n_33751;
assign n_33753 = ~n_33747 &  n_33752;
assign n_33754 = ~n_33746 &  n_33753;
assign n_33755 =  x_2129 & ~n_33754;
assign n_33756 = ~x_2129 &  n_33754;
assign n_33757 = ~n_33755 & ~n_33756;
assign n_33758 =  x_2128 &  n_33445;
assign n_33759 =  x_2064 &  n_26190;
assign n_33760 =  x_529 &  n_23812;
assign n_33761 =  x_721 &  n_26100;
assign n_33762 =  x_1904 &  n_27016;
assign n_33763 = ~n_33761 & ~n_33762;
assign n_33764 = ~n_33760 &  n_33763;
assign n_33765 = ~n_33759 &  n_33764;
assign n_33766 = ~n_33758 &  n_33765;
assign n_33767 =  x_2128 & ~n_33766;
assign n_33768 = ~x_2128 &  n_33766;
assign n_33769 = ~n_33767 & ~n_33768;
assign n_33770 =  x_2127 &  n_33445;
assign n_33771 =  x_2063 &  n_26190;
assign n_33772 =  x_528 &  n_23812;
assign n_33773 =  x_720 &  n_26100;
assign n_33774 =  x_1903 &  n_27016;
assign n_33775 = ~n_33773 & ~n_33774;
assign n_33776 = ~n_33772 &  n_33775;
assign n_33777 = ~n_33771 &  n_33776;
assign n_33778 = ~n_33770 &  n_33777;
assign n_33779 =  x_2127 & ~n_33778;
assign n_33780 = ~x_2127 &  n_33778;
assign n_33781 = ~n_33779 & ~n_33780;
assign n_33782 =  x_2126 &  n_33445;
assign n_33783 =  x_2062 &  n_26190;
assign n_33784 =  x_527 &  n_23812;
assign n_33785 =  x_719 &  n_26100;
assign n_33786 =  x_1902 &  n_27016;
assign n_33787 = ~n_33785 & ~n_33786;
assign n_33788 = ~n_33784 &  n_33787;
assign n_33789 = ~n_33783 &  n_33788;
assign n_33790 = ~n_33782 &  n_33789;
assign n_33791 =  x_2126 & ~n_33790;
assign n_33792 = ~x_2126 &  n_33790;
assign n_33793 = ~n_33791 & ~n_33792;
assign n_33794 =  x_2125 &  n_33445;
assign n_33795 =  x_2061 &  n_26190;
assign n_33796 =  x_526 &  n_23812;
assign n_33797 =  x_718 &  n_26100;
assign n_33798 =  x_1901 &  n_27016;
assign n_33799 = ~n_33797 & ~n_33798;
assign n_33800 = ~n_33796 &  n_33799;
assign n_33801 = ~n_33795 &  n_33800;
assign n_33802 = ~n_33794 &  n_33801;
assign n_33803 =  x_2125 & ~n_33802;
assign n_33804 = ~x_2125 &  n_33802;
assign n_33805 = ~n_33803 & ~n_33804;
assign n_33806 =  x_2124 &  n_33445;
assign n_33807 =  x_2060 &  n_26190;
assign n_33808 =  x_525 &  n_23812;
assign n_33809 =  x_717 &  n_26100;
assign n_33810 =  x_1900 &  n_27016;
assign n_33811 = ~n_33809 & ~n_33810;
assign n_33812 = ~n_33808 &  n_33811;
assign n_33813 = ~n_33807 &  n_33812;
assign n_33814 = ~n_33806 &  n_33813;
assign n_33815 =  x_2124 & ~n_33814;
assign n_33816 = ~x_2124 &  n_33814;
assign n_33817 = ~n_33815 & ~n_33816;
assign n_33818 =  x_2123 &  n_33445;
assign n_33819 =  x_2059 &  n_26190;
assign n_33820 =  x_524 &  n_23812;
assign n_33821 =  x_716 &  n_26100;
assign n_33822 =  x_1899 &  n_27016;
assign n_33823 = ~n_33821 & ~n_33822;
assign n_33824 = ~n_33820 &  n_33823;
assign n_33825 = ~n_33819 &  n_33824;
assign n_33826 = ~n_33818 &  n_33825;
assign n_33827 =  x_2123 & ~n_33826;
assign n_33828 = ~x_2123 &  n_33826;
assign n_33829 = ~n_33827 & ~n_33828;
assign n_33830 =  x_2122 & ~n_26411;
assign n_33831 =  i_32 &  n_26411;
assign n_33832 = ~n_33830 & ~n_33831;
assign n_33833 =  x_2122 & ~n_33832;
assign n_33834 = ~x_2122 &  n_33832;
assign n_33835 = ~n_33833 & ~n_33834;
assign n_33836 =  x_2121 & ~n_26411;
assign n_33837 =  i_31 &  n_26411;
assign n_33838 = ~n_33836 & ~n_33837;
assign n_33839 =  x_2121 & ~n_33838;
assign n_33840 = ~x_2121 &  n_33838;
assign n_33841 = ~n_33839 & ~n_33840;
assign n_33842 =  x_2120 & ~n_26411;
assign n_33843 =  i_30 &  n_26411;
assign n_33844 = ~n_33842 & ~n_33843;
assign n_33845 =  x_2120 & ~n_33844;
assign n_33846 = ~x_2120 &  n_33844;
assign n_33847 = ~n_33845 & ~n_33846;
assign n_33848 =  x_2119 & ~n_26411;
assign n_33849 =  i_29 &  n_26411;
assign n_33850 = ~n_33848 & ~n_33849;
assign n_33851 =  x_2119 & ~n_33850;
assign n_33852 = ~x_2119 &  n_33850;
assign n_33853 = ~n_33851 & ~n_33852;
assign n_33854 =  x_2118 & ~n_26411;
assign n_33855 =  i_28 &  n_26411;
assign n_33856 = ~n_33854 & ~n_33855;
assign n_33857 =  x_2118 & ~n_33856;
assign n_33858 = ~x_2118 &  n_33856;
assign n_33859 = ~n_33857 & ~n_33858;
assign n_33860 =  x_2117 & ~n_26411;
assign n_33861 =  i_27 &  n_26411;
assign n_33862 = ~n_33860 & ~n_33861;
assign n_33863 =  x_2117 & ~n_33862;
assign n_33864 = ~x_2117 &  n_33862;
assign n_33865 = ~n_33863 & ~n_33864;
assign n_33866 =  x_2116 & ~n_26411;
assign n_33867 =  i_26 &  n_26411;
assign n_33868 = ~n_33866 & ~n_33867;
assign n_33869 =  x_2116 & ~n_33868;
assign n_33870 = ~x_2116 &  n_33868;
assign n_33871 = ~n_33869 & ~n_33870;
assign n_33872 =  x_2115 & ~n_26411;
assign n_33873 =  i_25 &  n_26411;
assign n_33874 = ~n_33872 & ~n_33873;
assign n_33875 =  x_2115 & ~n_33874;
assign n_33876 = ~x_2115 &  n_33874;
assign n_33877 = ~n_33875 & ~n_33876;
assign n_33878 =  x_2114 & ~n_26411;
assign n_33879 =  i_24 &  n_26411;
assign n_33880 = ~n_33878 & ~n_33879;
assign n_33881 =  x_2114 & ~n_33880;
assign n_33882 = ~x_2114 &  n_33880;
assign n_33883 = ~n_33881 & ~n_33882;
assign n_33884 =  x_2113 & ~n_26411;
assign n_33885 =  i_23 &  n_26411;
assign n_33886 = ~n_33884 & ~n_33885;
assign n_33887 =  x_2113 & ~n_33886;
assign n_33888 = ~x_2113 &  n_33886;
assign n_33889 = ~n_33887 & ~n_33888;
assign n_33890 =  x_2112 & ~n_26411;
assign n_33891 =  i_22 &  n_26411;
assign n_33892 = ~n_33890 & ~n_33891;
assign n_33893 =  x_2112 & ~n_33892;
assign n_33894 = ~x_2112 &  n_33892;
assign n_33895 = ~n_33893 & ~n_33894;
assign n_33896 =  x_2111 & ~n_26411;
assign n_33897 =  i_21 &  n_26411;
assign n_33898 = ~n_33896 & ~n_33897;
assign n_33899 =  x_2111 & ~n_33898;
assign n_33900 = ~x_2111 &  n_33898;
assign n_33901 = ~n_33899 & ~n_33900;
assign n_33902 =  x_2110 & ~n_26411;
assign n_33903 =  i_20 &  n_26411;
assign n_33904 = ~n_33902 & ~n_33903;
assign n_33905 =  x_2110 & ~n_33904;
assign n_33906 = ~x_2110 &  n_33904;
assign n_33907 = ~n_33905 & ~n_33906;
assign n_33908 =  x_2109 & ~n_26411;
assign n_33909 =  i_19 &  n_26411;
assign n_33910 = ~n_33908 & ~n_33909;
assign n_33911 =  x_2109 & ~n_33910;
assign n_33912 = ~x_2109 &  n_33910;
assign n_33913 = ~n_33911 & ~n_33912;
assign n_33914 =  x_2108 & ~n_26411;
assign n_33915 =  i_18 &  n_26411;
assign n_33916 = ~n_33914 & ~n_33915;
assign n_33917 =  x_2108 & ~n_33916;
assign n_33918 = ~x_2108 &  n_33916;
assign n_33919 = ~n_33917 & ~n_33918;
assign n_33920 =  x_2107 & ~n_26411;
assign n_33921 =  i_17 &  n_26411;
assign n_33922 = ~n_33920 & ~n_33921;
assign n_33923 =  x_2107 & ~n_33922;
assign n_33924 = ~x_2107 &  n_33922;
assign n_33925 = ~n_33923 & ~n_33924;
assign n_33926 =  x_2106 & ~n_26411;
assign n_33927 =  i_16 &  n_26411;
assign n_33928 = ~n_33926 & ~n_33927;
assign n_33929 =  x_2106 & ~n_33928;
assign n_33930 = ~x_2106 &  n_33928;
assign n_33931 = ~n_33929 & ~n_33930;
assign n_33932 =  x_2105 & ~n_26411;
assign n_33933 =  i_15 &  n_26411;
assign n_33934 = ~n_33932 & ~n_33933;
assign n_33935 =  x_2105 & ~n_33934;
assign n_33936 = ~x_2105 &  n_33934;
assign n_33937 = ~n_33935 & ~n_33936;
assign n_33938 =  x_2104 & ~n_26411;
assign n_33939 =  i_14 &  n_26411;
assign n_33940 = ~n_33938 & ~n_33939;
assign n_33941 =  x_2104 & ~n_33940;
assign n_33942 = ~x_2104 &  n_33940;
assign n_33943 = ~n_33941 & ~n_33942;
assign n_33944 =  x_2103 & ~n_26411;
assign n_33945 =  i_13 &  n_26411;
assign n_33946 = ~n_33944 & ~n_33945;
assign n_33947 =  x_2103 & ~n_33946;
assign n_33948 = ~x_2103 &  n_33946;
assign n_33949 = ~n_33947 & ~n_33948;
assign n_33950 =  x_2102 & ~n_26411;
assign n_33951 =  i_12 &  n_26411;
assign n_33952 = ~n_33950 & ~n_33951;
assign n_33953 =  x_2102 & ~n_33952;
assign n_33954 = ~x_2102 &  n_33952;
assign n_33955 = ~n_33953 & ~n_33954;
assign n_33956 =  x_2101 & ~n_26411;
assign n_33957 =  i_11 &  n_26411;
assign n_33958 = ~n_33956 & ~n_33957;
assign n_33959 =  x_2101 & ~n_33958;
assign n_33960 = ~x_2101 &  n_33958;
assign n_33961 = ~n_33959 & ~n_33960;
assign n_33962 =  x_2100 & ~n_26411;
assign n_33963 =  i_10 &  n_26411;
assign n_33964 = ~n_33962 & ~n_33963;
assign n_33965 =  x_2100 & ~n_33964;
assign n_33966 = ~x_2100 &  n_33964;
assign n_33967 = ~n_33965 & ~n_33966;
assign n_33968 =  x_2099 & ~n_26411;
assign n_33969 =  i_9 &  n_26411;
assign n_33970 = ~n_33968 & ~n_33969;
assign n_33971 =  x_2099 & ~n_33970;
assign n_33972 = ~x_2099 &  n_33970;
assign n_33973 = ~n_33971 & ~n_33972;
assign n_33974 =  x_2098 & ~n_26411;
assign n_33975 =  i_8 &  n_26411;
assign n_33976 = ~n_33974 & ~n_33975;
assign n_33977 =  x_2098 & ~n_33976;
assign n_33978 = ~x_2098 &  n_33976;
assign n_33979 = ~n_33977 & ~n_33978;
assign n_33980 =  x_2097 & ~n_26411;
assign n_33981 =  i_7 &  n_26411;
assign n_33982 = ~n_33980 & ~n_33981;
assign n_33983 =  x_2097 & ~n_33982;
assign n_33984 = ~x_2097 &  n_33982;
assign n_33985 = ~n_33983 & ~n_33984;
assign n_33986 =  x_2096 & ~n_26411;
assign n_33987 =  i_6 &  n_26411;
assign n_33988 = ~n_33986 & ~n_33987;
assign n_33989 =  x_2096 & ~n_33988;
assign n_33990 = ~x_2096 &  n_33988;
assign n_33991 = ~n_33989 & ~n_33990;
assign n_33992 =  x_2095 & ~n_26411;
assign n_33993 =  i_5 &  n_26411;
assign n_33994 = ~n_33992 & ~n_33993;
assign n_33995 =  x_2095 & ~n_33994;
assign n_33996 = ~x_2095 &  n_33994;
assign n_33997 = ~n_33995 & ~n_33996;
assign n_33998 =  x_2094 & ~n_26411;
assign n_33999 =  i_4 &  n_26411;
assign n_34000 = ~n_33998 & ~n_33999;
assign n_34001 =  x_2094 & ~n_34000;
assign n_34002 = ~x_2094 &  n_34000;
assign n_34003 = ~n_34001 & ~n_34002;
assign n_34004 =  x_2093 & ~n_26411;
assign n_34005 =  i_3 &  n_26411;
assign n_34006 = ~n_34004 & ~n_34005;
assign n_34007 =  x_2093 & ~n_34006;
assign n_34008 = ~x_2093 &  n_34006;
assign n_34009 = ~n_34007 & ~n_34008;
assign n_34010 =  x_2092 & ~n_26411;
assign n_34011 =  i_2 &  n_26411;
assign n_34012 = ~n_34010 & ~n_34011;
assign n_34013 =  x_2092 & ~n_34012;
assign n_34014 = ~x_2092 &  n_34012;
assign n_34015 = ~n_34013 & ~n_34014;
assign n_34016 =  x_2091 & ~n_26411;
assign n_34017 =  i_1 &  n_26411;
assign n_34018 = ~n_34016 & ~n_34017;
assign n_34019 =  x_2091 & ~n_34018;
assign n_34020 = ~x_2091 &  n_34018;
assign n_34021 = ~n_34019 & ~n_34020;
assign n_34022 =  x_2090 & ~n_24504;
assign n_34023 =  i_32 &  n_24504;
assign n_34024 = ~n_34022 & ~n_34023;
assign n_34025 =  x_2090 & ~n_34024;
assign n_34026 = ~x_2090 &  n_34024;
assign n_34027 = ~n_34025 & ~n_34026;
assign n_34028 =  x_2089 & ~n_24504;
assign n_34029 =  i_31 &  n_24504;
assign n_34030 = ~n_34028 & ~n_34029;
assign n_34031 =  x_2089 & ~n_34030;
assign n_34032 = ~x_2089 &  n_34030;
assign n_34033 = ~n_34031 & ~n_34032;
assign n_34034 =  x_2088 & ~n_24504;
assign n_34035 =  i_30 &  n_24504;
assign n_34036 = ~n_34034 & ~n_34035;
assign n_34037 =  x_2088 & ~n_34036;
assign n_34038 = ~x_2088 &  n_34036;
assign n_34039 = ~n_34037 & ~n_34038;
assign n_34040 =  x_2087 & ~n_24504;
assign n_34041 =  i_29 &  n_24504;
assign n_34042 = ~n_34040 & ~n_34041;
assign n_34043 =  x_2087 & ~n_34042;
assign n_34044 = ~x_2087 &  n_34042;
assign n_34045 = ~n_34043 & ~n_34044;
assign n_34046 =  x_2086 & ~n_24504;
assign n_34047 =  i_28 &  n_24504;
assign n_34048 = ~n_34046 & ~n_34047;
assign n_34049 =  x_2086 & ~n_34048;
assign n_34050 = ~x_2086 &  n_34048;
assign n_34051 = ~n_34049 & ~n_34050;
assign n_34052 =  x_2085 & ~n_24504;
assign n_34053 =  i_27 &  n_24504;
assign n_34054 = ~n_34052 & ~n_34053;
assign n_34055 =  x_2085 & ~n_34054;
assign n_34056 = ~x_2085 &  n_34054;
assign n_34057 = ~n_34055 & ~n_34056;
assign n_34058 =  x_2084 & ~n_24504;
assign n_34059 =  i_26 &  n_24504;
assign n_34060 = ~n_34058 & ~n_34059;
assign n_34061 =  x_2084 & ~n_34060;
assign n_34062 = ~x_2084 &  n_34060;
assign n_34063 = ~n_34061 & ~n_34062;
assign n_34064 =  x_2083 & ~n_24504;
assign n_34065 =  i_25 &  n_24504;
assign n_34066 = ~n_34064 & ~n_34065;
assign n_34067 =  x_2083 & ~n_34066;
assign n_34068 = ~x_2083 &  n_34066;
assign n_34069 = ~n_34067 & ~n_34068;
assign n_34070 =  x_2082 & ~n_24504;
assign n_34071 =  i_24 &  n_24504;
assign n_34072 = ~n_34070 & ~n_34071;
assign n_34073 =  x_2082 & ~n_34072;
assign n_34074 = ~x_2082 &  n_34072;
assign n_34075 = ~n_34073 & ~n_34074;
assign n_34076 =  x_2081 & ~n_24504;
assign n_34077 =  i_23 &  n_24504;
assign n_34078 = ~n_34076 & ~n_34077;
assign n_34079 =  x_2081 & ~n_34078;
assign n_34080 = ~x_2081 &  n_34078;
assign n_34081 = ~n_34079 & ~n_34080;
assign n_34082 =  x_2080 & ~n_24504;
assign n_34083 =  i_22 &  n_24504;
assign n_34084 = ~n_34082 & ~n_34083;
assign n_34085 =  x_2080 & ~n_34084;
assign n_34086 = ~x_2080 &  n_34084;
assign n_34087 = ~n_34085 & ~n_34086;
assign n_34088 =  x_2079 & ~n_24504;
assign n_34089 =  i_21 &  n_24504;
assign n_34090 = ~n_34088 & ~n_34089;
assign n_34091 =  x_2079 & ~n_34090;
assign n_34092 = ~x_2079 &  n_34090;
assign n_34093 = ~n_34091 & ~n_34092;
assign n_34094 =  x_2078 & ~n_24504;
assign n_34095 =  i_20 &  n_24504;
assign n_34096 = ~n_34094 & ~n_34095;
assign n_34097 =  x_2078 & ~n_34096;
assign n_34098 = ~x_2078 &  n_34096;
assign n_34099 = ~n_34097 & ~n_34098;
assign n_34100 =  x_2077 & ~n_24504;
assign n_34101 =  i_19 &  n_24504;
assign n_34102 = ~n_34100 & ~n_34101;
assign n_34103 =  x_2077 & ~n_34102;
assign n_34104 = ~x_2077 &  n_34102;
assign n_34105 = ~n_34103 & ~n_34104;
assign n_34106 =  x_2076 & ~n_24504;
assign n_34107 =  i_18 &  n_24504;
assign n_34108 = ~n_34106 & ~n_34107;
assign n_34109 =  x_2076 & ~n_34108;
assign n_34110 = ~x_2076 &  n_34108;
assign n_34111 = ~n_34109 & ~n_34110;
assign n_34112 =  x_2075 & ~n_24504;
assign n_34113 =  i_17 &  n_24504;
assign n_34114 = ~n_34112 & ~n_34113;
assign n_34115 =  x_2075 & ~n_34114;
assign n_34116 = ~x_2075 &  n_34114;
assign n_34117 = ~n_34115 & ~n_34116;
assign n_34118 =  x_2074 & ~n_24504;
assign n_34119 =  i_16 &  n_24504;
assign n_34120 = ~n_34118 & ~n_34119;
assign n_34121 =  x_2074 & ~n_34120;
assign n_34122 = ~x_2074 &  n_34120;
assign n_34123 = ~n_34121 & ~n_34122;
assign n_34124 =  x_2073 & ~n_24504;
assign n_34125 =  i_15 &  n_24504;
assign n_34126 = ~n_34124 & ~n_34125;
assign n_34127 =  x_2073 & ~n_34126;
assign n_34128 = ~x_2073 &  n_34126;
assign n_34129 = ~n_34127 & ~n_34128;
assign n_34130 =  x_2072 & ~n_24504;
assign n_34131 =  i_14 &  n_24504;
assign n_34132 = ~n_34130 & ~n_34131;
assign n_34133 =  x_2072 & ~n_34132;
assign n_34134 = ~x_2072 &  n_34132;
assign n_34135 = ~n_34133 & ~n_34134;
assign n_34136 =  x_2071 & ~n_24504;
assign n_34137 =  i_13 &  n_24504;
assign n_34138 = ~n_34136 & ~n_34137;
assign n_34139 =  x_2071 & ~n_34138;
assign n_34140 = ~x_2071 &  n_34138;
assign n_34141 = ~n_34139 & ~n_34140;
assign n_34142 =  x_2070 & ~n_24504;
assign n_34143 =  i_12 &  n_24504;
assign n_34144 = ~n_34142 & ~n_34143;
assign n_34145 =  x_2070 & ~n_34144;
assign n_34146 = ~x_2070 &  n_34144;
assign n_34147 = ~n_34145 & ~n_34146;
assign n_34148 =  x_2069 & ~n_24504;
assign n_34149 =  i_11 &  n_24504;
assign n_34150 = ~n_34148 & ~n_34149;
assign n_34151 =  x_2069 & ~n_34150;
assign n_34152 = ~x_2069 &  n_34150;
assign n_34153 = ~n_34151 & ~n_34152;
assign n_34154 =  x_2068 & ~n_24504;
assign n_34155 =  i_10 &  n_24504;
assign n_34156 = ~n_34154 & ~n_34155;
assign n_34157 =  x_2068 & ~n_34156;
assign n_34158 = ~x_2068 &  n_34156;
assign n_34159 = ~n_34157 & ~n_34158;
assign n_34160 =  x_2067 & ~n_24504;
assign n_34161 =  i_9 &  n_24504;
assign n_34162 = ~n_34160 & ~n_34161;
assign n_34163 =  x_2067 & ~n_34162;
assign n_34164 = ~x_2067 &  n_34162;
assign n_34165 = ~n_34163 & ~n_34164;
assign n_34166 =  x_2066 & ~n_24504;
assign n_34167 =  i_8 &  n_24504;
assign n_34168 = ~n_34166 & ~n_34167;
assign n_34169 =  x_2066 & ~n_34168;
assign n_34170 = ~x_2066 &  n_34168;
assign n_34171 = ~n_34169 & ~n_34170;
assign n_34172 =  x_2065 & ~n_24504;
assign n_34173 =  i_7 &  n_24504;
assign n_34174 = ~n_34172 & ~n_34173;
assign n_34175 =  x_2065 & ~n_34174;
assign n_34176 = ~x_2065 &  n_34174;
assign n_34177 = ~n_34175 & ~n_34176;
assign n_34178 =  x_2064 & ~n_24504;
assign n_34179 =  i_6 &  n_24504;
assign n_34180 = ~n_34178 & ~n_34179;
assign n_34181 =  x_2064 & ~n_34180;
assign n_34182 = ~x_2064 &  n_34180;
assign n_34183 = ~n_34181 & ~n_34182;
assign n_34184 =  x_2063 & ~n_24504;
assign n_34185 =  i_5 &  n_24504;
assign n_34186 = ~n_34184 & ~n_34185;
assign n_34187 =  x_2063 & ~n_34186;
assign n_34188 = ~x_2063 &  n_34186;
assign n_34189 = ~n_34187 & ~n_34188;
assign n_34190 =  x_2062 & ~n_24504;
assign n_34191 =  i_4 &  n_24504;
assign n_34192 = ~n_34190 & ~n_34191;
assign n_34193 =  x_2062 & ~n_34192;
assign n_34194 = ~x_2062 &  n_34192;
assign n_34195 = ~n_34193 & ~n_34194;
assign n_34196 =  x_2061 & ~n_24504;
assign n_34197 =  i_3 &  n_24504;
assign n_34198 = ~n_34196 & ~n_34197;
assign n_34199 =  x_2061 & ~n_34198;
assign n_34200 = ~x_2061 &  n_34198;
assign n_34201 = ~n_34199 & ~n_34200;
assign n_34202 =  x_2060 & ~n_24504;
assign n_34203 =  i_2 &  n_24504;
assign n_34204 = ~n_34202 & ~n_34203;
assign n_34205 =  x_2060 & ~n_34204;
assign n_34206 = ~x_2060 &  n_34204;
assign n_34207 = ~n_34205 & ~n_34206;
assign n_34208 =  x_2059 & ~n_24504;
assign n_34209 =  i_1 &  n_24504;
assign n_34210 = ~n_34208 & ~n_34209;
assign n_34211 =  x_2059 & ~n_34210;
assign n_34212 = ~x_2059 &  n_34210;
assign n_34213 = ~n_34211 & ~n_34212;
assign n_34214 =  x_2058 & ~n_16882;
assign n_34215 =  x_4967 &  n_16882;
assign n_34216 = ~n_34214 & ~n_34215;
assign n_34217 =  x_2058 & ~n_34216;
assign n_34218 = ~x_2058 &  n_34216;
assign n_34219 = ~n_34217 & ~n_34218;
assign n_34220 =  x_2057 & ~n_16882;
assign n_34221 =  x_4966 &  n_16882;
assign n_34222 = ~n_34220 & ~n_34221;
assign n_34223 =  x_2057 & ~n_34222;
assign n_34224 = ~x_2057 &  n_34222;
assign n_34225 = ~n_34223 & ~n_34224;
assign n_34226 =  x_2056 & ~n_16882;
assign n_34227 =  x_4965 &  n_16882;
assign n_34228 = ~n_34226 & ~n_34227;
assign n_34229 =  x_2056 & ~n_34228;
assign n_34230 = ~x_2056 &  n_34228;
assign n_34231 = ~n_34229 & ~n_34230;
assign n_34232 =  x_2055 & ~n_16882;
assign n_34233 =  x_4964 &  n_16882;
assign n_34234 = ~n_34232 & ~n_34233;
assign n_34235 =  x_2055 & ~n_34234;
assign n_34236 = ~x_2055 &  n_34234;
assign n_34237 = ~n_34235 & ~n_34236;
assign n_34238 =  x_2054 & ~n_16882;
assign n_34239 =  x_4963 &  n_16882;
assign n_34240 = ~n_34238 & ~n_34239;
assign n_34241 =  x_2054 & ~n_34240;
assign n_34242 = ~x_2054 &  n_34240;
assign n_34243 = ~n_34241 & ~n_34242;
assign n_34244 =  x_2053 & ~n_16882;
assign n_34245 =  x_4962 &  n_16882;
assign n_34246 = ~n_34244 & ~n_34245;
assign n_34247 =  x_2053 & ~n_34246;
assign n_34248 = ~x_2053 &  n_34246;
assign n_34249 = ~n_34247 & ~n_34248;
assign n_34250 =  x_2052 & ~n_16882;
assign n_34251 =  x_4961 &  n_16882;
assign n_34252 = ~n_34250 & ~n_34251;
assign n_34253 =  x_2052 & ~n_34252;
assign n_34254 = ~x_2052 &  n_34252;
assign n_34255 = ~n_34253 & ~n_34254;
assign n_34256 =  x_2051 & ~n_16882;
assign n_34257 =  x_4960 &  n_16882;
assign n_34258 = ~n_34256 & ~n_34257;
assign n_34259 =  x_2051 & ~n_34258;
assign n_34260 = ~x_2051 &  n_34258;
assign n_34261 = ~n_34259 & ~n_34260;
assign n_34262 =  x_2050 & ~n_16882;
assign n_34263 =  x_4959 &  n_16882;
assign n_34264 = ~n_34262 & ~n_34263;
assign n_34265 =  x_2050 & ~n_34264;
assign n_34266 = ~x_2050 &  n_34264;
assign n_34267 = ~n_34265 & ~n_34266;
assign n_34268 =  x_2049 & ~n_16882;
assign n_34269 =  x_4958 &  n_16882;
assign n_34270 = ~n_34268 & ~n_34269;
assign n_34271 =  x_2049 & ~n_34270;
assign n_34272 = ~x_2049 &  n_34270;
assign n_34273 = ~n_34271 & ~n_34272;
assign n_34274 =  x_2048 & ~n_16882;
assign n_34275 =  x_4957 &  n_16882;
assign n_34276 = ~n_34274 & ~n_34275;
assign n_34277 =  x_2048 & ~n_34276;
assign n_34278 = ~x_2048 &  n_34276;
assign n_34279 = ~n_34277 & ~n_34278;
assign n_34280 =  x_2047 & ~n_16882;
assign n_34281 =  x_4956 &  n_16882;
assign n_34282 = ~n_34280 & ~n_34281;
assign n_34283 =  x_2047 & ~n_34282;
assign n_34284 = ~x_2047 &  n_34282;
assign n_34285 = ~n_34283 & ~n_34284;
assign n_34286 =  x_2046 & ~n_16882;
assign n_34287 =  x_4955 &  n_16882;
assign n_34288 = ~n_34286 & ~n_34287;
assign n_34289 =  x_2046 & ~n_34288;
assign n_34290 = ~x_2046 &  n_34288;
assign n_34291 = ~n_34289 & ~n_34290;
assign n_34292 =  x_2045 & ~n_16882;
assign n_34293 =  x_4954 &  n_16882;
assign n_34294 = ~n_34292 & ~n_34293;
assign n_34295 =  x_2045 & ~n_34294;
assign n_34296 = ~x_2045 &  n_34294;
assign n_34297 = ~n_34295 & ~n_34296;
assign n_34298 =  x_2044 & ~n_16882;
assign n_34299 =  x_4953 &  n_16882;
assign n_34300 = ~n_34298 & ~n_34299;
assign n_34301 =  x_2044 & ~n_34300;
assign n_34302 = ~x_2044 &  n_34300;
assign n_34303 = ~n_34301 & ~n_34302;
assign n_34304 =  x_2043 & ~n_16882;
assign n_34305 =  x_4952 &  n_16882;
assign n_34306 = ~n_34304 & ~n_34305;
assign n_34307 =  x_2043 & ~n_34306;
assign n_34308 = ~x_2043 &  n_34306;
assign n_34309 = ~n_34307 & ~n_34308;
assign n_34310 =  x_2042 & ~n_16882;
assign n_34311 =  x_4951 &  n_16882;
assign n_34312 = ~n_34310 & ~n_34311;
assign n_34313 =  x_2042 & ~n_34312;
assign n_34314 = ~x_2042 &  n_34312;
assign n_34315 = ~n_34313 & ~n_34314;
assign n_34316 =  x_2041 & ~n_16882;
assign n_34317 =  x_4950 &  n_16882;
assign n_34318 = ~n_34316 & ~n_34317;
assign n_34319 =  x_2041 & ~n_34318;
assign n_34320 = ~x_2041 &  n_34318;
assign n_34321 = ~n_34319 & ~n_34320;
assign n_34322 =  x_2040 & ~n_16882;
assign n_34323 =  x_4949 &  n_16882;
assign n_34324 = ~n_34322 & ~n_34323;
assign n_34325 =  x_2040 & ~n_34324;
assign n_34326 = ~x_2040 &  n_34324;
assign n_34327 = ~n_34325 & ~n_34326;
assign n_34328 =  x_2039 & ~n_16882;
assign n_34329 =  x_4948 &  n_16882;
assign n_34330 = ~n_34328 & ~n_34329;
assign n_34331 =  x_2039 & ~n_34330;
assign n_34332 = ~x_2039 &  n_34330;
assign n_34333 = ~n_34331 & ~n_34332;
assign n_34334 =  x_2038 & ~n_16882;
assign n_34335 =  x_4947 &  n_16882;
assign n_34336 = ~n_34334 & ~n_34335;
assign n_34337 =  x_2038 & ~n_34336;
assign n_34338 = ~x_2038 &  n_34336;
assign n_34339 = ~n_34337 & ~n_34338;
assign n_34340 =  x_2037 & ~n_16882;
assign n_34341 =  x_4946 &  n_16882;
assign n_34342 = ~n_34340 & ~n_34341;
assign n_34343 =  x_2037 & ~n_34342;
assign n_34344 = ~x_2037 &  n_34342;
assign n_34345 = ~n_34343 & ~n_34344;
assign n_34346 =  x_2036 & ~n_16882;
assign n_34347 =  x_4945 &  n_16882;
assign n_34348 = ~n_34346 & ~n_34347;
assign n_34349 =  x_2036 & ~n_34348;
assign n_34350 = ~x_2036 &  n_34348;
assign n_34351 = ~n_34349 & ~n_34350;
assign n_34352 =  x_2035 & ~n_16882;
assign n_34353 =  x_4944 &  n_16882;
assign n_34354 = ~n_34352 & ~n_34353;
assign n_34355 =  x_2035 & ~n_34354;
assign n_34356 = ~x_2035 &  n_34354;
assign n_34357 = ~n_34355 & ~n_34356;
assign n_34358 =  x_2034 & ~n_16882;
assign n_34359 =  x_4943 &  n_16882;
assign n_34360 = ~n_34358 & ~n_34359;
assign n_34361 =  x_2034 & ~n_34360;
assign n_34362 = ~x_2034 &  n_34360;
assign n_34363 = ~n_34361 & ~n_34362;
assign n_34364 =  x_2033 & ~n_16882;
assign n_34365 =  x_4942 &  n_16882;
assign n_34366 = ~n_34364 & ~n_34365;
assign n_34367 =  x_2033 & ~n_34366;
assign n_34368 = ~x_2033 &  n_34366;
assign n_34369 = ~n_34367 & ~n_34368;
assign n_34370 =  x_2032 & ~n_16882;
assign n_34371 =  x_4941 &  n_16882;
assign n_34372 = ~n_34370 & ~n_34371;
assign n_34373 =  x_2032 & ~n_34372;
assign n_34374 = ~x_2032 &  n_34372;
assign n_34375 = ~n_34373 & ~n_34374;
assign n_34376 =  x_2031 & ~n_16882;
assign n_34377 =  x_4940 &  n_16882;
assign n_34378 = ~n_34376 & ~n_34377;
assign n_34379 =  x_2031 & ~n_34378;
assign n_34380 = ~x_2031 &  n_34378;
assign n_34381 = ~n_34379 & ~n_34380;
assign n_34382 =  x_2030 & ~n_16882;
assign n_34383 =  x_4939 &  n_16882;
assign n_34384 = ~n_34382 & ~n_34383;
assign n_34385 =  x_2030 & ~n_34384;
assign n_34386 = ~x_2030 &  n_34384;
assign n_34387 = ~n_34385 & ~n_34386;
assign n_34388 =  x_2029 & ~n_16882;
assign n_34389 =  x_4938 &  n_16882;
assign n_34390 = ~n_34388 & ~n_34389;
assign n_34391 =  x_2029 & ~n_34390;
assign n_34392 = ~x_2029 &  n_34390;
assign n_34393 = ~n_34391 & ~n_34392;
assign n_34394 =  x_2028 & ~n_16882;
assign n_34395 =  x_4937 &  n_16882;
assign n_34396 = ~n_34394 & ~n_34395;
assign n_34397 =  x_2028 & ~n_34396;
assign n_34398 = ~x_2028 &  n_34396;
assign n_34399 = ~n_34397 & ~n_34398;
assign n_34400 =  x_2027 & ~n_16882;
assign n_34401 =  x_4936 &  n_16882;
assign n_34402 = ~n_34400 & ~n_34401;
assign n_34403 =  x_2027 & ~n_34402;
assign n_34404 = ~x_2027 &  n_34402;
assign n_34405 = ~n_34403 & ~n_34404;
assign n_34406 =  n_24994 & ~n_12344;
assign n_34407 =  x_2026 & ~n_24994;
assign n_34408 = ~n_34406 & ~n_34407;
assign n_34409 =  x_2026 & ~n_34408;
assign n_34410 = ~x_2026 &  n_34408;
assign n_34411 = ~n_34409 & ~n_34410;
assign n_34412 =  n_24994 & ~n_12362;
assign n_34413 =  x_2025 & ~n_24994;
assign n_34414 = ~n_34412 & ~n_34413;
assign n_34415 =  x_2025 & ~n_34414;
assign n_34416 = ~x_2025 &  n_34414;
assign n_34417 = ~n_34415 & ~n_34416;
assign n_34418 =  n_24994 & ~n_12380;
assign n_34419 =  x_2024 & ~n_24994;
assign n_34420 = ~n_34418 & ~n_34419;
assign n_34421 =  x_2024 & ~n_34420;
assign n_34422 = ~x_2024 &  n_34420;
assign n_34423 = ~n_34421 & ~n_34422;
assign n_34424 =  n_24994 & ~n_12398;
assign n_34425 =  x_2023 & ~n_24994;
assign n_34426 = ~n_34424 & ~n_34425;
assign n_34427 =  x_2023 & ~n_34426;
assign n_34428 = ~x_2023 &  n_34426;
assign n_34429 = ~n_34427 & ~n_34428;
assign n_34430 =  n_24994 & ~n_12416;
assign n_34431 =  x_2022 & ~n_24994;
assign n_34432 = ~n_34430 & ~n_34431;
assign n_34433 =  x_2022 & ~n_34432;
assign n_34434 = ~x_2022 &  n_34432;
assign n_34435 = ~n_34433 & ~n_34434;
assign n_34436 =  n_24994 & ~n_12434;
assign n_34437 =  x_2021 & ~n_24994;
assign n_34438 = ~n_34436 & ~n_34437;
assign n_34439 =  x_2021 & ~n_34438;
assign n_34440 = ~x_2021 &  n_34438;
assign n_34441 = ~n_34439 & ~n_34440;
assign n_34442 =  n_24994 & ~n_12452;
assign n_34443 =  x_2020 & ~n_24994;
assign n_34444 = ~n_34442 & ~n_34443;
assign n_34445 =  x_2020 & ~n_34444;
assign n_34446 = ~x_2020 &  n_34444;
assign n_34447 = ~n_34445 & ~n_34446;
assign n_34448 =  n_24994 & ~n_12470;
assign n_34449 =  x_2019 & ~n_24994;
assign n_34450 = ~n_34448 & ~n_34449;
assign n_34451 =  x_2019 & ~n_34450;
assign n_34452 = ~x_2019 &  n_34450;
assign n_34453 = ~n_34451 & ~n_34452;
assign n_34454 =  n_24994 & ~n_12488;
assign n_34455 =  x_2018 & ~n_24994;
assign n_34456 = ~n_34454 & ~n_34455;
assign n_34457 =  x_2018 & ~n_34456;
assign n_34458 = ~x_2018 &  n_34456;
assign n_34459 = ~n_34457 & ~n_34458;
assign n_34460 =  n_24994 & ~n_12506;
assign n_34461 =  x_2017 & ~n_24994;
assign n_34462 = ~n_34460 & ~n_34461;
assign n_34463 =  x_2017 & ~n_34462;
assign n_34464 = ~x_2017 &  n_34462;
assign n_34465 = ~n_34463 & ~n_34464;
assign n_34466 =  n_24994 & ~n_12524;
assign n_34467 =  x_2016 & ~n_24994;
assign n_34468 = ~n_34466 & ~n_34467;
assign n_34469 =  x_2016 & ~n_34468;
assign n_34470 = ~x_2016 &  n_34468;
assign n_34471 = ~n_34469 & ~n_34470;
assign n_34472 =  n_24994 & ~n_12542;
assign n_34473 =  x_2015 & ~n_24994;
assign n_34474 = ~n_34472 & ~n_34473;
assign n_34475 =  x_2015 & ~n_34474;
assign n_34476 = ~x_2015 &  n_34474;
assign n_34477 = ~n_34475 & ~n_34476;
assign n_34478 =  n_24994 & ~n_12560;
assign n_34479 =  x_2014 & ~n_24994;
assign n_34480 = ~n_34478 & ~n_34479;
assign n_34481 =  x_2014 & ~n_34480;
assign n_34482 = ~x_2014 &  n_34480;
assign n_34483 = ~n_34481 & ~n_34482;
assign n_34484 =  n_24994 & ~n_12578;
assign n_34485 =  x_2013 & ~n_24994;
assign n_34486 = ~n_34484 & ~n_34485;
assign n_34487 =  x_2013 & ~n_34486;
assign n_34488 = ~x_2013 &  n_34486;
assign n_34489 = ~n_34487 & ~n_34488;
assign n_34490 =  n_24994 & ~n_12596;
assign n_34491 =  x_2012 & ~n_24994;
assign n_34492 = ~n_34490 & ~n_34491;
assign n_34493 =  x_2012 & ~n_34492;
assign n_34494 = ~x_2012 &  n_34492;
assign n_34495 = ~n_34493 & ~n_34494;
assign n_34496 =  n_24994 & ~n_12614;
assign n_34497 =  x_2011 & ~n_24994;
assign n_34498 = ~n_34496 & ~n_34497;
assign n_34499 =  x_2011 & ~n_34498;
assign n_34500 = ~x_2011 &  n_34498;
assign n_34501 = ~n_34499 & ~n_34500;
assign n_34502 =  n_24994 & ~n_12632;
assign n_34503 =  x_2010 & ~n_24994;
assign n_34504 = ~n_34502 & ~n_34503;
assign n_34505 =  x_2010 & ~n_34504;
assign n_34506 = ~x_2010 &  n_34504;
assign n_34507 = ~n_34505 & ~n_34506;
assign n_34508 =  n_24994 & ~n_12650;
assign n_34509 =  x_2009 & ~n_24994;
assign n_34510 = ~n_34508 & ~n_34509;
assign n_34511 =  x_2009 & ~n_34510;
assign n_34512 = ~x_2009 &  n_34510;
assign n_34513 = ~n_34511 & ~n_34512;
assign n_34514 =  n_24994 & ~n_12668;
assign n_34515 =  x_2008 & ~n_24994;
assign n_34516 = ~n_34514 & ~n_34515;
assign n_34517 =  x_2008 & ~n_34516;
assign n_34518 = ~x_2008 &  n_34516;
assign n_34519 = ~n_34517 & ~n_34518;
assign n_34520 =  n_24994 & ~n_12686;
assign n_34521 =  x_2007 & ~n_24994;
assign n_34522 = ~n_34520 & ~n_34521;
assign n_34523 =  x_2007 & ~n_34522;
assign n_34524 = ~x_2007 &  n_34522;
assign n_34525 = ~n_34523 & ~n_34524;
assign n_34526 =  n_24994 & ~n_12704;
assign n_34527 =  x_2006 & ~n_24994;
assign n_34528 = ~n_34526 & ~n_34527;
assign n_34529 =  x_2006 & ~n_34528;
assign n_34530 = ~x_2006 &  n_34528;
assign n_34531 = ~n_34529 & ~n_34530;
assign n_34532 =  n_24994 & ~n_12722;
assign n_34533 =  x_2005 & ~n_24994;
assign n_34534 = ~n_34532 & ~n_34533;
assign n_34535 =  x_2005 & ~n_34534;
assign n_34536 = ~x_2005 &  n_34534;
assign n_34537 = ~n_34535 & ~n_34536;
assign n_34538 =  n_24994 & ~n_12740;
assign n_34539 =  x_2004 & ~n_24994;
assign n_34540 = ~n_34538 & ~n_34539;
assign n_34541 =  x_2004 & ~n_34540;
assign n_34542 = ~x_2004 &  n_34540;
assign n_34543 = ~n_34541 & ~n_34542;
assign n_34544 =  n_24994 & ~n_12758;
assign n_34545 =  x_2003 & ~n_24994;
assign n_34546 = ~n_34544 & ~n_34545;
assign n_34547 =  x_2003 & ~n_34546;
assign n_34548 = ~x_2003 &  n_34546;
assign n_34549 = ~n_34547 & ~n_34548;
assign n_34550 =  n_24994 & ~n_12776;
assign n_34551 =  x_2002 & ~n_24994;
assign n_34552 = ~n_34550 & ~n_34551;
assign n_34553 =  x_2002 & ~n_34552;
assign n_34554 = ~x_2002 &  n_34552;
assign n_34555 = ~n_34553 & ~n_34554;
assign n_34556 =  n_24994 & ~n_12794;
assign n_34557 =  x_2001 & ~n_24994;
assign n_34558 = ~n_34556 & ~n_34557;
assign n_34559 =  x_2001 & ~n_34558;
assign n_34560 = ~x_2001 &  n_34558;
assign n_34561 = ~n_34559 & ~n_34560;
assign n_34562 =  n_24994 & ~n_12812;
assign n_34563 =  x_2000 & ~n_24994;
assign n_34564 = ~n_34562 & ~n_34563;
assign n_34565 =  x_2000 & ~n_34564;
assign n_34566 = ~x_2000 &  n_34564;
assign n_34567 = ~n_34565 & ~n_34566;
assign n_34568 =  n_24994 & ~n_12830;
assign n_34569 =  x_1999 & ~n_24994;
assign n_34570 = ~n_34568 & ~n_34569;
assign n_34571 =  x_1999 & ~n_34570;
assign n_34572 = ~x_1999 &  n_34570;
assign n_34573 = ~n_34571 & ~n_34572;
assign n_34574 =  n_24994 & ~n_12848;
assign n_34575 =  x_1998 & ~n_24994;
assign n_34576 = ~n_34574 & ~n_34575;
assign n_34577 =  x_1998 & ~n_34576;
assign n_34578 = ~x_1998 &  n_34576;
assign n_34579 = ~n_34577 & ~n_34578;
assign n_34580 =  n_24994 & ~n_12866;
assign n_34581 =  x_1997 & ~n_24994;
assign n_34582 = ~n_34580 & ~n_34581;
assign n_34583 =  x_1997 & ~n_34582;
assign n_34584 = ~x_1997 &  n_34582;
assign n_34585 = ~n_34583 & ~n_34584;
assign n_34586 =  n_24994 & ~n_12884;
assign n_34587 =  x_1996 & ~n_24994;
assign n_34588 = ~n_34586 & ~n_34587;
assign n_34589 =  x_1996 & ~n_34588;
assign n_34590 = ~x_1996 &  n_34588;
assign n_34591 = ~n_34589 & ~n_34590;
assign n_34592 =  n_24994 & ~n_12902;
assign n_34593 =  x_1995 & ~n_24994;
assign n_34594 = ~n_34592 & ~n_34593;
assign n_34595 =  x_1995 & ~n_34594;
assign n_34596 = ~x_1995 &  n_34594;
assign n_34597 = ~n_34595 & ~n_34596;
assign n_34598 =  n_349 &  n_8348;
assign n_34599 =  x_1994 & ~n_34598;
assign n_34600 =  i_32 &  n_34598;
assign n_34601 = ~n_34599 & ~n_34600;
assign n_34602 =  x_1994 & ~n_34601;
assign n_34603 = ~x_1994 &  n_34601;
assign n_34604 = ~n_34602 & ~n_34603;
assign n_34605 =  x_1993 & ~n_34598;
assign n_34606 =  i_31 &  n_34598;
assign n_34607 = ~n_34605 & ~n_34606;
assign n_34608 =  x_1993 & ~n_34607;
assign n_34609 = ~x_1993 &  n_34607;
assign n_34610 = ~n_34608 & ~n_34609;
assign n_34611 =  x_1992 & ~n_34598;
assign n_34612 =  i_30 &  n_34598;
assign n_34613 = ~n_34611 & ~n_34612;
assign n_34614 =  x_1992 & ~n_34613;
assign n_34615 = ~x_1992 &  n_34613;
assign n_34616 = ~n_34614 & ~n_34615;
assign n_34617 =  x_1991 & ~n_34598;
assign n_34618 =  i_29 &  n_34598;
assign n_34619 = ~n_34617 & ~n_34618;
assign n_34620 =  x_1991 & ~n_34619;
assign n_34621 = ~x_1991 &  n_34619;
assign n_34622 = ~n_34620 & ~n_34621;
assign n_34623 =  x_1990 & ~n_34598;
assign n_34624 =  i_28 &  n_34598;
assign n_34625 = ~n_34623 & ~n_34624;
assign n_34626 =  x_1990 & ~n_34625;
assign n_34627 = ~x_1990 &  n_34625;
assign n_34628 = ~n_34626 & ~n_34627;
assign n_34629 =  x_1989 & ~n_34598;
assign n_34630 =  i_27 &  n_34598;
assign n_34631 = ~n_34629 & ~n_34630;
assign n_34632 =  x_1989 & ~n_34631;
assign n_34633 = ~x_1989 &  n_34631;
assign n_34634 = ~n_34632 & ~n_34633;
assign n_34635 =  x_1988 & ~n_34598;
assign n_34636 =  i_26 &  n_34598;
assign n_34637 = ~n_34635 & ~n_34636;
assign n_34638 =  x_1988 & ~n_34637;
assign n_34639 = ~x_1988 &  n_34637;
assign n_34640 = ~n_34638 & ~n_34639;
assign n_34641 =  x_1987 & ~n_34598;
assign n_34642 =  i_25 &  n_34598;
assign n_34643 = ~n_34641 & ~n_34642;
assign n_34644 =  x_1987 & ~n_34643;
assign n_34645 = ~x_1987 &  n_34643;
assign n_34646 = ~n_34644 & ~n_34645;
assign n_34647 =  x_1986 & ~n_34598;
assign n_34648 =  i_24 &  n_34598;
assign n_34649 = ~n_34647 & ~n_34648;
assign n_34650 =  x_1986 & ~n_34649;
assign n_34651 = ~x_1986 &  n_34649;
assign n_34652 = ~n_34650 & ~n_34651;
assign n_34653 =  x_1985 & ~n_34598;
assign n_34654 =  i_23 &  n_34598;
assign n_34655 = ~n_34653 & ~n_34654;
assign n_34656 =  x_1985 & ~n_34655;
assign n_34657 = ~x_1985 &  n_34655;
assign n_34658 = ~n_34656 & ~n_34657;
assign n_34659 =  x_1984 & ~n_34598;
assign n_34660 =  i_22 &  n_34598;
assign n_34661 = ~n_34659 & ~n_34660;
assign n_34662 =  x_1984 & ~n_34661;
assign n_34663 = ~x_1984 &  n_34661;
assign n_34664 = ~n_34662 & ~n_34663;
assign n_34665 =  x_1983 & ~n_34598;
assign n_34666 =  i_21 &  n_34598;
assign n_34667 = ~n_34665 & ~n_34666;
assign n_34668 =  x_1983 & ~n_34667;
assign n_34669 = ~x_1983 &  n_34667;
assign n_34670 = ~n_34668 & ~n_34669;
assign n_34671 =  x_1982 & ~n_34598;
assign n_34672 =  i_20 &  n_34598;
assign n_34673 = ~n_34671 & ~n_34672;
assign n_34674 =  x_1982 & ~n_34673;
assign n_34675 = ~x_1982 &  n_34673;
assign n_34676 = ~n_34674 & ~n_34675;
assign n_34677 =  x_1981 & ~n_34598;
assign n_34678 =  i_19 &  n_34598;
assign n_34679 = ~n_34677 & ~n_34678;
assign n_34680 =  x_1981 & ~n_34679;
assign n_34681 = ~x_1981 &  n_34679;
assign n_34682 = ~n_34680 & ~n_34681;
assign n_34683 =  x_1980 & ~n_34598;
assign n_34684 =  i_18 &  n_34598;
assign n_34685 = ~n_34683 & ~n_34684;
assign n_34686 =  x_1980 & ~n_34685;
assign n_34687 = ~x_1980 &  n_34685;
assign n_34688 = ~n_34686 & ~n_34687;
assign n_34689 =  x_1979 & ~n_34598;
assign n_34690 =  i_17 &  n_34598;
assign n_34691 = ~n_34689 & ~n_34690;
assign n_34692 =  x_1979 & ~n_34691;
assign n_34693 = ~x_1979 &  n_34691;
assign n_34694 = ~n_34692 & ~n_34693;
assign n_34695 =  x_1978 & ~n_34598;
assign n_34696 =  i_16 &  n_34598;
assign n_34697 = ~n_34695 & ~n_34696;
assign n_34698 =  x_1978 & ~n_34697;
assign n_34699 = ~x_1978 &  n_34697;
assign n_34700 = ~n_34698 & ~n_34699;
assign n_34701 =  x_1977 & ~n_34598;
assign n_34702 =  i_15 &  n_34598;
assign n_34703 = ~n_34701 & ~n_34702;
assign n_34704 =  x_1977 & ~n_34703;
assign n_34705 = ~x_1977 &  n_34703;
assign n_34706 = ~n_34704 & ~n_34705;
assign n_34707 =  x_1976 & ~n_34598;
assign n_34708 =  i_14 &  n_34598;
assign n_34709 = ~n_34707 & ~n_34708;
assign n_34710 =  x_1976 & ~n_34709;
assign n_34711 = ~x_1976 &  n_34709;
assign n_34712 = ~n_34710 & ~n_34711;
assign n_34713 =  x_1975 & ~n_34598;
assign n_34714 =  i_13 &  n_34598;
assign n_34715 = ~n_34713 & ~n_34714;
assign n_34716 =  x_1975 & ~n_34715;
assign n_34717 = ~x_1975 &  n_34715;
assign n_34718 = ~n_34716 & ~n_34717;
assign n_34719 =  x_1974 & ~n_34598;
assign n_34720 =  i_12 &  n_34598;
assign n_34721 = ~n_34719 & ~n_34720;
assign n_34722 =  x_1974 & ~n_34721;
assign n_34723 = ~x_1974 &  n_34721;
assign n_34724 = ~n_34722 & ~n_34723;
assign n_34725 =  x_1973 & ~n_34598;
assign n_34726 =  i_11 &  n_34598;
assign n_34727 = ~n_34725 & ~n_34726;
assign n_34728 =  x_1973 & ~n_34727;
assign n_34729 = ~x_1973 &  n_34727;
assign n_34730 = ~n_34728 & ~n_34729;
assign n_34731 =  x_1972 & ~n_34598;
assign n_34732 =  i_10 &  n_34598;
assign n_34733 = ~n_34731 & ~n_34732;
assign n_34734 =  x_1972 & ~n_34733;
assign n_34735 = ~x_1972 &  n_34733;
assign n_34736 = ~n_34734 & ~n_34735;
assign n_34737 =  x_1971 & ~n_34598;
assign n_34738 =  i_9 &  n_34598;
assign n_34739 = ~n_34737 & ~n_34738;
assign n_34740 =  x_1971 & ~n_34739;
assign n_34741 = ~x_1971 &  n_34739;
assign n_34742 = ~n_34740 & ~n_34741;
assign n_34743 =  x_1970 & ~n_34598;
assign n_34744 =  i_8 &  n_34598;
assign n_34745 = ~n_34743 & ~n_34744;
assign n_34746 =  x_1970 & ~n_34745;
assign n_34747 = ~x_1970 &  n_34745;
assign n_34748 = ~n_34746 & ~n_34747;
assign n_34749 =  x_1969 & ~n_34598;
assign n_34750 =  i_7 &  n_34598;
assign n_34751 = ~n_34749 & ~n_34750;
assign n_34752 =  x_1969 & ~n_34751;
assign n_34753 = ~x_1969 &  n_34751;
assign n_34754 = ~n_34752 & ~n_34753;
assign n_34755 =  x_1968 & ~n_34598;
assign n_34756 =  i_6 &  n_34598;
assign n_34757 = ~n_34755 & ~n_34756;
assign n_34758 =  x_1968 & ~n_34757;
assign n_34759 = ~x_1968 &  n_34757;
assign n_34760 = ~n_34758 & ~n_34759;
assign n_34761 =  x_1967 & ~n_34598;
assign n_34762 =  i_5 &  n_34598;
assign n_34763 = ~n_34761 & ~n_34762;
assign n_34764 =  x_1967 & ~n_34763;
assign n_34765 = ~x_1967 &  n_34763;
assign n_34766 = ~n_34764 & ~n_34765;
assign n_34767 =  x_1966 & ~n_34598;
assign n_34768 =  i_4 &  n_34598;
assign n_34769 = ~n_34767 & ~n_34768;
assign n_34770 =  x_1966 & ~n_34769;
assign n_34771 = ~x_1966 &  n_34769;
assign n_34772 = ~n_34770 & ~n_34771;
assign n_34773 =  x_1965 & ~n_34598;
assign n_34774 =  i_3 &  n_34598;
assign n_34775 = ~n_34773 & ~n_34774;
assign n_34776 =  x_1965 & ~n_34775;
assign n_34777 = ~x_1965 &  n_34775;
assign n_34778 = ~n_34776 & ~n_34777;
assign n_34779 =  x_1964 & ~n_34598;
assign n_34780 =  i_2 &  n_34598;
assign n_34781 = ~n_34779 & ~n_34780;
assign n_34782 =  x_1964 & ~n_34781;
assign n_34783 = ~x_1964 &  n_34781;
assign n_34784 = ~n_34782 & ~n_34783;
assign n_34785 =  x_1963 & ~n_34598;
assign n_34786 =  i_1 &  n_34598;
assign n_34787 = ~n_34785 & ~n_34786;
assign n_34788 =  x_1963 & ~n_34787;
assign n_34789 = ~x_1963 &  n_34787;
assign n_34790 = ~n_34788 & ~n_34789;
assign n_34791 =  n_28642 & ~n_12344;
assign n_34792 =  x_1962 & ~n_28642;
assign n_34793 = ~n_34791 & ~n_34792;
assign n_34794 =  x_1962 & ~n_34793;
assign n_34795 = ~x_1962 &  n_34793;
assign n_34796 = ~n_34794 & ~n_34795;
assign n_34797 =  n_28642 & ~n_12362;
assign n_34798 =  x_1961 & ~n_28642;
assign n_34799 = ~n_34797 & ~n_34798;
assign n_34800 =  x_1961 & ~n_34799;
assign n_34801 = ~x_1961 &  n_34799;
assign n_34802 = ~n_34800 & ~n_34801;
assign n_34803 =  n_28642 & ~n_12380;
assign n_34804 =  x_1960 & ~n_28642;
assign n_34805 = ~n_34803 & ~n_34804;
assign n_34806 =  x_1960 & ~n_34805;
assign n_34807 = ~x_1960 &  n_34805;
assign n_34808 = ~n_34806 & ~n_34807;
assign n_34809 =  n_28642 & ~n_12398;
assign n_34810 =  x_1959 & ~n_28642;
assign n_34811 = ~n_34809 & ~n_34810;
assign n_34812 =  x_1959 & ~n_34811;
assign n_34813 = ~x_1959 &  n_34811;
assign n_34814 = ~n_34812 & ~n_34813;
assign n_34815 =  n_28642 & ~n_12416;
assign n_34816 =  x_1958 & ~n_28642;
assign n_34817 = ~n_34815 & ~n_34816;
assign n_34818 =  x_1958 & ~n_34817;
assign n_34819 = ~x_1958 &  n_34817;
assign n_34820 = ~n_34818 & ~n_34819;
assign n_34821 =  n_28642 & ~n_12434;
assign n_34822 =  x_1957 & ~n_28642;
assign n_34823 = ~n_34821 & ~n_34822;
assign n_34824 =  x_1957 & ~n_34823;
assign n_34825 = ~x_1957 &  n_34823;
assign n_34826 = ~n_34824 & ~n_34825;
assign n_34827 =  n_28642 & ~n_12452;
assign n_34828 =  x_1956 & ~n_28642;
assign n_34829 = ~n_34827 & ~n_34828;
assign n_34830 =  x_1956 & ~n_34829;
assign n_34831 = ~x_1956 &  n_34829;
assign n_34832 = ~n_34830 & ~n_34831;
assign n_34833 =  n_28642 & ~n_12470;
assign n_34834 =  x_1955 & ~n_28642;
assign n_34835 = ~n_34833 & ~n_34834;
assign n_34836 =  x_1955 & ~n_34835;
assign n_34837 = ~x_1955 &  n_34835;
assign n_34838 = ~n_34836 & ~n_34837;
assign n_34839 =  n_28642 & ~n_12488;
assign n_34840 =  x_1954 & ~n_28642;
assign n_34841 = ~n_34839 & ~n_34840;
assign n_34842 =  x_1954 & ~n_34841;
assign n_34843 = ~x_1954 &  n_34841;
assign n_34844 = ~n_34842 & ~n_34843;
assign n_34845 =  n_28642 & ~n_12506;
assign n_34846 =  x_1953 & ~n_28642;
assign n_34847 = ~n_34845 & ~n_34846;
assign n_34848 =  x_1953 & ~n_34847;
assign n_34849 = ~x_1953 &  n_34847;
assign n_34850 = ~n_34848 & ~n_34849;
assign n_34851 =  n_28642 & ~n_12524;
assign n_34852 =  x_1952 & ~n_28642;
assign n_34853 = ~n_34851 & ~n_34852;
assign n_34854 =  x_1952 & ~n_34853;
assign n_34855 = ~x_1952 &  n_34853;
assign n_34856 = ~n_34854 & ~n_34855;
assign n_34857 =  n_28642 & ~n_12542;
assign n_34858 =  x_1951 & ~n_28642;
assign n_34859 = ~n_34857 & ~n_34858;
assign n_34860 =  x_1951 & ~n_34859;
assign n_34861 = ~x_1951 &  n_34859;
assign n_34862 = ~n_34860 & ~n_34861;
assign n_34863 =  n_28642 & ~n_12560;
assign n_34864 =  x_1950 & ~n_28642;
assign n_34865 = ~n_34863 & ~n_34864;
assign n_34866 =  x_1950 & ~n_34865;
assign n_34867 = ~x_1950 &  n_34865;
assign n_34868 = ~n_34866 & ~n_34867;
assign n_34869 =  n_28642 & ~n_12578;
assign n_34870 =  x_1949 & ~n_28642;
assign n_34871 = ~n_34869 & ~n_34870;
assign n_34872 =  x_1949 & ~n_34871;
assign n_34873 = ~x_1949 &  n_34871;
assign n_34874 = ~n_34872 & ~n_34873;
assign n_34875 =  n_28642 & ~n_12596;
assign n_34876 =  x_1948 & ~n_28642;
assign n_34877 = ~n_34875 & ~n_34876;
assign n_34878 =  x_1948 & ~n_34877;
assign n_34879 = ~x_1948 &  n_34877;
assign n_34880 = ~n_34878 & ~n_34879;
assign n_34881 =  n_28642 & ~n_12614;
assign n_34882 =  x_1947 & ~n_28642;
assign n_34883 = ~n_34881 & ~n_34882;
assign n_34884 =  x_1947 & ~n_34883;
assign n_34885 = ~x_1947 &  n_34883;
assign n_34886 = ~n_34884 & ~n_34885;
assign n_34887 =  n_28642 & ~n_12632;
assign n_34888 =  x_1946 & ~n_28642;
assign n_34889 = ~n_34887 & ~n_34888;
assign n_34890 =  x_1946 & ~n_34889;
assign n_34891 = ~x_1946 &  n_34889;
assign n_34892 = ~n_34890 & ~n_34891;
assign n_34893 =  n_28642 & ~n_12650;
assign n_34894 =  x_1945 & ~n_28642;
assign n_34895 = ~n_34893 & ~n_34894;
assign n_34896 =  x_1945 & ~n_34895;
assign n_34897 = ~x_1945 &  n_34895;
assign n_34898 = ~n_34896 & ~n_34897;
assign n_34899 =  n_28642 & ~n_12668;
assign n_34900 =  x_1944 & ~n_28642;
assign n_34901 = ~n_34899 & ~n_34900;
assign n_34902 =  x_1944 & ~n_34901;
assign n_34903 = ~x_1944 &  n_34901;
assign n_34904 = ~n_34902 & ~n_34903;
assign n_34905 =  n_28642 & ~n_12686;
assign n_34906 =  x_1943 & ~n_28642;
assign n_34907 = ~n_34905 & ~n_34906;
assign n_34908 =  x_1943 & ~n_34907;
assign n_34909 = ~x_1943 &  n_34907;
assign n_34910 = ~n_34908 & ~n_34909;
assign n_34911 =  n_28642 & ~n_12704;
assign n_34912 =  x_1942 & ~n_28642;
assign n_34913 = ~n_34911 & ~n_34912;
assign n_34914 =  x_1942 & ~n_34913;
assign n_34915 = ~x_1942 &  n_34913;
assign n_34916 = ~n_34914 & ~n_34915;
assign n_34917 =  n_28642 & ~n_12722;
assign n_34918 =  x_1941 & ~n_28642;
assign n_34919 = ~n_34917 & ~n_34918;
assign n_34920 =  x_1941 & ~n_34919;
assign n_34921 = ~x_1941 &  n_34919;
assign n_34922 = ~n_34920 & ~n_34921;
assign n_34923 =  n_28642 & ~n_12740;
assign n_34924 =  x_1940 & ~n_28642;
assign n_34925 = ~n_34923 & ~n_34924;
assign n_34926 =  x_1940 & ~n_34925;
assign n_34927 = ~x_1940 &  n_34925;
assign n_34928 = ~n_34926 & ~n_34927;
assign n_34929 =  n_28642 & ~n_12758;
assign n_34930 =  x_1939 & ~n_28642;
assign n_34931 = ~n_34929 & ~n_34930;
assign n_34932 =  x_1939 & ~n_34931;
assign n_34933 = ~x_1939 &  n_34931;
assign n_34934 = ~n_34932 & ~n_34933;
assign n_34935 =  n_28642 & ~n_12776;
assign n_34936 =  x_1938 & ~n_28642;
assign n_34937 = ~n_34935 & ~n_34936;
assign n_34938 =  x_1938 & ~n_34937;
assign n_34939 = ~x_1938 &  n_34937;
assign n_34940 = ~n_34938 & ~n_34939;
assign n_34941 =  n_28642 & ~n_12794;
assign n_34942 =  x_1937 & ~n_28642;
assign n_34943 = ~n_34941 & ~n_34942;
assign n_34944 =  x_1937 & ~n_34943;
assign n_34945 = ~x_1937 &  n_34943;
assign n_34946 = ~n_34944 & ~n_34945;
assign n_34947 =  n_28642 & ~n_12812;
assign n_34948 =  x_1936 & ~n_28642;
assign n_34949 = ~n_34947 & ~n_34948;
assign n_34950 =  x_1936 & ~n_34949;
assign n_34951 = ~x_1936 &  n_34949;
assign n_34952 = ~n_34950 & ~n_34951;
assign n_34953 =  n_28642 & ~n_12830;
assign n_34954 =  x_1935 & ~n_28642;
assign n_34955 = ~n_34953 & ~n_34954;
assign n_34956 =  x_1935 & ~n_34955;
assign n_34957 = ~x_1935 &  n_34955;
assign n_34958 = ~n_34956 & ~n_34957;
assign n_34959 =  n_28642 & ~n_12848;
assign n_34960 =  x_1934 & ~n_28642;
assign n_34961 = ~n_34959 & ~n_34960;
assign n_34962 =  x_1934 & ~n_34961;
assign n_34963 = ~x_1934 &  n_34961;
assign n_34964 = ~n_34962 & ~n_34963;
assign n_34965 =  n_28642 & ~n_12866;
assign n_34966 =  x_1933 & ~n_28642;
assign n_34967 = ~n_34965 & ~n_34966;
assign n_34968 =  x_1933 & ~n_34967;
assign n_34969 = ~x_1933 &  n_34967;
assign n_34970 = ~n_34968 & ~n_34969;
assign n_34971 =  n_28642 & ~n_12884;
assign n_34972 =  x_1932 & ~n_28642;
assign n_34973 = ~n_34971 & ~n_34972;
assign n_34974 =  x_1932 & ~n_34973;
assign n_34975 = ~x_1932 &  n_34973;
assign n_34976 = ~n_34974 & ~n_34975;
assign n_34977 =  n_28642 & ~n_12902;
assign n_34978 =  x_1931 & ~n_28642;
assign n_34979 = ~n_34977 & ~n_34978;
assign n_34980 =  x_1931 & ~n_34979;
assign n_34981 = ~x_1931 &  n_34979;
assign n_34982 = ~n_34980 & ~n_34981;
assign n_34983 =  x_1930 & ~n_26446;
assign n_34984 =  i_32 &  n_26446;
assign n_34985 = ~n_34983 & ~n_34984;
assign n_34986 =  x_1930 & ~n_34985;
assign n_34987 = ~x_1930 &  n_34985;
assign n_34988 = ~n_34986 & ~n_34987;
assign n_34989 =  x_1929 & ~n_26446;
assign n_34990 =  i_31 &  n_26446;
assign n_34991 = ~n_34989 & ~n_34990;
assign n_34992 =  x_1929 & ~n_34991;
assign n_34993 = ~x_1929 &  n_34991;
assign n_34994 = ~n_34992 & ~n_34993;
assign n_34995 =  x_1928 & ~n_26446;
assign n_34996 =  i_30 &  n_26446;
assign n_34997 = ~n_34995 & ~n_34996;
assign n_34998 =  x_1928 & ~n_34997;
assign n_34999 = ~x_1928 &  n_34997;
assign n_35000 = ~n_34998 & ~n_34999;
assign n_35001 =  x_1927 & ~n_26446;
assign n_35002 =  i_29 &  n_26446;
assign n_35003 = ~n_35001 & ~n_35002;
assign n_35004 =  x_1927 & ~n_35003;
assign n_35005 = ~x_1927 &  n_35003;
assign n_35006 = ~n_35004 & ~n_35005;
assign n_35007 =  x_1926 & ~n_26446;
assign n_35008 =  i_28 &  n_26446;
assign n_35009 = ~n_35007 & ~n_35008;
assign n_35010 =  x_1926 & ~n_35009;
assign n_35011 = ~x_1926 &  n_35009;
assign n_35012 = ~n_35010 & ~n_35011;
assign n_35013 =  x_1925 & ~n_26446;
assign n_35014 =  i_27 &  n_26446;
assign n_35015 = ~n_35013 & ~n_35014;
assign n_35016 =  x_1925 & ~n_35015;
assign n_35017 = ~x_1925 &  n_35015;
assign n_35018 = ~n_35016 & ~n_35017;
assign n_35019 =  x_1924 & ~n_26446;
assign n_35020 =  i_26 &  n_26446;
assign n_35021 = ~n_35019 & ~n_35020;
assign n_35022 =  x_1924 & ~n_35021;
assign n_35023 = ~x_1924 &  n_35021;
assign n_35024 = ~n_35022 & ~n_35023;
assign n_35025 =  x_1923 & ~n_26446;
assign n_35026 =  i_25 &  n_26446;
assign n_35027 = ~n_35025 & ~n_35026;
assign n_35028 =  x_1923 & ~n_35027;
assign n_35029 = ~x_1923 &  n_35027;
assign n_35030 = ~n_35028 & ~n_35029;
assign n_35031 =  x_1922 & ~n_26446;
assign n_35032 =  i_24 &  n_26446;
assign n_35033 = ~n_35031 & ~n_35032;
assign n_35034 =  x_1922 & ~n_35033;
assign n_35035 = ~x_1922 &  n_35033;
assign n_35036 = ~n_35034 & ~n_35035;
assign n_35037 =  x_1921 & ~n_26446;
assign n_35038 =  i_23 &  n_26446;
assign n_35039 = ~n_35037 & ~n_35038;
assign n_35040 =  x_1921 & ~n_35039;
assign n_35041 = ~x_1921 &  n_35039;
assign n_35042 = ~n_35040 & ~n_35041;
assign n_35043 =  x_1920 & ~n_26446;
assign n_35044 =  i_22 &  n_26446;
assign n_35045 = ~n_35043 & ~n_35044;
assign n_35046 =  x_1920 & ~n_35045;
assign n_35047 = ~x_1920 &  n_35045;
assign n_35048 = ~n_35046 & ~n_35047;
assign n_35049 =  x_1919 & ~n_26446;
assign n_35050 =  i_21 &  n_26446;
assign n_35051 = ~n_35049 & ~n_35050;
assign n_35052 =  x_1919 & ~n_35051;
assign n_35053 = ~x_1919 &  n_35051;
assign n_35054 = ~n_35052 & ~n_35053;
assign n_35055 =  x_1918 & ~n_26446;
assign n_35056 =  i_20 &  n_26446;
assign n_35057 = ~n_35055 & ~n_35056;
assign n_35058 =  x_1918 & ~n_35057;
assign n_35059 = ~x_1918 &  n_35057;
assign n_35060 = ~n_35058 & ~n_35059;
assign n_35061 =  x_1917 & ~n_26446;
assign n_35062 =  i_19 &  n_26446;
assign n_35063 = ~n_35061 & ~n_35062;
assign n_35064 =  x_1917 & ~n_35063;
assign n_35065 = ~x_1917 &  n_35063;
assign n_35066 = ~n_35064 & ~n_35065;
assign n_35067 =  x_1916 & ~n_26446;
assign n_35068 =  i_18 &  n_26446;
assign n_35069 = ~n_35067 & ~n_35068;
assign n_35070 =  x_1916 & ~n_35069;
assign n_35071 = ~x_1916 &  n_35069;
assign n_35072 = ~n_35070 & ~n_35071;
assign n_35073 =  x_1915 & ~n_26446;
assign n_35074 =  i_17 &  n_26446;
assign n_35075 = ~n_35073 & ~n_35074;
assign n_35076 =  x_1915 & ~n_35075;
assign n_35077 = ~x_1915 &  n_35075;
assign n_35078 = ~n_35076 & ~n_35077;
assign n_35079 =  x_1914 & ~n_26446;
assign n_35080 =  i_16 &  n_26446;
assign n_35081 = ~n_35079 & ~n_35080;
assign n_35082 =  x_1914 & ~n_35081;
assign n_35083 = ~x_1914 &  n_35081;
assign n_35084 = ~n_35082 & ~n_35083;
assign n_35085 =  x_1913 & ~n_26446;
assign n_35086 =  i_15 &  n_26446;
assign n_35087 = ~n_35085 & ~n_35086;
assign n_35088 =  x_1913 & ~n_35087;
assign n_35089 = ~x_1913 &  n_35087;
assign n_35090 = ~n_35088 & ~n_35089;
assign n_35091 =  x_1912 & ~n_26446;
assign n_35092 =  i_14 &  n_26446;
assign n_35093 = ~n_35091 & ~n_35092;
assign n_35094 =  x_1912 & ~n_35093;
assign n_35095 = ~x_1912 &  n_35093;
assign n_35096 = ~n_35094 & ~n_35095;
assign n_35097 =  x_1911 & ~n_26446;
assign n_35098 =  i_13 &  n_26446;
assign n_35099 = ~n_35097 & ~n_35098;
assign n_35100 =  x_1911 & ~n_35099;
assign n_35101 = ~x_1911 &  n_35099;
assign n_35102 = ~n_35100 & ~n_35101;
assign n_35103 =  x_1910 & ~n_26446;
assign n_35104 =  i_12 &  n_26446;
assign n_35105 = ~n_35103 & ~n_35104;
assign n_35106 =  x_1910 & ~n_35105;
assign n_35107 = ~x_1910 &  n_35105;
assign n_35108 = ~n_35106 & ~n_35107;
assign n_35109 =  x_1909 & ~n_26446;
assign n_35110 =  i_11 &  n_26446;
assign n_35111 = ~n_35109 & ~n_35110;
assign n_35112 =  x_1909 & ~n_35111;
assign n_35113 = ~x_1909 &  n_35111;
assign n_35114 = ~n_35112 & ~n_35113;
assign n_35115 =  x_1908 & ~n_26446;
assign n_35116 =  i_10 &  n_26446;
assign n_35117 = ~n_35115 & ~n_35116;
assign n_35118 =  x_1908 & ~n_35117;
assign n_35119 = ~x_1908 &  n_35117;
assign n_35120 = ~n_35118 & ~n_35119;
assign n_35121 =  x_1907 & ~n_26446;
assign n_35122 =  i_9 &  n_26446;
assign n_35123 = ~n_35121 & ~n_35122;
assign n_35124 =  x_1907 & ~n_35123;
assign n_35125 = ~x_1907 &  n_35123;
assign n_35126 = ~n_35124 & ~n_35125;
assign n_35127 =  x_1906 & ~n_26446;
assign n_35128 =  i_8 &  n_26446;
assign n_35129 = ~n_35127 & ~n_35128;
assign n_35130 =  x_1906 & ~n_35129;
assign n_35131 = ~x_1906 &  n_35129;
assign n_35132 = ~n_35130 & ~n_35131;
assign n_35133 =  x_1905 & ~n_26446;
assign n_35134 =  i_7 &  n_26446;
assign n_35135 = ~n_35133 & ~n_35134;
assign n_35136 =  x_1905 & ~n_35135;
assign n_35137 = ~x_1905 &  n_35135;
assign n_35138 = ~n_35136 & ~n_35137;
assign n_35139 =  x_1904 & ~n_26446;
assign n_35140 =  i_6 &  n_26446;
assign n_35141 = ~n_35139 & ~n_35140;
assign n_35142 =  x_1904 & ~n_35141;
assign n_35143 = ~x_1904 &  n_35141;
assign n_35144 = ~n_35142 & ~n_35143;
assign n_35145 =  x_1903 & ~n_26446;
assign n_35146 =  i_5 &  n_26446;
assign n_35147 = ~n_35145 & ~n_35146;
assign n_35148 =  x_1903 & ~n_35147;
assign n_35149 = ~x_1903 &  n_35147;
assign n_35150 = ~n_35148 & ~n_35149;
assign n_35151 =  x_1902 & ~n_26446;
assign n_35152 =  i_4 &  n_26446;
assign n_35153 = ~n_35151 & ~n_35152;
assign n_35154 =  x_1902 & ~n_35153;
assign n_35155 = ~x_1902 &  n_35153;
assign n_35156 = ~n_35154 & ~n_35155;
assign n_35157 =  x_1901 & ~n_26446;
assign n_35158 =  i_3 &  n_26446;
assign n_35159 = ~n_35157 & ~n_35158;
assign n_35160 =  x_1901 & ~n_35159;
assign n_35161 = ~x_1901 &  n_35159;
assign n_35162 = ~n_35160 & ~n_35161;
assign n_35163 =  x_1900 & ~n_26446;
assign n_35164 =  i_2 &  n_26446;
assign n_35165 = ~n_35163 & ~n_35164;
assign n_35166 =  x_1900 & ~n_35165;
assign n_35167 = ~x_1900 &  n_35165;
assign n_35168 = ~n_35166 & ~n_35167;
assign n_35169 =  x_1899 & ~n_26446;
assign n_35170 =  i_1 &  n_26446;
assign n_35171 = ~n_35169 & ~n_35170;
assign n_35172 =  x_1899 & ~n_35171;
assign n_35173 = ~x_1899 &  n_35171;
assign n_35174 = ~n_35172 & ~n_35173;
assign n_35175 =  x_1898 & ~n_24592;
assign n_35176 =  i_32 &  n_24592;
assign n_35177 = ~n_35175 & ~n_35176;
assign n_35178 =  x_1898 & ~n_35177;
assign n_35179 = ~x_1898 &  n_35177;
assign n_35180 = ~n_35178 & ~n_35179;
assign n_35181 =  x_1897 & ~n_24592;
assign n_35182 =  i_31 &  n_24592;
assign n_35183 = ~n_35181 & ~n_35182;
assign n_35184 =  x_1897 & ~n_35183;
assign n_35185 = ~x_1897 &  n_35183;
assign n_35186 = ~n_35184 & ~n_35185;
assign n_35187 =  x_1896 & ~n_24592;
assign n_35188 =  i_30 &  n_24592;
assign n_35189 = ~n_35187 & ~n_35188;
assign n_35190 =  x_1896 & ~n_35189;
assign n_35191 = ~x_1896 &  n_35189;
assign n_35192 = ~n_35190 & ~n_35191;
assign n_35193 =  x_1895 & ~n_24592;
assign n_35194 =  i_29 &  n_24592;
assign n_35195 = ~n_35193 & ~n_35194;
assign n_35196 =  x_1895 & ~n_35195;
assign n_35197 = ~x_1895 &  n_35195;
assign n_35198 = ~n_35196 & ~n_35197;
assign n_35199 =  x_1894 & ~n_24592;
assign n_35200 =  i_28 &  n_24592;
assign n_35201 = ~n_35199 & ~n_35200;
assign n_35202 =  x_1894 & ~n_35201;
assign n_35203 = ~x_1894 &  n_35201;
assign n_35204 = ~n_35202 & ~n_35203;
assign n_35205 =  x_1893 & ~n_24592;
assign n_35206 =  i_27 &  n_24592;
assign n_35207 = ~n_35205 & ~n_35206;
assign n_35208 =  x_1893 & ~n_35207;
assign n_35209 = ~x_1893 &  n_35207;
assign n_35210 = ~n_35208 & ~n_35209;
assign n_35211 =  x_1892 & ~n_24592;
assign n_35212 =  i_26 &  n_24592;
assign n_35213 = ~n_35211 & ~n_35212;
assign n_35214 =  x_1892 & ~n_35213;
assign n_35215 = ~x_1892 &  n_35213;
assign n_35216 = ~n_35214 & ~n_35215;
assign n_35217 =  x_1891 & ~n_24592;
assign n_35218 =  i_25 &  n_24592;
assign n_35219 = ~n_35217 & ~n_35218;
assign n_35220 =  x_1891 & ~n_35219;
assign n_35221 = ~x_1891 &  n_35219;
assign n_35222 = ~n_35220 & ~n_35221;
assign n_35223 =  x_1890 & ~n_24592;
assign n_35224 =  i_24 &  n_24592;
assign n_35225 = ~n_35223 & ~n_35224;
assign n_35226 =  x_1890 & ~n_35225;
assign n_35227 = ~x_1890 &  n_35225;
assign n_35228 = ~n_35226 & ~n_35227;
assign n_35229 =  x_1889 & ~n_24592;
assign n_35230 =  i_23 &  n_24592;
assign n_35231 = ~n_35229 & ~n_35230;
assign n_35232 =  x_1889 & ~n_35231;
assign n_35233 = ~x_1889 &  n_35231;
assign n_35234 = ~n_35232 & ~n_35233;
assign n_35235 =  x_1888 & ~n_24592;
assign n_35236 =  i_22 &  n_24592;
assign n_35237 = ~n_35235 & ~n_35236;
assign n_35238 =  x_1888 & ~n_35237;
assign n_35239 = ~x_1888 &  n_35237;
assign n_35240 = ~n_35238 & ~n_35239;
assign n_35241 =  x_1887 & ~n_24592;
assign n_35242 =  i_21 &  n_24592;
assign n_35243 = ~n_35241 & ~n_35242;
assign n_35244 =  x_1887 & ~n_35243;
assign n_35245 = ~x_1887 &  n_35243;
assign n_35246 = ~n_35244 & ~n_35245;
assign n_35247 =  x_1886 & ~n_24592;
assign n_35248 =  i_20 &  n_24592;
assign n_35249 = ~n_35247 & ~n_35248;
assign n_35250 =  x_1886 & ~n_35249;
assign n_35251 = ~x_1886 &  n_35249;
assign n_35252 = ~n_35250 & ~n_35251;
assign n_35253 =  x_1885 & ~n_24592;
assign n_35254 =  i_19 &  n_24592;
assign n_35255 = ~n_35253 & ~n_35254;
assign n_35256 =  x_1885 & ~n_35255;
assign n_35257 = ~x_1885 &  n_35255;
assign n_35258 = ~n_35256 & ~n_35257;
assign n_35259 =  x_1884 & ~n_24592;
assign n_35260 =  i_18 &  n_24592;
assign n_35261 = ~n_35259 & ~n_35260;
assign n_35262 =  x_1884 & ~n_35261;
assign n_35263 = ~x_1884 &  n_35261;
assign n_35264 = ~n_35262 & ~n_35263;
assign n_35265 =  x_1883 & ~n_24592;
assign n_35266 =  i_17 &  n_24592;
assign n_35267 = ~n_35265 & ~n_35266;
assign n_35268 =  x_1883 & ~n_35267;
assign n_35269 = ~x_1883 &  n_35267;
assign n_35270 = ~n_35268 & ~n_35269;
assign n_35271 =  x_1882 & ~n_24592;
assign n_35272 =  i_16 &  n_24592;
assign n_35273 = ~n_35271 & ~n_35272;
assign n_35274 =  x_1882 & ~n_35273;
assign n_35275 = ~x_1882 &  n_35273;
assign n_35276 = ~n_35274 & ~n_35275;
assign n_35277 =  x_1881 & ~n_24592;
assign n_35278 =  i_15 &  n_24592;
assign n_35279 = ~n_35277 & ~n_35278;
assign n_35280 =  x_1881 & ~n_35279;
assign n_35281 = ~x_1881 &  n_35279;
assign n_35282 = ~n_35280 & ~n_35281;
assign n_35283 =  x_1880 & ~n_24592;
assign n_35284 =  i_14 &  n_24592;
assign n_35285 = ~n_35283 & ~n_35284;
assign n_35286 =  x_1880 & ~n_35285;
assign n_35287 = ~x_1880 &  n_35285;
assign n_35288 = ~n_35286 & ~n_35287;
assign n_35289 =  x_1879 & ~n_24592;
assign n_35290 =  i_13 &  n_24592;
assign n_35291 = ~n_35289 & ~n_35290;
assign n_35292 =  x_1879 & ~n_35291;
assign n_35293 = ~x_1879 &  n_35291;
assign n_35294 = ~n_35292 & ~n_35293;
assign n_35295 =  x_1878 & ~n_24592;
assign n_35296 =  i_12 &  n_24592;
assign n_35297 = ~n_35295 & ~n_35296;
assign n_35298 =  x_1878 & ~n_35297;
assign n_35299 = ~x_1878 &  n_35297;
assign n_35300 = ~n_35298 & ~n_35299;
assign n_35301 =  x_1877 & ~n_24592;
assign n_35302 =  i_11 &  n_24592;
assign n_35303 = ~n_35301 & ~n_35302;
assign n_35304 =  x_1877 & ~n_35303;
assign n_35305 = ~x_1877 &  n_35303;
assign n_35306 = ~n_35304 & ~n_35305;
assign n_35307 =  x_1876 & ~n_24592;
assign n_35308 =  i_10 &  n_24592;
assign n_35309 = ~n_35307 & ~n_35308;
assign n_35310 =  x_1876 & ~n_35309;
assign n_35311 = ~x_1876 &  n_35309;
assign n_35312 = ~n_35310 & ~n_35311;
assign n_35313 =  x_1875 & ~n_24592;
assign n_35314 =  i_9 &  n_24592;
assign n_35315 = ~n_35313 & ~n_35314;
assign n_35316 =  x_1875 & ~n_35315;
assign n_35317 = ~x_1875 &  n_35315;
assign n_35318 = ~n_35316 & ~n_35317;
assign n_35319 =  x_1874 & ~n_24592;
assign n_35320 =  i_8 &  n_24592;
assign n_35321 = ~n_35319 & ~n_35320;
assign n_35322 =  x_1874 & ~n_35321;
assign n_35323 = ~x_1874 &  n_35321;
assign n_35324 = ~n_35322 & ~n_35323;
assign n_35325 =  x_1873 & ~n_24592;
assign n_35326 =  i_7 &  n_24592;
assign n_35327 = ~n_35325 & ~n_35326;
assign n_35328 =  x_1873 & ~n_35327;
assign n_35329 = ~x_1873 &  n_35327;
assign n_35330 = ~n_35328 & ~n_35329;
assign n_35331 =  x_1872 & ~n_24592;
assign n_35332 =  i_6 &  n_24592;
assign n_35333 = ~n_35331 & ~n_35332;
assign n_35334 =  x_1872 & ~n_35333;
assign n_35335 = ~x_1872 &  n_35333;
assign n_35336 = ~n_35334 & ~n_35335;
assign n_35337 =  x_1871 & ~n_24592;
assign n_35338 =  i_5 &  n_24592;
assign n_35339 = ~n_35337 & ~n_35338;
assign n_35340 =  x_1871 & ~n_35339;
assign n_35341 = ~x_1871 &  n_35339;
assign n_35342 = ~n_35340 & ~n_35341;
assign n_35343 =  x_1870 & ~n_24592;
assign n_35344 =  i_4 &  n_24592;
assign n_35345 = ~n_35343 & ~n_35344;
assign n_35346 =  x_1870 & ~n_35345;
assign n_35347 = ~x_1870 &  n_35345;
assign n_35348 = ~n_35346 & ~n_35347;
assign n_35349 =  x_1869 & ~n_24592;
assign n_35350 =  i_3 &  n_24592;
assign n_35351 = ~n_35349 & ~n_35350;
assign n_35352 =  x_1869 & ~n_35351;
assign n_35353 = ~x_1869 &  n_35351;
assign n_35354 = ~n_35352 & ~n_35353;
assign n_35355 =  x_1868 & ~n_24592;
assign n_35356 =  i_2 &  n_24592;
assign n_35357 = ~n_35355 & ~n_35356;
assign n_35358 =  x_1868 & ~n_35357;
assign n_35359 = ~x_1868 &  n_35357;
assign n_35360 = ~n_35358 & ~n_35359;
assign n_35361 =  x_1867 & ~n_24592;
assign n_35362 =  i_1 &  n_24592;
assign n_35363 = ~n_35361 & ~n_35362;
assign n_35364 =  x_1867 & ~n_35363;
assign n_35365 = ~x_1867 &  n_35363;
assign n_35366 = ~n_35364 & ~n_35365;
assign n_35367 =  x_1866 & ~n_25985;
assign n_35368 =  i_32 &  n_25985;
assign n_35369 = ~n_35367 & ~n_35368;
assign n_35370 =  x_1866 & ~n_35369;
assign n_35371 = ~x_1866 &  n_35369;
assign n_35372 = ~n_35370 & ~n_35371;
assign n_35373 =  x_1865 & ~n_25985;
assign n_35374 =  i_31 &  n_25985;
assign n_35375 = ~n_35373 & ~n_35374;
assign n_35376 =  x_1865 & ~n_35375;
assign n_35377 = ~x_1865 &  n_35375;
assign n_35378 = ~n_35376 & ~n_35377;
assign n_35379 =  x_1864 & ~n_25985;
assign n_35380 =  i_30 &  n_25985;
assign n_35381 = ~n_35379 & ~n_35380;
assign n_35382 =  x_1864 & ~n_35381;
assign n_35383 = ~x_1864 &  n_35381;
assign n_35384 = ~n_35382 & ~n_35383;
assign n_35385 =  x_1863 & ~n_25985;
assign n_35386 =  i_29 &  n_25985;
assign n_35387 = ~n_35385 & ~n_35386;
assign n_35388 =  x_1863 & ~n_35387;
assign n_35389 = ~x_1863 &  n_35387;
assign n_35390 = ~n_35388 & ~n_35389;
assign n_35391 =  x_1862 & ~n_25985;
assign n_35392 =  i_28 &  n_25985;
assign n_35393 = ~n_35391 & ~n_35392;
assign n_35394 =  x_1862 & ~n_35393;
assign n_35395 = ~x_1862 &  n_35393;
assign n_35396 = ~n_35394 & ~n_35395;
assign n_35397 =  x_1861 & ~n_25985;
assign n_35398 =  i_27 &  n_25985;
assign n_35399 = ~n_35397 & ~n_35398;
assign n_35400 =  x_1861 & ~n_35399;
assign n_35401 = ~x_1861 &  n_35399;
assign n_35402 = ~n_35400 & ~n_35401;
assign n_35403 =  x_1860 & ~n_25985;
assign n_35404 =  i_26 &  n_25985;
assign n_35405 = ~n_35403 & ~n_35404;
assign n_35406 =  x_1860 & ~n_35405;
assign n_35407 = ~x_1860 &  n_35405;
assign n_35408 = ~n_35406 & ~n_35407;
assign n_35409 =  x_1859 & ~n_25985;
assign n_35410 =  i_25 &  n_25985;
assign n_35411 = ~n_35409 & ~n_35410;
assign n_35412 =  x_1859 & ~n_35411;
assign n_35413 = ~x_1859 &  n_35411;
assign n_35414 = ~n_35412 & ~n_35413;
assign n_35415 =  x_1858 & ~n_25985;
assign n_35416 =  i_24 &  n_25985;
assign n_35417 = ~n_35415 & ~n_35416;
assign n_35418 =  x_1858 & ~n_35417;
assign n_35419 = ~x_1858 &  n_35417;
assign n_35420 = ~n_35418 & ~n_35419;
assign n_35421 =  x_1857 & ~n_25985;
assign n_35422 =  i_23 &  n_25985;
assign n_35423 = ~n_35421 & ~n_35422;
assign n_35424 =  x_1857 & ~n_35423;
assign n_35425 = ~x_1857 &  n_35423;
assign n_35426 = ~n_35424 & ~n_35425;
assign n_35427 =  x_1856 & ~n_25985;
assign n_35428 =  i_22 &  n_25985;
assign n_35429 = ~n_35427 & ~n_35428;
assign n_35430 =  x_1856 & ~n_35429;
assign n_35431 = ~x_1856 &  n_35429;
assign n_35432 = ~n_35430 & ~n_35431;
assign n_35433 =  x_1855 & ~n_25985;
assign n_35434 =  i_21 &  n_25985;
assign n_35435 = ~n_35433 & ~n_35434;
assign n_35436 =  x_1855 & ~n_35435;
assign n_35437 = ~x_1855 &  n_35435;
assign n_35438 = ~n_35436 & ~n_35437;
assign n_35439 =  x_1854 & ~n_25985;
assign n_35440 =  i_20 &  n_25985;
assign n_35441 = ~n_35439 & ~n_35440;
assign n_35442 =  x_1854 & ~n_35441;
assign n_35443 = ~x_1854 &  n_35441;
assign n_35444 = ~n_35442 & ~n_35443;
assign n_35445 =  x_1853 & ~n_25985;
assign n_35446 =  i_19 &  n_25985;
assign n_35447 = ~n_35445 & ~n_35446;
assign n_35448 =  x_1853 & ~n_35447;
assign n_35449 = ~x_1853 &  n_35447;
assign n_35450 = ~n_35448 & ~n_35449;
assign n_35451 =  x_1852 & ~n_25985;
assign n_35452 =  i_18 &  n_25985;
assign n_35453 = ~n_35451 & ~n_35452;
assign n_35454 =  x_1852 & ~n_35453;
assign n_35455 = ~x_1852 &  n_35453;
assign n_35456 = ~n_35454 & ~n_35455;
assign n_35457 =  x_1851 & ~n_25985;
assign n_35458 =  i_17 &  n_25985;
assign n_35459 = ~n_35457 & ~n_35458;
assign n_35460 =  x_1851 & ~n_35459;
assign n_35461 = ~x_1851 &  n_35459;
assign n_35462 = ~n_35460 & ~n_35461;
assign n_35463 =  x_1850 & ~n_25985;
assign n_35464 =  i_16 &  n_25985;
assign n_35465 = ~n_35463 & ~n_35464;
assign n_35466 =  x_1850 & ~n_35465;
assign n_35467 = ~x_1850 &  n_35465;
assign n_35468 = ~n_35466 & ~n_35467;
assign n_35469 =  x_1849 & ~n_25985;
assign n_35470 =  i_15 &  n_25985;
assign n_35471 = ~n_35469 & ~n_35470;
assign n_35472 =  x_1849 & ~n_35471;
assign n_35473 = ~x_1849 &  n_35471;
assign n_35474 = ~n_35472 & ~n_35473;
assign n_35475 =  x_1848 & ~n_25985;
assign n_35476 =  i_14 &  n_25985;
assign n_35477 = ~n_35475 & ~n_35476;
assign n_35478 =  x_1848 & ~n_35477;
assign n_35479 = ~x_1848 &  n_35477;
assign n_35480 = ~n_35478 & ~n_35479;
assign n_35481 =  x_1847 & ~n_25985;
assign n_35482 =  i_13 &  n_25985;
assign n_35483 = ~n_35481 & ~n_35482;
assign n_35484 =  x_1847 & ~n_35483;
assign n_35485 = ~x_1847 &  n_35483;
assign n_35486 = ~n_35484 & ~n_35485;
assign n_35487 =  x_1846 & ~n_25985;
assign n_35488 =  i_12 &  n_25985;
assign n_35489 = ~n_35487 & ~n_35488;
assign n_35490 =  x_1846 & ~n_35489;
assign n_35491 = ~x_1846 &  n_35489;
assign n_35492 = ~n_35490 & ~n_35491;
assign n_35493 =  x_1845 & ~n_25985;
assign n_35494 =  i_11 &  n_25985;
assign n_35495 = ~n_35493 & ~n_35494;
assign n_35496 =  x_1845 & ~n_35495;
assign n_35497 = ~x_1845 &  n_35495;
assign n_35498 = ~n_35496 & ~n_35497;
assign n_35499 =  x_1844 & ~n_25985;
assign n_35500 =  i_10 &  n_25985;
assign n_35501 = ~n_35499 & ~n_35500;
assign n_35502 =  x_1844 & ~n_35501;
assign n_35503 = ~x_1844 &  n_35501;
assign n_35504 = ~n_35502 & ~n_35503;
assign n_35505 =  x_1843 & ~n_25985;
assign n_35506 =  i_9 &  n_25985;
assign n_35507 = ~n_35505 & ~n_35506;
assign n_35508 =  x_1843 & ~n_35507;
assign n_35509 = ~x_1843 &  n_35507;
assign n_35510 = ~n_35508 & ~n_35509;
assign n_35511 =  x_1842 & ~n_25985;
assign n_35512 =  i_8 &  n_25985;
assign n_35513 = ~n_35511 & ~n_35512;
assign n_35514 =  x_1842 & ~n_35513;
assign n_35515 = ~x_1842 &  n_35513;
assign n_35516 = ~n_35514 & ~n_35515;
assign n_35517 =  x_1841 & ~n_25985;
assign n_35518 =  i_7 &  n_25985;
assign n_35519 = ~n_35517 & ~n_35518;
assign n_35520 =  x_1841 & ~n_35519;
assign n_35521 = ~x_1841 &  n_35519;
assign n_35522 = ~n_35520 & ~n_35521;
assign n_35523 =  x_1840 & ~n_25985;
assign n_35524 =  i_6 &  n_25985;
assign n_35525 = ~n_35523 & ~n_35524;
assign n_35526 =  x_1840 & ~n_35525;
assign n_35527 = ~x_1840 &  n_35525;
assign n_35528 = ~n_35526 & ~n_35527;
assign n_35529 =  x_1839 & ~n_25985;
assign n_35530 =  i_5 &  n_25985;
assign n_35531 = ~n_35529 & ~n_35530;
assign n_35532 =  x_1839 & ~n_35531;
assign n_35533 = ~x_1839 &  n_35531;
assign n_35534 = ~n_35532 & ~n_35533;
assign n_35535 =  x_1838 & ~n_25985;
assign n_35536 =  i_4 &  n_25985;
assign n_35537 = ~n_35535 & ~n_35536;
assign n_35538 =  x_1838 & ~n_35537;
assign n_35539 = ~x_1838 &  n_35537;
assign n_35540 = ~n_35538 & ~n_35539;
assign n_35541 =  x_1837 & ~n_25985;
assign n_35542 =  i_3 &  n_25985;
assign n_35543 = ~n_35541 & ~n_35542;
assign n_35544 =  x_1837 & ~n_35543;
assign n_35545 = ~x_1837 &  n_35543;
assign n_35546 = ~n_35544 & ~n_35545;
assign n_35547 =  x_1836 & ~n_25985;
assign n_35548 =  i_2 &  n_25985;
assign n_35549 = ~n_35547 & ~n_35548;
assign n_35550 =  x_1836 & ~n_35549;
assign n_35551 = ~x_1836 &  n_35549;
assign n_35552 = ~n_35550 & ~n_35551;
assign n_35553 =  x_1835 & ~n_25985;
assign n_35554 =  i_1 &  n_25985;
assign n_35555 = ~n_35553 & ~n_35554;
assign n_35556 =  x_1835 & ~n_35555;
assign n_35557 = ~x_1835 &  n_35555;
assign n_35558 = ~n_35556 & ~n_35557;
assign n_35559 = ~n_26262 & ~n_26436;
assign n_35560 =  x_1834 & ~n_26009;
assign n_35561 =  n_35559 & ~n_35560;
assign n_35562 =  x_1834 & ~n_35561;
assign n_35563 = ~x_1834 &  n_35561;
assign n_35564 = ~n_35562 & ~n_35563;
assign n_35565 = ~n_26009 &  n_35559;
assign n_35566 =  x_1833 &  n_35565;
assign n_35567 =  x_1833 &  n_35566;
assign n_35568 = ~x_1833 & ~n_35566;
assign n_35569 = ~n_35567 & ~n_35568;
assign n_35570 =  x_1832 &  n_35565;
assign n_35571 =  x_1832 &  n_35570;
assign n_35572 = ~x_1832 & ~n_35570;
assign n_35573 = ~n_35571 & ~n_35572;
assign n_35574 =  x_1831 &  n_35565;
assign n_35575 =  x_1831 &  n_35574;
assign n_35576 = ~x_1831 & ~n_35574;
assign n_35577 = ~n_35575 & ~n_35576;
assign n_35578 =  x_1830 &  n_35565;
assign n_35579 =  x_1830 &  n_35578;
assign n_35580 = ~x_1830 & ~n_35578;
assign n_35581 = ~n_35579 & ~n_35580;
assign n_35582 =  x_1829 &  n_35565;
assign n_35583 =  x_1829 &  n_35582;
assign n_35584 = ~x_1829 & ~n_35582;
assign n_35585 = ~n_35583 & ~n_35584;
assign n_35586 =  x_1828 &  n_35565;
assign n_35587 =  x_1828 &  n_35586;
assign n_35588 = ~x_1828 & ~n_35586;
assign n_35589 = ~n_35587 & ~n_35588;
assign n_35590 =  x_1827 &  n_35565;
assign n_35591 =  x_1827 &  n_35590;
assign n_35592 = ~x_1827 & ~n_35590;
assign n_35593 = ~n_35591 & ~n_35592;
assign n_35594 =  x_1826 &  n_35565;
assign n_35595 =  x_1826 &  n_35594;
assign n_35596 = ~x_1826 & ~n_35594;
assign n_35597 = ~n_35595 & ~n_35596;
assign n_35598 =  x_1825 &  n_35565;
assign n_35599 =  x_1825 &  n_35598;
assign n_35600 = ~x_1825 & ~n_35598;
assign n_35601 = ~n_35599 & ~n_35600;
assign n_35602 =  x_1824 &  n_35565;
assign n_35603 =  x_1824 &  n_35602;
assign n_35604 = ~x_1824 & ~n_35602;
assign n_35605 = ~n_35603 & ~n_35604;
assign n_35606 =  x_1823 &  n_35565;
assign n_35607 =  x_1823 &  n_35606;
assign n_35608 = ~x_1823 & ~n_35606;
assign n_35609 = ~n_35607 & ~n_35608;
assign n_35610 =  x_1822 &  n_35565;
assign n_35611 =  x_1822 &  n_35610;
assign n_35612 = ~x_1822 & ~n_35610;
assign n_35613 = ~n_35611 & ~n_35612;
assign n_35614 =  x_1821 &  n_35565;
assign n_35615 =  x_1821 &  n_35614;
assign n_35616 = ~x_1821 & ~n_35614;
assign n_35617 = ~n_35615 & ~n_35616;
assign n_35618 =  x_1820 &  n_35565;
assign n_35619 =  x_1820 &  n_35618;
assign n_35620 = ~x_1820 & ~n_35618;
assign n_35621 = ~n_35619 & ~n_35620;
assign n_35622 =  x_1819 &  n_35565;
assign n_35623 =  x_1819 &  n_35622;
assign n_35624 = ~x_1819 & ~n_35622;
assign n_35625 = ~n_35623 & ~n_35624;
assign n_35626 =  x_1818 &  n_35565;
assign n_35627 =  x_1818 &  n_35626;
assign n_35628 = ~x_1818 & ~n_35626;
assign n_35629 = ~n_35627 & ~n_35628;
assign n_35630 =  x_1817 &  n_35565;
assign n_35631 =  x_1817 &  n_35630;
assign n_35632 = ~x_1817 & ~n_35630;
assign n_35633 = ~n_35631 & ~n_35632;
assign n_35634 =  x_1816 &  n_35565;
assign n_35635 =  x_1816 &  n_35634;
assign n_35636 = ~x_1816 & ~n_35634;
assign n_35637 = ~n_35635 & ~n_35636;
assign n_35638 =  x_1815 &  n_35565;
assign n_35639 =  x_1815 &  n_35638;
assign n_35640 = ~x_1815 & ~n_35638;
assign n_35641 = ~n_35639 & ~n_35640;
assign n_35642 =  x_1814 &  n_35565;
assign n_35643 =  x_1814 &  n_35642;
assign n_35644 = ~x_1814 & ~n_35642;
assign n_35645 = ~n_35643 & ~n_35644;
assign n_35646 =  x_1813 &  n_35565;
assign n_35647 =  x_1813 &  n_35646;
assign n_35648 = ~x_1813 & ~n_35646;
assign n_35649 = ~n_35647 & ~n_35648;
assign n_35650 =  x_1812 &  n_35565;
assign n_35651 =  x_1812 &  n_35650;
assign n_35652 = ~x_1812 & ~n_35650;
assign n_35653 = ~n_35651 & ~n_35652;
assign n_35654 =  x_1811 &  n_35565;
assign n_35655 =  x_1811 &  n_35654;
assign n_35656 = ~x_1811 & ~n_35654;
assign n_35657 = ~n_35655 & ~n_35656;
assign n_35658 =  x_1810 &  n_35565;
assign n_35659 =  x_1810 &  n_35658;
assign n_35660 = ~x_1810 & ~n_35658;
assign n_35661 = ~n_35659 & ~n_35660;
assign n_35662 =  x_1809 &  n_35565;
assign n_35663 =  x_1809 &  n_35662;
assign n_35664 = ~x_1809 & ~n_35662;
assign n_35665 = ~n_35663 & ~n_35664;
assign n_35666 =  x_1808 &  n_35565;
assign n_35667 =  x_1808 &  n_35666;
assign n_35668 = ~x_1808 & ~n_35666;
assign n_35669 = ~n_35667 & ~n_35668;
assign n_35670 =  x_1807 &  n_35565;
assign n_35671 =  x_1807 &  n_35670;
assign n_35672 = ~x_1807 & ~n_35670;
assign n_35673 = ~n_35671 & ~n_35672;
assign n_35674 =  x_1806 &  n_35565;
assign n_35675 =  x_1806 &  n_35674;
assign n_35676 = ~x_1806 & ~n_35674;
assign n_35677 = ~n_35675 & ~n_35676;
assign n_35678 =  x_1805 &  n_35565;
assign n_35679 =  x_1805 &  n_35678;
assign n_35680 = ~x_1805 & ~n_35678;
assign n_35681 = ~n_35679 & ~n_35680;
assign n_35682 =  x_1804 &  n_35565;
assign n_35683 =  x_1804 &  n_35682;
assign n_35684 = ~x_1804 & ~n_35682;
assign n_35685 = ~n_35683 & ~n_35684;
assign n_35686 =  x_1803 &  n_35565;
assign n_35687 =  x_1803 &  n_35686;
assign n_35688 = ~x_1803 & ~n_35686;
assign n_35689 = ~n_35687 & ~n_35688;
assign n_35690 =  x_1802 & ~n_27955;
assign n_35691 =  x_1802 &  n_35690;
assign n_35692 = ~x_1802 & ~n_35690;
assign n_35693 = ~n_35691 & ~n_35692;
assign n_35694 =  x_1801 & ~n_27955;
assign n_35695 =  x_1801 &  n_35694;
assign n_35696 = ~x_1801 & ~n_35694;
assign n_35697 = ~n_35695 & ~n_35696;
assign n_35698 =  x_1800 & ~n_27955;
assign n_35699 =  x_1800 &  n_35698;
assign n_35700 = ~x_1800 & ~n_35698;
assign n_35701 = ~n_35699 & ~n_35700;
assign n_35702 =  x_1799 & ~n_27955;
assign n_35703 =  x_1799 &  n_35702;
assign n_35704 = ~x_1799 & ~n_35702;
assign n_35705 = ~n_35703 & ~n_35704;
assign n_35706 =  x_1798 & ~n_27955;
assign n_35707 =  x_1798 &  n_35706;
assign n_35708 = ~x_1798 & ~n_35706;
assign n_35709 = ~n_35707 & ~n_35708;
assign n_35710 =  x_1797 & ~n_27955;
assign n_35711 =  x_1797 &  n_35710;
assign n_35712 = ~x_1797 & ~n_35710;
assign n_35713 = ~n_35711 & ~n_35712;
assign n_35714 =  x_1796 & ~n_27955;
assign n_35715 =  x_1796 &  n_35714;
assign n_35716 = ~x_1796 & ~n_35714;
assign n_35717 = ~n_35715 & ~n_35716;
assign n_35718 =  x_1795 & ~n_27955;
assign n_35719 =  x_1795 &  n_35718;
assign n_35720 = ~x_1795 & ~n_35718;
assign n_35721 = ~n_35719 & ~n_35720;
assign n_35722 =  x_1794 & ~n_27955;
assign n_35723 =  x_1794 &  n_35722;
assign n_35724 = ~x_1794 & ~n_35722;
assign n_35725 = ~n_35723 & ~n_35724;
assign n_35726 =  x_1793 & ~n_27955;
assign n_35727 =  x_1793 &  n_35726;
assign n_35728 = ~x_1793 & ~n_35726;
assign n_35729 = ~n_35727 & ~n_35728;
assign n_35730 =  x_1792 & ~n_27955;
assign n_35731 =  x_1792 &  n_35730;
assign n_35732 = ~x_1792 & ~n_35730;
assign n_35733 = ~n_35731 & ~n_35732;
assign n_35734 =  x_1791 & ~n_27955;
assign n_35735 =  x_1791 &  n_35734;
assign n_35736 = ~x_1791 & ~n_35734;
assign n_35737 = ~n_35735 & ~n_35736;
assign n_35738 =  x_1790 & ~n_27955;
assign n_35739 =  x_1790 &  n_35738;
assign n_35740 = ~x_1790 & ~n_35738;
assign n_35741 = ~n_35739 & ~n_35740;
assign n_35742 =  x_1789 & ~n_27955;
assign n_35743 =  x_1789 &  n_35742;
assign n_35744 = ~x_1789 & ~n_35742;
assign n_35745 = ~n_35743 & ~n_35744;
assign n_35746 =  x_1788 & ~n_27955;
assign n_35747 =  x_1788 &  n_35746;
assign n_35748 = ~x_1788 & ~n_35746;
assign n_35749 = ~n_35747 & ~n_35748;
assign n_35750 =  x_1787 & ~n_27955;
assign n_35751 =  x_1787 &  n_35750;
assign n_35752 = ~x_1787 & ~n_35750;
assign n_35753 = ~n_35751 & ~n_35752;
assign n_35754 =  x_1786 & ~n_27955;
assign n_35755 =  x_1786 &  n_35754;
assign n_35756 = ~x_1786 & ~n_35754;
assign n_35757 = ~n_35755 & ~n_35756;
assign n_35758 =  x_1785 & ~n_27955;
assign n_35759 =  x_1785 &  n_35758;
assign n_35760 = ~x_1785 & ~n_35758;
assign n_35761 = ~n_35759 & ~n_35760;
assign n_35762 =  x_1784 & ~n_27955;
assign n_35763 =  x_1784 &  n_35762;
assign n_35764 = ~x_1784 & ~n_35762;
assign n_35765 = ~n_35763 & ~n_35764;
assign n_35766 =  x_1783 & ~n_27955;
assign n_35767 =  x_1783 &  n_35766;
assign n_35768 = ~x_1783 & ~n_35766;
assign n_35769 = ~n_35767 & ~n_35768;
assign n_35770 =  x_1782 & ~n_27955;
assign n_35771 =  x_1782 &  n_35770;
assign n_35772 = ~x_1782 & ~n_35770;
assign n_35773 = ~n_35771 & ~n_35772;
assign n_35774 =  x_1781 & ~n_27955;
assign n_35775 =  x_1781 &  n_35774;
assign n_35776 = ~x_1781 & ~n_35774;
assign n_35777 = ~n_35775 & ~n_35776;
assign n_35778 =  x_1780 & ~n_27955;
assign n_35779 =  x_1780 &  n_35778;
assign n_35780 = ~x_1780 & ~n_35778;
assign n_35781 = ~n_35779 & ~n_35780;
assign n_35782 =  x_1779 & ~n_27955;
assign n_35783 =  x_1779 &  n_35782;
assign n_35784 = ~x_1779 & ~n_35782;
assign n_35785 = ~n_35783 & ~n_35784;
assign n_35786 =  x_1778 & ~n_27955;
assign n_35787 =  x_1778 &  n_35786;
assign n_35788 = ~x_1778 & ~n_35786;
assign n_35789 = ~n_35787 & ~n_35788;
assign n_35790 =  x_1777 & ~n_27955;
assign n_35791 =  x_1777 &  n_35790;
assign n_35792 = ~x_1777 & ~n_35790;
assign n_35793 = ~n_35791 & ~n_35792;
assign n_35794 =  x_1776 & ~n_27955;
assign n_35795 =  x_1776 &  n_35794;
assign n_35796 = ~x_1776 & ~n_35794;
assign n_35797 = ~n_35795 & ~n_35796;
assign n_35798 =  x_1775 & ~n_27955;
assign n_35799 =  x_1775 &  n_35798;
assign n_35800 = ~x_1775 & ~n_35798;
assign n_35801 = ~n_35799 & ~n_35800;
assign n_35802 =  x_1774 & ~n_27955;
assign n_35803 =  x_1774 &  n_35802;
assign n_35804 = ~x_1774 & ~n_35802;
assign n_35805 = ~n_35803 & ~n_35804;
assign n_35806 =  x_1773 & ~n_27955;
assign n_35807 =  x_1773 &  n_35806;
assign n_35808 = ~x_1773 & ~n_35806;
assign n_35809 = ~n_35807 & ~n_35808;
assign n_35810 =  x_1772 & ~n_27955;
assign n_35811 =  x_1772 &  n_35810;
assign n_35812 = ~x_1772 & ~n_35810;
assign n_35813 = ~n_35811 & ~n_35812;
assign n_35814 =  x_1771 & ~n_27955;
assign n_35815 =  x_1771 &  n_35814;
assign n_35816 = ~x_1771 & ~n_35814;
assign n_35817 = ~n_35815 & ~n_35816;
assign n_35818 =  x_1770 & ~n_23856;
assign n_35819 =  x_874 &  n_23856;
assign n_35820 = ~n_35818 & ~n_35819;
assign n_35821 =  x_1770 & ~n_35820;
assign n_35822 = ~x_1770 &  n_35820;
assign n_35823 = ~n_35821 & ~n_35822;
assign n_35824 =  x_1769 & ~n_23856;
assign n_35825 =  x_873 &  n_23856;
assign n_35826 = ~n_35824 & ~n_35825;
assign n_35827 =  x_1769 & ~n_35826;
assign n_35828 = ~x_1769 &  n_35826;
assign n_35829 = ~n_35827 & ~n_35828;
assign n_35830 =  x_1768 & ~n_23856;
assign n_35831 =  x_872 &  n_23856;
assign n_35832 = ~n_35830 & ~n_35831;
assign n_35833 =  x_1768 & ~n_35832;
assign n_35834 = ~x_1768 &  n_35832;
assign n_35835 = ~n_35833 & ~n_35834;
assign n_35836 =  x_1767 & ~n_23856;
assign n_35837 =  x_871 &  n_23856;
assign n_35838 = ~n_35836 & ~n_35837;
assign n_35839 =  x_1767 & ~n_35838;
assign n_35840 = ~x_1767 &  n_35838;
assign n_35841 = ~n_35839 & ~n_35840;
assign n_35842 =  x_1766 & ~n_23856;
assign n_35843 =  x_870 &  n_23856;
assign n_35844 = ~n_35842 & ~n_35843;
assign n_35845 =  x_1766 & ~n_35844;
assign n_35846 = ~x_1766 &  n_35844;
assign n_35847 = ~n_35845 & ~n_35846;
assign n_35848 =  x_1765 & ~n_23856;
assign n_35849 =  x_869 &  n_23856;
assign n_35850 = ~n_35848 & ~n_35849;
assign n_35851 =  x_1765 & ~n_35850;
assign n_35852 = ~x_1765 &  n_35850;
assign n_35853 = ~n_35851 & ~n_35852;
assign n_35854 =  x_1764 & ~n_23856;
assign n_35855 =  x_868 &  n_23856;
assign n_35856 = ~n_35854 & ~n_35855;
assign n_35857 =  x_1764 & ~n_35856;
assign n_35858 = ~x_1764 &  n_35856;
assign n_35859 = ~n_35857 & ~n_35858;
assign n_35860 =  x_1763 & ~n_23856;
assign n_35861 =  x_867 &  n_23856;
assign n_35862 = ~n_35860 & ~n_35861;
assign n_35863 =  x_1763 & ~n_35862;
assign n_35864 = ~x_1763 &  n_35862;
assign n_35865 = ~n_35863 & ~n_35864;
assign n_35866 =  x_1762 & ~n_23856;
assign n_35867 =  x_866 &  n_23856;
assign n_35868 = ~n_35866 & ~n_35867;
assign n_35869 =  x_1762 & ~n_35868;
assign n_35870 = ~x_1762 &  n_35868;
assign n_35871 = ~n_35869 & ~n_35870;
assign n_35872 =  x_1761 & ~n_23856;
assign n_35873 =  x_865 &  n_23856;
assign n_35874 = ~n_35872 & ~n_35873;
assign n_35875 =  x_1761 & ~n_35874;
assign n_35876 = ~x_1761 &  n_35874;
assign n_35877 = ~n_35875 & ~n_35876;
assign n_35878 =  x_1760 & ~n_23856;
assign n_35879 =  x_864 &  n_23856;
assign n_35880 = ~n_35878 & ~n_35879;
assign n_35881 =  x_1760 & ~n_35880;
assign n_35882 = ~x_1760 &  n_35880;
assign n_35883 = ~n_35881 & ~n_35882;
assign n_35884 =  x_1759 & ~n_23856;
assign n_35885 =  x_863 &  n_23856;
assign n_35886 = ~n_35884 & ~n_35885;
assign n_35887 =  x_1759 & ~n_35886;
assign n_35888 = ~x_1759 &  n_35886;
assign n_35889 = ~n_35887 & ~n_35888;
assign n_35890 =  x_1758 & ~n_23856;
assign n_35891 =  x_862 &  n_23856;
assign n_35892 = ~n_35890 & ~n_35891;
assign n_35893 =  x_1758 & ~n_35892;
assign n_35894 = ~x_1758 &  n_35892;
assign n_35895 = ~n_35893 & ~n_35894;
assign n_35896 =  x_1757 & ~n_23856;
assign n_35897 =  x_861 &  n_23856;
assign n_35898 = ~n_35896 & ~n_35897;
assign n_35899 =  x_1757 & ~n_35898;
assign n_35900 = ~x_1757 &  n_35898;
assign n_35901 = ~n_35899 & ~n_35900;
assign n_35902 =  x_1756 & ~n_23856;
assign n_35903 =  x_860 &  n_23856;
assign n_35904 = ~n_35902 & ~n_35903;
assign n_35905 =  x_1756 & ~n_35904;
assign n_35906 = ~x_1756 &  n_35904;
assign n_35907 = ~n_35905 & ~n_35906;
assign n_35908 =  x_1755 & ~n_23856;
assign n_35909 =  x_859 &  n_23856;
assign n_35910 = ~n_35908 & ~n_35909;
assign n_35911 =  x_1755 & ~n_35910;
assign n_35912 = ~x_1755 &  n_35910;
assign n_35913 = ~n_35911 & ~n_35912;
assign n_35914 =  x_1754 & ~n_23856;
assign n_35915 =  x_858 &  n_23856;
assign n_35916 = ~n_35914 & ~n_35915;
assign n_35917 =  x_1754 & ~n_35916;
assign n_35918 = ~x_1754 &  n_35916;
assign n_35919 = ~n_35917 & ~n_35918;
assign n_35920 =  x_1753 & ~n_23856;
assign n_35921 =  x_857 &  n_23856;
assign n_35922 = ~n_35920 & ~n_35921;
assign n_35923 =  x_1753 & ~n_35922;
assign n_35924 = ~x_1753 &  n_35922;
assign n_35925 = ~n_35923 & ~n_35924;
assign n_35926 =  x_1752 & ~n_23856;
assign n_35927 =  x_856 &  n_23856;
assign n_35928 = ~n_35926 & ~n_35927;
assign n_35929 =  x_1752 & ~n_35928;
assign n_35930 = ~x_1752 &  n_35928;
assign n_35931 = ~n_35929 & ~n_35930;
assign n_35932 =  x_1751 & ~n_23856;
assign n_35933 =  x_855 &  n_23856;
assign n_35934 = ~n_35932 & ~n_35933;
assign n_35935 =  x_1751 & ~n_35934;
assign n_35936 = ~x_1751 &  n_35934;
assign n_35937 = ~n_35935 & ~n_35936;
assign n_35938 =  x_1750 & ~n_23856;
assign n_35939 =  x_854 &  n_23856;
assign n_35940 = ~n_35938 & ~n_35939;
assign n_35941 =  x_1750 & ~n_35940;
assign n_35942 = ~x_1750 &  n_35940;
assign n_35943 = ~n_35941 & ~n_35942;
assign n_35944 =  x_1749 & ~n_23856;
assign n_35945 =  x_853 &  n_23856;
assign n_35946 = ~n_35944 & ~n_35945;
assign n_35947 =  x_1749 & ~n_35946;
assign n_35948 = ~x_1749 &  n_35946;
assign n_35949 = ~n_35947 & ~n_35948;
assign n_35950 =  x_1748 & ~n_23856;
assign n_35951 =  x_852 &  n_23856;
assign n_35952 = ~n_35950 & ~n_35951;
assign n_35953 =  x_1748 & ~n_35952;
assign n_35954 = ~x_1748 &  n_35952;
assign n_35955 = ~n_35953 & ~n_35954;
assign n_35956 =  x_1747 & ~n_23856;
assign n_35957 =  x_851 &  n_23856;
assign n_35958 = ~n_35956 & ~n_35957;
assign n_35959 =  x_1747 & ~n_35958;
assign n_35960 = ~x_1747 &  n_35958;
assign n_35961 = ~n_35959 & ~n_35960;
assign n_35962 =  x_1746 & ~n_23856;
assign n_35963 =  x_850 &  n_23856;
assign n_35964 = ~n_35962 & ~n_35963;
assign n_35965 =  x_1746 & ~n_35964;
assign n_35966 = ~x_1746 &  n_35964;
assign n_35967 = ~n_35965 & ~n_35966;
assign n_35968 =  x_1745 & ~n_23856;
assign n_35969 =  x_849 &  n_23856;
assign n_35970 = ~n_35968 & ~n_35969;
assign n_35971 =  x_1745 & ~n_35970;
assign n_35972 = ~x_1745 &  n_35970;
assign n_35973 = ~n_35971 & ~n_35972;
assign n_35974 =  x_1744 & ~n_23856;
assign n_35975 =  x_848 &  n_23856;
assign n_35976 = ~n_35974 & ~n_35975;
assign n_35977 =  x_1744 & ~n_35976;
assign n_35978 = ~x_1744 &  n_35976;
assign n_35979 = ~n_35977 & ~n_35978;
assign n_35980 =  x_1743 & ~n_23856;
assign n_35981 =  x_847 &  n_23856;
assign n_35982 = ~n_35980 & ~n_35981;
assign n_35983 =  x_1743 & ~n_35982;
assign n_35984 = ~x_1743 &  n_35982;
assign n_35985 = ~n_35983 & ~n_35984;
assign n_35986 =  x_1742 & ~n_23856;
assign n_35987 =  x_846 &  n_23856;
assign n_35988 = ~n_35986 & ~n_35987;
assign n_35989 =  x_1742 & ~n_35988;
assign n_35990 = ~x_1742 &  n_35988;
assign n_35991 = ~n_35989 & ~n_35990;
assign n_35992 =  x_1741 & ~n_23856;
assign n_35993 =  x_845 &  n_23856;
assign n_35994 = ~n_35992 & ~n_35993;
assign n_35995 =  x_1741 & ~n_35994;
assign n_35996 = ~x_1741 &  n_35994;
assign n_35997 = ~n_35995 & ~n_35996;
assign n_35998 =  x_1740 & ~n_23856;
assign n_35999 =  x_844 &  n_23856;
assign n_36000 = ~n_35998 & ~n_35999;
assign n_36001 =  x_1740 & ~n_36000;
assign n_36002 = ~x_1740 &  n_36000;
assign n_36003 = ~n_36001 & ~n_36002;
assign n_36004 =  x_1739 & ~n_23856;
assign n_36005 =  x_1739 &  n_36004;
assign n_36006 = ~x_1739 & ~n_36004;
assign n_36007 = ~n_36005 & ~n_36006;
assign n_36008 = ~x_38 &  n_26264;
assign n_36009 = ~n_27730 & ~n_36008;
assign n_36010 =  i_32 & ~n_36009;
assign n_36011 =  x_1738 &  n_36009;
assign n_36012 = ~n_36010 & ~n_36011;
assign n_36013 =  x_1738 & ~n_36012;
assign n_36014 = ~x_1738 &  n_36012;
assign n_36015 = ~n_36013 & ~n_36014;
assign n_36016 =  i_31 & ~n_36009;
assign n_36017 =  x_1737 &  n_36009;
assign n_36018 = ~n_36016 & ~n_36017;
assign n_36019 =  x_1737 & ~n_36018;
assign n_36020 = ~x_1737 &  n_36018;
assign n_36021 = ~n_36019 & ~n_36020;
assign n_36022 =  i_30 & ~n_36009;
assign n_36023 =  x_1736 &  n_36009;
assign n_36024 = ~n_36022 & ~n_36023;
assign n_36025 =  x_1736 & ~n_36024;
assign n_36026 = ~x_1736 &  n_36024;
assign n_36027 = ~n_36025 & ~n_36026;
assign n_36028 =  i_29 & ~n_36009;
assign n_36029 =  x_1735 &  n_36009;
assign n_36030 = ~n_36028 & ~n_36029;
assign n_36031 =  x_1735 & ~n_36030;
assign n_36032 = ~x_1735 &  n_36030;
assign n_36033 = ~n_36031 & ~n_36032;
assign n_36034 =  i_28 & ~n_36009;
assign n_36035 =  x_1734 &  n_36009;
assign n_36036 = ~n_36034 & ~n_36035;
assign n_36037 =  x_1734 & ~n_36036;
assign n_36038 = ~x_1734 &  n_36036;
assign n_36039 = ~n_36037 & ~n_36038;
assign n_36040 =  i_27 & ~n_36009;
assign n_36041 =  x_1733 &  n_36009;
assign n_36042 = ~n_36040 & ~n_36041;
assign n_36043 =  x_1733 & ~n_36042;
assign n_36044 = ~x_1733 &  n_36042;
assign n_36045 = ~n_36043 & ~n_36044;
assign n_36046 =  i_26 & ~n_36009;
assign n_36047 =  x_1732 &  n_36009;
assign n_36048 = ~n_36046 & ~n_36047;
assign n_36049 =  x_1732 & ~n_36048;
assign n_36050 = ~x_1732 &  n_36048;
assign n_36051 = ~n_36049 & ~n_36050;
assign n_36052 =  i_25 & ~n_36009;
assign n_36053 =  x_1731 &  n_36009;
assign n_36054 = ~n_36052 & ~n_36053;
assign n_36055 =  x_1731 & ~n_36054;
assign n_36056 = ~x_1731 &  n_36054;
assign n_36057 = ~n_36055 & ~n_36056;
assign n_36058 =  i_24 & ~n_36009;
assign n_36059 =  x_1730 &  n_36009;
assign n_36060 = ~n_36058 & ~n_36059;
assign n_36061 =  x_1730 & ~n_36060;
assign n_36062 = ~x_1730 &  n_36060;
assign n_36063 = ~n_36061 & ~n_36062;
assign n_36064 =  i_23 & ~n_36009;
assign n_36065 =  x_1729 &  n_36009;
assign n_36066 = ~n_36064 & ~n_36065;
assign n_36067 =  x_1729 & ~n_36066;
assign n_36068 = ~x_1729 &  n_36066;
assign n_36069 = ~n_36067 & ~n_36068;
assign n_36070 =  i_22 & ~n_36009;
assign n_36071 =  x_1728 &  n_36009;
assign n_36072 = ~n_36070 & ~n_36071;
assign n_36073 =  x_1728 & ~n_36072;
assign n_36074 = ~x_1728 &  n_36072;
assign n_36075 = ~n_36073 & ~n_36074;
assign n_36076 =  i_21 & ~n_36009;
assign n_36077 =  x_1727 &  n_36009;
assign n_36078 = ~n_36076 & ~n_36077;
assign n_36079 =  x_1727 & ~n_36078;
assign n_36080 = ~x_1727 &  n_36078;
assign n_36081 = ~n_36079 & ~n_36080;
assign n_36082 =  i_20 & ~n_36009;
assign n_36083 =  x_1726 &  n_36009;
assign n_36084 = ~n_36082 & ~n_36083;
assign n_36085 =  x_1726 & ~n_36084;
assign n_36086 = ~x_1726 &  n_36084;
assign n_36087 = ~n_36085 & ~n_36086;
assign n_36088 =  i_19 & ~n_36009;
assign n_36089 =  x_1725 &  n_36009;
assign n_36090 = ~n_36088 & ~n_36089;
assign n_36091 =  x_1725 & ~n_36090;
assign n_36092 = ~x_1725 &  n_36090;
assign n_36093 = ~n_36091 & ~n_36092;
assign n_36094 =  i_18 & ~n_36009;
assign n_36095 =  x_1724 &  n_36009;
assign n_36096 = ~n_36094 & ~n_36095;
assign n_36097 =  x_1724 & ~n_36096;
assign n_36098 = ~x_1724 &  n_36096;
assign n_36099 = ~n_36097 & ~n_36098;
assign n_36100 =  i_17 & ~n_36009;
assign n_36101 =  x_1723 &  n_36009;
assign n_36102 = ~n_36100 & ~n_36101;
assign n_36103 =  x_1723 & ~n_36102;
assign n_36104 = ~x_1723 &  n_36102;
assign n_36105 = ~n_36103 & ~n_36104;
assign n_36106 =  i_16 & ~n_36009;
assign n_36107 =  x_1722 &  n_36009;
assign n_36108 = ~n_36106 & ~n_36107;
assign n_36109 =  x_1722 & ~n_36108;
assign n_36110 = ~x_1722 &  n_36108;
assign n_36111 = ~n_36109 & ~n_36110;
assign n_36112 =  i_15 & ~n_36009;
assign n_36113 =  x_1721 &  n_36009;
assign n_36114 = ~n_36112 & ~n_36113;
assign n_36115 =  x_1721 & ~n_36114;
assign n_36116 = ~x_1721 &  n_36114;
assign n_36117 = ~n_36115 & ~n_36116;
assign n_36118 =  i_14 & ~n_36009;
assign n_36119 =  x_1720 &  n_36009;
assign n_36120 = ~n_36118 & ~n_36119;
assign n_36121 =  x_1720 & ~n_36120;
assign n_36122 = ~x_1720 &  n_36120;
assign n_36123 = ~n_36121 & ~n_36122;
assign n_36124 =  i_13 & ~n_36009;
assign n_36125 =  x_1719 &  n_36009;
assign n_36126 = ~n_36124 & ~n_36125;
assign n_36127 =  x_1719 & ~n_36126;
assign n_36128 = ~x_1719 &  n_36126;
assign n_36129 = ~n_36127 & ~n_36128;
assign n_36130 =  i_12 & ~n_36009;
assign n_36131 =  x_1718 &  n_36009;
assign n_36132 = ~n_36130 & ~n_36131;
assign n_36133 =  x_1718 & ~n_36132;
assign n_36134 = ~x_1718 &  n_36132;
assign n_36135 = ~n_36133 & ~n_36134;
assign n_36136 =  i_11 & ~n_36009;
assign n_36137 =  x_1717 &  n_36009;
assign n_36138 = ~n_36136 & ~n_36137;
assign n_36139 =  x_1717 & ~n_36138;
assign n_36140 = ~x_1717 &  n_36138;
assign n_36141 = ~n_36139 & ~n_36140;
assign n_36142 =  i_10 & ~n_36009;
assign n_36143 =  x_1716 &  n_36009;
assign n_36144 = ~n_36142 & ~n_36143;
assign n_36145 =  x_1716 & ~n_36144;
assign n_36146 = ~x_1716 &  n_36144;
assign n_36147 = ~n_36145 & ~n_36146;
assign n_36148 =  i_9 & ~n_36009;
assign n_36149 =  x_1715 &  n_36009;
assign n_36150 = ~n_36148 & ~n_36149;
assign n_36151 =  x_1715 & ~n_36150;
assign n_36152 = ~x_1715 &  n_36150;
assign n_36153 = ~n_36151 & ~n_36152;
assign n_36154 =  i_8 & ~n_36009;
assign n_36155 =  x_1714 &  n_36009;
assign n_36156 = ~n_36154 & ~n_36155;
assign n_36157 =  x_1714 & ~n_36156;
assign n_36158 = ~x_1714 &  n_36156;
assign n_36159 = ~n_36157 & ~n_36158;
assign n_36160 =  i_7 & ~n_36009;
assign n_36161 =  x_1713 &  n_36009;
assign n_36162 = ~n_36160 & ~n_36161;
assign n_36163 =  x_1713 & ~n_36162;
assign n_36164 = ~x_1713 &  n_36162;
assign n_36165 = ~n_36163 & ~n_36164;
assign n_36166 =  i_6 & ~n_36009;
assign n_36167 =  x_1712 &  n_36009;
assign n_36168 = ~n_36166 & ~n_36167;
assign n_36169 =  x_1712 & ~n_36168;
assign n_36170 = ~x_1712 &  n_36168;
assign n_36171 = ~n_36169 & ~n_36170;
assign n_36172 =  i_5 & ~n_36009;
assign n_36173 =  x_1711 &  n_36009;
assign n_36174 = ~n_36172 & ~n_36173;
assign n_36175 =  x_1711 & ~n_36174;
assign n_36176 = ~x_1711 &  n_36174;
assign n_36177 = ~n_36175 & ~n_36176;
assign n_36178 =  i_4 & ~n_36009;
assign n_36179 =  x_1710 &  n_36009;
assign n_36180 = ~n_36178 & ~n_36179;
assign n_36181 =  x_1710 & ~n_36180;
assign n_36182 = ~x_1710 &  n_36180;
assign n_36183 = ~n_36181 & ~n_36182;
assign n_36184 =  i_3 & ~n_36009;
assign n_36185 =  x_1709 &  n_36009;
assign n_36186 = ~n_36184 & ~n_36185;
assign n_36187 =  x_1709 & ~n_36186;
assign n_36188 = ~x_1709 &  n_36186;
assign n_36189 = ~n_36187 & ~n_36188;
assign n_36190 =  i_2 & ~n_36009;
assign n_36191 =  x_1708 &  n_36009;
assign n_36192 = ~n_36190 & ~n_36191;
assign n_36193 =  x_1708 & ~n_36192;
assign n_36194 = ~x_1708 &  n_36192;
assign n_36195 = ~n_36193 & ~n_36194;
assign n_36196 =  i_1 & ~n_36009;
assign n_36197 =  x_1707 &  n_36009;
assign n_36198 = ~n_36196 & ~n_36197;
assign n_36199 =  x_1707 & ~n_36198;
assign n_36200 = ~x_1707 &  n_36198;
assign n_36201 = ~n_36199 & ~n_36200;
assign n_36202 = ~n_23251 & ~n_25975;
assign n_36203 =  i_32 & ~n_36202;
assign n_36204 =  x_1706 &  n_36202;
assign n_36205 = ~n_36203 & ~n_36204;
assign n_36206 =  x_1706 & ~n_36205;
assign n_36207 = ~x_1706 &  n_36205;
assign n_36208 = ~n_36206 & ~n_36207;
assign n_36209 =  i_31 & ~n_36202;
assign n_36210 =  x_1705 &  n_36202;
assign n_36211 = ~n_36209 & ~n_36210;
assign n_36212 =  x_1705 & ~n_36211;
assign n_36213 = ~x_1705 &  n_36211;
assign n_36214 = ~n_36212 & ~n_36213;
assign n_36215 =  i_30 & ~n_36202;
assign n_36216 =  x_1704 &  n_36202;
assign n_36217 = ~n_36215 & ~n_36216;
assign n_36218 =  x_1704 & ~n_36217;
assign n_36219 = ~x_1704 &  n_36217;
assign n_36220 = ~n_36218 & ~n_36219;
assign n_36221 =  i_29 & ~n_36202;
assign n_36222 =  x_1703 &  n_36202;
assign n_36223 = ~n_36221 & ~n_36222;
assign n_36224 =  x_1703 & ~n_36223;
assign n_36225 = ~x_1703 &  n_36223;
assign n_36226 = ~n_36224 & ~n_36225;
assign n_36227 =  i_28 & ~n_36202;
assign n_36228 =  x_1702 &  n_36202;
assign n_36229 = ~n_36227 & ~n_36228;
assign n_36230 =  x_1702 & ~n_36229;
assign n_36231 = ~x_1702 &  n_36229;
assign n_36232 = ~n_36230 & ~n_36231;
assign n_36233 =  i_27 & ~n_36202;
assign n_36234 =  x_1701 &  n_36202;
assign n_36235 = ~n_36233 & ~n_36234;
assign n_36236 =  x_1701 & ~n_36235;
assign n_36237 = ~x_1701 &  n_36235;
assign n_36238 = ~n_36236 & ~n_36237;
assign n_36239 =  i_26 & ~n_36202;
assign n_36240 =  x_1700 &  n_36202;
assign n_36241 = ~n_36239 & ~n_36240;
assign n_36242 =  x_1700 & ~n_36241;
assign n_36243 = ~x_1700 &  n_36241;
assign n_36244 = ~n_36242 & ~n_36243;
assign n_36245 =  i_25 & ~n_36202;
assign n_36246 =  x_1699 &  n_36202;
assign n_36247 = ~n_36245 & ~n_36246;
assign n_36248 =  x_1699 & ~n_36247;
assign n_36249 = ~x_1699 &  n_36247;
assign n_36250 = ~n_36248 & ~n_36249;
assign n_36251 =  i_24 & ~n_36202;
assign n_36252 =  x_1698 &  n_36202;
assign n_36253 = ~n_36251 & ~n_36252;
assign n_36254 =  x_1698 & ~n_36253;
assign n_36255 = ~x_1698 &  n_36253;
assign n_36256 = ~n_36254 & ~n_36255;
assign n_36257 =  i_23 & ~n_36202;
assign n_36258 =  x_1697 &  n_36202;
assign n_36259 = ~n_36257 & ~n_36258;
assign n_36260 =  x_1697 & ~n_36259;
assign n_36261 = ~x_1697 &  n_36259;
assign n_36262 = ~n_36260 & ~n_36261;
assign n_36263 =  i_22 & ~n_36202;
assign n_36264 =  x_1696 &  n_36202;
assign n_36265 = ~n_36263 & ~n_36264;
assign n_36266 =  x_1696 & ~n_36265;
assign n_36267 = ~x_1696 &  n_36265;
assign n_36268 = ~n_36266 & ~n_36267;
assign n_36269 =  i_21 & ~n_36202;
assign n_36270 =  x_1695 &  n_36202;
assign n_36271 = ~n_36269 & ~n_36270;
assign n_36272 =  x_1695 & ~n_36271;
assign n_36273 = ~x_1695 &  n_36271;
assign n_36274 = ~n_36272 & ~n_36273;
assign n_36275 =  i_20 & ~n_36202;
assign n_36276 =  x_1694 &  n_36202;
assign n_36277 = ~n_36275 & ~n_36276;
assign n_36278 =  x_1694 & ~n_36277;
assign n_36279 = ~x_1694 &  n_36277;
assign n_36280 = ~n_36278 & ~n_36279;
assign n_36281 =  i_19 & ~n_36202;
assign n_36282 =  x_1693 &  n_36202;
assign n_36283 = ~n_36281 & ~n_36282;
assign n_36284 =  x_1693 & ~n_36283;
assign n_36285 = ~x_1693 &  n_36283;
assign n_36286 = ~n_36284 & ~n_36285;
assign n_36287 =  i_18 & ~n_36202;
assign n_36288 =  x_1692 &  n_36202;
assign n_36289 = ~n_36287 & ~n_36288;
assign n_36290 =  x_1692 & ~n_36289;
assign n_36291 = ~x_1692 &  n_36289;
assign n_36292 = ~n_36290 & ~n_36291;
assign n_36293 =  i_17 & ~n_36202;
assign n_36294 =  x_1691 &  n_36202;
assign n_36295 = ~n_36293 & ~n_36294;
assign n_36296 =  x_1691 & ~n_36295;
assign n_36297 = ~x_1691 &  n_36295;
assign n_36298 = ~n_36296 & ~n_36297;
assign n_36299 =  i_16 & ~n_36202;
assign n_36300 =  x_1690 &  n_36202;
assign n_36301 = ~n_36299 & ~n_36300;
assign n_36302 =  x_1690 & ~n_36301;
assign n_36303 = ~x_1690 &  n_36301;
assign n_36304 = ~n_36302 & ~n_36303;
assign n_36305 =  i_15 & ~n_36202;
assign n_36306 =  x_1689 &  n_36202;
assign n_36307 = ~n_36305 & ~n_36306;
assign n_36308 =  x_1689 & ~n_36307;
assign n_36309 = ~x_1689 &  n_36307;
assign n_36310 = ~n_36308 & ~n_36309;
assign n_36311 =  i_14 & ~n_36202;
assign n_36312 =  x_1688 &  n_36202;
assign n_36313 = ~n_36311 & ~n_36312;
assign n_36314 =  x_1688 & ~n_36313;
assign n_36315 = ~x_1688 &  n_36313;
assign n_36316 = ~n_36314 & ~n_36315;
assign n_36317 =  i_13 & ~n_36202;
assign n_36318 =  x_1687 &  n_36202;
assign n_36319 = ~n_36317 & ~n_36318;
assign n_36320 =  x_1687 & ~n_36319;
assign n_36321 = ~x_1687 &  n_36319;
assign n_36322 = ~n_36320 & ~n_36321;
assign n_36323 =  i_12 & ~n_36202;
assign n_36324 =  x_1686 &  n_36202;
assign n_36325 = ~n_36323 & ~n_36324;
assign n_36326 =  x_1686 & ~n_36325;
assign n_36327 = ~x_1686 &  n_36325;
assign n_36328 = ~n_36326 & ~n_36327;
assign n_36329 =  i_11 & ~n_36202;
assign n_36330 =  x_1685 &  n_36202;
assign n_36331 = ~n_36329 & ~n_36330;
assign n_36332 =  x_1685 & ~n_36331;
assign n_36333 = ~x_1685 &  n_36331;
assign n_36334 = ~n_36332 & ~n_36333;
assign n_36335 =  i_10 & ~n_36202;
assign n_36336 =  x_1684 &  n_36202;
assign n_36337 = ~n_36335 & ~n_36336;
assign n_36338 =  x_1684 & ~n_36337;
assign n_36339 = ~x_1684 &  n_36337;
assign n_36340 = ~n_36338 & ~n_36339;
assign n_36341 =  i_9 & ~n_36202;
assign n_36342 =  x_1683 &  n_36202;
assign n_36343 = ~n_36341 & ~n_36342;
assign n_36344 =  x_1683 & ~n_36343;
assign n_36345 = ~x_1683 &  n_36343;
assign n_36346 = ~n_36344 & ~n_36345;
assign n_36347 =  i_8 & ~n_36202;
assign n_36348 =  x_1682 &  n_36202;
assign n_36349 = ~n_36347 & ~n_36348;
assign n_36350 =  x_1682 & ~n_36349;
assign n_36351 = ~x_1682 &  n_36349;
assign n_36352 = ~n_36350 & ~n_36351;
assign n_36353 =  i_7 & ~n_36202;
assign n_36354 =  x_1681 &  n_36202;
assign n_36355 = ~n_36353 & ~n_36354;
assign n_36356 =  x_1681 & ~n_36355;
assign n_36357 = ~x_1681 &  n_36355;
assign n_36358 = ~n_36356 & ~n_36357;
assign n_36359 =  i_6 & ~n_36202;
assign n_36360 =  x_1680 &  n_36202;
assign n_36361 = ~n_36359 & ~n_36360;
assign n_36362 =  x_1680 & ~n_36361;
assign n_36363 = ~x_1680 &  n_36361;
assign n_36364 = ~n_36362 & ~n_36363;
assign n_36365 =  i_5 & ~n_36202;
assign n_36366 =  x_1679 &  n_36202;
assign n_36367 = ~n_36365 & ~n_36366;
assign n_36368 =  x_1679 & ~n_36367;
assign n_36369 = ~x_1679 &  n_36367;
assign n_36370 = ~n_36368 & ~n_36369;
assign n_36371 =  i_4 & ~n_36202;
assign n_36372 =  x_1678 &  n_36202;
assign n_36373 = ~n_36371 & ~n_36372;
assign n_36374 =  x_1678 & ~n_36373;
assign n_36375 = ~x_1678 &  n_36373;
assign n_36376 = ~n_36374 & ~n_36375;
assign n_36377 =  i_3 & ~n_36202;
assign n_36378 =  x_1677 &  n_36202;
assign n_36379 = ~n_36377 & ~n_36378;
assign n_36380 =  x_1677 & ~n_36379;
assign n_36381 = ~x_1677 &  n_36379;
assign n_36382 = ~n_36380 & ~n_36381;
assign n_36383 =  i_2 & ~n_36202;
assign n_36384 =  x_1676 &  n_36202;
assign n_36385 = ~n_36383 & ~n_36384;
assign n_36386 =  x_1676 & ~n_36385;
assign n_36387 = ~x_1676 &  n_36385;
assign n_36388 = ~n_36386 & ~n_36387;
assign n_36389 =  i_1 & ~n_36202;
assign n_36390 =  x_1675 &  n_36202;
assign n_36391 = ~n_36389 & ~n_36390;
assign n_36392 =  x_1675 & ~n_36391;
assign n_36393 = ~x_1675 &  n_36391;
assign n_36394 = ~n_36392 & ~n_36393;
assign n_36395 =  x_1674 & ~n_27725;
assign n_36396 =  i_32 &  n_27725;
assign n_36397 = ~n_36395 & ~n_36396;
assign n_36398 =  x_1674 & ~n_36397;
assign n_36399 = ~x_1674 &  n_36397;
assign n_36400 = ~n_36398 & ~n_36399;
assign n_36401 =  x_1673 & ~n_27725;
assign n_36402 =  i_31 &  n_27725;
assign n_36403 = ~n_36401 & ~n_36402;
assign n_36404 =  x_1673 & ~n_36403;
assign n_36405 = ~x_1673 &  n_36403;
assign n_36406 = ~n_36404 & ~n_36405;
assign n_36407 =  x_1672 & ~n_27725;
assign n_36408 =  i_30 &  n_27725;
assign n_36409 = ~n_36407 & ~n_36408;
assign n_36410 =  x_1672 & ~n_36409;
assign n_36411 = ~x_1672 &  n_36409;
assign n_36412 = ~n_36410 & ~n_36411;
assign n_36413 =  x_1671 & ~n_27725;
assign n_36414 =  i_29 &  n_27725;
assign n_36415 = ~n_36413 & ~n_36414;
assign n_36416 =  x_1671 & ~n_36415;
assign n_36417 = ~x_1671 &  n_36415;
assign n_36418 = ~n_36416 & ~n_36417;
assign n_36419 =  x_1670 & ~n_27725;
assign n_36420 =  i_28 &  n_27725;
assign n_36421 = ~n_36419 & ~n_36420;
assign n_36422 =  x_1670 & ~n_36421;
assign n_36423 = ~x_1670 &  n_36421;
assign n_36424 = ~n_36422 & ~n_36423;
assign n_36425 =  x_1669 & ~n_27725;
assign n_36426 =  i_27 &  n_27725;
assign n_36427 = ~n_36425 & ~n_36426;
assign n_36428 =  x_1669 & ~n_36427;
assign n_36429 = ~x_1669 &  n_36427;
assign n_36430 = ~n_36428 & ~n_36429;
assign n_36431 =  x_1668 & ~n_27725;
assign n_36432 =  i_26 &  n_27725;
assign n_36433 = ~n_36431 & ~n_36432;
assign n_36434 =  x_1668 & ~n_36433;
assign n_36435 = ~x_1668 &  n_36433;
assign n_36436 = ~n_36434 & ~n_36435;
assign n_36437 =  x_1667 & ~n_27725;
assign n_36438 =  i_25 &  n_27725;
assign n_36439 = ~n_36437 & ~n_36438;
assign n_36440 =  x_1667 & ~n_36439;
assign n_36441 = ~x_1667 &  n_36439;
assign n_36442 = ~n_36440 & ~n_36441;
assign n_36443 =  x_1666 & ~n_27725;
assign n_36444 =  i_24 &  n_27725;
assign n_36445 = ~n_36443 & ~n_36444;
assign n_36446 =  x_1666 & ~n_36445;
assign n_36447 = ~x_1666 &  n_36445;
assign n_36448 = ~n_36446 & ~n_36447;
assign n_36449 =  x_1665 & ~n_27725;
assign n_36450 =  i_23 &  n_27725;
assign n_36451 = ~n_36449 & ~n_36450;
assign n_36452 =  x_1665 & ~n_36451;
assign n_36453 = ~x_1665 &  n_36451;
assign n_36454 = ~n_36452 & ~n_36453;
assign n_36455 =  x_1664 & ~n_27725;
assign n_36456 =  i_22 &  n_27725;
assign n_36457 = ~n_36455 & ~n_36456;
assign n_36458 =  x_1664 & ~n_36457;
assign n_36459 = ~x_1664 &  n_36457;
assign n_36460 = ~n_36458 & ~n_36459;
assign n_36461 =  x_1663 & ~n_27725;
assign n_36462 =  i_21 &  n_27725;
assign n_36463 = ~n_36461 & ~n_36462;
assign n_36464 =  x_1663 & ~n_36463;
assign n_36465 = ~x_1663 &  n_36463;
assign n_36466 = ~n_36464 & ~n_36465;
assign n_36467 =  x_1662 & ~n_27725;
assign n_36468 =  i_20 &  n_27725;
assign n_36469 = ~n_36467 & ~n_36468;
assign n_36470 =  x_1662 & ~n_36469;
assign n_36471 = ~x_1662 &  n_36469;
assign n_36472 = ~n_36470 & ~n_36471;
assign n_36473 =  x_1661 & ~n_27725;
assign n_36474 =  i_19 &  n_27725;
assign n_36475 = ~n_36473 & ~n_36474;
assign n_36476 =  x_1661 & ~n_36475;
assign n_36477 = ~x_1661 &  n_36475;
assign n_36478 = ~n_36476 & ~n_36477;
assign n_36479 =  x_1660 & ~n_27725;
assign n_36480 =  i_18 &  n_27725;
assign n_36481 = ~n_36479 & ~n_36480;
assign n_36482 =  x_1660 & ~n_36481;
assign n_36483 = ~x_1660 &  n_36481;
assign n_36484 = ~n_36482 & ~n_36483;
assign n_36485 =  x_1659 & ~n_27725;
assign n_36486 =  i_17 &  n_27725;
assign n_36487 = ~n_36485 & ~n_36486;
assign n_36488 =  x_1659 & ~n_36487;
assign n_36489 = ~x_1659 &  n_36487;
assign n_36490 = ~n_36488 & ~n_36489;
assign n_36491 =  x_1658 & ~n_27725;
assign n_36492 =  i_16 &  n_27725;
assign n_36493 = ~n_36491 & ~n_36492;
assign n_36494 =  x_1658 & ~n_36493;
assign n_36495 = ~x_1658 &  n_36493;
assign n_36496 = ~n_36494 & ~n_36495;
assign n_36497 =  x_1657 & ~n_27725;
assign n_36498 =  i_15 &  n_27725;
assign n_36499 = ~n_36497 & ~n_36498;
assign n_36500 =  x_1657 & ~n_36499;
assign n_36501 = ~x_1657 &  n_36499;
assign n_36502 = ~n_36500 & ~n_36501;
assign n_36503 =  x_1656 & ~n_27725;
assign n_36504 =  i_14 &  n_27725;
assign n_36505 = ~n_36503 & ~n_36504;
assign n_36506 =  x_1656 & ~n_36505;
assign n_36507 = ~x_1656 &  n_36505;
assign n_36508 = ~n_36506 & ~n_36507;
assign n_36509 =  x_1655 & ~n_27725;
assign n_36510 =  i_13 &  n_27725;
assign n_36511 = ~n_36509 & ~n_36510;
assign n_36512 =  x_1655 & ~n_36511;
assign n_36513 = ~x_1655 &  n_36511;
assign n_36514 = ~n_36512 & ~n_36513;
assign n_36515 =  x_1654 & ~n_27725;
assign n_36516 =  i_12 &  n_27725;
assign n_36517 = ~n_36515 & ~n_36516;
assign n_36518 =  x_1654 & ~n_36517;
assign n_36519 = ~x_1654 &  n_36517;
assign n_36520 = ~n_36518 & ~n_36519;
assign n_36521 =  x_1653 & ~n_27725;
assign n_36522 =  i_11 &  n_27725;
assign n_36523 = ~n_36521 & ~n_36522;
assign n_36524 =  x_1653 & ~n_36523;
assign n_36525 = ~x_1653 &  n_36523;
assign n_36526 = ~n_36524 & ~n_36525;
assign n_36527 =  x_1652 & ~n_27725;
assign n_36528 =  i_10 &  n_27725;
assign n_36529 = ~n_36527 & ~n_36528;
assign n_36530 =  x_1652 & ~n_36529;
assign n_36531 = ~x_1652 &  n_36529;
assign n_36532 = ~n_36530 & ~n_36531;
assign n_36533 =  x_1651 & ~n_27725;
assign n_36534 =  i_9 &  n_27725;
assign n_36535 = ~n_36533 & ~n_36534;
assign n_36536 =  x_1651 & ~n_36535;
assign n_36537 = ~x_1651 &  n_36535;
assign n_36538 = ~n_36536 & ~n_36537;
assign n_36539 =  x_1650 & ~n_27725;
assign n_36540 =  i_8 &  n_27725;
assign n_36541 = ~n_36539 & ~n_36540;
assign n_36542 =  x_1650 & ~n_36541;
assign n_36543 = ~x_1650 &  n_36541;
assign n_36544 = ~n_36542 & ~n_36543;
assign n_36545 =  x_1649 & ~n_27725;
assign n_36546 =  i_7 &  n_27725;
assign n_36547 = ~n_36545 & ~n_36546;
assign n_36548 =  x_1649 & ~n_36547;
assign n_36549 = ~x_1649 &  n_36547;
assign n_36550 = ~n_36548 & ~n_36549;
assign n_36551 =  x_1648 & ~n_27725;
assign n_36552 =  i_6 &  n_27725;
assign n_36553 = ~n_36551 & ~n_36552;
assign n_36554 =  x_1648 & ~n_36553;
assign n_36555 = ~x_1648 &  n_36553;
assign n_36556 = ~n_36554 & ~n_36555;
assign n_36557 =  x_1647 & ~n_27725;
assign n_36558 =  i_5 &  n_27725;
assign n_36559 = ~n_36557 & ~n_36558;
assign n_36560 =  x_1647 & ~n_36559;
assign n_36561 = ~x_1647 &  n_36559;
assign n_36562 = ~n_36560 & ~n_36561;
assign n_36563 =  x_1646 & ~n_27725;
assign n_36564 =  i_4 &  n_27725;
assign n_36565 = ~n_36563 & ~n_36564;
assign n_36566 =  x_1646 & ~n_36565;
assign n_36567 = ~x_1646 &  n_36565;
assign n_36568 = ~n_36566 & ~n_36567;
assign n_36569 =  x_1645 & ~n_27725;
assign n_36570 =  i_3 &  n_27725;
assign n_36571 = ~n_36569 & ~n_36570;
assign n_36572 =  x_1645 & ~n_36571;
assign n_36573 = ~x_1645 &  n_36571;
assign n_36574 = ~n_36572 & ~n_36573;
assign n_36575 =  x_1644 & ~n_27725;
assign n_36576 =  i_2 &  n_27725;
assign n_36577 = ~n_36575 & ~n_36576;
assign n_36578 =  x_1644 & ~n_36577;
assign n_36579 = ~x_1644 &  n_36577;
assign n_36580 = ~n_36578 & ~n_36579;
assign n_36581 =  x_1643 & ~n_27725;
assign n_36582 =  i_1 &  n_27725;
assign n_36583 = ~n_36581 & ~n_36582;
assign n_36584 =  x_1643 & ~n_36583;
assign n_36585 = ~x_1643 &  n_36583;
assign n_36586 = ~n_36584 & ~n_36585;
assign n_36587 =  i_32 & ~n_12324;
assign n_36588 =  x_3064 &  n_12324;
assign n_36589 = ~n_36587 & ~n_36588;
assign n_36590 = ~n_12331 & ~n_36589;
assign n_36591 =  x_2906 &  n_12331;
assign n_36592 = ~n_36590 & ~n_36591;
assign n_36593 = ~n_12332 & ~n_36592;
assign n_36594 =  x_2842 &  n_12332;
assign n_36595 = ~n_36593 & ~n_36594;
assign n_36596 =  n_28074 & ~n_36595;
assign n_36597 =  x_1642 & ~n_28074;
assign n_36598 = ~n_36596 & ~n_36597;
assign n_36599 =  x_1642 & ~n_36598;
assign n_36600 = ~x_1642 &  n_36598;
assign n_36601 = ~n_36599 & ~n_36600;
assign n_36602 =  i_31 & ~n_12324;
assign n_36603 =  x_3063 &  n_12324;
assign n_36604 = ~n_36602 & ~n_36603;
assign n_36605 = ~n_12331 & ~n_36604;
assign n_36606 =  x_2905 &  n_12331;
assign n_36607 = ~n_36605 & ~n_36606;
assign n_36608 = ~n_12332 & ~n_36607;
assign n_36609 =  x_2841 &  n_12332;
assign n_36610 = ~n_36608 & ~n_36609;
assign n_36611 =  n_28074 & ~n_36610;
assign n_36612 =  x_1641 & ~n_28074;
assign n_36613 = ~n_36611 & ~n_36612;
assign n_36614 =  x_1641 & ~n_36613;
assign n_36615 = ~x_1641 &  n_36613;
assign n_36616 = ~n_36614 & ~n_36615;
assign n_36617 =  i_30 & ~n_12324;
assign n_36618 =  x_3062 &  n_12324;
assign n_36619 = ~n_36617 & ~n_36618;
assign n_36620 = ~n_12331 & ~n_36619;
assign n_36621 =  x_2904 &  n_12331;
assign n_36622 = ~n_36620 & ~n_36621;
assign n_36623 = ~n_12332 & ~n_36622;
assign n_36624 =  x_2840 &  n_12332;
assign n_36625 = ~n_36623 & ~n_36624;
assign n_36626 =  n_28074 & ~n_36625;
assign n_36627 =  x_1640 & ~n_28074;
assign n_36628 = ~n_36626 & ~n_36627;
assign n_36629 =  x_1640 & ~n_36628;
assign n_36630 = ~x_1640 &  n_36628;
assign n_36631 = ~n_36629 & ~n_36630;
assign n_36632 =  i_29 & ~n_12324;
assign n_36633 =  x_3061 &  n_12324;
assign n_36634 = ~n_36632 & ~n_36633;
assign n_36635 = ~n_12331 & ~n_36634;
assign n_36636 =  x_2903 &  n_12331;
assign n_36637 = ~n_36635 & ~n_36636;
assign n_36638 = ~n_12332 & ~n_36637;
assign n_36639 =  x_2839 &  n_12332;
assign n_36640 = ~n_36638 & ~n_36639;
assign n_36641 =  n_28074 & ~n_36640;
assign n_36642 =  x_1639 & ~n_28074;
assign n_36643 = ~n_36641 & ~n_36642;
assign n_36644 =  x_1639 & ~n_36643;
assign n_36645 = ~x_1639 &  n_36643;
assign n_36646 = ~n_36644 & ~n_36645;
assign n_36647 =  i_28 & ~n_12324;
assign n_36648 =  x_3060 &  n_12324;
assign n_36649 = ~n_36647 & ~n_36648;
assign n_36650 = ~n_12331 & ~n_36649;
assign n_36651 =  x_2902 &  n_12331;
assign n_36652 = ~n_36650 & ~n_36651;
assign n_36653 = ~n_12332 & ~n_36652;
assign n_36654 =  x_2838 &  n_12332;
assign n_36655 = ~n_36653 & ~n_36654;
assign n_36656 =  n_28074 & ~n_36655;
assign n_36657 =  x_1638 & ~n_28074;
assign n_36658 = ~n_36656 & ~n_36657;
assign n_36659 =  x_1638 & ~n_36658;
assign n_36660 = ~x_1638 &  n_36658;
assign n_36661 = ~n_36659 & ~n_36660;
assign n_36662 =  i_27 & ~n_12324;
assign n_36663 =  x_3059 &  n_12324;
assign n_36664 = ~n_36662 & ~n_36663;
assign n_36665 = ~n_12331 & ~n_36664;
assign n_36666 =  x_2901 &  n_12331;
assign n_36667 = ~n_36665 & ~n_36666;
assign n_36668 = ~n_12332 & ~n_36667;
assign n_36669 =  x_2837 &  n_12332;
assign n_36670 = ~n_36668 & ~n_36669;
assign n_36671 =  n_28074 & ~n_36670;
assign n_36672 =  x_1637 & ~n_28074;
assign n_36673 = ~n_36671 & ~n_36672;
assign n_36674 =  x_1637 & ~n_36673;
assign n_36675 = ~x_1637 &  n_36673;
assign n_36676 = ~n_36674 & ~n_36675;
assign n_36677 =  i_26 & ~n_12324;
assign n_36678 =  x_3058 &  n_12324;
assign n_36679 = ~n_36677 & ~n_36678;
assign n_36680 = ~n_12331 & ~n_36679;
assign n_36681 =  x_2900 &  n_12331;
assign n_36682 = ~n_36680 & ~n_36681;
assign n_36683 = ~n_12332 & ~n_36682;
assign n_36684 =  x_2836 &  n_12332;
assign n_36685 = ~n_36683 & ~n_36684;
assign n_36686 =  n_28074 & ~n_36685;
assign n_36687 =  x_1636 & ~n_28074;
assign n_36688 = ~n_36686 & ~n_36687;
assign n_36689 =  x_1636 & ~n_36688;
assign n_36690 = ~x_1636 &  n_36688;
assign n_36691 = ~n_36689 & ~n_36690;
assign n_36692 =  i_25 & ~n_12324;
assign n_36693 =  x_3057 &  n_12324;
assign n_36694 = ~n_36692 & ~n_36693;
assign n_36695 = ~n_12331 & ~n_36694;
assign n_36696 =  x_2899 &  n_12331;
assign n_36697 = ~n_36695 & ~n_36696;
assign n_36698 = ~n_12332 & ~n_36697;
assign n_36699 =  x_2835 &  n_12332;
assign n_36700 = ~n_36698 & ~n_36699;
assign n_36701 =  n_28074 & ~n_36700;
assign n_36702 =  x_1635 & ~n_28074;
assign n_36703 = ~n_36701 & ~n_36702;
assign n_36704 =  x_1635 & ~n_36703;
assign n_36705 = ~x_1635 &  n_36703;
assign n_36706 = ~n_36704 & ~n_36705;
assign n_36707 =  i_24 & ~n_12324;
assign n_36708 =  x_3056 &  n_12324;
assign n_36709 = ~n_36707 & ~n_36708;
assign n_36710 = ~n_12331 & ~n_36709;
assign n_36711 =  x_2898 &  n_12331;
assign n_36712 = ~n_36710 & ~n_36711;
assign n_36713 = ~n_12332 & ~n_36712;
assign n_36714 =  x_2834 &  n_12332;
assign n_36715 = ~n_36713 & ~n_36714;
assign n_36716 =  n_28074 & ~n_36715;
assign n_36717 =  x_1634 & ~n_28074;
assign n_36718 = ~n_36716 & ~n_36717;
assign n_36719 =  x_1634 & ~n_36718;
assign n_36720 = ~x_1634 &  n_36718;
assign n_36721 = ~n_36719 & ~n_36720;
assign n_36722 =  i_23 & ~n_12324;
assign n_36723 =  x_3055 &  n_12324;
assign n_36724 = ~n_36722 & ~n_36723;
assign n_36725 = ~n_12331 & ~n_36724;
assign n_36726 =  x_2897 &  n_12331;
assign n_36727 = ~n_36725 & ~n_36726;
assign n_36728 = ~n_12332 & ~n_36727;
assign n_36729 =  x_2833 &  n_12332;
assign n_36730 = ~n_36728 & ~n_36729;
assign n_36731 =  n_28074 & ~n_36730;
assign n_36732 =  x_1633 & ~n_28074;
assign n_36733 = ~n_36731 & ~n_36732;
assign n_36734 =  x_1633 & ~n_36733;
assign n_36735 = ~x_1633 &  n_36733;
assign n_36736 = ~n_36734 & ~n_36735;
assign n_36737 =  i_22 & ~n_12324;
assign n_36738 =  x_3054 &  n_12324;
assign n_36739 = ~n_36737 & ~n_36738;
assign n_36740 = ~n_12331 & ~n_36739;
assign n_36741 =  x_2896 &  n_12331;
assign n_36742 = ~n_36740 & ~n_36741;
assign n_36743 = ~n_12332 & ~n_36742;
assign n_36744 =  x_2832 &  n_12332;
assign n_36745 = ~n_36743 & ~n_36744;
assign n_36746 =  n_28074 & ~n_36745;
assign n_36747 =  x_1632 & ~n_28074;
assign n_36748 = ~n_36746 & ~n_36747;
assign n_36749 =  x_1632 & ~n_36748;
assign n_36750 = ~x_1632 &  n_36748;
assign n_36751 = ~n_36749 & ~n_36750;
assign n_36752 =  i_21 & ~n_12324;
assign n_36753 =  x_3053 &  n_12324;
assign n_36754 = ~n_36752 & ~n_36753;
assign n_36755 = ~n_12331 & ~n_36754;
assign n_36756 =  x_2895 &  n_12331;
assign n_36757 = ~n_36755 & ~n_36756;
assign n_36758 = ~n_12332 & ~n_36757;
assign n_36759 =  x_2831 &  n_12332;
assign n_36760 = ~n_36758 & ~n_36759;
assign n_36761 =  n_28074 & ~n_36760;
assign n_36762 =  x_1631 & ~n_28074;
assign n_36763 = ~n_36761 & ~n_36762;
assign n_36764 =  x_1631 & ~n_36763;
assign n_36765 = ~x_1631 &  n_36763;
assign n_36766 = ~n_36764 & ~n_36765;
assign n_36767 =  i_20 & ~n_12324;
assign n_36768 =  x_3052 &  n_12324;
assign n_36769 = ~n_36767 & ~n_36768;
assign n_36770 = ~n_12331 & ~n_36769;
assign n_36771 =  x_2894 &  n_12331;
assign n_36772 = ~n_36770 & ~n_36771;
assign n_36773 = ~n_12332 & ~n_36772;
assign n_36774 =  x_2830 &  n_12332;
assign n_36775 = ~n_36773 & ~n_36774;
assign n_36776 =  n_28074 & ~n_36775;
assign n_36777 =  x_1630 & ~n_28074;
assign n_36778 = ~n_36776 & ~n_36777;
assign n_36779 =  x_1630 & ~n_36778;
assign n_36780 = ~x_1630 &  n_36778;
assign n_36781 = ~n_36779 & ~n_36780;
assign n_36782 =  i_19 & ~n_12324;
assign n_36783 =  x_3051 &  n_12324;
assign n_36784 = ~n_36782 & ~n_36783;
assign n_36785 = ~n_12331 & ~n_36784;
assign n_36786 =  x_2893 &  n_12331;
assign n_36787 = ~n_36785 & ~n_36786;
assign n_36788 = ~n_12332 & ~n_36787;
assign n_36789 =  x_2829 &  n_12332;
assign n_36790 = ~n_36788 & ~n_36789;
assign n_36791 =  n_28074 & ~n_36790;
assign n_36792 =  x_1629 & ~n_28074;
assign n_36793 = ~n_36791 & ~n_36792;
assign n_36794 =  x_1629 & ~n_36793;
assign n_36795 = ~x_1629 &  n_36793;
assign n_36796 = ~n_36794 & ~n_36795;
assign n_36797 =  i_18 & ~n_12324;
assign n_36798 =  x_3050 &  n_12324;
assign n_36799 = ~n_36797 & ~n_36798;
assign n_36800 = ~n_12331 & ~n_36799;
assign n_36801 =  x_2892 &  n_12331;
assign n_36802 = ~n_36800 & ~n_36801;
assign n_36803 = ~n_12332 & ~n_36802;
assign n_36804 =  x_2828 &  n_12332;
assign n_36805 = ~n_36803 & ~n_36804;
assign n_36806 =  n_28074 & ~n_36805;
assign n_36807 =  x_1628 & ~n_28074;
assign n_36808 = ~n_36806 & ~n_36807;
assign n_36809 =  x_1628 & ~n_36808;
assign n_36810 = ~x_1628 &  n_36808;
assign n_36811 = ~n_36809 & ~n_36810;
assign n_36812 =  i_17 & ~n_12324;
assign n_36813 =  x_3049 &  n_12324;
assign n_36814 = ~n_36812 & ~n_36813;
assign n_36815 = ~n_12331 & ~n_36814;
assign n_36816 =  x_2891 &  n_12331;
assign n_36817 = ~n_36815 & ~n_36816;
assign n_36818 = ~n_12332 & ~n_36817;
assign n_36819 =  x_2827 &  n_12332;
assign n_36820 = ~n_36818 & ~n_36819;
assign n_36821 =  n_28074 & ~n_36820;
assign n_36822 =  x_1627 & ~n_28074;
assign n_36823 = ~n_36821 & ~n_36822;
assign n_36824 =  x_1627 & ~n_36823;
assign n_36825 = ~x_1627 &  n_36823;
assign n_36826 = ~n_36824 & ~n_36825;
assign n_36827 =  i_16 & ~n_12324;
assign n_36828 =  x_3048 &  n_12324;
assign n_36829 = ~n_36827 & ~n_36828;
assign n_36830 = ~n_12331 & ~n_36829;
assign n_36831 =  x_2890 &  n_12331;
assign n_36832 = ~n_36830 & ~n_36831;
assign n_36833 = ~n_12332 & ~n_36832;
assign n_36834 =  x_2826 &  n_12332;
assign n_36835 = ~n_36833 & ~n_36834;
assign n_36836 =  n_28074 & ~n_36835;
assign n_36837 =  x_1626 & ~n_28074;
assign n_36838 = ~n_36836 & ~n_36837;
assign n_36839 =  x_1626 & ~n_36838;
assign n_36840 = ~x_1626 &  n_36838;
assign n_36841 = ~n_36839 & ~n_36840;
assign n_36842 =  i_15 & ~n_12324;
assign n_36843 =  x_3047 &  n_12324;
assign n_36844 = ~n_36842 & ~n_36843;
assign n_36845 = ~n_12331 & ~n_36844;
assign n_36846 =  x_2889 &  n_12331;
assign n_36847 = ~n_36845 & ~n_36846;
assign n_36848 = ~n_12332 & ~n_36847;
assign n_36849 =  x_2825 &  n_12332;
assign n_36850 = ~n_36848 & ~n_36849;
assign n_36851 =  n_28074 & ~n_36850;
assign n_36852 =  x_1625 & ~n_28074;
assign n_36853 = ~n_36851 & ~n_36852;
assign n_36854 =  x_1625 & ~n_36853;
assign n_36855 = ~x_1625 &  n_36853;
assign n_36856 = ~n_36854 & ~n_36855;
assign n_36857 =  i_14 & ~n_12324;
assign n_36858 =  x_3046 &  n_12324;
assign n_36859 = ~n_36857 & ~n_36858;
assign n_36860 = ~n_12331 & ~n_36859;
assign n_36861 =  x_2888 &  n_12331;
assign n_36862 = ~n_36860 & ~n_36861;
assign n_36863 = ~n_12332 & ~n_36862;
assign n_36864 =  x_2824 &  n_12332;
assign n_36865 = ~n_36863 & ~n_36864;
assign n_36866 =  n_28074 & ~n_36865;
assign n_36867 =  x_1624 & ~n_28074;
assign n_36868 = ~n_36866 & ~n_36867;
assign n_36869 =  x_1624 & ~n_36868;
assign n_36870 = ~x_1624 &  n_36868;
assign n_36871 = ~n_36869 & ~n_36870;
assign n_36872 =  i_13 & ~n_12324;
assign n_36873 =  x_3045 &  n_12324;
assign n_36874 = ~n_36872 & ~n_36873;
assign n_36875 = ~n_12331 & ~n_36874;
assign n_36876 =  x_2887 &  n_12331;
assign n_36877 = ~n_36875 & ~n_36876;
assign n_36878 = ~n_12332 & ~n_36877;
assign n_36879 =  x_2823 &  n_12332;
assign n_36880 = ~n_36878 & ~n_36879;
assign n_36881 =  n_28074 & ~n_36880;
assign n_36882 =  x_1623 & ~n_28074;
assign n_36883 = ~n_36881 & ~n_36882;
assign n_36884 =  x_1623 & ~n_36883;
assign n_36885 = ~x_1623 &  n_36883;
assign n_36886 = ~n_36884 & ~n_36885;
assign n_36887 =  i_12 & ~n_12324;
assign n_36888 =  x_3044 &  n_12324;
assign n_36889 = ~n_36887 & ~n_36888;
assign n_36890 = ~n_12331 & ~n_36889;
assign n_36891 =  x_2886 &  n_12331;
assign n_36892 = ~n_36890 & ~n_36891;
assign n_36893 = ~n_12332 & ~n_36892;
assign n_36894 =  x_2822 &  n_12332;
assign n_36895 = ~n_36893 & ~n_36894;
assign n_36896 =  n_28074 & ~n_36895;
assign n_36897 =  x_1622 & ~n_28074;
assign n_36898 = ~n_36896 & ~n_36897;
assign n_36899 =  x_1622 & ~n_36898;
assign n_36900 = ~x_1622 &  n_36898;
assign n_36901 = ~n_36899 & ~n_36900;
assign n_36902 =  i_11 & ~n_12324;
assign n_36903 =  x_3043 &  n_12324;
assign n_36904 = ~n_36902 & ~n_36903;
assign n_36905 = ~n_12331 & ~n_36904;
assign n_36906 =  x_2885 &  n_12331;
assign n_36907 = ~n_36905 & ~n_36906;
assign n_36908 = ~n_12332 & ~n_36907;
assign n_36909 =  x_2821 &  n_12332;
assign n_36910 = ~n_36908 & ~n_36909;
assign n_36911 =  n_28074 & ~n_36910;
assign n_36912 =  x_1621 & ~n_28074;
assign n_36913 = ~n_36911 & ~n_36912;
assign n_36914 =  x_1621 & ~n_36913;
assign n_36915 = ~x_1621 &  n_36913;
assign n_36916 = ~n_36914 & ~n_36915;
assign n_36917 =  i_10 & ~n_12324;
assign n_36918 =  x_3042 &  n_12324;
assign n_36919 = ~n_36917 & ~n_36918;
assign n_36920 = ~n_12331 & ~n_36919;
assign n_36921 =  x_2884 &  n_12331;
assign n_36922 = ~n_36920 & ~n_36921;
assign n_36923 = ~n_12332 & ~n_36922;
assign n_36924 =  x_2820 &  n_12332;
assign n_36925 = ~n_36923 & ~n_36924;
assign n_36926 =  n_28074 & ~n_36925;
assign n_36927 =  x_1620 & ~n_28074;
assign n_36928 = ~n_36926 & ~n_36927;
assign n_36929 =  x_1620 & ~n_36928;
assign n_36930 = ~x_1620 &  n_36928;
assign n_36931 = ~n_36929 & ~n_36930;
assign n_36932 =  i_9 & ~n_12324;
assign n_36933 =  x_3041 &  n_12324;
assign n_36934 = ~n_36932 & ~n_36933;
assign n_36935 = ~n_12331 & ~n_36934;
assign n_36936 =  x_2883 &  n_12331;
assign n_36937 = ~n_36935 & ~n_36936;
assign n_36938 = ~n_12332 & ~n_36937;
assign n_36939 =  x_2819 &  n_12332;
assign n_36940 = ~n_36938 & ~n_36939;
assign n_36941 =  n_28074 & ~n_36940;
assign n_36942 =  x_1619 & ~n_28074;
assign n_36943 = ~n_36941 & ~n_36942;
assign n_36944 =  x_1619 & ~n_36943;
assign n_36945 = ~x_1619 &  n_36943;
assign n_36946 = ~n_36944 & ~n_36945;
assign n_36947 =  i_8 & ~n_12324;
assign n_36948 =  x_3040 &  n_12324;
assign n_36949 = ~n_36947 & ~n_36948;
assign n_36950 = ~n_12331 & ~n_36949;
assign n_36951 =  x_2882 &  n_12331;
assign n_36952 = ~n_36950 & ~n_36951;
assign n_36953 = ~n_12332 & ~n_36952;
assign n_36954 =  x_2818 &  n_12332;
assign n_36955 = ~n_36953 & ~n_36954;
assign n_36956 =  n_28074 & ~n_36955;
assign n_36957 =  x_1618 & ~n_28074;
assign n_36958 = ~n_36956 & ~n_36957;
assign n_36959 =  x_1618 & ~n_36958;
assign n_36960 = ~x_1618 &  n_36958;
assign n_36961 = ~n_36959 & ~n_36960;
assign n_36962 =  i_7 & ~n_12324;
assign n_36963 =  x_3039 &  n_12324;
assign n_36964 = ~n_36962 & ~n_36963;
assign n_36965 = ~n_12331 & ~n_36964;
assign n_36966 =  x_2881 &  n_12331;
assign n_36967 = ~n_36965 & ~n_36966;
assign n_36968 = ~n_12332 & ~n_36967;
assign n_36969 =  x_2817 &  n_12332;
assign n_36970 = ~n_36968 & ~n_36969;
assign n_36971 =  n_28074 & ~n_36970;
assign n_36972 =  x_1617 & ~n_28074;
assign n_36973 = ~n_36971 & ~n_36972;
assign n_36974 =  x_1617 & ~n_36973;
assign n_36975 = ~x_1617 &  n_36973;
assign n_36976 = ~n_36974 & ~n_36975;
assign n_36977 =  i_6 & ~n_12324;
assign n_36978 =  x_3038 &  n_12324;
assign n_36979 = ~n_36977 & ~n_36978;
assign n_36980 = ~n_12331 & ~n_36979;
assign n_36981 =  x_2880 &  n_12331;
assign n_36982 = ~n_36980 & ~n_36981;
assign n_36983 = ~n_12332 & ~n_36982;
assign n_36984 =  x_2816 &  n_12332;
assign n_36985 = ~n_36983 & ~n_36984;
assign n_36986 =  n_28074 & ~n_36985;
assign n_36987 =  x_1616 & ~n_28074;
assign n_36988 = ~n_36986 & ~n_36987;
assign n_36989 =  x_1616 & ~n_36988;
assign n_36990 = ~x_1616 &  n_36988;
assign n_36991 = ~n_36989 & ~n_36990;
assign n_36992 =  i_5 & ~n_12324;
assign n_36993 =  x_3037 &  n_12324;
assign n_36994 = ~n_36992 & ~n_36993;
assign n_36995 = ~n_12331 & ~n_36994;
assign n_36996 =  x_2879 &  n_12331;
assign n_36997 = ~n_36995 & ~n_36996;
assign n_36998 = ~n_12332 & ~n_36997;
assign n_36999 =  x_2815 &  n_12332;
assign n_37000 = ~n_36998 & ~n_36999;
assign n_37001 =  n_28074 & ~n_37000;
assign n_37002 =  x_1615 & ~n_28074;
assign n_37003 = ~n_37001 & ~n_37002;
assign n_37004 =  x_1615 & ~n_37003;
assign n_37005 = ~x_1615 &  n_37003;
assign n_37006 = ~n_37004 & ~n_37005;
assign n_37007 =  i_4 & ~n_12324;
assign n_37008 =  x_3036 &  n_12324;
assign n_37009 = ~n_37007 & ~n_37008;
assign n_37010 = ~n_12331 & ~n_37009;
assign n_37011 =  x_2878 &  n_12331;
assign n_37012 = ~n_37010 & ~n_37011;
assign n_37013 = ~n_12332 & ~n_37012;
assign n_37014 =  x_2814 &  n_12332;
assign n_37015 = ~n_37013 & ~n_37014;
assign n_37016 =  n_28074 & ~n_37015;
assign n_37017 =  x_1614 & ~n_28074;
assign n_37018 = ~n_37016 & ~n_37017;
assign n_37019 =  x_1614 & ~n_37018;
assign n_37020 = ~x_1614 &  n_37018;
assign n_37021 = ~n_37019 & ~n_37020;
assign n_37022 =  i_3 & ~n_12324;
assign n_37023 =  x_3035 &  n_12324;
assign n_37024 = ~n_37022 & ~n_37023;
assign n_37025 = ~n_12331 & ~n_37024;
assign n_37026 =  x_2877 &  n_12331;
assign n_37027 = ~n_37025 & ~n_37026;
assign n_37028 = ~n_12332 & ~n_37027;
assign n_37029 =  x_2813 &  n_12332;
assign n_37030 = ~n_37028 & ~n_37029;
assign n_37031 =  n_28074 & ~n_37030;
assign n_37032 =  x_1613 & ~n_28074;
assign n_37033 = ~n_37031 & ~n_37032;
assign n_37034 =  x_1613 & ~n_37033;
assign n_37035 = ~x_1613 &  n_37033;
assign n_37036 = ~n_37034 & ~n_37035;
assign n_37037 =  i_2 & ~n_12324;
assign n_37038 =  x_3034 &  n_12324;
assign n_37039 = ~n_37037 & ~n_37038;
assign n_37040 = ~n_12331 & ~n_37039;
assign n_37041 =  x_2876 &  n_12331;
assign n_37042 = ~n_37040 & ~n_37041;
assign n_37043 = ~n_12332 & ~n_37042;
assign n_37044 =  x_2812 &  n_12332;
assign n_37045 = ~n_37043 & ~n_37044;
assign n_37046 =  n_28074 & ~n_37045;
assign n_37047 =  x_1612 & ~n_28074;
assign n_37048 = ~n_37046 & ~n_37047;
assign n_37049 =  x_1612 & ~n_37048;
assign n_37050 = ~x_1612 &  n_37048;
assign n_37051 = ~n_37049 & ~n_37050;
assign n_37052 =  i_1 & ~n_12324;
assign n_37053 =  x_3033 &  n_12324;
assign n_37054 = ~n_37052 & ~n_37053;
assign n_37055 = ~n_12331 & ~n_37054;
assign n_37056 =  x_2875 &  n_12331;
assign n_37057 = ~n_37055 & ~n_37056;
assign n_37058 = ~n_12332 & ~n_37057;
assign n_37059 =  x_2811 &  n_12332;
assign n_37060 = ~n_37058 & ~n_37059;
assign n_37061 =  n_28074 & ~n_37060;
assign n_37062 =  x_1611 & ~n_28074;
assign n_37063 = ~n_37061 & ~n_37062;
assign n_37064 =  x_1611 & ~n_37063;
assign n_37065 = ~x_1611 &  n_37063;
assign n_37066 = ~n_37064 & ~n_37065;
assign n_37067 =  x_1610 & ~n_16882;
assign n_37068 =  x_3096 &  n_16882;
assign n_37069 = ~n_37067 & ~n_37068;
assign n_37070 =  x_1610 & ~n_37069;
assign n_37071 = ~x_1610 &  n_37069;
assign n_37072 = ~n_37070 & ~n_37071;
assign n_37073 =  x_1609 & ~n_16882;
assign n_37074 =  x_3095 &  n_16882;
assign n_37075 = ~n_37073 & ~n_37074;
assign n_37076 =  x_1609 & ~n_37075;
assign n_37077 = ~x_1609 &  n_37075;
assign n_37078 = ~n_37076 & ~n_37077;
assign n_37079 =  x_1608 & ~n_16882;
assign n_37080 =  x_3094 &  n_16882;
assign n_37081 = ~n_37079 & ~n_37080;
assign n_37082 =  x_1608 & ~n_37081;
assign n_37083 = ~x_1608 &  n_37081;
assign n_37084 = ~n_37082 & ~n_37083;
assign n_37085 =  x_1607 & ~n_16882;
assign n_37086 =  x_3093 &  n_16882;
assign n_37087 = ~n_37085 & ~n_37086;
assign n_37088 =  x_1607 & ~n_37087;
assign n_37089 = ~x_1607 &  n_37087;
assign n_37090 = ~n_37088 & ~n_37089;
assign n_37091 =  x_1606 & ~n_16882;
assign n_37092 =  x_3092 &  n_16882;
assign n_37093 = ~n_37091 & ~n_37092;
assign n_37094 =  x_1606 & ~n_37093;
assign n_37095 = ~x_1606 &  n_37093;
assign n_37096 = ~n_37094 & ~n_37095;
assign n_37097 =  x_1605 & ~n_16882;
assign n_37098 =  x_3091 &  n_16882;
assign n_37099 = ~n_37097 & ~n_37098;
assign n_37100 =  x_1605 & ~n_37099;
assign n_37101 = ~x_1605 &  n_37099;
assign n_37102 = ~n_37100 & ~n_37101;
assign n_37103 =  x_1604 & ~n_16882;
assign n_37104 =  x_3090 &  n_16882;
assign n_37105 = ~n_37103 & ~n_37104;
assign n_37106 =  x_1604 & ~n_37105;
assign n_37107 = ~x_1604 &  n_37105;
assign n_37108 = ~n_37106 & ~n_37107;
assign n_37109 =  x_1603 & ~n_16882;
assign n_37110 =  x_3089 &  n_16882;
assign n_37111 = ~n_37109 & ~n_37110;
assign n_37112 =  x_1603 & ~n_37111;
assign n_37113 = ~x_1603 &  n_37111;
assign n_37114 = ~n_37112 & ~n_37113;
assign n_37115 =  x_1602 & ~n_16882;
assign n_37116 =  x_3088 &  n_16882;
assign n_37117 = ~n_37115 & ~n_37116;
assign n_37118 =  x_1602 & ~n_37117;
assign n_37119 = ~x_1602 &  n_37117;
assign n_37120 = ~n_37118 & ~n_37119;
assign n_37121 =  x_1601 & ~n_16882;
assign n_37122 =  x_3087 &  n_16882;
assign n_37123 = ~n_37121 & ~n_37122;
assign n_37124 =  x_1601 & ~n_37123;
assign n_37125 = ~x_1601 &  n_37123;
assign n_37126 = ~n_37124 & ~n_37125;
assign n_37127 =  x_1600 & ~n_16882;
assign n_37128 =  x_3086 &  n_16882;
assign n_37129 = ~n_37127 & ~n_37128;
assign n_37130 =  x_1600 & ~n_37129;
assign n_37131 = ~x_1600 &  n_37129;
assign n_37132 = ~n_37130 & ~n_37131;
assign n_37133 =  x_1599 & ~n_16882;
assign n_37134 =  x_3085 &  n_16882;
assign n_37135 = ~n_37133 & ~n_37134;
assign n_37136 =  x_1599 & ~n_37135;
assign n_37137 = ~x_1599 &  n_37135;
assign n_37138 = ~n_37136 & ~n_37137;
assign n_37139 =  x_1598 & ~n_16882;
assign n_37140 =  x_3084 &  n_16882;
assign n_37141 = ~n_37139 & ~n_37140;
assign n_37142 =  x_1598 & ~n_37141;
assign n_37143 = ~x_1598 &  n_37141;
assign n_37144 = ~n_37142 & ~n_37143;
assign n_37145 =  x_1597 & ~n_16882;
assign n_37146 =  x_3083 &  n_16882;
assign n_37147 = ~n_37145 & ~n_37146;
assign n_37148 =  x_1597 & ~n_37147;
assign n_37149 = ~x_1597 &  n_37147;
assign n_37150 = ~n_37148 & ~n_37149;
assign n_37151 =  x_1596 & ~n_16882;
assign n_37152 =  x_3082 &  n_16882;
assign n_37153 = ~n_37151 & ~n_37152;
assign n_37154 =  x_1596 & ~n_37153;
assign n_37155 = ~x_1596 &  n_37153;
assign n_37156 = ~n_37154 & ~n_37155;
assign n_37157 =  x_1595 & ~n_16882;
assign n_37158 =  x_3081 &  n_16882;
assign n_37159 = ~n_37157 & ~n_37158;
assign n_37160 =  x_1595 & ~n_37159;
assign n_37161 = ~x_1595 &  n_37159;
assign n_37162 = ~n_37160 & ~n_37161;
assign n_37163 =  x_1594 & ~n_16882;
assign n_37164 =  x_3080 &  n_16882;
assign n_37165 = ~n_37163 & ~n_37164;
assign n_37166 =  x_1594 & ~n_37165;
assign n_37167 = ~x_1594 &  n_37165;
assign n_37168 = ~n_37166 & ~n_37167;
assign n_37169 =  x_1593 & ~n_16882;
assign n_37170 =  x_3079 &  n_16882;
assign n_37171 = ~n_37169 & ~n_37170;
assign n_37172 =  x_1593 & ~n_37171;
assign n_37173 = ~x_1593 &  n_37171;
assign n_37174 = ~n_37172 & ~n_37173;
assign n_37175 =  x_1592 & ~n_16882;
assign n_37176 =  x_3078 &  n_16882;
assign n_37177 = ~n_37175 & ~n_37176;
assign n_37178 =  x_1592 & ~n_37177;
assign n_37179 = ~x_1592 &  n_37177;
assign n_37180 = ~n_37178 & ~n_37179;
assign n_37181 =  x_1591 & ~n_16882;
assign n_37182 =  x_3077 &  n_16882;
assign n_37183 = ~n_37181 & ~n_37182;
assign n_37184 =  x_1591 & ~n_37183;
assign n_37185 = ~x_1591 &  n_37183;
assign n_37186 = ~n_37184 & ~n_37185;
assign n_37187 =  x_1590 & ~n_16882;
assign n_37188 =  x_3076 &  n_16882;
assign n_37189 = ~n_37187 & ~n_37188;
assign n_37190 =  x_1590 & ~n_37189;
assign n_37191 = ~x_1590 &  n_37189;
assign n_37192 = ~n_37190 & ~n_37191;
assign n_37193 =  x_1589 & ~n_16882;
assign n_37194 =  x_3075 &  n_16882;
assign n_37195 = ~n_37193 & ~n_37194;
assign n_37196 =  x_1589 & ~n_37195;
assign n_37197 = ~x_1589 &  n_37195;
assign n_37198 = ~n_37196 & ~n_37197;
assign n_37199 =  x_1588 & ~n_16882;
assign n_37200 =  x_3074 &  n_16882;
assign n_37201 = ~n_37199 & ~n_37200;
assign n_37202 =  x_1588 & ~n_37201;
assign n_37203 = ~x_1588 &  n_37201;
assign n_37204 = ~n_37202 & ~n_37203;
assign n_37205 =  x_1587 & ~n_16882;
assign n_37206 =  x_3073 &  n_16882;
assign n_37207 = ~n_37205 & ~n_37206;
assign n_37208 =  x_1587 & ~n_37207;
assign n_37209 = ~x_1587 &  n_37207;
assign n_37210 = ~n_37208 & ~n_37209;
assign n_37211 =  x_1586 & ~n_16882;
assign n_37212 =  x_3072 &  n_16882;
assign n_37213 = ~n_37211 & ~n_37212;
assign n_37214 =  x_1586 & ~n_37213;
assign n_37215 = ~x_1586 &  n_37213;
assign n_37216 = ~n_37214 & ~n_37215;
assign n_37217 =  x_1585 & ~n_16882;
assign n_37218 =  x_3071 &  n_16882;
assign n_37219 = ~n_37217 & ~n_37218;
assign n_37220 =  x_1585 & ~n_37219;
assign n_37221 = ~x_1585 &  n_37219;
assign n_37222 = ~n_37220 & ~n_37221;
assign n_37223 =  x_1584 & ~n_16882;
assign n_37224 =  x_3070 &  n_16882;
assign n_37225 = ~n_37223 & ~n_37224;
assign n_37226 =  x_1584 & ~n_37225;
assign n_37227 = ~x_1584 &  n_37225;
assign n_37228 = ~n_37226 & ~n_37227;
assign n_37229 =  x_1583 & ~n_16882;
assign n_37230 =  x_3069 &  n_16882;
assign n_37231 = ~n_37229 & ~n_37230;
assign n_37232 =  x_1583 & ~n_37231;
assign n_37233 = ~x_1583 &  n_37231;
assign n_37234 = ~n_37232 & ~n_37233;
assign n_37235 =  x_1582 & ~n_16882;
assign n_37236 =  x_3068 &  n_16882;
assign n_37237 = ~n_37235 & ~n_37236;
assign n_37238 =  x_1582 & ~n_37237;
assign n_37239 = ~x_1582 &  n_37237;
assign n_37240 = ~n_37238 & ~n_37239;
assign n_37241 =  x_1581 & ~n_16882;
assign n_37242 =  x_3067 &  n_16882;
assign n_37243 = ~n_37241 & ~n_37242;
assign n_37244 =  x_1581 & ~n_37243;
assign n_37245 = ~x_1581 &  n_37243;
assign n_37246 = ~n_37244 & ~n_37245;
assign n_37247 =  x_1580 & ~n_16882;
assign n_37248 =  x_3066 &  n_16882;
assign n_37249 = ~n_37247 & ~n_37248;
assign n_37250 =  x_1580 & ~n_37249;
assign n_37251 = ~x_1580 &  n_37249;
assign n_37252 = ~n_37250 & ~n_37251;
assign n_37253 =  x_1579 & ~n_16882;
assign n_37254 =  x_3065 &  n_16882;
assign n_37255 = ~n_37253 & ~n_37254;
assign n_37256 =  x_1579 & ~n_37255;
assign n_37257 = ~x_1579 &  n_37255;
assign n_37258 = ~n_37256 & ~n_37257;
assign n_37259 = ~n_24051 & ~n_28364;
assign n_37260 =  x_1578 &  n_37259;
assign n_37261 =  x_1770 &  n_24051;
assign n_37262 =  x_3000 &  n_28364;
assign n_37263 = ~n_37261 & ~n_37262;
assign n_37264 = ~n_37260 &  n_37263;
assign n_37265 =  x_1578 & ~n_37264;
assign n_37266 = ~x_1578 &  n_37264;
assign n_37267 = ~n_37265 & ~n_37266;
assign n_37268 =  x_1577 &  n_37259;
assign n_37269 =  x_1769 &  n_24051;
assign n_37270 =  x_2999 &  n_28364;
assign n_37271 = ~n_37269 & ~n_37270;
assign n_37272 = ~n_37268 &  n_37271;
assign n_37273 =  x_1577 & ~n_37272;
assign n_37274 = ~x_1577 &  n_37272;
assign n_37275 = ~n_37273 & ~n_37274;
assign n_37276 =  x_1576 &  n_37259;
assign n_37277 =  x_1768 &  n_24051;
assign n_37278 =  x_2998 &  n_28364;
assign n_37279 = ~n_37277 & ~n_37278;
assign n_37280 = ~n_37276 &  n_37279;
assign n_37281 =  x_1576 & ~n_37280;
assign n_37282 = ~x_1576 &  n_37280;
assign n_37283 = ~n_37281 & ~n_37282;
assign n_37284 =  x_1575 &  n_37259;
assign n_37285 =  x_1767 &  n_24051;
assign n_37286 =  x_2997 &  n_28364;
assign n_37287 = ~n_37285 & ~n_37286;
assign n_37288 = ~n_37284 &  n_37287;
assign n_37289 =  x_1575 & ~n_37288;
assign n_37290 = ~x_1575 &  n_37288;
assign n_37291 = ~n_37289 & ~n_37290;
assign n_37292 =  x_1574 &  n_37259;
assign n_37293 =  x_1766 &  n_24051;
assign n_37294 =  x_2996 &  n_28364;
assign n_37295 = ~n_37293 & ~n_37294;
assign n_37296 = ~n_37292 &  n_37295;
assign n_37297 =  x_1574 & ~n_37296;
assign n_37298 = ~x_1574 &  n_37296;
assign n_37299 = ~n_37297 & ~n_37298;
assign n_37300 =  x_1573 &  n_37259;
assign n_37301 =  x_1765 &  n_24051;
assign n_37302 =  x_2995 &  n_28364;
assign n_37303 = ~n_37301 & ~n_37302;
assign n_37304 = ~n_37300 &  n_37303;
assign n_37305 =  x_1573 & ~n_37304;
assign n_37306 = ~x_1573 &  n_37304;
assign n_37307 = ~n_37305 & ~n_37306;
assign n_37308 =  x_1572 &  n_37259;
assign n_37309 =  x_1764 &  n_24051;
assign n_37310 =  x_2994 &  n_28364;
assign n_37311 = ~n_37309 & ~n_37310;
assign n_37312 = ~n_37308 &  n_37311;
assign n_37313 =  x_1572 & ~n_37312;
assign n_37314 = ~x_1572 &  n_37312;
assign n_37315 = ~n_37313 & ~n_37314;
assign n_37316 =  x_1571 &  n_37259;
assign n_37317 =  x_1763 &  n_24051;
assign n_37318 =  x_2993 &  n_28364;
assign n_37319 = ~n_37317 & ~n_37318;
assign n_37320 = ~n_37316 &  n_37319;
assign n_37321 =  x_1571 & ~n_37320;
assign n_37322 = ~x_1571 &  n_37320;
assign n_37323 = ~n_37321 & ~n_37322;
assign n_37324 =  x_1570 &  n_37259;
assign n_37325 =  x_1762 &  n_24051;
assign n_37326 =  x_2992 &  n_28364;
assign n_37327 = ~n_37325 & ~n_37326;
assign n_37328 = ~n_37324 &  n_37327;
assign n_37329 =  x_1570 & ~n_37328;
assign n_37330 = ~x_1570 &  n_37328;
assign n_37331 = ~n_37329 & ~n_37330;
assign n_37332 =  x_1569 &  n_37259;
assign n_37333 =  x_1761 &  n_24051;
assign n_37334 =  x_2991 &  n_28364;
assign n_37335 = ~n_37333 & ~n_37334;
assign n_37336 = ~n_37332 &  n_37335;
assign n_37337 =  x_1569 & ~n_37336;
assign n_37338 = ~x_1569 &  n_37336;
assign n_37339 = ~n_37337 & ~n_37338;
assign n_37340 =  x_1568 &  n_37259;
assign n_37341 =  x_1760 &  n_24051;
assign n_37342 =  x_2990 &  n_28364;
assign n_37343 = ~n_37341 & ~n_37342;
assign n_37344 = ~n_37340 &  n_37343;
assign n_37345 =  x_1568 & ~n_37344;
assign n_37346 = ~x_1568 &  n_37344;
assign n_37347 = ~n_37345 & ~n_37346;
assign n_37348 =  x_1567 &  n_37259;
assign n_37349 =  x_1759 &  n_24051;
assign n_37350 =  x_2989 &  n_28364;
assign n_37351 = ~n_37349 & ~n_37350;
assign n_37352 = ~n_37348 &  n_37351;
assign n_37353 =  x_1567 & ~n_37352;
assign n_37354 = ~x_1567 &  n_37352;
assign n_37355 = ~n_37353 & ~n_37354;
assign n_37356 =  x_1566 &  n_37259;
assign n_37357 =  x_1758 &  n_24051;
assign n_37358 =  x_2988 &  n_28364;
assign n_37359 = ~n_37357 & ~n_37358;
assign n_37360 = ~n_37356 &  n_37359;
assign n_37361 =  x_1566 & ~n_37360;
assign n_37362 = ~x_1566 &  n_37360;
assign n_37363 = ~n_37361 & ~n_37362;
assign n_37364 =  x_1565 &  n_37259;
assign n_37365 =  x_1757 &  n_24051;
assign n_37366 =  x_2987 &  n_28364;
assign n_37367 = ~n_37365 & ~n_37366;
assign n_37368 = ~n_37364 &  n_37367;
assign n_37369 =  x_1565 & ~n_37368;
assign n_37370 = ~x_1565 &  n_37368;
assign n_37371 = ~n_37369 & ~n_37370;
assign n_37372 =  x_1564 &  n_37259;
assign n_37373 =  x_1756 &  n_24051;
assign n_37374 =  x_2986 &  n_28364;
assign n_37375 = ~n_37373 & ~n_37374;
assign n_37376 = ~n_37372 &  n_37375;
assign n_37377 =  x_1564 & ~n_37376;
assign n_37378 = ~x_1564 &  n_37376;
assign n_37379 = ~n_37377 & ~n_37378;
assign n_37380 =  x_1563 &  n_37259;
assign n_37381 =  x_1755 &  n_24051;
assign n_37382 =  x_2985 &  n_28364;
assign n_37383 = ~n_37381 & ~n_37382;
assign n_37384 = ~n_37380 &  n_37383;
assign n_37385 =  x_1563 & ~n_37384;
assign n_37386 = ~x_1563 &  n_37384;
assign n_37387 = ~n_37385 & ~n_37386;
assign n_37388 =  x_1562 &  n_37259;
assign n_37389 =  x_1754 &  n_24051;
assign n_37390 =  x_2984 &  n_28364;
assign n_37391 = ~n_37389 & ~n_37390;
assign n_37392 = ~n_37388 &  n_37391;
assign n_37393 =  x_1562 & ~n_37392;
assign n_37394 = ~x_1562 &  n_37392;
assign n_37395 = ~n_37393 & ~n_37394;
assign n_37396 =  x_1561 &  n_37259;
assign n_37397 =  x_1753 &  n_24051;
assign n_37398 =  x_2983 &  n_28364;
assign n_37399 = ~n_37397 & ~n_37398;
assign n_37400 = ~n_37396 &  n_37399;
assign n_37401 =  x_1561 & ~n_37400;
assign n_37402 = ~x_1561 &  n_37400;
assign n_37403 = ~n_37401 & ~n_37402;
assign n_37404 =  x_1560 &  n_37259;
assign n_37405 =  x_1752 &  n_24051;
assign n_37406 =  x_2982 &  n_28364;
assign n_37407 = ~n_37405 & ~n_37406;
assign n_37408 = ~n_37404 &  n_37407;
assign n_37409 =  x_1560 & ~n_37408;
assign n_37410 = ~x_1560 &  n_37408;
assign n_37411 = ~n_37409 & ~n_37410;
assign n_37412 =  x_1559 &  n_37259;
assign n_37413 =  x_1751 &  n_24051;
assign n_37414 =  x_2981 &  n_28364;
assign n_37415 = ~n_37413 & ~n_37414;
assign n_37416 = ~n_37412 &  n_37415;
assign n_37417 =  x_1559 & ~n_37416;
assign n_37418 = ~x_1559 &  n_37416;
assign n_37419 = ~n_37417 & ~n_37418;
assign n_37420 =  x_1558 &  n_37259;
assign n_37421 =  x_1750 &  n_24051;
assign n_37422 =  x_2980 &  n_28364;
assign n_37423 = ~n_37421 & ~n_37422;
assign n_37424 = ~n_37420 &  n_37423;
assign n_37425 =  x_1558 & ~n_37424;
assign n_37426 = ~x_1558 &  n_37424;
assign n_37427 = ~n_37425 & ~n_37426;
assign n_37428 =  x_1557 &  n_37259;
assign n_37429 =  x_1749 &  n_24051;
assign n_37430 =  x_2979 &  n_28364;
assign n_37431 = ~n_37429 & ~n_37430;
assign n_37432 = ~n_37428 &  n_37431;
assign n_37433 =  x_1557 & ~n_37432;
assign n_37434 = ~x_1557 &  n_37432;
assign n_37435 = ~n_37433 & ~n_37434;
assign n_37436 =  x_1556 &  n_37259;
assign n_37437 =  x_1748 &  n_24051;
assign n_37438 =  x_2978 &  n_28364;
assign n_37439 = ~n_37437 & ~n_37438;
assign n_37440 = ~n_37436 &  n_37439;
assign n_37441 =  x_1556 & ~n_37440;
assign n_37442 = ~x_1556 &  n_37440;
assign n_37443 = ~n_37441 & ~n_37442;
assign n_37444 =  x_1555 &  n_37259;
assign n_37445 =  x_1747 &  n_24051;
assign n_37446 =  x_2977 &  n_28364;
assign n_37447 = ~n_37445 & ~n_37446;
assign n_37448 = ~n_37444 &  n_37447;
assign n_37449 =  x_1555 & ~n_37448;
assign n_37450 = ~x_1555 &  n_37448;
assign n_37451 = ~n_37449 & ~n_37450;
assign n_37452 =  x_1554 &  n_37259;
assign n_37453 =  x_1746 &  n_24051;
assign n_37454 =  x_2976 &  n_28364;
assign n_37455 = ~n_37453 & ~n_37454;
assign n_37456 = ~n_37452 &  n_37455;
assign n_37457 =  x_1554 & ~n_37456;
assign n_37458 = ~x_1554 &  n_37456;
assign n_37459 = ~n_37457 & ~n_37458;
assign n_37460 =  x_1553 &  n_37259;
assign n_37461 =  x_1745 &  n_24051;
assign n_37462 =  x_2975 &  n_28364;
assign n_37463 = ~n_37461 & ~n_37462;
assign n_37464 = ~n_37460 &  n_37463;
assign n_37465 =  x_1553 & ~n_37464;
assign n_37466 = ~x_1553 &  n_37464;
assign n_37467 = ~n_37465 & ~n_37466;
assign n_37468 =  x_1552 &  n_37259;
assign n_37469 =  x_1744 &  n_24051;
assign n_37470 =  x_2974 &  n_28364;
assign n_37471 = ~n_37469 & ~n_37470;
assign n_37472 = ~n_37468 &  n_37471;
assign n_37473 =  x_1552 & ~n_37472;
assign n_37474 = ~x_1552 &  n_37472;
assign n_37475 = ~n_37473 & ~n_37474;
assign n_37476 =  x_1551 &  n_37259;
assign n_37477 =  x_1743 &  n_24051;
assign n_37478 =  x_2973 &  n_28364;
assign n_37479 = ~n_37477 & ~n_37478;
assign n_37480 = ~n_37476 &  n_37479;
assign n_37481 =  x_1551 & ~n_37480;
assign n_37482 = ~x_1551 &  n_37480;
assign n_37483 = ~n_37481 & ~n_37482;
assign n_37484 =  x_1550 &  n_37259;
assign n_37485 =  x_1742 &  n_24051;
assign n_37486 =  x_2972 &  n_28364;
assign n_37487 = ~n_37485 & ~n_37486;
assign n_37488 = ~n_37484 &  n_37487;
assign n_37489 =  x_1550 & ~n_37488;
assign n_37490 = ~x_1550 &  n_37488;
assign n_37491 = ~n_37489 & ~n_37490;
assign n_37492 =  x_1549 &  n_37259;
assign n_37493 =  x_1741 &  n_24051;
assign n_37494 =  x_2971 &  n_28364;
assign n_37495 = ~n_37493 & ~n_37494;
assign n_37496 = ~n_37492 &  n_37495;
assign n_37497 =  x_1549 & ~n_37496;
assign n_37498 = ~x_1549 &  n_37496;
assign n_37499 = ~n_37497 & ~n_37498;
assign n_37500 =  x_1548 &  n_37259;
assign n_37501 =  x_1740 &  n_24051;
assign n_37502 =  x_2970 &  n_28364;
assign n_37503 = ~n_37501 & ~n_37502;
assign n_37504 = ~n_37500 &  n_37503;
assign n_37505 =  x_1548 & ~n_37504;
assign n_37506 = ~x_1548 &  n_37504;
assign n_37507 = ~n_37505 & ~n_37506;
assign n_37508 =  x_1739 &  n_24051;
assign n_37509 =  x_1547 &  n_37259;
assign n_37510 = ~n_37508 & ~n_37509;
assign n_37511 =  x_1547 & ~n_37510;
assign n_37512 = ~x_1547 &  n_37510;
assign n_37513 = ~n_37511 & ~n_37512;
assign n_37514 =  x_1546 & ~n_26173;
assign n_37515 =  i_32 &  n_26173;
assign n_37516 = ~n_37514 & ~n_37515;
assign n_37517 =  x_1546 & ~n_37516;
assign n_37518 = ~x_1546 &  n_37516;
assign n_37519 = ~n_37517 & ~n_37518;
assign n_37520 =  x_1545 & ~n_26173;
assign n_37521 =  i_31 &  n_26173;
assign n_37522 = ~n_37520 & ~n_37521;
assign n_37523 =  x_1545 & ~n_37522;
assign n_37524 = ~x_1545 &  n_37522;
assign n_37525 = ~n_37523 & ~n_37524;
assign n_37526 =  x_1544 & ~n_26173;
assign n_37527 =  i_30 &  n_26173;
assign n_37528 = ~n_37526 & ~n_37527;
assign n_37529 =  x_1544 & ~n_37528;
assign n_37530 = ~x_1544 &  n_37528;
assign n_37531 = ~n_37529 & ~n_37530;
assign n_37532 =  x_1543 & ~n_26173;
assign n_37533 =  i_29 &  n_26173;
assign n_37534 = ~n_37532 & ~n_37533;
assign n_37535 =  x_1543 & ~n_37534;
assign n_37536 = ~x_1543 &  n_37534;
assign n_37537 = ~n_37535 & ~n_37536;
assign n_37538 =  x_1542 & ~n_26173;
assign n_37539 =  i_28 &  n_26173;
assign n_37540 = ~n_37538 & ~n_37539;
assign n_37541 =  x_1542 & ~n_37540;
assign n_37542 = ~x_1542 &  n_37540;
assign n_37543 = ~n_37541 & ~n_37542;
assign n_37544 =  x_1541 & ~n_26173;
assign n_37545 =  i_27 &  n_26173;
assign n_37546 = ~n_37544 & ~n_37545;
assign n_37547 =  x_1541 & ~n_37546;
assign n_37548 = ~x_1541 &  n_37546;
assign n_37549 = ~n_37547 & ~n_37548;
assign n_37550 =  x_1540 & ~n_26173;
assign n_37551 =  i_26 &  n_26173;
assign n_37552 = ~n_37550 & ~n_37551;
assign n_37553 =  x_1540 & ~n_37552;
assign n_37554 = ~x_1540 &  n_37552;
assign n_37555 = ~n_37553 & ~n_37554;
assign n_37556 =  x_1539 & ~n_26173;
assign n_37557 =  i_25 &  n_26173;
assign n_37558 = ~n_37556 & ~n_37557;
assign n_37559 =  x_1539 & ~n_37558;
assign n_37560 = ~x_1539 &  n_37558;
assign n_37561 = ~n_37559 & ~n_37560;
assign n_37562 =  x_1538 & ~n_26173;
assign n_37563 =  i_24 &  n_26173;
assign n_37564 = ~n_37562 & ~n_37563;
assign n_37565 =  x_1538 & ~n_37564;
assign n_37566 = ~x_1538 &  n_37564;
assign n_37567 = ~n_37565 & ~n_37566;
assign n_37568 =  x_1537 & ~n_26173;
assign n_37569 =  i_23 &  n_26173;
assign n_37570 = ~n_37568 & ~n_37569;
assign n_37571 =  x_1537 & ~n_37570;
assign n_37572 = ~x_1537 &  n_37570;
assign n_37573 = ~n_37571 & ~n_37572;
assign n_37574 =  x_1536 & ~n_26173;
assign n_37575 =  i_22 &  n_26173;
assign n_37576 = ~n_37574 & ~n_37575;
assign n_37577 =  x_1536 & ~n_37576;
assign n_37578 = ~x_1536 &  n_37576;
assign n_37579 = ~n_37577 & ~n_37578;
assign n_37580 =  x_1535 & ~n_26173;
assign n_37581 =  i_21 &  n_26173;
assign n_37582 = ~n_37580 & ~n_37581;
assign n_37583 =  x_1535 & ~n_37582;
assign n_37584 = ~x_1535 &  n_37582;
assign n_37585 = ~n_37583 & ~n_37584;
assign n_37586 =  x_1534 & ~n_26173;
assign n_37587 =  i_20 &  n_26173;
assign n_37588 = ~n_37586 & ~n_37587;
assign n_37589 =  x_1534 & ~n_37588;
assign n_37590 = ~x_1534 &  n_37588;
assign n_37591 = ~n_37589 & ~n_37590;
assign n_37592 =  x_1533 & ~n_26173;
assign n_37593 =  i_19 &  n_26173;
assign n_37594 = ~n_37592 & ~n_37593;
assign n_37595 =  x_1533 & ~n_37594;
assign n_37596 = ~x_1533 &  n_37594;
assign n_37597 = ~n_37595 & ~n_37596;
assign n_37598 =  x_1532 & ~n_26173;
assign n_37599 =  i_18 &  n_26173;
assign n_37600 = ~n_37598 & ~n_37599;
assign n_37601 =  x_1532 & ~n_37600;
assign n_37602 = ~x_1532 &  n_37600;
assign n_37603 = ~n_37601 & ~n_37602;
assign n_37604 =  x_1531 & ~n_26173;
assign n_37605 =  i_17 &  n_26173;
assign n_37606 = ~n_37604 & ~n_37605;
assign n_37607 =  x_1531 & ~n_37606;
assign n_37608 = ~x_1531 &  n_37606;
assign n_37609 = ~n_37607 & ~n_37608;
assign n_37610 =  x_1530 & ~n_26173;
assign n_37611 =  i_16 &  n_26173;
assign n_37612 = ~n_37610 & ~n_37611;
assign n_37613 =  x_1530 & ~n_37612;
assign n_37614 = ~x_1530 &  n_37612;
assign n_37615 = ~n_37613 & ~n_37614;
assign n_37616 =  x_1529 & ~n_26173;
assign n_37617 =  i_15 &  n_26173;
assign n_37618 = ~n_37616 & ~n_37617;
assign n_37619 =  x_1529 & ~n_37618;
assign n_37620 = ~x_1529 &  n_37618;
assign n_37621 = ~n_37619 & ~n_37620;
assign n_37622 =  x_1528 & ~n_26173;
assign n_37623 =  i_14 &  n_26173;
assign n_37624 = ~n_37622 & ~n_37623;
assign n_37625 =  x_1528 & ~n_37624;
assign n_37626 = ~x_1528 &  n_37624;
assign n_37627 = ~n_37625 & ~n_37626;
assign n_37628 =  x_1527 & ~n_26173;
assign n_37629 =  i_13 &  n_26173;
assign n_37630 = ~n_37628 & ~n_37629;
assign n_37631 =  x_1527 & ~n_37630;
assign n_37632 = ~x_1527 &  n_37630;
assign n_37633 = ~n_37631 & ~n_37632;
assign n_37634 =  x_1526 & ~n_26173;
assign n_37635 =  i_12 &  n_26173;
assign n_37636 = ~n_37634 & ~n_37635;
assign n_37637 =  x_1526 & ~n_37636;
assign n_37638 = ~x_1526 &  n_37636;
assign n_37639 = ~n_37637 & ~n_37638;
assign n_37640 =  x_1525 & ~n_26173;
assign n_37641 =  i_11 &  n_26173;
assign n_37642 = ~n_37640 & ~n_37641;
assign n_37643 =  x_1525 & ~n_37642;
assign n_37644 = ~x_1525 &  n_37642;
assign n_37645 = ~n_37643 & ~n_37644;
assign n_37646 =  x_1524 & ~n_26173;
assign n_37647 =  i_10 &  n_26173;
assign n_37648 = ~n_37646 & ~n_37647;
assign n_37649 =  x_1524 & ~n_37648;
assign n_37650 = ~x_1524 &  n_37648;
assign n_37651 = ~n_37649 & ~n_37650;
assign n_37652 =  x_1523 & ~n_26173;
assign n_37653 =  i_9 &  n_26173;
assign n_37654 = ~n_37652 & ~n_37653;
assign n_37655 =  x_1523 & ~n_37654;
assign n_37656 = ~x_1523 &  n_37654;
assign n_37657 = ~n_37655 & ~n_37656;
assign n_37658 =  x_1522 & ~n_26173;
assign n_37659 =  i_8 &  n_26173;
assign n_37660 = ~n_37658 & ~n_37659;
assign n_37661 =  x_1522 & ~n_37660;
assign n_37662 = ~x_1522 &  n_37660;
assign n_37663 = ~n_37661 & ~n_37662;
assign n_37664 =  x_1521 & ~n_26173;
assign n_37665 =  i_7 &  n_26173;
assign n_37666 = ~n_37664 & ~n_37665;
assign n_37667 =  x_1521 & ~n_37666;
assign n_37668 = ~x_1521 &  n_37666;
assign n_37669 = ~n_37667 & ~n_37668;
assign n_37670 =  x_1520 & ~n_26173;
assign n_37671 =  i_6 &  n_26173;
assign n_37672 = ~n_37670 & ~n_37671;
assign n_37673 =  x_1520 & ~n_37672;
assign n_37674 = ~x_1520 &  n_37672;
assign n_37675 = ~n_37673 & ~n_37674;
assign n_37676 =  x_1519 & ~n_26173;
assign n_37677 =  i_5 &  n_26173;
assign n_37678 = ~n_37676 & ~n_37677;
assign n_37679 =  x_1519 & ~n_37678;
assign n_37680 = ~x_1519 &  n_37678;
assign n_37681 = ~n_37679 & ~n_37680;
assign n_37682 =  x_1518 & ~n_26173;
assign n_37683 =  i_4 &  n_26173;
assign n_37684 = ~n_37682 & ~n_37683;
assign n_37685 =  x_1518 & ~n_37684;
assign n_37686 = ~x_1518 &  n_37684;
assign n_37687 = ~n_37685 & ~n_37686;
assign n_37688 =  x_1517 & ~n_26173;
assign n_37689 =  i_3 &  n_26173;
assign n_37690 = ~n_37688 & ~n_37689;
assign n_37691 =  x_1517 & ~n_37690;
assign n_37692 = ~x_1517 &  n_37690;
assign n_37693 = ~n_37691 & ~n_37692;
assign n_37694 =  x_1516 & ~n_26173;
assign n_37695 =  i_2 &  n_26173;
assign n_37696 = ~n_37694 & ~n_37695;
assign n_37697 =  x_1516 & ~n_37696;
assign n_37698 = ~x_1516 &  n_37696;
assign n_37699 = ~n_37697 & ~n_37698;
assign n_37700 =  x_1515 & ~n_26173;
assign n_37701 =  i_1 &  n_26173;
assign n_37702 = ~n_37700 & ~n_37701;
assign n_37703 =  x_1515 & ~n_37702;
assign n_37704 = ~x_1515 &  n_37702;
assign n_37705 = ~n_37703 & ~n_37704;
assign n_37706 =  n_26156 & ~n_36595;
assign n_37707 =  x_1514 & ~n_26156;
assign n_37708 = ~n_37706 & ~n_37707;
assign n_37709 =  x_1514 & ~n_37708;
assign n_37710 = ~x_1514 &  n_37708;
assign n_37711 = ~n_37709 & ~n_37710;
assign n_37712 =  n_26156 & ~n_36610;
assign n_37713 =  x_1513 & ~n_26156;
assign n_37714 = ~n_37712 & ~n_37713;
assign n_37715 =  x_1513 & ~n_37714;
assign n_37716 = ~x_1513 &  n_37714;
assign n_37717 = ~n_37715 & ~n_37716;
assign n_37718 =  n_26156 & ~n_36625;
assign n_37719 =  x_1512 & ~n_26156;
assign n_37720 = ~n_37718 & ~n_37719;
assign n_37721 =  x_1512 & ~n_37720;
assign n_37722 = ~x_1512 &  n_37720;
assign n_37723 = ~n_37721 & ~n_37722;
assign n_37724 =  n_26156 & ~n_36640;
assign n_37725 =  x_1511 & ~n_26156;
assign n_37726 = ~n_37724 & ~n_37725;
assign n_37727 =  x_1511 & ~n_37726;
assign n_37728 = ~x_1511 &  n_37726;
assign n_37729 = ~n_37727 & ~n_37728;
assign n_37730 =  n_26156 & ~n_36655;
assign n_37731 =  x_1510 & ~n_26156;
assign n_37732 = ~n_37730 & ~n_37731;
assign n_37733 =  x_1510 & ~n_37732;
assign n_37734 = ~x_1510 &  n_37732;
assign n_37735 = ~n_37733 & ~n_37734;
assign n_37736 =  n_26156 & ~n_36670;
assign n_37737 =  x_1509 & ~n_26156;
assign n_37738 = ~n_37736 & ~n_37737;
assign n_37739 =  x_1509 & ~n_37738;
assign n_37740 = ~x_1509 &  n_37738;
assign n_37741 = ~n_37739 & ~n_37740;
assign n_37742 =  n_26156 & ~n_36685;
assign n_37743 =  x_1508 & ~n_26156;
assign n_37744 = ~n_37742 & ~n_37743;
assign n_37745 =  x_1508 & ~n_37744;
assign n_37746 = ~x_1508 &  n_37744;
assign n_37747 = ~n_37745 & ~n_37746;
assign n_37748 =  n_26156 & ~n_36700;
assign n_37749 =  x_1507 & ~n_26156;
assign n_37750 = ~n_37748 & ~n_37749;
assign n_37751 =  x_1507 & ~n_37750;
assign n_37752 = ~x_1507 &  n_37750;
assign n_37753 = ~n_37751 & ~n_37752;
assign n_37754 =  n_26156 & ~n_36715;
assign n_37755 =  x_1506 & ~n_26156;
assign n_37756 = ~n_37754 & ~n_37755;
assign n_37757 =  x_1506 & ~n_37756;
assign n_37758 = ~x_1506 &  n_37756;
assign n_37759 = ~n_37757 & ~n_37758;
assign n_37760 =  n_26156 & ~n_36730;
assign n_37761 =  x_1505 & ~n_26156;
assign n_37762 = ~n_37760 & ~n_37761;
assign n_37763 =  x_1505 & ~n_37762;
assign n_37764 = ~x_1505 &  n_37762;
assign n_37765 = ~n_37763 & ~n_37764;
assign n_37766 =  n_26156 & ~n_36745;
assign n_37767 =  x_1504 & ~n_26156;
assign n_37768 = ~n_37766 & ~n_37767;
assign n_37769 =  x_1504 & ~n_37768;
assign n_37770 = ~x_1504 &  n_37768;
assign n_37771 = ~n_37769 & ~n_37770;
assign n_37772 =  n_26156 & ~n_36760;
assign n_37773 =  x_1503 & ~n_26156;
assign n_37774 = ~n_37772 & ~n_37773;
assign n_37775 =  x_1503 & ~n_37774;
assign n_37776 = ~x_1503 &  n_37774;
assign n_37777 = ~n_37775 & ~n_37776;
assign n_37778 =  n_26156 & ~n_36775;
assign n_37779 =  x_1502 & ~n_26156;
assign n_37780 = ~n_37778 & ~n_37779;
assign n_37781 =  x_1502 & ~n_37780;
assign n_37782 = ~x_1502 &  n_37780;
assign n_37783 = ~n_37781 & ~n_37782;
assign n_37784 =  n_26156 & ~n_36790;
assign n_37785 =  x_1501 & ~n_26156;
assign n_37786 = ~n_37784 & ~n_37785;
assign n_37787 =  x_1501 & ~n_37786;
assign n_37788 = ~x_1501 &  n_37786;
assign n_37789 = ~n_37787 & ~n_37788;
assign n_37790 =  n_26156 & ~n_36805;
assign n_37791 =  x_1500 & ~n_26156;
assign n_37792 = ~n_37790 & ~n_37791;
assign n_37793 =  x_1500 & ~n_37792;
assign n_37794 = ~x_1500 &  n_37792;
assign n_37795 = ~n_37793 & ~n_37794;
assign n_37796 =  n_26156 & ~n_36820;
assign n_37797 =  x_1499 & ~n_26156;
assign n_37798 = ~n_37796 & ~n_37797;
assign n_37799 =  x_1499 & ~n_37798;
assign n_37800 = ~x_1499 &  n_37798;
assign n_37801 = ~n_37799 & ~n_37800;
assign n_37802 =  n_26156 & ~n_36835;
assign n_37803 =  x_1498 & ~n_26156;
assign n_37804 = ~n_37802 & ~n_37803;
assign n_37805 =  x_1498 & ~n_37804;
assign n_37806 = ~x_1498 &  n_37804;
assign n_37807 = ~n_37805 & ~n_37806;
assign n_37808 =  n_26156 & ~n_36850;
assign n_37809 =  x_1497 & ~n_26156;
assign n_37810 = ~n_37808 & ~n_37809;
assign n_37811 =  x_1497 & ~n_37810;
assign n_37812 = ~x_1497 &  n_37810;
assign n_37813 = ~n_37811 & ~n_37812;
assign n_37814 =  n_26156 & ~n_36865;
assign n_37815 =  x_1496 & ~n_26156;
assign n_37816 = ~n_37814 & ~n_37815;
assign n_37817 =  x_1496 & ~n_37816;
assign n_37818 = ~x_1496 &  n_37816;
assign n_37819 = ~n_37817 & ~n_37818;
assign n_37820 =  n_26156 & ~n_36880;
assign n_37821 =  x_1495 & ~n_26156;
assign n_37822 = ~n_37820 & ~n_37821;
assign n_37823 =  x_1495 & ~n_37822;
assign n_37824 = ~x_1495 &  n_37822;
assign n_37825 = ~n_37823 & ~n_37824;
assign n_37826 =  n_26156 & ~n_36895;
assign n_37827 =  x_1494 & ~n_26156;
assign n_37828 = ~n_37826 & ~n_37827;
assign n_37829 =  x_1494 & ~n_37828;
assign n_37830 = ~x_1494 &  n_37828;
assign n_37831 = ~n_37829 & ~n_37830;
assign n_37832 =  n_26156 & ~n_36910;
assign n_37833 =  x_1493 & ~n_26156;
assign n_37834 = ~n_37832 & ~n_37833;
assign n_37835 =  x_1493 & ~n_37834;
assign n_37836 = ~x_1493 &  n_37834;
assign n_37837 = ~n_37835 & ~n_37836;
assign n_37838 =  n_26156 & ~n_36925;
assign n_37839 =  x_1492 & ~n_26156;
assign n_37840 = ~n_37838 & ~n_37839;
assign n_37841 =  x_1492 & ~n_37840;
assign n_37842 = ~x_1492 &  n_37840;
assign n_37843 = ~n_37841 & ~n_37842;
assign n_37844 =  n_26156 & ~n_36940;
assign n_37845 =  x_1491 & ~n_26156;
assign n_37846 = ~n_37844 & ~n_37845;
assign n_37847 =  x_1491 & ~n_37846;
assign n_37848 = ~x_1491 &  n_37846;
assign n_37849 = ~n_37847 & ~n_37848;
assign n_37850 =  n_26156 & ~n_36955;
assign n_37851 =  x_1490 & ~n_26156;
assign n_37852 = ~n_37850 & ~n_37851;
assign n_37853 =  x_1490 & ~n_37852;
assign n_37854 = ~x_1490 &  n_37852;
assign n_37855 = ~n_37853 & ~n_37854;
assign n_37856 =  n_26156 & ~n_36970;
assign n_37857 =  x_1489 & ~n_26156;
assign n_37858 = ~n_37856 & ~n_37857;
assign n_37859 =  x_1489 & ~n_37858;
assign n_37860 = ~x_1489 &  n_37858;
assign n_37861 = ~n_37859 & ~n_37860;
assign n_37862 =  n_26156 & ~n_36985;
assign n_37863 =  x_1488 & ~n_26156;
assign n_37864 = ~n_37862 & ~n_37863;
assign n_37865 =  x_1488 & ~n_37864;
assign n_37866 = ~x_1488 &  n_37864;
assign n_37867 = ~n_37865 & ~n_37866;
assign n_37868 =  n_26156 & ~n_37000;
assign n_37869 =  x_1487 & ~n_26156;
assign n_37870 = ~n_37868 & ~n_37869;
assign n_37871 =  x_1487 & ~n_37870;
assign n_37872 = ~x_1487 &  n_37870;
assign n_37873 = ~n_37871 & ~n_37872;
assign n_37874 =  n_26156 & ~n_37015;
assign n_37875 =  x_1486 & ~n_26156;
assign n_37876 = ~n_37874 & ~n_37875;
assign n_37877 =  x_1486 & ~n_37876;
assign n_37878 = ~x_1486 &  n_37876;
assign n_37879 = ~n_37877 & ~n_37878;
assign n_37880 =  n_26156 & ~n_37030;
assign n_37881 =  x_1485 & ~n_26156;
assign n_37882 = ~n_37880 & ~n_37881;
assign n_37883 =  x_1485 & ~n_37882;
assign n_37884 = ~x_1485 &  n_37882;
assign n_37885 = ~n_37883 & ~n_37884;
assign n_37886 =  n_26156 & ~n_37045;
assign n_37887 =  x_1484 & ~n_26156;
assign n_37888 = ~n_37886 & ~n_37887;
assign n_37889 =  x_1484 & ~n_37888;
assign n_37890 = ~x_1484 &  n_37888;
assign n_37891 = ~n_37889 & ~n_37890;
assign n_37892 =  n_26156 & ~n_37060;
assign n_37893 =  x_1483 & ~n_26156;
assign n_37894 = ~n_37892 & ~n_37893;
assign n_37895 =  x_1483 & ~n_37894;
assign n_37896 = ~x_1483 &  n_37894;
assign n_37897 = ~n_37895 & ~n_37896;
assign n_37898 =  x_1482 & ~n_23255;
assign n_37899 =  i_32 &  n_23255;
assign n_37900 = ~n_37898 & ~n_37899;
assign n_37901 =  x_1482 & ~n_37900;
assign n_37902 = ~x_1482 &  n_37900;
assign n_37903 = ~n_37901 & ~n_37902;
assign n_37904 =  x_1481 & ~n_23255;
assign n_37905 =  i_31 &  n_23255;
assign n_37906 = ~n_37904 & ~n_37905;
assign n_37907 =  x_1481 & ~n_37906;
assign n_37908 = ~x_1481 &  n_37906;
assign n_37909 = ~n_37907 & ~n_37908;
assign n_37910 =  x_1480 & ~n_23255;
assign n_37911 =  i_30 &  n_23255;
assign n_37912 = ~n_37910 & ~n_37911;
assign n_37913 =  x_1480 & ~n_37912;
assign n_37914 = ~x_1480 &  n_37912;
assign n_37915 = ~n_37913 & ~n_37914;
assign n_37916 =  x_1479 & ~n_23255;
assign n_37917 =  i_29 &  n_23255;
assign n_37918 = ~n_37916 & ~n_37917;
assign n_37919 =  x_1479 & ~n_37918;
assign n_37920 = ~x_1479 &  n_37918;
assign n_37921 = ~n_37919 & ~n_37920;
assign n_37922 =  x_1478 & ~n_23255;
assign n_37923 =  i_28 &  n_23255;
assign n_37924 = ~n_37922 & ~n_37923;
assign n_37925 =  x_1478 & ~n_37924;
assign n_37926 = ~x_1478 &  n_37924;
assign n_37927 = ~n_37925 & ~n_37926;
assign n_37928 =  x_1477 & ~n_23255;
assign n_37929 =  i_27 &  n_23255;
assign n_37930 = ~n_37928 & ~n_37929;
assign n_37931 =  x_1477 & ~n_37930;
assign n_37932 = ~x_1477 &  n_37930;
assign n_37933 = ~n_37931 & ~n_37932;
assign n_37934 =  x_1476 & ~n_23255;
assign n_37935 =  i_26 &  n_23255;
assign n_37936 = ~n_37934 & ~n_37935;
assign n_37937 =  x_1476 & ~n_37936;
assign n_37938 = ~x_1476 &  n_37936;
assign n_37939 = ~n_37937 & ~n_37938;
assign n_37940 =  x_1475 & ~n_23255;
assign n_37941 =  i_25 &  n_23255;
assign n_37942 = ~n_37940 & ~n_37941;
assign n_37943 =  x_1475 & ~n_37942;
assign n_37944 = ~x_1475 &  n_37942;
assign n_37945 = ~n_37943 & ~n_37944;
assign n_37946 =  x_1474 & ~n_23255;
assign n_37947 =  i_24 &  n_23255;
assign n_37948 = ~n_37946 & ~n_37947;
assign n_37949 =  x_1474 & ~n_37948;
assign n_37950 = ~x_1474 &  n_37948;
assign n_37951 = ~n_37949 & ~n_37950;
assign n_37952 =  x_1473 & ~n_23255;
assign n_37953 =  i_23 &  n_23255;
assign n_37954 = ~n_37952 & ~n_37953;
assign n_37955 =  x_1473 & ~n_37954;
assign n_37956 = ~x_1473 &  n_37954;
assign n_37957 = ~n_37955 & ~n_37956;
assign n_37958 =  x_1472 & ~n_23255;
assign n_37959 =  i_22 &  n_23255;
assign n_37960 = ~n_37958 & ~n_37959;
assign n_37961 =  x_1472 & ~n_37960;
assign n_37962 = ~x_1472 &  n_37960;
assign n_37963 = ~n_37961 & ~n_37962;
assign n_37964 =  x_1471 & ~n_23255;
assign n_37965 =  i_21 &  n_23255;
assign n_37966 = ~n_37964 & ~n_37965;
assign n_37967 =  x_1471 & ~n_37966;
assign n_37968 = ~x_1471 &  n_37966;
assign n_37969 = ~n_37967 & ~n_37968;
assign n_37970 =  x_1470 & ~n_23255;
assign n_37971 =  i_20 &  n_23255;
assign n_37972 = ~n_37970 & ~n_37971;
assign n_37973 =  x_1470 & ~n_37972;
assign n_37974 = ~x_1470 &  n_37972;
assign n_37975 = ~n_37973 & ~n_37974;
assign n_37976 =  x_1469 & ~n_23255;
assign n_37977 =  i_19 &  n_23255;
assign n_37978 = ~n_37976 & ~n_37977;
assign n_37979 =  x_1469 & ~n_37978;
assign n_37980 = ~x_1469 &  n_37978;
assign n_37981 = ~n_37979 & ~n_37980;
assign n_37982 =  x_1468 & ~n_23255;
assign n_37983 =  i_18 &  n_23255;
assign n_37984 = ~n_37982 & ~n_37983;
assign n_37985 =  x_1468 & ~n_37984;
assign n_37986 = ~x_1468 &  n_37984;
assign n_37987 = ~n_37985 & ~n_37986;
assign n_37988 =  x_1467 & ~n_23255;
assign n_37989 =  i_17 &  n_23255;
assign n_37990 = ~n_37988 & ~n_37989;
assign n_37991 =  x_1467 & ~n_37990;
assign n_37992 = ~x_1467 &  n_37990;
assign n_37993 = ~n_37991 & ~n_37992;
assign n_37994 =  x_1466 & ~n_23255;
assign n_37995 =  i_16 &  n_23255;
assign n_37996 = ~n_37994 & ~n_37995;
assign n_37997 =  x_1466 & ~n_37996;
assign n_37998 = ~x_1466 &  n_37996;
assign n_37999 = ~n_37997 & ~n_37998;
assign n_38000 =  x_1465 & ~n_23255;
assign n_38001 =  i_15 &  n_23255;
assign n_38002 = ~n_38000 & ~n_38001;
assign n_38003 =  x_1465 & ~n_38002;
assign n_38004 = ~x_1465 &  n_38002;
assign n_38005 = ~n_38003 & ~n_38004;
assign n_38006 =  x_1464 & ~n_23255;
assign n_38007 =  i_14 &  n_23255;
assign n_38008 = ~n_38006 & ~n_38007;
assign n_38009 =  x_1464 & ~n_38008;
assign n_38010 = ~x_1464 &  n_38008;
assign n_38011 = ~n_38009 & ~n_38010;
assign n_38012 =  x_1463 & ~n_23255;
assign n_38013 =  i_13 &  n_23255;
assign n_38014 = ~n_38012 & ~n_38013;
assign n_38015 =  x_1463 & ~n_38014;
assign n_38016 = ~x_1463 &  n_38014;
assign n_38017 = ~n_38015 & ~n_38016;
assign n_38018 =  x_1462 & ~n_23255;
assign n_38019 =  i_12 &  n_23255;
assign n_38020 = ~n_38018 & ~n_38019;
assign n_38021 =  x_1462 & ~n_38020;
assign n_38022 = ~x_1462 &  n_38020;
assign n_38023 = ~n_38021 & ~n_38022;
assign n_38024 =  x_1461 & ~n_23255;
assign n_38025 =  i_11 &  n_23255;
assign n_38026 = ~n_38024 & ~n_38025;
assign n_38027 =  x_1461 & ~n_38026;
assign n_38028 = ~x_1461 &  n_38026;
assign n_38029 = ~n_38027 & ~n_38028;
assign n_38030 =  x_1460 & ~n_23255;
assign n_38031 =  i_10 &  n_23255;
assign n_38032 = ~n_38030 & ~n_38031;
assign n_38033 =  x_1460 & ~n_38032;
assign n_38034 = ~x_1460 &  n_38032;
assign n_38035 = ~n_38033 & ~n_38034;
assign n_38036 =  x_1459 & ~n_23255;
assign n_38037 =  i_9 &  n_23255;
assign n_38038 = ~n_38036 & ~n_38037;
assign n_38039 =  x_1459 & ~n_38038;
assign n_38040 = ~x_1459 &  n_38038;
assign n_38041 = ~n_38039 & ~n_38040;
assign n_38042 =  x_1458 & ~n_23255;
assign n_38043 =  i_8 &  n_23255;
assign n_38044 = ~n_38042 & ~n_38043;
assign n_38045 =  x_1458 & ~n_38044;
assign n_38046 = ~x_1458 &  n_38044;
assign n_38047 = ~n_38045 & ~n_38046;
assign n_38048 =  x_1457 & ~n_23255;
assign n_38049 =  i_7 &  n_23255;
assign n_38050 = ~n_38048 & ~n_38049;
assign n_38051 =  x_1457 & ~n_38050;
assign n_38052 = ~x_1457 &  n_38050;
assign n_38053 = ~n_38051 & ~n_38052;
assign n_38054 =  x_1456 & ~n_23255;
assign n_38055 =  i_6 &  n_23255;
assign n_38056 = ~n_38054 & ~n_38055;
assign n_38057 =  x_1456 & ~n_38056;
assign n_38058 = ~x_1456 &  n_38056;
assign n_38059 = ~n_38057 & ~n_38058;
assign n_38060 =  x_1455 & ~n_23255;
assign n_38061 =  i_5 &  n_23255;
assign n_38062 = ~n_38060 & ~n_38061;
assign n_38063 =  x_1455 & ~n_38062;
assign n_38064 = ~x_1455 &  n_38062;
assign n_38065 = ~n_38063 & ~n_38064;
assign n_38066 =  x_1454 & ~n_23255;
assign n_38067 =  i_4 &  n_23255;
assign n_38068 = ~n_38066 & ~n_38067;
assign n_38069 =  x_1454 & ~n_38068;
assign n_38070 = ~x_1454 &  n_38068;
assign n_38071 = ~n_38069 & ~n_38070;
assign n_38072 =  x_1453 & ~n_23255;
assign n_38073 =  i_3 &  n_23255;
assign n_38074 = ~n_38072 & ~n_38073;
assign n_38075 =  x_1453 & ~n_38074;
assign n_38076 = ~x_1453 &  n_38074;
assign n_38077 = ~n_38075 & ~n_38076;
assign n_38078 =  x_1452 & ~n_23255;
assign n_38079 =  i_2 &  n_23255;
assign n_38080 = ~n_38078 & ~n_38079;
assign n_38081 =  x_1452 & ~n_38080;
assign n_38082 = ~x_1452 &  n_38080;
assign n_38083 = ~n_38081 & ~n_38082;
assign n_38084 =  x_1451 & ~n_23255;
assign n_38085 =  i_1 &  n_23255;
assign n_38086 = ~n_38084 & ~n_38085;
assign n_38087 =  x_1451 & ~n_38086;
assign n_38088 = ~x_1451 &  n_38086;
assign n_38089 = ~n_38087 & ~n_38088;
assign n_38090 =  x_1450 & ~n_23946;
assign n_38091 =  i_32 &  n_23946;
assign n_38092 = ~n_38090 & ~n_38091;
assign n_38093 =  x_1450 & ~n_38092;
assign n_38094 = ~x_1450 &  n_38092;
assign n_38095 = ~n_38093 & ~n_38094;
assign n_38096 =  x_1449 & ~n_23946;
assign n_38097 =  i_31 &  n_23946;
assign n_38098 = ~n_38096 & ~n_38097;
assign n_38099 =  x_1449 & ~n_38098;
assign n_38100 = ~x_1449 &  n_38098;
assign n_38101 = ~n_38099 & ~n_38100;
assign n_38102 =  x_1448 & ~n_23946;
assign n_38103 =  i_30 &  n_23946;
assign n_38104 = ~n_38102 & ~n_38103;
assign n_38105 =  x_1448 & ~n_38104;
assign n_38106 = ~x_1448 &  n_38104;
assign n_38107 = ~n_38105 & ~n_38106;
assign n_38108 =  x_1447 & ~n_23946;
assign n_38109 =  i_29 &  n_23946;
assign n_38110 = ~n_38108 & ~n_38109;
assign n_38111 =  x_1447 & ~n_38110;
assign n_38112 = ~x_1447 &  n_38110;
assign n_38113 = ~n_38111 & ~n_38112;
assign n_38114 =  x_1446 & ~n_23946;
assign n_38115 =  i_28 &  n_23946;
assign n_38116 = ~n_38114 & ~n_38115;
assign n_38117 =  x_1446 & ~n_38116;
assign n_38118 = ~x_1446 &  n_38116;
assign n_38119 = ~n_38117 & ~n_38118;
assign n_38120 =  x_1445 & ~n_23946;
assign n_38121 =  i_27 &  n_23946;
assign n_38122 = ~n_38120 & ~n_38121;
assign n_38123 =  x_1445 & ~n_38122;
assign n_38124 = ~x_1445 &  n_38122;
assign n_38125 = ~n_38123 & ~n_38124;
assign n_38126 =  x_1444 & ~n_23946;
assign n_38127 =  i_26 &  n_23946;
assign n_38128 = ~n_38126 & ~n_38127;
assign n_38129 =  x_1444 & ~n_38128;
assign n_38130 = ~x_1444 &  n_38128;
assign n_38131 = ~n_38129 & ~n_38130;
assign n_38132 =  x_1443 & ~n_23946;
assign n_38133 =  i_25 &  n_23946;
assign n_38134 = ~n_38132 & ~n_38133;
assign n_38135 =  x_1443 & ~n_38134;
assign n_38136 = ~x_1443 &  n_38134;
assign n_38137 = ~n_38135 & ~n_38136;
assign n_38138 =  x_1442 & ~n_23946;
assign n_38139 =  i_24 &  n_23946;
assign n_38140 = ~n_38138 & ~n_38139;
assign n_38141 =  x_1442 & ~n_38140;
assign n_38142 = ~x_1442 &  n_38140;
assign n_38143 = ~n_38141 & ~n_38142;
assign n_38144 =  x_1441 & ~n_23946;
assign n_38145 =  i_23 &  n_23946;
assign n_38146 = ~n_38144 & ~n_38145;
assign n_38147 =  x_1441 & ~n_38146;
assign n_38148 = ~x_1441 &  n_38146;
assign n_38149 = ~n_38147 & ~n_38148;
assign n_38150 =  x_1440 & ~n_23946;
assign n_38151 =  i_22 &  n_23946;
assign n_38152 = ~n_38150 & ~n_38151;
assign n_38153 =  x_1440 & ~n_38152;
assign n_38154 = ~x_1440 &  n_38152;
assign n_38155 = ~n_38153 & ~n_38154;
assign n_38156 =  x_1439 & ~n_23946;
assign n_38157 =  i_21 &  n_23946;
assign n_38158 = ~n_38156 & ~n_38157;
assign n_38159 =  x_1439 & ~n_38158;
assign n_38160 = ~x_1439 &  n_38158;
assign n_38161 = ~n_38159 & ~n_38160;
assign n_38162 =  x_1438 & ~n_23946;
assign n_38163 =  i_20 &  n_23946;
assign n_38164 = ~n_38162 & ~n_38163;
assign n_38165 =  x_1438 & ~n_38164;
assign n_38166 = ~x_1438 &  n_38164;
assign n_38167 = ~n_38165 & ~n_38166;
assign n_38168 =  x_1437 & ~n_23946;
assign n_38169 =  i_19 &  n_23946;
assign n_38170 = ~n_38168 & ~n_38169;
assign n_38171 =  x_1437 & ~n_38170;
assign n_38172 = ~x_1437 &  n_38170;
assign n_38173 = ~n_38171 & ~n_38172;
assign n_38174 =  x_1436 & ~n_23946;
assign n_38175 =  i_18 &  n_23946;
assign n_38176 = ~n_38174 & ~n_38175;
assign n_38177 =  x_1436 & ~n_38176;
assign n_38178 = ~x_1436 &  n_38176;
assign n_38179 = ~n_38177 & ~n_38178;
assign n_38180 =  x_1435 & ~n_23946;
assign n_38181 =  i_17 &  n_23946;
assign n_38182 = ~n_38180 & ~n_38181;
assign n_38183 =  x_1435 & ~n_38182;
assign n_38184 = ~x_1435 &  n_38182;
assign n_38185 = ~n_38183 & ~n_38184;
assign n_38186 =  x_1434 & ~n_23946;
assign n_38187 =  i_16 &  n_23946;
assign n_38188 = ~n_38186 & ~n_38187;
assign n_38189 =  x_1434 & ~n_38188;
assign n_38190 = ~x_1434 &  n_38188;
assign n_38191 = ~n_38189 & ~n_38190;
assign n_38192 =  x_1433 & ~n_23946;
assign n_38193 =  i_15 &  n_23946;
assign n_38194 = ~n_38192 & ~n_38193;
assign n_38195 =  x_1433 & ~n_38194;
assign n_38196 = ~x_1433 &  n_38194;
assign n_38197 = ~n_38195 & ~n_38196;
assign n_38198 =  x_1432 & ~n_23946;
assign n_38199 =  i_14 &  n_23946;
assign n_38200 = ~n_38198 & ~n_38199;
assign n_38201 =  x_1432 & ~n_38200;
assign n_38202 = ~x_1432 &  n_38200;
assign n_38203 = ~n_38201 & ~n_38202;
assign n_38204 =  x_1431 & ~n_23946;
assign n_38205 =  i_13 &  n_23946;
assign n_38206 = ~n_38204 & ~n_38205;
assign n_38207 =  x_1431 & ~n_38206;
assign n_38208 = ~x_1431 &  n_38206;
assign n_38209 = ~n_38207 & ~n_38208;
assign n_38210 =  x_1430 & ~n_23946;
assign n_38211 =  i_12 &  n_23946;
assign n_38212 = ~n_38210 & ~n_38211;
assign n_38213 =  x_1430 & ~n_38212;
assign n_38214 = ~x_1430 &  n_38212;
assign n_38215 = ~n_38213 & ~n_38214;
assign n_38216 =  x_1429 & ~n_23946;
assign n_38217 =  i_11 &  n_23946;
assign n_38218 = ~n_38216 & ~n_38217;
assign n_38219 =  x_1429 & ~n_38218;
assign n_38220 = ~x_1429 &  n_38218;
assign n_38221 = ~n_38219 & ~n_38220;
assign n_38222 =  x_1428 & ~n_23946;
assign n_38223 =  i_10 &  n_23946;
assign n_38224 = ~n_38222 & ~n_38223;
assign n_38225 =  x_1428 & ~n_38224;
assign n_38226 = ~x_1428 &  n_38224;
assign n_38227 = ~n_38225 & ~n_38226;
assign n_38228 =  x_1427 & ~n_23946;
assign n_38229 =  i_9 &  n_23946;
assign n_38230 = ~n_38228 & ~n_38229;
assign n_38231 =  x_1427 & ~n_38230;
assign n_38232 = ~x_1427 &  n_38230;
assign n_38233 = ~n_38231 & ~n_38232;
assign n_38234 =  x_1426 & ~n_23946;
assign n_38235 =  i_8 &  n_23946;
assign n_38236 = ~n_38234 & ~n_38235;
assign n_38237 =  x_1426 & ~n_38236;
assign n_38238 = ~x_1426 &  n_38236;
assign n_38239 = ~n_38237 & ~n_38238;
assign n_38240 =  x_1425 & ~n_23946;
assign n_38241 =  i_7 &  n_23946;
assign n_38242 = ~n_38240 & ~n_38241;
assign n_38243 =  x_1425 & ~n_38242;
assign n_38244 = ~x_1425 &  n_38242;
assign n_38245 = ~n_38243 & ~n_38244;
assign n_38246 =  x_1424 & ~n_23946;
assign n_38247 =  i_6 &  n_23946;
assign n_38248 = ~n_38246 & ~n_38247;
assign n_38249 =  x_1424 & ~n_38248;
assign n_38250 = ~x_1424 &  n_38248;
assign n_38251 = ~n_38249 & ~n_38250;
assign n_38252 =  x_1423 & ~n_23946;
assign n_38253 =  i_5 &  n_23946;
assign n_38254 = ~n_38252 & ~n_38253;
assign n_38255 =  x_1423 & ~n_38254;
assign n_38256 = ~x_1423 &  n_38254;
assign n_38257 = ~n_38255 & ~n_38256;
assign n_38258 =  x_1422 & ~n_23946;
assign n_38259 =  i_4 &  n_23946;
assign n_38260 = ~n_38258 & ~n_38259;
assign n_38261 =  x_1422 & ~n_38260;
assign n_38262 = ~x_1422 &  n_38260;
assign n_38263 = ~n_38261 & ~n_38262;
assign n_38264 =  x_1421 & ~n_23946;
assign n_38265 =  i_3 &  n_23946;
assign n_38266 = ~n_38264 & ~n_38265;
assign n_38267 =  x_1421 & ~n_38266;
assign n_38268 = ~x_1421 &  n_38266;
assign n_38269 = ~n_38267 & ~n_38268;
assign n_38270 =  x_1420 & ~n_23946;
assign n_38271 =  i_2 &  n_23946;
assign n_38272 = ~n_38270 & ~n_38271;
assign n_38273 =  x_1420 & ~n_38272;
assign n_38274 = ~x_1420 &  n_38272;
assign n_38275 = ~n_38273 & ~n_38274;
assign n_38276 =  x_1419 & ~n_23946;
assign n_38277 =  i_1 &  n_23946;
assign n_38278 = ~n_38276 & ~n_38277;
assign n_38279 =  x_1419 & ~n_38278;
assign n_38280 = ~x_1419 &  n_38278;
assign n_38281 = ~n_38279 & ~n_38280;
assign n_38282 =  n_153 &  n_24581;
assign n_38283 = ~n_28296 & ~n_38282;
assign n_38284 =  n_24581 & ~n_25952;
assign n_38285 =  x_1418 & ~n_38284;
assign n_38286 =  n_38283 & ~n_38285;
assign n_38287 =  x_1418 & ~n_38286;
assign n_38288 = ~x_1418 &  n_38286;
assign n_38289 = ~n_38287 & ~n_38288;
assign n_38290 = ~n_38284 &  n_38283;
assign n_38291 =  x_1417 &  n_38290;
assign n_38292 =  x_1417 &  n_38291;
assign n_38293 = ~x_1417 & ~n_38291;
assign n_38294 = ~n_38292 & ~n_38293;
assign n_38295 =  x_1416 &  n_38290;
assign n_38296 =  x_1416 &  n_38295;
assign n_38297 = ~x_1416 & ~n_38295;
assign n_38298 = ~n_38296 & ~n_38297;
assign n_38299 =  x_1415 &  n_38290;
assign n_38300 =  x_1415 &  n_38299;
assign n_38301 = ~x_1415 & ~n_38299;
assign n_38302 = ~n_38300 & ~n_38301;
assign n_38303 =  x_1414 &  n_38290;
assign n_38304 =  x_1414 &  n_38303;
assign n_38305 = ~x_1414 & ~n_38303;
assign n_38306 = ~n_38304 & ~n_38305;
assign n_38307 =  x_1413 &  n_38290;
assign n_38308 =  x_1413 &  n_38307;
assign n_38309 = ~x_1413 & ~n_38307;
assign n_38310 = ~n_38308 & ~n_38309;
assign n_38311 =  x_1412 &  n_38290;
assign n_38312 =  x_1412 &  n_38311;
assign n_38313 = ~x_1412 & ~n_38311;
assign n_38314 = ~n_38312 & ~n_38313;
assign n_38315 =  x_1411 &  n_38290;
assign n_38316 =  x_1411 &  n_38315;
assign n_38317 = ~x_1411 & ~n_38315;
assign n_38318 = ~n_38316 & ~n_38317;
assign n_38319 =  x_1410 &  n_38290;
assign n_38320 =  x_1410 &  n_38319;
assign n_38321 = ~x_1410 & ~n_38319;
assign n_38322 = ~n_38320 & ~n_38321;
assign n_38323 =  x_1409 &  n_38290;
assign n_38324 =  x_1409 &  n_38323;
assign n_38325 = ~x_1409 & ~n_38323;
assign n_38326 = ~n_38324 & ~n_38325;
assign n_38327 =  x_1408 &  n_38290;
assign n_38328 =  x_1408 &  n_38327;
assign n_38329 = ~x_1408 & ~n_38327;
assign n_38330 = ~n_38328 & ~n_38329;
assign n_38331 =  x_1407 &  n_38290;
assign n_38332 =  x_1407 &  n_38331;
assign n_38333 = ~x_1407 & ~n_38331;
assign n_38334 = ~n_38332 & ~n_38333;
assign n_38335 =  x_1406 &  n_38290;
assign n_38336 =  x_1406 &  n_38335;
assign n_38337 = ~x_1406 & ~n_38335;
assign n_38338 = ~n_38336 & ~n_38337;
assign n_38339 =  x_1405 &  n_38290;
assign n_38340 =  x_1405 &  n_38339;
assign n_38341 = ~x_1405 & ~n_38339;
assign n_38342 = ~n_38340 & ~n_38341;
assign n_38343 =  x_1404 &  n_38290;
assign n_38344 =  x_1404 &  n_38343;
assign n_38345 = ~x_1404 & ~n_38343;
assign n_38346 = ~n_38344 & ~n_38345;
assign n_38347 =  x_1403 &  n_38290;
assign n_38348 =  x_1403 &  n_38347;
assign n_38349 = ~x_1403 & ~n_38347;
assign n_38350 = ~n_38348 & ~n_38349;
assign n_38351 =  x_1402 &  n_38290;
assign n_38352 =  x_1402 &  n_38351;
assign n_38353 = ~x_1402 & ~n_38351;
assign n_38354 = ~n_38352 & ~n_38353;
assign n_38355 =  x_1401 &  n_38290;
assign n_38356 =  x_1401 &  n_38355;
assign n_38357 = ~x_1401 & ~n_38355;
assign n_38358 = ~n_38356 & ~n_38357;
assign n_38359 =  x_1400 &  n_38290;
assign n_38360 =  x_1400 &  n_38359;
assign n_38361 = ~x_1400 & ~n_38359;
assign n_38362 = ~n_38360 & ~n_38361;
assign n_38363 =  x_1399 &  n_38290;
assign n_38364 =  x_1399 &  n_38363;
assign n_38365 = ~x_1399 & ~n_38363;
assign n_38366 = ~n_38364 & ~n_38365;
assign n_38367 =  x_1398 &  n_38290;
assign n_38368 =  x_1398 &  n_38367;
assign n_38369 = ~x_1398 & ~n_38367;
assign n_38370 = ~n_38368 & ~n_38369;
assign n_38371 =  x_1397 &  n_38290;
assign n_38372 =  x_1397 &  n_38371;
assign n_38373 = ~x_1397 & ~n_38371;
assign n_38374 = ~n_38372 & ~n_38373;
assign n_38375 =  x_1396 &  n_38290;
assign n_38376 =  x_1396 &  n_38375;
assign n_38377 = ~x_1396 & ~n_38375;
assign n_38378 = ~n_38376 & ~n_38377;
assign n_38379 =  x_1395 &  n_38290;
assign n_38380 =  x_1395 &  n_38379;
assign n_38381 = ~x_1395 & ~n_38379;
assign n_38382 = ~n_38380 & ~n_38381;
assign n_38383 =  x_1394 &  n_38290;
assign n_38384 =  x_1394 &  n_38383;
assign n_38385 = ~x_1394 & ~n_38383;
assign n_38386 = ~n_38384 & ~n_38385;
assign n_38387 =  x_1393 &  n_38290;
assign n_38388 =  x_1393 &  n_38387;
assign n_38389 = ~x_1393 & ~n_38387;
assign n_38390 = ~n_38388 & ~n_38389;
assign n_38391 =  x_1392 &  n_38290;
assign n_38392 =  x_1392 &  n_38391;
assign n_38393 = ~x_1392 & ~n_38391;
assign n_38394 = ~n_38392 & ~n_38393;
assign n_38395 =  x_1391 &  n_38290;
assign n_38396 =  x_1391 &  n_38395;
assign n_38397 = ~x_1391 & ~n_38395;
assign n_38398 = ~n_38396 & ~n_38397;
assign n_38399 =  x_1390 &  n_38290;
assign n_38400 =  x_1390 &  n_38399;
assign n_38401 = ~x_1390 & ~n_38399;
assign n_38402 = ~n_38400 & ~n_38401;
assign n_38403 =  x_1389 &  n_38290;
assign n_38404 =  x_1389 &  n_38403;
assign n_38405 = ~x_1389 & ~n_38403;
assign n_38406 = ~n_38404 & ~n_38405;
assign n_38407 =  x_1388 &  n_38290;
assign n_38408 =  x_1388 &  n_38407;
assign n_38409 = ~x_1388 & ~n_38407;
assign n_38410 = ~n_38408 & ~n_38409;
assign n_38411 =  x_1387 &  n_38290;
assign n_38412 =  x_1387 &  n_38411;
assign n_38413 = ~x_1387 & ~n_38411;
assign n_38414 = ~n_38412 & ~n_38413;
assign n_38415 =  x_1386 & ~n_26318;
assign n_38416 =  i_32 &  n_26318;
assign n_38417 = ~n_38415 & ~n_38416;
assign n_38418 =  x_1386 & ~n_38417;
assign n_38419 = ~x_1386 &  n_38417;
assign n_38420 = ~n_38418 & ~n_38419;
assign n_38421 =  x_1385 & ~n_26318;
assign n_38422 =  i_31 &  n_26318;
assign n_38423 = ~n_38421 & ~n_38422;
assign n_38424 =  x_1385 & ~n_38423;
assign n_38425 = ~x_1385 &  n_38423;
assign n_38426 = ~n_38424 & ~n_38425;
assign n_38427 =  x_1384 & ~n_26318;
assign n_38428 =  i_30 &  n_26318;
assign n_38429 = ~n_38427 & ~n_38428;
assign n_38430 =  x_1384 & ~n_38429;
assign n_38431 = ~x_1384 &  n_38429;
assign n_38432 = ~n_38430 & ~n_38431;
assign n_38433 =  x_1383 & ~n_26318;
assign n_38434 =  i_29 &  n_26318;
assign n_38435 = ~n_38433 & ~n_38434;
assign n_38436 =  x_1383 & ~n_38435;
assign n_38437 = ~x_1383 &  n_38435;
assign n_38438 = ~n_38436 & ~n_38437;
assign n_38439 =  x_1382 & ~n_26318;
assign n_38440 =  i_28 &  n_26318;
assign n_38441 = ~n_38439 & ~n_38440;
assign n_38442 =  x_1382 & ~n_38441;
assign n_38443 = ~x_1382 &  n_38441;
assign n_38444 = ~n_38442 & ~n_38443;
assign n_38445 =  x_1381 & ~n_26318;
assign n_38446 =  i_27 &  n_26318;
assign n_38447 = ~n_38445 & ~n_38446;
assign n_38448 =  x_1381 & ~n_38447;
assign n_38449 = ~x_1381 &  n_38447;
assign n_38450 = ~n_38448 & ~n_38449;
assign n_38451 =  x_1380 & ~n_26318;
assign n_38452 =  i_26 &  n_26318;
assign n_38453 = ~n_38451 & ~n_38452;
assign n_38454 =  x_1380 & ~n_38453;
assign n_38455 = ~x_1380 &  n_38453;
assign n_38456 = ~n_38454 & ~n_38455;
assign n_38457 =  x_1379 & ~n_26318;
assign n_38458 =  i_25 &  n_26318;
assign n_38459 = ~n_38457 & ~n_38458;
assign n_38460 =  x_1379 & ~n_38459;
assign n_38461 = ~x_1379 &  n_38459;
assign n_38462 = ~n_38460 & ~n_38461;
assign n_38463 =  x_1378 & ~n_26318;
assign n_38464 =  i_24 &  n_26318;
assign n_38465 = ~n_38463 & ~n_38464;
assign n_38466 =  x_1378 & ~n_38465;
assign n_38467 = ~x_1378 &  n_38465;
assign n_38468 = ~n_38466 & ~n_38467;
assign n_38469 =  x_1377 & ~n_26318;
assign n_38470 =  i_23 &  n_26318;
assign n_38471 = ~n_38469 & ~n_38470;
assign n_38472 =  x_1377 & ~n_38471;
assign n_38473 = ~x_1377 &  n_38471;
assign n_38474 = ~n_38472 & ~n_38473;
assign n_38475 =  x_1376 & ~n_26318;
assign n_38476 =  i_22 &  n_26318;
assign n_38477 = ~n_38475 & ~n_38476;
assign n_38478 =  x_1376 & ~n_38477;
assign n_38479 = ~x_1376 &  n_38477;
assign n_38480 = ~n_38478 & ~n_38479;
assign n_38481 =  x_1375 & ~n_26318;
assign n_38482 =  i_21 &  n_26318;
assign n_38483 = ~n_38481 & ~n_38482;
assign n_38484 =  x_1375 & ~n_38483;
assign n_38485 = ~x_1375 &  n_38483;
assign n_38486 = ~n_38484 & ~n_38485;
assign n_38487 =  x_1374 & ~n_26318;
assign n_38488 =  i_20 &  n_26318;
assign n_38489 = ~n_38487 & ~n_38488;
assign n_38490 =  x_1374 & ~n_38489;
assign n_38491 = ~x_1374 &  n_38489;
assign n_38492 = ~n_38490 & ~n_38491;
assign n_38493 =  x_1373 & ~n_26318;
assign n_38494 =  i_19 &  n_26318;
assign n_38495 = ~n_38493 & ~n_38494;
assign n_38496 =  x_1373 & ~n_38495;
assign n_38497 = ~x_1373 &  n_38495;
assign n_38498 = ~n_38496 & ~n_38497;
assign n_38499 =  x_1372 & ~n_26318;
assign n_38500 =  i_18 &  n_26318;
assign n_38501 = ~n_38499 & ~n_38500;
assign n_38502 =  x_1372 & ~n_38501;
assign n_38503 = ~x_1372 &  n_38501;
assign n_38504 = ~n_38502 & ~n_38503;
assign n_38505 =  x_1371 & ~n_26318;
assign n_38506 =  i_17 &  n_26318;
assign n_38507 = ~n_38505 & ~n_38506;
assign n_38508 =  x_1371 & ~n_38507;
assign n_38509 = ~x_1371 &  n_38507;
assign n_38510 = ~n_38508 & ~n_38509;
assign n_38511 =  x_1370 & ~n_26318;
assign n_38512 =  i_16 &  n_26318;
assign n_38513 = ~n_38511 & ~n_38512;
assign n_38514 =  x_1370 & ~n_38513;
assign n_38515 = ~x_1370 &  n_38513;
assign n_38516 = ~n_38514 & ~n_38515;
assign n_38517 =  x_1369 & ~n_26318;
assign n_38518 =  i_15 &  n_26318;
assign n_38519 = ~n_38517 & ~n_38518;
assign n_38520 =  x_1369 & ~n_38519;
assign n_38521 = ~x_1369 &  n_38519;
assign n_38522 = ~n_38520 & ~n_38521;
assign n_38523 =  x_1368 & ~n_26318;
assign n_38524 =  i_14 &  n_26318;
assign n_38525 = ~n_38523 & ~n_38524;
assign n_38526 =  x_1368 & ~n_38525;
assign n_38527 = ~x_1368 &  n_38525;
assign n_38528 = ~n_38526 & ~n_38527;
assign n_38529 =  x_1367 & ~n_26318;
assign n_38530 =  i_13 &  n_26318;
assign n_38531 = ~n_38529 & ~n_38530;
assign n_38532 =  x_1367 & ~n_38531;
assign n_38533 = ~x_1367 &  n_38531;
assign n_38534 = ~n_38532 & ~n_38533;
assign n_38535 =  x_1366 & ~n_26318;
assign n_38536 =  i_12 &  n_26318;
assign n_38537 = ~n_38535 & ~n_38536;
assign n_38538 =  x_1366 & ~n_38537;
assign n_38539 = ~x_1366 &  n_38537;
assign n_38540 = ~n_38538 & ~n_38539;
assign n_38541 =  x_1365 & ~n_26318;
assign n_38542 =  i_11 &  n_26318;
assign n_38543 = ~n_38541 & ~n_38542;
assign n_38544 =  x_1365 & ~n_38543;
assign n_38545 = ~x_1365 &  n_38543;
assign n_38546 = ~n_38544 & ~n_38545;
assign n_38547 =  x_1364 & ~n_26318;
assign n_38548 =  i_10 &  n_26318;
assign n_38549 = ~n_38547 & ~n_38548;
assign n_38550 =  x_1364 & ~n_38549;
assign n_38551 = ~x_1364 &  n_38549;
assign n_38552 = ~n_38550 & ~n_38551;
assign n_38553 =  x_1363 & ~n_26318;
assign n_38554 =  i_9 &  n_26318;
assign n_38555 = ~n_38553 & ~n_38554;
assign n_38556 =  x_1363 & ~n_38555;
assign n_38557 = ~x_1363 &  n_38555;
assign n_38558 = ~n_38556 & ~n_38557;
assign n_38559 =  x_1362 & ~n_26318;
assign n_38560 =  i_8 &  n_26318;
assign n_38561 = ~n_38559 & ~n_38560;
assign n_38562 =  x_1362 & ~n_38561;
assign n_38563 = ~x_1362 &  n_38561;
assign n_38564 = ~n_38562 & ~n_38563;
assign n_38565 =  x_1361 & ~n_26318;
assign n_38566 =  i_7 &  n_26318;
assign n_38567 = ~n_38565 & ~n_38566;
assign n_38568 =  x_1361 & ~n_38567;
assign n_38569 = ~x_1361 &  n_38567;
assign n_38570 = ~n_38568 & ~n_38569;
assign n_38571 =  x_1360 & ~n_26318;
assign n_38572 =  i_6 &  n_26318;
assign n_38573 = ~n_38571 & ~n_38572;
assign n_38574 =  x_1360 & ~n_38573;
assign n_38575 = ~x_1360 &  n_38573;
assign n_38576 = ~n_38574 & ~n_38575;
assign n_38577 =  x_1359 & ~n_26318;
assign n_38578 =  i_5 &  n_26318;
assign n_38579 = ~n_38577 & ~n_38578;
assign n_38580 =  x_1359 & ~n_38579;
assign n_38581 = ~x_1359 &  n_38579;
assign n_38582 = ~n_38580 & ~n_38581;
assign n_38583 =  x_1358 & ~n_26318;
assign n_38584 =  i_4 &  n_26318;
assign n_38585 = ~n_38583 & ~n_38584;
assign n_38586 =  x_1358 & ~n_38585;
assign n_38587 = ~x_1358 &  n_38585;
assign n_38588 = ~n_38586 & ~n_38587;
assign n_38589 =  x_1357 & ~n_26318;
assign n_38590 =  i_3 &  n_26318;
assign n_38591 = ~n_38589 & ~n_38590;
assign n_38592 =  x_1357 & ~n_38591;
assign n_38593 = ~x_1357 &  n_38591;
assign n_38594 = ~n_38592 & ~n_38593;
assign n_38595 =  x_1356 & ~n_26318;
assign n_38596 =  i_2 &  n_26318;
assign n_38597 = ~n_38595 & ~n_38596;
assign n_38598 =  x_1356 & ~n_38597;
assign n_38599 = ~x_1356 &  n_38597;
assign n_38600 = ~n_38598 & ~n_38599;
assign n_38601 =  x_1355 & ~n_26318;
assign n_38602 =  i_1 &  n_26318;
assign n_38603 = ~n_38601 & ~n_38602;
assign n_38604 =  x_1355 & ~n_38603;
assign n_38605 = ~x_1355 &  n_38603;
assign n_38606 = ~n_38604 & ~n_38605;
assign n_38607 =  x_1354 & ~n_13231;
assign n_38608 =  i_32 &  n_13231;
assign n_38609 = ~n_38607 & ~n_38608;
assign n_38610 =  x_1354 & ~n_38609;
assign n_38611 = ~x_1354 &  n_38609;
assign n_38612 = ~n_38610 & ~n_38611;
assign n_38613 =  x_1353 & ~n_13231;
assign n_38614 =  i_31 &  n_13231;
assign n_38615 = ~n_38613 & ~n_38614;
assign n_38616 =  x_1353 & ~n_38615;
assign n_38617 = ~x_1353 &  n_38615;
assign n_38618 = ~n_38616 & ~n_38617;
assign n_38619 =  x_1352 & ~n_13231;
assign n_38620 =  i_30 &  n_13231;
assign n_38621 = ~n_38619 & ~n_38620;
assign n_38622 =  x_1352 & ~n_38621;
assign n_38623 = ~x_1352 &  n_38621;
assign n_38624 = ~n_38622 & ~n_38623;
assign n_38625 =  x_1351 & ~n_13231;
assign n_38626 =  i_29 &  n_13231;
assign n_38627 = ~n_38625 & ~n_38626;
assign n_38628 =  x_1351 & ~n_38627;
assign n_38629 = ~x_1351 &  n_38627;
assign n_38630 = ~n_38628 & ~n_38629;
assign n_38631 =  x_1350 & ~n_13231;
assign n_38632 =  i_28 &  n_13231;
assign n_38633 = ~n_38631 & ~n_38632;
assign n_38634 =  x_1350 & ~n_38633;
assign n_38635 = ~x_1350 &  n_38633;
assign n_38636 = ~n_38634 & ~n_38635;
assign n_38637 =  x_1349 & ~n_13231;
assign n_38638 =  i_27 &  n_13231;
assign n_38639 = ~n_38637 & ~n_38638;
assign n_38640 =  x_1349 & ~n_38639;
assign n_38641 = ~x_1349 &  n_38639;
assign n_38642 = ~n_38640 & ~n_38641;
assign n_38643 =  x_1348 & ~n_13231;
assign n_38644 =  i_26 &  n_13231;
assign n_38645 = ~n_38643 & ~n_38644;
assign n_38646 =  x_1348 & ~n_38645;
assign n_38647 = ~x_1348 &  n_38645;
assign n_38648 = ~n_38646 & ~n_38647;
assign n_38649 =  x_1347 & ~n_13231;
assign n_38650 =  i_25 &  n_13231;
assign n_38651 = ~n_38649 & ~n_38650;
assign n_38652 =  x_1347 & ~n_38651;
assign n_38653 = ~x_1347 &  n_38651;
assign n_38654 = ~n_38652 & ~n_38653;
assign n_38655 =  x_1346 & ~n_13231;
assign n_38656 =  i_24 &  n_13231;
assign n_38657 = ~n_38655 & ~n_38656;
assign n_38658 =  x_1346 & ~n_38657;
assign n_38659 = ~x_1346 &  n_38657;
assign n_38660 = ~n_38658 & ~n_38659;
assign n_38661 =  x_1345 & ~n_13231;
assign n_38662 =  i_23 &  n_13231;
assign n_38663 = ~n_38661 & ~n_38662;
assign n_38664 =  x_1345 & ~n_38663;
assign n_38665 = ~x_1345 &  n_38663;
assign n_38666 = ~n_38664 & ~n_38665;
assign n_38667 =  x_1344 & ~n_13231;
assign n_38668 =  i_22 &  n_13231;
assign n_38669 = ~n_38667 & ~n_38668;
assign n_38670 =  x_1344 & ~n_38669;
assign n_38671 = ~x_1344 &  n_38669;
assign n_38672 = ~n_38670 & ~n_38671;
assign n_38673 =  x_1343 & ~n_13231;
assign n_38674 =  i_21 &  n_13231;
assign n_38675 = ~n_38673 & ~n_38674;
assign n_38676 =  x_1343 & ~n_38675;
assign n_38677 = ~x_1343 &  n_38675;
assign n_38678 = ~n_38676 & ~n_38677;
assign n_38679 =  x_1342 & ~n_13231;
assign n_38680 =  i_20 &  n_13231;
assign n_38681 = ~n_38679 & ~n_38680;
assign n_38682 =  x_1342 & ~n_38681;
assign n_38683 = ~x_1342 &  n_38681;
assign n_38684 = ~n_38682 & ~n_38683;
assign n_38685 =  x_1341 & ~n_13231;
assign n_38686 =  i_19 &  n_13231;
assign n_38687 = ~n_38685 & ~n_38686;
assign n_38688 =  x_1341 & ~n_38687;
assign n_38689 = ~x_1341 &  n_38687;
assign n_38690 = ~n_38688 & ~n_38689;
assign n_38691 =  x_1340 & ~n_13231;
assign n_38692 =  i_18 &  n_13231;
assign n_38693 = ~n_38691 & ~n_38692;
assign n_38694 =  x_1340 & ~n_38693;
assign n_38695 = ~x_1340 &  n_38693;
assign n_38696 = ~n_38694 & ~n_38695;
assign n_38697 =  x_1339 & ~n_13231;
assign n_38698 =  i_17 &  n_13231;
assign n_38699 = ~n_38697 & ~n_38698;
assign n_38700 =  x_1339 & ~n_38699;
assign n_38701 = ~x_1339 &  n_38699;
assign n_38702 = ~n_38700 & ~n_38701;
assign n_38703 =  x_1338 & ~n_13231;
assign n_38704 =  i_16 &  n_13231;
assign n_38705 = ~n_38703 & ~n_38704;
assign n_38706 =  x_1338 & ~n_38705;
assign n_38707 = ~x_1338 &  n_38705;
assign n_38708 = ~n_38706 & ~n_38707;
assign n_38709 =  x_1337 & ~n_13231;
assign n_38710 =  i_15 &  n_13231;
assign n_38711 = ~n_38709 & ~n_38710;
assign n_38712 =  x_1337 & ~n_38711;
assign n_38713 = ~x_1337 &  n_38711;
assign n_38714 = ~n_38712 & ~n_38713;
assign n_38715 =  x_1336 & ~n_13231;
assign n_38716 =  i_14 &  n_13231;
assign n_38717 = ~n_38715 & ~n_38716;
assign n_38718 =  x_1336 & ~n_38717;
assign n_38719 = ~x_1336 &  n_38717;
assign n_38720 = ~n_38718 & ~n_38719;
assign n_38721 =  x_1335 & ~n_13231;
assign n_38722 =  i_13 &  n_13231;
assign n_38723 = ~n_38721 & ~n_38722;
assign n_38724 =  x_1335 & ~n_38723;
assign n_38725 = ~x_1335 &  n_38723;
assign n_38726 = ~n_38724 & ~n_38725;
assign n_38727 =  x_1334 & ~n_13231;
assign n_38728 =  i_12 &  n_13231;
assign n_38729 = ~n_38727 & ~n_38728;
assign n_38730 =  x_1334 & ~n_38729;
assign n_38731 = ~x_1334 &  n_38729;
assign n_38732 = ~n_38730 & ~n_38731;
assign n_38733 =  x_1333 & ~n_13231;
assign n_38734 =  i_11 &  n_13231;
assign n_38735 = ~n_38733 & ~n_38734;
assign n_38736 =  x_1333 & ~n_38735;
assign n_38737 = ~x_1333 &  n_38735;
assign n_38738 = ~n_38736 & ~n_38737;
assign n_38739 =  x_1332 & ~n_13231;
assign n_38740 =  i_10 &  n_13231;
assign n_38741 = ~n_38739 & ~n_38740;
assign n_38742 =  x_1332 & ~n_38741;
assign n_38743 = ~x_1332 &  n_38741;
assign n_38744 = ~n_38742 & ~n_38743;
assign n_38745 =  x_4208 & ~n_6380;
assign n_38746 =  i_8 &  n_6380;
assign n_38747 = ~n_38745 & ~n_38746;
assign n_38748 =  x_4208 & ~n_38747;
assign n_38749 = ~x_4208 &  n_38747;
assign n_38750 = ~n_38748 & ~n_38749;
assign n_38751 =  x_4207 & ~n_6380;
assign n_38752 =  i_7 &  n_6380;
assign n_38753 = ~n_38751 & ~n_38752;
assign n_38754 =  x_4207 & ~n_38753;
assign n_38755 = ~x_4207 &  n_38753;
assign n_38756 = ~n_38754 & ~n_38755;
assign n_38757 =  x_4206 & ~n_6380;
assign n_38758 =  i_6 &  n_6380;
assign n_38759 = ~n_38757 & ~n_38758;
assign n_38760 =  x_4206 & ~n_38759;
assign n_38761 = ~x_4206 &  n_38759;
assign n_38762 = ~n_38760 & ~n_38761;
assign n_38763 =  x_4205 & ~n_6380;
assign n_38764 =  i_5 &  n_6380;
assign n_38765 = ~n_38763 & ~n_38764;
assign n_38766 =  x_4205 & ~n_38765;
assign n_38767 = ~x_4205 &  n_38765;
assign n_38768 = ~n_38766 & ~n_38767;
assign n_38769 =  x_4204 & ~n_6380;
assign n_38770 =  i_4 &  n_6380;
assign n_38771 = ~n_38769 & ~n_38770;
assign n_38772 =  x_4204 & ~n_38771;
assign n_38773 = ~x_4204 &  n_38771;
assign n_38774 = ~n_38772 & ~n_38773;
assign n_38775 =  x_4203 & ~n_6380;
assign n_38776 =  i_3 &  n_6380;
assign n_38777 = ~n_38775 & ~n_38776;
assign n_38778 =  x_4203 & ~n_38777;
assign n_38779 = ~x_4203 &  n_38777;
assign n_38780 = ~n_38778 & ~n_38779;
assign n_38781 =  x_4202 & ~n_6380;
assign n_38782 =  i_2 &  n_6380;
assign n_38783 = ~n_38781 & ~n_38782;
assign n_38784 =  x_4202 & ~n_38783;
assign n_38785 = ~x_4202 &  n_38783;
assign n_38786 = ~n_38784 & ~n_38785;
assign n_38787 =  x_4201 & ~n_6380;
assign n_38788 =  i_1 &  n_6380;
assign n_38789 = ~n_38787 & ~n_38788;
assign n_38790 =  x_4201 & ~n_38789;
assign n_38791 = ~x_4201 &  n_38789;
assign n_38792 = ~n_38790 & ~n_38791;
assign n_38793 =  x_4200 & ~n_25232;
assign n_38794 =  x_4200 &  n_38793;
assign n_38795 = ~x_4200 & ~n_38793;
assign n_38796 = ~n_38794 & ~n_38795;
assign n_38797 =  x_4199 & ~n_25232;
assign n_38798 =  x_4199 &  n_38797;
assign n_38799 = ~x_4199 & ~n_38797;
assign n_38800 = ~n_38798 & ~n_38799;
assign n_38801 =  x_4198 & ~n_25232;
assign n_38802 =  x_4198 &  n_38801;
assign n_38803 = ~x_4198 & ~n_38801;
assign n_38804 = ~n_38802 & ~n_38803;
assign n_38805 =  x_4197 & ~n_25232;
assign n_38806 =  x_4197 &  n_38805;
assign n_38807 = ~x_4197 & ~n_38805;
assign n_38808 = ~n_38806 & ~n_38807;
assign n_38809 =  x_4196 & ~n_25232;
assign n_38810 =  x_4196 &  n_38809;
assign n_38811 = ~x_4196 & ~n_38809;
assign n_38812 = ~n_38810 & ~n_38811;
assign n_38813 =  x_4195 & ~n_25232;
assign n_38814 =  x_4195 &  n_38813;
assign n_38815 = ~x_4195 & ~n_38813;
assign n_38816 = ~n_38814 & ~n_38815;
assign n_38817 =  x_4194 & ~n_25232;
assign n_38818 =  x_4194 &  n_38817;
assign n_38819 = ~x_4194 & ~n_38817;
assign n_38820 = ~n_38818 & ~n_38819;
assign n_38821 =  x_4193 & ~n_25232;
assign n_38822 =  x_4193 &  n_38821;
assign n_38823 = ~x_4193 & ~n_38821;
assign n_38824 = ~n_38822 & ~n_38823;
assign n_38825 =  x_4192 & ~n_25232;
assign n_38826 =  x_4192 &  n_38825;
assign n_38827 = ~x_4192 & ~n_38825;
assign n_38828 = ~n_38826 & ~n_38827;
assign n_38829 =  x_4191 & ~n_25232;
assign n_38830 =  x_4191 &  n_38829;
assign n_38831 = ~x_4191 & ~n_38829;
assign n_38832 = ~n_38830 & ~n_38831;
assign n_38833 =  x_4190 & ~n_25232;
assign n_38834 =  x_4190 &  n_38833;
assign n_38835 = ~x_4190 & ~n_38833;
assign n_38836 = ~n_38834 & ~n_38835;
assign n_38837 =  x_4189 & ~n_25232;
assign n_38838 =  x_4189 &  n_38837;
assign n_38839 = ~x_4189 & ~n_38837;
assign n_38840 = ~n_38838 & ~n_38839;
assign n_38841 =  x_4188 & ~n_25232;
assign n_38842 =  x_4188 &  n_38841;
assign n_38843 = ~x_4188 & ~n_38841;
assign n_38844 = ~n_38842 & ~n_38843;
assign n_38845 =  x_4187 & ~n_25232;
assign n_38846 =  x_4187 &  n_38845;
assign n_38847 = ~x_4187 & ~n_38845;
assign n_38848 = ~n_38846 & ~n_38847;
assign n_38849 =  x_4186 & ~n_25232;
assign n_38850 =  x_4186 &  n_38849;
assign n_38851 = ~x_4186 & ~n_38849;
assign n_38852 = ~n_38850 & ~n_38851;
assign n_38853 =  x_4185 & ~n_25232;
assign n_38854 =  x_4185 &  n_38853;
assign n_38855 = ~x_4185 & ~n_38853;
assign n_38856 = ~n_38854 & ~n_38855;
assign n_38857 =  x_4184 & ~n_25232;
assign n_38858 =  x_4184 &  n_38857;
assign n_38859 = ~x_4184 & ~n_38857;
assign n_38860 = ~n_38858 & ~n_38859;
assign n_38861 =  x_4183 & ~n_25232;
assign n_38862 =  x_4183 &  n_38861;
assign n_38863 = ~x_4183 & ~n_38861;
assign n_38864 = ~n_38862 & ~n_38863;
assign n_38865 =  x_4182 & ~n_25232;
assign n_38866 =  x_4182 &  n_38865;
assign n_38867 = ~x_4182 & ~n_38865;
assign n_38868 = ~n_38866 & ~n_38867;
assign n_38869 =  x_4181 & ~n_25232;
assign n_38870 =  x_4181 &  n_38869;
assign n_38871 = ~x_4181 & ~n_38869;
assign n_38872 = ~n_38870 & ~n_38871;
assign n_38873 =  x_4180 & ~n_25232;
assign n_38874 =  x_4180 &  n_38873;
assign n_38875 = ~x_4180 & ~n_38873;
assign n_38876 = ~n_38874 & ~n_38875;
assign n_38877 =  x_4179 & ~n_25232;
assign n_38878 =  x_4179 &  n_38877;
assign n_38879 = ~x_4179 & ~n_38877;
assign n_38880 = ~n_38878 & ~n_38879;
assign n_38881 =  x_4178 & ~n_25232;
assign n_38882 =  x_4178 &  n_38881;
assign n_38883 = ~x_4178 & ~n_38881;
assign n_38884 = ~n_38882 & ~n_38883;
assign n_38885 =  x_4177 & ~n_25232;
assign n_38886 =  x_4177 &  n_38885;
assign n_38887 = ~x_4177 & ~n_38885;
assign n_38888 = ~n_38886 & ~n_38887;
assign n_38889 =  x_4176 & ~n_25232;
assign n_38890 =  x_4176 &  n_38889;
assign n_38891 = ~x_4176 & ~n_38889;
assign n_38892 = ~n_38890 & ~n_38891;
assign n_38893 =  x_4175 & ~n_25232;
assign n_38894 =  x_4175 &  n_38893;
assign n_38895 = ~x_4175 & ~n_38893;
assign n_38896 = ~n_38894 & ~n_38895;
assign n_38897 =  x_4174 & ~n_25232;
assign n_38898 =  x_4174 &  n_38897;
assign n_38899 = ~x_4174 & ~n_38897;
assign n_38900 = ~n_38898 & ~n_38899;
assign n_38901 =  x_4173 & ~n_25232;
assign n_38902 =  x_4173 &  n_38901;
assign n_38903 = ~x_4173 & ~n_38901;
assign n_38904 = ~n_38902 & ~n_38903;
assign n_38905 =  x_4172 & ~n_25232;
assign n_38906 =  x_4172 &  n_38905;
assign n_38907 = ~x_4172 & ~n_38905;
assign n_38908 = ~n_38906 & ~n_38907;
assign n_38909 =  x_4171 & ~n_25232;
assign n_38910 =  x_4171 &  n_38909;
assign n_38911 = ~x_4171 & ~n_38909;
assign n_38912 = ~n_38910 & ~n_38911;
assign n_38913 =  x_4170 & ~n_25232;
assign n_38914 =  x_4170 &  n_38913;
assign n_38915 = ~x_4170 & ~n_38913;
assign n_38916 = ~n_38914 & ~n_38915;
assign n_38917 =  x_4169 & ~n_25232;
assign n_38918 =  x_4169 &  n_38917;
assign n_38919 = ~x_4169 & ~n_38917;
assign n_38920 = ~n_38918 & ~n_38919;
assign n_38921 =  x_4008 &  n_23768;
assign n_38922 =  n_23379 &  n_26416;
assign n_38923 =  x_4168 &  n_38922;
assign n_38924 = ~n_38921 & ~n_38923;
assign n_38925 =  x_4168 & ~n_38924;
assign n_38926 = ~x_4168 &  n_38924;
assign n_38927 = ~n_38925 & ~n_38926;
assign n_38928 =  x_4007 &  n_23768;
assign n_38929 =  x_4167 &  n_38922;
assign n_38930 = ~n_38928 & ~n_38929;
assign n_38931 =  x_4167 & ~n_38930;
assign n_38932 = ~x_4167 &  n_38930;
assign n_38933 = ~n_38931 & ~n_38932;
assign n_38934 =  x_4006 &  n_23768;
assign n_38935 =  x_4166 &  n_38922;
assign n_38936 = ~n_38934 & ~n_38935;
assign n_38937 =  x_4166 & ~n_38936;
assign n_38938 = ~x_4166 &  n_38936;
assign n_38939 = ~n_38937 & ~n_38938;
assign n_38940 =  x_4005 &  n_23768;
assign n_38941 =  x_4165 &  n_38922;
assign n_38942 = ~n_38940 & ~n_38941;
assign n_38943 =  x_4165 & ~n_38942;
assign n_38944 = ~x_4165 &  n_38942;
assign n_38945 = ~n_38943 & ~n_38944;
assign n_38946 =  x_4004 &  n_23768;
assign n_38947 =  x_4164 &  n_38922;
assign n_38948 = ~n_38946 & ~n_38947;
assign n_38949 =  x_4164 & ~n_38948;
assign n_38950 = ~x_4164 &  n_38948;
assign n_38951 = ~n_38949 & ~n_38950;
assign n_38952 =  x_4003 &  n_23768;
assign n_38953 =  x_4163 &  n_38922;
assign n_38954 = ~n_38952 & ~n_38953;
assign n_38955 =  x_4163 & ~n_38954;
assign n_38956 = ~x_4163 &  n_38954;
assign n_38957 = ~n_38955 & ~n_38956;
assign n_38958 =  x_4002 &  n_23768;
assign n_38959 =  x_4162 &  n_38922;
assign n_38960 = ~n_38958 & ~n_38959;
assign n_38961 =  x_4162 & ~n_38960;
assign n_38962 = ~x_4162 &  n_38960;
assign n_38963 = ~n_38961 & ~n_38962;
assign n_38964 =  x_4001 &  n_23768;
assign n_38965 =  x_4161 &  n_38922;
assign n_38966 = ~n_38964 & ~n_38965;
assign n_38967 =  x_4161 & ~n_38966;
assign n_38968 = ~x_4161 &  n_38966;
assign n_38969 = ~n_38967 & ~n_38968;
assign n_38970 =  x_4000 &  n_23768;
assign n_38971 =  x_4160 &  n_38922;
assign n_38972 = ~n_38970 & ~n_38971;
assign n_38973 =  x_4160 & ~n_38972;
assign n_38974 = ~x_4160 &  n_38972;
assign n_38975 = ~n_38973 & ~n_38974;
assign n_38976 =  x_3999 &  n_23768;
assign n_38977 =  x_4159 &  n_38922;
assign n_38978 = ~n_38976 & ~n_38977;
assign n_38979 =  x_4159 & ~n_38978;
assign n_38980 = ~x_4159 &  n_38978;
assign n_38981 = ~n_38979 & ~n_38980;
assign n_38982 =  x_3998 &  n_23768;
assign n_38983 =  x_4158 &  n_38922;
assign n_38984 = ~n_38982 & ~n_38983;
assign n_38985 =  x_4158 & ~n_38984;
assign n_38986 = ~x_4158 &  n_38984;
assign n_38987 = ~n_38985 & ~n_38986;
assign n_38988 =  x_3997 &  n_23768;
assign n_38989 =  x_4157 &  n_38922;
assign n_38990 = ~n_38988 & ~n_38989;
assign n_38991 =  x_4157 & ~n_38990;
assign n_38992 = ~x_4157 &  n_38990;
assign n_38993 = ~n_38991 & ~n_38992;
assign n_38994 =  x_3996 &  n_23768;
assign n_38995 =  x_4156 &  n_38922;
assign n_38996 = ~n_38994 & ~n_38995;
assign n_38997 =  x_4156 & ~n_38996;
assign n_38998 = ~x_4156 &  n_38996;
assign n_38999 = ~n_38997 & ~n_38998;
assign n_39000 =  x_3995 &  n_23768;
assign n_39001 =  x_4155 &  n_38922;
assign n_39002 = ~n_39000 & ~n_39001;
assign n_39003 =  x_4155 & ~n_39002;
assign n_39004 = ~x_4155 &  n_39002;
assign n_39005 = ~n_39003 & ~n_39004;
assign n_39006 =  x_3994 &  n_23768;
assign n_39007 =  x_4154 &  n_38922;
assign n_39008 = ~n_39006 & ~n_39007;
assign n_39009 =  x_4154 & ~n_39008;
assign n_39010 = ~x_4154 &  n_39008;
assign n_39011 = ~n_39009 & ~n_39010;
assign n_39012 =  x_3993 &  n_23768;
assign n_39013 =  x_4153 &  n_38922;
assign n_39014 = ~n_39012 & ~n_39013;
assign n_39015 =  x_4153 & ~n_39014;
assign n_39016 = ~x_4153 &  n_39014;
assign n_39017 = ~n_39015 & ~n_39016;
assign n_39018 =  x_3992 &  n_23768;
assign n_39019 =  x_4152 &  n_38922;
assign n_39020 = ~n_39018 & ~n_39019;
assign n_39021 =  x_4152 & ~n_39020;
assign n_39022 = ~x_4152 &  n_39020;
assign n_39023 = ~n_39021 & ~n_39022;
assign n_39024 =  x_3991 &  n_23768;
assign n_39025 =  x_4151 &  n_38922;
assign n_39026 = ~n_39024 & ~n_39025;
assign n_39027 =  x_4151 & ~n_39026;
assign n_39028 = ~x_4151 &  n_39026;
assign n_39029 = ~n_39027 & ~n_39028;
assign n_39030 =  x_3990 &  n_23768;
assign n_39031 =  x_4150 &  n_38922;
assign n_39032 = ~n_39030 & ~n_39031;
assign n_39033 =  x_4150 & ~n_39032;
assign n_39034 = ~x_4150 &  n_39032;
assign n_39035 = ~n_39033 & ~n_39034;
assign n_39036 =  x_3989 &  n_23768;
assign n_39037 =  x_4149 &  n_38922;
assign n_39038 = ~n_39036 & ~n_39037;
assign n_39039 =  x_4149 & ~n_39038;
assign n_39040 = ~x_4149 &  n_39038;
assign n_39041 = ~n_39039 & ~n_39040;
assign n_39042 =  x_3988 &  n_23768;
assign n_39043 =  x_4148 &  n_38922;
assign n_39044 = ~n_39042 & ~n_39043;
assign n_39045 =  x_4148 & ~n_39044;
assign n_39046 = ~x_4148 &  n_39044;
assign n_39047 = ~n_39045 & ~n_39046;
assign n_39048 =  x_3987 &  n_23768;
assign n_39049 =  x_4147 &  n_38922;
assign n_39050 = ~n_39048 & ~n_39049;
assign n_39051 =  x_4147 & ~n_39050;
assign n_39052 = ~x_4147 &  n_39050;
assign n_39053 = ~n_39051 & ~n_39052;
assign n_39054 =  x_3986 &  n_23768;
assign n_39055 =  x_4146 &  n_38922;
assign n_39056 = ~n_39054 & ~n_39055;
assign n_39057 =  x_4146 & ~n_39056;
assign n_39058 = ~x_4146 &  n_39056;
assign n_39059 = ~n_39057 & ~n_39058;
assign n_39060 =  x_3985 &  n_23768;
assign n_39061 =  x_4145 &  n_38922;
assign n_39062 = ~n_39060 & ~n_39061;
assign n_39063 =  x_4145 & ~n_39062;
assign n_39064 = ~x_4145 &  n_39062;
assign n_39065 = ~n_39063 & ~n_39064;
assign n_39066 =  x_3984 &  n_23768;
assign n_39067 =  x_4144 &  n_38922;
assign n_39068 = ~n_39066 & ~n_39067;
assign n_39069 =  x_4144 & ~n_39068;
assign n_39070 = ~x_4144 &  n_39068;
assign n_39071 = ~n_39069 & ~n_39070;
assign n_39072 =  x_3983 &  n_23768;
assign n_39073 =  x_4143 &  n_38922;
assign n_39074 = ~n_39072 & ~n_39073;
assign n_39075 =  x_4143 & ~n_39074;
assign n_39076 = ~x_4143 &  n_39074;
assign n_39077 = ~n_39075 & ~n_39076;
assign n_39078 =  x_3982 &  n_23768;
assign n_39079 =  x_4142 &  n_38922;
assign n_39080 = ~n_39078 & ~n_39079;
assign n_39081 =  x_4142 & ~n_39080;
assign n_39082 = ~x_4142 &  n_39080;
assign n_39083 = ~n_39081 & ~n_39082;
assign n_39084 =  x_3981 &  n_23768;
assign n_39085 =  x_4141 &  n_38922;
assign n_39086 = ~n_39084 & ~n_39085;
assign n_39087 =  x_4141 & ~n_39086;
assign n_39088 = ~x_4141 &  n_39086;
assign n_39089 = ~n_39087 & ~n_39088;
assign n_39090 =  x_3980 &  n_23768;
assign n_39091 =  x_4140 &  n_38922;
assign n_39092 = ~n_39090 & ~n_39091;
assign n_39093 =  x_4140 & ~n_39092;
assign n_39094 = ~x_4140 &  n_39092;
assign n_39095 = ~n_39093 & ~n_39094;
assign n_39096 =  x_3979 &  n_23768;
assign n_39097 =  x_4139 &  n_38922;
assign n_39098 = ~n_39096 & ~n_39097;
assign n_39099 =  x_4139 & ~n_39098;
assign n_39100 = ~x_4139 &  n_39098;
assign n_39101 = ~n_39099 & ~n_39100;
assign n_39102 =  x_3978 &  n_23768;
assign n_39103 =  x_4138 &  n_38922;
assign n_39104 = ~n_39102 & ~n_39103;
assign n_39105 =  x_4138 & ~n_39104;
assign n_39106 = ~x_4138 &  n_39104;
assign n_39107 = ~n_39105 & ~n_39106;
assign n_39108 =  x_3977 &  n_23768;
assign n_39109 =  x_4137 &  n_38922;
assign n_39110 = ~n_39108 & ~n_39109;
assign n_39111 =  x_4137 & ~n_39110;
assign n_39112 = ~x_4137 &  n_39110;
assign n_39113 = ~n_39111 & ~n_39112;
assign n_39114 =  x_4136 & ~n_26023;
assign n_39115 =  i_32 &  n_26023;
assign n_39116 = ~n_39114 & ~n_39115;
assign n_39117 =  x_4136 & ~n_39116;
assign n_39118 = ~x_4136 &  n_39116;
assign n_39119 = ~n_39117 & ~n_39118;
assign n_39120 =  x_4135 & ~n_26023;
assign n_39121 =  i_31 &  n_26023;
assign n_39122 = ~n_39120 & ~n_39121;
assign n_39123 =  x_4135 & ~n_39122;
assign n_39124 = ~x_4135 &  n_39122;
assign n_39125 = ~n_39123 & ~n_39124;
assign n_39126 =  x_4134 & ~n_26023;
assign n_39127 =  i_30 &  n_26023;
assign n_39128 = ~n_39126 & ~n_39127;
assign n_39129 =  x_4134 & ~n_39128;
assign n_39130 = ~x_4134 &  n_39128;
assign n_39131 = ~n_39129 & ~n_39130;
assign n_39132 =  x_4133 & ~n_26023;
assign n_39133 =  i_29 &  n_26023;
assign n_39134 = ~n_39132 & ~n_39133;
assign n_39135 =  x_4133 & ~n_39134;
assign n_39136 = ~x_4133 &  n_39134;
assign n_39137 = ~n_39135 & ~n_39136;
assign n_39138 =  x_4132 & ~n_26023;
assign n_39139 =  i_28 &  n_26023;
assign n_39140 = ~n_39138 & ~n_39139;
assign n_39141 =  x_4132 & ~n_39140;
assign n_39142 = ~x_4132 &  n_39140;
assign n_39143 = ~n_39141 & ~n_39142;
assign n_39144 =  x_4131 & ~n_26023;
assign n_39145 =  i_27 &  n_26023;
assign n_39146 = ~n_39144 & ~n_39145;
assign n_39147 =  x_4131 & ~n_39146;
assign n_39148 = ~x_4131 &  n_39146;
assign n_39149 = ~n_39147 & ~n_39148;
assign n_39150 =  x_4130 & ~n_26023;
assign n_39151 =  i_26 &  n_26023;
assign n_39152 = ~n_39150 & ~n_39151;
assign n_39153 =  x_4130 & ~n_39152;
assign n_39154 = ~x_4130 &  n_39152;
assign n_39155 = ~n_39153 & ~n_39154;
assign n_39156 =  x_4129 & ~n_26023;
assign n_39157 =  i_25 &  n_26023;
assign n_39158 = ~n_39156 & ~n_39157;
assign n_39159 =  x_4129 & ~n_39158;
assign n_39160 = ~x_4129 &  n_39158;
assign n_39161 = ~n_39159 & ~n_39160;
assign n_39162 =  x_4128 & ~n_26023;
assign n_39163 =  i_24 &  n_26023;
assign n_39164 = ~n_39162 & ~n_39163;
assign n_39165 =  x_4128 & ~n_39164;
assign n_39166 = ~x_4128 &  n_39164;
assign n_39167 = ~n_39165 & ~n_39166;
assign n_39168 =  x_4127 & ~n_26023;
assign n_39169 =  i_23 &  n_26023;
assign n_39170 = ~n_39168 & ~n_39169;
assign n_39171 =  x_4127 & ~n_39170;
assign n_39172 = ~x_4127 &  n_39170;
assign n_39173 = ~n_39171 & ~n_39172;
assign n_39174 =  x_4126 & ~n_26023;
assign n_39175 =  i_22 &  n_26023;
assign n_39176 = ~n_39174 & ~n_39175;
assign n_39177 =  x_4126 & ~n_39176;
assign n_39178 = ~x_4126 &  n_39176;
assign n_39179 = ~n_39177 & ~n_39178;
assign n_39180 =  x_4125 & ~n_26023;
assign n_39181 =  i_21 &  n_26023;
assign n_39182 = ~n_39180 & ~n_39181;
assign n_39183 =  x_4125 & ~n_39182;
assign n_39184 = ~x_4125 &  n_39182;
assign n_39185 = ~n_39183 & ~n_39184;
assign n_39186 =  x_4124 & ~n_26023;
assign n_39187 =  i_20 &  n_26023;
assign n_39188 = ~n_39186 & ~n_39187;
assign n_39189 =  x_4124 & ~n_39188;
assign n_39190 = ~x_4124 &  n_39188;
assign n_39191 = ~n_39189 & ~n_39190;
assign n_39192 =  x_4123 & ~n_26023;
assign n_39193 =  i_19 &  n_26023;
assign n_39194 = ~n_39192 & ~n_39193;
assign n_39195 =  x_4123 & ~n_39194;
assign n_39196 = ~x_4123 &  n_39194;
assign n_39197 = ~n_39195 & ~n_39196;
assign n_39198 =  x_4122 & ~n_26023;
assign n_39199 =  i_18 &  n_26023;
assign n_39200 = ~n_39198 & ~n_39199;
assign n_39201 =  x_4122 & ~n_39200;
assign n_39202 = ~x_4122 &  n_39200;
assign n_39203 = ~n_39201 & ~n_39202;
assign n_39204 =  x_4121 & ~n_26023;
assign n_39205 =  i_17 &  n_26023;
assign n_39206 = ~n_39204 & ~n_39205;
assign n_39207 =  x_4121 & ~n_39206;
assign n_39208 = ~x_4121 &  n_39206;
assign n_39209 = ~n_39207 & ~n_39208;
assign n_39210 =  x_4120 & ~n_26023;
assign n_39211 =  i_16 &  n_26023;
assign n_39212 = ~n_39210 & ~n_39211;
assign n_39213 =  x_4120 & ~n_39212;
assign n_39214 = ~x_4120 &  n_39212;
assign n_39215 = ~n_39213 & ~n_39214;
assign n_39216 =  x_4119 & ~n_26023;
assign n_39217 =  i_15 &  n_26023;
assign n_39218 = ~n_39216 & ~n_39217;
assign n_39219 =  x_4119 & ~n_39218;
assign n_39220 = ~x_4119 &  n_39218;
assign n_39221 = ~n_39219 & ~n_39220;
assign n_39222 =  x_4118 & ~n_26023;
assign n_39223 =  i_14 &  n_26023;
assign n_39224 = ~n_39222 & ~n_39223;
assign n_39225 =  x_4118 & ~n_39224;
assign n_39226 = ~x_4118 &  n_39224;
assign n_39227 = ~n_39225 & ~n_39226;
assign n_39228 =  x_4117 & ~n_26023;
assign n_39229 =  i_13 &  n_26023;
assign n_39230 = ~n_39228 & ~n_39229;
assign n_39231 =  x_4117 & ~n_39230;
assign n_39232 = ~x_4117 &  n_39230;
assign n_39233 = ~n_39231 & ~n_39232;
assign n_39234 =  x_4116 & ~n_26023;
assign n_39235 =  i_12 &  n_26023;
assign n_39236 = ~n_39234 & ~n_39235;
assign n_39237 =  x_4116 & ~n_39236;
assign n_39238 = ~x_4116 &  n_39236;
assign n_39239 = ~n_39237 & ~n_39238;
assign n_39240 =  x_4115 & ~n_26023;
assign n_39241 =  i_11 &  n_26023;
assign n_39242 = ~n_39240 & ~n_39241;
assign n_39243 =  x_4115 & ~n_39242;
assign n_39244 = ~x_4115 &  n_39242;
assign n_39245 = ~n_39243 & ~n_39244;
assign n_39246 =  x_4114 & ~n_26023;
assign n_39247 =  i_10 &  n_26023;
assign n_39248 = ~n_39246 & ~n_39247;
assign n_39249 =  x_4114 & ~n_39248;
assign n_39250 = ~x_4114 &  n_39248;
assign n_39251 = ~n_39249 & ~n_39250;
assign n_39252 =  x_4113 & ~n_26023;
assign n_39253 =  i_9 &  n_26023;
assign n_39254 = ~n_39252 & ~n_39253;
assign n_39255 =  x_4113 & ~n_39254;
assign n_39256 = ~x_4113 &  n_39254;
assign n_39257 = ~n_39255 & ~n_39256;
assign n_39258 =  x_4112 & ~n_26023;
assign n_39259 =  i_8 &  n_26023;
assign n_39260 = ~n_39258 & ~n_39259;
assign n_39261 =  x_4112 & ~n_39260;
assign n_39262 = ~x_4112 &  n_39260;
assign n_39263 = ~n_39261 & ~n_39262;
assign n_39264 =  x_4111 & ~n_26023;
assign n_39265 =  i_7 &  n_26023;
assign n_39266 = ~n_39264 & ~n_39265;
assign n_39267 =  x_4111 & ~n_39266;
assign n_39268 = ~x_4111 &  n_39266;
assign n_39269 = ~n_39267 & ~n_39268;
assign n_39270 =  x_4110 & ~n_26023;
assign n_39271 =  i_6 &  n_26023;
assign n_39272 = ~n_39270 & ~n_39271;
assign n_39273 =  x_4110 & ~n_39272;
assign n_39274 = ~x_4110 &  n_39272;
assign n_39275 = ~n_39273 & ~n_39274;
assign n_39276 =  x_4109 & ~n_26023;
assign n_39277 =  i_5 &  n_26023;
assign n_39278 = ~n_39276 & ~n_39277;
assign n_39279 =  x_4109 & ~n_39278;
assign n_39280 = ~x_4109 &  n_39278;
assign n_39281 = ~n_39279 & ~n_39280;
assign n_39282 =  x_4108 & ~n_26023;
assign n_39283 =  i_4 &  n_26023;
assign n_39284 = ~n_39282 & ~n_39283;
assign n_39285 =  x_4108 & ~n_39284;
assign n_39286 = ~x_4108 &  n_39284;
assign n_39287 = ~n_39285 & ~n_39286;
assign n_39288 =  x_4107 & ~n_26023;
assign n_39289 =  i_3 &  n_26023;
assign n_39290 = ~n_39288 & ~n_39289;
assign n_39291 =  x_4107 & ~n_39290;
assign n_39292 = ~x_4107 &  n_39290;
assign n_39293 = ~n_39291 & ~n_39292;
assign n_39294 =  x_4106 & ~n_26023;
assign n_39295 =  i_2 &  n_26023;
assign n_39296 = ~n_39294 & ~n_39295;
assign n_39297 =  x_4106 & ~n_39296;
assign n_39298 = ~x_4106 &  n_39296;
assign n_39299 = ~n_39297 & ~n_39298;
assign n_39300 =  x_4105 & ~n_26023;
assign n_39301 =  i_1 &  n_26023;
assign n_39302 = ~n_39300 & ~n_39301;
assign n_39303 =  x_4105 & ~n_39302;
assign n_39304 = ~x_4105 &  n_39302;
assign n_39305 = ~n_39303 & ~n_39304;
assign n_39306 =  x_4104 & ~n_28855;
assign n_39307 =  i_32 &  n_28855;
assign n_39308 = ~n_39306 & ~n_39307;
assign n_39309 =  x_4104 & ~n_39308;
assign n_39310 = ~x_4104 &  n_39308;
assign n_39311 = ~n_39309 & ~n_39310;
assign n_39312 =  x_4103 & ~n_28855;
assign n_39313 =  i_31 &  n_28855;
assign n_39314 = ~n_39312 & ~n_39313;
assign n_39315 =  x_4103 & ~n_39314;
assign n_39316 = ~x_4103 &  n_39314;
assign n_39317 = ~n_39315 & ~n_39316;
assign n_39318 =  x_4102 & ~n_28855;
assign n_39319 =  i_30 &  n_28855;
assign n_39320 = ~n_39318 & ~n_39319;
assign n_39321 =  x_4102 & ~n_39320;
assign n_39322 = ~x_4102 &  n_39320;
assign n_39323 = ~n_39321 & ~n_39322;
assign n_39324 =  x_4101 & ~n_28855;
assign n_39325 =  i_29 &  n_28855;
assign n_39326 = ~n_39324 & ~n_39325;
assign n_39327 =  x_4101 & ~n_39326;
assign n_39328 = ~x_4101 &  n_39326;
assign n_39329 = ~n_39327 & ~n_39328;
assign n_39330 =  x_4100 & ~n_28855;
assign n_39331 =  i_28 &  n_28855;
assign n_39332 = ~n_39330 & ~n_39331;
assign n_39333 =  x_4100 & ~n_39332;
assign n_39334 = ~x_4100 &  n_39332;
assign n_39335 = ~n_39333 & ~n_39334;
assign n_39336 =  x_4099 & ~n_28855;
assign n_39337 =  i_27 &  n_28855;
assign n_39338 = ~n_39336 & ~n_39337;
assign n_39339 =  x_4099 & ~n_39338;
assign n_39340 = ~x_4099 &  n_39338;
assign n_39341 = ~n_39339 & ~n_39340;
assign n_39342 =  x_4098 & ~n_28855;
assign n_39343 =  i_26 &  n_28855;
assign n_39344 = ~n_39342 & ~n_39343;
assign n_39345 =  x_4098 & ~n_39344;
assign n_39346 = ~x_4098 &  n_39344;
assign n_39347 = ~n_39345 & ~n_39346;
assign n_39348 =  x_4097 & ~n_28855;
assign n_39349 =  i_25 &  n_28855;
assign n_39350 = ~n_39348 & ~n_39349;
assign n_39351 =  x_4097 & ~n_39350;
assign n_39352 = ~x_4097 &  n_39350;
assign n_39353 = ~n_39351 & ~n_39352;
assign n_39354 =  x_4096 & ~n_28855;
assign n_39355 =  i_24 &  n_28855;
assign n_39356 = ~n_39354 & ~n_39355;
assign n_39357 =  x_4096 & ~n_39356;
assign n_39358 = ~x_4096 &  n_39356;
assign n_39359 = ~n_39357 & ~n_39358;
assign n_39360 =  x_4095 & ~n_28855;
assign n_39361 =  i_23 &  n_28855;
assign n_39362 = ~n_39360 & ~n_39361;
assign n_39363 =  x_4095 & ~n_39362;
assign n_39364 = ~x_4095 &  n_39362;
assign n_39365 = ~n_39363 & ~n_39364;
assign n_39366 =  x_4094 & ~n_28855;
assign n_39367 =  i_22 &  n_28855;
assign n_39368 = ~n_39366 & ~n_39367;
assign n_39369 =  x_4094 & ~n_39368;
assign n_39370 = ~x_4094 &  n_39368;
assign n_39371 = ~n_39369 & ~n_39370;
assign n_39372 =  x_4093 & ~n_28855;
assign n_39373 =  i_21 &  n_28855;
assign n_39374 = ~n_39372 & ~n_39373;
assign n_39375 =  x_4093 & ~n_39374;
assign n_39376 = ~x_4093 &  n_39374;
assign n_39377 = ~n_39375 & ~n_39376;
assign n_39378 =  x_4092 & ~n_28855;
assign n_39379 =  i_20 &  n_28855;
assign n_39380 = ~n_39378 & ~n_39379;
assign n_39381 =  x_4092 & ~n_39380;
assign n_39382 = ~x_4092 &  n_39380;
assign n_39383 = ~n_39381 & ~n_39382;
assign n_39384 =  x_4091 & ~n_28855;
assign n_39385 =  i_19 &  n_28855;
assign n_39386 = ~n_39384 & ~n_39385;
assign n_39387 =  x_4091 & ~n_39386;
assign n_39388 = ~x_4091 &  n_39386;
assign n_39389 = ~n_39387 & ~n_39388;
assign n_39390 =  x_4090 & ~n_28855;
assign n_39391 =  i_18 &  n_28855;
assign n_39392 = ~n_39390 & ~n_39391;
assign n_39393 =  x_4090 & ~n_39392;
assign n_39394 = ~x_4090 &  n_39392;
assign n_39395 = ~n_39393 & ~n_39394;
assign n_39396 =  x_4089 & ~n_28855;
assign n_39397 =  i_17 &  n_28855;
assign n_39398 = ~n_39396 & ~n_39397;
assign n_39399 =  x_4089 & ~n_39398;
assign n_39400 = ~x_4089 &  n_39398;
assign n_39401 = ~n_39399 & ~n_39400;
assign n_39402 =  x_4088 & ~n_28855;
assign n_39403 =  i_16 &  n_28855;
assign n_39404 = ~n_39402 & ~n_39403;
assign n_39405 =  x_4088 & ~n_39404;
assign n_39406 = ~x_4088 &  n_39404;
assign n_39407 = ~n_39405 & ~n_39406;
assign n_39408 =  x_4087 & ~n_28855;
assign n_39409 =  i_15 &  n_28855;
assign n_39410 = ~n_39408 & ~n_39409;
assign n_39411 =  x_4087 & ~n_39410;
assign n_39412 = ~x_4087 &  n_39410;
assign n_39413 = ~n_39411 & ~n_39412;
assign n_39414 =  x_4086 & ~n_28855;
assign n_39415 =  i_14 &  n_28855;
assign n_39416 = ~n_39414 & ~n_39415;
assign n_39417 =  x_4086 & ~n_39416;
assign n_39418 = ~x_4086 &  n_39416;
assign n_39419 = ~n_39417 & ~n_39418;
assign n_39420 =  x_4085 & ~n_28855;
assign n_39421 =  i_13 &  n_28855;
assign n_39422 = ~n_39420 & ~n_39421;
assign n_39423 =  x_4085 & ~n_39422;
assign n_39424 = ~x_4085 &  n_39422;
assign n_39425 = ~n_39423 & ~n_39424;
assign n_39426 =  x_4084 & ~n_28855;
assign n_39427 =  i_12 &  n_28855;
assign n_39428 = ~n_39426 & ~n_39427;
assign n_39429 =  x_4084 & ~n_39428;
assign n_39430 = ~x_4084 &  n_39428;
assign n_39431 = ~n_39429 & ~n_39430;
assign n_39432 =  x_4083 & ~n_28855;
assign n_39433 =  i_11 &  n_28855;
assign n_39434 = ~n_39432 & ~n_39433;
assign n_39435 =  x_4083 & ~n_39434;
assign n_39436 = ~x_4083 &  n_39434;
assign n_39437 = ~n_39435 & ~n_39436;
assign n_39438 =  x_4082 & ~n_28855;
assign n_39439 =  i_10 &  n_28855;
assign n_39440 = ~n_39438 & ~n_39439;
assign n_39441 =  x_4082 & ~n_39440;
assign n_39442 = ~x_4082 &  n_39440;
assign n_39443 = ~n_39441 & ~n_39442;
assign n_39444 =  x_4081 & ~n_28855;
assign n_39445 =  i_9 &  n_28855;
assign n_39446 = ~n_39444 & ~n_39445;
assign n_39447 =  x_4081 & ~n_39446;
assign n_39448 = ~x_4081 &  n_39446;
assign n_39449 = ~n_39447 & ~n_39448;
assign n_39450 =  x_4080 & ~n_28855;
assign n_39451 =  i_8 &  n_28855;
assign n_39452 = ~n_39450 & ~n_39451;
assign n_39453 =  x_4080 & ~n_39452;
assign n_39454 = ~x_4080 &  n_39452;
assign n_39455 = ~n_39453 & ~n_39454;
assign n_39456 =  x_4079 & ~n_28855;
assign n_39457 =  i_7 &  n_28855;
assign n_39458 = ~n_39456 & ~n_39457;
assign n_39459 =  x_4079 & ~n_39458;
assign n_39460 = ~x_4079 &  n_39458;
assign n_39461 = ~n_39459 & ~n_39460;
assign n_39462 =  x_4078 & ~n_28855;
assign n_39463 =  i_6 &  n_28855;
assign n_39464 = ~n_39462 & ~n_39463;
assign n_39465 =  x_4078 & ~n_39464;
assign n_39466 = ~x_4078 &  n_39464;
assign n_39467 = ~n_39465 & ~n_39466;
assign n_39468 =  x_4077 & ~n_28855;
assign n_39469 =  i_5 &  n_28855;
assign n_39470 = ~n_39468 & ~n_39469;
assign n_39471 =  x_4077 & ~n_39470;
assign n_39472 = ~x_4077 &  n_39470;
assign n_39473 = ~n_39471 & ~n_39472;
assign n_39474 =  x_4076 & ~n_28855;
assign n_39475 =  i_4 &  n_28855;
assign n_39476 = ~n_39474 & ~n_39475;
assign n_39477 =  x_4076 & ~n_39476;
assign n_39478 = ~x_4076 &  n_39476;
assign n_39479 = ~n_39477 & ~n_39478;
assign n_39480 =  x_4075 & ~n_28855;
assign n_39481 =  i_3 &  n_28855;
assign n_39482 = ~n_39480 & ~n_39481;
assign n_39483 =  x_4075 & ~n_39482;
assign n_39484 = ~x_4075 &  n_39482;
assign n_39485 = ~n_39483 & ~n_39484;
assign n_39486 =  x_4074 & ~n_28855;
assign n_39487 =  i_2 &  n_28855;
assign n_39488 = ~n_39486 & ~n_39487;
assign n_39489 =  x_4074 & ~n_39488;
assign n_39490 = ~x_4074 &  n_39488;
assign n_39491 = ~n_39489 & ~n_39490;
assign n_39492 =  x_4073 & ~n_28855;
assign n_39493 =  i_1 &  n_28855;
assign n_39494 = ~n_39492 & ~n_39493;
assign n_39495 =  x_4073 & ~n_39494;
assign n_39496 = ~x_4073 &  n_39494;
assign n_39497 = ~n_39495 & ~n_39496;
assign n_39498 =  n_13872 &  n_8365;
assign n_39499 =  x_4072 & ~n_39498;
assign n_39500 =  x_3160 &  n_39498;
assign n_39501 = ~n_39499 & ~n_39500;
assign n_39502 =  x_4072 & ~n_39501;
assign n_39503 = ~x_4072 &  n_39501;
assign n_39504 = ~n_39502 & ~n_39503;
assign n_39505 =  x_4071 & ~n_39498;
assign n_39506 =  x_3159 &  n_39498;
assign n_39507 = ~n_39505 & ~n_39506;
assign n_39508 =  x_4071 & ~n_39507;
assign n_39509 = ~x_4071 &  n_39507;
assign n_39510 = ~n_39508 & ~n_39509;
assign n_39511 =  x_4070 & ~n_39498;
assign n_39512 =  x_3158 &  n_39498;
assign n_39513 = ~n_39511 & ~n_39512;
assign n_39514 =  x_4070 & ~n_39513;
assign n_39515 = ~x_4070 &  n_39513;
assign n_39516 = ~n_39514 & ~n_39515;
assign n_39517 =  x_4069 & ~n_39498;
assign n_39518 =  x_3157 &  n_39498;
assign n_39519 = ~n_39517 & ~n_39518;
assign n_39520 =  x_4069 & ~n_39519;
assign n_39521 = ~x_4069 &  n_39519;
assign n_39522 = ~n_39520 & ~n_39521;
assign n_39523 =  x_4068 & ~n_39498;
assign n_39524 =  x_3156 &  n_39498;
assign n_39525 = ~n_39523 & ~n_39524;
assign n_39526 =  x_4068 & ~n_39525;
assign n_39527 = ~x_4068 &  n_39525;
assign n_39528 = ~n_39526 & ~n_39527;
assign n_39529 =  x_4067 & ~n_39498;
assign n_39530 =  x_3155 &  n_39498;
assign n_39531 = ~n_39529 & ~n_39530;
assign n_39532 =  x_4067 & ~n_39531;
assign n_39533 = ~x_4067 &  n_39531;
assign n_39534 = ~n_39532 & ~n_39533;
assign n_39535 =  x_4066 & ~n_39498;
assign n_39536 =  x_3154 &  n_39498;
assign n_39537 = ~n_39535 & ~n_39536;
assign n_39538 =  x_4066 & ~n_39537;
assign n_39539 = ~x_4066 &  n_39537;
assign n_39540 = ~n_39538 & ~n_39539;
assign n_39541 =  x_4065 & ~n_39498;
assign n_39542 =  x_3153 &  n_39498;
assign n_39543 = ~n_39541 & ~n_39542;
assign n_39544 =  x_4065 & ~n_39543;
assign n_39545 = ~x_4065 &  n_39543;
assign n_39546 = ~n_39544 & ~n_39545;
assign n_39547 =  x_4064 & ~n_39498;
assign n_39548 =  x_3152 &  n_39498;
assign n_39549 = ~n_39547 & ~n_39548;
assign n_39550 =  x_4064 & ~n_39549;
assign n_39551 = ~x_4064 &  n_39549;
assign n_39552 = ~n_39550 & ~n_39551;
assign n_39553 =  x_4063 & ~n_39498;
assign n_39554 =  x_3151 &  n_39498;
assign n_39555 = ~n_39553 & ~n_39554;
assign n_39556 =  x_4063 & ~n_39555;
assign n_39557 = ~x_4063 &  n_39555;
assign n_39558 = ~n_39556 & ~n_39557;
assign n_39559 =  x_4062 & ~n_39498;
assign n_39560 =  x_3150 &  n_39498;
assign n_39561 = ~n_39559 & ~n_39560;
assign n_39562 =  x_4062 & ~n_39561;
assign n_39563 = ~x_4062 &  n_39561;
assign n_39564 = ~n_39562 & ~n_39563;
assign n_39565 =  x_4061 & ~n_39498;
assign n_39566 =  x_3149 &  n_39498;
assign n_39567 = ~n_39565 & ~n_39566;
assign n_39568 =  x_4061 & ~n_39567;
assign n_39569 = ~x_4061 &  n_39567;
assign n_39570 = ~n_39568 & ~n_39569;
assign n_39571 =  x_4060 & ~n_39498;
assign n_39572 =  x_3148 &  n_39498;
assign n_39573 = ~n_39571 & ~n_39572;
assign n_39574 =  x_4060 & ~n_39573;
assign n_39575 = ~x_4060 &  n_39573;
assign n_39576 = ~n_39574 & ~n_39575;
assign n_39577 =  x_4059 & ~n_39498;
assign n_39578 =  x_3147 &  n_39498;
assign n_39579 = ~n_39577 & ~n_39578;
assign n_39580 =  x_4059 & ~n_39579;
assign n_39581 = ~x_4059 &  n_39579;
assign n_39582 = ~n_39580 & ~n_39581;
assign n_39583 =  x_4058 & ~n_39498;
assign n_39584 =  x_3146 &  n_39498;
assign n_39585 = ~n_39583 & ~n_39584;
assign n_39586 =  x_4058 & ~n_39585;
assign n_39587 = ~x_4058 &  n_39585;
assign n_39588 = ~n_39586 & ~n_39587;
assign n_39589 =  x_4057 & ~n_39498;
assign n_39590 =  x_3145 &  n_39498;
assign n_39591 = ~n_39589 & ~n_39590;
assign n_39592 =  x_4057 & ~n_39591;
assign n_39593 = ~x_4057 &  n_39591;
assign n_39594 = ~n_39592 & ~n_39593;
assign n_39595 =  x_4056 & ~n_39498;
assign n_39596 =  x_3144 &  n_39498;
assign n_39597 = ~n_39595 & ~n_39596;
assign n_39598 =  x_4056 & ~n_39597;
assign n_39599 = ~x_4056 &  n_39597;
assign n_39600 = ~n_39598 & ~n_39599;
assign n_39601 =  x_4055 & ~n_39498;
assign n_39602 =  x_3143 &  n_39498;
assign n_39603 = ~n_39601 & ~n_39602;
assign n_39604 =  x_4055 & ~n_39603;
assign n_39605 = ~x_4055 &  n_39603;
assign n_39606 = ~n_39604 & ~n_39605;
assign n_39607 =  x_4054 & ~n_39498;
assign n_39608 =  x_3142 &  n_39498;
assign n_39609 = ~n_39607 & ~n_39608;
assign n_39610 =  x_4054 & ~n_39609;
assign n_39611 = ~x_4054 &  n_39609;
assign n_39612 = ~n_39610 & ~n_39611;
assign n_39613 =  x_4053 & ~n_39498;
assign n_39614 =  x_3141 &  n_39498;
assign n_39615 = ~n_39613 & ~n_39614;
assign n_39616 =  x_4053 & ~n_39615;
assign n_39617 = ~x_4053 &  n_39615;
assign n_39618 = ~n_39616 & ~n_39617;
assign n_39619 =  x_4052 & ~n_39498;
assign n_39620 =  x_3140 &  n_39498;
assign n_39621 = ~n_39619 & ~n_39620;
assign n_39622 =  x_4052 & ~n_39621;
assign n_39623 = ~x_4052 &  n_39621;
assign n_39624 = ~n_39622 & ~n_39623;
assign n_39625 =  x_4051 & ~n_39498;
assign n_39626 =  x_3139 &  n_39498;
assign n_39627 = ~n_39625 & ~n_39626;
assign n_39628 =  x_4051 & ~n_39627;
assign n_39629 = ~x_4051 &  n_39627;
assign n_39630 = ~n_39628 & ~n_39629;
assign n_39631 =  x_4050 & ~n_39498;
assign n_39632 =  x_3138 &  n_39498;
assign n_39633 = ~n_39631 & ~n_39632;
assign n_39634 =  x_4050 & ~n_39633;
assign n_39635 = ~x_4050 &  n_39633;
assign n_39636 = ~n_39634 & ~n_39635;
assign n_39637 =  x_4049 & ~n_39498;
assign n_39638 =  x_3137 &  n_39498;
assign n_39639 = ~n_39637 & ~n_39638;
assign n_39640 =  x_4049 & ~n_39639;
assign n_39641 = ~x_4049 &  n_39639;
assign n_39642 = ~n_39640 & ~n_39641;
assign n_39643 =  x_4048 & ~n_39498;
assign n_39644 =  x_3136 &  n_39498;
assign n_39645 = ~n_39643 & ~n_39644;
assign n_39646 =  x_4048 & ~n_39645;
assign n_39647 = ~x_4048 &  n_39645;
assign n_39648 = ~n_39646 & ~n_39647;
assign n_39649 =  x_4047 & ~n_39498;
assign n_39650 =  x_3135 &  n_39498;
assign n_39651 = ~n_39649 & ~n_39650;
assign n_39652 =  x_4047 & ~n_39651;
assign n_39653 = ~x_4047 &  n_39651;
assign n_39654 = ~n_39652 & ~n_39653;
assign n_39655 =  x_4046 & ~n_39498;
assign n_39656 =  x_3134 &  n_39498;
assign n_39657 = ~n_39655 & ~n_39656;
assign n_39658 =  x_4046 & ~n_39657;
assign n_39659 = ~x_4046 &  n_39657;
assign n_39660 = ~n_39658 & ~n_39659;
assign n_39661 =  x_4045 & ~n_39498;
assign n_39662 =  x_3133 &  n_39498;
assign n_39663 = ~n_39661 & ~n_39662;
assign n_39664 =  x_4045 & ~n_39663;
assign n_39665 = ~x_4045 &  n_39663;
assign n_39666 = ~n_39664 & ~n_39665;
assign n_39667 =  x_4044 & ~n_39498;
assign n_39668 =  x_3132 &  n_39498;
assign n_39669 = ~n_39667 & ~n_39668;
assign n_39670 =  x_4044 & ~n_39669;
assign n_39671 = ~x_4044 &  n_39669;
assign n_39672 = ~n_39670 & ~n_39671;
assign n_39673 =  x_4043 & ~n_39498;
assign n_39674 =  x_3131 &  n_39498;
assign n_39675 = ~n_39673 & ~n_39674;
assign n_39676 =  x_4043 & ~n_39675;
assign n_39677 = ~x_4043 &  n_39675;
assign n_39678 = ~n_39676 & ~n_39677;
assign n_39679 =  x_4042 & ~n_39498;
assign n_39680 =  x_3130 &  n_39498;
assign n_39681 = ~n_39679 & ~n_39680;
assign n_39682 =  x_4042 & ~n_39681;
assign n_39683 = ~x_4042 &  n_39681;
assign n_39684 = ~n_39682 & ~n_39683;
assign n_39685 =  x_4041 & ~n_39498;
assign n_39686 =  x_3129 &  n_39498;
assign n_39687 = ~n_39685 & ~n_39686;
assign n_39688 =  x_4041 & ~n_39687;
assign n_39689 = ~x_4041 &  n_39687;
assign n_39690 = ~n_39688 & ~n_39689;
assign n_39691 =  x_4040 & ~n_24758;
assign n_39692 =  x_4040 &  n_39691;
assign n_39693 = ~x_4040 & ~n_39691;
assign n_39694 = ~n_39692 & ~n_39693;
assign n_39695 =  x_4039 & ~n_24758;
assign n_39696 =  x_4039 &  n_39695;
assign n_39697 = ~x_4039 & ~n_39695;
assign n_39698 = ~n_39696 & ~n_39697;
assign n_39699 =  x_4038 & ~n_24758;
assign n_39700 =  x_4038 &  n_39699;
assign n_39701 = ~x_4038 & ~n_39699;
assign n_39702 = ~n_39700 & ~n_39701;
assign n_39703 =  x_4037 & ~n_24758;
assign n_39704 =  x_4037 &  n_39703;
assign n_39705 = ~x_4037 & ~n_39703;
assign n_39706 = ~n_39704 & ~n_39705;
assign n_39707 =  x_4036 & ~n_24758;
assign n_39708 =  x_4036 &  n_39707;
assign n_39709 = ~x_4036 & ~n_39707;
assign n_39710 = ~n_39708 & ~n_39709;
assign n_39711 =  x_4035 & ~n_24758;
assign n_39712 =  x_4035 &  n_39711;
assign n_39713 = ~x_4035 & ~n_39711;
assign n_39714 = ~n_39712 & ~n_39713;
assign n_39715 =  x_4034 & ~n_24758;
assign n_39716 =  x_4034 &  n_39715;
assign n_39717 = ~x_4034 & ~n_39715;
assign n_39718 = ~n_39716 & ~n_39717;
assign n_39719 =  x_4033 & ~n_24758;
assign n_39720 =  x_4033 &  n_39719;
assign n_39721 = ~x_4033 & ~n_39719;
assign n_39722 = ~n_39720 & ~n_39721;
assign n_39723 =  x_4032 & ~n_24758;
assign n_39724 =  x_4032 &  n_39723;
assign n_39725 = ~x_4032 & ~n_39723;
assign n_39726 = ~n_39724 & ~n_39725;
assign n_39727 =  x_4031 & ~n_24758;
assign n_39728 =  x_4031 &  n_39727;
assign n_39729 = ~x_4031 & ~n_39727;
assign n_39730 = ~n_39728 & ~n_39729;
assign n_39731 =  x_4030 & ~n_24758;
assign n_39732 =  x_4030 &  n_39731;
assign n_39733 = ~x_4030 & ~n_39731;
assign n_39734 = ~n_39732 & ~n_39733;
assign n_39735 =  x_4029 & ~n_24758;
assign n_39736 =  x_4029 &  n_39735;
assign n_39737 = ~x_4029 & ~n_39735;
assign n_39738 = ~n_39736 & ~n_39737;
assign n_39739 =  x_4028 & ~n_24758;
assign n_39740 =  x_4028 &  n_39739;
assign n_39741 = ~x_4028 & ~n_39739;
assign n_39742 = ~n_39740 & ~n_39741;
assign n_39743 =  x_4027 & ~n_24758;
assign n_39744 =  x_4027 &  n_39743;
assign n_39745 = ~x_4027 & ~n_39743;
assign n_39746 = ~n_39744 & ~n_39745;
assign n_39747 =  x_4026 & ~n_24758;
assign n_39748 =  x_4026 &  n_39747;
assign n_39749 = ~x_4026 & ~n_39747;
assign n_39750 = ~n_39748 & ~n_39749;
assign n_39751 =  x_4025 & ~n_24758;
assign n_39752 =  x_4025 &  n_39751;
assign n_39753 = ~x_4025 & ~n_39751;
assign n_39754 = ~n_39752 & ~n_39753;
assign n_39755 =  x_4024 & ~n_24758;
assign n_39756 =  x_4024 &  n_39755;
assign n_39757 = ~x_4024 & ~n_39755;
assign n_39758 = ~n_39756 & ~n_39757;
assign n_39759 =  x_4023 & ~n_24758;
assign n_39760 =  x_4023 &  n_39759;
assign n_39761 = ~x_4023 & ~n_39759;
assign n_39762 = ~n_39760 & ~n_39761;
assign n_39763 =  x_4022 & ~n_24758;
assign n_39764 =  x_4022 &  n_39763;
assign n_39765 = ~x_4022 & ~n_39763;
assign n_39766 = ~n_39764 & ~n_39765;
assign n_39767 =  x_4021 & ~n_24758;
assign n_39768 =  x_4021 &  n_39767;
assign n_39769 = ~x_4021 & ~n_39767;
assign n_39770 = ~n_39768 & ~n_39769;
assign n_39771 =  x_4020 & ~n_24758;
assign n_39772 =  x_4020 &  n_39771;
assign n_39773 = ~x_4020 & ~n_39771;
assign n_39774 = ~n_39772 & ~n_39773;
assign n_39775 =  x_4019 & ~n_24758;
assign n_39776 =  x_4019 &  n_39775;
assign n_39777 = ~x_4019 & ~n_39775;
assign n_39778 = ~n_39776 & ~n_39777;
assign n_39779 =  x_4018 & ~n_24758;
assign n_39780 =  x_4018 &  n_39779;
assign n_39781 = ~x_4018 & ~n_39779;
assign n_39782 = ~n_39780 & ~n_39781;
assign n_39783 =  x_4017 & ~n_24758;
assign n_39784 =  x_4017 &  n_39783;
assign n_39785 = ~x_4017 & ~n_39783;
assign n_39786 = ~n_39784 & ~n_39785;
assign n_39787 =  x_4016 & ~n_24758;
assign n_39788 =  x_4016 &  n_39787;
assign n_39789 = ~x_4016 & ~n_39787;
assign n_39790 = ~n_39788 & ~n_39789;
assign n_39791 =  x_4015 & ~n_24758;
assign n_39792 =  x_4015 &  n_39791;
assign n_39793 = ~x_4015 & ~n_39791;
assign n_39794 = ~n_39792 & ~n_39793;
assign n_39795 =  x_4014 & ~n_24758;
assign n_39796 =  x_4014 &  n_39795;
assign n_39797 = ~x_4014 & ~n_39795;
assign n_39798 = ~n_39796 & ~n_39797;
assign n_39799 =  x_4013 & ~n_24758;
assign n_39800 =  x_4013 &  n_39799;
assign n_39801 = ~x_4013 & ~n_39799;
assign n_39802 = ~n_39800 & ~n_39801;
assign n_39803 =  x_4012 & ~n_24758;
assign n_39804 =  x_4012 &  n_39803;
assign n_39805 = ~x_4012 & ~n_39803;
assign n_39806 = ~n_39804 & ~n_39805;
assign n_39807 =  x_4011 & ~n_24758;
assign n_39808 =  x_4011 &  n_39807;
assign n_39809 = ~x_4011 & ~n_39807;
assign n_39810 = ~n_39808 & ~n_39809;
assign n_39811 =  x_4010 & ~n_24758;
assign n_39812 =  x_4010 &  n_39811;
assign n_39813 = ~x_4010 & ~n_39811;
assign n_39814 = ~n_39812 & ~n_39813;
assign n_39815 =  x_4009 & ~n_24758;
assign n_39816 =  x_4009 &  n_39815;
assign n_39817 = ~x_4009 & ~n_39815;
assign n_39818 = ~n_39816 & ~n_39817;
assign n_39819 =  x_4008 & ~n_27023;
assign n_39820 =  x_2937 &  n_27023;
assign n_39821 = ~n_39819 & ~n_39820;
assign n_39822 =  x_4008 & ~n_39821;
assign n_39823 = ~x_4008 &  n_39821;
assign n_39824 = ~n_39822 & ~n_39823;
assign n_39825 =  x_4007 & ~n_27023;
assign n_39826 =  x_2936 &  n_27023;
assign n_39827 = ~n_39825 & ~n_39826;
assign n_39828 =  x_4007 & ~n_39827;
assign n_39829 = ~x_4007 &  n_39827;
assign n_39830 = ~n_39828 & ~n_39829;
assign n_39831 =  x_4006 & ~n_27023;
assign n_39832 =  x_2935 &  n_27023;
assign n_39833 = ~n_39831 & ~n_39832;
assign n_39834 =  x_4006 & ~n_39833;
assign n_39835 = ~x_4006 &  n_39833;
assign n_39836 = ~n_39834 & ~n_39835;
assign n_39837 =  x_4005 & ~n_27023;
assign n_39838 =  x_2934 &  n_27023;
assign n_39839 = ~n_39837 & ~n_39838;
assign n_39840 =  x_4005 & ~n_39839;
assign n_39841 = ~x_4005 &  n_39839;
assign n_39842 = ~n_39840 & ~n_39841;
assign n_39843 =  x_4004 & ~n_27023;
assign n_39844 =  x_2933 &  n_27023;
assign n_39845 = ~n_39843 & ~n_39844;
assign n_39846 =  x_4004 & ~n_39845;
assign n_39847 = ~x_4004 &  n_39845;
assign n_39848 = ~n_39846 & ~n_39847;
assign n_39849 =  x_4003 & ~n_27023;
assign n_39850 =  x_2932 &  n_27023;
assign n_39851 = ~n_39849 & ~n_39850;
assign n_39852 =  x_4003 & ~n_39851;
assign n_39853 = ~x_4003 &  n_39851;
assign n_39854 = ~n_39852 & ~n_39853;
assign n_39855 =  x_4002 & ~n_27023;
assign n_39856 =  x_2931 &  n_27023;
assign n_39857 = ~n_39855 & ~n_39856;
assign n_39858 =  x_4002 & ~n_39857;
assign n_39859 = ~x_4002 &  n_39857;
assign n_39860 = ~n_39858 & ~n_39859;
assign n_39861 =  x_4001 & ~n_27023;
assign n_39862 =  x_2930 &  n_27023;
assign n_39863 = ~n_39861 & ~n_39862;
assign n_39864 =  x_4001 & ~n_39863;
assign n_39865 = ~x_4001 &  n_39863;
assign n_39866 = ~n_39864 & ~n_39865;
assign n_39867 =  x_4000 & ~n_27023;
assign n_39868 =  x_2929 &  n_27023;
assign n_39869 = ~n_39867 & ~n_39868;
assign n_39870 =  x_4000 & ~n_39869;
assign n_39871 = ~x_4000 &  n_39869;
assign n_39872 = ~n_39870 & ~n_39871;
assign n_39873 =  x_3999 & ~n_27023;
assign n_39874 =  x_2928 &  n_27023;
assign n_39875 = ~n_39873 & ~n_39874;
assign n_39876 =  x_3999 & ~n_39875;
assign n_39877 = ~x_3999 &  n_39875;
assign n_39878 = ~n_39876 & ~n_39877;
assign n_39879 =  x_3998 & ~n_27023;
assign n_39880 =  x_2927 &  n_27023;
assign n_39881 = ~n_39879 & ~n_39880;
assign n_39882 =  x_3998 & ~n_39881;
assign n_39883 = ~x_3998 &  n_39881;
assign n_39884 = ~n_39882 & ~n_39883;
assign n_39885 =  x_3997 & ~n_27023;
assign n_39886 =  x_2926 &  n_27023;
assign n_39887 = ~n_39885 & ~n_39886;
assign n_39888 =  x_3997 & ~n_39887;
assign n_39889 = ~x_3997 &  n_39887;
assign n_39890 = ~n_39888 & ~n_39889;
assign n_39891 =  x_3996 & ~n_27023;
assign n_39892 =  x_2925 &  n_27023;
assign n_39893 = ~n_39891 & ~n_39892;
assign n_39894 =  x_3996 & ~n_39893;
assign n_39895 = ~x_3996 &  n_39893;
assign n_39896 = ~n_39894 & ~n_39895;
assign n_39897 =  x_3995 & ~n_27023;
assign n_39898 =  x_2924 &  n_27023;
assign n_39899 = ~n_39897 & ~n_39898;
assign n_39900 =  x_3995 & ~n_39899;
assign n_39901 = ~x_3995 &  n_39899;
assign n_39902 = ~n_39900 & ~n_39901;
assign n_39903 =  x_3994 & ~n_27023;
assign n_39904 =  x_2923 &  n_27023;
assign n_39905 = ~n_39903 & ~n_39904;
assign n_39906 =  x_3994 & ~n_39905;
assign n_39907 = ~x_3994 &  n_39905;
assign n_39908 = ~n_39906 & ~n_39907;
assign n_39909 =  x_3993 & ~n_27023;
assign n_39910 =  x_2922 &  n_27023;
assign n_39911 = ~n_39909 & ~n_39910;
assign n_39912 =  x_3993 & ~n_39911;
assign n_39913 = ~x_3993 &  n_39911;
assign n_39914 = ~n_39912 & ~n_39913;
assign n_39915 =  x_3992 & ~n_27023;
assign n_39916 =  x_2921 &  n_27023;
assign n_39917 = ~n_39915 & ~n_39916;
assign n_39918 =  x_3992 & ~n_39917;
assign n_39919 = ~x_3992 &  n_39917;
assign n_39920 = ~n_39918 & ~n_39919;
assign n_39921 =  x_3991 & ~n_27023;
assign n_39922 =  x_2920 &  n_27023;
assign n_39923 = ~n_39921 & ~n_39922;
assign n_39924 =  x_3991 & ~n_39923;
assign n_39925 = ~x_3991 &  n_39923;
assign n_39926 = ~n_39924 & ~n_39925;
assign n_39927 =  x_3990 & ~n_27023;
assign n_39928 =  x_2919 &  n_27023;
assign n_39929 = ~n_39927 & ~n_39928;
assign n_39930 =  x_3990 & ~n_39929;
assign n_39931 = ~x_3990 &  n_39929;
assign n_39932 = ~n_39930 & ~n_39931;
assign n_39933 =  x_3989 & ~n_27023;
assign n_39934 =  x_2918 &  n_27023;
assign n_39935 = ~n_39933 & ~n_39934;
assign n_39936 =  x_3989 & ~n_39935;
assign n_39937 = ~x_3989 &  n_39935;
assign n_39938 = ~n_39936 & ~n_39937;
assign n_39939 =  x_3988 & ~n_27023;
assign n_39940 =  x_2917 &  n_27023;
assign n_39941 = ~n_39939 & ~n_39940;
assign n_39942 =  x_3988 & ~n_39941;
assign n_39943 = ~x_3988 &  n_39941;
assign n_39944 = ~n_39942 & ~n_39943;
assign n_39945 =  x_3987 & ~n_27023;
assign n_39946 =  x_2916 &  n_27023;
assign n_39947 = ~n_39945 & ~n_39946;
assign n_39948 =  x_3987 & ~n_39947;
assign n_39949 = ~x_3987 &  n_39947;
assign n_39950 = ~n_39948 & ~n_39949;
assign n_39951 =  x_3986 & ~n_27023;
assign n_39952 =  x_2915 &  n_27023;
assign n_39953 = ~n_39951 & ~n_39952;
assign n_39954 =  x_3986 & ~n_39953;
assign n_39955 = ~x_3986 &  n_39953;
assign n_39956 = ~n_39954 & ~n_39955;
assign n_39957 =  x_3985 & ~n_27023;
assign n_39958 =  x_2914 &  n_27023;
assign n_39959 = ~n_39957 & ~n_39958;
assign n_39960 =  x_3985 & ~n_39959;
assign n_39961 = ~x_3985 &  n_39959;
assign n_39962 = ~n_39960 & ~n_39961;
assign n_39963 =  x_3984 & ~n_27023;
assign n_39964 =  x_2913 &  n_27023;
assign n_39965 = ~n_39963 & ~n_39964;
assign n_39966 =  x_3984 & ~n_39965;
assign n_39967 = ~x_3984 &  n_39965;
assign n_39968 = ~n_39966 & ~n_39967;
assign n_39969 =  x_3983 & ~n_27023;
assign n_39970 =  x_2912 &  n_27023;
assign n_39971 = ~n_39969 & ~n_39970;
assign n_39972 =  x_3983 & ~n_39971;
assign n_39973 = ~x_3983 &  n_39971;
assign n_39974 = ~n_39972 & ~n_39973;
assign n_39975 =  x_3982 & ~n_27023;
assign n_39976 =  x_2911 &  n_27023;
assign n_39977 = ~n_39975 & ~n_39976;
assign n_39978 =  x_3982 & ~n_39977;
assign n_39979 = ~x_3982 &  n_39977;
assign n_39980 = ~n_39978 & ~n_39979;
assign n_39981 =  x_3981 & ~n_27023;
assign n_39982 =  x_2910 &  n_27023;
assign n_39983 = ~n_39981 & ~n_39982;
assign n_39984 =  x_3981 & ~n_39983;
assign n_39985 = ~x_3981 &  n_39983;
assign n_39986 = ~n_39984 & ~n_39985;
assign n_39987 =  x_3980 & ~n_27023;
assign n_39988 =  x_2909 &  n_27023;
assign n_39989 = ~n_39987 & ~n_39988;
assign n_39990 =  x_3980 & ~n_39989;
assign n_39991 = ~x_3980 &  n_39989;
assign n_39992 = ~n_39990 & ~n_39991;
assign n_39993 =  x_3979 & ~n_27023;
assign n_39994 =  x_2908 &  n_27023;
assign n_39995 = ~n_39993 & ~n_39994;
assign n_39996 =  x_3979 & ~n_39995;
assign n_39997 = ~x_3979 &  n_39995;
assign n_39998 = ~n_39996 & ~n_39997;
assign n_39999 =  x_3978 & ~n_27023;
assign n_40000 =  x_2907 &  n_27023;
assign n_40001 = ~n_39999 & ~n_40000;
assign n_40002 =  x_3978 & ~n_40001;
assign n_40003 = ~x_3978 &  n_40001;
assign n_40004 = ~n_40002 & ~n_40003;
assign n_40005 =  x_3977 & ~n_27023;
assign n_40006 =  x_3977 &  n_40005;
assign n_40007 = ~x_3977 & ~n_40005;
assign n_40008 = ~n_40006 & ~n_40007;
assign n_40009 =  x_3976 & ~n_25650;
assign n_40010 =  i_32 &  n_25650;
assign n_40011 = ~n_40009 & ~n_40010;
assign n_40012 =  x_3976 & ~n_40011;
assign n_40013 = ~x_3976 &  n_40011;
assign n_40014 = ~n_40012 & ~n_40013;
assign n_40015 =  x_3975 & ~n_25650;
assign n_40016 =  i_31 &  n_25650;
assign n_40017 = ~n_40015 & ~n_40016;
assign n_40018 =  x_3975 & ~n_40017;
assign n_40019 = ~x_3975 &  n_40017;
assign n_40020 = ~n_40018 & ~n_40019;
assign n_40021 =  x_3974 & ~n_25650;
assign n_40022 =  i_30 &  n_25650;
assign n_40023 = ~n_40021 & ~n_40022;
assign n_40024 =  x_3974 & ~n_40023;
assign n_40025 = ~x_3974 &  n_40023;
assign n_40026 = ~n_40024 & ~n_40025;
assign n_40027 =  x_3973 & ~n_25650;
assign n_40028 =  i_29 &  n_25650;
assign n_40029 = ~n_40027 & ~n_40028;
assign n_40030 =  x_3973 & ~n_40029;
assign n_40031 = ~x_3973 &  n_40029;
assign n_40032 = ~n_40030 & ~n_40031;
assign n_40033 =  x_3972 & ~n_25650;
assign n_40034 =  i_28 &  n_25650;
assign n_40035 = ~n_40033 & ~n_40034;
assign n_40036 =  x_3972 & ~n_40035;
assign n_40037 = ~x_3972 &  n_40035;
assign n_40038 = ~n_40036 & ~n_40037;
assign n_40039 =  x_3971 & ~n_25650;
assign n_40040 =  i_27 &  n_25650;
assign n_40041 = ~n_40039 & ~n_40040;
assign n_40042 =  x_3971 & ~n_40041;
assign n_40043 = ~x_3971 &  n_40041;
assign n_40044 = ~n_40042 & ~n_40043;
assign n_40045 =  x_3970 & ~n_25650;
assign n_40046 =  i_26 &  n_25650;
assign n_40047 = ~n_40045 & ~n_40046;
assign n_40048 =  x_3970 & ~n_40047;
assign n_40049 = ~x_3970 &  n_40047;
assign n_40050 = ~n_40048 & ~n_40049;
assign n_40051 =  x_3969 & ~n_25650;
assign n_40052 =  i_25 &  n_25650;
assign n_40053 = ~n_40051 & ~n_40052;
assign n_40054 =  x_3969 & ~n_40053;
assign n_40055 = ~x_3969 &  n_40053;
assign n_40056 = ~n_40054 & ~n_40055;
assign n_40057 =  x_3968 & ~n_25650;
assign n_40058 =  i_24 &  n_25650;
assign n_40059 = ~n_40057 & ~n_40058;
assign n_40060 =  x_3968 & ~n_40059;
assign n_40061 = ~x_3968 &  n_40059;
assign n_40062 = ~n_40060 & ~n_40061;
assign n_40063 =  x_3967 & ~n_25650;
assign n_40064 =  i_23 &  n_25650;
assign n_40065 = ~n_40063 & ~n_40064;
assign n_40066 =  x_3967 & ~n_40065;
assign n_40067 = ~x_3967 &  n_40065;
assign n_40068 = ~n_40066 & ~n_40067;
assign n_40069 =  x_3966 & ~n_25650;
assign n_40070 =  i_22 &  n_25650;
assign n_40071 = ~n_40069 & ~n_40070;
assign n_40072 =  x_3966 & ~n_40071;
assign n_40073 = ~x_3966 &  n_40071;
assign n_40074 = ~n_40072 & ~n_40073;
assign n_40075 =  x_3965 & ~n_25650;
assign n_40076 =  i_21 &  n_25650;
assign n_40077 = ~n_40075 & ~n_40076;
assign n_40078 =  x_3965 & ~n_40077;
assign n_40079 = ~x_3965 &  n_40077;
assign n_40080 = ~n_40078 & ~n_40079;
assign n_40081 =  x_3964 & ~n_25650;
assign n_40082 =  i_20 &  n_25650;
assign n_40083 = ~n_40081 & ~n_40082;
assign n_40084 =  x_3964 & ~n_40083;
assign n_40085 = ~x_3964 &  n_40083;
assign n_40086 = ~n_40084 & ~n_40085;
assign n_40087 =  x_3963 & ~n_25650;
assign n_40088 =  i_19 &  n_25650;
assign n_40089 = ~n_40087 & ~n_40088;
assign n_40090 =  x_3963 & ~n_40089;
assign n_40091 = ~x_3963 &  n_40089;
assign n_40092 = ~n_40090 & ~n_40091;
assign n_40093 =  x_3962 & ~n_25650;
assign n_40094 =  i_18 &  n_25650;
assign n_40095 = ~n_40093 & ~n_40094;
assign n_40096 =  x_3962 & ~n_40095;
assign n_40097 = ~x_3962 &  n_40095;
assign n_40098 = ~n_40096 & ~n_40097;
assign n_40099 =  x_3961 & ~n_25650;
assign n_40100 =  i_17 &  n_25650;
assign n_40101 = ~n_40099 & ~n_40100;
assign n_40102 =  x_3961 & ~n_40101;
assign n_40103 = ~x_3961 &  n_40101;
assign n_40104 = ~n_40102 & ~n_40103;
assign n_40105 =  x_3960 & ~n_25650;
assign n_40106 =  i_16 &  n_25650;
assign n_40107 = ~n_40105 & ~n_40106;
assign n_40108 =  x_3960 & ~n_40107;
assign n_40109 = ~x_3960 &  n_40107;
assign n_40110 = ~n_40108 & ~n_40109;
assign n_40111 =  x_3959 & ~n_25650;
assign n_40112 =  i_15 &  n_25650;
assign n_40113 = ~n_40111 & ~n_40112;
assign n_40114 =  x_3959 & ~n_40113;
assign n_40115 = ~x_3959 &  n_40113;
assign n_40116 = ~n_40114 & ~n_40115;
assign n_40117 =  x_3958 & ~n_25650;
assign n_40118 =  i_14 &  n_25650;
assign n_40119 = ~n_40117 & ~n_40118;
assign n_40120 =  x_3958 & ~n_40119;
assign n_40121 = ~x_3958 &  n_40119;
assign n_40122 = ~n_40120 & ~n_40121;
assign n_40123 =  x_3957 & ~n_25650;
assign n_40124 =  i_13 &  n_25650;
assign n_40125 = ~n_40123 & ~n_40124;
assign n_40126 =  x_3957 & ~n_40125;
assign n_40127 = ~x_3957 &  n_40125;
assign n_40128 = ~n_40126 & ~n_40127;
assign n_40129 =  x_3956 & ~n_25650;
assign n_40130 =  i_12 &  n_25650;
assign n_40131 = ~n_40129 & ~n_40130;
assign n_40132 =  x_3956 & ~n_40131;
assign n_40133 = ~x_3956 &  n_40131;
assign n_40134 = ~n_40132 & ~n_40133;
assign n_40135 =  x_3955 & ~n_25650;
assign n_40136 =  i_11 &  n_25650;
assign n_40137 = ~n_40135 & ~n_40136;
assign n_40138 =  x_3955 & ~n_40137;
assign n_40139 = ~x_3955 &  n_40137;
assign n_40140 = ~n_40138 & ~n_40139;
assign n_40141 =  x_3954 & ~n_25650;
assign n_40142 =  i_10 &  n_25650;
assign n_40143 = ~n_40141 & ~n_40142;
assign n_40144 =  x_3954 & ~n_40143;
assign n_40145 = ~x_3954 &  n_40143;
assign n_40146 = ~n_40144 & ~n_40145;
assign n_40147 =  x_3953 & ~n_25650;
assign n_40148 =  i_9 &  n_25650;
assign n_40149 = ~n_40147 & ~n_40148;
assign n_40150 =  x_3953 & ~n_40149;
assign n_40151 = ~x_3953 &  n_40149;
assign n_40152 = ~n_40150 & ~n_40151;
assign n_40153 =  x_3952 & ~n_25650;
assign n_40154 =  i_8 &  n_25650;
assign n_40155 = ~n_40153 & ~n_40154;
assign n_40156 =  x_3952 & ~n_40155;
assign n_40157 = ~x_3952 &  n_40155;
assign n_40158 = ~n_40156 & ~n_40157;
assign n_40159 =  x_3951 & ~n_25650;
assign n_40160 =  i_7 &  n_25650;
assign n_40161 = ~n_40159 & ~n_40160;
assign n_40162 =  x_3951 & ~n_40161;
assign n_40163 = ~x_3951 &  n_40161;
assign n_40164 = ~n_40162 & ~n_40163;
assign n_40165 =  x_3950 & ~n_25650;
assign n_40166 =  i_6 &  n_25650;
assign n_40167 = ~n_40165 & ~n_40166;
assign n_40168 =  x_3950 & ~n_40167;
assign n_40169 = ~x_3950 &  n_40167;
assign n_40170 = ~n_40168 & ~n_40169;
assign n_40171 =  x_3949 & ~n_25650;
assign n_40172 =  i_5 &  n_25650;
assign n_40173 = ~n_40171 & ~n_40172;
assign n_40174 =  x_3949 & ~n_40173;
assign n_40175 = ~x_3949 &  n_40173;
assign n_40176 = ~n_40174 & ~n_40175;
assign n_40177 =  x_3948 & ~n_25650;
assign n_40178 =  i_4 &  n_25650;
assign n_40179 = ~n_40177 & ~n_40178;
assign n_40180 =  x_3948 & ~n_40179;
assign n_40181 = ~x_3948 &  n_40179;
assign n_40182 = ~n_40180 & ~n_40181;
assign n_40183 =  x_3947 & ~n_25650;
assign n_40184 =  i_3 &  n_25650;
assign n_40185 = ~n_40183 & ~n_40184;
assign n_40186 =  x_3947 & ~n_40185;
assign n_40187 = ~x_3947 &  n_40185;
assign n_40188 = ~n_40186 & ~n_40187;
assign n_40189 =  x_3946 & ~n_25650;
assign n_40190 =  i_2 &  n_25650;
assign n_40191 = ~n_40189 & ~n_40190;
assign n_40192 =  x_3946 & ~n_40191;
assign n_40193 = ~x_3946 &  n_40191;
assign n_40194 = ~n_40192 & ~n_40193;
assign n_40195 =  x_3945 & ~n_25650;
assign n_40196 =  i_1 &  n_25650;
assign n_40197 = ~n_40195 & ~n_40196;
assign n_40198 =  x_3945 & ~n_40197;
assign n_40199 = ~x_3945 &  n_40197;
assign n_40200 = ~n_40198 & ~n_40199;
assign n_40201 = ~n_25236 & ~n_26458;
assign n_40202 =  x_43 & ~n_40201;
assign n_40203 =  x_3944 & ~n_40202;
assign n_40204 =  i_32 &  n_40202;
assign n_40205 = ~n_40203 & ~n_40204;
assign n_40206 =  x_3944 & ~n_40205;
assign n_40207 = ~x_3944 &  n_40205;
assign n_40208 = ~n_40206 & ~n_40207;
assign n_40209 =  x_3943 & ~n_40202;
assign n_40210 =  i_31 &  n_40202;
assign n_40211 = ~n_40209 & ~n_40210;
assign n_40212 =  x_3943 & ~n_40211;
assign n_40213 = ~x_3943 &  n_40211;
assign n_40214 = ~n_40212 & ~n_40213;
assign n_40215 =  x_3942 & ~n_40202;
assign n_40216 =  i_30 &  n_40202;
assign n_40217 = ~n_40215 & ~n_40216;
assign n_40218 =  x_3942 & ~n_40217;
assign n_40219 = ~x_3942 &  n_40217;
assign n_40220 = ~n_40218 & ~n_40219;
assign n_40221 =  x_3941 & ~n_40202;
assign n_40222 =  i_29 &  n_40202;
assign n_40223 = ~n_40221 & ~n_40222;
assign n_40224 =  x_3941 & ~n_40223;
assign n_40225 = ~x_3941 &  n_40223;
assign n_40226 = ~n_40224 & ~n_40225;
assign n_40227 =  x_3940 & ~n_40202;
assign n_40228 =  i_28 &  n_40202;
assign n_40229 = ~n_40227 & ~n_40228;
assign n_40230 =  x_3940 & ~n_40229;
assign n_40231 = ~x_3940 &  n_40229;
assign n_40232 = ~n_40230 & ~n_40231;
assign n_40233 =  x_3939 & ~n_40202;
assign n_40234 =  i_27 &  n_40202;
assign n_40235 = ~n_40233 & ~n_40234;
assign n_40236 =  x_3939 & ~n_40235;
assign n_40237 = ~x_3939 &  n_40235;
assign n_40238 = ~n_40236 & ~n_40237;
assign n_40239 =  x_3938 & ~n_40202;
assign n_40240 =  i_26 &  n_40202;
assign n_40241 = ~n_40239 & ~n_40240;
assign n_40242 =  x_3938 & ~n_40241;
assign n_40243 = ~x_3938 &  n_40241;
assign n_40244 = ~n_40242 & ~n_40243;
assign n_40245 =  x_3937 & ~n_40202;
assign n_40246 =  i_25 &  n_40202;
assign n_40247 = ~n_40245 & ~n_40246;
assign n_40248 =  x_3937 & ~n_40247;
assign n_40249 = ~x_3937 &  n_40247;
assign n_40250 = ~n_40248 & ~n_40249;
assign n_40251 =  x_3936 & ~n_40202;
assign n_40252 =  i_24 &  n_40202;
assign n_40253 = ~n_40251 & ~n_40252;
assign n_40254 =  x_3936 & ~n_40253;
assign n_40255 = ~x_3936 &  n_40253;
assign n_40256 = ~n_40254 & ~n_40255;
assign n_40257 =  x_3935 & ~n_40202;
assign n_40258 =  i_23 &  n_40202;
assign n_40259 = ~n_40257 & ~n_40258;
assign n_40260 =  x_3935 & ~n_40259;
assign n_40261 = ~x_3935 &  n_40259;
assign n_40262 = ~n_40260 & ~n_40261;
assign n_40263 =  x_3934 & ~n_40202;
assign n_40264 =  i_22 &  n_40202;
assign n_40265 = ~n_40263 & ~n_40264;
assign n_40266 =  x_3934 & ~n_40265;
assign n_40267 = ~x_3934 &  n_40265;
assign n_40268 = ~n_40266 & ~n_40267;
assign n_40269 =  x_3933 & ~n_40202;
assign n_40270 =  i_21 &  n_40202;
assign n_40271 = ~n_40269 & ~n_40270;
assign n_40272 =  x_3933 & ~n_40271;
assign n_40273 = ~x_3933 &  n_40271;
assign n_40274 = ~n_40272 & ~n_40273;
assign n_40275 =  x_3932 & ~n_40202;
assign n_40276 =  i_20 &  n_40202;
assign n_40277 = ~n_40275 & ~n_40276;
assign n_40278 =  x_3932 & ~n_40277;
assign n_40279 = ~x_3932 &  n_40277;
assign n_40280 = ~n_40278 & ~n_40279;
assign n_40281 =  x_3931 & ~n_40202;
assign n_40282 =  i_19 &  n_40202;
assign n_40283 = ~n_40281 & ~n_40282;
assign n_40284 =  x_3931 & ~n_40283;
assign n_40285 = ~x_3931 &  n_40283;
assign n_40286 = ~n_40284 & ~n_40285;
assign n_40287 =  x_3930 & ~n_40202;
assign n_40288 =  i_18 &  n_40202;
assign n_40289 = ~n_40287 & ~n_40288;
assign n_40290 =  x_3930 & ~n_40289;
assign n_40291 = ~x_3930 &  n_40289;
assign n_40292 = ~n_40290 & ~n_40291;
assign n_40293 =  x_3929 & ~n_40202;
assign n_40294 =  i_17 &  n_40202;
assign n_40295 = ~n_40293 & ~n_40294;
assign n_40296 =  x_3929 & ~n_40295;
assign n_40297 = ~x_3929 &  n_40295;
assign n_40298 = ~n_40296 & ~n_40297;
assign n_40299 =  x_3928 & ~n_40202;
assign n_40300 =  i_16 &  n_40202;
assign n_40301 = ~n_40299 & ~n_40300;
assign n_40302 =  x_3928 & ~n_40301;
assign n_40303 = ~x_3928 &  n_40301;
assign n_40304 = ~n_40302 & ~n_40303;
assign n_40305 =  x_3927 & ~n_40202;
assign n_40306 =  i_15 &  n_40202;
assign n_40307 = ~n_40305 & ~n_40306;
assign n_40308 =  x_3927 & ~n_40307;
assign n_40309 = ~x_3927 &  n_40307;
assign n_40310 = ~n_40308 & ~n_40309;
assign n_40311 =  x_3926 & ~n_40202;
assign n_40312 =  i_14 &  n_40202;
assign n_40313 = ~n_40311 & ~n_40312;
assign n_40314 =  x_3926 & ~n_40313;
assign n_40315 = ~x_3926 &  n_40313;
assign n_40316 = ~n_40314 & ~n_40315;
assign n_40317 =  x_3925 & ~n_40202;
assign n_40318 =  i_13 &  n_40202;
assign n_40319 = ~n_40317 & ~n_40318;
assign n_40320 =  x_3925 & ~n_40319;
assign n_40321 = ~x_3925 &  n_40319;
assign n_40322 = ~n_40320 & ~n_40321;
assign n_40323 =  x_3924 & ~n_40202;
assign n_40324 =  i_12 &  n_40202;
assign n_40325 = ~n_40323 & ~n_40324;
assign n_40326 =  x_3924 & ~n_40325;
assign n_40327 = ~x_3924 &  n_40325;
assign n_40328 = ~n_40326 & ~n_40327;
assign n_40329 =  x_3923 & ~n_40202;
assign n_40330 =  i_11 &  n_40202;
assign n_40331 = ~n_40329 & ~n_40330;
assign n_40332 =  x_3923 & ~n_40331;
assign n_40333 = ~x_3923 &  n_40331;
assign n_40334 = ~n_40332 & ~n_40333;
assign n_40335 =  x_3922 & ~n_40202;
assign n_40336 =  i_10 &  n_40202;
assign n_40337 = ~n_40335 & ~n_40336;
assign n_40338 =  x_3922 & ~n_40337;
assign n_40339 = ~x_3922 &  n_40337;
assign n_40340 = ~n_40338 & ~n_40339;
assign n_40341 =  x_3921 & ~n_40202;
assign n_40342 =  i_9 &  n_40202;
assign n_40343 = ~n_40341 & ~n_40342;
assign n_40344 =  x_3921 & ~n_40343;
assign n_40345 = ~x_3921 &  n_40343;
assign n_40346 = ~n_40344 & ~n_40345;
assign n_40347 =  x_3920 & ~n_40202;
assign n_40348 =  i_8 &  n_40202;
assign n_40349 = ~n_40347 & ~n_40348;
assign n_40350 =  x_3920 & ~n_40349;
assign n_40351 = ~x_3920 &  n_40349;
assign n_40352 = ~n_40350 & ~n_40351;
assign n_40353 =  x_3919 & ~n_40202;
assign n_40354 =  i_7 &  n_40202;
assign n_40355 = ~n_40353 & ~n_40354;
assign n_40356 =  x_3919 & ~n_40355;
assign n_40357 = ~x_3919 &  n_40355;
assign n_40358 = ~n_40356 & ~n_40357;
assign n_40359 =  x_3918 & ~n_40202;
assign n_40360 =  i_6 &  n_40202;
assign n_40361 = ~n_40359 & ~n_40360;
assign n_40362 =  x_3918 & ~n_40361;
assign n_40363 = ~x_3918 &  n_40361;
assign n_40364 = ~n_40362 & ~n_40363;
assign n_40365 =  x_3917 & ~n_40202;
assign n_40366 =  i_5 &  n_40202;
assign n_40367 = ~n_40365 & ~n_40366;
assign n_40368 =  x_3917 & ~n_40367;
assign n_40369 = ~x_3917 &  n_40367;
assign n_40370 = ~n_40368 & ~n_40369;
assign n_40371 =  x_3916 & ~n_40202;
assign n_40372 =  i_4 &  n_40202;
assign n_40373 = ~n_40371 & ~n_40372;
assign n_40374 =  x_3916 & ~n_40373;
assign n_40375 = ~x_3916 &  n_40373;
assign n_40376 = ~n_40374 & ~n_40375;
assign n_40377 =  x_3915 & ~n_40202;
assign n_40378 =  i_3 &  n_40202;
assign n_40379 = ~n_40377 & ~n_40378;
assign n_40380 =  x_3915 & ~n_40379;
assign n_40381 = ~x_3915 &  n_40379;
assign n_40382 = ~n_40380 & ~n_40381;
assign n_40383 =  x_3914 & ~n_40202;
assign n_40384 =  i_2 &  n_40202;
assign n_40385 = ~n_40383 & ~n_40384;
assign n_40386 =  x_3914 & ~n_40385;
assign n_40387 = ~x_3914 &  n_40385;
assign n_40388 = ~n_40386 & ~n_40387;
assign n_40389 =  x_3913 & ~n_40202;
assign n_40390 =  i_1 &  n_40202;
assign n_40391 = ~n_40389 & ~n_40390;
assign n_40392 =  x_3913 & ~n_40391;
assign n_40393 = ~x_3913 &  n_40391;
assign n_40394 = ~n_40392 & ~n_40393;
assign n_40395 =  x_3912 & ~n_23898;
assign n_40396 = ~n_23839 & ~n_23247;
assign n_40397 = ~n_40395 &  n_40396;
assign n_40398 =  x_3912 & ~n_40397;
assign n_40399 = ~x_3912 &  n_40397;
assign n_40400 = ~n_40398 & ~n_40399;
assign n_40401 = ~n_23898 & ~n_23247;
assign n_40402 =  x_3911 & ~n_23839;
assign n_40403 =  n_40401 & ~n_40402;
assign n_40404 =  x_3911 & ~n_40403;
assign n_40405 = ~x_3911 &  n_40403;
assign n_40406 = ~n_40404 & ~n_40405;
assign n_40407 = ~n_23839 &  n_40401;
assign n_40408 =  x_3910 &  n_40407;
assign n_40409 =  x_3910 &  n_40408;
assign n_40410 = ~x_3910 & ~n_40408;
assign n_40411 = ~n_40409 & ~n_40410;
assign n_40412 =  x_3909 &  n_40407;
assign n_40413 =  x_3909 &  n_40412;
assign n_40414 = ~x_3909 & ~n_40412;
assign n_40415 = ~n_40413 & ~n_40414;
assign n_40416 =  x_3908 &  n_40407;
assign n_40417 =  x_3908 &  n_40416;
assign n_40418 = ~x_3908 & ~n_40416;
assign n_40419 = ~n_40417 & ~n_40418;
assign n_40420 =  x_3907 &  n_40407;
assign n_40421 =  x_3907 &  n_40420;
assign n_40422 = ~x_3907 & ~n_40420;
assign n_40423 = ~n_40421 & ~n_40422;
assign n_40424 =  x_3906 &  n_40407;
assign n_40425 =  x_3906 &  n_40424;
assign n_40426 = ~x_3906 & ~n_40424;
assign n_40427 = ~n_40425 & ~n_40426;
assign n_40428 =  x_3905 &  n_40407;
assign n_40429 =  x_3905 &  n_40428;
assign n_40430 = ~x_3905 & ~n_40428;
assign n_40431 = ~n_40429 & ~n_40430;
assign n_40432 =  x_3904 &  n_40407;
assign n_40433 =  x_3904 &  n_40432;
assign n_40434 = ~x_3904 & ~n_40432;
assign n_40435 = ~n_40433 & ~n_40434;
assign n_40436 =  x_3903 &  n_40407;
assign n_40437 =  x_3903 &  n_40436;
assign n_40438 = ~x_3903 & ~n_40436;
assign n_40439 = ~n_40437 & ~n_40438;
assign n_40440 =  x_3902 &  n_40407;
assign n_40441 =  x_3902 &  n_40440;
assign n_40442 = ~x_3902 & ~n_40440;
assign n_40443 = ~n_40441 & ~n_40442;
assign n_40444 =  x_3901 &  n_40407;
assign n_40445 =  x_3901 &  n_40444;
assign n_40446 = ~x_3901 & ~n_40444;
assign n_40447 = ~n_40445 & ~n_40446;
assign n_40448 =  x_3900 &  n_40407;
assign n_40449 =  x_3900 &  n_40448;
assign n_40450 = ~x_3900 & ~n_40448;
assign n_40451 = ~n_40449 & ~n_40450;
assign n_40452 =  x_3899 &  n_40407;
assign n_40453 =  x_3899 &  n_40452;
assign n_40454 = ~x_3899 & ~n_40452;
assign n_40455 = ~n_40453 & ~n_40454;
assign n_40456 =  x_3898 &  n_40407;
assign n_40457 =  x_3898 &  n_40456;
assign n_40458 = ~x_3898 & ~n_40456;
assign n_40459 = ~n_40457 & ~n_40458;
assign n_40460 =  x_3897 &  n_40407;
assign n_40461 =  x_3897 &  n_40460;
assign n_40462 = ~x_3897 & ~n_40460;
assign n_40463 = ~n_40461 & ~n_40462;
assign n_40464 =  x_3896 &  n_40407;
assign n_40465 =  x_3896 &  n_40464;
assign n_40466 = ~x_3896 & ~n_40464;
assign n_40467 = ~n_40465 & ~n_40466;
assign n_40468 =  x_3895 & ~n_26301;
assign n_40469 =  x_2906 &  n_13142;
assign n_40470 = ~x_3064 &  n_13135;
assign n_40471 = ~n_13142 & ~n_40470;
assign n_40472 =  x_4775 & ~n_40471;
assign n_40473 = ~n_40469 &  n_40472;
assign n_40474 = ~n_13136 &  n_13147;
assign n_40475 = ~x_2842 &  n_13145;
assign n_40476 =  n_26301 & ~n_40475;
assign n_40477 = ~n_40474 &  n_40476;
assign n_40478 = ~n_40473 &  n_40477;
assign n_40479 = ~n_40468 & ~n_40478;
assign n_40480 =  x_3895 & ~n_40479;
assign n_40481 = ~x_3895 &  n_40479;
assign n_40482 = ~n_40480 & ~n_40481;
assign n_40483 =  x_3894 & ~n_26301;
assign n_40484 =  x_2905 &  n_13142;
assign n_40485 = ~x_3063 &  n_13135;
assign n_40486 = ~n_13142 & ~n_40485;
assign n_40487 =  x_4775 & ~n_40486;
assign n_40488 = ~n_40484 &  n_40487;
assign n_40489 = ~n_13136 &  n_13164;
assign n_40490 = ~x_2841 &  n_13145;
assign n_40491 =  n_26301 & ~n_40490;
assign n_40492 = ~n_40489 &  n_40491;
assign n_40493 = ~n_40488 &  n_40492;
assign n_40494 = ~n_40483 & ~n_40493;
assign n_40495 =  x_3894 & ~n_40494;
assign n_40496 = ~x_3894 &  n_40494;
assign n_40497 = ~n_40495 & ~n_40496;
assign n_40498 =  x_3893 & ~n_26301;
assign n_40499 =  x_2904 &  n_13142;
assign n_40500 = ~x_3062 &  n_13135;
assign n_40501 = ~n_13142 & ~n_40500;
assign n_40502 =  x_4775 & ~n_40501;
assign n_40503 = ~n_40499 &  n_40502;
assign n_40504 = ~n_13136 &  n_13181;
assign n_40505 = ~x_2840 &  n_13145;
assign n_40506 =  n_26301 & ~n_40505;
assign n_40507 = ~n_40504 &  n_40506;
assign n_40508 = ~n_40503 &  n_40507;
assign n_40509 = ~n_40498 & ~n_40508;
assign n_40510 =  x_3893 & ~n_40509;
assign n_40511 = ~x_3893 &  n_40509;
assign n_40512 = ~n_40510 & ~n_40511;
assign n_40513 =  x_3892 & ~n_26301;
assign n_40514 =  x_2903 &  n_13142;
assign n_40515 = ~x_3061 &  n_13135;
assign n_40516 = ~n_13142 & ~n_40515;
assign n_40517 =  x_4775 & ~n_40516;
assign n_40518 = ~n_40514 &  n_40517;
assign n_40519 = ~n_13136 &  n_13198;
assign n_40520 = ~x_2839 &  n_13145;
assign n_40521 =  n_26301 & ~n_40520;
assign n_40522 = ~n_40519 &  n_40521;
assign n_40523 = ~n_40518 &  n_40522;
assign n_40524 = ~n_40513 & ~n_40523;
assign n_40525 =  x_3892 & ~n_40524;
assign n_40526 = ~x_3892 &  n_40524;
assign n_40527 = ~n_40525 & ~n_40526;
assign n_40528 =  x_3891 & ~n_26301;
assign n_40529 =  x_2902 &  n_13142;
assign n_40530 = ~x_3060 &  n_13135;
assign n_40531 = ~n_13142 & ~n_40530;
assign n_40532 =  x_4775 & ~n_40531;
assign n_40533 = ~n_40529 &  n_40532;
assign n_40534 = ~n_13136 &  n_13215;
assign n_40535 = ~x_2838 &  n_13145;
assign n_40536 =  n_26301 & ~n_40535;
assign n_40537 = ~n_40534 &  n_40536;
assign n_40538 = ~n_40533 &  n_40537;
assign n_40539 = ~n_40528 & ~n_40538;
assign n_40540 =  x_3891 & ~n_40539;
assign n_40541 = ~x_3891 &  n_40539;
assign n_40542 = ~n_40540 & ~n_40541;
assign n_40543 =  x_3890 & ~n_26301;
assign n_40544 =  x_2901 &  n_13142;
assign n_40545 = ~x_3059 &  n_13135;
assign n_40546 = ~n_13142 & ~n_40545;
assign n_40547 =  x_4775 & ~n_40546;
assign n_40548 = ~n_40544 &  n_40547;
assign n_40549 = ~n_13136 &  n_29630;
assign n_40550 = ~x_2837 &  n_13145;
assign n_40551 =  n_26301 & ~n_40550;
assign n_40552 = ~n_40549 &  n_40551;
assign n_40553 = ~n_40548 &  n_40552;
assign n_40554 = ~n_40543 & ~n_40553;
assign n_40555 =  x_3890 & ~n_40554;
assign n_40556 = ~x_3890 &  n_40554;
assign n_40557 = ~n_40555 & ~n_40556;
assign n_40558 =  x_3889 & ~n_26301;
assign n_40559 =  x_2900 &  n_13142;
assign n_40560 = ~x_3058 &  n_13135;
assign n_40561 = ~n_13142 & ~n_40560;
assign n_40562 =  x_4775 & ~n_40561;
assign n_40563 = ~n_40559 &  n_40562;
assign n_40564 = ~n_13136 &  n_29647;
assign n_40565 = ~x_2836 &  n_13145;
assign n_40566 =  n_26301 & ~n_40565;
assign n_40567 = ~n_40564 &  n_40566;
assign n_40568 = ~n_40563 &  n_40567;
assign n_40569 = ~n_40558 & ~n_40568;
assign n_40570 =  x_3889 & ~n_40569;
assign n_40571 = ~x_3889 &  n_40569;
assign n_40572 = ~n_40570 & ~n_40571;
assign n_40573 =  x_3888 & ~n_26301;
assign n_40574 =  x_2899 &  n_13142;
assign n_40575 = ~x_3057 &  n_13135;
assign n_40576 = ~n_13142 & ~n_40575;
assign n_40577 =  x_4775 & ~n_40576;
assign n_40578 = ~n_40574 &  n_40577;
assign n_40579 = ~n_13136 &  n_29664;
assign n_40580 = ~x_2835 &  n_13145;
assign n_40581 =  n_26301 & ~n_40580;
assign n_40582 = ~n_40579 &  n_40581;
assign n_40583 = ~n_40578 &  n_40582;
assign n_40584 = ~n_40573 & ~n_40583;
assign n_40585 =  x_3888 & ~n_40584;
assign n_40586 = ~x_3888 &  n_40584;
assign n_40587 = ~n_40585 & ~n_40586;
assign n_40588 =  x_3887 & ~n_26301;
assign n_40589 =  x_2898 &  n_13142;
assign n_40590 = ~x_3056 &  n_13135;
assign n_40591 = ~n_13142 & ~n_40590;
assign n_40592 =  x_4775 & ~n_40591;
assign n_40593 = ~n_40589 &  n_40592;
assign n_40594 = ~n_13136 &  n_29681;
assign n_40595 = ~x_2834 &  n_13145;
assign n_40596 =  n_26301 & ~n_40595;
assign n_40597 = ~n_40594 &  n_40596;
assign n_40598 = ~n_40593 &  n_40597;
assign n_40599 = ~n_40588 & ~n_40598;
assign n_40600 =  x_3887 & ~n_40599;
assign n_40601 = ~x_3887 &  n_40599;
assign n_40602 = ~n_40600 & ~n_40601;
assign n_40603 =  x_3886 & ~n_26301;
assign n_40604 =  x_2897 &  n_13142;
assign n_40605 = ~x_3055 &  n_13135;
assign n_40606 = ~n_13142 & ~n_40605;
assign n_40607 =  x_4775 & ~n_40606;
assign n_40608 = ~n_40604 &  n_40607;
assign n_40609 = ~n_13136 &  n_29698;
assign n_40610 = ~x_2833 &  n_13145;
assign n_40611 =  n_26301 & ~n_40610;
assign n_40612 = ~n_40609 &  n_40611;
assign n_40613 = ~n_40608 &  n_40612;
assign n_40614 = ~n_40603 & ~n_40613;
assign n_40615 =  x_3886 & ~n_40614;
assign n_40616 = ~x_3886 &  n_40614;
assign n_40617 = ~n_40615 & ~n_40616;
assign n_40618 =  x_3885 & ~n_26301;
assign n_40619 =  x_2896 &  n_13142;
assign n_40620 = ~x_3054 &  n_13135;
assign n_40621 = ~n_13142 & ~n_40620;
assign n_40622 =  x_4775 & ~n_40621;
assign n_40623 = ~n_40619 &  n_40622;
assign n_40624 = ~n_13136 &  n_29715;
assign n_40625 = ~x_2832 &  n_13145;
assign n_40626 =  n_26301 & ~n_40625;
assign n_40627 = ~n_40624 &  n_40626;
assign n_40628 = ~n_40623 &  n_40627;
assign n_40629 = ~n_40618 & ~n_40628;
assign n_40630 =  x_3885 & ~n_40629;
assign n_40631 = ~x_3885 &  n_40629;
assign n_40632 = ~n_40630 & ~n_40631;
assign n_40633 =  x_3884 & ~n_26301;
assign n_40634 =  x_2895 &  n_13142;
assign n_40635 = ~x_3053 &  n_13135;
assign n_40636 = ~n_13142 & ~n_40635;
assign n_40637 =  x_4775 & ~n_40636;
assign n_40638 = ~n_40634 &  n_40637;
assign n_40639 = ~n_13136 &  n_29732;
assign n_40640 = ~x_2831 &  n_13145;
assign n_40641 =  n_26301 & ~n_40640;
assign n_40642 = ~n_40639 &  n_40641;
assign n_40643 = ~n_40638 &  n_40642;
assign n_40644 = ~n_40633 & ~n_40643;
assign n_40645 =  x_3884 & ~n_40644;
assign n_40646 = ~x_3884 &  n_40644;
assign n_40647 = ~n_40645 & ~n_40646;
assign n_40648 =  x_3883 & ~n_26301;
assign n_40649 =  x_2894 &  n_13142;
assign n_40650 = ~x_3052 &  n_13135;
assign n_40651 = ~n_13142 & ~n_40650;
assign n_40652 =  x_4775 & ~n_40651;
assign n_40653 = ~n_40649 &  n_40652;
assign n_40654 = ~n_13136 &  n_29749;
assign n_40655 = ~x_2830 &  n_13145;
assign n_40656 =  n_26301 & ~n_40655;
assign n_40657 = ~n_40654 &  n_40656;
assign n_40658 = ~n_40653 &  n_40657;
assign n_40659 = ~n_40648 & ~n_40658;
assign n_40660 =  x_3883 & ~n_40659;
assign n_40661 = ~x_3883 &  n_40659;
assign n_40662 = ~n_40660 & ~n_40661;
assign n_40663 =  x_3882 & ~n_26301;
assign n_40664 =  x_2893 &  n_13142;
assign n_40665 = ~x_3051 &  n_13135;
assign n_40666 = ~n_13142 & ~n_40665;
assign n_40667 =  x_4775 & ~n_40666;
assign n_40668 = ~n_40664 &  n_40667;
assign n_40669 = ~n_13136 &  n_29766;
assign n_40670 = ~x_2829 &  n_13145;
assign n_40671 =  n_26301 & ~n_40670;
assign n_40672 = ~n_40669 &  n_40671;
assign n_40673 = ~n_40668 &  n_40672;
assign n_40674 = ~n_40663 & ~n_40673;
assign n_40675 =  x_3882 & ~n_40674;
assign n_40676 = ~x_3882 &  n_40674;
assign n_40677 = ~n_40675 & ~n_40676;
assign n_40678 =  x_3881 & ~n_26301;
assign n_40679 =  x_2892 &  n_13142;
assign n_40680 = ~x_3050 &  n_13135;
assign n_40681 = ~n_13142 & ~n_40680;
assign n_40682 =  x_4775 & ~n_40681;
assign n_40683 = ~n_40679 &  n_40682;
assign n_40684 = ~n_13136 &  n_29783;
assign n_40685 = ~x_2828 &  n_13145;
assign n_40686 =  n_26301 & ~n_40685;
assign n_40687 = ~n_40684 &  n_40686;
assign n_40688 = ~n_40683 &  n_40687;
assign n_40689 = ~n_40678 & ~n_40688;
assign n_40690 =  x_3881 & ~n_40689;
assign n_40691 = ~x_3881 &  n_40689;
assign n_40692 = ~n_40690 & ~n_40691;
assign n_40693 =  x_3880 & ~n_26301;
assign n_40694 =  x_2891 &  n_13142;
assign n_40695 = ~x_3049 &  n_13135;
assign n_40696 = ~n_13142 & ~n_40695;
assign n_40697 =  x_4775 & ~n_40696;
assign n_40698 = ~n_40694 &  n_40697;
assign n_40699 = ~n_13136 &  n_29800;
assign n_40700 = ~x_2827 &  n_13145;
assign n_40701 =  n_26301 & ~n_40700;
assign n_40702 = ~n_40699 &  n_40701;
assign n_40703 = ~n_40698 &  n_40702;
assign n_40704 = ~n_40693 & ~n_40703;
assign n_40705 =  x_3880 & ~n_40704;
assign n_40706 = ~x_3880 &  n_40704;
assign n_40707 = ~n_40705 & ~n_40706;
assign n_40708 =  x_3879 & ~n_26301;
assign n_40709 =  x_2890 &  n_13142;
assign n_40710 = ~x_3048 &  n_13135;
assign n_40711 = ~n_13142 & ~n_40710;
assign n_40712 =  x_4775 & ~n_40711;
assign n_40713 = ~n_40709 &  n_40712;
assign n_40714 = ~n_13136 &  n_29817;
assign n_40715 = ~x_2826 &  n_13145;
assign n_40716 =  n_26301 & ~n_40715;
assign n_40717 = ~n_40714 &  n_40716;
assign n_40718 = ~n_40713 &  n_40717;
assign n_40719 = ~n_40708 & ~n_40718;
assign n_40720 =  x_3879 & ~n_40719;
assign n_40721 = ~x_3879 &  n_40719;
assign n_40722 = ~n_40720 & ~n_40721;
assign n_40723 =  x_3878 & ~n_26301;
assign n_40724 =  x_2889 &  n_13142;
assign n_40725 = ~x_3047 &  n_13135;
assign n_40726 = ~n_13142 & ~n_40725;
assign n_40727 =  x_4775 & ~n_40726;
assign n_40728 = ~n_40724 &  n_40727;
assign n_40729 = ~n_13136 &  n_29834;
assign n_40730 = ~x_2825 &  n_13145;
assign n_40731 =  n_26301 & ~n_40730;
assign n_40732 = ~n_40729 &  n_40731;
assign n_40733 = ~n_40728 &  n_40732;
assign n_40734 = ~n_40723 & ~n_40733;
assign n_40735 =  x_3878 & ~n_40734;
assign n_40736 = ~x_3878 &  n_40734;
assign n_40737 = ~n_40735 & ~n_40736;
assign n_40738 =  x_3877 & ~n_26301;
assign n_40739 =  x_2888 &  n_13142;
assign n_40740 = ~x_3046 &  n_13135;
assign n_40741 = ~n_13142 & ~n_40740;
assign n_40742 =  x_4775 & ~n_40741;
assign n_40743 = ~n_40739 &  n_40742;
assign n_40744 = ~n_13136 &  n_29851;
assign n_40745 = ~x_2824 &  n_13145;
assign n_40746 =  n_26301 & ~n_40745;
assign n_40747 = ~n_40744 &  n_40746;
assign n_40748 = ~n_40743 &  n_40747;
assign n_40749 = ~n_40738 & ~n_40748;
assign n_40750 =  x_3877 & ~n_40749;
assign n_40751 = ~x_3877 &  n_40749;
assign n_40752 = ~n_40750 & ~n_40751;
assign n_40753 =  x_3876 & ~n_26301;
assign n_40754 =  x_2887 &  n_13142;
assign n_40755 = ~x_3045 &  n_13135;
assign n_40756 = ~n_13142 & ~n_40755;
assign n_40757 =  x_4775 & ~n_40756;
assign n_40758 = ~n_40754 &  n_40757;
assign n_40759 = ~n_13136 &  n_29868;
assign n_40760 = ~x_2823 &  n_13145;
assign n_40761 =  n_26301 & ~n_40760;
assign n_40762 = ~n_40759 &  n_40761;
assign n_40763 = ~n_40758 &  n_40762;
assign n_40764 = ~n_40753 & ~n_40763;
assign n_40765 =  x_3876 & ~n_40764;
assign n_40766 = ~x_3876 &  n_40764;
assign n_40767 = ~n_40765 & ~n_40766;
assign n_40768 =  x_3875 & ~n_26301;
assign n_40769 =  x_2886 &  n_13142;
assign n_40770 = ~x_3044 &  n_13135;
assign n_40771 = ~n_13142 & ~n_40770;
assign n_40772 =  x_4775 & ~n_40771;
assign n_40773 = ~n_40769 &  n_40772;
assign n_40774 = ~n_13136 &  n_29885;
assign n_40775 = ~x_2822 &  n_13145;
assign n_40776 =  n_26301 & ~n_40775;
assign n_40777 = ~n_40774 &  n_40776;
assign n_40778 = ~n_40773 &  n_40777;
assign n_40779 = ~n_40768 & ~n_40778;
assign n_40780 =  x_3875 & ~n_40779;
assign n_40781 = ~x_3875 &  n_40779;
assign n_40782 = ~n_40780 & ~n_40781;
assign n_40783 =  x_3874 & ~n_26301;
assign n_40784 =  x_2885 &  n_13142;
assign n_40785 = ~x_3043 &  n_13135;
assign n_40786 = ~n_13142 & ~n_40785;
assign n_40787 =  x_4775 & ~n_40786;
assign n_40788 = ~n_40784 &  n_40787;
assign n_40789 = ~n_13136 &  n_29902;
assign n_40790 = ~x_2821 &  n_13145;
assign n_40791 =  n_26301 & ~n_40790;
assign n_40792 = ~n_40789 &  n_40791;
assign n_40793 = ~n_40788 &  n_40792;
assign n_40794 = ~n_40783 & ~n_40793;
assign n_40795 =  x_3874 & ~n_40794;
assign n_40796 = ~x_3874 &  n_40794;
assign n_40797 = ~n_40795 & ~n_40796;
assign n_40798 =  x_3873 & ~n_26301;
assign n_40799 =  x_2884 &  n_13142;
assign n_40800 = ~x_3042 &  n_13135;
assign n_40801 = ~n_13142 & ~n_40800;
assign n_40802 =  x_4775 & ~n_40801;
assign n_40803 = ~n_40799 &  n_40802;
assign n_40804 = ~n_13136 &  n_29919;
assign n_40805 = ~x_2820 &  n_13145;
assign n_40806 =  n_26301 & ~n_40805;
assign n_40807 = ~n_40804 &  n_40806;
assign n_40808 = ~n_40803 &  n_40807;
assign n_40809 = ~n_40798 & ~n_40808;
assign n_40810 =  x_3873 & ~n_40809;
assign n_40811 = ~x_3873 &  n_40809;
assign n_40812 = ~n_40810 & ~n_40811;
assign n_40813 =  x_3872 & ~n_26301;
assign n_40814 =  x_2883 &  n_13142;
assign n_40815 = ~x_3041 &  n_13135;
assign n_40816 = ~n_13142 & ~n_40815;
assign n_40817 =  x_4775 & ~n_40816;
assign n_40818 = ~n_40814 &  n_40817;
assign n_40819 = ~n_13136 &  n_29936;
assign n_40820 = ~x_2819 &  n_13145;
assign n_40821 =  n_26301 & ~n_40820;
assign n_40822 = ~n_40819 &  n_40821;
assign n_40823 = ~n_40818 &  n_40822;
assign n_40824 = ~n_40813 & ~n_40823;
assign n_40825 =  x_3872 & ~n_40824;
assign n_40826 = ~x_3872 &  n_40824;
assign n_40827 = ~n_40825 & ~n_40826;
assign n_40828 =  x_3871 & ~n_26301;
assign n_40829 =  x_2882 &  n_13142;
assign n_40830 = ~x_3040 &  n_13135;
assign n_40831 = ~n_13142 & ~n_40830;
assign n_40832 =  x_4775 & ~n_40831;
assign n_40833 = ~n_40829 &  n_40832;
assign n_40834 = ~n_13136 &  n_29953;
assign n_40835 = ~x_2818 &  n_13145;
assign n_40836 =  n_26301 & ~n_40835;
assign n_40837 = ~n_40834 &  n_40836;
assign n_40838 = ~n_40833 &  n_40837;
assign n_40839 = ~n_40828 & ~n_40838;
assign n_40840 =  x_3871 & ~n_40839;
assign n_40841 = ~x_3871 &  n_40839;
assign n_40842 = ~n_40840 & ~n_40841;
assign n_40843 =  x_3870 & ~n_26301;
assign n_40844 =  x_2881 &  n_13142;
assign n_40845 = ~x_3039 &  n_13135;
assign n_40846 = ~n_13142 & ~n_40845;
assign n_40847 =  x_4775 & ~n_40846;
assign n_40848 = ~n_40844 &  n_40847;
assign n_40849 = ~n_13136 &  n_29970;
assign n_40850 = ~x_2817 &  n_13145;
assign n_40851 =  n_26301 & ~n_40850;
assign n_40852 = ~n_40849 &  n_40851;
assign n_40853 = ~n_40848 &  n_40852;
assign n_40854 = ~n_40843 & ~n_40853;
assign n_40855 =  x_3870 & ~n_40854;
assign n_40856 = ~x_3870 &  n_40854;
assign n_40857 = ~n_40855 & ~n_40856;
assign n_40858 =  x_3869 & ~n_26301;
assign n_40859 =  x_2880 &  n_13142;
assign n_40860 = ~x_3038 &  n_13135;
assign n_40861 = ~n_13142 & ~n_40860;
assign n_40862 =  x_4775 & ~n_40861;
assign n_40863 = ~n_40859 &  n_40862;
assign n_40864 = ~n_13136 &  n_29987;
assign n_40865 = ~x_2816 &  n_13145;
assign n_40866 =  n_26301 & ~n_40865;
assign n_40867 = ~n_40864 &  n_40866;
assign n_40868 = ~n_40863 &  n_40867;
assign n_40869 = ~n_40858 & ~n_40868;
assign n_40870 =  x_3869 & ~n_40869;
assign n_40871 = ~x_3869 &  n_40869;
assign n_40872 = ~n_40870 & ~n_40871;
assign n_40873 =  x_3868 & ~n_26301;
assign n_40874 =  x_2879 &  n_13142;
assign n_40875 = ~x_3037 &  n_13135;
assign n_40876 = ~n_13142 & ~n_40875;
assign n_40877 =  x_4775 & ~n_40876;
assign n_40878 = ~n_40874 &  n_40877;
assign n_40879 = ~n_13136 &  n_30004;
assign n_40880 = ~x_2815 &  n_13145;
assign n_40881 =  n_26301 & ~n_40880;
assign n_40882 = ~n_40879 &  n_40881;
assign n_40883 = ~n_40878 &  n_40882;
assign n_40884 = ~n_40873 & ~n_40883;
assign n_40885 =  x_3868 & ~n_40884;
assign n_40886 = ~x_3868 &  n_40884;
assign n_40887 = ~n_40885 & ~n_40886;
assign n_40888 =  x_3867 & ~n_26301;
assign n_40889 =  x_2878 &  n_13142;
assign n_40890 = ~x_3036 &  n_13135;
assign n_40891 = ~n_13142 & ~n_40890;
assign n_40892 =  x_4775 & ~n_40891;
assign n_40893 = ~n_40889 &  n_40892;
assign n_40894 = ~n_13136 &  n_30021;
assign n_40895 = ~x_2814 &  n_13145;
assign n_40896 =  n_26301 & ~n_40895;
assign n_40897 = ~n_40894 &  n_40896;
assign n_40898 = ~n_40893 &  n_40897;
assign n_40899 = ~n_40888 & ~n_40898;
assign n_40900 =  x_3867 & ~n_40899;
assign n_40901 = ~x_3867 &  n_40899;
assign n_40902 = ~n_40900 & ~n_40901;
assign n_40903 =  x_3866 & ~n_26301;
assign n_40904 =  x_2877 &  n_13142;
assign n_40905 = ~x_3035 &  n_13135;
assign n_40906 = ~n_13142 & ~n_40905;
assign n_40907 =  x_4775 & ~n_40906;
assign n_40908 = ~n_40904 &  n_40907;
assign n_40909 = ~n_13136 &  n_30038;
assign n_40910 = ~x_2813 &  n_13145;
assign n_40911 =  n_26301 & ~n_40910;
assign n_40912 = ~n_40909 &  n_40911;
assign n_40913 = ~n_40908 &  n_40912;
assign n_40914 = ~n_40903 & ~n_40913;
assign n_40915 =  x_3866 & ~n_40914;
assign n_40916 = ~x_3866 &  n_40914;
assign n_40917 = ~n_40915 & ~n_40916;
assign n_40918 =  x_3865 & ~n_26301;
assign n_40919 =  x_2876 &  n_13142;
assign n_40920 = ~x_3034 &  n_13135;
assign n_40921 = ~n_13142 & ~n_40920;
assign n_40922 =  x_4775 & ~n_40921;
assign n_40923 = ~n_40919 &  n_40922;
assign n_40924 = ~n_13136 &  n_30055;
assign n_40925 = ~x_2812 &  n_13145;
assign n_40926 =  n_26301 & ~n_40925;
assign n_40927 = ~n_40924 &  n_40926;
assign n_40928 = ~n_40923 &  n_40927;
assign n_40929 = ~n_40918 & ~n_40928;
assign n_40930 =  x_3865 & ~n_40929;
assign n_40931 = ~x_3865 &  n_40929;
assign n_40932 = ~n_40930 & ~n_40931;
assign n_40933 =  x_3864 & ~n_26301;
assign n_40934 =  i_1 & ~n_13136;
assign n_40935 =  x_3033 &  n_13136;
assign n_40936 = ~n_13142 & ~n_40935;
assign n_40937 = ~n_40934 &  n_40936;
assign n_40938 = ~x_2811 & ~x_4775;
assign n_40939 = ~n_15903 & ~n_40938;
assign n_40940 =  n_13142 & ~n_40939;
assign n_40941 =  n_26301 & ~n_40940;
assign n_40942 = ~n_40937 &  n_40941;
assign n_40943 = ~n_40933 & ~n_40942;
assign n_40944 =  x_3864 & ~n_40943;
assign n_40945 = ~x_3864 &  n_40943;
assign n_40946 = ~n_40944 & ~n_40945;
assign n_40947 =  n_25230 & ~n_36595;
assign n_40948 =  x_3863 & ~n_25230;
assign n_40949 = ~n_40947 & ~n_40948;
assign n_40950 =  x_3863 & ~n_40949;
assign n_40951 = ~x_3863 &  n_40949;
assign n_40952 = ~n_40950 & ~n_40951;
assign n_40953 =  n_25230 & ~n_36610;
assign n_40954 =  x_3862 & ~n_25230;
assign n_40955 = ~n_40953 & ~n_40954;
assign n_40956 =  x_3862 & ~n_40955;
assign n_40957 = ~x_3862 &  n_40955;
assign n_40958 = ~n_40956 & ~n_40957;
assign n_40959 =  n_25230 & ~n_36625;
assign n_40960 =  x_3861 & ~n_25230;
assign n_40961 = ~n_40959 & ~n_40960;
assign n_40962 =  x_3861 & ~n_40961;
assign n_40963 = ~x_3861 &  n_40961;
assign n_40964 = ~n_40962 & ~n_40963;
assign n_40965 =  n_25230 & ~n_36640;
assign n_40966 =  x_3860 & ~n_25230;
assign n_40967 = ~n_40965 & ~n_40966;
assign n_40968 =  x_3860 & ~n_40967;
assign n_40969 = ~x_3860 &  n_40967;
assign n_40970 = ~n_40968 & ~n_40969;
assign n_40971 =  n_25230 & ~n_36655;
assign n_40972 =  x_3859 & ~n_25230;
assign n_40973 = ~n_40971 & ~n_40972;
assign n_40974 =  x_3859 & ~n_40973;
assign n_40975 = ~x_3859 &  n_40973;
assign n_40976 = ~n_40974 & ~n_40975;
assign n_40977 =  n_25230 & ~n_36670;
assign n_40978 =  x_3858 & ~n_25230;
assign n_40979 = ~n_40977 & ~n_40978;
assign n_40980 =  x_3858 & ~n_40979;
assign n_40981 = ~x_3858 &  n_40979;
assign n_40982 = ~n_40980 & ~n_40981;
assign n_40983 =  n_25230 & ~n_36685;
assign n_40984 =  x_3857 & ~n_25230;
assign n_40985 = ~n_40983 & ~n_40984;
assign n_40986 =  x_3857 & ~n_40985;
assign n_40987 = ~x_3857 &  n_40985;
assign n_40988 = ~n_40986 & ~n_40987;
assign n_40989 =  n_25230 & ~n_36700;
assign n_40990 =  x_3856 & ~n_25230;
assign n_40991 = ~n_40989 & ~n_40990;
assign n_40992 =  x_3856 & ~n_40991;
assign n_40993 = ~x_3856 &  n_40991;
assign n_40994 = ~n_40992 & ~n_40993;
assign n_40995 =  n_25230 & ~n_36715;
assign n_40996 =  x_3855 & ~n_25230;
assign n_40997 = ~n_40995 & ~n_40996;
assign n_40998 =  x_3855 & ~n_40997;
assign n_40999 = ~x_3855 &  n_40997;
assign n_41000 = ~n_40998 & ~n_40999;
assign n_41001 =  n_25230 & ~n_36730;
assign n_41002 =  x_3854 & ~n_25230;
assign n_41003 = ~n_41001 & ~n_41002;
assign n_41004 =  x_3854 & ~n_41003;
assign n_41005 = ~x_3854 &  n_41003;
assign n_41006 = ~n_41004 & ~n_41005;
assign n_41007 =  n_25230 & ~n_36745;
assign n_41008 =  x_3853 & ~n_25230;
assign n_41009 = ~n_41007 & ~n_41008;
assign n_41010 =  x_3853 & ~n_41009;
assign n_41011 = ~x_3853 &  n_41009;
assign n_41012 = ~n_41010 & ~n_41011;
assign n_41013 =  n_25230 & ~n_36760;
assign n_41014 =  x_3852 & ~n_25230;
assign n_41015 = ~n_41013 & ~n_41014;
assign n_41016 =  x_3852 & ~n_41015;
assign n_41017 = ~x_3852 &  n_41015;
assign n_41018 = ~n_41016 & ~n_41017;
assign n_41019 =  n_25230 & ~n_36775;
assign n_41020 =  x_3851 & ~n_25230;
assign n_41021 = ~n_41019 & ~n_41020;
assign n_41022 =  x_3851 & ~n_41021;
assign n_41023 = ~x_3851 &  n_41021;
assign n_41024 = ~n_41022 & ~n_41023;
assign n_41025 =  n_25230 & ~n_36790;
assign n_41026 =  x_3850 & ~n_25230;
assign n_41027 = ~n_41025 & ~n_41026;
assign n_41028 =  x_3850 & ~n_41027;
assign n_41029 = ~x_3850 &  n_41027;
assign n_41030 = ~n_41028 & ~n_41029;
assign n_41031 =  n_25230 & ~n_36805;
assign n_41032 =  x_3849 & ~n_25230;
assign n_41033 = ~n_41031 & ~n_41032;
assign n_41034 =  x_3849 & ~n_41033;
assign n_41035 = ~x_3849 &  n_41033;
assign n_41036 = ~n_41034 & ~n_41035;
assign n_41037 =  n_25230 & ~n_36820;
assign n_41038 =  x_3848 & ~n_25230;
assign n_41039 = ~n_41037 & ~n_41038;
assign n_41040 =  x_3848 & ~n_41039;
assign n_41041 = ~x_3848 &  n_41039;
assign n_41042 = ~n_41040 & ~n_41041;
assign n_41043 =  n_25230 & ~n_36835;
assign n_41044 =  x_3847 & ~n_25230;
assign n_41045 = ~n_41043 & ~n_41044;
assign n_41046 =  x_3847 & ~n_41045;
assign n_41047 = ~x_3847 &  n_41045;
assign n_41048 = ~n_41046 & ~n_41047;
assign n_41049 =  n_25230 & ~n_36850;
assign n_41050 =  x_3846 & ~n_25230;
assign n_41051 = ~n_41049 & ~n_41050;
assign n_41052 =  x_3846 & ~n_41051;
assign n_41053 = ~x_3846 &  n_41051;
assign n_41054 = ~n_41052 & ~n_41053;
assign n_41055 =  n_25230 & ~n_36865;
assign n_41056 =  x_3845 & ~n_25230;
assign n_41057 = ~n_41055 & ~n_41056;
assign n_41058 =  x_3845 & ~n_41057;
assign n_41059 = ~x_3845 &  n_41057;
assign n_41060 = ~n_41058 & ~n_41059;
assign n_41061 =  n_25230 & ~n_36880;
assign n_41062 =  x_3844 & ~n_25230;
assign n_41063 = ~n_41061 & ~n_41062;
assign n_41064 =  x_3844 & ~n_41063;
assign n_41065 = ~x_3844 &  n_41063;
assign n_41066 = ~n_41064 & ~n_41065;
assign n_41067 =  n_25230 & ~n_36895;
assign n_41068 =  x_3843 & ~n_25230;
assign n_41069 = ~n_41067 & ~n_41068;
assign n_41070 =  x_3843 & ~n_41069;
assign n_41071 = ~x_3843 &  n_41069;
assign n_41072 = ~n_41070 & ~n_41071;
assign n_41073 =  n_25230 & ~n_36910;
assign n_41074 =  x_3842 & ~n_25230;
assign n_41075 = ~n_41073 & ~n_41074;
assign n_41076 =  x_3842 & ~n_41075;
assign n_41077 = ~x_3842 &  n_41075;
assign n_41078 = ~n_41076 & ~n_41077;
assign n_41079 =  n_25230 & ~n_36925;
assign n_41080 =  x_3841 & ~n_25230;
assign n_41081 = ~n_41079 & ~n_41080;
assign n_41082 =  x_3841 & ~n_41081;
assign n_41083 = ~x_3841 &  n_41081;
assign n_41084 = ~n_41082 & ~n_41083;
assign n_41085 =  n_25230 & ~n_36940;
assign n_41086 =  x_3840 & ~n_25230;
assign n_41087 = ~n_41085 & ~n_41086;
assign n_41088 =  x_3840 & ~n_41087;
assign n_41089 = ~x_3840 &  n_41087;
assign n_41090 = ~n_41088 & ~n_41089;
assign n_41091 =  n_25230 & ~n_36955;
assign n_41092 =  x_3839 & ~n_25230;
assign n_41093 = ~n_41091 & ~n_41092;
assign n_41094 =  x_3839 & ~n_41093;
assign n_41095 = ~x_3839 &  n_41093;
assign n_41096 = ~n_41094 & ~n_41095;
assign n_41097 =  n_25230 & ~n_36970;
assign n_41098 =  x_3838 & ~n_25230;
assign n_41099 = ~n_41097 & ~n_41098;
assign n_41100 =  x_3838 & ~n_41099;
assign n_41101 = ~x_3838 &  n_41099;
assign n_41102 = ~n_41100 & ~n_41101;
assign n_41103 =  n_25230 & ~n_36985;
assign n_41104 =  x_3837 & ~n_25230;
assign n_41105 = ~n_41103 & ~n_41104;
assign n_41106 =  x_3837 & ~n_41105;
assign n_41107 = ~x_3837 &  n_41105;
assign n_41108 = ~n_41106 & ~n_41107;
assign n_41109 =  n_25230 & ~n_37000;
assign n_41110 =  x_3836 & ~n_25230;
assign n_41111 = ~n_41109 & ~n_41110;
assign n_41112 =  x_3836 & ~n_41111;
assign n_41113 = ~x_3836 &  n_41111;
assign n_41114 = ~n_41112 & ~n_41113;
assign n_41115 =  n_25230 & ~n_37015;
assign n_41116 =  x_3835 & ~n_25230;
assign n_41117 = ~n_41115 & ~n_41116;
assign n_41118 =  x_3835 & ~n_41117;
assign n_41119 = ~x_3835 &  n_41117;
assign n_41120 = ~n_41118 & ~n_41119;
assign n_41121 =  n_25230 & ~n_37030;
assign n_41122 =  x_3834 & ~n_25230;
assign n_41123 = ~n_41121 & ~n_41122;
assign n_41124 =  x_3834 & ~n_41123;
assign n_41125 = ~x_3834 &  n_41123;
assign n_41126 = ~n_41124 & ~n_41125;
assign n_41127 =  n_25230 & ~n_37045;
assign n_41128 =  x_3833 & ~n_25230;
assign n_41129 = ~n_41127 & ~n_41128;
assign n_41130 =  x_3833 & ~n_41129;
assign n_41131 = ~x_3833 &  n_41129;
assign n_41132 = ~n_41130 & ~n_41131;
assign n_41133 =  n_25230 & ~n_37060;
assign n_41134 =  x_3832 & ~n_25230;
assign n_41135 = ~n_41133 & ~n_41134;
assign n_41136 =  x_3832 & ~n_41135;
assign n_41137 = ~x_3832 &  n_41135;
assign n_41138 = ~n_41136 & ~n_41137;
assign n_41139 =  x_3831 & ~n_26992;
assign n_41140 =  x_3831 &  n_41139;
assign n_41141 = ~x_3831 & ~n_41139;
assign n_41142 = ~n_41140 & ~n_41141;
assign n_41143 =  x_3830 & ~n_26992;
assign n_41144 =  x_3830 &  n_41143;
assign n_41145 = ~x_3830 & ~n_41143;
assign n_41146 = ~n_41144 & ~n_41145;
assign n_41147 =  x_3829 & ~n_26992;
assign n_41148 =  x_3829 &  n_41147;
assign n_41149 = ~x_3829 & ~n_41147;
assign n_41150 = ~n_41148 & ~n_41149;
assign n_41151 =  x_3828 & ~n_26992;
assign n_41152 =  x_3828 &  n_41151;
assign n_41153 = ~x_3828 & ~n_41151;
assign n_41154 = ~n_41152 & ~n_41153;
assign n_41155 =  x_3827 & ~n_26992;
assign n_41156 =  x_3827 &  n_41155;
assign n_41157 = ~x_3827 & ~n_41155;
assign n_41158 = ~n_41156 & ~n_41157;
assign n_41159 =  x_3826 & ~n_26992;
assign n_41160 =  x_3826 &  n_41159;
assign n_41161 = ~x_3826 & ~n_41159;
assign n_41162 = ~n_41160 & ~n_41161;
assign n_41163 =  x_3825 & ~n_26992;
assign n_41164 =  x_3825 &  n_41163;
assign n_41165 = ~x_3825 & ~n_41163;
assign n_41166 = ~n_41164 & ~n_41165;
assign n_41167 =  x_3824 & ~n_26992;
assign n_41168 =  x_3824 &  n_41167;
assign n_41169 = ~x_3824 & ~n_41167;
assign n_41170 = ~n_41168 & ~n_41169;
assign n_41171 =  x_3823 & ~n_26992;
assign n_41172 =  x_3823 &  n_41171;
assign n_41173 = ~x_3823 & ~n_41171;
assign n_41174 = ~n_41172 & ~n_41173;
assign n_41175 =  x_3822 & ~n_26992;
assign n_41176 =  x_3822 &  n_41175;
assign n_41177 = ~x_3822 & ~n_41175;
assign n_41178 = ~n_41176 & ~n_41177;
assign n_41179 =  x_3821 & ~n_26992;
assign n_41180 =  x_3821 &  n_41179;
assign n_41181 = ~x_3821 & ~n_41179;
assign n_41182 = ~n_41180 & ~n_41181;
assign n_41183 =  x_3820 & ~n_26992;
assign n_41184 =  x_3820 &  n_41183;
assign n_41185 = ~x_3820 & ~n_41183;
assign n_41186 = ~n_41184 & ~n_41185;
assign n_41187 =  x_3819 & ~n_26992;
assign n_41188 =  x_3819 &  n_41187;
assign n_41189 = ~x_3819 & ~n_41187;
assign n_41190 = ~n_41188 & ~n_41189;
assign n_41191 =  x_3818 & ~n_26992;
assign n_41192 =  x_3818 &  n_41191;
assign n_41193 = ~x_3818 & ~n_41191;
assign n_41194 = ~n_41192 & ~n_41193;
assign n_41195 =  x_3817 & ~n_26992;
assign n_41196 =  x_3817 &  n_41195;
assign n_41197 = ~x_3817 & ~n_41195;
assign n_41198 = ~n_41196 & ~n_41197;
assign n_41199 =  x_3816 & ~n_26992;
assign n_41200 =  x_3816 &  n_41199;
assign n_41201 = ~x_3816 & ~n_41199;
assign n_41202 = ~n_41200 & ~n_41201;
assign n_41203 =  x_3815 & ~n_26992;
assign n_41204 =  x_3815 &  n_41203;
assign n_41205 = ~x_3815 & ~n_41203;
assign n_41206 = ~n_41204 & ~n_41205;
assign n_41207 =  x_3814 & ~n_26992;
assign n_41208 =  x_3814 &  n_41207;
assign n_41209 = ~x_3814 & ~n_41207;
assign n_41210 = ~n_41208 & ~n_41209;
assign n_41211 =  x_3813 & ~n_26992;
assign n_41212 =  x_3813 &  n_41211;
assign n_41213 = ~x_3813 & ~n_41211;
assign n_41214 = ~n_41212 & ~n_41213;
assign n_41215 =  x_3812 & ~n_26992;
assign n_41216 =  x_3812 &  n_41215;
assign n_41217 = ~x_3812 & ~n_41215;
assign n_41218 = ~n_41216 & ~n_41217;
assign n_41219 =  x_3811 & ~n_26992;
assign n_41220 =  x_3811 &  n_41219;
assign n_41221 = ~x_3811 & ~n_41219;
assign n_41222 = ~n_41220 & ~n_41221;
assign n_41223 =  x_3810 & ~n_26992;
assign n_41224 =  x_3810 &  n_41223;
assign n_41225 = ~x_3810 & ~n_41223;
assign n_41226 = ~n_41224 & ~n_41225;
assign n_41227 =  x_3809 & ~n_26992;
assign n_41228 =  x_3809 &  n_41227;
assign n_41229 = ~x_3809 & ~n_41227;
assign n_41230 = ~n_41228 & ~n_41229;
assign n_41231 =  x_3808 & ~n_26992;
assign n_41232 =  x_3808 &  n_41231;
assign n_41233 = ~x_3808 & ~n_41231;
assign n_41234 = ~n_41232 & ~n_41233;
assign n_41235 =  x_3807 & ~n_26992;
assign n_41236 =  x_3807 &  n_41235;
assign n_41237 = ~x_3807 & ~n_41235;
assign n_41238 = ~n_41236 & ~n_41237;
assign n_41239 =  x_3806 & ~n_26992;
assign n_41240 =  x_3806 &  n_41239;
assign n_41241 = ~x_3806 & ~n_41239;
assign n_41242 = ~n_41240 & ~n_41241;
assign n_41243 =  x_3805 & ~n_26992;
assign n_41244 =  x_3805 &  n_41243;
assign n_41245 = ~x_3805 & ~n_41243;
assign n_41246 = ~n_41244 & ~n_41245;
assign n_41247 =  x_3804 & ~n_26992;
assign n_41248 =  x_3804 &  n_41247;
assign n_41249 = ~x_3804 & ~n_41247;
assign n_41250 = ~n_41248 & ~n_41249;
assign n_41251 =  x_3803 & ~n_26992;
assign n_41252 =  x_3803 &  n_41251;
assign n_41253 = ~x_3803 & ~n_41251;
assign n_41254 = ~n_41252 & ~n_41253;
assign n_41255 =  x_3802 & ~n_26992;
assign n_41256 =  x_3802 &  n_41255;
assign n_41257 = ~x_3802 & ~n_41255;
assign n_41258 = ~n_41256 & ~n_41257;
assign n_41259 =  x_3801 & ~n_26992;
assign n_41260 =  x_3801 &  n_41259;
assign n_41261 = ~x_3801 & ~n_41259;
assign n_41262 = ~n_41260 & ~n_41261;
assign n_41263 =  x_3800 & ~n_26992;
assign n_41264 =  x_3800 &  n_41263;
assign n_41265 = ~x_3800 & ~n_41263;
assign n_41266 = ~n_41264 & ~n_41265;
assign n_41267 = ~n_26709 & ~n_26174;
assign n_41268 = ~n_25878 &  n_41267;
assign n_41269 = ~n_28543 &  n_41268;
assign n_41270 =  x_3799 &  n_41269;
assign n_41271 =  x_1130 &  n_28543;
assign n_41272 =  x_2650 &  n_26174;
assign n_41273 =  x_1642 &  n_25878;
assign n_41274 =  x_4999 &  n_26709;
assign n_41275 = ~n_41273 & ~n_41274;
assign n_41276 = ~n_41272 &  n_41275;
assign n_41277 = ~n_41271 &  n_41276;
assign n_41278 = ~n_41270 &  n_41277;
assign n_41279 =  x_3799 & ~n_41278;
assign n_41280 = ~x_3799 &  n_41278;
assign n_41281 = ~n_41279 & ~n_41280;
assign n_41282 =  x_3798 &  n_41269;
assign n_41283 =  x_1129 &  n_28543;
assign n_41284 =  x_2649 &  n_26174;
assign n_41285 =  x_1641 &  n_25878;
assign n_41286 =  x_4998 &  n_26709;
assign n_41287 = ~n_41285 & ~n_41286;
assign n_41288 = ~n_41284 &  n_41287;
assign n_41289 = ~n_41283 &  n_41288;
assign n_41290 = ~n_41282 &  n_41289;
assign n_41291 =  x_3798 & ~n_41290;
assign n_41292 = ~x_3798 &  n_41290;
assign n_41293 = ~n_41291 & ~n_41292;
assign n_41294 =  x_3797 &  n_41269;
assign n_41295 =  x_1128 &  n_28543;
assign n_41296 =  x_2648 &  n_26174;
assign n_41297 =  x_1640 &  n_25878;
assign n_41298 =  x_4997 &  n_26709;
assign n_41299 = ~n_41297 & ~n_41298;
assign n_41300 = ~n_41296 &  n_41299;
assign n_41301 = ~n_41295 &  n_41300;
assign n_41302 = ~n_41294 &  n_41301;
assign n_41303 =  x_3797 & ~n_41302;
assign n_41304 = ~x_3797 &  n_41302;
assign n_41305 = ~n_41303 & ~n_41304;
assign n_41306 =  x_3796 &  n_41269;
assign n_41307 =  x_1127 &  n_28543;
assign n_41308 =  x_2647 &  n_26174;
assign n_41309 =  x_1639 &  n_25878;
assign n_41310 =  x_4996 &  n_26709;
assign n_41311 = ~n_41309 & ~n_41310;
assign n_41312 = ~n_41308 &  n_41311;
assign n_41313 = ~n_41307 &  n_41312;
assign n_41314 = ~n_41306 &  n_41313;
assign n_41315 =  x_3796 & ~n_41314;
assign n_41316 = ~x_3796 &  n_41314;
assign n_41317 = ~n_41315 & ~n_41316;
assign n_41318 =  x_3795 &  n_41269;
assign n_41319 =  x_1126 &  n_28543;
assign n_41320 =  x_2646 &  n_26174;
assign n_41321 =  x_1638 &  n_25878;
assign n_41322 =  x_4995 &  n_26709;
assign n_41323 = ~n_41321 & ~n_41322;
assign n_41324 = ~n_41320 &  n_41323;
assign n_41325 = ~n_41319 &  n_41324;
assign n_41326 = ~n_41318 &  n_41325;
assign n_41327 =  x_3795 & ~n_41326;
assign n_41328 = ~x_3795 &  n_41326;
assign n_41329 = ~n_41327 & ~n_41328;
assign n_41330 =  x_3794 &  n_41269;
assign n_41331 =  x_1125 &  n_28543;
assign n_41332 =  x_2645 &  n_26174;
assign n_41333 =  x_1637 &  n_25878;
assign n_41334 =  x_4994 &  n_26709;
assign n_41335 = ~n_41333 & ~n_41334;
assign n_41336 = ~n_41332 &  n_41335;
assign n_41337 = ~n_41331 &  n_41336;
assign n_41338 = ~n_41330 &  n_41337;
assign n_41339 =  x_3794 & ~n_41338;
assign n_41340 = ~x_3794 &  n_41338;
assign n_41341 = ~n_41339 & ~n_41340;
assign n_41342 =  x_3793 &  n_41269;
assign n_41343 =  x_1124 &  n_28543;
assign n_41344 =  x_2644 &  n_26174;
assign n_41345 =  x_1636 &  n_25878;
assign n_41346 =  x_4993 &  n_26709;
assign n_41347 = ~n_41345 & ~n_41346;
assign n_41348 = ~n_41344 &  n_41347;
assign n_41349 = ~n_41343 &  n_41348;
assign n_41350 = ~n_41342 &  n_41349;
assign n_41351 =  x_3793 & ~n_41350;
assign n_41352 = ~x_3793 &  n_41350;
assign n_41353 = ~n_41351 & ~n_41352;
assign n_41354 =  x_3792 &  n_41269;
assign n_41355 =  x_1123 &  n_28543;
assign n_41356 =  x_2643 &  n_26174;
assign n_41357 =  x_1635 &  n_25878;
assign n_41358 =  x_4992 &  n_26709;
assign n_41359 = ~n_41357 & ~n_41358;
assign n_41360 = ~n_41356 &  n_41359;
assign n_41361 = ~n_41355 &  n_41360;
assign n_41362 = ~n_41354 &  n_41361;
assign n_41363 =  x_3792 & ~n_41362;
assign n_41364 = ~x_3792 &  n_41362;
assign n_41365 = ~n_41363 & ~n_41364;
assign n_41366 =  x_3791 &  n_41269;
assign n_41367 =  x_1122 &  n_28543;
assign n_41368 =  x_2642 &  n_26174;
assign n_41369 =  x_1634 &  n_25878;
assign n_41370 =  x_4991 &  n_26709;
assign n_41371 = ~n_41369 & ~n_41370;
assign n_41372 = ~n_41368 &  n_41371;
assign n_41373 = ~n_41367 &  n_41372;
assign n_41374 = ~n_41366 &  n_41373;
assign n_41375 =  x_3791 & ~n_41374;
assign n_41376 = ~x_3791 &  n_41374;
assign n_41377 = ~n_41375 & ~n_41376;
assign n_41378 =  x_3790 &  n_41269;
assign n_41379 =  x_1121 &  n_28543;
assign n_41380 =  x_2641 &  n_26174;
assign n_41381 =  x_1633 &  n_25878;
assign n_41382 =  x_4990 &  n_26709;
assign n_41383 = ~n_41381 & ~n_41382;
assign n_41384 = ~n_41380 &  n_41383;
assign n_41385 = ~n_41379 &  n_41384;
assign n_41386 = ~n_41378 &  n_41385;
assign n_41387 =  x_3790 & ~n_41386;
assign n_41388 = ~x_3790 &  n_41386;
assign n_41389 = ~n_41387 & ~n_41388;
assign n_41390 =  x_3789 &  n_41269;
assign n_41391 =  x_1120 &  n_28543;
assign n_41392 =  x_2640 &  n_26174;
assign n_41393 =  x_1632 &  n_25878;
assign n_41394 =  x_4989 &  n_26709;
assign n_41395 = ~n_41393 & ~n_41394;
assign n_41396 = ~n_41392 &  n_41395;
assign n_41397 = ~n_41391 &  n_41396;
assign n_41398 = ~n_41390 &  n_41397;
assign n_41399 =  x_3789 & ~n_41398;
assign n_41400 = ~x_3789 &  n_41398;
assign n_41401 = ~n_41399 & ~n_41400;
assign n_41402 =  x_3788 &  n_41269;
assign n_41403 =  x_1119 &  n_28543;
assign n_41404 =  x_2639 &  n_26174;
assign n_41405 =  x_1631 &  n_25878;
assign n_41406 =  x_4988 &  n_26709;
assign n_41407 = ~n_41405 & ~n_41406;
assign n_41408 = ~n_41404 &  n_41407;
assign n_41409 = ~n_41403 &  n_41408;
assign n_41410 = ~n_41402 &  n_41409;
assign n_41411 =  x_3788 & ~n_41410;
assign n_41412 = ~x_3788 &  n_41410;
assign n_41413 = ~n_41411 & ~n_41412;
assign n_41414 =  x_3787 &  n_41269;
assign n_41415 =  x_1118 &  n_28543;
assign n_41416 =  x_2638 &  n_26174;
assign n_41417 =  x_1630 &  n_25878;
assign n_41418 =  x_4987 &  n_26709;
assign n_41419 = ~n_41417 & ~n_41418;
assign n_41420 = ~n_41416 &  n_41419;
assign n_41421 = ~n_41415 &  n_41420;
assign n_41422 = ~n_41414 &  n_41421;
assign n_41423 =  x_3787 & ~n_41422;
assign n_41424 = ~x_3787 &  n_41422;
assign n_41425 = ~n_41423 & ~n_41424;
assign n_41426 =  x_3786 &  n_41269;
assign n_41427 =  x_1117 &  n_28543;
assign n_41428 =  x_2637 &  n_26174;
assign n_41429 =  x_1629 &  n_25878;
assign n_41430 =  x_4986 &  n_26709;
assign n_41431 = ~n_41429 & ~n_41430;
assign n_41432 = ~n_41428 &  n_41431;
assign n_41433 = ~n_41427 &  n_41432;
assign n_41434 = ~n_41426 &  n_41433;
assign n_41435 =  x_3786 & ~n_41434;
assign n_41436 = ~x_3786 &  n_41434;
assign n_41437 = ~n_41435 & ~n_41436;
assign n_41438 =  x_3785 &  n_41269;
assign n_41439 =  x_1116 &  n_28543;
assign n_41440 =  x_2636 &  n_26174;
assign n_41441 =  x_1628 &  n_25878;
assign n_41442 =  x_4985 &  n_26709;
assign n_41443 = ~n_41441 & ~n_41442;
assign n_41444 = ~n_41440 &  n_41443;
assign n_41445 = ~n_41439 &  n_41444;
assign n_41446 = ~n_41438 &  n_41445;
assign n_41447 =  x_3785 & ~n_41446;
assign n_41448 = ~x_3785 &  n_41446;
assign n_41449 = ~n_41447 & ~n_41448;
assign n_41450 =  x_3784 &  n_41269;
assign n_41451 =  x_1115 &  n_28543;
assign n_41452 =  x_2635 &  n_26174;
assign n_41453 =  x_1627 &  n_25878;
assign n_41454 =  x_4984 &  n_26709;
assign n_41455 = ~n_41453 & ~n_41454;
assign n_41456 = ~n_41452 &  n_41455;
assign n_41457 = ~n_41451 &  n_41456;
assign n_41458 = ~n_41450 &  n_41457;
assign n_41459 =  x_3784 & ~n_41458;
assign n_41460 = ~x_3784 &  n_41458;
assign n_41461 = ~n_41459 & ~n_41460;
assign n_41462 =  x_3783 &  n_41269;
assign n_41463 =  x_1114 &  n_28543;
assign n_41464 =  x_2634 &  n_26174;
assign n_41465 =  x_1626 &  n_25878;
assign n_41466 =  x_4983 &  n_26709;
assign n_41467 = ~n_41465 & ~n_41466;
assign n_41468 = ~n_41464 &  n_41467;
assign n_41469 = ~n_41463 &  n_41468;
assign n_41470 = ~n_41462 &  n_41469;
assign n_41471 =  x_3783 & ~n_41470;
assign n_41472 = ~x_3783 &  n_41470;
assign n_41473 = ~n_41471 & ~n_41472;
assign n_41474 =  x_3782 &  n_41269;
assign n_41475 =  x_1113 &  n_28543;
assign n_41476 =  x_2633 &  n_26174;
assign n_41477 =  x_1625 &  n_25878;
assign n_41478 =  x_4982 &  n_26709;
assign n_41479 = ~n_41477 & ~n_41478;
assign n_41480 = ~n_41476 &  n_41479;
assign n_41481 = ~n_41475 &  n_41480;
assign n_41482 = ~n_41474 &  n_41481;
assign n_41483 =  x_3782 & ~n_41482;
assign n_41484 = ~x_3782 &  n_41482;
assign n_41485 = ~n_41483 & ~n_41484;
assign n_41486 =  x_3781 &  n_41269;
assign n_41487 =  x_1112 &  n_28543;
assign n_41488 =  x_2632 &  n_26174;
assign n_41489 =  x_1624 &  n_25878;
assign n_41490 =  x_4981 &  n_26709;
assign n_41491 = ~n_41489 & ~n_41490;
assign n_41492 = ~n_41488 &  n_41491;
assign n_41493 = ~n_41487 &  n_41492;
assign n_41494 = ~n_41486 &  n_41493;
assign n_41495 =  x_3781 & ~n_41494;
assign n_41496 = ~x_3781 &  n_41494;
assign n_41497 = ~n_41495 & ~n_41496;
assign n_41498 =  x_3780 &  n_41269;
assign n_41499 =  x_1111 &  n_28543;
assign n_41500 =  x_2631 &  n_26174;
assign n_41501 =  x_1623 &  n_25878;
assign n_41502 =  x_4980 &  n_26709;
assign n_41503 = ~n_41501 & ~n_41502;
assign n_41504 = ~n_41500 &  n_41503;
assign n_41505 = ~n_41499 &  n_41504;
assign n_41506 = ~n_41498 &  n_41505;
assign n_41507 =  x_3780 & ~n_41506;
assign n_41508 = ~x_3780 &  n_41506;
assign n_41509 = ~n_41507 & ~n_41508;
assign n_41510 =  x_3779 &  n_41269;
assign n_41511 =  x_1110 &  n_28543;
assign n_41512 =  x_2630 &  n_26174;
assign n_41513 =  x_1622 &  n_25878;
assign n_41514 =  x_4979 &  n_26709;
assign n_41515 = ~n_41513 & ~n_41514;
assign n_41516 = ~n_41512 &  n_41515;
assign n_41517 = ~n_41511 &  n_41516;
assign n_41518 = ~n_41510 &  n_41517;
assign n_41519 =  x_3779 & ~n_41518;
assign n_41520 = ~x_3779 &  n_41518;
assign n_41521 = ~n_41519 & ~n_41520;
assign n_41522 =  x_3778 &  n_41269;
assign n_41523 =  x_1109 &  n_28543;
assign n_41524 =  x_2629 &  n_26174;
assign n_41525 =  x_1621 &  n_25878;
assign n_41526 =  x_4978 &  n_26709;
assign n_41527 = ~n_41525 & ~n_41526;
assign n_41528 = ~n_41524 &  n_41527;
assign n_41529 = ~n_41523 &  n_41528;
assign n_41530 = ~n_41522 &  n_41529;
assign n_41531 =  x_3778 & ~n_41530;
assign n_41532 = ~x_3778 &  n_41530;
assign n_41533 = ~n_41531 & ~n_41532;
assign n_41534 =  x_3777 &  n_41269;
assign n_41535 =  x_1108 &  n_28543;
assign n_41536 =  x_2628 &  n_26174;
assign n_41537 =  x_1620 &  n_25878;
assign n_41538 =  x_4977 &  n_26709;
assign n_41539 = ~n_41537 & ~n_41538;
assign n_41540 = ~n_41536 &  n_41539;
assign n_41541 = ~n_41535 &  n_41540;
assign n_41542 = ~n_41534 &  n_41541;
assign n_41543 =  x_3777 & ~n_41542;
assign n_41544 = ~x_3777 &  n_41542;
assign n_41545 = ~n_41543 & ~n_41544;
assign n_41546 =  x_3776 &  n_41269;
assign n_41547 =  x_1107 &  n_28543;
assign n_41548 =  x_2627 &  n_26174;
assign n_41549 =  x_1619 &  n_25878;
assign n_41550 =  x_4976 &  n_26709;
assign n_41551 = ~n_41549 & ~n_41550;
assign n_41552 = ~n_41548 &  n_41551;
assign n_41553 = ~n_41547 &  n_41552;
assign n_41554 = ~n_41546 &  n_41553;
assign n_41555 =  x_3776 & ~n_41554;
assign n_41556 = ~x_3776 &  n_41554;
assign n_41557 = ~n_41555 & ~n_41556;
assign n_41558 =  x_3775 &  n_41269;
assign n_41559 =  x_1106 &  n_28543;
assign n_41560 =  x_2626 &  n_26174;
assign n_41561 =  x_1618 &  n_25878;
assign n_41562 =  x_4975 &  n_26709;
assign n_41563 = ~n_41561 & ~n_41562;
assign n_41564 = ~n_41560 &  n_41563;
assign n_41565 = ~n_41559 &  n_41564;
assign n_41566 = ~n_41558 &  n_41565;
assign n_41567 =  x_3775 & ~n_41566;
assign n_41568 = ~x_3775 &  n_41566;
assign n_41569 = ~n_41567 & ~n_41568;
assign n_41570 =  x_3774 &  n_41269;
assign n_41571 =  x_1105 &  n_28543;
assign n_41572 =  x_2625 &  n_26174;
assign n_41573 =  x_1617 &  n_25878;
assign n_41574 =  x_4974 &  n_26709;
assign n_41575 = ~n_41573 & ~n_41574;
assign n_41576 = ~n_41572 &  n_41575;
assign n_41577 = ~n_41571 &  n_41576;
assign n_41578 = ~n_41570 &  n_41577;
assign n_41579 =  x_3774 & ~n_41578;
assign n_41580 = ~x_3774 &  n_41578;
assign n_41581 = ~n_41579 & ~n_41580;
assign n_41582 =  x_3773 &  n_41269;
assign n_41583 =  x_1104 &  n_28543;
assign n_41584 =  x_2624 &  n_26174;
assign n_41585 =  x_1616 &  n_25878;
assign n_41586 =  x_4973 &  n_26709;
assign n_41587 = ~n_41585 & ~n_41586;
assign n_41588 = ~n_41584 &  n_41587;
assign n_41589 = ~n_41583 &  n_41588;
assign n_41590 = ~n_41582 &  n_41589;
assign n_41591 =  x_3773 & ~n_41590;
assign n_41592 = ~x_3773 &  n_41590;
assign n_41593 = ~n_41591 & ~n_41592;
assign n_41594 =  x_3772 &  n_41269;
assign n_41595 =  x_1103 &  n_28543;
assign n_41596 =  x_2623 &  n_26174;
assign n_41597 =  x_1615 &  n_25878;
assign n_41598 =  x_4972 &  n_26709;
assign n_41599 = ~n_41597 & ~n_41598;
assign n_41600 = ~n_41596 &  n_41599;
assign n_41601 = ~n_41595 &  n_41600;
assign n_41602 = ~n_41594 &  n_41601;
assign n_41603 =  x_3772 & ~n_41602;
assign n_41604 = ~x_3772 &  n_41602;
assign n_41605 = ~n_41603 & ~n_41604;
assign n_41606 =  x_3771 &  n_41269;
assign n_41607 =  x_1102 &  n_28543;
assign n_41608 =  x_2622 &  n_26174;
assign n_41609 =  x_1614 &  n_25878;
assign n_41610 =  x_4971 &  n_26709;
assign n_41611 = ~n_41609 & ~n_41610;
assign n_41612 = ~n_41608 &  n_41611;
assign n_41613 = ~n_41607 &  n_41612;
assign n_41614 = ~n_41606 &  n_41613;
assign n_41615 =  x_3771 & ~n_41614;
assign n_41616 = ~x_3771 &  n_41614;
assign n_41617 = ~n_41615 & ~n_41616;
assign n_41618 =  x_3770 &  n_41269;
assign n_41619 =  x_1101 &  n_28543;
assign n_41620 =  x_2621 &  n_26174;
assign n_41621 =  x_1613 &  n_25878;
assign n_41622 =  x_4970 &  n_26709;
assign n_41623 = ~n_41621 & ~n_41622;
assign n_41624 = ~n_41620 &  n_41623;
assign n_41625 = ~n_41619 &  n_41624;
assign n_41626 = ~n_41618 &  n_41625;
assign n_41627 =  x_3770 & ~n_41626;
assign n_41628 = ~x_3770 &  n_41626;
assign n_41629 = ~n_41627 & ~n_41628;
assign n_41630 =  x_3769 &  n_41269;
assign n_41631 =  x_1100 &  n_28543;
assign n_41632 =  x_2620 &  n_26174;
assign n_41633 =  x_1612 &  n_25878;
assign n_41634 =  x_4969 &  n_26709;
assign n_41635 = ~n_41633 & ~n_41634;
assign n_41636 = ~n_41632 &  n_41635;
assign n_41637 = ~n_41631 &  n_41636;
assign n_41638 = ~n_41630 &  n_41637;
assign n_41639 =  x_3769 & ~n_41638;
assign n_41640 = ~x_3769 &  n_41638;
assign n_41641 = ~n_41639 & ~n_41640;
assign n_41642 =  x_3768 &  n_41269;
assign n_41643 =  x_1099 &  n_28543;
assign n_41644 =  x_2619 &  n_26174;
assign n_41645 =  x_1611 &  n_25878;
assign n_41646 =  x_4968 &  n_26709;
assign n_41647 = ~n_41645 & ~n_41646;
assign n_41648 = ~n_41644 &  n_41647;
assign n_41649 = ~n_41643 &  n_41648;
assign n_41650 = ~n_41642 &  n_41649;
assign n_41651 =  x_3768 & ~n_41650;
assign n_41652 = ~x_3768 &  n_41650;
assign n_41653 = ~n_41651 & ~n_41652;
assign n_41654 =  n_26824 & ~n_14801;
assign n_41655 =  x_3767 & ~n_26824;
assign n_41656 = ~n_41654 & ~n_41655;
assign n_41657 =  x_3767 & ~n_41656;
assign n_41658 = ~x_3767 &  n_41656;
assign n_41659 = ~n_41657 & ~n_41658;
assign n_41660 =  n_26824 & ~n_14819;
assign n_41661 =  x_3766 & ~n_26824;
assign n_41662 = ~n_41660 & ~n_41661;
assign n_41663 =  x_3766 & ~n_41662;
assign n_41664 = ~x_3766 &  n_41662;
assign n_41665 = ~n_41663 & ~n_41664;
assign n_41666 =  n_26824 & ~n_14837;
assign n_41667 =  x_3765 & ~n_26824;
assign n_41668 = ~n_41666 & ~n_41667;
assign n_41669 =  x_3765 & ~n_41668;
assign n_41670 = ~x_3765 &  n_41668;
assign n_41671 = ~n_41669 & ~n_41670;
assign n_41672 =  n_26824 & ~n_14855;
assign n_41673 =  x_3764 & ~n_26824;
assign n_41674 = ~n_41672 & ~n_41673;
assign n_41675 =  x_3764 & ~n_41674;
assign n_41676 = ~x_3764 &  n_41674;
assign n_41677 = ~n_41675 & ~n_41676;
assign n_41678 =  n_26824 & ~n_14873;
assign n_41679 =  x_3763 & ~n_26824;
assign n_41680 = ~n_41678 & ~n_41679;
assign n_41681 =  x_3763 & ~n_41680;
assign n_41682 = ~x_3763 &  n_41680;
assign n_41683 = ~n_41681 & ~n_41682;
assign n_41684 =  n_26824 & ~n_14891;
assign n_41685 =  x_3762 & ~n_26824;
assign n_41686 = ~n_41684 & ~n_41685;
assign n_41687 =  x_3762 & ~n_41686;
assign n_41688 = ~x_3762 &  n_41686;
assign n_41689 = ~n_41687 & ~n_41688;
assign n_41690 =  n_26824 & ~n_14909;
assign n_41691 =  x_3761 & ~n_26824;
assign n_41692 = ~n_41690 & ~n_41691;
assign n_41693 =  x_3761 & ~n_41692;
assign n_41694 = ~x_3761 &  n_41692;
assign n_41695 = ~n_41693 & ~n_41694;
assign n_41696 =  n_26824 & ~n_14927;
assign n_41697 =  x_3760 & ~n_26824;
assign n_41698 = ~n_41696 & ~n_41697;
assign n_41699 =  x_3760 & ~n_41698;
assign n_41700 = ~x_3760 &  n_41698;
assign n_41701 = ~n_41699 & ~n_41700;
assign n_41702 =  n_26824 & ~n_14945;
assign n_41703 =  x_3759 & ~n_26824;
assign n_41704 = ~n_41702 & ~n_41703;
assign n_41705 =  x_3759 & ~n_41704;
assign n_41706 = ~x_3759 &  n_41704;
assign n_41707 = ~n_41705 & ~n_41706;
assign n_41708 =  n_26824 & ~n_14963;
assign n_41709 =  x_3758 & ~n_26824;
assign n_41710 = ~n_41708 & ~n_41709;
assign n_41711 =  x_3758 & ~n_41710;
assign n_41712 = ~x_3758 &  n_41710;
assign n_41713 = ~n_41711 & ~n_41712;
assign n_41714 =  n_26824 & ~n_14981;
assign n_41715 =  x_3757 & ~n_26824;
assign n_41716 = ~n_41714 & ~n_41715;
assign n_41717 =  x_3757 & ~n_41716;
assign n_41718 = ~x_3757 &  n_41716;
assign n_41719 = ~n_41717 & ~n_41718;
assign n_41720 =  n_26824 & ~n_14999;
assign n_41721 =  x_3756 & ~n_26824;
assign n_41722 = ~n_41720 & ~n_41721;
assign n_41723 =  x_3756 & ~n_41722;
assign n_41724 = ~x_3756 &  n_41722;
assign n_41725 = ~n_41723 & ~n_41724;
assign n_41726 =  n_26824 & ~n_15017;
assign n_41727 =  x_3755 & ~n_26824;
assign n_41728 = ~n_41726 & ~n_41727;
assign n_41729 =  x_3755 & ~n_41728;
assign n_41730 = ~x_3755 &  n_41728;
assign n_41731 = ~n_41729 & ~n_41730;
assign n_41732 =  n_26824 & ~n_15035;
assign n_41733 =  x_3754 & ~n_26824;
assign n_41734 = ~n_41732 & ~n_41733;
assign n_41735 =  x_3754 & ~n_41734;
assign n_41736 = ~x_3754 &  n_41734;
assign n_41737 = ~n_41735 & ~n_41736;
assign n_41738 =  n_26824 & ~n_15053;
assign n_41739 =  x_3753 & ~n_26824;
assign n_41740 = ~n_41738 & ~n_41739;
assign n_41741 =  x_3753 & ~n_41740;
assign n_41742 = ~x_3753 &  n_41740;
assign n_41743 = ~n_41741 & ~n_41742;
assign n_41744 =  n_26824 & ~n_15071;
assign n_41745 =  x_3752 & ~n_26824;
assign n_41746 = ~n_41744 & ~n_41745;
assign n_41747 =  x_3752 & ~n_41746;
assign n_41748 = ~x_3752 &  n_41746;
assign n_41749 = ~n_41747 & ~n_41748;
assign n_41750 =  n_26824 & ~n_15089;
assign n_41751 =  x_3751 & ~n_26824;
assign n_41752 = ~n_41750 & ~n_41751;
assign n_41753 =  x_3751 & ~n_41752;
assign n_41754 = ~x_3751 &  n_41752;
assign n_41755 = ~n_41753 & ~n_41754;
assign n_41756 =  n_26824 & ~n_15107;
assign n_41757 =  x_3750 & ~n_26824;
assign n_41758 = ~n_41756 & ~n_41757;
assign n_41759 =  x_3750 & ~n_41758;
assign n_41760 = ~x_3750 &  n_41758;
assign n_41761 = ~n_41759 & ~n_41760;
assign n_41762 =  n_26824 & ~n_15125;
assign n_41763 =  x_3749 & ~n_26824;
assign n_41764 = ~n_41762 & ~n_41763;
assign n_41765 =  x_3749 & ~n_41764;
assign n_41766 = ~x_3749 &  n_41764;
assign n_41767 = ~n_41765 & ~n_41766;
assign n_41768 =  n_26824 & ~n_15143;
assign n_41769 =  x_3748 & ~n_26824;
assign n_41770 = ~n_41768 & ~n_41769;
assign n_41771 =  x_3748 & ~n_41770;
assign n_41772 = ~x_3748 &  n_41770;
assign n_41773 = ~n_41771 & ~n_41772;
assign n_41774 =  n_26824 & ~n_15161;
assign n_41775 =  x_3747 & ~n_26824;
assign n_41776 = ~n_41774 & ~n_41775;
assign n_41777 =  x_3747 & ~n_41776;
assign n_41778 = ~x_3747 &  n_41776;
assign n_41779 = ~n_41777 & ~n_41778;
assign n_41780 =  n_26824 & ~n_15179;
assign n_41781 =  x_3746 & ~n_26824;
assign n_41782 = ~n_41780 & ~n_41781;
assign n_41783 =  x_3746 & ~n_41782;
assign n_41784 = ~x_3746 &  n_41782;
assign n_41785 = ~n_41783 & ~n_41784;
assign n_41786 =  n_26824 & ~n_15197;
assign n_41787 =  x_3745 & ~n_26824;
assign n_41788 = ~n_41786 & ~n_41787;
assign n_41789 =  x_3745 & ~n_41788;
assign n_41790 = ~x_3745 &  n_41788;
assign n_41791 = ~n_41789 & ~n_41790;
assign n_41792 =  n_26824 & ~n_15215;
assign n_41793 =  x_3744 & ~n_26824;
assign n_41794 = ~n_41792 & ~n_41793;
assign n_41795 =  x_3744 & ~n_41794;
assign n_41796 = ~x_3744 &  n_41794;
assign n_41797 = ~n_41795 & ~n_41796;
assign n_41798 =  n_26824 & ~n_15233;
assign n_41799 =  x_3743 & ~n_26824;
assign n_41800 = ~n_41798 & ~n_41799;
assign n_41801 =  x_3743 & ~n_41800;
assign n_41802 = ~x_3743 &  n_41800;
assign n_41803 = ~n_41801 & ~n_41802;
assign n_41804 =  n_26824 & ~n_15251;
assign n_41805 =  x_3742 & ~n_26824;
assign n_41806 = ~n_41804 & ~n_41805;
assign n_41807 =  x_3742 & ~n_41806;
assign n_41808 = ~x_3742 &  n_41806;
assign n_41809 = ~n_41807 & ~n_41808;
assign n_41810 =  n_26824 & ~n_15269;
assign n_41811 =  x_3741 & ~n_26824;
assign n_41812 = ~n_41810 & ~n_41811;
assign n_41813 =  x_3741 & ~n_41812;
assign n_41814 = ~x_3741 &  n_41812;
assign n_41815 = ~n_41813 & ~n_41814;
assign n_41816 =  n_26824 & ~n_15287;
assign n_41817 =  x_3740 & ~n_26824;
assign n_41818 = ~n_41816 & ~n_41817;
assign n_41819 =  x_3740 & ~n_41818;
assign n_41820 = ~x_3740 &  n_41818;
assign n_41821 = ~n_41819 & ~n_41820;
assign n_41822 =  n_26824 & ~n_15305;
assign n_41823 =  x_3739 & ~n_26824;
assign n_41824 = ~n_41822 & ~n_41823;
assign n_41825 =  x_3739 & ~n_41824;
assign n_41826 = ~x_3739 &  n_41824;
assign n_41827 = ~n_41825 & ~n_41826;
assign n_41828 =  n_26824 & ~n_15323;
assign n_41829 =  x_3738 & ~n_26824;
assign n_41830 = ~n_41828 & ~n_41829;
assign n_41831 =  x_3738 & ~n_41830;
assign n_41832 = ~x_3738 &  n_41830;
assign n_41833 = ~n_41831 & ~n_41832;
assign n_41834 =  n_26824 & ~n_15341;
assign n_41835 =  x_3737 & ~n_26824;
assign n_41836 = ~n_41834 & ~n_41835;
assign n_41837 =  x_3737 & ~n_41836;
assign n_41838 = ~x_3737 &  n_41836;
assign n_41839 = ~n_41837 & ~n_41838;
assign n_41840 =  n_26824 & ~n_15359;
assign n_41841 =  x_3736 & ~n_26824;
assign n_41842 = ~n_41840 & ~n_41841;
assign n_41843 =  x_3736 & ~n_41842;
assign n_41844 = ~x_3736 &  n_41842;
assign n_41845 = ~n_41843 & ~n_41844;
assign n_41846 =  x_3735 & ~n_25969;
assign n_41847 =  i_32 &  n_25969;
assign n_41848 = ~n_41846 & ~n_41847;
assign n_41849 =  x_3735 & ~n_41848;
assign n_41850 = ~x_3735 &  n_41848;
assign n_41851 = ~n_41849 & ~n_41850;
assign n_41852 =  x_3734 & ~n_25969;
assign n_41853 =  i_31 &  n_25969;
assign n_41854 = ~n_41852 & ~n_41853;
assign n_41855 =  x_3734 & ~n_41854;
assign n_41856 = ~x_3734 &  n_41854;
assign n_41857 = ~n_41855 & ~n_41856;
assign n_41858 =  x_3733 & ~n_25969;
assign n_41859 =  i_30 &  n_25969;
assign n_41860 = ~n_41858 & ~n_41859;
assign n_41861 =  x_3733 & ~n_41860;
assign n_41862 = ~x_3733 &  n_41860;
assign n_41863 = ~n_41861 & ~n_41862;
assign n_41864 =  x_3732 & ~n_25969;
assign n_41865 =  i_29 &  n_25969;
assign n_41866 = ~n_41864 & ~n_41865;
assign n_41867 =  x_3732 & ~n_41866;
assign n_41868 = ~x_3732 &  n_41866;
assign n_41869 = ~n_41867 & ~n_41868;
assign n_41870 =  x_3731 & ~n_25969;
assign n_41871 =  i_28 &  n_25969;
assign n_41872 = ~n_41870 & ~n_41871;
assign n_41873 =  x_3731 & ~n_41872;
assign n_41874 = ~x_3731 &  n_41872;
assign n_41875 = ~n_41873 & ~n_41874;
assign n_41876 =  x_3730 & ~n_25969;
assign n_41877 =  i_27 &  n_25969;
assign n_41878 = ~n_41876 & ~n_41877;
assign n_41879 =  x_3730 & ~n_41878;
assign n_41880 = ~x_3730 &  n_41878;
assign n_41881 = ~n_41879 & ~n_41880;
assign n_41882 =  x_3729 & ~n_25969;
assign n_41883 =  i_26 &  n_25969;
assign n_41884 = ~n_41882 & ~n_41883;
assign n_41885 =  x_3729 & ~n_41884;
assign n_41886 = ~x_3729 &  n_41884;
assign n_41887 = ~n_41885 & ~n_41886;
assign n_41888 =  x_3728 & ~n_25969;
assign n_41889 =  i_25 &  n_25969;
assign n_41890 = ~n_41888 & ~n_41889;
assign n_41891 =  x_3728 & ~n_41890;
assign n_41892 = ~x_3728 &  n_41890;
assign n_41893 = ~n_41891 & ~n_41892;
assign n_41894 =  x_3727 & ~n_25969;
assign n_41895 =  i_24 &  n_25969;
assign n_41896 = ~n_41894 & ~n_41895;
assign n_41897 =  x_3727 & ~n_41896;
assign n_41898 = ~x_3727 &  n_41896;
assign n_41899 = ~n_41897 & ~n_41898;
assign n_41900 =  x_3726 & ~n_25969;
assign n_41901 =  i_23 &  n_25969;
assign n_41902 = ~n_41900 & ~n_41901;
assign n_41903 =  x_3726 & ~n_41902;
assign n_41904 = ~x_3726 &  n_41902;
assign n_41905 = ~n_41903 & ~n_41904;
assign n_41906 =  x_3725 & ~n_25969;
assign n_41907 =  i_22 &  n_25969;
assign n_41908 = ~n_41906 & ~n_41907;
assign n_41909 =  x_3725 & ~n_41908;
assign n_41910 = ~x_3725 &  n_41908;
assign n_41911 = ~n_41909 & ~n_41910;
assign n_41912 =  x_3724 & ~n_25969;
assign n_41913 =  i_21 &  n_25969;
assign n_41914 = ~n_41912 & ~n_41913;
assign n_41915 =  x_3724 & ~n_41914;
assign n_41916 = ~x_3724 &  n_41914;
assign n_41917 = ~n_41915 & ~n_41916;
assign n_41918 =  x_3723 & ~n_25969;
assign n_41919 =  i_20 &  n_25969;
assign n_41920 = ~n_41918 & ~n_41919;
assign n_41921 =  x_3723 & ~n_41920;
assign n_41922 = ~x_3723 &  n_41920;
assign n_41923 = ~n_41921 & ~n_41922;
assign n_41924 =  x_3722 & ~n_25969;
assign n_41925 =  i_19 &  n_25969;
assign n_41926 = ~n_41924 & ~n_41925;
assign n_41927 =  x_3722 & ~n_41926;
assign n_41928 = ~x_3722 &  n_41926;
assign n_41929 = ~n_41927 & ~n_41928;
assign n_41930 =  x_3721 & ~n_25969;
assign n_41931 =  i_18 &  n_25969;
assign n_41932 = ~n_41930 & ~n_41931;
assign n_41933 =  x_3721 & ~n_41932;
assign n_41934 = ~x_3721 &  n_41932;
assign n_41935 = ~n_41933 & ~n_41934;
assign n_41936 =  x_3720 & ~n_25969;
assign n_41937 =  i_17 &  n_25969;
assign n_41938 = ~n_41936 & ~n_41937;
assign n_41939 =  x_3720 & ~n_41938;
assign n_41940 = ~x_3720 &  n_41938;
assign n_41941 = ~n_41939 & ~n_41940;
assign n_41942 =  x_3719 & ~n_25969;
assign n_41943 =  i_16 &  n_25969;
assign n_41944 = ~n_41942 & ~n_41943;
assign n_41945 =  x_3719 & ~n_41944;
assign n_41946 = ~x_3719 &  n_41944;
assign n_41947 = ~n_41945 & ~n_41946;
assign n_41948 =  x_3718 & ~n_25969;
assign n_41949 =  i_15 &  n_25969;
assign n_41950 = ~n_41948 & ~n_41949;
assign n_41951 =  x_3718 & ~n_41950;
assign n_41952 = ~x_3718 &  n_41950;
assign n_41953 = ~n_41951 & ~n_41952;
assign n_41954 =  x_3717 & ~n_25969;
assign n_41955 =  i_14 &  n_25969;
assign n_41956 = ~n_41954 & ~n_41955;
assign n_41957 =  x_3717 & ~n_41956;
assign n_41958 = ~x_3717 &  n_41956;
assign n_41959 = ~n_41957 & ~n_41958;
assign n_41960 =  x_3716 & ~n_25969;
assign n_41961 =  i_13 &  n_25969;
assign n_41962 = ~n_41960 & ~n_41961;
assign n_41963 =  x_3716 & ~n_41962;
assign n_41964 = ~x_3716 &  n_41962;
assign n_41965 = ~n_41963 & ~n_41964;
assign n_41966 =  x_3715 & ~n_25969;
assign n_41967 =  i_12 &  n_25969;
assign n_41968 = ~n_41966 & ~n_41967;
assign n_41969 =  x_3715 & ~n_41968;
assign n_41970 = ~x_3715 &  n_41968;
assign n_41971 = ~n_41969 & ~n_41970;
assign n_41972 =  x_3714 & ~n_25969;
assign n_41973 =  i_11 &  n_25969;
assign n_41974 = ~n_41972 & ~n_41973;
assign n_41975 =  x_3714 & ~n_41974;
assign n_41976 = ~x_3714 &  n_41974;
assign n_41977 = ~n_41975 & ~n_41976;
assign n_41978 =  x_3713 & ~n_25969;
assign n_41979 =  i_10 &  n_25969;
assign n_41980 = ~n_41978 & ~n_41979;
assign n_41981 =  x_3713 & ~n_41980;
assign n_41982 = ~x_3713 &  n_41980;
assign n_41983 = ~n_41981 & ~n_41982;
assign n_41984 =  x_3712 & ~n_25969;
assign n_41985 =  i_9 &  n_25969;
assign n_41986 = ~n_41984 & ~n_41985;
assign n_41987 =  x_3712 & ~n_41986;
assign n_41988 = ~x_3712 &  n_41986;
assign n_41989 = ~n_41987 & ~n_41988;
assign n_41990 =  x_3711 & ~n_25969;
assign n_41991 =  i_8 &  n_25969;
assign n_41992 = ~n_41990 & ~n_41991;
assign n_41993 =  x_3711 & ~n_41992;
assign n_41994 = ~x_3711 &  n_41992;
assign n_41995 = ~n_41993 & ~n_41994;
assign n_41996 =  x_3710 & ~n_25969;
assign n_41997 =  i_7 &  n_25969;
assign n_41998 = ~n_41996 & ~n_41997;
assign n_41999 =  x_3710 & ~n_41998;
assign n_42000 = ~x_3710 &  n_41998;
assign n_42001 = ~n_41999 & ~n_42000;
assign n_42002 =  x_3709 & ~n_25969;
assign n_42003 =  i_6 &  n_25969;
assign n_42004 = ~n_42002 & ~n_42003;
assign n_42005 =  x_3709 & ~n_42004;
assign n_42006 = ~x_3709 &  n_42004;
assign n_42007 = ~n_42005 & ~n_42006;
assign n_42008 =  x_3708 & ~n_25969;
assign n_42009 =  i_5 &  n_25969;
assign n_42010 = ~n_42008 & ~n_42009;
assign n_42011 =  x_3708 & ~n_42010;
assign n_42012 = ~x_3708 &  n_42010;
assign n_42013 = ~n_42011 & ~n_42012;
assign n_42014 =  x_3707 & ~n_25969;
assign n_42015 =  i_4 &  n_25969;
assign n_42016 = ~n_42014 & ~n_42015;
assign n_42017 =  x_3707 & ~n_42016;
assign n_42018 = ~x_3707 &  n_42016;
assign n_42019 = ~n_42017 & ~n_42018;
assign n_42020 =  x_3706 & ~n_25969;
assign n_42021 =  i_3 &  n_25969;
assign n_42022 = ~n_42020 & ~n_42021;
assign n_42023 =  x_3706 & ~n_42022;
assign n_42024 = ~x_3706 &  n_42022;
assign n_42025 = ~n_42023 & ~n_42024;
assign n_42026 =  x_3705 & ~n_25969;
assign n_42027 =  i_2 &  n_25969;
assign n_42028 = ~n_42026 & ~n_42027;
assign n_42029 =  x_3705 & ~n_42028;
assign n_42030 = ~x_3705 &  n_42028;
assign n_42031 = ~n_42029 & ~n_42030;
assign n_42032 =  x_3704 & ~n_25969;
assign n_42033 =  i_1 &  n_25969;
assign n_42034 = ~n_42032 & ~n_42033;
assign n_42035 =  x_3704 & ~n_42034;
assign n_42036 = ~x_3704 &  n_42034;
assign n_42037 = ~n_42035 & ~n_42036;
assign n_42038 = ~n_24005 & ~n_28297;
assign n_42039 = ~n_24036 &  n_42038;
assign n_42040 = ~n_27857 &  n_42039;
assign n_42041 =  x_3703 &  n_42040;
assign n_42042 =  x_203 &  n_27857;
assign n_42043 =  x_2586 &  n_24036;
assign n_42044 =  x_1098 &  n_24005;
assign n_42045 =  x_3895 &  n_28297;
assign n_42046 = ~n_42044 & ~n_42045;
assign n_42047 = ~n_42043 &  n_42046;
assign n_42048 = ~n_42042 &  n_42047;
assign n_42049 = ~n_42041 &  n_42048;
assign n_42050 =  x_3703 & ~n_42049;
assign n_42051 = ~x_3703 &  n_42049;
assign n_42052 = ~n_42050 & ~n_42051;
assign n_42053 =  x_3702 &  n_42040;
assign n_42054 =  x_202 &  n_27857;
assign n_42055 =  x_2585 &  n_24036;
assign n_42056 =  x_1097 &  n_24005;
assign n_42057 =  x_3894 &  n_28297;
assign n_42058 = ~n_42056 & ~n_42057;
assign n_42059 = ~n_42055 &  n_42058;
assign n_42060 = ~n_42054 &  n_42059;
assign n_42061 = ~n_42053 &  n_42060;
assign n_42062 =  x_3702 & ~n_42061;
assign n_42063 = ~x_3702 &  n_42061;
assign n_42064 = ~n_42062 & ~n_42063;
assign n_42065 =  x_3701 &  n_42040;
assign n_42066 =  x_201 &  n_27857;
assign n_42067 =  x_2584 &  n_24036;
assign n_42068 =  x_1096 &  n_24005;
assign n_42069 =  x_3893 &  n_28297;
assign n_42070 = ~n_42068 & ~n_42069;
assign n_42071 = ~n_42067 &  n_42070;
assign n_42072 = ~n_42066 &  n_42071;
assign n_42073 = ~n_42065 &  n_42072;
assign n_42074 =  x_3701 & ~n_42073;
assign n_42075 = ~x_3701 &  n_42073;
assign n_42076 = ~n_42074 & ~n_42075;
assign n_42077 =  x_3700 &  n_42040;
assign n_42078 =  x_200 &  n_27857;
assign n_42079 =  x_2583 &  n_24036;
assign n_42080 =  x_1095 &  n_24005;
assign n_42081 =  x_3892 &  n_28297;
assign n_42082 = ~n_42080 & ~n_42081;
assign n_42083 = ~n_42079 &  n_42082;
assign n_42084 = ~n_42078 &  n_42083;
assign n_42085 = ~n_42077 &  n_42084;
assign n_42086 =  x_3700 & ~n_42085;
assign n_42087 = ~x_3700 &  n_42085;
assign n_42088 = ~n_42086 & ~n_42087;
assign n_42089 =  x_3699 &  n_42040;
assign n_42090 =  x_199 &  n_27857;
assign n_42091 =  x_2582 &  n_24036;
assign n_42092 =  x_1094 &  n_24005;
assign n_42093 =  x_3891 &  n_28297;
assign n_42094 = ~n_42092 & ~n_42093;
assign n_42095 = ~n_42091 &  n_42094;
assign n_42096 = ~n_42090 &  n_42095;
assign n_42097 = ~n_42089 &  n_42096;
assign n_42098 =  x_3699 & ~n_42097;
assign n_42099 = ~x_3699 &  n_42097;
assign n_42100 = ~n_42098 & ~n_42099;
assign n_42101 =  x_3698 &  n_42040;
assign n_42102 =  x_198 &  n_27857;
assign n_42103 =  x_2581 &  n_24036;
assign n_42104 =  x_1093 &  n_24005;
assign n_42105 =  x_3890 &  n_28297;
assign n_42106 = ~n_42104 & ~n_42105;
assign n_42107 = ~n_42103 &  n_42106;
assign n_42108 = ~n_42102 &  n_42107;
assign n_42109 = ~n_42101 &  n_42108;
assign n_42110 =  x_3698 & ~n_42109;
assign n_42111 = ~x_3698 &  n_42109;
assign n_42112 = ~n_42110 & ~n_42111;
assign n_42113 =  x_3697 &  n_42040;
assign n_42114 =  x_197 &  n_27857;
assign n_42115 =  x_2580 &  n_24036;
assign n_42116 =  x_1092 &  n_24005;
assign n_42117 =  x_3889 &  n_28297;
assign n_42118 = ~n_42116 & ~n_42117;
assign n_42119 = ~n_42115 &  n_42118;
assign n_42120 = ~n_42114 &  n_42119;
assign n_42121 = ~n_42113 &  n_42120;
assign n_42122 =  x_3697 & ~n_42121;
assign n_42123 = ~x_3697 &  n_42121;
assign n_42124 = ~n_42122 & ~n_42123;
assign n_42125 =  x_3696 &  n_42040;
assign n_42126 =  x_196 &  n_27857;
assign n_42127 =  x_2579 &  n_24036;
assign n_42128 =  x_1091 &  n_24005;
assign n_42129 =  x_3888 &  n_28297;
assign n_42130 = ~n_42128 & ~n_42129;
assign n_42131 = ~n_42127 &  n_42130;
assign n_42132 = ~n_42126 &  n_42131;
assign n_42133 = ~n_42125 &  n_42132;
assign n_42134 =  x_3696 & ~n_42133;
assign n_42135 = ~x_3696 &  n_42133;
assign n_42136 = ~n_42134 & ~n_42135;
assign n_42137 =  x_3695 &  n_42040;
assign n_42138 =  x_195 &  n_27857;
assign n_42139 =  x_2578 &  n_24036;
assign n_42140 =  x_1090 &  n_24005;
assign n_42141 =  x_3887 &  n_28297;
assign n_42142 = ~n_42140 & ~n_42141;
assign n_42143 = ~n_42139 &  n_42142;
assign n_42144 = ~n_42138 &  n_42143;
assign n_42145 = ~n_42137 &  n_42144;
assign n_42146 =  x_3695 & ~n_42145;
assign n_42147 = ~x_3695 &  n_42145;
assign n_42148 = ~n_42146 & ~n_42147;
assign n_42149 =  x_3694 &  n_42040;
assign n_42150 =  x_194 &  n_27857;
assign n_42151 =  x_2577 &  n_24036;
assign n_42152 =  x_1089 &  n_24005;
assign n_42153 =  x_3886 &  n_28297;
assign n_42154 = ~n_42152 & ~n_42153;
assign n_42155 = ~n_42151 &  n_42154;
assign n_42156 = ~n_42150 &  n_42155;
assign n_42157 = ~n_42149 &  n_42156;
assign n_42158 =  x_3694 & ~n_42157;
assign n_42159 = ~x_3694 &  n_42157;
assign n_42160 = ~n_42158 & ~n_42159;
assign n_42161 =  x_3693 &  n_42040;
assign n_42162 =  x_193 &  n_27857;
assign n_42163 =  x_2576 &  n_24036;
assign n_42164 =  x_1088 &  n_24005;
assign n_42165 =  x_3885 &  n_28297;
assign n_42166 = ~n_42164 & ~n_42165;
assign n_42167 = ~n_42163 &  n_42166;
assign n_42168 = ~n_42162 &  n_42167;
assign n_42169 = ~n_42161 &  n_42168;
assign n_42170 =  x_3693 & ~n_42169;
assign n_42171 = ~x_3693 &  n_42169;
assign n_42172 = ~n_42170 & ~n_42171;
assign n_42173 =  x_3692 &  n_42040;
assign n_42174 =  x_192 &  n_27857;
assign n_42175 =  x_2575 &  n_24036;
assign n_42176 =  x_1087 &  n_24005;
assign n_42177 =  x_3884 &  n_28297;
assign n_42178 = ~n_42176 & ~n_42177;
assign n_42179 = ~n_42175 &  n_42178;
assign n_42180 = ~n_42174 &  n_42179;
assign n_42181 = ~n_42173 &  n_42180;
assign n_42182 =  x_3692 & ~n_42181;
assign n_42183 = ~x_3692 &  n_42181;
assign n_42184 = ~n_42182 & ~n_42183;
assign n_42185 =  x_3691 &  n_42040;
assign n_42186 =  x_191 &  n_27857;
assign n_42187 =  x_2574 &  n_24036;
assign n_42188 =  x_1086 &  n_24005;
assign n_42189 =  x_3883 &  n_28297;
assign n_42190 = ~n_42188 & ~n_42189;
assign n_42191 = ~n_42187 &  n_42190;
assign n_42192 = ~n_42186 &  n_42191;
assign n_42193 = ~n_42185 &  n_42192;
assign n_42194 =  x_3691 & ~n_42193;
assign n_42195 = ~x_3691 &  n_42193;
assign n_42196 = ~n_42194 & ~n_42195;
assign n_42197 =  x_3690 &  n_42040;
assign n_42198 =  x_190 &  n_27857;
assign n_42199 =  x_2573 &  n_24036;
assign n_42200 =  x_1085 &  n_24005;
assign n_42201 =  x_3882 &  n_28297;
assign n_42202 = ~n_42200 & ~n_42201;
assign n_42203 = ~n_42199 &  n_42202;
assign n_42204 = ~n_42198 &  n_42203;
assign n_42205 = ~n_42197 &  n_42204;
assign n_42206 =  x_3690 & ~n_42205;
assign n_42207 = ~x_3690 &  n_42205;
assign n_42208 = ~n_42206 & ~n_42207;
assign n_42209 =  x_3689 &  n_42040;
assign n_42210 =  x_189 &  n_27857;
assign n_42211 =  x_2572 &  n_24036;
assign n_42212 =  x_1084 &  n_24005;
assign n_42213 =  x_3881 &  n_28297;
assign n_42214 = ~n_42212 & ~n_42213;
assign n_42215 = ~n_42211 &  n_42214;
assign n_42216 = ~n_42210 &  n_42215;
assign n_42217 = ~n_42209 &  n_42216;
assign n_42218 =  x_3689 & ~n_42217;
assign n_42219 = ~x_3689 &  n_42217;
assign n_42220 = ~n_42218 & ~n_42219;
assign n_42221 =  x_3688 &  n_42040;
assign n_42222 =  x_188 &  n_27857;
assign n_42223 =  x_2571 &  n_24036;
assign n_42224 =  x_1083 &  n_24005;
assign n_42225 =  x_3880 &  n_28297;
assign n_42226 = ~n_42224 & ~n_42225;
assign n_42227 = ~n_42223 &  n_42226;
assign n_42228 = ~n_42222 &  n_42227;
assign n_42229 = ~n_42221 &  n_42228;
assign n_42230 =  x_3688 & ~n_42229;
assign n_42231 = ~x_3688 &  n_42229;
assign n_42232 = ~n_42230 & ~n_42231;
assign n_42233 =  x_3687 &  n_42040;
assign n_42234 =  x_187 &  n_27857;
assign n_42235 =  x_2570 &  n_24036;
assign n_42236 =  x_1082 &  n_24005;
assign n_42237 =  x_3879 &  n_28297;
assign n_42238 = ~n_42236 & ~n_42237;
assign n_42239 = ~n_42235 &  n_42238;
assign n_42240 = ~n_42234 &  n_42239;
assign n_42241 = ~n_42233 &  n_42240;
assign n_42242 =  x_3687 & ~n_42241;
assign n_42243 = ~x_3687 &  n_42241;
assign n_42244 = ~n_42242 & ~n_42243;
assign n_42245 =  x_3686 &  n_42040;
assign n_42246 =  x_186 &  n_27857;
assign n_42247 =  x_2569 &  n_24036;
assign n_42248 =  x_1081 &  n_24005;
assign n_42249 =  x_3878 &  n_28297;
assign n_42250 = ~n_42248 & ~n_42249;
assign n_42251 = ~n_42247 &  n_42250;
assign n_42252 = ~n_42246 &  n_42251;
assign n_42253 = ~n_42245 &  n_42252;
assign n_42254 =  x_3686 & ~n_42253;
assign n_42255 = ~x_3686 &  n_42253;
assign n_42256 = ~n_42254 & ~n_42255;
assign n_42257 =  x_3685 &  n_42040;
assign n_42258 =  x_185 &  n_27857;
assign n_42259 =  x_2568 &  n_24036;
assign n_42260 =  x_1080 &  n_24005;
assign n_42261 =  x_3877 &  n_28297;
assign n_42262 = ~n_42260 & ~n_42261;
assign n_42263 = ~n_42259 &  n_42262;
assign n_42264 = ~n_42258 &  n_42263;
assign n_42265 = ~n_42257 &  n_42264;
assign n_42266 =  x_3685 & ~n_42265;
assign n_42267 = ~x_3685 &  n_42265;
assign n_42268 = ~n_42266 & ~n_42267;
assign n_42269 =  x_3684 &  n_42040;
assign n_42270 =  x_184 &  n_27857;
assign n_42271 =  x_2567 &  n_24036;
assign n_42272 =  x_1079 &  n_24005;
assign n_42273 =  x_3876 &  n_28297;
assign n_42274 = ~n_42272 & ~n_42273;
assign n_42275 = ~n_42271 &  n_42274;
assign n_42276 = ~n_42270 &  n_42275;
assign n_42277 = ~n_42269 &  n_42276;
assign n_42278 =  x_3684 & ~n_42277;
assign n_42279 = ~x_3684 &  n_42277;
assign n_42280 = ~n_42278 & ~n_42279;
assign n_42281 =  x_3683 &  n_42040;
assign n_42282 =  x_183 &  n_27857;
assign n_42283 =  x_2566 &  n_24036;
assign n_42284 =  x_1078 &  n_24005;
assign n_42285 =  x_3875 &  n_28297;
assign n_42286 = ~n_42284 & ~n_42285;
assign n_42287 = ~n_42283 &  n_42286;
assign n_42288 = ~n_42282 &  n_42287;
assign n_42289 = ~n_42281 &  n_42288;
assign n_42290 =  x_3683 & ~n_42289;
assign n_42291 = ~x_3683 &  n_42289;
assign n_42292 = ~n_42290 & ~n_42291;
assign n_42293 =  x_3682 &  n_42040;
assign n_42294 =  x_182 &  n_27857;
assign n_42295 =  x_2565 &  n_24036;
assign n_42296 =  x_1077 &  n_24005;
assign n_42297 =  x_3874 &  n_28297;
assign n_42298 = ~n_42296 & ~n_42297;
assign n_42299 = ~n_42295 &  n_42298;
assign n_42300 = ~n_42294 &  n_42299;
assign n_42301 = ~n_42293 &  n_42300;
assign n_42302 =  x_3682 & ~n_42301;
assign n_42303 = ~x_3682 &  n_42301;
assign n_42304 = ~n_42302 & ~n_42303;
assign n_42305 =  x_3681 &  n_42040;
assign n_42306 =  x_181 &  n_27857;
assign n_42307 =  x_2564 &  n_24036;
assign n_42308 =  x_1076 &  n_24005;
assign n_42309 =  x_3873 &  n_28297;
assign n_42310 = ~n_42308 & ~n_42309;
assign n_42311 = ~n_42307 &  n_42310;
assign n_42312 = ~n_42306 &  n_42311;
assign n_42313 = ~n_42305 &  n_42312;
assign n_42314 =  x_3681 & ~n_42313;
assign n_42315 = ~x_3681 &  n_42313;
assign n_42316 = ~n_42314 & ~n_42315;
assign n_42317 =  x_3680 &  n_42040;
assign n_42318 =  x_180 &  n_27857;
assign n_42319 =  x_2563 &  n_24036;
assign n_42320 =  x_1075 &  n_24005;
assign n_42321 =  x_3872 &  n_28297;
assign n_42322 = ~n_42320 & ~n_42321;
assign n_42323 = ~n_42319 &  n_42322;
assign n_42324 = ~n_42318 &  n_42323;
assign n_42325 = ~n_42317 &  n_42324;
assign n_42326 =  x_3680 & ~n_42325;
assign n_42327 = ~x_3680 &  n_42325;
assign n_42328 = ~n_42326 & ~n_42327;
assign n_42329 =  x_3679 &  n_42040;
assign n_42330 =  x_179 &  n_27857;
assign n_42331 =  x_2562 &  n_24036;
assign n_42332 =  x_1074 &  n_24005;
assign n_42333 =  x_3871 &  n_28297;
assign n_42334 = ~n_42332 & ~n_42333;
assign n_42335 = ~n_42331 &  n_42334;
assign n_42336 = ~n_42330 &  n_42335;
assign n_42337 = ~n_42329 &  n_42336;
assign n_42338 =  x_3679 & ~n_42337;
assign n_42339 = ~x_3679 &  n_42337;
assign n_42340 = ~n_42338 & ~n_42339;
assign n_42341 =  x_3678 &  n_42040;
assign n_42342 =  x_178 &  n_27857;
assign n_42343 =  x_2561 &  n_24036;
assign n_42344 =  x_1073 &  n_24005;
assign n_42345 =  x_3870 &  n_28297;
assign n_42346 = ~n_42344 & ~n_42345;
assign n_42347 = ~n_42343 &  n_42346;
assign n_42348 = ~n_42342 &  n_42347;
assign n_42349 = ~n_42341 &  n_42348;
assign n_42350 =  x_3678 & ~n_42349;
assign n_42351 = ~x_3678 &  n_42349;
assign n_42352 = ~n_42350 & ~n_42351;
assign n_42353 =  x_3677 &  n_42040;
assign n_42354 =  x_177 &  n_27857;
assign n_42355 =  x_2560 &  n_24036;
assign n_42356 =  x_1072 &  n_24005;
assign n_42357 =  x_3869 &  n_28297;
assign n_42358 = ~n_42356 & ~n_42357;
assign n_42359 = ~n_42355 &  n_42358;
assign n_42360 = ~n_42354 &  n_42359;
assign n_42361 = ~n_42353 &  n_42360;
assign n_42362 =  x_3677 & ~n_42361;
assign n_42363 = ~x_3677 &  n_42361;
assign n_42364 = ~n_42362 & ~n_42363;
assign n_42365 =  x_3676 &  n_42040;
assign n_42366 =  x_176 &  n_27857;
assign n_42367 =  x_2559 &  n_24036;
assign n_42368 =  x_1071 &  n_24005;
assign n_42369 =  x_3868 &  n_28297;
assign n_42370 = ~n_42368 & ~n_42369;
assign n_42371 = ~n_42367 &  n_42370;
assign n_42372 = ~n_42366 &  n_42371;
assign n_42373 = ~n_42365 &  n_42372;
assign n_42374 =  x_3676 & ~n_42373;
assign n_42375 = ~x_3676 &  n_42373;
assign n_42376 = ~n_42374 & ~n_42375;
assign n_42377 =  x_3675 &  n_42040;
assign n_42378 =  x_175 &  n_27857;
assign n_42379 =  x_2558 &  n_24036;
assign n_42380 =  x_1070 &  n_24005;
assign n_42381 =  x_3867 &  n_28297;
assign n_42382 = ~n_42380 & ~n_42381;
assign n_42383 = ~n_42379 &  n_42382;
assign n_42384 = ~n_42378 &  n_42383;
assign n_42385 = ~n_42377 &  n_42384;
assign n_42386 =  x_3675 & ~n_42385;
assign n_42387 = ~x_3675 &  n_42385;
assign n_42388 = ~n_42386 & ~n_42387;
assign n_42389 =  x_3674 &  n_42040;
assign n_42390 =  x_174 &  n_27857;
assign n_42391 =  x_2557 &  n_24036;
assign n_42392 =  x_1069 &  n_24005;
assign n_42393 =  x_3866 &  n_28297;
assign n_42394 = ~n_42392 & ~n_42393;
assign n_42395 = ~n_42391 &  n_42394;
assign n_42396 = ~n_42390 &  n_42395;
assign n_42397 = ~n_42389 &  n_42396;
assign n_42398 =  x_3674 & ~n_42397;
assign n_42399 = ~x_3674 &  n_42397;
assign n_42400 = ~n_42398 & ~n_42399;
assign n_42401 =  x_3673 &  n_42040;
assign n_42402 =  x_173 &  n_27857;
assign n_42403 =  x_2556 &  n_24036;
assign n_42404 =  x_1068 &  n_24005;
assign n_42405 =  x_3865 &  n_28297;
assign n_42406 = ~n_42404 & ~n_42405;
assign n_42407 = ~n_42403 &  n_42406;
assign n_42408 = ~n_42402 &  n_42407;
assign n_42409 = ~n_42401 &  n_42408;
assign n_42410 =  x_3673 & ~n_42409;
assign n_42411 = ~x_3673 &  n_42409;
assign n_42412 = ~n_42410 & ~n_42411;
assign n_42413 =  x_3672 &  n_42040;
assign n_42414 =  x_172 &  n_27857;
assign n_42415 =  x_2555 &  n_24036;
assign n_42416 =  x_1067 &  n_24005;
assign n_42417 =  x_3864 &  n_28297;
assign n_42418 = ~n_42416 & ~n_42417;
assign n_42419 = ~n_42415 &  n_42418;
assign n_42420 = ~n_42414 &  n_42419;
assign n_42421 = ~n_42413 &  n_42420;
assign n_42422 =  x_3672 & ~n_42421;
assign n_42423 = ~x_3672 &  n_42421;
assign n_42424 = ~n_42422 & ~n_42423;
assign n_42425 = ~n_26345 & ~n_25980;
assign n_42426 = ~n_26261 &  n_42425;
assign n_42427 = ~n_26368 & ~n_26071;
assign n_42428 = ~n_26171 &  n_42427;
assign n_42429 = ~n_28790 &  n_42428;
assign n_42430 =  n_42426 &  n_42429;
assign n_42431 =  x_3671 &  n_42430;
assign n_42432 =  i_32 & ~n_42426;
assign n_42433 =  x_3607 &  n_26171;
assign n_42434 =  x_4328 &  n_28790;
assign n_42435 =  x_3575 &  n_26368;
assign n_42436 =  x_4360 &  n_26071;
assign n_42437 = ~n_42435 & ~n_42436;
assign n_42438 = ~n_42434 &  n_42437;
assign n_42439 = ~n_42433 &  n_42438;
assign n_42440 = ~n_42432 &  n_42439;
assign n_42441 = ~n_42431 &  n_42440;
assign n_42442 =  x_3671 & ~n_42441;
assign n_42443 = ~x_3671 &  n_42441;
assign n_42444 = ~n_42442 & ~n_42443;
assign n_42445 =  x_3670 &  n_42430;
assign n_42446 =  i_31 & ~n_42426;
assign n_42447 =  x_3606 &  n_26171;
assign n_42448 =  x_4327 &  n_28790;
assign n_42449 =  x_3574 &  n_26368;
assign n_42450 =  x_4359 &  n_26071;
assign n_42451 = ~n_42449 & ~n_42450;
assign n_42452 = ~n_42448 &  n_42451;
assign n_42453 = ~n_42447 &  n_42452;
assign n_42454 = ~n_42446 &  n_42453;
assign n_42455 = ~n_42445 &  n_42454;
assign n_42456 =  x_3670 & ~n_42455;
assign n_42457 = ~x_3670 &  n_42455;
assign n_42458 = ~n_42456 & ~n_42457;
assign n_42459 =  x_3669 &  n_42430;
assign n_42460 =  i_30 & ~n_42426;
assign n_42461 =  x_3605 &  n_26171;
assign n_42462 =  x_4326 &  n_28790;
assign n_42463 =  x_3573 &  n_26368;
assign n_42464 =  x_4358 &  n_26071;
assign n_42465 = ~n_42463 & ~n_42464;
assign n_42466 = ~n_42462 &  n_42465;
assign n_42467 = ~n_42461 &  n_42466;
assign n_42468 = ~n_42460 &  n_42467;
assign n_42469 = ~n_42459 &  n_42468;
assign n_42470 =  x_3669 & ~n_42469;
assign n_42471 = ~x_3669 &  n_42469;
assign n_42472 = ~n_42470 & ~n_42471;
assign n_42473 =  x_3668 &  n_42430;
assign n_42474 =  i_29 & ~n_42426;
assign n_42475 =  x_3604 &  n_26171;
assign n_42476 =  x_4325 &  n_28790;
assign n_42477 =  x_3572 &  n_26368;
assign n_42478 =  x_4357 &  n_26071;
assign n_42479 = ~n_42477 & ~n_42478;
assign n_42480 = ~n_42476 &  n_42479;
assign n_42481 = ~n_42475 &  n_42480;
assign n_42482 = ~n_42474 &  n_42481;
assign n_42483 = ~n_42473 &  n_42482;
assign n_42484 =  x_3668 & ~n_42483;
assign n_42485 = ~x_3668 &  n_42483;
assign n_42486 = ~n_42484 & ~n_42485;
assign n_42487 =  x_3667 &  n_42430;
assign n_42488 =  i_28 & ~n_42426;
assign n_42489 =  x_3603 &  n_26171;
assign n_42490 =  x_4324 &  n_28790;
assign n_42491 =  x_3571 &  n_26368;
assign n_42492 =  x_4356 &  n_26071;
assign n_42493 = ~n_42491 & ~n_42492;
assign n_42494 = ~n_42490 &  n_42493;
assign n_42495 = ~n_42489 &  n_42494;
assign n_42496 = ~n_42488 &  n_42495;
assign n_42497 = ~n_42487 &  n_42496;
assign n_42498 =  x_3667 & ~n_42497;
assign n_42499 = ~x_3667 &  n_42497;
assign n_42500 = ~n_42498 & ~n_42499;
assign n_42501 =  x_3666 &  n_42430;
assign n_42502 =  i_27 & ~n_42426;
assign n_42503 =  x_3602 &  n_26171;
assign n_42504 =  x_4323 &  n_28790;
assign n_42505 =  x_3570 &  n_26368;
assign n_42506 =  x_4355 &  n_26071;
assign n_42507 = ~n_42505 & ~n_42506;
assign n_42508 = ~n_42504 &  n_42507;
assign n_42509 = ~n_42503 &  n_42508;
assign n_42510 = ~n_42502 &  n_42509;
assign n_42511 = ~n_42501 &  n_42510;
assign n_42512 =  x_3666 & ~n_42511;
assign n_42513 = ~x_3666 &  n_42511;
assign n_42514 = ~n_42512 & ~n_42513;
assign n_42515 =  x_3665 &  n_42430;
assign n_42516 =  i_26 & ~n_42426;
assign n_42517 =  x_3601 &  n_26171;
assign n_42518 =  x_4322 &  n_28790;
assign n_42519 =  x_3569 &  n_26368;
assign n_42520 =  x_4354 &  n_26071;
assign n_42521 = ~n_42519 & ~n_42520;
assign n_42522 = ~n_42518 &  n_42521;
assign n_42523 = ~n_42517 &  n_42522;
assign n_42524 = ~n_42516 &  n_42523;
assign n_42525 = ~n_42515 &  n_42524;
assign n_42526 =  x_3665 & ~n_42525;
assign n_42527 = ~x_3665 &  n_42525;
assign n_42528 = ~n_42526 & ~n_42527;
assign n_42529 =  x_3664 &  n_42430;
assign n_42530 =  i_25 & ~n_42426;
assign n_42531 =  x_3600 &  n_26171;
assign n_42532 =  x_4321 &  n_28790;
assign n_42533 =  x_3568 &  n_26368;
assign n_42534 =  x_4353 &  n_26071;
assign n_42535 = ~n_42533 & ~n_42534;
assign n_42536 = ~n_42532 &  n_42535;
assign n_42537 = ~n_42531 &  n_42536;
assign n_42538 = ~n_42530 &  n_42537;
assign n_42539 = ~n_42529 &  n_42538;
assign n_42540 =  x_3664 & ~n_42539;
assign n_42541 = ~x_3664 &  n_42539;
assign n_42542 = ~n_42540 & ~n_42541;
assign n_42543 =  x_3663 &  n_42430;
assign n_42544 =  i_24 & ~n_42426;
assign n_42545 =  x_3599 &  n_26171;
assign n_42546 =  x_4320 &  n_28790;
assign n_42547 =  x_3567 &  n_26368;
assign n_42548 =  x_4352 &  n_26071;
assign n_42549 = ~n_42547 & ~n_42548;
assign n_42550 = ~n_42546 &  n_42549;
assign n_42551 = ~n_42545 &  n_42550;
assign n_42552 = ~n_42544 &  n_42551;
assign n_42553 = ~n_42543 &  n_42552;
assign n_42554 =  x_3663 & ~n_42553;
assign n_42555 = ~x_3663 &  n_42553;
assign n_42556 = ~n_42554 & ~n_42555;
assign n_42557 =  x_3662 &  n_42430;
assign n_42558 =  i_23 & ~n_42426;
assign n_42559 =  x_3598 &  n_26171;
assign n_42560 =  x_4319 &  n_28790;
assign n_42561 =  x_3566 &  n_26368;
assign n_42562 =  x_4351 &  n_26071;
assign n_42563 = ~n_42561 & ~n_42562;
assign n_42564 = ~n_42560 &  n_42563;
assign n_42565 = ~n_42559 &  n_42564;
assign n_42566 = ~n_42558 &  n_42565;
assign n_42567 = ~n_42557 &  n_42566;
assign n_42568 =  x_3662 & ~n_42567;
assign n_42569 = ~x_3662 &  n_42567;
assign n_42570 = ~n_42568 & ~n_42569;
assign n_42571 =  x_3661 &  n_42430;
assign n_42572 =  i_22 & ~n_42426;
assign n_42573 =  x_3597 &  n_26171;
assign n_42574 =  x_4318 &  n_28790;
assign n_42575 =  x_3565 &  n_26368;
assign n_42576 =  x_4350 &  n_26071;
assign n_42577 = ~n_42575 & ~n_42576;
assign n_42578 = ~n_42574 &  n_42577;
assign n_42579 = ~n_42573 &  n_42578;
assign n_42580 = ~n_42572 &  n_42579;
assign n_42581 = ~n_42571 &  n_42580;
assign n_42582 =  x_3661 & ~n_42581;
assign n_42583 = ~x_3661 &  n_42581;
assign n_42584 = ~n_42582 & ~n_42583;
assign n_42585 =  x_3660 &  n_42430;
assign n_42586 =  i_21 & ~n_42426;
assign n_42587 =  x_3596 &  n_26171;
assign n_42588 =  x_4317 &  n_28790;
assign n_42589 =  x_3564 &  n_26368;
assign n_42590 =  x_4349 &  n_26071;
assign n_42591 = ~n_42589 & ~n_42590;
assign n_42592 = ~n_42588 &  n_42591;
assign n_42593 = ~n_42587 &  n_42592;
assign n_42594 = ~n_42586 &  n_42593;
assign n_42595 = ~n_42585 &  n_42594;
assign n_42596 =  x_3660 & ~n_42595;
assign n_42597 = ~x_3660 &  n_42595;
assign n_42598 = ~n_42596 & ~n_42597;
assign n_42599 =  x_3659 &  n_42430;
assign n_42600 =  i_20 & ~n_42426;
assign n_42601 =  x_3595 &  n_26171;
assign n_42602 =  x_4316 &  n_28790;
assign n_42603 =  x_3563 &  n_26368;
assign n_42604 =  x_4348 &  n_26071;
assign n_42605 = ~n_42603 & ~n_42604;
assign n_42606 = ~n_42602 &  n_42605;
assign n_42607 = ~n_42601 &  n_42606;
assign n_42608 = ~n_42600 &  n_42607;
assign n_42609 = ~n_42599 &  n_42608;
assign n_42610 =  x_3659 & ~n_42609;
assign n_42611 = ~x_3659 &  n_42609;
assign n_42612 = ~n_42610 & ~n_42611;
assign n_42613 =  x_3658 &  n_42430;
assign n_42614 =  i_19 & ~n_42426;
assign n_42615 =  x_3594 &  n_26171;
assign n_42616 =  x_4315 &  n_28790;
assign n_42617 =  x_3562 &  n_26368;
assign n_42618 =  x_4347 &  n_26071;
assign n_42619 = ~n_42617 & ~n_42618;
assign n_42620 = ~n_42616 &  n_42619;
assign n_42621 = ~n_42615 &  n_42620;
assign n_42622 = ~n_42614 &  n_42621;
assign n_42623 = ~n_42613 &  n_42622;
assign n_42624 =  x_3658 & ~n_42623;
assign n_42625 = ~x_3658 &  n_42623;
assign n_42626 = ~n_42624 & ~n_42625;
assign n_42627 =  x_3657 &  n_42430;
assign n_42628 =  i_18 & ~n_42426;
assign n_42629 =  x_3593 &  n_26171;
assign n_42630 =  x_4314 &  n_28790;
assign n_42631 =  x_3561 &  n_26368;
assign n_42632 =  x_4346 &  n_26071;
assign n_42633 = ~n_42631 & ~n_42632;
assign n_42634 = ~n_42630 &  n_42633;
assign n_42635 = ~n_42629 &  n_42634;
assign n_42636 = ~n_42628 &  n_42635;
assign n_42637 = ~n_42627 &  n_42636;
assign n_42638 =  x_3657 & ~n_42637;
assign n_42639 = ~x_3657 &  n_42637;
assign n_42640 = ~n_42638 & ~n_42639;
assign n_42641 =  x_3656 &  n_42430;
assign n_42642 =  i_17 & ~n_42426;
assign n_42643 =  x_3592 &  n_26171;
assign n_42644 =  x_4313 &  n_28790;
assign n_42645 =  x_3560 &  n_26368;
assign n_42646 =  x_4345 &  n_26071;
assign n_42647 = ~n_42645 & ~n_42646;
assign n_42648 = ~n_42644 &  n_42647;
assign n_42649 = ~n_42643 &  n_42648;
assign n_42650 = ~n_42642 &  n_42649;
assign n_42651 = ~n_42641 &  n_42650;
assign n_42652 =  x_3656 & ~n_42651;
assign n_42653 = ~x_3656 &  n_42651;
assign n_42654 = ~n_42652 & ~n_42653;
assign n_42655 =  x_3655 &  n_42430;
assign n_42656 =  i_16 & ~n_42426;
assign n_42657 =  x_3591 &  n_26171;
assign n_42658 =  x_4312 &  n_28790;
assign n_42659 =  x_3559 &  n_26368;
assign n_42660 =  x_4344 &  n_26071;
assign n_42661 = ~n_42659 & ~n_42660;
assign n_42662 = ~n_42658 &  n_42661;
assign n_42663 = ~n_42657 &  n_42662;
assign n_42664 = ~n_42656 &  n_42663;
assign n_42665 = ~n_42655 &  n_42664;
assign n_42666 =  x_3655 & ~n_42665;
assign n_42667 = ~x_3655 &  n_42665;
assign n_42668 = ~n_42666 & ~n_42667;
assign n_42669 =  x_3654 &  n_42430;
assign n_42670 =  i_15 & ~n_42426;
assign n_42671 =  x_3590 &  n_26171;
assign n_42672 =  x_4311 &  n_28790;
assign n_42673 =  x_3558 &  n_26368;
assign n_42674 =  x_4343 &  n_26071;
assign n_42675 = ~n_42673 & ~n_42674;
assign n_42676 = ~n_42672 &  n_42675;
assign n_42677 = ~n_42671 &  n_42676;
assign n_42678 = ~n_42670 &  n_42677;
assign n_42679 = ~n_42669 &  n_42678;
assign n_42680 =  x_3654 & ~n_42679;
assign n_42681 = ~x_3654 &  n_42679;
assign n_42682 = ~n_42680 & ~n_42681;
assign n_42683 =  x_3653 &  n_42430;
assign n_42684 =  i_14 & ~n_42426;
assign n_42685 =  x_3589 &  n_26171;
assign n_42686 =  x_4310 &  n_28790;
assign n_42687 =  x_3557 &  n_26368;
assign n_42688 =  x_4342 &  n_26071;
assign n_42689 = ~n_42687 & ~n_42688;
assign n_42690 = ~n_42686 &  n_42689;
assign n_42691 = ~n_42685 &  n_42690;
assign n_42692 = ~n_42684 &  n_42691;
assign n_42693 = ~n_42683 &  n_42692;
assign n_42694 =  x_3653 & ~n_42693;
assign n_42695 = ~x_3653 &  n_42693;
assign n_42696 = ~n_42694 & ~n_42695;
assign n_42697 =  x_3652 &  n_42430;
assign n_42698 =  i_13 & ~n_42426;
assign n_42699 =  x_3588 &  n_26171;
assign n_42700 =  x_4309 &  n_28790;
assign n_42701 =  x_3556 &  n_26368;
assign n_42702 =  x_4341 &  n_26071;
assign n_42703 = ~n_42701 & ~n_42702;
assign n_42704 = ~n_42700 &  n_42703;
assign n_42705 = ~n_42699 &  n_42704;
assign n_42706 = ~n_42698 &  n_42705;
assign n_42707 = ~n_42697 &  n_42706;
assign n_42708 =  x_3652 & ~n_42707;
assign n_42709 = ~x_3652 &  n_42707;
assign n_42710 = ~n_42708 & ~n_42709;
assign n_42711 =  x_3651 &  n_42430;
assign n_42712 =  i_12 & ~n_42426;
assign n_42713 =  x_3587 &  n_26171;
assign n_42714 =  x_4308 &  n_28790;
assign n_42715 =  x_3555 &  n_26368;
assign n_42716 =  x_4340 &  n_26071;
assign n_42717 = ~n_42715 & ~n_42716;
assign n_42718 = ~n_42714 &  n_42717;
assign n_42719 = ~n_42713 &  n_42718;
assign n_42720 = ~n_42712 &  n_42719;
assign n_42721 = ~n_42711 &  n_42720;
assign n_42722 =  x_3651 & ~n_42721;
assign n_42723 = ~x_3651 &  n_42721;
assign n_42724 = ~n_42722 & ~n_42723;
assign n_42725 =  x_3650 &  n_42430;
assign n_42726 =  i_11 & ~n_42426;
assign n_42727 =  x_3586 &  n_26171;
assign n_42728 =  x_4307 &  n_28790;
assign n_42729 =  x_3554 &  n_26368;
assign n_42730 =  x_4339 &  n_26071;
assign n_42731 = ~n_42729 & ~n_42730;
assign n_42732 = ~n_42728 &  n_42731;
assign n_42733 = ~n_42727 &  n_42732;
assign n_42734 = ~n_42726 &  n_42733;
assign n_42735 = ~n_42725 &  n_42734;
assign n_42736 =  x_3650 & ~n_42735;
assign n_42737 = ~x_3650 &  n_42735;
assign n_42738 = ~n_42736 & ~n_42737;
assign n_42739 =  x_3649 &  n_42430;
assign n_42740 =  i_10 & ~n_42426;
assign n_42741 =  x_3585 &  n_26171;
assign n_42742 =  x_4306 &  n_28790;
assign n_42743 =  x_3553 &  n_26368;
assign n_42744 =  x_4338 &  n_26071;
assign n_42745 = ~n_42743 & ~n_42744;
assign n_42746 = ~n_42742 &  n_42745;
assign n_42747 = ~n_42741 &  n_42746;
assign n_42748 = ~n_42740 &  n_42747;
assign n_42749 = ~n_42739 &  n_42748;
assign n_42750 =  x_3649 & ~n_42749;
assign n_42751 = ~x_3649 &  n_42749;
assign n_42752 = ~n_42750 & ~n_42751;
assign n_42753 =  x_3648 &  n_42430;
assign n_42754 =  i_9 & ~n_42426;
assign n_42755 =  x_3584 &  n_26171;
assign n_42756 =  x_4305 &  n_28790;
assign n_42757 =  x_3552 &  n_26368;
assign n_42758 =  x_4337 &  n_26071;
assign n_42759 = ~n_42757 & ~n_42758;
assign n_42760 = ~n_42756 &  n_42759;
assign n_42761 = ~n_42755 &  n_42760;
assign n_42762 = ~n_42754 &  n_42761;
assign n_42763 = ~n_42753 &  n_42762;
assign n_42764 =  x_3648 & ~n_42763;
assign n_42765 = ~x_3648 &  n_42763;
assign n_42766 = ~n_42764 & ~n_42765;
assign n_42767 =  x_3647 &  n_42430;
assign n_42768 =  i_8 & ~n_42426;
assign n_42769 =  x_3583 &  n_26171;
assign n_42770 =  x_4304 &  n_28790;
assign n_42771 =  x_3551 &  n_26368;
assign n_42772 =  x_4336 &  n_26071;
assign n_42773 = ~n_42771 & ~n_42772;
assign n_42774 = ~n_42770 &  n_42773;
assign n_42775 = ~n_42769 &  n_42774;
assign n_42776 = ~n_42768 &  n_42775;
assign n_42777 = ~n_42767 &  n_42776;
assign n_42778 =  x_3647 & ~n_42777;
assign n_42779 = ~x_3647 &  n_42777;
assign n_42780 = ~n_42778 & ~n_42779;
assign n_42781 =  x_3646 &  n_42430;
assign n_42782 =  i_7 & ~n_42426;
assign n_42783 =  x_3582 &  n_26171;
assign n_42784 =  x_4303 &  n_28790;
assign n_42785 =  x_3550 &  n_26368;
assign n_42786 =  x_4335 &  n_26071;
assign n_42787 = ~n_42785 & ~n_42786;
assign n_42788 = ~n_42784 &  n_42787;
assign n_42789 = ~n_42783 &  n_42788;
assign n_42790 = ~n_42782 &  n_42789;
assign n_42791 = ~n_42781 &  n_42790;
assign n_42792 =  x_3646 & ~n_42791;
assign n_42793 = ~x_3646 &  n_42791;
assign n_42794 = ~n_42792 & ~n_42793;
assign n_42795 =  x_3645 &  n_42430;
assign n_42796 =  i_6 & ~n_42426;
assign n_42797 =  x_3581 &  n_26171;
assign n_42798 =  x_4302 &  n_28790;
assign n_42799 =  x_3549 &  n_26368;
assign n_42800 =  x_4334 &  n_26071;
assign n_42801 = ~n_42799 & ~n_42800;
assign n_42802 = ~n_42798 &  n_42801;
assign n_42803 = ~n_42797 &  n_42802;
assign n_42804 = ~n_42796 &  n_42803;
assign n_42805 = ~n_42795 &  n_42804;
assign n_42806 =  x_3645 & ~n_42805;
assign n_42807 = ~x_3645 &  n_42805;
assign n_42808 = ~n_42806 & ~n_42807;
assign n_42809 =  x_3644 &  n_42430;
assign n_42810 =  i_5 & ~n_42426;
assign n_42811 =  x_3580 &  n_26171;
assign n_42812 =  x_4301 &  n_28790;
assign n_42813 =  x_3548 &  n_26368;
assign n_42814 =  x_4333 &  n_26071;
assign n_42815 = ~n_42813 & ~n_42814;
assign n_42816 = ~n_42812 &  n_42815;
assign n_42817 = ~n_42811 &  n_42816;
assign n_42818 = ~n_42810 &  n_42817;
assign n_42819 = ~n_42809 &  n_42818;
assign n_42820 =  x_3644 & ~n_42819;
assign n_42821 = ~x_3644 &  n_42819;
assign n_42822 = ~n_42820 & ~n_42821;
assign n_42823 =  x_3643 &  n_42430;
assign n_42824 =  i_4 & ~n_42426;
assign n_42825 =  x_3579 &  n_26171;
assign n_42826 =  x_4300 &  n_28790;
assign n_42827 =  x_3547 &  n_26368;
assign n_42828 =  x_4332 &  n_26071;
assign n_42829 = ~n_42827 & ~n_42828;
assign n_42830 = ~n_42826 &  n_42829;
assign n_42831 = ~n_42825 &  n_42830;
assign n_42832 = ~n_42824 &  n_42831;
assign n_42833 = ~n_42823 &  n_42832;
assign n_42834 =  x_3643 & ~n_42833;
assign n_42835 = ~x_3643 &  n_42833;
assign n_42836 = ~n_42834 & ~n_42835;
assign n_42837 =  x_3642 &  n_42430;
assign n_42838 =  i_3 & ~n_42426;
assign n_42839 =  x_3578 &  n_26171;
assign n_42840 =  x_4299 &  n_28790;
assign n_42841 =  x_3546 &  n_26368;
assign n_42842 =  x_4331 &  n_26071;
assign n_42843 = ~n_42841 & ~n_42842;
assign n_42844 = ~n_42840 &  n_42843;
assign n_42845 = ~n_42839 &  n_42844;
assign n_42846 = ~n_42838 &  n_42845;
assign n_42847 = ~n_42837 &  n_42846;
assign n_42848 =  x_3642 & ~n_42847;
assign n_42849 = ~x_3642 &  n_42847;
assign n_42850 = ~n_42848 & ~n_42849;
assign n_42851 =  x_3641 &  n_42430;
assign n_42852 =  i_2 & ~n_42426;
assign n_42853 =  x_3577 &  n_26171;
assign n_42854 =  x_4298 &  n_28790;
assign n_42855 =  x_3545 &  n_26368;
assign n_42856 =  x_4330 &  n_26071;
assign n_42857 = ~n_42855 & ~n_42856;
assign n_42858 = ~n_42854 &  n_42857;
assign n_42859 = ~n_42853 &  n_42858;
assign n_42860 = ~n_42852 &  n_42859;
assign n_42861 = ~n_42851 &  n_42860;
assign n_42862 =  x_3641 & ~n_42861;
assign n_42863 = ~x_3641 &  n_42861;
assign n_42864 = ~n_42862 & ~n_42863;
assign n_42865 =  x_3640 &  n_42430;
assign n_42866 =  i_1 & ~n_42426;
assign n_42867 =  x_3576 &  n_26171;
assign n_42868 =  x_4297 &  n_28790;
assign n_42869 =  x_3544 &  n_26368;
assign n_42870 =  x_4329 &  n_26071;
assign n_42871 = ~n_42869 & ~n_42870;
assign n_42872 = ~n_42868 &  n_42871;
assign n_42873 = ~n_42867 &  n_42872;
assign n_42874 = ~n_42866 &  n_42873;
assign n_42875 = ~n_42865 &  n_42874;
assign n_42876 =  x_3640 & ~n_42875;
assign n_42877 = ~x_3640 &  n_42875;
assign n_42878 = ~n_42876 & ~n_42877;
assign n_42879 =  n_25638 & ~n_14801;
assign n_42880 =  x_3639 & ~n_25638;
assign n_42881 = ~n_42879 & ~n_42880;
assign n_42882 =  x_3639 & ~n_42881;
assign n_42883 = ~x_3639 &  n_42881;
assign n_42884 = ~n_42882 & ~n_42883;
assign n_42885 =  n_25638 & ~n_14819;
assign n_42886 =  x_3638 & ~n_25638;
assign n_42887 = ~n_42885 & ~n_42886;
assign n_42888 =  x_3638 & ~n_42887;
assign n_42889 = ~x_3638 &  n_42887;
assign n_42890 = ~n_42888 & ~n_42889;
assign n_42891 =  n_25638 & ~n_14837;
assign n_42892 =  x_3637 & ~n_25638;
assign n_42893 = ~n_42891 & ~n_42892;
assign n_42894 =  x_3637 & ~n_42893;
assign n_42895 = ~x_3637 &  n_42893;
assign n_42896 = ~n_42894 & ~n_42895;
assign n_42897 =  n_25638 & ~n_14855;
assign n_42898 =  x_3636 & ~n_25638;
assign n_42899 = ~n_42897 & ~n_42898;
assign n_42900 =  x_3636 & ~n_42899;
assign n_42901 = ~x_3636 &  n_42899;
assign n_42902 = ~n_42900 & ~n_42901;
assign n_42903 =  n_25638 & ~n_14873;
assign n_42904 =  x_3635 & ~n_25638;
assign n_42905 = ~n_42903 & ~n_42904;
assign n_42906 =  x_3635 & ~n_42905;
assign n_42907 = ~x_3635 &  n_42905;
assign n_42908 = ~n_42906 & ~n_42907;
assign n_42909 =  n_25638 & ~n_14891;
assign n_42910 =  x_3634 & ~n_25638;
assign n_42911 = ~n_42909 & ~n_42910;
assign n_42912 =  x_3634 & ~n_42911;
assign n_42913 = ~x_3634 &  n_42911;
assign n_42914 = ~n_42912 & ~n_42913;
assign n_42915 =  n_25638 & ~n_14909;
assign n_42916 =  x_3633 & ~n_25638;
assign n_42917 = ~n_42915 & ~n_42916;
assign n_42918 =  x_3633 & ~n_42917;
assign n_42919 = ~x_3633 &  n_42917;
assign n_42920 = ~n_42918 & ~n_42919;
assign n_42921 =  n_25638 & ~n_14927;
assign n_42922 =  x_3632 & ~n_25638;
assign n_42923 = ~n_42921 & ~n_42922;
assign n_42924 =  x_3632 & ~n_42923;
assign n_42925 = ~x_3632 &  n_42923;
assign n_42926 = ~n_42924 & ~n_42925;
assign n_42927 =  n_25638 & ~n_14945;
assign n_42928 =  x_3631 & ~n_25638;
assign n_42929 = ~n_42927 & ~n_42928;
assign n_42930 =  x_3631 & ~n_42929;
assign n_42931 = ~x_3631 &  n_42929;
assign n_42932 = ~n_42930 & ~n_42931;
assign n_42933 =  n_25638 & ~n_14963;
assign n_42934 =  x_3630 & ~n_25638;
assign n_42935 = ~n_42933 & ~n_42934;
assign n_42936 =  x_3630 & ~n_42935;
assign n_42937 = ~x_3630 &  n_42935;
assign n_42938 = ~n_42936 & ~n_42937;
assign n_42939 =  n_25638 & ~n_14981;
assign n_42940 =  x_3629 & ~n_25638;
assign n_42941 = ~n_42939 & ~n_42940;
assign n_42942 =  x_3629 & ~n_42941;
assign n_42943 = ~x_3629 &  n_42941;
assign n_42944 = ~n_42942 & ~n_42943;
assign n_42945 =  n_25638 & ~n_14999;
assign n_42946 =  x_3628 & ~n_25638;
assign n_42947 = ~n_42945 & ~n_42946;
assign n_42948 =  x_3628 & ~n_42947;
assign n_42949 = ~x_3628 &  n_42947;
assign n_42950 = ~n_42948 & ~n_42949;
assign n_42951 =  n_25638 & ~n_15017;
assign n_42952 =  x_3627 & ~n_25638;
assign n_42953 = ~n_42951 & ~n_42952;
assign n_42954 =  x_3627 & ~n_42953;
assign n_42955 = ~x_3627 &  n_42953;
assign n_42956 = ~n_42954 & ~n_42955;
assign n_42957 =  n_25638 & ~n_15035;
assign n_42958 =  x_3626 & ~n_25638;
assign n_42959 = ~n_42957 & ~n_42958;
assign n_42960 =  x_3626 & ~n_42959;
assign n_42961 = ~x_3626 &  n_42959;
assign n_42962 = ~n_42960 & ~n_42961;
assign n_42963 =  n_25638 & ~n_15053;
assign n_42964 =  x_3625 & ~n_25638;
assign n_42965 = ~n_42963 & ~n_42964;
assign n_42966 =  x_3625 & ~n_42965;
assign n_42967 = ~x_3625 &  n_42965;
assign n_42968 = ~n_42966 & ~n_42967;
assign n_42969 =  n_25638 & ~n_15071;
assign n_42970 =  x_3624 & ~n_25638;
assign n_42971 = ~n_42969 & ~n_42970;
assign n_42972 =  x_3624 & ~n_42971;
assign n_42973 = ~x_3624 &  n_42971;
assign n_42974 = ~n_42972 & ~n_42973;
assign n_42975 =  n_25638 & ~n_15089;
assign n_42976 =  x_3623 & ~n_25638;
assign n_42977 = ~n_42975 & ~n_42976;
assign n_42978 =  x_3623 & ~n_42977;
assign n_42979 = ~x_3623 &  n_42977;
assign n_42980 = ~n_42978 & ~n_42979;
assign n_42981 =  n_25638 & ~n_15107;
assign n_42982 =  x_3622 & ~n_25638;
assign n_42983 = ~n_42981 & ~n_42982;
assign n_42984 =  x_3622 & ~n_42983;
assign n_42985 = ~x_3622 &  n_42983;
assign n_42986 = ~n_42984 & ~n_42985;
assign n_42987 =  n_25638 & ~n_15125;
assign n_42988 =  x_3621 & ~n_25638;
assign n_42989 = ~n_42987 & ~n_42988;
assign n_42990 =  x_3621 & ~n_42989;
assign n_42991 = ~x_3621 &  n_42989;
assign n_42992 = ~n_42990 & ~n_42991;
assign n_42993 =  n_25638 & ~n_15143;
assign n_42994 =  x_3620 & ~n_25638;
assign n_42995 = ~n_42993 & ~n_42994;
assign n_42996 =  x_3620 & ~n_42995;
assign n_42997 = ~x_3620 &  n_42995;
assign n_42998 = ~n_42996 & ~n_42997;
assign n_42999 =  n_25638 & ~n_15161;
assign n_43000 =  x_3619 & ~n_25638;
assign n_43001 = ~n_42999 & ~n_43000;
assign n_43002 =  x_3619 & ~n_43001;
assign n_43003 = ~x_3619 &  n_43001;
assign n_43004 = ~n_43002 & ~n_43003;
assign n_43005 =  n_25638 & ~n_15179;
assign n_43006 =  x_3618 & ~n_25638;
assign n_43007 = ~n_43005 & ~n_43006;
assign n_43008 =  x_3618 & ~n_43007;
assign n_43009 = ~x_3618 &  n_43007;
assign n_43010 = ~n_43008 & ~n_43009;
assign n_43011 =  n_25638 & ~n_15197;
assign n_43012 =  x_3617 & ~n_25638;
assign n_43013 = ~n_43011 & ~n_43012;
assign n_43014 =  x_3617 & ~n_43013;
assign n_43015 = ~x_3617 &  n_43013;
assign n_43016 = ~n_43014 & ~n_43015;
assign n_43017 =  n_25638 & ~n_15215;
assign n_43018 =  x_3616 & ~n_25638;
assign n_43019 = ~n_43017 & ~n_43018;
assign n_43020 =  x_3616 & ~n_43019;
assign n_43021 = ~x_3616 &  n_43019;
assign n_43022 = ~n_43020 & ~n_43021;
assign n_43023 =  n_25638 & ~n_15233;
assign n_43024 =  x_3615 & ~n_25638;
assign n_43025 = ~n_43023 & ~n_43024;
assign n_43026 =  x_3615 & ~n_43025;
assign n_43027 = ~x_3615 &  n_43025;
assign n_43028 = ~n_43026 & ~n_43027;
assign n_43029 =  n_25638 & ~n_15251;
assign n_43030 =  x_3614 & ~n_25638;
assign n_43031 = ~n_43029 & ~n_43030;
assign n_43032 =  x_3614 & ~n_43031;
assign n_43033 = ~x_3614 &  n_43031;
assign n_43034 = ~n_43032 & ~n_43033;
assign n_43035 =  n_25638 & ~n_15269;
assign n_43036 =  x_3613 & ~n_25638;
assign n_43037 = ~n_43035 & ~n_43036;
assign n_43038 =  x_3613 & ~n_43037;
assign n_43039 = ~x_3613 &  n_43037;
assign n_43040 = ~n_43038 & ~n_43039;
assign n_43041 =  n_25638 & ~n_15287;
assign n_43042 =  x_3612 & ~n_25638;
assign n_43043 = ~n_43041 & ~n_43042;
assign n_43044 =  x_3612 & ~n_43043;
assign n_43045 = ~x_3612 &  n_43043;
assign n_43046 = ~n_43044 & ~n_43045;
assign n_43047 =  n_25638 & ~n_15305;
assign n_43048 =  x_3611 & ~n_25638;
assign n_43049 = ~n_43047 & ~n_43048;
assign n_43050 =  x_3611 & ~n_43049;
assign n_43051 = ~x_3611 &  n_43049;
assign n_43052 = ~n_43050 & ~n_43051;
assign n_43053 =  n_25638 & ~n_15323;
assign n_43054 =  x_3610 & ~n_25638;
assign n_43055 = ~n_43053 & ~n_43054;
assign n_43056 =  x_3610 & ~n_43055;
assign n_43057 = ~x_3610 &  n_43055;
assign n_43058 = ~n_43056 & ~n_43057;
assign n_43059 =  n_25638 & ~n_15341;
assign n_43060 =  x_3609 & ~n_25638;
assign n_43061 = ~n_43059 & ~n_43060;
assign n_43062 =  x_3609 & ~n_43061;
assign n_43063 = ~x_3609 &  n_43061;
assign n_43064 = ~n_43062 & ~n_43063;
assign n_43065 =  n_25638 & ~n_15359;
assign n_43066 =  x_3608 & ~n_25638;
assign n_43067 = ~n_43065 & ~n_43066;
assign n_43068 =  x_3608 & ~n_43067;
assign n_43069 = ~x_3608 &  n_43067;
assign n_43070 = ~n_43068 & ~n_43069;
assign n_43071 = ~n_23851 & ~n_25653;
assign n_43072 =  n_28564 &  n_43071;
assign n_43073 =  x_3607 &  n_43072;
assign n_43074 =  x_1002 &  n_25653;
assign n_43075 =  x_3351 &  n_23851;
assign n_43076 =  x_4264 &  n_27122;
assign n_43077 = ~n_43075 & ~n_43076;
assign n_43078 = ~n_43074 &  n_43077;
assign n_43079 = ~n_43073 &  n_43078;
assign n_43080 =  x_3607 & ~n_43079;
assign n_43081 = ~x_3607 &  n_43079;
assign n_43082 = ~n_43080 & ~n_43081;
assign n_43083 =  x_3606 &  n_43072;
assign n_43084 =  x_1001 &  n_25653;
assign n_43085 =  x_3350 &  n_23851;
assign n_43086 =  x_4263 &  n_27122;
assign n_43087 = ~n_43085 & ~n_43086;
assign n_43088 = ~n_43084 &  n_43087;
assign n_43089 = ~n_43083 &  n_43088;
assign n_43090 =  x_3606 & ~n_43089;
assign n_43091 = ~x_3606 &  n_43089;
assign n_43092 = ~n_43090 & ~n_43091;
assign n_43093 =  x_3605 &  n_43072;
assign n_43094 =  x_1000 &  n_25653;
assign n_43095 =  x_3349 &  n_23851;
assign n_43096 =  x_4262 &  n_27122;
assign n_43097 = ~n_43095 & ~n_43096;
assign n_43098 = ~n_43094 &  n_43097;
assign n_43099 = ~n_43093 &  n_43098;
assign n_43100 =  x_3605 & ~n_43099;
assign n_43101 = ~x_3605 &  n_43099;
assign n_43102 = ~n_43100 & ~n_43101;
assign n_43103 =  x_3604 &  n_43072;
assign n_43104 =  x_999 &  n_25653;
assign n_43105 =  x_3348 &  n_23851;
assign n_43106 =  x_4261 &  n_27122;
assign n_43107 = ~n_43105 & ~n_43106;
assign n_43108 = ~n_43104 &  n_43107;
assign n_43109 = ~n_43103 &  n_43108;
assign n_43110 =  x_3604 & ~n_43109;
assign n_43111 = ~x_3604 &  n_43109;
assign n_43112 = ~n_43110 & ~n_43111;
assign n_43113 =  x_3603 &  n_43072;
assign n_43114 =  x_998 &  n_25653;
assign n_43115 =  x_3347 &  n_23851;
assign n_43116 =  x_4260 &  n_27122;
assign n_43117 = ~n_43115 & ~n_43116;
assign n_43118 = ~n_43114 &  n_43117;
assign n_43119 = ~n_43113 &  n_43118;
assign n_43120 =  x_3603 & ~n_43119;
assign n_43121 = ~x_3603 &  n_43119;
assign n_43122 = ~n_43120 & ~n_43121;
assign n_43123 =  x_3602 &  n_43072;
assign n_43124 =  x_997 &  n_25653;
assign n_43125 =  x_3346 &  n_23851;
assign n_43126 =  x_4259 &  n_27122;
assign n_43127 = ~n_43125 & ~n_43126;
assign n_43128 = ~n_43124 &  n_43127;
assign n_43129 = ~n_43123 &  n_43128;
assign n_43130 =  x_3602 & ~n_43129;
assign n_43131 = ~x_3602 &  n_43129;
assign n_43132 = ~n_43130 & ~n_43131;
assign n_43133 =  x_3601 &  n_43072;
assign n_43134 =  x_996 &  n_25653;
assign n_43135 =  x_3345 &  n_23851;
assign n_43136 =  x_4258 &  n_27122;
assign n_43137 = ~n_43135 & ~n_43136;
assign n_43138 = ~n_43134 &  n_43137;
assign n_43139 = ~n_43133 &  n_43138;
assign n_43140 =  x_3601 & ~n_43139;
assign n_43141 = ~x_3601 &  n_43139;
assign n_43142 = ~n_43140 & ~n_43141;
assign n_43143 =  x_3600 &  n_43072;
assign n_43144 =  x_995 &  n_25653;
assign n_43145 =  x_3344 &  n_23851;
assign n_43146 =  x_4257 &  n_27122;
assign n_43147 = ~n_43145 & ~n_43146;
assign n_43148 = ~n_43144 &  n_43147;
assign n_43149 = ~n_43143 &  n_43148;
assign n_43150 =  x_3600 & ~n_43149;
assign n_43151 = ~x_3600 &  n_43149;
assign n_43152 = ~n_43150 & ~n_43151;
assign n_43153 =  x_3599 &  n_43072;
assign n_43154 =  x_994 &  n_25653;
assign n_43155 =  x_3343 &  n_23851;
assign n_43156 =  x_4256 &  n_27122;
assign n_43157 = ~n_43155 & ~n_43156;
assign n_43158 = ~n_43154 &  n_43157;
assign n_43159 = ~n_43153 &  n_43158;
assign n_43160 =  x_3599 & ~n_43159;
assign n_43161 = ~x_3599 &  n_43159;
assign n_43162 = ~n_43160 & ~n_43161;
assign n_43163 =  x_3598 &  n_43072;
assign n_43164 =  x_993 &  n_25653;
assign n_43165 =  x_3342 &  n_23851;
assign n_43166 =  x_4255 &  n_27122;
assign n_43167 = ~n_43165 & ~n_43166;
assign n_43168 = ~n_43164 &  n_43167;
assign n_43169 = ~n_43163 &  n_43168;
assign n_43170 =  x_3598 & ~n_43169;
assign n_43171 = ~x_3598 &  n_43169;
assign n_43172 = ~n_43170 & ~n_43171;
assign n_43173 =  x_3597 &  n_43072;
assign n_43174 =  x_992 &  n_25653;
assign n_43175 =  x_3341 &  n_23851;
assign n_43176 =  x_4254 &  n_27122;
assign n_43177 = ~n_43175 & ~n_43176;
assign n_43178 = ~n_43174 &  n_43177;
assign n_43179 = ~n_43173 &  n_43178;
assign n_43180 =  x_3597 & ~n_43179;
assign n_43181 = ~x_3597 &  n_43179;
assign n_43182 = ~n_43180 & ~n_43181;
assign n_43183 =  x_3596 &  n_43072;
assign n_43184 =  x_991 &  n_25653;
assign n_43185 =  x_3340 &  n_23851;
assign n_43186 =  x_4253 &  n_27122;
assign n_43187 = ~n_43185 & ~n_43186;
assign n_43188 = ~n_43184 &  n_43187;
assign n_43189 = ~n_43183 &  n_43188;
assign n_43190 =  x_3596 & ~n_43189;
assign n_43191 = ~x_3596 &  n_43189;
assign n_43192 = ~n_43190 & ~n_43191;
assign n_43193 =  x_3595 &  n_43072;
assign n_43194 =  x_990 &  n_25653;
assign n_43195 =  x_3339 &  n_23851;
assign n_43196 =  x_4252 &  n_27122;
assign n_43197 = ~n_43195 & ~n_43196;
assign n_43198 = ~n_43194 &  n_43197;
assign n_43199 = ~n_43193 &  n_43198;
assign n_43200 =  x_3595 & ~n_43199;
assign n_43201 = ~x_3595 &  n_43199;
assign n_43202 = ~n_43200 & ~n_43201;
assign n_43203 =  x_3594 &  n_43072;
assign n_43204 =  x_989 &  n_25653;
assign n_43205 =  x_3338 &  n_23851;
assign n_43206 =  x_4251 &  n_27122;
assign n_43207 = ~n_43205 & ~n_43206;
assign n_43208 = ~n_43204 &  n_43207;
assign n_43209 = ~n_43203 &  n_43208;
assign n_43210 =  x_3594 & ~n_43209;
assign n_43211 = ~x_3594 &  n_43209;
assign n_43212 = ~n_43210 & ~n_43211;
assign n_43213 =  x_3593 &  n_43072;
assign n_43214 =  x_988 &  n_25653;
assign n_43215 =  x_3337 &  n_23851;
assign n_43216 =  x_4250 &  n_27122;
assign n_43217 = ~n_43215 & ~n_43216;
assign n_43218 = ~n_43214 &  n_43217;
assign n_43219 = ~n_43213 &  n_43218;
assign n_43220 =  x_3593 & ~n_43219;
assign n_43221 = ~x_3593 &  n_43219;
assign n_43222 = ~n_43220 & ~n_43221;
assign n_43223 =  x_3592 &  n_43072;
assign n_43224 =  x_987 &  n_25653;
assign n_43225 =  x_3336 &  n_23851;
assign n_43226 =  x_4249 &  n_27122;
assign n_43227 = ~n_43225 & ~n_43226;
assign n_43228 = ~n_43224 &  n_43227;
assign n_43229 = ~n_43223 &  n_43228;
assign n_43230 =  x_3592 & ~n_43229;
assign n_43231 = ~x_3592 &  n_43229;
assign n_43232 = ~n_43230 & ~n_43231;
assign n_43233 =  x_3591 &  n_43072;
assign n_43234 =  x_986 &  n_25653;
assign n_43235 =  x_3335 &  n_23851;
assign n_43236 =  x_4248 &  n_27122;
assign n_43237 = ~n_43235 & ~n_43236;
assign n_43238 = ~n_43234 &  n_43237;
assign n_43239 = ~n_43233 &  n_43238;
assign n_43240 =  x_3591 & ~n_43239;
assign n_43241 = ~x_3591 &  n_43239;
assign n_43242 = ~n_43240 & ~n_43241;
assign n_43243 =  x_3590 &  n_43072;
assign n_43244 =  x_985 &  n_25653;
assign n_43245 =  x_3334 &  n_23851;
assign n_43246 =  x_4247 &  n_27122;
assign n_43247 = ~n_43245 & ~n_43246;
assign n_43248 = ~n_43244 &  n_43247;
assign n_43249 = ~n_43243 &  n_43248;
assign n_43250 =  x_3590 & ~n_43249;
assign n_43251 = ~x_3590 &  n_43249;
assign n_43252 = ~n_43250 & ~n_43251;
assign n_43253 =  x_3589 &  n_43072;
assign n_43254 =  x_984 &  n_25653;
assign n_43255 =  x_3333 &  n_23851;
assign n_43256 =  x_4246 &  n_27122;
assign n_43257 = ~n_43255 & ~n_43256;
assign n_43258 = ~n_43254 &  n_43257;
assign n_43259 = ~n_43253 &  n_43258;
assign n_43260 =  x_3589 & ~n_43259;
assign n_43261 = ~x_3589 &  n_43259;
assign n_43262 = ~n_43260 & ~n_43261;
assign n_43263 =  x_3588 &  n_43072;
assign n_43264 =  x_983 &  n_25653;
assign n_43265 =  x_3332 &  n_23851;
assign n_43266 =  x_4245 &  n_27122;
assign n_43267 = ~n_43265 & ~n_43266;
assign n_43268 = ~n_43264 &  n_43267;
assign n_43269 = ~n_43263 &  n_43268;
assign n_43270 =  x_3588 & ~n_43269;
assign n_43271 = ~x_3588 &  n_43269;
assign n_43272 = ~n_43270 & ~n_43271;
assign n_43273 =  x_3587 &  n_43072;
assign n_43274 =  x_982 &  n_25653;
assign n_43275 =  x_3331 &  n_23851;
assign n_43276 =  x_4244 &  n_27122;
assign n_43277 = ~n_43275 & ~n_43276;
assign n_43278 = ~n_43274 &  n_43277;
assign n_43279 = ~n_43273 &  n_43278;
assign n_43280 =  x_3587 & ~n_43279;
assign n_43281 = ~x_3587 &  n_43279;
assign n_43282 = ~n_43280 & ~n_43281;
assign n_43283 =  x_3586 &  n_43072;
assign n_43284 =  x_981 &  n_25653;
assign n_43285 =  x_3330 &  n_23851;
assign n_43286 =  x_4243 &  n_27122;
assign n_43287 = ~n_43285 & ~n_43286;
assign n_43288 = ~n_43284 &  n_43287;
assign n_43289 = ~n_43283 &  n_43288;
assign n_43290 =  x_3586 & ~n_43289;
assign n_43291 = ~x_3586 &  n_43289;
assign n_43292 = ~n_43290 & ~n_43291;
assign n_43293 =  x_3585 &  n_43072;
assign n_43294 =  x_980 &  n_25653;
assign n_43295 =  x_3329 &  n_23851;
assign n_43296 =  x_4242 &  n_27122;
assign n_43297 = ~n_43295 & ~n_43296;
assign n_43298 = ~n_43294 &  n_43297;
assign n_43299 = ~n_43293 &  n_43298;
assign n_43300 =  x_3585 & ~n_43299;
assign n_43301 = ~x_3585 &  n_43299;
assign n_43302 = ~n_43300 & ~n_43301;
assign n_43303 =  x_3584 &  n_43072;
assign n_43304 =  x_979 &  n_25653;
assign n_43305 =  x_3328 &  n_23851;
assign n_43306 =  x_4241 &  n_27122;
assign n_43307 = ~n_43305 & ~n_43306;
assign n_43308 = ~n_43304 &  n_43307;
assign n_43309 = ~n_43303 &  n_43308;
assign n_43310 =  x_3584 & ~n_43309;
assign n_43311 = ~x_3584 &  n_43309;
assign n_43312 = ~n_43310 & ~n_43311;
assign n_43313 =  x_3583 &  n_43072;
assign n_43314 =  x_978 &  n_25653;
assign n_43315 =  x_3327 &  n_23851;
assign n_43316 =  x_4240 &  n_27122;
assign n_43317 = ~n_43315 & ~n_43316;
assign n_43318 = ~n_43314 &  n_43317;
assign n_43319 = ~n_43313 &  n_43318;
assign n_43320 =  x_3583 & ~n_43319;
assign n_43321 = ~x_3583 &  n_43319;
assign n_43322 = ~n_43320 & ~n_43321;
assign n_43323 =  x_3582 &  n_43072;
assign n_43324 =  x_977 &  n_25653;
assign n_43325 =  x_3326 &  n_23851;
assign n_43326 =  x_4239 &  n_27122;
assign n_43327 = ~n_43325 & ~n_43326;
assign n_43328 = ~n_43324 &  n_43327;
assign n_43329 = ~n_43323 &  n_43328;
assign n_43330 =  x_3582 & ~n_43329;
assign n_43331 = ~x_3582 &  n_43329;
assign n_43332 = ~n_43330 & ~n_43331;
assign n_43333 =  x_3581 &  n_43072;
assign n_43334 =  x_976 &  n_25653;
assign n_43335 =  x_3325 &  n_23851;
assign n_43336 =  x_4238 &  n_27122;
assign n_43337 = ~n_43335 & ~n_43336;
assign n_43338 = ~n_43334 &  n_43337;
assign n_43339 = ~n_43333 &  n_43338;
assign n_43340 =  x_3581 & ~n_43339;
assign n_43341 = ~x_3581 &  n_43339;
assign n_43342 = ~n_43340 & ~n_43341;
assign n_43343 =  x_3580 &  n_43072;
assign n_43344 =  x_975 &  n_25653;
assign n_43345 =  x_3324 &  n_23851;
assign n_43346 =  x_4237 &  n_27122;
assign n_43347 = ~n_43345 & ~n_43346;
assign n_43348 = ~n_43344 &  n_43347;
assign n_43349 = ~n_43343 &  n_43348;
assign n_43350 =  x_3580 & ~n_43349;
assign n_43351 = ~x_3580 &  n_43349;
assign n_43352 = ~n_43350 & ~n_43351;
assign n_43353 =  x_3579 &  n_43072;
assign n_43354 =  x_974 &  n_25653;
assign n_43355 =  x_3323 &  n_23851;
assign n_43356 =  x_4236 &  n_27122;
assign n_43357 = ~n_43355 & ~n_43356;
assign n_43358 = ~n_43354 &  n_43357;
assign n_43359 = ~n_43353 &  n_43358;
assign n_43360 =  x_3579 & ~n_43359;
assign n_43361 = ~x_3579 &  n_43359;
assign n_43362 = ~n_43360 & ~n_43361;
assign n_43363 =  x_3578 &  n_43072;
assign n_43364 =  x_973 &  n_25653;
assign n_43365 =  x_3322 &  n_23851;
assign n_43366 =  x_4235 &  n_27122;
assign n_43367 = ~n_43365 & ~n_43366;
assign n_43368 = ~n_43364 &  n_43367;
assign n_43369 = ~n_43363 &  n_43368;
assign n_43370 =  x_3578 & ~n_43369;
assign n_43371 = ~x_3578 &  n_43369;
assign n_43372 = ~n_43370 & ~n_43371;
assign n_43373 =  x_3577 &  n_43072;
assign n_43374 =  x_972 &  n_25653;
assign n_43375 =  x_3321 &  n_23851;
assign n_43376 =  x_4234 &  n_27122;
assign n_43377 = ~n_43375 & ~n_43376;
assign n_43378 = ~n_43374 &  n_43377;
assign n_43379 = ~n_43373 &  n_43378;
assign n_43380 =  x_3577 & ~n_43379;
assign n_43381 = ~x_3577 &  n_43379;
assign n_43382 = ~n_43380 & ~n_43381;
assign n_43383 =  x_3576 &  n_43072;
assign n_43384 =  x_971 &  n_25653;
assign n_43385 =  x_3320 &  n_23851;
assign n_43386 =  x_4233 &  n_27122;
assign n_43387 = ~n_43385 & ~n_43386;
assign n_43388 = ~n_43384 &  n_43387;
assign n_43389 = ~n_43383 &  n_43388;
assign n_43390 =  x_3576 & ~n_43389;
assign n_43391 = ~x_3576 &  n_43389;
assign n_43392 = ~n_43390 & ~n_43391;
assign n_43393 = ~n_26889 & ~n_25660;
assign n_43394 =  n_29021 &  n_43393;
assign n_43395 =  x_3575 &  n_43394;
assign n_43396 =  x_4232 &  n_25660;
assign n_43397 =  x_2490 &  n_26889;
assign n_43398 =  x_970 &  n_26426;
assign n_43399 = ~n_43397 & ~n_43398;
assign n_43400 = ~n_43396 &  n_43399;
assign n_43401 = ~n_43395 &  n_43400;
assign n_43402 =  x_3575 & ~n_43401;
assign n_43403 = ~x_3575 &  n_43401;
assign n_43404 = ~n_43402 & ~n_43403;
assign n_43405 =  x_3574 &  n_43394;
assign n_43406 =  x_4231 &  n_25660;
assign n_43407 =  x_2489 &  n_26889;
assign n_43408 =  x_969 &  n_26426;
assign n_43409 = ~n_43407 & ~n_43408;
assign n_43410 = ~n_43406 &  n_43409;
assign n_43411 = ~n_43405 &  n_43410;
assign n_43412 =  x_3574 & ~n_43411;
assign n_43413 = ~x_3574 &  n_43411;
assign n_43414 = ~n_43412 & ~n_43413;
assign n_43415 =  x_3573 &  n_43394;
assign n_43416 =  x_4230 &  n_25660;
assign n_43417 =  x_2488 &  n_26889;
assign n_43418 =  x_968 &  n_26426;
assign n_43419 = ~n_43417 & ~n_43418;
assign n_43420 = ~n_43416 &  n_43419;
assign n_43421 = ~n_43415 &  n_43420;
assign n_43422 =  x_3573 & ~n_43421;
assign n_43423 = ~x_3573 &  n_43421;
assign n_43424 = ~n_43422 & ~n_43423;
assign n_43425 =  x_3572 &  n_43394;
assign n_43426 =  x_4229 &  n_25660;
assign n_43427 =  x_2487 &  n_26889;
assign n_43428 =  x_967 &  n_26426;
assign n_43429 = ~n_43427 & ~n_43428;
assign n_43430 = ~n_43426 &  n_43429;
assign n_43431 = ~n_43425 &  n_43430;
assign n_43432 =  x_3572 & ~n_43431;
assign n_43433 = ~x_3572 &  n_43431;
assign n_43434 = ~n_43432 & ~n_43433;
assign n_43435 =  x_3571 &  n_43394;
assign n_43436 =  x_4228 &  n_25660;
assign n_43437 =  x_2486 &  n_26889;
assign n_43438 =  x_966 &  n_26426;
assign n_43439 = ~n_43437 & ~n_43438;
assign n_43440 = ~n_43436 &  n_43439;
assign n_43441 = ~n_43435 &  n_43440;
assign n_43442 =  x_3571 & ~n_43441;
assign n_43443 = ~x_3571 &  n_43441;
assign n_43444 = ~n_43442 & ~n_43443;
assign n_43445 =  x_3570 &  n_43394;
assign n_43446 =  x_4227 &  n_25660;
assign n_43447 =  x_2485 &  n_26889;
assign n_43448 =  x_965 &  n_26426;
assign n_43449 = ~n_43447 & ~n_43448;
assign n_43450 = ~n_43446 &  n_43449;
assign n_43451 = ~n_43445 &  n_43450;
assign n_43452 =  x_3570 & ~n_43451;
assign n_43453 = ~x_3570 &  n_43451;
assign n_43454 = ~n_43452 & ~n_43453;
assign n_43455 =  x_3569 &  n_43394;
assign n_43456 =  x_4226 &  n_25660;
assign n_43457 =  x_2484 &  n_26889;
assign n_43458 =  x_964 &  n_26426;
assign n_43459 = ~n_43457 & ~n_43458;
assign n_43460 = ~n_43456 &  n_43459;
assign n_43461 = ~n_43455 &  n_43460;
assign n_43462 =  x_3569 & ~n_43461;
assign n_43463 = ~x_3569 &  n_43461;
assign n_43464 = ~n_43462 & ~n_43463;
assign n_43465 =  x_3568 &  n_43394;
assign n_43466 =  x_4225 &  n_25660;
assign n_43467 =  x_2483 &  n_26889;
assign n_43468 =  x_963 &  n_26426;
assign n_43469 = ~n_43467 & ~n_43468;
assign n_43470 = ~n_43466 &  n_43469;
assign n_43471 = ~n_43465 &  n_43470;
assign n_43472 =  x_3568 & ~n_43471;
assign n_43473 = ~x_3568 &  n_43471;
assign n_43474 = ~n_43472 & ~n_43473;
assign n_43475 =  x_3567 &  n_43394;
assign n_43476 =  x_4224 &  n_25660;
assign n_43477 =  x_2482 &  n_26889;
assign n_43478 =  x_962 &  n_26426;
assign n_43479 = ~n_43477 & ~n_43478;
assign n_43480 = ~n_43476 &  n_43479;
assign n_43481 = ~n_43475 &  n_43480;
assign n_43482 =  x_3567 & ~n_43481;
assign n_43483 = ~x_3567 &  n_43481;
assign n_43484 = ~n_43482 & ~n_43483;
assign n_43485 =  x_3566 &  n_43394;
assign n_43486 =  x_4223 &  n_25660;
assign n_43487 =  x_2481 &  n_26889;
assign n_43488 =  x_961 &  n_26426;
assign n_43489 = ~n_43487 & ~n_43488;
assign n_43490 = ~n_43486 &  n_43489;
assign n_43491 = ~n_43485 &  n_43490;
assign n_43492 =  x_3566 & ~n_43491;
assign n_43493 = ~x_3566 &  n_43491;
assign n_43494 = ~n_43492 & ~n_43493;
assign n_43495 =  x_3565 &  n_43394;
assign n_43496 =  x_4222 &  n_25660;
assign n_43497 =  x_2480 &  n_26889;
assign n_43498 =  x_960 &  n_26426;
assign n_43499 = ~n_43497 & ~n_43498;
assign n_43500 = ~n_43496 &  n_43499;
assign n_43501 = ~n_43495 &  n_43500;
assign n_43502 =  x_3565 & ~n_43501;
assign n_43503 = ~x_3565 &  n_43501;
assign n_43504 = ~n_43502 & ~n_43503;
assign n_43505 =  x_3564 &  n_43394;
assign n_43506 =  x_4221 &  n_25660;
assign n_43507 =  x_2479 &  n_26889;
assign n_43508 =  x_959 &  n_26426;
assign n_43509 = ~n_43507 & ~n_43508;
assign n_43510 = ~n_43506 &  n_43509;
assign n_43511 = ~n_43505 &  n_43510;
assign n_43512 =  x_3564 & ~n_43511;
assign n_43513 = ~x_3564 &  n_43511;
assign n_43514 = ~n_43512 & ~n_43513;
assign n_43515 =  x_3563 &  n_43394;
assign n_43516 =  x_4220 &  n_25660;
assign n_43517 =  x_2478 &  n_26889;
assign n_43518 =  x_958 &  n_26426;
assign n_43519 = ~n_43517 & ~n_43518;
assign n_43520 = ~n_43516 &  n_43519;
assign n_43521 = ~n_43515 &  n_43520;
assign n_43522 =  x_3563 & ~n_43521;
assign n_43523 = ~x_3563 &  n_43521;
assign n_43524 = ~n_43522 & ~n_43523;
assign n_43525 =  x_3562 &  n_43394;
assign n_43526 =  x_4219 &  n_25660;
assign n_43527 =  x_2477 &  n_26889;
assign n_43528 =  x_957 &  n_26426;
assign n_43529 = ~n_43527 & ~n_43528;
assign n_43530 = ~n_43526 &  n_43529;
assign n_43531 = ~n_43525 &  n_43530;
assign n_43532 =  x_3562 & ~n_43531;
assign n_43533 = ~x_3562 &  n_43531;
assign n_43534 = ~n_43532 & ~n_43533;
assign n_43535 =  x_3561 &  n_43394;
assign n_43536 =  x_4218 &  n_25660;
assign n_43537 =  x_2476 &  n_26889;
assign n_43538 =  x_956 &  n_26426;
assign n_43539 = ~n_43537 & ~n_43538;
assign n_43540 = ~n_43536 &  n_43539;
assign n_43541 = ~n_43535 &  n_43540;
assign n_43542 =  x_3561 & ~n_43541;
assign n_43543 = ~x_3561 &  n_43541;
assign n_43544 = ~n_43542 & ~n_43543;
assign n_43545 =  x_3560 &  n_43394;
assign n_43546 =  x_4217 &  n_25660;
assign n_43547 =  x_2475 &  n_26889;
assign n_43548 =  x_955 &  n_26426;
assign n_43549 = ~n_43547 & ~n_43548;
assign n_43550 = ~n_43546 &  n_43549;
assign n_43551 = ~n_43545 &  n_43550;
assign n_43552 =  x_3560 & ~n_43551;
assign n_43553 = ~x_3560 &  n_43551;
assign n_43554 = ~n_43552 & ~n_43553;
assign n_43555 =  x_3559 &  n_43394;
assign n_43556 =  x_4216 &  n_25660;
assign n_43557 =  x_2474 &  n_26889;
assign n_43558 =  x_954 &  n_26426;
assign n_43559 = ~n_43557 & ~n_43558;
assign n_43560 = ~n_43556 &  n_43559;
assign n_43561 = ~n_43555 &  n_43560;
assign n_43562 =  x_3559 & ~n_43561;
assign n_43563 = ~x_3559 &  n_43561;
assign n_43564 = ~n_43562 & ~n_43563;
assign n_43565 =  x_3558 &  n_43394;
assign n_43566 =  x_4215 &  n_25660;
assign n_43567 =  x_2473 &  n_26889;
assign n_43568 =  x_953 &  n_26426;
assign n_43569 = ~n_43567 & ~n_43568;
assign n_43570 = ~n_43566 &  n_43569;
assign n_43571 = ~n_43565 &  n_43570;
assign n_43572 =  x_3558 & ~n_43571;
assign n_43573 = ~x_3558 &  n_43571;
assign n_43574 = ~n_43572 & ~n_43573;
assign n_43575 =  x_3557 &  n_43394;
assign n_43576 =  x_4214 &  n_25660;
assign n_43577 =  x_2472 &  n_26889;
assign n_43578 =  x_952 &  n_26426;
assign n_43579 = ~n_43577 & ~n_43578;
assign n_43580 = ~n_43576 &  n_43579;
assign n_43581 = ~n_43575 &  n_43580;
assign n_43582 =  x_3557 & ~n_43581;
assign n_43583 = ~x_3557 &  n_43581;
assign n_43584 = ~n_43582 & ~n_43583;
assign n_43585 =  x_3556 &  n_43394;
assign n_43586 =  x_4213 &  n_25660;
assign n_43587 =  x_2471 &  n_26889;
assign n_43588 =  x_951 &  n_26426;
assign n_43589 = ~n_43587 & ~n_43588;
assign n_43590 = ~n_43586 &  n_43589;
assign n_43591 = ~n_43585 &  n_43590;
assign n_43592 =  x_3556 & ~n_43591;
assign n_43593 = ~x_3556 &  n_43591;
assign n_43594 = ~n_43592 & ~n_43593;
assign n_43595 =  x_3555 &  n_43394;
assign n_43596 =  x_4212 &  n_25660;
assign n_43597 =  x_2470 &  n_26889;
assign n_43598 =  x_950 &  n_26426;
assign n_43599 = ~n_43597 & ~n_43598;
assign n_43600 = ~n_43596 &  n_43599;
assign n_43601 = ~n_43595 &  n_43600;
assign n_43602 =  x_3555 & ~n_43601;
assign n_43603 = ~x_3555 &  n_43601;
assign n_43604 = ~n_43602 & ~n_43603;
assign n_43605 =  x_3554 &  n_43394;
assign n_43606 =  x_4211 &  n_25660;
assign n_43607 =  x_2469 &  n_26889;
assign n_43608 =  x_949 &  n_26426;
assign n_43609 = ~n_43607 & ~n_43608;
assign n_43610 = ~n_43606 &  n_43609;
assign n_43611 = ~n_43605 &  n_43610;
assign n_43612 =  x_3554 & ~n_43611;
assign n_43613 = ~x_3554 &  n_43611;
assign n_43614 = ~n_43612 & ~n_43613;
assign n_43615 =  x_3553 &  n_43394;
assign n_43616 =  x_4210 &  n_25660;
assign n_43617 =  x_2468 &  n_26889;
assign n_43618 =  x_948 &  n_26426;
assign n_43619 = ~n_43617 & ~n_43618;
assign n_43620 = ~n_43616 &  n_43619;
assign n_43621 = ~n_43615 &  n_43620;
assign n_43622 =  x_3553 & ~n_43621;
assign n_43623 = ~x_3553 &  n_43621;
assign n_43624 = ~n_43622 & ~n_43623;
assign n_43625 =  x_3552 &  n_43394;
assign n_43626 =  x_4209 &  n_25660;
assign n_43627 =  x_2467 &  n_26889;
assign n_43628 =  x_947 &  n_26426;
assign n_43629 = ~n_43627 & ~n_43628;
assign n_43630 = ~n_43626 &  n_43629;
assign n_43631 = ~n_43625 &  n_43630;
assign n_43632 =  x_3552 & ~n_43631;
assign n_43633 = ~x_3552 &  n_43631;
assign n_43634 = ~n_43632 & ~n_43633;
assign n_43635 =  x_3551 &  n_43394;
assign n_43636 =  x_4208 &  n_25660;
assign n_43637 =  x_2466 &  n_26889;
assign n_43638 =  x_946 &  n_26426;
assign n_43639 = ~n_43637 & ~n_43638;
assign n_43640 = ~n_43636 &  n_43639;
assign n_43641 = ~n_43635 &  n_43640;
assign n_43642 =  x_3551 & ~n_43641;
assign n_43643 = ~x_3551 &  n_43641;
assign n_43644 = ~n_43642 & ~n_43643;
assign n_43645 =  x_3550 &  n_43394;
assign n_43646 =  x_4207 &  n_25660;
assign n_43647 =  x_2465 &  n_26889;
assign n_43648 =  x_945 &  n_26426;
assign n_43649 = ~n_43647 & ~n_43648;
assign n_43650 = ~n_43646 &  n_43649;
assign n_43651 = ~n_43645 &  n_43650;
assign n_43652 =  x_3550 & ~n_43651;
assign n_43653 = ~x_3550 &  n_43651;
assign n_43654 = ~n_43652 & ~n_43653;
assign n_43655 =  x_3549 &  n_43394;
assign n_43656 =  x_4206 &  n_25660;
assign n_43657 =  x_2464 &  n_26889;
assign n_43658 =  x_944 &  n_26426;
assign n_43659 = ~n_43657 & ~n_43658;
assign n_43660 = ~n_43656 &  n_43659;
assign n_43661 = ~n_43655 &  n_43660;
assign n_43662 =  x_3549 & ~n_43661;
assign n_43663 = ~x_3549 &  n_43661;
assign n_43664 = ~n_43662 & ~n_43663;
assign n_43665 =  x_3548 &  n_43394;
assign n_43666 =  x_4205 &  n_25660;
assign n_43667 =  x_2463 &  n_26889;
assign n_43668 =  x_943 &  n_26426;
assign n_43669 = ~n_43667 & ~n_43668;
assign n_43670 = ~n_43666 &  n_43669;
assign n_43671 = ~n_43665 &  n_43670;
assign n_43672 =  x_3548 & ~n_43671;
assign n_43673 = ~x_3548 &  n_43671;
assign n_43674 = ~n_43672 & ~n_43673;
assign n_43675 =  x_3547 &  n_43394;
assign n_43676 =  x_4204 &  n_25660;
assign n_43677 =  x_2462 &  n_26889;
assign n_43678 =  x_942 &  n_26426;
assign n_43679 = ~n_43677 & ~n_43678;
assign n_43680 = ~n_43676 &  n_43679;
assign n_43681 = ~n_43675 &  n_43680;
assign n_43682 =  x_3547 & ~n_43681;
assign n_43683 = ~x_3547 &  n_43681;
assign n_43684 = ~n_43682 & ~n_43683;
assign n_43685 =  x_3546 &  n_43394;
assign n_43686 =  x_4203 &  n_25660;
assign n_43687 =  x_2461 &  n_26889;
assign n_43688 =  x_941 &  n_26426;
assign n_43689 = ~n_43687 & ~n_43688;
assign n_43690 = ~n_43686 &  n_43689;
assign n_43691 = ~n_43685 &  n_43690;
assign n_43692 =  x_3546 & ~n_43691;
assign n_43693 = ~x_3546 &  n_43691;
assign n_43694 = ~n_43692 & ~n_43693;
assign n_43695 =  x_3545 &  n_43394;
assign n_43696 =  x_4202 &  n_25660;
assign n_43697 =  x_2460 &  n_26889;
assign n_43698 =  x_940 &  n_26426;
assign n_43699 = ~n_43697 & ~n_43698;
assign n_43700 = ~n_43696 &  n_43699;
assign n_43701 = ~n_43695 &  n_43700;
assign n_43702 =  x_3545 & ~n_43701;
assign n_43703 = ~x_3545 &  n_43701;
assign n_43704 = ~n_43702 & ~n_43703;
assign n_43705 =  x_3544 &  n_43394;
assign n_43706 =  x_4201 &  n_25660;
assign n_43707 =  x_2459 &  n_26889;
assign n_43708 =  x_939 &  n_26426;
assign n_43709 = ~n_43707 & ~n_43708;
assign n_43710 = ~n_43706 &  n_43709;
assign n_43711 = ~n_43705 &  n_43710;
assign n_43712 =  x_3544 & ~n_43711;
assign n_43713 = ~x_3544 &  n_43711;
assign n_43714 = ~n_43712 & ~n_43713;
assign n_43715 =  x_3543 & ~n_26240;
assign n_43716 =  i_32 &  n_26240;
assign n_43717 = ~n_43715 & ~n_43716;
assign n_43718 =  x_3543 & ~n_43717;
assign n_43719 = ~x_3543 &  n_43717;
assign n_43720 = ~n_43718 & ~n_43719;
assign n_43721 =  x_3542 & ~n_26240;
assign n_43722 =  i_31 &  n_26240;
assign n_43723 = ~n_43721 & ~n_43722;
assign n_43724 =  x_3542 & ~n_43723;
assign n_43725 = ~x_3542 &  n_43723;
assign n_43726 = ~n_43724 & ~n_43725;
assign n_43727 =  x_3541 & ~n_26240;
assign n_43728 =  i_30 &  n_26240;
assign n_43729 = ~n_43727 & ~n_43728;
assign n_43730 =  x_3541 & ~n_43729;
assign n_43731 = ~x_3541 &  n_43729;
assign n_43732 = ~n_43730 & ~n_43731;
assign n_43733 =  x_3540 & ~n_26240;
assign n_43734 =  i_29 &  n_26240;
assign n_43735 = ~n_43733 & ~n_43734;
assign n_43736 =  x_3540 & ~n_43735;
assign n_43737 = ~x_3540 &  n_43735;
assign n_43738 = ~n_43736 & ~n_43737;
assign n_43739 =  x_3539 & ~n_26240;
assign n_43740 =  i_28 &  n_26240;
assign n_43741 = ~n_43739 & ~n_43740;
assign n_43742 =  x_3539 & ~n_43741;
assign n_43743 = ~x_3539 &  n_43741;
assign n_43744 = ~n_43742 & ~n_43743;
assign n_43745 =  x_3538 & ~n_26240;
assign n_43746 =  i_27 &  n_26240;
assign n_43747 = ~n_43745 & ~n_43746;
assign n_43748 =  x_3538 & ~n_43747;
assign n_43749 = ~x_3538 &  n_43747;
assign n_43750 = ~n_43748 & ~n_43749;
assign n_43751 =  x_3537 & ~n_26240;
assign n_43752 =  i_26 &  n_26240;
assign n_43753 = ~n_43751 & ~n_43752;
assign n_43754 =  x_3537 & ~n_43753;
assign n_43755 = ~x_3537 &  n_43753;
assign n_43756 = ~n_43754 & ~n_43755;
assign n_43757 =  x_3536 & ~n_26240;
assign n_43758 =  i_25 &  n_26240;
assign n_43759 = ~n_43757 & ~n_43758;
assign n_43760 =  x_3536 & ~n_43759;
assign n_43761 = ~x_3536 &  n_43759;
assign n_43762 = ~n_43760 & ~n_43761;
assign n_43763 =  x_3535 & ~n_26240;
assign n_43764 =  i_24 &  n_26240;
assign n_43765 = ~n_43763 & ~n_43764;
assign n_43766 =  x_3535 & ~n_43765;
assign n_43767 = ~x_3535 &  n_43765;
assign n_43768 = ~n_43766 & ~n_43767;
assign n_43769 =  x_3534 & ~n_26240;
assign n_43770 =  i_23 &  n_26240;
assign n_43771 = ~n_43769 & ~n_43770;
assign n_43772 =  x_3534 & ~n_43771;
assign n_43773 = ~x_3534 &  n_43771;
assign n_43774 = ~n_43772 & ~n_43773;
assign n_43775 =  x_3533 & ~n_26240;
assign n_43776 =  i_22 &  n_26240;
assign n_43777 = ~n_43775 & ~n_43776;
assign n_43778 =  x_3533 & ~n_43777;
assign n_43779 = ~x_3533 &  n_43777;
assign n_43780 = ~n_43778 & ~n_43779;
assign n_43781 =  x_3532 & ~n_26240;
assign n_43782 =  i_21 &  n_26240;
assign n_43783 = ~n_43781 & ~n_43782;
assign n_43784 =  x_3532 & ~n_43783;
assign n_43785 = ~x_3532 &  n_43783;
assign n_43786 = ~n_43784 & ~n_43785;
assign n_43787 =  x_3531 & ~n_26240;
assign n_43788 =  i_20 &  n_26240;
assign n_43789 = ~n_43787 & ~n_43788;
assign n_43790 =  x_3531 & ~n_43789;
assign n_43791 = ~x_3531 &  n_43789;
assign n_43792 = ~n_43790 & ~n_43791;
assign n_43793 =  x_3530 & ~n_26240;
assign n_43794 =  i_19 &  n_26240;
assign n_43795 = ~n_43793 & ~n_43794;
assign n_43796 =  x_3530 & ~n_43795;
assign n_43797 = ~x_3530 &  n_43795;
assign n_43798 = ~n_43796 & ~n_43797;
assign n_43799 =  x_3529 & ~n_26240;
assign n_43800 =  i_18 &  n_26240;
assign n_43801 = ~n_43799 & ~n_43800;
assign n_43802 =  x_3529 & ~n_43801;
assign n_43803 = ~x_3529 &  n_43801;
assign n_43804 = ~n_43802 & ~n_43803;
assign n_43805 =  x_3528 & ~n_26240;
assign n_43806 =  i_17 &  n_26240;
assign n_43807 = ~n_43805 & ~n_43806;
assign n_43808 =  x_3528 & ~n_43807;
assign n_43809 = ~x_3528 &  n_43807;
assign n_43810 = ~n_43808 & ~n_43809;
assign n_43811 =  x_3527 & ~n_26240;
assign n_43812 =  i_16 &  n_26240;
assign n_43813 = ~n_43811 & ~n_43812;
assign n_43814 =  x_3527 & ~n_43813;
assign n_43815 = ~x_3527 &  n_43813;
assign n_43816 = ~n_43814 & ~n_43815;
assign n_43817 =  x_3526 & ~n_26240;
assign n_43818 =  i_15 &  n_26240;
assign n_43819 = ~n_43817 & ~n_43818;
assign n_43820 =  x_3526 & ~n_43819;
assign n_43821 = ~x_3526 &  n_43819;
assign n_43822 = ~n_43820 & ~n_43821;
assign n_43823 =  x_3525 & ~n_26240;
assign n_43824 =  i_14 &  n_26240;
assign n_43825 = ~n_43823 & ~n_43824;
assign n_43826 =  x_3525 & ~n_43825;
assign n_43827 = ~x_3525 &  n_43825;
assign n_43828 = ~n_43826 & ~n_43827;
assign n_43829 =  x_3524 & ~n_26240;
assign n_43830 =  i_13 &  n_26240;
assign n_43831 = ~n_43829 & ~n_43830;
assign n_43832 =  x_3524 & ~n_43831;
assign n_43833 = ~x_3524 &  n_43831;
assign n_43834 = ~n_43832 & ~n_43833;
assign n_43835 =  x_3523 & ~n_26240;
assign n_43836 =  i_12 &  n_26240;
assign n_43837 = ~n_43835 & ~n_43836;
assign n_43838 =  x_3523 & ~n_43837;
assign n_43839 = ~x_3523 &  n_43837;
assign n_43840 = ~n_43838 & ~n_43839;
assign n_43841 =  x_3522 & ~n_26240;
assign n_43842 =  i_11 &  n_26240;
assign n_43843 = ~n_43841 & ~n_43842;
assign n_43844 =  x_3522 & ~n_43843;
assign n_43845 = ~x_3522 &  n_43843;
assign n_43846 = ~n_43844 & ~n_43845;
assign n_43847 =  x_3521 & ~n_26240;
assign n_43848 =  i_10 &  n_26240;
assign n_43849 = ~n_43847 & ~n_43848;
assign n_43850 =  x_3521 & ~n_43849;
assign n_43851 = ~x_3521 &  n_43849;
assign n_43852 = ~n_43850 & ~n_43851;
assign n_43853 =  x_3520 & ~n_26240;
assign n_43854 =  i_9 &  n_26240;
assign n_43855 = ~n_43853 & ~n_43854;
assign n_43856 =  x_3520 & ~n_43855;
assign n_43857 = ~x_3520 &  n_43855;
assign n_43858 = ~n_43856 & ~n_43857;
assign n_43859 =  x_3519 & ~n_26240;
assign n_43860 =  i_8 &  n_26240;
assign n_43861 = ~n_43859 & ~n_43860;
assign n_43862 =  x_3519 & ~n_43861;
assign n_43863 = ~x_3519 &  n_43861;
assign n_43864 = ~n_43862 & ~n_43863;
assign n_43865 =  x_3518 & ~n_26240;
assign n_43866 =  i_7 &  n_26240;
assign n_43867 = ~n_43865 & ~n_43866;
assign n_43868 =  x_3518 & ~n_43867;
assign n_43869 = ~x_3518 &  n_43867;
assign n_43870 = ~n_43868 & ~n_43869;
assign n_43871 =  x_3517 & ~n_26240;
assign n_43872 =  i_6 &  n_26240;
assign n_43873 = ~n_43871 & ~n_43872;
assign n_43874 =  x_3517 & ~n_43873;
assign n_43875 = ~x_3517 &  n_43873;
assign n_43876 = ~n_43874 & ~n_43875;
assign n_43877 =  x_3516 & ~n_26240;
assign n_43878 =  i_5 &  n_26240;
assign n_43879 = ~n_43877 & ~n_43878;
assign n_43880 =  x_3516 & ~n_43879;
assign n_43881 = ~x_3516 &  n_43879;
assign n_43882 = ~n_43880 & ~n_43881;
assign n_43883 =  x_3515 & ~n_26240;
assign n_43884 =  i_4 &  n_26240;
assign n_43885 = ~n_43883 & ~n_43884;
assign n_43886 =  x_3515 & ~n_43885;
assign n_43887 = ~x_3515 &  n_43885;
assign n_43888 = ~n_43886 & ~n_43887;
assign n_43889 =  x_3514 & ~n_26240;
assign n_43890 =  i_3 &  n_26240;
assign n_43891 = ~n_43889 & ~n_43890;
assign n_43892 =  x_3514 & ~n_43891;
assign n_43893 = ~x_3514 &  n_43891;
assign n_43894 = ~n_43892 & ~n_43893;
assign n_43895 =  x_3513 & ~n_26240;
assign n_43896 =  i_2 &  n_26240;
assign n_43897 = ~n_43895 & ~n_43896;
assign n_43898 =  x_3513 & ~n_43897;
assign n_43899 = ~x_3513 &  n_43897;
assign n_43900 = ~n_43898 & ~n_43899;
assign n_43901 =  x_3512 & ~n_26240;
assign n_43902 =  i_1 &  n_26240;
assign n_43903 = ~n_43901 & ~n_43902;
assign n_43904 =  x_3512 & ~n_43903;
assign n_43905 = ~x_3512 &  n_43903;
assign n_43906 = ~n_43904 & ~n_43905;
assign n_43907 =  x_3511 & ~n_6527;
assign n_43908 =  i_32 &  n_6527;
assign n_43909 = ~n_43907 & ~n_43908;
assign n_43910 =  x_3511 & ~n_43909;
assign n_43911 = ~x_3511 &  n_43909;
assign n_43912 = ~n_43910 & ~n_43911;
assign n_43913 =  x_3510 & ~n_6527;
assign n_43914 =  i_31 &  n_6527;
assign n_43915 = ~n_43913 & ~n_43914;
assign n_43916 =  x_3510 & ~n_43915;
assign n_43917 = ~x_3510 &  n_43915;
assign n_43918 = ~n_43916 & ~n_43917;
assign n_43919 =  x_3509 & ~n_6527;
assign n_43920 =  i_30 &  n_6527;
assign n_43921 = ~n_43919 & ~n_43920;
assign n_43922 =  x_3509 & ~n_43921;
assign n_43923 = ~x_3509 &  n_43921;
assign n_43924 = ~n_43922 & ~n_43923;
assign n_43925 =  x_3508 & ~n_6527;
assign n_43926 =  i_29 &  n_6527;
assign n_43927 = ~n_43925 & ~n_43926;
assign n_43928 =  x_3508 & ~n_43927;
assign n_43929 = ~x_3508 &  n_43927;
assign n_43930 = ~n_43928 & ~n_43929;
assign n_43931 =  x_3506 & ~n_6527;
assign n_43932 =  i_27 &  n_6527;
assign n_43933 = ~n_43931 & ~n_43932;
assign n_43934 =  x_3506 & ~n_43933;
assign n_43935 = ~x_3506 &  n_43933;
assign n_43936 = ~n_43934 & ~n_43935;
assign n_43937 =  x_3507 & ~n_6527;
assign n_43938 =  i_28 &  n_6527;
assign n_43939 = ~n_43937 & ~n_43938;
assign n_43940 =  x_3507 & ~n_43939;
assign n_43941 = ~x_3507 &  n_43939;
assign n_43942 = ~n_43940 & ~n_43941;
assign n_43943 = ~n_43936 & ~n_43942;
assign n_43944 = ~n_43930 &  n_43943;
assign n_43945 = ~n_43924 &  n_43944;
assign n_43946 = ~n_43918 &  n_43945;
assign n_43947 = ~n_43912 &  n_43946;
assign n_43948 = ~n_43906 &  n_43947;
assign n_43949 = ~n_43900 &  n_43948;
assign n_43950 = ~n_43894 &  n_43949;
assign n_43951 = ~n_43888 &  n_43950;
assign n_43952 = ~n_43882 &  n_43951;
assign n_43953 = ~n_43876 &  n_43952;
assign n_43954 = ~n_43870 &  n_43953;
assign n_43955 = ~n_43864 &  n_43954;
assign n_43956 = ~n_43858 &  n_43955;
assign n_43957 = ~n_43852 &  n_43956;
assign n_43958 = ~n_43846 &  n_43957;
assign n_43959 = ~n_43840 &  n_43958;
assign n_43960 = ~n_43834 &  n_43959;
assign n_43961 = ~n_43828 &  n_43960;
assign n_43962 = ~n_43822 &  n_43961;
assign n_43963 = ~n_43816 &  n_43962;
assign n_43964 = ~n_43810 &  n_43963;
assign n_43965 = ~n_43804 &  n_43964;
assign n_43966 = ~n_43798 &  n_43965;
assign n_43967 = ~n_43792 &  n_43966;
assign n_43968 = ~n_43786 &  n_43967;
assign n_43969 = ~n_43780 &  n_43968;
assign n_43970 = ~n_43774 &  n_43969;
assign n_43971 = ~n_43768 &  n_43970;
assign n_43972 = ~n_43762 &  n_43971;
assign n_43973 = ~n_43756 &  n_43972;
assign n_43974 = ~n_43750 &  n_43973;
assign n_43975 = ~n_43744 &  n_43974;
assign n_43976 = ~n_43738 &  n_43975;
assign n_43977 = ~n_43732 &  n_43976;
assign n_43978 = ~n_43726 &  n_43977;
assign n_43979 = ~n_43720 &  n_43978;
assign n_43980 = ~n_43714 &  n_43979;
assign n_43981 = ~n_43704 &  n_43980;
assign n_43982 = ~n_43694 &  n_43981;
assign n_43983 = ~n_43684 &  n_43982;
assign n_43984 = ~n_43674 &  n_43983;
assign n_43985 = ~n_43664 &  n_43984;
assign n_43986 = ~n_43654 &  n_43985;
assign n_43987 = ~n_43644 &  n_43986;
assign n_43988 = ~n_43634 &  n_43987;
assign n_43989 = ~n_43624 &  n_43988;
assign n_43990 = ~n_43614 &  n_43989;
assign n_43991 = ~n_43604 &  n_43990;
assign n_43992 = ~n_43594 &  n_43991;
assign n_43993 = ~n_43584 &  n_43992;
assign n_43994 = ~n_43574 &  n_43993;
assign n_43995 = ~n_43564 &  n_43994;
assign n_43996 = ~n_43554 &  n_43995;
assign n_43997 = ~n_43544 &  n_43996;
assign n_43998 = ~n_43534 &  n_43997;
assign n_43999 = ~n_43524 &  n_43998;
assign n_44000 = ~n_43514 &  n_43999;
assign n_44001 = ~n_43504 &  n_44000;
assign n_44002 = ~n_43494 &  n_44001;
assign n_44003 = ~n_43484 &  n_44002;
assign n_44004 = ~n_43474 &  n_44003;
assign n_44005 = ~n_43464 &  n_44004;
assign n_44006 = ~n_43454 &  n_44005;
assign n_44007 = ~n_43444 &  n_44006;
assign n_44008 = ~n_43434 &  n_44007;
assign n_44009 = ~n_43424 &  n_44008;
assign n_44010 = ~n_43414 &  n_44009;
assign n_44011 = ~n_43404 &  n_44010;
assign n_44012 = ~n_43392 &  n_44011;
assign n_44013 = ~n_43382 &  n_44012;
assign n_44014 = ~n_43372 &  n_44013;
assign n_44015 = ~n_43362 &  n_44014;
assign n_44016 = ~n_43352 &  n_44015;
assign n_44017 = ~n_43342 &  n_44016;
assign n_44018 = ~n_43332 &  n_44017;
assign n_44019 = ~n_43322 &  n_44018;
assign n_44020 = ~n_43312 &  n_44019;
assign n_44021 = ~n_43302 &  n_44020;
assign n_44022 = ~n_43292 &  n_44021;
assign n_44023 = ~n_43282 &  n_44022;
assign n_44024 = ~n_43272 &  n_44023;
assign n_44025 = ~n_43262 &  n_44024;
assign n_44026 = ~n_43252 &  n_44025;
assign n_44027 = ~n_43242 &  n_44026;
assign n_44028 = ~n_43232 &  n_44027;
assign n_44029 = ~n_43222 &  n_44028;
assign n_44030 = ~n_43212 &  n_44029;
assign n_44031 = ~n_43202 &  n_44030;
assign n_44032 = ~n_43192 &  n_44031;
assign n_44033 = ~n_43182 &  n_44032;
assign n_44034 = ~n_43172 &  n_44033;
assign n_44035 = ~n_43162 &  n_44034;
assign n_44036 = ~n_43152 &  n_44035;
assign n_44037 = ~n_43142 &  n_44036;
assign n_44038 = ~n_43132 &  n_44037;
assign n_44039 = ~n_43122 &  n_44038;
assign n_44040 = ~n_43112 &  n_44039;
assign n_44041 = ~n_43102 &  n_44040;
assign n_44042 = ~n_43092 &  n_44041;
assign n_44043 = ~n_43082 &  n_44042;
assign n_44044 = ~n_43070 &  n_44043;
assign n_44045 = ~n_43064 &  n_44044;
assign n_44046 = ~n_43058 &  n_44045;
assign n_44047 = ~n_43052 &  n_44046;
assign n_44048 = ~n_43046 &  n_44047;
assign n_44049 = ~n_43040 &  n_44048;
assign n_44050 = ~n_43034 &  n_44049;
assign n_44051 = ~n_43028 &  n_44050;
assign n_44052 = ~n_43022 &  n_44051;
assign n_44053 = ~n_43016 &  n_44052;
assign n_44054 = ~n_43010 &  n_44053;
assign n_44055 = ~n_43004 &  n_44054;
assign n_44056 = ~n_42998 &  n_44055;
assign n_44057 = ~n_42992 &  n_44056;
assign n_44058 = ~n_42986 &  n_44057;
assign n_44059 = ~n_42980 &  n_44058;
assign n_44060 = ~n_42974 &  n_44059;
assign n_44061 = ~n_42968 &  n_44060;
assign n_44062 = ~n_42962 &  n_44061;
assign n_44063 = ~n_42956 &  n_44062;
assign n_44064 = ~n_42950 &  n_44063;
assign n_44065 = ~n_42944 &  n_44064;
assign n_44066 = ~n_42938 &  n_44065;
assign n_44067 = ~n_42932 &  n_44066;
assign n_44068 = ~n_42926 &  n_44067;
assign n_44069 = ~n_42920 &  n_44068;
assign n_44070 = ~n_42914 &  n_44069;
assign n_44071 = ~n_42908 &  n_44070;
assign n_44072 = ~n_42902 &  n_44071;
assign n_44073 = ~n_42896 &  n_44072;
assign n_44074 = ~n_42890 &  n_44073;
assign n_44075 = ~n_42884 &  n_44074;
assign n_44076 = ~n_42878 &  n_44075;
assign n_44077 = ~n_42864 &  n_44076;
assign n_44078 = ~n_42850 &  n_44077;
assign n_44079 = ~n_42836 &  n_44078;
assign n_44080 = ~n_42822 &  n_44079;
assign n_44081 = ~n_42808 &  n_44080;
assign n_44082 = ~n_42794 &  n_44081;
assign n_44083 = ~n_42780 &  n_44082;
assign n_44084 = ~n_42766 &  n_44083;
assign n_44085 = ~n_42752 &  n_44084;
assign n_44086 = ~n_42738 &  n_44085;
assign n_44087 = ~n_42724 &  n_44086;
assign n_44088 = ~n_42710 &  n_44087;
assign n_44089 = ~n_42696 &  n_44088;
assign n_44090 = ~n_42682 &  n_44089;
assign n_44091 = ~n_42668 &  n_44090;
assign n_44092 = ~n_42654 &  n_44091;
assign n_44093 = ~n_42640 &  n_44092;
assign n_44094 = ~n_42626 &  n_44093;
assign n_44095 = ~n_42612 &  n_44094;
assign n_44096 = ~n_42598 &  n_44095;
assign n_44097 = ~n_42584 &  n_44096;
assign n_44098 = ~n_42570 &  n_44097;
assign n_44099 = ~n_42556 &  n_44098;
assign n_44100 = ~n_42542 &  n_44099;
assign n_44101 = ~n_42528 &  n_44100;
assign n_44102 = ~n_42514 &  n_44101;
assign n_44103 = ~n_42500 &  n_44102;
assign n_44104 = ~n_42486 &  n_44103;
assign n_44105 = ~n_42472 &  n_44104;
assign n_44106 = ~n_42458 &  n_44105;
assign n_44107 = ~n_42444 &  n_44106;
assign n_44108 = ~n_42424 &  n_44107;
assign n_44109 = ~n_42412 &  n_44108;
assign n_44110 = ~n_42400 &  n_44109;
assign n_44111 = ~n_42388 &  n_44110;
assign n_44112 = ~n_42376 &  n_44111;
assign n_44113 = ~n_42364 &  n_44112;
assign n_44114 = ~n_42352 &  n_44113;
assign n_44115 = ~n_42340 &  n_44114;
assign n_44116 = ~n_42328 &  n_44115;
assign n_44117 = ~n_42316 &  n_44116;
assign n_44118 = ~n_42304 &  n_44117;
assign n_44119 = ~n_42292 &  n_44118;
assign n_44120 = ~n_42280 &  n_44119;
assign n_44121 = ~n_42268 &  n_44120;
assign n_44122 = ~n_42256 &  n_44121;
assign n_44123 = ~n_42244 &  n_44122;
assign n_44124 = ~n_42232 &  n_44123;
assign n_44125 = ~n_42220 &  n_44124;
assign n_44126 = ~n_42208 &  n_44125;
assign n_44127 = ~n_42196 &  n_44126;
assign n_44128 = ~n_42184 &  n_44127;
assign n_44129 = ~n_42172 &  n_44128;
assign n_44130 = ~n_42160 &  n_44129;
assign n_44131 = ~n_42148 &  n_44130;
assign n_44132 = ~n_42136 &  n_44131;
assign n_44133 = ~n_42124 &  n_44132;
assign n_44134 = ~n_42112 &  n_44133;
assign n_44135 = ~n_42100 &  n_44134;
assign n_44136 = ~n_42088 &  n_44135;
assign n_44137 = ~n_42076 &  n_44136;
assign n_44138 = ~n_42064 &  n_44137;
assign n_44139 = ~n_42052 &  n_44138;
assign n_44140 = ~n_42037 &  n_44139;
assign n_44141 = ~n_42031 &  n_44140;
assign n_44142 = ~n_42025 &  n_44141;
assign n_44143 = ~n_42019 &  n_44142;
assign n_44144 = ~n_42013 &  n_44143;
assign n_44145 = ~n_42007 &  n_44144;
assign n_44146 = ~n_42001 &  n_44145;
assign n_44147 = ~n_41995 &  n_44146;
assign n_44148 = ~n_41989 &  n_44147;
assign n_44149 = ~n_41983 &  n_44148;
assign n_44150 = ~n_41977 &  n_44149;
assign n_44151 = ~n_41971 &  n_44150;
assign n_44152 = ~n_41965 &  n_44151;
assign n_44153 = ~n_41959 &  n_44152;
assign n_44154 = ~n_41953 &  n_44153;
assign n_44155 = ~n_41947 &  n_44154;
assign n_44156 = ~n_41941 &  n_44155;
assign n_44157 = ~n_41935 &  n_44156;
assign n_44158 = ~n_41929 &  n_44157;
assign n_44159 = ~n_41923 &  n_44158;
assign n_44160 = ~n_41917 &  n_44159;
assign n_44161 = ~n_41911 &  n_44160;
assign n_44162 = ~n_41905 &  n_44161;
assign n_44163 = ~n_41899 &  n_44162;
assign n_44164 = ~n_41893 &  n_44163;
assign n_44165 = ~n_41887 &  n_44164;
assign n_44166 = ~n_41881 &  n_44165;
assign n_44167 = ~n_41875 &  n_44166;
assign n_44168 = ~n_41869 &  n_44167;
assign n_44169 = ~n_41863 &  n_44168;
assign n_44170 = ~n_41857 &  n_44169;
assign n_44171 = ~n_41851 &  n_44170;
assign n_44172 = ~n_41845 &  n_44171;
assign n_44173 = ~n_41839 &  n_44172;
assign n_44174 = ~n_41833 &  n_44173;
assign n_44175 = ~n_41827 &  n_44174;
assign n_44176 = ~n_41821 &  n_44175;
assign n_44177 = ~n_41815 &  n_44176;
assign n_44178 = ~n_41809 &  n_44177;
assign n_44179 = ~n_41803 &  n_44178;
assign n_44180 = ~n_41797 &  n_44179;
assign n_44181 = ~n_41791 &  n_44180;
assign n_44182 = ~n_41785 &  n_44181;
assign n_44183 = ~n_41779 &  n_44182;
assign n_44184 = ~n_41773 &  n_44183;
assign n_44185 = ~n_41767 &  n_44184;
assign n_44186 = ~n_41761 &  n_44185;
assign n_44187 = ~n_41755 &  n_44186;
assign n_44188 = ~n_41749 &  n_44187;
assign n_44189 = ~n_41743 &  n_44188;
assign n_44190 = ~n_41737 &  n_44189;
assign n_44191 = ~n_41731 &  n_44190;
assign n_44192 = ~n_41725 &  n_44191;
assign n_44193 = ~n_41719 &  n_44192;
assign n_44194 = ~n_41713 &  n_44193;
assign n_44195 = ~n_41707 &  n_44194;
assign n_44196 = ~n_41701 &  n_44195;
assign n_44197 = ~n_41695 &  n_44196;
assign n_44198 = ~n_41689 &  n_44197;
assign n_44199 = ~n_41683 &  n_44198;
assign n_44200 = ~n_41677 &  n_44199;
assign n_44201 = ~n_41671 &  n_44200;
assign n_44202 = ~n_41665 &  n_44201;
assign n_44203 = ~n_41659 &  n_44202;
assign n_44204 = ~n_41653 &  n_44203;
assign n_44205 = ~n_41641 &  n_44204;
assign n_44206 = ~n_41629 &  n_44205;
assign n_44207 = ~n_41617 &  n_44206;
assign n_44208 = ~n_41605 &  n_44207;
assign n_44209 = ~n_41593 &  n_44208;
assign n_44210 = ~n_41581 &  n_44209;
assign n_44211 = ~n_41569 &  n_44210;
assign n_44212 = ~n_41557 &  n_44211;
assign n_44213 = ~n_41545 &  n_44212;
assign n_44214 = ~n_41533 &  n_44213;
assign n_44215 = ~n_41521 &  n_44214;
assign n_44216 = ~n_41509 &  n_44215;
assign n_44217 = ~n_41497 &  n_44216;
assign n_44218 = ~n_41485 &  n_44217;
assign n_44219 = ~n_41473 &  n_44218;
assign n_44220 = ~n_41461 &  n_44219;
assign n_44221 = ~n_41449 &  n_44220;
assign n_44222 = ~n_41437 &  n_44221;
assign n_44223 = ~n_41425 &  n_44222;
assign n_44224 = ~n_41413 &  n_44223;
assign n_44225 = ~n_41401 &  n_44224;
assign n_44226 = ~n_41389 &  n_44225;
assign n_44227 = ~n_41377 &  n_44226;
assign n_44228 = ~n_41365 &  n_44227;
assign n_44229 = ~n_41353 &  n_44228;
assign n_44230 = ~n_41341 &  n_44229;
assign n_44231 = ~n_41329 &  n_44230;
assign n_44232 = ~n_41317 &  n_44231;
assign n_44233 = ~n_41305 &  n_44232;
assign n_44234 = ~n_41293 &  n_44233;
assign n_44235 = ~n_41281 &  n_44234;
assign n_44236 = ~n_41266 &  n_44235;
assign n_44237 = ~n_41262 &  n_44236;
assign n_44238 = ~n_41258 &  n_44237;
assign n_44239 = ~n_41254 &  n_44238;
assign n_44240 = ~n_41250 &  n_44239;
assign n_44241 = ~n_41246 &  n_44240;
assign n_44242 = ~n_41242 &  n_44241;
assign n_44243 = ~n_41238 &  n_44242;
assign n_44244 = ~n_41234 &  n_44243;
assign n_44245 = ~n_41230 &  n_44244;
assign n_44246 = ~n_41226 &  n_44245;
assign n_44247 = ~n_41222 &  n_44246;
assign n_44248 = ~n_41218 &  n_44247;
assign n_44249 = ~n_41214 &  n_44248;
assign n_44250 = ~n_41210 &  n_44249;
assign n_44251 = ~n_41206 &  n_44250;
assign n_44252 = ~n_41202 &  n_44251;
assign n_44253 = ~n_41198 &  n_44252;
assign n_44254 = ~n_41194 &  n_44253;
assign n_44255 = ~n_41190 &  n_44254;
assign n_44256 = ~n_41186 &  n_44255;
assign n_44257 = ~n_41182 &  n_44256;
assign n_44258 = ~n_41178 &  n_44257;
assign n_44259 = ~n_41174 &  n_44258;
assign n_44260 = ~n_41170 &  n_44259;
assign n_44261 = ~n_41166 &  n_44260;
assign n_44262 = ~n_41162 &  n_44261;
assign n_44263 = ~n_41158 &  n_44262;
assign n_44264 = ~n_41154 &  n_44263;
assign n_44265 = ~n_41150 &  n_44264;
assign n_44266 = ~n_41146 &  n_44265;
assign n_44267 = ~n_41142 &  n_44266;
assign n_44268 = ~n_41138 &  n_44267;
assign n_44269 = ~n_41132 &  n_44268;
assign n_44270 = ~n_41126 &  n_44269;
assign n_44271 = ~n_41120 &  n_44270;
assign n_44272 = ~n_41114 &  n_44271;
assign n_44273 = ~n_41108 &  n_44272;
assign n_44274 = ~n_41102 &  n_44273;
assign n_44275 = ~n_41096 &  n_44274;
assign n_44276 = ~n_41090 &  n_44275;
assign n_44277 = ~n_41084 &  n_44276;
assign n_44278 = ~n_41078 &  n_44277;
assign n_44279 = ~n_41072 &  n_44278;
assign n_44280 = ~n_41066 &  n_44279;
assign n_44281 = ~n_41060 &  n_44280;
assign n_44282 = ~n_41054 &  n_44281;
assign n_44283 = ~n_41048 &  n_44282;
assign n_44284 = ~n_41042 &  n_44283;
assign n_44285 = ~n_41036 &  n_44284;
assign n_44286 = ~n_41030 &  n_44285;
assign n_44287 = ~n_41024 &  n_44286;
assign n_44288 = ~n_41018 &  n_44287;
assign n_44289 = ~n_41012 &  n_44288;
assign n_44290 = ~n_41006 &  n_44289;
assign n_44291 = ~n_41000 &  n_44290;
assign n_44292 = ~n_40994 &  n_44291;
assign n_44293 = ~n_40988 &  n_44292;
assign n_44294 = ~n_40982 &  n_44293;
assign n_44295 = ~n_40976 &  n_44294;
assign n_44296 = ~n_40970 &  n_44295;
assign n_44297 = ~n_40964 &  n_44296;
assign n_44298 = ~n_40958 &  n_44297;
assign n_44299 = ~n_40952 &  n_44298;
assign n_44300 = ~n_40946 &  n_44299;
assign n_44301 = ~n_40932 &  n_44300;
assign n_44302 = ~n_40917 &  n_44301;
assign n_44303 = ~n_40902 &  n_44302;
assign n_44304 = ~n_40887 &  n_44303;
assign n_44305 = ~n_40872 &  n_44304;
assign n_44306 = ~n_40857 &  n_44305;
assign n_44307 = ~n_40842 &  n_44306;
assign n_44308 = ~n_40827 &  n_44307;
assign n_44309 = ~n_40812 &  n_44308;
assign n_44310 = ~n_40797 &  n_44309;
assign n_44311 = ~n_40782 &  n_44310;
assign n_44312 = ~n_40767 &  n_44311;
assign n_44313 = ~n_40752 &  n_44312;
assign n_44314 = ~n_40737 &  n_44313;
assign n_44315 = ~n_40722 &  n_44314;
assign n_44316 = ~n_40707 &  n_44315;
assign n_44317 = ~n_40692 &  n_44316;
assign n_44318 = ~n_40677 &  n_44317;
assign n_44319 = ~n_40662 &  n_44318;
assign n_44320 = ~n_40647 &  n_44319;
assign n_44321 = ~n_40632 &  n_44320;
assign n_44322 = ~n_40617 &  n_44321;
assign n_44323 = ~n_40602 &  n_44322;
assign n_44324 = ~n_40587 &  n_44323;
assign n_44325 = ~n_40572 &  n_44324;
assign n_44326 = ~n_40557 &  n_44325;
assign n_44327 = ~n_40542 &  n_44326;
assign n_44328 = ~n_40527 &  n_44327;
assign n_44329 = ~n_40512 &  n_44328;
assign n_44330 = ~n_40497 &  n_44329;
assign n_44331 = ~n_40482 &  n_44330;
assign n_44332 = ~n_40467 &  n_44331;
assign n_44333 = ~n_40463 &  n_44332;
assign n_44334 = ~n_40459 &  n_44333;
assign n_44335 = ~n_40455 &  n_44334;
assign n_44336 = ~n_40451 &  n_44335;
assign n_44337 = ~n_40447 &  n_44336;
assign n_44338 = ~n_40443 &  n_44337;
assign n_44339 = ~n_40439 &  n_44338;
assign n_44340 = ~n_40435 &  n_44339;
assign n_44341 = ~n_40431 &  n_44340;
assign n_44342 = ~n_40427 &  n_44341;
assign n_44343 = ~n_40423 &  n_44342;
assign n_44344 = ~n_40419 &  n_44343;
assign n_44345 = ~n_40415 &  n_44344;
assign n_44346 = ~n_40411 &  n_44345;
assign n_44347 = ~n_40406 &  n_44346;
assign n_44348 = ~n_40400 &  n_44347;
assign n_44349 = ~n_40394 &  n_44348;
assign n_44350 = ~n_40388 &  n_44349;
assign n_44351 = ~n_40382 &  n_44350;
assign n_44352 = ~n_40376 &  n_44351;
assign n_44353 = ~n_40370 &  n_44352;
assign n_44354 = ~n_40364 &  n_44353;
assign n_44355 = ~n_40358 &  n_44354;
assign n_44356 = ~n_40352 &  n_44355;
assign n_44357 = ~n_40346 &  n_44356;
assign n_44358 = ~n_40340 &  n_44357;
assign n_44359 = ~n_40334 &  n_44358;
assign n_44360 = ~n_40328 &  n_44359;
assign n_44361 = ~n_40322 &  n_44360;
assign n_44362 = ~n_40316 &  n_44361;
assign n_44363 = ~n_40310 &  n_44362;
assign n_44364 = ~n_40304 &  n_44363;
assign n_44365 = ~n_40298 &  n_44364;
assign n_44366 = ~n_40292 &  n_44365;
assign n_44367 = ~n_40286 &  n_44366;
assign n_44368 = ~n_40280 &  n_44367;
assign n_44369 = ~n_40274 &  n_44368;
assign n_44370 = ~n_40268 &  n_44369;
assign n_44371 = ~n_40262 &  n_44370;
assign n_44372 = ~n_40256 &  n_44371;
assign n_44373 = ~n_40250 &  n_44372;
assign n_44374 = ~n_40244 &  n_44373;
assign n_44375 = ~n_40238 &  n_44374;
assign n_44376 = ~n_40232 &  n_44375;
assign n_44377 = ~n_40226 &  n_44376;
assign n_44378 = ~n_40220 &  n_44377;
assign n_44379 = ~n_40214 &  n_44378;
assign n_44380 = ~n_40208 &  n_44379;
assign n_44381 = ~n_40200 &  n_44380;
assign n_44382 = ~n_40194 &  n_44381;
assign n_44383 = ~n_40188 &  n_44382;
assign n_44384 = ~n_40182 &  n_44383;
assign n_44385 = ~n_40176 &  n_44384;
assign n_44386 = ~n_40170 &  n_44385;
assign n_44387 = ~n_40164 &  n_44386;
assign n_44388 = ~n_40158 &  n_44387;
assign n_44389 = ~n_40152 &  n_44388;
assign n_44390 = ~n_40146 &  n_44389;
assign n_44391 = ~n_40140 &  n_44390;
assign n_44392 = ~n_40134 &  n_44391;
assign n_44393 = ~n_40128 &  n_44392;
assign n_44394 = ~n_40122 &  n_44393;
assign n_44395 = ~n_40116 &  n_44394;
assign n_44396 = ~n_40110 &  n_44395;
assign n_44397 = ~n_40104 &  n_44396;
assign n_44398 = ~n_40098 &  n_44397;
assign n_44399 = ~n_40092 &  n_44398;
assign n_44400 = ~n_40086 &  n_44399;
assign n_44401 = ~n_40080 &  n_44400;
assign n_44402 = ~n_40074 &  n_44401;
assign n_44403 = ~n_40068 &  n_44402;
assign n_44404 = ~n_40062 &  n_44403;
assign n_44405 = ~n_40056 &  n_44404;
assign n_44406 = ~n_40050 &  n_44405;
assign n_44407 = ~n_40044 &  n_44406;
assign n_44408 = ~n_40038 &  n_44407;
assign n_44409 = ~n_40032 &  n_44408;
assign n_44410 = ~n_40026 &  n_44409;
assign n_44411 = ~n_40020 &  n_44410;
assign n_44412 = ~n_40014 &  n_44411;
assign n_44413 = ~n_40008 &  n_44412;
assign n_44414 = ~n_40004 &  n_44413;
assign n_44415 = ~n_39998 &  n_44414;
assign n_44416 = ~n_39992 &  n_44415;
assign n_44417 = ~n_39986 &  n_44416;
assign n_44418 = ~n_39980 &  n_44417;
assign n_44419 = ~n_39974 &  n_44418;
assign n_44420 = ~n_39968 &  n_44419;
assign n_44421 = ~n_39962 &  n_44420;
assign n_44422 = ~n_39956 &  n_44421;
assign n_44423 = ~n_39950 &  n_44422;
assign n_44424 = ~n_39944 &  n_44423;
assign n_44425 = ~n_39938 &  n_44424;
assign n_44426 = ~n_39932 &  n_44425;
assign n_44427 = ~n_39926 &  n_44426;
assign n_44428 = ~n_39920 &  n_44427;
assign n_44429 = ~n_39914 &  n_44428;
assign n_44430 = ~n_39908 &  n_44429;
assign n_44431 = ~n_39902 &  n_44430;
assign n_44432 = ~n_39896 &  n_44431;
assign n_44433 = ~n_39890 &  n_44432;
assign n_44434 = ~n_39884 &  n_44433;
assign n_44435 = ~n_39878 &  n_44434;
assign n_44436 = ~n_39872 &  n_44435;
assign n_44437 = ~n_39866 &  n_44436;
assign n_44438 = ~n_39860 &  n_44437;
assign n_44439 = ~n_39854 &  n_44438;
assign n_44440 = ~n_39848 &  n_44439;
assign n_44441 = ~n_39842 &  n_44440;
assign n_44442 = ~n_39836 &  n_44441;
assign n_44443 = ~n_39830 &  n_44442;
assign n_44444 = ~n_39824 &  n_44443;
assign n_44445 = ~n_39818 &  n_44444;
assign n_44446 = ~n_39814 &  n_44445;
assign n_44447 = ~n_39810 &  n_44446;
assign n_44448 = ~n_39806 &  n_44447;
assign n_44449 = ~n_39802 &  n_44448;
assign n_44450 = ~n_39798 &  n_44449;
assign n_44451 = ~n_39794 &  n_44450;
assign n_44452 = ~n_39790 &  n_44451;
assign n_44453 = ~n_39786 &  n_44452;
assign n_44454 = ~n_39782 &  n_44453;
assign n_44455 = ~n_39778 &  n_44454;
assign n_44456 = ~n_39774 &  n_44455;
assign n_44457 = ~n_39770 &  n_44456;
assign n_44458 = ~n_39766 &  n_44457;
assign n_44459 = ~n_39762 &  n_44458;
assign n_44460 = ~n_39758 &  n_44459;
assign n_44461 = ~n_39754 &  n_44460;
assign n_44462 = ~n_39750 &  n_44461;
assign n_44463 = ~n_39746 &  n_44462;
assign n_44464 = ~n_39742 &  n_44463;
assign n_44465 = ~n_39738 &  n_44464;
assign n_44466 = ~n_39734 &  n_44465;
assign n_44467 = ~n_39730 &  n_44466;
assign n_44468 = ~n_39726 &  n_44467;
assign n_44469 = ~n_39722 &  n_44468;
assign n_44470 = ~n_39718 &  n_44469;
assign n_44471 = ~n_39714 &  n_44470;
assign n_44472 = ~n_39710 &  n_44471;
assign n_44473 = ~n_39706 &  n_44472;
assign n_44474 = ~n_39702 &  n_44473;
assign n_44475 = ~n_39698 &  n_44474;
assign n_44476 = ~n_39694 &  n_44475;
assign n_44477 = ~n_39690 &  n_44476;
assign n_44478 = ~n_39684 &  n_44477;
assign n_44479 = ~n_39678 &  n_44478;
assign n_44480 = ~n_39672 &  n_44479;
assign n_44481 = ~n_39666 &  n_44480;
assign n_44482 = ~n_39660 &  n_44481;
assign n_44483 = ~n_39654 &  n_44482;
assign n_44484 = ~n_39648 &  n_44483;
assign n_44485 = ~n_39642 &  n_44484;
assign n_44486 = ~n_39636 &  n_44485;
assign n_44487 = ~n_39630 &  n_44486;
assign n_44488 = ~n_39624 &  n_44487;
assign n_44489 = ~n_39618 &  n_44488;
assign n_44490 = ~n_39612 &  n_44489;
assign n_44491 = ~n_39606 &  n_44490;
assign n_44492 = ~n_39600 &  n_44491;
assign n_44493 = ~n_39594 &  n_44492;
assign n_44494 = ~n_39588 &  n_44493;
assign n_44495 = ~n_39582 &  n_44494;
assign n_44496 = ~n_39576 &  n_44495;
assign n_44497 = ~n_39570 &  n_44496;
assign n_44498 = ~n_39564 &  n_44497;
assign n_44499 = ~n_39558 &  n_44498;
assign n_44500 = ~n_39552 &  n_44499;
assign n_44501 = ~n_39546 &  n_44500;
assign n_44502 = ~n_39540 &  n_44501;
assign n_44503 = ~n_39534 &  n_44502;
assign n_44504 = ~n_39528 &  n_44503;
assign n_44505 = ~n_39522 &  n_44504;
assign n_44506 = ~n_39516 &  n_44505;
assign n_44507 = ~n_39510 &  n_44506;
assign n_44508 = ~n_39504 &  n_44507;
assign n_44509 = ~n_39497 &  n_44508;
assign n_44510 = ~n_39491 &  n_44509;
assign n_44511 = ~n_39485 &  n_44510;
assign n_44512 = ~n_39479 &  n_44511;
assign n_44513 = ~n_39473 &  n_44512;
assign n_44514 = ~n_39467 &  n_44513;
assign n_44515 = ~n_39461 &  n_44514;
assign n_44516 = ~n_39455 &  n_44515;
assign n_44517 = ~n_39449 &  n_44516;
assign n_44518 = ~n_39443 &  n_44517;
assign n_44519 = ~n_39437 &  n_44518;
assign n_44520 = ~n_39431 &  n_44519;
assign n_44521 = ~n_39425 &  n_44520;
assign n_44522 = ~n_39419 &  n_44521;
assign n_44523 = ~n_39413 &  n_44522;
assign n_44524 = ~n_39407 &  n_44523;
assign n_44525 = ~n_39401 &  n_44524;
assign n_44526 = ~n_39395 &  n_44525;
assign n_44527 = ~n_39389 &  n_44526;
assign n_44528 = ~n_39383 &  n_44527;
assign n_44529 = ~n_39377 &  n_44528;
assign n_44530 = ~n_39371 &  n_44529;
assign n_44531 = ~n_39365 &  n_44530;
assign n_44532 = ~n_39359 &  n_44531;
assign n_44533 = ~n_39353 &  n_44532;
assign n_44534 = ~n_39347 &  n_44533;
assign n_44535 = ~n_39341 &  n_44534;
assign n_44536 = ~n_39335 &  n_44535;
assign n_44537 = ~n_39329 &  n_44536;
assign n_44538 = ~n_39323 &  n_44537;
assign n_44539 = ~n_39317 &  n_44538;
assign n_44540 = ~n_39311 &  n_44539;
assign n_44541 = ~n_39305 &  n_44540;
assign n_44542 = ~n_39299 &  n_44541;
assign n_44543 = ~n_39293 &  n_44542;
assign n_44544 = ~n_39287 &  n_44543;
assign n_44545 = ~n_39281 &  n_44544;
assign n_44546 = ~n_39275 &  n_44545;
assign n_44547 = ~n_39269 &  n_44546;
assign n_44548 = ~n_39263 &  n_44547;
assign n_44549 = ~n_39257 &  n_44548;
assign n_44550 = ~n_39251 &  n_44549;
assign n_44551 = ~n_39245 &  n_44550;
assign n_44552 = ~n_39239 &  n_44551;
assign n_44553 = ~n_39233 &  n_44552;
assign n_44554 = ~n_39227 &  n_44553;
assign n_44555 = ~n_39221 &  n_44554;
assign n_44556 = ~n_39215 &  n_44555;
assign n_44557 = ~n_39209 &  n_44556;
assign n_44558 = ~n_39203 &  n_44557;
assign n_44559 = ~n_39197 &  n_44558;
assign n_44560 = ~n_39191 &  n_44559;
assign n_44561 = ~n_39185 &  n_44560;
assign n_44562 = ~n_39179 &  n_44561;
assign n_44563 = ~n_39173 &  n_44562;
assign n_44564 = ~n_39167 &  n_44563;
assign n_44565 = ~n_39161 &  n_44564;
assign n_44566 = ~n_39155 &  n_44565;
assign n_44567 = ~n_39149 &  n_44566;
assign n_44568 = ~n_39143 &  n_44567;
assign n_44569 = ~n_39137 &  n_44568;
assign n_44570 = ~n_39131 &  n_44569;
assign n_44571 = ~n_39125 &  n_44570;
assign n_44572 = ~n_39119 &  n_44571;
assign n_44573 = ~n_39113 &  n_44572;
assign n_44574 = ~n_39107 &  n_44573;
assign n_44575 = ~n_39101 &  n_44574;
assign n_44576 = ~n_39095 &  n_44575;
assign n_44577 = ~n_39089 &  n_44576;
assign n_44578 = ~n_39083 &  n_44577;
assign n_44579 = ~n_39077 &  n_44578;
assign n_44580 = ~n_39071 &  n_44579;
assign n_44581 = ~n_39065 &  n_44580;
assign n_44582 = ~n_39059 &  n_44581;
assign n_44583 = ~n_39053 &  n_44582;
assign n_44584 = ~n_39047 &  n_44583;
assign n_44585 = ~n_39041 &  n_44584;
assign n_44586 = ~n_39035 &  n_44585;
assign n_44587 = ~n_39029 &  n_44586;
assign n_44588 = ~n_39023 &  n_44587;
assign n_44589 = ~n_39017 &  n_44588;
assign n_44590 = ~n_39011 &  n_44589;
assign n_44591 = ~n_39005 &  n_44590;
assign n_44592 = ~n_38999 &  n_44591;
assign n_44593 = ~n_38993 &  n_44592;
assign n_44594 = ~n_38987 &  n_44593;
assign n_44595 = ~n_38981 &  n_44594;
assign n_44596 = ~n_38975 &  n_44595;
assign n_44597 = ~n_38969 &  n_44596;
assign n_44598 = ~n_38963 &  n_44597;
assign n_44599 = ~n_38957 &  n_44598;
assign n_44600 = ~n_38951 &  n_44599;
assign n_44601 = ~n_38945 &  n_44600;
assign n_44602 = ~n_38939 &  n_44601;
assign n_44603 = ~n_38933 &  n_44602;
assign n_44604 = ~n_38927 &  n_44603;
assign n_44605 = ~n_38920 &  n_44604;
assign n_44606 = ~n_38916 &  n_44605;
assign n_44607 = ~n_38912 &  n_44606;
assign n_44608 = ~n_38908 &  n_44607;
assign n_44609 = ~n_38904 &  n_44608;
assign n_44610 = ~n_38900 &  n_44609;
assign n_44611 = ~n_38896 &  n_44610;
assign n_44612 = ~n_38892 &  n_44611;
assign n_44613 = ~n_38888 &  n_44612;
assign n_44614 = ~n_38884 &  n_44613;
assign n_44615 = ~n_38880 &  n_44614;
assign n_44616 = ~n_38876 &  n_44615;
assign n_44617 = ~n_38872 &  n_44616;
assign n_44618 = ~n_38868 &  n_44617;
assign n_44619 = ~n_38864 &  n_44618;
assign n_44620 = ~n_38860 &  n_44619;
assign n_44621 = ~n_38856 &  n_44620;
assign n_44622 = ~n_38852 &  n_44621;
assign n_44623 = ~n_38848 &  n_44622;
assign n_44624 = ~n_38844 &  n_44623;
assign n_44625 = ~n_38840 &  n_44624;
assign n_44626 = ~n_38836 &  n_44625;
assign n_44627 = ~n_38832 &  n_44626;
assign n_44628 = ~n_38828 &  n_44627;
assign n_44629 = ~n_38824 &  n_44628;
assign n_44630 = ~n_38820 &  n_44629;
assign n_44631 = ~n_38816 &  n_44630;
assign n_44632 = ~n_38812 &  n_44631;
assign n_44633 = ~n_38808 &  n_44632;
assign n_44634 = ~n_38804 &  n_44633;
assign n_44635 = ~n_38800 &  n_44634;
assign n_44636 = ~n_38796 &  n_44635;
assign n_44637 = ~n_38792 &  n_44636;
assign n_44638 = ~n_38786 &  n_44637;
assign n_44639 = ~n_38780 &  n_44638;
assign n_44640 = ~n_38774 &  n_44639;
assign n_44641 = ~n_38768 &  n_44640;
assign n_44642 = ~n_38762 &  n_44641;
assign n_44643 = ~n_38756 &  n_44642;
assign n_44644 = ~n_38750 &  n_44643;
assign n_44645 = ~n_38744 &  n_44644;
assign n_44646 = ~n_38738 &  n_44645;
assign n_44647 = ~n_38732 &  n_44646;
assign n_44648 = ~n_38726 &  n_44647;
assign n_44649 = ~n_38720 &  n_44648;
assign n_44650 = ~n_38714 &  n_44649;
assign n_44651 = ~n_38708 &  n_44650;
assign n_44652 = ~n_38702 &  n_44651;
assign n_44653 = ~n_38696 &  n_44652;
assign n_44654 = ~n_38690 &  n_44653;
assign n_44655 = ~n_38684 &  n_44654;
assign n_44656 = ~n_38678 &  n_44655;
assign n_44657 = ~n_38672 &  n_44656;
assign n_44658 = ~n_38666 &  n_44657;
assign n_44659 = ~n_38660 &  n_44658;
assign n_44660 = ~n_38654 &  n_44659;
assign n_44661 = ~n_38648 &  n_44660;
assign n_44662 = ~n_38642 &  n_44661;
assign n_44663 = ~n_38636 &  n_44662;
assign n_44664 = ~n_38630 &  n_44663;
assign n_44665 = ~n_38624 &  n_44664;
assign n_44666 = ~n_38618 &  n_44665;
assign n_44667 = ~n_38612 &  n_44666;
assign n_44668 = ~n_38606 &  n_44667;
assign n_44669 = ~n_38600 &  n_44668;
assign n_44670 = ~n_38594 &  n_44669;
assign n_44671 = ~n_38588 &  n_44670;
assign n_44672 = ~n_38582 &  n_44671;
assign n_44673 = ~n_38576 &  n_44672;
assign n_44674 = ~n_38570 &  n_44673;
assign n_44675 = ~n_38564 &  n_44674;
assign n_44676 = ~n_38558 &  n_44675;
assign n_44677 = ~n_38552 &  n_44676;
assign n_44678 = ~n_38546 &  n_44677;
assign n_44679 = ~n_38540 &  n_44678;
assign n_44680 = ~n_38534 &  n_44679;
assign n_44681 = ~n_38528 &  n_44680;
assign n_44682 = ~n_38522 &  n_44681;
assign n_44683 = ~n_38516 &  n_44682;
assign n_44684 = ~n_38510 &  n_44683;
assign n_44685 = ~n_38504 &  n_44684;
assign n_44686 = ~n_38498 &  n_44685;
assign n_44687 = ~n_38492 &  n_44686;
assign n_44688 = ~n_38486 &  n_44687;
assign n_44689 = ~n_38480 &  n_44688;
assign n_44690 = ~n_38474 &  n_44689;
assign n_44691 = ~n_38468 &  n_44690;
assign n_44692 = ~n_38462 &  n_44691;
assign n_44693 = ~n_38456 &  n_44692;
assign n_44694 = ~n_38450 &  n_44693;
assign n_44695 = ~n_38444 &  n_44694;
assign n_44696 = ~n_38438 &  n_44695;
assign n_44697 = ~n_38432 &  n_44696;
assign n_44698 = ~n_38426 &  n_44697;
assign n_44699 = ~n_38420 &  n_44698;
assign n_44700 = ~n_38414 &  n_44699;
assign n_44701 = ~n_38410 &  n_44700;
assign n_44702 = ~n_38406 &  n_44701;
assign n_44703 = ~n_38402 &  n_44702;
assign n_44704 = ~n_38398 &  n_44703;
assign n_44705 = ~n_38394 &  n_44704;
assign n_44706 = ~n_38390 &  n_44705;
assign n_44707 = ~n_38386 &  n_44706;
assign n_44708 = ~n_38382 &  n_44707;
assign n_44709 = ~n_38378 &  n_44708;
assign n_44710 = ~n_38374 &  n_44709;
assign n_44711 = ~n_38370 &  n_44710;
assign n_44712 = ~n_38366 &  n_44711;
assign n_44713 = ~n_38362 &  n_44712;
assign n_44714 = ~n_38358 &  n_44713;
assign n_44715 = ~n_38354 &  n_44714;
assign n_44716 = ~n_38350 &  n_44715;
assign n_44717 = ~n_38346 &  n_44716;
assign n_44718 = ~n_38342 &  n_44717;
assign n_44719 = ~n_38338 &  n_44718;
assign n_44720 = ~n_38334 &  n_44719;
assign n_44721 = ~n_38330 &  n_44720;
assign n_44722 = ~n_38326 &  n_44721;
assign n_44723 = ~n_38322 &  n_44722;
assign n_44724 = ~n_38318 &  n_44723;
assign n_44725 = ~n_38314 &  n_44724;
assign n_44726 = ~n_38310 &  n_44725;
assign n_44727 = ~n_38306 &  n_44726;
assign n_44728 = ~n_38302 &  n_44727;
assign n_44729 = ~n_38298 &  n_44728;
assign n_44730 = ~n_38294 &  n_44729;
assign n_44731 = ~n_38289 &  n_44730;
assign n_44732 = ~n_38281 &  n_44731;
assign n_44733 = ~n_38275 &  n_44732;
assign n_44734 = ~n_38269 &  n_44733;
assign n_44735 = ~n_38263 &  n_44734;
assign n_44736 = ~n_38257 &  n_44735;
assign n_44737 = ~n_38251 &  n_44736;
assign n_44738 = ~n_38245 &  n_44737;
assign n_44739 = ~n_38239 &  n_44738;
assign n_44740 = ~n_38233 &  n_44739;
assign n_44741 = ~n_38227 &  n_44740;
assign n_44742 = ~n_38221 &  n_44741;
assign n_44743 = ~n_38215 &  n_44742;
assign n_44744 = ~n_38209 &  n_44743;
assign n_44745 = ~n_38203 &  n_44744;
assign n_44746 = ~n_38197 &  n_44745;
assign n_44747 = ~n_38191 &  n_44746;
assign n_44748 = ~n_38185 &  n_44747;
assign n_44749 = ~n_38179 &  n_44748;
assign n_44750 = ~n_38173 &  n_44749;
assign n_44751 = ~n_38167 &  n_44750;
assign n_44752 = ~n_38161 &  n_44751;
assign n_44753 = ~n_38155 &  n_44752;
assign n_44754 = ~n_38149 &  n_44753;
assign n_44755 = ~n_38143 &  n_44754;
assign n_44756 = ~n_38137 &  n_44755;
assign n_44757 = ~n_38131 &  n_44756;
assign n_44758 = ~n_38125 &  n_44757;
assign n_44759 = ~n_38119 &  n_44758;
assign n_44760 = ~n_38113 &  n_44759;
assign n_44761 = ~n_38107 &  n_44760;
assign n_44762 = ~n_38101 &  n_44761;
assign n_44763 = ~n_38095 &  n_44762;
assign n_44764 = ~n_38089 &  n_44763;
assign n_44765 = ~n_38083 &  n_44764;
assign n_44766 = ~n_38077 &  n_44765;
assign n_44767 = ~n_38071 &  n_44766;
assign n_44768 = ~n_38065 &  n_44767;
assign n_44769 = ~n_38059 &  n_44768;
assign n_44770 = ~n_38053 &  n_44769;
assign n_44771 = ~n_38047 &  n_44770;
assign n_44772 = ~n_38041 &  n_44771;
assign n_44773 = ~n_38035 &  n_44772;
assign n_44774 = ~n_38029 &  n_44773;
assign n_44775 = ~n_38023 &  n_44774;
assign n_44776 = ~n_38017 &  n_44775;
assign n_44777 = ~n_38011 &  n_44776;
assign n_44778 = ~n_38005 &  n_44777;
assign n_44779 = ~n_37999 &  n_44778;
assign n_44780 = ~n_37993 &  n_44779;
assign n_44781 = ~n_37987 &  n_44780;
assign n_44782 = ~n_37981 &  n_44781;
assign n_44783 = ~n_37975 &  n_44782;
assign n_44784 = ~n_37969 &  n_44783;
assign n_44785 = ~n_37963 &  n_44784;
assign n_44786 = ~n_37957 &  n_44785;
assign n_44787 = ~n_37951 &  n_44786;
assign n_44788 = ~n_37945 &  n_44787;
assign n_44789 = ~n_37939 &  n_44788;
assign n_44790 = ~n_37933 &  n_44789;
assign n_44791 = ~n_37927 &  n_44790;
assign n_44792 = ~n_37921 &  n_44791;
assign n_44793 = ~n_37915 &  n_44792;
assign n_44794 = ~n_37909 &  n_44793;
assign n_44795 = ~n_37903 &  n_44794;
assign n_44796 = ~n_37897 &  n_44795;
assign n_44797 = ~n_37891 &  n_44796;
assign n_44798 = ~n_37885 &  n_44797;
assign n_44799 = ~n_37879 &  n_44798;
assign n_44800 = ~n_37873 &  n_44799;
assign n_44801 = ~n_37867 &  n_44800;
assign n_44802 = ~n_37861 &  n_44801;
assign n_44803 = ~n_37855 &  n_44802;
assign n_44804 = ~n_37849 &  n_44803;
assign n_44805 = ~n_37843 &  n_44804;
assign n_44806 = ~n_37837 &  n_44805;
assign n_44807 = ~n_37831 &  n_44806;
assign n_44808 = ~n_37825 &  n_44807;
assign n_44809 = ~n_37819 &  n_44808;
assign n_44810 = ~n_37813 &  n_44809;
assign n_44811 = ~n_37807 &  n_44810;
assign n_44812 = ~n_37801 &  n_44811;
assign n_44813 = ~n_37795 &  n_44812;
assign n_44814 = ~n_37789 &  n_44813;
assign n_44815 = ~n_37783 &  n_44814;
assign n_44816 = ~n_37777 &  n_44815;
assign n_44817 = ~n_37771 &  n_44816;
assign n_44818 = ~n_37765 &  n_44817;
assign n_44819 = ~n_37759 &  n_44818;
assign n_44820 = ~n_37753 &  n_44819;
assign n_44821 = ~n_37747 &  n_44820;
assign n_44822 = ~n_37741 &  n_44821;
assign n_44823 = ~n_37735 &  n_44822;
assign n_44824 = ~n_37729 &  n_44823;
assign n_44825 = ~n_37723 &  n_44824;
assign n_44826 = ~n_37717 &  n_44825;
assign n_44827 = ~n_37711 &  n_44826;
assign n_44828 = ~n_37705 &  n_44827;
assign n_44829 = ~n_37699 &  n_44828;
assign n_44830 = ~n_37693 &  n_44829;
assign n_44831 = ~n_37687 &  n_44830;
assign n_44832 = ~n_37681 &  n_44831;
assign n_44833 = ~n_37675 &  n_44832;
assign n_44834 = ~n_37669 &  n_44833;
assign n_44835 = ~n_37663 &  n_44834;
assign n_44836 = ~n_37657 &  n_44835;
assign n_44837 = ~n_37651 &  n_44836;
assign n_44838 = ~n_37645 &  n_44837;
assign n_44839 = ~n_37639 &  n_44838;
assign n_44840 = ~n_37633 &  n_44839;
assign n_44841 = ~n_37627 &  n_44840;
assign n_44842 = ~n_37621 &  n_44841;
assign n_44843 = ~n_37615 &  n_44842;
assign n_44844 = ~n_37609 &  n_44843;
assign n_44845 = ~n_37603 &  n_44844;
assign n_44846 = ~n_37597 &  n_44845;
assign n_44847 = ~n_37591 &  n_44846;
assign n_44848 = ~n_37585 &  n_44847;
assign n_44849 = ~n_37579 &  n_44848;
assign n_44850 = ~n_37573 &  n_44849;
assign n_44851 = ~n_37567 &  n_44850;
assign n_44852 = ~n_37561 &  n_44851;
assign n_44853 = ~n_37555 &  n_44852;
assign n_44854 = ~n_37549 &  n_44853;
assign n_44855 = ~n_37543 &  n_44854;
assign n_44856 = ~n_37537 &  n_44855;
assign n_44857 = ~n_37531 &  n_44856;
assign n_44858 = ~n_37525 &  n_44857;
assign n_44859 = ~n_37519 &  n_44858;
assign n_44860 = ~n_37513 &  n_44859;
assign n_44861 = ~n_37507 &  n_44860;
assign n_44862 = ~n_37499 &  n_44861;
assign n_44863 = ~n_37491 &  n_44862;
assign n_44864 = ~n_37483 &  n_44863;
assign n_44865 = ~n_37475 &  n_44864;
assign n_44866 = ~n_37467 &  n_44865;
assign n_44867 = ~n_37459 &  n_44866;
assign n_44868 = ~n_37451 &  n_44867;
assign n_44869 = ~n_37443 &  n_44868;
assign n_44870 = ~n_37435 &  n_44869;
assign n_44871 = ~n_37427 &  n_44870;
assign n_44872 = ~n_37419 &  n_44871;
assign n_44873 = ~n_37411 &  n_44872;
assign n_44874 = ~n_37403 &  n_44873;
assign n_44875 = ~n_37395 &  n_44874;
assign n_44876 = ~n_37387 &  n_44875;
assign n_44877 = ~n_37379 &  n_44876;
assign n_44878 = ~n_37371 &  n_44877;
assign n_44879 = ~n_37363 &  n_44878;
assign n_44880 = ~n_37355 &  n_44879;
assign n_44881 = ~n_37347 &  n_44880;
assign n_44882 = ~n_37339 &  n_44881;
assign n_44883 = ~n_37331 &  n_44882;
assign n_44884 = ~n_37323 &  n_44883;
assign n_44885 = ~n_37315 &  n_44884;
assign n_44886 = ~n_37307 &  n_44885;
assign n_44887 = ~n_37299 &  n_44886;
assign n_44888 = ~n_37291 &  n_44887;
assign n_44889 = ~n_37283 &  n_44888;
assign n_44890 = ~n_37275 &  n_44889;
assign n_44891 = ~n_37267 &  n_44890;
assign n_44892 = ~n_37258 &  n_44891;
assign n_44893 = ~n_37252 &  n_44892;
assign n_44894 = ~n_37246 &  n_44893;
assign n_44895 = ~n_37240 &  n_44894;
assign n_44896 = ~n_37234 &  n_44895;
assign n_44897 = ~n_37228 &  n_44896;
assign n_44898 = ~n_37222 &  n_44897;
assign n_44899 = ~n_37216 &  n_44898;
assign n_44900 = ~n_37210 &  n_44899;
assign n_44901 = ~n_37204 &  n_44900;
assign n_44902 = ~n_37198 &  n_44901;
assign n_44903 = ~n_37192 &  n_44902;
assign n_44904 = ~n_37186 &  n_44903;
assign n_44905 = ~n_37180 &  n_44904;
assign n_44906 = ~n_37174 &  n_44905;
assign n_44907 = ~n_37168 &  n_44906;
assign n_44908 = ~n_37162 &  n_44907;
assign n_44909 = ~n_37156 &  n_44908;
assign n_44910 = ~n_37150 &  n_44909;
assign n_44911 = ~n_37144 &  n_44910;
assign n_44912 = ~n_37138 &  n_44911;
assign n_44913 = ~n_37132 &  n_44912;
assign n_44914 = ~n_37126 &  n_44913;
assign n_44915 = ~n_37120 &  n_44914;
assign n_44916 = ~n_37114 &  n_44915;
assign n_44917 = ~n_37108 &  n_44916;
assign n_44918 = ~n_37102 &  n_44917;
assign n_44919 = ~n_37096 &  n_44918;
assign n_44920 = ~n_37090 &  n_44919;
assign n_44921 = ~n_37084 &  n_44920;
assign n_44922 = ~n_37078 &  n_44921;
assign n_44923 = ~n_37072 &  n_44922;
assign n_44924 = ~n_37066 &  n_44923;
assign n_44925 = ~n_37051 &  n_44924;
assign n_44926 = ~n_37036 &  n_44925;
assign n_44927 = ~n_37021 &  n_44926;
assign n_44928 = ~n_37006 &  n_44927;
assign n_44929 = ~n_36991 &  n_44928;
assign n_44930 = ~n_36976 &  n_44929;
assign n_44931 = ~n_36961 &  n_44930;
assign n_44932 = ~n_36946 &  n_44931;
assign n_44933 = ~n_36931 &  n_44932;
assign n_44934 = ~n_36916 &  n_44933;
assign n_44935 = ~n_36901 &  n_44934;
assign n_44936 = ~n_36886 &  n_44935;
assign n_44937 = ~n_36871 &  n_44936;
assign n_44938 = ~n_36856 &  n_44937;
assign n_44939 = ~n_36841 &  n_44938;
assign n_44940 = ~n_36826 &  n_44939;
assign n_44941 = ~n_36811 &  n_44940;
assign n_44942 = ~n_36796 &  n_44941;
assign n_44943 = ~n_36781 &  n_44942;
assign n_44944 = ~n_36766 &  n_44943;
assign n_44945 = ~n_36751 &  n_44944;
assign n_44946 = ~n_36736 &  n_44945;
assign n_44947 = ~n_36721 &  n_44946;
assign n_44948 = ~n_36706 &  n_44947;
assign n_44949 = ~n_36691 &  n_44948;
assign n_44950 = ~n_36676 &  n_44949;
assign n_44951 = ~n_36661 &  n_44950;
assign n_44952 = ~n_36646 &  n_44951;
assign n_44953 = ~n_36631 &  n_44952;
assign n_44954 = ~n_36616 &  n_44953;
assign n_44955 = ~n_36601 &  n_44954;
assign n_44956 = ~n_36586 &  n_44955;
assign n_44957 = ~n_36580 &  n_44956;
assign n_44958 = ~n_36574 &  n_44957;
assign n_44959 = ~n_36568 &  n_44958;
assign n_44960 = ~n_36562 &  n_44959;
assign n_44961 = ~n_36556 &  n_44960;
assign n_44962 = ~n_36550 &  n_44961;
assign n_44963 = ~n_36544 &  n_44962;
assign n_44964 = ~n_36538 &  n_44963;
assign n_44965 = ~n_36532 &  n_44964;
assign n_44966 = ~n_36526 &  n_44965;
assign n_44967 = ~n_36520 &  n_44966;
assign n_44968 = ~n_36514 &  n_44967;
assign n_44969 = ~n_36508 &  n_44968;
assign n_44970 = ~n_36502 &  n_44969;
assign n_44971 = ~n_36496 &  n_44970;
assign n_44972 = ~n_36490 &  n_44971;
assign n_44973 = ~n_36484 &  n_44972;
assign n_44974 = ~n_36478 &  n_44973;
assign n_44975 = ~n_36472 &  n_44974;
assign n_44976 = ~n_36466 &  n_44975;
assign n_44977 = ~n_36460 &  n_44976;
assign n_44978 = ~n_36454 &  n_44977;
assign n_44979 = ~n_36448 &  n_44978;
assign n_44980 = ~n_36442 &  n_44979;
assign n_44981 = ~n_36436 &  n_44980;
assign n_44982 = ~n_36430 &  n_44981;
assign n_44983 = ~n_36424 &  n_44982;
assign n_44984 = ~n_36418 &  n_44983;
assign n_44985 = ~n_36412 &  n_44984;
assign n_44986 = ~n_36406 &  n_44985;
assign n_44987 = ~n_36400 &  n_44986;
assign n_44988 = ~n_36394 &  n_44987;
assign n_44989 = ~n_36388 &  n_44988;
assign n_44990 = ~n_36382 &  n_44989;
assign n_44991 = ~n_36376 &  n_44990;
assign n_44992 = ~n_36370 &  n_44991;
assign n_44993 = ~n_36364 &  n_44992;
assign n_44994 = ~n_36358 &  n_44993;
assign n_44995 = ~n_36352 &  n_44994;
assign n_44996 = ~n_36346 &  n_44995;
assign n_44997 = ~n_36340 &  n_44996;
assign n_44998 = ~n_36334 &  n_44997;
assign n_44999 = ~n_36328 &  n_44998;
assign n_45000 = ~n_36322 &  n_44999;
assign n_45001 = ~n_36316 &  n_45000;
assign n_45002 = ~n_36310 &  n_45001;
assign n_45003 = ~n_36304 &  n_45002;
assign n_45004 = ~n_36298 &  n_45003;
assign n_45005 = ~n_36292 &  n_45004;
assign n_45006 = ~n_36286 &  n_45005;
assign n_45007 = ~n_36280 &  n_45006;
assign n_45008 = ~n_36274 &  n_45007;
assign n_45009 = ~n_36268 &  n_45008;
assign n_45010 = ~n_36262 &  n_45009;
assign n_45011 = ~n_36256 &  n_45010;
assign n_45012 = ~n_36250 &  n_45011;
assign n_45013 = ~n_36244 &  n_45012;
assign n_45014 = ~n_36238 &  n_45013;
assign n_45015 = ~n_36232 &  n_45014;
assign n_45016 = ~n_36226 &  n_45015;
assign n_45017 = ~n_36220 &  n_45016;
assign n_45018 = ~n_36214 &  n_45017;
assign n_45019 = ~n_36208 &  n_45018;
assign n_45020 = ~n_36201 &  n_45019;
assign n_45021 = ~n_36195 &  n_45020;
assign n_45022 = ~n_36189 &  n_45021;
assign n_45023 = ~n_36183 &  n_45022;
assign n_45024 = ~n_36177 &  n_45023;
assign n_45025 = ~n_36171 &  n_45024;
assign n_45026 = ~n_36165 &  n_45025;
assign n_45027 = ~n_36159 &  n_45026;
assign n_45028 = ~n_36153 &  n_45027;
assign n_45029 = ~n_36147 &  n_45028;
assign n_45030 = ~n_36141 &  n_45029;
assign n_45031 = ~n_36135 &  n_45030;
assign n_45032 = ~n_36129 &  n_45031;
assign n_45033 = ~n_36123 &  n_45032;
assign n_45034 = ~n_36117 &  n_45033;
assign n_45035 = ~n_36111 &  n_45034;
assign n_45036 = ~n_36105 &  n_45035;
assign n_45037 = ~n_36099 &  n_45036;
assign n_45038 = ~n_36093 &  n_45037;
assign n_45039 = ~n_36087 &  n_45038;
assign n_45040 = ~n_36081 &  n_45039;
assign n_45041 = ~n_36075 &  n_45040;
assign n_45042 = ~n_36069 &  n_45041;
assign n_45043 = ~n_36063 &  n_45042;
assign n_45044 = ~n_36057 &  n_45043;
assign n_45045 = ~n_36051 &  n_45044;
assign n_45046 = ~n_36045 &  n_45045;
assign n_45047 = ~n_36039 &  n_45046;
assign n_45048 = ~n_36033 &  n_45047;
assign n_45049 = ~n_36027 &  n_45048;
assign n_45050 = ~n_36021 &  n_45049;
assign n_45051 = ~n_36015 &  n_45050;
assign n_45052 = ~n_36007 &  n_45051;
assign n_45053 = ~n_36003 &  n_45052;
assign n_45054 = ~n_35997 &  n_45053;
assign n_45055 = ~n_35991 &  n_45054;
assign n_45056 = ~n_35985 &  n_45055;
assign n_45057 = ~n_35979 &  n_45056;
assign n_45058 = ~n_35973 &  n_45057;
assign n_45059 = ~n_35967 &  n_45058;
assign n_45060 = ~n_35961 &  n_45059;
assign n_45061 = ~n_35955 &  n_45060;
assign n_45062 = ~n_35949 &  n_45061;
assign n_45063 = ~n_35943 &  n_45062;
assign n_45064 = ~n_35937 &  n_45063;
assign n_45065 = ~n_35931 &  n_45064;
assign n_45066 = ~n_35925 &  n_45065;
assign n_45067 = ~n_35919 &  n_45066;
assign n_45068 = ~n_35913 &  n_45067;
assign n_45069 = ~n_35907 &  n_45068;
assign n_45070 = ~n_35901 &  n_45069;
assign n_45071 = ~n_35895 &  n_45070;
assign n_45072 = ~n_35889 &  n_45071;
assign n_45073 = ~n_35883 &  n_45072;
assign n_45074 = ~n_35877 &  n_45073;
assign n_45075 = ~n_35871 &  n_45074;
assign n_45076 = ~n_35865 &  n_45075;
assign n_45077 = ~n_35859 &  n_45076;
assign n_45078 = ~n_35853 &  n_45077;
assign n_45079 = ~n_35847 &  n_45078;
assign n_45080 = ~n_35841 &  n_45079;
assign n_45081 = ~n_35835 &  n_45080;
assign n_45082 = ~n_35829 &  n_45081;
assign n_45083 = ~n_35823 &  n_45082;
assign n_45084 = ~n_35817 &  n_45083;
assign n_45085 = ~n_35813 &  n_45084;
assign n_45086 = ~n_35809 &  n_45085;
assign n_45087 = ~n_35805 &  n_45086;
assign n_45088 = ~n_35801 &  n_45087;
assign n_45089 = ~n_35797 &  n_45088;
assign n_45090 = ~n_35793 &  n_45089;
assign n_45091 = ~n_35789 &  n_45090;
assign n_45092 = ~n_35785 &  n_45091;
assign n_45093 = ~n_35781 &  n_45092;
assign n_45094 = ~n_35777 &  n_45093;
assign n_45095 = ~n_35773 &  n_45094;
assign n_45096 = ~n_35769 &  n_45095;
assign n_45097 = ~n_35765 &  n_45096;
assign n_45098 = ~n_35761 &  n_45097;
assign n_45099 = ~n_35757 &  n_45098;
assign n_45100 = ~n_35753 &  n_45099;
assign n_45101 = ~n_35749 &  n_45100;
assign n_45102 = ~n_35745 &  n_45101;
assign n_45103 = ~n_35741 &  n_45102;
assign n_45104 = ~n_35737 &  n_45103;
assign n_45105 = ~n_35733 &  n_45104;
assign n_45106 = ~n_35729 &  n_45105;
assign n_45107 = ~n_35725 &  n_45106;
assign n_45108 = ~n_35721 &  n_45107;
assign n_45109 = ~n_35717 &  n_45108;
assign n_45110 = ~n_35713 &  n_45109;
assign n_45111 = ~n_35709 &  n_45110;
assign n_45112 = ~n_35705 &  n_45111;
assign n_45113 = ~n_35701 &  n_45112;
assign n_45114 = ~n_35697 &  n_45113;
assign n_45115 = ~n_35693 &  n_45114;
assign n_45116 = ~n_35689 &  n_45115;
assign n_45117 = ~n_35685 &  n_45116;
assign n_45118 = ~n_35681 &  n_45117;
assign n_45119 = ~n_35677 &  n_45118;
assign n_45120 = ~n_35673 &  n_45119;
assign n_45121 = ~n_35669 &  n_45120;
assign n_45122 = ~n_35665 &  n_45121;
assign n_45123 = ~n_35661 &  n_45122;
assign n_45124 = ~n_35657 &  n_45123;
assign n_45125 = ~n_35653 &  n_45124;
assign n_45126 = ~n_35649 &  n_45125;
assign n_45127 = ~n_35645 &  n_45126;
assign n_45128 = ~n_35641 &  n_45127;
assign n_45129 = ~n_35637 &  n_45128;
assign n_45130 = ~n_35633 &  n_45129;
assign n_45131 = ~n_35629 &  n_45130;
assign n_45132 = ~n_35625 &  n_45131;
assign n_45133 = ~n_35621 &  n_45132;
assign n_45134 = ~n_35617 &  n_45133;
assign n_45135 = ~n_35613 &  n_45134;
assign n_45136 = ~n_35609 &  n_45135;
assign n_45137 = ~n_35605 &  n_45136;
assign n_45138 = ~n_35601 &  n_45137;
assign n_45139 = ~n_35597 &  n_45138;
assign n_45140 = ~n_35593 &  n_45139;
assign n_45141 = ~n_35589 &  n_45140;
assign n_45142 = ~n_35585 &  n_45141;
assign n_45143 = ~n_35581 &  n_45142;
assign n_45144 = ~n_35577 &  n_45143;
assign n_45145 = ~n_35573 &  n_45144;
assign n_45146 = ~n_35569 &  n_45145;
assign n_45147 = ~n_35564 &  n_45146;
assign n_45148 = ~n_35558 &  n_45147;
assign n_45149 = ~n_35552 &  n_45148;
assign n_45150 = ~n_35546 &  n_45149;
assign n_45151 = ~n_35540 &  n_45150;
assign n_45152 = ~n_35534 &  n_45151;
assign n_45153 = ~n_35528 &  n_45152;
assign n_45154 = ~n_35522 &  n_45153;
assign n_45155 = ~n_35516 &  n_45154;
assign n_45156 = ~n_35510 &  n_45155;
assign n_45157 = ~n_35504 &  n_45156;
assign n_45158 = ~n_35498 &  n_45157;
assign n_45159 = ~n_35492 &  n_45158;
assign n_45160 = ~n_35486 &  n_45159;
assign n_45161 = ~n_35480 &  n_45160;
assign n_45162 = ~n_35474 &  n_45161;
assign n_45163 = ~n_35468 &  n_45162;
assign n_45164 = ~n_35462 &  n_45163;
assign n_45165 = ~n_35456 &  n_45164;
assign n_45166 = ~n_35450 &  n_45165;
assign n_45167 = ~n_35444 &  n_45166;
assign n_45168 = ~n_35438 &  n_45167;
assign n_45169 = ~n_35432 &  n_45168;
assign n_45170 = ~n_35426 &  n_45169;
assign n_45171 = ~n_35420 &  n_45170;
assign n_45172 = ~n_35414 &  n_45171;
assign n_45173 = ~n_35408 &  n_45172;
assign n_45174 = ~n_35402 &  n_45173;
assign n_45175 = ~n_35396 &  n_45174;
assign n_45176 = ~n_35390 &  n_45175;
assign n_45177 = ~n_35384 &  n_45176;
assign n_45178 = ~n_35378 &  n_45177;
assign n_45179 = ~n_35372 &  n_45178;
assign n_45180 = ~n_35366 &  n_45179;
assign n_45181 = ~n_35360 &  n_45180;
assign n_45182 = ~n_35354 &  n_45181;
assign n_45183 = ~n_35348 &  n_45182;
assign n_45184 = ~n_35342 &  n_45183;
assign n_45185 = ~n_35336 &  n_45184;
assign n_45186 = ~n_35330 &  n_45185;
assign n_45187 = ~n_35324 &  n_45186;
assign n_45188 = ~n_35318 &  n_45187;
assign n_45189 = ~n_35312 &  n_45188;
assign n_45190 = ~n_35306 &  n_45189;
assign n_45191 = ~n_35300 &  n_45190;
assign n_45192 = ~n_35294 &  n_45191;
assign n_45193 = ~n_35288 &  n_45192;
assign n_45194 = ~n_35282 &  n_45193;
assign n_45195 = ~n_35276 &  n_45194;
assign n_45196 = ~n_35270 &  n_45195;
assign n_45197 = ~n_35264 &  n_45196;
assign n_45198 = ~n_35258 &  n_45197;
assign n_45199 = ~n_35252 &  n_45198;
assign n_45200 = ~n_35246 &  n_45199;
assign n_45201 = ~n_35240 &  n_45200;
assign n_45202 = ~n_35234 &  n_45201;
assign n_45203 = ~n_35228 &  n_45202;
assign n_45204 = ~n_35222 &  n_45203;
assign n_45205 = ~n_35216 &  n_45204;
assign n_45206 = ~n_35210 &  n_45205;
assign n_45207 = ~n_35204 &  n_45206;
assign n_45208 = ~n_35198 &  n_45207;
assign n_45209 = ~n_35192 &  n_45208;
assign n_45210 = ~n_35186 &  n_45209;
assign n_45211 = ~n_35180 &  n_45210;
assign n_45212 = ~n_35174 &  n_45211;
assign n_45213 = ~n_35168 &  n_45212;
assign n_45214 = ~n_35162 &  n_45213;
assign n_45215 = ~n_35156 &  n_45214;
assign n_45216 = ~n_35150 &  n_45215;
assign n_45217 = ~n_35144 &  n_45216;
assign n_45218 = ~n_35138 &  n_45217;
assign n_45219 = ~n_35132 &  n_45218;
assign n_45220 = ~n_35126 &  n_45219;
assign n_45221 = ~n_35120 &  n_45220;
assign n_45222 = ~n_35114 &  n_45221;
assign n_45223 = ~n_35108 &  n_45222;
assign n_45224 = ~n_35102 &  n_45223;
assign n_45225 = ~n_35096 &  n_45224;
assign n_45226 = ~n_35090 &  n_45225;
assign n_45227 = ~n_35084 &  n_45226;
assign n_45228 = ~n_35078 &  n_45227;
assign n_45229 = ~n_35072 &  n_45228;
assign n_45230 = ~n_35066 &  n_45229;
assign n_45231 = ~n_35060 &  n_45230;
assign n_45232 = ~n_35054 &  n_45231;
assign n_45233 = ~n_35048 &  n_45232;
assign n_45234 = ~n_35042 &  n_45233;
assign n_45235 = ~n_35036 &  n_45234;
assign n_45236 = ~n_35030 &  n_45235;
assign n_45237 = ~n_35024 &  n_45236;
assign n_45238 = ~n_35018 &  n_45237;
assign n_45239 = ~n_35012 &  n_45238;
assign n_45240 = ~n_35006 &  n_45239;
assign n_45241 = ~n_35000 &  n_45240;
assign n_45242 = ~n_34994 &  n_45241;
assign n_45243 = ~n_34988 &  n_45242;
assign n_45244 = ~n_34982 &  n_45243;
assign n_45245 = ~n_34976 &  n_45244;
assign n_45246 = ~n_34970 &  n_45245;
assign n_45247 = ~n_34964 &  n_45246;
assign n_45248 = ~n_34958 &  n_45247;
assign n_45249 = ~n_34952 &  n_45248;
assign n_45250 = ~n_34946 &  n_45249;
assign n_45251 = ~n_34940 &  n_45250;
assign n_45252 = ~n_34934 &  n_45251;
assign n_45253 = ~n_34928 &  n_45252;
assign n_45254 = ~n_34922 &  n_45253;
assign n_45255 = ~n_34916 &  n_45254;
assign n_45256 = ~n_34910 &  n_45255;
assign n_45257 = ~n_34904 &  n_45256;
assign n_45258 = ~n_34898 &  n_45257;
assign n_45259 = ~n_34892 &  n_45258;
assign n_45260 = ~n_34886 &  n_45259;
assign n_45261 = ~n_34880 &  n_45260;
assign n_45262 = ~n_34874 &  n_45261;
assign n_45263 = ~n_34868 &  n_45262;
assign n_45264 = ~n_34862 &  n_45263;
assign n_45265 = ~n_34856 &  n_45264;
assign n_45266 = ~n_34850 &  n_45265;
assign n_45267 = ~n_34844 &  n_45266;
assign n_45268 = ~n_34838 &  n_45267;
assign n_45269 = ~n_34832 &  n_45268;
assign n_45270 = ~n_34826 &  n_45269;
assign n_45271 = ~n_34820 &  n_45270;
assign n_45272 = ~n_34814 &  n_45271;
assign n_45273 = ~n_34808 &  n_45272;
assign n_45274 = ~n_34802 &  n_45273;
assign n_45275 = ~n_34796 &  n_45274;
assign n_45276 = ~n_34790 &  n_45275;
assign n_45277 = ~n_34784 &  n_45276;
assign n_45278 = ~n_34778 &  n_45277;
assign n_45279 = ~n_34772 &  n_45278;
assign n_45280 = ~n_34766 &  n_45279;
assign n_45281 = ~n_34760 &  n_45280;
assign n_45282 = ~n_34754 &  n_45281;
assign n_45283 = ~n_34748 &  n_45282;
assign n_45284 = ~n_34742 &  n_45283;
assign n_45285 = ~n_34736 &  n_45284;
assign n_45286 = ~n_34730 &  n_45285;
assign n_45287 = ~n_34724 &  n_45286;
assign n_45288 = ~n_34718 &  n_45287;
assign n_45289 = ~n_34712 &  n_45288;
assign n_45290 = ~n_34706 &  n_45289;
assign n_45291 = ~n_34700 &  n_45290;
assign n_45292 = ~n_34694 &  n_45291;
assign n_45293 = ~n_34688 &  n_45292;
assign n_45294 = ~n_34682 &  n_45293;
assign n_45295 = ~n_34676 &  n_45294;
assign n_45296 = ~n_34670 &  n_45295;
assign n_45297 = ~n_34664 &  n_45296;
assign n_45298 = ~n_34658 &  n_45297;
assign n_45299 = ~n_34652 &  n_45298;
assign n_45300 = ~n_34646 &  n_45299;
assign n_45301 = ~n_34640 &  n_45300;
assign n_45302 = ~n_34634 &  n_45301;
assign n_45303 = ~n_34628 &  n_45302;
assign n_45304 = ~n_34622 &  n_45303;
assign n_45305 = ~n_34616 &  n_45304;
assign n_45306 = ~n_34610 &  n_45305;
assign n_45307 = ~n_34604 &  n_45306;
assign n_45308 = ~n_34597 &  n_45307;
assign n_45309 = ~n_34591 &  n_45308;
assign n_45310 = ~n_34585 &  n_45309;
assign n_45311 = ~n_34579 &  n_45310;
assign n_45312 = ~n_34573 &  n_45311;
assign n_45313 = ~n_34567 &  n_45312;
assign n_45314 = ~n_34561 &  n_45313;
assign n_45315 = ~n_34555 &  n_45314;
assign n_45316 = ~n_34549 &  n_45315;
assign n_45317 = ~n_34543 &  n_45316;
assign n_45318 = ~n_34537 &  n_45317;
assign n_45319 = ~n_34531 &  n_45318;
assign n_45320 = ~n_34525 &  n_45319;
assign n_45321 = ~n_34519 &  n_45320;
assign n_45322 = ~n_34513 &  n_45321;
assign n_45323 = ~n_34507 &  n_45322;
assign n_45324 = ~n_34501 &  n_45323;
assign n_45325 = ~n_34495 &  n_45324;
assign n_45326 = ~n_34489 &  n_45325;
assign n_45327 = ~n_34483 &  n_45326;
assign n_45328 = ~n_34477 &  n_45327;
assign n_45329 = ~n_34471 &  n_45328;
assign n_45330 = ~n_34465 &  n_45329;
assign n_45331 = ~n_34459 &  n_45330;
assign n_45332 = ~n_34453 &  n_45331;
assign n_45333 = ~n_34447 &  n_45332;
assign n_45334 = ~n_34441 &  n_45333;
assign n_45335 = ~n_34435 &  n_45334;
assign n_45336 = ~n_34429 &  n_45335;
assign n_45337 = ~n_34423 &  n_45336;
assign n_45338 = ~n_34417 &  n_45337;
assign n_45339 = ~n_34411 &  n_45338;
assign n_45340 = ~n_34405 &  n_45339;
assign n_45341 = ~n_34399 &  n_45340;
assign n_45342 = ~n_34393 &  n_45341;
assign n_45343 = ~n_34387 &  n_45342;
assign n_45344 = ~n_34381 &  n_45343;
assign n_45345 = ~n_34375 &  n_45344;
assign n_45346 = ~n_34369 &  n_45345;
assign n_45347 = ~n_34363 &  n_45346;
assign n_45348 = ~n_34357 &  n_45347;
assign n_45349 = ~n_34351 &  n_45348;
assign n_45350 = ~n_34345 &  n_45349;
assign n_45351 = ~n_34339 &  n_45350;
assign n_45352 = ~n_34333 &  n_45351;
assign n_45353 = ~n_34327 &  n_45352;
assign n_45354 = ~n_34321 &  n_45353;
assign n_45355 = ~n_34315 &  n_45354;
assign n_45356 = ~n_34309 &  n_45355;
assign n_45357 = ~n_34303 &  n_45356;
assign n_45358 = ~n_34297 &  n_45357;
assign n_45359 = ~n_34291 &  n_45358;
assign n_45360 = ~n_34285 &  n_45359;
assign n_45361 = ~n_34279 &  n_45360;
assign n_45362 = ~n_34273 &  n_45361;
assign n_45363 = ~n_34267 &  n_45362;
assign n_45364 = ~n_34261 &  n_45363;
assign n_45365 = ~n_34255 &  n_45364;
assign n_45366 = ~n_34249 &  n_45365;
assign n_45367 = ~n_34243 &  n_45366;
assign n_45368 = ~n_34237 &  n_45367;
assign n_45369 = ~n_34231 &  n_45368;
assign n_45370 = ~n_34225 &  n_45369;
assign n_45371 = ~n_34219 &  n_45370;
assign n_45372 = ~n_34213 &  n_45371;
assign n_45373 = ~n_34207 &  n_45372;
assign n_45374 = ~n_34201 &  n_45373;
assign n_45375 = ~n_34195 &  n_45374;
assign n_45376 = ~n_34189 &  n_45375;
assign n_45377 = ~n_34183 &  n_45376;
assign n_45378 = ~n_34177 &  n_45377;
assign n_45379 = ~n_34171 &  n_45378;
assign n_45380 = ~n_34165 &  n_45379;
assign n_45381 = ~n_34159 &  n_45380;
assign n_45382 = ~n_34153 &  n_45381;
assign n_45383 = ~n_34147 &  n_45382;
assign n_45384 = ~n_34141 &  n_45383;
assign n_45385 = ~n_34135 &  n_45384;
assign n_45386 = ~n_34129 &  n_45385;
assign n_45387 = ~n_34123 &  n_45386;
assign n_45388 = ~n_34117 &  n_45387;
assign n_45389 = ~n_34111 &  n_45388;
assign n_45390 = ~n_34105 &  n_45389;
assign n_45391 = ~n_34099 &  n_45390;
assign n_45392 = ~n_34093 &  n_45391;
assign n_45393 = ~n_34087 &  n_45392;
assign n_45394 = ~n_34081 &  n_45393;
assign n_45395 = ~n_34075 &  n_45394;
assign n_45396 = ~n_34069 &  n_45395;
assign n_45397 = ~n_34063 &  n_45396;
assign n_45398 = ~n_34057 &  n_45397;
assign n_45399 = ~n_34051 &  n_45398;
assign n_45400 = ~n_34045 &  n_45399;
assign n_45401 = ~n_34039 &  n_45400;
assign n_45402 = ~n_34033 &  n_45401;
assign n_45403 = ~n_34027 &  n_45402;
assign n_45404 = ~n_34021 &  n_45403;
assign n_45405 = ~n_34015 &  n_45404;
assign n_45406 = ~n_34009 &  n_45405;
assign n_45407 = ~n_34003 &  n_45406;
assign n_45408 = ~n_33997 &  n_45407;
assign n_45409 = ~n_33991 &  n_45408;
assign n_45410 = ~n_33985 &  n_45409;
assign n_45411 = ~n_33979 &  n_45410;
assign n_45412 = ~n_33973 &  n_45411;
assign n_45413 = ~n_33967 &  n_45412;
assign n_45414 = ~n_33961 &  n_45413;
assign n_45415 = ~n_33955 &  n_45414;
assign n_45416 = ~n_33949 &  n_45415;
assign n_45417 = ~n_33943 &  n_45416;
assign n_45418 = ~n_33937 &  n_45417;
assign n_45419 = ~n_33931 &  n_45418;
assign n_45420 = ~n_33925 &  n_45419;
assign n_45421 = ~n_33919 &  n_45420;
assign n_45422 = ~n_33913 &  n_45421;
assign n_45423 = ~n_33907 &  n_45422;
assign n_45424 = ~n_33901 &  n_45423;
assign n_45425 = ~n_33895 &  n_45424;
assign n_45426 = ~n_33889 &  n_45425;
assign n_45427 = ~n_33883 &  n_45426;
assign n_45428 = ~n_33877 &  n_45427;
assign n_45429 = ~n_33871 &  n_45428;
assign n_45430 = ~n_33865 &  n_45429;
assign n_45431 = ~n_33859 &  n_45430;
assign n_45432 = ~n_33853 &  n_45431;
assign n_45433 = ~n_33847 &  n_45432;
assign n_45434 = ~n_33841 &  n_45433;
assign n_45435 = ~n_33835 &  n_45434;
assign n_45436 = ~n_33829 &  n_45435;
assign n_45437 = ~n_33817 &  n_45436;
assign n_45438 = ~n_33805 &  n_45437;
assign n_45439 = ~n_33793 &  n_45438;
assign n_45440 = ~n_33781 &  n_45439;
assign n_45441 = ~n_33769 &  n_45440;
assign n_45442 = ~n_33757 &  n_45441;
assign n_45443 = ~n_33745 &  n_45442;
assign n_45444 = ~n_33733 &  n_45443;
assign n_45445 = ~n_33721 &  n_45444;
assign n_45446 = ~n_33709 &  n_45445;
assign n_45447 = ~n_33697 &  n_45446;
assign n_45448 = ~n_33685 &  n_45447;
assign n_45449 = ~n_33673 &  n_45448;
assign n_45450 = ~n_33661 &  n_45449;
assign n_45451 = ~n_33649 &  n_45450;
assign n_45452 = ~n_33637 &  n_45451;
assign n_45453 = ~n_33625 &  n_45452;
assign n_45454 = ~n_33613 &  n_45453;
assign n_45455 = ~n_33601 &  n_45454;
assign n_45456 = ~n_33589 &  n_45455;
assign n_45457 = ~n_33577 &  n_45456;
assign n_45458 = ~n_33565 &  n_45457;
assign n_45459 = ~n_33553 &  n_45458;
assign n_45460 = ~n_33541 &  n_45459;
assign n_45461 = ~n_33529 &  n_45460;
assign n_45462 = ~n_33517 &  n_45461;
assign n_45463 = ~n_33505 &  n_45462;
assign n_45464 = ~n_33493 &  n_45463;
assign n_45465 = ~n_33481 &  n_45464;
assign n_45466 = ~n_33469 &  n_45465;
assign n_45467 = ~n_33457 &  n_45466;
assign n_45468 = ~n_33442 &  n_45467;
assign n_45469 = ~n_33434 &  n_45468;
assign n_45470 = ~n_33426 &  n_45469;
assign n_45471 = ~n_33418 &  n_45470;
assign n_45472 = ~n_33410 &  n_45471;
assign n_45473 = ~n_33402 &  n_45472;
assign n_45474 = ~n_33394 &  n_45473;
assign n_45475 = ~n_33386 &  n_45474;
assign n_45476 = ~n_33378 &  n_45475;
assign n_45477 = ~n_33370 &  n_45476;
assign n_45478 = ~n_33362 &  n_45477;
assign n_45479 = ~n_33354 &  n_45478;
assign n_45480 = ~n_33346 &  n_45479;
assign n_45481 = ~n_33338 &  n_45480;
assign n_45482 = ~n_33330 &  n_45481;
assign n_45483 = ~n_33322 &  n_45482;
assign n_45484 = ~n_33314 &  n_45483;
assign n_45485 = ~n_33306 &  n_45484;
assign n_45486 = ~n_33298 &  n_45485;
assign n_45487 = ~n_33290 &  n_45486;
assign n_45488 = ~n_33282 &  n_45487;
assign n_45489 = ~n_33274 &  n_45488;
assign n_45490 = ~n_33266 &  n_45489;
assign n_45491 = ~n_33258 &  n_45490;
assign n_45492 = ~n_33250 &  n_45491;
assign n_45493 = ~n_33242 &  n_45492;
assign n_45494 = ~n_33234 &  n_45493;
assign n_45495 = ~n_33226 &  n_45494;
assign n_45496 = ~n_33218 &  n_45495;
assign n_45497 = ~n_33210 &  n_45496;
assign n_45498 = ~n_33202 &  n_45497;
assign n_45499 = ~n_33194 &  n_45498;
assign n_45500 = ~n_33184 &  n_45499;
assign n_45501 = ~n_33180 &  n_45500;
assign n_45502 = ~n_33176 &  n_45501;
assign n_45503 = ~n_33172 &  n_45502;
assign n_45504 = ~n_33168 &  n_45503;
assign n_45505 = ~n_33164 &  n_45504;
assign n_45506 = ~n_33160 &  n_45505;
assign n_45507 = ~n_33156 &  n_45506;
assign n_45508 = ~n_33152 &  n_45507;
assign n_45509 = ~n_33148 &  n_45508;
assign n_45510 = ~n_33144 &  n_45509;
assign n_45511 = ~n_33140 &  n_45510;
assign n_45512 = ~n_33136 &  n_45511;
assign n_45513 = ~n_33132 &  n_45512;
assign n_45514 = ~n_33128 &  n_45513;
assign n_45515 = ~n_33124 &  n_45514;
assign n_45516 = ~n_33120 &  n_45515;
assign n_45517 = ~n_33116 &  n_45516;
assign n_45518 = ~n_33112 &  n_45517;
assign n_45519 = ~n_33108 &  n_45518;
assign n_45520 = ~n_33104 &  n_45519;
assign n_45521 = ~n_33100 &  n_45520;
assign n_45522 = ~n_33096 &  n_45521;
assign n_45523 = ~n_33092 &  n_45522;
assign n_45524 = ~n_33088 &  n_45523;
assign n_45525 = ~n_33084 &  n_45524;
assign n_45526 = ~n_33080 &  n_45525;
assign n_45527 = ~n_33076 &  n_45526;
assign n_45528 = ~n_33072 &  n_45527;
assign n_45529 = ~n_33068 &  n_45528;
assign n_45530 = ~n_33064 &  n_45529;
assign n_45531 = ~n_33060 &  n_45530;
assign n_45532 = ~n_33056 &  n_45531;
assign n_45533 = ~n_33052 &  n_45532;
assign n_45534 = ~n_33048 &  n_45533;
assign n_45535 = ~n_33044 &  n_45534;
assign n_45536 = ~n_33040 &  n_45535;
assign n_45537 = ~n_33036 &  n_45536;
assign n_45538 = ~n_33032 &  n_45537;
assign n_45539 = ~n_33028 &  n_45538;
assign n_45540 = ~n_33024 &  n_45539;
assign n_45541 = ~n_33020 &  n_45540;
assign n_45542 = ~n_33016 &  n_45541;
assign n_45543 = ~n_33012 &  n_45542;
assign n_45544 = ~n_33008 &  n_45543;
assign n_45545 = ~n_33004 &  n_45544;
assign n_45546 = ~n_33000 &  n_45545;
assign n_45547 = ~n_32996 &  n_45546;
assign n_45548 = ~n_32992 &  n_45547;
assign n_45549 = ~n_32988 &  n_45548;
assign n_45550 = ~n_32984 &  n_45549;
assign n_45551 = ~n_32980 &  n_45550;
assign n_45552 = ~n_32976 &  n_45551;
assign n_45553 = ~n_32972 &  n_45552;
assign n_45554 = ~n_32968 &  n_45553;
assign n_45555 = ~n_32964 &  n_45554;
assign n_45556 = ~n_32960 &  n_45555;
assign n_45557 = ~n_32956 &  n_45556;
assign n_45558 = ~n_32952 &  n_45557;
assign n_45559 = ~n_32948 &  n_45558;
assign n_45560 = ~n_32944 &  n_45559;
assign n_45561 = ~n_32940 &  n_45560;
assign n_45562 = ~n_32936 &  n_45561;
assign n_45563 = ~n_32932 &  n_45562;
assign n_45564 = ~n_32928 &  n_45563;
assign n_45565 = ~n_32886 &  n_45564;
assign n_45566 = ~n_32841 &  n_45565;
assign n_45567 = ~n_32796 &  n_45566;
assign n_45568 = ~n_32751 &  n_45567;
assign n_45569 = ~n_32706 &  n_45568;
assign n_45570 = ~n_32661 &  n_45569;
assign n_45571 = ~n_32616 &  n_45570;
assign n_45572 = ~n_32571 &  n_45571;
assign n_45573 = ~n_32526 &  n_45572;
assign n_45574 = ~n_32481 &  n_45573;
assign n_45575 = ~n_32436 &  n_45574;
assign n_45576 = ~n_32391 &  n_45575;
assign n_45577 = ~n_32346 &  n_45576;
assign n_45578 = ~n_32301 &  n_45577;
assign n_45579 = ~n_32256 &  n_45578;
assign n_45580 = ~n_32211 &  n_45579;
assign n_45581 = ~n_32166 &  n_45580;
assign n_45582 = ~n_32121 &  n_45581;
assign n_45583 = ~n_32076 &  n_45582;
assign n_45584 = ~n_32031 &  n_45583;
assign n_45585 = ~n_31986 &  n_45584;
assign n_45586 = ~n_31941 &  n_45585;
assign n_45587 = ~n_31896 &  n_45586;
assign n_45588 = ~n_31851 &  n_45587;
assign n_45589 = ~n_31806 &  n_45588;
assign n_45590 = ~n_31761 &  n_45589;
assign n_45591 = ~n_31716 &  n_45590;
assign n_45592 = ~n_31671 &  n_45591;
assign n_45593 = ~n_31626 &  n_45592;
assign n_45594 = ~n_31575 &  n_45593;
assign n_45595 = ~n_31536 &  n_45594;
assign n_45596 = ~n_31512 &  n_45595;
assign n_45597 = ~n_31506 &  n_45596;
assign n_45598 = ~n_31500 &  n_45597;
assign n_45599 = ~n_31494 &  n_45598;
assign n_45600 = ~n_31488 &  n_45599;
assign n_45601 = ~n_31482 &  n_45600;
assign n_45602 = ~n_31476 &  n_45601;
assign n_45603 = ~n_31470 &  n_45602;
assign n_45604 = ~n_31464 &  n_45603;
assign n_45605 = ~n_31458 &  n_45604;
assign n_45606 = ~n_31452 &  n_45605;
assign n_45607 = ~n_31446 &  n_45606;
assign n_45608 = ~n_31440 &  n_45607;
assign n_45609 = ~n_31434 &  n_45608;
assign n_45610 = ~n_31428 &  n_45609;
assign n_45611 = ~n_31422 &  n_45610;
assign n_45612 = ~n_31416 &  n_45611;
assign n_45613 = ~n_31410 &  n_45612;
assign n_45614 = ~n_31404 &  n_45613;
assign n_45615 = ~n_31398 &  n_45614;
assign n_45616 = ~n_31392 &  n_45615;
assign n_45617 = ~n_31386 &  n_45616;
assign n_45618 = ~n_31380 &  n_45617;
assign n_45619 = ~n_31374 &  n_45618;
assign n_45620 = ~n_31368 &  n_45619;
assign n_45621 = ~n_31362 &  n_45620;
assign n_45622 = ~n_31356 &  n_45621;
assign n_45623 = ~n_31350 &  n_45622;
assign n_45624 = ~n_31344 &  n_45623;
assign n_45625 = ~n_31338 &  n_45624;
assign n_45626 = ~n_31332 &  n_45625;
assign n_45627 = ~n_31326 &  n_45626;
assign n_45628 = ~n_31320 &  n_45627;
assign n_45629 = ~n_31314 &  n_45628;
assign n_45630 = ~n_31308 &  n_45629;
assign n_45631 = ~n_31302 &  n_45630;
assign n_45632 = ~n_31296 &  n_45631;
assign n_45633 = ~n_31290 &  n_45632;
assign n_45634 = ~n_31284 &  n_45633;
assign n_45635 = ~n_31278 &  n_45634;
assign n_45636 = ~n_31272 &  n_45635;
assign n_45637 = ~n_31266 &  n_45636;
assign n_45638 = ~n_31260 &  n_45637;
assign n_45639 = ~n_31254 &  n_45638;
assign n_45640 = ~n_31248 &  n_45639;
assign n_45641 = ~n_31242 &  n_45640;
assign n_45642 = ~n_31236 &  n_45641;
assign n_45643 = ~n_31230 &  n_45642;
assign n_45644 = ~n_31224 &  n_45643;
assign n_45645 = ~n_31218 &  n_45644;
assign n_45646 = ~n_31212 &  n_45645;
assign n_45647 = ~n_31206 &  n_45646;
assign n_45648 = ~n_31200 &  n_45647;
assign n_45649 = ~n_31194 &  n_45648;
assign n_45650 = ~n_31188 &  n_45649;
assign n_45651 = ~n_31182 &  n_45650;
assign n_45652 = ~n_31176 &  n_45651;
assign n_45653 = ~n_31170 &  n_45652;
assign n_45654 = ~n_31164 &  n_45653;
assign n_45655 = ~n_31158 &  n_45654;
assign n_45656 = ~n_31152 &  n_45655;
assign n_45657 = ~n_31146 &  n_45656;
assign n_45658 = ~n_31140 &  n_45657;
assign n_45659 = ~n_31134 &  n_45658;
assign n_45660 = ~n_31124 &  n_45659;
assign n_45661 = ~n_31118 &  n_45660;
assign n_45662 = ~n_31112 &  n_45661;
assign n_45663 = ~n_31106 &  n_45662;
assign n_45664 = ~n_31100 &  n_45663;
assign n_45665 = ~n_31094 &  n_45664;
assign n_45666 = ~n_31088 &  n_45665;
assign n_45667 = ~n_31082 &  n_45666;
assign n_45668 = ~n_31076 &  n_45667;
assign n_45669 = ~n_31070 &  n_45668;
assign n_45670 = ~n_31064 &  n_45669;
assign n_45671 = ~n_31058 &  n_45670;
assign n_45672 = ~n_31052 &  n_45671;
assign n_45673 = ~n_31046 &  n_45672;
assign n_45674 = ~n_31040 &  n_45673;
assign n_45675 = ~n_31034 &  n_45674;
assign n_45676 = ~n_31028 &  n_45675;
assign n_45677 = ~n_31022 &  n_45676;
assign n_45678 = ~n_31016 &  n_45677;
assign n_45679 = ~n_31010 &  n_45678;
assign n_45680 = ~n_31004 &  n_45679;
assign n_45681 = ~n_30998 &  n_45680;
assign n_45682 = ~n_30992 &  n_45681;
assign n_45683 = ~n_30986 &  n_45682;
assign n_45684 = ~n_30980 &  n_45683;
assign n_45685 = ~n_30974 &  n_45684;
assign n_45686 = ~n_30968 &  n_45685;
assign n_45687 = ~n_30962 &  n_45686;
assign n_45688 = ~n_30956 &  n_45687;
assign n_45689 = ~n_30950 &  n_45688;
assign n_45690 = ~n_30944 &  n_45689;
assign n_45691 = ~n_30938 &  n_45690;
assign n_45692 = ~n_30932 &  n_45691;
assign n_45693 = ~n_30928 &  n_45692;
assign n_45694 = ~n_30924 &  n_45693;
assign n_45695 = ~n_30920 &  n_45694;
assign n_45696 = ~n_30916 &  n_45695;
assign n_45697 = ~n_30912 &  n_45696;
assign n_45698 = ~n_30908 &  n_45697;
assign n_45699 = ~n_30904 &  n_45698;
assign n_45700 = ~n_30900 &  n_45699;
assign n_45701 = ~n_30896 &  n_45700;
assign n_45702 = ~n_30892 &  n_45701;
assign n_45703 = ~n_30888 &  n_45702;
assign n_45704 = ~n_30884 &  n_45703;
assign n_45705 = ~n_30880 &  n_45704;
assign n_45706 = ~n_30876 &  n_45705;
assign n_45707 = ~n_30869 &  n_45706;
assign n_45708 = ~n_30864 &  n_45707;
assign n_45709 = ~n_30855 &  n_45708;
assign n_45710 = ~n_30849 &  n_45709;
assign n_45711 = ~n_30843 &  n_45710;
assign n_45712 = ~n_30837 &  n_45711;
assign n_45713 = ~n_30831 &  n_45712;
assign n_45714 = ~n_30825 &  n_45713;
assign n_45715 = ~n_30819 &  n_45714;
assign n_45716 = ~n_30813 &  n_45715;
assign n_45717 = ~n_30807 &  n_45716;
assign n_45718 = ~n_30801 &  n_45717;
assign n_45719 = ~n_30795 &  n_45718;
assign n_45720 = ~n_30789 &  n_45719;
assign n_45721 = ~n_30783 &  n_45720;
assign n_45722 = ~n_30777 &  n_45721;
assign n_45723 = ~n_30771 &  n_45722;
assign n_45724 = ~n_30765 &  n_45723;
assign n_45725 = ~n_30759 &  n_45724;
assign n_45726 = ~n_30753 &  n_45725;
assign n_45727 = ~n_30747 &  n_45726;
assign n_45728 = ~n_30741 &  n_45727;
assign n_45729 = ~n_30735 &  n_45728;
assign n_45730 = ~n_30729 &  n_45729;
assign n_45731 = ~n_30723 &  n_45730;
assign n_45732 = ~n_30717 &  n_45731;
assign n_45733 = ~n_30711 &  n_45732;
assign n_45734 = ~n_30705 &  n_45733;
assign n_45735 = ~n_30699 &  n_45734;
assign n_45736 = ~n_30693 &  n_45735;
assign n_45737 = ~n_30687 &  n_45736;
assign n_45738 = ~n_30681 &  n_45737;
assign n_45739 = ~n_30675 &  n_45738;
assign n_45740 = ~n_30669 &  n_45739;
assign n_45741 = ~n_30663 &  n_45740;
assign n_45742 = ~n_30657 &  n_45741;
assign n_45743 = ~n_30651 &  n_45742;
assign n_45744 = ~n_30645 &  n_45743;
assign n_45745 = ~n_30639 &  n_45744;
assign n_45746 = ~n_30633 &  n_45745;
assign n_45747 = ~n_30627 &  n_45746;
assign n_45748 = ~n_30621 &  n_45747;
assign n_45749 = ~n_30615 &  n_45748;
assign n_45750 = ~n_30609 &  n_45749;
assign n_45751 = ~n_30603 &  n_45750;
assign n_45752 = ~n_30597 &  n_45751;
assign n_45753 = ~n_30591 &  n_45752;
assign n_45754 = ~n_30585 &  n_45753;
assign n_45755 = ~n_30579 &  n_45754;
assign n_45756 = ~n_30573 &  n_45755;
assign n_45757 = ~n_30567 &  n_45756;
assign n_45758 = ~n_30561 &  n_45757;
assign n_45759 = ~n_30555 &  n_45758;
assign n_45760 = ~n_30549 &  n_45759;
assign n_45761 = ~n_30543 &  n_45760;
assign n_45762 = ~n_30537 &  n_45761;
assign n_45763 = ~n_30531 &  n_45762;
assign n_45764 = ~n_30525 &  n_45763;
assign n_45765 = ~n_30519 &  n_45764;
assign n_45766 = ~n_30513 &  n_45765;
assign n_45767 = ~n_30507 &  n_45766;
assign n_45768 = ~n_30501 &  n_45767;
assign n_45769 = ~n_30495 &  n_45768;
assign n_45770 = ~n_30489 &  n_45769;
assign n_45771 = ~n_30483 &  n_45770;
assign n_45772 = ~n_30477 &  n_45771;
assign n_45773 = ~n_30471 &  n_45772;
assign n_45774 = ~n_30465 &  n_45773;
assign n_45775 = ~n_30459 &  n_45774;
assign n_45776 = ~n_30453 &  n_45775;
assign n_45777 = ~n_30447 &  n_45776;
assign n_45778 = ~n_30441 &  n_45777;
assign n_45779 = ~n_30435 &  n_45778;
assign n_45780 = ~n_30429 &  n_45779;
assign n_45781 = ~n_30423 &  n_45780;
assign n_45782 = ~n_30417 &  n_45781;
assign n_45783 = ~n_30411 &  n_45782;
assign n_45784 = ~n_30405 &  n_45783;
assign n_45785 = ~n_30399 &  n_45784;
assign n_45786 = ~n_30393 &  n_45785;
assign n_45787 = ~n_30387 &  n_45786;
assign n_45788 = ~n_30381 &  n_45787;
assign n_45789 = ~n_30375 &  n_45788;
assign n_45790 = ~n_30369 &  n_45789;
assign n_45791 = ~n_30363 &  n_45790;
assign n_45792 = ~n_30357 &  n_45791;
assign n_45793 = ~n_30351 &  n_45792;
assign n_45794 = ~n_30345 &  n_45793;
assign n_45795 = ~n_30339 &  n_45794;
assign n_45796 = ~n_30333 &  n_45795;
assign n_45797 = ~n_30327 &  n_45796;
assign n_45798 = ~n_30321 &  n_45797;
assign n_45799 = ~n_30315 &  n_45798;
assign n_45800 = ~n_30309 &  n_45799;
assign n_45801 = ~n_30303 &  n_45800;
assign n_45802 = ~n_30297 &  n_45801;
assign n_45803 = ~n_30291 &  n_45802;
assign n_45804 = ~n_30285 &  n_45803;
assign n_45805 = ~n_30279 &  n_45804;
assign n_45806 = ~n_30273 &  n_45805;
assign n_45807 = ~n_30267 &  n_45806;
assign n_45808 = ~n_30261 &  n_45807;
assign n_45809 = ~n_30255 &  n_45808;
assign n_45810 = ~n_30249 &  n_45809;
assign n_45811 = ~n_30243 &  n_45810;
assign n_45812 = ~n_30237 &  n_45811;
assign n_45813 = ~n_30231 &  n_45812;
assign n_45814 = ~n_30225 &  n_45813;
assign n_45815 = ~n_30219 &  n_45814;
assign n_45816 = ~n_30213 &  n_45815;
assign n_45817 = ~n_30207 &  n_45816;
assign n_45818 = ~n_30201 &  n_45817;
assign n_45819 = ~n_30195 &  n_45818;
assign n_45820 = ~n_30189 &  n_45819;
assign n_45821 = ~n_30183 &  n_45820;
assign n_45822 = ~n_30177 &  n_45821;
assign n_45823 = ~n_30171 &  n_45822;
assign n_45824 = ~n_30165 &  n_45823;
assign n_45825 = ~n_30159 &  n_45824;
assign n_45826 = ~n_30153 &  n_45825;
assign n_45827 = ~n_30147 &  n_45826;
assign n_45828 = ~n_30141 &  n_45827;
assign n_45829 = ~n_30135 &  n_45828;
assign n_45830 = ~n_30129 &  n_45829;
assign n_45831 = ~n_30123 &  n_45830;
assign n_45832 = ~n_30117 &  n_45831;
assign n_45833 = ~n_30111 &  n_45832;
assign n_45834 = ~n_30105 &  n_45833;
assign n_45835 = ~n_30099 &  n_45834;
assign n_45836 = ~n_30093 &  n_45835;
assign n_45837 = ~n_30087 &  n_45836;
assign n_45838 = ~n_30069 &  n_45837;
assign n_45839 = ~n_30052 &  n_45838;
assign n_45840 = ~n_30035 &  n_45839;
assign n_45841 = ~n_30018 &  n_45840;
assign n_45842 = ~n_30001 &  n_45841;
assign n_45843 = ~n_29984 &  n_45842;
assign n_45844 = ~n_29967 &  n_45843;
assign n_45845 = ~n_29950 &  n_45844;
assign n_45846 = ~n_29933 &  n_45845;
assign n_45847 = ~n_29916 &  n_45846;
assign n_45848 = ~n_29899 &  n_45847;
assign n_45849 = ~n_29882 &  n_45848;
assign n_45850 = ~n_29865 &  n_45849;
assign n_45851 = ~n_29848 &  n_45850;
assign n_45852 = ~n_29831 &  n_45851;
assign n_45853 = ~n_29814 &  n_45852;
assign n_45854 = ~n_29797 &  n_45853;
assign n_45855 = ~n_29780 &  n_45854;
assign n_45856 = ~n_29763 &  n_45855;
assign n_45857 = ~n_29746 &  n_45856;
assign n_45858 = ~n_29729 &  n_45857;
assign n_45859 = ~n_29712 &  n_45858;
assign n_45860 = ~n_29695 &  n_45859;
assign n_45861 = ~n_29678 &  n_45860;
assign n_45862 = ~n_29661 &  n_45861;
assign n_45863 = ~n_29644 &  n_45862;
assign n_45864 = ~n_29627 &  n_45863;
assign n_45865 = ~n_29487 &  n_45864;
assign n_45866 = ~n_29362 &  n_45865;
assign n_45867 = ~n_29178 &  n_45866;
assign n_45868 = ~n_28977 &  n_45867;
assign n_45869 = ~n_28695 &  n_45868;
assign n_45870 = ~n_28357 &  n_45869;
assign n_45871 = ~n_28029 &  n_45870;
assign n_45872 = ~n_27362 &  n_45871;
assign n_45873 = ~n_26507 &  n_45872;
assign n_45874 = ~n_25716 &  n_45873;
assign n_45875 = ~n_21951 &  n_45874;
assign n_45876 = ~n_21945 &  n_45875;
assign n_45877 = ~n_21939 &  n_45876;
assign n_45878 = ~n_21933 &  n_45877;
assign n_45879 = ~n_21927 &  n_45878;
assign n_45880 = ~n_21921 &  n_45879;
assign n_45881 = ~n_21915 &  n_45880;
assign n_45882 = ~n_21909 &  n_45881;
assign n_45883 = ~n_21903 &  n_45882;
assign n_45884 = ~n_21897 &  n_45883;
assign n_45885 = ~n_21891 &  n_45884;
assign n_45886 = ~n_21885 &  n_45885;
assign n_45887 = ~n_21879 &  n_45886;
assign n_45888 = ~n_21873 &  n_45887;
assign n_45889 = ~n_21867 &  n_45888;
assign n_45890 = ~n_21861 &  n_45889;
assign n_45891 = ~n_21855 &  n_45890;
assign n_45892 = ~n_21849 &  n_45891;
assign n_45893 = ~n_21843 &  n_45892;
assign n_45894 = ~n_21837 &  n_45893;
assign n_45895 = ~n_21831 &  n_45894;
assign n_45896 = ~n_21825 &  n_45895;
assign n_45897 = ~n_21819 &  n_45896;
assign n_45898 = ~n_21813 &  n_45897;
assign n_45899 = ~n_21807 &  n_45898;
assign n_45900 = ~n_21801 &  n_45899;
assign n_45901 = ~n_21795 &  n_45900;
assign n_45902 = ~n_21789 &  n_45901;
assign n_45903 = ~n_21783 &  n_45902;
assign n_45904 = ~n_21777 &  n_45903;
assign n_45905 = ~n_21771 &  n_45904;
assign n_45906 = ~n_21765 &  n_45905;
assign n_45907 = ~n_21757 &  n_45906;
assign n_45908 = ~n_21751 &  n_45907;
assign n_45909 = ~n_21745 &  n_45908;
assign n_45910 = ~n_21739 &  n_45909;
assign n_45911 = ~n_21733 &  n_45910;
assign n_45912 = ~n_21727 &  n_45911;
assign n_45913 = ~n_21721 &  n_45912;
assign n_45914 = ~n_21715 &  n_45913;
assign n_45915 = ~n_21709 &  n_45914;
assign n_45916 = ~n_21703 &  n_45915;
assign n_45917 = ~n_21697 &  n_45916;
assign n_45918 = ~n_21691 &  n_45917;
assign n_45919 = ~n_21685 &  n_45918;
assign n_45920 = ~n_21679 &  n_45919;
assign n_45921 = ~n_21673 &  n_45920;
assign n_45922 = ~n_21667 &  n_45921;
assign n_45923 = ~n_21661 &  n_45922;
assign n_45924 = ~n_21655 &  n_45923;
assign n_45925 = ~n_21649 &  n_45924;
assign n_45926 = ~n_21643 &  n_45925;
assign n_45927 = ~n_21637 &  n_45926;
assign n_45928 = ~n_21631 &  n_45927;
assign n_45929 = ~n_21625 &  n_45928;
assign n_45930 = ~n_21619 &  n_45929;
assign n_45931 = ~n_21613 &  n_45930;
assign n_45932 = ~n_21607 &  n_45931;
assign n_45933 = ~n_21601 &  n_45932;
assign n_45934 = ~n_21595 &  n_45933;
assign n_45935 = ~n_21589 &  n_45934;
assign n_45936 = ~n_21583 &  n_45935;
assign n_45937 = ~n_21577 &  n_45936;
assign n_45938 = ~n_21571 &  n_45937;
assign n_45939 = ~n_21563 &  n_45938;
assign n_45940 = ~n_21557 &  n_45939;
assign n_45941 = ~n_21551 &  n_45940;
assign n_45942 = ~n_21545 &  n_45941;
assign n_45943 = ~n_21539 &  n_45942;
assign n_45944 = ~n_21533 &  n_45943;
assign n_45945 = ~n_21527 &  n_45944;
assign n_45946 = ~n_21521 &  n_45945;
assign n_45947 = ~n_21515 &  n_45946;
assign n_45948 = ~n_21509 &  n_45947;
assign n_45949 = ~n_21503 &  n_45948;
assign n_45950 = ~n_21497 &  n_45949;
assign n_45951 = ~n_21491 &  n_45950;
assign n_45952 = ~n_21485 &  n_45951;
assign n_45953 = ~n_21479 &  n_45952;
assign n_45954 = ~n_21473 &  n_45953;
assign n_45955 = ~n_21467 &  n_45954;
assign n_45956 = ~n_21461 &  n_45955;
assign n_45957 = ~n_21455 &  n_45956;
assign n_45958 = ~n_21449 &  n_45957;
assign n_45959 = ~n_21443 &  n_45958;
assign n_45960 = ~n_21437 &  n_45959;
assign n_45961 = ~n_21431 &  n_45960;
assign n_45962 = ~n_21425 &  n_45961;
assign n_45963 = ~n_21419 &  n_45962;
assign n_45964 = ~n_21413 &  n_45963;
assign n_45965 = ~n_21407 &  n_45964;
assign n_45966 = ~n_21401 &  n_45965;
assign n_45967 = ~n_21395 &  n_45966;
assign n_45968 = ~n_21389 &  n_45967;
assign n_45969 = ~n_21383 &  n_45968;
assign n_45970 = ~n_21377 &  n_45969;
assign n_45971 = ~n_21370 &  n_45970;
assign n_45972 = ~n_21364 &  n_45971;
assign n_45973 = ~n_21358 &  n_45972;
assign n_45974 = ~n_21352 &  n_45973;
assign n_45975 = ~n_21346 &  n_45974;
assign n_45976 = ~n_21340 &  n_45975;
assign n_45977 = ~n_21334 &  n_45976;
assign n_45978 = ~n_21328 &  n_45977;
assign n_45979 = ~n_21322 &  n_45978;
assign n_45980 = ~n_21316 &  n_45979;
assign n_45981 = ~n_21310 &  n_45980;
assign n_45982 = ~n_21304 &  n_45981;
assign n_45983 = ~n_21298 &  n_45982;
assign n_45984 = ~n_21292 &  n_45983;
assign n_45985 = ~n_21286 &  n_45984;
assign n_45986 = ~n_21280 &  n_45985;
assign n_45987 = ~n_21274 &  n_45986;
assign n_45988 = ~n_21268 &  n_45987;
assign n_45989 = ~n_21262 &  n_45988;
assign n_45990 = ~n_21256 &  n_45989;
assign n_45991 = ~n_21250 &  n_45990;
assign n_45992 = ~n_21244 &  n_45991;
assign n_45993 = ~n_21238 &  n_45992;
assign n_45994 = ~n_21232 &  n_45993;
assign n_45995 = ~n_21226 &  n_45994;
assign n_45996 = ~n_21220 &  n_45995;
assign n_45997 = ~n_21214 &  n_45996;
assign n_45998 = ~n_21208 &  n_45997;
assign n_45999 = ~n_21202 &  n_45998;
assign n_46000 = ~n_21196 &  n_45999;
assign n_46001 = ~n_21190 &  n_46000;
assign n_46002 = ~n_21184 &  n_46001;
assign n_46003 = ~n_21177 &  n_46002;
assign n_46004 = ~n_21171 &  n_46003;
assign n_46005 = ~n_21165 &  n_46004;
assign n_46006 = ~n_21159 &  n_46005;
assign n_46007 = ~n_21153 &  n_46006;
assign n_46008 = ~n_21147 &  n_46007;
assign n_46009 = ~n_21141 &  n_46008;
assign n_46010 = ~n_21135 &  n_46009;
assign n_46011 = ~n_21129 &  n_46010;
assign n_46012 = ~n_21123 &  n_46011;
assign n_46013 = ~n_21117 &  n_46012;
assign n_46014 = ~n_21111 &  n_46013;
assign n_46015 = ~n_21105 &  n_46014;
assign n_46016 = ~n_21099 &  n_46015;
assign n_46017 = ~n_21093 &  n_46016;
assign n_46018 = ~n_21087 &  n_46017;
assign n_46019 = ~n_21081 &  n_46018;
assign n_46020 = ~n_21075 &  n_46019;
assign n_46021 = ~n_21069 &  n_46020;
assign n_46022 = ~n_21063 &  n_46021;
assign n_46023 = ~n_21057 &  n_46022;
assign n_46024 = ~n_21051 &  n_46023;
assign n_46025 = ~n_21045 &  n_46024;
assign n_46026 = ~n_21039 &  n_46025;
assign n_46027 = ~n_21033 &  n_46026;
assign n_46028 = ~n_21027 &  n_46027;
assign n_46029 = ~n_21021 &  n_46028;
assign n_46030 = ~n_21015 &  n_46029;
assign n_46031 = ~n_21009 &  n_46030;
assign n_46032 = ~n_21003 &  n_46031;
assign n_46033 = ~n_20997 &  n_46032;
assign n_46034 = ~n_20991 &  n_46033;
assign n_46035 = ~n_20983 &  n_46034;
assign n_46036 = ~n_20977 &  n_46035;
assign n_46037 = ~n_20971 &  n_46036;
assign n_46038 = ~n_20965 &  n_46037;
assign n_46039 = ~n_20959 &  n_46038;
assign n_46040 = ~n_20953 &  n_46039;
assign n_46041 = ~n_20947 &  n_46040;
assign n_46042 = ~n_20941 &  n_46041;
assign n_46043 = ~n_20935 &  n_46042;
assign n_46044 = ~n_20929 &  n_46043;
assign n_46045 = ~n_20923 &  n_46044;
assign n_46046 = ~n_20917 &  n_46045;
assign n_46047 = ~n_20911 &  n_46046;
assign n_46048 = ~n_20905 &  n_46047;
assign n_46049 = ~n_20899 &  n_46048;
assign n_46050 = ~n_20893 &  n_46049;
assign n_46051 = ~n_20887 &  n_46050;
assign n_46052 = ~n_20881 &  n_46051;
assign n_46053 = ~n_20875 &  n_46052;
assign n_46054 = ~n_20869 &  n_46053;
assign n_46055 = ~n_20863 &  n_46054;
assign n_46056 = ~n_20857 &  n_46055;
assign n_46057 = ~n_20851 &  n_46056;
assign n_46058 = ~n_20845 &  n_46057;
assign n_46059 = ~n_20839 &  n_46058;
assign n_46060 = ~n_20833 &  n_46059;
assign n_46061 = ~n_20827 &  n_46060;
assign n_46062 = ~n_20821 &  n_46061;
assign n_46063 = ~n_20815 &  n_46062;
assign n_46064 = ~n_20809 &  n_46063;
assign n_46065 = ~n_20803 &  n_46064;
assign n_46066 = ~n_20797 &  n_46065;
assign n_46067 = ~n_20789 &  n_46066;
assign n_46068 = ~n_20783 &  n_46067;
assign n_46069 = ~n_20777 &  n_46068;
assign n_46070 = ~n_20771 &  n_46069;
assign n_46071 = ~n_20765 &  n_46070;
assign n_46072 = ~n_20759 &  n_46071;
assign n_46073 = ~n_20753 &  n_46072;
assign n_46074 = ~n_20747 &  n_46073;
assign n_46075 = ~n_20741 &  n_46074;
assign n_46076 = ~n_20735 &  n_46075;
assign n_46077 = ~n_20729 &  n_46076;
assign n_46078 = ~n_20723 &  n_46077;
assign n_46079 = ~n_20717 &  n_46078;
assign n_46080 = ~n_20711 &  n_46079;
assign n_46081 = ~n_20705 &  n_46080;
assign n_46082 = ~n_20699 &  n_46081;
assign n_46083 = ~n_20693 &  n_46082;
assign n_46084 = ~n_20687 &  n_46083;
assign n_46085 = ~n_20681 &  n_46084;
assign n_46086 = ~n_20675 &  n_46085;
assign n_46087 = ~n_20669 &  n_46086;
assign n_46088 = ~n_20663 &  n_46087;
assign n_46089 = ~n_20657 &  n_46088;
assign n_46090 = ~n_20651 &  n_46089;
assign n_46091 = ~n_20645 &  n_46090;
assign n_46092 = ~n_20639 &  n_46091;
assign n_46093 = ~n_20633 &  n_46092;
assign n_46094 = ~n_20627 &  n_46093;
assign n_46095 = ~n_20621 &  n_46094;
assign n_46096 = ~n_20615 &  n_46095;
assign n_46097 = ~n_20609 &  n_46096;
assign n_46098 = ~n_20603 &  n_46097;
assign n_46099 = ~n_20595 &  n_46098;
assign n_46100 = ~n_20589 &  n_46099;
assign n_46101 = ~n_20583 &  n_46100;
assign n_46102 = ~n_20577 &  n_46101;
assign n_46103 = ~n_20571 &  n_46102;
assign n_46104 = ~n_20565 &  n_46103;
assign n_46105 = ~n_20559 &  n_46104;
assign n_46106 = ~n_20553 &  n_46105;
assign n_46107 = ~n_20547 &  n_46106;
assign n_46108 = ~n_20541 &  n_46107;
assign n_46109 = ~n_20535 &  n_46108;
assign n_46110 = ~n_20529 &  n_46109;
assign n_46111 = ~n_20523 &  n_46110;
assign n_46112 = ~n_20517 &  n_46111;
assign n_46113 = ~n_20511 &  n_46112;
assign n_46114 = ~n_20505 &  n_46113;
assign n_46115 = ~n_20499 &  n_46114;
assign n_46116 = ~n_20493 &  n_46115;
assign n_46117 = ~n_20487 &  n_46116;
assign n_46118 = ~n_20481 &  n_46117;
assign n_46119 = ~n_20475 &  n_46118;
assign n_46120 = ~n_20469 &  n_46119;
assign n_46121 = ~n_20463 &  n_46120;
assign n_46122 = ~n_20457 &  n_46121;
assign n_46123 = ~n_20451 &  n_46122;
assign n_46124 = ~n_20445 &  n_46123;
assign n_46125 = ~n_20439 &  n_46124;
assign n_46126 = ~n_20433 &  n_46125;
assign n_46127 = ~n_20427 &  n_46126;
assign n_46128 = ~n_20421 &  n_46127;
assign n_46129 = ~n_20415 &  n_46128;
assign n_46130 = ~n_20409 &  n_46129;
assign n_46131 = ~n_20400 &  n_46130;
assign n_46132 = ~n_20394 &  n_46131;
assign n_46133 = ~n_20388 &  n_46132;
assign n_46134 = ~n_20382 &  n_46133;
assign n_46135 = ~n_20376 &  n_46134;
assign n_46136 = ~n_20370 &  n_46135;
assign n_46137 = ~n_20364 &  n_46136;
assign n_46138 = ~n_20358 &  n_46137;
assign n_46139 = ~n_20352 &  n_46138;
assign n_46140 = ~n_20346 &  n_46139;
assign n_46141 = ~n_20340 &  n_46140;
assign n_46142 = ~n_20334 &  n_46141;
assign n_46143 = ~n_20328 &  n_46142;
assign n_46144 = ~n_20322 &  n_46143;
assign n_46145 = ~n_20316 &  n_46144;
assign n_46146 = ~n_20310 &  n_46145;
assign n_46147 = ~n_20304 &  n_46146;
assign n_46148 = ~n_20298 &  n_46147;
assign n_46149 = ~n_20292 &  n_46148;
assign n_46150 = ~n_20286 &  n_46149;
assign n_46151 = ~n_20280 &  n_46150;
assign n_46152 = ~n_20274 &  n_46151;
assign n_46153 = ~n_20268 &  n_46152;
assign n_46154 = ~n_20262 &  n_46153;
assign n_46155 = ~n_20256 &  n_46154;
assign n_46156 = ~n_20250 &  n_46155;
assign n_46157 = ~n_20244 &  n_46156;
assign n_46158 = ~n_20238 &  n_46157;
assign n_46159 = ~n_20232 &  n_46158;
assign n_46160 = ~n_20226 &  n_46159;
assign n_46161 = ~n_20220 &  n_46160;
assign n_46162 = ~n_20214 &  n_46161;
assign n_46163 = ~n_20206 &  n_46162;
assign n_46164 = ~n_20202 &  n_46163;
assign n_46165 = ~n_20198 &  n_46164;
assign n_46166 = ~n_20194 &  n_46165;
assign n_46167 = ~n_20190 &  n_46166;
assign n_46168 = ~n_20186 &  n_46167;
assign n_46169 = ~n_20182 &  n_46168;
assign n_46170 = ~n_20178 &  n_46169;
assign n_46171 = ~n_20174 &  n_46170;
assign n_46172 = ~n_20170 &  n_46171;
assign n_46173 = ~n_20166 &  n_46172;
assign n_46174 = ~n_20162 &  n_46173;
assign n_46175 = ~n_20158 &  n_46174;
assign n_46176 = ~n_20154 &  n_46175;
assign n_46177 = ~n_20150 &  n_46176;
assign n_46178 = ~n_20146 &  n_46177;
assign n_46179 = ~n_20142 &  n_46178;
assign n_46180 = ~n_20138 &  n_46179;
assign n_46181 = ~n_20134 &  n_46180;
assign n_46182 = ~n_20130 &  n_46181;
assign n_46183 = ~n_20126 &  n_46182;
assign n_46184 = ~n_20122 &  n_46183;
assign n_46185 = ~n_20118 &  n_46184;
assign n_46186 = ~n_20114 &  n_46185;
assign n_46187 = ~n_20110 &  n_46186;
assign n_46188 = ~n_20106 &  n_46187;
assign n_46189 = ~n_20102 &  n_46188;
assign n_46190 = ~n_20098 &  n_46189;
assign n_46191 = ~n_20094 &  n_46190;
assign n_46192 = ~n_20090 &  n_46191;
assign n_46193 = ~n_20086 &  n_46192;
assign n_46194 = ~n_20082 &  n_46193;
assign n_46195 = ~n_20076 &  n_46194;
assign n_46196 = ~n_20070 &  n_46195;
assign n_46197 = ~n_20064 &  n_46196;
assign n_46198 = ~n_20058 &  n_46197;
assign n_46199 = ~n_20052 &  n_46198;
assign n_46200 = ~n_20046 &  n_46199;
assign n_46201 = ~n_20040 &  n_46200;
assign n_46202 = ~n_20034 &  n_46201;
assign n_46203 = ~n_20028 &  n_46202;
assign n_46204 = ~n_20022 &  n_46203;
assign n_46205 = ~n_20016 &  n_46204;
assign n_46206 = ~n_20010 &  n_46205;
assign n_46207 = ~n_20004 &  n_46206;
assign n_46208 = ~n_19998 &  n_46207;
assign n_46209 = ~n_19992 &  n_46208;
assign n_46210 = ~n_19986 &  n_46209;
assign n_46211 = ~n_19980 &  n_46210;
assign n_46212 = ~n_19974 &  n_46211;
assign n_46213 = ~n_19968 &  n_46212;
assign n_46214 = ~n_19962 &  n_46213;
assign n_46215 = ~n_19956 &  n_46214;
assign n_46216 = ~n_19950 &  n_46215;
assign n_46217 = ~n_19944 &  n_46216;
assign n_46218 = ~n_19938 &  n_46217;
assign n_46219 = ~n_19932 &  n_46218;
assign n_46220 = ~n_19926 &  n_46219;
assign n_46221 = ~n_19920 &  n_46220;
assign n_46222 = ~n_19914 &  n_46221;
assign n_46223 = ~n_19908 &  n_46222;
assign n_46224 = ~n_19902 &  n_46223;
assign n_46225 = ~n_19896 &  n_46224;
assign n_46226 = ~n_19890 &  n_46225;
assign n_46227 = ~n_19884 &  n_46226;
assign n_46228 = ~n_19880 &  n_46227;
assign n_46229 = ~n_19874 &  n_46228;
assign n_46230 = ~n_19868 &  n_46229;
assign n_46231 = ~n_19862 &  n_46230;
assign n_46232 = ~n_19856 &  n_46231;
assign n_46233 = ~n_19850 &  n_46232;
assign n_46234 = ~n_19844 &  n_46233;
assign n_46235 = ~n_19838 &  n_46234;
assign n_46236 = ~n_19832 &  n_46235;
assign n_46237 = ~n_19826 &  n_46236;
assign n_46238 = ~n_19820 &  n_46237;
assign n_46239 = ~n_19814 &  n_46238;
assign n_46240 = ~n_19808 &  n_46239;
assign n_46241 = ~n_19802 &  n_46240;
assign n_46242 = ~n_19796 &  n_46241;
assign n_46243 = ~n_19790 &  n_46242;
assign n_46244 = ~n_19784 &  n_46243;
assign n_46245 = ~n_19778 &  n_46244;
assign n_46246 = ~n_19772 &  n_46245;
assign n_46247 = ~n_19766 &  n_46246;
assign n_46248 = ~n_19760 &  n_46247;
assign n_46249 = ~n_19754 &  n_46248;
assign n_46250 = ~n_19748 &  n_46249;
assign n_46251 = ~n_19742 &  n_46250;
assign n_46252 = ~n_19736 &  n_46251;
assign n_46253 = ~n_19730 &  n_46252;
assign n_46254 = ~n_19724 &  n_46253;
assign n_46255 = ~n_19718 &  n_46254;
assign n_46256 = ~n_19712 &  n_46255;
assign n_46257 = ~n_19706 &  n_46256;
assign n_46258 = ~n_19700 &  n_46257;
assign n_46259 = ~n_19693 &  n_46258;
assign n_46260 = ~n_19687 &  n_46259;
assign n_46261 = ~n_19681 &  n_46260;
assign n_46262 = ~n_19675 &  n_46261;
assign n_46263 = ~n_19669 &  n_46262;
assign n_46264 = ~n_19663 &  n_46263;
assign n_46265 = ~n_19657 &  n_46264;
assign n_46266 = ~n_19651 &  n_46265;
assign n_46267 = ~n_19645 &  n_46266;
assign n_46268 = ~n_19639 &  n_46267;
assign n_46269 = ~n_19633 &  n_46268;
assign n_46270 = ~n_19627 &  n_46269;
assign n_46271 = ~n_19621 &  n_46270;
assign n_46272 = ~n_19615 &  n_46271;
assign n_46273 = ~n_19609 &  n_46272;
assign n_46274 = ~n_19603 &  n_46273;
assign n_46275 = ~n_19597 &  n_46274;
assign n_46276 = ~n_19591 &  n_46275;
assign n_46277 = ~n_19585 &  n_46276;
assign n_46278 = ~n_19579 &  n_46277;
assign n_46279 = ~n_19573 &  n_46278;
assign n_46280 = ~n_19567 &  n_46279;
assign n_46281 = ~n_19561 &  n_46280;
assign n_46282 = ~n_19555 &  n_46281;
assign n_46283 = ~n_19549 &  n_46282;
assign n_46284 = ~n_19543 &  n_46283;
assign n_46285 = ~n_19537 &  n_46284;
assign n_46286 = ~n_19531 &  n_46285;
assign n_46287 = ~n_19525 &  n_46286;
assign n_46288 = ~n_19519 &  n_46287;
assign n_46289 = ~n_19513 &  n_46288;
assign n_46290 = ~n_19507 &  n_46289;
assign n_46291 = ~n_19492 &  n_46290;
assign n_46292 = ~n_19486 &  n_46291;
assign n_46293 = ~n_19480 &  n_46292;
assign n_46294 = ~n_19474 &  n_46293;
assign n_46295 = ~n_19468 &  n_46294;
assign n_46296 = ~n_19462 &  n_46295;
assign n_46297 = ~n_19456 &  n_46296;
assign n_46298 = ~n_19450 &  n_46297;
assign n_46299 = ~n_19444 &  n_46298;
assign n_46300 = ~n_19438 &  n_46299;
assign n_46301 = ~n_19432 &  n_46300;
assign n_46302 = ~n_19426 &  n_46301;
assign n_46303 = ~n_19420 &  n_46302;
assign n_46304 = ~n_19414 &  n_46303;
assign n_46305 = ~n_19408 &  n_46304;
assign n_46306 = ~n_19402 &  n_46305;
assign n_46307 = ~n_19396 &  n_46306;
assign n_46308 = ~n_19390 &  n_46307;
assign n_46309 = ~n_19384 &  n_46308;
assign n_46310 = ~n_19378 &  n_46309;
assign n_46311 = ~n_19372 &  n_46310;
assign n_46312 = ~n_19366 &  n_46311;
assign n_46313 = ~n_19360 &  n_46312;
assign n_46314 = ~n_19354 &  n_46313;
assign n_46315 = ~n_19348 &  n_46314;
assign n_46316 = ~n_19342 &  n_46315;
assign n_46317 = ~n_19336 &  n_46316;
assign n_46318 = ~n_19330 &  n_46317;
assign n_46319 = ~n_19324 &  n_46318;
assign n_46320 = ~n_19318 &  n_46319;
assign n_46321 = ~n_19312 &  n_46320;
assign n_46322 = ~n_19306 &  n_46321;
assign n_46323 = ~n_19300 &  n_46322;
assign n_46324 = ~n_19294 &  n_46323;
assign n_46325 = ~n_19288 &  n_46324;
assign n_46326 = ~n_19282 &  n_46325;
assign n_46327 = ~n_19276 &  n_46326;
assign n_46328 = ~n_19270 &  n_46327;
assign n_46329 = ~n_19264 &  n_46328;
assign n_46330 = ~n_19258 &  n_46329;
assign n_46331 = ~n_19252 &  n_46330;
assign n_46332 = ~n_19246 &  n_46331;
assign n_46333 = ~n_19240 &  n_46332;
assign n_46334 = ~n_19234 &  n_46333;
assign n_46335 = ~n_19228 &  n_46334;
assign n_46336 = ~n_19222 &  n_46335;
assign n_46337 = ~n_19216 &  n_46336;
assign n_46338 = ~n_19210 &  n_46337;
assign n_46339 = ~n_19204 &  n_46338;
assign n_46340 = ~n_19198 &  n_46339;
assign n_46341 = ~n_19192 &  n_46340;
assign n_46342 = ~n_19186 &  n_46341;
assign n_46343 = ~n_19180 &  n_46342;
assign n_46344 = ~n_19174 &  n_46343;
assign n_46345 = ~n_19168 &  n_46344;
assign n_46346 = ~n_19162 &  n_46345;
assign n_46347 = ~n_19156 &  n_46346;
assign n_46348 = ~n_19150 &  n_46347;
assign n_46349 = ~n_19144 &  n_46348;
assign n_46350 = ~n_19138 &  n_46349;
assign n_46351 = ~n_19132 &  n_46350;
assign n_46352 = ~n_19126 &  n_46351;
assign n_46353 = ~n_19120 &  n_46352;
assign n_46354 = ~n_19114 &  n_46353;
assign n_46355 = ~n_19107 &  n_46354;
assign n_46356 = ~n_19101 &  n_46355;
assign n_46357 = ~n_19095 &  n_46356;
assign n_46358 = ~n_19089 &  n_46357;
assign n_46359 = ~n_19083 &  n_46358;
assign n_46360 = ~n_19077 &  n_46359;
assign n_46361 = ~n_19071 &  n_46360;
assign n_46362 = ~n_19065 &  n_46361;
assign n_46363 = ~n_19059 &  n_46362;
assign n_46364 = ~n_19053 &  n_46363;
assign n_46365 = ~n_19047 &  n_46364;
assign n_46366 = ~n_19041 &  n_46365;
assign n_46367 = ~n_19035 &  n_46366;
assign n_46368 = ~n_19029 &  n_46367;
assign n_46369 = ~n_19023 &  n_46368;
assign n_46370 = ~n_19017 &  n_46369;
assign n_46371 = ~n_19011 &  n_46370;
assign n_46372 = ~n_19005 &  n_46371;
assign n_46373 = ~n_18999 &  n_46372;
assign n_46374 = ~n_18993 &  n_46373;
assign n_46375 = ~n_18987 &  n_46374;
assign n_46376 = ~n_18981 &  n_46375;
assign n_46377 = ~n_18975 &  n_46376;
assign n_46378 = ~n_18969 &  n_46377;
assign n_46379 = ~n_18963 &  n_46378;
assign n_46380 = ~n_18957 &  n_46379;
assign n_46381 = ~n_18951 &  n_46380;
assign n_46382 = ~n_18945 &  n_46381;
assign n_46383 = ~n_18939 &  n_46382;
assign n_46384 = ~n_18933 &  n_46383;
assign n_46385 = ~n_18927 &  n_46384;
assign n_46386 = ~n_18921 &  n_46385;
assign n_46387 = ~n_18913 &  n_46386;
assign n_46388 = ~n_18908 &  n_46387;
assign n_46389 = ~n_18903 &  n_46388;
assign n_46390 = ~n_18898 &  n_46389;
assign n_46391 = ~n_18893 &  n_46390;
assign n_46392 = ~n_18888 &  n_46391;
assign n_46393 = ~n_18883 &  n_46392;
assign n_46394 = ~n_18878 &  n_46393;
assign n_46395 = ~n_18873 &  n_46394;
assign n_46396 = ~n_18868 &  n_46395;
assign n_46397 = ~n_18863 &  n_46396;
assign n_46398 = ~n_18858 &  n_46397;
assign n_46399 = ~n_18853 &  n_46398;
assign n_46400 = ~n_18848 &  n_46399;
assign n_46401 = ~n_18843 &  n_46400;
assign n_46402 = ~n_18838 &  n_46401;
assign n_46403 = ~n_18833 &  n_46402;
assign n_46404 = ~n_18828 &  n_46403;
assign n_46405 = ~n_18823 &  n_46404;
assign n_46406 = ~n_18818 &  n_46405;
assign n_46407 = ~n_18813 &  n_46406;
assign n_46408 = ~n_18808 &  n_46407;
assign n_46409 = ~n_18803 &  n_46408;
assign n_46410 = ~n_18798 &  n_46409;
assign n_46411 = ~n_18793 &  n_46410;
assign n_46412 = ~n_18788 &  n_46411;
assign n_46413 = ~n_18783 &  n_46412;
assign n_46414 = ~n_18778 &  n_46413;
assign n_46415 = ~n_18773 &  n_46414;
assign n_46416 = ~n_18768 &  n_46415;
assign n_46417 = ~n_18763 &  n_46416;
assign n_46418 = ~n_18758 &  n_46417;
assign n_46419 = ~n_18753 &  n_46418;
assign n_46420 = ~n_18749 &  n_46419;
assign n_46421 = ~n_18745 &  n_46420;
assign n_46422 = ~n_18741 &  n_46421;
assign n_46423 = ~n_18737 &  n_46422;
assign n_46424 = ~n_18733 &  n_46423;
assign n_46425 = ~n_18729 &  n_46424;
assign n_46426 = ~n_18725 &  n_46425;
assign n_46427 = ~n_18721 &  n_46426;
assign n_46428 = ~n_18717 &  n_46427;
assign n_46429 = ~n_18713 &  n_46428;
assign n_46430 = ~n_18709 &  n_46429;
assign n_46431 = ~n_18705 &  n_46430;
assign n_46432 = ~n_18701 &  n_46431;
assign n_46433 = ~n_18697 &  n_46432;
assign n_46434 = ~n_18693 &  n_46433;
assign n_46435 = ~n_18689 &  n_46434;
assign n_46436 = ~n_18685 &  n_46435;
assign n_46437 = ~n_18681 &  n_46436;
assign n_46438 = ~n_18677 &  n_46437;
assign n_46439 = ~n_18673 &  n_46438;
assign n_46440 = ~n_18669 &  n_46439;
assign n_46441 = ~n_18665 &  n_46440;
assign n_46442 = ~n_18661 &  n_46441;
assign n_46443 = ~n_18657 &  n_46442;
assign n_46444 = ~n_18653 &  n_46443;
assign n_46445 = ~n_18649 &  n_46444;
assign n_46446 = ~n_18645 &  n_46445;
assign n_46447 = ~n_18641 &  n_46446;
assign n_46448 = ~n_18637 &  n_46447;
assign n_46449 = ~n_18633 &  n_46448;
assign n_46450 = ~n_18629 &  n_46449;
assign n_46451 = ~n_18623 &  n_46450;
assign n_46452 = ~n_18619 &  n_46451;
assign n_46453 = ~n_18615 &  n_46452;
assign n_46454 = ~n_18611 &  n_46453;
assign n_46455 = ~n_18607 &  n_46454;
assign n_46456 = ~n_18603 &  n_46455;
assign n_46457 = ~n_18599 &  n_46456;
assign n_46458 = ~n_18595 &  n_46457;
assign n_46459 = ~n_18591 &  n_46458;
assign n_46460 = ~n_18587 &  n_46459;
assign n_46461 = ~n_18583 &  n_46460;
assign n_46462 = ~n_18579 &  n_46461;
assign n_46463 = ~n_18575 &  n_46462;
assign n_46464 = ~n_18571 &  n_46463;
assign n_46465 = ~n_18567 &  n_46464;
assign n_46466 = ~n_18563 &  n_46465;
assign n_46467 = ~n_18559 &  n_46466;
assign n_46468 = ~n_18555 &  n_46467;
assign n_46469 = ~n_18551 &  n_46468;
assign n_46470 = ~n_18547 &  n_46469;
assign n_46471 = ~n_18543 &  n_46470;
assign n_46472 = ~n_18539 &  n_46471;
assign n_46473 = ~n_18535 &  n_46472;
assign n_46474 = ~n_18531 &  n_46473;
assign n_46475 = ~n_18527 &  n_46474;
assign n_46476 = ~n_18523 &  n_46475;
assign n_46477 = ~n_18519 &  n_46476;
assign n_46478 = ~n_18515 &  n_46477;
assign n_46479 = ~n_18511 &  n_46478;
assign n_46480 = ~n_18507 &  n_46479;
assign n_46481 = ~n_18503 &  n_46480;
assign n_46482 = ~n_18499 &  n_46481;
assign n_46483 = ~n_18494 &  n_46482;
assign n_46484 = ~n_18488 &  n_46483;
assign n_46485 = ~n_18482 &  n_46484;
assign n_46486 = ~n_18476 &  n_46485;
assign n_46487 = ~n_18470 &  n_46486;
assign n_46488 = ~n_18464 &  n_46487;
assign n_46489 = ~n_18458 &  n_46488;
assign n_46490 = ~n_18452 &  n_46489;
assign n_46491 = ~n_18446 &  n_46490;
assign n_46492 = ~n_18440 &  n_46491;
assign n_46493 = ~n_18434 &  n_46492;
assign n_46494 = ~n_18428 &  n_46493;
assign n_46495 = ~n_18422 &  n_46494;
assign n_46496 = ~n_18416 &  n_46495;
assign n_46497 = ~n_18410 &  n_46496;
assign n_46498 = ~n_18404 &  n_46497;
assign n_46499 = ~n_18398 &  n_46498;
assign n_46500 = ~n_18392 &  n_46499;
assign n_46501 = ~n_18386 &  n_46500;
assign n_46502 = ~n_18380 &  n_46501;
assign n_46503 = ~n_18374 &  n_46502;
assign n_46504 = ~n_18368 &  n_46503;
assign n_46505 = ~n_18362 &  n_46504;
assign n_46506 = ~n_18356 &  n_46505;
assign n_46507 = ~n_18350 &  n_46506;
assign n_46508 = ~n_18344 &  n_46507;
assign n_46509 = ~n_18338 &  n_46508;
assign n_46510 = ~n_18332 &  n_46509;
assign n_46511 = ~n_18326 &  n_46510;
assign n_46512 = ~n_18320 &  n_46511;
assign n_46513 = ~n_18314 &  n_46512;
assign n_46514 = ~n_18308 &  n_46513;
assign n_46515 = ~n_18301 &  n_46514;
assign n_46516 = ~n_18295 &  n_46515;
assign n_46517 = ~n_18289 &  n_46516;
assign n_46518 = ~n_18283 &  n_46517;
assign n_46519 = ~n_18277 &  n_46518;
assign n_46520 = ~n_18271 &  n_46519;
assign n_46521 = ~n_18265 &  n_46520;
assign n_46522 = ~n_18259 &  n_46521;
assign n_46523 = ~n_18253 &  n_46522;
assign n_46524 = ~n_18247 &  n_46523;
assign n_46525 = ~n_18241 &  n_46524;
assign n_46526 = ~n_18235 &  n_46525;
assign n_46527 = ~n_18229 &  n_46526;
assign n_46528 = ~n_18223 &  n_46527;
assign n_46529 = ~n_18217 &  n_46528;
assign n_46530 = ~n_18211 &  n_46529;
assign n_46531 = ~n_18205 &  n_46530;
assign n_46532 = ~n_18199 &  n_46531;
assign n_46533 = ~n_18193 &  n_46532;
assign n_46534 = ~n_18187 &  n_46533;
assign n_46535 = ~n_18181 &  n_46534;
assign n_46536 = ~n_18175 &  n_46535;
assign n_46537 = ~n_18169 &  n_46536;
assign n_46538 = ~n_18163 &  n_46537;
assign n_46539 = ~n_18157 &  n_46538;
assign n_46540 = ~n_18151 &  n_46539;
assign n_46541 = ~n_18145 &  n_46540;
assign n_46542 = ~n_18139 &  n_46541;
assign n_46543 = ~n_18133 &  n_46542;
assign n_46544 = ~n_18127 &  n_46543;
assign n_46545 = ~n_18121 &  n_46544;
assign n_46546 = ~n_18115 &  n_46545;
assign n_46547 = ~n_18108 &  n_46546;
assign n_46548 = ~n_18104 &  n_46547;
assign n_46549 = ~n_18100 &  n_46548;
assign n_46550 = ~n_18096 &  n_46549;
assign n_46551 = ~n_18092 &  n_46550;
assign n_46552 = ~n_18088 &  n_46551;
assign n_46553 = ~n_18084 &  n_46552;
assign n_46554 = ~n_18080 &  n_46553;
assign n_46555 = ~n_18076 &  n_46554;
assign n_46556 = ~n_18072 &  n_46555;
assign n_46557 = ~n_18068 &  n_46556;
assign n_46558 = ~n_18064 &  n_46557;
assign n_46559 = ~n_18060 &  n_46558;
assign n_46560 = ~n_18056 &  n_46559;
assign n_46561 = ~n_18052 &  n_46560;
assign n_46562 = ~n_18048 &  n_46561;
assign n_46563 = ~n_18044 &  n_46562;
assign n_46564 = ~n_18040 &  n_46563;
assign n_46565 = ~n_18036 &  n_46564;
assign n_46566 = ~n_18032 &  n_46565;
assign n_46567 = ~n_18028 &  n_46566;
assign n_46568 = ~n_18024 &  n_46567;
assign n_46569 = ~n_18020 &  n_46568;
assign n_46570 = ~n_18016 &  n_46569;
assign n_46571 = ~n_18012 &  n_46570;
assign n_46572 = ~n_18008 &  n_46571;
assign n_46573 = ~n_18004 &  n_46572;
assign n_46574 = ~n_18000 &  n_46573;
assign n_46575 = ~n_17996 &  n_46574;
assign n_46576 = ~n_17992 &  n_46575;
assign n_46577 = ~n_17988 &  n_46576;
assign n_46578 = ~n_17984 &  n_46577;
assign n_46579 = ~n_17979 &  n_46578;
assign n_46580 = ~n_17973 &  n_46579;
assign n_46581 = ~n_17967 &  n_46580;
assign n_46582 = ~n_17961 &  n_46581;
assign n_46583 = ~n_17955 &  n_46582;
assign n_46584 = ~n_17949 &  n_46583;
assign n_46585 = ~n_17943 &  n_46584;
assign n_46586 = ~n_17937 &  n_46585;
assign n_46587 = ~n_17931 &  n_46586;
assign n_46588 = ~n_17925 &  n_46587;
assign n_46589 = ~n_17919 &  n_46588;
assign n_46590 = ~n_17913 &  n_46589;
assign n_46591 = ~n_17907 &  n_46590;
assign n_46592 = ~n_17901 &  n_46591;
assign n_46593 = ~n_17895 &  n_46592;
assign n_46594 = ~n_17889 &  n_46593;
assign n_46595 = ~n_17883 &  n_46594;
assign n_46596 = ~n_17877 &  n_46595;
assign n_46597 = ~n_17871 &  n_46596;
assign n_46598 = ~n_17865 &  n_46597;
assign n_46599 = ~n_17859 &  n_46598;
assign n_46600 = ~n_17853 &  n_46599;
assign n_46601 = ~n_17847 &  n_46600;
assign n_46602 = ~n_17841 &  n_46601;
assign n_46603 = ~n_17835 &  n_46602;
assign n_46604 = ~n_17829 &  n_46603;
assign n_46605 = ~n_17823 &  n_46604;
assign n_46606 = ~n_17817 &  n_46605;
assign n_46607 = ~n_17811 &  n_46606;
assign n_46608 = ~n_17805 &  n_46607;
assign n_46609 = ~n_17799 &  n_46608;
assign n_46610 = ~n_17793 &  n_46609;
assign n_46611 = ~n_17781 &  n_46610;
assign n_46612 = ~n_17764 &  n_46611;
assign n_46613 = ~n_17747 &  n_46612;
assign n_46614 = ~n_17730 &  n_46613;
assign n_46615 = ~n_17713 &  n_46614;
assign n_46616 = ~n_17696 &  n_46615;
assign n_46617 = ~n_17679 &  n_46616;
assign n_46618 = ~n_17662 &  n_46617;
assign n_46619 = ~n_17645 &  n_46618;
assign n_46620 = ~n_17628 &  n_46619;
assign n_46621 = ~n_17611 &  n_46620;
assign n_46622 = ~n_17594 &  n_46621;
assign n_46623 = ~n_17577 &  n_46622;
assign n_46624 = ~n_17560 &  n_46623;
assign n_46625 = ~n_17543 &  n_46624;
assign n_46626 = ~n_17526 &  n_46625;
assign n_46627 = ~n_17509 &  n_46626;
assign n_46628 = ~n_17492 &  n_46627;
assign n_46629 = ~n_17475 &  n_46628;
assign n_46630 = ~n_17458 &  n_46629;
assign n_46631 = ~n_17441 &  n_46630;
assign n_46632 = ~n_17424 &  n_46631;
assign n_46633 = ~n_17407 &  n_46632;
assign n_46634 = ~n_17390 &  n_46633;
assign n_46635 = ~n_17373 &  n_46634;
assign n_46636 = ~n_17356 &  n_46635;
assign n_46637 = ~n_17339 &  n_46636;
assign n_46638 = ~n_17322 &  n_46637;
assign n_46639 = ~n_17305 &  n_46638;
assign n_46640 = ~n_17288 &  n_46639;
assign n_46641 = ~n_17271 &  n_46640;
assign n_46642 = ~n_17254 &  n_46641;
assign n_46643 = ~n_17205 &  n_46642;
assign n_46644 = ~n_17201 &  n_46643;
assign n_46645 = ~n_17197 &  n_46644;
assign n_46646 = ~n_17193 &  n_46645;
assign n_46647 = ~n_17189 &  n_46646;
assign n_46648 = ~n_17185 &  n_46647;
assign n_46649 = ~n_17181 &  n_46648;
assign n_46650 = ~n_17177 &  n_46649;
assign n_46651 = ~n_17173 &  n_46650;
assign n_46652 = ~n_17169 &  n_46651;
assign n_46653 = ~n_17165 &  n_46652;
assign n_46654 = ~n_17161 &  n_46653;
assign n_46655 = ~n_17157 &  n_46654;
assign n_46656 = ~n_17153 &  n_46655;
assign n_46657 = ~n_17149 &  n_46656;
assign n_46658 = ~n_17145 &  n_46657;
assign n_46659 = ~n_17141 &  n_46658;
assign n_46660 = ~n_17137 &  n_46659;
assign n_46661 = ~n_17133 &  n_46660;
assign n_46662 = ~n_17129 &  n_46661;
assign n_46663 = ~n_17125 &  n_46662;
assign n_46664 = ~n_17121 &  n_46663;
assign n_46665 = ~n_17117 &  n_46664;
assign n_46666 = ~n_17113 &  n_46665;
assign n_46667 = ~n_17109 &  n_46666;
assign n_46668 = ~n_17105 &  n_46667;
assign n_46669 = ~n_17101 &  n_46668;
assign n_46670 = ~n_17097 &  n_46669;
assign n_46671 = ~n_17093 &  n_46670;
assign n_46672 = ~n_17089 &  n_46671;
assign n_46673 = ~n_17085 &  n_46672;
assign n_46674 = ~n_17081 &  n_46673;
assign n_46675 = ~n_17075 &  n_46674;
assign n_46676 = ~n_17069 &  n_46675;
assign n_46677 = ~n_17063 &  n_46676;
assign n_46678 = ~n_17057 &  n_46677;
assign n_46679 = ~n_17051 &  n_46678;
assign n_46680 = ~n_17045 &  n_46679;
assign n_46681 = ~n_17039 &  n_46680;
assign n_46682 = ~n_17033 &  n_46681;
assign n_46683 = ~n_17027 &  n_46682;
assign n_46684 = ~n_17021 &  n_46683;
assign n_46685 = ~n_17015 &  n_46684;
assign n_46686 = ~n_17009 &  n_46685;
assign n_46687 = ~n_17003 &  n_46686;
assign n_46688 = ~n_16997 &  n_46687;
assign n_46689 = ~n_16991 &  n_46688;
assign n_46690 = ~n_16985 &  n_46689;
assign n_46691 = ~n_16979 &  n_46690;
assign n_46692 = ~n_16973 &  n_46691;
assign n_46693 = ~n_16967 &  n_46692;
assign n_46694 = ~n_16961 &  n_46693;
assign n_46695 = ~n_16955 &  n_46694;
assign n_46696 = ~n_16949 &  n_46695;
assign n_46697 = ~n_16943 &  n_46696;
assign n_46698 = ~n_16937 &  n_46697;
assign n_46699 = ~n_16931 &  n_46698;
assign n_46700 = ~n_16925 &  n_46699;
assign n_46701 = ~n_16919 &  n_46700;
assign n_46702 = ~n_16913 &  n_46701;
assign n_46703 = ~n_16907 &  n_46702;
assign n_46704 = ~n_16901 &  n_46703;
assign n_46705 = ~n_16895 &  n_46704;
assign n_46706 = ~n_16889 &  n_46705;
assign n_46707 = ~n_16881 &  n_46706;
assign n_46708 = ~n_16875 &  n_46707;
assign n_46709 = ~n_16869 &  n_46708;
assign n_46710 = ~n_16863 &  n_46709;
assign n_46711 = ~n_16857 &  n_46710;
assign n_46712 = ~n_16851 &  n_46711;
assign n_46713 = ~n_16845 &  n_46712;
assign n_46714 = ~n_16839 &  n_46713;
assign n_46715 = ~n_16833 &  n_46714;
assign n_46716 = ~n_16827 &  n_46715;
assign n_46717 = ~n_16821 &  n_46716;
assign n_46718 = ~n_16815 &  n_46717;
assign n_46719 = ~n_16809 &  n_46718;
assign n_46720 = ~n_16803 &  n_46719;
assign n_46721 = ~n_16797 &  n_46720;
assign n_46722 = ~n_16791 &  n_46721;
assign n_46723 = ~n_16785 &  n_46722;
assign n_46724 = ~n_16779 &  n_46723;
assign n_46725 = ~n_16773 &  n_46724;
assign n_46726 = ~n_16767 &  n_46725;
assign n_46727 = ~n_16761 &  n_46726;
assign n_46728 = ~n_16755 &  n_46727;
assign n_46729 = ~n_16749 &  n_46728;
assign n_46730 = ~n_16743 &  n_46729;
assign n_46731 = ~n_16737 &  n_46730;
assign n_46732 = ~n_16731 &  n_46731;
assign n_46733 = ~n_16725 &  n_46732;
assign n_46734 = ~n_16719 &  n_46733;
assign n_46735 = ~n_16713 &  n_46734;
assign n_46736 = ~n_16707 &  n_46735;
assign n_46737 = ~n_16701 &  n_46736;
assign n_46738 = ~n_16695 &  n_46737;
assign n_46739 = ~n_16688 &  n_46738;
assign n_46740 = ~n_16682 &  n_46739;
assign n_46741 = ~n_16676 &  n_46740;
assign n_46742 = ~n_16670 &  n_46741;
assign n_46743 = ~n_16664 &  n_46742;
assign n_46744 = ~n_16658 &  n_46743;
assign n_46745 = ~n_16652 &  n_46744;
assign n_46746 = ~n_16646 &  n_46745;
assign n_46747 = ~n_16640 &  n_46746;
assign n_46748 = ~n_16634 &  n_46747;
assign n_46749 = ~n_16628 &  n_46748;
assign n_46750 = ~n_16622 &  n_46749;
assign n_46751 = ~n_16616 &  n_46750;
assign n_46752 = ~n_16610 &  n_46751;
assign n_46753 = ~n_16604 &  n_46752;
assign n_46754 = ~n_16598 &  n_46753;
assign n_46755 = ~n_16592 &  n_46754;
assign n_46756 = ~n_16586 &  n_46755;
assign n_46757 = ~n_16580 &  n_46756;
assign n_46758 = ~n_16574 &  n_46757;
assign n_46759 = ~n_16568 &  n_46758;
assign n_46760 = ~n_16562 &  n_46759;
assign n_46761 = ~n_16556 &  n_46760;
assign n_46762 = ~n_16550 &  n_46761;
assign n_46763 = ~n_16544 &  n_46762;
assign n_46764 = ~n_16538 &  n_46763;
assign n_46765 = ~n_16532 &  n_46764;
assign n_46766 = ~n_16526 &  n_46765;
assign n_46767 = ~n_16520 &  n_46766;
assign n_46768 = ~n_16514 &  n_46767;
assign n_46769 = ~n_16508 &  n_46768;
assign n_46770 = ~n_16502 &  n_46769;
assign n_46771 = ~n_16494 &  n_46770;
assign n_46772 = ~n_16488 &  n_46771;
assign n_46773 = ~n_16482 &  n_46772;
assign n_46774 = ~n_16476 &  n_46773;
assign n_46775 = ~n_16470 &  n_46774;
assign n_46776 = ~n_16464 &  n_46775;
assign n_46777 = ~n_16458 &  n_46776;
assign n_46778 = ~n_16452 &  n_46777;
assign n_46779 = ~n_16446 &  n_46778;
assign n_46780 = ~n_16440 &  n_46779;
assign n_46781 = ~n_16434 &  n_46780;
assign n_46782 = ~n_16428 &  n_46781;
assign n_46783 = ~n_16422 &  n_46782;
assign n_46784 = ~n_16416 &  n_46783;
assign n_46785 = ~n_16410 &  n_46784;
assign n_46786 = ~n_16404 &  n_46785;
assign n_46787 = ~n_16398 &  n_46786;
assign n_46788 = ~n_16392 &  n_46787;
assign n_46789 = ~n_16386 &  n_46788;
assign n_46790 = ~n_16380 &  n_46789;
assign n_46791 = ~n_16374 &  n_46790;
assign n_46792 = ~n_16368 &  n_46791;
assign n_46793 = ~n_16362 &  n_46792;
assign n_46794 = ~n_16356 &  n_46793;
assign n_46795 = ~n_16350 &  n_46794;
assign n_46796 = ~n_16344 &  n_46795;
assign n_46797 = ~n_16338 &  n_46796;
assign n_46798 = ~n_16332 &  n_46797;
assign n_46799 = ~n_16326 &  n_46798;
assign n_46800 = ~n_16320 &  n_46799;
assign n_46801 = ~n_16314 &  n_46800;
assign n_46802 = ~n_16308 &  n_46801;
assign n_46803 = ~n_16301 &  n_46802;
assign n_46804 = ~n_16297 &  n_46803;
assign n_46805 = ~n_16291 &  n_46804;
assign n_46806 = ~n_16285 &  n_46805;
assign n_46807 = ~n_16279 &  n_46806;
assign n_46808 = ~n_16273 &  n_46807;
assign n_46809 = ~n_16267 &  n_46808;
assign n_46810 = ~n_16261 &  n_46809;
assign n_46811 = ~n_16255 &  n_46810;
assign n_46812 = ~n_16249 &  n_46811;
assign n_46813 = ~n_16243 &  n_46812;
assign n_46814 = ~n_16237 &  n_46813;
assign n_46815 = ~n_16231 &  n_46814;
assign n_46816 = ~n_16225 &  n_46815;
assign n_46817 = ~n_16219 &  n_46816;
assign n_46818 = ~n_16213 &  n_46817;
assign n_46819 = ~n_16207 &  n_46818;
assign n_46820 = ~n_16201 &  n_46819;
assign n_46821 = ~n_16195 &  n_46820;
assign n_46822 = ~n_16189 &  n_46821;
assign n_46823 = ~n_16183 &  n_46822;
assign n_46824 = ~n_16177 &  n_46823;
assign n_46825 = ~n_16171 &  n_46824;
assign n_46826 = ~n_16165 &  n_46825;
assign n_46827 = ~n_16159 &  n_46826;
assign n_46828 = ~n_16153 &  n_46827;
assign n_46829 = ~n_16147 &  n_46828;
assign n_46830 = ~n_16141 &  n_46829;
assign n_46831 = ~n_16135 &  n_46830;
assign n_46832 = ~n_16129 &  n_46831;
assign n_46833 = ~n_16123 &  n_46832;
assign n_46834 = ~n_16117 &  n_46833;
assign n_46835 = ~n_16109 &  n_46834;
assign n_46836 = ~n_16105 &  n_46835;
assign n_46837 = ~n_16099 &  n_46836;
assign n_46838 = ~n_16093 &  n_46837;
assign n_46839 = ~n_16087 &  n_46838;
assign n_46840 = ~n_16081 &  n_46839;
assign n_46841 = ~n_16075 &  n_46840;
assign n_46842 = ~n_16069 &  n_46841;
assign n_46843 = ~n_16063 &  n_46842;
assign n_46844 = ~n_16057 &  n_46843;
assign n_46845 = ~n_16051 &  n_46844;
assign n_46846 = ~n_16045 &  n_46845;
assign n_46847 = ~n_16039 &  n_46846;
assign n_46848 = ~n_16033 &  n_46847;
assign n_46849 = ~n_16027 &  n_46848;
assign n_46850 = ~n_16021 &  n_46849;
assign n_46851 = ~n_16015 &  n_46850;
assign n_46852 = ~n_16009 &  n_46851;
assign n_46853 = ~n_16003 &  n_46852;
assign n_46854 = ~n_15997 &  n_46853;
assign n_46855 = ~n_15991 &  n_46854;
assign n_46856 = ~n_15985 &  n_46855;
assign n_46857 = ~n_15979 &  n_46856;
assign n_46858 = ~n_15973 &  n_46857;
assign n_46859 = ~n_15967 &  n_46858;
assign n_46860 = ~n_15961 &  n_46859;
assign n_46861 = ~n_15955 &  n_46860;
assign n_46862 = ~n_15949 &  n_46861;
assign n_46863 = ~n_15943 &  n_46862;
assign n_46864 = ~n_15937 &  n_46863;
assign n_46865 = ~n_15931 &  n_46864;
assign n_46866 = ~n_15925 &  n_46865;
assign n_46867 = ~n_15915 &  n_46866;
assign n_46868 = ~n_15896 &  n_46867;
assign n_46869 = ~n_15879 &  n_46868;
assign n_46870 = ~n_15862 &  n_46869;
assign n_46871 = ~n_15845 &  n_46870;
assign n_46872 = ~n_15828 &  n_46871;
assign n_46873 = ~n_15811 &  n_46872;
assign n_46874 = ~n_15794 &  n_46873;
assign n_46875 = ~n_15777 &  n_46874;
assign n_46876 = ~n_15760 &  n_46875;
assign n_46877 = ~n_15743 &  n_46876;
assign n_46878 = ~n_15726 &  n_46877;
assign n_46879 = ~n_15709 &  n_46878;
assign n_46880 = ~n_15692 &  n_46879;
assign n_46881 = ~n_15675 &  n_46880;
assign n_46882 = ~n_15658 &  n_46881;
assign n_46883 = ~n_15641 &  n_46882;
assign n_46884 = ~n_15624 &  n_46883;
assign n_46885 = ~n_15607 &  n_46884;
assign n_46886 = ~n_15590 &  n_46885;
assign n_46887 = ~n_15573 &  n_46886;
assign n_46888 = ~n_15556 &  n_46887;
assign n_46889 = ~n_15539 &  n_46888;
assign n_46890 = ~n_15522 &  n_46889;
assign n_46891 = ~n_15505 &  n_46890;
assign n_46892 = ~n_15488 &  n_46891;
assign n_46893 = ~n_15471 &  n_46892;
assign n_46894 = ~n_15454 &  n_46893;
assign n_46895 = ~n_15437 &  n_46894;
assign n_46896 = ~n_15420 &  n_46895;
assign n_46897 = ~n_15403 &  n_46896;
assign n_46898 = ~n_15386 &  n_46897;
assign n_46899 = ~n_15365 &  n_46898;
assign n_46900 = ~n_15347 &  n_46899;
assign n_46901 = ~n_15329 &  n_46900;
assign n_46902 = ~n_15311 &  n_46901;
assign n_46903 = ~n_15293 &  n_46902;
assign n_46904 = ~n_15275 &  n_46903;
assign n_46905 = ~n_15257 &  n_46904;
assign n_46906 = ~n_15239 &  n_46905;
assign n_46907 = ~n_15221 &  n_46906;
assign n_46908 = ~n_15203 &  n_46907;
assign n_46909 = ~n_15185 &  n_46908;
assign n_46910 = ~n_15167 &  n_46909;
assign n_46911 = ~n_15149 &  n_46910;
assign n_46912 = ~n_15131 &  n_46911;
assign n_46913 = ~n_15113 &  n_46912;
assign n_46914 = ~n_15095 &  n_46913;
assign n_46915 = ~n_15077 &  n_46914;
assign n_46916 = ~n_15059 &  n_46915;
assign n_46917 = ~n_15041 &  n_46916;
assign n_46918 = ~n_15023 &  n_46917;
assign n_46919 = ~n_15005 &  n_46918;
assign n_46920 = ~n_14987 &  n_46919;
assign n_46921 = ~n_14969 &  n_46920;
assign n_46922 = ~n_14951 &  n_46921;
assign n_46923 = ~n_14933 &  n_46922;
assign n_46924 = ~n_14915 &  n_46923;
assign n_46925 = ~n_14897 &  n_46924;
assign n_46926 = ~n_14879 &  n_46925;
assign n_46927 = ~n_14861 &  n_46926;
assign n_46928 = ~n_14843 &  n_46927;
assign n_46929 = ~n_14825 &  n_46928;
assign n_46930 = ~n_14807 &  n_46929;
assign n_46931 = ~n_14784 &  n_46930;
assign n_46932 = ~n_14780 &  n_46931;
assign n_46933 = ~n_14776 &  n_46932;
assign n_46934 = ~n_14772 &  n_46933;
assign n_46935 = ~n_14768 &  n_46934;
assign n_46936 = ~n_14764 &  n_46935;
assign n_46937 = ~n_14760 &  n_46936;
assign n_46938 = ~n_14756 &  n_46937;
assign n_46939 = ~n_14752 &  n_46938;
assign n_46940 = ~n_14748 &  n_46939;
assign n_46941 = ~n_14744 &  n_46940;
assign n_46942 = ~n_14740 &  n_46941;
assign n_46943 = ~n_14736 &  n_46942;
assign n_46944 = ~n_14732 &  n_46943;
assign n_46945 = ~n_14728 &  n_46944;
assign n_46946 = ~n_14724 &  n_46945;
assign n_46947 = ~n_14720 &  n_46946;
assign n_46948 = ~n_14716 &  n_46947;
assign n_46949 = ~n_14712 &  n_46948;
assign n_46950 = ~n_14708 &  n_46949;
assign n_46951 = ~n_14704 &  n_46950;
assign n_46952 = ~n_14700 &  n_46951;
assign n_46953 = ~n_14696 &  n_46952;
assign n_46954 = ~n_14692 &  n_46953;
assign n_46955 = ~n_14688 &  n_46954;
assign n_46956 = ~n_14684 &  n_46955;
assign n_46957 = ~n_14680 &  n_46956;
assign n_46958 = ~n_14676 &  n_46957;
assign n_46959 = ~n_14672 &  n_46958;
assign n_46960 = ~n_14668 &  n_46959;
assign n_46961 = ~n_14664 &  n_46960;
assign n_46962 = ~n_14660 &  n_46961;
assign n_46963 = ~n_14654 &  n_46962;
assign n_46964 = ~n_14642 &  n_46963;
assign n_46965 = ~n_14630 &  n_46964;
assign n_46966 = ~n_14618 &  n_46965;
assign n_46967 = ~n_14606 &  n_46966;
assign n_46968 = ~n_14594 &  n_46967;
assign n_46969 = ~n_14582 &  n_46968;
assign n_46970 = ~n_14570 &  n_46969;
assign n_46971 = ~n_14558 &  n_46970;
assign n_46972 = ~n_14546 &  n_46971;
assign n_46973 = ~n_14534 &  n_46972;
assign n_46974 = ~n_14522 &  n_46973;
assign n_46975 = ~n_14510 &  n_46974;
assign n_46976 = ~n_14498 &  n_46975;
assign n_46977 = ~n_14486 &  n_46976;
assign n_46978 = ~n_14474 &  n_46977;
assign n_46979 = ~n_14462 &  n_46978;
assign n_46980 = ~n_14450 &  n_46979;
assign n_46981 = ~n_14438 &  n_46980;
assign n_46982 = ~n_14426 &  n_46981;
assign n_46983 = ~n_14414 &  n_46982;
assign n_46984 = ~n_14402 &  n_46983;
assign n_46985 = ~n_14390 &  n_46984;
assign n_46986 = ~n_14378 &  n_46985;
assign n_46987 = ~n_14366 &  n_46986;
assign n_46988 = ~n_14354 &  n_46987;
assign n_46989 = ~n_14342 &  n_46988;
assign n_46990 = ~n_14330 &  n_46989;
assign n_46991 = ~n_14318 &  n_46990;
assign n_46992 = ~n_14306 &  n_46991;
assign n_46993 = ~n_14294 &  n_46992;
assign n_46994 = ~n_14282 &  n_46993;
assign n_46995 = ~n_14259 &  n_46994;
assign n_46996 = ~n_14247 &  n_46995;
assign n_46997 = ~n_14235 &  n_46996;
assign n_46998 = ~n_14223 &  n_46997;
assign n_46999 = ~n_14211 &  n_46998;
assign n_47000 = ~n_14199 &  n_46999;
assign n_47001 = ~n_14187 &  n_47000;
assign n_47002 = ~n_14175 &  n_47001;
assign n_47003 = ~n_14163 &  n_47002;
assign n_47004 = ~n_14151 &  n_47003;
assign n_47005 = ~n_14139 &  n_47004;
assign n_47006 = ~n_14127 &  n_47005;
assign n_47007 = ~n_14115 &  n_47006;
assign n_47008 = ~n_14103 &  n_47007;
assign n_47009 = ~n_14091 &  n_47008;
assign n_47010 = ~n_14079 &  n_47009;
assign n_47011 = ~n_14067 &  n_47010;
assign n_47012 = ~n_14055 &  n_47011;
assign n_47013 = ~n_14043 &  n_47012;
assign n_47014 = ~n_14031 &  n_47013;
assign n_47015 = ~n_14019 &  n_47014;
assign n_47016 = ~n_14007 &  n_47015;
assign n_47017 = ~n_13995 &  n_47016;
assign n_47018 = ~n_13983 &  n_47017;
assign n_47019 = ~n_13971 &  n_47018;
assign n_47020 = ~n_13959 &  n_47019;
assign n_47021 = ~n_13947 &  n_47020;
assign n_47022 = ~n_13935 &  n_47021;
assign n_47023 = ~n_13923 &  n_47022;
assign n_47024 = ~n_13911 &  n_47023;
assign n_47025 = ~n_13899 &  n_47024;
assign n_47026 = ~n_13887 &  n_47025;
assign n_47027 = ~n_13865 &  n_47026;
assign n_47028 = ~n_13859 &  n_47027;
assign n_47029 = ~n_13853 &  n_47028;
assign n_47030 = ~n_13847 &  n_47029;
assign n_47031 = ~n_13841 &  n_47030;
assign n_47032 = ~n_13835 &  n_47031;
assign n_47033 = ~n_13829 &  n_47032;
assign n_47034 = ~n_13823 &  n_47033;
assign n_47035 = ~n_13817 &  n_47034;
assign n_47036 = ~n_13811 &  n_47035;
assign n_47037 = ~n_13805 &  n_47036;
assign n_47038 = ~n_13799 &  n_47037;
assign n_47039 = ~n_13793 &  n_47038;
assign n_47040 = ~n_13787 &  n_47039;
assign n_47041 = ~n_13781 &  n_47040;
assign n_47042 = ~n_13775 &  n_47041;
assign n_47043 = ~n_13769 &  n_47042;
assign n_47044 = ~n_13763 &  n_47043;
assign n_47045 = ~n_13757 &  n_47044;
assign n_47046 = ~n_13751 &  n_47045;
assign n_47047 = ~n_13745 &  n_47046;
assign n_47048 = ~n_13739 &  n_47047;
assign n_47049 = ~n_13733 &  n_47048;
assign n_47050 = ~n_13727 &  n_47049;
assign n_47051 = ~n_13721 &  n_47050;
assign n_47052 = ~n_13715 &  n_47051;
assign n_47053 = ~n_13709 &  n_47052;
assign n_47054 = ~n_13703 &  n_47053;
assign n_47055 = ~n_13697 &  n_47054;
assign n_47056 = ~n_13691 &  n_47055;
assign n_47057 = ~n_13685 &  n_47056;
assign n_47058 = ~n_13679 &  n_47057;
assign n_47059 = ~n_13671 &  n_47058;
assign n_47060 = ~n_13665 &  n_47059;
assign n_47061 = ~n_13659 &  n_47060;
assign n_47062 = ~n_13653 &  n_47061;
assign n_47063 = ~n_13647 &  n_47062;
assign n_47064 = ~n_13641 &  n_47063;
assign n_47065 = ~n_13635 &  n_47064;
assign n_47066 = ~n_13629 &  n_47065;
assign n_47067 = ~n_13623 &  n_47066;
assign n_47068 = ~n_13617 &  n_47067;
assign n_47069 = ~n_13611 &  n_47068;
assign n_47070 = ~n_13605 &  n_47069;
assign n_47071 = ~n_13599 &  n_47070;
assign n_47072 = ~n_13593 &  n_47071;
assign n_47073 = ~n_13587 &  n_47072;
assign n_47074 = ~n_13581 &  n_47073;
assign n_47075 = ~n_13575 &  n_47074;
assign n_47076 = ~n_13569 &  n_47075;
assign n_47077 = ~n_13563 &  n_47076;
assign n_47078 = ~n_13557 &  n_47077;
assign n_47079 = ~n_13551 &  n_47078;
assign n_47080 = ~n_13545 &  n_47079;
assign n_47081 = ~n_13539 &  n_47080;
assign n_47082 = ~n_13533 &  n_47081;
assign n_47083 = ~n_13527 &  n_47082;
assign n_47084 = ~n_13521 &  n_47083;
assign n_47085 = ~n_13515 &  n_47084;
assign n_47086 = ~n_13509 &  n_47085;
assign n_47087 = ~n_13503 &  n_47086;
assign n_47088 = ~n_13497 &  n_47087;
assign n_47089 = ~n_13491 &  n_47088;
assign n_47090 = ~n_13485 &  n_47089;
assign n_47091 = ~n_13478 &  n_47090;
assign n_47092 = ~n_13472 &  n_47091;
assign n_47093 = ~n_13466 &  n_47092;
assign n_47094 = ~n_13460 &  n_47093;
assign n_47095 = ~n_13454 &  n_47094;
assign n_47096 = ~n_13448 &  n_47095;
assign n_47097 = ~n_13442 &  n_47096;
assign n_47098 = ~n_13436 &  n_47097;
assign n_47099 = ~n_13430 &  n_47098;
assign n_47100 = ~n_13424 &  n_47099;
assign n_47101 = ~n_13418 &  n_47100;
assign n_47102 = ~n_13412 &  n_47101;
assign n_47103 = ~n_13406 &  n_47102;
assign n_47104 = ~n_13400 &  n_47103;
assign n_47105 = ~n_13394 &  n_47104;
assign n_47106 = ~n_13388 &  n_47105;
assign n_47107 = ~n_13382 &  n_47106;
assign n_47108 = ~n_13376 &  n_47107;
assign n_47109 = ~n_13370 &  n_47108;
assign n_47110 = ~n_13364 &  n_47109;
assign n_47111 = ~n_13358 &  n_47110;
assign n_47112 = ~n_13352 &  n_47111;
assign n_47113 = ~n_13346 &  n_47112;
assign n_47114 = ~n_13340 &  n_47113;
assign n_47115 = ~n_13334 &  n_47114;
assign n_47116 = ~n_13328 &  n_47115;
assign n_47117 = ~n_13322 &  n_47116;
assign n_47118 = ~n_13316 &  n_47117;
assign n_47119 = ~n_13310 &  n_47118;
assign n_47120 = ~n_13304 &  n_47119;
assign n_47121 = ~n_13298 &  n_47120;
assign n_47122 = ~n_13292 &  n_47121;
assign n_47123 = ~n_13285 &  n_47122;
assign n_47124 = ~n_13279 &  n_47123;
assign n_47125 = ~n_13273 &  n_47124;
assign n_47126 = ~n_13267 &  n_47125;
assign n_47127 = ~n_13261 &  n_47126;
assign n_47128 = ~n_13255 &  n_47127;
assign n_47129 = ~n_13249 &  n_47128;
assign n_47130 = ~n_13243 &  n_47129;
assign n_47131 = ~n_13237 &  n_47130;
assign n_47132 = ~n_13229 &  n_47131;
assign n_47133 = ~n_13212 &  n_47132;
assign n_47134 = ~n_13195 &  n_47133;
assign n_47135 = ~n_13178 &  n_47134;
assign n_47136 = ~n_13161 &  n_47135;
assign n_47137 = ~n_13103 &  n_47136;
assign n_47138 = ~n_13097 &  n_47137;
assign n_47139 = ~n_13091 &  n_47138;
assign n_47140 = ~n_13085 &  n_47139;
assign n_47141 = ~n_13079 &  n_47140;
assign n_47142 = ~n_13073 &  n_47141;
assign n_47143 = ~n_13067 &  n_47142;
assign n_47144 = ~n_13061 &  n_47143;
assign n_47145 = ~n_13055 &  n_47144;
assign n_47146 = ~n_13049 &  n_47145;
assign n_47147 = ~n_13043 &  n_47146;
assign n_47148 = ~n_13037 &  n_47147;
assign n_47149 = ~n_13031 &  n_47148;
assign n_47150 = ~n_13025 &  n_47149;
assign n_47151 = ~n_13019 &  n_47150;
assign n_47152 = ~n_13013 &  n_47151;
assign n_47153 = ~n_13007 &  n_47152;
assign n_47154 = ~n_13001 &  n_47153;
assign n_47155 = ~n_12995 &  n_47154;
assign n_47156 = ~n_12989 &  n_47155;
assign n_47157 = ~n_12983 &  n_47156;
assign n_47158 = ~n_12977 &  n_47157;
assign n_47159 = ~n_12971 &  n_47158;
assign n_47160 = ~n_12965 &  n_47159;
assign n_47161 = ~n_12959 &  n_47160;
assign n_47162 = ~n_12953 &  n_47161;
assign n_47163 = ~n_12947 &  n_47162;
assign n_47164 = ~n_12941 &  n_47163;
assign n_47165 = ~n_12935 &  n_47164;
assign n_47166 = ~n_12929 &  n_47165;
assign n_47167 = ~n_12923 &  n_47166;
assign n_47168 = ~n_12917 &  n_47167;
assign n_47169 = ~n_12908 &  n_47168;
assign n_47170 = ~n_12890 &  n_47169;
assign n_47171 = ~n_12872 &  n_47170;
assign n_47172 = ~n_12854 &  n_47171;
assign n_47173 = ~n_12836 &  n_47172;
assign n_47174 = ~n_12818 &  n_47173;
assign n_47175 = ~n_12800 &  n_47174;
assign n_47176 = ~n_12782 &  n_47175;
assign n_47177 = ~n_12764 &  n_47176;
assign n_47178 = ~n_12746 &  n_47177;
assign n_47179 = ~n_12728 &  n_47178;
assign n_47180 = ~n_12710 &  n_47179;
assign n_47181 = ~n_12692 &  n_47180;
assign n_47182 = ~n_12674 &  n_47181;
assign n_47183 = ~n_12656 &  n_47182;
assign n_47184 = ~n_12638 &  n_47183;
assign n_47185 = ~n_12620 &  n_47184;
assign n_47186 = ~n_12602 &  n_47185;
assign n_47187 = ~n_12584 &  n_47186;
assign n_47188 = ~n_12566 &  n_47187;
assign n_47189 = ~n_12548 &  n_47188;
assign n_47190 = ~n_12530 &  n_47189;
assign n_47191 = ~n_12512 &  n_47190;
assign n_47192 = ~n_12494 &  n_47191;
assign n_47193 = ~n_12476 &  n_47192;
assign n_47194 = ~n_12458 &  n_47193;
assign n_47195 = ~n_12440 &  n_47194;
assign n_47196 = ~n_12422 &  n_47195;
assign n_47197 = ~n_12404 &  n_47196;
assign n_47198 = ~n_12386 &  n_47197;
assign n_47199 = ~n_12368 &  n_47198;
assign n_47200 = ~n_12350 &  n_47199;
assign n_47201 = ~n_12291 &  n_47200;
assign n_47202 = ~n_12249 &  n_47201;
assign n_47203 = ~n_12204 &  n_47202;
assign n_47204 = ~n_12159 &  n_47203;
assign n_47205 = ~n_12114 &  n_47204;
assign n_47206 = ~n_12069 &  n_47205;
assign n_47207 = ~n_12024 &  n_47206;
assign n_47208 = ~n_11979 &  n_47207;
assign n_47209 = ~n_11934 &  n_47208;
assign n_47210 = ~n_11889 &  n_47209;
assign n_47211 = ~n_11844 &  n_47210;
assign n_47212 = ~n_11799 &  n_47211;
assign n_47213 = ~n_11754 &  n_47212;
assign n_47214 = ~n_11709 &  n_47213;
assign n_47215 = ~n_11664 &  n_47214;
assign n_47216 = ~n_11619 &  n_47215;
assign n_47217 = ~n_11574 &  n_47216;
assign n_47218 = ~n_11529 &  n_47217;
assign n_47219 = ~n_11484 &  n_47218;
assign n_47220 = ~n_11439 &  n_47219;
assign n_47221 = ~n_11394 &  n_47220;
assign n_47222 = ~n_11349 &  n_47221;
assign n_47223 = ~n_11304 &  n_47222;
assign n_47224 = ~n_11259 &  n_47223;
assign n_47225 = ~n_11214 &  n_47224;
assign n_47226 = ~n_11169 &  n_47225;
assign n_47227 = ~n_11124 &  n_47226;
assign n_47228 = ~n_11079 &  n_47227;
assign n_47229 = ~n_11034 &  n_47228;
assign n_47230 = ~n_10988 &  n_47229;
assign n_47231 = ~n_10938 &  n_47230;
assign n_47232 = ~n_10899 &  n_47231;
assign n_47233 = ~n_10866 &  n_47232;
assign n_47234 = ~n_10854 &  n_47233;
assign n_47235 = ~n_10842 &  n_47234;
assign n_47236 = ~n_10830 &  n_47235;
assign n_47237 = ~n_10818 &  n_47236;
assign n_47238 = ~n_10806 &  n_47237;
assign n_47239 = ~n_10794 &  n_47238;
assign n_47240 = ~n_10782 &  n_47239;
assign n_47241 = ~n_10770 &  n_47240;
assign n_47242 = ~n_10758 &  n_47241;
assign n_47243 = ~n_10746 &  n_47242;
assign n_47244 = ~n_10734 &  n_47243;
assign n_47245 = ~n_10722 &  n_47244;
assign n_47246 = ~n_10710 &  n_47245;
assign n_47247 = ~n_10698 &  n_47246;
assign n_47248 = ~n_10686 &  n_47247;
assign n_47249 = ~n_10674 &  n_47248;
assign n_47250 = ~n_10662 &  n_47249;
assign n_47251 = ~n_10650 &  n_47250;
assign n_47252 = ~n_10638 &  n_47251;
assign n_47253 = ~n_10626 &  n_47252;
assign n_47254 = ~n_10614 &  n_47253;
assign n_47255 = ~n_10602 &  n_47254;
assign n_47256 = ~n_10590 &  n_47255;
assign n_47257 = ~n_10578 &  n_47256;
assign n_47258 = ~n_10566 &  n_47257;
assign n_47259 = ~n_10554 &  n_47258;
assign n_47260 = ~n_10542 &  n_47259;
assign n_47261 = ~n_10530 &  n_47260;
assign n_47262 = ~n_10518 &  n_47261;
assign n_47263 = ~n_10506 &  n_47262;
assign n_47264 = ~n_10494 &  n_47263;
assign n_47265 = ~n_10469 &  n_47264;
assign n_47266 = ~n_10463 &  n_47265;
assign n_47267 = ~n_10457 &  n_47266;
assign n_47268 = ~n_10451 &  n_47267;
assign n_47269 = ~n_10445 &  n_47268;
assign n_47270 = ~n_10439 &  n_47269;
assign n_47271 = ~n_10433 &  n_47270;
assign n_47272 = ~n_10427 &  n_47271;
assign n_47273 = ~n_10421 &  n_47272;
assign n_47274 = ~n_10415 &  n_47273;
assign n_47275 = ~n_10409 &  n_47274;
assign n_47276 = ~n_10403 &  n_47275;
assign n_47277 = ~n_10397 &  n_47276;
assign n_47278 = ~n_10391 &  n_47277;
assign n_47279 = ~n_10385 &  n_47278;
assign n_47280 = ~n_10379 &  n_47279;
assign n_47281 = ~n_10373 &  n_47280;
assign n_47282 = ~n_10367 &  n_47281;
assign n_47283 = ~n_10361 &  n_47282;
assign n_47284 = ~n_10355 &  n_47283;
assign n_47285 = ~n_10349 &  n_47284;
assign n_47286 = ~n_10343 &  n_47285;
assign n_47287 = ~n_10337 &  n_47286;
assign n_47288 = ~n_10331 &  n_47287;
assign n_47289 = ~n_10325 &  n_47288;
assign n_47290 = ~n_10319 &  n_47289;
assign n_47291 = ~n_10313 &  n_47290;
assign n_47292 = ~n_10307 &  n_47291;
assign n_47293 = ~n_10301 &  n_47292;
assign n_47294 = ~n_10295 &  n_47293;
assign n_47295 = ~n_10289 &  n_47294;
assign n_47296 = ~n_10283 &  n_47295;
assign n_47297 = ~n_10273 &  n_47296;
assign n_47298 = ~n_10267 &  n_47297;
assign n_47299 = ~n_10261 &  n_47298;
assign n_47300 = ~n_10255 &  n_47299;
assign n_47301 = ~n_10249 &  n_47300;
assign n_47302 = ~n_10243 &  n_47301;
assign n_47303 = ~n_10237 &  n_47302;
assign n_47304 = ~n_10231 &  n_47303;
assign n_47305 = ~n_10225 &  n_47304;
assign n_47306 = ~n_10219 &  n_47305;
assign n_47307 = ~n_10213 &  n_47306;
assign n_47308 = ~n_10207 &  n_47307;
assign n_47309 = ~n_10201 &  n_47308;
assign n_47310 = ~n_10195 &  n_47309;
assign n_47311 = ~n_10189 &  n_47310;
assign n_47312 = ~n_10183 &  n_47311;
assign n_47313 = ~n_10177 &  n_47312;
assign n_47314 = ~n_10171 &  n_47313;
assign n_47315 = ~n_10165 &  n_47314;
assign n_47316 = ~n_10159 &  n_47315;
assign n_47317 = ~n_10153 &  n_47316;
assign n_47318 = ~n_10147 &  n_47317;
assign n_47319 = ~n_10141 &  n_47318;
assign n_47320 = ~n_10135 &  n_47319;
assign n_47321 = ~n_10129 &  n_47320;
assign n_47322 = ~n_10123 &  n_47321;
assign n_47323 = ~n_10117 &  n_47322;
assign n_47324 = ~n_10111 &  n_47323;
assign n_47325 = ~n_10105 &  n_47324;
assign n_47326 = ~n_10099 &  n_47325;
assign n_47327 = ~n_10093 &  n_47326;
assign n_47328 = ~n_10087 &  n_47327;
assign n_47329 = ~n_10077 &  n_47328;
assign n_47330 = ~n_10071 &  n_47329;
assign n_47331 = ~n_10065 &  n_47330;
assign n_47332 = ~n_10059 &  n_47331;
assign n_47333 = ~n_10053 &  n_47332;
assign n_47334 = ~n_10047 &  n_47333;
assign n_47335 = ~n_10041 &  n_47334;
assign n_47336 = ~n_10035 &  n_47335;
assign n_47337 = ~n_10029 &  n_47336;
assign n_47338 = ~n_10023 &  n_47337;
assign n_47339 = ~n_10017 &  n_47338;
assign n_47340 = ~n_10011 &  n_47339;
assign n_47341 = ~n_10005 &  n_47340;
assign n_47342 = ~n_9999 &  n_47341;
assign n_47343 = ~n_9993 &  n_47342;
assign n_47344 = ~n_9987 &  n_47343;
assign n_47345 = ~n_9981 &  n_47344;
assign n_47346 = ~n_9975 &  n_47345;
assign n_47347 = ~n_9969 &  n_47346;
assign n_47348 = ~n_9963 &  n_47347;
assign n_47349 = ~n_9957 &  n_47348;
assign n_47350 = ~n_9951 &  n_47349;
assign n_47351 = ~n_9945 &  n_47350;
assign n_47352 = ~n_9939 &  n_47351;
assign n_47353 = ~n_9933 &  n_47352;
assign n_47354 = ~n_9927 &  n_47353;
assign n_47355 = ~n_9921 &  n_47354;
assign n_47356 = ~n_9915 &  n_47355;
assign n_47357 = ~n_9909 &  n_47356;
assign n_47358 = ~n_9903 &  n_47357;
assign n_47359 = ~n_9897 &  n_47358;
assign n_47360 = ~n_9891 &  n_47359;
assign n_47361 = ~n_9883 &  n_47360;
assign n_47362 = ~n_9877 &  n_47361;
assign n_47363 = ~n_9871 &  n_47362;
assign n_47364 = ~n_9865 &  n_47363;
assign n_47365 = ~n_9859 &  n_47364;
assign n_47366 = ~n_9853 &  n_47365;
assign n_47367 = ~n_9847 &  n_47366;
assign n_47368 = ~n_9841 &  n_47367;
assign n_47369 = ~n_9835 &  n_47368;
assign n_47370 = ~n_9829 &  n_47369;
assign n_47371 = ~n_9823 &  n_47370;
assign n_47372 = ~n_9817 &  n_47371;
assign n_47373 = ~n_9811 &  n_47372;
assign n_47374 = ~n_9805 &  n_47373;
assign n_47375 = ~n_9799 &  n_47374;
assign n_47376 = ~n_9793 &  n_47375;
assign n_47377 = ~n_9787 &  n_47376;
assign n_47378 = ~n_9781 &  n_47377;
assign n_47379 = ~n_9775 &  n_47378;
assign n_47380 = ~n_9769 &  n_47379;
assign n_47381 = ~n_9763 &  n_47380;
assign n_47382 = ~n_9757 &  n_47381;
assign n_47383 = ~n_9751 &  n_47382;
assign n_47384 = ~n_9745 &  n_47383;
assign n_47385 = ~n_9739 &  n_47384;
assign n_47386 = ~n_9733 &  n_47385;
assign n_47387 = ~n_9727 &  n_47386;
assign n_47388 = ~n_9721 &  n_47387;
assign n_47389 = ~n_9715 &  n_47388;
assign n_47390 = ~n_9709 &  n_47389;
assign n_47391 = ~n_9703 &  n_47390;
assign n_47392 = ~n_9697 &  n_47391;
assign n_47393 = ~n_9688 &  n_47392;
assign n_47394 = ~n_9680 &  n_47393;
assign n_47395 = ~n_9672 &  n_47394;
assign n_47396 = ~n_9664 &  n_47395;
assign n_47397 = ~n_9656 &  n_47396;
assign n_47398 = ~n_9648 &  n_47397;
assign n_47399 = ~n_9640 &  n_47398;
assign n_47400 = ~n_9632 &  n_47399;
assign n_47401 = ~n_9624 &  n_47400;
assign n_47402 = ~n_9616 &  n_47401;
assign n_47403 = ~n_9608 &  n_47402;
assign n_47404 = ~n_9600 &  n_47403;
assign n_47405 = ~n_9592 &  n_47404;
assign n_47406 = ~n_9584 &  n_47405;
assign n_47407 = ~n_9576 &  n_47406;
assign n_47408 = ~n_9568 &  n_47407;
assign n_47409 = ~n_9560 &  n_47408;
assign n_47410 = ~n_9552 &  n_47409;
assign n_47411 = ~n_9544 &  n_47410;
assign n_47412 = ~n_9536 &  n_47411;
assign n_47413 = ~n_9528 &  n_47412;
assign n_47414 = ~n_9520 &  n_47413;
assign n_47415 = ~n_9512 &  n_47414;
assign n_47416 = ~n_9504 &  n_47415;
assign n_47417 = ~n_9496 &  n_47416;
assign n_47418 = ~n_9488 &  n_47417;
assign n_47419 = ~n_9480 &  n_47418;
assign n_47420 = ~n_9472 &  n_47419;
assign n_47421 = ~n_9464 &  n_47420;
assign n_47422 = ~n_9456 &  n_47421;
assign n_47423 = ~n_9448 &  n_47422;
assign n_47424 = ~n_9440 &  n_47423;
assign n_47425 = ~n_9299 &  n_47424;
assign n_47426 = ~n_9293 &  n_47425;
assign n_47427 = ~n_9287 &  n_47426;
assign n_47428 = ~n_9281 &  n_47427;
assign n_47429 = ~n_9275 &  n_47428;
assign n_47430 = ~n_9269 &  n_47429;
assign n_47431 = ~n_9263 &  n_47430;
assign n_47432 = ~n_9257 &  n_47431;
assign n_47433 = ~n_9251 &  n_47432;
assign n_47434 = ~n_9245 &  n_47433;
assign n_47435 = ~n_9239 &  n_47434;
assign n_47436 = ~n_9233 &  n_47435;
assign n_47437 = ~n_9227 &  n_47436;
assign n_47438 = ~n_9221 &  n_47437;
assign n_47439 = ~n_9215 &  n_47438;
assign n_47440 = ~n_9209 &  n_47439;
assign n_47441 = ~n_9203 &  n_47440;
assign n_47442 = ~n_9197 &  n_47441;
assign n_47443 = ~n_9191 &  n_47442;
assign n_47444 = ~n_9185 &  n_47443;
assign n_47445 = ~n_9179 &  n_47444;
assign n_47446 = ~n_9173 &  n_47445;
assign n_47447 = ~n_9167 &  n_47446;
assign n_47448 = ~n_9161 &  n_47447;
assign n_47449 = ~n_9155 &  n_47448;
assign n_47450 = ~n_9149 &  n_47449;
assign n_47451 = ~n_9143 &  n_47450;
assign n_47452 = ~n_9137 &  n_47451;
assign n_47453 = ~n_9131 &  n_47452;
assign n_47454 = ~n_9125 &  n_47453;
assign n_47455 = ~n_9119 &  n_47454;
assign n_47456 = ~n_9113 &  n_47455;
assign n_47457 = ~n_9107 &  n_47456;
assign n_47458 = ~n_9102 &  n_47457;
assign n_47459 = ~n_9097 &  n_47458;
assign n_47460 = ~n_9092 &  n_47459;
assign n_47461 = ~n_9087 &  n_47460;
assign n_47462 = ~n_9082 &  n_47461;
assign n_47463 = ~n_9077 &  n_47462;
assign n_47464 = ~n_9072 &  n_47463;
assign n_47465 = ~n_9067 &  n_47464;
assign n_47466 = ~n_9062 &  n_47465;
assign n_47467 = ~n_9057 &  n_47466;
assign n_47468 = ~n_9052 &  n_47467;
assign n_47469 = ~n_9047 &  n_47468;
assign n_47470 = ~n_9042 &  n_47469;
assign n_47471 = ~n_9037 &  n_47470;
assign n_47472 = ~n_9032 &  n_47471;
assign n_47473 = ~n_9027 &  n_47472;
assign n_47474 = ~n_9022 &  n_47473;
assign n_47475 = ~n_9017 &  n_47474;
assign n_47476 = ~n_9012 &  n_47475;
assign n_47477 = ~n_9007 &  n_47476;
assign n_47478 = ~n_9002 &  n_47477;
assign n_47479 = ~n_8997 &  n_47478;
assign n_47480 = ~n_8992 &  n_47479;
assign n_47481 = ~n_8987 &  n_47480;
assign n_47482 = ~n_8982 &  n_47481;
assign n_47483 = ~n_8977 &  n_47482;
assign n_47484 = ~n_8972 &  n_47483;
assign n_47485 = ~n_8967 &  n_47484;
assign n_47486 = ~n_8962 &  n_47485;
assign n_47487 = ~n_8957 &  n_47486;
assign n_47488 = ~n_8952 &  n_47487;
assign n_47489 = ~n_8947 &  n_47488;
assign n_47490 = ~n_8943 &  n_47489;
assign n_47491 = ~n_8939 &  n_47490;
assign n_47492 = ~n_8935 &  n_47491;
assign n_47493 = ~n_8931 &  n_47492;
assign n_47494 = ~n_8927 &  n_47493;
assign n_47495 = ~n_8923 &  n_47494;
assign n_47496 = ~n_8919 &  n_47495;
assign n_47497 = ~n_8915 &  n_47496;
assign n_47498 = ~n_8911 &  n_47497;
assign n_47499 = ~n_8907 &  n_47498;
assign n_47500 = ~n_8903 &  n_47499;
assign n_47501 = ~n_8899 &  n_47500;
assign n_47502 = ~n_8895 &  n_47501;
assign n_47503 = ~n_8891 &  n_47502;
assign n_47504 = ~n_8887 &  n_47503;
assign n_47505 = ~n_8883 &  n_47504;
assign n_47506 = ~n_8879 &  n_47505;
assign n_47507 = ~n_8875 &  n_47506;
assign n_47508 = ~n_8871 &  n_47507;
assign n_47509 = ~n_8867 &  n_47508;
assign n_47510 = ~n_8863 &  n_47509;
assign n_47511 = ~n_8859 &  n_47510;
assign n_47512 = ~n_8855 &  n_47511;
assign n_47513 = ~n_8851 &  n_47512;
assign n_47514 = ~n_8847 &  n_47513;
assign n_47515 = ~n_8843 &  n_47514;
assign n_47516 = ~n_8839 &  n_47515;
assign n_47517 = ~n_8835 &  n_47516;
assign n_47518 = ~n_8831 &  n_47517;
assign n_47519 = ~n_8827 &  n_47518;
assign n_47520 = ~n_8823 &  n_47519;
assign n_47521 = ~n_8817 &  n_47520;
assign n_47522 = ~n_8803 &  n_47521;
assign n_47523 = ~n_8789 &  n_47522;
assign n_47524 = ~n_8775 &  n_47523;
assign n_47525 = ~n_8761 &  n_47524;
assign n_47526 = ~n_8747 &  n_47525;
assign n_47527 = ~n_8733 &  n_47526;
assign n_47528 = ~n_8719 &  n_47527;
assign n_47529 = ~n_8705 &  n_47528;
assign n_47530 = ~n_8691 &  n_47529;
assign n_47531 = ~n_8677 &  n_47530;
assign n_47532 = ~n_8663 &  n_47531;
assign n_47533 = ~n_8649 &  n_47532;
assign n_47534 = ~n_8635 &  n_47533;
assign n_47535 = ~n_8621 &  n_47534;
assign n_47536 = ~n_8607 &  n_47535;
assign n_47537 = ~n_8593 &  n_47536;
assign n_47538 = ~n_8579 &  n_47537;
assign n_47539 = ~n_8565 &  n_47538;
assign n_47540 = ~n_8551 &  n_47539;
assign n_47541 = ~n_8537 &  n_47540;
assign n_47542 = ~n_8523 &  n_47541;
assign n_47543 = ~n_8509 &  n_47542;
assign n_47544 = ~n_8495 &  n_47543;
assign n_47545 = ~n_8481 &  n_47544;
assign n_47546 = ~n_8467 &  n_47545;
assign n_47547 = ~n_8453 &  n_47546;
assign n_47548 = ~n_8439 &  n_47547;
assign n_47549 = ~n_8425 &  n_47548;
assign n_47550 = ~n_8411 &  n_47549;
assign n_47551 = ~n_8397 &  n_47550;
assign n_47552 = ~n_8383 &  n_47551;
assign n_47553 = ~n_8343 &  n_47552;
assign n_47554 = ~n_8336 &  n_47553;
assign n_47555 = ~n_8327 &  n_47554;
assign n_47556 = ~n_8318 &  n_47555;
assign n_47557 = ~n_8309 &  n_47556;
assign n_47558 = ~n_8300 &  n_47557;
assign n_47559 = ~n_8291 &  n_47558;
assign n_47560 = ~n_8282 &  n_47559;
assign n_47561 = ~n_8273 &  n_47560;
assign n_47562 = ~n_8264 &  n_47561;
assign n_47563 = ~n_8255 &  n_47562;
assign n_47564 = ~n_8246 &  n_47563;
assign n_47565 = ~n_8237 &  n_47564;
assign n_47566 = ~n_8228 &  n_47565;
assign n_47567 = ~n_8219 &  n_47566;
assign n_47568 = ~n_8210 &  n_47567;
assign n_47569 = ~n_8201 &  n_47568;
assign n_47570 = ~n_8192 &  n_47569;
assign n_47571 = ~n_8183 &  n_47570;
assign n_47572 = ~n_8174 &  n_47571;
assign n_47573 = ~n_8165 &  n_47572;
assign n_47574 = ~n_8156 &  n_47573;
assign n_47575 = ~n_8146 &  n_47574;
assign n_47576 = ~n_8137 &  n_47575;
assign n_47577 = ~n_8127 &  n_47576;
assign n_47578 = ~n_8118 &  n_47577;
assign n_47579 = ~n_8107 &  n_47578;
assign n_47580 = ~n_8098 &  n_47579;
assign n_47581 = ~n_8088 &  n_47580;
assign n_47582 = ~n_8079 &  n_47581;
assign n_47583 = ~n_8069 &  n_47582;
assign n_47584 = ~n_8061 &  n_47583;
assign n_47585 = ~n_8048 &  n_47584;
assign n_47586 = ~n_8042 &  n_47585;
assign n_47587 = ~n_8036 &  n_47586;
assign n_47588 = ~n_8030 &  n_47587;
assign n_47589 = ~n_8024 &  n_47588;
assign n_47590 = ~n_8018 &  n_47589;
assign n_47591 = ~n_8012 &  n_47590;
assign n_47592 = ~n_8006 &  n_47591;
assign n_47593 = ~n_8000 &  n_47592;
assign n_47594 = ~n_7994 &  n_47593;
assign n_47595 = ~n_7988 &  n_47594;
assign n_47596 = ~n_7982 &  n_47595;
assign n_47597 = ~n_7976 &  n_47596;
assign n_47598 = ~n_7970 &  n_47597;
assign n_47599 = ~n_7964 &  n_47598;
assign n_47600 = ~n_7958 &  n_47599;
assign n_47601 = ~n_7952 &  n_47600;
assign n_47602 = ~n_7946 &  n_47601;
assign n_47603 = ~n_7940 &  n_47602;
assign n_47604 = ~n_7934 &  n_47603;
assign n_47605 = ~n_7928 &  n_47604;
assign n_47606 = ~n_7922 &  n_47605;
assign n_47607 = ~n_7916 &  n_47606;
assign n_47608 = ~n_7910 &  n_47607;
assign n_47609 = ~n_7904 &  n_47608;
assign n_47610 = ~n_7898 &  n_47609;
assign n_47611 = ~n_7892 &  n_47610;
assign n_47612 = ~n_7886 &  n_47611;
assign n_47613 = ~n_7880 &  n_47612;
assign n_47614 = ~n_7874 &  n_47613;
assign n_47615 = ~n_7868 &  n_47614;
assign n_47616 = ~n_7862 &  n_47615;
assign n_47617 = ~n_7854 &  n_47616;
assign n_47618 = ~n_7848 &  n_47617;
assign n_47619 = ~n_7842 &  n_47618;
assign n_47620 = ~n_7836 &  n_47619;
assign n_47621 = ~n_7830 &  n_47620;
assign n_47622 = ~n_7824 &  n_47621;
assign n_47623 = ~n_7818 &  n_47622;
assign n_47624 = ~n_7812 &  n_47623;
assign n_47625 = ~n_7806 &  n_47624;
assign n_47626 = ~n_7800 &  n_47625;
assign n_47627 = ~n_7794 &  n_47626;
assign n_47628 = ~n_7788 &  n_47627;
assign n_47629 = ~n_7782 &  n_47628;
assign n_47630 = ~n_7776 &  n_47629;
assign n_47631 = ~n_7770 &  n_47630;
assign n_47632 = ~n_7764 &  n_47631;
assign n_47633 = ~n_7758 &  n_47632;
assign n_47634 = ~n_7752 &  n_47633;
assign n_47635 = ~n_7746 &  n_47634;
assign n_47636 = ~n_7740 &  n_47635;
assign n_47637 = ~n_7734 &  n_47636;
assign n_47638 = ~n_7728 &  n_47637;
assign n_47639 = ~n_7722 &  n_47638;
assign n_47640 = ~n_7716 &  n_47639;
assign n_47641 = ~n_7710 &  n_47640;
assign n_47642 = ~n_7704 &  n_47641;
assign n_47643 = ~n_7698 &  n_47642;
assign n_47644 = ~n_7692 &  n_47643;
assign n_47645 = ~n_7686 &  n_47644;
assign n_47646 = ~n_7680 &  n_47645;
assign n_47647 = ~n_7674 &  n_47646;
assign n_47648 = ~n_7668 &  n_47647;
assign n_47649 = ~n_7660 &  n_47648;
assign n_47650 = ~n_7654 &  n_47649;
assign n_47651 = ~n_7648 &  n_47650;
assign n_47652 = ~n_7642 &  n_47651;
assign n_47653 = ~n_7636 &  n_47652;
assign n_47654 = ~n_7630 &  n_47653;
assign n_47655 = ~n_7624 &  n_47654;
assign n_47656 = ~n_7618 &  n_47655;
assign n_47657 = ~n_7612 &  n_47656;
assign n_47658 = ~n_7606 &  n_47657;
assign n_47659 = ~n_7600 &  n_47658;
assign n_47660 = ~n_7594 &  n_47659;
assign n_47661 = ~n_7588 &  n_47660;
assign n_47662 = ~n_7582 &  n_47661;
assign n_47663 = ~n_7576 &  n_47662;
assign n_47664 = ~n_7570 &  n_47663;
assign n_47665 = ~n_7564 &  n_47664;
assign n_47666 = ~n_7558 &  n_47665;
assign n_47667 = ~n_7552 &  n_47666;
assign n_47668 = ~n_7546 &  n_47667;
assign n_47669 = ~n_7540 &  n_47668;
assign n_47670 = ~n_7534 &  n_47669;
assign n_47671 = ~n_7528 &  n_47670;
assign n_47672 = ~n_7522 &  n_47671;
assign n_47673 = ~n_7516 &  n_47672;
assign n_47674 = ~n_7510 &  n_47673;
assign n_47675 = ~n_7504 &  n_47674;
assign n_47676 = ~n_7498 &  n_47675;
assign n_47677 = ~n_7492 &  n_47676;
assign n_47678 = ~n_7486 &  n_47677;
assign n_47679 = ~n_7480 &  n_47678;
assign n_47680 = ~n_7474 &  n_47679;
assign n_47681 = ~n_7466 &  n_47680;
assign n_47682 = ~n_7460 &  n_47681;
assign n_47683 = ~n_7454 &  n_47682;
assign n_47684 = ~n_7448 &  n_47683;
assign n_47685 = ~n_7442 &  n_47684;
assign n_47686 = ~n_7436 &  n_47685;
assign n_47687 = ~n_7430 &  n_47686;
assign n_47688 = ~n_7424 &  n_47687;
assign n_47689 = ~n_7418 &  n_47688;
assign n_47690 = ~n_7412 &  n_47689;
assign n_47691 = ~n_7406 &  n_47690;
assign n_47692 = ~n_7400 &  n_47691;
assign n_47693 = ~n_7394 &  n_47692;
assign n_47694 = ~n_7388 &  n_47693;
assign n_47695 = ~n_7382 &  n_47694;
assign n_47696 = ~n_7376 &  n_47695;
assign n_47697 = ~n_7370 &  n_47696;
assign n_47698 = ~n_7364 &  n_47697;
assign n_47699 = ~n_7358 &  n_47698;
assign n_47700 = ~n_7352 &  n_47699;
assign n_47701 = ~n_7346 &  n_47700;
assign n_47702 = ~n_7340 &  n_47701;
assign n_47703 = ~n_7334 &  n_47702;
assign n_47704 = ~n_7328 &  n_47703;
assign n_47705 = ~n_7322 &  n_47704;
assign n_47706 = ~n_7316 &  n_47705;
assign n_47707 = ~n_7310 &  n_47706;
assign n_47708 = ~n_7304 &  n_47707;
assign n_47709 = ~n_7298 &  n_47708;
assign n_47710 = ~n_7292 &  n_47709;
assign n_47711 = ~n_7286 &  n_47710;
assign n_47712 = ~n_7280 &  n_47711;
assign n_47713 = ~n_7272 &  n_47712;
assign n_47714 = ~n_7266 &  n_47713;
assign n_47715 = ~n_7260 &  n_47714;
assign n_47716 = ~n_7254 &  n_47715;
assign n_47717 = ~n_7248 &  n_47716;
assign n_47718 = ~n_7242 &  n_47717;
assign n_47719 = ~n_7236 &  n_47718;
assign n_47720 = ~n_7230 &  n_47719;
assign n_47721 = ~n_7224 &  n_47720;
assign n_47722 = ~n_7218 &  n_47721;
assign n_47723 = ~n_7212 &  n_47722;
assign n_47724 = ~n_7206 &  n_47723;
assign n_47725 = ~n_7200 &  n_47724;
assign n_47726 = ~n_7194 &  n_47725;
assign n_47727 = ~n_7188 &  n_47726;
assign n_47728 = ~n_7182 &  n_47727;
assign n_47729 = ~n_7176 &  n_47728;
assign n_47730 = ~n_7170 &  n_47729;
assign n_47731 = ~n_7164 &  n_47730;
assign n_47732 = ~n_7158 &  n_47731;
assign n_47733 = ~n_7152 &  n_47732;
assign n_47734 = ~n_7146 &  n_47733;
assign n_47735 = ~n_7140 &  n_47734;
assign n_47736 = ~n_7134 &  n_47735;
assign n_47737 = ~n_7128 &  n_47736;
assign n_47738 = ~n_7122 &  n_47737;
assign n_47739 = ~n_7116 &  n_47738;
assign n_47740 = ~n_7110 &  n_47739;
assign n_47741 = ~n_7104 &  n_47740;
assign n_47742 = ~n_7098 &  n_47741;
assign n_47743 = ~n_7092 &  n_47742;
assign n_47744 = ~n_7086 &  n_47743;
assign n_47745 = ~n_7077 &  n_47744;
assign n_47746 = ~n_7071 &  n_47745;
assign n_47747 = ~n_7065 &  n_47746;
assign n_47748 = ~n_7059 &  n_47747;
assign n_47749 = ~n_7053 &  n_47748;
assign n_47750 = ~n_7047 &  n_47749;
assign n_47751 = ~n_7041 &  n_47750;
assign n_47752 = ~n_7035 &  n_47751;
assign n_47753 = ~n_7029 &  n_47752;
assign n_47754 = ~n_7023 &  n_47753;
assign n_47755 = ~n_7017 &  n_47754;
assign n_47756 = ~n_7011 &  n_47755;
assign n_47757 = ~n_7005 &  n_47756;
assign n_47758 = ~n_6999 &  n_47757;
assign n_47759 = ~n_6993 &  n_47758;
assign n_47760 = ~n_6987 &  n_47759;
assign n_47761 = ~n_6981 &  n_47760;
assign n_47762 = ~n_6975 &  n_47761;
assign n_47763 = ~n_6969 &  n_47762;
assign n_47764 = ~n_6963 &  n_47763;
assign n_47765 = ~n_6957 &  n_47764;
assign n_47766 = ~n_6951 &  n_47765;
assign n_47767 = ~n_6945 &  n_47766;
assign n_47768 = ~n_6939 &  n_47767;
assign n_47769 = ~n_6933 &  n_47768;
assign n_47770 = ~n_6927 &  n_47769;
assign n_47771 = ~n_6921 &  n_47770;
assign n_47772 = ~n_6915 &  n_47771;
assign n_47773 = ~n_6909 &  n_47772;
assign n_47774 = ~n_6903 &  n_47773;
assign n_47775 = ~n_6897 &  n_47774;
assign n_47776 = ~n_6891 &  n_47775;
assign n_47777 = ~n_6875 &  n_47776;
assign n_47778 = ~n_6869 &  n_47777;
assign n_47779 = ~n_6863 &  n_47778;
assign n_47780 = ~n_6857 &  n_47779;
assign n_47781 = ~n_6851 &  n_47780;
assign n_47782 = ~n_6845 &  n_47781;
assign n_47783 = ~n_6839 &  n_47782;
assign n_47784 = ~n_6833 &  n_47783;
assign n_47785 = ~n_6827 &  n_47784;
assign n_47786 = ~n_6821 &  n_47785;
assign n_47787 = ~n_6815 &  n_47786;
assign n_47788 = ~n_6809 &  n_47787;
assign n_47789 = ~n_6803 &  n_47788;
assign n_47790 = ~n_6797 &  n_47789;
assign n_47791 = ~n_6791 &  n_47790;
assign n_47792 = ~n_6785 &  n_47791;
assign n_47793 = ~n_6779 &  n_47792;
assign n_47794 = ~n_6773 &  n_47793;
assign n_47795 = ~n_6767 &  n_47794;
assign n_47796 = ~n_6761 &  n_47795;
assign n_47797 = ~n_6755 &  n_47796;
assign n_47798 = ~n_6749 &  n_47797;
assign n_47799 = ~n_6743 &  n_47798;
assign n_47800 = ~n_6737 &  n_47799;
assign n_47801 = ~n_6731 &  n_47800;
assign n_47802 = ~n_6725 &  n_47801;
assign n_47803 = ~n_6719 &  n_47802;
assign n_47804 = ~n_6713 &  n_47803;
assign n_47805 = ~n_6707 &  n_47804;
assign n_47806 = ~n_6701 &  n_47805;
assign n_47807 = ~n_6695 &  n_47806;
assign n_47808 = ~n_6689 &  n_47807;
assign n_47809 = ~n_6683 &  n_47808;
assign n_47810 = ~n_6677 &  n_47809;
assign n_47811 = ~n_6671 &  n_47810;
assign n_47812 = ~n_6665 &  n_47811;
assign n_47813 = ~n_6659 &  n_47812;
assign n_47814 = ~n_6653 &  n_47813;
assign n_47815 = ~n_6647 &  n_47814;
assign n_47816 = ~n_6641 &  n_47815;
assign n_47817 = ~n_6635 &  n_47816;
assign n_47818 = ~n_6629 &  n_47817;
assign n_47819 = ~n_6623 &  n_47818;
assign n_47820 = ~n_6617 &  n_47819;
assign n_47821 = ~n_6611 &  n_47820;
assign n_47822 = ~n_6605 &  n_47821;
assign n_47823 = ~n_6599 &  n_47822;
assign n_47824 = ~n_6593 &  n_47823;
assign n_47825 = ~n_6587 &  n_47824;
assign n_47826 = ~n_6581 &  n_47825;
assign n_47827 = ~n_6575 &  n_47826;
assign n_47828 = ~n_6569 &  n_47827;
assign n_47829 = ~n_6563 &  n_47828;
assign n_47830 = ~n_6557 &  n_47829;
assign n_47831 = ~n_6551 &  n_47830;
assign n_47832 = ~n_6545 &  n_47831;
assign n_47833 = ~n_6539 &  n_47832;
assign n_47834 = ~n_6533 &  n_47833;
assign n_47835 = ~n_6524 &  n_47834;
assign n_47836 = ~n_6518 &  n_47835;
assign n_47837 = ~n_6512 &  n_47836;
assign n_47838 = ~n_6506 &  n_47837;
assign n_47839 = ~n_6500 &  n_47838;
assign n_47840 = ~n_6494 &  n_47839;
assign n_47841 = ~n_6488 &  n_47840;
assign n_47842 = ~n_6482 &  n_47841;
assign n_47843 = ~n_6476 &  n_47842;
assign n_47844 = ~n_6470 &  n_47843;
assign n_47845 = ~n_6464 &  n_47844;
assign n_47846 = ~n_6458 &  n_47845;
assign n_47847 = ~n_6452 &  n_47846;
assign n_47848 = ~n_6446 &  n_47847;
assign n_47849 = ~n_6440 &  n_47848;
assign n_47850 = ~n_6434 &  n_47849;
assign n_47851 = ~n_6428 &  n_47850;
assign n_47852 = ~n_6422 &  n_47851;
assign n_47853 = ~n_6416 &  n_47852;
assign n_47854 = ~n_6410 &  n_47853;
assign n_47855 = ~n_6404 &  n_47854;
assign n_47856 = ~n_6398 &  n_47855;
assign n_47857 = ~n_6392 &  n_47856;
assign n_47858 = ~n_6386 &  n_47857;
assign n_47859 = ~n_6376 &  n_47858;
assign n_47860 = ~n_6370 &  n_47859;
assign n_47861 = ~n_6364 &  n_47860;
assign n_47862 = ~n_6358 &  n_47861;
assign n_47863 = ~n_6352 &  n_47862;
assign n_47864 = ~n_6346 &  n_47863;
assign n_47865 = ~n_6340 &  n_47864;
assign n_47866 = ~n_6334 &  n_47865;
assign n_47867 = ~n_6328 &  n_47866;
assign n_47868 = ~n_6322 &  n_47867;
assign n_47869 = ~n_6316 &  n_47868;
assign n_47870 = ~n_6310 &  n_47869;
assign n_47871 = ~n_6304 &  n_47870;
assign n_47872 = ~n_6298 &  n_47871;
assign n_47873 = ~n_6292 &  n_47872;
assign n_47874 = ~n_6286 &  n_47873;
assign n_47875 = ~n_6280 &  n_47874;
assign n_47876 = ~n_6274 &  n_47875;
assign n_47877 = ~n_6268 &  n_47876;
assign n_47878 = ~n_6262 &  n_47877;
assign n_47879 = ~n_6256 &  n_47878;
assign n_47880 = ~n_6250 &  n_47879;
assign n_47881 = ~n_6244 &  n_47880;
assign n_47882 = ~n_6238 &  n_47881;
assign n_47883 = ~n_6232 &  n_47882;
assign n_47884 = ~n_6226 &  n_47883;
assign n_47885 = ~n_6220 &  n_47884;
assign n_47886 = ~n_6214 &  n_47885;
assign n_47887 = ~n_6208 &  n_47886;
assign n_47888 = ~n_6202 &  n_47887;
assign n_47889 = ~n_6196 &  n_47888;
assign n_47890 = ~n_6190 &  n_47889;
assign n_47891 = ~n_6179 &  n_47890;
assign n_47892 = ~n_6173 &  n_47891;
assign n_47893 = ~n_6167 &  n_47892;
assign n_47894 = ~n_6161 &  n_47893;
assign n_47895 = ~n_6155 &  n_47894;
assign n_47896 = ~n_6149 &  n_47895;
assign n_47897 = ~n_6143 &  n_47896;
assign n_47898 = ~n_6137 &  n_47897;
assign n_47899 = ~n_6131 &  n_47898;
assign n_47900 = ~n_6125 &  n_47899;
assign n_47901 = ~n_6119 &  n_47900;
assign n_47902 = ~n_6113 &  n_47901;
assign n_47903 = ~n_6107 &  n_47902;
assign n_47904 = ~n_6101 &  n_47903;
assign n_47905 = ~n_6095 &  n_47904;
assign n_47906 = ~n_6089 &  n_47905;
assign n_47907 = ~n_6083 &  n_47906;
assign n_47908 = ~n_6077 &  n_47907;
assign n_47909 = ~n_6071 &  n_47908;
assign n_47910 = ~n_6065 &  n_47909;
assign n_47911 = ~n_6059 &  n_47910;
assign n_47912 = ~n_6053 &  n_47911;
assign n_47913 = ~n_6047 &  n_47912;
assign n_47914 = ~n_6041 &  n_47913;
assign n_47915 = ~n_6035 &  n_47914;
assign n_47916 = ~n_6029 &  n_47915;
assign n_47917 = ~n_6023 &  n_47916;
assign n_47918 = ~n_6017 &  n_47917;
assign n_47919 = ~n_6011 &  n_47918;
assign n_47920 = ~n_6005 &  n_47919;
assign n_47921 = ~n_5999 &  n_47920;
assign n_47922 = ~n_5993 &  n_47921;
assign n_47923 = ~n_5980 &  n_47922;
assign n_47924 = ~n_5970 &  n_47923;
assign n_47925 = ~n_5960 &  n_47924;
assign n_47926 = ~n_5950 &  n_47925;
assign n_47927 = ~n_5940 &  n_47926;
assign n_47928 = ~n_5930 &  n_47927;
assign n_47929 = ~n_5920 &  n_47928;
assign n_47930 = ~n_5910 &  n_47929;
assign n_47931 = ~n_5900 &  n_47930;
assign n_47932 = ~n_5890 &  n_47931;
assign n_47933 = ~n_5880 &  n_47932;
assign n_47934 = ~n_5870 &  n_47933;
assign n_47935 = ~n_5860 &  n_47934;
assign n_47936 = ~n_5850 &  n_47935;
assign n_47937 = ~n_5840 &  n_47936;
assign n_47938 = ~n_5830 &  n_47937;
assign n_47939 = ~n_5820 &  n_47938;
assign n_47940 = ~n_5810 &  n_47939;
assign n_47941 = ~n_5800 &  n_47940;
assign n_47942 = ~n_5790 &  n_47941;
assign n_47943 = ~n_5780 &  n_47942;
assign n_47944 = ~n_5770 &  n_47943;
assign n_47945 = ~n_5760 &  n_47944;
assign n_47946 = ~n_5750 &  n_47945;
assign n_47947 = ~n_5740 &  n_47946;
assign n_47948 = ~n_5730 &  n_47947;
assign n_47949 = ~n_5720 &  n_47948;
assign n_47950 = ~n_5710 &  n_47949;
assign n_47951 = ~n_5700 &  n_47950;
assign n_47952 = ~n_5690 &  n_47951;
assign n_47953 = ~n_5680 &  n_47952;
assign n_47954 = ~n_5670 &  n_47953;
assign n_47955 = ~n_5644 &  n_47954;
assign n_47956 = ~n_5604 &  n_47955;
assign n_47957 = ~n_5561 &  n_47956;
assign n_47958 = ~n_5518 &  n_47957;
assign n_47959 = ~n_5475 &  n_47958;
assign n_47960 = ~n_5432 &  n_47959;
assign n_47961 = ~n_5389 &  n_47960;
assign n_47962 = ~n_5346 &  n_47961;
assign n_47963 = ~n_5303 &  n_47962;
assign n_47964 = ~n_5260 &  n_47963;
assign n_47965 = ~n_5217 &  n_47964;
assign n_47966 = ~n_5174 &  n_47965;
assign n_47967 = ~n_5131 &  n_47966;
assign n_47968 = ~n_5088 &  n_47967;
assign n_47969 = ~n_5045 &  n_47968;
assign n_47970 = ~n_5002 &  n_47969;
assign n_47971 = ~n_4959 &  n_47970;
assign n_47972 = ~n_4916 &  n_47971;
assign n_47973 = ~n_4873 &  n_47972;
assign n_47974 = ~n_4830 &  n_47973;
assign n_47975 = ~n_4787 &  n_47974;
assign n_47976 = ~n_4744 &  n_47975;
assign n_47977 = ~n_4701 &  n_47976;
assign n_47978 = ~n_4658 &  n_47977;
assign n_47979 = ~n_4615 &  n_47978;
assign n_47980 = ~n_4572 &  n_47979;
assign n_47981 = ~n_4529 &  n_47980;
assign n_47982 = ~n_4486 &  n_47981;
assign n_47983 = ~n_4443 &  n_47982;
assign n_47984 = ~n_4400 &  n_47983;
assign n_47985 = ~n_4351 &  n_47984;
assign n_47986 = ~n_4314 &  n_47985;
assign n_47987 = ~n_4282 &  n_47986;
assign n_47988 = ~n_4276 &  n_47987;
assign n_47989 = ~n_4270 &  n_47988;
assign n_47990 = ~n_4264 &  n_47989;
assign n_47991 = ~n_4258 &  n_47990;
assign n_47992 = ~n_4252 &  n_47991;
assign n_47993 = ~n_4246 &  n_47992;
assign n_47994 = ~n_4240 &  n_47993;
assign n_47995 = ~n_4234 &  n_47994;
assign n_47996 = ~n_4228 &  n_47995;
assign n_47997 = ~n_4222 &  n_47996;
assign n_47998 = ~n_4216 &  n_47997;
assign n_47999 = ~n_4210 &  n_47998;
assign n_48000 = ~n_4204 &  n_47999;
assign n_48001 = ~n_4198 &  n_48000;
assign n_48002 = ~n_4192 &  n_48001;
assign n_48003 = ~n_4186 &  n_48002;
assign n_48004 = ~n_4180 &  n_48003;
assign n_48005 = ~n_4174 &  n_48004;
assign n_48006 = ~n_4168 &  n_48005;
assign n_48007 = ~n_4162 &  n_48006;
assign n_48008 = ~n_4156 &  n_48007;
assign n_48009 = ~n_4150 &  n_48008;
assign n_48010 = ~n_4144 &  n_48009;
assign n_48011 = ~n_4138 &  n_48010;
assign n_48012 = ~n_4132 &  n_48011;
assign n_48013 = ~n_4126 &  n_48012;
assign n_48014 = ~n_4120 &  n_48013;
assign n_48015 = ~n_4114 &  n_48014;
assign n_48016 = ~n_4108 &  n_48015;
assign n_48017 = ~n_4102 &  n_48016;
assign n_48018 = ~n_4096 &  n_48017;
assign n_48019 = ~n_4087 &  n_48018;
assign n_48020 = ~n_4073 &  n_48019;
assign n_48021 = ~n_4059 &  n_48020;
assign n_48022 = ~n_4045 &  n_48021;
assign n_48023 = ~n_4031 &  n_48022;
assign n_48024 = ~n_4017 &  n_48023;
assign n_48025 = ~n_4003 &  n_48024;
assign n_48026 = ~n_3989 &  n_48025;
assign n_48027 = ~n_3975 &  n_48026;
assign n_48028 = ~n_3961 &  n_48027;
assign n_48029 = ~n_3947 &  n_48028;
assign n_48030 = ~n_3933 &  n_48029;
assign n_48031 = ~n_3919 &  n_48030;
assign n_48032 = ~n_3905 &  n_48031;
assign n_48033 = ~n_3891 &  n_48032;
assign n_48034 = ~n_3877 &  n_48033;
assign n_48035 = ~n_3863 &  n_48034;
assign n_48036 = ~n_3849 &  n_48035;
assign n_48037 = ~n_3835 &  n_48036;
assign n_48038 = ~n_3821 &  n_48037;
assign n_48039 = ~n_3807 &  n_48038;
assign n_48040 = ~n_3793 &  n_48039;
assign n_48041 = ~n_3779 &  n_48040;
assign n_48042 = ~n_3765 &  n_48041;
assign n_48043 = ~n_3751 &  n_48042;
assign n_48044 = ~n_3737 &  n_48043;
assign n_48045 = ~n_3723 &  n_48044;
assign n_48046 = ~n_3709 &  n_48045;
assign n_48047 = ~n_3695 &  n_48046;
assign n_48048 = ~n_3681 &  n_48047;
assign n_48049 = ~n_3667 &  n_48048;
assign n_48050 = ~n_3653 &  n_48049;
assign n_48051 = ~n_3614 &  n_48050;
assign n_48052 = ~n_3610 &  n_48051;
assign n_48053 = ~n_3606 &  n_48052;
assign n_48054 = ~n_3602 &  n_48053;
assign n_48055 = ~n_3598 &  n_48054;
assign n_48056 = ~n_3594 &  n_48055;
assign n_48057 = ~n_3590 &  n_48056;
assign n_48058 = ~n_3586 &  n_48057;
assign n_48059 = ~n_3582 &  n_48058;
assign n_48060 = ~n_3578 &  n_48059;
assign n_48061 = ~n_3574 &  n_48060;
assign n_48062 = ~n_3570 &  n_48061;
assign n_48063 = ~n_3566 &  n_48062;
assign n_48064 = ~n_3562 &  n_48063;
assign n_48065 = ~n_3558 &  n_48064;
assign n_48066 = ~n_3554 &  n_48065;
assign n_48067 = ~n_3550 &  n_48066;
assign n_48068 = ~n_3546 &  n_48067;
assign n_48069 = ~n_3542 &  n_48068;
assign n_48070 = ~n_3538 &  n_48069;
assign n_48071 = ~n_3534 &  n_48070;
assign n_48072 = ~n_3530 &  n_48071;
assign n_48073 = ~n_3525 &  n_48072;
assign n_48074 = ~n_3521 &  n_48073;
assign n_48075 = ~n_3516 &  n_48074;
assign n_48076 = ~n_3512 &  n_48075;
assign n_48077 = ~n_3507 &  n_48076;
assign n_48078 = ~n_3502 &  n_48077;
assign n_48079 = ~n_3497 &  n_48078;
assign n_48080 = ~n_3493 &  n_48079;
assign n_48081 = ~n_3489 &  n_48080;
assign n_48082 = ~n_3485 &  n_48081;
assign n_48083 = ~n_3480 &  n_48082;
assign n_48084 = ~n_3476 &  n_48083;
assign n_48085 = ~n_3472 &  n_48084;
assign n_48086 = ~n_3468 &  n_48085;
assign n_48087 = ~n_3464 &  n_48086;
assign n_48088 = ~n_3460 &  n_48087;
assign n_48089 = ~n_3456 &  n_48088;
assign n_48090 = ~n_3452 &  n_48089;
assign n_48091 = ~n_3448 &  n_48090;
assign n_48092 = ~n_3444 &  n_48091;
assign n_48093 = ~n_3440 &  n_48092;
assign n_48094 = ~n_3436 &  n_48093;
assign n_48095 = ~n_3432 &  n_48094;
assign n_48096 = ~n_3428 &  n_48095;
assign n_48097 = ~n_3424 &  n_48096;
assign n_48098 = ~n_3420 &  n_48097;
assign n_48099 = ~n_3416 &  n_48098;
assign n_48100 = ~n_3412 &  n_48099;
assign n_48101 = ~n_3408 &  n_48100;
assign n_48102 = ~n_3404 &  n_48101;
assign n_48103 = ~n_3400 &  n_48102;
assign n_48104 = ~n_3396 &  n_48103;
assign n_48105 = ~n_3392 &  n_48104;
assign n_48106 = ~n_3388 &  n_48105;
assign n_48107 = ~n_3384 &  n_48106;
assign n_48108 = ~n_3380 &  n_48107;
assign n_48109 = ~n_3376 &  n_48108;
assign n_48110 = ~n_3372 &  n_48109;
assign n_48111 = ~n_3368 &  n_48110;
assign n_48112 = ~n_3364 &  n_48111;
assign n_48113 = ~n_3360 &  n_48112;
assign n_48114 = ~n_3355 &  n_48113;
assign n_48115 = ~n_3337 &  n_48114;
assign n_48116 = ~n_3331 &  n_48115;
assign n_48117 = ~n_3325 &  n_48116;
assign n_48118 = ~n_3319 &  n_48117;
assign n_48119 = ~n_3313 &  n_48118;
assign n_48120 = ~n_3307 &  n_48119;
assign n_48121 = ~n_3301 &  n_48120;
assign n_48122 = ~n_3295 &  n_48121;
assign n_48123 = ~n_3289 &  n_48122;
assign n_48124 = ~n_3283 &  n_48123;
assign n_48125 = ~n_3277 &  n_48124;
assign n_48126 = ~n_3271 &  n_48125;
assign n_48127 = ~n_3265 &  n_48126;
assign n_48128 = ~n_3259 &  n_48127;
assign n_48129 = ~n_3253 &  n_48128;
assign n_48130 = ~n_3247 &  n_48129;
assign n_48131 = ~n_3241 &  n_48130;
assign n_48132 = ~n_3235 &  n_48131;
assign n_48133 = ~n_3229 &  n_48132;
assign n_48134 = ~n_3223 &  n_48133;
assign n_48135 = ~n_3217 &  n_48134;
assign n_48136 = ~n_3211 &  n_48135;
assign n_48137 = ~n_3205 &  n_48136;
assign n_48138 = ~n_3199 &  n_48137;
assign n_48139 = ~n_3193 &  n_48138;
assign n_48140 = ~n_3187 &  n_48139;
assign n_48141 = ~n_3181 &  n_48140;
assign n_48142 = ~n_3175 &  n_48141;
assign n_48143 = ~n_3169 &  n_48142;
assign n_48144 = ~n_3163 &  n_48143;
assign n_48145 = ~n_3157 &  n_48144;
assign n_48146 = ~n_3151 &  n_48145;
assign n_48147 = ~n_3140 &  n_48146;
assign n_48148 = ~n_3132 &  n_48147;
assign n_48149 = ~n_3124 &  n_48148;
assign n_48150 = ~n_3116 &  n_48149;
assign n_48151 = ~n_3108 &  n_48150;
assign n_48152 = ~n_3100 &  n_48151;
assign n_48153 = ~n_3092 &  n_48152;
assign n_48154 = ~n_3084 &  n_48153;
assign n_48155 = ~n_3076 &  n_48154;
assign n_48156 = ~n_3068 &  n_48155;
assign n_48157 = ~n_3060 &  n_48156;
assign n_48158 = ~n_3052 &  n_48157;
assign n_48159 = ~n_3044 &  n_48158;
assign n_48160 = ~n_3036 &  n_48159;
assign n_48161 = ~n_3028 &  n_48160;
assign n_48162 = ~n_3020 &  n_48161;
assign n_48163 = ~n_3012 &  n_48162;
assign n_48164 = ~n_3004 &  n_48163;
assign n_48165 = ~n_2996 &  n_48164;
assign n_48166 = ~n_2988 &  n_48165;
assign n_48167 = ~n_2980 &  n_48166;
assign n_48168 = ~n_2972 &  n_48167;
assign n_48169 = ~n_2964 &  n_48168;
assign n_48170 = ~n_2956 &  n_48169;
assign n_48171 = ~n_2948 &  n_48170;
assign n_48172 = ~n_2940 &  n_48171;
assign n_48173 = ~n_2932 &  n_48172;
assign n_48174 = ~n_2924 &  n_48173;
assign n_48175 = ~n_2916 &  n_48174;
assign n_48176 = ~n_2908 &  n_48175;
assign n_48177 = ~n_2900 &  n_48176;
assign n_48178 = ~n_2892 &  n_48177;
assign n_48179 = ~n_2878 &  n_48178;
assign n_48180 = ~n_2872 &  n_48179;
assign n_48181 = ~n_2866 &  n_48180;
assign n_48182 = ~n_2860 &  n_48181;
assign n_48183 = ~n_2854 &  n_48182;
assign n_48184 = ~n_2848 &  n_48183;
assign n_48185 = ~n_2842 &  n_48184;
assign n_48186 = ~n_2836 &  n_48185;
assign n_48187 = ~n_2830 &  n_48186;
assign n_48188 = ~n_2824 &  n_48187;
assign n_48189 = ~n_2818 &  n_48188;
assign n_48190 = ~n_2812 &  n_48189;
assign n_48191 = ~n_2806 &  n_48190;
assign n_48192 = ~n_2800 &  n_48191;
assign n_48193 = ~n_2794 &  n_48192;
assign n_48194 = ~n_2788 &  n_48193;
assign n_48195 = ~n_2782 &  n_48194;
assign n_48196 = ~n_2776 &  n_48195;
assign n_48197 = ~n_2770 &  n_48196;
assign n_48198 = ~n_2764 &  n_48197;
assign n_48199 = ~n_2758 &  n_48198;
assign n_48200 = ~n_2752 &  n_48199;
assign n_48201 = ~n_2746 &  n_48200;
assign n_48202 = ~n_2740 &  n_48201;
assign n_48203 = ~n_2734 &  n_48202;
assign n_48204 = ~n_2728 &  n_48203;
assign n_48205 = ~n_2722 &  n_48204;
assign n_48206 = ~n_2716 &  n_48205;
assign n_48207 = ~n_2710 &  n_48206;
assign n_48208 = ~n_2704 &  n_48207;
assign n_48209 = ~n_2698 &  n_48208;
assign n_48210 = ~n_2692 &  n_48209;
assign n_48211 = ~n_2680 &  n_48210;
assign n_48212 = ~n_2674 &  n_48211;
assign n_48213 = ~n_2668 &  n_48212;
assign n_48214 = ~n_2662 &  n_48213;
assign n_48215 = ~n_2656 &  n_48214;
assign n_48216 = ~n_2650 &  n_48215;
assign n_48217 = ~n_2644 &  n_48216;
assign n_48218 = ~n_2638 &  n_48217;
assign n_48219 = ~n_2632 &  n_48218;
assign n_48220 = ~n_2626 &  n_48219;
assign n_48221 = ~n_2620 &  n_48220;
assign n_48222 = ~n_2614 &  n_48221;
assign n_48223 = ~n_2608 &  n_48222;
assign n_48224 = ~n_2602 &  n_48223;
assign n_48225 = ~n_2596 &  n_48224;
assign n_48226 = ~n_2590 &  n_48225;
assign n_48227 = ~n_2584 &  n_48226;
assign n_48228 = ~n_2578 &  n_48227;
assign n_48229 = ~n_2572 &  n_48228;
assign n_48230 = ~n_2566 &  n_48229;
assign n_48231 = ~n_2560 &  n_48230;
assign n_48232 = ~n_2554 &  n_48231;
assign n_48233 = ~n_2548 &  n_48232;
assign n_48234 = ~n_2542 &  n_48233;
assign n_48235 = ~n_2536 &  n_48234;
assign n_48236 = ~n_2530 &  n_48235;
assign n_48237 = ~n_2524 &  n_48236;
assign n_48238 = ~n_2518 &  n_48237;
assign n_48239 = ~n_2512 &  n_48238;
assign n_48240 = ~n_2506 &  n_48239;
assign n_48241 = ~n_2500 &  n_48240;
assign n_48242 = ~n_2494 &  n_48241;
assign n_48243 = ~n_2484 &  n_48242;
assign n_48244 = ~n_2478 &  n_48243;
assign n_48245 = ~n_2472 &  n_48244;
assign n_48246 = ~n_2466 &  n_48245;
assign n_48247 = ~n_2460 &  n_48246;
assign n_48248 = ~n_2454 &  n_48247;
assign n_48249 = ~n_2448 &  n_48248;
assign n_48250 = ~n_2442 &  n_48249;
assign n_48251 = ~n_2436 &  n_48250;
assign n_48252 = ~n_2430 &  n_48251;
assign n_48253 = ~n_2424 &  n_48252;
assign n_48254 = ~n_2418 &  n_48253;
assign n_48255 = ~n_2412 &  n_48254;
assign n_48256 = ~n_2406 &  n_48255;
assign n_48257 = ~n_2400 &  n_48256;
assign n_48258 = ~n_2394 &  n_48257;
assign n_48259 = ~n_2388 &  n_48258;
assign n_48260 = ~n_2382 &  n_48259;
assign n_48261 = ~n_2376 &  n_48260;
assign n_48262 = ~n_2370 &  n_48261;
assign n_48263 = ~n_2364 &  n_48262;
assign n_48264 = ~n_2358 &  n_48263;
assign n_48265 = ~n_2352 &  n_48264;
assign n_48266 = ~n_2346 &  n_48265;
assign n_48267 = ~n_2340 &  n_48266;
assign n_48268 = ~n_2334 &  n_48267;
assign n_48269 = ~n_2328 &  n_48268;
assign n_48270 = ~n_2322 &  n_48269;
assign n_48271 = ~n_2316 &  n_48270;
assign n_48272 = ~n_2310 &  n_48271;
assign n_48273 = ~n_2304 &  n_48272;
assign n_48274 = ~n_2298 &  n_48273;
assign n_48275 = ~n_2289 &  n_48274;
assign n_48276 = ~n_2283 &  n_48275;
assign n_48277 = ~n_2277 &  n_48276;
assign n_48278 = ~n_2271 &  n_48277;
assign n_48279 = ~n_2265 &  n_48278;
assign n_48280 = ~n_2259 &  n_48279;
assign n_48281 = ~n_2253 &  n_48280;
assign n_48282 = ~n_2247 &  n_48281;
assign n_48283 = ~n_2241 &  n_48282;
assign n_48284 = ~n_2235 &  n_48283;
assign n_48285 = ~n_2229 &  n_48284;
assign n_48286 = ~n_2223 &  n_48285;
assign n_48287 = ~n_2217 &  n_48286;
assign n_48288 = ~n_2211 &  n_48287;
assign n_48289 = ~n_2205 &  n_48288;
assign n_48290 = ~n_2199 &  n_48289;
assign n_48291 = ~n_2193 &  n_48290;
assign n_48292 = ~n_2187 &  n_48291;
assign n_48293 = ~n_2181 &  n_48292;
assign n_48294 = ~n_2175 &  n_48293;
assign n_48295 = ~n_2169 &  n_48294;
assign n_48296 = ~n_2163 &  n_48295;
assign n_48297 = ~n_2157 &  n_48296;
assign n_48298 = ~n_2151 &  n_48297;
assign n_48299 = ~n_2145 &  n_48298;
assign n_48300 = ~n_2139 &  n_48299;
assign n_48301 = ~n_2133 &  n_48300;
assign n_48302 = ~n_2127 &  n_48301;
assign n_48303 = ~n_2121 &  n_48302;
assign n_48304 = ~n_2115 &  n_48303;
assign n_48305 = ~n_2109 &  n_48304;
assign n_48306 = ~n_2103 &  n_48305;
assign n_48307 = ~n_2093 &  n_48306;
assign n_48308 = ~n_2087 &  n_48307;
assign n_48309 = ~n_2081 &  n_48308;
assign n_48310 = ~n_2075 &  n_48309;
assign n_48311 = ~n_2069 &  n_48310;
assign n_48312 = ~n_2063 &  n_48311;
assign n_48313 = ~n_2057 &  n_48312;
assign n_48314 = ~n_2051 &  n_48313;
assign n_48315 = ~n_2045 &  n_48314;
assign n_48316 = ~n_2039 &  n_48315;
assign n_48317 = ~n_2033 &  n_48316;
assign n_48318 = ~n_2027 &  n_48317;
assign n_48319 = ~n_2021 &  n_48318;
assign n_48320 = ~n_2015 &  n_48319;
assign n_48321 = ~n_2009 &  n_48320;
assign n_48322 = ~n_2003 &  n_48321;
assign n_48323 = ~n_1997 &  n_48322;
assign n_48324 = ~n_1991 &  n_48323;
assign n_48325 = ~n_1985 &  n_48324;
assign n_48326 = ~n_1979 &  n_48325;
assign n_48327 = ~n_1973 &  n_48326;
assign n_48328 = ~n_1967 &  n_48327;
assign n_48329 = ~n_1961 &  n_48328;
assign n_48330 = ~n_1955 &  n_48329;
assign n_48331 = ~n_1949 &  n_48330;
assign n_48332 = ~n_1943 &  n_48331;
assign n_48333 = ~n_1937 &  n_48332;
assign n_48334 = ~n_1931 &  n_48333;
assign n_48335 = ~n_1925 &  n_48334;
assign n_48336 = ~n_1919 &  n_48335;
assign n_48337 = ~n_1913 &  n_48336;
assign n_48338 = ~n_1907 &  n_48337;
assign n_48339 = ~n_1893 &  n_48338;
assign n_48340 = ~n_1887 &  n_48339;
assign n_48341 = ~n_1881 &  n_48340;
assign n_48342 = ~n_1875 &  n_48341;
assign n_48343 = ~n_1869 &  n_48342;
assign n_48344 = ~n_1863 &  n_48343;
assign n_48345 = ~n_1857 &  n_48344;
assign n_48346 = ~n_1851 &  n_48345;
assign n_48347 = ~n_1845 &  n_48346;
assign n_48348 = ~n_1839 &  n_48347;
assign n_48349 = ~n_1833 &  n_48348;
assign n_48350 = ~n_1827 &  n_48349;
assign n_48351 = ~n_1821 &  n_48350;
assign n_48352 = ~n_1815 &  n_48351;
assign n_48353 = ~n_1809 &  n_48352;
assign n_48354 = ~n_1803 &  n_48353;
assign n_48355 = ~n_1797 &  n_48354;
assign n_48356 = ~n_1791 &  n_48355;
assign n_48357 = ~n_1785 &  n_48356;
assign n_48358 = ~n_1779 &  n_48357;
assign n_48359 = ~n_1773 &  n_48358;
assign n_48360 = ~n_1767 &  n_48359;
assign n_48361 = ~n_1761 &  n_48360;
assign n_48362 = ~n_1755 &  n_48361;
assign n_48363 = ~n_1749 &  n_48362;
assign n_48364 = ~n_1743 &  n_48363;
assign n_48365 = ~n_1737 &  n_48364;
assign n_48366 = ~n_1731 &  n_48365;
assign n_48367 = ~n_1725 &  n_48366;
assign n_48368 = ~n_1719 &  n_48367;
assign n_48369 = ~n_1713 &  n_48368;
assign n_48370 = ~n_1707 &  n_48369;
assign n_48371 = ~n_1697 &  n_48370;
assign n_48372 = ~n_1691 &  n_48371;
assign n_48373 = ~n_1685 &  n_48372;
assign n_48374 = ~n_1679 &  n_48373;
assign n_48375 = ~n_1673 &  n_48374;
assign n_48376 = ~n_1667 &  n_48375;
assign n_48377 = ~n_1661 &  n_48376;
assign n_48378 = ~n_1655 &  n_48377;
assign n_48379 = ~n_1649 &  n_48378;
assign n_48380 = ~n_1643 &  n_48379;
assign n_48381 = ~n_1637 &  n_48380;
assign n_48382 = ~n_1631 &  n_48381;
assign n_48383 = ~n_1625 &  n_48382;
assign n_48384 = ~n_1619 &  n_48383;
assign n_48385 = ~n_1613 &  n_48384;
assign n_48386 = ~n_1607 &  n_48385;
assign n_48387 = ~n_1601 &  n_48386;
assign n_48388 = ~n_1595 &  n_48387;
assign n_48389 = ~n_1589 &  n_48388;
assign n_48390 = ~n_1583 &  n_48389;
assign n_48391 = ~n_1577 &  n_48390;
assign n_48392 = ~n_1571 &  n_48391;
assign n_48393 = ~n_1565 &  n_48392;
assign n_48394 = ~n_1559 &  n_48393;
assign n_48395 = ~n_1553 &  n_48394;
assign n_48396 = ~n_1547 &  n_48395;
assign n_48397 = ~n_1541 &  n_48396;
assign n_48398 = ~n_1535 &  n_48397;
assign n_48399 = ~n_1529 &  n_48398;
assign n_48400 = ~n_1523 &  n_48399;
assign n_48401 = ~n_1517 &  n_48400;
assign n_48402 = ~n_1511 &  n_48401;
assign n_48403 = ~n_1500 &  n_48402;
assign n_48404 = ~n_1494 &  n_48403;
assign n_48405 = ~n_1488 &  n_48404;
assign n_48406 = ~n_1482 &  n_48405;
assign n_48407 = ~n_1476 &  n_48406;
assign n_48408 = ~n_1470 &  n_48407;
assign n_48409 = ~n_1464 &  n_48408;
assign n_48410 = ~n_1458 &  n_48409;
assign n_48411 = ~n_1452 &  n_48410;
assign n_48412 = ~n_1446 &  n_48411;
assign n_48413 = ~n_1440 &  n_48412;
assign n_48414 = ~n_1434 &  n_48413;
assign n_48415 = ~n_1428 &  n_48414;
assign n_48416 = ~n_1422 &  n_48415;
assign n_48417 = ~n_1416 &  n_48416;
assign n_48418 = ~n_1410 &  n_48417;
assign n_48419 = ~n_1404 &  n_48418;
assign n_48420 = ~n_1398 &  n_48419;
assign n_48421 = ~n_1392 &  n_48420;
assign n_48422 = ~n_1386 &  n_48421;
assign n_48423 = ~n_1380 &  n_48422;
assign n_48424 = ~n_1374 &  n_48423;
assign n_48425 = ~n_1368 &  n_48424;
assign n_48426 = ~n_1362 &  n_48425;
assign n_48427 = ~n_1356 &  n_48426;
assign n_48428 = ~n_1350 &  n_48427;
assign n_48429 = ~n_1344 &  n_48428;
assign n_48430 = ~n_1338 &  n_48429;
assign n_48431 = ~n_1332 &  n_48430;
assign n_48432 = ~n_1326 &  n_48431;
assign n_48433 = ~n_1320 &  n_48432;
assign n_48434 = ~n_1314 &  n_48433;
assign n_48435 = ~n_1304 &  n_48434;
assign n_48436 = ~n_1300 &  n_48435;
assign n_48437 = ~n_1296 &  n_48436;
assign n_48438 = ~n_1292 &  n_48437;
assign n_48439 = ~n_1288 &  n_48438;
assign n_48440 = ~n_1284 &  n_48439;
assign n_48441 = ~n_1280 &  n_48440;
assign n_48442 = ~n_1276 &  n_48441;
assign n_48443 = ~n_1272 &  n_48442;
assign n_48444 = ~n_1268 &  n_48443;
assign n_48445 = ~n_1264 &  n_48444;
assign n_48446 = ~n_1260 &  n_48445;
assign n_48447 = ~n_1256 &  n_48446;
assign n_48448 = ~n_1252 &  n_48447;
assign n_48449 = ~n_1248 &  n_48448;
assign n_48450 = ~n_1244 &  n_48449;
assign n_48451 = ~n_1240 &  n_48450;
assign n_48452 = ~n_1236 &  n_48451;
assign n_48453 = ~n_1232 &  n_48452;
assign n_48454 = ~n_1228 &  n_48453;
assign n_48455 = ~n_1224 &  n_48454;
assign n_48456 = ~n_1220 &  n_48455;
assign n_48457 = ~n_1216 &  n_48456;
assign n_48458 = ~n_1212 &  n_48457;
assign n_48459 = ~n_1208 &  n_48458;
assign n_48460 = ~n_1204 &  n_48459;
assign n_48461 = ~n_1200 &  n_48460;
assign n_48462 = ~n_1196 &  n_48461;
assign n_48463 = ~n_1192 &  n_48462;
assign n_48464 = ~n_1188 &  n_48463;
assign n_48465 = ~n_1184 &  n_48464;
assign n_48466 = ~n_1180 &  n_48465;
assign n_48467 = ~n_1172 &  n_48466;
assign n_48468 = ~n_1168 &  n_48467;
assign n_48469 = ~n_1164 &  n_48468;
assign n_48470 = ~n_1160 &  n_48469;
assign n_48471 = ~n_1156 &  n_48470;
assign n_48472 = ~n_1152 &  n_48471;
assign n_48473 = ~n_1148 &  n_48472;
assign n_48474 = ~n_1144 &  n_48473;
assign n_48475 = ~n_1140 &  n_48474;
assign n_48476 = ~n_1136 &  n_48475;
assign n_48477 = ~n_1132 &  n_48476;
assign n_48478 = ~n_1128 &  n_48477;
assign n_48479 = ~n_1124 &  n_48478;
assign n_48480 = ~n_1120 &  n_48479;
assign n_48481 = ~n_1116 &  n_48480;
assign n_48482 = ~n_1112 &  n_48481;
assign n_48483 = ~n_1108 &  n_48482;
assign n_48484 = ~n_1104 &  n_48483;
assign n_48485 = ~n_1100 &  n_48484;
assign n_48486 = ~n_1096 &  n_48485;
assign n_48487 = ~n_1092 &  n_48486;
assign n_48488 = ~n_1088 &  n_48487;
assign n_48489 = ~n_1084 &  n_48488;
assign n_48490 = ~n_1080 &  n_48489;
assign n_48491 = ~n_1076 &  n_48490;
assign n_48492 = ~n_1072 &  n_48491;
assign n_48493 = ~n_1068 &  n_48492;
assign n_48494 = ~n_1064 &  n_48493;
assign n_48495 = ~n_1060 &  n_48494;
assign n_48496 = ~n_1056 &  n_48495;
assign n_48497 = ~n_1052 &  n_48496;
assign n_48498 = ~n_1048 &  n_48497;
assign n_48499 = ~n_1036 &  n_48498;
assign n_48500 = ~n_1032 &  n_48499;
assign n_48501 = ~n_1028 &  n_48500;
assign n_48502 = ~n_1024 &  n_48501;
assign n_48503 = ~n_1020 &  n_48502;
assign n_48504 = ~n_1016 &  n_48503;
assign n_48505 = ~n_1012 &  n_48504;
assign n_48506 = ~n_1008 &  n_48505;
assign n_48507 = ~n_1004 &  n_48506;
assign n_48508 = ~n_1000 &  n_48507;
assign n_48509 = ~n_996 &  n_48508;
assign n_48510 = ~n_992 &  n_48509;
assign n_48511 = ~n_988 &  n_48510;
assign n_48512 = ~n_984 &  n_48511;
assign n_48513 = ~n_980 &  n_48512;
assign n_48514 = ~n_976 &  n_48513;
assign n_48515 = ~n_972 &  n_48514;
assign n_48516 = ~n_968 &  n_48515;
assign n_48517 = ~n_964 &  n_48516;
assign n_48518 = ~n_960 &  n_48517;
assign n_48519 = ~n_956 &  n_48518;
assign n_48520 = ~n_952 &  n_48519;
assign n_48521 = ~n_947 &  n_48520;
assign n_48522 = ~n_943 &  n_48521;
assign n_48523 = ~n_938 &  n_48522;
assign n_48524 = ~n_934 &  n_48523;
assign n_48525 = ~n_929 &  n_48524;
assign n_48526 = ~n_924 &  n_48525;
assign n_48527 = ~n_919 &  n_48526;
assign n_48528 = ~n_914 &  n_48527;
assign n_48529 = ~n_910 &  n_48528;
assign n_48530 = ~n_905 &  n_48529;
assign n_48531 = ~n_755 &  n_48530;
assign n_48532 = ~n_749 &  n_48531;
assign n_48533 = ~n_743 &  n_48532;
assign n_48534 = ~n_737 &  n_48533;
assign n_48535 = ~n_731 &  n_48534;
assign n_48536 = ~n_725 &  n_48535;
assign n_48537 = ~n_719 &  n_48536;
assign n_48538 = ~n_713 &  n_48537;
assign n_48539 = ~n_707 &  n_48538;
assign n_48540 = ~n_701 &  n_48539;
assign n_48541 = ~n_695 &  n_48540;
assign n_48542 = ~n_689 &  n_48541;
assign n_48543 = ~n_683 &  n_48542;
assign n_48544 = ~n_677 &  n_48543;
assign n_48545 = ~n_671 &  n_48544;
assign n_48546 = ~n_665 &  n_48545;
assign n_48547 = ~n_659 &  n_48546;
assign n_48548 = ~n_653 &  n_48547;
assign n_48549 = ~n_647 &  n_48548;
assign n_48550 = ~n_641 &  n_48549;
assign n_48551 = ~n_635 &  n_48550;
assign n_48552 = ~n_629 &  n_48551;
assign n_48553 = ~n_623 &  n_48552;
assign n_48554 = ~n_617 &  n_48553;
assign n_48555 = ~n_611 &  n_48554;
assign n_48556 = ~n_605 &  n_48555;
assign n_48557 = ~n_599 &  n_48556;
assign n_48558 = ~n_593 &  n_48557;
assign n_48559 = ~n_587 &  n_48558;
assign n_48560 = ~n_581 &  n_48559;
assign n_48561 = ~n_575 &  n_48560;
assign n_48562 = ~n_569 &  n_48561;
assign n_48563 = ~n_550 &  n_48562;
assign n_48564 = ~n_544 &  n_48563;
assign n_48565 = ~n_538 &  n_48564;
assign n_48566 = ~n_532 &  n_48565;
assign n_48567 = ~n_526 &  n_48566;
assign n_48568 = ~n_520 &  n_48567;
assign n_48569 = ~n_514 &  n_48568;
assign n_48570 = ~n_508 &  n_48569;
assign n_48571 = ~n_502 &  n_48570;
assign n_48572 = ~n_496 &  n_48571;
assign n_48573 = ~n_490 &  n_48572;
assign n_48574 = ~n_484 &  n_48573;
assign n_48575 = ~n_478 &  n_48574;
assign n_48576 = ~n_472 &  n_48575;
assign n_48577 = ~n_466 &  n_48576;
assign n_48578 = ~n_460 &  n_48577;
assign n_48579 = ~n_454 &  n_48578;
assign n_48580 = ~n_448 &  n_48579;
assign n_48581 = ~n_442 &  n_48580;
assign n_48582 = ~n_436 &  n_48581;
assign n_48583 = ~n_430 &  n_48582;
assign n_48584 = ~n_424 &  n_48583;
assign n_48585 = ~n_418 &  n_48584;
assign n_48586 = ~n_412 &  n_48585;
assign n_48587 = ~n_406 &  n_48586;
assign n_48588 = ~n_400 &  n_48587;
assign n_48589 = ~n_394 &  n_48588;
assign n_48590 = ~n_388 &  n_48589;
assign n_48591 = ~n_382 &  n_48590;
assign n_48592 = ~n_376 &  n_48591;
assign n_48593 = ~n_370 &  n_48592;
assign n_48594 = ~n_364 &  n_48593;
assign n_48595 = ~n_348 &  n_48594;
assign n_48596 = ~n_342 &  n_48595;
assign n_48597 = ~n_336 &  n_48596;
assign n_48598 = ~n_330 &  n_48597;
assign n_48599 = ~n_324 &  n_48598;
assign n_48600 = ~n_318 &  n_48599;
assign n_48601 = ~n_312 &  n_48600;
assign n_48602 = ~n_306 &  n_48601;
assign n_48603 = ~n_300 &  n_48602;
assign n_48604 = ~n_294 &  n_48603;
assign n_48605 = ~n_288 &  n_48604;
assign n_48606 = ~n_282 &  n_48605;
assign n_48607 = ~n_276 &  n_48606;
assign n_48608 = ~n_270 &  n_48607;
assign n_48609 = ~n_264 &  n_48608;
assign n_48610 = ~n_258 &  n_48609;
assign n_48611 = ~n_252 &  n_48610;
assign n_48612 = ~n_246 &  n_48611;
assign n_48613 = ~n_240 &  n_48612;
assign n_48614 = ~n_234 &  n_48613;
assign n_48615 = ~n_228 &  n_48614;
assign n_48616 = ~n_222 &  n_48615;
assign n_48617 = ~n_216 &  n_48616;
assign n_48618 = ~n_210 &  n_48617;
assign n_48619 = ~n_204 &  n_48618;
assign n_48620 = ~n_198 &  n_48619;
assign n_48621 = ~n_192 &  n_48620;
assign n_48622 = ~n_186 &  n_48621;
assign n_48623 = ~n_180 &  n_48622;
assign n_48624 = ~n_174 &  n_48623;
assign n_48625 = ~n_168 &  n_48624;
assign n_48626 = ~n_162 &  n_48625;
assign n_48627 = ~n_146 &  n_48626;
assign n_48628 = ~n_142 &  n_48627;
assign n_48629 = ~n_138 &  n_48628;
assign n_48630 = ~n_134 &  n_48629;
assign n_48631 = ~n_130 &  n_48630;
assign n_48632 = ~n_126 &  n_48631;
assign n_48633 = ~n_122 &  n_48632;
assign n_48634 = ~n_118 &  n_48633;
assign n_48635 = ~n_114 &  n_48634;
assign n_48636 = ~n_110 &  n_48635;
assign n_48637 = ~n_106 &  n_48636;
assign n_48638 = ~n_102 &  n_48637;
assign n_48639 = ~n_98 &  n_48638;
assign n_48640 = ~n_94 &  n_48639;
assign n_48641 = ~n_90 &  n_48640;
assign n_48642 = ~n_86 &  n_48641;
assign n_48643 = ~n_82 &  n_48642;
assign n_48644 = ~n_78 &  n_48643;
assign n_48645 = ~n_74 &  n_48644;
assign n_48646 = ~n_70 &  n_48645;
assign n_48647 = ~n_66 &  n_48646;
assign n_48648 = ~n_62 &  n_48647;
assign n_48649 = ~n_58 &  n_48648;
assign n_48650 = ~n_54 &  n_48649;
assign n_48651 = ~n_50 &  n_48650;
assign n_48652 = ~n_46 &  n_48651;
assign n_48653 = ~n_42 &  n_48652;
assign n_48654 = ~n_38 &  n_48653;
assign n_48655 = ~n_34 &  n_48654;
assign n_48656 = ~n_30 &  n_48655;
assign n_48657 = ~n_26 &  n_48656;
assign n_48658 = ~n_22 &  n_48657;
assign o_1 = ~n_48658;
endmodule

