// test verilog file
module factorization8_simplified (x1,x2);
input x1;
input x2;
output o1;
assign o1 =  ~x1 & x2;
endmodule
