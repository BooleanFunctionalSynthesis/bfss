// Generated using findDep.cpp 
module small-swap2-fixpoint-6 (v_1, v_2, v_3, v_4, v_5, v_6, v_7, v_8, v_9, v_10, v_11, v_12, v_13, v_14, v_15, v_16, v_17, v_18, v_19, v_20, v_21, v_22, v_23, v_24, v_25, v_26, v_27, v_28, v_29, v_30, v_31, v_32, v_33, v_34, v_35, v_36, v_37, v_38, v_39, v_40, v_41, v_42, v_43, v_44, v_45, v_46, v_47, v_48, v_49, v_50, v_51, v_52, v_53, v_54, v_55, v_56, v_57, v_58, v_59, v_60, v_61, v_62, v_63, v_64, v_65, v_66, v_67, v_68, v_69, v_70, v_71, v_72, v_73, v_74, v_75, v_76, v_77, v_78, v_79, v_80, v_81, v_82, v_83, v_84, v_85, v_86, v_87, v_88, v_89, v_90, v_91, v_92, v_93, v_94, v_95, v_96, v_97, v_98, v_99, v_100, v_101, v_102, v_103, v_104, v_105, v_106, v_107, v_108, v_109, v_110, v_111, v_112, v_113, v_114, v_115, v_116, v_117, v_118, v_119, v_120, v_121, v_122, v_123, v_124, v_125, v_126, v_127, v_128, v_129, v_130, v_131, v_132, v_133, v_134, v_135, v_136, v_137, v_138, v_139, v_140, v_141, v_142, v_143, v_144, v_145, v_146, v_147, v_148, v_149, v_150, v_151, v_152, v_153, v_154, v_155, v_156, v_157, v_158, v_159, v_160, v_161, v_162, v_163, v_164, v_165, v_166, v_167, v_168, v_169, v_170, v_171, v_172, v_173, v_174, v_175, v_176, v_177, v_178, v_179, v_180, v_181, v_182, v_183, v_184, v_185, v_186, v_187, v_188, v_189, v_190, v_191, v_192, v_193, v_194, v_195, v_196, v_197, v_198, v_199, v_200, v_201, v_202, v_203, v_204, v_205, v_206, v_207, v_208, v_209, v_210, v_211, v_212, v_213, v_214, v_215, v_216, v_217, v_218, v_219, v_220, v_221, v_222, v_223, v_224, v_225, v_226, v_227, v_228, v_229, v_230, v_231, v_232, v_233, v_234, v_235, v_236, v_237, v_238, v_239, v_240, v_241, v_242, v_243, v_244, v_245, v_246, v_247, v_248, v_249, v_250, v_251, v_252, v_253, v_254, v_255, v_256, v_257, v_258, v_259, v_260, v_261, v_262, v_263, v_264, v_265, v_266, v_267, v_268, v_269, v_270, v_271, v_272, v_273, v_274, v_275, v_276, v_277, v_278, v_279, v_280, v_281, v_282, v_283, v_284, v_285, v_286, v_287, v_288, v_289, v_290, v_291, v_292, v_293, v_294, v_295, v_296, v_297, v_298, v_299, v_300, v_301, v_302, v_303, v_304, v_305, v_306, v_307, v_308, v_309, v_310, v_311, v_312, v_313, v_314, v_315, v_316, v_317, v_318, v_319, v_320, v_321, v_322, v_323, v_324, v_325, v_326, v_327, v_328, v_329, v_330, v_331, v_332, v_333, v_334, v_335, v_336, v_337, v_338, v_339, v_340, v_341, v_342, v_343, v_344, v_345, v_346, v_347, v_348, v_349, v_350, v_351, v_352, v_353, v_354, v_355, v_356, v_357, v_358, v_359, v_360, v_361, v_362, v_363, v_364, v_365, v_366, v_367, v_368, v_369, v_370, v_371, v_372, v_373, v_374, v_375, v_376, v_377, v_378, v_379, v_380, v_381, v_382, v_383, v_384, v_385, v_386, v_387, v_388, v_389, v_390, v_391, v_392, v_393, v_394, v_395, v_396, v_397, v_398, v_399, v_400, v_401, v_402, v_403, v_404, v_405, v_406, v_407, v_408, v_409, v_410, v_411, v_412, v_413, v_414, v_415, v_416, v_417, v_418, v_419, v_420, v_421, v_422, v_423, v_424, v_425, v_426, v_427, v_428, v_429, v_430, v_431, v_432, v_433, v_434, v_435, v_436, v_437, v_438, v_439, v_440, v_441, v_442, v_443, v_444, v_445, v_446, v_447, v_448, v_449, v_450, v_451, v_452, v_453, v_454, v_455, v_456, v_457, v_458, v_459, v_460, v_461, v_462, v_463, v_464, v_465, v_466, v_467, v_468, v_469, v_470, v_471, v_472, v_473, v_474, v_475, v_476, v_477, v_478, v_479, v_480, v_481, v_482, v_483, v_484, v_485, v_486, v_487, v_488, v_489, v_490, v_491, v_492, v_493, v_494, v_495, v_496, v_497, v_498, v_499, v_500, v_501, v_502, v_503, v_504, v_505, v_506, v_507, v_508, v_509, v_510, v_511, v_512, v_513, v_514, v_515, v_516, v_517, v_518, v_519, v_520, v_521, v_522, v_523, v_524, v_525, v_526, v_527, v_528, v_529, v_530, v_531, v_532, v_533, v_534, v_535, v_536, v_537, v_538, v_539, v_540, v_541, v_542, v_543, v_544, v_545, v_546, v_547, v_548, v_549, v_550, v_551, v_552, v_553, v_554, v_555, v_556, v_557, v_558, v_559, v_560, v_561, v_562, v_563, v_564, v_565, v_566, v_567, v_568, v_569, v_570, v_571, v_572, v_573, v_574, v_575, v_576, v_577, v_578, v_579, v_580, v_581, v_582, v_583, v_584, v_585, v_586, v_587, v_588, v_589, v_590, v_591, v_592, v_593, v_594, v_595, v_596, v_597, v_598, v_599, v_600, v_601, v_602, v_603, v_604, v_605, v_606, v_607, v_608, v_609, v_610, v_611, v_612, v_613, v_614, v_615, v_616, v_617, v_618, v_619, v_620, v_621, v_622, v_623, v_624, v_625, v_626, v_627, v_628, v_629, v_630, v_631, v_632, v_633, v_634, v_635, v_636, v_637, v_638, v_639, v_640, v_641, v_642, v_643, v_644, v_645, v_646, v_647, v_648, v_649, v_650, v_651, v_652, v_653, v_654, v_655, v_656, v_657, v_658, v_659, v_660, v_661, v_662, v_663, v_664, v_665, v_666, v_667, v_668, v_669, v_670, v_671, v_672, v_673, v_674, v_675, v_676, v_677, v_678, v_679, v_680, v_681, v_682, v_683, v_684, v_685, v_686, v_687, v_688, v_689, v_690, v_691, v_692, v_693, v_694, v_695, v_696, v_697, v_698, v_699, v_700, v_701, v_702, v_703, v_704, v_705, v_706, v_707, v_708, v_709, v_710, v_711, v_712, v_713, v_714, v_715, v_716, v_717, v_718, v_719, v_720, v_721, v_722, v_723, v_724, v_725, v_726, v_727, v_728, v_729, v_730, v_731, v_732, v_733, v_734, v_735, v_736, v_737, v_738, v_739, v_740, v_741, v_742, v_743, v_744, v_745, v_746, v_747, v_748, v_749, v_750, v_751, v_752, v_753, v_754, v_755, v_756, v_757, v_758, v_759, v_760, v_761, v_762, v_763, v_764, v_765, v_766, v_767, v_768, v_769, v_770, v_771, v_772, v_773, v_774, v_775, v_776, v_777, v_778, v_779, v_780, o_1);
input v_1;
input v_2;
input v_3;
input v_4;
input v_5;
input v_6;
input v_7;
input v_8;
input v_9;
input v_10;
input v_11;
input v_12;
input v_13;
input v_14;
input v_15;
input v_16;
input v_17;
input v_18;
input v_19;
input v_20;
input v_21;
input v_22;
input v_23;
input v_24;
input v_25;
input v_26;
input v_27;
input v_28;
input v_29;
input v_30;
input v_31;
input v_32;
input v_33;
input v_34;
input v_35;
input v_36;
input v_37;
input v_38;
input v_39;
input v_40;
input v_41;
input v_42;
input v_43;
input v_44;
input v_45;
input v_46;
input v_47;
input v_48;
input v_49;
input v_50;
input v_51;
input v_52;
input v_53;
input v_54;
input v_55;
input v_56;
input v_57;
input v_58;
input v_59;
input v_60;
input v_61;
input v_62;
input v_63;
input v_64;
input v_65;
input v_66;
input v_67;
input v_68;
input v_69;
input v_70;
input v_71;
input v_72;
input v_73;
input v_74;
input v_75;
input v_76;
input v_77;
input v_78;
input v_79;
input v_80;
input v_81;
input v_82;
input v_83;
input v_84;
input v_85;
input v_86;
input v_87;
input v_88;
input v_89;
input v_90;
input v_91;
input v_92;
input v_93;
input v_94;
input v_95;
input v_96;
input v_97;
input v_98;
input v_99;
input v_100;
input v_101;
input v_102;
input v_103;
input v_104;
input v_105;
input v_106;
input v_107;
input v_108;
input v_109;
input v_110;
input v_111;
input v_112;
input v_113;
input v_114;
input v_115;
input v_116;
input v_117;
input v_118;
input v_119;
input v_120;
input v_121;
input v_122;
input v_123;
input v_124;
input v_125;
input v_126;
input v_127;
input v_128;
input v_129;
input v_130;
input v_131;
input v_132;
input v_133;
input v_134;
input v_135;
input v_136;
input v_137;
input v_138;
input v_139;
input v_140;
input v_141;
input v_142;
input v_143;
input v_144;
input v_145;
input v_146;
input v_147;
input v_148;
input v_149;
input v_150;
input v_151;
input v_152;
input v_153;
input v_154;
input v_155;
input v_156;
input v_157;
input v_158;
input v_159;
input v_160;
input v_161;
input v_162;
input v_163;
input v_164;
input v_165;
input v_166;
input v_167;
input v_168;
input v_169;
input v_170;
input v_171;
input v_172;
input v_173;
input v_174;
input v_175;
input v_176;
input v_177;
input v_178;
input v_179;
input v_180;
input v_181;
input v_182;
input v_183;
input v_184;
input v_185;
input v_186;
input v_187;
input v_188;
input v_189;
input v_190;
input v_191;
input v_192;
input v_193;
input v_194;
input v_195;
input v_196;
input v_197;
input v_198;
input v_199;
input v_200;
input v_201;
input v_202;
input v_203;
input v_204;
input v_205;
input v_206;
input v_207;
input v_208;
input v_209;
input v_210;
input v_211;
input v_212;
input v_213;
input v_214;
input v_215;
input v_216;
input v_217;
input v_218;
input v_219;
input v_220;
input v_221;
input v_222;
input v_223;
input v_224;
input v_225;
input v_226;
input v_227;
input v_228;
input v_229;
input v_230;
input v_231;
input v_232;
input v_233;
input v_234;
input v_235;
input v_236;
input v_237;
input v_238;
input v_239;
input v_240;
input v_241;
input v_242;
input v_243;
input v_244;
input v_245;
input v_246;
input v_247;
input v_248;
input v_249;
input v_250;
input v_251;
input v_252;
input v_253;
input v_254;
input v_255;
input v_256;
input v_257;
input v_258;
input v_259;
input v_260;
input v_261;
input v_262;
input v_263;
input v_264;
input v_265;
input v_266;
input v_267;
input v_268;
input v_269;
input v_270;
input v_271;
input v_272;
input v_273;
input v_274;
input v_275;
input v_276;
input v_277;
input v_278;
input v_279;
input v_280;
input v_281;
input v_282;
input v_283;
input v_284;
input v_285;
input v_286;
input v_287;
input v_288;
input v_289;
input v_290;
input v_291;
input v_292;
input v_293;
input v_294;
input v_295;
input v_296;
input v_297;
input v_298;
input v_299;
input v_300;
input v_301;
input v_302;
input v_303;
input v_304;
input v_305;
input v_306;
input v_307;
input v_308;
input v_309;
input v_310;
input v_311;
input v_312;
input v_313;
input v_314;
input v_315;
input v_316;
input v_317;
input v_318;
input v_319;
input v_320;
input v_321;
input v_322;
input v_323;
input v_324;
input v_325;
input v_326;
input v_327;
input v_328;
input v_329;
input v_330;
input v_331;
input v_332;
input v_333;
input v_334;
input v_335;
input v_336;
input v_337;
input v_338;
input v_339;
input v_340;
input v_341;
input v_342;
input v_343;
input v_344;
input v_345;
input v_346;
input v_347;
input v_348;
input v_349;
input v_350;
input v_351;
input v_352;
input v_353;
input v_354;
input v_355;
input v_356;
input v_357;
input v_358;
input v_359;
input v_360;
input v_361;
input v_362;
input v_363;
input v_364;
input v_365;
input v_366;
input v_367;
input v_368;
input v_369;
input v_370;
input v_371;
input v_372;
input v_373;
input v_374;
input v_375;
input v_376;
input v_377;
input v_378;
input v_379;
input v_380;
input v_381;
input v_382;
input v_383;
input v_384;
input v_385;
input v_386;
input v_387;
input v_388;
input v_389;
input v_390;
input v_391;
input v_392;
input v_393;
input v_394;
input v_395;
input v_396;
input v_397;
input v_398;
input v_399;
input v_400;
input v_401;
input v_402;
input v_403;
input v_404;
input v_405;
input v_406;
input v_407;
input v_408;
input v_409;
input v_410;
input v_411;
input v_412;
input v_413;
input v_414;
input v_415;
input v_416;
input v_417;
input v_418;
input v_419;
input v_420;
input v_421;
input v_422;
input v_423;
input v_424;
input v_425;
input v_426;
input v_427;
input v_428;
input v_429;
input v_430;
input v_431;
input v_432;
input v_433;
input v_434;
input v_435;
input v_436;
input v_437;
input v_438;
input v_439;
input v_440;
input v_441;
input v_442;
input v_443;
input v_444;
input v_445;
input v_446;
input v_447;
input v_448;
input v_449;
input v_450;
input v_451;
input v_452;
input v_453;
input v_454;
input v_455;
input v_456;
input v_457;
input v_458;
input v_459;
input v_460;
input v_461;
input v_462;
input v_463;
input v_464;
input v_465;
input v_466;
input v_467;
input v_468;
input v_469;
input v_470;
input v_471;
input v_472;
input v_473;
input v_474;
input v_475;
input v_476;
input v_477;
input v_478;
input v_479;
input v_480;
input v_481;
input v_482;
input v_483;
input v_484;
input v_485;
input v_486;
input v_487;
input v_488;
input v_489;
input v_490;
input v_491;
input v_492;
input v_493;
input v_494;
input v_495;
input v_496;
input v_497;
input v_498;
input v_499;
input v_500;
input v_501;
input v_502;
input v_503;
input v_504;
input v_505;
input v_506;
input v_507;
input v_508;
input v_509;
input v_510;
input v_511;
input v_512;
input v_513;
input v_514;
input v_515;
input v_516;
input v_517;
input v_518;
input v_519;
input v_520;
input v_521;
input v_522;
input v_523;
input v_524;
input v_525;
input v_526;
input v_527;
input v_528;
input v_529;
input v_530;
input v_531;
input v_532;
input v_533;
input v_534;
input v_535;
input v_536;
input v_537;
input v_538;
input v_539;
input v_540;
input v_541;
input v_542;
input v_543;
input v_544;
input v_545;
input v_546;
input v_547;
input v_548;
input v_549;
input v_550;
input v_551;
input v_552;
input v_553;
input v_554;
input v_555;
input v_556;
input v_557;
input v_558;
input v_559;
input v_560;
input v_561;
input v_562;
input v_563;
input v_564;
input v_565;
input v_566;
input v_567;
input v_568;
input v_569;
input v_570;
input v_571;
input v_572;
input v_573;
input v_574;
input v_575;
input v_576;
input v_577;
input v_578;
input v_579;
input v_580;
input v_581;
input v_582;
input v_583;
input v_584;
input v_585;
input v_586;
input v_587;
input v_588;
input v_589;
input v_590;
input v_591;
input v_592;
input v_593;
input v_594;
input v_595;
input v_596;
input v_597;
input v_598;
input v_599;
input v_600;
input v_601;
input v_602;
input v_603;
input v_604;
input v_605;
input v_606;
input v_607;
input v_608;
input v_609;
input v_610;
input v_611;
input v_612;
input v_613;
input v_614;
input v_615;
input v_616;
input v_617;
input v_618;
input v_619;
input v_620;
input v_621;
input v_622;
input v_623;
input v_624;
input v_625;
input v_626;
input v_627;
input v_628;
input v_629;
input v_630;
input v_631;
input v_632;
input v_633;
input v_634;
input v_635;
input v_636;
input v_637;
input v_638;
input v_639;
input v_640;
input v_641;
input v_642;
input v_643;
input v_644;
input v_645;
input v_646;
input v_647;
input v_648;
input v_649;
input v_650;
input v_651;
input v_652;
input v_653;
input v_654;
input v_655;
input v_656;
input v_657;
input v_658;
input v_659;
input v_660;
input v_661;
input v_662;
input v_663;
input v_664;
input v_665;
input v_666;
input v_667;
input v_668;
input v_669;
input v_670;
input v_671;
input v_672;
input v_673;
input v_674;
input v_675;
input v_676;
input v_677;
input v_678;
input v_679;
input v_680;
input v_681;
input v_682;
input v_683;
input v_684;
input v_685;
input v_686;
input v_687;
input v_688;
input v_689;
input v_690;
input v_691;
input v_692;
input v_693;
input v_694;
input v_695;
input v_696;
input v_697;
input v_698;
input v_699;
input v_700;
input v_701;
input v_702;
input v_703;
input v_704;
input v_705;
input v_706;
input v_707;
input v_708;
input v_709;
input v_710;
input v_711;
input v_712;
input v_713;
input v_714;
input v_715;
input v_716;
input v_717;
input v_718;
input v_719;
input v_720;
input v_721;
input v_722;
input v_723;
input v_724;
input v_725;
input v_726;
input v_727;
input v_728;
input v_729;
input v_730;
input v_731;
input v_732;
input v_733;
input v_734;
input v_735;
input v_736;
input v_737;
input v_738;
input v_739;
input v_740;
input v_741;
input v_742;
input v_743;
input v_744;
input v_745;
input v_746;
input v_747;
input v_748;
input v_749;
input v_750;
input v_751;
input v_752;
input v_753;
input v_754;
input v_755;
input v_756;
input v_757;
input v_758;
input v_759;
input v_760;
input v_761;
input v_762;
input v_763;
input v_764;
input v_765;
input v_766;
input v_767;
input v_768;
input v_769;
input v_770;
input v_771;
input v_772;
input v_773;
input v_774;
input v_775;
input v_776;
input v_777;
input v_778;
input v_779;
input v_780;
output o_1;
wire v_781;
wire v_782;
wire v_783;
wire v_784;
wire v_785;
wire v_786;
wire v_787;
wire v_788;
wire v_789;
wire v_790;
wire v_791;
wire v_792;
wire v_793;
wire v_794;
wire v_795;
wire v_796;
wire v_797;
wire v_798;
wire v_799;
wire v_800;
wire v_801;
wire v_802;
wire v_803;
wire v_804;
wire v_805;
wire v_806;
wire v_807;
wire v_808;
wire v_809;
wire v_810;
wire v_811;
wire v_812;
wire v_813;
wire v_814;
wire v_815;
wire v_816;
wire v_817;
wire v_818;
wire v_819;
wire v_820;
wire v_821;
wire v_822;
wire v_823;
wire v_824;
wire v_825;
wire v_826;
wire v_827;
wire v_828;
wire v_829;
wire v_830;
wire v_831;
wire v_832;
wire v_833;
wire v_834;
wire v_835;
wire v_836;
wire v_837;
wire v_838;
wire v_839;
wire v_840;
wire v_841;
wire v_842;
wire v_843;
wire v_844;
wire v_845;
wire v_846;
wire v_847;
wire v_848;
wire v_849;
wire v_850;
wire v_851;
wire v_852;
wire v_853;
wire v_854;
wire v_855;
wire v_856;
wire v_857;
wire v_858;
wire v_859;
wire v_860;
wire v_861;
wire v_862;
wire v_863;
wire v_864;
wire v_865;
wire v_866;
wire v_867;
wire v_868;
wire v_869;
wire v_870;
wire v_871;
wire v_872;
wire v_873;
wire v_874;
wire v_875;
wire v_876;
wire v_877;
wire v_878;
wire v_879;
wire v_880;
wire v_881;
wire v_882;
wire v_883;
wire v_884;
wire v_885;
wire v_886;
wire v_887;
wire v_888;
wire v_889;
wire v_890;
wire v_891;
wire v_892;
wire v_893;
wire v_894;
wire v_895;
wire v_896;
wire v_897;
wire v_898;
wire v_899;
wire v_900;
wire v_901;
wire v_902;
wire v_903;
wire v_904;
wire v_905;
wire v_906;
wire v_907;
wire v_908;
wire v_909;
wire v_910;
wire v_911;
wire v_912;
wire v_913;
wire v_914;
wire v_915;
wire v_916;
wire v_917;
wire v_918;
wire v_919;
wire v_920;
wire v_921;
wire v_922;
wire v_923;
wire v_924;
wire v_925;
wire v_926;
wire v_927;
wire v_928;
wire v_929;
wire v_930;
wire v_931;
wire v_932;
wire v_933;
wire v_934;
wire v_935;
wire v_936;
wire v_937;
wire v_938;
wire v_939;
wire v_940;
wire v_941;
wire v_942;
wire v_943;
wire v_944;
wire v_945;
wire v_946;
wire v_947;
wire v_948;
wire v_949;
wire v_950;
wire v_951;
wire v_952;
wire v_953;
wire v_954;
wire v_955;
wire v_956;
wire v_957;
wire v_958;
wire v_959;
wire v_960;
wire v_961;
wire v_962;
wire v_963;
wire v_964;
wire v_965;
wire v_966;
wire v_967;
wire v_968;
wire v_969;
wire v_970;
wire v_971;
wire v_972;
wire v_973;
wire v_974;
wire v_975;
wire v_976;
wire v_977;
wire v_978;
wire v_979;
wire v_980;
wire v_981;
wire v_982;
wire v_983;
wire v_984;
wire v_985;
wire v_986;
wire v_987;
wire v_988;
wire v_989;
wire v_990;
wire v_991;
wire v_992;
wire v_993;
wire v_994;
wire v_995;
wire v_996;
wire v_997;
wire v_998;
wire v_999;
wire v_1000;
wire v_1001;
wire v_1002;
wire v_1003;
wire v_1004;
wire v_1005;
wire v_1006;
wire v_1007;
wire v_1008;
wire v_1009;
wire v_1010;
wire v_1011;
wire v_1012;
wire v_1013;
wire v_1014;
wire v_1015;
wire v_1016;
wire v_1017;
wire v_1018;
wire v_1019;
wire v_1020;
wire v_1021;
wire v_1022;
wire v_1023;
wire v_1024;
wire v_1025;
wire v_1026;
wire v_1027;
wire v_1028;
wire v_1029;
wire v_1030;
wire v_1031;
wire v_1032;
wire v_1033;
wire v_1034;
wire v_1035;
wire v_1036;
wire v_1037;
wire v_1038;
wire v_1039;
wire v_1040;
wire v_1041;
wire v_1042;
wire v_1043;
wire v_1044;
wire v_1045;
wire v_1046;
wire v_1047;
wire v_1048;
wire v_1049;
wire v_1050;
wire v_1051;
wire v_1052;
wire v_1053;
wire v_1054;
wire v_1055;
wire v_1056;
wire v_1057;
wire v_1058;
wire v_1059;
wire v_1060;
wire v_1061;
wire v_1062;
wire v_1063;
wire v_1064;
wire v_1065;
wire v_1066;
wire v_1067;
wire v_1068;
wire v_1069;
wire v_1070;
wire v_1071;
wire v_1072;
wire v_1073;
wire v_1074;
wire v_1075;
wire v_1076;
wire v_1077;
wire v_1078;
wire v_1079;
wire v_1080;
wire v_1081;
wire v_1082;
wire v_1083;
wire v_1084;
wire v_1085;
wire v_1086;
wire v_1087;
wire v_1088;
wire v_1089;
wire v_1090;
wire v_1091;
wire v_1092;
wire v_1093;
wire v_1094;
wire v_1095;
wire v_1096;
wire v_1097;
wire v_1098;
wire v_1099;
wire v_1100;
wire v_1101;
wire v_1102;
wire v_1103;
wire v_1104;
wire v_1105;
wire v_1106;
wire v_1107;
wire v_1108;
wire v_1109;
wire v_1110;
wire v_1111;
wire v_1112;
wire v_1113;
wire v_1114;
wire v_1115;
wire v_1116;
wire v_1117;
wire v_1118;
wire v_1119;
wire v_1120;
wire v_1121;
wire v_1122;
wire v_1123;
wire v_1124;
wire v_1125;
wire v_1126;
wire v_1127;
wire v_1128;
wire v_1129;
wire v_1130;
wire v_1131;
wire v_1132;
wire v_1133;
wire v_1134;
wire v_1135;
wire v_1136;
wire v_1137;
wire v_1138;
wire v_1139;
wire v_1140;
wire v_1141;
wire v_1142;
wire v_1143;
wire v_1144;
wire v_1145;
wire v_1146;
wire v_1147;
wire v_1148;
wire v_1149;
wire v_1150;
wire v_1151;
wire v_1152;
wire v_1153;
wire v_1154;
wire v_1155;
wire v_1156;
wire v_1157;
wire v_1158;
wire v_1159;
wire v_1160;
wire v_1161;
wire v_1162;
wire v_1163;
wire v_1164;
wire v_1165;
wire v_1166;
wire v_1167;
wire v_1168;
wire v_1169;
wire v_1170;
wire v_1171;
wire v_1172;
wire v_1173;
wire v_1174;
wire v_1175;
wire v_1176;
wire v_1177;
wire v_1178;
wire v_1179;
wire v_1180;
wire v_1181;
wire v_1182;
wire v_1183;
wire v_1184;
wire v_1185;
wire v_1186;
wire v_1187;
wire v_1188;
wire v_1189;
wire v_1190;
wire v_1191;
wire v_1192;
wire v_1193;
wire v_1194;
wire v_1195;
wire v_1196;
wire v_1197;
wire v_1198;
wire v_1199;
wire v_1200;
wire v_1201;
wire v_1202;
wire v_1203;
wire v_1204;
wire v_1205;
wire v_1206;
wire v_1207;
wire v_1208;
wire v_1209;
wire v_1210;
wire v_1211;
wire v_1212;
wire v_1213;
wire v_1214;
wire v_1215;
wire v_1216;
wire v_1217;
wire v_1218;
wire v_1219;
wire v_1220;
wire v_1221;
wire v_1222;
wire v_1223;
wire v_1224;
wire v_1225;
wire v_1226;
wire v_1227;
wire v_1228;
wire v_1229;
wire v_1230;
wire v_1231;
wire v_1232;
wire v_1233;
wire v_1234;
wire v_1235;
wire v_1236;
wire v_1237;
wire v_1238;
wire v_1239;
wire v_1240;
wire v_1241;
wire v_1242;
wire v_1243;
wire v_1244;
wire v_1245;
wire v_1246;
wire v_1247;
wire v_1248;
wire v_1249;
wire v_1250;
wire v_1251;
wire v_1252;
wire v_1253;
wire v_1254;
wire v_1255;
wire v_1256;
wire v_1257;
wire v_1258;
wire v_1259;
wire v_1260;
wire v_1261;
wire v_1262;
wire v_1263;
wire v_1264;
wire v_1265;
wire v_1266;
wire v_1267;
wire v_1268;
wire v_1269;
wire v_1270;
wire v_1271;
wire v_1272;
wire v_1273;
wire v_1274;
wire v_1275;
wire v_1276;
wire v_1277;
wire v_1278;
wire v_1279;
wire v_1280;
wire v_1281;
wire v_1282;
wire v_1283;
wire v_1284;
wire v_1285;
wire v_1286;
wire v_1287;
wire v_1288;
wire v_1289;
wire v_1290;
wire v_1291;
wire v_1292;
wire v_1293;
wire v_1294;
wire v_1295;
wire v_1296;
wire v_1297;
wire v_1298;
wire v_1299;
wire v_1300;
wire v_1301;
wire v_1302;
wire v_1303;
wire v_1304;
wire v_1305;
wire v_1306;
wire v_1307;
wire v_1308;
wire v_1309;
wire v_1310;
wire v_1311;
wire v_1312;
wire v_1313;
wire v_1314;
wire v_1315;
wire v_1316;
wire v_1317;
wire v_1318;
wire v_1319;
wire v_1320;
wire v_1321;
wire v_1322;
wire v_1323;
wire v_1324;
wire v_1325;
wire v_1326;
wire v_1327;
wire v_1328;
wire v_1329;
wire v_1330;
wire v_1331;
wire v_1332;
wire v_1333;
wire v_1334;
wire v_1335;
wire v_1336;
wire v_1337;
wire v_1338;
wire v_1339;
wire v_1340;
wire v_1341;
wire v_1342;
wire v_1343;
wire v_1344;
wire v_1345;
wire v_1346;
wire v_1347;
wire v_1348;
wire v_1349;
wire v_1350;
wire v_1351;
wire v_1352;
wire v_1353;
wire v_1354;
wire v_1355;
wire v_1356;
wire v_1357;
wire v_1358;
wire v_1359;
wire v_1360;
wire v_1361;
wire v_1362;
wire v_1363;
wire v_1364;
wire v_1365;
wire v_1366;
wire v_1367;
wire v_1368;
wire v_1369;
wire v_1370;
wire v_1371;
wire v_1372;
wire v_1373;
wire v_1374;
wire v_1375;
wire v_1376;
wire v_1377;
wire v_1378;
wire v_1379;
wire v_1380;
wire v_1381;
wire v_1382;
wire v_1383;
wire v_1384;
wire v_1385;
wire v_1386;
wire v_1387;
wire v_1388;
wire v_1389;
wire v_1390;
wire v_1391;
wire v_1392;
wire v_1393;
wire v_1394;
wire v_1395;
wire v_1396;
wire v_1397;
wire v_1398;
wire v_1399;
wire v_1400;
wire v_1401;
wire v_1402;
wire v_1403;
wire v_1404;
wire v_1405;
wire v_1406;
wire v_1407;
wire v_1408;
wire v_1409;
wire v_1410;
wire v_1411;
wire v_1412;
wire v_1413;
wire v_1414;
wire v_1415;
wire v_1416;
wire v_1417;
wire v_1418;
wire v_1419;
wire v_1420;
wire v_1421;
wire v_1422;
wire v_1423;
wire v_1424;
wire v_1425;
wire v_1426;
wire v_1427;
wire v_1428;
wire v_1429;
wire v_1430;
wire v_1431;
wire v_1432;
wire v_1433;
wire v_1434;
wire v_1435;
wire v_1436;
wire v_1437;
wire v_1438;
wire v_1439;
wire v_1440;
wire v_1441;
wire v_1442;
wire v_1443;
wire v_1444;
wire v_1445;
wire v_1446;
wire v_1447;
wire v_1448;
wire v_1449;
wire v_1450;
wire v_1451;
wire v_1452;
wire v_1453;
wire v_1454;
wire v_1455;
wire v_1456;
wire v_1457;
wire v_1458;
wire v_1459;
wire v_1460;
wire v_1461;
wire v_1462;
wire v_1463;
wire v_1464;
wire v_1465;
wire v_1466;
wire v_1467;
wire v_1468;
wire v_1469;
wire v_1470;
wire v_1471;
wire v_1472;
wire v_1473;
wire v_1474;
wire v_1475;
wire v_1476;
wire v_1477;
wire v_1478;
wire v_1479;
wire v_1480;
wire v_1481;
wire v_1482;
wire v_1483;
wire v_1484;
wire v_1485;
wire v_1486;
wire v_1487;
wire v_1488;
wire v_1489;
wire v_1490;
wire v_1491;
wire v_1492;
wire v_1493;
wire v_1494;
wire v_1495;
wire v_1496;
wire v_1497;
wire v_1498;
wire v_1499;
wire v_1500;
wire v_1501;
wire v_1502;
wire v_1503;
wire v_1504;
wire v_1505;
wire v_1506;
wire v_1507;
wire v_1508;
wire v_1509;
wire v_1510;
wire v_1511;
wire v_1512;
wire v_1513;
wire v_1514;
wire v_1515;
wire v_1516;
wire v_1517;
wire v_1518;
wire v_1519;
wire v_1520;
wire v_1521;
wire v_1522;
wire v_1523;
wire v_1524;
wire v_1525;
wire v_1526;
wire v_1527;
wire v_1528;
wire v_1529;
wire v_1530;
wire v_1531;
wire v_1532;
wire v_1533;
wire v_1534;
wire v_1535;
wire v_1536;
wire v_1537;
wire v_1538;
wire v_1539;
wire v_1540;
wire v_1541;
wire v_1542;
wire v_1543;
wire v_1544;
wire v_1545;
wire v_1546;
wire v_1547;
wire v_1548;
wire v_1549;
wire v_1550;
wire v_1551;
wire v_1552;
wire v_1553;
wire v_1554;
wire v_1555;
wire v_1556;
wire v_1557;
wire v_1558;
wire v_1559;
wire v_1560;
wire v_1561;
wire v_1562;
wire v_1563;
wire v_1564;
wire v_1565;
wire v_1566;
wire v_1567;
wire v_1568;
wire v_1569;
wire v_1570;
wire v_1571;
wire v_1572;
wire v_1573;
wire v_1574;
wire v_1575;
wire v_1576;
wire v_1577;
wire v_1578;
wire v_1579;
wire v_1580;
wire v_1581;
wire v_1582;
wire v_1583;
wire v_1584;
wire v_1585;
wire v_1586;
wire v_1587;
wire v_1588;
wire v_1589;
wire v_1590;
wire v_1591;
wire v_1592;
wire v_1593;
wire v_1594;
wire v_1595;
wire v_1596;
wire v_1597;
wire v_1598;
wire v_1599;
wire v_1600;
wire v_1601;
wire v_1602;
wire v_1603;
wire v_1604;
wire v_1605;
wire v_1606;
wire v_1607;
wire v_1608;
wire v_1609;
wire v_1610;
wire v_1611;
wire v_1612;
wire v_1613;
wire v_1614;
wire v_1615;
wire v_1616;
wire v_1617;
wire v_1618;
wire v_1619;
wire v_1620;
wire v_1621;
wire v_1622;
wire v_1623;
wire v_1624;
wire v_1625;
wire v_1626;
wire v_1627;
wire v_1628;
wire v_1629;
wire v_1630;
wire v_1631;
wire v_1632;
wire v_1633;
wire v_1634;
wire v_1635;
wire v_1636;
wire v_1637;
wire v_1638;
wire v_1639;
wire v_1640;
wire v_1641;
wire v_1642;
wire v_1643;
wire v_1644;
wire v_1645;
wire v_1646;
wire v_1647;
wire v_1648;
wire v_1649;
wire v_1650;
wire v_1651;
wire v_1652;
wire v_1653;
wire v_1654;
wire v_1655;
wire v_1656;
wire v_1657;
wire v_1658;
wire v_1659;
wire v_1660;
wire v_1661;
wire v_1662;
wire v_1663;
wire v_1664;
wire v_1665;
wire v_1666;
wire v_1667;
wire v_1668;
wire v_1669;
wire v_1670;
wire v_1671;
wire v_1672;
wire v_1673;
wire v_1674;
wire v_1675;
wire v_1676;
wire v_1677;
wire v_1678;
wire v_1679;
wire v_1680;
wire v_1681;
wire v_1682;
wire v_1683;
wire v_1684;
wire v_1685;
wire v_1686;
wire v_1687;
wire v_1688;
wire v_1689;
wire v_1690;
wire v_1691;
wire v_1692;
wire v_1693;
wire v_1694;
wire v_1695;
wire v_1696;
wire v_1697;
wire v_1698;
wire v_1699;
wire v_1700;
wire v_1701;
wire v_1702;
wire v_1703;
wire v_1704;
wire v_1705;
wire v_1706;
wire v_1707;
wire v_1708;
wire v_1709;
wire v_1710;
wire v_1711;
wire v_1712;
wire v_1713;
wire v_1714;
wire v_1715;
wire v_1716;
wire v_1717;
wire v_1718;
wire v_1719;
wire v_1720;
wire v_1721;
wire v_1722;
wire v_1723;
wire v_1724;
wire v_1725;
wire v_1726;
wire v_1727;
wire v_1728;
wire v_1729;
wire v_1730;
wire v_1731;
wire v_1732;
wire v_1733;
wire v_1734;
wire v_1735;
wire v_1736;
wire v_1737;
wire v_1738;
wire v_1739;
wire v_1740;
wire v_1741;
wire v_1742;
wire v_1743;
wire v_1744;
wire v_1745;
wire v_1746;
wire v_1747;
wire v_1748;
wire v_1749;
wire v_1750;
wire v_1751;
wire v_1752;
wire v_1753;
wire v_1754;
wire v_1755;
wire v_1756;
wire v_1757;
wire v_1758;
wire v_1759;
wire v_1760;
wire v_1761;
wire v_1762;
wire v_1763;
wire v_1764;
wire v_1765;
wire v_1766;
wire v_1767;
wire v_1768;
wire v_1769;
wire v_1770;
wire v_1771;
wire v_1772;
wire v_1773;
wire v_1774;
wire v_1775;
wire v_1776;
wire v_1777;
wire v_1778;
wire v_1779;
wire v_1780;
wire v_1781;
wire v_1782;
wire v_1783;
wire v_1784;
wire v_1785;
wire v_1786;
wire v_1787;
wire v_1788;
wire v_1789;
wire v_1790;
wire v_1791;
wire v_1792;
wire v_1793;
wire v_1794;
wire v_1795;
wire v_1796;
wire v_1797;
wire v_1798;
wire v_1799;
wire v_1800;
wire v_1801;
wire v_1802;
wire v_1803;
wire v_1804;
wire v_1805;
wire v_1806;
wire v_1807;
wire v_1808;
wire v_1809;
wire v_1810;
wire v_1811;
wire v_1812;
wire v_1813;
wire v_1814;
wire v_1815;
wire v_1816;
wire v_1817;
wire v_1818;
wire v_1819;
wire v_1820;
wire v_1821;
wire v_1822;
wire v_1823;
wire v_1824;
wire v_1825;
wire v_1826;
wire v_1827;
wire v_1828;
wire v_1829;
wire v_1830;
wire v_1831;
wire v_1832;
wire v_1833;
wire v_1834;
wire v_1835;
wire v_1836;
wire v_1837;
wire v_1838;
wire v_1839;
wire v_1840;
wire v_1841;
wire v_1842;
wire v_1843;
wire v_1844;
wire v_1845;
wire v_1846;
wire v_1847;
wire v_1848;
wire v_1849;
wire v_1850;
wire v_1851;
wire v_1852;
wire v_1853;
wire v_1854;
wire v_1855;
wire v_1856;
wire v_1857;
wire v_1858;
wire v_1859;
wire v_1860;
wire v_1861;
wire v_1862;
wire v_1863;
wire v_1864;
wire v_1865;
wire v_1866;
wire v_1867;
wire v_1868;
wire v_1869;
wire v_1870;
wire v_1871;
wire v_1872;
wire v_1873;
wire v_1874;
wire v_1875;
wire v_1876;
wire v_1877;
wire v_1878;
wire v_1879;
wire v_1880;
wire v_1881;
wire v_1882;
wire v_1883;
wire v_1884;
wire v_1885;
wire v_1886;
wire v_1887;
wire v_1888;
wire v_1889;
wire v_1890;
wire v_1891;
wire v_1892;
wire v_1893;
wire v_1894;
wire v_1895;
wire v_1896;
wire v_1897;
wire v_1898;
wire v_1899;
wire v_1900;
wire v_1901;
wire v_1902;
wire v_1903;
wire v_1904;
wire v_1905;
wire v_1906;
wire v_1907;
wire v_1908;
wire v_1909;
wire v_1910;
wire v_1911;
wire v_1912;
wire v_1913;
wire v_1914;
wire v_1915;
wire v_1916;
wire v_1917;
wire v_1918;
wire v_1919;
wire v_1920;
wire v_1921;
wire v_1922;
wire v_1923;
wire v_1924;
wire v_1925;
wire v_1926;
wire v_1927;
wire v_1928;
wire v_1929;
wire v_1930;
wire v_1931;
wire v_1932;
wire v_1933;
wire v_1934;
wire v_1935;
wire v_1936;
wire v_1937;
wire v_1938;
wire v_1939;
wire v_1940;
wire v_1941;
wire v_1942;
wire v_1943;
wire v_1944;
wire v_1945;
wire v_1946;
wire v_1947;
wire v_1948;
wire v_1949;
wire v_1950;
wire v_1951;
wire v_1952;
wire v_1953;
wire v_1954;
wire v_1955;
wire v_1956;
wire v_1957;
wire v_1958;
wire v_1959;
wire v_1960;
wire v_1961;
wire v_1962;
wire v_1963;
wire v_1964;
wire v_1965;
wire v_1966;
wire v_1967;
wire v_1968;
wire v_1969;
wire v_1970;
wire v_1971;
wire v_1972;
wire v_1973;
wire v_1974;
wire v_1975;
wire v_1976;
wire v_1977;
wire v_1978;
wire v_1979;
wire v_1980;
wire v_1981;
wire v_1982;
wire v_1983;
wire v_1984;
wire v_1985;
wire v_1986;
wire v_1987;
wire v_1988;
wire v_1989;
wire v_1990;
wire v_1991;
wire v_1992;
wire v_1993;
wire v_1994;
wire v_1995;
wire v_1996;
wire v_1997;
wire v_1998;
wire v_1999;
wire v_2000;
wire v_2001;
wire v_2002;
wire v_2003;
wire v_2004;
wire v_2005;
wire v_2006;
wire v_2007;
wire v_2008;
wire v_2009;
wire v_2010;
wire v_2011;
wire v_2012;
wire v_2013;
wire v_2014;
wire v_2015;
wire v_2016;
wire v_2017;
wire v_2018;
wire v_2019;
wire v_2020;
wire v_2021;
wire v_2022;
wire v_2023;
wire v_2024;
wire v_2025;
wire v_2026;
wire v_2027;
wire v_2028;
wire v_2029;
wire v_2030;
wire v_2031;
wire v_2032;
wire v_2033;
wire v_2034;
wire v_2035;
wire v_2036;
wire v_2037;
wire v_2038;
wire v_2039;
wire v_2040;
wire v_2041;
wire v_2042;
wire v_2043;
wire v_2044;
wire v_2045;
wire v_2046;
wire v_2047;
wire v_2048;
wire v_2049;
wire v_2050;
wire v_2051;
wire v_2052;
wire v_2053;
wire v_2054;
wire v_2055;
wire v_2056;
wire v_2057;
wire v_2058;
wire v_2059;
wire v_2060;
wire v_2061;
wire v_2062;
wire v_2063;
wire v_2064;
wire v_2065;
wire v_2066;
wire v_2067;
wire v_2068;
wire v_2069;
wire v_2070;
wire v_2071;
wire v_2072;
wire v_2073;
wire v_2074;
wire v_2075;
wire v_2076;
wire v_2077;
wire v_2078;
wire v_2079;
wire v_2080;
wire v_2081;
wire v_2082;
wire v_2083;
wire v_2084;
wire v_2085;
wire v_2086;
wire v_2087;
wire v_2088;
wire v_2089;
wire v_2090;
wire v_2091;
wire v_2092;
wire v_2093;
wire v_2094;
wire v_2095;
wire v_2096;
wire v_2097;
wire v_2098;
wire v_2099;
wire v_2100;
wire v_2101;
wire v_2102;
wire v_2103;
wire v_2104;
wire v_2105;
wire v_2106;
wire v_2107;
wire v_2108;
wire v_2109;
wire v_2110;
wire v_2111;
wire v_2112;
wire v_2113;
wire v_2114;
wire x_1;
assign v_781 = v_1881 & v_1882 & v_1883 & v_1884;
assign v_782 = v_1885 & v_1886 & v_1887 & v_1888;
assign v_783 = v_1889 & v_1890 & v_1891 & v_1892;
assign v_784 = v_781 & v_782 & v_783;
assign v_805 = v_1893 & v_1894 & v_1895 & v_1896;
assign v_826 = v_1897 & v_1898 & v_1899 & v_1900;
assign v_847 = v_1901 & v_1902 & v_1903 & v_1904;
assign v_848 = v_805 & v_826 & v_847;
assign v_869 = v_1905 & v_1906 & v_1907 & v_1908;
assign v_890 = v_1909 & v_1910 & v_1911 & v_1912;
assign v_911 = v_1913 & v_1914 & v_1915 & v_1916;
assign v_912 = v_869 & v_890 & v_911;
assign v_933 = v_1917 & v_1918 & v_1919 & v_1920;
assign v_954 = v_1921 & v_1922 & v_1923 & v_1924;
assign v_975 = v_1925 & v_1926 & v_1927 & v_1928;
assign v_976 = v_933 & v_954 & v_975;
assign v_997 = v_1929 & v_1930 & v_1931 & v_1932;
assign v_1018 = v_1933 & v_1934 & v_1935 & v_1936;
assign v_1039 = v_1937 & v_1938 & v_1939 & v_1940;
assign v_1040 = v_997 & v_1018 & v_1039;
assign v_1061 = v_1941 & v_1942 & v_1943 & v_1944;
assign v_1082 = v_1945 & v_1946 & v_1947 & v_1948;
assign v_1103 = v_1949 & v_1950 & v_1951 & v_1952;
assign v_1104 = v_1061 & v_1082 & v_1103;
assign v_1125 = v_1953 & v_1954 & v_1955 & v_1956;
assign v_1146 = v_1957 & v_1958 & v_1959 & v_1960;
assign v_1167 = v_1961 & v_1962 & v_1963 & v_1964;
assign v_1168 = v_1125 & v_1146 & v_1167;
assign v_1169 = v_1965 & v_1966;
assign v_1170 = v_1967 & v_1968 & v_1969 & v_1970;
assign v_1171 = v_1971 & v_1972 & v_1973 & v_1974;
assign v_1172 = v_1975 & v_1976 & v_1977 & v_1978;
assign v_1173 = v_1170 & v_1171 & v_1172;
assign v_1194 = v_1979 & v_1980 & v_1981 & v_1982;
assign v_1215 = v_1983 & v_1984 & v_1985 & v_1986;
assign v_1236 = v_1987 & v_1988 & v_1989 & v_1990;
assign v_1237 = v_1194 & v_1215 & v_1236;
assign v_1258 = v_1991 & v_1992 & v_1993 & v_1994;
assign v_1279 = v_1995 & v_1996 & v_1997 & v_1998;
assign v_1300 = v_1999 & v_2000 & v_2001 & v_2002;
assign v_1301 = v_1258 & v_1279 & v_1300;
assign v_1322 = v_2003 & v_2004 & v_2005 & v_2006;
assign v_1343 = v_2007 & v_2008 & v_2009 & v_2010;
assign v_1364 = v_2011 & v_2012 & v_2013 & v_2014;
assign v_1365 = v_1322 & v_1343 & v_1364;
assign v_1386 = v_2015 & v_2016 & v_2017 & v_2018;
assign v_1407 = v_2019 & v_2020 & v_2021 & v_2022;
assign v_1428 = v_2023 & v_2024 & v_2025 & v_2026;
assign v_1429 = v_1386 & v_1407 & v_1428;
assign v_1450 = v_2027 & v_2028 & v_2029 & v_2030;
assign v_1471 = v_2031 & v_2032 & v_2033 & v_2034;
assign v_1492 = v_2035 & v_2036 & v_2037 & v_2038;
assign v_1493 = v_1450 & v_1471 & v_1492;
assign v_1494 = v_2039 & v_2040;
assign v_1515 = v_2041 & v_2042 & v_2043 & v_2044;
assign v_1536 = v_2045 & v_2046 & v_2047 & v_2048;
assign v_1557 = v_2049 & v_2050 & v_2051 & v_2052;
assign v_1558 = v_1515 & v_1536 & v_1557;
assign v_1579 = v_2053 & v_2054 & v_2055 & v_2056;
assign v_1600 = v_2057 & v_2058 & v_2059 & v_2060;
assign v_1621 = v_2061 & v_2062 & v_2063 & v_2064;
assign v_1622 = v_1579 & v_1600 & v_1621;
assign v_1643 = v_2065 & v_2066 & v_2067 & v_2068;
assign v_1664 = v_2069 & v_2070 & v_2071 & v_2072;
assign v_1685 = v_2073 & v_2074 & v_2075 & v_2076;
assign v_1686 = v_1643 & v_1664 & v_1685;
assign v_1707 = v_2077 & v_2078 & v_2079 & v_2080;
assign v_1728 = v_2081 & v_2082 & v_2083 & v_2084;
assign v_1749 = v_2085 & v_2086 & v_2087 & v_2088;
assign v_1750 = v_1707 & v_1728 & v_1749;
assign v_1771 = v_2089 & v_2090 & v_2091 & v_2092;
assign v_1792 = v_2093 & v_2094 & v_2095 & v_2096;
assign v_1813 = v_2097 & v_2098 & v_2099 & v_2100;
assign v_1814 = v_1771 & v_1792 & v_1813;
assign v_1835 = v_2101 & v_2102 & v_2103 & v_2104;
assign v_1856 = v_2105 & v_2106 & v_2107 & v_2108;
assign v_1877 = v_2109 & v_2110 & v_2111 & v_2112;
assign v_1878 = v_1835 & v_1856 & v_1877;
assign v_1880 = v_1494 & v_1879;
assign v_1881 = ~v_2 & ~v_3 & ~v_4 & ~v_5 & ~v_6;
assign v_1882 = ~v_7 & ~v_8 & ~v_9 & ~v_10 & ~v_11;
assign v_1883 = ~v_12 & ~v_13 & ~v_14 & ~v_15 & ~v_16;
assign v_1884 = ~v_17 & ~v_18 & ~v_19 & ~v_20 & v_1;
assign v_1885 = ~v_22 & ~v_24 & ~v_25 & ~v_26 & ~v_27;
assign v_1886 = ~v_28 & ~v_29 & ~v_30 & ~v_31 & ~v_32;
assign v_1887 = ~v_33 & ~v_34 & ~v_35 & ~v_36 & ~v_37;
assign v_1888 = ~v_38 & ~v_39 & ~v_40 & v_21 & v_23;
assign v_1889 = ~v_44 & ~v_45 & ~v_46 & ~v_47 & ~v_48;
assign v_1890 = ~v_49 & ~v_50 & ~v_51 & ~v_52 & ~v_53;
assign v_1891 = ~v_54 & ~v_55 & ~v_56 & ~v_57 & ~v_58;
assign v_1892 = ~v_59 & ~v_60 & v_41 & v_42 & v_43;
assign v_1893 = ~v_785 & ~v_786 & ~v_787 & ~v_788 & ~v_789;
assign v_1894 = ~v_790 & ~v_791 & ~v_792 & ~v_793 & ~v_794;
assign v_1895 = ~v_795 & ~v_796 & ~v_797 & ~v_798 & ~v_799;
assign v_1896 = ~v_800 & ~v_801 & ~v_802 & ~v_803 & ~v_804;
assign v_1897 = ~v_806 & ~v_807 & ~v_808 & ~v_809 & ~v_810;
assign v_1898 = ~v_811 & ~v_812 & ~v_813 & ~v_814 & ~v_815;
assign v_1899 = ~v_816 & ~v_817 & ~v_818 & ~v_819 & ~v_820;
assign v_1900 = ~v_821 & ~v_822 & ~v_823 & ~v_824 & ~v_825;
assign v_1901 = ~v_827 & ~v_828 & ~v_829 & ~v_830 & ~v_831;
assign v_1902 = ~v_832 & ~v_833 & ~v_834 & ~v_835 & ~v_836;
assign v_1903 = ~v_837 & ~v_838 & ~v_839 & ~v_840 & ~v_841;
assign v_1904 = ~v_842 & ~v_843 & ~v_844 & ~v_845 & ~v_846;
assign v_1905 = ~v_849 & ~v_850 & ~v_851 & ~v_852 & ~v_853;
assign v_1906 = ~v_854 & ~v_855 & ~v_856 & ~v_857 & ~v_858;
assign v_1907 = ~v_859 & ~v_860 & ~v_861 & ~v_862 & ~v_863;
assign v_1908 = ~v_864 & ~v_865 & ~v_866 & ~v_867 & ~v_868;
assign v_1909 = ~v_870 & ~v_871 & ~v_872 & ~v_873 & ~v_874;
assign v_1910 = ~v_875 & ~v_876 & ~v_877 & ~v_878 & ~v_879;
assign v_1911 = ~v_880 & ~v_881 & ~v_882 & ~v_883 & ~v_884;
assign v_1912 = ~v_885 & ~v_886 & ~v_887 & ~v_888 & ~v_889;
assign v_1913 = ~v_891 & ~v_892 & ~v_893 & ~v_894 & ~v_895;
assign v_1914 = ~v_896 & ~v_897 & ~v_898 & ~v_899 & ~v_900;
assign v_1915 = ~v_901 & ~v_902 & ~v_903 & ~v_904 & ~v_905;
assign v_1916 = ~v_906 & ~v_907 & ~v_908 & ~v_909 & ~v_910;
assign v_1917 = ~v_913 & ~v_914 & ~v_915 & ~v_916 & ~v_917;
assign v_1918 = ~v_918 & ~v_919 & ~v_920 & ~v_921 & ~v_922;
assign v_1919 = ~v_923 & ~v_924 & ~v_925 & ~v_926 & ~v_927;
assign v_1920 = ~v_928 & ~v_929 & ~v_930 & ~v_931 & ~v_932;
assign v_1921 = ~v_934 & ~v_935 & ~v_936 & ~v_937 & ~v_938;
assign v_1922 = ~v_939 & ~v_940 & ~v_941 & ~v_942 & ~v_943;
assign v_1923 = ~v_944 & ~v_945 & ~v_946 & ~v_947 & ~v_948;
assign v_1924 = ~v_949 & ~v_950 & ~v_951 & ~v_952 & ~v_953;
assign v_1925 = ~v_955 & ~v_956 & ~v_957 & ~v_958 & ~v_959;
assign v_1926 = ~v_960 & ~v_961 & ~v_962 & ~v_963 & ~v_964;
assign v_1927 = ~v_965 & ~v_966 & ~v_967 & ~v_968 & ~v_969;
assign v_1928 = ~v_970 & ~v_971 & ~v_972 & ~v_973 & ~v_974;
assign v_1929 = ~v_977 & ~v_978 & ~v_979 & ~v_980 & ~v_981;
assign v_1930 = ~v_982 & ~v_983 & ~v_984 & ~v_985 & ~v_986;
assign v_1931 = ~v_987 & ~v_988 & ~v_989 & ~v_990 & ~v_991;
assign v_1932 = ~v_992 & ~v_993 & ~v_994 & ~v_995 & ~v_996;
assign v_1933 = ~v_998 & ~v_999 & ~v_1000 & ~v_1001 & ~v_1002;
assign v_1934 = ~v_1003 & ~v_1004 & ~v_1005 & ~v_1006 & ~v_1007;
assign v_1935 = ~v_1008 & ~v_1009 & ~v_1010 & ~v_1011 & ~v_1012;
assign v_1936 = ~v_1013 & ~v_1014 & ~v_1015 & ~v_1016 & ~v_1017;
assign v_1937 = ~v_1019 & ~v_1020 & ~v_1021 & ~v_1022 & ~v_1023;
assign v_1938 = ~v_1024 & ~v_1025 & ~v_1026 & ~v_1027 & ~v_1028;
assign v_1939 = ~v_1029 & ~v_1030 & ~v_1031 & ~v_1032 & ~v_1033;
assign v_1940 = ~v_1034 & ~v_1035 & ~v_1036 & ~v_1037 & ~v_1038;
assign v_1941 = ~v_1041 & ~v_1042 & ~v_1043 & ~v_1044 & ~v_1045;
assign v_1942 = ~v_1046 & ~v_1047 & ~v_1048 & ~v_1049 & ~v_1050;
assign v_1943 = ~v_1051 & ~v_1052 & ~v_1053 & ~v_1054 & ~v_1055;
assign v_1944 = ~v_1056 & ~v_1057 & ~v_1058 & ~v_1059 & ~v_1060;
assign v_1945 = ~v_1062 & ~v_1063 & ~v_1064 & ~v_1065 & ~v_1066;
assign v_1946 = ~v_1067 & ~v_1068 & ~v_1069 & ~v_1070 & ~v_1071;
assign v_1947 = ~v_1072 & ~v_1073 & ~v_1074 & ~v_1075 & ~v_1076;
assign v_1948 = ~v_1077 & ~v_1078 & ~v_1079 & ~v_1080 & ~v_1081;
assign v_1949 = ~v_1083 & ~v_1084 & ~v_1085 & ~v_1086 & ~v_1087;
assign v_1950 = ~v_1088 & ~v_1089 & ~v_1090 & ~v_1091 & ~v_1092;
assign v_1951 = ~v_1093 & ~v_1094 & ~v_1095 & ~v_1096 & ~v_1097;
assign v_1952 = ~v_1098 & ~v_1099 & ~v_1100 & ~v_1101 & ~v_1102;
assign v_1953 = ~v_1105 & ~v_1106 & ~v_1107 & ~v_1108 & ~v_1109;
assign v_1954 = ~v_1110 & ~v_1111 & ~v_1112 & ~v_1113 & ~v_1114;
assign v_1955 = ~v_1115 & ~v_1116 & ~v_1117 & ~v_1118 & ~v_1119;
assign v_1956 = ~v_1120 & ~v_1121 & ~v_1122 & ~v_1123 & ~v_1124;
assign v_1957 = ~v_1126 & ~v_1127 & ~v_1128 & ~v_1129 & ~v_1130;
assign v_1958 = ~v_1131 & ~v_1132 & ~v_1133 & ~v_1134 & ~v_1135;
assign v_1959 = ~v_1136 & ~v_1137 & ~v_1138 & ~v_1139 & ~v_1140;
assign v_1960 = ~v_1141 & ~v_1142 & ~v_1143 & ~v_1144 & ~v_1145;
assign v_1961 = ~v_1147 & ~v_1148 & ~v_1149 & ~v_1150 & ~v_1151;
assign v_1962 = ~v_1152 & ~v_1153 & ~v_1154 & ~v_1155 & ~v_1156;
assign v_1963 = ~v_1157 & ~v_1158 & ~v_1159 & ~v_1160 & ~v_1161;
assign v_1964 = ~v_1162 & ~v_1163 & ~v_1164 & ~v_1165 & ~v_1166;
assign v_1965 = v_784 & v_848 & v_912 & v_976 & v_1040;
assign v_1966 = v_1104 & v_1168;
assign v_1967 = ~v_422 & ~v_423 & ~v_424 & ~v_425 & ~v_426;
assign v_1968 = ~v_427 & ~v_428 & ~v_429 & ~v_430 & ~v_431;
assign v_1969 = ~v_432 & ~v_433 & ~v_434 & ~v_435 & ~v_436;
assign v_1970 = ~v_437 & ~v_438 & ~v_439 & ~v_440 & v_421;
assign v_1971 = ~v_442 & ~v_444 & ~v_445 & ~v_446 & ~v_447;
assign v_1972 = ~v_448 & ~v_449 & ~v_450 & ~v_451 & ~v_452;
assign v_1973 = ~v_453 & ~v_454 & ~v_455 & ~v_456 & ~v_457;
assign v_1974 = ~v_458 & ~v_459 & ~v_460 & v_441 & v_443;
assign v_1975 = ~v_464 & ~v_465 & ~v_466 & ~v_467 & ~v_468;
assign v_1976 = ~v_469 & ~v_470 & ~v_471 & ~v_472 & ~v_473;
assign v_1977 = ~v_474 & ~v_475 & ~v_476 & ~v_477 & ~v_478;
assign v_1978 = ~v_479 & ~v_480 & v_461 & v_462 & v_463;
assign v_1979 = ~v_1174 & ~v_1175 & ~v_1176 & ~v_1177 & ~v_1178;
assign v_1980 = ~v_1179 & ~v_1180 & ~v_1181 & ~v_1182 & ~v_1183;
assign v_1981 = ~v_1184 & ~v_1185 & ~v_1186 & ~v_1187 & ~v_1188;
assign v_1982 = ~v_1189 & ~v_1190 & ~v_1191 & ~v_1192 & ~v_1193;
assign v_1983 = ~v_1195 & ~v_1196 & ~v_1197 & ~v_1198 & ~v_1199;
assign v_1984 = ~v_1200 & ~v_1201 & ~v_1202 & ~v_1203 & ~v_1204;
assign v_1985 = ~v_1205 & ~v_1206 & ~v_1207 & ~v_1208 & ~v_1209;
assign v_1986 = ~v_1210 & ~v_1211 & ~v_1212 & ~v_1213 & ~v_1214;
assign v_1987 = ~v_1216 & ~v_1217 & ~v_1218 & ~v_1219 & ~v_1220;
assign v_1988 = ~v_1221 & ~v_1222 & ~v_1223 & ~v_1224 & ~v_1225;
assign v_1989 = ~v_1226 & ~v_1227 & ~v_1228 & ~v_1229 & ~v_1230;
assign v_1990 = ~v_1231 & ~v_1232 & ~v_1233 & ~v_1234 & ~v_1235;
assign v_1991 = ~v_1238 & ~v_1239 & ~v_1240 & ~v_1241 & ~v_1242;
assign v_1992 = ~v_1243 & ~v_1244 & ~v_1245 & ~v_1246 & ~v_1247;
assign v_1993 = ~v_1248 & ~v_1249 & ~v_1250 & ~v_1251 & ~v_1252;
assign v_1994 = ~v_1253 & ~v_1254 & ~v_1255 & ~v_1256 & ~v_1257;
assign v_1995 = ~v_1259 & ~v_1260 & ~v_1261 & ~v_1262 & ~v_1263;
assign v_1996 = ~v_1264 & ~v_1265 & ~v_1266 & ~v_1267 & ~v_1268;
assign v_1997 = ~v_1269 & ~v_1270 & ~v_1271 & ~v_1272 & ~v_1273;
assign v_1998 = ~v_1274 & ~v_1275 & ~v_1276 & ~v_1277 & ~v_1278;
assign v_1999 = ~v_1280 & ~v_1281 & ~v_1282 & ~v_1283 & ~v_1284;
assign v_2000 = ~v_1285 & ~v_1286 & ~v_1287 & ~v_1288 & ~v_1289;
assign v_2001 = ~v_1290 & ~v_1291 & ~v_1292 & ~v_1293 & ~v_1294;
assign v_2002 = ~v_1295 & ~v_1296 & ~v_1297 & ~v_1298 & ~v_1299;
assign v_2003 = ~v_1302 & ~v_1303 & ~v_1304 & ~v_1305 & ~v_1306;
assign v_2004 = ~v_1307 & ~v_1308 & ~v_1309 & ~v_1310 & ~v_1311;
assign v_2005 = ~v_1312 & ~v_1313 & ~v_1314 & ~v_1315 & ~v_1316;
assign v_2006 = ~v_1317 & ~v_1318 & ~v_1319 & ~v_1320 & ~v_1321;
assign v_2007 = ~v_1323 & ~v_1324 & ~v_1325 & ~v_1326 & ~v_1327;
assign v_2008 = ~v_1328 & ~v_1329 & ~v_1330 & ~v_1331 & ~v_1332;
assign v_2009 = ~v_1333 & ~v_1334 & ~v_1335 & ~v_1336 & ~v_1337;
assign v_2010 = ~v_1338 & ~v_1339 & ~v_1340 & ~v_1341 & ~v_1342;
assign v_2011 = ~v_1344 & ~v_1345 & ~v_1346 & ~v_1347 & ~v_1348;
assign v_2012 = ~v_1349 & ~v_1350 & ~v_1351 & ~v_1352 & ~v_1353;
assign v_2013 = ~v_1354 & ~v_1355 & ~v_1356 & ~v_1357 & ~v_1358;
assign v_2014 = ~v_1359 & ~v_1360 & ~v_1361 & ~v_1362 & ~v_1363;
assign v_2015 = ~v_1366 & ~v_1367 & ~v_1368 & ~v_1369 & ~v_1370;
assign v_2016 = ~v_1371 & ~v_1372 & ~v_1373 & ~v_1374 & ~v_1375;
assign v_2017 = ~v_1376 & ~v_1377 & ~v_1378 & ~v_1379 & ~v_1380;
assign v_2018 = ~v_1381 & ~v_1382 & ~v_1383 & ~v_1384 & ~v_1385;
assign v_2019 = ~v_1387 & ~v_1388 & ~v_1389 & ~v_1390 & ~v_1391;
assign v_2020 = ~v_1392 & ~v_1393 & ~v_1394 & ~v_1395 & ~v_1396;
assign v_2021 = ~v_1397 & ~v_1398 & ~v_1399 & ~v_1400 & ~v_1401;
assign v_2022 = ~v_1402 & ~v_1403 & ~v_1404 & ~v_1405 & ~v_1406;
assign v_2023 = ~v_1408 & ~v_1409 & ~v_1410 & ~v_1411 & ~v_1412;
assign v_2024 = ~v_1413 & ~v_1414 & ~v_1415 & ~v_1416 & ~v_1417;
assign v_2025 = ~v_1418 & ~v_1419 & ~v_1420 & ~v_1421 & ~v_1422;
assign v_2026 = ~v_1423 & ~v_1424 & ~v_1425 & ~v_1426 & ~v_1427;
assign v_2027 = ~v_1430 & ~v_1431 & ~v_1432 & ~v_1433 & ~v_1434;
assign v_2028 = ~v_1435 & ~v_1436 & ~v_1437 & ~v_1438 & ~v_1439;
assign v_2029 = ~v_1440 & ~v_1441 & ~v_1442 & ~v_1443 & ~v_1444;
assign v_2030 = ~v_1445 & ~v_1446 & ~v_1447 & ~v_1448 & ~v_1449;
assign v_2031 = ~v_1451 & ~v_1452 & ~v_1453 & ~v_1454 & ~v_1455;
assign v_2032 = ~v_1456 & ~v_1457 & ~v_1458 & ~v_1459 & ~v_1460;
assign v_2033 = ~v_1461 & ~v_1462 & ~v_1463 & ~v_1464 & ~v_1465;
assign v_2034 = ~v_1466 & ~v_1467 & ~v_1468 & ~v_1469 & ~v_1470;
assign v_2035 = ~v_1472 & ~v_1473 & ~v_1474 & ~v_1475 & ~v_1476;
assign v_2036 = ~v_1477 & ~v_1478 & ~v_1479 & ~v_1480 & ~v_1481;
assign v_2037 = ~v_1482 & ~v_1483 & ~v_1484 & ~v_1485 & ~v_1486;
assign v_2038 = ~v_1487 & ~v_1488 & ~v_1489 & ~v_1490 & ~v_1491;
assign v_2039 = v_1173 & v_1237 & v_1301 & v_1365 & v_1429;
assign v_2040 = v_1493;
assign v_2041 = ~v_1495 & ~v_1496 & ~v_1497 & ~v_1498 & ~v_1499;
assign v_2042 = ~v_1500 & ~v_1501 & ~v_1502 & ~v_1503 & ~v_1504;
assign v_2043 = ~v_1505 & ~v_1506 & ~v_1507 & ~v_1508 & ~v_1509;
assign v_2044 = ~v_1510 & ~v_1511 & ~v_1512 & ~v_1513 & ~v_1514;
assign v_2045 = ~v_1516 & ~v_1517 & ~v_1518 & ~v_1519 & ~v_1520;
assign v_2046 = ~v_1521 & ~v_1522 & ~v_1523 & ~v_1524 & ~v_1525;
assign v_2047 = ~v_1526 & ~v_1527 & ~v_1528 & ~v_1529 & ~v_1530;
assign v_2048 = ~v_1531 & ~v_1532 & ~v_1533 & ~v_1534 & ~v_1535;
assign v_2049 = ~v_1537 & ~v_1538 & ~v_1539 & ~v_1540 & ~v_1541;
assign v_2050 = ~v_1542 & ~v_1543 & ~v_1544 & ~v_1545 & ~v_1546;
assign v_2051 = ~v_1547 & ~v_1548 & ~v_1549 & ~v_1550 & ~v_1551;
assign v_2052 = ~v_1552 & ~v_1553 & ~v_1554 & ~v_1555 & ~v_1556;
assign v_2053 = ~v_1559 & ~v_1560 & ~v_1561 & ~v_1562 & ~v_1563;
assign v_2054 = ~v_1564 & ~v_1565 & ~v_1566 & ~v_1567 & ~v_1568;
assign v_2055 = ~v_1569 & ~v_1570 & ~v_1571 & ~v_1572 & ~v_1573;
assign v_2056 = ~v_1574 & ~v_1575 & ~v_1576 & ~v_1577 & ~v_1578;
assign v_2057 = ~v_1580 & ~v_1581 & ~v_1582 & ~v_1583 & ~v_1584;
assign v_2058 = ~v_1585 & ~v_1586 & ~v_1587 & ~v_1588 & ~v_1589;
assign v_2059 = ~v_1590 & ~v_1591 & ~v_1592 & ~v_1593 & ~v_1594;
assign v_2060 = ~v_1595 & ~v_1596 & ~v_1597 & ~v_1598 & ~v_1599;
assign v_2061 = ~v_1601 & ~v_1602 & ~v_1603 & ~v_1604 & ~v_1605;
assign v_2062 = ~v_1606 & ~v_1607 & ~v_1608 & ~v_1609 & ~v_1610;
assign v_2063 = ~v_1611 & ~v_1612 & ~v_1613 & ~v_1614 & ~v_1615;
assign v_2064 = ~v_1616 & ~v_1617 & ~v_1618 & ~v_1619 & ~v_1620;
assign v_2065 = ~v_1623 & ~v_1624 & ~v_1625 & ~v_1626 & ~v_1627;
assign v_2066 = ~v_1628 & ~v_1629 & ~v_1630 & ~v_1631 & ~v_1632;
assign v_2067 = ~v_1633 & ~v_1634 & ~v_1635 & ~v_1636 & ~v_1637;
assign v_2068 = ~v_1638 & ~v_1639 & ~v_1640 & ~v_1641 & ~v_1642;
assign v_2069 = ~v_1644 & ~v_1645 & ~v_1646 & ~v_1647 & ~v_1648;
assign v_2070 = ~v_1649 & ~v_1650 & ~v_1651 & ~v_1652 & ~v_1653;
assign v_2071 = ~v_1654 & ~v_1655 & ~v_1656 & ~v_1657 & ~v_1658;
assign v_2072 = ~v_1659 & ~v_1660 & ~v_1661 & ~v_1662 & ~v_1663;
assign v_2073 = ~v_1665 & ~v_1666 & ~v_1667 & ~v_1668 & ~v_1669;
assign v_2074 = ~v_1670 & ~v_1671 & ~v_1672 & ~v_1673 & ~v_1674;
assign v_2075 = ~v_1675 & ~v_1676 & ~v_1677 & ~v_1678 & ~v_1679;
assign v_2076 = ~v_1680 & ~v_1681 & ~v_1682 & ~v_1683 & ~v_1684;
assign v_2077 = ~v_1687 & ~v_1688 & ~v_1689 & ~v_1690 & ~v_1691;
assign v_2078 = ~v_1692 & ~v_1693 & ~v_1694 & ~v_1695 & ~v_1696;
assign v_2079 = ~v_1697 & ~v_1698 & ~v_1699 & ~v_1700 & ~v_1701;
assign v_2080 = ~v_1702 & ~v_1703 & ~v_1704 & ~v_1705 & ~v_1706;
assign v_2081 = ~v_1708 & ~v_1709 & ~v_1710 & ~v_1711 & ~v_1712;
assign v_2082 = ~v_1713 & ~v_1714 & ~v_1715 & ~v_1716 & ~v_1717;
assign v_2083 = ~v_1718 & ~v_1719 & ~v_1720 & ~v_1721 & ~v_1722;
assign v_2084 = ~v_1723 & ~v_1724 & ~v_1725 & ~v_1726 & ~v_1727;
assign v_2085 = ~v_1729 & ~v_1730 & ~v_1731 & ~v_1732 & ~v_1733;
assign v_2086 = ~v_1734 & ~v_1735 & ~v_1736 & ~v_1737 & ~v_1738;
assign v_2087 = ~v_1739 & ~v_1740 & ~v_1741 & ~v_1742 & ~v_1743;
assign v_2088 = ~v_1744 & ~v_1745 & ~v_1746 & ~v_1747 & ~v_1748;
assign v_2089 = ~v_1751 & ~v_1752 & ~v_1753 & ~v_1754 & ~v_1755;
assign v_2090 = ~v_1756 & ~v_1757 & ~v_1758 & ~v_1759 & ~v_1760;
assign v_2091 = ~v_1761 & ~v_1762 & ~v_1763 & ~v_1764 & ~v_1765;
assign v_2092 = ~v_1766 & ~v_1767 & ~v_1768 & ~v_1769 & ~v_1770;
assign v_2093 = ~v_1772 & ~v_1773 & ~v_1774 & ~v_1775 & ~v_1776;
assign v_2094 = ~v_1777 & ~v_1778 & ~v_1779 & ~v_1780 & ~v_1781;
assign v_2095 = ~v_1782 & ~v_1783 & ~v_1784 & ~v_1785 & ~v_1786;
assign v_2096 = ~v_1787 & ~v_1788 & ~v_1789 & ~v_1790 & ~v_1791;
assign v_2097 = ~v_1793 & ~v_1794 & ~v_1795 & ~v_1796 & ~v_1797;
assign v_2098 = ~v_1798 & ~v_1799 & ~v_1800 & ~v_1801 & ~v_1802;
assign v_2099 = ~v_1803 & ~v_1804 & ~v_1805 & ~v_1806 & ~v_1807;
assign v_2100 = ~v_1808 & ~v_1809 & ~v_1810 & ~v_1811 & ~v_1812;
assign v_2101 = ~v_1815 & ~v_1816 & ~v_1817 & ~v_1818 & ~v_1819;
assign v_2102 = ~v_1820 & ~v_1821 & ~v_1822 & ~v_1823 & ~v_1824;
assign v_2103 = ~v_1825 & ~v_1826 & ~v_1827 & ~v_1828 & ~v_1829;
assign v_2104 = ~v_1830 & ~v_1831 & ~v_1832 & ~v_1833 & ~v_1834;
assign v_2105 = ~v_1836 & ~v_1837 & ~v_1838 & ~v_1839 & ~v_1840;
assign v_2106 = ~v_1841 & ~v_1842 & ~v_1843 & ~v_1844 & ~v_1845;
assign v_2107 = ~v_1846 & ~v_1847 & ~v_1848 & ~v_1849 & ~v_1850;
assign v_2108 = ~v_1851 & ~v_1852 & ~v_1853 & ~v_1854 & ~v_1855;
assign v_2109 = ~v_1857 & ~v_1858 & ~v_1859 & ~v_1860 & ~v_1861;
assign v_2110 = ~v_1862 & ~v_1863 & ~v_1864 & ~v_1865 & ~v_1866;
assign v_2111 = ~v_1867 & ~v_1868 & ~v_1869 & ~v_1870 & ~v_1871;
assign v_2112 = ~v_1872 & ~v_1873 & ~v_1874 & ~v_1875 & ~v_1876;
assign v_1879 = v_2113 | v_2114;
assign v_2113 = v_1558 | v_1622 | v_1686 | v_1750 | v_1814;
assign v_2114 = v_1878;
assign v_785 = v_21 ^ v_61;
assign v_786 = v_22 ^ v_62;
assign v_787 = v_23 ^ v_63;
assign v_788 = v_24 ^ v_64;
assign v_789 = v_25 ^ v_65;
assign v_790 = v_26 ^ v_66;
assign v_791 = v_27 ^ v_67;
assign v_792 = v_28 ^ v_68;
assign v_793 = v_29 ^ v_69;
assign v_794 = v_30 ^ v_70;
assign v_795 = v_31 ^ v_71;
assign v_796 = v_32 ^ v_72;
assign v_797 = v_33 ^ v_73;
assign v_798 = v_34 ^ v_74;
assign v_799 = v_35 ^ v_75;
assign v_800 = v_36 ^ v_76;
assign v_801 = v_37 ^ v_77;
assign v_802 = v_38 ^ v_78;
assign v_803 = v_39 ^ v_79;
assign v_804 = v_40 ^ v_80;
assign v_806 = v_41 ^ v_81;
assign v_807 = v_42 ^ v_82;
assign v_808 = v_43 ^ v_83;
assign v_809 = v_44 ^ v_84;
assign v_810 = v_45 ^ v_85;
assign v_811 = v_46 ^ v_86;
assign v_812 = v_47 ^ v_87;
assign v_813 = v_48 ^ v_88;
assign v_814 = v_49 ^ v_89;
assign v_815 = v_50 ^ v_90;
assign v_816 = v_51 ^ v_91;
assign v_817 = v_52 ^ v_92;
assign v_818 = v_53 ^ v_93;
assign v_819 = v_54 ^ v_94;
assign v_820 = v_55 ^ v_95;
assign v_821 = v_56 ^ v_96;
assign v_822 = v_57 ^ v_97;
assign v_823 = v_58 ^ v_98;
assign v_824 = v_59 ^ v_99;
assign v_825 = v_60 ^ v_100;
assign v_827 = v_1 ^ v_101;
assign v_828 = v_2 ^ v_102;
assign v_829 = v_3 ^ v_103;
assign v_830 = v_4 ^ v_104;
assign v_831 = v_5 ^ v_105;
assign v_832 = v_6 ^ v_106;
assign v_833 = v_7 ^ v_107;
assign v_834 = v_8 ^ v_108;
assign v_835 = v_9 ^ v_109;
assign v_836 = v_10 ^ v_110;
assign v_837 = v_11 ^ v_111;
assign v_838 = v_12 ^ v_112;
assign v_839 = v_13 ^ v_113;
assign v_840 = v_14 ^ v_114;
assign v_841 = v_15 ^ v_115;
assign v_842 = v_16 ^ v_116;
assign v_843 = v_17 ^ v_117;
assign v_844 = v_18 ^ v_118;
assign v_845 = v_19 ^ v_119;
assign v_846 = v_20 ^ v_120;
assign v_849 = v_81 ^ v_121;
assign v_850 = v_82 ^ v_122;
assign v_851 = v_83 ^ v_123;
assign v_852 = v_84 ^ v_124;
assign v_853 = v_85 ^ v_125;
assign v_854 = v_86 ^ v_126;
assign v_855 = v_87 ^ v_127;
assign v_856 = v_88 ^ v_128;
assign v_857 = v_89 ^ v_129;
assign v_858 = v_90 ^ v_130;
assign v_859 = v_91 ^ v_131;
assign v_860 = v_92 ^ v_132;
assign v_861 = v_93 ^ v_133;
assign v_862 = v_94 ^ v_134;
assign v_863 = v_95 ^ v_135;
assign v_864 = v_96 ^ v_136;
assign v_865 = v_97 ^ v_137;
assign v_866 = v_98 ^ v_138;
assign v_867 = v_99 ^ v_139;
assign v_868 = v_100 ^ v_140;
assign v_870 = v_101 ^ v_141;
assign v_871 = v_102 ^ v_142;
assign v_872 = v_103 ^ v_143;
assign v_873 = v_104 ^ v_144;
assign v_874 = v_105 ^ v_145;
assign v_875 = v_106 ^ v_146;
assign v_876 = v_107 ^ v_147;
assign v_877 = v_108 ^ v_148;
assign v_878 = v_109 ^ v_149;
assign v_879 = v_110 ^ v_150;
assign v_880 = v_111 ^ v_151;
assign v_881 = v_112 ^ v_152;
assign v_882 = v_113 ^ v_153;
assign v_883 = v_114 ^ v_154;
assign v_884 = v_115 ^ v_155;
assign v_885 = v_116 ^ v_156;
assign v_886 = v_117 ^ v_157;
assign v_887 = v_118 ^ v_158;
assign v_888 = v_119 ^ v_159;
assign v_889 = v_120 ^ v_160;
assign v_891 = v_61 ^ v_161;
assign v_892 = v_62 ^ v_162;
assign v_893 = v_63 ^ v_163;
assign v_894 = v_64 ^ v_164;
assign v_895 = v_65 ^ v_165;
assign v_896 = v_66 ^ v_166;
assign v_897 = v_67 ^ v_167;
assign v_898 = v_68 ^ v_168;
assign v_899 = v_69 ^ v_169;
assign v_900 = v_70 ^ v_170;
assign v_901 = v_71 ^ v_171;
assign v_902 = v_72 ^ v_172;
assign v_903 = v_73 ^ v_173;
assign v_904 = v_74 ^ v_174;
assign v_905 = v_75 ^ v_175;
assign v_906 = v_76 ^ v_176;
assign v_907 = v_77 ^ v_177;
assign v_908 = v_78 ^ v_178;
assign v_909 = v_79 ^ v_179;
assign v_910 = v_80 ^ v_180;
assign v_913 = v_141 ^ v_181;
assign v_914 = v_142 ^ v_182;
assign v_915 = v_143 ^ v_183;
assign v_916 = v_144 ^ v_184;
assign v_917 = v_145 ^ v_185;
assign v_918 = v_146 ^ v_186;
assign v_919 = v_147 ^ v_187;
assign v_920 = v_148 ^ v_188;
assign v_921 = v_149 ^ v_189;
assign v_922 = v_150 ^ v_190;
assign v_923 = v_151 ^ v_191;
assign v_924 = v_152 ^ v_192;
assign v_925 = v_153 ^ v_193;
assign v_926 = v_154 ^ v_194;
assign v_927 = v_155 ^ v_195;
assign v_928 = v_156 ^ v_196;
assign v_929 = v_157 ^ v_197;
assign v_930 = v_158 ^ v_198;
assign v_931 = v_159 ^ v_199;
assign v_932 = v_160 ^ v_200;
assign v_934 = v_161 ^ v_201;
assign v_935 = v_162 ^ v_202;
assign v_936 = v_163 ^ v_203;
assign v_937 = v_164 ^ v_204;
assign v_938 = v_165 ^ v_205;
assign v_939 = v_166 ^ v_206;
assign v_940 = v_167 ^ v_207;
assign v_941 = v_168 ^ v_208;
assign v_942 = v_169 ^ v_209;
assign v_943 = v_170 ^ v_210;
assign v_944 = v_171 ^ v_211;
assign v_945 = v_172 ^ v_212;
assign v_946 = v_173 ^ v_213;
assign v_947 = v_174 ^ v_214;
assign v_948 = v_175 ^ v_215;
assign v_949 = v_176 ^ v_216;
assign v_950 = v_177 ^ v_217;
assign v_951 = v_178 ^ v_218;
assign v_952 = v_179 ^ v_219;
assign v_953 = v_180 ^ v_220;
assign v_955 = v_121 ^ v_221;
assign v_956 = v_122 ^ v_222;
assign v_957 = v_123 ^ v_223;
assign v_958 = v_124 ^ v_224;
assign v_959 = v_125 ^ v_225;
assign v_960 = v_126 ^ v_226;
assign v_961 = v_127 ^ v_227;
assign v_962 = v_128 ^ v_228;
assign v_963 = v_129 ^ v_229;
assign v_964 = v_130 ^ v_230;
assign v_965 = v_131 ^ v_231;
assign v_966 = v_132 ^ v_232;
assign v_967 = v_133 ^ v_233;
assign v_968 = v_134 ^ v_234;
assign v_969 = v_135 ^ v_235;
assign v_970 = v_136 ^ v_236;
assign v_971 = v_137 ^ v_237;
assign v_972 = v_138 ^ v_238;
assign v_973 = v_139 ^ v_239;
assign v_974 = v_140 ^ v_240;
assign v_977 = v_201 ^ v_241;
assign v_978 = v_202 ^ v_242;
assign v_979 = v_203 ^ v_243;
assign v_980 = v_204 ^ v_244;
assign v_981 = v_205 ^ v_245;
assign v_982 = v_206 ^ v_246;
assign v_983 = v_207 ^ v_247;
assign v_984 = v_208 ^ v_248;
assign v_985 = v_209 ^ v_249;
assign v_986 = v_210 ^ v_250;
assign v_987 = v_211 ^ v_251;
assign v_988 = v_212 ^ v_252;
assign v_989 = v_213 ^ v_253;
assign v_990 = v_214 ^ v_254;
assign v_991 = v_215 ^ v_255;
assign v_992 = v_216 ^ v_256;
assign v_993 = v_217 ^ v_257;
assign v_994 = v_218 ^ v_258;
assign v_995 = v_219 ^ v_259;
assign v_996 = v_220 ^ v_260;
assign v_998 = v_221 ^ v_261;
assign v_999 = v_222 ^ v_262;
assign v_1000 = v_223 ^ v_263;
assign v_1001 = v_224 ^ v_264;
assign v_1002 = v_225 ^ v_265;
assign v_1003 = v_226 ^ v_266;
assign v_1004 = v_227 ^ v_267;
assign v_1005 = v_228 ^ v_268;
assign v_1006 = v_229 ^ v_269;
assign v_1007 = v_230 ^ v_270;
assign v_1008 = v_231 ^ v_271;
assign v_1009 = v_232 ^ v_272;
assign v_1010 = v_233 ^ v_273;
assign v_1011 = v_234 ^ v_274;
assign v_1012 = v_235 ^ v_275;
assign v_1013 = v_236 ^ v_276;
assign v_1014 = v_237 ^ v_277;
assign v_1015 = v_238 ^ v_278;
assign v_1016 = v_239 ^ v_279;
assign v_1017 = v_240 ^ v_280;
assign v_1019 = v_181 ^ v_281;
assign v_1020 = v_182 ^ v_282;
assign v_1021 = v_183 ^ v_283;
assign v_1022 = v_184 ^ v_284;
assign v_1023 = v_185 ^ v_285;
assign v_1024 = v_186 ^ v_286;
assign v_1025 = v_187 ^ v_287;
assign v_1026 = v_188 ^ v_288;
assign v_1027 = v_189 ^ v_289;
assign v_1028 = v_190 ^ v_290;
assign v_1029 = v_191 ^ v_291;
assign v_1030 = v_192 ^ v_292;
assign v_1031 = v_193 ^ v_293;
assign v_1032 = v_194 ^ v_294;
assign v_1033 = v_195 ^ v_295;
assign v_1034 = v_196 ^ v_296;
assign v_1035 = v_197 ^ v_297;
assign v_1036 = v_198 ^ v_298;
assign v_1037 = v_199 ^ v_299;
assign v_1038 = v_200 ^ v_300;
assign v_1041 = v_261 ^ v_301;
assign v_1042 = v_262 ^ v_302;
assign v_1043 = v_263 ^ v_303;
assign v_1044 = v_264 ^ v_304;
assign v_1045 = v_265 ^ v_305;
assign v_1046 = v_266 ^ v_306;
assign v_1047 = v_267 ^ v_307;
assign v_1048 = v_268 ^ v_308;
assign v_1049 = v_269 ^ v_309;
assign v_1050 = v_270 ^ v_310;
assign v_1051 = v_271 ^ v_311;
assign v_1052 = v_272 ^ v_312;
assign v_1053 = v_273 ^ v_313;
assign v_1054 = v_274 ^ v_314;
assign v_1055 = v_275 ^ v_315;
assign v_1056 = v_276 ^ v_316;
assign v_1057 = v_277 ^ v_317;
assign v_1058 = v_278 ^ v_318;
assign v_1059 = v_279 ^ v_319;
assign v_1060 = v_280 ^ v_320;
assign v_1062 = v_281 ^ v_321;
assign v_1063 = v_282 ^ v_322;
assign v_1064 = v_283 ^ v_323;
assign v_1065 = v_284 ^ v_324;
assign v_1066 = v_285 ^ v_325;
assign v_1067 = v_286 ^ v_326;
assign v_1068 = v_287 ^ v_327;
assign v_1069 = v_288 ^ v_328;
assign v_1070 = v_289 ^ v_329;
assign v_1071 = v_290 ^ v_330;
assign v_1072 = v_291 ^ v_331;
assign v_1073 = v_292 ^ v_332;
assign v_1074 = v_293 ^ v_333;
assign v_1075 = v_294 ^ v_334;
assign v_1076 = v_295 ^ v_335;
assign v_1077 = v_296 ^ v_336;
assign v_1078 = v_297 ^ v_337;
assign v_1079 = v_298 ^ v_338;
assign v_1080 = v_299 ^ v_339;
assign v_1081 = v_300 ^ v_340;
assign v_1083 = v_241 ^ v_341;
assign v_1084 = v_242 ^ v_342;
assign v_1085 = v_243 ^ v_343;
assign v_1086 = v_244 ^ v_344;
assign v_1087 = v_245 ^ v_345;
assign v_1088 = v_246 ^ v_346;
assign v_1089 = v_247 ^ v_347;
assign v_1090 = v_248 ^ v_348;
assign v_1091 = v_249 ^ v_349;
assign v_1092 = v_250 ^ v_350;
assign v_1093 = v_251 ^ v_351;
assign v_1094 = v_252 ^ v_352;
assign v_1095 = v_253 ^ v_353;
assign v_1096 = v_254 ^ v_354;
assign v_1097 = v_255 ^ v_355;
assign v_1098 = v_256 ^ v_356;
assign v_1099 = v_257 ^ v_357;
assign v_1100 = v_258 ^ v_358;
assign v_1101 = v_259 ^ v_359;
assign v_1102 = v_260 ^ v_360;
assign v_1105 = v_321 ^ v_361;
assign v_1106 = v_322 ^ v_362;
assign v_1107 = v_323 ^ v_363;
assign v_1108 = v_324 ^ v_364;
assign v_1109 = v_325 ^ v_365;
assign v_1110 = v_326 ^ v_366;
assign v_1111 = v_327 ^ v_367;
assign v_1112 = v_328 ^ v_368;
assign v_1113 = v_329 ^ v_369;
assign v_1114 = v_330 ^ v_370;
assign v_1115 = v_331 ^ v_371;
assign v_1116 = v_332 ^ v_372;
assign v_1117 = v_333 ^ v_373;
assign v_1118 = v_334 ^ v_374;
assign v_1119 = v_335 ^ v_375;
assign v_1120 = v_336 ^ v_376;
assign v_1121 = v_337 ^ v_377;
assign v_1122 = v_338 ^ v_378;
assign v_1123 = v_339 ^ v_379;
assign v_1124 = v_340 ^ v_380;
assign v_1126 = v_341 ^ v_381;
assign v_1127 = v_342 ^ v_382;
assign v_1128 = v_343 ^ v_383;
assign v_1129 = v_344 ^ v_384;
assign v_1130 = v_345 ^ v_385;
assign v_1131 = v_346 ^ v_386;
assign v_1132 = v_347 ^ v_387;
assign v_1133 = v_348 ^ v_388;
assign v_1134 = v_349 ^ v_389;
assign v_1135 = v_350 ^ v_390;
assign v_1136 = v_351 ^ v_391;
assign v_1137 = v_352 ^ v_392;
assign v_1138 = v_353 ^ v_393;
assign v_1139 = v_354 ^ v_394;
assign v_1140 = v_355 ^ v_395;
assign v_1141 = v_356 ^ v_396;
assign v_1142 = v_357 ^ v_397;
assign v_1143 = v_358 ^ v_398;
assign v_1144 = v_359 ^ v_399;
assign v_1145 = v_360 ^ v_400;
assign v_1147 = v_301 ^ v_401;
assign v_1148 = v_302 ^ v_402;
assign v_1149 = v_303 ^ v_403;
assign v_1150 = v_304 ^ v_404;
assign v_1151 = v_305 ^ v_405;
assign v_1152 = v_306 ^ v_406;
assign v_1153 = v_307 ^ v_407;
assign v_1154 = v_308 ^ v_408;
assign v_1155 = v_309 ^ v_409;
assign v_1156 = v_310 ^ v_410;
assign v_1157 = v_311 ^ v_411;
assign v_1158 = v_312 ^ v_412;
assign v_1159 = v_313 ^ v_413;
assign v_1160 = v_314 ^ v_414;
assign v_1161 = v_315 ^ v_415;
assign v_1162 = v_316 ^ v_416;
assign v_1163 = v_317 ^ v_417;
assign v_1164 = v_318 ^ v_418;
assign v_1165 = v_319 ^ v_419;
assign v_1166 = v_320 ^ v_420;
assign v_1174 = v_441 ^ v_481;
assign v_1175 = v_442 ^ v_482;
assign v_1176 = v_443 ^ v_483;
assign v_1177 = v_444 ^ v_484;
assign v_1178 = v_445 ^ v_485;
assign v_1179 = v_446 ^ v_486;
assign v_1180 = v_447 ^ v_487;
assign v_1181 = v_448 ^ v_488;
assign v_1182 = v_449 ^ v_489;
assign v_1183 = v_450 ^ v_490;
assign v_1184 = v_451 ^ v_491;
assign v_1185 = v_452 ^ v_492;
assign v_1186 = v_453 ^ v_493;
assign v_1187 = v_454 ^ v_494;
assign v_1188 = v_455 ^ v_495;
assign v_1189 = v_456 ^ v_496;
assign v_1190 = v_457 ^ v_497;
assign v_1191 = v_458 ^ v_498;
assign v_1192 = v_459 ^ v_499;
assign v_1193 = v_460 ^ v_500;
assign v_1195 = v_461 ^ v_501;
assign v_1196 = v_462 ^ v_502;
assign v_1197 = v_463 ^ v_503;
assign v_1198 = v_464 ^ v_504;
assign v_1199 = v_465 ^ v_505;
assign v_1200 = v_466 ^ v_506;
assign v_1201 = v_467 ^ v_507;
assign v_1202 = v_468 ^ v_508;
assign v_1203 = v_469 ^ v_509;
assign v_1204 = v_470 ^ v_510;
assign v_1205 = v_471 ^ v_511;
assign v_1206 = v_472 ^ v_512;
assign v_1207 = v_473 ^ v_513;
assign v_1208 = v_474 ^ v_514;
assign v_1209 = v_475 ^ v_515;
assign v_1210 = v_476 ^ v_516;
assign v_1211 = v_477 ^ v_517;
assign v_1212 = v_478 ^ v_518;
assign v_1213 = v_479 ^ v_519;
assign v_1214 = v_480 ^ v_520;
assign v_1216 = v_421 ^ v_521;
assign v_1217 = v_422 ^ v_522;
assign v_1218 = v_423 ^ v_523;
assign v_1219 = v_424 ^ v_524;
assign v_1220 = v_425 ^ v_525;
assign v_1221 = v_426 ^ v_526;
assign v_1222 = v_427 ^ v_527;
assign v_1223 = v_428 ^ v_528;
assign v_1224 = v_429 ^ v_529;
assign v_1225 = v_430 ^ v_530;
assign v_1226 = v_431 ^ v_531;
assign v_1227 = v_432 ^ v_532;
assign v_1228 = v_433 ^ v_533;
assign v_1229 = v_434 ^ v_534;
assign v_1230 = v_435 ^ v_535;
assign v_1231 = v_436 ^ v_536;
assign v_1232 = v_437 ^ v_537;
assign v_1233 = v_438 ^ v_538;
assign v_1234 = v_439 ^ v_539;
assign v_1235 = v_440 ^ v_540;
assign v_1238 = v_501 ^ v_541;
assign v_1239 = v_502 ^ v_542;
assign v_1240 = v_503 ^ v_543;
assign v_1241 = v_504 ^ v_544;
assign v_1242 = v_505 ^ v_545;
assign v_1243 = v_506 ^ v_546;
assign v_1244 = v_507 ^ v_547;
assign v_1245 = v_508 ^ v_548;
assign v_1246 = v_509 ^ v_549;
assign v_1247 = v_510 ^ v_550;
assign v_1248 = v_511 ^ v_551;
assign v_1249 = v_512 ^ v_552;
assign v_1250 = v_513 ^ v_553;
assign v_1251 = v_514 ^ v_554;
assign v_1252 = v_515 ^ v_555;
assign v_1253 = v_516 ^ v_556;
assign v_1254 = v_517 ^ v_557;
assign v_1255 = v_518 ^ v_558;
assign v_1256 = v_519 ^ v_559;
assign v_1257 = v_520 ^ v_560;
assign v_1259 = v_521 ^ v_561;
assign v_1260 = v_522 ^ v_562;
assign v_1261 = v_523 ^ v_563;
assign v_1262 = v_524 ^ v_564;
assign v_1263 = v_525 ^ v_565;
assign v_1264 = v_526 ^ v_566;
assign v_1265 = v_527 ^ v_567;
assign v_1266 = v_528 ^ v_568;
assign v_1267 = v_529 ^ v_569;
assign v_1268 = v_530 ^ v_570;
assign v_1269 = v_531 ^ v_571;
assign v_1270 = v_532 ^ v_572;
assign v_1271 = v_533 ^ v_573;
assign v_1272 = v_534 ^ v_574;
assign v_1273 = v_535 ^ v_575;
assign v_1274 = v_536 ^ v_576;
assign v_1275 = v_537 ^ v_577;
assign v_1276 = v_538 ^ v_578;
assign v_1277 = v_539 ^ v_579;
assign v_1278 = v_540 ^ v_580;
assign v_1280 = v_481 ^ v_581;
assign v_1281 = v_482 ^ v_582;
assign v_1282 = v_483 ^ v_583;
assign v_1283 = v_484 ^ v_584;
assign v_1284 = v_485 ^ v_585;
assign v_1285 = v_486 ^ v_586;
assign v_1286 = v_487 ^ v_587;
assign v_1287 = v_488 ^ v_588;
assign v_1288 = v_489 ^ v_589;
assign v_1289 = v_490 ^ v_590;
assign v_1290 = v_491 ^ v_591;
assign v_1291 = v_492 ^ v_592;
assign v_1292 = v_493 ^ v_593;
assign v_1293 = v_494 ^ v_594;
assign v_1294 = v_495 ^ v_595;
assign v_1295 = v_496 ^ v_596;
assign v_1296 = v_497 ^ v_597;
assign v_1297 = v_498 ^ v_598;
assign v_1298 = v_499 ^ v_599;
assign v_1299 = v_500 ^ v_600;
assign v_1302 = v_561 ^ v_601;
assign v_1303 = v_562 ^ v_602;
assign v_1304 = v_563 ^ v_603;
assign v_1305 = v_564 ^ v_604;
assign v_1306 = v_565 ^ v_605;
assign v_1307 = v_566 ^ v_606;
assign v_1308 = v_567 ^ v_607;
assign v_1309 = v_568 ^ v_608;
assign v_1310 = v_569 ^ v_609;
assign v_1311 = v_570 ^ v_610;
assign v_1312 = v_571 ^ v_611;
assign v_1313 = v_572 ^ v_612;
assign v_1314 = v_573 ^ v_613;
assign v_1315 = v_574 ^ v_614;
assign v_1316 = v_575 ^ v_615;
assign v_1317 = v_576 ^ v_616;
assign v_1318 = v_577 ^ v_617;
assign v_1319 = v_578 ^ v_618;
assign v_1320 = v_579 ^ v_619;
assign v_1321 = v_580 ^ v_620;
assign v_1323 = v_581 ^ v_621;
assign v_1324 = v_582 ^ v_622;
assign v_1325 = v_583 ^ v_623;
assign v_1326 = v_584 ^ v_624;
assign v_1327 = v_585 ^ v_625;
assign v_1328 = v_586 ^ v_626;
assign v_1329 = v_587 ^ v_627;
assign v_1330 = v_588 ^ v_628;
assign v_1331 = v_589 ^ v_629;
assign v_1332 = v_590 ^ v_630;
assign v_1333 = v_591 ^ v_631;
assign v_1334 = v_592 ^ v_632;
assign v_1335 = v_593 ^ v_633;
assign v_1336 = v_594 ^ v_634;
assign v_1337 = v_595 ^ v_635;
assign v_1338 = v_596 ^ v_636;
assign v_1339 = v_597 ^ v_637;
assign v_1340 = v_598 ^ v_638;
assign v_1341 = v_599 ^ v_639;
assign v_1342 = v_600 ^ v_640;
assign v_1344 = v_541 ^ v_641;
assign v_1345 = v_542 ^ v_642;
assign v_1346 = v_543 ^ v_643;
assign v_1347 = v_544 ^ v_644;
assign v_1348 = v_545 ^ v_645;
assign v_1349 = v_546 ^ v_646;
assign v_1350 = v_547 ^ v_647;
assign v_1351 = v_548 ^ v_648;
assign v_1352 = v_549 ^ v_649;
assign v_1353 = v_550 ^ v_650;
assign v_1354 = v_551 ^ v_651;
assign v_1355 = v_552 ^ v_652;
assign v_1356 = v_553 ^ v_653;
assign v_1357 = v_554 ^ v_654;
assign v_1358 = v_555 ^ v_655;
assign v_1359 = v_556 ^ v_656;
assign v_1360 = v_557 ^ v_657;
assign v_1361 = v_558 ^ v_658;
assign v_1362 = v_559 ^ v_659;
assign v_1363 = v_560 ^ v_660;
assign v_1366 = v_621 ^ v_661;
assign v_1367 = v_622 ^ v_662;
assign v_1368 = v_623 ^ v_663;
assign v_1369 = v_624 ^ v_664;
assign v_1370 = v_625 ^ v_665;
assign v_1371 = v_626 ^ v_666;
assign v_1372 = v_627 ^ v_667;
assign v_1373 = v_628 ^ v_668;
assign v_1374 = v_629 ^ v_669;
assign v_1375 = v_630 ^ v_670;
assign v_1376 = v_631 ^ v_671;
assign v_1377 = v_632 ^ v_672;
assign v_1378 = v_633 ^ v_673;
assign v_1379 = v_634 ^ v_674;
assign v_1380 = v_635 ^ v_675;
assign v_1381 = v_636 ^ v_676;
assign v_1382 = v_637 ^ v_677;
assign v_1383 = v_638 ^ v_678;
assign v_1384 = v_639 ^ v_679;
assign v_1385 = v_640 ^ v_680;
assign v_1387 = v_641 ^ v_681;
assign v_1388 = v_642 ^ v_682;
assign v_1389 = v_643 ^ v_683;
assign v_1390 = v_644 ^ v_684;
assign v_1391 = v_645 ^ v_685;
assign v_1392 = v_646 ^ v_686;
assign v_1393 = v_647 ^ v_687;
assign v_1394 = v_648 ^ v_688;
assign v_1395 = v_649 ^ v_689;
assign v_1396 = v_650 ^ v_690;
assign v_1397 = v_651 ^ v_691;
assign v_1398 = v_652 ^ v_692;
assign v_1399 = v_653 ^ v_693;
assign v_1400 = v_654 ^ v_694;
assign v_1401 = v_655 ^ v_695;
assign v_1402 = v_656 ^ v_696;
assign v_1403 = v_657 ^ v_697;
assign v_1404 = v_658 ^ v_698;
assign v_1405 = v_659 ^ v_699;
assign v_1406 = v_660 ^ v_700;
assign v_1408 = v_601 ^ v_701;
assign v_1409 = v_602 ^ v_702;
assign v_1410 = v_603 ^ v_703;
assign v_1411 = v_604 ^ v_704;
assign v_1412 = v_605 ^ v_705;
assign v_1413 = v_606 ^ v_706;
assign v_1414 = v_607 ^ v_707;
assign v_1415 = v_608 ^ v_708;
assign v_1416 = v_609 ^ v_709;
assign v_1417 = v_610 ^ v_710;
assign v_1418 = v_611 ^ v_711;
assign v_1419 = v_612 ^ v_712;
assign v_1420 = v_613 ^ v_713;
assign v_1421 = v_614 ^ v_714;
assign v_1422 = v_615 ^ v_715;
assign v_1423 = v_616 ^ v_716;
assign v_1424 = v_617 ^ v_717;
assign v_1425 = v_618 ^ v_718;
assign v_1426 = v_619 ^ v_719;
assign v_1427 = v_620 ^ v_720;
assign v_1430 = v_681 ^ v_721;
assign v_1431 = v_682 ^ v_722;
assign v_1432 = v_683 ^ v_723;
assign v_1433 = v_684 ^ v_724;
assign v_1434 = v_685 ^ v_725;
assign v_1435 = v_686 ^ v_726;
assign v_1436 = v_687 ^ v_727;
assign v_1437 = v_688 ^ v_728;
assign v_1438 = v_689 ^ v_729;
assign v_1439 = v_690 ^ v_730;
assign v_1440 = v_691 ^ v_731;
assign v_1441 = v_692 ^ v_732;
assign v_1442 = v_693 ^ v_733;
assign v_1443 = v_694 ^ v_734;
assign v_1444 = v_695 ^ v_735;
assign v_1445 = v_696 ^ v_736;
assign v_1446 = v_697 ^ v_737;
assign v_1447 = v_698 ^ v_738;
assign v_1448 = v_699 ^ v_739;
assign v_1449 = v_700 ^ v_740;
assign v_1451 = v_701 ^ v_741;
assign v_1452 = v_702 ^ v_742;
assign v_1453 = v_703 ^ v_743;
assign v_1454 = v_704 ^ v_744;
assign v_1455 = v_705 ^ v_745;
assign v_1456 = v_706 ^ v_746;
assign v_1457 = v_707 ^ v_747;
assign v_1458 = v_708 ^ v_748;
assign v_1459 = v_709 ^ v_749;
assign v_1460 = v_710 ^ v_750;
assign v_1461 = v_711 ^ v_751;
assign v_1462 = v_712 ^ v_752;
assign v_1463 = v_713 ^ v_753;
assign v_1464 = v_714 ^ v_754;
assign v_1465 = v_715 ^ v_755;
assign v_1466 = v_716 ^ v_756;
assign v_1467 = v_717 ^ v_757;
assign v_1468 = v_718 ^ v_758;
assign v_1469 = v_719 ^ v_759;
assign v_1470 = v_720 ^ v_760;
assign v_1472 = v_661 ^ v_761;
assign v_1473 = v_662 ^ v_762;
assign v_1474 = v_663 ^ v_763;
assign v_1475 = v_664 ^ v_764;
assign v_1476 = v_665 ^ v_765;
assign v_1477 = v_666 ^ v_766;
assign v_1478 = v_667 ^ v_767;
assign v_1479 = v_668 ^ v_768;
assign v_1480 = v_669 ^ v_769;
assign v_1481 = v_670 ^ v_770;
assign v_1482 = v_671 ^ v_771;
assign v_1483 = v_672 ^ v_772;
assign v_1484 = v_673 ^ v_773;
assign v_1485 = v_674 ^ v_774;
assign v_1486 = v_675 ^ v_775;
assign v_1487 = v_676 ^ v_776;
assign v_1488 = v_677 ^ v_777;
assign v_1489 = v_678 ^ v_778;
assign v_1490 = v_679 ^ v_779;
assign v_1491 = v_680 ^ v_780;
assign v_1495 = v_421 ^ v_361;
assign v_1496 = v_422 ^ v_362;
assign v_1497 = v_423 ^ v_363;
assign v_1498 = v_424 ^ v_364;
assign v_1499 = v_425 ^ v_365;
assign v_1500 = v_426 ^ v_366;
assign v_1501 = v_427 ^ v_367;
assign v_1502 = v_428 ^ v_368;
assign v_1503 = v_429 ^ v_369;
assign v_1504 = v_430 ^ v_370;
assign v_1505 = v_431 ^ v_371;
assign v_1506 = v_432 ^ v_372;
assign v_1507 = v_433 ^ v_373;
assign v_1508 = v_434 ^ v_374;
assign v_1509 = v_435 ^ v_375;
assign v_1510 = v_436 ^ v_376;
assign v_1511 = v_437 ^ v_377;
assign v_1512 = v_438 ^ v_378;
assign v_1513 = v_439 ^ v_379;
assign v_1514 = v_440 ^ v_380;
assign v_1516 = v_441 ^ v_381;
assign v_1517 = v_442 ^ v_382;
assign v_1518 = v_443 ^ v_383;
assign v_1519 = v_444 ^ v_384;
assign v_1520 = v_445 ^ v_385;
assign v_1521 = v_446 ^ v_386;
assign v_1522 = v_447 ^ v_387;
assign v_1523 = v_448 ^ v_388;
assign v_1524 = v_449 ^ v_389;
assign v_1525 = v_450 ^ v_390;
assign v_1526 = v_451 ^ v_391;
assign v_1527 = v_452 ^ v_392;
assign v_1528 = v_453 ^ v_393;
assign v_1529 = v_454 ^ v_394;
assign v_1530 = v_455 ^ v_395;
assign v_1531 = v_456 ^ v_396;
assign v_1532 = v_457 ^ v_397;
assign v_1533 = v_458 ^ v_398;
assign v_1534 = v_459 ^ v_399;
assign v_1535 = v_460 ^ v_400;
assign v_1537 = v_461 ^ v_401;
assign v_1538 = v_462 ^ v_402;
assign v_1539 = v_463 ^ v_403;
assign v_1540 = v_464 ^ v_404;
assign v_1541 = v_465 ^ v_405;
assign v_1542 = v_466 ^ v_406;
assign v_1543 = v_467 ^ v_407;
assign v_1544 = v_468 ^ v_408;
assign v_1545 = v_469 ^ v_409;
assign v_1546 = v_470 ^ v_410;
assign v_1547 = v_471 ^ v_411;
assign v_1548 = v_472 ^ v_412;
assign v_1549 = v_473 ^ v_413;
assign v_1550 = v_474 ^ v_414;
assign v_1551 = v_475 ^ v_415;
assign v_1552 = v_476 ^ v_416;
assign v_1553 = v_477 ^ v_417;
assign v_1554 = v_478 ^ v_418;
assign v_1555 = v_479 ^ v_419;
assign v_1556 = v_480 ^ v_420;
assign v_1559 = v_481 ^ v_361;
assign v_1560 = v_482 ^ v_362;
assign v_1561 = v_483 ^ v_363;
assign v_1562 = v_484 ^ v_364;
assign v_1563 = v_485 ^ v_365;
assign v_1564 = v_486 ^ v_366;
assign v_1565 = v_487 ^ v_367;
assign v_1566 = v_488 ^ v_368;
assign v_1567 = v_489 ^ v_369;
assign v_1568 = v_490 ^ v_370;
assign v_1569 = v_491 ^ v_371;
assign v_1570 = v_492 ^ v_372;
assign v_1571 = v_493 ^ v_373;
assign v_1572 = v_494 ^ v_374;
assign v_1573 = v_495 ^ v_375;
assign v_1574 = v_496 ^ v_376;
assign v_1575 = v_497 ^ v_377;
assign v_1576 = v_498 ^ v_378;
assign v_1577 = v_499 ^ v_379;
assign v_1578 = v_500 ^ v_380;
assign v_1580 = v_501 ^ v_381;
assign v_1581 = v_502 ^ v_382;
assign v_1582 = v_503 ^ v_383;
assign v_1583 = v_504 ^ v_384;
assign v_1584 = v_505 ^ v_385;
assign v_1585 = v_506 ^ v_386;
assign v_1586 = v_507 ^ v_387;
assign v_1587 = v_508 ^ v_388;
assign v_1588 = v_509 ^ v_389;
assign v_1589 = v_510 ^ v_390;
assign v_1590 = v_511 ^ v_391;
assign v_1591 = v_512 ^ v_392;
assign v_1592 = v_513 ^ v_393;
assign v_1593 = v_514 ^ v_394;
assign v_1594 = v_515 ^ v_395;
assign v_1595 = v_516 ^ v_396;
assign v_1596 = v_517 ^ v_397;
assign v_1597 = v_518 ^ v_398;
assign v_1598 = v_519 ^ v_399;
assign v_1599 = v_520 ^ v_400;
assign v_1601 = v_521 ^ v_401;
assign v_1602 = v_522 ^ v_402;
assign v_1603 = v_523 ^ v_403;
assign v_1604 = v_524 ^ v_404;
assign v_1605 = v_525 ^ v_405;
assign v_1606 = v_526 ^ v_406;
assign v_1607 = v_527 ^ v_407;
assign v_1608 = v_528 ^ v_408;
assign v_1609 = v_529 ^ v_409;
assign v_1610 = v_530 ^ v_410;
assign v_1611 = v_531 ^ v_411;
assign v_1612 = v_532 ^ v_412;
assign v_1613 = v_533 ^ v_413;
assign v_1614 = v_534 ^ v_414;
assign v_1615 = v_535 ^ v_415;
assign v_1616 = v_536 ^ v_416;
assign v_1617 = v_537 ^ v_417;
assign v_1618 = v_538 ^ v_418;
assign v_1619 = v_539 ^ v_419;
assign v_1620 = v_540 ^ v_420;
assign v_1623 = v_541 ^ v_361;
assign v_1624 = v_542 ^ v_362;
assign v_1625 = v_543 ^ v_363;
assign v_1626 = v_544 ^ v_364;
assign v_1627 = v_545 ^ v_365;
assign v_1628 = v_546 ^ v_366;
assign v_1629 = v_547 ^ v_367;
assign v_1630 = v_548 ^ v_368;
assign v_1631 = v_549 ^ v_369;
assign v_1632 = v_550 ^ v_370;
assign v_1633 = v_551 ^ v_371;
assign v_1634 = v_552 ^ v_372;
assign v_1635 = v_553 ^ v_373;
assign v_1636 = v_554 ^ v_374;
assign v_1637 = v_555 ^ v_375;
assign v_1638 = v_556 ^ v_376;
assign v_1639 = v_557 ^ v_377;
assign v_1640 = v_558 ^ v_378;
assign v_1641 = v_559 ^ v_379;
assign v_1642 = v_560 ^ v_380;
assign v_1644 = v_561 ^ v_381;
assign v_1645 = v_562 ^ v_382;
assign v_1646 = v_563 ^ v_383;
assign v_1647 = v_564 ^ v_384;
assign v_1648 = v_565 ^ v_385;
assign v_1649 = v_566 ^ v_386;
assign v_1650 = v_567 ^ v_387;
assign v_1651 = v_568 ^ v_388;
assign v_1652 = v_569 ^ v_389;
assign v_1653 = v_570 ^ v_390;
assign v_1654 = v_571 ^ v_391;
assign v_1655 = v_572 ^ v_392;
assign v_1656 = v_573 ^ v_393;
assign v_1657 = v_574 ^ v_394;
assign v_1658 = v_575 ^ v_395;
assign v_1659 = v_576 ^ v_396;
assign v_1660 = v_577 ^ v_397;
assign v_1661 = v_578 ^ v_398;
assign v_1662 = v_579 ^ v_399;
assign v_1663 = v_580 ^ v_400;
assign v_1665 = v_581 ^ v_401;
assign v_1666 = v_582 ^ v_402;
assign v_1667 = v_583 ^ v_403;
assign v_1668 = v_584 ^ v_404;
assign v_1669 = v_585 ^ v_405;
assign v_1670 = v_586 ^ v_406;
assign v_1671 = v_587 ^ v_407;
assign v_1672 = v_588 ^ v_408;
assign v_1673 = v_589 ^ v_409;
assign v_1674 = v_590 ^ v_410;
assign v_1675 = v_591 ^ v_411;
assign v_1676 = v_592 ^ v_412;
assign v_1677 = v_593 ^ v_413;
assign v_1678 = v_594 ^ v_414;
assign v_1679 = v_595 ^ v_415;
assign v_1680 = v_596 ^ v_416;
assign v_1681 = v_597 ^ v_417;
assign v_1682 = v_598 ^ v_418;
assign v_1683 = v_599 ^ v_419;
assign v_1684 = v_600 ^ v_420;
assign v_1687 = v_601 ^ v_361;
assign v_1688 = v_602 ^ v_362;
assign v_1689 = v_603 ^ v_363;
assign v_1690 = v_604 ^ v_364;
assign v_1691 = v_605 ^ v_365;
assign v_1692 = v_606 ^ v_366;
assign v_1693 = v_607 ^ v_367;
assign v_1694 = v_608 ^ v_368;
assign v_1695 = v_609 ^ v_369;
assign v_1696 = v_610 ^ v_370;
assign v_1697 = v_611 ^ v_371;
assign v_1698 = v_612 ^ v_372;
assign v_1699 = v_613 ^ v_373;
assign v_1700 = v_614 ^ v_374;
assign v_1701 = v_615 ^ v_375;
assign v_1702 = v_616 ^ v_376;
assign v_1703 = v_617 ^ v_377;
assign v_1704 = v_618 ^ v_378;
assign v_1705 = v_619 ^ v_379;
assign v_1706 = v_620 ^ v_380;
assign v_1708 = v_621 ^ v_381;
assign v_1709 = v_622 ^ v_382;
assign v_1710 = v_623 ^ v_383;
assign v_1711 = v_624 ^ v_384;
assign v_1712 = v_625 ^ v_385;
assign v_1713 = v_626 ^ v_386;
assign v_1714 = v_627 ^ v_387;
assign v_1715 = v_628 ^ v_388;
assign v_1716 = v_629 ^ v_389;
assign v_1717 = v_630 ^ v_390;
assign v_1718 = v_631 ^ v_391;
assign v_1719 = v_632 ^ v_392;
assign v_1720 = v_633 ^ v_393;
assign v_1721 = v_634 ^ v_394;
assign v_1722 = v_635 ^ v_395;
assign v_1723 = v_636 ^ v_396;
assign v_1724 = v_637 ^ v_397;
assign v_1725 = v_638 ^ v_398;
assign v_1726 = v_639 ^ v_399;
assign v_1727 = v_640 ^ v_400;
assign v_1729 = v_641 ^ v_401;
assign v_1730 = v_642 ^ v_402;
assign v_1731 = v_643 ^ v_403;
assign v_1732 = v_644 ^ v_404;
assign v_1733 = v_645 ^ v_405;
assign v_1734 = v_646 ^ v_406;
assign v_1735 = v_647 ^ v_407;
assign v_1736 = v_648 ^ v_408;
assign v_1737 = v_649 ^ v_409;
assign v_1738 = v_650 ^ v_410;
assign v_1739 = v_651 ^ v_411;
assign v_1740 = v_652 ^ v_412;
assign v_1741 = v_653 ^ v_413;
assign v_1742 = v_654 ^ v_414;
assign v_1743 = v_655 ^ v_415;
assign v_1744 = v_656 ^ v_416;
assign v_1745 = v_657 ^ v_417;
assign v_1746 = v_658 ^ v_418;
assign v_1747 = v_659 ^ v_419;
assign v_1748 = v_660 ^ v_420;
assign v_1751 = v_661 ^ v_361;
assign v_1752 = v_662 ^ v_362;
assign v_1753 = v_663 ^ v_363;
assign v_1754 = v_664 ^ v_364;
assign v_1755 = v_665 ^ v_365;
assign v_1756 = v_666 ^ v_366;
assign v_1757 = v_667 ^ v_367;
assign v_1758 = v_668 ^ v_368;
assign v_1759 = v_669 ^ v_369;
assign v_1760 = v_670 ^ v_370;
assign v_1761 = v_671 ^ v_371;
assign v_1762 = v_672 ^ v_372;
assign v_1763 = v_673 ^ v_373;
assign v_1764 = v_674 ^ v_374;
assign v_1765 = v_675 ^ v_375;
assign v_1766 = v_676 ^ v_376;
assign v_1767 = v_677 ^ v_377;
assign v_1768 = v_678 ^ v_378;
assign v_1769 = v_679 ^ v_379;
assign v_1770 = v_680 ^ v_380;
assign v_1772 = v_681 ^ v_381;
assign v_1773 = v_682 ^ v_382;
assign v_1774 = v_683 ^ v_383;
assign v_1775 = v_684 ^ v_384;
assign v_1776 = v_685 ^ v_385;
assign v_1777 = v_686 ^ v_386;
assign v_1778 = v_687 ^ v_387;
assign v_1779 = v_688 ^ v_388;
assign v_1780 = v_689 ^ v_389;
assign v_1781 = v_690 ^ v_390;
assign v_1782 = v_691 ^ v_391;
assign v_1783 = v_692 ^ v_392;
assign v_1784 = v_693 ^ v_393;
assign v_1785 = v_694 ^ v_394;
assign v_1786 = v_695 ^ v_395;
assign v_1787 = v_696 ^ v_396;
assign v_1788 = v_697 ^ v_397;
assign v_1789 = v_698 ^ v_398;
assign v_1790 = v_699 ^ v_399;
assign v_1791 = v_700 ^ v_400;
assign v_1793 = v_701 ^ v_401;
assign v_1794 = v_702 ^ v_402;
assign v_1795 = v_703 ^ v_403;
assign v_1796 = v_704 ^ v_404;
assign v_1797 = v_705 ^ v_405;
assign v_1798 = v_706 ^ v_406;
assign v_1799 = v_707 ^ v_407;
assign v_1800 = v_708 ^ v_408;
assign v_1801 = v_709 ^ v_409;
assign v_1802 = v_710 ^ v_410;
assign v_1803 = v_711 ^ v_411;
assign v_1804 = v_712 ^ v_412;
assign v_1805 = v_713 ^ v_413;
assign v_1806 = v_714 ^ v_414;
assign v_1807 = v_715 ^ v_415;
assign v_1808 = v_716 ^ v_416;
assign v_1809 = v_717 ^ v_417;
assign v_1810 = v_718 ^ v_418;
assign v_1811 = v_719 ^ v_419;
assign v_1812 = v_720 ^ v_420;
assign v_1815 = v_721 ^ v_361;
assign v_1816 = v_722 ^ v_362;
assign v_1817 = v_723 ^ v_363;
assign v_1818 = v_724 ^ v_364;
assign v_1819 = v_725 ^ v_365;
assign v_1820 = v_726 ^ v_366;
assign v_1821 = v_727 ^ v_367;
assign v_1822 = v_728 ^ v_368;
assign v_1823 = v_729 ^ v_369;
assign v_1824 = v_730 ^ v_370;
assign v_1825 = v_731 ^ v_371;
assign v_1826 = v_732 ^ v_372;
assign v_1827 = v_733 ^ v_373;
assign v_1828 = v_734 ^ v_374;
assign v_1829 = v_735 ^ v_375;
assign v_1830 = v_736 ^ v_376;
assign v_1831 = v_737 ^ v_377;
assign v_1832 = v_738 ^ v_378;
assign v_1833 = v_739 ^ v_379;
assign v_1834 = v_740 ^ v_380;
assign v_1836 = v_741 ^ v_381;
assign v_1837 = v_742 ^ v_382;
assign v_1838 = v_743 ^ v_383;
assign v_1839 = v_744 ^ v_384;
assign v_1840 = v_745 ^ v_385;
assign v_1841 = v_746 ^ v_386;
assign v_1842 = v_747 ^ v_387;
assign v_1843 = v_748 ^ v_388;
assign v_1844 = v_749 ^ v_389;
assign v_1845 = v_750 ^ v_390;
assign v_1846 = v_751 ^ v_391;
assign v_1847 = v_752 ^ v_392;
assign v_1848 = v_753 ^ v_393;
assign v_1849 = v_754 ^ v_394;
assign v_1850 = v_755 ^ v_395;
assign v_1851 = v_756 ^ v_396;
assign v_1852 = v_757 ^ v_397;
assign v_1853 = v_758 ^ v_398;
assign v_1854 = v_759 ^ v_399;
assign v_1855 = v_760 ^ v_400;
assign v_1857 = v_761 ^ v_401;
assign v_1858 = v_762 ^ v_402;
assign v_1859 = v_763 ^ v_403;
assign v_1860 = v_764 ^ v_404;
assign v_1861 = v_765 ^ v_405;
assign v_1862 = v_766 ^ v_406;
assign v_1863 = v_767 ^ v_407;
assign v_1864 = v_768 ^ v_408;
assign v_1865 = v_769 ^ v_409;
assign v_1866 = v_770 ^ v_410;
assign v_1867 = v_771 ^ v_411;
assign v_1868 = v_772 ^ v_412;
assign v_1869 = v_773 ^ v_413;
assign v_1870 = v_774 ^ v_414;
assign v_1871 = v_775 ^ v_415;
assign v_1872 = v_776 ^ v_416;
assign v_1873 = v_777 ^ v_417;
assign v_1874 = v_778 ^ v_418;
assign v_1875 = v_779 ^ v_419;
assign v_1876 = v_780 ^ v_420;
assign x_1 = v_1880 | ~v_1169;
assign o_1 = x_1;
endmodule
