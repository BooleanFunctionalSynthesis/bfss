// Generated using findDep.cpp 
module small-bug1-fixpoint-3 (v_1, v_2, v_3, v_4, v_5, v_6, v_7, v_8, v_9, v_10, v_11, v_12, v_13, v_14, v_15, v_16, v_17, v_18, v_19, o_1);
input v_1;
input v_2;
input v_3;
input v_4;
input v_5;
input v_6;
input v_7;
input v_8;
input v_9;
input v_10;
input v_11;
input v_12;
input v_13;
input v_14;
input v_15;
input v_16;
input v_17;
input v_18;
input v_19;
output o_1;
wire v_20;
wire v_21;
wire v_22;
wire v_23;
wire v_24;
wire v_25;
wire v_26;
wire v_27;
wire v_28;
wire v_29;
wire v_30;
wire v_31;
wire v_32;
wire v_33;
wire v_34;
wire v_35;
wire v_36;
wire v_37;
wire v_38;
wire v_39;
wire v_40;
wire v_41;
wire v_42;
wire v_43;
wire v_44;
wire v_45;
wire v_46;
wire v_47;
wire v_48;
wire v_49;
wire v_50;
wire v_51;
wire v_52;
wire v_53;
wire v_54;
wire x_1;
assign v_20 = ~v_1 & v_7;
assign v_21 = ~v_6 & v_20;
assign v_24 = ~v_2 & v_5;
assign v_25 = ~v_9 & v_24;
assign v_28 = ~v_3 & v_8;
assign v_29 = ~v_11 & v_28;
assign v_32 = v_53 & v_54;
assign v_33 = ~v_12 & v_17;
assign v_34 = ~v_16 & v_33;
assign v_37 = ~v_13 & v_15;
assign v_38 = ~v_19 & v_37;
assign v_41 = ~v_12 & ~v_13 & ~v_14 & ~v_36 & ~v_40;
assign v_44 = ~v_42 & ~v_43;
assign v_47 = ~v_45 & ~v_46;
assign v_50 = ~v_48 & ~v_49;
assign v_52 = v_41 & v_51;
assign v_53 = ~v_1 & ~v_2 & ~v_3 & ~v_4 & ~v_23;
assign v_54 = ~v_27 & ~v_31;
assign v_22 = v_6 | v_21;
assign v_26 = v_9 | v_25;
assign v_30 = v_11 | v_29;
assign v_35 = v_16 | v_34;
assign v_39 = v_19 | v_38;
assign v_51 = v_44 | v_47 | v_50;
assign v_23 = v_22 ^ v_5;
assign v_27 = v_26 ^ v_8;
assign v_31 = v_30 ^ v_10;
assign v_36 = v_35 ^ v_15;
assign v_40 = v_39 ^ v_18;
assign v_42 = v_12 ^ v_4;
assign v_43 = v_17 ^ v_10;
assign v_45 = v_13 ^ v_4;
assign v_46 = v_15 ^ v_10;
assign v_48 = v_14 ^ v_4;
assign v_49 = v_18 ^ v_10;
assign x_1 = v_52 | ~v_32;
assign o_1 = x_1;
endmodule
