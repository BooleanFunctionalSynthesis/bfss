// Verilog file written by procedure writeCombinationalCircuitInVerilog
//Skolem functions to be generated for i_ variables
module neclaftp4001_all_bit_differing_from_cycle ( i_1, i_2, i_3, i_4, i_5, i_6, i_7, i_8, i_9, i_10, i_11, i_12, i_13, i_14, i_15, i_16, i_17, i_18, i_19, i_20, i_21, i_22, i_23, i_24, i_25, i_26, i_27, i_28, i_29, i_30, i_31, i_32, x_33, x_34, x_35, x_36, x_37, x_38, x_39, x_40, x_41, x_42, x_43, x_44, x_45, x_46, x_47, x_48, x_49, x_50, x_51, x_52, x_53, x_54, x_55, x_56, x_57, x_58, x_59, x_60, x_61, x_62, x_63, x_64, x_65, x_66, x_67, x_68, x_69, x_70, x_71, x_72, x_73, x_74, x_75, x_76, x_77, x_78, x_79, x_80, x_81, x_82, x_83, x_84, x_85, x_86, x_87, x_88, x_89, x_90, x_91, x_92, x_93, x_94, x_95, x_96, x_97, x_98, x_99, x_100, x_101, x_102, x_103, x_104, x_105, x_106, x_107, x_108, x_109, x_110, x_111, x_112, x_113, x_114, x_115, x_116, x_117, x_118, x_119, x_120, x_121, x_122, x_123, x_124, x_125, x_126, x_127, x_128, x_129, x_130, x_131, x_132, x_133, x_134, x_135, x_136, x_137, x_138, x_139, x_140, x_141, x_142, x_143, x_144, x_145, x_146, x_147, x_148, x_149, x_150, x_151, x_152, x_153, x_154, x_155, x_156, x_157, x_158, x_159, x_160, x_161, x_162, x_163, x_164, x_165, x_166, x_167, x_168, x_169, x_170, x_171, x_172, x_173, x_174, x_175, x_176, x_177, x_178, x_179, x_180, x_181, x_182, x_183, x_184, x_185, x_186, x_187, x_188, x_189, x_190, x_191, x_192, x_193, x_194, x_195, x_196, x_197, x_198, x_199, x_200, x_201, x_202, x_203, x_204, x_205, x_206, x_207, x_208, x_209, x_210, x_211, x_212, x_213, x_214, x_215, x_216, x_217, x_218, x_219, x_220, x_221, x_222, x_223, x_224, x_225, x_226, x_227, x_228, x_229, x_230, x_231, x_232, x_233, x_234, x_235, x_236, x_237, x_238, x_239, x_240, x_241, x_242, x_243, x_244, x_245, x_246, x_247, x_248, x_249, x_250, x_251, x_252, x_253, x_254, x_255, x_256, x_257, x_258, x_259, x_260, x_261, x_262, x_263, x_264, x_265, x_266, x_267, x_268, x_269, x_270, x_271, x_272, x_273, x_274, x_275, x_276, x_277, x_278, x_279, x_280, x_281, x_282, x_283, x_284, x_285, x_286, x_287, x_288, x_289, x_290, x_291, x_292, x_293, x_294, x_295, x_296, x_297, x_298, x_299, x_300, x_301, x_302, x_303, x_304, x_305, x_306, x_307, x_308, x_309, x_310, x_311, x_312, x_313, x_314, x_315, x_316, x_317, x_318, x_319, x_320, x_321, x_322, x_323, x_324, x_325, x_326, x_327, x_328, x_329, x_330, x_331, x_332, x_333, x_334, x_335, x_336, x_337, x_338, x_339, x_340, x_341, x_342, x_343, x_344, x_345, x_346, x_347, x_348, x_349, x_350, x_351, x_352, x_353, x_354, x_355, x_356, x_357, x_358, x_359, x_360, x_361, x_362, x_363, x_364, x_365, x_366, x_367, x_368, x_369, x_370, x_371, x_372, x_373, x_374, x_375, x_376, x_377, x_378, x_379, x_380, x_381, x_382, x_383, x_384, x_385, x_386, x_387, x_388, x_389, x_390, x_391, x_392, x_393, x_394, x_395, x_396, x_397, x_398, x_399, x_400, x_401, x_402, x_403, x_404, x_405, x_406, x_407, x_408, x_409, x_410, x_411, x_412, x_413, x_414, x_415, x_416, x_417, x_418, x_419, x_420, x_421, x_422, x_423, x_424, x_425, x_426, x_427, x_428, x_429, x_430, x_431, x_432, x_433, x_434, x_435, x_436, x_437, x_438, x_439, x_440, x_441, x_442, x_443, x_444, x_445, x_446, x_447, x_448, x_449, x_450, x_451, x_452, x_453, x_454, x_455, x_456, x_457, x_458, x_459, x_460, x_461, x_462, x_463, x_464, x_465, x_466, x_467, x_468, x_469, x_470, x_471, x_472, x_473, x_474, x_475, x_476, x_477, x_478, x_479, x_480, x_481, x_482, x_483, x_484, x_485, x_486, x_487, x_488, x_489, x_490, x_491, x_492, x_493, x_494, x_495, x_496, x_497, x_498, x_499, x_500, x_501, x_502, x_503, x_504, x_505, x_506, x_507, x_508, x_509, x_510, x_511, x_512, x_513, x_514, x_515, x_516, x_517, x_518, x_519, x_520, x_521, x_522, x_523, x_524, x_525, x_526, x_527, x_528, x_529, x_530, x_531, x_532, x_533, x_534, x_535, x_536, x_537, x_538, x_539, x_540, x_541, x_542, x_543, x_544, x_545, x_546, x_547, x_548, x_549, x_550, x_551, x_552, x_553, x_554, x_555, x_556, x_557, x_558, x_559, x_560, x_561, x_562, x_563, x_564, x_565, x_566, x_567, x_568, x_569, x_570, x_571, x_572, x_573, x_574, x_575, x_576, x_577, x_578, x_579, x_580, x_581, x_582, x_583, x_584, x_585, x_586, x_587, x_588, x_589, x_590, x_591, x_592, x_593, x_594, x_595, x_596, x_597, x_598, x_599, x_600, x_601, x_602, x_603, x_604, x_605, x_606, x_607, x_608, x_609, x_610, x_611, x_612, x_613, x_614, x_615, x_616, x_617, x_618, x_619, x_620, x_621, x_622, x_623, x_624, x_625, x_626, x_627, x_628, x_629, x_630, x_631, x_632, x_633, x_634, x_635, x_636, x_637, x_638, x_639, x_640, x_641, x_642, x_643, x_644, x_645, x_646, x_647, x_648, x_649, x_650, x_651, x_652, x_653, x_654, x_655, x_656, x_657, x_658, x_659, x_660, x_661, x_662, x_663, x_664, x_665, x_666, x_667, x_668, x_669, x_670, x_671, x_672, x_673, x_674, x_675, x_676, x_677, x_678, x_679, x_680, x_681, x_682, x_683, x_684, x_685, x_686, x_687, x_688, x_689, x_690, x_691, x_692, x_693, x_694, x_695, x_696, x_697, x_698, x_699, x_700, x_701, x_702, x_703, x_704, x_705, x_706, x_707, x_708, x_709, x_710, x_711, x_712, x_713, x_714, x_715, x_716, x_717, x_718, x_719, x_720, x_721, x_722, x_723, x_724, x_725, x_726, x_727, x_728, x_729, x_730, x_731, x_732, x_733, x_734, x_735, x_736, x_737, x_738, x_739, x_740, x_741, x_742, x_743, x_744, x_745, x_746, x_747, x_748, x_749, x_750, x_751, x_752, x_753, x_754, x_755, x_756, x_757, x_758, x_759, x_760, x_761, x_762, x_763, x_764, x_765, x_766, x_767, x_768, x_769, x_770, x_771, x_772, x_773, x_774, x_775, x_776, x_777, x_778, x_779, x_780, x_781, x_782, x_783, x_784, x_785, x_786, x_787, x_788, x_789, x_790, x_791, x_792, x_793, x_794, x_795, x_796, x_797, x_798, x_799, x_800, x_801, x_802, x_803, x_804, x_805, x_806, x_807, x_808, x_809, x_810, x_811, x_812, x_813, x_814, x_815, x_816, x_817, x_818, x_819, x_820, x_821, x_822, x_823, x_824, x_825, x_826, x_827, x_828, x_829, x_830, x_831, x_832, x_833, x_834, x_835, x_836, x_837, x_838, x_839, x_840, x_841, x_842, x_843, x_844, x_845, x_846, x_847, x_848, x_849, x_850, x_851, x_852, x_853, x_854, x_855, x_856, x_857, x_858, x_859, x_860, x_861, x_862, x_863, x_864, x_865, x_866, x_867, x_868, x_869, x_870, x_871, x_872, x_873, x_874, x_875, x_876, x_877, x_878, x_879, x_880, x_881, x_882, x_883, x_884, x_885, x_886, x_887, x_888, x_889, x_890, x_891, x_892, x_893, x_894, x_895, x_896, x_897, x_898, x_899, x_900, x_901, x_902, x_903, x_904, x_905, x_906, x_907, x_908, x_909, x_910, x_911, x_912, x_913, x_914, x_915, x_916, x_917, x_918, x_919, x_920, x_921, x_922, x_923, x_924, x_925, x_926, x_927, x_928, x_929, x_930, x_931, x_932, x_933, x_934, x_935, x_936, x_937, x_938, x_939, x_940, x_941, x_942, x_943, x_944, x_945, x_946, x_947, x_948, x_949, x_950, x_951, x_952, x_953, x_954, x_955, x_956, x_957, x_958, x_959, x_960, x_961, x_962, x_963, x_964, x_965, x_966, x_967, x_968, x_969, x_970, x_971, x_972, x_973, x_974, x_975, x_976, x_977, x_978, x_979, x_980, x_981, x_982, x_983, x_984, x_985, x_986, x_987, x_988, x_989, x_990, x_991, x_992, x_993, x_994, x_995, x_996, x_997, x_998, x_999, x_1000, x_1001, x_1002, x_1003, x_1004, x_1005, x_1006, x_1007, x_1008, x_1009, x_1010, x_1011, x_1012, x_1013, x_1014, x_1015, x_1016, x_1017, x_1018, x_1019, x_1020, x_1021, x_1022, x_1023, x_1024, x_1025, x_1026, x_1027, x_1028, x_1029, x_1030, x_1031, x_1032, x_1033, x_1034, x_1035, x_1036, x_1037, x_1038, x_1039, x_1040, x_1041, x_1042, x_1043, x_1044, x_1045, x_1046, x_1047, x_1048, x_1049, x_1050, x_1051, x_1052, x_1053, x_1054, x_1055, x_1056, x_1057, x_1058, x_1059, x_1060, x_1061, x_1062, x_1063, x_1064, x_1065, x_1066, x_1067, x_1068, x_1069, x_1070, x_1071, x_1072, x_1073, x_1074, x_1075, x_1076, x_1077, x_1078, x_1079, x_1080, x_1081, x_1082, x_1083, x_1084, x_1085, x_1086, x_1087, x_1088, x_1089, x_1090, x_1091, x_1092, x_1093, x_1094, x_1095, x_1096, x_1097, x_1098, x_1099, x_1100, x_1101, x_1102, x_1103, x_1104, x_1105, x_1106, x_1107, x_1108, x_1109, x_1110, x_1111, x_1112, x_1113, x_1114, x_1115, x_1116, x_1117, x_1118, x_1119, x_1120, x_1121, x_1122, x_1123, x_1124, x_1125, x_1126, x_1127, x_1128, x_1129, x_1130, x_1131, x_1132, x_1133, x_1134, x_1135, x_1136, x_1137, x_1138, x_1139, x_1140, x_1141, x_1142, x_1143, x_1144, x_1145, x_1146, x_1147, x_1148, x_1149, x_1150, x_1151, x_1152, x_1153, x_1154, x_1155, x_1156, x_1157, x_1158, x_1159, x_1160, x_1161, x_1162, x_1163, x_1164, x_1165, x_1166, x_1167, x_1168, x_1169, x_1170, x_1171, x_1172, x_1173, x_1174, x_1175, x_1176, x_1177, x_1178, x_1179, x_1180, x_1181, x_1182, x_1183, x_1184, x_1185, x_1186, x_1187, x_1188, x_1189, x_1190, x_1191, x_1192, x_1193, x_1194, x_1195, x_1196, x_1197, x_1198, x_1199, x_1200, x_1201, x_1202, x_1203, x_1204, x_1205, x_1206, x_1207, x_1208, x_1209, x_1210, x_1211, x_1212, x_1213, x_1214, x_1215, x_1216, x_1217, x_1218, x_1219, x_1220, x_1221, x_1222, x_1223, x_1224, x_1225, x_1226, x_1227, x_1228, x_1229, x_1230, x_1231, x_1232, x_1233, x_1234, x_1235, x_1236, x_1237, x_1238, x_1239, x_1240, x_1241, x_1242, x_1243, x_1244, x_1245, x_1246, x_1247, x_1248, x_1249, x_1250, x_1251, x_1252, x_1253, x_1254, x_1255, x_1256, x_1257, x_1258, x_1259, x_1260, x_1261, x_1262, x_1263, x_1264, x_1265, x_1266, x_1267, x_1268, x_1269, x_1270, x_1271, x_1272, x_1273, x_1274, x_1275, x_1276, x_1277, x_1278, x_1279, x_1280, x_1281, x_1282, x_1283, x_1284, x_1285, x_1286, x_1287, x_1288, x_1289, x_1290, x_1291, x_1292, x_1293, x_1294, x_1295, x_1296, x_1297, x_1298, x_1299, x_1300, x_1301, x_1302, x_1303, x_1304, x_1305, x_1306, x_1307, x_1308, x_1309, x_1310, x_1311, x_1312, x_1313, x_1314, x_1315, x_1316, x_1317, x_1318, x_1319, x_1320, x_1321, x_1322, x_1323, x_1324, x_1325, x_1326, x_1327, x_1328, x_1329, x_1330, x_1331, x_1332, x_1333, x_1334, x_1335, x_1336, x_1337, x_1338, x_1339, x_1340, x_1341, x_1342, x_1343, x_1344, x_1345, x_1346, x_1347, x_1348, x_1349, x_1350, x_1351, x_1352, x_1353, x_1354, x_1355, x_1356, x_1357, x_1358, x_1359, x_1360, x_1361, x_1362, x_1363, x_1364, x_1365, x_1366, x_1367, x_1368, x_1369, x_1370, x_1371, x_1372, x_1373, x_1374, x_1375, x_1376, x_1377, x_1378, x_1379, x_1380, x_1381, x_1382, x_1383, x_1384, x_1385, x_1386, x_1387, x_1388, x_1389, x_1390, x_1391, x_1392, x_1393, x_1394, x_1395, x_1396, x_1397, x_1398, x_1399, x_1400, x_1401, x_1402, x_1403, x_1404, x_1405, x_1406, x_1407, x_1408, x_1409, x_1410, x_1411, x_1412, x_1413, x_1414, x_1415, x_1416, x_1417, x_1418, x_1419, x_1420, x_1421, x_1422, x_1423, x_1424, x_1425, x_1426, x_1427, x_1428, x_1429, x_1430, x_1431, x_1432, x_1433, x_1434, x_1435, x_1436, x_1437, x_1438, x_1439, x_1440, x_1441, x_1442, x_1443, x_1444, x_1445, x_1446, x_1447, x_1448, x_1449, x_1450, x_1451, x_1452, x_1453, x_1454, x_1455, x_1456, x_1457, x_1458, x_1459, x_1460, x_1461, x_1462, x_1463, x_1464, x_1465, x_1466, x_1467, x_1468, x_1469, x_1470, x_1471, x_1472, x_1473, x_1474, x_1475, x_1476, x_1477, x_1478, x_1479, x_1480, x_1481, x_1482, x_1483, x_1484, x_1485, x_1486, x_1487, x_1488, x_1489, x_1490, x_1491, x_1492, x_1493, x_1494, x_1495, x_1496, x_1497, x_1498, x_1499, x_1500, x_1501, x_1502, x_1503, x_1504, x_1505, x_1506, x_1507, x_1508, x_1509, x_1510, x_1511, x_1512, x_1513, x_1514, x_1515, x_1516, x_1517, x_1518, x_1519, x_1520, x_1521, x_1522, x_1523, x_1524, x_1525, x_1526, x_1527, x_1528, x_1529, x_1530, x_1531, x_1532, x_1533, x_1534, x_1535, x_1536, x_1537, x_1538, x_1539, x_1540, x_1541, x_1542, x_1543, x_1544, x_1545, x_1546, x_1547, x_1548, x_1549, x_1550, x_1551, x_1552, x_1553, x_1554, x_1555, x_1556, x_1557, x_1558, x_1559, x_1560, x_1561, x_1562, x_1563, x_1564, x_1565, x_1566, x_1567, x_1568, x_1569, x_1570, x_1571, x_1572, x_1573, x_1574, x_1575, x_1576, x_1577, x_1578, x_1579, x_1580, x_1581, x_1582, x_1583, x_1584, x_1585, x_1586, x_1587, x_1588, x_1589, x_1590, x_1591, x_1592, x_1593, x_1594, x_1595, x_1596, x_1597, x_1598, x_1599, x_1600, x_1601, x_1602, x_1603, x_1604, x_1605, x_1606, x_1607, x_1608, x_1609, x_1610, x_1611, x_1612, x_1613, x_1614, x_1615, x_1616, x_1617, x_1618, x_1619, x_1620, x_1621, x_1622, x_1623, x_1624, x_1625, x_1626, x_1627, x_1628, x_1629, x_1630, x_1631, x_1632, x_1633, x_1634, x_1635, x_1636, x_1637, x_1638, x_1639, x_1640, x_1641, x_1642, x_1643, x_1644, x_1645, x_1646, x_1647, x_1648, x_1649, x_1650, x_1651, x_1652, x_1653, x_1654, x_1655, x_1656, x_1657, x_1658, x_1659, x_1660, x_1661, x_1662, x_1663, x_1664, x_1665, x_1666, x_1667, x_1668, x_1669, x_1670, x_1671, x_1672, x_1673, x_1674, x_1675, x_1676, x_1677, x_1678, x_1679, x_1680, x_1681, x_1682, x_1683, x_1684, x_1685, x_1686, x_1687, x_1688, x_1689, x_1690, x_1691, x_1692, x_1693, x_1694, x_1695, x_1696, x_1697, x_1698, x_1699, x_1700, x_1701, x_1702, x_1703, x_1704, x_1705, x_1706, x_1707, x_1708, x_1709, x_1710, x_1711, x_1712, x_1713, x_1714, x_1715, x_1716, x_1717, x_1718, x_1719, x_1720, x_1721, x_1722, x_1723, x_1724, x_1725, x_1726, x_1727, x_1728, x_1729, x_1730, x_1731, x_1732, x_1733, x_1734, x_1735, x_1736, x_1737, x_1738, x_1739, x_1740, x_1741, x_1742, x_1743, x_1744, x_1745, x_1746, x_1747, x_1748, x_1749, x_1750, x_1751, x_1752, x_1753, x_1754, x_1755, x_1756, x_1757, x_1758, x_1759, x_1760, x_1761, x_1762, x_1763, x_1764, x_1765, x_1766, x_1767, x_1768, x_1769, x_1770, x_1771, x_1772, x_1773, x_1774, x_1775, x_1776, x_1777, x_1778, x_1779, x_1780, x_1781, x_1782, x_1783, x_1784, x_1785, x_1786, x_1787, x_1788, x_1789, x_1790, x_1791, x_1792, x_1793, x_1794, x_1795, x_1796, x_1797, x_1798, x_1799, x_1800, x_1801, x_1802, x_1803, x_1804, x_1805, x_1806, x_1807, x_1808, x_1809, x_1810, x_1811, x_1812, x_1813, x_1814, x_1815, x_1816, x_1817, x_1818, x_1819, x_1820, x_1821, x_1822, x_1823, x_1824, x_1825, x_1826, x_1827, x_1828, x_1829, x_1830, x_1831, x_1832, x_1833, x_1834, x_1835, x_1836, x_1837, x_1838, x_1839, x_1840, x_1841, x_1842, x_1843, x_1844, x_1845, x_1846, x_1847, x_1848, x_1849, x_1850, x_1851, x_1852, x_1853, x_1854, x_1855, x_1856, x_1857, x_1858, x_1859, x_1860, x_1861, x_1862, x_1863, x_1864, x_1865, x_1866, x_1867, x_1868, x_1869, x_1870, x_1871, x_1872, x_1873, x_1874, x_1875, x_1876, x_1877, x_1878, x_1879, x_1880, x_1881, x_1882, x_1883, x_1884, x_1885, x_1886, x_1887, x_1888, x_1889, x_1890, x_1891, x_1892, x_1893, x_1894, x_1895, x_1896, x_1897, x_1898, x_1899, x_1900, x_1901, x_1902, x_1903, x_1904, x_1905, x_1906, x_1907, x_1908, x_1909, x_1910, x_1911, x_1912, x_1913, x_1914, x_1915, x_1916, x_1917, x_1918, x_1919, x_1920, x_1921, x_1922, x_1923, x_1924, x_1925, x_1926, x_1927, x_1928, x_1929, x_1930, x_1931, x_1932, x_1933, x_1934, x_1935, x_1936, x_1937, x_1938, x_1939, x_1940, x_1941, x_1942, x_1943, x_1944, x_1945, x_1946, x_1947, x_1948, x_1949, x_1950, x_1951, x_1952, x_1953, x_1954, x_1955, x_1956, x_1957, x_1958, x_1959, x_1960, x_1961, x_1962, x_1963, x_1964, x_1965, x_1966, x_1967, x_1968, x_1969, x_1970, x_1971, x_1972, x_1973, x_1974, x_1975, x_1976, x_1977, x_1978, x_1979, x_1980, x_1981, x_1982, x_1983, x_1984, x_1985, x_1986, x_1987, x_1988, x_1989, x_1990, x_1991, x_1992, x_1993, x_1994, x_1995, x_1996, x_1997, x_1998, x_1999, x_2000, x_2001, x_2002, x_2003, x_2004, x_2005, x_2006, x_2007, x_2008, x_2009, x_2010, x_2011, x_2012, x_2013, x_2014, x_2015, x_2016, x_2017, x_2018, x_2019, x_2020, x_2021, x_2022, x_2023, x_2024, x_2025, x_2026, x_2027, x_2028, x_2029, x_2030, x_2031, x_2032, x_2033, x_2034, x_2035, x_2036, x_2037, x_2038, x_2039, x_2040, x_2041, x_2042, x_2043, x_2044, x_2045, x_2046, x_2047, x_2048, x_2049, x_2050, x_2051, x_2052, x_2053, x_2054, x_2055, x_2056, x_2057, x_2058, x_2059, x_2060, x_2061, x_2062, x_2063, x_2064, x_2065, x_2066, x_2067, x_2068, x_2069, x_2070, x_2071, x_2072, x_2073, x_2074, x_2075, x_2076, x_2077, x_2078, x_2079, x_2080, x_2081, x_2082, x_2083, x_2084, x_2085, x_2086, x_2087, x_2088, x_2089, x_2090, x_2091, x_2092, x_2093, x_2094, x_2095, x_2096, x_2097, x_2098, x_2099, x_2100, x_2101, x_2102, x_2103, x_2104, x_2105, x_2106, x_2107, x_2108, x_2109, x_2110, x_2111, x_2112, x_2113, x_2114, x_2115, x_2116, x_2117, x_2118, x_2119, x_2120, x_2121, x_2122, x_2123, x_2124, x_2125, x_2126, x_2127, x_2128, x_2129, x_2130, x_2131, x_2132, x_2133, x_2134, x_2135, x_2136, x_2137, x_2138, x_2139, x_2140, x_2141, x_2142, x_2143, x_2144, x_2145, x_2146, x_2147, x_2148, x_2149, x_2150, x_2151, x_2152, x_2153, x_2154, x_2155, x_2156, x_2157, x_2158, x_2159, x_2160, x_2161, x_2162, x_2163, x_2164, x_2165, x_2166, x_2167, x_2168, x_2169, x_2170, x_2171, x_2172, x_2173, x_2174, x_2175, x_2176, x_2177, x_2178, x_2179, x_2180, x_2181, x_2182, x_2183, x_2184, x_2185, x_2186, x_2187, x_2188, x_2189, x_2190, x_2191, x_2192, x_2193, x_2194, x_2195, x_2196, x_2197, x_2198, x_2199, x_2200, x_2201, x_2202, x_2203, x_2204, x_2205, x_2206, x_2207, x_2208, x_2209, x_2210, x_2211, x_2212, x_2213, x_2214, x_2215, x_2216, x_2217, x_2218, x_2219, x_2220, o_1 );
input i_1;
input i_2;
input i_3;
input i_4;
input i_5;
input i_6;
input i_7;
input i_8;
input i_9;
input i_10;
input i_11;
input i_12;
input i_13;
input i_14;
input i_15;
input i_16;
input i_17;
input i_18;
input i_19;
input i_20;
input i_21;
input i_22;
input i_23;
input i_24;
input i_25;
input i_26;
input i_27;
input i_28;
input i_29;
input i_30;
input i_31;
input i_32;
input x_33;
input x_34;
input x_35;
input x_36;
input x_37;
input x_38;
input x_39;
input x_40;
input x_41;
input x_42;
input x_43;
input x_44;
input x_45;
input x_46;
input x_47;
input x_48;
input x_49;
input x_50;
input x_51;
input x_52;
input x_53;
input x_54;
input x_55;
input x_56;
input x_57;
input x_58;
input x_59;
input x_60;
input x_61;
input x_62;
input x_63;
input x_64;
input x_65;
input x_66;
input x_67;
input x_68;
input x_69;
input x_70;
input x_71;
input x_72;
input x_73;
input x_74;
input x_75;
input x_76;
input x_77;
input x_78;
input x_79;
input x_80;
input x_81;
input x_82;
input x_83;
input x_84;
input x_85;
input x_86;
input x_87;
input x_88;
input x_89;
input x_90;
input x_91;
input x_92;
input x_93;
input x_94;
input x_95;
input x_96;
input x_97;
input x_98;
input x_99;
input x_100;
input x_101;
input x_102;
input x_103;
input x_104;
input x_105;
input x_106;
input x_107;
input x_108;
input x_109;
input x_110;
input x_111;
input x_112;
input x_113;
input x_114;
input x_115;
input x_116;
input x_117;
input x_118;
input x_119;
input x_120;
input x_121;
input x_122;
input x_123;
input x_124;
input x_125;
input x_126;
input x_127;
input x_128;
input x_129;
input x_130;
input x_131;
input x_132;
input x_133;
input x_134;
input x_135;
input x_136;
input x_137;
input x_138;
input x_139;
input x_140;
input x_141;
input x_142;
input x_143;
input x_144;
input x_145;
input x_146;
input x_147;
input x_148;
input x_149;
input x_150;
input x_151;
input x_152;
input x_153;
input x_154;
input x_155;
input x_156;
input x_157;
input x_158;
input x_159;
input x_160;
input x_161;
input x_162;
input x_163;
input x_164;
input x_165;
input x_166;
input x_167;
input x_168;
input x_169;
input x_170;
input x_171;
input x_172;
input x_173;
input x_174;
input x_175;
input x_176;
input x_177;
input x_178;
input x_179;
input x_180;
input x_181;
input x_182;
input x_183;
input x_184;
input x_185;
input x_186;
input x_187;
input x_188;
input x_189;
input x_190;
input x_191;
input x_192;
input x_193;
input x_194;
input x_195;
input x_196;
input x_197;
input x_198;
input x_199;
input x_200;
input x_201;
input x_202;
input x_203;
input x_204;
input x_205;
input x_206;
input x_207;
input x_208;
input x_209;
input x_210;
input x_211;
input x_212;
input x_213;
input x_214;
input x_215;
input x_216;
input x_217;
input x_218;
input x_219;
input x_220;
input x_221;
input x_222;
input x_223;
input x_224;
input x_225;
input x_226;
input x_227;
input x_228;
input x_229;
input x_230;
input x_231;
input x_232;
input x_233;
input x_234;
input x_235;
input x_236;
input x_237;
input x_238;
input x_239;
input x_240;
input x_241;
input x_242;
input x_243;
input x_244;
input x_245;
input x_246;
input x_247;
input x_248;
input x_249;
input x_250;
input x_251;
input x_252;
input x_253;
input x_254;
input x_255;
input x_256;
input x_257;
input x_258;
input x_259;
input x_260;
input x_261;
input x_262;
input x_263;
input x_264;
input x_265;
input x_266;
input x_267;
input x_268;
input x_269;
input x_270;
input x_271;
input x_272;
input x_273;
input x_274;
input x_275;
input x_276;
input x_277;
input x_278;
input x_279;
input x_280;
input x_281;
input x_282;
input x_283;
input x_284;
input x_285;
input x_286;
input x_287;
input x_288;
input x_289;
input x_290;
input x_291;
input x_292;
input x_293;
input x_294;
input x_295;
input x_296;
input x_297;
input x_298;
input x_299;
input x_300;
input x_301;
input x_302;
input x_303;
input x_304;
input x_305;
input x_306;
input x_307;
input x_308;
input x_309;
input x_310;
input x_311;
input x_312;
input x_313;
input x_314;
input x_315;
input x_316;
input x_317;
input x_318;
input x_319;
input x_320;
input x_321;
input x_322;
input x_323;
input x_324;
input x_325;
input x_326;
input x_327;
input x_328;
input x_329;
input x_330;
input x_331;
input x_332;
input x_333;
input x_334;
input x_335;
input x_336;
input x_337;
input x_338;
input x_339;
input x_340;
input x_341;
input x_342;
input x_343;
input x_344;
input x_345;
input x_346;
input x_347;
input x_348;
input x_349;
input x_350;
input x_351;
input x_352;
input x_353;
input x_354;
input x_355;
input x_356;
input x_357;
input x_358;
input x_359;
input x_360;
input x_361;
input x_362;
input x_363;
input x_364;
input x_365;
input x_366;
input x_367;
input x_368;
input x_369;
input x_370;
input x_371;
input x_372;
input x_373;
input x_374;
input x_375;
input x_376;
input x_377;
input x_378;
input x_379;
input x_380;
input x_381;
input x_382;
input x_383;
input x_384;
input x_385;
input x_386;
input x_387;
input x_388;
input x_389;
input x_390;
input x_391;
input x_392;
input x_393;
input x_394;
input x_395;
input x_396;
input x_397;
input x_398;
input x_399;
input x_400;
input x_401;
input x_402;
input x_403;
input x_404;
input x_405;
input x_406;
input x_407;
input x_408;
input x_409;
input x_410;
input x_411;
input x_412;
input x_413;
input x_414;
input x_415;
input x_416;
input x_417;
input x_418;
input x_419;
input x_420;
input x_421;
input x_422;
input x_423;
input x_424;
input x_425;
input x_426;
input x_427;
input x_428;
input x_429;
input x_430;
input x_431;
input x_432;
input x_433;
input x_434;
input x_435;
input x_436;
input x_437;
input x_438;
input x_439;
input x_440;
input x_441;
input x_442;
input x_443;
input x_444;
input x_445;
input x_446;
input x_447;
input x_448;
input x_449;
input x_450;
input x_451;
input x_452;
input x_453;
input x_454;
input x_455;
input x_456;
input x_457;
input x_458;
input x_459;
input x_460;
input x_461;
input x_462;
input x_463;
input x_464;
input x_465;
input x_466;
input x_467;
input x_468;
input x_469;
input x_470;
input x_471;
input x_472;
input x_473;
input x_474;
input x_475;
input x_476;
input x_477;
input x_478;
input x_479;
input x_480;
input x_481;
input x_482;
input x_483;
input x_484;
input x_485;
input x_486;
input x_487;
input x_488;
input x_489;
input x_490;
input x_491;
input x_492;
input x_493;
input x_494;
input x_495;
input x_496;
input x_497;
input x_498;
input x_499;
input x_500;
input x_501;
input x_502;
input x_503;
input x_504;
input x_505;
input x_506;
input x_507;
input x_508;
input x_509;
input x_510;
input x_511;
input x_512;
input x_513;
input x_514;
input x_515;
input x_516;
input x_517;
input x_518;
input x_519;
input x_520;
input x_521;
input x_522;
input x_523;
input x_524;
input x_525;
input x_526;
input x_527;
input x_528;
input x_529;
input x_530;
input x_531;
input x_532;
input x_533;
input x_534;
input x_535;
input x_536;
input x_537;
input x_538;
input x_539;
input x_540;
input x_541;
input x_542;
input x_543;
input x_544;
input x_545;
input x_546;
input x_547;
input x_548;
input x_549;
input x_550;
input x_551;
input x_552;
input x_553;
input x_554;
input x_555;
input x_556;
input x_557;
input x_558;
input x_559;
input x_560;
input x_561;
input x_562;
input x_563;
input x_564;
input x_565;
input x_566;
input x_567;
input x_568;
input x_569;
input x_570;
input x_571;
input x_572;
input x_573;
input x_574;
input x_575;
input x_576;
input x_577;
input x_578;
input x_579;
input x_580;
input x_581;
input x_582;
input x_583;
input x_584;
input x_585;
input x_586;
input x_587;
input x_588;
input x_589;
input x_590;
input x_591;
input x_592;
input x_593;
input x_594;
input x_595;
input x_596;
input x_597;
input x_598;
input x_599;
input x_600;
input x_601;
input x_602;
input x_603;
input x_604;
input x_605;
input x_606;
input x_607;
input x_608;
input x_609;
input x_610;
input x_611;
input x_612;
input x_613;
input x_614;
input x_615;
input x_616;
input x_617;
input x_618;
input x_619;
input x_620;
input x_621;
input x_622;
input x_623;
input x_624;
input x_625;
input x_626;
input x_627;
input x_628;
input x_629;
input x_630;
input x_631;
input x_632;
input x_633;
input x_634;
input x_635;
input x_636;
input x_637;
input x_638;
input x_639;
input x_640;
input x_641;
input x_642;
input x_643;
input x_644;
input x_645;
input x_646;
input x_647;
input x_648;
input x_649;
input x_650;
input x_651;
input x_652;
input x_653;
input x_654;
input x_655;
input x_656;
input x_657;
input x_658;
input x_659;
input x_660;
input x_661;
input x_662;
input x_663;
input x_664;
input x_665;
input x_666;
input x_667;
input x_668;
input x_669;
input x_670;
input x_671;
input x_672;
input x_673;
input x_674;
input x_675;
input x_676;
input x_677;
input x_678;
input x_679;
input x_680;
input x_681;
input x_682;
input x_683;
input x_684;
input x_685;
input x_686;
input x_687;
input x_688;
input x_689;
input x_690;
input x_691;
input x_692;
input x_693;
input x_694;
input x_695;
input x_696;
input x_697;
input x_698;
input x_699;
input x_700;
input x_701;
input x_702;
input x_703;
input x_704;
input x_705;
input x_706;
input x_707;
input x_708;
input x_709;
input x_710;
input x_711;
input x_712;
input x_713;
input x_714;
input x_715;
input x_716;
input x_717;
input x_718;
input x_719;
input x_720;
input x_721;
input x_722;
input x_723;
input x_724;
input x_725;
input x_726;
input x_727;
input x_728;
input x_729;
input x_730;
input x_731;
input x_732;
input x_733;
input x_734;
input x_735;
input x_736;
input x_737;
input x_738;
input x_739;
input x_740;
input x_741;
input x_742;
input x_743;
input x_744;
input x_745;
input x_746;
input x_747;
input x_748;
input x_749;
input x_750;
input x_751;
input x_752;
input x_753;
input x_754;
input x_755;
input x_756;
input x_757;
input x_758;
input x_759;
input x_760;
input x_761;
input x_762;
input x_763;
input x_764;
input x_765;
input x_766;
input x_767;
input x_768;
input x_769;
input x_770;
input x_771;
input x_772;
input x_773;
input x_774;
input x_775;
input x_776;
input x_777;
input x_778;
input x_779;
input x_780;
input x_781;
input x_782;
input x_783;
input x_784;
input x_785;
input x_786;
input x_787;
input x_788;
input x_789;
input x_790;
input x_791;
input x_792;
input x_793;
input x_794;
input x_795;
input x_796;
input x_797;
input x_798;
input x_799;
input x_800;
input x_801;
input x_802;
input x_803;
input x_804;
input x_805;
input x_806;
input x_807;
input x_808;
input x_809;
input x_810;
input x_811;
input x_812;
input x_813;
input x_814;
input x_815;
input x_816;
input x_817;
input x_818;
input x_819;
input x_820;
input x_821;
input x_822;
input x_823;
input x_824;
input x_825;
input x_826;
input x_827;
input x_828;
input x_829;
input x_830;
input x_831;
input x_832;
input x_833;
input x_834;
input x_835;
input x_836;
input x_837;
input x_838;
input x_839;
input x_840;
input x_841;
input x_842;
input x_843;
input x_844;
input x_845;
input x_846;
input x_847;
input x_848;
input x_849;
input x_850;
input x_851;
input x_852;
input x_853;
input x_854;
input x_855;
input x_856;
input x_857;
input x_858;
input x_859;
input x_860;
input x_861;
input x_862;
input x_863;
input x_864;
input x_865;
input x_866;
input x_867;
input x_868;
input x_869;
input x_870;
input x_871;
input x_872;
input x_873;
input x_874;
input x_875;
input x_876;
input x_877;
input x_878;
input x_879;
input x_880;
input x_881;
input x_882;
input x_883;
input x_884;
input x_885;
input x_886;
input x_887;
input x_888;
input x_889;
input x_890;
input x_891;
input x_892;
input x_893;
input x_894;
input x_895;
input x_896;
input x_897;
input x_898;
input x_899;
input x_900;
input x_901;
input x_902;
input x_903;
input x_904;
input x_905;
input x_906;
input x_907;
input x_908;
input x_909;
input x_910;
input x_911;
input x_912;
input x_913;
input x_914;
input x_915;
input x_916;
input x_917;
input x_918;
input x_919;
input x_920;
input x_921;
input x_922;
input x_923;
input x_924;
input x_925;
input x_926;
input x_927;
input x_928;
input x_929;
input x_930;
input x_931;
input x_932;
input x_933;
input x_934;
input x_935;
input x_936;
input x_937;
input x_938;
input x_939;
input x_940;
input x_941;
input x_942;
input x_943;
input x_944;
input x_945;
input x_946;
input x_947;
input x_948;
input x_949;
input x_950;
input x_951;
input x_952;
input x_953;
input x_954;
input x_955;
input x_956;
input x_957;
input x_958;
input x_959;
input x_960;
input x_961;
input x_962;
input x_963;
input x_964;
input x_965;
input x_966;
input x_967;
input x_968;
input x_969;
input x_970;
input x_971;
input x_972;
input x_973;
input x_974;
input x_975;
input x_976;
input x_977;
input x_978;
input x_979;
input x_980;
input x_981;
input x_982;
input x_983;
input x_984;
input x_985;
input x_986;
input x_987;
input x_988;
input x_989;
input x_990;
input x_991;
input x_992;
input x_993;
input x_994;
input x_995;
input x_996;
input x_997;
input x_998;
input x_999;
input x_1000;
input x_1001;
input x_1002;
input x_1003;
input x_1004;
input x_1005;
input x_1006;
input x_1007;
input x_1008;
input x_1009;
input x_1010;
input x_1011;
input x_1012;
input x_1013;
input x_1014;
input x_1015;
input x_1016;
input x_1017;
input x_1018;
input x_1019;
input x_1020;
input x_1021;
input x_1022;
input x_1023;
input x_1024;
input x_1025;
input x_1026;
input x_1027;
input x_1028;
input x_1029;
input x_1030;
input x_1031;
input x_1032;
input x_1033;
input x_1034;
input x_1035;
input x_1036;
input x_1037;
input x_1038;
input x_1039;
input x_1040;
input x_1041;
input x_1042;
input x_1043;
input x_1044;
input x_1045;
input x_1046;
input x_1047;
input x_1048;
input x_1049;
input x_1050;
input x_1051;
input x_1052;
input x_1053;
input x_1054;
input x_1055;
input x_1056;
input x_1057;
input x_1058;
input x_1059;
input x_1060;
input x_1061;
input x_1062;
input x_1063;
input x_1064;
input x_1065;
input x_1066;
input x_1067;
input x_1068;
input x_1069;
input x_1070;
input x_1071;
input x_1072;
input x_1073;
input x_1074;
input x_1075;
input x_1076;
input x_1077;
input x_1078;
input x_1079;
input x_1080;
input x_1081;
input x_1082;
input x_1083;
input x_1084;
input x_1085;
input x_1086;
input x_1087;
input x_1088;
input x_1089;
input x_1090;
input x_1091;
input x_1092;
input x_1093;
input x_1094;
input x_1095;
input x_1096;
input x_1097;
input x_1098;
input x_1099;
input x_1100;
input x_1101;
input x_1102;
input x_1103;
input x_1104;
input x_1105;
input x_1106;
input x_1107;
input x_1108;
input x_1109;
input x_1110;
input x_1111;
input x_1112;
input x_1113;
input x_1114;
input x_1115;
input x_1116;
input x_1117;
input x_1118;
input x_1119;
input x_1120;
input x_1121;
input x_1122;
input x_1123;
input x_1124;
input x_1125;
input x_1126;
input x_1127;
input x_1128;
input x_1129;
input x_1130;
input x_1131;
input x_1132;
input x_1133;
input x_1134;
input x_1135;
input x_1136;
input x_1137;
input x_1138;
input x_1139;
input x_1140;
input x_1141;
input x_1142;
input x_1143;
input x_1144;
input x_1145;
input x_1146;
input x_1147;
input x_1148;
input x_1149;
input x_1150;
input x_1151;
input x_1152;
input x_1153;
input x_1154;
input x_1155;
input x_1156;
input x_1157;
input x_1158;
input x_1159;
input x_1160;
input x_1161;
input x_1162;
input x_1163;
input x_1164;
input x_1165;
input x_1166;
input x_1167;
input x_1168;
input x_1169;
input x_1170;
input x_1171;
input x_1172;
input x_1173;
input x_1174;
input x_1175;
input x_1176;
input x_1177;
input x_1178;
input x_1179;
input x_1180;
input x_1181;
input x_1182;
input x_1183;
input x_1184;
input x_1185;
input x_1186;
input x_1187;
input x_1188;
input x_1189;
input x_1190;
input x_1191;
input x_1192;
input x_1193;
input x_1194;
input x_1195;
input x_1196;
input x_1197;
input x_1198;
input x_1199;
input x_1200;
input x_1201;
input x_1202;
input x_1203;
input x_1204;
input x_1205;
input x_1206;
input x_1207;
input x_1208;
input x_1209;
input x_1210;
input x_1211;
input x_1212;
input x_1213;
input x_1214;
input x_1215;
input x_1216;
input x_1217;
input x_1218;
input x_1219;
input x_1220;
input x_1221;
input x_1222;
input x_1223;
input x_1224;
input x_1225;
input x_1226;
input x_1227;
input x_1228;
input x_1229;
input x_1230;
input x_1231;
input x_1232;
input x_1233;
input x_1234;
input x_1235;
input x_1236;
input x_1237;
input x_1238;
input x_1239;
input x_1240;
input x_1241;
input x_1242;
input x_1243;
input x_1244;
input x_1245;
input x_1246;
input x_1247;
input x_1248;
input x_1249;
input x_1250;
input x_1251;
input x_1252;
input x_1253;
input x_1254;
input x_1255;
input x_1256;
input x_1257;
input x_1258;
input x_1259;
input x_1260;
input x_1261;
input x_1262;
input x_1263;
input x_1264;
input x_1265;
input x_1266;
input x_1267;
input x_1268;
input x_1269;
input x_1270;
input x_1271;
input x_1272;
input x_1273;
input x_1274;
input x_1275;
input x_1276;
input x_1277;
input x_1278;
input x_1279;
input x_1280;
input x_1281;
input x_1282;
input x_1283;
input x_1284;
input x_1285;
input x_1286;
input x_1287;
input x_1288;
input x_1289;
input x_1290;
input x_1291;
input x_1292;
input x_1293;
input x_1294;
input x_1295;
input x_1296;
input x_1297;
input x_1298;
input x_1299;
input x_1300;
input x_1301;
input x_1302;
input x_1303;
input x_1304;
input x_1305;
input x_1306;
input x_1307;
input x_1308;
input x_1309;
input x_1310;
input x_1311;
input x_1312;
input x_1313;
input x_1314;
input x_1315;
input x_1316;
input x_1317;
input x_1318;
input x_1319;
input x_1320;
input x_1321;
input x_1322;
input x_1323;
input x_1324;
input x_1325;
input x_1326;
input x_1327;
input x_1328;
input x_1329;
input x_1330;
input x_1331;
input x_1332;
input x_1333;
input x_1334;
input x_1335;
input x_1336;
input x_1337;
input x_1338;
input x_1339;
input x_1340;
input x_1341;
input x_1342;
input x_1343;
input x_1344;
input x_1345;
input x_1346;
input x_1347;
input x_1348;
input x_1349;
input x_1350;
input x_1351;
input x_1352;
input x_1353;
input x_1354;
input x_1355;
input x_1356;
input x_1357;
input x_1358;
input x_1359;
input x_1360;
input x_1361;
input x_1362;
input x_1363;
input x_1364;
input x_1365;
input x_1366;
input x_1367;
input x_1368;
input x_1369;
input x_1370;
input x_1371;
input x_1372;
input x_1373;
input x_1374;
input x_1375;
input x_1376;
input x_1377;
input x_1378;
input x_1379;
input x_1380;
input x_1381;
input x_1382;
input x_1383;
input x_1384;
input x_1385;
input x_1386;
input x_1387;
input x_1388;
input x_1389;
input x_1390;
input x_1391;
input x_1392;
input x_1393;
input x_1394;
input x_1395;
input x_1396;
input x_1397;
input x_1398;
input x_1399;
input x_1400;
input x_1401;
input x_1402;
input x_1403;
input x_1404;
input x_1405;
input x_1406;
input x_1407;
input x_1408;
input x_1409;
input x_1410;
input x_1411;
input x_1412;
input x_1413;
input x_1414;
input x_1415;
input x_1416;
input x_1417;
input x_1418;
input x_1419;
input x_1420;
input x_1421;
input x_1422;
input x_1423;
input x_1424;
input x_1425;
input x_1426;
input x_1427;
input x_1428;
input x_1429;
input x_1430;
input x_1431;
input x_1432;
input x_1433;
input x_1434;
input x_1435;
input x_1436;
input x_1437;
input x_1438;
input x_1439;
input x_1440;
input x_1441;
input x_1442;
input x_1443;
input x_1444;
input x_1445;
input x_1446;
input x_1447;
input x_1448;
input x_1449;
input x_1450;
input x_1451;
input x_1452;
input x_1453;
input x_1454;
input x_1455;
input x_1456;
input x_1457;
input x_1458;
input x_1459;
input x_1460;
input x_1461;
input x_1462;
input x_1463;
input x_1464;
input x_1465;
input x_1466;
input x_1467;
input x_1468;
input x_1469;
input x_1470;
input x_1471;
input x_1472;
input x_1473;
input x_1474;
input x_1475;
input x_1476;
input x_1477;
input x_1478;
input x_1479;
input x_1480;
input x_1481;
input x_1482;
input x_1483;
input x_1484;
input x_1485;
input x_1486;
input x_1487;
input x_1488;
input x_1489;
input x_1490;
input x_1491;
input x_1492;
input x_1493;
input x_1494;
input x_1495;
input x_1496;
input x_1497;
input x_1498;
input x_1499;
input x_1500;
input x_1501;
input x_1502;
input x_1503;
input x_1504;
input x_1505;
input x_1506;
input x_1507;
input x_1508;
input x_1509;
input x_1510;
input x_1511;
input x_1512;
input x_1513;
input x_1514;
input x_1515;
input x_1516;
input x_1517;
input x_1518;
input x_1519;
input x_1520;
input x_1521;
input x_1522;
input x_1523;
input x_1524;
input x_1525;
input x_1526;
input x_1527;
input x_1528;
input x_1529;
input x_1530;
input x_1531;
input x_1532;
input x_1533;
input x_1534;
input x_1535;
input x_1536;
input x_1537;
input x_1538;
input x_1539;
input x_1540;
input x_1541;
input x_1542;
input x_1543;
input x_1544;
input x_1545;
input x_1546;
input x_1547;
input x_1548;
input x_1549;
input x_1550;
input x_1551;
input x_1552;
input x_1553;
input x_1554;
input x_1555;
input x_1556;
input x_1557;
input x_1558;
input x_1559;
input x_1560;
input x_1561;
input x_1562;
input x_1563;
input x_1564;
input x_1565;
input x_1566;
input x_1567;
input x_1568;
input x_1569;
input x_1570;
input x_1571;
input x_1572;
input x_1573;
input x_1574;
input x_1575;
input x_1576;
input x_1577;
input x_1578;
input x_1579;
input x_1580;
input x_1581;
input x_1582;
input x_1583;
input x_1584;
input x_1585;
input x_1586;
input x_1587;
input x_1588;
input x_1589;
input x_1590;
input x_1591;
input x_1592;
input x_1593;
input x_1594;
input x_1595;
input x_1596;
input x_1597;
input x_1598;
input x_1599;
input x_1600;
input x_1601;
input x_1602;
input x_1603;
input x_1604;
input x_1605;
input x_1606;
input x_1607;
input x_1608;
input x_1609;
input x_1610;
input x_1611;
input x_1612;
input x_1613;
input x_1614;
input x_1615;
input x_1616;
input x_1617;
input x_1618;
input x_1619;
input x_1620;
input x_1621;
input x_1622;
input x_1623;
input x_1624;
input x_1625;
input x_1626;
input x_1627;
input x_1628;
input x_1629;
input x_1630;
input x_1631;
input x_1632;
input x_1633;
input x_1634;
input x_1635;
input x_1636;
input x_1637;
input x_1638;
input x_1639;
input x_1640;
input x_1641;
input x_1642;
input x_1643;
input x_1644;
input x_1645;
input x_1646;
input x_1647;
input x_1648;
input x_1649;
input x_1650;
input x_1651;
input x_1652;
input x_1653;
input x_1654;
input x_1655;
input x_1656;
input x_1657;
input x_1658;
input x_1659;
input x_1660;
input x_1661;
input x_1662;
input x_1663;
input x_1664;
input x_1665;
input x_1666;
input x_1667;
input x_1668;
input x_1669;
input x_1670;
input x_1671;
input x_1672;
input x_1673;
input x_1674;
input x_1675;
input x_1676;
input x_1677;
input x_1678;
input x_1679;
input x_1680;
input x_1681;
input x_1682;
input x_1683;
input x_1684;
input x_1685;
input x_1686;
input x_1687;
input x_1688;
input x_1689;
input x_1690;
input x_1691;
input x_1692;
input x_1693;
input x_1694;
input x_1695;
input x_1696;
input x_1697;
input x_1698;
input x_1699;
input x_1700;
input x_1701;
input x_1702;
input x_1703;
input x_1704;
input x_1705;
input x_1706;
input x_1707;
input x_1708;
input x_1709;
input x_1710;
input x_1711;
input x_1712;
input x_1713;
input x_1714;
input x_1715;
input x_1716;
input x_1717;
input x_1718;
input x_1719;
input x_1720;
input x_1721;
input x_1722;
input x_1723;
input x_1724;
input x_1725;
input x_1726;
input x_1727;
input x_1728;
input x_1729;
input x_1730;
input x_1731;
input x_1732;
input x_1733;
input x_1734;
input x_1735;
input x_1736;
input x_1737;
input x_1738;
input x_1739;
input x_1740;
input x_1741;
input x_1742;
input x_1743;
input x_1744;
input x_1745;
input x_1746;
input x_1747;
input x_1748;
input x_1749;
input x_1750;
input x_1751;
input x_1752;
input x_1753;
input x_1754;
input x_1755;
input x_1756;
input x_1757;
input x_1758;
input x_1759;
input x_1760;
input x_1761;
input x_1762;
input x_1763;
input x_1764;
input x_1765;
input x_1766;
input x_1767;
input x_1768;
input x_1769;
input x_1770;
input x_1771;
input x_1772;
input x_1773;
input x_1774;
input x_1775;
input x_1776;
input x_1777;
input x_1778;
input x_1779;
input x_1780;
input x_1781;
input x_1782;
input x_1783;
input x_1784;
input x_1785;
input x_1786;
input x_1787;
input x_1788;
input x_1789;
input x_1790;
input x_1791;
input x_1792;
input x_1793;
input x_1794;
input x_1795;
input x_1796;
input x_1797;
input x_1798;
input x_1799;
input x_1800;
input x_1801;
input x_1802;
input x_1803;
input x_1804;
input x_1805;
input x_1806;
input x_1807;
input x_1808;
input x_1809;
input x_1810;
input x_1811;
input x_1812;
input x_1813;
input x_1814;
input x_1815;
input x_1816;
input x_1817;
input x_1818;
input x_1819;
input x_1820;
input x_1821;
input x_1822;
input x_1823;
input x_1824;
input x_1825;
input x_1826;
input x_1827;
input x_1828;
input x_1829;
input x_1830;
input x_1831;
input x_1832;
input x_1833;
input x_1834;
input x_1835;
input x_1836;
input x_1837;
input x_1838;
input x_1839;
input x_1840;
input x_1841;
input x_1842;
input x_1843;
input x_1844;
input x_1845;
input x_1846;
input x_1847;
input x_1848;
input x_1849;
input x_1850;
input x_1851;
input x_1852;
input x_1853;
input x_1854;
input x_1855;
input x_1856;
input x_1857;
input x_1858;
input x_1859;
input x_1860;
input x_1861;
input x_1862;
input x_1863;
input x_1864;
input x_1865;
input x_1866;
input x_1867;
input x_1868;
input x_1869;
input x_1870;
input x_1871;
input x_1872;
input x_1873;
input x_1874;
input x_1875;
input x_1876;
input x_1877;
input x_1878;
input x_1879;
input x_1880;
input x_1881;
input x_1882;
input x_1883;
input x_1884;
input x_1885;
input x_1886;
input x_1887;
input x_1888;
input x_1889;
input x_1890;
input x_1891;
input x_1892;
input x_1893;
input x_1894;
input x_1895;
input x_1896;
input x_1897;
input x_1898;
input x_1899;
input x_1900;
input x_1901;
input x_1902;
input x_1903;
input x_1904;
input x_1905;
input x_1906;
input x_1907;
input x_1908;
input x_1909;
input x_1910;
input x_1911;
input x_1912;
input x_1913;
input x_1914;
input x_1915;
input x_1916;
input x_1917;
input x_1918;
input x_1919;
input x_1920;
input x_1921;
input x_1922;
input x_1923;
input x_1924;
input x_1925;
input x_1926;
input x_1927;
input x_1928;
input x_1929;
input x_1930;
input x_1931;
input x_1932;
input x_1933;
input x_1934;
input x_1935;
input x_1936;
input x_1937;
input x_1938;
input x_1939;
input x_1940;
input x_1941;
input x_1942;
input x_1943;
input x_1944;
input x_1945;
input x_1946;
input x_1947;
input x_1948;
input x_1949;
input x_1950;
input x_1951;
input x_1952;
input x_1953;
input x_1954;
input x_1955;
input x_1956;
input x_1957;
input x_1958;
input x_1959;
input x_1960;
input x_1961;
input x_1962;
input x_1963;
input x_1964;
input x_1965;
input x_1966;
input x_1967;
input x_1968;
input x_1969;
input x_1970;
input x_1971;
input x_1972;
input x_1973;
input x_1974;
input x_1975;
input x_1976;
input x_1977;
input x_1978;
input x_1979;
input x_1980;
input x_1981;
input x_1982;
input x_1983;
input x_1984;
input x_1985;
input x_1986;
input x_1987;
input x_1988;
input x_1989;
input x_1990;
input x_1991;
input x_1992;
input x_1993;
input x_1994;
input x_1995;
input x_1996;
input x_1997;
input x_1998;
input x_1999;
input x_2000;
input x_2001;
input x_2002;
input x_2003;
input x_2004;
input x_2005;
input x_2006;
input x_2007;
input x_2008;
input x_2009;
input x_2010;
input x_2011;
input x_2012;
input x_2013;
input x_2014;
input x_2015;
input x_2016;
input x_2017;
input x_2018;
input x_2019;
input x_2020;
input x_2021;
input x_2022;
input x_2023;
input x_2024;
input x_2025;
input x_2026;
input x_2027;
input x_2028;
input x_2029;
input x_2030;
input x_2031;
input x_2032;
input x_2033;
input x_2034;
input x_2035;
input x_2036;
input x_2037;
input x_2038;
input x_2039;
input x_2040;
input x_2041;
input x_2042;
input x_2043;
input x_2044;
input x_2045;
input x_2046;
input x_2047;
input x_2048;
input x_2049;
input x_2050;
input x_2051;
input x_2052;
input x_2053;
input x_2054;
input x_2055;
input x_2056;
input x_2057;
input x_2058;
input x_2059;
input x_2060;
input x_2061;
input x_2062;
input x_2063;
input x_2064;
input x_2065;
input x_2066;
input x_2067;
input x_2068;
input x_2069;
input x_2070;
input x_2071;
input x_2072;
input x_2073;
input x_2074;
input x_2075;
input x_2076;
input x_2077;
input x_2078;
input x_2079;
input x_2080;
input x_2081;
input x_2082;
input x_2083;
input x_2084;
input x_2085;
input x_2086;
input x_2087;
input x_2088;
input x_2089;
input x_2090;
input x_2091;
input x_2092;
input x_2093;
input x_2094;
input x_2095;
input x_2096;
input x_2097;
input x_2098;
input x_2099;
input x_2100;
input x_2101;
input x_2102;
input x_2103;
input x_2104;
input x_2105;
input x_2106;
input x_2107;
input x_2108;
input x_2109;
input x_2110;
input x_2111;
input x_2112;
input x_2113;
input x_2114;
input x_2115;
input x_2116;
input x_2117;
input x_2118;
input x_2119;
input x_2120;
input x_2121;
input x_2122;
input x_2123;
input x_2124;
input x_2125;
input x_2126;
input x_2127;
input x_2128;
input x_2129;
input x_2130;
input x_2131;
input x_2132;
input x_2133;
input x_2134;
input x_2135;
input x_2136;
input x_2137;
input x_2138;
input x_2139;
input x_2140;
input x_2141;
input x_2142;
input x_2143;
input x_2144;
input x_2145;
input x_2146;
input x_2147;
input x_2148;
input x_2149;
input x_2150;
input x_2151;
input x_2152;
input x_2153;
input x_2154;
input x_2155;
input x_2156;
input x_2157;
input x_2158;
input x_2159;
input x_2160;
input x_2161;
input x_2162;
input x_2163;
input x_2164;
input x_2165;
input x_2166;
input x_2167;
input x_2168;
input x_2169;
input x_2170;
input x_2171;
input x_2172;
input x_2173;
input x_2174;
input x_2175;
input x_2176;
input x_2177;
input x_2178;
input x_2179;
input x_2180;
input x_2181;
input x_2182;
input x_2183;
input x_2184;
input x_2185;
input x_2186;
input x_2187;
input x_2188;
input x_2189;
input x_2190;
input x_2191;
input x_2192;
input x_2193;
input x_2194;
input x_2195;
input x_2196;
input x_2197;
input x_2198;
input x_2199;
input x_2200;
input x_2201;
input x_2202;
input x_2203;
input x_2204;
input x_2205;
input x_2206;
input x_2207;
input x_2208;
input x_2209;
input x_2210;
input x_2211;
input x_2212;
input x_2213;
input x_2214;
input x_2215;
input x_2216;
input x_2217;
input x_2218;
input x_2219;
input x_2220;
output o_1;
wire n_1;
wire n_2;
wire n_3;
wire n_4;
wire n_5;
wire n_6;
wire n_7;
wire n_8;
wire n_9;
wire n_10;
wire n_11;
wire n_12;
wire n_13;
wire n_14;
wire n_15;
wire n_16;
wire n_17;
wire n_18;
wire n_19;
wire n_20;
wire n_21;
wire n_22;
wire n_23;
wire n_24;
wire n_25;
wire n_26;
wire n_27;
wire n_28;
wire n_29;
wire n_30;
wire n_31;
wire n_32;
wire n_33;
wire n_34;
wire n_35;
wire n_36;
wire n_37;
wire n_38;
wire n_39;
wire n_40;
wire n_41;
wire n_42;
wire n_43;
wire n_44;
wire n_45;
wire n_46;
wire n_47;
wire n_48;
wire n_49;
wire n_50;
wire n_51;
wire n_52;
wire n_53;
wire n_54;
wire n_55;
wire n_56;
wire n_57;
wire n_58;
wire n_59;
wire n_60;
wire n_61;
wire n_62;
wire n_63;
wire n_64;
wire n_65;
wire n_66;
wire n_67;
wire n_68;
wire n_69;
wire n_70;
wire n_71;
wire n_72;
wire n_73;
wire n_74;
wire n_75;
wire n_76;
wire n_77;
wire n_78;
wire n_79;
wire n_80;
wire n_81;
wire n_82;
wire n_83;
wire n_84;
wire n_85;
wire n_86;
wire n_87;
wire n_88;
wire n_89;
wire n_90;
wire n_91;
wire n_92;
wire n_93;
wire n_94;
wire n_95;
wire n_96;
wire n_97;
wire n_98;
wire n_99;
wire n_100;
wire n_101;
wire n_102;
wire n_103;
wire n_104;
wire n_105;
wire n_106;
wire n_107;
wire n_108;
wire n_109;
wire n_110;
wire n_111;
wire n_112;
wire n_113;
wire n_114;
wire n_115;
wire n_116;
wire n_117;
wire n_118;
wire n_119;
wire n_120;
wire n_121;
wire n_122;
wire n_123;
wire n_124;
wire n_125;
wire n_126;
wire n_127;
wire n_128;
wire n_129;
wire n_130;
wire n_131;
wire n_132;
wire n_133;
wire n_134;
wire n_135;
wire n_136;
wire n_137;
wire n_138;
wire n_139;
wire n_140;
wire n_141;
wire n_142;
wire n_143;
wire n_144;
wire n_145;
wire n_146;
wire n_147;
wire n_148;
wire n_149;
wire n_150;
wire n_151;
wire n_152;
wire n_153;
wire n_154;
wire n_155;
wire n_156;
wire n_157;
wire n_158;
wire n_159;
wire n_160;
wire n_161;
wire n_162;
wire n_163;
wire n_164;
wire n_165;
wire n_166;
wire n_167;
wire n_168;
wire n_169;
wire n_170;
wire n_171;
wire n_172;
wire n_173;
wire n_174;
wire n_175;
wire n_176;
wire n_177;
wire n_178;
wire n_179;
wire n_180;
wire n_181;
wire n_182;
wire n_183;
wire n_184;
wire n_185;
wire n_186;
wire n_187;
wire n_188;
wire n_189;
wire n_190;
wire n_191;
wire n_192;
wire n_193;
wire n_194;
wire n_195;
wire n_196;
wire n_197;
wire n_198;
wire n_199;
wire n_200;
wire n_201;
wire n_202;
wire n_203;
wire n_204;
wire n_205;
wire n_206;
wire n_207;
wire n_208;
wire n_209;
wire n_210;
wire n_211;
wire n_212;
wire n_213;
wire n_214;
wire n_215;
wire n_216;
wire n_217;
wire n_218;
wire n_219;
wire n_220;
wire n_221;
wire n_222;
wire n_223;
wire n_224;
wire n_225;
wire n_226;
wire n_227;
wire n_228;
wire n_229;
wire n_230;
wire n_231;
wire n_232;
wire n_233;
wire n_234;
wire n_235;
wire n_236;
wire n_237;
wire n_238;
wire n_239;
wire n_240;
wire n_241;
wire n_242;
wire n_243;
wire n_244;
wire n_245;
wire n_246;
wire n_247;
wire n_248;
wire n_249;
wire n_250;
wire n_251;
wire n_252;
wire n_253;
wire n_254;
wire n_255;
wire n_256;
wire n_257;
wire n_258;
wire n_259;
wire n_260;
wire n_261;
wire n_262;
wire n_263;
wire n_264;
wire n_265;
wire n_266;
wire n_267;
wire n_268;
wire n_269;
wire n_270;
wire n_271;
wire n_272;
wire n_273;
wire n_274;
wire n_275;
wire n_276;
wire n_277;
wire n_278;
wire n_279;
wire n_280;
wire n_281;
wire n_282;
wire n_283;
wire n_284;
wire n_285;
wire n_286;
wire n_287;
wire n_288;
wire n_289;
wire n_290;
wire n_291;
wire n_292;
wire n_293;
wire n_294;
wire n_295;
wire n_296;
wire n_297;
wire n_298;
wire n_299;
wire n_300;
wire n_301;
wire n_302;
wire n_303;
wire n_304;
wire n_305;
wire n_306;
wire n_307;
wire n_308;
wire n_309;
wire n_310;
wire n_311;
wire n_312;
wire n_313;
wire n_314;
wire n_315;
wire n_316;
wire n_317;
wire n_318;
wire n_319;
wire n_320;
wire n_321;
wire n_322;
wire n_323;
wire n_324;
wire n_325;
wire n_326;
wire n_327;
wire n_328;
wire n_329;
wire n_330;
wire n_331;
wire n_332;
wire n_333;
wire n_334;
wire n_335;
wire n_336;
wire n_337;
wire n_338;
wire n_339;
wire n_340;
wire n_341;
wire n_342;
wire n_343;
wire n_344;
wire n_345;
wire n_346;
wire n_347;
wire n_348;
wire n_349;
wire n_350;
wire n_351;
wire n_352;
wire n_353;
wire n_354;
wire n_355;
wire n_356;
wire n_357;
wire n_358;
wire n_359;
wire n_360;
wire n_361;
wire n_362;
wire n_363;
wire n_364;
wire n_365;
wire n_366;
wire n_367;
wire n_368;
wire n_369;
wire n_370;
wire n_371;
wire n_372;
wire n_373;
wire n_374;
wire n_375;
wire n_376;
wire n_377;
wire n_378;
wire n_379;
wire n_380;
wire n_381;
wire n_382;
wire n_383;
wire n_384;
wire n_385;
wire n_386;
wire n_387;
wire n_388;
wire n_389;
wire n_390;
wire n_391;
wire n_392;
wire n_393;
wire n_394;
wire n_395;
wire n_396;
wire n_397;
wire n_398;
wire n_399;
wire n_400;
wire n_401;
wire n_402;
wire n_403;
wire n_404;
wire n_405;
wire n_406;
wire n_407;
wire n_408;
wire n_409;
wire n_410;
wire n_411;
wire n_412;
wire n_413;
wire n_414;
wire n_415;
wire n_416;
wire n_417;
wire n_418;
wire n_419;
wire n_420;
wire n_421;
wire n_422;
wire n_423;
wire n_424;
wire n_425;
wire n_426;
wire n_427;
wire n_428;
wire n_429;
wire n_430;
wire n_431;
wire n_432;
wire n_433;
wire n_434;
wire n_435;
wire n_436;
wire n_437;
wire n_438;
wire n_439;
wire n_440;
wire n_441;
wire n_442;
wire n_443;
wire n_444;
wire n_445;
wire n_446;
wire n_447;
wire n_448;
wire n_449;
wire n_450;
wire n_451;
wire n_452;
wire n_453;
wire n_454;
wire n_455;
wire n_456;
wire n_457;
wire n_458;
wire n_459;
wire n_460;
wire n_461;
wire n_462;
wire n_463;
wire n_464;
wire n_465;
wire n_466;
wire n_467;
wire n_468;
wire n_469;
wire n_470;
wire n_471;
wire n_472;
wire n_473;
wire n_474;
wire n_475;
wire n_476;
wire n_477;
wire n_478;
wire n_479;
wire n_480;
wire n_481;
wire n_482;
wire n_483;
wire n_484;
wire n_485;
wire n_486;
wire n_487;
wire n_488;
wire n_489;
wire n_490;
wire n_491;
wire n_492;
wire n_493;
wire n_494;
wire n_495;
wire n_496;
wire n_497;
wire n_498;
wire n_499;
wire n_500;
wire n_501;
wire n_502;
wire n_503;
wire n_504;
wire n_505;
wire n_506;
wire n_507;
wire n_508;
wire n_509;
wire n_510;
wire n_511;
wire n_512;
wire n_513;
wire n_514;
wire n_515;
wire n_516;
wire n_517;
wire n_518;
wire n_519;
wire n_520;
wire n_521;
wire n_522;
wire n_523;
wire n_524;
wire n_525;
wire n_526;
wire n_527;
wire n_528;
wire n_529;
wire n_530;
wire n_531;
wire n_532;
wire n_533;
wire n_534;
wire n_535;
wire n_536;
wire n_537;
wire n_538;
wire n_539;
wire n_540;
wire n_541;
wire n_542;
wire n_543;
wire n_544;
wire n_545;
wire n_546;
wire n_547;
wire n_548;
wire n_549;
wire n_550;
wire n_551;
wire n_552;
wire n_553;
wire n_554;
wire n_555;
wire n_556;
wire n_557;
wire n_558;
wire n_559;
wire n_560;
wire n_561;
wire n_562;
wire n_563;
wire n_564;
wire n_565;
wire n_566;
wire n_567;
wire n_568;
wire n_569;
wire n_570;
wire n_571;
wire n_572;
wire n_573;
wire n_574;
wire n_575;
wire n_576;
wire n_577;
wire n_578;
wire n_579;
wire n_580;
wire n_581;
wire n_582;
wire n_583;
wire n_584;
wire n_585;
wire n_586;
wire n_587;
wire n_588;
wire n_589;
wire n_590;
wire n_591;
wire n_592;
wire n_593;
wire n_594;
wire n_595;
wire n_596;
wire n_597;
wire n_598;
wire n_599;
wire n_600;
wire n_601;
wire n_602;
wire n_603;
wire n_604;
wire n_605;
wire n_606;
wire n_607;
wire n_608;
wire n_609;
wire n_610;
wire n_611;
wire n_612;
wire n_613;
wire n_614;
wire n_615;
wire n_616;
wire n_617;
wire n_618;
wire n_619;
wire n_620;
wire n_621;
wire n_622;
wire n_623;
wire n_624;
wire n_625;
wire n_626;
wire n_627;
wire n_628;
wire n_629;
wire n_630;
wire n_631;
wire n_632;
wire n_633;
wire n_634;
wire n_635;
wire n_636;
wire n_637;
wire n_638;
wire n_639;
wire n_640;
wire n_641;
wire n_642;
wire n_643;
wire n_644;
wire n_645;
wire n_646;
wire n_647;
wire n_648;
wire n_649;
wire n_650;
wire n_651;
wire n_652;
wire n_653;
wire n_654;
wire n_655;
wire n_656;
wire n_657;
wire n_658;
wire n_659;
wire n_660;
wire n_661;
wire n_662;
wire n_663;
wire n_664;
wire n_665;
wire n_666;
wire n_667;
wire n_668;
wire n_669;
wire n_670;
wire n_671;
wire n_672;
wire n_673;
wire n_674;
wire n_675;
wire n_676;
wire n_677;
wire n_678;
wire n_679;
wire n_680;
wire n_681;
wire n_682;
wire n_683;
wire n_684;
wire n_685;
wire n_686;
wire n_687;
wire n_688;
wire n_689;
wire n_690;
wire n_691;
wire n_692;
wire n_693;
wire n_694;
wire n_695;
wire n_696;
wire n_697;
wire n_698;
wire n_699;
wire n_700;
wire n_701;
wire n_702;
wire n_703;
wire n_704;
wire n_705;
wire n_706;
wire n_707;
wire n_708;
wire n_709;
wire n_710;
wire n_711;
wire n_712;
wire n_713;
wire n_714;
wire n_715;
wire n_716;
wire n_717;
wire n_718;
wire n_719;
wire n_720;
wire n_721;
wire n_722;
wire n_723;
wire n_724;
wire n_725;
wire n_726;
wire n_727;
wire n_728;
wire n_729;
wire n_730;
wire n_731;
wire n_732;
wire n_733;
wire n_734;
wire n_735;
wire n_736;
wire n_737;
wire n_738;
wire n_739;
wire n_740;
wire n_741;
wire n_742;
wire n_743;
wire n_744;
wire n_745;
wire n_746;
wire n_747;
wire n_748;
wire n_749;
wire n_750;
wire n_751;
wire n_752;
wire n_753;
wire n_754;
wire n_755;
wire n_756;
wire n_757;
wire n_758;
wire n_759;
wire n_760;
wire n_761;
wire n_762;
wire n_763;
wire n_764;
wire n_765;
wire n_766;
wire n_767;
wire n_768;
wire n_769;
wire n_770;
wire n_771;
wire n_772;
wire n_773;
wire n_774;
wire n_775;
wire n_776;
wire n_777;
wire n_778;
wire n_779;
wire n_780;
wire n_781;
wire n_782;
wire n_783;
wire n_784;
wire n_785;
wire n_786;
wire n_787;
wire n_788;
wire n_789;
wire n_790;
wire n_791;
wire n_792;
wire n_793;
wire n_794;
wire n_795;
wire n_796;
wire n_797;
wire n_798;
wire n_799;
wire n_800;
wire n_801;
wire n_802;
wire n_803;
wire n_804;
wire n_805;
wire n_806;
wire n_807;
wire n_808;
wire n_809;
wire n_810;
wire n_811;
wire n_812;
wire n_813;
wire n_814;
wire n_815;
wire n_816;
wire n_817;
wire n_818;
wire n_819;
wire n_820;
wire n_821;
wire n_822;
wire n_823;
wire n_824;
wire n_825;
wire n_826;
wire n_827;
wire n_828;
wire n_829;
wire n_830;
wire n_831;
wire n_832;
wire n_833;
wire n_834;
wire n_835;
wire n_836;
wire n_837;
wire n_838;
wire n_839;
wire n_840;
wire n_841;
wire n_842;
wire n_843;
wire n_844;
wire n_845;
wire n_846;
wire n_847;
wire n_848;
wire n_849;
wire n_850;
wire n_851;
wire n_852;
wire n_853;
wire n_854;
wire n_855;
wire n_856;
wire n_857;
wire n_858;
wire n_859;
wire n_860;
wire n_861;
wire n_862;
wire n_863;
wire n_864;
wire n_865;
wire n_866;
wire n_867;
wire n_868;
wire n_869;
wire n_870;
wire n_871;
wire n_872;
wire n_873;
wire n_874;
wire n_875;
wire n_876;
wire n_877;
wire n_878;
wire n_879;
wire n_880;
wire n_881;
wire n_882;
wire n_883;
wire n_884;
wire n_885;
wire n_886;
wire n_887;
wire n_888;
wire n_889;
wire n_890;
wire n_891;
wire n_892;
wire n_893;
wire n_894;
wire n_895;
wire n_896;
wire n_897;
wire n_898;
wire n_899;
wire n_900;
wire n_901;
wire n_902;
wire n_903;
wire n_904;
wire n_905;
wire n_906;
wire n_907;
wire n_908;
wire n_909;
wire n_910;
wire n_911;
wire n_912;
wire n_913;
wire n_914;
wire n_915;
wire n_916;
wire n_917;
wire n_918;
wire n_919;
wire n_920;
wire n_921;
wire n_922;
wire n_923;
wire n_924;
wire n_925;
wire n_926;
wire n_927;
wire n_928;
wire n_929;
wire n_930;
wire n_931;
wire n_932;
wire n_933;
wire n_934;
wire n_935;
wire n_936;
wire n_937;
wire n_938;
wire n_939;
wire n_940;
wire n_941;
wire n_942;
wire n_943;
wire n_944;
wire n_945;
wire n_946;
wire n_947;
wire n_948;
wire n_949;
wire n_950;
wire n_951;
wire n_952;
wire n_953;
wire n_954;
wire n_955;
wire n_956;
wire n_957;
wire n_958;
wire n_959;
wire n_960;
wire n_961;
wire n_962;
wire n_963;
wire n_964;
wire n_965;
wire n_966;
wire n_967;
wire n_968;
wire n_969;
wire n_970;
wire n_971;
wire n_972;
wire n_973;
wire n_974;
wire n_975;
wire n_976;
wire n_977;
wire n_978;
wire n_979;
wire n_980;
wire n_981;
wire n_982;
wire n_983;
wire n_984;
wire n_985;
wire n_986;
wire n_987;
wire n_988;
wire n_989;
wire n_990;
wire n_991;
wire n_992;
wire n_993;
wire n_994;
wire n_995;
wire n_996;
wire n_997;
wire n_998;
wire n_999;
wire n_1000;
wire n_1001;
wire n_1002;
wire n_1003;
wire n_1004;
wire n_1005;
wire n_1006;
wire n_1007;
wire n_1008;
wire n_1009;
wire n_1010;
wire n_1011;
wire n_1012;
wire n_1013;
wire n_1014;
wire n_1015;
wire n_1016;
wire n_1017;
wire n_1018;
wire n_1019;
wire n_1020;
wire n_1021;
wire n_1022;
wire n_1023;
wire n_1024;
wire n_1025;
wire n_1026;
wire n_1027;
wire n_1028;
wire n_1029;
wire n_1030;
wire n_1031;
wire n_1032;
wire n_1033;
wire n_1034;
wire n_1035;
wire n_1036;
wire n_1037;
wire n_1038;
wire n_1039;
wire n_1040;
wire n_1041;
wire n_1042;
wire n_1043;
wire n_1044;
wire n_1045;
wire n_1046;
wire n_1047;
wire n_1048;
wire n_1049;
wire n_1050;
wire n_1051;
wire n_1052;
wire n_1053;
wire n_1054;
wire n_1055;
wire n_1056;
wire n_1057;
wire n_1058;
wire n_1059;
wire n_1060;
wire n_1061;
wire n_1062;
wire n_1063;
wire n_1064;
wire n_1065;
wire n_1066;
wire n_1067;
wire n_1068;
wire n_1069;
wire n_1070;
wire n_1071;
wire n_1072;
wire n_1073;
wire n_1074;
wire n_1075;
wire n_1076;
wire n_1077;
wire n_1078;
wire n_1079;
wire n_1080;
wire n_1081;
wire n_1082;
wire n_1083;
wire n_1084;
wire n_1085;
wire n_1086;
wire n_1087;
wire n_1088;
wire n_1089;
wire n_1090;
wire n_1091;
wire n_1092;
wire n_1093;
wire n_1094;
wire n_1095;
wire n_1096;
wire n_1097;
wire n_1098;
wire n_1099;
wire n_1100;
wire n_1101;
wire n_1102;
wire n_1103;
wire n_1104;
wire n_1105;
wire n_1106;
wire n_1107;
wire n_1108;
wire n_1109;
wire n_1110;
wire n_1111;
wire n_1112;
wire n_1113;
wire n_1114;
wire n_1115;
wire n_1116;
wire n_1117;
wire n_1118;
wire n_1119;
wire n_1120;
wire n_1121;
wire n_1122;
wire n_1123;
wire n_1124;
wire n_1125;
wire n_1126;
wire n_1127;
wire n_1128;
wire n_1129;
wire n_1130;
wire n_1131;
wire n_1132;
wire n_1133;
wire n_1134;
wire n_1135;
wire n_1136;
wire n_1137;
wire n_1138;
wire n_1139;
wire n_1140;
wire n_1141;
wire n_1142;
wire n_1143;
wire n_1144;
wire n_1145;
wire n_1146;
wire n_1147;
wire n_1148;
wire n_1149;
wire n_1150;
wire n_1151;
wire n_1152;
wire n_1153;
wire n_1154;
wire n_1155;
wire n_1156;
wire n_1157;
wire n_1158;
wire n_1159;
wire n_1160;
wire n_1161;
wire n_1162;
wire n_1163;
wire n_1164;
wire n_1165;
wire n_1166;
wire n_1167;
wire n_1168;
wire n_1169;
wire n_1170;
wire n_1171;
wire n_1172;
wire n_1173;
wire n_1174;
wire n_1175;
wire n_1176;
wire n_1177;
wire n_1178;
wire n_1179;
wire n_1180;
wire n_1181;
wire n_1182;
wire n_1183;
wire n_1184;
wire n_1185;
wire n_1186;
wire n_1187;
wire n_1188;
wire n_1189;
wire n_1190;
wire n_1191;
wire n_1192;
wire n_1193;
wire n_1194;
wire n_1195;
wire n_1196;
wire n_1197;
wire n_1198;
wire n_1199;
wire n_1200;
wire n_1201;
wire n_1202;
wire n_1203;
wire n_1204;
wire n_1205;
wire n_1206;
wire n_1207;
wire n_1208;
wire n_1209;
wire n_1210;
wire n_1211;
wire n_1212;
wire n_1213;
wire n_1214;
wire n_1215;
wire n_1216;
wire n_1217;
wire n_1218;
wire n_1219;
wire n_1220;
wire n_1221;
wire n_1222;
wire n_1223;
wire n_1224;
wire n_1225;
wire n_1226;
wire n_1227;
wire n_1228;
wire n_1229;
wire n_1230;
wire n_1231;
wire n_1232;
wire n_1233;
wire n_1234;
wire n_1235;
wire n_1236;
wire n_1237;
wire n_1238;
wire n_1239;
wire n_1240;
wire n_1241;
wire n_1242;
wire n_1243;
wire n_1244;
wire n_1245;
wire n_1246;
wire n_1247;
wire n_1248;
wire n_1249;
wire n_1250;
wire n_1251;
wire n_1252;
wire n_1253;
wire n_1254;
wire n_1255;
wire n_1256;
wire n_1257;
wire n_1258;
wire n_1259;
wire n_1260;
wire n_1261;
wire n_1262;
wire n_1263;
wire n_1264;
wire n_1265;
wire n_1266;
wire n_1267;
wire n_1268;
wire n_1269;
wire n_1270;
wire n_1271;
wire n_1272;
wire n_1273;
wire n_1274;
wire n_1275;
wire n_1276;
wire n_1277;
wire n_1278;
wire n_1279;
wire n_1280;
wire n_1281;
wire n_1282;
wire n_1283;
wire n_1284;
wire n_1285;
wire n_1286;
wire n_1287;
wire n_1288;
wire n_1289;
wire n_1290;
wire n_1291;
wire n_1292;
wire n_1293;
wire n_1294;
wire n_1295;
wire n_1296;
wire n_1297;
wire n_1298;
wire n_1299;
wire n_1300;
wire n_1301;
wire n_1302;
wire n_1303;
wire n_1304;
wire n_1305;
wire n_1306;
wire n_1307;
wire n_1308;
wire n_1309;
wire n_1310;
wire n_1311;
wire n_1312;
wire n_1313;
wire n_1314;
wire n_1315;
wire n_1316;
wire n_1317;
wire n_1318;
wire n_1319;
wire n_1320;
wire n_1321;
wire n_1322;
wire n_1323;
wire n_1324;
wire n_1325;
wire n_1326;
wire n_1327;
wire n_1328;
wire n_1329;
wire n_1330;
wire n_1331;
wire n_1332;
wire n_1333;
wire n_1334;
wire n_1335;
wire n_1336;
wire n_1337;
wire n_1338;
wire n_1339;
wire n_1340;
wire n_1341;
wire n_1342;
wire n_1343;
wire n_1344;
wire n_1345;
wire n_1346;
wire n_1347;
wire n_1348;
wire n_1349;
wire n_1350;
wire n_1351;
wire n_1352;
wire n_1353;
wire n_1354;
wire n_1355;
wire n_1356;
wire n_1357;
wire n_1358;
wire n_1359;
wire n_1360;
wire n_1361;
wire n_1362;
wire n_1363;
wire n_1364;
wire n_1365;
wire n_1366;
wire n_1367;
wire n_1368;
wire n_1369;
wire n_1370;
wire n_1371;
wire n_1372;
wire n_1373;
wire n_1374;
wire n_1375;
wire n_1376;
wire n_1377;
wire n_1378;
wire n_1379;
wire n_1380;
wire n_1381;
wire n_1382;
wire n_1383;
wire n_1384;
wire n_1385;
wire n_1386;
wire n_1387;
wire n_1388;
wire n_1389;
wire n_1390;
wire n_1391;
wire n_1392;
wire n_1393;
wire n_1394;
wire n_1395;
wire n_1396;
wire n_1397;
wire n_1398;
wire n_1399;
wire n_1400;
wire n_1401;
wire n_1402;
wire n_1403;
wire n_1404;
wire n_1405;
wire n_1406;
wire n_1407;
wire n_1408;
wire n_1409;
wire n_1410;
wire n_1411;
wire n_1412;
wire n_1413;
wire n_1414;
wire n_1415;
wire n_1416;
wire n_1417;
wire n_1418;
wire n_1419;
wire n_1420;
wire n_1421;
wire n_1422;
wire n_1423;
wire n_1424;
wire n_1425;
wire n_1426;
wire n_1427;
wire n_1428;
wire n_1429;
wire n_1430;
wire n_1431;
wire n_1432;
wire n_1433;
wire n_1434;
wire n_1435;
wire n_1436;
wire n_1437;
wire n_1438;
wire n_1439;
wire n_1440;
wire n_1441;
wire n_1442;
wire n_1443;
wire n_1444;
wire n_1445;
wire n_1446;
wire n_1447;
wire n_1448;
wire n_1449;
wire n_1450;
wire n_1451;
wire n_1452;
wire n_1453;
wire n_1454;
wire n_1455;
wire n_1456;
wire n_1457;
wire n_1458;
wire n_1459;
wire n_1460;
wire n_1461;
wire n_1462;
wire n_1463;
wire n_1464;
wire n_1465;
wire n_1466;
wire n_1467;
wire n_1468;
wire n_1469;
wire n_1470;
wire n_1471;
wire n_1472;
wire n_1473;
wire n_1474;
wire n_1475;
wire n_1476;
wire n_1477;
wire n_1478;
wire n_1479;
wire n_1480;
wire n_1481;
wire n_1482;
wire n_1483;
wire n_1484;
wire n_1485;
wire n_1486;
wire n_1487;
wire n_1488;
wire n_1489;
wire n_1490;
wire n_1491;
wire n_1492;
wire n_1493;
wire n_1494;
wire n_1495;
wire n_1496;
wire n_1497;
wire n_1498;
wire n_1499;
wire n_1500;
wire n_1501;
wire n_1502;
wire n_1503;
wire n_1504;
wire n_1505;
wire n_1506;
wire n_1507;
wire n_1508;
wire n_1509;
wire n_1510;
wire n_1511;
wire n_1512;
wire n_1513;
wire n_1514;
wire n_1515;
wire n_1516;
wire n_1517;
wire n_1518;
wire n_1519;
wire n_1520;
wire n_1521;
wire n_1522;
wire n_1523;
wire n_1524;
wire n_1525;
wire n_1526;
wire n_1527;
wire n_1528;
wire n_1529;
wire n_1530;
wire n_1531;
wire n_1532;
wire n_1533;
wire n_1534;
wire n_1535;
wire n_1536;
wire n_1537;
wire n_1538;
wire n_1539;
wire n_1540;
wire n_1541;
wire n_1542;
wire n_1543;
wire n_1544;
wire n_1545;
wire n_1546;
wire n_1547;
wire n_1548;
wire n_1549;
wire n_1550;
wire n_1551;
wire n_1552;
wire n_1553;
wire n_1554;
wire n_1555;
wire n_1556;
wire n_1557;
wire n_1558;
wire n_1559;
wire n_1560;
wire n_1561;
wire n_1562;
wire n_1563;
wire n_1564;
wire n_1565;
wire n_1566;
wire n_1567;
wire n_1568;
wire n_1569;
wire n_1570;
wire n_1571;
wire n_1572;
wire n_1573;
wire n_1574;
wire n_1575;
wire n_1576;
wire n_1577;
wire n_1578;
wire n_1579;
wire n_1580;
wire n_1581;
wire n_1582;
wire n_1583;
wire n_1584;
wire n_1585;
wire n_1586;
wire n_1587;
wire n_1588;
wire n_1589;
wire n_1590;
wire n_1591;
wire n_1592;
wire n_1593;
wire n_1594;
wire n_1595;
wire n_1596;
wire n_1597;
wire n_1598;
wire n_1599;
wire n_1600;
wire n_1601;
wire n_1602;
wire n_1603;
wire n_1604;
wire n_1605;
wire n_1606;
wire n_1607;
wire n_1608;
wire n_1609;
wire n_1610;
wire n_1611;
wire n_1612;
wire n_1613;
wire n_1614;
wire n_1615;
wire n_1616;
wire n_1617;
wire n_1618;
wire n_1619;
wire n_1620;
wire n_1621;
wire n_1622;
wire n_1623;
wire n_1624;
wire n_1625;
wire n_1626;
wire n_1627;
wire n_1628;
wire n_1629;
wire n_1630;
wire n_1631;
wire n_1632;
wire n_1633;
wire n_1634;
wire n_1635;
wire n_1636;
wire n_1637;
wire n_1638;
wire n_1639;
wire n_1640;
wire n_1641;
wire n_1642;
wire n_1643;
wire n_1644;
wire n_1645;
wire n_1646;
wire n_1647;
wire n_1648;
wire n_1649;
wire n_1650;
wire n_1651;
wire n_1652;
wire n_1653;
wire n_1654;
wire n_1655;
wire n_1656;
wire n_1657;
wire n_1658;
wire n_1659;
wire n_1660;
wire n_1661;
wire n_1662;
wire n_1663;
wire n_1664;
wire n_1665;
wire n_1666;
wire n_1667;
wire n_1668;
wire n_1669;
wire n_1670;
wire n_1671;
wire n_1672;
wire n_1673;
wire n_1674;
wire n_1675;
wire n_1676;
wire n_1677;
wire n_1678;
wire n_1679;
wire n_1680;
wire n_1681;
wire n_1682;
wire n_1683;
wire n_1684;
wire n_1685;
wire n_1686;
wire n_1687;
wire n_1688;
wire n_1689;
wire n_1690;
wire n_1691;
wire n_1692;
wire n_1693;
wire n_1694;
wire n_1695;
wire n_1696;
wire n_1697;
wire n_1698;
wire n_1699;
wire n_1700;
wire n_1701;
wire n_1702;
wire n_1703;
wire n_1704;
wire n_1705;
wire n_1706;
wire n_1707;
wire n_1708;
wire n_1709;
wire n_1710;
wire n_1711;
wire n_1712;
wire n_1713;
wire n_1714;
wire n_1715;
wire n_1716;
wire n_1717;
wire n_1718;
wire n_1719;
wire n_1720;
wire n_1721;
wire n_1722;
wire n_1723;
wire n_1724;
wire n_1725;
wire n_1726;
wire n_1727;
wire n_1728;
wire n_1729;
wire n_1730;
wire n_1731;
wire n_1732;
wire n_1733;
wire n_1734;
wire n_1735;
wire n_1736;
wire n_1737;
wire n_1738;
wire n_1739;
wire n_1740;
wire n_1741;
wire n_1742;
wire n_1743;
wire n_1744;
wire n_1745;
wire n_1746;
wire n_1747;
wire n_1748;
wire n_1749;
wire n_1750;
wire n_1751;
wire n_1752;
wire n_1753;
wire n_1754;
wire n_1755;
wire n_1756;
wire n_1757;
wire n_1758;
wire n_1759;
wire n_1760;
wire n_1761;
wire n_1762;
wire n_1763;
wire n_1764;
wire n_1765;
wire n_1766;
wire n_1767;
wire n_1768;
wire n_1769;
wire n_1770;
wire n_1771;
wire n_1772;
wire n_1773;
wire n_1774;
wire n_1775;
wire n_1776;
wire n_1777;
wire n_1778;
wire n_1779;
wire n_1780;
wire n_1781;
wire n_1782;
wire n_1783;
wire n_1784;
wire n_1785;
wire n_1786;
wire n_1787;
wire n_1788;
wire n_1789;
wire n_1790;
wire n_1791;
wire n_1792;
wire n_1793;
wire n_1794;
wire n_1795;
wire n_1796;
wire n_1797;
wire n_1798;
wire n_1799;
wire n_1800;
wire n_1801;
wire n_1802;
wire n_1803;
wire n_1804;
wire n_1805;
wire n_1806;
wire n_1807;
wire n_1808;
wire n_1809;
wire n_1810;
wire n_1811;
wire n_1812;
wire n_1813;
wire n_1814;
wire n_1815;
wire n_1816;
wire n_1817;
wire n_1818;
wire n_1819;
wire n_1820;
wire n_1821;
wire n_1822;
wire n_1823;
wire n_1824;
wire n_1825;
wire n_1826;
wire n_1827;
wire n_1828;
wire n_1829;
wire n_1830;
wire n_1831;
wire n_1832;
wire n_1833;
wire n_1834;
wire n_1835;
wire n_1836;
wire n_1837;
wire n_1838;
wire n_1839;
wire n_1840;
wire n_1841;
wire n_1842;
wire n_1843;
wire n_1844;
wire n_1845;
wire n_1846;
wire n_1847;
wire n_1848;
wire n_1849;
wire n_1850;
wire n_1851;
wire n_1852;
wire n_1853;
wire n_1854;
wire n_1855;
wire n_1856;
wire n_1857;
wire n_1858;
wire n_1859;
wire n_1860;
wire n_1861;
wire n_1862;
wire n_1863;
wire n_1864;
wire n_1865;
wire n_1866;
wire n_1867;
wire n_1868;
wire n_1869;
wire n_1870;
wire n_1871;
wire n_1872;
wire n_1873;
wire n_1874;
wire n_1875;
wire n_1876;
wire n_1877;
wire n_1878;
wire n_1879;
wire n_1880;
wire n_1881;
wire n_1882;
wire n_1883;
wire n_1884;
wire n_1885;
wire n_1886;
wire n_1887;
wire n_1888;
wire n_1889;
wire n_1890;
wire n_1891;
wire n_1892;
wire n_1893;
wire n_1894;
wire n_1895;
wire n_1896;
wire n_1897;
wire n_1898;
wire n_1899;
wire n_1900;
wire n_1901;
wire n_1902;
wire n_1903;
wire n_1904;
wire n_1905;
wire n_1906;
wire n_1907;
wire n_1908;
wire n_1909;
wire n_1910;
wire n_1911;
wire n_1912;
wire n_1913;
wire n_1914;
wire n_1915;
wire n_1916;
wire n_1917;
wire n_1918;
wire n_1919;
wire n_1920;
wire n_1921;
wire n_1922;
wire n_1923;
wire n_1924;
wire n_1925;
wire n_1926;
wire n_1927;
wire n_1928;
wire n_1929;
wire n_1930;
wire n_1931;
wire n_1932;
wire n_1933;
wire n_1934;
wire n_1935;
wire n_1936;
wire n_1937;
wire n_1938;
wire n_1939;
wire n_1940;
wire n_1941;
wire n_1942;
wire n_1943;
wire n_1944;
wire n_1945;
wire n_1946;
wire n_1947;
wire n_1948;
wire n_1949;
wire n_1950;
wire n_1951;
wire n_1952;
wire n_1953;
wire n_1954;
wire n_1955;
wire n_1956;
wire n_1957;
wire n_1958;
wire n_1959;
wire n_1960;
wire n_1961;
wire n_1962;
wire n_1963;
wire n_1964;
wire n_1965;
wire n_1966;
wire n_1967;
wire n_1968;
wire n_1969;
wire n_1970;
wire n_1971;
wire n_1972;
wire n_1973;
wire n_1974;
wire n_1975;
wire n_1976;
wire n_1977;
wire n_1978;
wire n_1979;
wire n_1980;
wire n_1981;
wire n_1982;
wire n_1983;
wire n_1984;
wire n_1985;
wire n_1986;
wire n_1987;
wire n_1988;
wire n_1989;
wire n_1990;
wire n_1991;
wire n_1992;
wire n_1993;
wire n_1994;
wire n_1995;
wire n_1996;
wire n_1997;
wire n_1998;
wire n_1999;
wire n_2000;
wire n_2001;
wire n_2002;
wire n_2003;
wire n_2004;
wire n_2005;
wire n_2006;
wire n_2007;
wire n_2008;
wire n_2009;
wire n_2010;
wire n_2011;
wire n_2012;
wire n_2013;
wire n_2014;
wire n_2015;
wire n_2016;
wire n_2017;
wire n_2018;
wire n_2019;
wire n_2020;
wire n_2021;
wire n_2022;
wire n_2023;
wire n_2024;
wire n_2025;
wire n_2026;
wire n_2027;
wire n_2028;
wire n_2029;
wire n_2030;
wire n_2031;
wire n_2032;
wire n_2033;
wire n_2034;
wire n_2035;
wire n_2036;
wire n_2037;
wire n_2038;
wire n_2039;
wire n_2040;
wire n_2041;
wire n_2042;
wire n_2043;
wire n_2044;
wire n_2045;
wire n_2046;
wire n_2047;
wire n_2048;
wire n_2049;
wire n_2050;
wire n_2051;
wire n_2052;
wire n_2053;
wire n_2054;
wire n_2055;
wire n_2056;
wire n_2057;
wire n_2058;
wire n_2059;
wire n_2060;
wire n_2061;
wire n_2062;
wire n_2063;
wire n_2064;
wire n_2065;
wire n_2066;
wire n_2067;
wire n_2068;
wire n_2069;
wire n_2070;
wire n_2071;
wire n_2072;
wire n_2073;
wire n_2074;
wire n_2075;
wire n_2076;
wire n_2077;
wire n_2078;
wire n_2079;
wire n_2080;
wire n_2081;
wire n_2082;
wire n_2083;
wire n_2084;
wire n_2085;
wire n_2086;
wire n_2087;
wire n_2088;
wire n_2089;
wire n_2090;
wire n_2091;
wire n_2092;
wire n_2093;
wire n_2094;
wire n_2095;
wire n_2096;
wire n_2097;
wire n_2098;
wire n_2099;
wire n_2100;
wire n_2101;
wire n_2102;
wire n_2103;
wire n_2104;
wire n_2105;
wire n_2106;
wire n_2107;
wire n_2108;
wire n_2109;
wire n_2110;
wire n_2111;
wire n_2112;
wire n_2113;
wire n_2114;
wire n_2115;
wire n_2116;
wire n_2117;
wire n_2118;
wire n_2119;
wire n_2120;
wire n_2121;
wire n_2122;
wire n_2123;
wire n_2124;
wire n_2125;
wire n_2126;
wire n_2127;
wire n_2128;
wire n_2129;
wire n_2130;
wire n_2131;
wire n_2132;
wire n_2133;
wire n_2134;
wire n_2135;
wire n_2136;
wire n_2137;
wire n_2138;
wire n_2139;
wire n_2140;
wire n_2141;
wire n_2142;
wire n_2143;
wire n_2144;
wire n_2145;
wire n_2146;
wire n_2147;
wire n_2148;
wire n_2149;
wire n_2150;
wire n_2151;
wire n_2152;
wire n_2153;
wire n_2154;
wire n_2155;
wire n_2156;
wire n_2157;
wire n_2158;
wire n_2159;
wire n_2160;
wire n_2161;
wire n_2162;
wire n_2163;
wire n_2164;
wire n_2165;
wire n_2166;
wire n_2167;
wire n_2168;
wire n_2169;
wire n_2170;
wire n_2171;
wire n_2172;
wire n_2173;
wire n_2174;
wire n_2175;
wire n_2176;
wire n_2177;
wire n_2178;
wire n_2179;
wire n_2180;
wire n_2181;
wire n_2182;
wire n_2183;
wire n_2184;
wire n_2185;
wire n_2186;
wire n_2187;
wire n_2188;
wire n_2189;
wire n_2190;
wire n_2191;
wire n_2192;
wire n_2193;
wire n_2194;
wire n_2195;
wire n_2196;
wire n_2197;
wire n_2198;
wire n_2199;
wire n_2200;
wire n_2201;
wire n_2202;
wire n_2203;
wire n_2204;
wire n_2205;
wire n_2206;
wire n_2207;
wire n_2208;
wire n_2209;
wire n_2210;
wire n_2211;
wire n_2212;
wire n_2213;
wire n_2214;
wire n_2215;
wire n_2216;
wire n_2217;
wire n_2218;
wire n_2219;
wire n_2220;
wire n_2221;
wire n_2222;
wire n_2223;
wire n_2224;
wire n_2225;
wire n_2226;
wire n_2227;
wire n_2228;
wire n_2229;
wire n_2230;
wire n_2231;
wire n_2232;
wire n_2233;
wire n_2234;
wire n_2235;
wire n_2236;
wire n_2237;
wire n_2238;
wire n_2239;
wire n_2240;
wire n_2241;
wire n_2242;
wire n_2243;
wire n_2244;
wire n_2245;
wire n_2246;
wire n_2247;
wire n_2248;
wire n_2249;
wire n_2250;
wire n_2251;
wire n_2252;
wire n_2253;
wire n_2254;
wire n_2255;
wire n_2256;
wire n_2257;
wire n_2258;
wire n_2259;
wire n_2260;
wire n_2261;
wire n_2262;
wire n_2263;
wire n_2264;
wire n_2265;
wire n_2266;
wire n_2267;
wire n_2268;
wire n_2269;
wire n_2270;
wire n_2271;
wire n_2272;
wire n_2273;
wire n_2274;
wire n_2275;
wire n_2276;
wire n_2277;
wire n_2278;
wire n_2279;
wire n_2280;
wire n_2281;
wire n_2282;
wire n_2283;
wire n_2284;
wire n_2285;
wire n_2286;
wire n_2287;
wire n_2288;
wire n_2289;
wire n_2290;
wire n_2291;
wire n_2292;
wire n_2293;
wire n_2294;
wire n_2295;
wire n_2296;
wire n_2297;
wire n_2298;
wire n_2299;
wire n_2300;
wire n_2301;
wire n_2302;
wire n_2303;
wire n_2304;
wire n_2305;
wire n_2306;
wire n_2307;
wire n_2308;
wire n_2309;
wire n_2310;
wire n_2311;
wire n_2312;
wire n_2313;
wire n_2314;
wire n_2315;
wire n_2316;
wire n_2317;
wire n_2318;
wire n_2319;
wire n_2320;
wire n_2321;
wire n_2322;
wire n_2323;
wire n_2324;
wire n_2325;
wire n_2326;
wire n_2327;
wire n_2328;
wire n_2329;
wire n_2330;
wire n_2331;
wire n_2332;
wire n_2333;
wire n_2334;
wire n_2335;
wire n_2336;
wire n_2337;
wire n_2338;
wire n_2339;
wire n_2340;
wire n_2341;
wire n_2342;
wire n_2343;
wire n_2344;
wire n_2345;
wire n_2346;
wire n_2347;
wire n_2348;
wire n_2349;
wire n_2350;
wire n_2351;
wire n_2352;
wire n_2353;
wire n_2354;
wire n_2355;
wire n_2356;
wire n_2357;
wire n_2358;
wire n_2359;
wire n_2360;
wire n_2361;
wire n_2362;
wire n_2363;
wire n_2364;
wire n_2365;
wire n_2366;
wire n_2367;
wire n_2368;
wire n_2369;
wire n_2370;
wire n_2371;
wire n_2372;
wire n_2373;
wire n_2374;
wire n_2375;
wire n_2376;
wire n_2377;
wire n_2378;
wire n_2379;
wire n_2380;
wire n_2381;
wire n_2382;
wire n_2383;
wire n_2384;
wire n_2385;
wire n_2386;
wire n_2387;
wire n_2388;
wire n_2389;
wire n_2390;
wire n_2391;
wire n_2392;
wire n_2393;
wire n_2394;
wire n_2395;
wire n_2396;
wire n_2397;
wire n_2398;
wire n_2399;
wire n_2400;
wire n_2401;
wire n_2402;
wire n_2403;
wire n_2404;
wire n_2405;
wire n_2406;
wire n_2407;
wire n_2408;
wire n_2409;
wire n_2410;
wire n_2411;
wire n_2412;
wire n_2413;
wire n_2414;
wire n_2415;
wire n_2416;
wire n_2417;
wire n_2418;
wire n_2419;
wire n_2420;
wire n_2421;
wire n_2422;
wire n_2423;
wire n_2424;
wire n_2425;
wire n_2426;
wire n_2427;
wire n_2428;
wire n_2429;
wire n_2430;
wire n_2431;
wire n_2432;
wire n_2433;
wire n_2434;
wire n_2435;
wire n_2436;
wire n_2437;
wire n_2438;
wire n_2439;
wire n_2440;
wire n_2441;
wire n_2442;
wire n_2443;
wire n_2444;
wire n_2445;
wire n_2446;
wire n_2447;
wire n_2448;
wire n_2449;
wire n_2450;
wire n_2451;
wire n_2452;
wire n_2453;
wire n_2454;
wire n_2455;
wire n_2456;
wire n_2457;
wire n_2458;
wire n_2459;
wire n_2460;
wire n_2461;
wire n_2462;
wire n_2463;
wire n_2464;
wire n_2465;
wire n_2466;
wire n_2467;
wire n_2468;
wire n_2469;
wire n_2470;
wire n_2471;
wire n_2472;
wire n_2473;
wire n_2474;
wire n_2475;
wire n_2476;
wire n_2477;
wire n_2478;
wire n_2479;
wire n_2480;
wire n_2481;
wire n_2482;
wire n_2483;
wire n_2484;
wire n_2485;
wire n_2486;
wire n_2487;
wire n_2488;
wire n_2489;
wire n_2490;
wire n_2491;
wire n_2492;
wire n_2493;
wire n_2494;
wire n_2495;
wire n_2496;
wire n_2497;
wire n_2498;
wire n_2499;
wire n_2500;
wire n_2501;
wire n_2502;
wire n_2503;
wire n_2504;
wire n_2505;
wire n_2506;
wire n_2507;
wire n_2508;
wire n_2509;
wire n_2510;
wire n_2511;
wire n_2512;
wire n_2513;
wire n_2514;
wire n_2515;
wire n_2516;
wire n_2517;
wire n_2518;
wire n_2519;
wire n_2520;
wire n_2521;
wire n_2522;
wire n_2523;
wire n_2524;
wire n_2525;
wire n_2526;
wire n_2527;
wire n_2528;
wire n_2529;
wire n_2530;
wire n_2531;
wire n_2532;
wire n_2533;
wire n_2534;
wire n_2535;
wire n_2536;
wire n_2537;
wire n_2538;
wire n_2539;
wire n_2540;
wire n_2541;
wire n_2542;
wire n_2543;
wire n_2544;
wire n_2545;
wire n_2546;
wire n_2547;
wire n_2548;
wire n_2549;
wire n_2550;
wire n_2551;
wire n_2552;
wire n_2553;
wire n_2554;
wire n_2555;
wire n_2556;
wire n_2557;
wire n_2558;
wire n_2559;
wire n_2560;
wire n_2561;
wire n_2562;
wire n_2563;
wire n_2564;
wire n_2565;
wire n_2566;
wire n_2567;
wire n_2568;
wire n_2569;
wire n_2570;
wire n_2571;
wire n_2572;
wire n_2573;
wire n_2574;
wire n_2575;
wire n_2576;
wire n_2577;
wire n_2578;
wire n_2579;
wire n_2580;
wire n_2581;
wire n_2582;
wire n_2583;
wire n_2584;
wire n_2585;
wire n_2586;
wire n_2587;
wire n_2588;
wire n_2589;
wire n_2590;
wire n_2591;
wire n_2592;
wire n_2593;
wire n_2594;
wire n_2595;
wire n_2596;
wire n_2597;
wire n_2598;
wire n_2599;
wire n_2600;
wire n_2601;
wire n_2602;
wire n_2603;
wire n_2604;
wire n_2605;
wire n_2606;
wire n_2607;
wire n_2608;
wire n_2609;
wire n_2610;
wire n_2611;
wire n_2612;
wire n_2613;
wire n_2614;
wire n_2615;
wire n_2616;
wire n_2617;
wire n_2618;
wire n_2619;
wire n_2620;
wire n_2621;
wire n_2622;
wire n_2623;
wire n_2624;
wire n_2625;
wire n_2626;
wire n_2627;
wire n_2628;
wire n_2629;
wire n_2630;
wire n_2631;
wire n_2632;
wire n_2633;
wire n_2634;
wire n_2635;
wire n_2636;
wire n_2637;
wire n_2638;
wire n_2639;
wire n_2640;
wire n_2641;
wire n_2642;
wire n_2643;
wire n_2644;
wire n_2645;
wire n_2646;
wire n_2647;
wire n_2648;
wire n_2649;
wire n_2650;
wire n_2651;
wire n_2652;
wire n_2653;
wire n_2654;
wire n_2655;
wire n_2656;
wire n_2657;
wire n_2658;
wire n_2659;
wire n_2660;
wire n_2661;
wire n_2662;
wire n_2663;
wire n_2664;
wire n_2665;
wire n_2666;
wire n_2667;
wire n_2668;
wire n_2669;
wire n_2670;
wire n_2671;
wire n_2672;
wire n_2673;
wire n_2674;
wire n_2675;
wire n_2676;
wire n_2677;
wire n_2678;
wire n_2679;
wire n_2680;
wire n_2681;
wire n_2682;
wire n_2683;
wire n_2684;
wire n_2685;
wire n_2686;
wire n_2687;
wire n_2688;
wire n_2689;
wire n_2690;
wire n_2691;
wire n_2692;
wire n_2693;
wire n_2694;
wire n_2695;
wire n_2696;
wire n_2697;
wire n_2698;
wire n_2699;
wire n_2700;
wire n_2701;
wire n_2702;
wire n_2703;
wire n_2704;
wire n_2705;
wire n_2706;
wire n_2707;
wire n_2708;
wire n_2709;
wire n_2710;
wire n_2711;
wire n_2712;
wire n_2713;
wire n_2714;
wire n_2715;
wire n_2716;
wire n_2717;
wire n_2718;
wire n_2719;
wire n_2720;
wire n_2721;
wire n_2722;
wire n_2723;
wire n_2724;
wire n_2725;
wire n_2726;
wire n_2727;
wire n_2728;
wire n_2729;
wire n_2730;
wire n_2731;
wire n_2732;
wire n_2733;
wire n_2734;
wire n_2735;
wire n_2736;
wire n_2737;
wire n_2738;
wire n_2739;
wire n_2740;
wire n_2741;
wire n_2742;
wire n_2743;
wire n_2744;
wire n_2745;
wire n_2746;
wire n_2747;
wire n_2748;
wire n_2749;
wire n_2750;
wire n_2751;
wire n_2752;
wire n_2753;
wire n_2754;
wire n_2755;
wire n_2756;
wire n_2757;
wire n_2758;
wire n_2759;
wire n_2760;
wire n_2761;
wire n_2762;
wire n_2763;
wire n_2764;
wire n_2765;
wire n_2766;
wire n_2767;
wire n_2768;
wire n_2769;
wire n_2770;
wire n_2771;
wire n_2772;
wire n_2773;
wire n_2774;
wire n_2775;
wire n_2776;
wire n_2777;
wire n_2778;
wire n_2779;
wire n_2780;
wire n_2781;
wire n_2782;
wire n_2783;
wire n_2784;
wire n_2785;
wire n_2786;
wire n_2787;
wire n_2788;
wire n_2789;
wire n_2790;
wire n_2791;
wire n_2792;
wire n_2793;
wire n_2794;
wire n_2795;
wire n_2796;
wire n_2797;
wire n_2798;
wire n_2799;
wire n_2800;
wire n_2801;
wire n_2802;
wire n_2803;
wire n_2804;
wire n_2805;
wire n_2806;
wire n_2807;
wire n_2808;
wire n_2809;
wire n_2810;
wire n_2811;
wire n_2812;
wire n_2813;
wire n_2814;
wire n_2815;
wire n_2816;
wire n_2817;
wire n_2818;
wire n_2819;
wire n_2820;
wire n_2821;
wire n_2822;
wire n_2823;
wire n_2824;
wire n_2825;
wire n_2826;
wire n_2827;
wire n_2828;
wire n_2829;
wire n_2830;
wire n_2831;
wire n_2832;
wire n_2833;
wire n_2834;
wire n_2835;
wire n_2836;
wire n_2837;
wire n_2838;
wire n_2839;
wire n_2840;
wire n_2841;
wire n_2842;
wire n_2843;
wire n_2844;
wire n_2845;
wire n_2846;
wire n_2847;
wire n_2848;
wire n_2849;
wire n_2850;
wire n_2851;
wire n_2852;
wire n_2853;
wire n_2854;
wire n_2855;
wire n_2856;
wire n_2857;
wire n_2858;
wire n_2859;
wire n_2860;
wire n_2861;
wire n_2862;
wire n_2863;
wire n_2864;
wire n_2865;
wire n_2866;
wire n_2867;
wire n_2868;
wire n_2869;
wire n_2870;
wire n_2871;
wire n_2872;
wire n_2873;
wire n_2874;
wire n_2875;
wire n_2876;
wire n_2877;
wire n_2878;
wire n_2879;
wire n_2880;
wire n_2881;
wire n_2882;
wire n_2883;
wire n_2884;
wire n_2885;
wire n_2886;
wire n_2887;
wire n_2888;
wire n_2889;
wire n_2890;
wire n_2891;
wire n_2892;
wire n_2893;
wire n_2894;
wire n_2895;
wire n_2896;
wire n_2897;
wire n_2898;
wire n_2899;
wire n_2900;
wire n_2901;
wire n_2902;
wire n_2903;
wire n_2904;
wire n_2905;
wire n_2906;
wire n_2907;
wire n_2908;
wire n_2909;
wire n_2910;
wire n_2911;
wire n_2912;
wire n_2913;
wire n_2914;
wire n_2915;
wire n_2916;
wire n_2917;
wire n_2918;
wire n_2919;
wire n_2920;
wire n_2921;
wire n_2922;
wire n_2923;
wire n_2924;
wire n_2925;
wire n_2926;
wire n_2927;
wire n_2928;
wire n_2929;
wire n_2930;
wire n_2931;
wire n_2932;
wire n_2933;
wire n_2934;
wire n_2935;
wire n_2936;
wire n_2937;
wire n_2938;
wire n_2939;
wire n_2940;
wire n_2941;
wire n_2942;
wire n_2943;
wire n_2944;
wire n_2945;
wire n_2946;
wire n_2947;
wire n_2948;
wire n_2949;
wire n_2950;
wire n_2951;
wire n_2952;
wire n_2953;
wire n_2954;
wire n_2955;
wire n_2956;
wire n_2957;
wire n_2958;
wire n_2959;
wire n_2960;
wire n_2961;
wire n_2962;
wire n_2963;
wire n_2964;
wire n_2965;
wire n_2966;
wire n_2967;
wire n_2968;
wire n_2969;
wire n_2970;
wire n_2971;
wire n_2972;
wire n_2973;
wire n_2974;
wire n_2975;
wire n_2976;
wire n_2977;
wire n_2978;
wire n_2979;
wire n_2980;
wire n_2981;
wire n_2982;
wire n_2983;
wire n_2984;
wire n_2985;
wire n_2986;
wire n_2987;
wire n_2988;
wire n_2989;
wire n_2990;
wire n_2991;
wire n_2992;
wire n_2993;
wire n_2994;
wire n_2995;
wire n_2996;
wire n_2997;
wire n_2998;
wire n_2999;
wire n_3000;
wire n_3001;
wire n_3002;
wire n_3003;
wire n_3004;
wire n_3005;
wire n_3006;
wire n_3007;
wire n_3008;
wire n_3009;
wire n_3010;
wire n_3011;
wire n_3012;
wire n_3013;
wire n_3014;
wire n_3015;
wire n_3016;
wire n_3017;
wire n_3018;
wire n_3019;
wire n_3020;
wire n_3021;
wire n_3022;
wire n_3023;
wire n_3024;
wire n_3025;
wire n_3026;
wire n_3027;
wire n_3028;
wire n_3029;
wire n_3030;
wire n_3031;
wire n_3032;
wire n_3033;
wire n_3034;
wire n_3035;
wire n_3036;
wire n_3037;
wire n_3038;
wire n_3039;
wire n_3040;
wire n_3041;
wire n_3042;
wire n_3043;
wire n_3044;
wire n_3045;
wire n_3046;
wire n_3047;
wire n_3048;
wire n_3049;
wire n_3050;
wire n_3051;
wire n_3052;
wire n_3053;
wire n_3054;
wire n_3055;
wire n_3056;
wire n_3057;
wire n_3058;
wire n_3059;
wire n_3060;
wire n_3061;
wire n_3062;
wire n_3063;
wire n_3064;
wire n_3065;
wire n_3066;
wire n_3067;
wire n_3068;
wire n_3069;
wire n_3070;
wire n_3071;
wire n_3072;
wire n_3073;
wire n_3074;
wire n_3075;
wire n_3076;
wire n_3077;
wire n_3078;
wire n_3079;
wire n_3080;
wire n_3081;
wire n_3082;
wire n_3083;
wire n_3084;
wire n_3085;
wire n_3086;
wire n_3087;
wire n_3088;
wire n_3089;
wire n_3090;
wire n_3091;
wire n_3092;
wire n_3093;
wire n_3094;
wire n_3095;
wire n_3096;
wire n_3097;
wire n_3098;
wire n_3099;
wire n_3100;
wire n_3101;
wire n_3102;
wire n_3103;
wire n_3104;
wire n_3105;
wire n_3106;
wire n_3107;
wire n_3108;
wire n_3109;
wire n_3110;
wire n_3111;
wire n_3112;
wire n_3113;
wire n_3114;
wire n_3115;
wire n_3116;
wire n_3117;
wire n_3118;
wire n_3119;
wire n_3120;
wire n_3121;
wire n_3122;
wire n_3123;
wire n_3124;
wire n_3125;
wire n_3126;
wire n_3127;
wire n_3128;
wire n_3129;
wire n_3130;
wire n_3131;
wire n_3132;
wire n_3133;
wire n_3134;
wire n_3135;
wire n_3136;
wire n_3137;
wire n_3138;
wire n_3139;
wire n_3140;
wire n_3141;
wire n_3142;
wire n_3143;
wire n_3144;
wire n_3145;
wire n_3146;
wire n_3147;
wire n_3148;
wire n_3149;
wire n_3150;
wire n_3151;
wire n_3152;
wire n_3153;
wire n_3154;
wire n_3155;
wire n_3156;
wire n_3157;
wire n_3158;
wire n_3159;
wire n_3160;
wire n_3161;
wire n_3162;
wire n_3163;
wire n_3164;
wire n_3165;
wire n_3166;
wire n_3167;
wire n_3168;
wire n_3169;
wire n_3170;
wire n_3171;
wire n_3172;
wire n_3173;
wire n_3174;
wire n_3175;
wire n_3176;
wire n_3177;
wire n_3178;
wire n_3179;
wire n_3180;
wire n_3181;
wire n_3182;
wire n_3183;
wire n_3184;
wire n_3185;
wire n_3186;
wire n_3187;
wire n_3188;
wire n_3189;
wire n_3190;
wire n_3191;
wire n_3192;
wire n_3193;
wire n_3194;
wire n_3195;
wire n_3196;
wire n_3197;
wire n_3198;
wire n_3199;
wire n_3200;
wire n_3201;
wire n_3202;
wire n_3203;
wire n_3204;
wire n_3205;
wire n_3206;
wire n_3207;
wire n_3208;
wire n_3209;
wire n_3210;
wire n_3211;
wire n_3212;
wire n_3213;
wire n_3214;
wire n_3215;
wire n_3216;
wire n_3217;
wire n_3218;
wire n_3219;
wire n_3220;
wire n_3221;
wire n_3222;
wire n_3223;
wire n_3224;
wire n_3225;
wire n_3226;
wire n_3227;
wire n_3228;
wire n_3229;
wire n_3230;
wire n_3231;
wire n_3232;
wire n_3233;
wire n_3234;
wire n_3235;
wire n_3236;
wire n_3237;
wire n_3238;
wire n_3239;
wire n_3240;
wire n_3241;
wire n_3242;
wire n_3243;
wire n_3244;
wire n_3245;
wire n_3246;
wire n_3247;
wire n_3248;
wire n_3249;
wire n_3250;
wire n_3251;
wire n_3252;
wire n_3253;
wire n_3254;
wire n_3255;
wire n_3256;
wire n_3257;
wire n_3258;
wire n_3259;
wire n_3260;
wire n_3261;
wire n_3262;
wire n_3263;
wire n_3264;
wire n_3265;
wire n_3266;
wire n_3267;
wire n_3268;
wire n_3269;
wire n_3270;
wire n_3271;
wire n_3272;
wire n_3273;
wire n_3274;
wire n_3275;
wire n_3276;
wire n_3277;
wire n_3278;
wire n_3279;
wire n_3280;
wire n_3281;
wire n_3282;
wire n_3283;
wire n_3284;
wire n_3285;
wire n_3286;
wire n_3287;
wire n_3288;
wire n_3289;
wire n_3290;
wire n_3291;
wire n_3292;
wire n_3293;
wire n_3294;
wire n_3295;
wire n_3296;
wire n_3297;
wire n_3298;
wire n_3299;
wire n_3300;
wire n_3301;
wire n_3302;
wire n_3303;
wire n_3304;
wire n_3305;
wire n_3306;
wire n_3307;
wire n_3308;
wire n_3309;
wire n_3310;
wire n_3311;
wire n_3312;
wire n_3313;
wire n_3314;
wire n_3315;
wire n_3316;
wire n_3317;
wire n_3318;
wire n_3319;
wire n_3320;
wire n_3321;
wire n_3322;
wire n_3323;
wire n_3324;
wire n_3325;
wire n_3326;
wire n_3327;
wire n_3328;
wire n_3329;
wire n_3330;
wire n_3331;
wire n_3332;
wire n_3333;
wire n_3334;
wire n_3335;
wire n_3336;
wire n_3337;
wire n_3338;
wire n_3339;
wire n_3340;
wire n_3341;
wire n_3342;
wire n_3343;
wire n_3344;
wire n_3345;
wire n_3346;
wire n_3347;
wire n_3348;
wire n_3349;
wire n_3350;
wire n_3351;
wire n_3352;
wire n_3353;
wire n_3354;
wire n_3355;
wire n_3356;
wire n_3357;
wire n_3358;
wire n_3359;
wire n_3360;
wire n_3361;
wire n_3362;
wire n_3363;
wire n_3364;
wire n_3365;
wire n_3366;
wire n_3367;
wire n_3368;
wire n_3369;
wire n_3370;
wire n_3371;
wire n_3372;
wire n_3373;
wire n_3374;
wire n_3375;
wire n_3376;
wire n_3377;
wire n_3378;
wire n_3379;
wire n_3380;
wire n_3381;
wire n_3382;
wire n_3383;
wire n_3384;
wire n_3385;
wire n_3386;
wire n_3387;
wire n_3388;
wire n_3389;
wire n_3390;
wire n_3391;
wire n_3392;
wire n_3393;
wire n_3394;
wire n_3395;
wire n_3396;
wire n_3397;
wire n_3398;
wire n_3399;
wire n_3400;
wire n_3401;
wire n_3402;
wire n_3403;
wire n_3404;
wire n_3405;
wire n_3406;
wire n_3407;
wire n_3408;
wire n_3409;
wire n_3410;
wire n_3411;
wire n_3412;
wire n_3413;
wire n_3414;
wire n_3415;
wire n_3416;
wire n_3417;
wire n_3418;
wire n_3419;
wire n_3420;
wire n_3421;
wire n_3422;
wire n_3423;
wire n_3424;
wire n_3425;
wire n_3426;
wire n_3427;
wire n_3428;
wire n_3429;
wire n_3430;
wire n_3431;
wire n_3432;
wire n_3433;
wire n_3434;
wire n_3435;
wire n_3436;
wire n_3437;
wire n_3438;
wire n_3439;
wire n_3440;
wire n_3441;
wire n_3442;
wire n_3443;
wire n_3444;
wire n_3445;
wire n_3446;
wire n_3447;
wire n_3448;
wire n_3449;
wire n_3450;
wire n_3451;
wire n_3452;
wire n_3453;
wire n_3454;
wire n_3455;
wire n_3456;
wire n_3457;
wire n_3458;
wire n_3459;
wire n_3460;
wire n_3461;
wire n_3462;
wire n_3463;
wire n_3464;
wire n_3465;
wire n_3466;
wire n_3467;
wire n_3468;
wire n_3469;
wire n_3470;
wire n_3471;
wire n_3472;
wire n_3473;
wire n_3474;
wire n_3475;
wire n_3476;
wire n_3477;
wire n_3478;
wire n_3479;
wire n_3480;
wire n_3481;
wire n_3482;
wire n_3483;
wire n_3484;
wire n_3485;
wire n_3486;
wire n_3487;
wire n_3488;
wire n_3489;
wire n_3490;
wire n_3491;
wire n_3492;
wire n_3493;
wire n_3494;
wire n_3495;
wire n_3496;
wire n_3497;
wire n_3498;
wire n_3499;
wire n_3500;
wire n_3501;
wire n_3502;
wire n_3503;
wire n_3504;
wire n_3505;
wire n_3506;
wire n_3507;
wire n_3508;
wire n_3509;
wire n_3510;
wire n_3511;
wire n_3512;
wire n_3513;
wire n_3514;
wire n_3515;
wire n_3516;
wire n_3517;
wire n_3518;
wire n_3519;
wire n_3520;
wire n_3521;
wire n_3522;
wire n_3523;
wire n_3524;
wire n_3525;
wire n_3526;
wire n_3527;
wire n_3528;
wire n_3529;
wire n_3530;
wire n_3531;
wire n_3532;
wire n_3533;
wire n_3534;
wire n_3535;
wire n_3536;
wire n_3537;
wire n_3538;
wire n_3539;
wire n_3540;
wire n_3541;
wire n_3542;
wire n_3543;
wire n_3544;
wire n_3545;
wire n_3546;
wire n_3547;
wire n_3548;
wire n_3549;
wire n_3550;
wire n_3551;
wire n_3552;
wire n_3553;
wire n_3554;
wire n_3555;
wire n_3556;
wire n_3557;
wire n_3558;
wire n_3559;
wire n_3560;
wire n_3561;
wire n_3562;
wire n_3563;
wire n_3564;
wire n_3565;
wire n_3566;
wire n_3567;
wire n_3568;
wire n_3569;
wire n_3570;
wire n_3571;
wire n_3572;
wire n_3573;
wire n_3574;
wire n_3575;
wire n_3576;
wire n_3577;
wire n_3578;
wire n_3579;
wire n_3580;
wire n_3581;
wire n_3582;
wire n_3583;
wire n_3584;
wire n_3585;
wire n_3586;
wire n_3587;
wire n_3588;
wire n_3589;
wire n_3590;
wire n_3591;
wire n_3592;
wire n_3593;
wire n_3594;
wire n_3595;
wire n_3596;
wire n_3597;
wire n_3598;
wire n_3599;
wire n_3600;
wire n_3601;
wire n_3602;
wire n_3603;
wire n_3604;
wire n_3605;
wire n_3606;
wire n_3607;
wire n_3608;
wire n_3609;
wire n_3610;
wire n_3611;
wire n_3612;
wire n_3613;
wire n_3614;
wire n_3615;
wire n_3616;
wire n_3617;
wire n_3618;
wire n_3619;
wire n_3620;
wire n_3621;
wire n_3622;
wire n_3623;
wire n_3624;
wire n_3625;
wire n_3626;
wire n_3627;
wire n_3628;
wire n_3629;
wire n_3630;
wire n_3631;
wire n_3632;
wire n_3633;
wire n_3634;
wire n_3635;
wire n_3636;
wire n_3637;
wire n_3638;
wire n_3639;
wire n_3640;
wire n_3641;
wire n_3642;
wire n_3643;
wire n_3644;
wire n_3645;
wire n_3646;
wire n_3647;
wire n_3648;
wire n_3649;
wire n_3650;
wire n_3651;
wire n_3652;
wire n_3653;
wire n_3654;
wire n_3655;
wire n_3656;
wire n_3657;
wire n_3658;
wire n_3659;
wire n_3660;
wire n_3661;
wire n_3662;
wire n_3663;
wire n_3664;
wire n_3665;
wire n_3666;
wire n_3667;
wire n_3668;
wire n_3669;
wire n_3670;
wire n_3671;
wire n_3672;
wire n_3673;
wire n_3674;
wire n_3675;
wire n_3676;
wire n_3677;
wire n_3678;
wire n_3679;
wire n_3680;
wire n_3681;
wire n_3682;
wire n_3683;
wire n_3684;
wire n_3685;
wire n_3686;
wire n_3687;
wire n_3688;
wire n_3689;
wire n_3690;
wire n_3691;
wire n_3692;
wire n_3693;
wire n_3694;
wire n_3695;
wire n_3696;
wire n_3697;
wire n_3698;
wire n_3699;
wire n_3700;
wire n_3701;
wire n_3702;
wire n_3703;
wire n_3704;
wire n_3705;
wire n_3706;
wire n_3707;
wire n_3708;
wire n_3709;
wire n_3710;
wire n_3711;
wire n_3712;
wire n_3713;
wire n_3714;
wire n_3715;
wire n_3716;
wire n_3717;
wire n_3718;
wire n_3719;
wire n_3720;
wire n_3721;
wire n_3722;
wire n_3723;
wire n_3724;
wire n_3725;
wire n_3726;
wire n_3727;
wire n_3728;
wire n_3729;
wire n_3730;
wire n_3731;
wire n_3732;
wire n_3733;
wire n_3734;
wire n_3735;
wire n_3736;
wire n_3737;
wire n_3738;
wire n_3739;
wire n_3740;
wire n_3741;
wire n_3742;
wire n_3743;
wire n_3744;
wire n_3745;
wire n_3746;
wire n_3747;
wire n_3748;
wire n_3749;
wire n_3750;
wire n_3751;
wire n_3752;
wire n_3753;
wire n_3754;
wire n_3755;
wire n_3756;
wire n_3757;
wire n_3758;
wire n_3759;
wire n_3760;
wire n_3761;
wire n_3762;
wire n_3763;
wire n_3764;
wire n_3765;
wire n_3766;
wire n_3767;
wire n_3768;
wire n_3769;
wire n_3770;
wire n_3771;
wire n_3772;
wire n_3773;
wire n_3774;
wire n_3775;
wire n_3776;
wire n_3777;
wire n_3778;
wire n_3779;
wire n_3780;
wire n_3781;
wire n_3782;
wire n_3783;
wire n_3784;
wire n_3785;
wire n_3786;
wire n_3787;
wire n_3788;
wire n_3789;
wire n_3790;
wire n_3791;
wire n_3792;
wire n_3793;
wire n_3794;
wire n_3795;
wire n_3796;
wire n_3797;
wire n_3798;
wire n_3799;
wire n_3800;
wire n_3801;
wire n_3802;
wire n_3803;
wire n_3804;
wire n_3805;
wire n_3806;
wire n_3807;
wire n_3808;
wire n_3809;
wire n_3810;
wire n_3811;
wire n_3812;
wire n_3813;
wire n_3814;
wire n_3815;
wire n_3816;
wire n_3817;
wire n_3818;
wire n_3819;
wire n_3820;
wire n_3821;
wire n_3822;
wire n_3823;
wire n_3824;
wire n_3825;
wire n_3826;
wire n_3827;
wire n_3828;
wire n_3829;
wire n_3830;
wire n_3831;
wire n_3832;
wire n_3833;
wire n_3834;
wire n_3835;
wire n_3836;
wire n_3837;
wire n_3838;
wire n_3839;
wire n_3840;
wire n_3841;
wire n_3842;
wire n_3843;
wire n_3844;
wire n_3845;
wire n_3846;
wire n_3847;
wire n_3848;
wire n_3849;
wire n_3850;
wire n_3851;
wire n_3852;
wire n_3853;
wire n_3854;
wire n_3855;
wire n_3856;
wire n_3857;
wire n_3858;
wire n_3859;
wire n_3860;
wire n_3861;
wire n_3862;
wire n_3863;
wire n_3864;
wire n_3865;
wire n_3866;
wire n_3867;
wire n_3868;
wire n_3869;
wire n_3870;
wire n_3871;
wire n_3872;
wire n_3873;
wire n_3874;
wire n_3875;
wire n_3876;
wire n_3877;
wire n_3878;
wire n_3879;
wire n_3880;
wire n_3881;
wire n_3882;
wire n_3883;
wire n_3884;
wire n_3885;
wire n_3886;
wire n_3887;
wire n_3888;
wire n_3889;
wire n_3890;
wire n_3891;
wire n_3892;
wire n_3893;
wire n_3894;
wire n_3895;
wire n_3896;
wire n_3897;
wire n_3898;
wire n_3899;
wire n_3900;
wire n_3901;
wire n_3902;
wire n_3903;
wire n_3904;
wire n_3905;
wire n_3906;
wire n_3907;
wire n_3908;
wire n_3909;
wire n_3910;
wire n_3911;
wire n_3912;
wire n_3913;
wire n_3914;
wire n_3915;
wire n_3916;
wire n_3917;
wire n_3918;
wire n_3919;
wire n_3920;
wire n_3921;
wire n_3922;
wire n_3923;
wire n_3924;
wire n_3925;
wire n_3926;
wire n_3927;
wire n_3928;
wire n_3929;
wire n_3930;
wire n_3931;
wire n_3932;
wire n_3933;
wire n_3934;
wire n_3935;
wire n_3936;
wire n_3937;
wire n_3938;
wire n_3939;
wire n_3940;
wire n_3941;
wire n_3942;
wire n_3943;
wire n_3944;
wire n_3945;
wire n_3946;
wire n_3947;
wire n_3948;
wire n_3949;
wire n_3950;
wire n_3951;
wire n_3952;
wire n_3953;
wire n_3954;
wire n_3955;
wire n_3956;
wire n_3957;
wire n_3958;
wire n_3959;
wire n_3960;
wire n_3961;
wire n_3962;
wire n_3963;
wire n_3964;
wire n_3965;
wire n_3966;
wire n_3967;
wire n_3968;
wire n_3969;
wire n_3970;
wire n_3971;
wire n_3972;
wire n_3973;
wire n_3974;
wire n_3975;
wire n_3976;
wire n_3977;
wire n_3978;
wire n_3979;
wire n_3980;
wire n_3981;
wire n_3982;
wire n_3983;
wire n_3984;
wire n_3985;
wire n_3986;
wire n_3987;
wire n_3988;
wire n_3989;
wire n_3990;
wire n_3991;
wire n_3992;
wire n_3993;
wire n_3994;
wire n_3995;
wire n_3996;
wire n_3997;
wire n_3998;
wire n_3999;
wire n_4000;
wire n_4001;
wire n_4002;
wire n_4003;
wire n_4004;
wire n_4005;
wire n_4006;
wire n_4007;
wire n_4008;
wire n_4009;
wire n_4010;
wire n_4011;
wire n_4012;
wire n_4013;
wire n_4014;
wire n_4015;
wire n_4016;
wire n_4017;
wire n_4018;
wire n_4019;
wire n_4020;
wire n_4021;
wire n_4022;
wire n_4023;
wire n_4024;
wire n_4025;
wire n_4026;
wire n_4027;
wire n_4028;
wire n_4029;
wire n_4030;
wire n_4031;
wire n_4032;
wire n_4033;
wire n_4034;
wire n_4035;
wire n_4036;
wire n_4037;
wire n_4038;
wire n_4039;
wire n_4040;
wire n_4041;
wire n_4042;
wire n_4043;
wire n_4044;
wire n_4045;
wire n_4046;
wire n_4047;
wire n_4048;
wire n_4049;
wire n_4050;
wire n_4051;
wire n_4052;
wire n_4053;
wire n_4054;
wire n_4055;
wire n_4056;
wire n_4057;
wire n_4058;
wire n_4059;
wire n_4060;
wire n_4061;
wire n_4062;
wire n_4063;
wire n_4064;
wire n_4065;
wire n_4066;
wire n_4067;
wire n_4068;
wire n_4069;
wire n_4070;
wire n_4071;
wire n_4072;
wire n_4073;
wire n_4074;
wire n_4075;
wire n_4076;
wire n_4077;
wire n_4078;
wire n_4079;
wire n_4080;
wire n_4081;
wire n_4082;
wire n_4083;
wire n_4084;
wire n_4085;
wire n_4086;
wire n_4087;
wire n_4088;
wire n_4089;
wire n_4090;
wire n_4091;
wire n_4092;
wire n_4093;
wire n_4094;
wire n_4095;
wire n_4096;
wire n_4097;
wire n_4098;
wire n_4099;
wire n_4100;
wire n_4101;
wire n_4102;
wire n_4103;
wire n_4104;
wire n_4105;
wire n_4106;
wire n_4107;
wire n_4108;
wire n_4109;
wire n_4110;
wire n_4111;
wire n_4112;
wire n_4113;
wire n_4114;
wire n_4115;
wire n_4116;
wire n_4117;
wire n_4118;
wire n_4119;
wire n_4120;
wire n_4121;
wire n_4122;
wire n_4123;
wire n_4124;
wire n_4125;
wire n_4126;
wire n_4127;
wire n_4128;
wire n_4129;
wire n_4130;
wire n_4131;
wire n_4132;
wire n_4133;
wire n_4134;
wire n_4135;
wire n_4136;
wire n_4137;
wire n_4138;
wire n_4139;
wire n_4140;
wire n_4141;
wire n_4142;
wire n_4143;
wire n_4144;
wire n_4145;
wire n_4146;
wire n_4147;
wire n_4148;
wire n_4149;
wire n_4150;
wire n_4151;
wire n_4152;
wire n_4153;
wire n_4154;
wire n_4155;
wire n_4156;
wire n_4157;
wire n_4158;
wire n_4159;
wire n_4160;
wire n_4161;
wire n_4162;
wire n_4163;
wire n_4164;
wire n_4165;
wire n_4166;
wire n_4167;
wire n_4168;
wire n_4169;
wire n_4170;
wire n_4171;
wire n_4172;
wire n_4173;
wire n_4174;
wire n_4175;
wire n_4176;
wire n_4177;
wire n_4178;
wire n_4179;
wire n_4180;
wire n_4181;
wire n_4182;
wire n_4183;
wire n_4184;
wire n_4185;
wire n_4186;
wire n_4187;
wire n_4188;
wire n_4189;
wire n_4190;
wire n_4191;
wire n_4192;
wire n_4193;
wire n_4194;
wire n_4195;
wire n_4196;
wire n_4197;
wire n_4198;
wire n_4199;
wire n_4200;
wire n_4201;
wire n_4202;
wire n_4203;
wire n_4204;
wire n_4205;
wire n_4206;
wire n_4207;
wire n_4208;
wire n_4209;
wire n_4210;
wire n_4211;
wire n_4212;
wire n_4213;
wire n_4214;
wire n_4215;
wire n_4216;
wire n_4217;
wire n_4218;
wire n_4219;
wire n_4220;
wire n_4221;
wire n_4222;
wire n_4223;
wire n_4224;
wire n_4225;
wire n_4226;
wire n_4227;
wire n_4228;
wire n_4229;
wire n_4230;
wire n_4231;
wire n_4232;
wire n_4233;
wire n_4234;
wire n_4235;
wire n_4236;
wire n_4237;
wire n_4238;
wire n_4239;
wire n_4240;
wire n_4241;
wire n_4242;
wire n_4243;
wire n_4244;
wire n_4245;
wire n_4246;
wire n_4247;
wire n_4248;
wire n_4249;
wire n_4250;
wire n_4251;
wire n_4252;
wire n_4253;
wire n_4254;
wire n_4255;
wire n_4256;
wire n_4257;
wire n_4258;
wire n_4259;
wire n_4260;
wire n_4261;
wire n_4262;
wire n_4263;
wire n_4264;
wire n_4265;
wire n_4266;
wire n_4267;
wire n_4268;
wire n_4269;
wire n_4270;
wire n_4271;
wire n_4272;
wire n_4273;
wire n_4274;
wire n_4275;
wire n_4276;
wire n_4277;
wire n_4278;
wire n_4279;
wire n_4280;
wire n_4281;
wire n_4282;
wire n_4283;
wire n_4284;
wire n_4285;
wire n_4286;
wire n_4287;
wire n_4288;
wire n_4289;
wire n_4290;
wire n_4291;
wire n_4292;
wire n_4293;
wire n_4294;
wire n_4295;
wire n_4296;
wire n_4297;
wire n_4298;
wire n_4299;
wire n_4300;
wire n_4301;
wire n_4302;
wire n_4303;
wire n_4304;
wire n_4305;
wire n_4306;
wire n_4307;
wire n_4308;
wire n_4309;
wire n_4310;
wire n_4311;
wire n_4312;
wire n_4313;
wire n_4314;
wire n_4315;
wire n_4316;
wire n_4317;
wire n_4318;
wire n_4319;
wire n_4320;
wire n_4321;
wire n_4322;
wire n_4323;
wire n_4324;
wire n_4325;
wire n_4326;
wire n_4327;
wire n_4328;
wire n_4329;
wire n_4330;
wire n_4331;
wire n_4332;
wire n_4333;
wire n_4334;
wire n_4335;
wire n_4336;
wire n_4337;
wire n_4338;
wire n_4339;
wire n_4340;
wire n_4341;
wire n_4342;
wire n_4343;
wire n_4344;
wire n_4345;
wire n_4346;
wire n_4347;
wire n_4348;
wire n_4349;
wire n_4350;
wire n_4351;
wire n_4352;
wire n_4353;
wire n_4354;
wire n_4355;
wire n_4356;
wire n_4357;
wire n_4358;
wire n_4359;
wire n_4360;
wire n_4361;
wire n_4362;
wire n_4363;
wire n_4364;
wire n_4365;
wire n_4366;
wire n_4367;
wire n_4368;
wire n_4369;
wire n_4370;
wire n_4371;
wire n_4372;
wire n_4373;
wire n_4374;
wire n_4375;
wire n_4376;
wire n_4377;
wire n_4378;
wire n_4379;
wire n_4380;
wire n_4381;
wire n_4382;
wire n_4383;
wire n_4384;
wire n_4385;
wire n_4386;
wire n_4387;
wire n_4388;
wire n_4389;
wire n_4390;
wire n_4391;
wire n_4392;
wire n_4393;
wire n_4394;
wire n_4395;
wire n_4396;
wire n_4397;
wire n_4398;
wire n_4399;
wire n_4400;
wire n_4401;
wire n_4402;
wire n_4403;
wire n_4404;
wire n_4405;
wire n_4406;
wire n_4407;
wire n_4408;
wire n_4409;
wire n_4410;
wire n_4411;
wire n_4412;
wire n_4413;
wire n_4414;
wire n_4415;
wire n_4416;
wire n_4417;
wire n_4418;
wire n_4419;
wire n_4420;
wire n_4421;
wire n_4422;
wire n_4423;
wire n_4424;
wire n_4425;
wire n_4426;
wire n_4427;
wire n_4428;
wire n_4429;
wire n_4430;
wire n_4431;
wire n_4432;
wire n_4433;
wire n_4434;
wire n_4435;
wire n_4436;
wire n_4437;
wire n_4438;
wire n_4439;
wire n_4440;
wire n_4441;
wire n_4442;
wire n_4443;
wire n_4444;
wire n_4445;
wire n_4446;
wire n_4447;
wire n_4448;
wire n_4449;
wire n_4450;
wire n_4451;
wire n_4452;
wire n_4453;
wire n_4454;
wire n_4455;
wire n_4456;
wire n_4457;
wire n_4458;
wire n_4459;
wire n_4460;
wire n_4461;
wire n_4462;
wire n_4463;
wire n_4464;
wire n_4465;
wire n_4466;
wire n_4467;
wire n_4468;
wire n_4469;
wire n_4470;
wire n_4471;
wire n_4472;
wire n_4473;
wire n_4474;
wire n_4475;
wire n_4476;
wire n_4477;
wire n_4478;
wire n_4479;
wire n_4480;
wire n_4481;
wire n_4482;
wire n_4483;
wire n_4484;
wire n_4485;
wire n_4486;
wire n_4487;
wire n_4488;
wire n_4489;
wire n_4490;
wire n_4491;
wire n_4492;
wire n_4493;
wire n_4494;
wire n_4495;
wire n_4496;
wire n_4497;
wire n_4498;
wire n_4499;
wire n_4500;
wire n_4501;
wire n_4502;
wire n_4503;
wire n_4504;
wire n_4505;
wire n_4506;
wire n_4507;
wire n_4508;
wire n_4509;
wire n_4510;
wire n_4511;
wire n_4512;
wire n_4513;
wire n_4514;
wire n_4515;
wire n_4516;
wire n_4517;
wire n_4518;
wire n_4519;
wire n_4520;
wire n_4521;
wire n_4522;
wire n_4523;
wire n_4524;
wire n_4525;
wire n_4526;
wire n_4527;
wire n_4528;
wire n_4529;
wire n_4530;
wire n_4531;
wire n_4532;
wire n_4533;
wire n_4534;
wire n_4535;
wire n_4536;
wire n_4537;
wire n_4538;
wire n_4539;
wire n_4540;
wire n_4541;
wire n_4542;
wire n_4543;
wire n_4544;
wire n_4545;
wire n_4546;
wire n_4547;
wire n_4548;
wire n_4549;
wire n_4550;
wire n_4551;
wire n_4552;
wire n_4553;
wire n_4554;
wire n_4555;
wire n_4556;
wire n_4557;
wire n_4558;
wire n_4559;
wire n_4560;
wire n_4561;
wire n_4562;
wire n_4563;
wire n_4564;
wire n_4565;
wire n_4566;
wire n_4567;
wire n_4568;
wire n_4569;
wire n_4570;
wire n_4571;
wire n_4572;
wire n_4573;
wire n_4574;
wire n_4575;
wire n_4576;
wire n_4577;
wire n_4578;
wire n_4579;
wire n_4580;
wire n_4581;
wire n_4582;
wire n_4583;
wire n_4584;
wire n_4585;
wire n_4586;
wire n_4587;
wire n_4588;
wire n_4589;
wire n_4590;
wire n_4591;
wire n_4592;
wire n_4593;
wire n_4594;
wire n_4595;
wire n_4596;
wire n_4597;
wire n_4598;
wire n_4599;
wire n_4600;
wire n_4601;
wire n_4602;
wire n_4603;
wire n_4604;
wire n_4605;
wire n_4606;
wire n_4607;
wire n_4608;
wire n_4609;
wire n_4610;
wire n_4611;
wire n_4612;
wire n_4613;
wire n_4614;
wire n_4615;
wire n_4616;
wire n_4617;
wire n_4618;
wire n_4619;
wire n_4620;
wire n_4621;
wire n_4622;
wire n_4623;
wire n_4624;
wire n_4625;
wire n_4626;
wire n_4627;
wire n_4628;
wire n_4629;
wire n_4630;
wire n_4631;
wire n_4632;
wire n_4633;
wire n_4634;
wire n_4635;
wire n_4636;
wire n_4637;
wire n_4638;
wire n_4639;
wire n_4640;
wire n_4641;
wire n_4642;
wire n_4643;
wire n_4644;
wire n_4645;
wire n_4646;
wire n_4647;
wire n_4648;
wire n_4649;
wire n_4650;
wire n_4651;
wire n_4652;
wire n_4653;
wire n_4654;
wire n_4655;
wire n_4656;
wire n_4657;
wire n_4658;
wire n_4659;
wire n_4660;
wire n_4661;
wire n_4662;
wire n_4663;
wire n_4664;
wire n_4665;
wire n_4666;
wire n_4667;
wire n_4668;
wire n_4669;
wire n_4670;
wire n_4671;
wire n_4672;
wire n_4673;
wire n_4674;
wire n_4675;
wire n_4676;
wire n_4677;
wire n_4678;
wire n_4679;
wire n_4680;
wire n_4681;
wire n_4682;
wire n_4683;
wire n_4684;
wire n_4685;
wire n_4686;
wire n_4687;
wire n_4688;
wire n_4689;
wire n_4690;
wire n_4691;
wire n_4692;
wire n_4693;
wire n_4694;
wire n_4695;
wire n_4696;
wire n_4697;
wire n_4698;
wire n_4699;
wire n_4700;
wire n_4701;
wire n_4702;
wire n_4703;
wire n_4704;
wire n_4705;
wire n_4706;
wire n_4707;
wire n_4708;
wire n_4709;
wire n_4710;
wire n_4711;
wire n_4712;
wire n_4713;
wire n_4714;
wire n_4715;
wire n_4716;
wire n_4717;
wire n_4718;
wire n_4719;
wire n_4720;
wire n_4721;
wire n_4722;
wire n_4723;
wire n_4724;
wire n_4725;
wire n_4726;
wire n_4727;
wire n_4728;
wire n_4729;
wire n_4730;
wire n_4731;
wire n_4732;
wire n_4733;
wire n_4734;
wire n_4735;
wire n_4736;
wire n_4737;
wire n_4738;
wire n_4739;
wire n_4740;
wire n_4741;
wire n_4742;
wire n_4743;
wire n_4744;
wire n_4745;
wire n_4746;
wire n_4747;
wire n_4748;
wire n_4749;
wire n_4750;
wire n_4751;
wire n_4752;
wire n_4753;
wire n_4754;
wire n_4755;
wire n_4756;
wire n_4757;
wire n_4758;
wire n_4759;
wire n_4760;
wire n_4761;
wire n_4762;
wire n_4763;
wire n_4764;
wire n_4765;
wire n_4766;
wire n_4767;
wire n_4768;
wire n_4769;
wire n_4770;
wire n_4771;
wire n_4772;
wire n_4773;
wire n_4774;
wire n_4775;
wire n_4776;
wire n_4777;
wire n_4778;
wire n_4779;
wire n_4780;
wire n_4781;
wire n_4782;
wire n_4783;
wire n_4784;
wire n_4785;
wire n_4786;
wire n_4787;
wire n_4788;
wire n_4789;
wire n_4790;
wire n_4791;
wire n_4792;
wire n_4793;
wire n_4794;
wire n_4795;
wire n_4796;
wire n_4797;
wire n_4798;
wire n_4799;
wire n_4800;
wire n_4801;
wire n_4802;
wire n_4803;
wire n_4804;
wire n_4805;
wire n_4806;
wire n_4807;
wire n_4808;
wire n_4809;
wire n_4810;
wire n_4811;
wire n_4812;
wire n_4813;
wire n_4814;
wire n_4815;
wire n_4816;
wire n_4817;
wire n_4818;
wire n_4819;
wire n_4820;
wire n_4821;
wire n_4822;
wire n_4823;
wire n_4824;
wire n_4825;
wire n_4826;
wire n_4827;
wire n_4828;
wire n_4829;
wire n_4830;
wire n_4831;
wire n_4832;
wire n_4833;
wire n_4834;
wire n_4835;
wire n_4836;
wire n_4837;
wire n_4838;
wire n_4839;
wire n_4840;
wire n_4841;
wire n_4842;
wire n_4843;
wire n_4844;
wire n_4845;
wire n_4846;
wire n_4847;
wire n_4848;
wire n_4849;
wire n_4850;
wire n_4851;
wire n_4852;
wire n_4853;
wire n_4854;
wire n_4855;
wire n_4856;
wire n_4857;
wire n_4858;
wire n_4859;
wire n_4860;
wire n_4861;
wire n_4862;
wire n_4863;
wire n_4864;
wire n_4865;
wire n_4866;
wire n_4867;
wire n_4868;
wire n_4869;
wire n_4870;
wire n_4871;
wire n_4872;
wire n_4873;
wire n_4874;
wire n_4875;
wire n_4876;
wire n_4877;
wire n_4878;
wire n_4879;
wire n_4880;
wire n_4881;
wire n_4882;
wire n_4883;
wire n_4884;
wire n_4885;
wire n_4886;
wire n_4887;
wire n_4888;
wire n_4889;
wire n_4890;
wire n_4891;
wire n_4892;
wire n_4893;
wire n_4894;
wire n_4895;
wire n_4896;
wire n_4897;
wire n_4898;
wire n_4899;
wire n_4900;
wire n_4901;
wire n_4902;
wire n_4903;
wire n_4904;
wire n_4905;
wire n_4906;
wire n_4907;
wire n_4908;
wire n_4909;
wire n_4910;
wire n_4911;
wire n_4912;
wire n_4913;
wire n_4914;
wire n_4915;
wire n_4916;
wire n_4917;
wire n_4918;
wire n_4919;
wire n_4920;
wire n_4921;
wire n_4922;
wire n_4923;
wire n_4924;
wire n_4925;
wire n_4926;
wire n_4927;
wire n_4928;
wire n_4929;
wire n_4930;
wire n_4931;
wire n_4932;
wire n_4933;
wire n_4934;
wire n_4935;
wire n_4936;
wire n_4937;
wire n_4938;
wire n_4939;
wire n_4940;
wire n_4941;
wire n_4942;
wire n_4943;
wire n_4944;
wire n_4945;
wire n_4946;
wire n_4947;
wire n_4948;
wire n_4949;
wire n_4950;
wire n_4951;
wire n_4952;
wire n_4953;
wire n_4954;
wire n_4955;
wire n_4956;
wire n_4957;
wire n_4958;
wire n_4959;
wire n_4960;
wire n_4961;
wire n_4962;
wire n_4963;
wire n_4964;
wire n_4965;
wire n_4966;
wire n_4967;
wire n_4968;
wire n_4969;
wire n_4970;
wire n_4971;
wire n_4972;
wire n_4973;
wire n_4974;
wire n_4975;
wire n_4976;
wire n_4977;
wire n_4978;
wire n_4979;
wire n_4980;
wire n_4981;
wire n_4982;
wire n_4983;
wire n_4984;
wire n_4985;
wire n_4986;
wire n_4987;
wire n_4988;
wire n_4989;
wire n_4990;
wire n_4991;
wire n_4992;
wire n_4993;
wire n_4994;
wire n_4995;
wire n_4996;
wire n_4997;
wire n_4998;
wire n_4999;
wire n_5000;
wire n_5001;
wire n_5002;
wire n_5003;
wire n_5004;
wire n_5005;
wire n_5006;
wire n_5007;
wire n_5008;
wire n_5009;
wire n_5010;
wire n_5011;
wire n_5012;
wire n_5013;
wire n_5014;
wire n_5015;
wire n_5016;
wire n_5017;
wire n_5018;
wire n_5019;
wire n_5020;
wire n_5021;
wire n_5022;
wire n_5023;
wire n_5024;
wire n_5025;
wire n_5026;
wire n_5027;
wire n_5028;
wire n_5029;
wire n_5030;
wire n_5031;
wire n_5032;
wire n_5033;
wire n_5034;
wire n_5035;
wire n_5036;
wire n_5037;
wire n_5038;
wire n_5039;
wire n_5040;
wire n_5041;
wire n_5042;
wire n_5043;
wire n_5044;
wire n_5045;
wire n_5046;
wire n_5047;
wire n_5048;
wire n_5049;
wire n_5050;
wire n_5051;
wire n_5052;
wire n_5053;
wire n_5054;
wire n_5055;
wire n_5056;
wire n_5057;
wire n_5058;
wire n_5059;
wire n_5060;
wire n_5061;
wire n_5062;
wire n_5063;
wire n_5064;
wire n_5065;
wire n_5066;
wire n_5067;
wire n_5068;
wire n_5069;
wire n_5070;
wire n_5071;
wire n_5072;
wire n_5073;
wire n_5074;
wire n_5075;
wire n_5076;
wire n_5077;
wire n_5078;
wire n_5079;
wire n_5080;
wire n_5081;
wire n_5082;
wire n_5083;
wire n_5084;
wire n_5085;
wire n_5086;
wire n_5087;
wire n_5088;
wire n_5089;
wire n_5090;
wire n_5091;
wire n_5092;
wire n_5093;
wire n_5094;
wire n_5095;
wire n_5096;
wire n_5097;
wire n_5098;
wire n_5099;
wire n_5100;
wire n_5101;
wire n_5102;
wire n_5103;
wire n_5104;
wire n_5105;
wire n_5106;
wire n_5107;
wire n_5108;
wire n_5109;
wire n_5110;
wire n_5111;
wire n_5112;
wire n_5113;
wire n_5114;
wire n_5115;
wire n_5116;
wire n_5117;
wire n_5118;
wire n_5119;
wire n_5120;
wire n_5121;
wire n_5122;
wire n_5123;
wire n_5124;
wire n_5125;
wire n_5126;
wire n_5127;
wire n_5128;
wire n_5129;
wire n_5130;
wire n_5131;
wire n_5132;
wire n_5133;
wire n_5134;
wire n_5135;
wire n_5136;
wire n_5137;
wire n_5138;
wire n_5139;
wire n_5140;
wire n_5141;
wire n_5142;
wire n_5143;
wire n_5144;
wire n_5145;
wire n_5146;
wire n_5147;
wire n_5148;
wire n_5149;
wire n_5150;
wire n_5151;
wire n_5152;
wire n_5153;
wire n_5154;
wire n_5155;
wire n_5156;
wire n_5157;
wire n_5158;
wire n_5159;
wire n_5160;
wire n_5161;
wire n_5162;
wire n_5163;
wire n_5164;
wire n_5165;
wire n_5166;
wire n_5167;
wire n_5168;
wire n_5169;
wire n_5170;
wire n_5171;
wire n_5172;
wire n_5173;
wire n_5174;
wire n_5175;
wire n_5176;
wire n_5177;
wire n_5178;
wire n_5179;
wire n_5180;
wire n_5181;
wire n_5182;
wire n_5183;
wire n_5184;
wire n_5185;
wire n_5186;
wire n_5187;
wire n_5188;
wire n_5189;
wire n_5190;
wire n_5191;
wire n_5192;
wire n_5193;
wire n_5194;
wire n_5195;
wire n_5196;
wire n_5197;
wire n_5198;
wire n_5199;
wire n_5200;
wire n_5201;
wire n_5202;
wire n_5203;
wire n_5204;
wire n_5205;
wire n_5206;
wire n_5207;
wire n_5208;
wire n_5209;
wire n_5210;
wire n_5211;
wire n_5212;
wire n_5213;
wire n_5214;
wire n_5215;
wire n_5216;
wire n_5217;
wire n_5218;
wire n_5219;
wire n_5220;
wire n_5221;
wire n_5222;
wire n_5223;
wire n_5224;
wire n_5225;
wire n_5226;
wire n_5227;
wire n_5228;
wire n_5229;
wire n_5230;
wire n_5231;
wire n_5232;
wire n_5233;
wire n_5234;
wire n_5235;
wire n_5236;
wire n_5237;
wire n_5238;
wire n_5239;
wire n_5240;
wire n_5241;
wire n_5242;
wire n_5243;
wire n_5244;
wire n_5245;
wire n_5246;
wire n_5247;
wire n_5248;
wire n_5249;
wire n_5250;
wire n_5251;
wire n_5252;
wire n_5253;
wire n_5254;
wire n_5255;
wire n_5256;
wire n_5257;
wire n_5258;
wire n_5259;
wire n_5260;
wire n_5261;
wire n_5262;
wire n_5263;
wire n_5264;
wire n_5265;
wire n_5266;
wire n_5267;
wire n_5268;
wire n_5269;
wire n_5270;
wire n_5271;
wire n_5272;
wire n_5273;
wire n_5274;
wire n_5275;
wire n_5276;
wire n_5277;
wire n_5278;
wire n_5279;
wire n_5280;
wire n_5281;
wire n_5282;
wire n_5283;
wire n_5284;
wire n_5285;
wire n_5286;
wire n_5287;
wire n_5288;
wire n_5289;
wire n_5290;
wire n_5291;
wire n_5292;
wire n_5293;
wire n_5294;
wire n_5295;
wire n_5296;
wire n_5297;
wire n_5298;
wire n_5299;
wire n_5300;
wire n_5301;
wire n_5302;
wire n_5303;
wire n_5304;
wire n_5305;
wire n_5306;
wire n_5307;
wire n_5308;
wire n_5309;
wire n_5310;
wire n_5311;
wire n_5312;
wire n_5313;
wire n_5314;
wire n_5315;
wire n_5316;
wire n_5317;
wire n_5318;
wire n_5319;
wire n_5320;
wire n_5321;
wire n_5322;
wire n_5323;
wire n_5324;
wire n_5325;
wire n_5326;
wire n_5327;
wire n_5328;
wire n_5329;
wire n_5330;
wire n_5331;
wire n_5332;
wire n_5333;
wire n_5334;
wire n_5335;
wire n_5336;
wire n_5337;
wire n_5338;
wire n_5339;
wire n_5340;
wire n_5341;
wire n_5342;
wire n_5343;
wire n_5344;
wire n_5345;
wire n_5346;
wire n_5347;
wire n_5348;
wire n_5349;
wire n_5350;
wire n_5351;
wire n_5352;
wire n_5353;
wire n_5354;
wire n_5355;
wire n_5356;
wire n_5357;
wire n_5358;
wire n_5359;
wire n_5360;
wire n_5361;
wire n_5362;
wire n_5363;
wire n_5364;
wire n_5365;
wire n_5366;
wire n_5367;
wire n_5368;
wire n_5369;
wire n_5370;
wire n_5371;
wire n_5372;
wire n_5373;
wire n_5374;
wire n_5375;
wire n_5376;
wire n_5377;
wire n_5378;
wire n_5379;
wire n_5380;
wire n_5381;
wire n_5382;
wire n_5383;
wire n_5384;
wire n_5385;
wire n_5386;
wire n_5387;
wire n_5388;
wire n_5389;
wire n_5390;
wire n_5391;
wire n_5392;
wire n_5393;
wire n_5394;
wire n_5395;
wire n_5396;
wire n_5397;
wire n_5398;
wire n_5399;
wire n_5400;
wire n_5401;
wire n_5402;
wire n_5403;
wire n_5404;
wire n_5405;
wire n_5406;
wire n_5407;
wire n_5408;
wire n_5409;
wire n_5410;
wire n_5411;
wire n_5412;
wire n_5413;
wire n_5414;
wire n_5415;
wire n_5416;
wire n_5417;
wire n_5418;
wire n_5419;
wire n_5420;
wire n_5421;
wire n_5422;
wire n_5423;
wire n_5424;
wire n_5425;
wire n_5426;
wire n_5427;
wire n_5428;
wire n_5429;
wire n_5430;
wire n_5431;
wire n_5432;
wire n_5433;
wire n_5434;
wire n_5435;
wire n_5436;
wire n_5437;
wire n_5438;
wire n_5439;
wire n_5440;
wire n_5441;
wire n_5442;
wire n_5443;
wire n_5444;
wire n_5445;
wire n_5446;
wire n_5447;
wire n_5448;
wire n_5449;
wire n_5450;
wire n_5451;
wire n_5452;
wire n_5453;
wire n_5454;
wire n_5455;
wire n_5456;
wire n_5457;
wire n_5458;
wire n_5459;
wire n_5460;
wire n_5461;
wire n_5462;
wire n_5463;
wire n_5464;
wire n_5465;
wire n_5466;
wire n_5467;
wire n_5468;
wire n_5469;
wire n_5470;
wire n_5471;
wire n_5472;
wire n_5473;
wire n_5474;
wire n_5475;
wire n_5476;
wire n_5477;
wire n_5478;
wire n_5479;
wire n_5480;
wire n_5481;
wire n_5482;
wire n_5483;
wire n_5484;
wire n_5485;
wire n_5486;
wire n_5487;
wire n_5488;
wire n_5489;
wire n_5490;
wire n_5491;
wire n_5492;
wire n_5493;
wire n_5494;
wire n_5495;
wire n_5496;
wire n_5497;
wire n_5498;
wire n_5499;
wire n_5500;
wire n_5501;
wire n_5502;
wire n_5503;
wire n_5504;
wire n_5505;
wire n_5506;
wire n_5507;
wire n_5508;
wire n_5509;
wire n_5510;
wire n_5511;
wire n_5512;
wire n_5513;
wire n_5514;
wire n_5515;
wire n_5516;
wire n_5517;
wire n_5518;
wire n_5519;
wire n_5520;
wire n_5521;
wire n_5522;
wire n_5523;
wire n_5524;
wire n_5525;
wire n_5526;
wire n_5527;
wire n_5528;
wire n_5529;
wire n_5530;
wire n_5531;
wire n_5532;
wire n_5533;
wire n_5534;
wire n_5535;
wire n_5536;
wire n_5537;
wire n_5538;
wire n_5539;
wire n_5540;
wire n_5541;
wire n_5542;
wire n_5543;
wire n_5544;
wire n_5545;
wire n_5546;
wire n_5547;
wire n_5548;
wire n_5549;
wire n_5550;
wire n_5551;
wire n_5552;
wire n_5553;
wire n_5554;
wire n_5555;
wire n_5556;
wire n_5557;
wire n_5558;
wire n_5559;
wire n_5560;
wire n_5561;
wire n_5562;
wire n_5563;
wire n_5564;
wire n_5565;
wire n_5566;
wire n_5567;
wire n_5568;
wire n_5569;
wire n_5570;
wire n_5571;
wire n_5572;
wire n_5573;
wire n_5574;
wire n_5575;
wire n_5576;
wire n_5577;
wire n_5578;
wire n_5579;
wire n_5580;
wire n_5581;
wire n_5582;
wire n_5583;
wire n_5584;
wire n_5585;
wire n_5586;
wire n_5587;
wire n_5588;
wire n_5589;
wire n_5590;
wire n_5591;
wire n_5592;
wire n_5593;
wire n_5594;
wire n_5595;
wire n_5596;
wire n_5597;
wire n_5598;
wire n_5599;
wire n_5600;
wire n_5601;
wire n_5602;
wire n_5603;
wire n_5604;
wire n_5605;
wire n_5606;
wire n_5607;
wire n_5608;
wire n_5609;
wire n_5610;
wire n_5611;
wire n_5612;
wire n_5613;
wire n_5614;
wire n_5615;
wire n_5616;
wire n_5617;
wire n_5618;
wire n_5619;
wire n_5620;
wire n_5621;
wire n_5622;
wire n_5623;
wire n_5624;
wire n_5625;
wire n_5626;
wire n_5627;
wire n_5628;
wire n_5629;
wire n_5630;
wire n_5631;
wire n_5632;
wire n_5633;
wire n_5634;
wire n_5635;
wire n_5636;
wire n_5637;
wire n_5638;
wire n_5639;
wire n_5640;
wire n_5641;
wire n_5642;
wire n_5643;
wire n_5644;
wire n_5645;
wire n_5646;
wire n_5647;
wire n_5648;
wire n_5649;
wire n_5650;
wire n_5651;
wire n_5652;
wire n_5653;
wire n_5654;
wire n_5655;
wire n_5656;
wire n_5657;
wire n_5658;
wire n_5659;
wire n_5660;
wire n_5661;
wire n_5662;
wire n_5663;
wire n_5664;
wire n_5665;
wire n_5666;
wire n_5667;
wire n_5668;
wire n_5669;
wire n_5670;
wire n_5671;
wire n_5672;
wire n_5673;
wire n_5674;
wire n_5675;
wire n_5676;
wire n_5677;
wire n_5678;
wire n_5679;
wire n_5680;
wire n_5681;
wire n_5682;
wire n_5683;
wire n_5684;
wire n_5685;
wire n_5686;
wire n_5687;
wire n_5688;
wire n_5689;
wire n_5690;
wire n_5691;
wire n_5692;
wire n_5693;
wire n_5694;
wire n_5695;
wire n_5696;
wire n_5697;
wire n_5698;
wire n_5699;
wire n_5700;
wire n_5701;
wire n_5702;
wire n_5703;
wire n_5704;
wire n_5705;
wire n_5706;
wire n_5707;
wire n_5708;
wire n_5709;
wire n_5710;
wire n_5711;
wire n_5712;
wire n_5713;
wire n_5714;
wire n_5715;
wire n_5716;
wire n_5717;
wire n_5718;
wire n_5719;
wire n_5720;
wire n_5721;
wire n_5722;
wire n_5723;
wire n_5724;
wire n_5725;
wire n_5726;
wire n_5727;
wire n_5728;
wire n_5729;
wire n_5730;
wire n_5731;
wire n_5732;
wire n_5733;
wire n_5734;
wire n_5735;
wire n_5736;
wire n_5737;
wire n_5738;
wire n_5739;
wire n_5740;
wire n_5741;
wire n_5742;
wire n_5743;
wire n_5744;
wire n_5745;
wire n_5746;
wire n_5747;
wire n_5748;
wire n_5749;
wire n_5750;
wire n_5751;
wire n_5752;
wire n_5753;
wire n_5754;
wire n_5755;
wire n_5756;
wire n_5757;
wire n_5758;
wire n_5759;
wire n_5760;
wire n_5761;
wire n_5762;
wire n_5763;
wire n_5764;
wire n_5765;
wire n_5766;
wire n_5767;
wire n_5768;
wire n_5769;
wire n_5770;
wire n_5771;
wire n_5772;
wire n_5773;
wire n_5774;
wire n_5775;
wire n_5776;
wire n_5777;
wire n_5778;
wire n_5779;
wire n_5780;
wire n_5781;
wire n_5782;
wire n_5783;
wire n_5784;
wire n_5785;
wire n_5786;
wire n_5787;
wire n_5788;
wire n_5789;
wire n_5790;
wire n_5791;
wire n_5792;
wire n_5793;
wire n_5794;
wire n_5795;
wire n_5796;
wire n_5797;
wire n_5798;
wire n_5799;
wire n_5800;
wire n_5801;
wire n_5802;
wire n_5803;
wire n_5804;
wire n_5805;
wire n_5806;
wire n_5807;
wire n_5808;
wire n_5809;
wire n_5810;
wire n_5811;
wire n_5812;
wire n_5813;
wire n_5814;
wire n_5815;
wire n_5816;
wire n_5817;
wire n_5818;
wire n_5819;
wire n_5820;
wire n_5821;
wire n_5822;
wire n_5823;
wire n_5824;
wire n_5825;
wire n_5826;
wire n_5827;
wire n_5828;
wire n_5829;
wire n_5830;
wire n_5831;
wire n_5832;
wire n_5833;
wire n_5834;
wire n_5835;
wire n_5836;
wire n_5837;
wire n_5838;
wire n_5839;
wire n_5840;
wire n_5841;
wire n_5842;
wire n_5843;
wire n_5844;
wire n_5845;
wire n_5846;
wire n_5847;
wire n_5848;
wire n_5849;
wire n_5850;
wire n_5851;
wire n_5852;
wire n_5853;
wire n_5854;
wire n_5855;
wire n_5856;
wire n_5857;
wire n_5858;
wire n_5859;
wire n_5860;
wire n_5861;
wire n_5862;
wire n_5863;
wire n_5864;
wire n_5865;
wire n_5866;
wire n_5867;
wire n_5868;
wire n_5869;
wire n_5870;
wire n_5871;
wire n_5872;
wire n_5873;
wire n_5874;
wire n_5875;
wire n_5876;
wire n_5877;
wire n_5878;
wire n_5879;
wire n_5880;
wire n_5881;
wire n_5882;
wire n_5883;
wire n_5884;
wire n_5885;
wire n_5886;
wire n_5887;
wire n_5888;
wire n_5889;
wire n_5890;
wire n_5891;
wire n_5892;
wire n_5893;
wire n_5894;
wire n_5895;
wire n_5896;
wire n_5897;
wire n_5898;
wire n_5899;
wire n_5900;
wire n_5901;
wire n_5902;
wire n_5903;
wire n_5904;
wire n_5905;
wire n_5906;
wire n_5907;
wire n_5908;
wire n_5909;
wire n_5910;
wire n_5911;
wire n_5912;
wire n_5913;
wire n_5914;
wire n_5915;
wire n_5916;
wire n_5917;
wire n_5918;
wire n_5919;
wire n_5920;
wire n_5921;
wire n_5922;
wire n_5923;
wire n_5924;
wire n_5925;
wire n_5926;
wire n_5927;
wire n_5928;
wire n_5929;
wire n_5930;
wire n_5931;
wire n_5932;
wire n_5933;
wire n_5934;
wire n_5935;
wire n_5936;
wire n_5937;
wire n_5938;
wire n_5939;
wire n_5940;
wire n_5941;
wire n_5942;
wire n_5943;
wire n_5944;
wire n_5945;
wire n_5946;
wire n_5947;
wire n_5948;
wire n_5949;
wire n_5950;
wire n_5951;
wire n_5952;
wire n_5953;
wire n_5954;
wire n_5955;
wire n_5956;
wire n_5957;
wire n_5958;
wire n_5959;
wire n_5960;
wire n_5961;
wire n_5962;
wire n_5963;
wire n_5964;
wire n_5965;
wire n_5966;
wire n_5967;
wire n_5968;
wire n_5969;
wire n_5970;
wire n_5971;
wire n_5972;
wire n_5973;
wire n_5974;
wire n_5975;
wire n_5976;
wire n_5977;
wire n_5978;
wire n_5979;
wire n_5980;
wire n_5981;
wire n_5982;
wire n_5983;
wire n_5984;
wire n_5985;
wire n_5986;
wire n_5987;
wire n_5988;
wire n_5989;
wire n_5990;
wire n_5991;
wire n_5992;
wire n_5993;
wire n_5994;
wire n_5995;
wire n_5996;
wire n_5997;
wire n_5998;
wire n_5999;
wire n_6000;
wire n_6001;
wire n_6002;
wire n_6003;
wire n_6004;
wire n_6005;
wire n_6006;
wire n_6007;
wire n_6008;
wire n_6009;
wire n_6010;
wire n_6011;
wire n_6012;
wire n_6013;
wire n_6014;
wire n_6015;
wire n_6016;
wire n_6017;
wire n_6018;
wire n_6019;
wire n_6020;
wire n_6021;
wire n_6022;
wire n_6023;
wire n_6024;
wire n_6025;
wire n_6026;
wire n_6027;
wire n_6028;
wire n_6029;
wire n_6030;
wire n_6031;
wire n_6032;
wire n_6033;
wire n_6034;
wire n_6035;
wire n_6036;
wire n_6037;
wire n_6038;
wire n_6039;
wire n_6040;
wire n_6041;
wire n_6042;
wire n_6043;
wire n_6044;
wire n_6045;
wire n_6046;
wire n_6047;
wire n_6048;
wire n_6049;
wire n_6050;
wire n_6051;
wire n_6052;
wire n_6053;
wire n_6054;
wire n_6055;
wire n_6056;
wire n_6057;
wire n_6058;
wire n_6059;
wire n_6060;
wire n_6061;
wire n_6062;
wire n_6063;
wire n_6064;
wire n_6065;
wire n_6066;
wire n_6067;
wire n_6068;
wire n_6069;
wire n_6070;
wire n_6071;
wire n_6072;
wire n_6073;
wire n_6074;
wire n_6075;
wire n_6076;
wire n_6077;
wire n_6078;
wire n_6079;
wire n_6080;
wire n_6081;
wire n_6082;
wire n_6083;
wire n_6084;
wire n_6085;
wire n_6086;
wire n_6087;
wire n_6088;
wire n_6089;
wire n_6090;
wire n_6091;
wire n_6092;
wire n_6093;
wire n_6094;
wire n_6095;
wire n_6096;
wire n_6097;
wire n_6098;
wire n_6099;
wire n_6100;
wire n_6101;
wire n_6102;
wire n_6103;
wire n_6104;
wire n_6105;
wire n_6106;
wire n_6107;
wire n_6108;
wire n_6109;
wire n_6110;
wire n_6111;
wire n_6112;
wire n_6113;
wire n_6114;
wire n_6115;
wire n_6116;
wire n_6117;
wire n_6118;
wire n_6119;
wire n_6120;
wire n_6121;
wire n_6122;
wire n_6123;
wire n_6124;
wire n_6125;
wire n_6126;
wire n_6127;
wire n_6128;
wire n_6129;
wire n_6130;
wire n_6131;
wire n_6132;
wire n_6133;
wire n_6134;
wire n_6135;
wire n_6136;
wire n_6137;
wire n_6138;
wire n_6139;
wire n_6140;
wire n_6141;
wire n_6142;
wire n_6143;
wire n_6144;
wire n_6145;
wire n_6146;
wire n_6147;
wire n_6148;
wire n_6149;
wire n_6150;
wire n_6151;
wire n_6152;
wire n_6153;
wire n_6154;
wire n_6155;
wire n_6156;
wire n_6157;
wire n_6158;
wire n_6159;
wire n_6160;
wire n_6161;
wire n_6162;
wire n_6163;
wire n_6164;
wire n_6165;
wire n_6166;
wire n_6167;
wire n_6168;
wire n_6169;
wire n_6170;
wire n_6171;
wire n_6172;
wire n_6173;
wire n_6174;
wire n_6175;
wire n_6176;
wire n_6177;
wire n_6178;
wire n_6179;
wire n_6180;
wire n_6181;
wire n_6182;
wire n_6183;
wire n_6184;
wire n_6185;
wire n_6186;
wire n_6187;
wire n_6188;
wire n_6189;
wire n_6190;
wire n_6191;
wire n_6192;
wire n_6193;
wire n_6194;
wire n_6195;
wire n_6196;
wire n_6197;
wire n_6198;
wire n_6199;
wire n_6200;
wire n_6201;
wire n_6202;
wire n_6203;
wire n_6204;
wire n_6205;
wire n_6206;
wire n_6207;
wire n_6208;
wire n_6209;
wire n_6210;
wire n_6211;
wire n_6212;
wire n_6213;
wire n_6214;
wire n_6215;
wire n_6216;
wire n_6217;
wire n_6218;
wire n_6219;
wire n_6220;
wire n_6221;
wire n_6222;
wire n_6223;
wire n_6224;
wire n_6225;
wire n_6226;
wire n_6227;
wire n_6228;
wire n_6229;
wire n_6230;
wire n_6231;
wire n_6232;
wire n_6233;
wire n_6234;
wire n_6235;
wire n_6236;
wire n_6237;
wire n_6238;
wire n_6239;
wire n_6240;
wire n_6241;
wire n_6242;
wire n_6243;
wire n_6244;
wire n_6245;
wire n_6246;
wire n_6247;
wire n_6248;
wire n_6249;
wire n_6250;
wire n_6251;
wire n_6252;
wire n_6253;
wire n_6254;
wire n_6255;
wire n_6256;
wire n_6257;
wire n_6258;
wire n_6259;
wire n_6260;
wire n_6261;
wire n_6262;
wire n_6263;
wire n_6264;
wire n_6265;
wire n_6266;
wire n_6267;
wire n_6268;
wire n_6269;
wire n_6270;
wire n_6271;
wire n_6272;
wire n_6273;
wire n_6274;
wire n_6275;
wire n_6276;
wire n_6277;
wire n_6278;
wire n_6279;
wire n_6280;
wire n_6281;
wire n_6282;
wire n_6283;
wire n_6284;
wire n_6285;
wire n_6286;
wire n_6287;
wire n_6288;
wire n_6289;
wire n_6290;
wire n_6291;
wire n_6292;
wire n_6293;
wire n_6294;
wire n_6295;
wire n_6296;
wire n_6297;
wire n_6298;
wire n_6299;
wire n_6300;
wire n_6301;
wire n_6302;
wire n_6303;
wire n_6304;
wire n_6305;
wire n_6306;
wire n_6307;
wire n_6308;
wire n_6309;
wire n_6310;
wire n_6311;
wire n_6312;
wire n_6313;
wire n_6314;
wire n_6315;
wire n_6316;
wire n_6317;
wire n_6318;
wire n_6319;
wire n_6320;
wire n_6321;
wire n_6322;
wire n_6323;
wire n_6324;
wire n_6325;
wire n_6326;
wire n_6327;
wire n_6328;
wire n_6329;
wire n_6330;
wire n_6331;
wire n_6332;
wire n_6333;
wire n_6334;
wire n_6335;
wire n_6336;
wire n_6337;
wire n_6338;
wire n_6339;
wire n_6340;
wire n_6341;
wire n_6342;
wire n_6343;
wire n_6344;
wire n_6345;
wire n_6346;
wire n_6347;
wire n_6348;
wire n_6349;
wire n_6350;
wire n_6351;
wire n_6352;
wire n_6353;
wire n_6354;
wire n_6355;
wire n_6356;
wire n_6357;
wire n_6358;
wire n_6359;
wire n_6360;
wire n_6361;
wire n_6362;
wire n_6363;
wire n_6364;
wire n_6365;
wire n_6366;
wire n_6367;
wire n_6368;
wire n_6369;
wire n_6370;
wire n_6371;
wire n_6372;
wire n_6373;
wire n_6374;
wire n_6375;
wire n_6376;
wire n_6377;
wire n_6378;
wire n_6379;
wire n_6380;
wire n_6381;
wire n_6382;
wire n_6383;
wire n_6384;
wire n_6385;
wire n_6386;
wire n_6387;
wire n_6388;
wire n_6389;
wire n_6390;
wire n_6391;
wire n_6392;
wire n_6393;
wire n_6394;
wire n_6395;
wire n_6396;
wire n_6397;
wire n_6398;
wire n_6399;
wire n_6400;
wire n_6401;
wire n_6402;
wire n_6403;
wire n_6404;
wire n_6405;
wire n_6406;
wire n_6407;
wire n_6408;
wire n_6409;
wire n_6410;
wire n_6411;
wire n_6412;
wire n_6413;
wire n_6414;
wire n_6415;
wire n_6416;
wire n_6417;
wire n_6418;
wire n_6419;
wire n_6420;
wire n_6421;
wire n_6422;
wire n_6423;
wire n_6424;
wire n_6425;
wire n_6426;
wire n_6427;
wire n_6428;
wire n_6429;
wire n_6430;
wire n_6431;
wire n_6432;
wire n_6433;
wire n_6434;
wire n_6435;
wire n_6436;
wire n_6437;
wire n_6438;
wire n_6439;
wire n_6440;
wire n_6441;
wire n_6442;
wire n_6443;
wire n_6444;
wire n_6445;
wire n_6446;
wire n_6447;
wire n_6448;
wire n_6449;
wire n_6450;
wire n_6451;
wire n_6452;
wire n_6453;
wire n_6454;
wire n_6455;
wire n_6456;
wire n_6457;
wire n_6458;
wire n_6459;
wire n_6460;
wire n_6461;
wire n_6462;
wire n_6463;
wire n_6464;
wire n_6465;
wire n_6466;
wire n_6467;
wire n_6468;
wire n_6469;
wire n_6470;
wire n_6471;
wire n_6472;
wire n_6473;
wire n_6474;
wire n_6475;
wire n_6476;
wire n_6477;
wire n_6478;
wire n_6479;
wire n_6480;
wire n_6481;
wire n_6482;
wire n_6483;
wire n_6484;
wire n_6485;
wire n_6486;
wire n_6487;
wire n_6488;
wire n_6489;
wire n_6490;
wire n_6491;
wire n_6492;
wire n_6493;
wire n_6494;
wire n_6495;
wire n_6496;
wire n_6497;
wire n_6498;
wire n_6499;
wire n_6500;
wire n_6501;
wire n_6502;
wire n_6503;
wire n_6504;
wire n_6505;
wire n_6506;
wire n_6507;
wire n_6508;
wire n_6509;
wire n_6510;
wire n_6511;
wire n_6512;
wire n_6513;
wire n_6514;
wire n_6515;
wire n_6516;
wire n_6517;
wire n_6518;
wire n_6519;
wire n_6520;
wire n_6521;
wire n_6522;
wire n_6523;
wire n_6524;
wire n_6525;
wire n_6526;
wire n_6527;
wire n_6528;
wire n_6529;
wire n_6530;
wire n_6531;
wire n_6532;
wire n_6533;
wire n_6534;
wire n_6535;
wire n_6536;
wire n_6537;
wire n_6538;
wire n_6539;
wire n_6540;
wire n_6541;
wire n_6542;
wire n_6543;
wire n_6544;
wire n_6545;
wire n_6546;
wire n_6547;
wire n_6548;
wire n_6549;
wire n_6550;
wire n_6551;
wire n_6552;
wire n_6553;
wire n_6554;
wire n_6555;
wire n_6556;
wire n_6557;
wire n_6558;
wire n_6559;
wire n_6560;
wire n_6561;
wire n_6562;
wire n_6563;
wire n_6564;
wire n_6565;
wire n_6566;
wire n_6567;
wire n_6568;
wire n_6569;
wire n_6570;
wire n_6571;
wire n_6572;
wire n_6573;
wire n_6574;
wire n_6575;
wire n_6576;
wire n_6577;
wire n_6578;
wire n_6579;
wire n_6580;
wire n_6581;
wire n_6582;
wire n_6583;
wire n_6584;
wire n_6585;
wire n_6586;
wire n_6587;
wire n_6588;
wire n_6589;
wire n_6590;
wire n_6591;
wire n_6592;
wire n_6593;
wire n_6594;
wire n_6595;
wire n_6596;
wire n_6597;
wire n_6598;
wire n_6599;
wire n_6600;
wire n_6601;
wire n_6602;
wire n_6603;
wire n_6604;
wire n_6605;
wire n_6606;
wire n_6607;
wire n_6608;
wire n_6609;
wire n_6610;
wire n_6611;
wire n_6612;
wire n_6613;
wire n_6614;
wire n_6615;
wire n_6616;
wire n_6617;
wire n_6618;
wire n_6619;
wire n_6620;
wire n_6621;
wire n_6622;
wire n_6623;
wire n_6624;
wire n_6625;
wire n_6626;
wire n_6627;
wire n_6628;
wire n_6629;
wire n_6630;
wire n_6631;
wire n_6632;
wire n_6633;
wire n_6634;
wire n_6635;
wire n_6636;
wire n_6637;
wire n_6638;
wire n_6639;
wire n_6640;
wire n_6641;
wire n_6642;
wire n_6643;
wire n_6644;
wire n_6645;
wire n_6646;
wire n_6647;
wire n_6648;
wire n_6649;
wire n_6650;
wire n_6651;
wire n_6652;
wire n_6653;
wire n_6654;
wire n_6655;
wire n_6656;
wire n_6657;
wire n_6658;
wire n_6659;
wire n_6660;
wire n_6661;
wire n_6662;
wire n_6663;
wire n_6664;
wire n_6665;
wire n_6666;
wire n_6667;
wire n_6668;
wire n_6669;
wire n_6670;
wire n_6671;
wire n_6672;
wire n_6673;
wire n_6674;
wire n_6675;
wire n_6676;
wire n_6677;
wire n_6678;
wire n_6679;
wire n_6680;
wire n_6681;
wire n_6682;
wire n_6683;
wire n_6684;
wire n_6685;
wire n_6686;
wire n_6687;
wire n_6688;
wire n_6689;
wire n_6690;
wire n_6691;
wire n_6692;
wire n_6693;
wire n_6694;
wire n_6695;
wire n_6696;
wire n_6697;
wire n_6698;
wire n_6699;
wire n_6700;
wire n_6701;
wire n_6702;
wire n_6703;
wire n_6704;
wire n_6705;
wire n_6706;
wire n_6707;
wire n_6708;
wire n_6709;
wire n_6710;
wire n_6711;
wire n_6712;
wire n_6713;
wire n_6714;
wire n_6715;
wire n_6716;
wire n_6717;
wire n_6718;
wire n_6719;
wire n_6720;
wire n_6721;
wire n_6722;
wire n_6723;
wire n_6724;
wire n_6725;
wire n_6726;
wire n_6727;
wire n_6728;
wire n_6729;
wire n_6730;
wire n_6731;
wire n_6732;
wire n_6733;
wire n_6734;
wire n_6735;
wire n_6736;
wire n_6737;
wire n_6738;
wire n_6739;
wire n_6740;
wire n_6741;
wire n_6742;
wire n_6743;
wire n_6744;
wire n_6745;
wire n_6746;
wire n_6747;
wire n_6748;
wire n_6749;
wire n_6750;
wire n_6751;
wire n_6752;
wire n_6753;
wire n_6754;
wire n_6755;
wire n_6756;
wire n_6757;
wire n_6758;
wire n_6759;
wire n_6760;
wire n_6761;
wire n_6762;
wire n_6763;
wire n_6764;
wire n_6765;
wire n_6766;
wire n_6767;
wire n_6768;
wire n_6769;
wire n_6770;
wire n_6771;
wire n_6772;
wire n_6773;
wire n_6774;
wire n_6775;
wire n_6776;
wire n_6777;
wire n_6778;
wire n_6779;
wire n_6780;
wire n_6781;
wire n_6782;
wire n_6783;
wire n_6784;
wire n_6785;
wire n_6786;
wire n_6787;
wire n_6788;
wire n_6789;
wire n_6790;
wire n_6791;
wire n_6792;
wire n_6793;
wire n_6794;
wire n_6795;
wire n_6796;
wire n_6797;
wire n_6798;
wire n_6799;
wire n_6800;
wire n_6801;
wire n_6802;
wire n_6803;
wire n_6804;
wire n_6805;
wire n_6806;
wire n_6807;
wire n_6808;
wire n_6809;
wire n_6810;
wire n_6811;
wire n_6812;
wire n_6813;
wire n_6814;
wire n_6815;
wire n_6816;
wire n_6817;
wire n_6818;
wire n_6819;
wire n_6820;
wire n_6821;
wire n_6822;
wire n_6823;
wire n_6824;
wire n_6825;
wire n_6826;
wire n_6827;
wire n_6828;
wire n_6829;
wire n_6830;
wire n_6831;
wire n_6832;
wire n_6833;
wire n_6834;
wire n_6835;
wire n_6836;
wire n_6837;
wire n_6838;
wire n_6839;
wire n_6840;
wire n_6841;
wire n_6842;
wire n_6843;
wire n_6844;
wire n_6845;
wire n_6846;
wire n_6847;
wire n_6848;
wire n_6849;
wire n_6850;
wire n_6851;
wire n_6852;
wire n_6853;
wire n_6854;
wire n_6855;
wire n_6856;
wire n_6857;
wire n_6858;
wire n_6859;
wire n_6860;
wire n_6861;
wire n_6862;
wire n_6863;
wire n_6864;
wire n_6865;
wire n_6866;
wire n_6867;
wire n_6868;
wire n_6869;
wire n_6870;
wire n_6871;
wire n_6872;
wire n_6873;
wire n_6874;
wire n_6875;
wire n_6876;
wire n_6877;
wire n_6878;
wire n_6879;
wire n_6880;
wire n_6881;
wire n_6882;
wire n_6883;
wire n_6884;
wire n_6885;
wire n_6886;
wire n_6887;
wire n_6888;
wire n_6889;
wire n_6890;
wire n_6891;
wire n_6892;
wire n_6893;
wire n_6894;
wire n_6895;
wire n_6896;
wire n_6897;
wire n_6898;
wire n_6899;
wire n_6900;
wire n_6901;
wire n_6902;
wire n_6903;
wire n_6904;
wire n_6905;
wire n_6906;
wire n_6907;
wire n_6908;
wire n_6909;
wire n_6910;
wire n_6911;
wire n_6912;
wire n_6913;
wire n_6914;
wire n_6915;
wire n_6916;
wire n_6917;
wire n_6918;
wire n_6919;
wire n_6920;
wire n_6921;
wire n_6922;
wire n_6923;
wire n_6924;
wire n_6925;
wire n_6926;
wire n_6927;
wire n_6928;
wire n_6929;
wire n_6930;
wire n_6931;
wire n_6932;
wire n_6933;
wire n_6934;
wire n_6935;
wire n_6936;
wire n_6937;
wire n_6938;
wire n_6939;
wire n_6940;
wire n_6941;
wire n_6942;
wire n_6943;
wire n_6944;
wire n_6945;
wire n_6946;
wire n_6947;
wire n_6948;
wire n_6949;
wire n_6950;
wire n_6951;
wire n_6952;
wire n_6953;
wire n_6954;
wire n_6955;
wire n_6956;
wire n_6957;
wire n_6958;
wire n_6959;
wire n_6960;
wire n_6961;
wire n_6962;
wire n_6963;
wire n_6964;
wire n_6965;
wire n_6966;
wire n_6967;
wire n_6968;
wire n_6969;
wire n_6970;
wire n_6971;
wire n_6972;
wire n_6973;
wire n_6974;
wire n_6975;
wire n_6976;
wire n_6977;
wire n_6978;
wire n_6979;
wire n_6980;
wire n_6981;
wire n_6982;
wire n_6983;
wire n_6984;
wire n_6985;
wire n_6986;
wire n_6987;
wire n_6988;
wire n_6989;
wire n_6990;
wire n_6991;
wire n_6992;
wire n_6993;
wire n_6994;
wire n_6995;
wire n_6996;
wire n_6997;
wire n_6998;
wire n_6999;
wire n_7000;
wire n_7001;
wire n_7002;
wire n_7003;
wire n_7004;
wire n_7005;
wire n_7006;
wire n_7007;
wire n_7008;
wire n_7009;
wire n_7010;
wire n_7011;
wire n_7012;
wire n_7013;
wire n_7014;
wire n_7015;
wire n_7016;
wire n_7017;
wire n_7018;
wire n_7019;
wire n_7020;
wire n_7021;
wire n_7022;
wire n_7023;
wire n_7024;
wire n_7025;
wire n_7026;
wire n_7027;
wire n_7028;
wire n_7029;
wire n_7030;
wire n_7031;
wire n_7032;
wire n_7033;
wire n_7034;
wire n_7035;
wire n_7036;
wire n_7037;
wire n_7038;
wire n_7039;
wire n_7040;
wire n_7041;
wire n_7042;
wire n_7043;
wire n_7044;
wire n_7045;
wire n_7046;
wire n_7047;
wire n_7048;
wire n_7049;
wire n_7050;
wire n_7051;
wire n_7052;
wire n_7053;
wire n_7054;
wire n_7055;
wire n_7056;
wire n_7057;
wire n_7058;
wire n_7059;
wire n_7060;
wire n_7061;
wire n_7062;
wire n_7063;
wire n_7064;
wire n_7065;
wire n_7066;
wire n_7067;
wire n_7068;
wire n_7069;
wire n_7070;
wire n_7071;
wire n_7072;
wire n_7073;
wire n_7074;
wire n_7075;
wire n_7076;
wire n_7077;
wire n_7078;
wire n_7079;
wire n_7080;
wire n_7081;
wire n_7082;
wire n_7083;
wire n_7084;
wire n_7085;
wire n_7086;
wire n_7087;
wire n_7088;
wire n_7089;
wire n_7090;
wire n_7091;
wire n_7092;
wire n_7093;
wire n_7094;
wire n_7095;
wire n_7096;
wire n_7097;
wire n_7098;
wire n_7099;
wire n_7100;
wire n_7101;
wire n_7102;
wire n_7103;
wire n_7104;
wire n_7105;
wire n_7106;
wire n_7107;
wire n_7108;
wire n_7109;
wire n_7110;
wire n_7111;
wire n_7112;
wire n_7113;
wire n_7114;
wire n_7115;
wire n_7116;
wire n_7117;
wire n_7118;
wire n_7119;
wire n_7120;
wire n_7121;
wire n_7122;
wire n_7123;
wire n_7124;
wire n_7125;
wire n_7126;
wire n_7127;
wire n_7128;
wire n_7129;
wire n_7130;
wire n_7131;
wire n_7132;
wire n_7133;
wire n_7134;
wire n_7135;
wire n_7136;
wire n_7137;
wire n_7138;
wire n_7139;
wire n_7140;
wire n_7141;
wire n_7142;
wire n_7143;
wire n_7144;
wire n_7145;
wire n_7146;
wire n_7147;
wire n_7148;
wire n_7149;
wire n_7150;
wire n_7151;
wire n_7152;
wire n_7153;
wire n_7154;
wire n_7155;
wire n_7156;
wire n_7157;
wire n_7158;
wire n_7159;
wire n_7160;
wire n_7161;
wire n_7162;
wire n_7163;
wire n_7164;
wire n_7165;
wire n_7166;
wire n_7167;
wire n_7168;
wire n_7169;
wire n_7170;
wire n_7171;
wire n_7172;
wire n_7173;
wire n_7174;
wire n_7175;
wire n_7176;
wire n_7177;
wire n_7178;
wire n_7179;
wire n_7180;
wire n_7181;
wire n_7182;
wire n_7183;
wire n_7184;
wire n_7185;
wire n_7186;
wire n_7187;
wire n_7188;
wire n_7189;
wire n_7190;
wire n_7191;
wire n_7192;
wire n_7193;
wire n_7194;
wire n_7195;
wire n_7196;
wire n_7197;
wire n_7198;
wire n_7199;
wire n_7200;
wire n_7201;
wire n_7202;
wire n_7203;
wire n_7204;
wire n_7205;
wire n_7206;
wire n_7207;
wire n_7208;
wire n_7209;
wire n_7210;
wire n_7211;
wire n_7212;
wire n_7213;
wire n_7214;
wire n_7215;
wire n_7216;
wire n_7217;
wire n_7218;
wire n_7219;
wire n_7220;
wire n_7221;
wire n_7222;
wire n_7223;
wire n_7224;
wire n_7225;
wire n_7226;
wire n_7227;
wire n_7228;
wire n_7229;
wire n_7230;
wire n_7231;
wire n_7232;
wire n_7233;
wire n_7234;
wire n_7235;
wire n_7236;
wire n_7237;
wire n_7238;
wire n_7239;
wire n_7240;
wire n_7241;
wire n_7242;
wire n_7243;
wire n_7244;
wire n_7245;
wire n_7246;
wire n_7247;
wire n_7248;
wire n_7249;
wire n_7250;
wire n_7251;
wire n_7252;
wire n_7253;
wire n_7254;
wire n_7255;
wire n_7256;
wire n_7257;
wire n_7258;
wire n_7259;
wire n_7260;
wire n_7261;
wire n_7262;
wire n_7263;
wire n_7264;
wire n_7265;
wire n_7266;
wire n_7267;
wire n_7268;
wire n_7269;
wire n_7270;
wire n_7271;
wire n_7272;
wire n_7273;
wire n_7274;
wire n_7275;
wire n_7276;
wire n_7277;
wire n_7278;
wire n_7279;
wire n_7280;
wire n_7281;
wire n_7282;
wire n_7283;
wire n_7284;
wire n_7285;
wire n_7286;
wire n_7287;
wire n_7288;
wire n_7289;
wire n_7290;
wire n_7291;
wire n_7292;
wire n_7293;
wire n_7294;
wire n_7295;
wire n_7296;
wire n_7297;
wire n_7298;
wire n_7299;
wire n_7300;
wire n_7301;
wire n_7302;
wire n_7303;
wire n_7304;
wire n_7305;
wire n_7306;
wire n_7307;
wire n_7308;
wire n_7309;
wire n_7310;
wire n_7311;
wire n_7312;
wire n_7313;
wire n_7314;
wire n_7315;
wire n_7316;
wire n_7317;
wire n_7318;
wire n_7319;
wire n_7320;
wire n_7321;
wire n_7322;
wire n_7323;
wire n_7324;
wire n_7325;
wire n_7326;
wire n_7327;
wire n_7328;
wire n_7329;
wire n_7330;
wire n_7331;
wire n_7332;
wire n_7333;
wire n_7334;
wire n_7335;
wire n_7336;
wire n_7337;
wire n_7338;
wire n_7339;
wire n_7340;
wire n_7341;
wire n_7342;
wire n_7343;
wire n_7344;
wire n_7345;
wire n_7346;
wire n_7347;
wire n_7348;
wire n_7349;
wire n_7350;
wire n_7351;
wire n_7352;
wire n_7353;
wire n_7354;
wire n_7355;
wire n_7356;
wire n_7357;
wire n_7358;
wire n_7359;
wire n_7360;
wire n_7361;
wire n_7362;
wire n_7363;
wire n_7364;
wire n_7365;
wire n_7366;
wire n_7367;
wire n_7368;
wire n_7369;
wire n_7370;
wire n_7371;
wire n_7372;
wire n_7373;
wire n_7374;
wire n_7375;
wire n_7376;
wire n_7377;
wire n_7378;
wire n_7379;
wire n_7380;
wire n_7381;
wire n_7382;
wire n_7383;
wire n_7384;
wire n_7385;
wire n_7386;
wire n_7387;
wire n_7388;
wire n_7389;
wire n_7390;
wire n_7391;
wire n_7392;
wire n_7393;
wire n_7394;
wire n_7395;
wire n_7396;
wire n_7397;
wire n_7398;
wire n_7399;
wire n_7400;
wire n_7401;
wire n_7402;
wire n_7403;
wire n_7404;
wire n_7405;
wire n_7406;
wire n_7407;
wire n_7408;
wire n_7409;
wire n_7410;
wire n_7411;
wire n_7412;
wire n_7413;
wire n_7414;
wire n_7415;
wire n_7416;
wire n_7417;
wire n_7418;
wire n_7419;
wire n_7420;
wire n_7421;
wire n_7422;
wire n_7423;
wire n_7424;
wire n_7425;
wire n_7426;
wire n_7427;
wire n_7428;
wire n_7429;
wire n_7430;
wire n_7431;
wire n_7432;
wire n_7433;
wire n_7434;
wire n_7435;
wire n_7436;
wire n_7437;
wire n_7438;
wire n_7439;
wire n_7440;
wire n_7441;
wire n_7442;
wire n_7443;
wire n_7444;
wire n_7445;
wire n_7446;
wire n_7447;
wire n_7448;
wire n_7449;
wire n_7450;
wire n_7451;
wire n_7452;
wire n_7453;
wire n_7454;
wire n_7455;
wire n_7456;
wire n_7457;
wire n_7458;
wire n_7459;
wire n_7460;
wire n_7461;
wire n_7462;
wire n_7463;
wire n_7464;
wire n_7465;
wire n_7466;
wire n_7467;
wire n_7468;
wire n_7469;
wire n_7470;
wire n_7471;
wire n_7472;
wire n_7473;
wire n_7474;
wire n_7475;
wire n_7476;
wire n_7477;
wire n_7478;
wire n_7479;
wire n_7480;
wire n_7481;
wire n_7482;
wire n_7483;
wire n_7484;
wire n_7485;
wire n_7486;
wire n_7487;
wire n_7488;
wire n_7489;
wire n_7490;
wire n_7491;
wire n_7492;
wire n_7493;
wire n_7494;
wire n_7495;
wire n_7496;
wire n_7497;
wire n_7498;
wire n_7499;
wire n_7500;
wire n_7501;
wire n_7502;
wire n_7503;
wire n_7504;
wire n_7505;
wire n_7506;
wire n_7507;
wire n_7508;
wire n_7509;
wire n_7510;
wire n_7511;
wire n_7512;
wire n_7513;
wire n_7514;
wire n_7515;
wire n_7516;
wire n_7517;
wire n_7518;
wire n_7519;
wire n_7520;
wire n_7521;
wire n_7522;
wire n_7523;
wire n_7524;
wire n_7525;
wire n_7526;
wire n_7527;
wire n_7528;
wire n_7529;
wire n_7530;
wire n_7531;
wire n_7532;
wire n_7533;
wire n_7534;
wire n_7535;
wire n_7536;
wire n_7537;
wire n_7538;
wire n_7539;
wire n_7540;
wire n_7541;
wire n_7542;
wire n_7543;
wire n_7544;
wire n_7545;
wire n_7546;
wire n_7547;
wire n_7548;
wire n_7549;
wire n_7550;
wire n_7551;
wire n_7552;
wire n_7553;
wire n_7554;
wire n_7555;
wire n_7556;
wire n_7557;
wire n_7558;
wire n_7559;
wire n_7560;
wire n_7561;
wire n_7562;
wire n_7563;
wire n_7564;
wire n_7565;
wire n_7566;
wire n_7567;
wire n_7568;
wire n_7569;
wire n_7570;
wire n_7571;
wire n_7572;
wire n_7573;
wire n_7574;
wire n_7575;
wire n_7576;
wire n_7577;
wire n_7578;
wire n_7579;
wire n_7580;
wire n_7581;
wire n_7582;
wire n_7583;
wire n_7584;
wire n_7585;
wire n_7586;
wire n_7587;
wire n_7588;
wire n_7589;
wire n_7590;
wire n_7591;
wire n_7592;
wire n_7593;
wire n_7594;
wire n_7595;
wire n_7596;
wire n_7597;
wire n_7598;
wire n_7599;
wire n_7600;
wire n_7601;
wire n_7602;
wire n_7603;
wire n_7604;
wire n_7605;
wire n_7606;
wire n_7607;
wire n_7608;
wire n_7609;
wire n_7610;
wire n_7611;
wire n_7612;
wire n_7613;
wire n_7614;
wire n_7615;
wire n_7616;
wire n_7617;
wire n_7618;
wire n_7619;
wire n_7620;
wire n_7621;
wire n_7622;
wire n_7623;
wire n_7624;
wire n_7625;
wire n_7626;
wire n_7627;
wire n_7628;
wire n_7629;
wire n_7630;
wire n_7631;
wire n_7632;
wire n_7633;
wire n_7634;
wire n_7635;
wire n_7636;
wire n_7637;
wire n_7638;
wire n_7639;
wire n_7640;
wire n_7641;
wire n_7642;
wire n_7643;
wire n_7644;
wire n_7645;
wire n_7646;
wire n_7647;
wire n_7648;
wire n_7649;
wire n_7650;
wire n_7651;
wire n_7652;
wire n_7653;
wire n_7654;
wire n_7655;
wire n_7656;
wire n_7657;
wire n_7658;
wire n_7659;
wire n_7660;
wire n_7661;
wire n_7662;
wire n_7663;
wire n_7664;
wire n_7665;
wire n_7666;
wire n_7667;
wire n_7668;
wire n_7669;
wire n_7670;
wire n_7671;
wire n_7672;
wire n_7673;
wire n_7674;
wire n_7675;
wire n_7676;
wire n_7677;
wire n_7678;
wire n_7679;
wire n_7680;
wire n_7681;
wire n_7682;
wire n_7683;
wire n_7684;
wire n_7685;
wire n_7686;
wire n_7687;
wire n_7688;
wire n_7689;
wire n_7690;
wire n_7691;
wire n_7692;
wire n_7693;
wire n_7694;
wire n_7695;
wire n_7696;
wire n_7697;
wire n_7698;
wire n_7699;
wire n_7700;
wire n_7701;
wire n_7702;
wire n_7703;
wire n_7704;
wire n_7705;
wire n_7706;
wire n_7707;
wire n_7708;
wire n_7709;
wire n_7710;
wire n_7711;
wire n_7712;
wire n_7713;
wire n_7714;
wire n_7715;
wire n_7716;
wire n_7717;
wire n_7718;
wire n_7719;
wire n_7720;
wire n_7721;
wire n_7722;
wire n_7723;
wire n_7724;
wire n_7725;
wire n_7726;
wire n_7727;
wire n_7728;
wire n_7729;
wire n_7730;
wire n_7731;
wire n_7732;
wire n_7733;
wire n_7734;
wire n_7735;
wire n_7736;
wire n_7737;
wire n_7738;
wire n_7739;
wire n_7740;
wire n_7741;
wire n_7742;
wire n_7743;
wire n_7744;
wire n_7745;
wire n_7746;
wire n_7747;
wire n_7748;
wire n_7749;
wire n_7750;
wire n_7751;
wire n_7752;
wire n_7753;
wire n_7754;
wire n_7755;
wire n_7756;
wire n_7757;
wire n_7758;
wire n_7759;
wire n_7760;
wire n_7761;
wire n_7762;
wire n_7763;
wire n_7764;
wire n_7765;
wire n_7766;
wire n_7767;
wire n_7768;
wire n_7769;
wire n_7770;
wire n_7771;
wire n_7772;
wire n_7773;
wire n_7774;
wire n_7775;
wire n_7776;
wire n_7777;
wire n_7778;
wire n_7779;
wire n_7780;
wire n_7781;
wire n_7782;
wire n_7783;
wire n_7784;
wire n_7785;
wire n_7786;
wire n_7787;
wire n_7788;
wire n_7789;
wire n_7790;
wire n_7791;
wire n_7792;
wire n_7793;
wire n_7794;
wire n_7795;
wire n_7796;
wire n_7797;
wire n_7798;
wire n_7799;
wire n_7800;
wire n_7801;
wire n_7802;
wire n_7803;
wire n_7804;
wire n_7805;
wire n_7806;
wire n_7807;
wire n_7808;
wire n_7809;
wire n_7810;
wire n_7811;
wire n_7812;
wire n_7813;
wire n_7814;
wire n_7815;
wire n_7816;
wire n_7817;
wire n_7818;
wire n_7819;
wire n_7820;
wire n_7821;
wire n_7822;
wire n_7823;
wire n_7824;
wire n_7825;
wire n_7826;
wire n_7827;
wire n_7828;
wire n_7829;
wire n_7830;
wire n_7831;
wire n_7832;
wire n_7833;
wire n_7834;
wire n_7835;
wire n_7836;
wire n_7837;
wire n_7838;
wire n_7839;
wire n_7840;
wire n_7841;
wire n_7842;
wire n_7843;
wire n_7844;
wire n_7845;
wire n_7846;
wire n_7847;
wire n_7848;
wire n_7849;
wire n_7850;
wire n_7851;
wire n_7852;
wire n_7853;
wire n_7854;
wire n_7855;
wire n_7856;
wire n_7857;
wire n_7858;
wire n_7859;
wire n_7860;
wire n_7861;
wire n_7862;
wire n_7863;
wire n_7864;
wire n_7865;
wire n_7866;
wire n_7867;
wire n_7868;
wire n_7869;
wire n_7870;
wire n_7871;
wire n_7872;
wire n_7873;
wire n_7874;
wire n_7875;
wire n_7876;
wire n_7877;
wire n_7878;
wire n_7879;
wire n_7880;
wire n_7881;
wire n_7882;
wire n_7883;
wire n_7884;
wire n_7885;
wire n_7886;
wire n_7887;
wire n_7888;
wire n_7889;
wire n_7890;
wire n_7891;
wire n_7892;
wire n_7893;
wire n_7894;
wire n_7895;
wire n_7896;
wire n_7897;
wire n_7898;
wire n_7899;
wire n_7900;
wire n_7901;
wire n_7902;
wire n_7903;
wire n_7904;
wire n_7905;
wire n_7906;
wire n_7907;
wire n_7908;
wire n_7909;
wire n_7910;
wire n_7911;
wire n_7912;
wire n_7913;
wire n_7914;
wire n_7915;
wire n_7916;
wire n_7917;
wire n_7918;
wire n_7919;
wire n_7920;
wire n_7921;
wire n_7922;
wire n_7923;
wire n_7924;
wire n_7925;
wire n_7926;
wire n_7927;
wire n_7928;
wire n_7929;
wire n_7930;
wire n_7931;
wire n_7932;
wire n_7933;
wire n_7934;
wire n_7935;
wire n_7936;
wire n_7937;
wire n_7938;
wire n_7939;
wire n_7940;
wire n_7941;
wire n_7942;
wire n_7943;
wire n_7944;
wire n_7945;
wire n_7946;
wire n_7947;
wire n_7948;
wire n_7949;
wire n_7950;
wire n_7951;
wire n_7952;
wire n_7953;
wire n_7954;
wire n_7955;
wire n_7956;
wire n_7957;
wire n_7958;
wire n_7959;
wire n_7960;
wire n_7961;
wire n_7962;
wire n_7963;
wire n_7964;
wire n_7965;
wire n_7966;
wire n_7967;
wire n_7968;
wire n_7969;
wire n_7970;
wire n_7971;
wire n_7972;
wire n_7973;
wire n_7974;
wire n_7975;
wire n_7976;
wire n_7977;
wire n_7978;
wire n_7979;
wire n_7980;
wire n_7981;
wire n_7982;
wire n_7983;
wire n_7984;
wire n_7985;
wire n_7986;
wire n_7987;
wire n_7988;
wire n_7989;
wire n_7990;
wire n_7991;
wire n_7992;
wire n_7993;
wire n_7994;
wire n_7995;
wire n_7996;
wire n_7997;
wire n_7998;
wire n_7999;
wire n_8000;
wire n_8001;
wire n_8002;
wire n_8003;
wire n_8004;
wire n_8005;
wire n_8006;
wire n_8007;
wire n_8008;
wire n_8009;
wire n_8010;
wire n_8011;
wire n_8012;
wire n_8013;
wire n_8014;
wire n_8015;
wire n_8016;
wire n_8017;
wire n_8018;
wire n_8019;
wire n_8020;
wire n_8021;
wire n_8022;
wire n_8023;
wire n_8024;
wire n_8025;
wire n_8026;
wire n_8027;
wire n_8028;
wire n_8029;
wire n_8030;
wire n_8031;
wire n_8032;
wire n_8033;
wire n_8034;
wire n_8035;
wire n_8036;
wire n_8037;
wire n_8038;
wire n_8039;
wire n_8040;
wire n_8041;
wire n_8042;
wire n_8043;
wire n_8044;
wire n_8045;
wire n_8046;
wire n_8047;
wire n_8048;
wire n_8049;
wire n_8050;
wire n_8051;
wire n_8052;
wire n_8053;
wire n_8054;
wire n_8055;
wire n_8056;
wire n_8057;
wire n_8058;
wire n_8059;
wire n_8060;
wire n_8061;
wire n_8062;
wire n_8063;
wire n_8064;
wire n_8065;
wire n_8066;
wire n_8067;
wire n_8068;
wire n_8069;
wire n_8070;
wire n_8071;
wire n_8072;
wire n_8073;
wire n_8074;
wire n_8075;
wire n_8076;
wire n_8077;
wire n_8078;
wire n_8079;
wire n_8080;
wire n_8081;
wire n_8082;
wire n_8083;
wire n_8084;
wire n_8085;
wire n_8086;
wire n_8087;
wire n_8088;
wire n_8089;
wire n_8090;
wire n_8091;
wire n_8092;
wire n_8093;
wire n_8094;
wire n_8095;
wire n_8096;
wire n_8097;
wire n_8098;
wire n_8099;
wire n_8100;
wire n_8101;
wire n_8102;
wire n_8103;
wire n_8104;
wire n_8105;
wire n_8106;
wire n_8107;
wire n_8108;
wire n_8109;
wire n_8110;
wire n_8111;
wire n_8112;
wire n_8113;
wire n_8114;
wire n_8115;
wire n_8116;
wire n_8117;
wire n_8118;
wire n_8119;
wire n_8120;
wire n_8121;
wire n_8122;
wire n_8123;
wire n_8124;
wire n_8125;
wire n_8126;
wire n_8127;
wire n_8128;
wire n_8129;
wire n_8130;
wire n_8131;
wire n_8132;
wire n_8133;
wire n_8134;
wire n_8135;
wire n_8136;
wire n_8137;
wire n_8138;
wire n_8139;
wire n_8140;
wire n_8141;
wire n_8142;
wire n_8143;
wire n_8144;
wire n_8145;
wire n_8146;
wire n_8147;
wire n_8148;
wire n_8149;
wire n_8150;
wire n_8151;
wire n_8152;
wire n_8153;
wire n_8154;
wire n_8155;
wire n_8156;
wire n_8157;
wire n_8158;
wire n_8159;
wire n_8160;
wire n_8161;
wire n_8162;
wire n_8163;
wire n_8164;
wire n_8165;
wire n_8166;
wire n_8167;
wire n_8168;
wire n_8169;
wire n_8170;
wire n_8171;
wire n_8172;
wire n_8173;
wire n_8174;
wire n_8175;
wire n_8176;
wire n_8177;
wire n_8178;
wire n_8179;
wire n_8180;
wire n_8181;
wire n_8182;
wire n_8183;
wire n_8184;
wire n_8185;
wire n_8186;
wire n_8187;
wire n_8188;
wire n_8189;
wire n_8190;
wire n_8191;
wire n_8192;
wire n_8193;
wire n_8194;
wire n_8195;
wire n_8196;
wire n_8197;
wire n_8198;
wire n_8199;
wire n_8200;
wire n_8201;
wire n_8202;
wire n_8203;
wire n_8204;
wire n_8205;
wire n_8206;
wire n_8207;
wire n_8208;
wire n_8209;
wire n_8210;
wire n_8211;
wire n_8212;
wire n_8213;
wire n_8214;
wire n_8215;
wire n_8216;
wire n_8217;
wire n_8218;
wire n_8219;
wire n_8220;
wire n_8221;
wire n_8222;
wire n_8223;
wire n_8224;
wire n_8225;
wire n_8226;
wire n_8227;
wire n_8228;
wire n_8229;
wire n_8230;
wire n_8231;
wire n_8232;
wire n_8233;
wire n_8234;
wire n_8235;
wire n_8236;
wire n_8237;
wire n_8238;
wire n_8239;
wire n_8240;
wire n_8241;
wire n_8242;
wire n_8243;
wire n_8244;
wire n_8245;
wire n_8246;
wire n_8247;
wire n_8248;
wire n_8249;
wire n_8250;
wire n_8251;
wire n_8252;
wire n_8253;
wire n_8254;
wire n_8255;
wire n_8256;
wire n_8257;
wire n_8258;
wire n_8259;
wire n_8260;
wire n_8261;
wire n_8262;
wire n_8263;
wire n_8264;
wire n_8265;
wire n_8266;
wire n_8267;
wire n_8268;
wire n_8269;
wire n_8270;
wire n_8271;
wire n_8272;
wire n_8273;
wire n_8274;
wire n_8275;
wire n_8276;
wire n_8277;
wire n_8278;
wire n_8279;
wire n_8280;
wire n_8281;
wire n_8282;
wire n_8283;
wire n_8284;
wire n_8285;
wire n_8286;
wire n_8287;
wire n_8288;
wire n_8289;
wire n_8290;
wire n_8291;
wire n_8292;
wire n_8293;
wire n_8294;
wire n_8295;
wire n_8296;
wire n_8297;
wire n_8298;
wire n_8299;
wire n_8300;
wire n_8301;
wire n_8302;
wire n_8303;
wire n_8304;
wire n_8305;
wire n_8306;
wire n_8307;
wire n_8308;
wire n_8309;
wire n_8310;
wire n_8311;
wire n_8312;
wire n_8313;
wire n_8314;
wire n_8315;
wire n_8316;
wire n_8317;
wire n_8318;
wire n_8319;
wire n_8320;
wire n_8321;
wire n_8322;
wire n_8323;
wire n_8324;
wire n_8325;
wire n_8326;
wire n_8327;
wire n_8328;
wire n_8329;
wire n_8330;
wire n_8331;
wire n_8332;
wire n_8333;
wire n_8334;
wire n_8335;
wire n_8336;
wire n_8337;
wire n_8338;
wire n_8339;
wire n_8340;
wire n_8341;
wire n_8342;
wire n_8343;
wire n_8344;
wire n_8345;
wire n_8346;
wire n_8347;
wire n_8348;
wire n_8349;
wire n_8350;
wire n_8351;
wire n_8352;
wire n_8353;
wire n_8354;
wire n_8355;
wire n_8356;
wire n_8357;
wire n_8358;
wire n_8359;
wire n_8360;
wire n_8361;
wire n_8362;
wire n_8363;
wire n_8364;
wire n_8365;
wire n_8366;
wire n_8367;
wire n_8368;
wire n_8369;
wire n_8370;
wire n_8371;
wire n_8372;
wire n_8373;
wire n_8374;
wire n_8375;
wire n_8376;
wire n_8377;
wire n_8378;
wire n_8379;
wire n_8380;
wire n_8381;
wire n_8382;
wire n_8383;
wire n_8384;
wire n_8385;
wire n_8386;
wire n_8387;
wire n_8388;
wire n_8389;
wire n_8390;
wire n_8391;
wire n_8392;
wire n_8393;
wire n_8394;
wire n_8395;
wire n_8396;
wire n_8397;
wire n_8398;
wire n_8399;
wire n_8400;
wire n_8401;
wire n_8402;
wire n_8403;
wire n_8404;
wire n_8405;
wire n_8406;
wire n_8407;
wire n_8408;
wire n_8409;
wire n_8410;
wire n_8411;
wire n_8412;
wire n_8413;
wire n_8414;
wire n_8415;
wire n_8416;
wire n_8417;
wire n_8418;
wire n_8419;
wire n_8420;
wire n_8421;
wire n_8422;
wire n_8423;
wire n_8424;
wire n_8425;
wire n_8426;
wire n_8427;
wire n_8428;
wire n_8429;
wire n_8430;
wire n_8431;
wire n_8432;
wire n_8433;
wire n_8434;
wire n_8435;
wire n_8436;
wire n_8437;
wire n_8438;
wire n_8439;
wire n_8440;
wire n_8441;
wire n_8442;
wire n_8443;
wire n_8444;
wire n_8445;
wire n_8446;
wire n_8447;
wire n_8448;
wire n_8449;
wire n_8450;
wire n_8451;
wire n_8452;
wire n_8453;
wire n_8454;
wire n_8455;
wire n_8456;
wire n_8457;
wire n_8458;
wire n_8459;
wire n_8460;
wire n_8461;
wire n_8462;
wire n_8463;
wire n_8464;
wire n_8465;
wire n_8466;
wire n_8467;
wire n_8468;
wire n_8469;
wire n_8470;
wire n_8471;
wire n_8472;
wire n_8473;
wire n_8474;
wire n_8475;
wire n_8476;
wire n_8477;
wire n_8478;
wire n_8479;
wire n_8480;
wire n_8481;
wire n_8482;
wire n_8483;
wire n_8484;
wire n_8485;
wire n_8486;
wire n_8487;
wire n_8488;
wire n_8489;
wire n_8490;
wire n_8491;
wire n_8492;
wire n_8493;
wire n_8494;
wire n_8495;
wire n_8496;
wire n_8497;
wire n_8498;
wire n_8499;
wire n_8500;
wire n_8501;
wire n_8502;
wire n_8503;
wire n_8504;
wire n_8505;
wire n_8506;
wire n_8507;
wire n_8508;
wire n_8509;
wire n_8510;
wire n_8511;
wire n_8512;
wire n_8513;
wire n_8514;
wire n_8515;
wire n_8516;
wire n_8517;
wire n_8518;
wire n_8519;
wire n_8520;
wire n_8521;
wire n_8522;
wire n_8523;
wire n_8524;
wire n_8525;
wire n_8526;
wire n_8527;
wire n_8528;
wire n_8529;
wire n_8530;
wire n_8531;
wire n_8532;
wire n_8533;
wire n_8534;
wire n_8535;
wire n_8536;
wire n_8537;
wire n_8538;
wire n_8539;
wire n_8540;
wire n_8541;
wire n_8542;
wire n_8543;
wire n_8544;
wire n_8545;
wire n_8546;
wire n_8547;
wire n_8548;
wire n_8549;
wire n_8550;
wire n_8551;
wire n_8552;
wire n_8553;
wire n_8554;
wire n_8555;
wire n_8556;
wire n_8557;
wire n_8558;
wire n_8559;
wire n_8560;
wire n_8561;
wire n_8562;
wire n_8563;
wire n_8564;
wire n_8565;
wire n_8566;
wire n_8567;
wire n_8568;
wire n_8569;
wire n_8570;
wire n_8571;
wire n_8572;
wire n_8573;
wire n_8574;
wire n_8575;
wire n_8576;
wire n_8577;
wire n_8578;
wire n_8579;
wire n_8580;
wire n_8581;
wire n_8582;
wire n_8583;
wire n_8584;
wire n_8585;
wire n_8586;
wire n_8587;
wire n_8588;
wire n_8589;
wire n_8590;
wire n_8591;
wire n_8592;
wire n_8593;
wire n_8594;
wire n_8595;
wire n_8596;
wire n_8597;
wire n_8598;
wire n_8599;
wire n_8600;
wire n_8601;
wire n_8602;
wire n_8603;
wire n_8604;
wire n_8605;
wire n_8606;
wire n_8607;
wire n_8608;
wire n_8609;
wire n_8610;
wire n_8611;
wire n_8612;
wire n_8613;
wire n_8614;
wire n_8615;
wire n_8616;
wire n_8617;
wire n_8618;
wire n_8619;
wire n_8620;
wire n_8621;
wire n_8622;
wire n_8623;
wire n_8624;
wire n_8625;
wire n_8626;
wire n_8627;
wire n_8628;
wire n_8629;
wire n_8630;
wire n_8631;
wire n_8632;
wire n_8633;
wire n_8634;
wire n_8635;
wire n_8636;
wire n_8637;
wire n_8638;
wire n_8639;
wire n_8640;
wire n_8641;
wire n_8642;
wire n_8643;
wire n_8644;
wire n_8645;
wire n_8646;
wire n_8647;
wire n_8648;
wire n_8649;
wire n_8650;
wire n_8651;
wire n_8652;
wire n_8653;
wire n_8654;
wire n_8655;
wire n_8656;
wire n_8657;
wire n_8658;
wire n_8659;
wire n_8660;
wire n_8661;
wire n_8662;
wire n_8663;
wire n_8664;
wire n_8665;
wire n_8666;
wire n_8667;
wire n_8668;
wire n_8669;
wire n_8670;
wire n_8671;
wire n_8672;
wire n_8673;
wire n_8674;
wire n_8675;
wire n_8676;
wire n_8677;
wire n_8678;
wire n_8679;
wire n_8680;
wire n_8681;
wire n_8682;
wire n_8683;
wire n_8684;
wire n_8685;
wire n_8686;
wire n_8687;
wire n_8688;
wire n_8689;
wire n_8690;
wire n_8691;
wire n_8692;
wire n_8693;
wire n_8694;
wire n_8695;
wire n_8696;
wire n_8697;
wire n_8698;
wire n_8699;
wire n_8700;
wire n_8701;
wire n_8702;
wire n_8703;
wire n_8704;
wire n_8705;
wire n_8706;
wire n_8707;
wire n_8708;
wire n_8709;
wire n_8710;
wire n_8711;
wire n_8712;
wire n_8713;
wire n_8714;
wire n_8715;
wire n_8716;
wire n_8717;
wire n_8718;
wire n_8719;
wire n_8720;
wire n_8721;
wire n_8722;
wire n_8723;
wire n_8724;
wire n_8725;
wire n_8726;
wire n_8727;
wire n_8728;
wire n_8729;
wire n_8730;
wire n_8731;
wire n_8732;
wire n_8733;
wire n_8734;
wire n_8735;
wire n_8736;
wire n_8737;
wire n_8738;
wire n_8739;
wire n_8740;
wire n_8741;
wire n_8742;
wire n_8743;
wire n_8744;
wire n_8745;
wire n_8746;
wire n_8747;
wire n_8748;
wire n_8749;
wire n_8750;
wire n_8751;
wire n_8752;
wire n_8753;
wire n_8754;
wire n_8755;
wire n_8756;
wire n_8757;
wire n_8758;
wire n_8759;
wire n_8760;
wire n_8761;
wire n_8762;
wire n_8763;
wire n_8764;
wire n_8765;
wire n_8766;
wire n_8767;
wire n_8768;
wire n_8769;
wire n_8770;
wire n_8771;
wire n_8772;
wire n_8773;
wire n_8774;
wire n_8775;
wire n_8776;
wire n_8777;
wire n_8778;
wire n_8779;
wire n_8780;
wire n_8781;
wire n_8782;
wire n_8783;
wire n_8784;
wire n_8785;
wire n_8786;
wire n_8787;
wire n_8788;
wire n_8789;
wire n_8790;
wire n_8791;
wire n_8792;
wire n_8793;
wire n_8794;
wire n_8795;
wire n_8796;
wire n_8797;
wire n_8798;
wire n_8799;
wire n_8800;
wire n_8801;
wire n_8802;
wire n_8803;
wire n_8804;
wire n_8805;
wire n_8806;
wire n_8807;
wire n_8808;
wire n_8809;
wire n_8810;
wire n_8811;
wire n_8812;
wire n_8813;
wire n_8814;
wire n_8815;
wire n_8816;
wire n_8817;
wire n_8818;
wire n_8819;
wire n_8820;
wire n_8821;
wire n_8822;
wire n_8823;
wire n_8824;
wire n_8825;
wire n_8826;
wire n_8827;
wire n_8828;
wire n_8829;
wire n_8830;
wire n_8831;
wire n_8832;
wire n_8833;
wire n_8834;
wire n_8835;
wire n_8836;
wire n_8837;
wire n_8838;
wire n_8839;
wire n_8840;
wire n_8841;
wire n_8842;
wire n_8843;
wire n_8844;
wire n_8845;
wire n_8846;
wire n_8847;
wire n_8848;
wire n_8849;
wire n_8850;
wire n_8851;
wire n_8852;
wire n_8853;
wire n_8854;
wire n_8855;
wire n_8856;
wire n_8857;
wire n_8858;
wire n_8859;
wire n_8860;
wire n_8861;
wire n_8862;
wire n_8863;
wire n_8864;
wire n_8865;
wire n_8866;
wire n_8867;
wire n_8868;
wire n_8869;
wire n_8870;
wire n_8871;
wire n_8872;
wire n_8873;
wire n_8874;
wire n_8875;
wire n_8876;
wire n_8877;
wire n_8878;
wire n_8879;
wire n_8880;
wire n_8881;
wire n_8882;
wire n_8883;
wire n_8884;
wire n_8885;
wire n_8886;
wire n_8887;
wire n_8888;
wire n_8889;
wire n_8890;
wire n_8891;
wire n_8892;
wire n_8893;
wire n_8894;
wire n_8895;
wire n_8896;
wire n_8897;
wire n_8898;
wire n_8899;
wire n_8900;
wire n_8901;
wire n_8902;
wire n_8903;
wire n_8904;
wire n_8905;
wire n_8906;
wire n_8907;
wire n_8908;
wire n_8909;
wire n_8910;
wire n_8911;
wire n_8912;
wire n_8913;
wire n_8914;
wire n_8915;
wire n_8916;
wire n_8917;
wire n_8918;
wire n_8919;
wire n_8920;
wire n_8921;
wire n_8922;
wire n_8923;
wire n_8924;
wire n_8925;
wire n_8926;
wire n_8927;
wire n_8928;
wire n_8929;
wire n_8930;
wire n_8931;
wire n_8932;
wire n_8933;
wire n_8934;
wire n_8935;
wire n_8936;
wire n_8937;
wire n_8938;
wire n_8939;
wire n_8940;
wire n_8941;
wire n_8942;
wire n_8943;
wire n_8944;
wire n_8945;
wire n_8946;
wire n_8947;
wire n_8948;
wire n_8949;
wire n_8950;
wire n_8951;
wire n_8952;
wire n_8953;
wire n_8954;
wire n_8955;
wire n_8956;
wire n_8957;
wire n_8958;
wire n_8959;
wire n_8960;
wire n_8961;
wire n_8962;
wire n_8963;
wire n_8964;
wire n_8965;
wire n_8966;
wire n_8967;
wire n_8968;
wire n_8969;
wire n_8970;
wire n_8971;
wire n_8972;
wire n_8973;
wire n_8974;
wire n_8975;
wire n_8976;
wire n_8977;
wire n_8978;
wire n_8979;
wire n_8980;
wire n_8981;
wire n_8982;
wire n_8983;
wire n_8984;
wire n_8985;
wire n_8986;
wire n_8987;
wire n_8988;
wire n_8989;
wire n_8990;
wire n_8991;
wire n_8992;
wire n_8993;
wire n_8994;
wire n_8995;
wire n_8996;
wire n_8997;
wire n_8998;
wire n_8999;
wire n_9000;
wire n_9001;
wire n_9002;
wire n_9003;
wire n_9004;
wire n_9005;
wire n_9006;
wire n_9007;
wire n_9008;
wire n_9009;
wire n_9010;
wire n_9011;
wire n_9012;
wire n_9013;
wire n_9014;
wire n_9015;
wire n_9016;
wire n_9017;
wire n_9018;
wire n_9019;
wire n_9020;
wire n_9021;
wire n_9022;
wire n_9023;
wire n_9024;
wire n_9025;
wire n_9026;
wire n_9027;
wire n_9028;
wire n_9029;
wire n_9030;
wire n_9031;
wire n_9032;
wire n_9033;
wire n_9034;
wire n_9035;
wire n_9036;
wire n_9037;
wire n_9038;
wire n_9039;
wire n_9040;
wire n_9041;
wire n_9042;
wire n_9043;
wire n_9044;
wire n_9045;
wire n_9046;
wire n_9047;
wire n_9048;
wire n_9049;
wire n_9050;
wire n_9051;
wire n_9052;
wire n_9053;
wire n_9054;
wire n_9055;
wire n_9056;
wire n_9057;
wire n_9058;
wire n_9059;
wire n_9060;
wire n_9061;
wire n_9062;
wire n_9063;
wire n_9064;
wire n_9065;
wire n_9066;
wire n_9067;
wire n_9068;
wire n_9069;
wire n_9070;
wire n_9071;
wire n_9072;
wire n_9073;
wire n_9074;
wire n_9075;
wire n_9076;
wire n_9077;
wire n_9078;
wire n_9079;
wire n_9080;
wire n_9081;
wire n_9082;
wire n_9083;
wire n_9084;
wire n_9085;
wire n_9086;
wire n_9087;
wire n_9088;
wire n_9089;
wire n_9090;
wire n_9091;
wire n_9092;
wire n_9093;
wire n_9094;
wire n_9095;
wire n_9096;
wire n_9097;
wire n_9098;
wire n_9099;
wire n_9100;
wire n_9101;
wire n_9102;
wire n_9103;
wire n_9104;
wire n_9105;
wire n_9106;
wire n_9107;
wire n_9108;
wire n_9109;
wire n_9110;
wire n_9111;
wire n_9112;
wire n_9113;
wire n_9114;
wire n_9115;
wire n_9116;
wire n_9117;
wire n_9118;
wire n_9119;
wire n_9120;
wire n_9121;
wire n_9122;
wire n_9123;
wire n_9124;
wire n_9125;
wire n_9126;
wire n_9127;
wire n_9128;
wire n_9129;
wire n_9130;
wire n_9131;
wire n_9132;
wire n_9133;
wire n_9134;
wire n_9135;
wire n_9136;
wire n_9137;
wire n_9138;
wire n_9139;
wire n_9140;
wire n_9141;
wire n_9142;
wire n_9143;
wire n_9144;
wire n_9145;
wire n_9146;
wire n_9147;
wire n_9148;
wire n_9149;
wire n_9150;
wire n_9151;
wire n_9152;
wire n_9153;
wire n_9154;
wire n_9155;
wire n_9156;
wire n_9157;
wire n_9158;
wire n_9159;
wire n_9160;
wire n_9161;
wire n_9162;
wire n_9163;
wire n_9164;
wire n_9165;
wire n_9166;
wire n_9167;
wire n_9168;
wire n_9169;
wire n_9170;
wire n_9171;
wire n_9172;
wire n_9173;
wire n_9174;
wire n_9175;
wire n_9176;
wire n_9177;
wire n_9178;
wire n_9179;
wire n_9180;
wire n_9181;
wire n_9182;
wire n_9183;
wire n_9184;
wire n_9185;
wire n_9186;
wire n_9187;
wire n_9188;
wire n_9189;
wire n_9190;
wire n_9191;
wire n_9192;
wire n_9193;
wire n_9194;
wire n_9195;
wire n_9196;
wire n_9197;
wire n_9198;
wire n_9199;
wire n_9200;
wire n_9201;
wire n_9202;
wire n_9203;
wire n_9204;
wire n_9205;
wire n_9206;
wire n_9207;
wire n_9208;
wire n_9209;
wire n_9210;
wire n_9211;
wire n_9212;
wire n_9213;
wire n_9214;
wire n_9215;
wire n_9216;
wire n_9217;
wire n_9218;
wire n_9219;
wire n_9220;
wire n_9221;
wire n_9222;
wire n_9223;
wire n_9224;
wire n_9225;
wire n_9226;
wire n_9227;
wire n_9228;
wire n_9229;
wire n_9230;
wire n_9231;
wire n_9232;
wire n_9233;
wire n_9234;
wire n_9235;
wire n_9236;
wire n_9237;
wire n_9238;
wire n_9239;
wire n_9240;
wire n_9241;
wire n_9242;
wire n_9243;
wire n_9244;
wire n_9245;
wire n_9246;
wire n_9247;
wire n_9248;
wire n_9249;
wire n_9250;
wire n_9251;
wire n_9252;
wire n_9253;
wire n_9254;
wire n_9255;
wire n_9256;
wire n_9257;
wire n_9258;
wire n_9259;
wire n_9260;
wire n_9261;
wire n_9262;
wire n_9263;
wire n_9264;
wire n_9265;
wire n_9266;
wire n_9267;
wire n_9268;
wire n_9269;
wire n_9270;
wire n_9271;
wire n_9272;
wire n_9273;
wire n_9274;
wire n_9275;
wire n_9276;
wire n_9277;
wire n_9278;
wire n_9279;
wire n_9280;
wire n_9281;
wire n_9282;
wire n_9283;
wire n_9284;
wire n_9285;
wire n_9286;
wire n_9287;
wire n_9288;
wire n_9289;
wire n_9290;
wire n_9291;
wire n_9292;
wire n_9293;
wire n_9294;
wire n_9295;
wire n_9296;
wire n_9297;
wire n_9298;
wire n_9299;
wire n_9300;
wire n_9301;
wire n_9302;
wire n_9303;
wire n_9304;
wire n_9305;
wire n_9306;
wire n_9307;
wire n_9308;
wire n_9309;
wire n_9310;
wire n_9311;
wire n_9312;
wire n_9313;
wire n_9314;
wire n_9315;
wire n_9316;
wire n_9317;
wire n_9318;
wire n_9319;
wire n_9320;
wire n_9321;
wire n_9322;
wire n_9323;
wire n_9324;
wire n_9325;
wire n_9326;
wire n_9327;
wire n_9328;
wire n_9329;
wire n_9330;
wire n_9331;
wire n_9332;
wire n_9333;
wire n_9334;
wire n_9335;
wire n_9336;
wire n_9337;
wire n_9338;
wire n_9339;
wire n_9340;
wire n_9341;
wire n_9342;
wire n_9343;
wire n_9344;
wire n_9345;
wire n_9346;
wire n_9347;
wire n_9348;
wire n_9349;
wire n_9350;
wire n_9351;
wire n_9352;
wire n_9353;
wire n_9354;
wire n_9355;
wire n_9356;
wire n_9357;
wire n_9358;
wire n_9359;
wire n_9360;
wire n_9361;
wire n_9362;
wire n_9363;
wire n_9364;
wire n_9365;
wire n_9366;
wire n_9367;
wire n_9368;
wire n_9369;
wire n_9370;
wire n_9371;
wire n_9372;
wire n_9373;
wire n_9374;
wire n_9375;
wire n_9376;
wire n_9377;
wire n_9378;
wire n_9379;
wire n_9380;
wire n_9381;
wire n_9382;
wire n_9383;
wire n_9384;
wire n_9385;
wire n_9386;
wire n_9387;
wire n_9388;
wire n_9389;
wire n_9390;
wire n_9391;
wire n_9392;
wire n_9393;
wire n_9394;
wire n_9395;
wire n_9396;
wire n_9397;
wire n_9398;
wire n_9399;
wire n_9400;
wire n_9401;
wire n_9402;
wire n_9403;
wire n_9404;
wire n_9405;
wire n_9406;
wire n_9407;
wire n_9408;
wire n_9409;
wire n_9410;
wire n_9411;
wire n_9412;
wire n_9413;
wire n_9414;
wire n_9415;
wire n_9416;
wire n_9417;
wire n_9418;
wire n_9419;
wire n_9420;
wire n_9421;
wire n_9422;
wire n_9423;
wire n_9424;
wire n_9425;
wire n_9426;
wire n_9427;
wire n_9428;
wire n_9429;
wire n_9430;
wire n_9431;
wire n_9432;
wire n_9433;
wire n_9434;
wire n_9435;
wire n_9436;
wire n_9437;
wire n_9438;
wire n_9439;
wire n_9440;
wire n_9441;
wire n_9442;
wire n_9443;
wire n_9444;
wire n_9445;
wire n_9446;
wire n_9447;
wire n_9448;
wire n_9449;
wire n_9450;
wire n_9451;
wire n_9452;
wire n_9453;
wire n_9454;
wire n_9455;
wire n_9456;
wire n_9457;
wire n_9458;
wire n_9459;
wire n_9460;
wire n_9461;
wire n_9462;
wire n_9463;
wire n_9464;
wire n_9465;
wire n_9466;
wire n_9467;
wire n_9468;
wire n_9469;
wire n_9470;
wire n_9471;
wire n_9472;
wire n_9473;
wire n_9474;
wire n_9475;
wire n_9476;
wire n_9477;
wire n_9478;
wire n_9479;
wire n_9480;
wire n_9481;
wire n_9482;
wire n_9483;
wire n_9484;
wire n_9485;
wire n_9486;
wire n_9487;
wire n_9488;
wire n_9489;
wire n_9490;
wire n_9491;
wire n_9492;
wire n_9493;
wire n_9494;
wire n_9495;
wire n_9496;
wire n_9497;
wire n_9498;
wire n_9499;
wire n_9500;
wire n_9501;
wire n_9502;
wire n_9503;
wire n_9504;
wire n_9505;
wire n_9506;
wire n_9507;
wire n_9508;
wire n_9509;
wire n_9510;
wire n_9511;
wire n_9512;
wire n_9513;
wire n_9514;
wire n_9515;
wire n_9516;
wire n_9517;
wire n_9518;
wire n_9519;
wire n_9520;
wire n_9521;
wire n_9522;
wire n_9523;
wire n_9524;
wire n_9525;
wire n_9526;
wire n_9527;
wire n_9528;
wire n_9529;
wire n_9530;
wire n_9531;
wire n_9532;
wire n_9533;
wire n_9534;
wire n_9535;
wire n_9536;
wire n_9537;
wire n_9538;
wire n_9539;
wire n_9540;
wire n_9541;
wire n_9542;
wire n_9543;
wire n_9544;
wire n_9545;
wire n_9546;
wire n_9547;
wire n_9548;
wire n_9549;
wire n_9550;
wire n_9551;
wire n_9552;
wire n_9553;
wire n_9554;
wire n_9555;
wire n_9556;
wire n_9557;
wire n_9558;
wire n_9559;
wire n_9560;
wire n_9561;
wire n_9562;
wire n_9563;
wire n_9564;
wire n_9565;
wire n_9566;
wire n_9567;
wire n_9568;
wire n_9569;
wire n_9570;
wire n_9571;
wire n_9572;
wire n_9573;
wire n_9574;
wire n_9575;
wire n_9576;
wire n_9577;
wire n_9578;
wire n_9579;
wire n_9580;
wire n_9581;
wire n_9582;
wire n_9583;
wire n_9584;
wire n_9585;
wire n_9586;
wire n_9587;
wire n_9588;
wire n_9589;
wire n_9590;
wire n_9591;
wire n_9592;
wire n_9593;
wire n_9594;
wire n_9595;
wire n_9596;
wire n_9597;
wire n_9598;
wire n_9599;
wire n_9600;
wire n_9601;
wire n_9602;
wire n_9603;
wire n_9604;
wire n_9605;
wire n_9606;
wire n_9607;
wire n_9608;
wire n_9609;
wire n_9610;
wire n_9611;
wire n_9612;
wire n_9613;
wire n_9614;
wire n_9615;
wire n_9616;
wire n_9617;
wire n_9618;
wire n_9619;
wire n_9620;
wire n_9621;
wire n_9622;
wire n_9623;
wire n_9624;
wire n_9625;
wire n_9626;
wire n_9627;
wire n_9628;
wire n_9629;
wire n_9630;
wire n_9631;
wire n_9632;
wire n_9633;
wire n_9634;
wire n_9635;
wire n_9636;
wire n_9637;
wire n_9638;
wire n_9639;
wire n_9640;
wire n_9641;
wire n_9642;
wire n_9643;
wire n_9644;
wire n_9645;
wire n_9646;
wire n_9647;
wire n_9648;
wire n_9649;
wire n_9650;
wire n_9651;
wire n_9652;
wire n_9653;
wire n_9654;
wire n_9655;
wire n_9656;
wire n_9657;
assign n_1 = ~x_40 & ~x_41;
assign n_2 = ~x_42 &  n_1;
assign n_3 =  x_39 &  n_2;
assign n_4 = ~x_36 &  x_37;
assign n_5 = ~x_33 &  x_34;
assign n_6 = ~x_35 &  n_5;
assign n_7 =  n_4 &  n_6;
assign n_8 = ~x_38 &  n_7;
assign n_9 =  n_3 &  n_8;
assign n_10 =  x_66 & ~n_9;
assign n_11 =  x_258 &  n_9;
assign n_12 = ~n_10 & ~n_11;
assign n_13 =  x_66 & ~n_12;
assign n_14 = ~x_66 &  n_12;
assign n_15 = ~n_13 & ~n_14;
assign n_16 =  x_65 & ~n_9;
assign n_17 =  x_257 &  n_9;
assign n_18 = ~n_16 & ~n_17;
assign n_19 =  x_65 & ~n_18;
assign n_20 = ~x_65 &  n_18;
assign n_21 = ~n_19 & ~n_20;
assign n_22 =  x_64 & ~n_9;
assign n_23 =  x_256 &  n_9;
assign n_24 = ~n_22 & ~n_23;
assign n_25 =  x_64 & ~n_24;
assign n_26 = ~x_64 &  n_24;
assign n_27 = ~n_25 & ~n_26;
assign n_28 =  x_63 & ~n_9;
assign n_29 =  x_255 &  n_9;
assign n_30 = ~n_28 & ~n_29;
assign n_31 =  x_63 & ~n_30;
assign n_32 = ~x_63 &  n_30;
assign n_33 = ~n_31 & ~n_32;
assign n_34 =  x_62 & ~n_9;
assign n_35 =  x_254 &  n_9;
assign n_36 = ~n_34 & ~n_35;
assign n_37 =  x_62 & ~n_36;
assign n_38 = ~x_62 &  n_36;
assign n_39 = ~n_37 & ~n_38;
assign n_40 =  x_61 & ~n_9;
assign n_41 =  x_253 &  n_9;
assign n_42 = ~n_40 & ~n_41;
assign n_43 =  x_61 & ~n_42;
assign n_44 = ~x_61 &  n_42;
assign n_45 = ~n_43 & ~n_44;
assign n_46 =  x_60 & ~n_9;
assign n_47 =  x_252 &  n_9;
assign n_48 = ~n_46 & ~n_47;
assign n_49 =  x_60 & ~n_48;
assign n_50 = ~x_60 &  n_48;
assign n_51 = ~n_49 & ~n_50;
assign n_52 =  x_59 & ~n_9;
assign n_53 =  x_251 &  n_9;
assign n_54 = ~n_52 & ~n_53;
assign n_55 =  x_59 & ~n_54;
assign n_56 = ~x_59 &  n_54;
assign n_57 = ~n_55 & ~n_56;
assign n_58 =  x_58 & ~n_9;
assign n_59 =  x_250 &  n_9;
assign n_60 = ~n_58 & ~n_59;
assign n_61 =  x_58 & ~n_60;
assign n_62 = ~x_58 &  n_60;
assign n_63 = ~n_61 & ~n_62;
assign n_64 =  x_57 & ~n_9;
assign n_65 =  x_249 &  n_9;
assign n_66 = ~n_64 & ~n_65;
assign n_67 =  x_57 & ~n_66;
assign n_68 = ~x_57 &  n_66;
assign n_69 = ~n_67 & ~n_68;
assign n_70 =  x_56 & ~n_9;
assign n_71 =  x_248 &  n_9;
assign n_72 = ~n_70 & ~n_71;
assign n_73 =  x_56 & ~n_72;
assign n_74 = ~x_56 &  n_72;
assign n_75 = ~n_73 & ~n_74;
assign n_76 =  x_55 & ~n_9;
assign n_77 =  x_247 &  n_9;
assign n_78 = ~n_76 & ~n_77;
assign n_79 =  x_55 & ~n_78;
assign n_80 = ~x_55 &  n_78;
assign n_81 = ~n_79 & ~n_80;
assign n_82 =  x_54 & ~n_9;
assign n_83 =  x_246 &  n_9;
assign n_84 = ~n_82 & ~n_83;
assign n_85 =  x_54 & ~n_84;
assign n_86 = ~x_54 &  n_84;
assign n_87 = ~n_85 & ~n_86;
assign n_88 =  x_53 & ~n_9;
assign n_89 =  x_245 &  n_9;
assign n_90 = ~n_88 & ~n_89;
assign n_91 =  x_53 & ~n_90;
assign n_92 = ~x_53 &  n_90;
assign n_93 = ~n_91 & ~n_92;
assign n_94 =  x_52 & ~n_9;
assign n_95 =  x_244 &  n_9;
assign n_96 = ~n_94 & ~n_95;
assign n_97 =  x_52 & ~n_96;
assign n_98 = ~x_52 &  n_96;
assign n_99 = ~n_97 & ~n_98;
assign n_100 =  x_51 & ~n_9;
assign n_101 =  x_243 &  n_9;
assign n_102 = ~n_100 & ~n_101;
assign n_103 =  x_51 & ~n_102;
assign n_104 = ~x_51 &  n_102;
assign n_105 = ~n_103 & ~n_104;
assign n_106 =  x_50 & ~n_9;
assign n_107 =  x_242 &  n_9;
assign n_108 = ~n_106 & ~n_107;
assign n_109 =  x_50 & ~n_108;
assign n_110 = ~x_50 &  n_108;
assign n_111 = ~n_109 & ~n_110;
assign n_112 =  x_49 & ~n_9;
assign n_113 =  x_241 &  n_9;
assign n_114 = ~n_112 & ~n_113;
assign n_115 =  x_49 & ~n_114;
assign n_116 = ~x_49 &  n_114;
assign n_117 = ~n_115 & ~n_116;
assign n_118 =  x_48 & ~n_9;
assign n_119 =  x_240 &  n_9;
assign n_120 = ~n_118 & ~n_119;
assign n_121 =  x_48 & ~n_120;
assign n_122 = ~x_48 &  n_120;
assign n_123 = ~n_121 & ~n_122;
assign n_124 =  x_47 & ~n_9;
assign n_125 =  x_239 &  n_9;
assign n_126 = ~n_124 & ~n_125;
assign n_127 =  x_47 & ~n_126;
assign n_128 = ~x_47 &  n_126;
assign n_129 = ~n_127 & ~n_128;
assign n_130 =  x_46 & ~n_9;
assign n_131 =  x_238 &  n_9;
assign n_132 = ~n_130 & ~n_131;
assign n_133 =  x_46 & ~n_132;
assign n_134 = ~x_46 &  n_132;
assign n_135 = ~n_133 & ~n_134;
assign n_136 =  x_45 & ~n_9;
assign n_137 =  x_237 &  n_9;
assign n_138 = ~n_136 & ~n_137;
assign n_139 =  x_45 & ~n_138;
assign n_140 = ~x_45 &  n_138;
assign n_141 = ~n_139 & ~n_140;
assign n_142 =  x_44 & ~n_9;
assign n_143 =  x_236 &  n_9;
assign n_144 = ~n_142 & ~n_143;
assign n_145 =  x_44 & ~n_144;
assign n_146 = ~x_44 &  n_144;
assign n_147 = ~n_145 & ~n_146;
assign n_148 =  x_43 & ~n_9;
assign n_149 =  x_235 &  n_9;
assign n_150 = ~n_148 & ~n_149;
assign n_151 =  x_43 & ~n_150;
assign n_152 = ~x_43 &  n_150;
assign n_153 = ~n_151 & ~n_152;
assign n_154 = ~x_139 &  x_935;
assign n_155 =  x_139 & ~x_935;
assign n_156 =  x_140 & ~x_936;
assign n_157 = ~x_140 &  x_936;
assign n_158 =  x_141 & ~x_937;
assign n_159 = ~x_141 &  x_937;
assign n_160 =  x_142 & ~x_938;
assign n_161 = ~x_142 &  x_938;
assign n_162 =  x_143 & ~x_939;
assign n_163 = ~x_143 &  x_939;
assign n_164 =  x_144 & ~x_940;
assign n_165 = ~x_144 &  x_940;
assign n_166 =  x_145 & ~x_941;
assign n_167 = ~x_145 &  x_941;
assign n_168 =  x_146 & ~x_942;
assign n_169 = ~x_146 &  x_942;
assign n_170 =  x_147 & ~x_943;
assign n_171 = ~x_147 &  x_943;
assign n_172 =  x_148 & ~x_944;
assign n_173 = ~x_148 &  x_944;
assign n_174 =  x_149 & ~x_945;
assign n_175 = ~x_149 &  x_945;
assign n_176 =  x_150 & ~x_946;
assign n_177 = ~x_150 &  x_946;
assign n_178 =  x_151 & ~x_947;
assign n_179 = ~x_151 &  x_947;
assign n_180 =  x_152 & ~x_948;
assign n_181 = ~x_152 &  x_948;
assign n_182 =  x_153 & ~x_949;
assign n_183 = ~x_153 &  x_949;
assign n_184 =  x_154 & ~x_950;
assign n_185 = ~x_154 &  x_950;
assign n_186 =  x_155 & ~x_951;
assign n_187 = ~x_155 &  x_951;
assign n_188 =  x_156 & ~x_952;
assign n_189 = ~x_156 &  x_952;
assign n_190 =  x_157 & ~x_953;
assign n_191 = ~x_157 &  x_953;
assign n_192 =  x_158 & ~x_954;
assign n_193 = ~x_158 &  x_954;
assign n_194 =  x_159 & ~x_955;
assign n_195 = ~x_159 &  x_955;
assign n_196 =  x_160 & ~x_956;
assign n_197 = ~x_160 &  x_956;
assign n_198 =  x_161 & ~x_957;
assign n_199 = ~x_161 &  x_957;
assign n_200 =  x_162 & ~x_958;
assign n_201 = ~x_162 &  x_958;
assign n_202 =  x_163 & ~x_959;
assign n_203 = ~x_163 &  x_959;
assign n_204 =  x_164 & ~x_960;
assign n_205 = ~x_164 &  x_960;
assign n_206 =  x_165 & ~x_961;
assign n_207 = ~x_165 &  x_961;
assign n_208 =  x_166 & ~x_962;
assign n_209 = ~x_166 &  x_962;
assign n_210 =  x_167 & ~x_963;
assign n_211 = ~x_167 &  x_963;
assign n_212 =  x_168 & ~x_964;
assign n_213 = ~x_168 &  x_964;
assign n_214 =  x_169 & ~x_965;
assign n_215 = ~x_169 &  x_965;
assign n_216 =  x_170 & ~x_966;
assign n_217 = ~n_215 &  n_216;
assign n_218 = ~n_214 & ~n_217;
assign n_219 = ~n_213 & ~n_218;
assign n_220 = ~n_212 & ~n_219;
assign n_221 = ~n_211 & ~n_220;
assign n_222 = ~n_210 & ~n_221;
assign n_223 = ~n_209 & ~n_222;
assign n_224 = ~n_208 & ~n_223;
assign n_225 = ~n_207 & ~n_224;
assign n_226 = ~n_206 & ~n_225;
assign n_227 = ~n_205 & ~n_226;
assign n_228 = ~n_204 & ~n_227;
assign n_229 = ~n_203 & ~n_228;
assign n_230 = ~n_202 & ~n_229;
assign n_231 = ~n_201 & ~n_230;
assign n_232 = ~n_200 & ~n_231;
assign n_233 = ~n_199 & ~n_232;
assign n_234 = ~n_198 & ~n_233;
assign n_235 = ~n_197 & ~n_234;
assign n_236 = ~n_196 & ~n_235;
assign n_237 = ~n_195 & ~n_236;
assign n_238 = ~n_194 & ~n_237;
assign n_239 = ~n_193 & ~n_238;
assign n_240 = ~n_192 & ~n_239;
assign n_241 = ~n_191 & ~n_240;
assign n_242 = ~n_190 & ~n_241;
assign n_243 = ~n_189 & ~n_242;
assign n_244 = ~n_188 & ~n_243;
assign n_245 = ~n_187 & ~n_244;
assign n_246 = ~n_186 & ~n_245;
assign n_247 = ~n_185 & ~n_246;
assign n_248 = ~n_184 & ~n_247;
assign n_249 = ~n_183 & ~n_248;
assign n_250 = ~n_182 & ~n_249;
assign n_251 = ~n_181 & ~n_250;
assign n_252 = ~n_180 & ~n_251;
assign n_253 = ~n_179 & ~n_252;
assign n_254 = ~n_178 & ~n_253;
assign n_255 = ~n_177 & ~n_254;
assign n_256 = ~n_176 & ~n_255;
assign n_257 = ~n_175 & ~n_256;
assign n_258 = ~n_174 & ~n_257;
assign n_259 = ~n_173 & ~n_258;
assign n_260 = ~n_172 & ~n_259;
assign n_261 = ~n_171 & ~n_260;
assign n_262 = ~n_170 & ~n_261;
assign n_263 = ~n_169 & ~n_262;
assign n_264 = ~n_168 & ~n_263;
assign n_265 = ~n_167 & ~n_264;
assign n_266 = ~n_166 & ~n_265;
assign n_267 = ~n_165 & ~n_266;
assign n_268 = ~n_164 & ~n_267;
assign n_269 = ~n_163 & ~n_268;
assign n_270 = ~n_162 & ~n_269;
assign n_271 = ~n_161 & ~n_270;
assign n_272 = ~n_160 & ~n_271;
assign n_273 = ~n_159 & ~n_272;
assign n_274 = ~n_158 & ~n_273;
assign n_275 = ~n_157 & ~n_274;
assign n_276 = ~n_156 & ~n_275;
assign n_277 = ~n_155 & ~n_276;
assign n_278 = ~n_154 & ~n_277;
assign n_279 = ~x_40 &  x_41;
assign n_280 =  x_42 &  n_279;
assign n_281 =  x_39 &  n_280;
assign n_282 =  x_33 & ~x_34;
assign n_283 =  x_35 & ~x_36;
assign n_284 =  n_282 &  n_283;
assign n_285 =  x_37 &  n_284;
assign n_286 = ~x_38 &  n_285;
assign n_287 =  n_281 &  n_286;
assign n_288 =  n_278 &  n_287;
assign n_289 = ~x_41 &  x_42;
assign n_290 = ~x_39 &  x_40;
assign n_291 =  n_289 &  n_290;
assign n_292 = ~x_38 &  n_291;
assign n_293 = ~x_107 &  x_935;
assign n_294 =  x_107 & ~x_935;
assign n_295 =  x_108 & ~x_936;
assign n_296 = ~x_108 &  x_936;
assign n_297 =  x_109 & ~x_937;
assign n_298 = ~x_109 &  x_937;
assign n_299 =  x_110 & ~x_938;
assign n_300 = ~x_110 &  x_938;
assign n_301 =  x_111 & ~x_939;
assign n_302 = ~x_111 &  x_939;
assign n_303 =  x_112 & ~x_940;
assign n_304 = ~x_112 &  x_940;
assign n_305 =  x_113 & ~x_941;
assign n_306 = ~x_113 &  x_941;
assign n_307 =  x_114 & ~x_942;
assign n_308 = ~x_114 &  x_942;
assign n_309 =  x_115 & ~x_943;
assign n_310 = ~x_115 &  x_943;
assign n_311 =  x_116 & ~x_944;
assign n_312 = ~x_116 &  x_944;
assign n_313 =  x_117 & ~x_945;
assign n_314 = ~x_117 &  x_945;
assign n_315 =  x_118 & ~x_946;
assign n_316 = ~x_118 &  x_946;
assign n_317 =  x_119 & ~x_947;
assign n_318 = ~x_119 &  x_947;
assign n_319 =  x_120 & ~x_948;
assign n_320 = ~x_120 &  x_948;
assign n_321 =  x_121 & ~x_949;
assign n_322 = ~x_121 &  x_949;
assign n_323 =  x_122 & ~x_950;
assign n_324 = ~x_122 &  x_950;
assign n_325 =  x_123 & ~x_951;
assign n_326 = ~x_123 &  x_951;
assign n_327 =  x_124 & ~x_952;
assign n_328 = ~x_124 &  x_952;
assign n_329 =  x_125 & ~x_953;
assign n_330 = ~x_125 &  x_953;
assign n_331 =  x_126 & ~x_954;
assign n_332 = ~x_126 &  x_954;
assign n_333 =  x_127 & ~x_955;
assign n_334 = ~x_127 &  x_955;
assign n_335 =  x_128 & ~x_956;
assign n_336 = ~x_128 &  x_956;
assign n_337 =  x_129 & ~x_957;
assign n_338 = ~x_129 &  x_957;
assign n_339 =  x_130 & ~x_958;
assign n_340 = ~x_130 &  x_958;
assign n_341 =  x_131 & ~x_959;
assign n_342 = ~x_131 &  x_959;
assign n_343 =  x_132 & ~x_960;
assign n_344 = ~x_132 &  x_960;
assign n_345 =  x_133 & ~x_961;
assign n_346 = ~x_133 &  x_961;
assign n_347 =  x_134 & ~x_962;
assign n_348 = ~x_134 &  x_962;
assign n_349 =  x_135 & ~x_963;
assign n_350 = ~x_135 &  x_963;
assign n_351 =  x_136 & ~x_964;
assign n_352 = ~x_136 &  x_964;
assign n_353 =  x_137 & ~x_965;
assign n_354 = ~x_137 &  x_965;
assign n_355 =  x_138 & ~x_966;
assign n_356 = ~n_354 &  n_355;
assign n_357 = ~n_353 & ~n_356;
assign n_358 = ~n_352 & ~n_357;
assign n_359 = ~n_351 & ~n_358;
assign n_360 = ~n_350 & ~n_359;
assign n_361 = ~n_349 & ~n_360;
assign n_362 = ~n_348 & ~n_361;
assign n_363 = ~n_347 & ~n_362;
assign n_364 = ~n_346 & ~n_363;
assign n_365 = ~n_345 & ~n_364;
assign n_366 = ~n_344 & ~n_365;
assign n_367 = ~n_343 & ~n_366;
assign n_368 = ~n_342 & ~n_367;
assign n_369 = ~n_341 & ~n_368;
assign n_370 = ~n_340 & ~n_369;
assign n_371 = ~n_339 & ~n_370;
assign n_372 = ~n_338 & ~n_371;
assign n_373 = ~n_337 & ~n_372;
assign n_374 = ~n_336 & ~n_373;
assign n_375 = ~n_335 & ~n_374;
assign n_376 = ~n_334 & ~n_375;
assign n_377 = ~n_333 & ~n_376;
assign n_378 = ~n_332 & ~n_377;
assign n_379 = ~n_331 & ~n_378;
assign n_380 = ~n_330 & ~n_379;
assign n_381 = ~n_329 & ~n_380;
assign n_382 = ~n_328 & ~n_381;
assign n_383 = ~n_327 & ~n_382;
assign n_384 = ~n_326 & ~n_383;
assign n_385 = ~n_325 & ~n_384;
assign n_386 = ~n_324 & ~n_385;
assign n_387 = ~n_323 & ~n_386;
assign n_388 = ~n_322 & ~n_387;
assign n_389 = ~n_321 & ~n_388;
assign n_390 = ~n_320 & ~n_389;
assign n_391 = ~n_319 & ~n_390;
assign n_392 = ~n_318 & ~n_391;
assign n_393 = ~n_317 & ~n_392;
assign n_394 = ~n_316 & ~n_393;
assign n_395 = ~n_315 & ~n_394;
assign n_396 = ~n_314 & ~n_395;
assign n_397 = ~n_313 & ~n_396;
assign n_398 = ~n_312 & ~n_397;
assign n_399 = ~n_311 & ~n_398;
assign n_400 = ~n_310 & ~n_399;
assign n_401 = ~n_309 & ~n_400;
assign n_402 = ~n_308 & ~n_401;
assign n_403 = ~n_307 & ~n_402;
assign n_404 = ~n_306 & ~n_403;
assign n_405 = ~n_305 & ~n_404;
assign n_406 = ~n_304 & ~n_405;
assign n_407 = ~n_303 & ~n_406;
assign n_408 = ~n_302 & ~n_407;
assign n_409 = ~n_301 & ~n_408;
assign n_410 = ~n_300 & ~n_409;
assign n_411 = ~n_299 & ~n_410;
assign n_412 = ~n_298 & ~n_411;
assign n_413 = ~n_297 & ~n_412;
assign n_414 = ~n_296 & ~n_413;
assign n_415 = ~n_295 & ~n_414;
assign n_416 = ~n_294 & ~n_415;
assign n_417 = ~n_293 & ~n_416;
assign n_418 = ~n_417 &  n_285;
assign n_419 =  n_292 &  n_418;
assign n_420 = ~n_288 & ~n_419;
assign n_421 =  x_40 &  x_41;
assign n_422 =  x_42 &  n_421;
assign n_423 = ~x_37 &  x_38;
assign n_424 = ~x_39 &  n_423;
assign n_425 =  n_422 &  n_424;
assign n_426 =  x_75 & ~x_1063;
assign n_427 = ~x_75 &  x_1063;
assign n_428 = ~x_76 &  x_1064;
assign n_429 =  x_76 & ~x_1064;
assign n_430 = ~x_77 &  x_1065;
assign n_431 =  x_77 & ~x_1065;
assign n_432 = ~x_78 &  x_1066;
assign n_433 =  x_78 & ~x_1066;
assign n_434 = ~x_79 &  x_1067;
assign n_435 =  x_79 & ~x_1067;
assign n_436 = ~x_80 &  x_1068;
assign n_437 =  x_80 & ~x_1068;
assign n_438 = ~x_81 &  x_1069;
assign n_439 =  x_81 & ~x_1069;
assign n_440 = ~x_82 &  x_1070;
assign n_441 =  x_82 & ~x_1070;
assign n_442 = ~x_83 &  x_1071;
assign n_443 =  x_83 & ~x_1071;
assign n_444 = ~x_84 &  x_1072;
assign n_445 =  x_84 & ~x_1072;
assign n_446 = ~x_85 &  x_1073;
assign n_447 =  x_85 & ~x_1073;
assign n_448 = ~x_86 &  x_1074;
assign n_449 =  x_86 & ~x_1074;
assign n_450 = ~x_87 &  x_1075;
assign n_451 =  x_87 & ~x_1075;
assign n_452 = ~x_88 &  x_1076;
assign n_453 =  x_88 & ~x_1076;
assign n_454 = ~x_89 &  x_1077;
assign n_455 =  x_89 & ~x_1077;
assign n_456 = ~x_90 &  x_1078;
assign n_457 =  x_90 & ~x_1078;
assign n_458 = ~x_91 &  x_1079;
assign n_459 =  x_91 & ~x_1079;
assign n_460 = ~x_92 &  x_1080;
assign n_461 =  x_92 & ~x_1080;
assign n_462 = ~x_93 &  x_1081;
assign n_463 =  x_93 & ~x_1081;
assign n_464 = ~x_94 &  x_1082;
assign n_465 =  x_94 & ~x_1082;
assign n_466 = ~x_95 &  x_1083;
assign n_467 =  x_95 & ~x_1083;
assign n_468 = ~x_96 &  x_1084;
assign n_469 =  x_96 & ~x_1084;
assign n_470 = ~x_97 &  x_1085;
assign n_471 =  x_97 & ~x_1085;
assign n_472 = ~x_98 &  x_1086;
assign n_473 =  x_98 & ~x_1086;
assign n_474 = ~x_99 &  x_1087;
assign n_475 =  x_99 & ~x_1087;
assign n_476 = ~x_100 &  x_1088;
assign n_477 =  x_100 & ~x_1088;
assign n_478 = ~x_101 &  x_1089;
assign n_479 =  x_101 & ~x_1089;
assign n_480 = ~x_102 &  x_1090;
assign n_481 =  x_102 & ~x_1090;
assign n_482 = ~x_103 &  x_1091;
assign n_483 =  x_103 & ~x_1091;
assign n_484 = ~x_104 &  x_1092;
assign n_485 =  x_104 & ~x_1092;
assign n_486 = ~x_105 &  x_1093;
assign n_487 =  x_105 & ~x_1093;
assign n_488 = ~x_106 &  x_1094;
assign n_489 = ~n_487 &  n_488;
assign n_490 = ~n_486 & ~n_489;
assign n_491 = ~n_485 & ~n_490;
assign n_492 = ~n_484 & ~n_491;
assign n_493 = ~n_483 & ~n_492;
assign n_494 = ~n_482 & ~n_493;
assign n_495 = ~n_481 & ~n_494;
assign n_496 = ~n_480 & ~n_495;
assign n_497 = ~n_479 & ~n_496;
assign n_498 = ~n_478 & ~n_497;
assign n_499 = ~n_477 & ~n_498;
assign n_500 = ~n_476 & ~n_499;
assign n_501 = ~n_475 & ~n_500;
assign n_502 = ~n_474 & ~n_501;
assign n_503 = ~n_473 & ~n_502;
assign n_504 = ~n_472 & ~n_503;
assign n_505 = ~n_471 & ~n_504;
assign n_506 = ~n_470 & ~n_505;
assign n_507 = ~n_469 & ~n_506;
assign n_508 = ~n_468 & ~n_507;
assign n_509 = ~n_467 & ~n_508;
assign n_510 = ~n_466 & ~n_509;
assign n_511 = ~n_465 & ~n_510;
assign n_512 = ~n_464 & ~n_511;
assign n_513 = ~n_463 & ~n_512;
assign n_514 = ~n_462 & ~n_513;
assign n_515 = ~n_461 & ~n_514;
assign n_516 = ~n_460 & ~n_515;
assign n_517 = ~n_459 & ~n_516;
assign n_518 = ~n_458 & ~n_517;
assign n_519 = ~n_457 & ~n_518;
assign n_520 = ~n_456 & ~n_519;
assign n_521 = ~n_455 & ~n_520;
assign n_522 = ~n_454 & ~n_521;
assign n_523 = ~n_453 & ~n_522;
assign n_524 = ~n_452 & ~n_523;
assign n_525 = ~n_451 & ~n_524;
assign n_526 = ~n_450 & ~n_525;
assign n_527 = ~n_449 & ~n_526;
assign n_528 = ~n_448 & ~n_527;
assign n_529 = ~n_447 & ~n_528;
assign n_530 = ~n_446 & ~n_529;
assign n_531 = ~n_445 & ~n_530;
assign n_532 = ~n_444 & ~n_531;
assign n_533 = ~n_443 & ~n_532;
assign n_534 = ~n_442 & ~n_533;
assign n_535 = ~n_441 & ~n_534;
assign n_536 = ~n_440 & ~n_535;
assign n_537 = ~n_439 & ~n_536;
assign n_538 = ~n_438 & ~n_537;
assign n_539 = ~n_437 & ~n_538;
assign n_540 = ~n_436 & ~n_539;
assign n_541 = ~n_435 & ~n_540;
assign n_542 = ~n_434 & ~n_541;
assign n_543 = ~n_433 & ~n_542;
assign n_544 = ~n_432 & ~n_543;
assign n_545 = ~n_431 & ~n_544;
assign n_546 = ~n_430 & ~n_545;
assign n_547 = ~n_429 & ~n_546;
assign n_548 = ~n_428 & ~n_547;
assign n_549 = ~n_427 & ~n_548;
assign n_550 = ~n_426 & ~n_549;
assign n_551 =  n_550 &  n_284;
assign n_552 =  n_425 &  n_551;
assign n_553 =  x_37 &  x_38;
assign n_554 =  n_291 &  n_553;
assign n_555 =  x_33 &  x_34;
assign n_556 = ~x_35 &  n_555;
assign n_557 = ~x_36 &  n_556;
assign n_558 = ~n_417 &  n_557;
assign n_559 =  n_554 &  n_558;
assign n_560 = ~n_552 & ~n_559;
assign n_561 =  n_420 &  n_560;
assign n_562 =  x_38 & ~x_39;
assign n_563 =  x_40 &  n_562;
assign n_564 =  n_289 &  n_563;
assign n_565 =  x_35 &  x_36;
assign n_566 =  n_282 &  n_565;
assign n_567 = ~x_37 &  n_566;
assign n_568 =  x_75 & ~x_967;
assign n_569 = ~x_75 &  x_967;
assign n_570 = ~x_76 &  x_968;
assign n_571 =  x_76 & ~x_968;
assign n_572 = ~x_77 &  x_969;
assign n_573 =  x_77 & ~x_969;
assign n_574 = ~x_78 &  x_970;
assign n_575 =  x_78 & ~x_970;
assign n_576 = ~x_79 &  x_971;
assign n_577 =  x_79 & ~x_971;
assign n_578 = ~x_80 &  x_972;
assign n_579 =  x_80 & ~x_972;
assign n_580 = ~x_81 &  x_973;
assign n_581 =  x_81 & ~x_973;
assign n_582 = ~x_82 &  x_974;
assign n_583 =  x_82 & ~x_974;
assign n_584 = ~x_83 &  x_975;
assign n_585 =  x_83 & ~x_975;
assign n_586 = ~x_84 &  x_976;
assign n_587 =  x_84 & ~x_976;
assign n_588 = ~x_85 &  x_977;
assign n_589 =  x_85 & ~x_977;
assign n_590 = ~x_86 &  x_978;
assign n_591 =  x_86 & ~x_978;
assign n_592 = ~x_87 &  x_979;
assign n_593 =  x_87 & ~x_979;
assign n_594 = ~x_88 &  x_980;
assign n_595 =  x_88 & ~x_980;
assign n_596 = ~x_89 &  x_981;
assign n_597 =  x_89 & ~x_981;
assign n_598 = ~x_90 &  x_982;
assign n_599 =  x_90 & ~x_982;
assign n_600 = ~x_91 &  x_983;
assign n_601 =  x_91 & ~x_983;
assign n_602 = ~x_92 &  x_984;
assign n_603 =  x_92 & ~x_984;
assign n_604 = ~x_93 &  x_985;
assign n_605 =  x_93 & ~x_985;
assign n_606 = ~x_94 &  x_986;
assign n_607 =  x_94 & ~x_986;
assign n_608 = ~x_95 &  x_987;
assign n_609 =  x_95 & ~x_987;
assign n_610 = ~x_96 &  x_988;
assign n_611 =  x_96 & ~x_988;
assign n_612 = ~x_97 &  x_989;
assign n_613 =  x_97 & ~x_989;
assign n_614 = ~x_98 &  x_990;
assign n_615 =  x_98 & ~x_990;
assign n_616 = ~x_99 &  x_991;
assign n_617 =  x_99 & ~x_991;
assign n_618 = ~x_100 &  x_992;
assign n_619 =  x_100 & ~x_992;
assign n_620 = ~x_101 &  x_993;
assign n_621 =  x_101 & ~x_993;
assign n_622 = ~x_102 &  x_994;
assign n_623 =  x_102 & ~x_994;
assign n_624 = ~x_103 &  x_995;
assign n_625 =  x_103 & ~x_995;
assign n_626 = ~x_104 &  x_996;
assign n_627 =  x_104 & ~x_996;
assign n_628 = ~x_105 &  x_997;
assign n_629 =  x_105 & ~x_997;
assign n_630 = ~x_106 &  x_998;
assign n_631 = ~n_629 &  n_630;
assign n_632 = ~n_628 & ~n_631;
assign n_633 = ~n_627 & ~n_632;
assign n_634 = ~n_626 & ~n_633;
assign n_635 = ~n_625 & ~n_634;
assign n_636 = ~n_624 & ~n_635;
assign n_637 = ~n_623 & ~n_636;
assign n_638 = ~n_622 & ~n_637;
assign n_639 = ~n_621 & ~n_638;
assign n_640 = ~n_620 & ~n_639;
assign n_641 = ~n_619 & ~n_640;
assign n_642 = ~n_618 & ~n_641;
assign n_643 = ~n_617 & ~n_642;
assign n_644 = ~n_616 & ~n_643;
assign n_645 = ~n_615 & ~n_644;
assign n_646 = ~n_614 & ~n_645;
assign n_647 = ~n_613 & ~n_646;
assign n_648 = ~n_612 & ~n_647;
assign n_649 = ~n_611 & ~n_648;
assign n_650 = ~n_610 & ~n_649;
assign n_651 = ~n_609 & ~n_650;
assign n_652 = ~n_608 & ~n_651;
assign n_653 = ~n_607 & ~n_652;
assign n_654 = ~n_606 & ~n_653;
assign n_655 = ~n_605 & ~n_654;
assign n_656 = ~n_604 & ~n_655;
assign n_657 = ~n_603 & ~n_656;
assign n_658 = ~n_602 & ~n_657;
assign n_659 = ~n_601 & ~n_658;
assign n_660 = ~n_600 & ~n_659;
assign n_661 = ~n_599 & ~n_660;
assign n_662 = ~n_598 & ~n_661;
assign n_663 = ~n_597 & ~n_662;
assign n_664 = ~n_596 & ~n_663;
assign n_665 = ~n_595 & ~n_664;
assign n_666 = ~n_594 & ~n_665;
assign n_667 = ~n_593 & ~n_666;
assign n_668 = ~n_592 & ~n_667;
assign n_669 = ~n_591 & ~n_668;
assign n_670 = ~n_590 & ~n_669;
assign n_671 = ~n_589 & ~n_670;
assign n_672 = ~n_588 & ~n_671;
assign n_673 = ~n_587 & ~n_672;
assign n_674 = ~n_586 & ~n_673;
assign n_675 = ~n_585 & ~n_674;
assign n_676 = ~n_584 & ~n_675;
assign n_677 = ~n_583 & ~n_676;
assign n_678 = ~n_582 & ~n_677;
assign n_679 = ~n_581 & ~n_678;
assign n_680 = ~n_580 & ~n_679;
assign n_681 = ~n_579 & ~n_680;
assign n_682 = ~n_578 & ~n_681;
assign n_683 = ~n_577 & ~n_682;
assign n_684 = ~n_576 & ~n_683;
assign n_685 = ~n_575 & ~n_684;
assign n_686 = ~n_574 & ~n_685;
assign n_687 = ~n_573 & ~n_686;
assign n_688 = ~n_572 & ~n_687;
assign n_689 = ~n_571 & ~n_688;
assign n_690 = ~n_570 & ~n_689;
assign n_691 = ~n_569 & ~n_690;
assign n_692 = ~n_568 & ~n_691;
assign n_693 =  n_567 & ~n_692;
assign n_694 =  n_564 &  n_693;
assign n_695 = ~x_38 &  x_39;
assign n_696 =  n_280 &  n_695;
assign n_697 =  n_567 &  n_696;
assign n_698 =  n_550 &  n_697;
assign n_699 = ~n_694 & ~n_698;
assign n_700 = ~x_39 &  n_280;
assign n_701 =  n_700 &  n_286;
assign n_702 = ~x_35 &  x_36;
assign n_703 =  n_282 &  n_702;
assign n_704 =  x_39 &  n_553;
assign n_705 =  n_280 &  n_704;
assign n_706 =  n_703 &  n_705;
assign n_707 = ~n_701 & ~n_706;
assign n_708 =  x_36 & ~x_37;
assign n_709 =  n_556 &  n_708;
assign n_710 =  n_696 &  n_709;
assign n_711 =  n_425 &  n_557;
assign n_712 = ~n_710 & ~n_711;
assign n_713 = ~x_35 &  n_282;
assign n_714 = ~x_36 & ~x_37;
assign n_715 =  n_695 &  n_714;
assign n_716 =  n_713 &  n_715;
assign n_717 =  n_422 &  n_716;
assign n_718 = ~x_38 & ~x_39;
assign n_719 =  n_718 &  n_422;
assign n_720 =  n_567 &  n_719;
assign n_721 = ~n_717 & ~n_720;
assign n_722 =  n_712 &  n_721;
assign n_723 =  n_707 &  n_722;
assign n_724 =  x_38 &  x_39;
assign n_725 = ~x_36 &  n_713;
assign n_726 = ~x_37 &  n_725;
assign n_727 =  n_724 &  n_726;
assign n_728 =  n_422 &  n_727;
assign n_729 = ~x_37 &  n_284;
assign n_730 =  x_38 &  n_281;
assign n_731 =  n_729 &  n_730;
assign n_732 =  x_37 &  n_703;
assign n_733 =  n_732 &  n_562;
assign n_734 =  n_422 &  n_733;
assign n_735 = ~n_731 & ~n_734;
assign n_736 = ~n_728 &  n_735;
assign n_737 =  n_723 &  n_736;
assign n_738 =  n_278 & ~n_737;
assign n_739 = ~x_37 & ~x_38;
assign n_740 =  n_284 &  n_739;
assign n_741 =  n_291 &  n_740;
assign n_742 = ~n_417 &  n_741;
assign n_743 =  n_566 &  n_705;
assign n_744 =  x_41 &  x_42;
assign n_745 =  n_290 &  n_744;
assign n_746 =  n_739 &  n_557;
assign n_747 =  n_745 &  n_746;
assign n_748 = ~n_743 & ~n_747;
assign n_749 =  n_703 &  n_423;
assign n_750 = ~x_39 &  n_749;
assign n_751 =  n_744 &  n_750;
assign n_752 =  n_565 &  n_5;
assign n_753 =  n_553 &  n_752;
assign n_754 = ~x_39 &  n_753;
assign n_755 =  n_744 &  n_754;
assign n_756 = ~n_751 & ~n_755;
assign n_757 =  n_748 &  n_756;
assign n_758 =  n_550 & ~n_757;
assign n_759 = ~n_742 & ~n_758;
assign n_760 = ~n_738 &  n_759;
assign n_761 =  n_699 &  n_760;
assign n_762 =  n_561 &  n_761;
assign n_763 =  x_39 &  x_40;
assign n_764 =  n_744 &  n_763;
assign n_765 =  n_764 &  n_553;
assign n_766 = ~x_39 & ~x_40;
assign n_767 =  n_766 &  n_423;
assign n_768 =  n_744 &  n_767;
assign n_769 = ~n_765 & ~n_768;
assign n_770 =  n_551 & ~n_769;
assign n_771 = ~n_417 &  n_709;
assign n_772 =  n_564 &  n_771;
assign n_773 = ~n_770 & ~n_772;
assign n_774 = ~n_692 &  n_284;
assign n_775 =  x_42 &  n_1;
assign n_776 =  x_39 &  n_775;
assign n_777 =  n_776 &  n_553;
assign n_778 =  n_774 &  n_777;
assign n_779 =  n_291 &  n_746;
assign n_780 = ~n_692 &  n_779;
assign n_781 =  n_289 &  n_766;
assign n_782 =  n_781 &  n_749;
assign n_783 = ~n_692 &  n_782;
assign n_784 = ~n_780 & ~n_783;
assign n_785 = ~n_778 &  n_784;
assign n_786 =  n_773 &  n_785;
assign n_787 =  n_289 &  n_763;
assign n_788 =  n_787 &  n_753;
assign n_789 = ~n_692 &  n_788;
assign n_790 =  n_556 &  n_4;
assign n_791 = ~x_38 &  n_790;
assign n_792 =  n_791 &  n_787;
assign n_793 = ~n_692 &  n_792;
assign n_794 = ~n_789 & ~n_793;
assign n_795 =  n_775 &  n_754;
assign n_796 = ~n_692 &  n_795;
assign n_797 =  n_790 &  n_696;
assign n_798 =  n_278 &  n_797;
assign n_799 = ~n_796 & ~n_798;
assign n_800 =  n_794 &  n_799;
assign n_801 =  n_700 &  n_791;
assign n_802 =  n_550 &  n_801;
assign n_803 =  n_790 &  n_730;
assign n_804 =  n_278 &  n_803;
assign n_805 = ~n_802 & ~n_804;
assign n_806 = ~x_38 &  n_732;
assign n_807 =  n_745 &  n_806;
assign n_808 =  n_807 &  n_278;
assign n_809 =  x_41 & ~x_42;
assign n_810 = ~x_33 & ~x_34;
assign n_811 = ~x_35 &  n_810;
assign n_812 = ~x_36 &  n_811;
assign n_813 =  n_424 &  n_812;
assign n_814 =  x_40 &  n_813;
assign n_815 =  x_37 & ~x_38;
assign n_816 = ~x_39 &  n_815;
assign n_817 =  n_812 &  n_816;
assign n_818 =  x_40 &  n_817;
assign n_819 = ~n_814 & ~n_818;
assign n_820 =  n_809 & ~n_819;
assign n_821 =  n_283 &  n_5;
assign n_822 =  n_739 &  n_821;
assign n_823 =  n_822 &  n_281;
assign n_824 =  n_766 &  n_809;
assign n_825 = ~x_38 &  n_824;
assign n_826 =  n_285 &  n_825;
assign n_827 = ~n_823 & ~n_826;
assign n_828 = ~x_42 &  n_421;
assign n_829 =  n_562 &  n_828;
assign n_830 =  n_790 &  n_829;
assign n_831 =  n_827 & ~n_830;
assign n_832 = ~n_820 &  n_831;
assign n_833 =  n_746 &  n_824;
assign n_834 = ~x_41 & ~x_42;
assign n_835 =  n_763 &  n_834;
assign n_836 =  n_835 &  n_753;
assign n_837 =  x_37 &  n_5;
assign n_838 =  n_702 &  n_837;
assign n_839 = ~x_38 &  n_838;
assign n_840 = ~x_39 &  n_279;
assign n_841 =  n_839 &  n_840;
assign n_842 = ~n_836 & ~n_841;
assign n_843 = ~n_833 &  n_842;
assign n_844 =  n_806 &  n_776;
assign n_845 =  x_1095 &  n_844;
assign n_846 =  n_806 &  n_764;
assign n_847 = ~x_1095 &  n_846;
assign n_848 = ~n_845 & ~n_847;
assign n_849 =  n_843 &  n_848;
assign n_850 =  n_2 &  n_727;
assign n_851 =  n_557 &  n_767;
assign n_852 =  n_834 &  n_851;
assign n_853 =  n_835 &  n_749;
assign n_854 =  n_2 &  n_733;
assign n_855 = ~n_853 & ~n_854;
assign n_856 = ~n_852 &  n_855;
assign n_857 = ~n_850 &  n_856;
assign n_858 =  n_849 &  n_857;
assign n_859 =  n_832 &  n_858;
assign n_860 =  n_725 &  n_553;
assign n_861 =  n_700 &  n_860;
assign n_862 = ~x_776 &  n_861;
assign n_863 = ~x_40 &  n_817;
assign n_864 =  n_834 &  n_863;
assign n_865 =  n_739 &  n_812;
assign n_866 =  n_290 &  n_865;
assign n_867 =  x_42 &  n_866;
assign n_868 = ~n_864 & ~n_867;
assign n_869 = ~n_862 &  n_868;
assign n_870 =  n_860 &  n_787;
assign n_871 =  x_776 &  n_870;
assign n_872 =  n_745 &  n_822;
assign n_873 =  n_708 &  n_6;
assign n_874 =  n_421 &  n_562;
assign n_875 =  n_873 &  n_874;
assign n_876 = ~x_42 &  n_875;
assign n_877 = ~n_872 & ~n_876;
assign n_878 = ~n_871 &  n_877;
assign n_879 = ~x_42 &  n_279;
assign n_880 =  x_39 &  n_879;
assign n_881 =  n_423 &  n_812;
assign n_882 =  n_880 &  n_881;
assign n_883 =  n_752 &  n_815;
assign n_884 =  n_291 &  n_883;
assign n_885 = ~x_39 &  n_2;
assign n_886 =  n_822 &  n_885;
assign n_887 = ~n_884 & ~n_886;
assign n_888 = ~n_882 &  n_887;
assign n_889 =  x_40 & ~x_41;
assign n_890 = ~x_42 &  n_889;
assign n_891 =  n_695 &  n_7;
assign n_892 =  n_718 &  n_708;
assign n_893 =  n_6 &  n_892;
assign n_894 = ~n_891 & ~n_893;
assign n_895 =  n_890 & ~n_894;
assign n_896 =  n_888 & ~n_895;
assign n_897 =  n_878 &  n_896;
assign n_898 =  n_869 &  n_897;
assign n_899 =  n_806 &  n_885;
assign n_900 =  n_763 &  n_809;
assign n_901 =  n_900 &  n_753;
assign n_902 = ~n_899 & ~n_901;
assign n_903 =  n_284 &  n_553;
assign n_904 =  n_903 &  n_880;
assign n_905 = ~x_39 &  n_746;
assign n_906 =  n_2 &  n_905;
assign n_907 = ~n_904 & ~n_906;
assign n_908 =  n_902 &  n_907;
assign n_909 =  n_890 &  n_905;
assign n_910 =  n_2 &  n_750;
assign n_911 =  n_567 &  n_718;
assign n_912 =  n_911 &  n_890;
assign n_913 =  n_562 &  n_890;
assign n_914 =  n_790 &  n_913;
assign n_915 =  n_749 &  n_824;
assign n_916 = ~n_914 & ~n_915;
assign n_917 = ~n_912 &  n_916;
assign n_918 = ~n_910 &  n_917;
assign n_919 = ~n_909 &  n_918;
assign n_920 =  n_908 &  n_919;
assign n_921 =  n_898 &  n_920;
assign n_922 =  n_566 &  n_423;
assign n_923 = ~x_42 &  n_290;
assign n_924 =  n_922 &  n_923;
assign n_925 =  n_567 &  n_825;
assign n_926 = ~n_924 & ~n_925;
assign n_927 =  n_7 &  n_825;
assign n_928 =  n_740 &  n_880;
assign n_929 = ~n_927 & ~n_928;
assign n_930 =  n_926 &  n_929;
assign n_931 =  n_2 &  n_911;
assign n_932 =  x_38 &  n_763;
assign n_933 =  n_834 &  n_932;
assign n_934 =  n_729 &  n_933;
assign n_935 = ~x_38 &  n_835;
assign n_936 =  n_935 &  n_873;
assign n_937 = ~n_934 & ~n_936;
assign n_938 = ~n_931 &  n_937;
assign n_939 =  n_930 &  n_938;
assign n_940 =  x_39 &  n_922;
assign n_941 =  n_940 &  n_890;
assign n_942 =  n_695 &  n_729;
assign n_943 =  n_2 &  n_942;
assign n_944 = ~n_941 & ~n_943;
assign n_945 =  n_715 &  n_811;
assign n_946 = ~x_42 & ~n_889;
assign n_947 =  n_945 &  n_946;
assign n_948 =  n_709 &  n_829;
assign n_949 =  n_889 &  n_811;
assign n_950 =  n_892 &  n_949;
assign n_951 = ~n_948 & ~n_950;
assign n_952 = ~n_947 &  n_951;
assign n_953 =  n_944 &  n_952;
assign n_954 =  n_939 &  n_953;
assign n_955 =  n_822 &  n_880;
assign n_956 =  n_696 &  n_838;
assign n_957 = ~n_955 & ~n_956;
assign n_958 = ~x_38 &  n_3;
assign n_959 =  n_873 &  n_958;
assign n_960 =  n_957 & ~n_959;
assign n_961 =  n_3 &  n_286;
assign n_962 =  n_828 &  n_940;
assign n_963 = ~n_961 & ~n_962;
assign n_964 =  n_960 &  n_963;
assign n_965 =  n_835 &  n_286;
assign n_966 = ~x_41 &  n_923;
assign n_967 =  n_966 &  n_286;
assign n_968 = ~n_965 & ~n_967;
assign n_969 =  n_708 &  n_696;
assign n_970 = ~x_776 &  n_713;
assign n_971 =  n_969 &  n_970;
assign n_972 =  n_283 &  n_837;
assign n_973 = ~x_38 &  n_972;
assign n_974 =  n_764 &  n_973;
assign n_975 = ~n_971 & ~n_974;
assign n_976 =  n_968 &  n_975;
assign n_977 =  n_964 &  n_976;
assign n_978 =  n_954 &  n_977;
assign n_979 =  n_709 &  n_913;
assign n_980 =  n_791 &  n_835;
assign n_981 = ~n_979 & ~n_980;
assign n_982 =  x_776 &  n_922;
assign n_983 =  n_787 &  n_982;
assign n_984 =  n_806 &  n_880;
assign n_985 = ~n_983 & ~n_984;
assign n_986 =  n_981 &  n_985;
assign n_987 =  x_42 &  n_875;
assign n_988 =  n_828 &  n_911;
assign n_989 = ~n_987 & ~n_988;
assign n_990 = ~x_36 &  n_6;
assign n_991 =  n_423 &  n_990;
assign n_992 =  n_835 &  n_991;
assign n_993 =  n_806 &  n_824;
assign n_994 = ~n_992 & ~n_993;
assign n_995 =  n_989 &  n_994;
assign n_996 =  n_986 &  n_995;
assign n_997 =  n_966 &  n_749;
assign n_998 =  n_806 &  n_3;
assign n_999 = ~n_997 & ~n_998;
assign n_1000 = ~x_604 & ~x_605;
assign n_1001 = ~x_606 & ~x_607;
assign n_1002 =  n_1000 &  n_1001;
assign n_1003 = ~x_600 & ~x_601;
assign n_1004 = ~x_602 & ~x_603;
assign n_1005 =  n_1003 &  n_1004;
assign n_1006 =  n_1002 &  n_1005;
assign n_1007 = ~x_612 & ~x_613;
assign n_1008 = ~x_614 & ~x_615;
assign n_1009 =  n_1007 &  n_1008;
assign n_1010 = ~x_608 & ~x_609;
assign n_1011 = ~x_610 & ~x_611;
assign n_1012 =  n_1010 &  n_1011;
assign n_1013 =  n_1009 &  n_1012;
assign n_1014 =  n_1006 &  n_1013;
assign n_1015 = ~x_588 & ~x_589;
assign n_1016 = ~x_590 & ~x_591;
assign n_1017 =  n_1015 &  n_1016;
assign n_1018 = ~x_584 & ~x_585;
assign n_1019 = ~x_586 & ~x_587;
assign n_1020 =  n_1018 &  n_1019;
assign n_1021 =  n_1017 &  n_1020;
assign n_1022 = ~x_596 & ~x_597;
assign n_1023 = ~x_598 & ~x_599;
assign n_1024 =  n_1022 &  n_1023;
assign n_1025 = ~x_592 & ~x_593;
assign n_1026 = ~x_594 & ~x_595;
assign n_1027 =  n_1025 &  n_1026;
assign n_1028 =  n_1024 &  n_1027;
assign n_1029 =  n_1021 &  n_1028;
assign n_1030 =  n_1014 &  n_1029;
assign n_1031 =  n_553 &  n_900;
assign n_1032 =  n_812 &  n_1031;
assign n_1033 =  n_1030 &  n_1032;
assign n_1034 =  n_999 & ~n_1033;
assign n_1035 = ~x_776 &  n_940;
assign n_1036 =  n_422 &  n_1035;
assign n_1037 =  n_835 &  n_860;
assign n_1038 =  n_838 &  n_913;
assign n_1039 =  n_725 &  n_1031;
assign n_1040 = ~n_1038 & ~n_1039;
assign n_1041 = ~n_1037 &  n_1040;
assign n_1042 = ~n_1036 &  n_1041;
assign n_1043 =  n_1034 &  n_1042;
assign n_1044 =  n_996 &  n_1043;
assign n_1045 =  n_978 &  n_1044;
assign n_1046 =  n_921 &  n_1045;
assign n_1047 =  n_859 &  n_1046;
assign n_1048 =  n_822 &  n_835;
assign n_1049 = ~x_700 & ~x_701;
assign n_1050 = ~x_702 & ~x_703;
assign n_1051 =  n_1049 &  n_1050;
assign n_1052 = ~x_696 & ~x_697;
assign n_1053 = ~x_698 & ~x_699;
assign n_1054 =  n_1052 &  n_1053;
assign n_1055 =  n_1051 &  n_1054;
assign n_1056 = ~x_708 & ~x_709;
assign n_1057 = ~x_710 & ~x_711;
assign n_1058 =  n_1056 &  n_1057;
assign n_1059 = ~x_704 & ~x_705;
assign n_1060 = ~x_706 & ~x_707;
assign n_1061 =  n_1059 &  n_1060;
assign n_1062 =  n_1058 &  n_1061;
assign n_1063 =  n_1055 &  n_1062;
assign n_1064 = ~x_684 & ~x_685;
assign n_1065 = ~x_686 & ~x_687;
assign n_1066 =  n_1064 &  n_1065;
assign n_1067 = ~x_680 & ~x_681;
assign n_1068 = ~x_682 & ~x_683;
assign n_1069 =  n_1067 &  n_1068;
assign n_1070 =  n_1066 &  n_1069;
assign n_1071 = ~x_692 & ~x_693;
assign n_1072 = ~x_694 & ~x_695;
assign n_1073 =  n_1071 &  n_1072;
assign n_1074 = ~x_688 & ~x_689;
assign n_1075 = ~x_690 & ~x_691;
assign n_1076 =  n_1074 &  n_1075;
assign n_1077 =  n_1073 &  n_1076;
assign n_1078 =  n_1070 &  n_1077;
assign n_1079 =  n_1063 &  n_1078;
assign n_1080 =  n_1048 &  n_1079;
assign n_1081 =  n_839 &  n_787;
assign n_1082 = ~x_636 & ~x_637;
assign n_1083 = ~x_638 & ~x_639;
assign n_1084 =  n_1082 &  n_1083;
assign n_1085 = ~x_632 & ~x_633;
assign n_1086 = ~x_634 & ~x_635;
assign n_1087 =  n_1085 &  n_1086;
assign n_1088 =  n_1084 &  n_1087;
assign n_1089 = ~x_644 & ~x_645;
assign n_1090 = ~x_646 & ~x_647;
assign n_1091 =  n_1089 &  n_1090;
assign n_1092 = ~x_640 & ~x_641;
assign n_1093 = ~x_642 & ~x_643;
assign n_1094 =  n_1092 &  n_1093;
assign n_1095 =  n_1091 &  n_1094;
assign n_1096 =  n_1088 &  n_1095;
assign n_1097 = ~x_620 & ~x_621;
assign n_1098 = ~x_622 & ~x_623;
assign n_1099 =  n_1097 &  n_1098;
assign n_1100 = ~x_616 & ~x_617;
assign n_1101 = ~x_618 & ~x_619;
assign n_1102 =  n_1100 &  n_1101;
assign n_1103 =  n_1099 &  n_1102;
assign n_1104 = ~x_628 & ~x_629;
assign n_1105 = ~x_630 & ~x_631;
assign n_1106 =  n_1104 &  n_1105;
assign n_1107 = ~x_624 & ~x_625;
assign n_1108 = ~x_626 & ~x_627;
assign n_1109 =  n_1107 &  n_1108;
assign n_1110 =  n_1106 &  n_1109;
assign n_1111 =  n_1103 &  n_1110;
assign n_1112 =  n_1096 &  n_1111;
assign n_1113 =  n_1081 &  n_1112;
assign n_1114 =  n_775 &  n_718;
assign n_1115 =  n_1114 &  n_972;
assign n_1116 = ~x_732 & ~x_733;
assign n_1117 = ~x_734 & ~x_735;
assign n_1118 =  n_1116 &  n_1117;
assign n_1119 = ~x_728 & ~x_729;
assign n_1120 = ~x_730 & ~x_731;
assign n_1121 =  n_1119 &  n_1120;
assign n_1122 =  n_1118 &  n_1121;
assign n_1123 = ~x_740 & ~x_741;
assign n_1124 = ~x_742 & ~x_743;
assign n_1125 =  n_1123 &  n_1124;
assign n_1126 = ~x_736 & ~x_737;
assign n_1127 = ~x_738 & ~x_739;
assign n_1128 =  n_1126 &  n_1127;
assign n_1129 =  n_1125 &  n_1128;
assign n_1130 =  n_1122 &  n_1129;
assign n_1131 = ~x_716 & ~x_717;
assign n_1132 = ~x_718 & ~x_719;
assign n_1133 =  n_1131 &  n_1132;
assign n_1134 = ~x_712 & ~x_713;
assign n_1135 = ~x_714 & ~x_715;
assign n_1136 =  n_1134 &  n_1135;
assign n_1137 =  n_1133 &  n_1136;
assign n_1138 = ~x_724 & ~x_725;
assign n_1139 = ~x_726 & ~x_727;
assign n_1140 =  n_1138 &  n_1139;
assign n_1141 = ~x_720 & ~x_721;
assign n_1142 = ~x_722 & ~x_723;
assign n_1143 =  n_1141 &  n_1142;
assign n_1144 =  n_1140 &  n_1143;
assign n_1145 =  n_1137 &  n_1144;
assign n_1146 =  n_1130 &  n_1145;
assign n_1147 =  n_1115 & ~n_1146;
assign n_1148 =  n_1048 & ~n_1079;
assign n_1149 = ~n_1147 & ~n_1148;
assign n_1150 = ~n_1113 &  n_1149;
assign n_1151 = ~n_1080 &  n_1150;
assign n_1152 = ~x_95 & ~x_96;
assign n_1153 = ~x_97 & ~x_98;
assign n_1154 =  n_1152 &  n_1153;
assign n_1155 = ~x_91 & ~x_92;
assign n_1156 = ~x_93 & ~x_94;
assign n_1157 =  n_1155 &  n_1156;
assign n_1158 =  n_1154 &  n_1157;
assign n_1159 = ~x_103 & ~x_104;
assign n_1160 = ~x_105 & ~x_106;
assign n_1161 =  n_1159 &  n_1160;
assign n_1162 = ~x_99 & ~x_100;
assign n_1163 = ~x_101 & ~x_102;
assign n_1164 =  n_1162 &  n_1163;
assign n_1165 =  n_1161 &  n_1164;
assign n_1166 =  n_1158 &  n_1165;
assign n_1167 = ~x_79 & ~x_80;
assign n_1168 = ~x_81 & ~x_82;
assign n_1169 =  n_1167 &  n_1168;
assign n_1170 = ~x_75 & ~x_76;
assign n_1171 = ~x_77 & ~x_78;
assign n_1172 =  n_1170 &  n_1171;
assign n_1173 =  n_1169 &  n_1172;
assign n_1174 = ~x_87 & ~x_88;
assign n_1175 = ~x_89 & ~x_90;
assign n_1176 =  n_1174 &  n_1175;
assign n_1177 = ~x_83 & ~x_84;
assign n_1178 = ~x_85 & ~x_86;
assign n_1179 =  n_1177 &  n_1178;
assign n_1180 =  n_1176 &  n_1179;
assign n_1181 =  n_1173 &  n_1180;
assign n_1182 =  n_1166 &  n_1181;
assign n_1183 =  n_991 & ~n_1182;
assign n_1184 =  n_745 &  n_1183;
assign n_1185 =  n_922 &  n_3;
assign n_1186 = ~n_1184 & ~n_1185;
assign n_1187 =  n_281 &  n_1183;
assign n_1188 =  n_421 &  n_891;
assign n_1189 = ~n_1188 & ~n_9;
assign n_1190 = ~n_1187 &  n_1189;
assign n_1191 =  n_1186 &  n_1190;
assign n_1192 =  n_1151 &  n_1191;
assign n_1193 =  n_1081 & ~n_1112;
assign n_1194 =  n_553 &  n_812;
assign n_1195 =  n_824 &  n_1194;
assign n_1196 = ~x_540 & ~x_541;
assign n_1197 = ~x_542 & ~x_543;
assign n_1198 =  n_1196 &  n_1197;
assign n_1199 = ~x_536 & ~x_537;
assign n_1200 = ~x_538 & ~x_539;
assign n_1201 =  n_1199 &  n_1200;
assign n_1202 =  n_1198 &  n_1201;
assign n_1203 = ~x_548 & ~x_549;
assign n_1204 = ~x_550 & ~x_551;
assign n_1205 =  n_1203 &  n_1204;
assign n_1206 = ~x_544 & ~x_545;
assign n_1207 = ~x_546 & ~x_547;
assign n_1208 =  n_1206 &  n_1207;
assign n_1209 =  n_1205 &  n_1208;
assign n_1210 =  n_1202 &  n_1209;
assign n_1211 = ~x_524 & ~x_525;
assign n_1212 = ~x_526 & ~x_527;
assign n_1213 =  n_1211 &  n_1212;
assign n_1214 = ~x_520 & ~x_521;
assign n_1215 = ~x_522 & ~x_523;
assign n_1216 =  n_1214 &  n_1215;
assign n_1217 =  n_1213 &  n_1216;
assign n_1218 = ~x_532 & ~x_533;
assign n_1219 = ~x_534 & ~x_535;
assign n_1220 =  n_1218 &  n_1219;
assign n_1221 = ~x_528 & ~x_529;
assign n_1222 = ~x_530 & ~x_531;
assign n_1223 =  n_1221 &  n_1222;
assign n_1224 =  n_1220 &  n_1223;
assign n_1225 =  n_1217 &  n_1224;
assign n_1226 =  n_1210 &  n_1225;
assign n_1227 =  n_1195 & ~n_1226;
assign n_1228 = ~n_1193 & ~n_1227;
assign n_1229 = ~x_39 &  n_883;
assign n_1230 =  n_828 &  n_1229;
assign n_1231 =  n_7 &  n_719;
assign n_1232 = ~x_318 & ~x_319;
assign n_1233 = ~x_320 & ~x_321;
assign n_1234 =  n_1232 &  n_1233;
assign n_1235 = ~x_314 & ~x_315;
assign n_1236 = ~x_316 & ~x_317;
assign n_1237 =  n_1235 &  n_1236;
assign n_1238 =  n_1234 &  n_1237;
assign n_1239 = ~x_326 & ~x_327;
assign n_1240 = ~x_328 & ~x_329;
assign n_1241 =  n_1239 &  n_1240;
assign n_1242 = ~x_322 & ~x_323;
assign n_1243 = ~x_324 & ~x_325;
assign n_1244 =  n_1242 &  n_1243;
assign n_1245 =  n_1241 &  n_1244;
assign n_1246 =  n_1238 &  n_1245;
assign n_1247 = ~x_302 & ~x_303;
assign n_1248 = ~x_304 & ~x_305;
assign n_1249 =  n_1247 &  n_1248;
assign n_1250 = ~x_298 & ~x_299;
assign n_1251 = ~x_300 & ~x_301;
assign n_1252 =  n_1250 &  n_1251;
assign n_1253 =  n_1249 &  n_1252;
assign n_1254 = ~x_310 & ~x_311;
assign n_1255 = ~x_312 & ~x_313;
assign n_1256 =  n_1254 &  n_1255;
assign n_1257 = ~x_306 & ~x_307;
assign n_1258 = ~x_308 & ~x_309;
assign n_1259 =  n_1257 &  n_1258;
assign n_1260 =  n_1256 &  n_1259;
assign n_1261 =  n_1253 &  n_1260;
assign n_1262 =  n_1246 &  n_1261;
assign n_1263 =  n_1231 &  n_1262;
assign n_1264 = ~n_1230 & ~n_1263;
assign n_1265 =  n_809 &  n_863;
assign n_1266 =  n_767 &  n_990;
assign n_1267 =  n_715 &  n_6;
assign n_1268 =  x_40 &  n_1267;
assign n_1269 = ~n_1266 & ~n_1268;
assign n_1270 =  n_809 & ~n_1269;
assign n_1271 = ~n_1265 & ~n_1270;
assign n_1272 =  n_1264 &  n_1271;
assign n_1273 =  n_1228 &  n_1272;
assign n_1274 =  x_39 &  n_881;
assign n_1275 = ~n_893 & ~n_1274;
assign n_1276 = ~n_279 & ~n_889;
assign n_1277 = ~n_1275 &  n_1276;
assign n_1278 =  n_840 &  n_881;
assign n_1279 =  x_39 &  n_889;
assign n_1280 = ~n_766 & ~n_1279;
assign n_1281 =  n_865 & ~n_1280;
assign n_1282 = ~n_1278 & ~n_1281;
assign n_1283 = ~n_1277 &  n_1282;
assign n_1284 = ~x_42 & ~n_1283;
assign n_1285 =  n_1273 & ~n_1284;
assign n_1286 =  n_1192 &  n_1285;
assign n_1287 =  n_739 &  n_752;
assign n_1288 = ~x_39 &  n_1287;
assign n_1289 =  n_828 &  n_1288;
assign n_1290 = ~x_764 & ~x_765;
assign n_1291 = ~x_766 & ~x_767;
assign n_1292 =  n_1290 &  n_1291;
assign n_1293 = ~x_760 & ~x_761;
assign n_1294 = ~x_762 & ~x_763;
assign n_1295 =  n_1293 &  n_1294;
assign n_1296 =  n_1292 &  n_1295;
assign n_1297 = ~x_772 & ~x_773;
assign n_1298 = ~x_774 & ~x_775;
assign n_1299 =  n_1297 &  n_1298;
assign n_1300 = ~x_768 & ~x_769;
assign n_1301 = ~x_770 & ~x_771;
assign n_1302 =  n_1300 &  n_1301;
assign n_1303 =  n_1299 &  n_1302;
assign n_1304 =  n_1296 &  n_1303;
assign n_1305 = ~x_748 & ~x_749;
assign n_1306 = ~x_750 & ~x_751;
assign n_1307 =  n_1305 &  n_1306;
assign n_1308 = ~x_744 & ~x_745;
assign n_1309 = ~x_746 & ~x_747;
assign n_1310 =  n_1308 &  n_1309;
assign n_1311 =  n_1307 &  n_1310;
assign n_1312 = ~x_756 & ~x_757;
assign n_1313 = ~x_758 & ~x_759;
assign n_1314 =  n_1312 &  n_1313;
assign n_1315 = ~x_752 & ~x_753;
assign n_1316 = ~x_754 & ~x_755;
assign n_1317 =  n_1315 &  n_1316;
assign n_1318 =  n_1314 &  n_1317;
assign n_1319 =  n_1311 &  n_1318;
assign n_1320 =  n_1304 &  n_1319;
assign n_1321 =  n_1289 & ~n_1320;
assign n_1322 =  n_1115 &  n_1146;
assign n_1323 = ~n_1321 & ~n_1322;
assign n_1324 =  n_879 &  n_754;
assign n_1325 = ~x_39 &  n_828;
assign n_1326 =  n_746 &  n_1325;
assign n_1327 = ~n_1324 & ~n_1326;
assign n_1328 =  n_745 &  n_973;
assign n_1329 =  n_885 &  n_753;
assign n_1330 = ~n_1328 & ~n_1329;
assign n_1331 =  n_1327 &  n_1330;
assign n_1332 =  n_1323 &  n_1331;
assign n_1333 =  x_39 &  n_991;
assign n_1334 =  n_1 &  n_1333;
assign n_1335 = ~x_39 &  n_889;
assign n_1336 =  n_991 &  n_1335;
assign n_1337 = ~n_1334 & ~n_1336;
assign n_1338 =  n_563 &  n_7;
assign n_1339 = ~x_42 &  n_1338;
assign n_1340 =  n_879 & ~n_894;
assign n_1341 = ~n_1339 & ~n_1340;
assign n_1342 =  n_1337 &  n_1341;
assign n_1343 =  n_1332 &  n_1342;
assign n_1344 = ~n_766 & ~n_763;
assign n_1345 =  n_834 & ~n_1344;
assign n_1346 =  n_881 &  n_1345;
assign n_1347 = ~x_40 & ~x_42;
assign n_1348 =  n_1229 &  n_1347;
assign n_1349 = ~n_1346 & ~n_1348;
assign n_1350 =  n_562 &  n_7;
assign n_1351 =  n_2 &  n_1350;
assign n_1352 =  n_923 &  n_740;
assign n_1353 = ~x_41 &  n_1352;
assign n_1354 = ~n_1351 & ~n_1353;
assign n_1355 =  n_1349 &  n_1354;
assign n_1356 =  n_1 &  n_1267;
assign n_1357 = ~x_42 &  n_1356;
assign n_1358 =  n_739 &  n_990;
assign n_1359 =  n_700 &  n_1358;
assign n_1360 = ~n_1357 & ~n_1359;
assign n_1361 =  n_973 &  n_1325;
assign n_1362 =  n_724 &  n_7;
assign n_1363 =  n_1 &  n_1362;
assign n_1364 = ~n_1361 & ~n_1363;
assign n_1365 =  n_1360 &  n_1364;
assign n_1366 =  n_1355 &  n_1365;
assign n_1367 = ~x_776 &  n_942;
assign n_1368 =  n_422 &  n_1367;
assign n_1369 =  n_700 &  n_922;
assign n_1370 = ~x_776 &  n_1369;
assign n_1371 = ~n_1368 & ~n_1370;
assign n_1372 = ~x_38 &  n_709;
assign n_1373 =  n_1372 &  n_966;
assign n_1374 =  n_1287 &  n_835;
assign n_1375 = ~n_1373 & ~n_1374;
assign n_1376 =  x_776 &  n_942;
assign n_1377 =  n_775 &  n_1376;
assign n_1378 =  n_1375 & ~n_1377;
assign n_1379 =  n_1371 &  n_1378;
assign n_1380 =  n_1366 &  n_1379;
assign n_1381 =  n_1343 &  n_1380;
assign n_1382 =  n_834 & ~n_819;
assign n_1383 =  n_727 &  n_879;
assign n_1384 =  n_1372 &  n_900;
assign n_1385 = ~n_1383 & ~n_1384;
assign n_1386 =  n_1289 &  n_1320;
assign n_1387 =  n_726 &  n_958;
assign n_1388 =  x_40 &  n_695;
assign n_1389 =  n_1388 &  n_809;
assign n_1390 =  n_790 &  n_1389;
assign n_1391 =  n_740 &  n_1325;
assign n_1392 = ~n_1390 & ~n_1391;
assign n_1393 = ~n_1387 &  n_1392;
assign n_1394 = ~n_1386 &  n_1393;
assign n_1395 =  n_1385 &  n_1394;
assign n_1396 = ~n_1382 &  n_1395;
assign n_1397 =  n_280 &  n_1350;
assign n_1398 =  n_809 &  n_1362;
assign n_1399 = ~x_40 &  n_1398;
assign n_1400 = ~n_1397 & ~n_1399;
assign n_1401 =  n_990 &  n_1031;
assign n_1402 =  n_880 &  n_1194;
assign n_1403 = ~n_1401 & ~n_1402;
assign n_1404 =  n_285 &  n_913;
assign n_1405 =  n_3 &  n_903;
assign n_1406 = ~n_1404 & ~n_1405;
assign n_1407 =  n_1403 &  n_1406;
assign n_1408 =  n_1400 &  n_1407;
assign n_1409 =  n_284 &  n_767;
assign n_1410 =  n_834 &  n_1409;
assign n_1411 =  n_286 &  n_880;
assign n_1412 = ~n_1410 & ~n_1411;
assign n_1413 =  n_705 &  n_812;
assign n_1414 =  n_286 &  n_1325;
assign n_1415 = ~n_1413 & ~n_1414;
assign n_1416 =  n_1412 &  n_1415;
assign n_1417 =  n_828 &  n_1333;
assign n_1418 =  n_879 &  n_1267;
assign n_1419 = ~n_1417 & ~n_1418;
assign n_1420 =  n_1416 &  n_1419;
assign n_1421 =  n_1408 &  n_1420;
assign n_1422 =  n_1396 &  n_1421;
assign n_1423 =  n_1381 &  n_1422;
assign n_1424 =  n_1286 &  n_1423;
assign n_1425 =  n_1047 &  n_1424;
assign n_1426 = ~n_808 &  n_1425;
assign n_1427 =  n_805 &  n_1426;
assign n_1428 =  n_800 &  n_1427;
assign n_1429 =  n_786 &  n_1428;
assign n_1430 =  n_732 & ~n_417;
assign n_1431 =  n_1114 &  n_1430;
assign n_1432 =  n_775 &  n_727;
assign n_1433 = ~n_417 &  n_1432;
assign n_1434 = ~n_1431 & ~n_1433;
assign n_1435 =  n_292 &  n_693;
assign n_1436 =  n_744 &  n_1388;
assign n_1437 =  n_285 &  n_1436;
assign n_1438 =  n_278 &  n_1437;
assign n_1439 = ~n_1435 & ~n_1438;
assign n_1440 =  n_1434 &  n_1439;
assign n_1441 =  n_551 &  n_705;
assign n_1442 = ~x_38 &  n_776;
assign n_1443 =  n_1442 &  n_418;
assign n_1444 =  n_775 &  n_905;
assign n_1445 = ~n_692 &  n_1444;
assign n_1446 =  n_567 &  n_1114;
assign n_1447 = ~n_417 &  n_1446;
assign n_1448 = ~n_1445 & ~n_1447;
assign n_1449 = ~n_1443 &  n_1448;
assign n_1450 = ~n_1441 &  n_1449;
assign n_1451 =  n_1440 &  n_1450;
assign n_1452 =  n_1429 &  n_1451;
assign n_1453 =  n_762 &  n_1452;
assign n_1454 =  x_42 & ~n_1453;
assign n_1455 = ~x_42 &  n_1453;
assign n_1456 = ~n_1454 & ~n_1455;
assign n_1457 =  n_567 &  n_692;
assign n_1458 =  n_1457 &  n_564;
assign n_1459 =  n_417 &  n_1432;
assign n_1460 = ~n_1458 & ~n_1459;
assign n_1461 =  n_289 &  n_1388;
assign n_1462 =  n_417 &  n_1461;
assign n_1463 = ~n_1462 & ~n_1442;
assign n_1464 =  n_285 & ~n_1463;
assign n_1465 =  n_1460 & ~n_1464;
assign n_1466 =  n_775 &  n_716;
assign n_1467 =  n_417 &  n_1466;
assign n_1468 = ~n_782 & ~n_789;
assign n_1469 = ~n_1467 &  n_1468;
assign n_1470 =  n_692 &  n_905;
assign n_1471 =  n_289 &  n_1470;
assign n_1472 =  n_417 &  n_709;
assign n_1473 =  n_291 &  n_1472;
assign n_1474 = ~n_1471 & ~n_1473;
assign n_1475 =  n_1469 &  n_1474;
assign n_1476 =  n_1465 &  n_1475;
assign n_1477 =  n_417 &  n_557;
assign n_1478 =  n_1477 &  n_554;
assign n_1479 =  n_775 &  n_424;
assign n_1480 =  n_1477 &  n_1479;
assign n_1481 = ~n_1478 & ~n_1480;
assign n_1482 = ~n_780 & ~n_1445;
assign n_1483 =  n_1481 &  n_1482;
assign n_1484 = ~n_417 &  n_1466;
assign n_1485 = ~n_694 & ~n_1484;
assign n_1486 =  n_1434 &  n_1485;
assign n_1487 =  n_1483 &  n_1486;
assign n_1488 =  n_1476 &  n_1487;
assign n_1489 =  n_1457 &  n_292;
assign n_1490 =  n_732 &  n_417;
assign n_1491 =  x_38 &  n_781;
assign n_1492 =  n_1490 &  n_1491;
assign n_1493 = ~n_1489 & ~n_1492;
assign n_1494 =  n_692 &  n_792;
assign n_1495 =  n_289 &  n_1035;
assign n_1496 = ~x_40 &  n_1495;
assign n_1497 = ~x_223 & ~x_224;
assign n_1498 = ~x_225 & ~x_226;
assign n_1499 =  n_1497 &  n_1498;
assign n_1500 = ~x_219 & ~x_220;
assign n_1501 = ~x_221 & ~x_222;
assign n_1502 =  n_1500 &  n_1501;
assign n_1503 =  n_1499 &  n_1502;
assign n_1504 = ~x_231 & ~x_232;
assign n_1505 = ~x_233 & ~x_234;
assign n_1506 =  n_1504 &  n_1505;
assign n_1507 = ~x_227 & ~x_228;
assign n_1508 = ~x_229 & ~x_230;
assign n_1509 =  n_1507 &  n_1508;
assign n_1510 =  n_1506 &  n_1509;
assign n_1511 =  n_1503 &  n_1510;
assign n_1512 = ~x_207 & ~x_208;
assign n_1513 = ~x_209 & ~x_210;
assign n_1514 =  n_1512 &  n_1513;
assign n_1515 = ~x_203 & ~x_204;
assign n_1516 = ~x_205 & ~x_206;
assign n_1517 =  n_1515 &  n_1516;
assign n_1518 =  n_1514 &  n_1517;
assign n_1519 = ~x_215 & ~x_216;
assign n_1520 = ~x_217 & ~x_218;
assign n_1521 =  n_1519 &  n_1520;
assign n_1522 = ~x_211 & ~x_212;
assign n_1523 = ~x_213 & ~x_214;
assign n_1524 =  n_1522 &  n_1523;
assign n_1525 =  n_1521 &  n_1524;
assign n_1526 =  n_1518 &  n_1525;
assign n_1527 =  n_1511 &  n_1526;
assign n_1528 =  n_959 &  n_1527;
assign n_1529 = ~n_1386 & ~n_1528;
assign n_1530 = ~n_1496 &  n_1529;
assign n_1531 =  n_1288 &  n_890;
assign n_1532 = ~n_1361 & ~n_1531;
assign n_1533 =  n_1327 &  n_1532;
assign n_1534 =  n_972 &  n_935;
assign n_1535 = ~n_974 & ~n_1534;
assign n_1536 =  x_37 &  n_935;
assign n_1537 =  n_812 &  n_1536;
assign n_1538 =  n_1535 & ~n_1537;
assign n_1539 =  n_1533 &  n_1538;
assign n_1540 =  n_1530 &  n_1539;
assign n_1541 = ~n_870 &  n_1040;
assign n_1542 =  n_776 &  n_8;
assign n_1543 = ~n_987 & ~n_1542;
assign n_1544 =  n_1541 &  n_1543;
assign n_1545 =  n_695 &  n_873;
assign n_1546 =  n_280 &  n_1545;
assign n_1547 = ~n_1411 & ~n_1546;
assign n_1548 =  n_708 &  n_564;
assign n_1549 =  n_970 &  n_1548;
assign n_1550 = ~n_1549 & ~n_1188;
assign n_1551 =  n_1547 &  n_1550;
assign n_1552 =  n_1544 &  n_1551;
assign n_1553 =  x_40 &  n_893;
assign n_1554 = ~n_289 & ~n_809;
assign n_1555 =  n_1553 & ~n_1554;
assign n_1556 = ~n_775 & ~n_879;
assign n_1557 =  n_945 & ~n_1556;
assign n_1558 =  n_879 &  n_893;
assign n_1559 = ~n_1557 & ~n_1558;
assign n_1560 =  n_766 & ~n_1554;
assign n_1561 =  n_1560 &  n_865;
assign n_1562 =  n_1559 & ~n_1561;
assign n_1563 = ~n_1555 &  n_1562;
assign n_1564 = ~n_993 & ~n_833;
assign n_1565 =  n_289 &  n_1338;
assign n_1566 =  n_990 &  n_777;
assign n_1567 = ~n_1565 & ~n_1566;
assign n_1568 =  n_1564 &  n_1567;
assign n_1569 =  n_1563 &  n_1568;
assign n_1570 =  n_1552 &  n_1569;
assign n_1571 =  n_1540 &  n_1570;
assign n_1572 =  n_781 &  n_1287;
assign n_1573 = ~n_1572 & ~n_1374;
assign n_1574 =  n_877 &  n_1573;
assign n_1575 =  n_289 & ~n_819;
assign n_1576 =  n_1574 & ~n_1575;
assign n_1577 = ~n_1333 & ~n_1274;
assign n_1578 =  n_828 & ~n_1577;
assign n_1579 =  n_1 &  n_1350;
assign n_1580 = ~n_1336 & ~n_1579;
assign n_1581 =  x_42 & ~n_1580;
assign n_1582 = ~n_1578 & ~n_1581;
assign n_1583 =  n_1576 &  n_1582;
assign n_1584 =  n_1273 &  n_1583;
assign n_1585 =  n_1571 &  n_1584;
assign n_1586 =  n_991 &  n_1279;
assign n_1587 = ~n_1356 & ~n_1586;
assign n_1588 =  x_42 & ~n_1587;
assign n_1589 = ~n_1588 & ~n_1418;
assign n_1590 =  n_289 &  n_863;
assign n_1591 =  n_775 &  n_1333;
assign n_1592 = ~n_1590 & ~n_1591;
assign n_1593 =  n_289 &  n_866;
assign n_1594 =  n_1274 & ~n_1556;
assign n_1595 = ~n_1593 & ~n_1594;
assign n_1596 =  n_1592 &  n_1595;
assign n_1597 =  n_1589 &  n_1596;
assign n_1598 = ~x_508 & ~x_509;
assign n_1599 = ~x_510 & ~x_511;
assign n_1600 =  n_1598 &  n_1599;
assign n_1601 = ~x_504 & ~x_505;
assign n_1602 = ~x_506 & ~x_507;
assign n_1603 =  n_1601 &  n_1602;
assign n_1604 =  n_1600 &  n_1603;
assign n_1605 = ~x_516 & ~x_517;
assign n_1606 = ~x_518 &  x_519;
assign n_1607 =  n_1605 &  n_1606;
assign n_1608 = ~x_512 & ~x_513;
assign n_1609 = ~x_514 & ~x_515;
assign n_1610 =  n_1608 &  n_1609;
assign n_1611 =  n_1607 &  n_1610;
assign n_1612 =  n_1604 &  n_1611;
assign n_1613 = ~x_492 & ~x_493;
assign n_1614 = ~x_494 & ~x_495;
assign n_1615 =  n_1613 &  n_1614;
assign n_1616 = ~x_488 & ~x_489;
assign n_1617 = ~x_490 & ~x_491;
assign n_1618 =  n_1616 &  n_1617;
assign n_1619 =  n_1615 &  n_1618;
assign n_1620 = ~x_500 & ~x_501;
assign n_1621 = ~x_502 & ~x_503;
assign n_1622 =  n_1620 &  n_1621;
assign n_1623 = ~x_496 & ~x_497;
assign n_1624 = ~x_498 & ~x_499;
assign n_1625 =  n_1623 &  n_1624;
assign n_1626 =  n_1622 &  n_1625;
assign n_1627 =  n_1619 &  n_1626;
assign n_1628 =  n_1612 &  n_1627;
assign n_1629 = ~n_1628 &  n_927;
assign n_1630 =  x_42 &  n_889;
assign n_1631 =  n_1362 &  n_1630;
assign n_1632 =  n_1631 &  n_1628;
assign n_1633 = ~n_1629 & ~n_1632;
assign n_1634 =  n_828 &  n_750;
assign n_1635 =  n_1628 &  n_927;
assign n_1636 = ~n_1634 & ~n_1635;
assign n_1637 =  n_1633 &  n_1636;
assign n_1638 =  n_729 &  n_809;
assign n_1639 =  n_563 &  n_1638;
assign n_1640 =  n_883 &  n_1560;
assign n_1641 =  x_776 &  n_713;
assign n_1642 =  n_1548 &  n_1641;
assign n_1643 = ~n_1640 & ~n_1642;
assign n_1644 = ~n_1639 &  n_1643;
assign n_1645 = ~n_1321 &  n_1644;
assign n_1646 =  n_1637 &  n_1645;
assign n_1647 =  n_1597 &  n_1646;
assign n_1648 =  n_775 &  n_1367;
assign n_1649 = ~n_1113 & ~n_1648;
assign n_1650 = ~x_1095 &  n_844;
assign n_1651 = ~n_1413 & ~n_884;
assign n_1652 =  n_957 &  n_1651;
assign n_1653 = ~n_1650 &  n_1652;
assign n_1654 =  n_1649 &  n_1653;
assign n_1655 =  n_764 &  n_822;
assign n_1656 =  n_922 &  n_1325;
assign n_1657 = ~n_1655 & ~n_1656;
assign n_1658 = ~n_936 & ~n_886;
assign n_1659 =  n_1657 &  n_1658;
assign n_1660 = ~n_1048 & ~n_1115;
assign n_1661 =  n_776 &  n_903;
assign n_1662 = ~n_1661 & ~n_915;
assign n_1663 =  n_1660 &  n_1662;
assign n_1664 =  n_1659 &  n_1663;
assign n_1665 =  n_828 &  n_945;
assign n_1666 = ~x_37 &  n_787;
assign n_1667 =  n_812 &  n_1666;
assign n_1668 =  n_7 &  n_1461;
assign n_1669 = ~n_1667 & ~n_1668;
assign n_1670 = ~n_1665 &  n_1669;
assign n_1671 =  n_716 &  n_879;
assign n_1672 = ~n_904 & ~n_1671;
assign n_1673 =  n_702 &  n_555;
assign n_1674 =  n_815 &  n_1673;
assign n_1675 =  n_900 &  n_1674;
assign n_1676 = ~n_1675 & ~n_1391;
assign n_1677 =  n_1672 &  n_1676;
assign n_1678 =  n_1670 &  n_1677;
assign n_1679 =  n_1664 &  n_1678;
assign n_1680 =  n_1654 &  n_1679;
assign n_1681 =  n_885 &  n_1194;
assign n_1682 = ~n_700 & ~n_835;
assign n_1683 =  n_1194 & ~n_1682;
assign n_1684 = ~n_1681 & ~n_1683;
assign n_1685 =  n_1684 &  n_1403;
assign n_1686 = ~n_1030 &  n_1032;
assign n_1687 =  x_41 &  n_1339;
assign n_1688 = ~n_1686 & ~n_1687;
assign n_1689 =  n_1685 &  n_1688;
assign n_1690 =  n_1631 & ~n_1628;
assign n_1691 =  n_289 &  n_1268;
assign n_1692 =  x_42 &  n_950;
assign n_1693 = ~n_1691 & ~n_1692;
assign n_1694 = ~n_1690 &  n_1693;
assign n_1695 =  n_781 &  n_822;
assign n_1696 = ~n_1414 & ~n_1695;
assign n_1697 =  n_1696 & ~n_1399;
assign n_1698 =  n_1694 &  n_1697;
assign n_1699 =  n_1689 &  n_1698;
assign n_1700 =  n_1680 &  n_1699;
assign n_1701 =  n_1647 &  n_1700;
assign n_1702 =  n_851 &  n_809;
assign n_1703 =  n_752 &  n_1536;
assign n_1704 = ~n_1702 & ~n_1703;
assign n_1705 =  n_839 &  n_3;
assign n_1706 = ~n_901 & ~n_9;
assign n_1707 = ~n_1705 &  n_1706;
assign n_1708 =  n_1704 &  n_1707;
assign n_1709 =  n_889 &  n_1545;
assign n_1710 =  x_42 &  n_1709;
assign n_1711 =  n_879 &  n_1350;
assign n_1712 = ~n_1710 & ~n_1711;
assign n_1713 =  x_40 &  n_1495;
assign n_1714 = ~n_745 & ~n_281;
assign n_1715 =  n_1183 & ~n_1714;
assign n_1716 = ~n_1713 & ~n_1715;
assign n_1717 =  n_1712 &  n_1716;
assign n_1718 =  n_1708 &  n_1717;
assign n_1719 = ~n_983 & ~n_962;
assign n_1720 = ~n_1033 &  n_1719;
assign n_1721 =  n_959 & ~n_1527;
assign n_1722 =  n_885 &  n_8;
assign n_1723 =  n_839 &  n_824;
assign n_1724 = ~n_1722 & ~n_1723;
assign n_1725 = ~n_1721 &  n_1724;
assign n_1726 =  n_1720 &  n_1725;
assign n_1727 =  n_1560 &  n_881;
assign n_1728 =  n_1114 &  n_873;
assign n_1729 =  n_880 &  n_8;
assign n_1730 = ~n_1728 & ~n_1729;
assign n_1731 = ~n_1727 &  n_1730;
assign n_1732 =  n_1385 &  n_1731;
assign n_1733 =  n_1726 &  n_1732;
assign n_1734 =  n_832 &  n_1733;
assign n_1735 =  n_1718 &  n_1734;
assign n_1736 =  n_1701 &  n_1735;
assign n_1737 =  n_1585 &  n_1736;
assign n_1738 = ~n_1494 &  n_1737;
assign n_1739 =  n_692 &  n_795;
assign n_1740 =  n_417 &  n_741;
assign n_1741 = ~n_1739 & ~n_1740;
assign n_1742 =  n_1738 &  n_1741;
assign n_1743 =  n_1493 &  n_1742;
assign n_1744 =  n_692 &  n_284;
assign n_1745 =  n_423 &  n_787;
assign n_1746 =  n_1744 &  n_1745;
assign n_1747 =  n_1479 &  n_1744;
assign n_1748 = ~n_1746 & ~n_1747;
assign n_1749 =  n_1490 &  n_1114;
assign n_1750 = ~n_1749 & ~n_742;
assign n_1751 =  n_1748 &  n_1750;
assign n_1752 =  n_1743 &  n_1751;
assign n_1753 =  n_703 &  n_1745;
assign n_1754 =  n_692 &  n_1753;
assign n_1755 =  n_417 &  n_1446;
assign n_1756 = ~n_1754 & ~n_1755;
assign n_1757 =  n_692 &  n_788;
assign n_1758 = ~n_1757 & ~n_796;
assign n_1759 =  n_1479 &  n_558;
assign n_1760 =  n_1758 & ~n_1759;
assign n_1761 =  n_1756 &  n_1760;
assign n_1762 =  n_417 &  n_285;
assign n_1763 =  n_564 &  n_1762;
assign n_1764 =  n_292 &  n_1762;
assign n_1765 = ~n_1763 & ~n_1764;
assign n_1766 = ~n_559 & ~n_419;
assign n_1767 =  n_1765 &  n_1766;
assign n_1768 =  n_1761 &  n_1767;
assign n_1769 =  n_1752 &  n_1768;
assign n_1770 =  n_1488 &  n_1769;
assign n_1771 =  x_41 & ~n_1770;
assign n_1772 = ~x_41 &  n_1770;
assign n_1773 = ~n_1771 & ~n_1772;
assign n_1774 =  n_278 &  n_717;
assign n_1775 = ~n_1437 & ~n_728;
assign n_1776 = ~n_1467 &  n_1775;
assign n_1777 = ~n_1774 &  n_1776;
assign n_1778 = ~n_419 &  n_1777;
assign n_1779 =  n_291 &  n_693;
assign n_1780 =  n_692 &  n_1661;
assign n_1781 = ~n_789 & ~n_1780;
assign n_1782 =  n_775 &  n_1470;
assign n_1783 =  n_1781 & ~n_1782;
assign n_1784 = ~n_1779 &  n_1783;
assign n_1785 =  n_1745 &  n_774;
assign n_1786 =  n_564 &  n_418;
assign n_1787 = ~n_1785 & ~n_1786;
assign n_1788 =  n_1461 &  n_418;
assign n_1789 =  n_692 &  n_782;
assign n_1790 = ~n_793 & ~n_1789;
assign n_1791 = ~n_1788 &  n_1790;
assign n_1792 =  n_1787 &  n_1791;
assign n_1793 =  n_1784 &  n_1792;
assign n_1794 =  n_1778 &  n_1793;
assign n_1795 = ~n_692 &  n_1753;
assign n_1796 =  n_292 &  n_771;
assign n_1797 = ~n_1795 & ~n_1796;
assign n_1798 = ~n_1759 & ~n_1447;
assign n_1799 =  n_1797 &  n_1798;
assign n_1800 =  n_1750 &  n_1799;
assign n_1801 =  n_278 &  n_711;
assign n_1802 =  n_828 &  n_1545;
assign n_1803 = ~n_1695 & ~n_1802;
assign n_1804 =  n_1330 &  n_1803;
assign n_1805 = ~n_425 & ~n_765;
assign n_1806 =  n_284 & ~n_1805;
assign n_1807 = ~n_1579 & ~n_1806;
assign n_1808 =  n_776 &  n_286;
assign n_1809 =  n_1559 & ~n_1808;
assign n_1810 =  n_1807 &  n_1809;
assign n_1811 =  n_1804 &  n_1810;
assign n_1812 =  n_932 &  n_1638;
assign n_1813 = ~n_1690 & ~n_1812;
assign n_1814 =  n_1813 &  n_1323;
assign n_1815 =  n_1811 &  n_1814;
assign n_1816 = ~n_807 & ~n_998;
assign n_1817 =  n_809 &  n_1266;
assign n_1818 = ~n_734 & ~n_1817;
assign n_1819 =  n_1816 &  n_1818;
assign n_1820 = ~n_1374 & ~n_1038;
assign n_1821 = ~n_872 & ~n_884;
assign n_1822 =  n_1820 &  n_1821;
assign n_1823 = ~n_943 & ~n_910;
assign n_1824 =  n_1822 &  n_1823;
assign n_1825 =  n_1819 &  n_1824;
assign n_1826 =  n_764 &  n_991;
assign n_1827 = ~n_1826 & ~n_1681;
assign n_1828 =  n_749 &  n_900;
assign n_1829 = ~n_925 & ~n_1828;
assign n_1830 = ~n_1402 &  n_1829;
assign n_1831 =  n_1827 &  n_1830;
assign n_1832 = ~n_422 & ~n_2;
assign n_1833 =  n_1229 & ~n_1832;
assign n_1834 =  n_286 &  n_900;
assign n_1835 = ~n_1833 & ~n_1834;
assign n_1836 = ~n_1692 & ~n_833;
assign n_1837 =  n_1835 &  n_1836;
assign n_1838 =  n_1831 &  n_1837;
assign n_1839 =  n_1825 &  n_1838;
assign n_1840 =  n_1815 &  n_1839;
assign n_1841 = ~x_40 &  n_1362;
assign n_1842 = ~x_42 &  n_1841;
assign n_1843 = ~n_1566 & ~n_1842;
assign n_1844 =  n_1372 &  n_1325;
assign n_1845 = ~n_745 & ~n_885;
assign n_1846 =  n_881 & ~n_1845;
assign n_1847 = ~n_1844 & ~n_1846;
assign n_1848 = ~n_1187 &  n_1847;
assign n_1849 =  n_1843 &  n_1848;
assign n_1850 =  x_40 &  n_755;
assign n_1851 =  n_423 &  n_752;
assign n_1852 =  n_3 &  n_1851;
assign n_1853 = ~n_1850 & ~n_1852;
assign n_1854 =  n_766 &  n_865;
assign n_1855 = ~n_863 & ~n_1854;
assign n_1856 = ~n_744 & ~n_1855;
assign n_1857 =  n_1853 & ~n_1856;
assign n_1858 =  x_41 &  n_818;
assign n_1859 =  x_42 &  n_1858;
assign n_1860 =  n_1394 & ~n_1859;
assign n_1861 =  n_1857 &  n_1860;
assign n_1862 =  n_1849 &  n_1861;
assign n_1863 =  n_1840 &  n_1862;
assign n_1864 =  n_2 &  n_893;
assign n_1865 = ~n_1542 & ~n_1864;
assign n_1866 = ~n_1414 &  n_1865;
assign n_1867 =  n_989 &  n_1866;
assign n_1868 = ~x_191 & ~x_192;
assign n_1869 = ~x_193 & ~x_194;
assign n_1870 =  n_1868 &  n_1869;
assign n_1871 = ~x_187 & ~x_188;
assign n_1872 = ~x_189 & ~x_190;
assign n_1873 =  n_1871 &  n_1872;
assign n_1874 =  n_1870 &  n_1873;
assign n_1875 = ~x_199 & ~x_200;
assign n_1876 = ~x_201 & ~x_202;
assign n_1877 =  n_1875 &  n_1876;
assign n_1878 = ~x_195 & ~x_196;
assign n_1879 = ~x_197 & ~x_198;
assign n_1880 =  n_1878 &  n_1879;
assign n_1881 =  n_1877 &  n_1880;
assign n_1882 =  n_1874 &  n_1881;
assign n_1883 = ~x_175 & ~x_176;
assign n_1884 = ~x_177 & ~x_178;
assign n_1885 =  n_1883 &  n_1884;
assign n_1886 = ~x_171 & ~x_172;
assign n_1887 = ~x_173 & ~x_174;
assign n_1888 =  n_1886 &  n_1887;
assign n_1889 =  n_1885 &  n_1888;
assign n_1890 = ~x_183 & ~x_184;
assign n_1891 = ~x_185 & ~x_186;
assign n_1892 =  n_1890 &  n_1891;
assign n_1893 = ~x_179 & ~x_180;
assign n_1894 = ~x_181 & ~x_182;
assign n_1895 =  n_1893 &  n_1894;
assign n_1896 =  n_1892 &  n_1895;
assign n_1897 =  n_1889 &  n_1896;
assign n_1898 =  n_1882 &  n_1897;
assign n_1899 =  n_1691 &  n_1898;
assign n_1900 = ~n_1188 & ~n_961;
assign n_1901 = ~n_1899 &  n_1900;
assign n_1902 = ~n_893 & ~n_945;
assign n_1903 = ~n_750 &  n_1902;
assign n_1904 =  n_422 & ~n_1903;
assign n_1905 = ~n_1338 & ~n_1268;
assign n_1906 =  n_744 & ~n_1905;
assign n_1907 = ~n_1904 & ~n_1906;
assign n_1908 =  n_1901 &  n_1907;
assign n_1909 =  n_1867 &  n_1908;
assign n_1910 = ~n_931 & ~n_1496;
assign n_1911 = ~x_796 & ~x_797;
assign n_1912 = ~x_798 & ~x_799;
assign n_1913 =  n_1911 &  n_1912;
assign n_1914 = ~x_792 & ~x_793;
assign n_1915 = ~x_794 & ~x_795;
assign n_1916 =  n_1914 &  n_1915;
assign n_1917 =  n_1913 &  n_1916;
assign n_1918 = ~x_804 & ~x_805;
assign n_1919 = ~x_806 & ~x_807;
assign n_1920 =  n_1918 &  n_1919;
assign n_1921 = ~x_800 & ~x_801;
assign n_1922 = ~x_802 & ~x_803;
assign n_1923 =  n_1921 &  n_1922;
assign n_1924 =  n_1920 &  n_1923;
assign n_1925 =  n_1917 &  n_1924;
assign n_1926 = ~x_780 & ~x_781;
assign n_1927 = ~x_782 & ~x_783;
assign n_1928 =  n_1926 &  n_1927;
assign n_1929 = ~x_776 & ~x_777;
assign n_1930 = ~x_778 & ~x_779;
assign n_1931 =  n_1929 &  n_1930;
assign n_1932 =  n_1928 &  n_1931;
assign n_1933 = ~x_788 & ~x_789;
assign n_1934 = ~x_790 & ~x_791;
assign n_1935 =  n_1933 &  n_1934;
assign n_1936 = ~x_784 & ~x_785;
assign n_1937 = ~x_786 & ~x_787;
assign n_1938 =  n_1936 &  n_1937;
assign n_1939 =  n_1935 &  n_1938;
assign n_1940 =  n_1932 &  n_1939;
assign n_1941 =  n_1925 &  n_1940;
assign n_1942 =  x_34 &  x_37;
assign n_1943 =  n_565 &  n_1942;
assign n_1944 = ~x_34 & ~x_35;
assign n_1945 =  n_4 &  n_1944;
assign n_1946 = ~n_1943 & ~n_1945;
assign n_1947 = ~x_33 &  n_695;
assign n_1948 =  n_828 &  n_1947;
assign n_1949 = ~n_1946 &  n_1948;
assign n_1950 = ~n_1941 &  n_1949;
assign n_1951 =  n_1287 &  n_787;
assign n_1952 =  n_991 & ~n_1714;
assign n_1953 =  n_1182 &  n_1952;
assign n_1954 = ~n_1951 & ~n_1953;
assign n_1955 = ~n_1950 &  n_1954;
assign n_1956 =  n_1910 &  n_1955;
assign n_1957 =  n_1909 &  n_1956;
assign n_1958 = ~n_850 & ~n_1033;
assign n_1959 = ~n_876 & ~n_854;
assign n_1960 =  n_902 &  n_1959;
assign n_1961 =  n_1958 &  n_1960;
assign n_1962 =  n_2 &  n_945;
assign n_1963 =  n_285 &  n_829;
assign n_1964 =  n_990 &  n_765;
assign n_1965 = ~n_1963 & ~n_1964;
assign n_1966 = ~n_1962 &  n_1965;
assign n_1967 = ~n_1356 & ~n_1418;
assign n_1968 = ~n_1656 & ~n_1231;
assign n_1969 =  n_1967 &  n_1968;
assign n_1970 =  n_1966 &  n_1969;
assign n_1971 = ~n_1148 &  n_1535;
assign n_1972 =  n_1970 &  n_1971;
assign n_1973 =  n_1961 &  n_1972;
assign n_1974 = ~n_1702 & ~n_1640;
assign n_1975 = ~n_1334 &  n_1974;
assign n_1976 =  n_1724 &  n_1412;
assign n_1977 =  n_1975 &  n_1976;
assign n_1978 = ~n_906 & ~n_1432;
assign n_1979 = ~n_852 & ~n_747;
assign n_1980 = ~n_1635 &  n_1979;
assign n_1981 =  n_1978 &  n_1980;
assign n_1982 =  n_1977 &  n_1981;
assign n_1983 =  n_1973 &  n_1982;
assign n_1984 =  n_1957 &  n_1983;
assign n_1985 =  n_764 &  n_982;
assign n_1986 = ~n_1036 & ~n_1985;
assign n_1987 =  n_1186 &  n_1986;
assign n_1988 = ~n_1 & ~n_422;
assign n_1989 = ~n_879 &  n_1988;
assign n_1990 =  n_1274 & ~n_1989;
assign n_1991 =  n_1987 & ~n_1990;
assign n_1992 = ~n_1686 &  n_1228;
assign n_1993 = ~n_846 & ~n_1650;
assign n_1994 =  n_1993 & ~n_1675;
assign n_1995 =  n_1992 &  n_1994;
assign n_1996 =  n_422 &  n_1376;
assign n_1997 = ~n_1648 & ~n_1996;
assign n_1998 = ~n_1368 & ~n_1405;
assign n_1999 =  n_1997 &  n_1998;
assign n_2000 =  n_1999 &  n_1732;
assign n_2001 =  n_1995 &  n_2000;
assign n_2002 =  n_1991 &  n_2001;
assign n_2003 =  n_1984 &  n_2002;
assign n_2004 =  n_1863 &  n_2003;
assign n_2005 = ~n_1801 &  n_2004;
assign n_2006 = ~n_1492 &  n_2005;
assign n_2007 = ~n_1480 & ~n_1747;
assign n_2008 =  n_2006 &  n_2007;
assign n_2009 = ~n_278 &  n_711;
assign n_2010 = ~n_1755 & ~n_720;
assign n_2011 = ~n_2009 &  n_2010;
assign n_2012 = ~n_278 &  n_717;
assign n_2013 = ~n_1445 & ~n_1739;
assign n_2014 = ~n_2012 &  n_2013;
assign n_2015 =  n_2011 &  n_2014;
assign n_2016 =  n_2008 &  n_2015;
assign n_2017 =  n_1800 &  n_2016;
assign n_2018 =  n_1794 &  n_2017;
assign n_2019 =  x_40 &  n_2018;
assign n_2020 = ~x_40 & ~n_2018;
assign n_2021 = ~n_2019 & ~n_2020;
assign n_2022 =  n_1797 & ~n_772;
assign n_2023 = ~n_1746 &  n_1758;
assign n_2024 = ~n_550 &  n_284;
assign n_2025 =  n_2024 & ~n_769;
assign n_2026 = ~n_2025 &  n_1448;
assign n_2027 =  n_2023 &  n_2026;
assign n_2028 =  n_2022 &  n_2027;
assign n_2029 =  n_1778 &  n_2028;
assign n_2030 = ~n_1464 & ~n_1788;
assign n_2031 =  n_1479 &  n_774;
assign n_2032 = ~n_701 & ~n_2031;
assign n_2033 = ~n_1786 &  n_2032;
assign n_2034 =  n_2030 &  n_2033;
assign n_2035 = ~n_801 & ~n_1494;
assign n_2036 = ~n_1780 &  n_2035;
assign n_2037 =  n_280 &  n_750;
assign n_2038 = ~n_2012 & ~n_2037;
assign n_2039 =  n_1986 & ~n_1413;
assign n_2040 = ~n_1148 & ~n_1721;
assign n_2041 =  n_2039 &  n_2040;
assign n_2042 =  n_1 & ~n_1577;
assign n_2043 = ~n_2042 &  n_1574;
assign n_2044 =  n_1419 &  n_1385;
assign n_2045 =  n_2043 &  n_2044;
assign n_2046 = ~n_1377 & ~n_1802;
assign n_2047 =  n_2046 &  n_1712;
assign n_2048 = ~n_1542 & ~n_836;
assign n_2049 =  n_8 &  n_1279;
assign n_2050 =  n_700 &  n_839;
assign n_2051 = ~n_2049 & ~n_2050;
assign n_2052 =  n_2048 &  n_2051;
assign n_2053 =  n_2052 &  n_1843;
assign n_2054 =  n_2047 &  n_2053;
assign n_2055 =  n_2045 &  n_2054;
assign n_2056 =  n_2041 &  n_2055;
assign n_2057 = ~n_861 &  n_1829;
assign n_2058 =  n_1041 &  n_2057;
assign n_2059 = ~n_1686 &  n_2058;
assign n_2060 =  n_744 &  n_863;
assign n_2061 =  n_1900 & ~n_2060;
assign n_2062 =  n_1691 & ~n_1898;
assign n_2063 = ~n_2062 &  n_888;
assign n_2064 =  n_2061 &  n_2063;
assign n_2065 =  n_2059 &  n_2064;
assign n_2066 =  n_1994 &  n_1999;
assign n_2067 =  n_2065 &  n_2066;
assign n_2068 = ~n_936 & ~n_1387;
assign n_2069 =  n_2068 & ~n_1432;
assign n_2070 =  n_700 &  n_8;
assign n_2071 = ~n_2070 & ~n_1963;
assign n_2072 = ~n_1690 &  n_2071;
assign n_2073 =  n_2069 &  n_2072;
assign n_2074 = ~n_1080 & ~n_1495;
assign n_2075 =  n_944 & ~n_1322;
assign n_2076 =  n_2074 &  n_2075;
assign n_2077 =  n_2073 &  n_2076;
assign n_2078 = ~n_1185 & ~n_998;
assign n_2079 =  n_2078 &  n_1403;
assign n_2080 =  n_1195 &  n_1226;
assign n_2081 =  n_744 &  n_1854;
assign n_2082 = ~n_2080 & ~n_2081;
assign n_2083 =  n_2079 &  n_2082;
assign n_2084 =  n_809 &  n_1268;
assign n_2085 =  n_280 &  n_1229;
assign n_2086 = ~n_2084 & ~n_2085;
assign n_2087 = ~n_928 & ~n_833;
assign n_2088 =  n_2086 &  n_2087;
assign n_2089 = ~n_1397 & ~n_1826;
assign n_2090 = ~n_1359 & ~n_1703;
assign n_2091 =  n_2089 &  n_2090;
assign n_2092 =  n_2088 &  n_2091;
assign n_2093 =  n_2083 &  n_2092;
assign n_2094 =  n_2077 &  n_2093;
assign n_2095 = ~n_934 & ~n_1655;
assign n_2096 = ~n_1705 &  n_2095;
assign n_2097 = ~n_850 &  n_2096;
assign n_2098 = ~n_1729 & ~n_1537;
assign n_2099 =  n_763 &  n_881;
assign n_2100 =  n_280 &  n_813;
assign n_2101 = ~n_2099 & ~n_2100;
assign n_2102 =  n_2098 &  n_2101;
assign n_2103 =  n_2097 &  n_2102;
assign n_2104 =  n_744 & ~n_1269;
assign n_2105 =  n_1409 &  n_809;
assign n_2106 = ~n_2105 & ~n_1834;
assign n_2107 = ~n_2104 &  n_2106;
assign n_2108 =  n_2107 &  n_1633;
assign n_2109 =  n_2103 &  n_2108;
assign n_2110 = ~n_870 & ~n_965;
assign n_2111 = ~n_1289 & ~n_980;
assign n_2112 =  n_2110 &  n_2111;
assign n_2113 = ~n_1356 & ~n_826;
assign n_2114 = ~n_280 &  n_945;
assign n_2115 = ~n_1964 & ~n_2114;
assign n_2116 =  n_2113 &  n_2115;
assign n_2117 = ~n_1369 & ~n_955;
assign n_2118 =  n_700 &  n_753;
assign n_2119 = ~n_853 & ~n_2118;
assign n_2120 =  n_2117 &  n_2119;
assign n_2121 =  n_2116 &  n_2120;
assign n_2122 =  n_2112 &  n_2121;
assign n_2123 =  n_716 &  n_828;
assign n_2124 = ~n_2123 & ~n_948;
assign n_2125 =  n_822 &  n_824;
assign n_2126 =  n_280 &  n_893;
assign n_2127 = ~n_2125 & ~n_2126;
assign n_2128 =  n_2124 &  n_2127;
assign n_2129 = ~n_1324 & ~n_1683;
assign n_2130 =  n_2128 &  n_2129;
assign n_2131 = ~n_1411 & ~n_1586;
assign n_2132 = ~n_1844 & ~n_1414;
assign n_2133 =  n_2131 &  n_2132;
assign n_2134 =  n_2130 &  n_2133;
assign n_2135 =  n_2122 &  n_2134;
assign n_2136 =  n_2109 &  n_2135;
assign n_2137 =  n_2094 &  n_2136;
assign n_2138 =  n_2067 &  n_2137;
assign n_2139 =  n_2056 &  n_2138;
assign n_2140 = ~n_1754 &  n_2139;
assign n_2141 = ~n_770 &  n_2140;
assign n_2142 =  n_2038 &  n_2141;
assign n_2143 =  n_2036 &  n_2142;
assign n_2144 =  n_2034 &  n_2143;
assign n_2145 =  n_2029 &  n_2144;
assign n_2146 =  x_39 & ~n_2145;
assign n_2147 = ~x_39 &  n_2145;
assign n_2148 = ~n_2146 & ~n_2147;
assign n_2149 =  n_564 &  n_1472;
assign n_2150 = ~n_278 &  n_797;
assign n_2151 = ~n_780 & ~n_2150;
assign n_2152 = ~n_2149 &  n_2151;
assign n_2153 =  n_1781 & ~n_1443;
assign n_2154 =  n_2152 &  n_2153;
assign n_2155 = ~n_278 &  n_287;
assign n_2156 =  n_421 &  n_1362;
assign n_2157 =  n_281 &  n_1358;
assign n_2158 = ~n_2156 & ~n_2157;
assign n_2159 = ~n_1417 &  n_2158;
assign n_2160 =  n_2089 &  n_2159;
assign n_2161 =  n_1337 &  n_2160;
assign n_2162 = ~n_1326 & ~n_1329;
assign n_2163 = ~n_941 & ~n_997;
assign n_2164 =  n_2162 &  n_2163;
assign n_2165 =  n_2164 &  n_1416;
assign n_2166 =  n_1853 &  n_2165;
assign n_2167 =  n_2161 &  n_2166;
assign n_2168 =  n_1684 &  n_1955;
assign n_2169 =  n_2168 &  n_1849;
assign n_2170 =  n_2167 &  n_2169;
assign n_2171 = ~n_744 &  n_2099;
assign n_2172 = ~x_776 &  n_870;
assign n_2173 = ~n_2080 & ~n_2172;
assign n_2174 = ~n_2171 &  n_2173;
assign n_2175 =  n_879 &  n_733;
assign n_2176 = ~n_2175 & ~n_1631;
assign n_2177 =  n_2176 & ~n_1263;
assign n_2178 = ~n_744 &  n_814;
assign n_2179 = ~n_2178 & ~n_1899;
assign n_2180 =  n_2177 &  n_2179;
assign n_2181 =  n_2174 &  n_2180;
assign n_2182 = ~n_1404 & ~n_1713;
assign n_2183 = ~n_1033 & ~n_959;
assign n_2184 = ~n_1496 &  n_2183;
assign n_2185 =  n_2182 &  n_2184;
assign n_2186 =  n_2181 &  n_2185;
assign n_2187 = ~n_934 & ~n_915;
assign n_2188 =  n_2187 & ~n_1402;
assign n_2189 = ~n_872 & ~n_914;
assign n_2190 =  n_2189 & ~n_1727;
assign n_2191 =  n_2188 &  n_2190;
assign n_2192 = ~n_861 & ~n_1037;
assign n_2193 =  n_280 &  n_891;
assign n_2194 = ~n_1586 & ~n_2193;
assign n_2195 =  n_2192 &  n_2194;
assign n_2196 =  n_2191 &  n_2195;
assign n_2197 =  x_41 &  n_1266;
assign n_2198 = ~n_2197 & ~n_1579;
assign n_2199 =  n_281 &  n_865;
assign n_2200 = ~n_2199 & ~n_2100;
assign n_2201 =  n_2198 &  n_2200;
assign n_2202 =  n_1149 &  n_2201;
assign n_2203 =  n_2196 &  n_2202;
assign n_2204 = ~n_971 & ~n_1549;
assign n_2205 = ~n_1639 & ~n_836;
assign n_2206 =  n_2204 &  n_2205;
assign n_2207 = ~n_956 & ~n_910;
assign n_2208 = ~n_751 & ~n_697;
assign n_2209 =  n_2207 &  n_2208;
assign n_2210 =  n_2206 &  n_2209;
assign n_2211 = ~n_955 & ~n_710;
assign n_2212 = ~n_782 & ~n_1338;
assign n_2213 =  n_2211 &  n_2212;
assign n_2214 = ~n_1369 & ~n_1038;
assign n_2215 = ~n_901 & ~n_979;
assign n_2216 =  n_2214 &  n_2215;
assign n_2217 =  n_2213 &  n_2216;
assign n_2218 = ~n_1405 & ~n_1546;
assign n_2219 =  n_922 &  n_966;
assign n_2220 = ~n_830 & ~n_2219;
assign n_2221 = ~n_1391 &  n_2220;
assign n_2222 =  n_2218 &  n_2221;
assign n_2223 =  n_2217 &  n_2222;
assign n_2224 =  n_2210 &  n_2223;
assign n_2225 =  n_2203 &  n_2224;
assign n_2226 =  n_2186 &  n_2225;
assign n_2227 =  n_969 &  n_1641;
assign n_2228 = ~n_1322 & ~n_2227;
assign n_2229 = ~n_728 & ~n_1386;
assign n_2230 =  n_2228 &  n_2229;
assign n_2231 =  n_2230 &  n_857;
assign n_2232 =  n_1992 &  n_2231;
assign n_2233 =  n_1991 &  n_2232;
assign n_2234 =  n_2226 &  n_2233;
assign n_2235 =  n_2170 &  n_2234;
assign n_2236 = ~n_2155 &  n_2235;
assign n_2237 = ~n_2009 & ~n_742;
assign n_2238 =  n_2236 &  n_2237;
assign n_2239 =  n_1491 &  n_1430;
assign n_2240 = ~n_1796 & ~n_2239;
assign n_2241 =  n_2238 &  n_2240;
assign n_2242 =  n_2154 &  n_2241;
assign n_2243 =  n_2024 &  n_765;
assign n_2244 = ~n_2243 & ~n_1763;
assign n_2245 = ~n_425 & ~n_768;
assign n_2246 =  n_2024 & ~n_2245;
assign n_2247 = ~n_2246 & ~n_770;
assign n_2248 =  n_2244 &  n_2247;
assign n_2249 =  n_550 &  n_2118;
assign n_2250 = ~n_550 &  n_2118;
assign n_2251 = ~n_1739 & ~n_2250;
assign n_2252 = ~n_1757 &  n_2251;
assign n_2253 = ~n_2249 &  n_2252;
assign n_2254 =  n_2248 &  n_2253;
assign n_2255 =  n_2242 &  n_2254;
assign n_2256 = ~n_1801 & ~n_734;
assign n_2257 = ~n_1754 &  n_2256;
assign n_2258 =  n_1748 &  n_2257;
assign n_2259 =  n_1481 &  n_2258;
assign n_2260 = ~n_1492 & ~n_798;
assign n_2261 =  n_1460 &  n_2260;
assign n_2262 =  n_2261 &  n_561;
assign n_2263 =  n_2259 &  n_2262;
assign n_2264 =  n_2255 &  n_2263;
assign n_2265 =  x_38 & ~n_2264;
assign n_2266 = ~x_38 &  n_2264;
assign n_2267 = ~n_2265 & ~n_2266;
assign n_2268 = ~n_2155 & ~n_1764;
assign n_2269 =  n_2268 & ~n_419;
assign n_2270 =  n_551 &  n_765;
assign n_2271 = ~n_278 &  n_1437;
assign n_2272 = ~n_288 & ~n_2271;
assign n_2273 =  n_2272 &  n_2151;
assign n_2274 = ~n_2270 &  n_2273;
assign n_2275 = ~n_1478 & ~n_694;
assign n_2276 = ~n_550 &  n_1850;
assign n_2277 = ~n_2249 & ~n_2276;
assign n_2278 =  n_2277 & ~n_2239;
assign n_2279 =  n_2275 &  n_2278;
assign n_2280 =  n_2274 &  n_2279;
assign n_2281 =  n_2269 &  n_2280;
assign n_2282 =  n_2252 &  n_2036;
assign n_2283 =  n_2260 &  n_2282;
assign n_2284 =  n_550 &  n_1850;
assign n_2285 = ~n_1795 & ~n_2284;
assign n_2286 = ~n_1438 &  n_2285;
assign n_2287 =  n_806 &  n_2;
assign n_2288 = ~n_2287 &  n_2189;
assign n_2289 = ~n_1729 & ~n_1363;
assign n_2290 =  n_2288 &  n_2289;
assign n_2291 =  n_1993 &  n_2290;
assign n_2292 = ~n_1193 & ~n_1231;
assign n_2293 =  n_2292 &  n_2052;
assign n_2294 =  n_2291 &  n_2293;
assign n_2295 = ~n_956 & ~n_927;
assign n_2296 =  n_827 &  n_2295;
assign n_2297 =  n_2296 &  n_2110;
assign n_2298 = ~n_817 & ~n_1964;
assign n_2299 =  n_1436 &  n_7;
assign n_2300 = ~n_2299 & ~n_1852;
assign n_2301 =  n_2298 &  n_2300;
assign n_2302 = ~n_1113 &  n_2301;
assign n_2303 =  n_2297 &  n_2302;
assign n_2304 =  n_1350 & ~n_1988;
assign n_2305 = ~n_1339 & ~n_2304;
assign n_2306 = ~n_889 &  n_1229;
assign n_2307 = ~n_2306 & ~n_1195;
assign n_2308 =  n_2305 &  n_2307;
assign n_2309 = ~n_807 & ~n_1328;
assign n_2310 = ~n_1414 & ~n_1642;
assign n_2311 =  n_2309 &  n_2310;
assign n_2312 =  n_2308 &  n_2311;
assign n_2313 =  n_2303 &  n_2312;
assign n_2314 =  n_2294 &  n_2313;
assign n_2315 =  n_1538 &  n_1408;
assign n_2316 =  n_2168 &  n_2315;
assign n_2317 =  n_2314 &  n_2316;
assign n_2318 = ~n_886 & ~n_961;
assign n_2319 = ~n_1361 & ~n_1671;
assign n_2320 =  n_2318 &  n_2319;
assign n_2321 = ~n_1634 & ~n_984;
assign n_2322 =  n_2106 &  n_2321;
assign n_2323 =  n_2320 &  n_2322;
assign n_2324 =  n_2323 &  n_1726;
assign n_2325 =  n_2059 &  n_2324;
assign n_2326 = ~n_980 &  n_1657;
assign n_2327 =  n_2326 &  n_2071;
assign n_2328 = ~n_1565 & ~n_2193;
assign n_2329 = ~n_845 &  n_2328;
assign n_2330 =  n_2327 &  n_2329;
assign n_2331 = ~n_967 & ~n_1411;
assign n_2332 = ~n_1148 &  n_2331;
assign n_2333 = ~n_1386 &  n_1959;
assign n_2334 =  n_2332 &  n_2333;
assign n_2335 =  n_2330 &  n_2334;
assign n_2336 =  n_280 &  n_1274;
assign n_2337 = ~x_42 &  n_1188;
assign n_2338 =  n_2176 & ~n_2337;
assign n_2339 = ~n_2336 &  n_2338;
assign n_2340 =  n_2162 &  n_1704;
assign n_2341 = ~n_987 & ~n_1384;
assign n_2342 =  n_2341 &  n_735;
assign n_2343 =  n_2340 &  n_2342;
assign n_2344 =  n_2339 &  n_2343;
assign n_2345 =  n_2335 &  n_2344;
assign n_2346 =  n_2325 &  n_2345;
assign n_2347 =  n_2317 &  n_2346;
assign n_2348 = ~n_1484 &  n_2347;
assign n_2349 = ~n_1749 &  n_2348;
assign n_2350 =  n_2286 &  n_2349;
assign n_2351 =  n_2244 &  n_1798;
assign n_2352 =  n_2350 &  n_2351;
assign n_2353 =  n_2283 &  n_2352;
assign n_2354 =  n_2034 &  n_2353;
assign n_2355 =  n_2281 &  n_2354;
assign n_2356 =  x_37 & ~n_2355;
assign n_2357 = ~x_37 &  n_2355;
assign n_2358 = ~n_2356 & ~n_2357;
assign n_2359 = ~n_1749 & ~n_808;
assign n_2360 =  n_1493 &  n_2359;
assign n_2361 = ~n_2149 &  n_1756;
assign n_2362 =  n_292 &  n_1472;
assign n_2363 = ~n_2362 &  n_1790;
assign n_2364 =  n_2361 &  n_2363;
assign n_2365 =  n_2360 &  n_2364;
assign n_2366 =  n_2253 &  n_2365;
assign n_2367 = ~n_559 &  n_2022;
assign n_2368 =  n_807 & ~n_278;
assign n_2369 = ~n_2368 & ~n_710;
assign n_2370 = ~n_912 & ~n_2219;
assign n_2371 =  n_1910 &  n_2370;
assign n_2372 = ~n_979 & ~n_803;
assign n_2373 = ~n_2175 &  n_2372;
assign n_2374 =  n_3 &  n_973;
assign n_2375 = ~n_1844 & ~n_2374;
assign n_2376 = ~n_1230 & ~n_1833;
assign n_2377 =  n_2375 &  n_2376;
assign n_2378 =  n_2373 &  n_2377;
assign n_2379 =  n_2164 &  n_2046;
assign n_2380 =  n_2378 &  n_2379;
assign n_2381 =  n_730 &  n_972;
assign n_2382 = ~n_734 & ~n_2381;
assign n_2383 = ~n_1828 & ~n_830;
assign n_2384 = ~n_2085 &  n_2383;
assign n_2385 =  n_2382 &  n_2384;
assign n_2386 = ~n_2227 &  n_1040;
assign n_2387 = ~n_853 & ~n_872;
assign n_2388 =  n_2387 & ~n_899;
assign n_2389 =  n_2386 &  n_2388;
assign n_2390 =  n_2385 &  n_2389;
assign n_2391 =  x_776 &  n_1369;
assign n_2392 =  n_2204 & ~n_2391;
assign n_2393 =  n_776 &  n_982;
assign n_2394 =  n_940 &  n_879;
assign n_2395 = ~n_1531 & ~n_2394;
assign n_2396 = ~n_2393 &  n_2395;
assign n_2397 =  n_2392 &  n_2396;
assign n_2398 =  n_2390 &  n_2397;
assign n_2399 =  n_2380 &  n_2398;
assign n_2400 =  n_2371 &  n_2399;
assign n_2401 =  n_1150 &  n_2039;
assign n_2402 =  n_1645 &  n_849;
assign n_2403 =  n_2401 &  n_2402;
assign n_2404 = ~n_1650 & ~n_1850;
assign n_2405 =  n_2124 & ~n_1390;
assign n_2406 =  n_2405 & ~n_1193;
assign n_2407 =  n_2404 &  n_2406;
assign n_2408 = ~n_1655 & ~n_893;
assign n_2409 =  n_903 &  n_281;
assign n_2410 = ~n_884 & ~n_2409;
assign n_2411 =  n_2408 &  n_2410;
assign n_2412 = ~n_1370 & ~n_854;
assign n_2413 =  n_2411 &  n_2412;
assign n_2414 =  n_705 &  n_990;
assign n_2415 = ~n_720 & ~n_928;
assign n_2416 = ~n_2414 &  n_2415;
assign n_2417 =  n_1375 &  n_2416;
assign n_2418 =  n_2413 &  n_2417;
assign n_2419 =  n_2407 &  n_2418;
assign n_2420 =  n_744 &  n_866;
assign n_2421 = ~n_2420 &  n_2207;
assign n_2422 =  n_2078 & ~n_871;
assign n_2423 =  n_2421 &  n_2422;
assign n_2424 =  n_2321 &  n_2208;
assign n_2425 =  x_1095 &  n_846;
assign n_2426 = ~n_2425 &  n_2341;
assign n_2427 =  n_2424 &  n_2426;
assign n_2428 =  n_2423 &  n_2427;
assign n_2429 =  n_2419 &  n_2428;
assign n_2430 =  n_2403 &  n_2429;
assign n_2431 =  n_1718 &  n_2430;
assign n_2432 =  n_2400 &  n_2431;
assign n_2433 = ~n_789 &  n_2432;
assign n_2434 =  n_2369 &  n_2433;
assign n_2435 = ~n_1458 &  n_1482;
assign n_2436 = ~n_1759 & ~n_2239;
assign n_2437 =  n_2435 &  n_2436;
assign n_2438 =  n_2434 &  n_2437;
assign n_2439 =  n_2367 &  n_2438;
assign n_2440 =  n_2366 &  n_2439;
assign n_2441 =  x_36 & ~n_2440;
assign n_2442 = ~x_36 &  n_2440;
assign n_2443 = ~n_2441 & ~n_2442;
assign n_2444 =  n_2277 & ~n_1785;
assign n_2445 = ~n_2031 &  n_2444;
assign n_2446 =  n_2445 &  n_2269;
assign n_2447 =  n_2030 &  n_1440;
assign n_2448 =  n_2446 &  n_2447;
assign n_2449 =  n_2248 & ~n_2409;
assign n_2450 =  n_1758 &  n_2251;
assign n_2451 = ~n_1383 &  n_2405;
assign n_2452 = ~n_1675 & ~n_2381;
assign n_2453 = ~n_845 &  n_2452;
assign n_2454 =  n_2451 &  n_2453;
assign n_2455 =  n_2454 &  n_1332;
assign n_2456 =  n_1191 &  n_2455;
assign n_2457 =  n_2041 &  n_2371;
assign n_2458 =  n_2456 &  n_2457;
assign n_2459 = ~n_1352 & ~n_1410;
assign n_2460 = ~n_965 &  n_2459;
assign n_2461 =  n_944 &  n_2460;
assign n_2462 =  n_2461 &  n_1997;
assign n_2463 =  n_1371 &  n_2462;
assign n_2464 =  n_2331 &  n_2218;
assign n_2465 =  n_1535 &  n_2464;
assign n_2466 =  n_2182 &  n_2465;
assign n_2467 =  n_2463 &  n_2466;
assign n_2468 = ~n_741 & ~n_936;
assign n_2469 = ~n_731 &  n_2468;
assign n_2470 = ~n_2391 & ~n_988;
assign n_2471 =  n_2469 &  n_2470;
assign n_2472 = ~n_697 & ~n_2125;
assign n_2473 = ~n_836 &  n_2472;
assign n_2474 =  n_707 &  n_2473;
assign n_2475 =  n_2471 &  n_2474;
assign n_2476 = ~n_1531 & ~n_993;
assign n_2477 = ~n_2306 &  n_2187;
assign n_2478 =  n_2476 &  n_2477;
assign n_2479 = ~n_1812 & ~n_1642;
assign n_2480 = ~n_1703 &  n_827;
assign n_2481 =  n_2479 &  n_2480;
assign n_2482 =  n_2478 &  n_2481;
assign n_2483 =  n_2475 &  n_2482;
assign n_2484 =  n_2375 & ~n_1193;
assign n_2485 =  n_1696 &  n_2484;
assign n_2486 =  n_2323 &  n_2485;
assign n_2487 =  n_2483 &  n_2486;
assign n_2488 =  n_2467 &  n_2487;
assign n_2489 =  n_2458 &  n_2488;
assign n_2490 = ~n_1484 &  n_2489;
assign n_2491 = ~n_1780 &  n_2490;
assign n_2492 =  n_1748 &  n_2491;
assign n_2493 =  n_2450 &  n_2492;
assign n_2494 = ~n_2284 & ~n_793;
assign n_2495 =  n_291 &  n_771;
assign n_2496 =  n_2494 & ~n_2495;
assign n_2497 =  n_2272 &  n_784;
assign n_2498 =  n_2496 &  n_2497;
assign n_2499 = ~n_1489 & ~n_552;
assign n_2500 = ~n_1458 &  n_2010;
assign n_2501 =  n_2499 &  n_2500;
assign n_2502 =  n_2498 &  n_2501;
assign n_2503 =  n_2493 &  n_2502;
assign n_2504 =  n_2449 &  n_2503;
assign n_2505 =  n_2448 &  n_2504;
assign n_2506 =  x_35 & ~n_2505;
assign n_2507 = ~x_35 &  n_2505;
assign n_2508 = ~n_2506 & ~n_2507;
assign n_2509 =  n_2445 &  n_1486;
assign n_2510 =  n_1483 &  n_2509;
assign n_2511 =  n_1341 &  n_2451;
assign n_2512 =  n_2453 &  n_1533;
assign n_2513 =  n_2511 &  n_2512;
assign n_2514 =  n_1813 &  n_2107;
assign n_2515 =  n_2378 &  n_2514;
assign n_2516 =  n_2513 &  n_2515;
assign n_2517 =  n_2161 &  n_2516;
assign n_2518 =  n_2328 &  n_1693;
assign n_2519 = ~n_1710 &  n_2518;
assign n_2520 =  n_1589 &  n_2519;
assign n_2521 =  n_1867 &  n_1637;
assign n_2522 =  n_2520 &  n_2521;
assign n_2523 = ~n_1671 & ~n_1728;
assign n_2524 = ~n_925 &  n_2523;
assign n_2525 = ~n_909 &  n_2524;
assign n_2526 =  n_1979 &  n_985;
assign n_2527 =  n_2525 &  n_2526;
assign n_2528 = ~n_801 & ~n_962;
assign n_2529 = ~n_1357 & ~n_1841;
assign n_2530 =  n_2528 &  n_2529;
assign n_2531 = ~n_797 & ~n_914;
assign n_2532 = ~n_743 & ~n_1553;
assign n_2533 =  n_2531 &  n_2532;
assign n_2534 = ~n_1705 & ~n_876;
assign n_2535 =  n_2533 &  n_2534;
assign n_2536 =  n_2530 &  n_2535;
assign n_2537 =  n_2527 &  n_2536;
assign n_2538 =  n_2086 &  n_1974;
assign n_2539 =  n_2090 &  n_994;
assign n_2540 =  n_2538 &  n_2539;
assign n_2541 =  n_2087 &  n_2205;
assign n_2542 =  n_2327 &  n_2541;
assign n_2543 =  n_2540 &  n_2542;
assign n_2544 =  n_2537 &  n_2543;
assign n_2545 =  n_2292 &  n_1529;
assign n_2546 =  n_1378 &  n_1804;
assign n_2547 =  n_2545 &  n_2546;
assign n_2548 = ~n_1711 & ~n_1642;
assign n_2549 = ~n_1722 & ~n_1384;
assign n_2550 =  n_2548 &  n_2549;
assign n_2551 = ~n_1817 & ~n_841;
assign n_2552 =  n_2127 &  n_712;
assign n_2553 =  n_2551 &  n_2552;
assign n_2554 =  n_2550 &  n_2553;
assign n_2555 =  n_827 & ~n_2049;
assign n_2556 = ~n_2304 &  n_2383;
assign n_2557 =  n_2555 &  n_2556;
assign n_2558 =  n_907 &  n_2557;
assign n_2559 =  n_2554 &  n_2558;
assign n_2560 =  n_2547 &  n_2559;
assign n_2561 =  n_2544 &  n_2560;
assign n_2562 =  n_2522 &  n_2561;
assign n_2563 =  n_2517 &  n_2562;
assign n_2564 = ~n_1494 &  n_2563;
assign n_2565 = ~n_1471 &  n_2564;
assign n_2566 =  n_1798 &  n_2565;
assign n_2567 =  n_2450 &  n_2566;
assign n_2568 = ~n_778 & ~n_1786;
assign n_2569 = ~n_1788 & ~n_2239;
assign n_2570 =  n_2568 &  n_2569;
assign n_2571 = ~n_1473 & ~n_1435;
assign n_2572 = ~n_419 &  n_2494;
assign n_2573 =  n_2571 &  n_2572;
assign n_2574 =  n_2570 &  n_2573;
assign n_2575 =  n_2567 &  n_2574;
assign n_2576 =  n_2367 &  n_2575;
assign n_2577 =  n_2510 &  n_2576;
assign n_2578 =  x_34 & ~n_2577;
assign n_2579 = ~x_34 &  n_2577;
assign n_2580 = ~n_2578 & ~n_2579;
assign n_2581 = ~n_550 &  n_801;
assign n_2582 =  n_2392 &  n_2097;
assign n_2583 =  n_1993 &  n_2582;
assign n_2584 = ~n_717 & ~n_743;
assign n_2585 = ~n_1437 & ~n_924;
assign n_2586 =  n_2584 &  n_2585;
assign n_2587 = ~n_1661 & ~n_741;
assign n_2588 = ~n_797 & ~n_1572;
assign n_2589 =  n_2587 &  n_2588;
assign n_2590 =  n_2586 &  n_2589;
assign n_2591 =  n_1375 & ~n_1321;
assign n_2592 =  n_2590 &  n_2591;
assign n_2593 = ~n_870 & ~n_861;
assign n_2594 =  n_2387 & ~n_852;
assign n_2595 =  n_2593 &  n_2594;
assign n_2596 = ~n_931 & ~n_747;
assign n_2597 = ~n_731 & ~n_751;
assign n_2598 =  n_2596 &  n_2597;
assign n_2599 =  n_2595 &  n_2598;
assign n_2600 =  n_2592 &  n_2599;
assign n_2601 =  n_2583 &  n_2600;
assign n_2602 =  n_1151 &  n_1987;
assign n_2603 =  n_2601 &  n_2602;
assign n_2604 =  n_1190 &  n_2230;
assign n_2605 =  n_908 &  n_2604;
assign n_2606 =  n_981 &  n_2068;
assign n_2607 =  n_1652 &  n_2318;
assign n_2608 =  n_2606 &  n_2607;
assign n_2609 =  n_707 &  n_999;
assign n_2610 =  n_1959 &  n_1041;
assign n_2611 =  n_2609 &  n_2610;
assign n_2612 =  n_2608 &  n_2611;
assign n_2613 =  n_919 &  n_2184;
assign n_2614 =  n_2612 &  n_2613;
assign n_2615 =  n_2605 &  n_2614;
assign n_2616 =  n_2467 &  n_2615;
assign n_2617 =  n_2603 &  n_2616;
assign n_2618 = ~n_2581 &  n_2617;
assign n_2619 = ~n_552 &  n_2618;
assign n_2620 =  n_2369 &  n_805;
assign n_2621 =  n_2619 &  n_2620;
assign n_2622 =  n_2360 &  n_2621;
assign n_2623 =  n_2622 &  n_1476;
assign n_2624 = ~n_550 &  n_697;
assign n_2625 = ~n_288 & ~n_2624;
assign n_2626 = ~n_278 &  n_803;
assign n_2627 = ~n_1494 & ~n_2626;
assign n_2628 =  n_2625 &  n_2627;
assign n_2629 =  n_2268 &  n_2628;
assign n_2630 =  n_2011 &  n_699;
assign n_2631 =  n_2629 &  n_2630;
assign n_2632 =  n_2449 &  n_2631;
assign n_2633 =  n_2259 &  n_2632;
assign n_2634 =  n_2623 &  n_2633;
assign n_2635 =  x_33 & ~n_2634;
assign n_2636 = ~x_33 &  n_2634;
assign n_2637 = ~n_2635 & ~n_2636;
assign n_2638 =  x_1126 & ~n_1590;
assign n_2639 =  x_297 &  n_1590;
assign n_2640 = ~n_2638 & ~n_2639;
assign n_2641 =  x_1126 & ~n_2640;
assign n_2642 = ~x_1126 &  n_2640;
assign n_2643 = ~n_2641 & ~n_2642;
assign n_2644 =  x_1125 & ~n_1590;
assign n_2645 =  x_296 &  n_1590;
assign n_2646 = ~n_2644 & ~n_2645;
assign n_2647 =  x_1125 & ~n_2646;
assign n_2648 = ~x_1125 &  n_2646;
assign n_2649 = ~n_2647 & ~n_2648;
assign n_2650 =  x_1124 & ~n_1590;
assign n_2651 =  x_295 &  n_1590;
assign n_2652 = ~n_2650 & ~n_2651;
assign n_2653 =  x_1124 & ~n_2652;
assign n_2654 = ~x_1124 &  n_2652;
assign n_2655 = ~n_2653 & ~n_2654;
assign n_2656 =  x_1123 & ~n_1590;
assign n_2657 =  x_294 &  n_1590;
assign n_2658 = ~n_2656 & ~n_2657;
assign n_2659 =  x_1123 & ~n_2658;
assign n_2660 = ~x_1123 &  n_2658;
assign n_2661 = ~n_2659 & ~n_2660;
assign n_2662 =  x_1122 & ~n_1590;
assign n_2663 =  x_293 &  n_1590;
assign n_2664 = ~n_2662 & ~n_2663;
assign n_2665 =  x_1122 & ~n_2664;
assign n_2666 = ~x_1122 &  n_2664;
assign n_2667 = ~n_2665 & ~n_2666;
assign n_2668 =  x_1121 & ~n_1590;
assign n_2669 =  x_292 &  n_1590;
assign n_2670 = ~n_2668 & ~n_2669;
assign n_2671 =  x_1121 & ~n_2670;
assign n_2672 = ~x_1121 &  n_2670;
assign n_2673 = ~n_2671 & ~n_2672;
assign n_2674 =  x_1120 & ~n_1590;
assign n_2675 =  x_291 &  n_1590;
assign n_2676 = ~n_2674 & ~n_2675;
assign n_2677 =  x_1120 & ~n_2676;
assign n_2678 = ~x_1120 &  n_2676;
assign n_2679 = ~n_2677 & ~n_2678;
assign n_2680 =  x_1119 & ~n_1590;
assign n_2681 =  x_290 &  n_1590;
assign n_2682 = ~n_2680 & ~n_2681;
assign n_2683 =  x_1119 & ~n_2682;
assign n_2684 = ~x_1119 &  n_2682;
assign n_2685 = ~n_2683 & ~n_2684;
assign n_2686 =  x_1118 & ~n_1590;
assign n_2687 =  x_289 &  n_1590;
assign n_2688 = ~n_2686 & ~n_2687;
assign n_2689 =  x_1118 & ~n_2688;
assign n_2690 = ~x_1118 &  n_2688;
assign n_2691 = ~n_2689 & ~n_2690;
assign n_2692 =  x_1117 & ~n_1590;
assign n_2693 =  x_288 &  n_1590;
assign n_2694 = ~n_2692 & ~n_2693;
assign n_2695 =  x_1117 & ~n_2694;
assign n_2696 = ~x_1117 &  n_2694;
assign n_2697 = ~n_2695 & ~n_2696;
assign n_2698 =  x_1116 & ~n_1590;
assign n_2699 =  x_287 &  n_1590;
assign n_2700 = ~n_2698 & ~n_2699;
assign n_2701 =  x_1116 & ~n_2700;
assign n_2702 = ~x_1116 &  n_2700;
assign n_2703 = ~n_2701 & ~n_2702;
assign n_2704 =  x_1115 & ~n_1590;
assign n_2705 =  x_286 &  n_1590;
assign n_2706 = ~n_2704 & ~n_2705;
assign n_2707 =  x_1115 & ~n_2706;
assign n_2708 = ~x_1115 &  n_2706;
assign n_2709 = ~n_2707 & ~n_2708;
assign n_2710 =  x_1114 & ~n_1590;
assign n_2711 =  x_285 &  n_1590;
assign n_2712 = ~n_2710 & ~n_2711;
assign n_2713 =  x_1114 & ~n_2712;
assign n_2714 = ~x_1114 &  n_2712;
assign n_2715 = ~n_2713 & ~n_2714;
assign n_2716 =  x_1113 & ~n_1590;
assign n_2717 =  x_284 &  n_1590;
assign n_2718 = ~n_2716 & ~n_2717;
assign n_2719 =  x_1113 & ~n_2718;
assign n_2720 = ~x_1113 &  n_2718;
assign n_2721 = ~n_2719 & ~n_2720;
assign n_2722 =  x_1112 & ~n_1590;
assign n_2723 =  x_283 &  n_1590;
assign n_2724 = ~n_2722 & ~n_2723;
assign n_2725 =  x_1112 & ~n_2724;
assign n_2726 = ~x_1112 &  n_2724;
assign n_2727 = ~n_2725 & ~n_2726;
assign n_2728 =  x_1111 & ~n_1590;
assign n_2729 =  x_282 &  n_1590;
assign n_2730 = ~n_2728 & ~n_2729;
assign n_2731 =  x_1111 & ~n_2730;
assign n_2732 = ~x_1111 &  n_2730;
assign n_2733 = ~n_2731 & ~n_2732;
assign n_2734 =  x_1110 & ~n_1590;
assign n_2735 =  x_281 &  n_1590;
assign n_2736 = ~n_2734 & ~n_2735;
assign n_2737 =  x_1110 & ~n_2736;
assign n_2738 = ~x_1110 &  n_2736;
assign n_2739 = ~n_2737 & ~n_2738;
assign n_2740 =  x_1109 & ~n_1590;
assign n_2741 =  x_280 &  n_1590;
assign n_2742 = ~n_2740 & ~n_2741;
assign n_2743 =  x_1109 & ~n_2742;
assign n_2744 = ~x_1109 &  n_2742;
assign n_2745 = ~n_2743 & ~n_2744;
assign n_2746 =  x_1108 & ~n_1590;
assign n_2747 =  x_279 &  n_1590;
assign n_2748 = ~n_2746 & ~n_2747;
assign n_2749 =  x_1108 & ~n_2748;
assign n_2750 = ~x_1108 &  n_2748;
assign n_2751 = ~n_2749 & ~n_2750;
assign n_2752 =  x_1107 & ~n_1590;
assign n_2753 =  x_278 &  n_1590;
assign n_2754 = ~n_2752 & ~n_2753;
assign n_2755 =  x_1107 & ~n_2754;
assign n_2756 = ~x_1107 &  n_2754;
assign n_2757 = ~n_2755 & ~n_2756;
assign n_2758 =  x_1106 & ~n_1590;
assign n_2759 =  x_277 &  n_1590;
assign n_2760 = ~n_2758 & ~n_2759;
assign n_2761 =  x_1106 & ~n_2760;
assign n_2762 = ~x_1106 &  n_2760;
assign n_2763 = ~n_2761 & ~n_2762;
assign n_2764 =  x_1105 & ~n_1590;
assign n_2765 =  x_276 &  n_1590;
assign n_2766 = ~n_2764 & ~n_2765;
assign n_2767 =  x_1105 & ~n_2766;
assign n_2768 = ~x_1105 &  n_2766;
assign n_2769 = ~n_2767 & ~n_2768;
assign n_2770 =  x_1104 & ~n_1590;
assign n_2771 =  x_275 &  n_1590;
assign n_2772 = ~n_2770 & ~n_2771;
assign n_2773 =  x_1104 & ~n_2772;
assign n_2774 = ~x_1104 &  n_2772;
assign n_2775 = ~n_2773 & ~n_2774;
assign n_2776 =  x_1103 & ~n_1590;
assign n_2777 =  x_274 &  n_1590;
assign n_2778 = ~n_2776 & ~n_2777;
assign n_2779 =  x_1103 & ~n_2778;
assign n_2780 = ~x_1103 &  n_2778;
assign n_2781 = ~n_2779 & ~n_2780;
assign n_2782 =  x_1102 & ~n_1590;
assign n_2783 =  x_273 &  n_1590;
assign n_2784 = ~n_2782 & ~n_2783;
assign n_2785 =  x_1102 & ~n_2784;
assign n_2786 = ~x_1102 &  n_2784;
assign n_2787 = ~n_2785 & ~n_2786;
assign n_2788 =  x_1101 & ~n_1590;
assign n_2789 =  x_272 &  n_1590;
assign n_2790 = ~n_2788 & ~n_2789;
assign n_2791 =  x_1101 & ~n_2790;
assign n_2792 = ~x_1101 &  n_2790;
assign n_2793 = ~n_2791 & ~n_2792;
assign n_2794 =  x_1100 & ~n_1590;
assign n_2795 =  x_271 &  n_1590;
assign n_2796 = ~n_2794 & ~n_2795;
assign n_2797 =  x_1100 & ~n_2796;
assign n_2798 = ~x_1100 &  n_2796;
assign n_2799 = ~n_2797 & ~n_2798;
assign n_2800 =  x_1099 & ~n_1590;
assign n_2801 =  x_270 &  n_1590;
assign n_2802 = ~n_2800 & ~n_2801;
assign n_2803 =  x_1099 & ~n_2802;
assign n_2804 = ~x_1099 &  n_2802;
assign n_2805 = ~n_2803 & ~n_2804;
assign n_2806 =  x_1098 & ~n_1590;
assign n_2807 =  x_269 &  n_1590;
assign n_2808 = ~n_2806 & ~n_2807;
assign n_2809 =  x_1098 & ~n_2808;
assign n_2810 = ~x_1098 &  n_2808;
assign n_2811 = ~n_2809 & ~n_2810;
assign n_2812 =  x_1097 & ~n_1590;
assign n_2813 =  x_268 &  n_1590;
assign n_2814 = ~n_2812 & ~n_2813;
assign n_2815 =  x_1097 & ~n_2814;
assign n_2816 = ~x_1097 &  n_2814;
assign n_2817 = ~n_2815 & ~n_2816;
assign n_2818 =  x_1096 & ~n_1590;
assign n_2819 =  x_267 &  n_1590;
assign n_2820 = ~n_2818 & ~n_2819;
assign n_2821 =  x_1096 & ~n_2820;
assign n_2822 = ~x_1096 &  n_2820;
assign n_2823 = ~n_2821 & ~n_2822;
assign n_2824 =  x_1095 & ~n_1590;
assign n_2825 =  x_1095 &  n_2824;
assign n_2826 = ~x_1095 & ~n_2824;
assign n_2827 = ~n_2825 & ~n_2826;
assign n_2828 =  i_32 &  n_1270;
assign n_2829 =  x_1094 & ~n_1270;
assign n_2830 = ~n_2828 & ~n_2829;
assign n_2831 =  x_1094 & ~n_2830;
assign n_2832 = ~x_1094 &  n_2830;
assign n_2833 = ~n_2831 & ~n_2832;
assign n_2834 =  i_31 &  n_1270;
assign n_2835 =  x_1093 & ~n_1270;
assign n_2836 = ~n_2834 & ~n_2835;
assign n_2837 =  x_1093 & ~n_2836;
assign n_2838 = ~x_1093 &  n_2836;
assign n_2839 = ~n_2837 & ~n_2838;
assign n_2840 =  i_30 &  n_1270;
assign n_2841 =  x_1092 & ~n_1270;
assign n_2842 = ~n_2840 & ~n_2841;
assign n_2843 =  x_1092 & ~n_2842;
assign n_2844 = ~x_1092 &  n_2842;
assign n_2845 = ~n_2843 & ~n_2844;
assign n_2846 =  i_29 &  n_1270;
assign n_2847 =  x_1091 & ~n_1270;
assign n_2848 = ~n_2846 & ~n_2847;
assign n_2849 =  x_1091 & ~n_2848;
assign n_2850 = ~x_1091 &  n_2848;
assign n_2851 = ~n_2849 & ~n_2850;
assign n_2852 =  i_28 &  n_1270;
assign n_2853 =  x_1090 & ~n_1270;
assign n_2854 = ~n_2852 & ~n_2853;
assign n_2855 =  x_1090 & ~n_2854;
assign n_2856 = ~x_1090 &  n_2854;
assign n_2857 = ~n_2855 & ~n_2856;
assign n_2858 =  i_27 &  n_1270;
assign n_2859 =  x_1089 & ~n_1270;
assign n_2860 = ~n_2858 & ~n_2859;
assign n_2861 =  x_1089 & ~n_2860;
assign n_2862 = ~x_1089 &  n_2860;
assign n_2863 = ~n_2861 & ~n_2862;
assign n_2864 =  i_26 &  n_1270;
assign n_2865 =  x_1088 & ~n_1270;
assign n_2866 = ~n_2864 & ~n_2865;
assign n_2867 =  x_1088 & ~n_2866;
assign n_2868 = ~x_1088 &  n_2866;
assign n_2869 = ~n_2867 & ~n_2868;
assign n_2870 =  i_25 &  n_1270;
assign n_2871 =  x_1087 & ~n_1270;
assign n_2872 = ~n_2870 & ~n_2871;
assign n_2873 =  x_1087 & ~n_2872;
assign n_2874 = ~x_1087 &  n_2872;
assign n_2875 = ~n_2873 & ~n_2874;
assign n_2876 =  i_24 &  n_1270;
assign n_2877 =  x_1086 & ~n_1270;
assign n_2878 = ~n_2876 & ~n_2877;
assign n_2879 =  x_1086 & ~n_2878;
assign n_2880 = ~x_1086 &  n_2878;
assign n_2881 = ~n_2879 & ~n_2880;
assign n_2882 =  i_23 &  n_1270;
assign n_2883 =  x_1085 & ~n_1270;
assign n_2884 = ~n_2882 & ~n_2883;
assign n_2885 =  x_1085 & ~n_2884;
assign n_2886 = ~x_1085 &  n_2884;
assign n_2887 = ~n_2885 & ~n_2886;
assign n_2888 =  i_22 &  n_1270;
assign n_2889 =  x_1084 & ~n_1270;
assign n_2890 = ~n_2888 & ~n_2889;
assign n_2891 =  x_1084 & ~n_2890;
assign n_2892 = ~x_1084 &  n_2890;
assign n_2893 = ~n_2891 & ~n_2892;
assign n_2894 =  i_21 &  n_1270;
assign n_2895 =  x_1083 & ~n_1270;
assign n_2896 = ~n_2894 & ~n_2895;
assign n_2897 =  x_1083 & ~n_2896;
assign n_2898 = ~x_1083 &  n_2896;
assign n_2899 = ~n_2897 & ~n_2898;
assign n_2900 =  i_20 &  n_1270;
assign n_2901 =  x_1082 & ~n_1270;
assign n_2902 = ~n_2900 & ~n_2901;
assign n_2903 =  x_1082 & ~n_2902;
assign n_2904 = ~x_1082 &  n_2902;
assign n_2905 = ~n_2903 & ~n_2904;
assign n_2906 =  i_19 &  n_1270;
assign n_2907 =  x_1081 & ~n_1270;
assign n_2908 = ~n_2906 & ~n_2907;
assign n_2909 =  x_1081 & ~n_2908;
assign n_2910 = ~x_1081 &  n_2908;
assign n_2911 = ~n_2909 & ~n_2910;
assign n_2912 =  i_18 &  n_1270;
assign n_2913 =  x_1080 & ~n_1270;
assign n_2914 = ~n_2912 & ~n_2913;
assign n_2915 =  x_1080 & ~n_2914;
assign n_2916 = ~x_1080 &  n_2914;
assign n_2917 = ~n_2915 & ~n_2916;
assign n_2918 =  i_17 &  n_1270;
assign n_2919 =  x_1079 & ~n_1270;
assign n_2920 = ~n_2918 & ~n_2919;
assign n_2921 =  x_1079 & ~n_2920;
assign n_2922 = ~x_1079 &  n_2920;
assign n_2923 = ~n_2921 & ~n_2922;
assign n_2924 =  i_16 &  n_1270;
assign n_2925 =  x_1078 & ~n_1270;
assign n_2926 = ~n_2924 & ~n_2925;
assign n_2927 =  x_1078 & ~n_2926;
assign n_2928 = ~x_1078 &  n_2926;
assign n_2929 = ~n_2927 & ~n_2928;
assign n_2930 =  i_15 &  n_1270;
assign n_2931 =  x_1077 & ~n_1270;
assign n_2932 = ~n_2930 & ~n_2931;
assign n_2933 =  x_1077 & ~n_2932;
assign n_2934 = ~x_1077 &  n_2932;
assign n_2935 = ~n_2933 & ~n_2934;
assign n_2936 =  i_14 &  n_1270;
assign n_2937 =  x_1076 & ~n_1270;
assign n_2938 = ~n_2936 & ~n_2937;
assign n_2939 =  x_1076 & ~n_2938;
assign n_2940 = ~x_1076 &  n_2938;
assign n_2941 = ~n_2939 & ~n_2940;
assign n_2942 =  i_13 &  n_1270;
assign n_2943 =  x_1075 & ~n_1270;
assign n_2944 = ~n_2942 & ~n_2943;
assign n_2945 =  x_1075 & ~n_2944;
assign n_2946 = ~x_1075 &  n_2944;
assign n_2947 = ~n_2945 & ~n_2946;
assign n_2948 =  i_12 &  n_1270;
assign n_2949 =  x_1074 & ~n_1270;
assign n_2950 = ~n_2948 & ~n_2949;
assign n_2951 =  x_1074 & ~n_2950;
assign n_2952 = ~x_1074 &  n_2950;
assign n_2953 = ~n_2951 & ~n_2952;
assign n_2954 =  i_11 &  n_1270;
assign n_2955 =  x_1073 & ~n_1270;
assign n_2956 = ~n_2954 & ~n_2955;
assign n_2957 =  x_1073 & ~n_2956;
assign n_2958 = ~x_1073 &  n_2956;
assign n_2959 = ~n_2957 & ~n_2958;
assign n_2960 =  i_10 &  n_1270;
assign n_2961 =  x_1072 & ~n_1270;
assign n_2962 = ~n_2960 & ~n_2961;
assign n_2963 =  x_1072 & ~n_2962;
assign n_2964 = ~x_1072 &  n_2962;
assign n_2965 = ~n_2963 & ~n_2964;
assign n_2966 =  i_9 &  n_1270;
assign n_2967 =  x_1071 & ~n_1270;
assign n_2968 = ~n_2966 & ~n_2967;
assign n_2969 =  x_1071 & ~n_2968;
assign n_2970 = ~x_1071 &  n_2968;
assign n_2971 = ~n_2969 & ~n_2970;
assign n_2972 =  i_8 &  n_1270;
assign n_2973 =  x_1070 & ~n_1270;
assign n_2974 = ~n_2972 & ~n_2973;
assign n_2975 =  x_1070 & ~n_2974;
assign n_2976 = ~x_1070 &  n_2974;
assign n_2977 = ~n_2975 & ~n_2976;
assign n_2978 =  i_7 &  n_1270;
assign n_2979 =  x_1069 & ~n_1270;
assign n_2980 = ~n_2978 & ~n_2979;
assign n_2981 =  x_1069 & ~n_2980;
assign n_2982 = ~x_1069 &  n_2980;
assign n_2983 = ~n_2981 & ~n_2982;
assign n_2984 =  i_6 &  n_1270;
assign n_2985 =  x_1068 & ~n_1270;
assign n_2986 = ~n_2984 & ~n_2985;
assign n_2987 =  x_1068 & ~n_2986;
assign n_2988 = ~x_1068 &  n_2986;
assign n_2989 = ~n_2987 & ~n_2988;
assign n_2990 =  i_5 &  n_1270;
assign n_2991 =  x_1067 & ~n_1270;
assign n_2992 = ~n_2990 & ~n_2991;
assign n_2993 =  x_1067 & ~n_2992;
assign n_2994 = ~x_1067 &  n_2992;
assign n_2995 = ~n_2993 & ~n_2994;
assign n_2996 =  i_4 &  n_1270;
assign n_2997 =  x_1066 & ~n_1270;
assign n_2998 = ~n_2996 & ~n_2997;
assign n_2999 =  x_1066 & ~n_2998;
assign n_3000 = ~x_1066 &  n_2998;
assign n_3001 = ~n_2999 & ~n_3000;
assign n_3002 =  i_3 &  n_1270;
assign n_3003 =  x_1065 & ~n_1270;
assign n_3004 = ~n_3002 & ~n_3003;
assign n_3005 =  x_1065 & ~n_3004;
assign n_3006 = ~x_1065 &  n_3004;
assign n_3007 = ~n_3005 & ~n_3006;
assign n_3008 =  i_2 &  n_1270;
assign n_3009 =  x_1064 & ~n_1270;
assign n_3010 = ~n_3008 & ~n_3009;
assign n_3011 =  x_1064 & ~n_3010;
assign n_3012 = ~x_1064 &  n_3010;
assign n_3013 = ~n_3011 & ~n_3012;
assign n_3014 =  i_1 &  n_1270;
assign n_3015 =  x_1063 & ~n_1270;
assign n_3016 = ~n_3014 & ~n_3015;
assign n_3017 =  x_1063 & ~n_3016;
assign n_3018 = ~x_1063 &  n_3016;
assign n_3019 = ~n_3017 & ~n_3018;
assign n_3020 =  x_1062 & ~n_9;
assign n_3021 =  x_361 &  n_9;
assign n_3022 = ~n_3020 & ~n_3021;
assign n_3023 =  x_1062 & ~n_3022;
assign n_3024 = ~x_1062 &  n_3022;
assign n_3025 = ~n_3023 & ~n_3024;
assign n_3026 =  x_1061 & ~n_9;
assign n_3027 =  x_360 &  n_9;
assign n_3028 = ~n_3026 & ~n_3027;
assign n_3029 =  x_1061 & ~n_3028;
assign n_3030 = ~x_1061 &  n_3028;
assign n_3031 = ~n_3029 & ~n_3030;
assign n_3032 =  x_1060 & ~n_9;
assign n_3033 =  x_359 &  n_9;
assign n_3034 = ~n_3032 & ~n_3033;
assign n_3035 =  x_1060 & ~n_3034;
assign n_3036 = ~x_1060 &  n_3034;
assign n_3037 = ~n_3035 & ~n_3036;
assign n_3038 =  x_1059 & ~n_9;
assign n_3039 =  x_358 &  n_9;
assign n_3040 = ~n_3038 & ~n_3039;
assign n_3041 =  x_1059 & ~n_3040;
assign n_3042 = ~x_1059 &  n_3040;
assign n_3043 = ~n_3041 & ~n_3042;
assign n_3044 =  x_1058 & ~n_9;
assign n_3045 =  x_357 &  n_9;
assign n_3046 = ~n_3044 & ~n_3045;
assign n_3047 =  x_1058 & ~n_3046;
assign n_3048 = ~x_1058 &  n_3046;
assign n_3049 = ~n_3047 & ~n_3048;
assign n_3050 =  x_1057 & ~n_9;
assign n_3051 =  x_356 &  n_9;
assign n_3052 = ~n_3050 & ~n_3051;
assign n_3053 =  x_1057 & ~n_3052;
assign n_3054 = ~x_1057 &  n_3052;
assign n_3055 = ~n_3053 & ~n_3054;
assign n_3056 =  x_1056 & ~n_9;
assign n_3057 =  x_355 &  n_9;
assign n_3058 = ~n_3056 & ~n_3057;
assign n_3059 =  x_1056 & ~n_3058;
assign n_3060 = ~x_1056 &  n_3058;
assign n_3061 = ~n_3059 & ~n_3060;
assign n_3062 =  x_1055 & ~n_9;
assign n_3063 =  x_354 &  n_9;
assign n_3064 = ~n_3062 & ~n_3063;
assign n_3065 =  x_1055 & ~n_3064;
assign n_3066 = ~x_1055 &  n_3064;
assign n_3067 = ~n_3065 & ~n_3066;
assign n_3068 =  x_1054 & ~n_9;
assign n_3069 =  x_353 &  n_9;
assign n_3070 = ~n_3068 & ~n_3069;
assign n_3071 =  x_1054 & ~n_3070;
assign n_3072 = ~x_1054 &  n_3070;
assign n_3073 = ~n_3071 & ~n_3072;
assign n_3074 =  x_1053 & ~n_9;
assign n_3075 =  x_352 &  n_9;
assign n_3076 = ~n_3074 & ~n_3075;
assign n_3077 =  x_1053 & ~n_3076;
assign n_3078 = ~x_1053 &  n_3076;
assign n_3079 = ~n_3077 & ~n_3078;
assign n_3080 =  x_1052 & ~n_9;
assign n_3081 =  x_351 &  n_9;
assign n_3082 = ~n_3080 & ~n_3081;
assign n_3083 =  x_1052 & ~n_3082;
assign n_3084 = ~x_1052 &  n_3082;
assign n_3085 = ~n_3083 & ~n_3084;
assign n_3086 =  x_1051 & ~n_9;
assign n_3087 =  x_350 &  n_9;
assign n_3088 = ~n_3086 & ~n_3087;
assign n_3089 =  x_1051 & ~n_3088;
assign n_3090 = ~x_1051 &  n_3088;
assign n_3091 = ~n_3089 & ~n_3090;
assign n_3092 =  x_1050 & ~n_9;
assign n_3093 =  x_349 &  n_9;
assign n_3094 = ~n_3092 & ~n_3093;
assign n_3095 =  x_1050 & ~n_3094;
assign n_3096 = ~x_1050 &  n_3094;
assign n_3097 = ~n_3095 & ~n_3096;
assign n_3098 =  x_1049 & ~n_9;
assign n_3099 =  x_348 &  n_9;
assign n_3100 = ~n_3098 & ~n_3099;
assign n_3101 =  x_1049 & ~n_3100;
assign n_3102 = ~x_1049 &  n_3100;
assign n_3103 = ~n_3101 & ~n_3102;
assign n_3104 =  x_1048 & ~n_9;
assign n_3105 =  x_347 &  n_9;
assign n_3106 = ~n_3104 & ~n_3105;
assign n_3107 =  x_1048 & ~n_3106;
assign n_3108 = ~x_1048 &  n_3106;
assign n_3109 = ~n_3107 & ~n_3108;
assign n_3110 =  x_1047 & ~n_9;
assign n_3111 =  x_346 &  n_9;
assign n_3112 = ~n_3110 & ~n_3111;
assign n_3113 =  x_1047 & ~n_3112;
assign n_3114 = ~x_1047 &  n_3112;
assign n_3115 = ~n_3113 & ~n_3114;
assign n_3116 =  x_1046 & ~n_9;
assign n_3117 =  x_345 &  n_9;
assign n_3118 = ~n_3116 & ~n_3117;
assign n_3119 =  x_1046 & ~n_3118;
assign n_3120 = ~x_1046 &  n_3118;
assign n_3121 = ~n_3119 & ~n_3120;
assign n_3122 =  x_1045 & ~n_9;
assign n_3123 =  x_344 &  n_9;
assign n_3124 = ~n_3122 & ~n_3123;
assign n_3125 =  x_1045 & ~n_3124;
assign n_3126 = ~x_1045 &  n_3124;
assign n_3127 = ~n_3125 & ~n_3126;
assign n_3128 =  x_1044 & ~n_9;
assign n_3129 =  x_343 &  n_9;
assign n_3130 = ~n_3128 & ~n_3129;
assign n_3131 =  x_1044 & ~n_3130;
assign n_3132 = ~x_1044 &  n_3130;
assign n_3133 = ~n_3131 & ~n_3132;
assign n_3134 =  x_1043 & ~n_9;
assign n_3135 =  x_342 &  n_9;
assign n_3136 = ~n_3134 & ~n_3135;
assign n_3137 =  x_1043 & ~n_3136;
assign n_3138 = ~x_1043 &  n_3136;
assign n_3139 = ~n_3137 & ~n_3138;
assign n_3140 =  x_1042 & ~n_9;
assign n_3141 =  x_341 &  n_9;
assign n_3142 = ~n_3140 & ~n_3141;
assign n_3143 =  x_1042 & ~n_3142;
assign n_3144 = ~x_1042 &  n_3142;
assign n_3145 = ~n_3143 & ~n_3144;
assign n_3146 =  x_1041 & ~n_9;
assign n_3147 =  x_340 &  n_9;
assign n_3148 = ~n_3146 & ~n_3147;
assign n_3149 =  x_1041 & ~n_3148;
assign n_3150 = ~x_1041 &  n_3148;
assign n_3151 = ~n_3149 & ~n_3150;
assign n_3152 =  x_1040 & ~n_9;
assign n_3153 =  x_339 &  n_9;
assign n_3154 = ~n_3152 & ~n_3153;
assign n_3155 =  x_1040 & ~n_3154;
assign n_3156 = ~x_1040 &  n_3154;
assign n_3157 = ~n_3155 & ~n_3156;
assign n_3158 =  x_1039 & ~n_9;
assign n_3159 =  x_338 &  n_9;
assign n_3160 = ~n_3158 & ~n_3159;
assign n_3161 =  x_1039 & ~n_3160;
assign n_3162 = ~x_1039 &  n_3160;
assign n_3163 = ~n_3161 & ~n_3162;
assign n_3164 =  x_1038 & ~n_9;
assign n_3165 =  x_337 &  n_9;
assign n_3166 = ~n_3164 & ~n_3165;
assign n_3167 =  x_1038 & ~n_3166;
assign n_3168 = ~x_1038 &  n_3166;
assign n_3169 = ~n_3167 & ~n_3168;
assign n_3170 =  x_1037 & ~n_9;
assign n_3171 =  x_336 &  n_9;
assign n_3172 = ~n_3170 & ~n_3171;
assign n_3173 =  x_1037 & ~n_3172;
assign n_3174 = ~x_1037 &  n_3172;
assign n_3175 = ~n_3173 & ~n_3174;
assign n_3176 =  x_1036 & ~n_9;
assign n_3177 =  x_335 &  n_9;
assign n_3178 = ~n_3176 & ~n_3177;
assign n_3179 =  x_1036 & ~n_3178;
assign n_3180 = ~x_1036 &  n_3178;
assign n_3181 = ~n_3179 & ~n_3180;
assign n_3182 =  x_1035 & ~n_9;
assign n_3183 =  x_334 &  n_9;
assign n_3184 = ~n_3182 & ~n_3183;
assign n_3185 =  x_1035 & ~n_3184;
assign n_3186 = ~x_1035 &  n_3184;
assign n_3187 = ~n_3185 & ~n_3186;
assign n_3188 =  x_1034 & ~n_9;
assign n_3189 =  x_333 &  n_9;
assign n_3190 = ~n_3188 & ~n_3189;
assign n_3191 =  x_1034 & ~n_3190;
assign n_3192 = ~x_1034 &  n_3190;
assign n_3193 = ~n_3191 & ~n_3192;
assign n_3194 =  x_1033 & ~n_9;
assign n_3195 =  x_332 &  n_9;
assign n_3196 = ~n_3194 & ~n_3195;
assign n_3197 =  x_1033 & ~n_3196;
assign n_3198 = ~x_1033 &  n_3196;
assign n_3199 = ~n_3197 & ~n_3198;
assign n_3200 =  x_1032 & ~n_9;
assign n_3201 =  x_331 &  n_9;
assign n_3202 = ~n_3200 & ~n_3201;
assign n_3203 =  x_1032 & ~n_3202;
assign n_3204 = ~x_1032 &  n_3202;
assign n_3205 = ~n_3203 & ~n_3204;
assign n_3206 =  x_1031 & ~n_9;
assign n_3207 =  x_330 &  n_9;
assign n_3208 = ~n_3206 & ~n_3207;
assign n_3209 =  x_1031 & ~n_3208;
assign n_3210 = ~x_1031 &  n_3208;
assign n_3211 = ~n_3209 & ~n_3210;
assign n_3212 =  x_902 &  n_1566;
assign n_3213 = ~n_1398 & ~n_1566;
assign n_3214 =  x_1030 &  n_3213;
assign n_3215 = ~n_3212 & ~n_3214;
assign n_3216 =  x_1030 & ~n_3215;
assign n_3217 = ~x_1030 &  n_3215;
assign n_3218 = ~n_3216 & ~n_3217;
assign n_3219 =  x_1029 &  n_3213;
assign n_3220 =  x_901 &  n_1566;
assign n_3221 = ~n_1401 & ~n_3220;
assign n_3222 = ~n_3219 &  n_3221;
assign n_3223 =  x_1029 & ~n_3222;
assign n_3224 = ~x_1029 &  n_3222;
assign n_3225 = ~n_3223 & ~n_3224;
assign n_3226 =  x_900 &  n_1566;
assign n_3227 =  x_1028 &  n_3213;
assign n_3228 = ~n_3226 & ~n_3227;
assign n_3229 =  x_1028 & ~n_3228;
assign n_3230 = ~x_1028 &  n_3228;
assign n_3231 = ~n_3229 & ~n_3230;
assign n_3232 =  x_899 &  n_1566;
assign n_3233 =  x_1027 &  n_3213;
assign n_3234 = ~n_3232 & ~n_3233;
assign n_3235 =  x_1027 & ~n_3234;
assign n_3236 = ~x_1027 &  n_3234;
assign n_3237 = ~n_3235 & ~n_3236;
assign n_3238 =  x_898 &  n_1566;
assign n_3239 =  x_1026 &  n_3213;
assign n_3240 = ~n_3238 & ~n_3239;
assign n_3241 =  x_1026 & ~n_3240;
assign n_3242 = ~x_1026 &  n_3240;
assign n_3243 = ~n_3241 & ~n_3242;
assign n_3244 =  x_1025 &  n_3213;
assign n_3245 =  x_897 &  n_1566;
assign n_3246 = ~n_1401 & ~n_3245;
assign n_3247 = ~n_3244 &  n_3246;
assign n_3248 =  x_1025 & ~n_3247;
assign n_3249 = ~x_1025 &  n_3247;
assign n_3250 = ~n_3248 & ~n_3249;
assign n_3251 =  x_896 &  n_1566;
assign n_3252 =  x_1024 &  n_3213;
assign n_3253 = ~n_3251 & ~n_3252;
assign n_3254 =  x_1024 & ~n_3253;
assign n_3255 = ~x_1024 &  n_3253;
assign n_3256 = ~n_3254 & ~n_3255;
assign n_3257 =  x_895 &  n_1566;
assign n_3258 =  x_1023 &  n_3213;
assign n_3259 = ~n_3257 & ~n_3258;
assign n_3260 =  x_1023 & ~n_3259;
assign n_3261 = ~x_1023 &  n_3259;
assign n_3262 = ~n_3260 & ~n_3261;
assign n_3263 =  x_894 &  n_1566;
assign n_3264 =  x_1022 &  n_3213;
assign n_3265 = ~n_3263 & ~n_3264;
assign n_3266 =  x_1022 & ~n_3265;
assign n_3267 = ~x_1022 &  n_3265;
assign n_3268 = ~n_3266 & ~n_3267;
assign n_3269 =  x_893 &  n_1566;
assign n_3270 =  x_1021 &  n_3213;
assign n_3271 = ~n_3269 & ~n_3270;
assign n_3272 =  x_1021 & ~n_3271;
assign n_3273 = ~x_1021 &  n_3271;
assign n_3274 = ~n_3272 & ~n_3273;
assign n_3275 =  x_1020 &  n_3213;
assign n_3276 =  x_892 &  n_1566;
assign n_3277 = ~n_1401 & ~n_3276;
assign n_3278 = ~n_3275 &  n_3277;
assign n_3279 =  x_1020 & ~n_3278;
assign n_3280 = ~x_1020 &  n_3278;
assign n_3281 = ~n_3279 & ~n_3280;
assign n_3282 =  x_891 &  n_1566;
assign n_3283 =  x_1019 &  n_3213;
assign n_3284 = ~n_3282 & ~n_3283;
assign n_3285 =  x_1019 & ~n_3284;
assign n_3286 = ~x_1019 &  n_3284;
assign n_3287 = ~n_3285 & ~n_3286;
assign n_3288 =  x_890 &  n_1566;
assign n_3289 =  x_1018 &  n_3213;
assign n_3290 = ~n_3288 & ~n_3289;
assign n_3291 =  x_1018 & ~n_3290;
assign n_3292 = ~x_1018 &  n_3290;
assign n_3293 = ~n_3291 & ~n_3292;
assign n_3294 =  x_889 &  n_1566;
assign n_3295 =  x_1017 &  n_3213;
assign n_3296 = ~n_3294 & ~n_3295;
assign n_3297 =  x_1017 & ~n_3296;
assign n_3298 = ~x_1017 &  n_3296;
assign n_3299 = ~n_3297 & ~n_3298;
assign n_3300 =  x_888 &  n_1566;
assign n_3301 =  x_1016 &  n_3213;
assign n_3302 = ~n_3300 & ~n_3301;
assign n_3303 =  x_1016 & ~n_3302;
assign n_3304 = ~x_1016 &  n_3302;
assign n_3305 = ~n_3303 & ~n_3304;
assign n_3306 =  x_887 &  n_1566;
assign n_3307 =  x_1015 &  n_3213;
assign n_3308 = ~n_3306 & ~n_3307;
assign n_3309 =  x_1015 & ~n_3308;
assign n_3310 = ~x_1015 &  n_3308;
assign n_3311 = ~n_3309 & ~n_3310;
assign n_3312 =  x_886 &  n_1566;
assign n_3313 =  x_1014 &  n_3213;
assign n_3314 = ~n_3312 & ~n_3313;
assign n_3315 =  x_1014 & ~n_3314;
assign n_3316 = ~x_1014 &  n_3314;
assign n_3317 = ~n_3315 & ~n_3316;
assign n_3318 =  x_885 &  n_1566;
assign n_3319 =  x_1013 &  n_3213;
assign n_3320 = ~n_3318 & ~n_3319;
assign n_3321 =  x_1013 & ~n_3320;
assign n_3322 = ~x_1013 &  n_3320;
assign n_3323 = ~n_3321 & ~n_3322;
assign n_3324 =  x_884 &  n_1566;
assign n_3325 =  x_1012 &  n_3213;
assign n_3326 = ~n_3324 & ~n_3325;
assign n_3327 =  x_1012 & ~n_3326;
assign n_3328 = ~x_1012 &  n_3326;
assign n_3329 = ~n_3327 & ~n_3328;
assign n_3330 =  x_883 &  n_1566;
assign n_3331 =  x_1011 &  n_3213;
assign n_3332 = ~n_3330 & ~n_3331;
assign n_3333 =  x_1011 & ~n_3332;
assign n_3334 = ~x_1011 &  n_3332;
assign n_3335 = ~n_3333 & ~n_3334;
assign n_3336 =  x_882 &  n_1566;
assign n_3337 =  x_1010 &  n_3213;
assign n_3338 = ~n_3336 & ~n_3337;
assign n_3339 =  x_1010 & ~n_3338;
assign n_3340 = ~x_1010 &  n_3338;
assign n_3341 = ~n_3339 & ~n_3340;
assign n_3342 =  x_881 &  n_1566;
assign n_3343 =  x_1009 &  n_3213;
assign n_3344 = ~n_3342 & ~n_3343;
assign n_3345 =  x_1009 & ~n_3344;
assign n_3346 = ~x_1009 &  n_3344;
assign n_3347 = ~n_3345 & ~n_3346;
assign n_3348 =  x_880 &  n_1566;
assign n_3349 =  x_1008 &  n_3213;
assign n_3350 = ~n_3348 & ~n_3349;
assign n_3351 =  x_1008 & ~n_3350;
assign n_3352 = ~x_1008 &  n_3350;
assign n_3353 = ~n_3351 & ~n_3352;
assign n_3354 =  x_879 &  n_1566;
assign n_3355 =  x_1007 &  n_3213;
assign n_3356 = ~n_3354 & ~n_3355;
assign n_3357 =  x_1007 & ~n_3356;
assign n_3358 = ~x_1007 &  n_3356;
assign n_3359 = ~n_3357 & ~n_3358;
assign n_3360 =  x_878 &  n_1566;
assign n_3361 =  x_1006 &  n_3213;
assign n_3362 = ~n_3360 & ~n_3361;
assign n_3363 =  x_1006 & ~n_3362;
assign n_3364 = ~x_1006 &  n_3362;
assign n_3365 = ~n_3363 & ~n_3364;
assign n_3366 =  x_877 &  n_1566;
assign n_3367 =  x_1005 &  n_3213;
assign n_3368 = ~n_3366 & ~n_3367;
assign n_3369 =  x_1005 & ~n_3368;
assign n_3370 = ~x_1005 &  n_3368;
assign n_3371 = ~n_3369 & ~n_3370;
assign n_3372 =  x_876 &  n_1566;
assign n_3373 =  x_1004 &  n_3213;
assign n_3374 = ~n_3372 & ~n_3373;
assign n_3375 =  x_1004 & ~n_3374;
assign n_3376 = ~x_1004 &  n_3374;
assign n_3377 = ~n_3375 & ~n_3376;
assign n_3378 =  x_875 &  n_1566;
assign n_3379 =  x_1003 &  n_3213;
assign n_3380 = ~n_3378 & ~n_3379;
assign n_3381 =  x_1003 & ~n_3380;
assign n_3382 = ~x_1003 &  n_3380;
assign n_3383 = ~n_3381 & ~n_3382;
assign n_3384 =  x_874 &  n_1566;
assign n_3385 =  x_1002 &  n_3213;
assign n_3386 = ~n_3384 & ~n_3385;
assign n_3387 =  x_1002 & ~n_3386;
assign n_3388 = ~x_1002 &  n_3386;
assign n_3389 = ~n_3387 & ~n_3388;
assign n_3390 =  x_873 &  n_1566;
assign n_3391 =  x_1001 &  n_3213;
assign n_3392 = ~n_3390 & ~n_3391;
assign n_3393 =  x_1001 & ~n_3392;
assign n_3394 = ~x_1001 &  n_3392;
assign n_3395 = ~n_3393 & ~n_3394;
assign n_3396 =  x_872 &  n_1566;
assign n_3397 =  x_1000 &  n_3213;
assign n_3398 = ~n_3396 & ~n_3397;
assign n_3399 =  x_1000 & ~n_3398;
assign n_3400 = ~x_1000 &  n_3398;
assign n_3401 = ~n_3399 & ~n_3400;
assign n_3402 =  x_871 &  n_1566;
assign n_3403 =  x_999 &  n_3213;
assign n_3404 = ~n_3402 & ~n_3403;
assign n_3405 =  x_999 & ~n_3404;
assign n_3406 = ~x_999 &  n_3404;
assign n_3407 = ~n_3405 & ~n_3406;
assign n_3408 =  x_998 & ~n_1270;
assign n_3409 = ~n_2828 & ~n_3408;
assign n_3410 =  x_998 & ~n_3409;
assign n_3411 = ~x_998 &  n_3409;
assign n_3412 = ~n_3410 & ~n_3411;
assign n_3413 =  x_997 & ~n_1270;
assign n_3414 = ~n_2834 & ~n_3413;
assign n_3415 =  x_997 & ~n_3414;
assign n_3416 = ~x_997 &  n_3414;
assign n_3417 = ~n_3415 & ~n_3416;
assign n_3418 =  x_996 & ~n_1270;
assign n_3419 = ~n_2840 & ~n_3418;
assign n_3420 =  x_996 & ~n_3419;
assign n_3421 = ~x_996 &  n_3419;
assign n_3422 = ~n_3420 & ~n_3421;
assign n_3423 =  x_995 & ~n_1270;
assign n_3424 = ~n_2846 & ~n_3423;
assign n_3425 =  x_995 & ~n_3424;
assign n_3426 = ~x_995 &  n_3424;
assign n_3427 = ~n_3425 & ~n_3426;
assign n_3428 =  x_994 & ~n_1270;
assign n_3429 = ~n_2852 & ~n_3428;
assign n_3430 =  x_994 & ~n_3429;
assign n_3431 = ~x_994 &  n_3429;
assign n_3432 = ~n_3430 & ~n_3431;
assign n_3433 =  x_993 & ~n_1270;
assign n_3434 = ~n_2858 & ~n_3433;
assign n_3435 =  x_993 & ~n_3434;
assign n_3436 = ~x_993 &  n_3434;
assign n_3437 = ~n_3435 & ~n_3436;
assign n_3438 =  x_992 & ~n_1270;
assign n_3439 = ~n_2864 & ~n_3438;
assign n_3440 =  x_992 & ~n_3439;
assign n_3441 = ~x_992 &  n_3439;
assign n_3442 = ~n_3440 & ~n_3441;
assign n_3443 =  x_991 & ~n_1270;
assign n_3444 = ~n_2870 & ~n_3443;
assign n_3445 =  x_991 & ~n_3444;
assign n_3446 = ~x_991 &  n_3444;
assign n_3447 = ~n_3445 & ~n_3446;
assign n_3448 =  x_990 & ~n_1270;
assign n_3449 = ~n_2876 & ~n_3448;
assign n_3450 =  x_990 & ~n_3449;
assign n_3451 = ~x_990 &  n_3449;
assign n_3452 = ~n_3450 & ~n_3451;
assign n_3453 =  x_989 & ~n_1270;
assign n_3454 = ~n_2882 & ~n_3453;
assign n_3455 =  x_989 & ~n_3454;
assign n_3456 = ~x_989 &  n_3454;
assign n_3457 = ~n_3455 & ~n_3456;
assign n_3458 =  x_988 & ~n_1270;
assign n_3459 = ~n_2888 & ~n_3458;
assign n_3460 =  x_988 & ~n_3459;
assign n_3461 = ~x_988 &  n_3459;
assign n_3462 = ~n_3460 & ~n_3461;
assign n_3463 =  x_987 & ~n_1270;
assign n_3464 = ~n_2894 & ~n_3463;
assign n_3465 =  x_987 & ~n_3464;
assign n_3466 = ~x_987 &  n_3464;
assign n_3467 = ~n_3465 & ~n_3466;
assign n_3468 =  x_986 & ~n_1270;
assign n_3469 = ~n_2900 & ~n_3468;
assign n_3470 =  x_986 & ~n_3469;
assign n_3471 = ~x_986 &  n_3469;
assign n_3472 = ~n_3470 & ~n_3471;
assign n_3473 =  x_985 & ~n_1270;
assign n_3474 = ~n_2906 & ~n_3473;
assign n_3475 =  x_985 & ~n_3474;
assign n_3476 = ~x_985 &  n_3474;
assign n_3477 = ~n_3475 & ~n_3476;
assign n_3478 =  x_984 & ~n_1270;
assign n_3479 = ~n_2912 & ~n_3478;
assign n_3480 =  x_984 & ~n_3479;
assign n_3481 = ~x_984 &  n_3479;
assign n_3482 = ~n_3480 & ~n_3481;
assign n_3483 =  x_983 & ~n_1270;
assign n_3484 = ~n_2918 & ~n_3483;
assign n_3485 =  x_983 & ~n_3484;
assign n_3486 = ~x_983 &  n_3484;
assign n_3487 = ~n_3485 & ~n_3486;
assign n_3488 =  x_982 & ~n_1270;
assign n_3489 = ~n_2924 & ~n_3488;
assign n_3490 =  x_982 & ~n_3489;
assign n_3491 = ~x_982 &  n_3489;
assign n_3492 = ~n_3490 & ~n_3491;
assign n_3493 =  x_981 & ~n_1270;
assign n_3494 = ~n_2930 & ~n_3493;
assign n_3495 =  x_981 & ~n_3494;
assign n_3496 = ~x_981 &  n_3494;
assign n_3497 = ~n_3495 & ~n_3496;
assign n_3498 =  x_980 & ~n_1270;
assign n_3499 = ~n_2936 & ~n_3498;
assign n_3500 =  x_980 & ~n_3499;
assign n_3501 = ~x_980 &  n_3499;
assign n_3502 = ~n_3500 & ~n_3501;
assign n_3503 =  x_979 & ~n_1270;
assign n_3504 = ~n_2942 & ~n_3503;
assign n_3505 =  x_979 & ~n_3504;
assign n_3506 = ~x_979 &  n_3504;
assign n_3507 = ~n_3505 & ~n_3506;
assign n_3508 =  x_978 & ~n_1270;
assign n_3509 = ~n_2948 & ~n_3508;
assign n_3510 =  x_978 & ~n_3509;
assign n_3511 = ~x_978 &  n_3509;
assign n_3512 = ~n_3510 & ~n_3511;
assign n_3513 =  x_977 & ~n_1270;
assign n_3514 = ~n_2954 & ~n_3513;
assign n_3515 =  x_977 & ~n_3514;
assign n_3516 = ~x_977 &  n_3514;
assign n_3517 = ~n_3515 & ~n_3516;
assign n_3518 =  x_976 & ~n_1270;
assign n_3519 = ~n_2960 & ~n_3518;
assign n_3520 =  x_976 & ~n_3519;
assign n_3521 = ~x_976 &  n_3519;
assign n_3522 = ~n_3520 & ~n_3521;
assign n_3523 =  x_747 & ~n_1531;
assign n_3524 =  i_4 &  n_1531;
assign n_3525 = ~n_3523 & ~n_3524;
assign n_3526 =  x_747 & ~n_3525;
assign n_3527 = ~x_747 &  n_3525;
assign n_3528 = ~n_3526 & ~n_3527;
assign n_3529 =  x_746 & ~n_1531;
assign n_3530 =  i_3 &  n_1531;
assign n_3531 = ~n_3529 & ~n_3530;
assign n_3532 =  x_746 & ~n_3531;
assign n_3533 = ~x_746 &  n_3531;
assign n_3534 = ~n_3532 & ~n_3533;
assign n_3535 =  x_745 & ~n_1531;
assign n_3536 =  i_2 &  n_1531;
assign n_3537 = ~n_3535 & ~n_3536;
assign n_3538 =  x_745 & ~n_3537;
assign n_3539 = ~x_745 &  n_3537;
assign n_3540 = ~n_3538 & ~n_3539;
assign n_3541 =  x_744 & ~n_1531;
assign n_3542 =  i_1 &  n_1531;
assign n_3543 = ~n_3541 & ~n_3542;
assign n_3544 =  x_744 & ~n_3543;
assign n_3545 = ~x_744 &  n_3543;
assign n_3546 = ~n_3544 & ~n_3545;
assign n_3547 =  x_743 & ~n_1328;
assign n_3548 =  i_32 &  n_1328;
assign n_3549 = ~n_3547 & ~n_3548;
assign n_3550 =  x_743 & ~n_3549;
assign n_3551 = ~x_743 &  n_3549;
assign n_3552 = ~n_3550 & ~n_3551;
assign n_3553 =  x_742 & ~n_1328;
assign n_3554 =  i_31 &  n_1328;
assign n_3555 = ~n_3553 & ~n_3554;
assign n_3556 =  x_742 & ~n_3555;
assign n_3557 = ~x_742 &  n_3555;
assign n_3558 = ~n_3556 & ~n_3557;
assign n_3559 =  x_741 & ~n_1328;
assign n_3560 =  i_30 &  n_1328;
assign n_3561 = ~n_3559 & ~n_3560;
assign n_3562 =  x_741 & ~n_3561;
assign n_3563 = ~x_741 &  n_3561;
assign n_3564 = ~n_3562 & ~n_3563;
assign n_3565 =  x_740 & ~n_1328;
assign n_3566 =  i_29 &  n_1328;
assign n_3567 = ~n_3565 & ~n_3566;
assign n_3568 =  x_740 & ~n_3567;
assign n_3569 = ~x_740 &  n_3567;
assign n_3570 = ~n_3568 & ~n_3569;
assign n_3571 =  x_739 & ~n_1328;
assign n_3572 =  i_28 &  n_1328;
assign n_3573 = ~n_3571 & ~n_3572;
assign n_3574 =  x_739 & ~n_3573;
assign n_3575 = ~x_739 &  n_3573;
assign n_3576 = ~n_3574 & ~n_3575;
assign n_3577 =  x_738 & ~n_1328;
assign n_3578 =  i_27 &  n_1328;
assign n_3579 = ~n_3577 & ~n_3578;
assign n_3580 =  x_738 & ~n_3579;
assign n_3581 = ~x_738 &  n_3579;
assign n_3582 = ~n_3580 & ~n_3581;
assign n_3583 =  x_737 & ~n_1328;
assign n_3584 =  i_26 &  n_1328;
assign n_3585 = ~n_3583 & ~n_3584;
assign n_3586 =  x_737 & ~n_3585;
assign n_3587 = ~x_737 &  n_3585;
assign n_3588 = ~n_3586 & ~n_3587;
assign n_3589 =  x_736 & ~n_1328;
assign n_3590 =  i_25 &  n_1328;
assign n_3591 = ~n_3589 & ~n_3590;
assign n_3592 =  x_736 & ~n_3591;
assign n_3593 = ~x_736 &  n_3591;
assign n_3594 = ~n_3592 & ~n_3593;
assign n_3595 =  x_735 & ~n_1328;
assign n_3596 =  i_24 &  n_1328;
assign n_3597 = ~n_3595 & ~n_3596;
assign n_3598 =  x_735 & ~n_3597;
assign n_3599 = ~x_735 &  n_3597;
assign n_3600 = ~n_3598 & ~n_3599;
assign n_3601 =  x_734 & ~n_1328;
assign n_3602 =  i_23 &  n_1328;
assign n_3603 = ~n_3601 & ~n_3602;
assign n_3604 =  x_734 & ~n_3603;
assign n_3605 = ~x_734 &  n_3603;
assign n_3606 = ~n_3604 & ~n_3605;
assign n_3607 =  x_733 & ~n_1328;
assign n_3608 =  i_22 &  n_1328;
assign n_3609 = ~n_3607 & ~n_3608;
assign n_3610 =  x_733 & ~n_3609;
assign n_3611 = ~x_733 &  n_3609;
assign n_3612 = ~n_3610 & ~n_3611;
assign n_3613 =  x_732 & ~n_1328;
assign n_3614 =  i_21 &  n_1328;
assign n_3615 = ~n_3613 & ~n_3614;
assign n_3616 =  x_732 & ~n_3615;
assign n_3617 = ~x_732 &  n_3615;
assign n_3618 = ~n_3616 & ~n_3617;
assign n_3619 =  x_731 & ~n_1328;
assign n_3620 =  i_20 &  n_1328;
assign n_3621 = ~n_3619 & ~n_3620;
assign n_3622 =  x_731 & ~n_3621;
assign n_3623 = ~x_731 &  n_3621;
assign n_3624 = ~n_3622 & ~n_3623;
assign n_3625 =  x_730 & ~n_1328;
assign n_3626 =  i_19 &  n_1328;
assign n_3627 = ~n_3625 & ~n_3626;
assign n_3628 =  x_730 & ~n_3627;
assign n_3629 = ~x_730 &  n_3627;
assign n_3630 = ~n_3628 & ~n_3629;
assign n_3631 =  x_729 & ~n_1328;
assign n_3632 =  i_18 &  n_1328;
assign n_3633 = ~n_3631 & ~n_3632;
assign n_3634 =  x_729 & ~n_3633;
assign n_3635 = ~x_729 &  n_3633;
assign n_3636 = ~n_3634 & ~n_3635;
assign n_3637 =  x_728 & ~n_1328;
assign n_3638 =  i_17 &  n_1328;
assign n_3639 = ~n_3637 & ~n_3638;
assign n_3640 =  x_728 & ~n_3639;
assign n_3641 = ~x_728 &  n_3639;
assign n_3642 = ~n_3640 & ~n_3641;
assign n_3643 =  x_727 & ~n_1328;
assign n_3644 =  i_16 &  n_1328;
assign n_3645 = ~n_3643 & ~n_3644;
assign n_3646 =  x_727 & ~n_3645;
assign n_3647 = ~x_727 &  n_3645;
assign n_3648 = ~n_3646 & ~n_3647;
assign n_3649 =  x_726 & ~n_1328;
assign n_3650 =  i_15 &  n_1328;
assign n_3651 = ~n_3649 & ~n_3650;
assign n_3652 =  x_726 & ~n_3651;
assign n_3653 = ~x_726 &  n_3651;
assign n_3654 = ~n_3652 & ~n_3653;
assign n_3655 =  x_725 & ~n_1328;
assign n_3656 =  i_14 &  n_1328;
assign n_3657 = ~n_3655 & ~n_3656;
assign n_3658 =  x_725 & ~n_3657;
assign n_3659 = ~x_725 &  n_3657;
assign n_3660 = ~n_3658 & ~n_3659;
assign n_3661 =  x_724 & ~n_1328;
assign n_3662 =  i_13 &  n_1328;
assign n_3663 = ~n_3661 & ~n_3662;
assign n_3664 =  x_724 & ~n_3663;
assign n_3665 = ~x_724 &  n_3663;
assign n_3666 = ~n_3664 & ~n_3665;
assign n_3667 =  x_723 & ~n_1328;
assign n_3668 =  i_12 &  n_1328;
assign n_3669 = ~n_3667 & ~n_3668;
assign n_3670 =  x_723 & ~n_3669;
assign n_3671 = ~x_723 &  n_3669;
assign n_3672 = ~n_3670 & ~n_3671;
assign n_3673 =  x_722 & ~n_1328;
assign n_3674 =  i_11 &  n_1328;
assign n_3675 = ~n_3673 & ~n_3674;
assign n_3676 =  x_722 & ~n_3675;
assign n_3677 = ~x_722 &  n_3675;
assign n_3678 = ~n_3676 & ~n_3677;
assign n_3679 =  x_721 & ~n_1328;
assign n_3680 =  i_10 &  n_1328;
assign n_3681 = ~n_3679 & ~n_3680;
assign n_3682 =  x_721 & ~n_3681;
assign n_3683 = ~x_721 &  n_3681;
assign n_3684 = ~n_3682 & ~n_3683;
assign n_3685 =  x_720 & ~n_1328;
assign n_3686 =  i_9 &  n_1328;
assign n_3687 = ~n_3685 & ~n_3686;
assign n_3688 =  x_720 & ~n_3687;
assign n_3689 = ~x_720 &  n_3687;
assign n_3690 = ~n_3688 & ~n_3689;
assign n_3691 =  x_719 & ~n_1328;
assign n_3692 =  i_8 &  n_1328;
assign n_3693 = ~n_3691 & ~n_3692;
assign n_3694 =  x_719 & ~n_3693;
assign n_3695 = ~x_719 &  n_3693;
assign n_3696 = ~n_3694 & ~n_3695;
assign n_3697 =  x_718 & ~n_1328;
assign n_3698 =  i_7 &  n_1328;
assign n_3699 = ~n_3697 & ~n_3698;
assign n_3700 =  x_718 & ~n_3699;
assign n_3701 = ~x_718 &  n_3699;
assign n_3702 = ~n_3700 & ~n_3701;
assign n_3703 =  x_717 & ~n_1328;
assign n_3704 =  i_6 &  n_1328;
assign n_3705 = ~n_3703 & ~n_3704;
assign n_3706 =  x_717 & ~n_3705;
assign n_3707 = ~x_717 &  n_3705;
assign n_3708 = ~n_3706 & ~n_3707;
assign n_3709 =  x_716 & ~n_1328;
assign n_3710 =  i_5 &  n_1328;
assign n_3711 = ~n_3709 & ~n_3710;
assign n_3712 =  x_716 & ~n_3711;
assign n_3713 = ~x_716 &  n_3711;
assign n_3714 = ~n_3712 & ~n_3713;
assign n_3715 =  x_715 & ~n_1328;
assign n_3716 =  i_4 &  n_1328;
assign n_3717 = ~n_3715 & ~n_3716;
assign n_3718 =  x_715 & ~n_3717;
assign n_3719 = ~x_715 &  n_3717;
assign n_3720 = ~n_3718 & ~n_3719;
assign n_3721 =  x_714 & ~n_1328;
assign n_3722 =  i_3 &  n_1328;
assign n_3723 = ~n_3721 & ~n_3722;
assign n_3724 =  x_714 & ~n_3723;
assign n_3725 = ~x_714 &  n_3723;
assign n_3726 = ~n_3724 & ~n_3725;
assign n_3727 =  x_713 & ~n_1328;
assign n_3728 =  i_2 &  n_1328;
assign n_3729 = ~n_3727 & ~n_3728;
assign n_3730 =  x_713 & ~n_3729;
assign n_3731 = ~x_713 &  n_3729;
assign n_3732 = ~n_3730 & ~n_3731;
assign n_3733 =  x_712 & ~n_1328;
assign n_3734 =  i_1 &  n_1328;
assign n_3735 = ~n_3733 & ~n_3734;
assign n_3736 =  x_712 & ~n_3735;
assign n_3737 = ~x_712 &  n_3735;
assign n_3738 = ~n_3736 & ~n_3737;
assign n_3739 =  x_711 & ~n_2125;
assign n_3740 =  i_32 &  n_2125;
assign n_3741 = ~n_3739 & ~n_3740;
assign n_3742 =  x_711 & ~n_3741;
assign n_3743 = ~x_711 &  n_3741;
assign n_3744 = ~n_3742 & ~n_3743;
assign n_3745 =  x_710 & ~n_2125;
assign n_3746 =  i_31 &  n_2125;
assign n_3747 = ~n_3745 & ~n_3746;
assign n_3748 =  x_710 & ~n_3747;
assign n_3749 = ~x_710 &  n_3747;
assign n_3750 = ~n_3748 & ~n_3749;
assign n_3751 =  x_709 & ~n_2125;
assign n_3752 =  i_30 &  n_2125;
assign n_3753 = ~n_3751 & ~n_3752;
assign n_3754 =  x_709 & ~n_3753;
assign n_3755 = ~x_709 &  n_3753;
assign n_3756 = ~n_3754 & ~n_3755;
assign n_3757 =  x_708 & ~n_2125;
assign n_3758 =  i_29 &  n_2125;
assign n_3759 = ~n_3757 & ~n_3758;
assign n_3760 =  x_708 & ~n_3759;
assign n_3761 = ~x_708 &  n_3759;
assign n_3762 = ~n_3760 & ~n_3761;
assign n_3763 =  x_707 & ~n_2125;
assign n_3764 =  i_28 &  n_2125;
assign n_3765 = ~n_3763 & ~n_3764;
assign n_3766 =  x_707 & ~n_3765;
assign n_3767 = ~x_707 &  n_3765;
assign n_3768 = ~n_3766 & ~n_3767;
assign n_3769 =  x_706 & ~n_2125;
assign n_3770 =  i_27 &  n_2125;
assign n_3771 = ~n_3769 & ~n_3770;
assign n_3772 =  x_706 & ~n_3771;
assign n_3773 = ~x_706 &  n_3771;
assign n_3774 = ~n_3772 & ~n_3773;
assign n_3775 =  x_705 & ~n_2125;
assign n_3776 =  i_26 &  n_2125;
assign n_3777 = ~n_3775 & ~n_3776;
assign n_3778 =  x_705 & ~n_3777;
assign n_3779 = ~x_705 &  n_3777;
assign n_3780 = ~n_3778 & ~n_3779;
assign n_3781 =  x_704 & ~n_2125;
assign n_3782 =  i_25 &  n_2125;
assign n_3783 = ~n_3781 & ~n_3782;
assign n_3784 =  x_704 & ~n_3783;
assign n_3785 = ~x_704 &  n_3783;
assign n_3786 = ~n_3784 & ~n_3785;
assign n_3787 =  x_703 & ~n_2125;
assign n_3788 =  i_24 &  n_2125;
assign n_3789 = ~n_3787 & ~n_3788;
assign n_3790 =  x_703 & ~n_3789;
assign n_3791 = ~x_703 &  n_3789;
assign n_3792 = ~n_3790 & ~n_3791;
assign n_3793 =  x_702 & ~n_2125;
assign n_3794 =  i_23 &  n_2125;
assign n_3795 = ~n_3793 & ~n_3794;
assign n_3796 =  x_702 & ~n_3795;
assign n_3797 = ~x_702 &  n_3795;
assign n_3798 = ~n_3796 & ~n_3797;
assign n_3799 =  x_701 & ~n_2125;
assign n_3800 =  i_22 &  n_2125;
assign n_3801 = ~n_3799 & ~n_3800;
assign n_3802 =  x_701 & ~n_3801;
assign n_3803 = ~x_701 &  n_3801;
assign n_3804 = ~n_3802 & ~n_3803;
assign n_3805 =  x_700 & ~n_2125;
assign n_3806 =  i_21 &  n_2125;
assign n_3807 = ~n_3805 & ~n_3806;
assign n_3808 =  x_700 & ~n_3807;
assign n_3809 = ~x_700 &  n_3807;
assign n_3810 = ~n_3808 & ~n_3809;
assign n_3811 =  x_699 & ~n_2125;
assign n_3812 =  i_20 &  n_2125;
assign n_3813 = ~n_3811 & ~n_3812;
assign n_3814 =  x_699 & ~n_3813;
assign n_3815 = ~x_699 &  n_3813;
assign n_3816 = ~n_3814 & ~n_3815;
assign n_3817 =  x_698 & ~n_2125;
assign n_3818 =  i_19 &  n_2125;
assign n_3819 = ~n_3817 & ~n_3818;
assign n_3820 =  x_698 & ~n_3819;
assign n_3821 = ~x_698 &  n_3819;
assign n_3822 = ~n_3820 & ~n_3821;
assign n_3823 =  x_697 & ~n_2125;
assign n_3824 =  i_18 &  n_2125;
assign n_3825 = ~n_3823 & ~n_3824;
assign n_3826 =  x_697 & ~n_3825;
assign n_3827 = ~x_697 &  n_3825;
assign n_3828 = ~n_3826 & ~n_3827;
assign n_3829 =  x_696 & ~n_2125;
assign n_3830 =  i_17 &  n_2125;
assign n_3831 = ~n_3829 & ~n_3830;
assign n_3832 =  x_696 & ~n_3831;
assign n_3833 = ~x_696 &  n_3831;
assign n_3834 = ~n_3832 & ~n_3833;
assign n_3835 =  x_695 & ~n_2125;
assign n_3836 =  i_16 &  n_2125;
assign n_3837 = ~n_3835 & ~n_3836;
assign n_3838 =  x_695 & ~n_3837;
assign n_3839 = ~x_695 &  n_3837;
assign n_3840 = ~n_3838 & ~n_3839;
assign n_3841 =  x_694 & ~n_2125;
assign n_3842 =  i_15 &  n_2125;
assign n_3843 = ~n_3841 & ~n_3842;
assign n_3844 =  x_694 & ~n_3843;
assign n_3845 = ~x_694 &  n_3843;
assign n_3846 = ~n_3844 & ~n_3845;
assign n_3847 =  x_693 & ~n_2125;
assign n_3848 =  i_14 &  n_2125;
assign n_3849 = ~n_3847 & ~n_3848;
assign n_3850 =  x_693 & ~n_3849;
assign n_3851 = ~x_693 &  n_3849;
assign n_3852 = ~n_3850 & ~n_3851;
assign n_3853 =  x_692 & ~n_2125;
assign n_3854 =  i_13 &  n_2125;
assign n_3855 = ~n_3853 & ~n_3854;
assign n_3856 =  x_692 & ~n_3855;
assign n_3857 = ~x_692 &  n_3855;
assign n_3858 = ~n_3856 & ~n_3857;
assign n_3859 =  x_691 & ~n_2125;
assign n_3860 =  i_12 &  n_2125;
assign n_3861 = ~n_3859 & ~n_3860;
assign n_3862 =  x_691 & ~n_3861;
assign n_3863 = ~x_691 &  n_3861;
assign n_3864 = ~n_3862 & ~n_3863;
assign n_3865 =  x_690 & ~n_2125;
assign n_3866 =  i_11 &  n_2125;
assign n_3867 = ~n_3865 & ~n_3866;
assign n_3868 =  x_690 & ~n_3867;
assign n_3869 = ~x_690 &  n_3867;
assign n_3870 = ~n_3868 & ~n_3869;
assign n_3871 =  x_689 & ~n_2125;
assign n_3872 =  i_10 &  n_2125;
assign n_3873 = ~n_3871 & ~n_3872;
assign n_3874 =  x_689 & ~n_3873;
assign n_3875 = ~x_689 &  n_3873;
assign n_3876 = ~n_3874 & ~n_3875;
assign n_3877 =  x_688 & ~n_2125;
assign n_3878 =  i_9 &  n_2125;
assign n_3879 = ~n_3877 & ~n_3878;
assign n_3880 =  x_688 & ~n_3879;
assign n_3881 = ~x_688 &  n_3879;
assign n_3882 = ~n_3880 & ~n_3881;
assign n_3883 =  x_687 & ~n_2125;
assign n_3884 =  i_8 &  n_2125;
assign n_3885 = ~n_3883 & ~n_3884;
assign n_3886 =  x_687 & ~n_3885;
assign n_3887 = ~x_687 &  n_3885;
assign n_3888 = ~n_3886 & ~n_3887;
assign n_3889 =  x_686 & ~n_2125;
assign n_3890 =  i_7 &  n_2125;
assign n_3891 = ~n_3889 & ~n_3890;
assign n_3892 =  x_686 & ~n_3891;
assign n_3893 = ~x_686 &  n_3891;
assign n_3894 = ~n_3892 & ~n_3893;
assign n_3895 =  x_685 & ~n_2125;
assign n_3896 =  i_6 &  n_2125;
assign n_3897 = ~n_3895 & ~n_3896;
assign n_3898 =  x_685 & ~n_3897;
assign n_3899 = ~x_685 &  n_3897;
assign n_3900 = ~n_3898 & ~n_3899;
assign n_3901 =  x_684 & ~n_2125;
assign n_3902 =  i_5 &  n_2125;
assign n_3903 = ~n_3901 & ~n_3902;
assign n_3904 =  x_684 & ~n_3903;
assign n_3905 = ~x_684 &  n_3903;
assign n_3906 = ~n_3904 & ~n_3905;
assign n_3907 =  x_683 & ~n_2125;
assign n_3908 =  i_4 &  n_2125;
assign n_3909 = ~n_3907 & ~n_3908;
assign n_3910 =  x_683 & ~n_3909;
assign n_3911 = ~x_683 &  n_3909;
assign n_3912 = ~n_3910 & ~n_3911;
assign n_3913 =  x_682 & ~n_2125;
assign n_3914 =  i_3 &  n_2125;
assign n_3915 = ~n_3913 & ~n_3914;
assign n_3916 =  x_682 & ~n_3915;
assign n_3917 = ~x_682 &  n_3915;
assign n_3918 = ~n_3916 & ~n_3917;
assign n_3919 =  x_681 & ~n_2125;
assign n_3920 =  i_2 &  n_2125;
assign n_3921 = ~n_3919 & ~n_3920;
assign n_3922 =  x_681 & ~n_3921;
assign n_3923 = ~x_681 &  n_3921;
assign n_3924 = ~n_3922 & ~n_3923;
assign n_3925 =  x_680 & ~n_2125;
assign n_3926 =  i_1 &  n_2125;
assign n_3927 = ~n_3925 & ~n_3926;
assign n_3928 =  x_680 & ~n_3927;
assign n_3929 = ~x_680 &  n_3927;
assign n_3930 = ~n_3928 & ~n_3929;
assign n_3931 =  x_870 &  n_2070;
assign n_3932 =  n_744 & ~n_1344;
assign n_3933 =  n_8 &  n_3932;
assign n_3934 =  x_679 & ~n_3933;
assign n_3935 = ~n_3931 & ~n_3934;
assign n_3936 =  x_679 & ~n_3935;
assign n_3937 = ~x_679 &  n_3935;
assign n_3938 = ~n_3936 & ~n_3937;
assign n_3939 =  x_869 &  n_2070;
assign n_3940 =  x_678 & ~n_3933;
assign n_3941 = ~n_3939 & ~n_3940;
assign n_3942 =  x_678 & ~n_3941;
assign n_3943 = ~x_678 &  n_3941;
assign n_3944 = ~n_3942 & ~n_3943;
assign n_3945 =  x_868 &  n_2070;
assign n_3946 =  x_677 & ~n_3933;
assign n_3947 = ~n_3945 & ~n_3946;
assign n_3948 =  x_677 & ~n_3947;
assign n_3949 = ~x_677 &  n_3947;
assign n_3950 = ~n_3948 & ~n_3949;
assign n_3951 =  x_867 &  n_2070;
assign n_3952 =  x_676 & ~n_3933;
assign n_3953 = ~n_3951 & ~n_3952;
assign n_3954 =  x_676 & ~n_3953;
assign n_3955 = ~x_676 &  n_3953;
assign n_3956 = ~n_3954 & ~n_3955;
assign n_3957 =  x_866 &  n_2070;
assign n_3958 =  x_675 & ~n_3933;
assign n_3959 = ~n_3957 & ~n_3958;
assign n_3960 =  x_675 & ~n_3959;
assign n_3961 = ~x_675 &  n_3959;
assign n_3962 = ~n_3960 & ~n_3961;
assign n_3963 =  x_865 &  n_2070;
assign n_3964 =  x_674 & ~n_3933;
assign n_3965 = ~n_3963 & ~n_3964;
assign n_3966 =  x_674 & ~n_3965;
assign n_3967 = ~x_674 &  n_3965;
assign n_3968 = ~n_3966 & ~n_3967;
assign n_3969 =  x_864 &  n_2070;
assign n_3970 =  x_673 & ~n_3933;
assign n_3971 = ~n_3969 & ~n_3970;
assign n_3972 =  x_673 & ~n_3971;
assign n_3973 = ~x_673 &  n_3971;
assign n_3974 = ~n_3972 & ~n_3973;
assign n_3975 =  x_863 &  n_2070;
assign n_3976 =  x_672 & ~n_3933;
assign n_3977 = ~n_3975 & ~n_3976;
assign n_3978 =  x_672 & ~n_3977;
assign n_3979 = ~x_672 &  n_3977;
assign n_3980 = ~n_3978 & ~n_3979;
assign n_3981 =  x_862 &  n_2070;
assign n_3982 =  x_671 & ~n_3933;
assign n_3983 = ~n_3981 & ~n_3982;
assign n_3984 =  x_671 & ~n_3983;
assign n_3985 = ~x_671 &  n_3983;
assign n_3986 = ~n_3984 & ~n_3985;
assign n_3987 =  x_861 &  n_2070;
assign n_3988 =  x_670 & ~n_3933;
assign n_3989 = ~n_3987 & ~n_3988;
assign n_3990 =  x_670 & ~n_3989;
assign n_3991 = ~x_670 &  n_3989;
assign n_3992 = ~n_3990 & ~n_3991;
assign n_3993 =  x_860 &  n_2070;
assign n_3994 =  x_669 & ~n_3933;
assign n_3995 = ~n_3993 & ~n_3994;
assign n_3996 =  x_669 & ~n_3995;
assign n_3997 = ~x_669 &  n_3995;
assign n_3998 = ~n_3996 & ~n_3997;
assign n_3999 =  x_859 &  n_2070;
assign n_4000 =  x_668 & ~n_3933;
assign n_4001 = ~n_3999 & ~n_4000;
assign n_4002 =  x_668 & ~n_4001;
assign n_4003 = ~x_668 &  n_4001;
assign n_4004 = ~n_4002 & ~n_4003;
assign n_4005 =  x_858 &  n_2070;
assign n_4006 =  x_667 & ~n_3933;
assign n_4007 = ~n_4005 & ~n_4006;
assign n_4008 =  x_667 & ~n_4007;
assign n_4009 = ~x_667 &  n_4007;
assign n_4010 = ~n_4008 & ~n_4009;
assign n_4011 =  x_857 &  n_2070;
assign n_4012 =  x_666 & ~n_3933;
assign n_4013 = ~n_4011 & ~n_4012;
assign n_4014 =  x_666 & ~n_4013;
assign n_4015 = ~x_666 &  n_4013;
assign n_4016 = ~n_4014 & ~n_4015;
assign n_4017 =  x_856 &  n_2070;
assign n_4018 =  x_665 & ~n_3933;
assign n_4019 = ~n_4017 & ~n_4018;
assign n_4020 =  x_665 & ~n_4019;
assign n_4021 = ~x_665 &  n_4019;
assign n_4022 = ~n_4020 & ~n_4021;
assign n_4023 =  x_855 &  n_2070;
assign n_4024 =  x_664 & ~n_3933;
assign n_4025 = ~n_4023 & ~n_4024;
assign n_4026 =  x_664 & ~n_4025;
assign n_4027 = ~x_664 &  n_4025;
assign n_4028 = ~n_4026 & ~n_4027;
assign n_4029 =  x_854 &  n_2070;
assign n_4030 =  x_663 & ~n_3933;
assign n_4031 = ~n_4029 & ~n_4030;
assign n_4032 =  x_663 & ~n_4031;
assign n_4033 = ~x_663 &  n_4031;
assign n_4034 = ~n_4032 & ~n_4033;
assign n_4035 =  x_853 &  n_2070;
assign n_4036 =  x_662 & ~n_3933;
assign n_4037 = ~n_4035 & ~n_4036;
assign n_4038 =  x_662 & ~n_4037;
assign n_4039 = ~x_662 &  n_4037;
assign n_4040 = ~n_4038 & ~n_4039;
assign n_4041 =  x_852 &  n_2070;
assign n_4042 =  x_661 & ~n_3933;
assign n_4043 = ~n_4041 & ~n_4042;
assign n_4044 =  x_661 & ~n_4043;
assign n_4045 = ~x_661 &  n_4043;
assign n_4046 = ~n_4044 & ~n_4045;
assign n_4047 =  x_851 &  n_2070;
assign n_4048 =  x_660 & ~n_3933;
assign n_4049 = ~n_4047 & ~n_4048;
assign n_4050 =  x_660 & ~n_4049;
assign n_4051 = ~x_660 &  n_4049;
assign n_4052 = ~n_4050 & ~n_4051;
assign n_4053 =  x_850 &  n_2070;
assign n_4054 =  x_659 & ~n_3933;
assign n_4055 = ~n_4053 & ~n_4054;
assign n_4056 =  x_659 & ~n_4055;
assign n_4057 = ~x_659 &  n_4055;
assign n_4058 = ~n_4056 & ~n_4057;
assign n_4059 =  x_849 &  n_2070;
assign n_4060 =  x_658 & ~n_3933;
assign n_4061 = ~n_4059 & ~n_4060;
assign n_4062 =  x_658 & ~n_4061;
assign n_4063 = ~x_658 &  n_4061;
assign n_4064 = ~n_4062 & ~n_4063;
assign n_4065 =  x_848 &  n_2070;
assign n_4066 =  x_657 & ~n_3933;
assign n_4067 = ~n_4065 & ~n_4066;
assign n_4068 =  x_657 & ~n_4067;
assign n_4069 = ~x_657 &  n_4067;
assign n_4070 = ~n_4068 & ~n_4069;
assign n_4071 =  x_847 &  n_2070;
assign n_4072 =  x_656 & ~n_3933;
assign n_4073 = ~n_4071 & ~n_4072;
assign n_4074 =  x_656 & ~n_4073;
assign n_4075 = ~x_656 &  n_4073;
assign n_4076 = ~n_4074 & ~n_4075;
assign n_4077 =  x_846 &  n_2070;
assign n_4078 =  x_655 & ~n_3933;
assign n_4079 = ~n_4077 & ~n_4078;
assign n_4080 =  x_655 & ~n_4079;
assign n_4081 = ~x_655 &  n_4079;
assign n_4082 = ~n_4080 & ~n_4081;
assign n_4083 =  x_845 &  n_2070;
assign n_4084 =  x_654 & ~n_3933;
assign n_4085 = ~n_4083 & ~n_4084;
assign n_4086 =  x_654 & ~n_4085;
assign n_4087 = ~x_654 &  n_4085;
assign n_4088 = ~n_4086 & ~n_4087;
assign n_4089 =  x_844 &  n_2070;
assign n_4090 =  x_653 & ~n_3933;
assign n_4091 = ~n_4089 & ~n_4090;
assign n_4092 =  x_653 & ~n_4091;
assign n_4093 = ~x_653 &  n_4091;
assign n_4094 = ~n_4092 & ~n_4093;
assign n_4095 =  x_843 &  n_2070;
assign n_4096 =  x_652 & ~n_3933;
assign n_4097 = ~n_4095 & ~n_4096;
assign n_4098 =  x_652 & ~n_4097;
assign n_4099 = ~x_652 &  n_4097;
assign n_4100 = ~n_4098 & ~n_4099;
assign n_4101 =  x_842 &  n_2070;
assign n_4102 =  x_651 & ~n_3933;
assign n_4103 = ~n_4101 & ~n_4102;
assign n_4104 =  x_651 & ~n_4103;
assign n_4105 = ~x_651 &  n_4103;
assign n_4106 = ~n_4104 & ~n_4105;
assign n_4107 =  x_841 &  n_2070;
assign n_4108 =  x_650 & ~n_3933;
assign n_4109 = ~n_4107 & ~n_4108;
assign n_4110 =  x_650 & ~n_4109;
assign n_4111 = ~x_650 &  n_4109;
assign n_4112 = ~n_4110 & ~n_4111;
assign n_4113 =  x_840 &  n_2070;
assign n_4114 =  x_649 & ~n_3933;
assign n_4115 = ~n_4113 & ~n_4114;
assign n_4116 =  x_649 & ~n_4115;
assign n_4117 = ~x_649 &  n_4115;
assign n_4118 = ~n_4116 & ~n_4117;
assign n_4119 =  x_839 &  n_2070;
assign n_4120 =  x_648 & ~n_3933;
assign n_4121 = ~n_4119 & ~n_4120;
assign n_4122 =  x_648 & ~n_4121;
assign n_4123 = ~x_648 &  n_4121;
assign n_4124 = ~n_4122 & ~n_4123;
assign n_4125 =  x_647 & ~n_2050;
assign n_4126 =  i_32 &  n_2050;
assign n_4127 = ~n_4125 & ~n_4126;
assign n_4128 =  x_647 & ~n_4127;
assign n_4129 = ~x_647 &  n_4127;
assign n_4130 = ~n_4128 & ~n_4129;
assign n_4131 =  x_646 & ~n_2050;
assign n_4132 =  i_31 &  n_2050;
assign n_4133 = ~n_4131 & ~n_4132;
assign n_4134 =  x_646 & ~n_4133;
assign n_4135 = ~x_646 &  n_4133;
assign n_4136 = ~n_4134 & ~n_4135;
assign n_4137 =  x_645 & ~n_2050;
assign n_4138 =  i_30 &  n_2050;
assign n_4139 = ~n_4137 & ~n_4138;
assign n_4140 =  x_645 & ~n_4139;
assign n_4141 = ~x_645 &  n_4139;
assign n_4142 = ~n_4140 & ~n_4141;
assign n_4143 =  x_644 & ~n_2050;
assign n_4144 =  i_29 &  n_2050;
assign n_4145 = ~n_4143 & ~n_4144;
assign n_4146 =  x_644 & ~n_4145;
assign n_4147 = ~x_644 &  n_4145;
assign n_4148 = ~n_4146 & ~n_4147;
assign n_4149 =  x_643 & ~n_2050;
assign n_4150 =  i_28 &  n_2050;
assign n_4151 = ~n_4149 & ~n_4150;
assign n_4152 =  x_643 & ~n_4151;
assign n_4153 = ~x_643 &  n_4151;
assign n_4154 = ~n_4152 & ~n_4153;
assign n_4155 =  x_642 & ~n_2050;
assign n_4156 =  i_27 &  n_2050;
assign n_4157 = ~n_4155 & ~n_4156;
assign n_4158 =  x_642 & ~n_4157;
assign n_4159 = ~x_642 &  n_4157;
assign n_4160 = ~n_4158 & ~n_4159;
assign n_4161 =  x_641 & ~n_2050;
assign n_4162 =  i_26 &  n_2050;
assign n_4163 = ~n_4161 & ~n_4162;
assign n_4164 =  x_641 & ~n_4163;
assign n_4165 = ~x_641 &  n_4163;
assign n_4166 = ~n_4164 & ~n_4165;
assign n_4167 =  x_640 & ~n_2050;
assign n_4168 =  i_25 &  n_2050;
assign n_4169 = ~n_4167 & ~n_4168;
assign n_4170 =  x_640 & ~n_4169;
assign n_4171 = ~x_640 &  n_4169;
assign n_4172 = ~n_4170 & ~n_4171;
assign n_4173 =  x_639 & ~n_2050;
assign n_4174 =  i_24 &  n_2050;
assign n_4175 = ~n_4173 & ~n_4174;
assign n_4176 =  x_639 & ~n_4175;
assign n_4177 = ~x_639 &  n_4175;
assign n_4178 = ~n_4176 & ~n_4177;
assign n_4179 =  x_638 & ~n_2050;
assign n_4180 =  i_23 &  n_2050;
assign n_4181 = ~n_4179 & ~n_4180;
assign n_4182 =  x_638 & ~n_4181;
assign n_4183 = ~x_638 &  n_4181;
assign n_4184 = ~n_4182 & ~n_4183;
assign n_4185 =  x_637 & ~n_2050;
assign n_4186 =  i_22 &  n_2050;
assign n_4187 = ~n_4185 & ~n_4186;
assign n_4188 =  x_637 & ~n_4187;
assign n_4189 = ~x_637 &  n_4187;
assign n_4190 = ~n_4188 & ~n_4189;
assign n_4191 =  x_636 & ~n_2050;
assign n_4192 =  i_21 &  n_2050;
assign n_4193 = ~n_4191 & ~n_4192;
assign n_4194 =  x_636 & ~n_4193;
assign n_4195 = ~x_636 &  n_4193;
assign n_4196 = ~n_4194 & ~n_4195;
assign n_4197 =  x_635 & ~n_2050;
assign n_4198 =  i_20 &  n_2050;
assign n_4199 = ~n_4197 & ~n_4198;
assign n_4200 =  x_635 & ~n_4199;
assign n_4201 = ~x_635 &  n_4199;
assign n_4202 = ~n_4200 & ~n_4201;
assign n_4203 =  x_634 & ~n_2050;
assign n_4204 =  i_19 &  n_2050;
assign n_4205 = ~n_4203 & ~n_4204;
assign n_4206 =  x_634 & ~n_4205;
assign n_4207 = ~x_634 &  n_4205;
assign n_4208 = ~n_4206 & ~n_4207;
assign n_4209 =  x_633 & ~n_2050;
assign n_4210 =  i_18 &  n_2050;
assign n_4211 = ~n_4209 & ~n_4210;
assign n_4212 =  x_633 & ~n_4211;
assign n_4213 = ~x_633 &  n_4211;
assign n_4214 = ~n_4212 & ~n_4213;
assign n_4215 =  x_632 & ~n_2050;
assign n_4216 =  i_17 &  n_2050;
assign n_4217 = ~n_4215 & ~n_4216;
assign n_4218 =  x_632 & ~n_4217;
assign n_4219 = ~x_632 &  n_4217;
assign n_4220 = ~n_4218 & ~n_4219;
assign n_4221 =  x_631 & ~n_2050;
assign n_4222 =  i_16 &  n_2050;
assign n_4223 = ~n_4221 & ~n_4222;
assign n_4224 =  x_631 & ~n_4223;
assign n_4225 = ~x_631 &  n_4223;
assign n_4226 = ~n_4224 & ~n_4225;
assign n_4227 =  x_630 & ~n_2050;
assign n_4228 =  i_15 &  n_2050;
assign n_4229 = ~n_4227 & ~n_4228;
assign n_4230 =  x_630 & ~n_4229;
assign n_4231 = ~x_630 &  n_4229;
assign n_4232 = ~n_4230 & ~n_4231;
assign n_4233 =  x_629 & ~n_2050;
assign n_4234 =  i_14 &  n_2050;
assign n_4235 = ~n_4233 & ~n_4234;
assign n_4236 =  x_629 & ~n_4235;
assign n_4237 = ~x_629 &  n_4235;
assign n_4238 = ~n_4236 & ~n_4237;
assign n_4239 =  x_628 & ~n_2050;
assign n_4240 =  i_13 &  n_2050;
assign n_4241 = ~n_4239 & ~n_4240;
assign n_4242 =  x_628 & ~n_4241;
assign n_4243 = ~x_628 &  n_4241;
assign n_4244 = ~n_4242 & ~n_4243;
assign n_4245 =  x_627 & ~n_2050;
assign n_4246 =  i_12 &  n_2050;
assign n_4247 = ~n_4245 & ~n_4246;
assign n_4248 =  x_627 & ~n_4247;
assign n_4249 = ~x_627 &  n_4247;
assign n_4250 = ~n_4248 & ~n_4249;
assign n_4251 =  x_626 & ~n_2050;
assign n_4252 =  i_11 &  n_2050;
assign n_4253 = ~n_4251 & ~n_4252;
assign n_4254 =  x_626 & ~n_4253;
assign n_4255 = ~x_626 &  n_4253;
assign n_4256 = ~n_4254 & ~n_4255;
assign n_4257 =  x_625 & ~n_2050;
assign n_4258 =  i_10 &  n_2050;
assign n_4259 = ~n_4257 & ~n_4258;
assign n_4260 =  x_625 & ~n_4259;
assign n_4261 = ~x_625 &  n_4259;
assign n_4262 = ~n_4260 & ~n_4261;
assign n_4263 =  x_624 & ~n_2050;
assign n_4264 =  i_9 &  n_2050;
assign n_4265 = ~n_4263 & ~n_4264;
assign n_4266 =  x_624 & ~n_4265;
assign n_4267 = ~x_624 &  n_4265;
assign n_4268 = ~n_4266 & ~n_4267;
assign n_4269 =  x_623 & ~n_2050;
assign n_4270 =  i_8 &  n_2050;
assign n_4271 = ~n_4269 & ~n_4270;
assign n_4272 =  x_623 & ~n_4271;
assign n_4273 = ~x_623 &  n_4271;
assign n_4274 = ~n_4272 & ~n_4273;
assign n_4275 =  x_622 & ~n_2050;
assign n_4276 =  i_7 &  n_2050;
assign n_4277 = ~n_4275 & ~n_4276;
assign n_4278 =  x_622 & ~n_4277;
assign n_4279 = ~x_622 &  n_4277;
assign n_4280 = ~n_4278 & ~n_4279;
assign n_4281 =  x_621 & ~n_2050;
assign n_4282 =  i_6 &  n_2050;
assign n_4283 = ~n_4281 & ~n_4282;
assign n_4284 =  x_621 & ~n_4283;
assign n_4285 = ~x_621 &  n_4283;
assign n_4286 = ~n_4284 & ~n_4285;
assign n_4287 =  x_620 & ~n_2050;
assign n_4288 =  i_5 &  n_2050;
assign n_4289 = ~n_4287 & ~n_4288;
assign n_4290 =  x_620 & ~n_4289;
assign n_4291 = ~x_620 &  n_4289;
assign n_4292 = ~n_4290 & ~n_4291;
assign n_4293 =  x_619 & ~n_2050;
assign n_4294 =  i_4 &  n_2050;
assign n_4295 = ~n_4293 & ~n_4294;
assign n_4296 =  x_619 & ~n_4295;
assign n_4297 = ~x_619 &  n_4295;
assign n_4298 = ~n_4296 & ~n_4297;
assign n_4299 =  x_618 & ~n_2050;
assign n_4300 =  i_3 &  n_2050;
assign n_4301 = ~n_4299 & ~n_4300;
assign n_4302 =  x_618 & ~n_4301;
assign n_4303 = ~x_618 &  n_4301;
assign n_4304 = ~n_4302 & ~n_4303;
assign n_4305 =  x_617 & ~n_2050;
assign n_4306 =  i_2 &  n_2050;
assign n_4307 = ~n_4305 & ~n_4306;
assign n_4308 =  x_617 & ~n_4307;
assign n_4309 = ~x_617 &  n_4307;
assign n_4310 = ~n_4308 & ~n_4309;
assign n_4311 =  x_616 & ~n_2050;
assign n_4312 =  i_1 &  n_2050;
assign n_4313 = ~n_4311 & ~n_4312;
assign n_4314 =  x_616 & ~n_4313;
assign n_4315 = ~x_616 &  n_4313;
assign n_4316 = ~n_4314 & ~n_4315;
assign n_4317 =  x_615 & ~n_1683;
assign n_4318 =  i_32 &  n_1683;
assign n_4319 = ~n_4317 & ~n_4318;
assign n_4320 =  x_615 & ~n_4319;
assign n_4321 = ~x_615 &  n_4319;
assign n_4322 = ~n_4320 & ~n_4321;
assign n_4323 =  x_614 & ~n_1683;
assign n_4324 =  i_31 &  n_1683;
assign n_4325 = ~n_4323 & ~n_4324;
assign n_4326 =  x_614 & ~n_4325;
assign n_4327 = ~x_614 &  n_4325;
assign n_4328 = ~n_4326 & ~n_4327;
assign n_4329 =  x_613 & ~n_1683;
assign n_4330 =  i_30 &  n_1683;
assign n_4331 = ~n_4329 & ~n_4330;
assign n_4332 =  x_613 & ~n_4331;
assign n_4333 = ~x_613 &  n_4331;
assign n_4334 = ~n_4332 & ~n_4333;
assign n_4335 =  x_612 & ~n_1683;
assign n_4336 =  i_29 &  n_1683;
assign n_4337 = ~n_4335 & ~n_4336;
assign n_4338 =  x_612 & ~n_4337;
assign n_4339 = ~x_612 &  n_4337;
assign n_4340 = ~n_4338 & ~n_4339;
assign n_4341 =  x_611 & ~n_1683;
assign n_4342 =  i_28 &  n_1683;
assign n_4343 = ~n_4341 & ~n_4342;
assign n_4344 =  x_611 & ~n_4343;
assign n_4345 = ~x_611 &  n_4343;
assign n_4346 = ~n_4344 & ~n_4345;
assign n_4347 =  x_610 & ~n_1683;
assign n_4348 =  i_27 &  n_1683;
assign n_4349 = ~n_4347 & ~n_4348;
assign n_4350 =  x_610 & ~n_4349;
assign n_4351 = ~x_610 &  n_4349;
assign n_4352 = ~n_4350 & ~n_4351;
assign n_4353 =  x_609 & ~n_1683;
assign n_4354 =  i_26 &  n_1683;
assign n_4355 = ~n_4353 & ~n_4354;
assign n_4356 =  x_609 & ~n_4355;
assign n_4357 = ~x_609 &  n_4355;
assign n_4358 = ~n_4356 & ~n_4357;
assign n_4359 =  x_608 & ~n_1683;
assign n_4360 =  i_25 &  n_1683;
assign n_4361 = ~n_4359 & ~n_4360;
assign n_4362 =  x_608 & ~n_4361;
assign n_4363 = ~x_608 &  n_4361;
assign n_4364 = ~n_4362 & ~n_4363;
assign n_4365 =  x_607 & ~n_1683;
assign n_4366 =  i_24 &  n_1683;
assign n_4367 = ~n_4365 & ~n_4366;
assign n_4368 =  x_607 & ~n_4367;
assign n_4369 = ~x_607 &  n_4367;
assign n_4370 = ~n_4368 & ~n_4369;
assign n_4371 =  x_606 & ~n_1683;
assign n_4372 =  i_23 &  n_1683;
assign n_4373 = ~n_4371 & ~n_4372;
assign n_4374 =  x_606 & ~n_4373;
assign n_4375 = ~x_606 &  n_4373;
assign n_4376 = ~n_4374 & ~n_4375;
assign n_4377 =  x_605 & ~n_1683;
assign n_4378 =  i_22 &  n_1683;
assign n_4379 = ~n_4377 & ~n_4378;
assign n_4380 =  x_605 & ~n_4379;
assign n_4381 = ~x_605 &  n_4379;
assign n_4382 = ~n_4380 & ~n_4381;
assign n_4383 =  x_604 & ~n_1683;
assign n_4384 =  i_21 &  n_1683;
assign n_4385 = ~n_4383 & ~n_4384;
assign n_4386 =  x_604 & ~n_4385;
assign n_4387 = ~x_604 &  n_4385;
assign n_4388 = ~n_4386 & ~n_4387;
assign n_4389 =  x_603 & ~n_1683;
assign n_4390 =  i_20 &  n_1683;
assign n_4391 = ~n_4389 & ~n_4390;
assign n_4392 =  x_603 & ~n_4391;
assign n_4393 = ~x_603 &  n_4391;
assign n_4394 = ~n_4392 & ~n_4393;
assign n_4395 =  x_602 & ~n_1683;
assign n_4396 =  i_19 &  n_1683;
assign n_4397 = ~n_4395 & ~n_4396;
assign n_4398 =  x_602 & ~n_4397;
assign n_4399 = ~x_602 &  n_4397;
assign n_4400 = ~n_4398 & ~n_4399;
assign n_4401 =  x_601 & ~n_1683;
assign n_4402 =  i_18 &  n_1683;
assign n_4403 = ~n_4401 & ~n_4402;
assign n_4404 =  x_601 & ~n_4403;
assign n_4405 = ~x_601 &  n_4403;
assign n_4406 = ~n_4404 & ~n_4405;
assign n_4407 =  x_600 & ~n_1683;
assign n_4408 =  i_17 &  n_1683;
assign n_4409 = ~n_4407 & ~n_4408;
assign n_4410 =  x_600 & ~n_4409;
assign n_4411 = ~x_600 &  n_4409;
assign n_4412 = ~n_4410 & ~n_4411;
assign n_4413 =  x_599 & ~n_1683;
assign n_4414 =  i_16 &  n_1683;
assign n_4415 = ~n_4413 & ~n_4414;
assign n_4416 =  x_599 & ~n_4415;
assign n_4417 = ~x_599 &  n_4415;
assign n_4418 = ~n_4416 & ~n_4417;
assign n_4419 =  x_598 & ~n_1683;
assign n_4420 =  i_15 &  n_1683;
assign n_4421 = ~n_4419 & ~n_4420;
assign n_4422 =  x_598 & ~n_4421;
assign n_4423 = ~x_598 &  n_4421;
assign n_4424 = ~n_4422 & ~n_4423;
assign n_4425 =  x_597 & ~n_1683;
assign n_4426 =  i_14 &  n_1683;
assign n_4427 = ~n_4425 & ~n_4426;
assign n_4428 =  x_597 & ~n_4427;
assign n_4429 = ~x_597 &  n_4427;
assign n_4430 = ~n_4428 & ~n_4429;
assign n_4431 =  x_596 & ~n_1683;
assign n_4432 =  i_13 &  n_1683;
assign n_4433 = ~n_4431 & ~n_4432;
assign n_4434 =  x_596 & ~n_4433;
assign n_4435 = ~x_596 &  n_4433;
assign n_4436 = ~n_4434 & ~n_4435;
assign n_4437 =  x_595 & ~n_1683;
assign n_4438 =  i_12 &  n_1683;
assign n_4439 = ~n_4437 & ~n_4438;
assign n_4440 =  x_595 & ~n_4439;
assign n_4441 = ~x_595 &  n_4439;
assign n_4442 = ~n_4440 & ~n_4441;
assign n_4443 =  x_594 & ~n_1683;
assign n_4444 =  i_11 &  n_1683;
assign n_4445 = ~n_4443 & ~n_4444;
assign n_4446 =  x_594 & ~n_4445;
assign n_4447 = ~x_594 &  n_4445;
assign n_4448 = ~n_4446 & ~n_4447;
assign n_4449 =  x_593 & ~n_1683;
assign n_4450 =  i_10 &  n_1683;
assign n_4451 = ~n_4449 & ~n_4450;
assign n_4452 =  x_593 & ~n_4451;
assign n_4453 = ~x_593 &  n_4451;
assign n_4454 = ~n_4452 & ~n_4453;
assign n_4455 =  x_592 & ~n_1683;
assign n_4456 =  i_9 &  n_1683;
assign n_4457 = ~n_4455 & ~n_4456;
assign n_4458 =  x_592 & ~n_4457;
assign n_4459 = ~x_592 &  n_4457;
assign n_4460 = ~n_4458 & ~n_4459;
assign n_4461 =  x_591 & ~n_1683;
assign n_4462 =  i_8 &  n_1683;
assign n_4463 = ~n_4461 & ~n_4462;
assign n_4464 =  x_591 & ~n_4463;
assign n_4465 = ~x_591 &  n_4463;
assign n_4466 = ~n_4464 & ~n_4465;
assign n_4467 =  x_590 & ~n_1683;
assign n_4468 =  i_7 &  n_1683;
assign n_4469 = ~n_4467 & ~n_4468;
assign n_4470 =  x_590 & ~n_4469;
assign n_4471 = ~x_590 &  n_4469;
assign n_4472 = ~n_4470 & ~n_4471;
assign n_4473 =  x_589 & ~n_1683;
assign n_4474 =  i_6 &  n_1683;
assign n_4475 = ~n_4473 & ~n_4474;
assign n_4476 =  x_589 & ~n_4475;
assign n_4477 = ~x_589 &  n_4475;
assign n_4478 = ~n_4476 & ~n_4477;
assign n_4479 =  x_588 & ~n_1683;
assign n_4480 =  i_5 &  n_1683;
assign n_4481 = ~n_4479 & ~n_4480;
assign n_4482 =  x_588 & ~n_4481;
assign n_4483 = ~x_588 &  n_4481;
assign n_4484 = ~n_4482 & ~n_4483;
assign n_4485 =  x_587 & ~n_1683;
assign n_4486 =  i_4 &  n_1683;
assign n_4487 = ~n_4485 & ~n_4486;
assign n_4488 =  x_587 & ~n_4487;
assign n_4489 = ~x_587 &  n_4487;
assign n_4490 = ~n_4488 & ~n_4489;
assign n_4491 =  x_586 & ~n_1683;
assign n_4492 =  i_3 &  n_1683;
assign n_4493 = ~n_4491 & ~n_4492;
assign n_4494 =  x_586 & ~n_4493;
assign n_4495 = ~x_586 &  n_4493;
assign n_4496 = ~n_4494 & ~n_4495;
assign n_4497 =  x_585 & ~n_1683;
assign n_4498 =  i_2 &  n_1683;
assign n_4499 = ~n_4497 & ~n_4498;
assign n_4500 =  x_585 & ~n_4499;
assign n_4501 = ~x_585 &  n_4499;
assign n_4502 = ~n_4500 & ~n_4501;
assign n_4503 =  x_584 & ~n_1683;
assign n_4504 =  i_1 &  n_1683;
assign n_4505 = ~n_4503 & ~n_4504;
assign n_4506 =  x_584 & ~n_4505;
assign n_4507 = ~x_584 &  n_4505;
assign n_4508 = ~n_4506 & ~n_4507;
assign n_4509 =  x_583 & ~n_1398;
assign n_4510 =  x_902 &  n_1401;
assign n_4511 = ~n_4509 & ~n_4510;
assign n_4512 =  x_583 & ~n_4511;
assign n_4513 = ~x_583 &  n_4511;
assign n_4514 = ~n_4512 & ~n_4513;
assign n_4515 =  x_582 & ~n_1398;
assign n_4516 =  x_901 &  n_1401;
assign n_4517 = ~n_4515 & ~n_4516;
assign n_4518 =  x_582 & ~n_4517;
assign n_4519 = ~x_582 &  n_4517;
assign n_4520 = ~n_4518 & ~n_4519;
assign n_4521 =  x_581 & ~n_1398;
assign n_4522 =  x_900 &  n_1401;
assign n_4523 = ~n_4521 & ~n_4522;
assign n_4524 =  x_581 & ~n_4523;
assign n_4525 = ~x_581 &  n_4523;
assign n_4526 = ~n_4524 & ~n_4525;
assign n_4527 =  x_580 & ~n_1398;
assign n_4528 =  x_899 &  n_1401;
assign n_4529 = ~n_4527 & ~n_4528;
assign n_4530 =  x_580 & ~n_4529;
assign n_4531 = ~x_580 &  n_4529;
assign n_4532 = ~n_4530 & ~n_4531;
assign n_4533 =  x_579 & ~n_1398;
assign n_4534 =  x_898 &  n_1401;
assign n_4535 = ~n_4533 & ~n_4534;
assign n_4536 =  x_579 & ~n_4535;
assign n_4537 = ~x_579 &  n_4535;
assign n_4538 = ~n_4536 & ~n_4537;
assign n_4539 =  x_578 & ~n_1398;
assign n_4540 =  x_897 &  n_1401;
assign n_4541 = ~n_4539 & ~n_4540;
assign n_4542 =  x_578 & ~n_4541;
assign n_4543 = ~x_578 &  n_4541;
assign n_4544 = ~n_4542 & ~n_4543;
assign n_4545 =  x_577 & ~n_1398;
assign n_4546 =  x_896 &  n_1401;
assign n_4547 = ~n_4545 & ~n_4546;
assign n_4548 =  x_577 & ~n_4547;
assign n_4549 = ~x_577 &  n_4547;
assign n_4550 = ~n_4548 & ~n_4549;
assign n_4551 =  x_576 & ~n_1398;
assign n_4552 =  x_895 &  n_1401;
assign n_4553 = ~n_4551 & ~n_4552;
assign n_4554 =  x_576 & ~n_4553;
assign n_4555 = ~x_576 &  n_4553;
assign n_4556 = ~n_4554 & ~n_4555;
assign n_4557 =  x_575 & ~n_1398;
assign n_4558 =  x_894 &  n_1401;
assign n_4559 = ~n_4557 & ~n_4558;
assign n_4560 =  x_575 & ~n_4559;
assign n_4561 = ~x_575 &  n_4559;
assign n_4562 = ~n_4560 & ~n_4561;
assign n_4563 =  x_574 & ~n_1398;
assign n_4564 =  x_893 &  n_1401;
assign n_4565 = ~n_4563 & ~n_4564;
assign n_4566 =  x_574 & ~n_4565;
assign n_4567 = ~x_574 &  n_4565;
assign n_4568 = ~n_4566 & ~n_4567;
assign n_4569 =  x_573 & ~n_1398;
assign n_4570 =  x_892 &  n_1401;
assign n_4571 = ~n_4569 & ~n_4570;
assign n_4572 =  x_573 & ~n_4571;
assign n_4573 = ~x_573 &  n_4571;
assign n_4574 = ~n_4572 & ~n_4573;
assign n_4575 =  x_572 & ~n_1398;
assign n_4576 =  x_891 &  n_1401;
assign n_4577 = ~n_4575 & ~n_4576;
assign n_4578 =  x_572 & ~n_4577;
assign n_4579 = ~x_572 &  n_4577;
assign n_4580 = ~n_4578 & ~n_4579;
assign n_4581 =  x_571 & ~n_1398;
assign n_4582 =  x_890 &  n_1401;
assign n_4583 = ~n_4581 & ~n_4582;
assign n_4584 =  x_571 & ~n_4583;
assign n_4585 = ~x_571 &  n_4583;
assign n_4586 = ~n_4584 & ~n_4585;
assign n_4587 =  x_570 & ~n_1398;
assign n_4588 =  x_889 &  n_1401;
assign n_4589 = ~n_4587 & ~n_4588;
assign n_4590 =  x_570 & ~n_4589;
assign n_4591 = ~x_570 &  n_4589;
assign n_4592 = ~n_4590 & ~n_4591;
assign n_4593 =  x_569 & ~n_1398;
assign n_4594 =  x_888 &  n_1401;
assign n_4595 = ~n_4593 & ~n_4594;
assign n_4596 =  x_569 & ~n_4595;
assign n_4597 = ~x_569 &  n_4595;
assign n_4598 = ~n_4596 & ~n_4597;
assign n_4599 =  x_568 & ~n_1398;
assign n_4600 =  x_887 &  n_1401;
assign n_4601 = ~n_4599 & ~n_4600;
assign n_4602 =  x_568 & ~n_4601;
assign n_4603 = ~x_568 &  n_4601;
assign n_4604 = ~n_4602 & ~n_4603;
assign n_4605 =  x_567 & ~n_1398;
assign n_4606 =  x_886 &  n_1401;
assign n_4607 = ~n_4605 & ~n_4606;
assign n_4608 =  x_567 & ~n_4607;
assign n_4609 = ~x_567 &  n_4607;
assign n_4610 = ~n_4608 & ~n_4609;
assign n_4611 =  x_566 & ~n_1398;
assign n_4612 =  x_885 &  n_1401;
assign n_4613 = ~n_4611 & ~n_4612;
assign n_4614 =  x_566 & ~n_4613;
assign n_4615 = ~x_566 &  n_4613;
assign n_4616 = ~n_4614 & ~n_4615;
assign n_4617 =  x_565 & ~n_1398;
assign n_4618 =  x_884 &  n_1401;
assign n_4619 = ~n_4617 & ~n_4618;
assign n_4620 =  x_565 & ~n_4619;
assign n_4621 = ~x_565 &  n_4619;
assign n_4622 = ~n_4620 & ~n_4621;
assign n_4623 =  x_564 & ~n_1398;
assign n_4624 =  x_883 &  n_1401;
assign n_4625 = ~n_4623 & ~n_4624;
assign n_4626 =  x_564 & ~n_4625;
assign n_4627 = ~x_564 &  n_4625;
assign n_4628 = ~n_4626 & ~n_4627;
assign n_4629 =  x_563 & ~n_1398;
assign n_4630 =  x_882 &  n_1401;
assign n_4631 = ~n_4629 & ~n_4630;
assign n_4632 =  x_563 & ~n_4631;
assign n_4633 = ~x_563 &  n_4631;
assign n_4634 = ~n_4632 & ~n_4633;
assign n_4635 =  x_562 & ~n_1398;
assign n_4636 =  x_881 &  n_1401;
assign n_4637 = ~n_4635 & ~n_4636;
assign n_4638 =  x_562 & ~n_4637;
assign n_4639 = ~x_562 &  n_4637;
assign n_4640 = ~n_4638 & ~n_4639;
assign n_4641 =  x_561 & ~n_1398;
assign n_4642 =  x_880 &  n_1401;
assign n_4643 = ~n_4641 & ~n_4642;
assign n_4644 =  x_561 & ~n_4643;
assign n_4645 = ~x_561 &  n_4643;
assign n_4646 = ~n_4644 & ~n_4645;
assign n_4647 =  x_560 & ~n_1398;
assign n_4648 =  x_879 &  n_1401;
assign n_4649 = ~n_4647 & ~n_4648;
assign n_4650 =  x_560 & ~n_4649;
assign n_4651 = ~x_560 &  n_4649;
assign n_4652 = ~n_4650 & ~n_4651;
assign n_4653 =  x_559 & ~n_1398;
assign n_4654 =  x_878 &  n_1401;
assign n_4655 = ~n_4653 & ~n_4654;
assign n_4656 =  x_559 & ~n_4655;
assign n_4657 = ~x_559 &  n_4655;
assign n_4658 = ~n_4656 & ~n_4657;
assign n_4659 =  x_558 & ~n_1398;
assign n_4660 =  x_877 &  n_1401;
assign n_4661 = ~n_4659 & ~n_4660;
assign n_4662 =  x_558 & ~n_4661;
assign n_4663 = ~x_558 &  n_4661;
assign n_4664 = ~n_4662 & ~n_4663;
assign n_4665 =  x_557 & ~n_1398;
assign n_4666 =  x_876 &  n_1401;
assign n_4667 = ~n_4665 & ~n_4666;
assign n_4668 =  x_557 & ~n_4667;
assign n_4669 = ~x_557 &  n_4667;
assign n_4670 = ~n_4668 & ~n_4669;
assign n_4671 =  x_556 & ~n_1398;
assign n_4672 =  x_875 &  n_1401;
assign n_4673 = ~n_4671 & ~n_4672;
assign n_4674 =  x_556 & ~n_4673;
assign n_4675 = ~x_556 &  n_4673;
assign n_4676 = ~n_4674 & ~n_4675;
assign n_4677 =  x_555 & ~n_1398;
assign n_4678 =  x_874 &  n_1401;
assign n_4679 = ~n_4677 & ~n_4678;
assign n_4680 =  x_555 & ~n_4679;
assign n_4681 = ~x_555 &  n_4679;
assign n_4682 = ~n_4680 & ~n_4681;
assign n_4683 =  x_554 & ~n_1398;
assign n_4684 =  x_873 &  n_1401;
assign n_4685 = ~n_4683 & ~n_4684;
assign n_4686 =  x_554 & ~n_4685;
assign n_4687 = ~x_554 &  n_4685;
assign n_4688 = ~n_4686 & ~n_4687;
assign n_4689 =  x_553 & ~n_1398;
assign n_4690 =  x_872 &  n_1401;
assign n_4691 = ~n_4689 & ~n_4690;
assign n_4692 =  x_553 & ~n_4691;
assign n_4693 = ~x_553 &  n_4691;
assign n_4694 = ~n_4692 & ~n_4693;
assign n_4695 =  x_552 & ~n_1398;
assign n_4696 =  x_871 &  n_1401;
assign n_4697 = ~n_4695 & ~n_4696;
assign n_4698 =  x_552 & ~n_4697;
assign n_4699 = ~x_552 &  n_4697;
assign n_4700 = ~n_4698 & ~n_4699;
assign n_4701 =  x_551 & ~n_1681;
assign n_4702 =  i_32 &  n_1681;
assign n_4703 = ~n_4701 & ~n_4702;
assign n_4704 =  x_551 & ~n_4703;
assign n_4705 = ~x_551 &  n_4703;
assign n_4706 = ~n_4704 & ~n_4705;
assign n_4707 =  x_550 & ~n_1681;
assign n_4708 =  i_31 &  n_1681;
assign n_4709 = ~n_4707 & ~n_4708;
assign n_4710 =  x_550 & ~n_4709;
assign n_4711 = ~x_550 &  n_4709;
assign n_4712 = ~n_4710 & ~n_4711;
assign n_4713 =  x_549 & ~n_1681;
assign n_4714 =  i_30 &  n_1681;
assign n_4715 = ~n_4713 & ~n_4714;
assign n_4716 =  x_549 & ~n_4715;
assign n_4717 = ~x_549 &  n_4715;
assign n_4718 = ~n_4716 & ~n_4717;
assign n_4719 =  x_548 & ~n_1681;
assign n_4720 =  i_29 &  n_1681;
assign n_4721 = ~n_4719 & ~n_4720;
assign n_4722 =  x_548 & ~n_4721;
assign n_4723 = ~x_548 &  n_4721;
assign n_4724 = ~n_4722 & ~n_4723;
assign n_4725 =  x_547 & ~n_1681;
assign n_4726 =  i_28 &  n_1681;
assign n_4727 = ~n_4725 & ~n_4726;
assign n_4728 =  x_547 & ~n_4727;
assign n_4729 = ~x_547 &  n_4727;
assign n_4730 = ~n_4728 & ~n_4729;
assign n_4731 =  x_546 & ~n_1681;
assign n_4732 =  i_27 &  n_1681;
assign n_4733 = ~n_4731 & ~n_4732;
assign n_4734 =  x_546 & ~n_4733;
assign n_4735 = ~x_546 &  n_4733;
assign n_4736 = ~n_4734 & ~n_4735;
assign n_4737 =  x_545 & ~n_1681;
assign n_4738 =  i_26 &  n_1681;
assign n_4739 = ~n_4737 & ~n_4738;
assign n_4740 =  x_545 & ~n_4739;
assign n_4741 = ~x_545 &  n_4739;
assign n_4742 = ~n_4740 & ~n_4741;
assign n_4743 =  x_544 & ~n_1681;
assign n_4744 =  i_25 &  n_1681;
assign n_4745 = ~n_4743 & ~n_4744;
assign n_4746 =  x_544 & ~n_4745;
assign n_4747 = ~x_544 &  n_4745;
assign n_4748 = ~n_4746 & ~n_4747;
assign n_4749 =  x_543 & ~n_1681;
assign n_4750 =  i_24 &  n_1681;
assign n_4751 = ~n_4749 & ~n_4750;
assign n_4752 =  x_543 & ~n_4751;
assign n_4753 = ~x_543 &  n_4751;
assign n_4754 = ~n_4752 & ~n_4753;
assign n_4755 =  x_542 & ~n_1681;
assign n_4756 =  i_23 &  n_1681;
assign n_4757 = ~n_4755 & ~n_4756;
assign n_4758 =  x_542 & ~n_4757;
assign n_4759 = ~x_542 &  n_4757;
assign n_4760 = ~n_4758 & ~n_4759;
assign n_4761 =  x_541 & ~n_1681;
assign n_4762 =  i_22 &  n_1681;
assign n_4763 = ~n_4761 & ~n_4762;
assign n_4764 =  x_541 & ~n_4763;
assign n_4765 = ~x_541 &  n_4763;
assign n_4766 = ~n_4764 & ~n_4765;
assign n_4767 =  x_540 & ~n_1681;
assign n_4768 =  i_21 &  n_1681;
assign n_4769 = ~n_4767 & ~n_4768;
assign n_4770 =  x_540 & ~n_4769;
assign n_4771 = ~x_540 &  n_4769;
assign n_4772 = ~n_4770 & ~n_4771;
assign n_4773 =  x_539 & ~n_1681;
assign n_4774 =  i_20 &  n_1681;
assign n_4775 = ~n_4773 & ~n_4774;
assign n_4776 =  x_539 & ~n_4775;
assign n_4777 = ~x_539 &  n_4775;
assign n_4778 = ~n_4776 & ~n_4777;
assign n_4779 =  x_538 & ~n_1681;
assign n_4780 =  i_19 &  n_1681;
assign n_4781 = ~n_4779 & ~n_4780;
assign n_4782 =  x_538 & ~n_4781;
assign n_4783 = ~x_538 &  n_4781;
assign n_4784 = ~n_4782 & ~n_4783;
assign n_4785 =  x_537 & ~n_1681;
assign n_4786 =  i_18 &  n_1681;
assign n_4787 = ~n_4785 & ~n_4786;
assign n_4788 =  x_537 & ~n_4787;
assign n_4789 = ~x_537 &  n_4787;
assign n_4790 = ~n_4788 & ~n_4789;
assign n_4791 =  x_536 & ~n_1681;
assign n_4792 =  i_17 &  n_1681;
assign n_4793 = ~n_4791 & ~n_4792;
assign n_4794 =  x_536 & ~n_4793;
assign n_4795 = ~x_536 &  n_4793;
assign n_4796 = ~n_4794 & ~n_4795;
assign n_4797 =  x_535 & ~n_1681;
assign n_4798 =  i_16 &  n_1681;
assign n_4799 = ~n_4797 & ~n_4798;
assign n_4800 =  x_535 & ~n_4799;
assign n_4801 = ~x_535 &  n_4799;
assign n_4802 = ~n_4800 & ~n_4801;
assign n_4803 =  x_534 & ~n_1681;
assign n_4804 =  i_15 &  n_1681;
assign n_4805 = ~n_4803 & ~n_4804;
assign n_4806 =  x_534 & ~n_4805;
assign n_4807 = ~x_534 &  n_4805;
assign n_4808 = ~n_4806 & ~n_4807;
assign n_4809 =  x_533 & ~n_1681;
assign n_4810 =  i_14 &  n_1681;
assign n_4811 = ~n_4809 & ~n_4810;
assign n_4812 =  x_533 & ~n_4811;
assign n_4813 = ~x_533 &  n_4811;
assign n_4814 = ~n_4812 & ~n_4813;
assign n_4815 =  x_532 & ~n_1681;
assign n_4816 =  i_13 &  n_1681;
assign n_4817 = ~n_4815 & ~n_4816;
assign n_4818 =  x_532 & ~n_4817;
assign n_4819 = ~x_532 &  n_4817;
assign n_4820 = ~n_4818 & ~n_4819;
assign n_4821 =  x_531 & ~n_1681;
assign n_4822 =  i_12 &  n_1681;
assign n_4823 = ~n_4821 & ~n_4822;
assign n_4824 =  x_531 & ~n_4823;
assign n_4825 = ~x_531 &  n_4823;
assign n_4826 = ~n_4824 & ~n_4825;
assign n_4827 =  x_530 & ~n_1681;
assign n_4828 =  i_11 &  n_1681;
assign n_4829 = ~n_4827 & ~n_4828;
assign n_4830 =  x_530 & ~n_4829;
assign n_4831 = ~x_530 &  n_4829;
assign n_4832 = ~n_4830 & ~n_4831;
assign n_4833 =  x_529 & ~n_1681;
assign n_4834 =  i_10 &  n_1681;
assign n_4835 = ~n_4833 & ~n_4834;
assign n_4836 =  x_529 & ~n_4835;
assign n_4837 = ~x_529 &  n_4835;
assign n_4838 = ~n_4836 & ~n_4837;
assign n_4839 =  x_528 & ~n_1681;
assign n_4840 =  i_9 &  n_1681;
assign n_4841 = ~n_4839 & ~n_4840;
assign n_4842 =  x_528 & ~n_4841;
assign n_4843 = ~x_528 &  n_4841;
assign n_4844 = ~n_4842 & ~n_4843;
assign n_4845 =  x_527 & ~n_1681;
assign n_4846 =  i_8 &  n_1681;
assign n_4847 = ~n_4845 & ~n_4846;
assign n_4848 =  x_527 & ~n_4847;
assign n_4849 = ~x_527 &  n_4847;
assign n_4850 = ~n_4848 & ~n_4849;
assign n_4851 =  x_526 & ~n_1681;
assign n_4852 =  i_7 &  n_1681;
assign n_4853 = ~n_4851 & ~n_4852;
assign n_4854 =  x_526 & ~n_4853;
assign n_4855 = ~x_526 &  n_4853;
assign n_4856 = ~n_4854 & ~n_4855;
assign n_4857 =  x_525 & ~n_1681;
assign n_4858 =  i_6 &  n_1681;
assign n_4859 = ~n_4857 & ~n_4858;
assign n_4860 =  x_525 & ~n_4859;
assign n_4861 = ~x_525 &  n_4859;
assign n_4862 = ~n_4860 & ~n_4861;
assign n_4863 =  x_524 & ~n_1681;
assign n_4864 =  i_5 &  n_1681;
assign n_4865 = ~n_4863 & ~n_4864;
assign n_4866 =  x_524 & ~n_4865;
assign n_4867 = ~x_524 &  n_4865;
assign n_4868 = ~n_4866 & ~n_4867;
assign n_4869 =  x_523 & ~n_1681;
assign n_4870 =  i_4 &  n_1681;
assign n_4871 = ~n_4869 & ~n_4870;
assign n_4872 =  x_523 & ~n_4871;
assign n_4873 = ~x_523 &  n_4871;
assign n_4874 = ~n_4872 & ~n_4873;
assign n_4875 =  x_522 & ~n_1681;
assign n_4876 =  i_3 &  n_1681;
assign n_4877 = ~n_4875 & ~n_4876;
assign n_4878 =  x_522 & ~n_4877;
assign n_4879 = ~x_522 &  n_4877;
assign n_4880 = ~n_4878 & ~n_4879;
assign n_4881 =  x_521 & ~n_1681;
assign n_4882 =  i_2 &  n_1681;
assign n_4883 = ~n_4881 & ~n_4882;
assign n_4884 =  x_521 & ~n_4883;
assign n_4885 = ~x_521 &  n_4883;
assign n_4886 = ~n_4884 & ~n_4885;
assign n_4887 =  x_520 & ~n_1681;
assign n_4888 =  i_1 &  n_1681;
assign n_4889 = ~n_4887 & ~n_4888;
assign n_4890 =  x_520 & ~n_4889;
assign n_4891 = ~x_520 &  n_4889;
assign n_4892 = ~n_4890 & ~n_4891;
assign n_4893 = ~n_1397 & ~n_1722;
assign n_4894 =  i_32 & ~n_4893;
assign n_4895 =  x_519 &  n_4893;
assign n_4896 = ~n_4894 & ~n_4895;
assign n_4897 =  x_519 & ~n_4896;
assign n_4898 = ~x_519 &  n_4896;
assign n_4899 = ~n_4897 & ~n_4898;
assign n_4900 =  i_31 & ~n_4893;
assign n_4901 =  x_518 &  n_4893;
assign n_4902 = ~n_4900 & ~n_4901;
assign n_4903 =  x_518 & ~n_4902;
assign n_4904 = ~x_518 &  n_4902;
assign n_4905 = ~n_4903 & ~n_4904;
assign n_4906 =  i_30 & ~n_4893;
assign n_4907 =  x_517 &  n_4893;
assign n_4908 = ~n_4906 & ~n_4907;
assign n_4909 =  x_517 & ~n_4908;
assign n_4910 = ~x_517 &  n_4908;
assign n_4911 = ~n_4909 & ~n_4910;
assign n_4912 =  i_29 & ~n_4893;
assign n_4913 =  x_516 &  n_4893;
assign n_4914 = ~n_4912 & ~n_4913;
assign n_4915 =  x_516 & ~n_4914;
assign n_4916 = ~x_516 &  n_4914;
assign n_4917 = ~n_4915 & ~n_4916;
assign n_4918 =  i_28 & ~n_4893;
assign n_4919 =  x_515 &  n_4893;
assign n_4920 = ~n_4918 & ~n_4919;
assign n_4921 =  x_515 & ~n_4920;
assign n_4922 = ~x_515 &  n_4920;
assign n_4923 = ~n_4921 & ~n_4922;
assign n_4924 =  i_27 & ~n_4893;
assign n_4925 =  x_514 &  n_4893;
assign n_4926 = ~n_4924 & ~n_4925;
assign n_4927 =  x_514 & ~n_4926;
assign n_4928 = ~x_514 &  n_4926;
assign n_4929 = ~n_4927 & ~n_4928;
assign n_4930 =  i_26 & ~n_4893;
assign n_4931 =  x_513 &  n_4893;
assign n_4932 = ~n_4930 & ~n_4931;
assign n_4933 =  x_513 & ~n_4932;
assign n_4934 = ~x_513 &  n_4932;
assign n_4935 = ~n_4933 & ~n_4934;
assign n_4936 =  i_25 & ~n_4893;
assign n_4937 =  x_512 &  n_4893;
assign n_4938 = ~n_4936 & ~n_4937;
assign n_4939 =  x_512 & ~n_4938;
assign n_4940 = ~x_512 &  n_4938;
assign n_4941 = ~n_4939 & ~n_4940;
assign n_4942 =  i_24 & ~n_4893;
assign n_4943 =  x_511 &  n_4893;
assign n_4944 = ~n_4942 & ~n_4943;
assign n_4945 =  x_511 & ~n_4944;
assign n_4946 = ~x_511 &  n_4944;
assign n_4947 = ~n_4945 & ~n_4946;
assign n_4948 =  i_23 & ~n_4893;
assign n_4949 =  x_510 &  n_4893;
assign n_4950 = ~n_4948 & ~n_4949;
assign n_4951 =  x_510 & ~n_4950;
assign n_4952 = ~x_510 &  n_4950;
assign n_4953 = ~n_4951 & ~n_4952;
assign n_4954 =  i_22 & ~n_4893;
assign n_4955 =  x_509 &  n_4893;
assign n_4956 = ~n_4954 & ~n_4955;
assign n_4957 =  x_509 & ~n_4956;
assign n_4958 = ~x_509 &  n_4956;
assign n_4959 = ~n_4957 & ~n_4958;
assign n_4960 =  i_21 & ~n_4893;
assign n_4961 =  x_508 &  n_4893;
assign n_4962 = ~n_4960 & ~n_4961;
assign n_4963 =  x_508 & ~n_4962;
assign n_4964 = ~x_508 &  n_4962;
assign n_4965 = ~n_4963 & ~n_4964;
assign n_4966 =  i_20 & ~n_4893;
assign n_4967 =  x_507 &  n_4893;
assign n_4968 = ~n_4966 & ~n_4967;
assign n_4969 =  x_507 & ~n_4968;
assign n_4970 = ~x_507 &  n_4968;
assign n_4971 = ~n_4969 & ~n_4970;
assign n_4972 =  i_19 & ~n_4893;
assign n_4973 =  x_506 &  n_4893;
assign n_4974 = ~n_4972 & ~n_4973;
assign n_4975 =  x_506 & ~n_4974;
assign n_4976 = ~x_506 &  n_4974;
assign n_4977 = ~n_4975 & ~n_4976;
assign n_4978 =  i_18 & ~n_4893;
assign n_4979 =  x_505 &  n_4893;
assign n_4980 = ~n_4978 & ~n_4979;
assign n_4981 =  x_505 & ~n_4980;
assign n_4982 = ~x_505 &  n_4980;
assign n_4983 = ~n_4981 & ~n_4982;
assign n_4984 =  i_17 & ~n_4893;
assign n_4985 =  x_504 &  n_4893;
assign n_4986 = ~n_4984 & ~n_4985;
assign n_4987 =  x_504 & ~n_4986;
assign n_4988 = ~x_504 &  n_4986;
assign n_4989 = ~n_4987 & ~n_4988;
assign n_4990 =  i_16 & ~n_4893;
assign n_4991 =  x_503 &  n_4893;
assign n_4992 = ~n_4990 & ~n_4991;
assign n_4993 =  x_503 & ~n_4992;
assign n_4994 = ~x_503 &  n_4992;
assign n_4995 = ~n_4993 & ~n_4994;
assign n_4996 =  i_15 & ~n_4893;
assign n_4997 =  x_502 &  n_4893;
assign n_4998 = ~n_4996 & ~n_4997;
assign n_4999 =  x_502 & ~n_4998;
assign n_5000 = ~x_502 &  n_4998;
assign n_5001 = ~n_4999 & ~n_5000;
assign n_5002 =  i_14 & ~n_4893;
assign n_5003 =  x_501 &  n_4893;
assign n_5004 = ~n_5002 & ~n_5003;
assign n_5005 =  x_501 & ~n_5004;
assign n_5006 = ~x_501 &  n_5004;
assign n_5007 = ~n_5005 & ~n_5006;
assign n_5008 =  i_13 & ~n_4893;
assign n_5009 =  x_500 &  n_4893;
assign n_5010 = ~n_5008 & ~n_5009;
assign n_5011 =  x_500 & ~n_5010;
assign n_5012 = ~x_500 &  n_5010;
assign n_5013 = ~n_5011 & ~n_5012;
assign n_5014 =  i_12 & ~n_4893;
assign n_5015 =  x_499 &  n_4893;
assign n_5016 = ~n_5014 & ~n_5015;
assign n_5017 =  x_499 & ~n_5016;
assign n_5018 = ~x_499 &  n_5016;
assign n_5019 = ~n_5017 & ~n_5018;
assign n_5020 =  i_11 & ~n_4893;
assign n_5021 =  x_498 &  n_4893;
assign n_5022 = ~n_5020 & ~n_5021;
assign n_5023 =  x_498 & ~n_5022;
assign n_5024 = ~x_498 &  n_5022;
assign n_5025 = ~n_5023 & ~n_5024;
assign n_5026 =  i_10 & ~n_4893;
assign n_5027 =  x_497 &  n_4893;
assign n_5028 = ~n_5026 & ~n_5027;
assign n_5029 =  x_497 & ~n_5028;
assign n_5030 = ~x_497 &  n_5028;
assign n_5031 = ~n_5029 & ~n_5030;
assign n_5032 =  i_9 & ~n_4893;
assign n_5033 =  x_496 &  n_4893;
assign n_5034 = ~n_5032 & ~n_5033;
assign n_5035 =  x_496 & ~n_5034;
assign n_5036 = ~x_496 &  n_5034;
assign n_5037 = ~n_5035 & ~n_5036;
assign n_5038 =  i_8 & ~n_4893;
assign n_5039 =  x_495 &  n_4893;
assign n_5040 = ~n_5038 & ~n_5039;
assign n_5041 =  x_495 & ~n_5040;
assign n_5042 = ~x_495 &  n_5040;
assign n_5043 = ~n_5041 & ~n_5042;
assign n_5044 =  i_7 & ~n_4893;
assign n_5045 =  x_494 &  n_4893;
assign n_5046 = ~n_5044 & ~n_5045;
assign n_5047 =  x_494 & ~n_5046;
assign n_5048 = ~x_494 &  n_5046;
assign n_5049 = ~n_5047 & ~n_5048;
assign n_5050 =  i_6 & ~n_4893;
assign n_5051 =  x_493 &  n_4893;
assign n_5052 = ~n_5050 & ~n_5051;
assign n_5053 =  x_493 & ~n_5052;
assign n_5054 = ~x_493 &  n_5052;
assign n_5055 = ~n_5053 & ~n_5054;
assign n_5056 =  i_5 & ~n_4893;
assign n_5057 =  x_492 &  n_4893;
assign n_5058 = ~n_5056 & ~n_5057;
assign n_5059 =  x_492 & ~n_5058;
assign n_5060 = ~x_492 &  n_5058;
assign n_5061 = ~n_5059 & ~n_5060;
assign n_5062 =  i_4 & ~n_4893;
assign n_5063 =  x_491 &  n_4893;
assign n_5064 = ~n_5062 & ~n_5063;
assign n_5065 =  x_491 & ~n_5064;
assign n_5066 = ~x_491 &  n_5064;
assign n_5067 = ~n_5065 & ~n_5066;
assign n_5068 =  i_3 & ~n_4893;
assign n_5069 =  x_490 &  n_4893;
assign n_5070 = ~n_5068 & ~n_5069;
assign n_5071 =  x_490 & ~n_5070;
assign n_5072 = ~x_490 &  n_5070;
assign n_5073 = ~n_5071 & ~n_5072;
assign n_5074 =  i_2 & ~n_4893;
assign n_5075 =  x_489 &  n_4893;
assign n_5076 = ~n_5074 & ~n_5075;
assign n_5077 =  x_489 & ~n_5076;
assign n_5078 = ~x_489 &  n_5076;
assign n_5079 = ~n_5077 & ~n_5078;
assign n_5080 =  i_1 & ~n_4893;
assign n_5081 =  x_488 &  n_4893;
assign n_5082 = ~n_5080 & ~n_5081;
assign n_5083 =  x_488 & ~n_5082;
assign n_5084 = ~x_488 &  n_5082;
assign n_5085 = ~n_5083 & ~n_5084;
assign n_5086 =  x_456 & ~n_9;
assign n_5087 =  x_679 &  n_9;
assign n_5088 = ~n_5086 & ~n_5087;
assign n_5089 =  x_456 & ~n_5088;
assign n_5090 = ~x_456 &  n_5088;
assign n_5091 = ~n_5089 & ~n_5090;
assign n_5092 =  x_455 & ~n_9;
assign n_5093 =  x_678 &  n_9;
assign n_5094 = ~n_5092 & ~n_5093;
assign n_5095 =  x_455 & ~n_5094;
assign n_5096 = ~x_455 &  n_5094;
assign n_5097 = ~n_5095 & ~n_5096;
assign n_5098 =  x_454 & ~n_9;
assign n_5099 =  x_677 &  n_9;
assign n_5100 = ~n_5098 & ~n_5099;
assign n_5101 =  x_454 & ~n_5100;
assign n_5102 = ~x_454 &  n_5100;
assign n_5103 = ~n_5101 & ~n_5102;
assign n_5104 =  x_453 & ~n_9;
assign n_5105 =  x_676 &  n_9;
assign n_5106 = ~n_5104 & ~n_5105;
assign n_5107 =  x_453 & ~n_5106;
assign n_5108 = ~x_453 &  n_5106;
assign n_5109 = ~n_5107 & ~n_5108;
assign n_5110 =  x_452 & ~n_9;
assign n_5111 =  x_675 &  n_9;
assign n_5112 = ~n_5110 & ~n_5111;
assign n_5113 =  x_452 & ~n_5112;
assign n_5114 = ~x_452 &  n_5112;
assign n_5115 = ~n_5113 & ~n_5114;
assign n_5116 =  x_451 & ~n_9;
assign n_5117 =  x_674 &  n_9;
assign n_5118 = ~n_5116 & ~n_5117;
assign n_5119 =  x_451 & ~n_5118;
assign n_5120 = ~x_451 &  n_5118;
assign n_5121 = ~n_5119 & ~n_5120;
assign n_5122 =  x_450 & ~n_9;
assign n_5123 =  x_673 &  n_9;
assign n_5124 = ~n_5122 & ~n_5123;
assign n_5125 =  x_450 & ~n_5124;
assign n_5126 = ~x_450 &  n_5124;
assign n_5127 = ~n_5125 & ~n_5126;
assign n_5128 =  x_449 & ~n_9;
assign n_5129 =  x_672 &  n_9;
assign n_5130 = ~n_5128 & ~n_5129;
assign n_5131 =  x_449 & ~n_5130;
assign n_5132 = ~x_449 &  n_5130;
assign n_5133 = ~n_5131 & ~n_5132;
assign n_5134 =  x_448 & ~n_9;
assign n_5135 =  x_671 &  n_9;
assign n_5136 = ~n_5134 & ~n_5135;
assign n_5137 =  x_448 & ~n_5136;
assign n_5138 = ~x_448 &  n_5136;
assign n_5139 = ~n_5137 & ~n_5138;
assign n_5140 =  x_447 & ~n_9;
assign n_5141 =  x_670 &  n_9;
assign n_5142 = ~n_5140 & ~n_5141;
assign n_5143 =  x_447 & ~n_5142;
assign n_5144 = ~x_447 &  n_5142;
assign n_5145 = ~n_5143 & ~n_5144;
assign n_5146 =  x_446 & ~n_9;
assign n_5147 =  x_669 &  n_9;
assign n_5148 = ~n_5146 & ~n_5147;
assign n_5149 =  x_446 & ~n_5148;
assign n_5150 = ~x_446 &  n_5148;
assign n_5151 = ~n_5149 & ~n_5150;
assign n_5152 =  x_445 & ~n_9;
assign n_5153 =  x_668 &  n_9;
assign n_5154 = ~n_5152 & ~n_5153;
assign n_5155 =  x_445 & ~n_5154;
assign n_5156 = ~x_445 &  n_5154;
assign n_5157 = ~n_5155 & ~n_5156;
assign n_5158 =  x_444 & ~n_9;
assign n_5159 =  x_667 &  n_9;
assign n_5160 = ~n_5158 & ~n_5159;
assign n_5161 =  x_444 & ~n_5160;
assign n_5162 = ~x_444 &  n_5160;
assign n_5163 = ~n_5161 & ~n_5162;
assign n_5164 =  x_443 & ~n_9;
assign n_5165 =  x_666 &  n_9;
assign n_5166 = ~n_5164 & ~n_5165;
assign n_5167 =  x_443 & ~n_5166;
assign n_5168 = ~x_443 &  n_5166;
assign n_5169 = ~n_5167 & ~n_5168;
assign n_5170 =  x_442 & ~n_9;
assign n_5171 =  x_665 &  n_9;
assign n_5172 = ~n_5170 & ~n_5171;
assign n_5173 =  x_442 & ~n_5172;
assign n_5174 = ~x_442 &  n_5172;
assign n_5175 = ~n_5173 & ~n_5174;
assign n_5176 =  x_441 & ~n_9;
assign n_5177 =  x_664 &  n_9;
assign n_5178 = ~n_5176 & ~n_5177;
assign n_5179 =  x_441 & ~n_5178;
assign n_5180 = ~x_441 &  n_5178;
assign n_5181 = ~n_5179 & ~n_5180;
assign n_5182 =  x_440 & ~n_9;
assign n_5183 =  x_663 &  n_9;
assign n_5184 = ~n_5182 & ~n_5183;
assign n_5185 =  x_440 & ~n_5184;
assign n_5186 = ~x_440 &  n_5184;
assign n_5187 = ~n_5185 & ~n_5186;
assign n_5188 =  x_439 & ~n_9;
assign n_5189 =  x_662 &  n_9;
assign n_5190 = ~n_5188 & ~n_5189;
assign n_5191 =  x_439 & ~n_5190;
assign n_5192 = ~x_439 &  n_5190;
assign n_5193 = ~n_5191 & ~n_5192;
assign n_5194 =  x_438 & ~n_9;
assign n_5195 =  x_661 &  n_9;
assign n_5196 = ~n_5194 & ~n_5195;
assign n_5197 =  x_438 & ~n_5196;
assign n_5198 = ~x_438 &  n_5196;
assign n_5199 = ~n_5197 & ~n_5198;
assign n_5200 =  x_437 & ~n_9;
assign n_5201 =  x_660 &  n_9;
assign n_5202 = ~n_5200 & ~n_5201;
assign n_5203 =  x_437 & ~n_5202;
assign n_5204 = ~x_437 &  n_5202;
assign n_5205 = ~n_5203 & ~n_5204;
assign n_5206 =  x_436 & ~n_9;
assign n_5207 =  x_659 &  n_9;
assign n_5208 = ~n_5206 & ~n_5207;
assign n_5209 =  x_436 & ~n_5208;
assign n_5210 = ~x_436 &  n_5208;
assign n_5211 = ~n_5209 & ~n_5210;
assign n_5212 =  x_435 & ~n_9;
assign n_5213 =  x_658 &  n_9;
assign n_5214 = ~n_5212 & ~n_5213;
assign n_5215 =  x_435 & ~n_5214;
assign n_5216 = ~x_435 &  n_5214;
assign n_5217 = ~n_5215 & ~n_5216;
assign n_5218 =  x_434 & ~n_9;
assign n_5219 =  x_657 &  n_9;
assign n_5220 = ~n_5218 & ~n_5219;
assign n_5221 =  x_434 & ~n_5220;
assign n_5222 = ~x_434 &  n_5220;
assign n_5223 = ~n_5221 & ~n_5222;
assign n_5224 =  x_433 & ~n_9;
assign n_5225 =  x_656 &  n_9;
assign n_5226 = ~n_5224 & ~n_5225;
assign n_5227 =  x_433 & ~n_5226;
assign n_5228 = ~x_433 &  n_5226;
assign n_5229 = ~n_5227 & ~n_5228;
assign n_5230 =  x_432 & ~n_9;
assign n_5231 =  x_655 &  n_9;
assign n_5232 = ~n_5230 & ~n_5231;
assign n_5233 =  x_432 & ~n_5232;
assign n_5234 = ~x_432 &  n_5232;
assign n_5235 = ~n_5233 & ~n_5234;
assign n_5236 =  x_431 & ~n_9;
assign n_5237 =  x_654 &  n_9;
assign n_5238 = ~n_5236 & ~n_5237;
assign n_5239 =  x_431 & ~n_5238;
assign n_5240 = ~x_431 &  n_5238;
assign n_5241 = ~n_5239 & ~n_5240;
assign n_5242 =  x_430 & ~n_9;
assign n_5243 =  x_653 &  n_9;
assign n_5244 = ~n_5242 & ~n_5243;
assign n_5245 =  x_430 & ~n_5244;
assign n_5246 = ~x_430 &  n_5244;
assign n_5247 = ~n_5245 & ~n_5246;
assign n_5248 =  x_429 & ~n_9;
assign n_5249 =  x_652 &  n_9;
assign n_5250 = ~n_5248 & ~n_5249;
assign n_5251 =  x_429 & ~n_5250;
assign n_5252 = ~x_429 &  n_5250;
assign n_5253 = ~n_5251 & ~n_5252;
assign n_5254 =  x_428 & ~n_9;
assign n_5255 =  x_651 &  n_9;
assign n_5256 = ~n_5254 & ~n_5255;
assign n_5257 =  x_428 & ~n_5256;
assign n_5258 = ~x_428 &  n_5256;
assign n_5259 = ~n_5257 & ~n_5258;
assign n_5260 =  x_427 & ~n_9;
assign n_5261 =  x_650 &  n_9;
assign n_5262 = ~n_5260 & ~n_5261;
assign n_5263 =  x_427 & ~n_5262;
assign n_5264 = ~x_427 &  n_5262;
assign n_5265 = ~n_5263 & ~n_5264;
assign n_5266 =  x_426 & ~n_9;
assign n_5267 =  x_649 &  n_9;
assign n_5268 = ~n_5266 & ~n_5267;
assign n_5269 =  x_426 & ~n_5268;
assign n_5270 = ~x_426 &  n_5268;
assign n_5271 = ~n_5269 & ~n_5270;
assign n_5272 =  x_425 & ~n_9;
assign n_5273 =  x_648 &  n_9;
assign n_5274 = ~n_5272 & ~n_5273;
assign n_5275 =  x_425 & ~n_5274;
assign n_5276 = ~x_425 &  n_5274;
assign n_5277 = ~n_5275 & ~n_5276;
assign n_5278 =  x_424 & ~n_1537;
assign n_5279 =  x_838 &  n_1537;
assign n_5280 = ~n_5278 & ~n_5279;
assign n_5281 =  x_424 & ~n_5280;
assign n_5282 = ~x_424 &  n_5280;
assign n_5283 = ~n_5281 & ~n_5282;
assign n_5284 =  x_423 & ~n_1537;
assign n_5285 =  x_837 &  n_1537;
assign n_5286 = ~n_5284 & ~n_5285;
assign n_5287 =  x_423 & ~n_5286;
assign n_5288 = ~x_423 &  n_5286;
assign n_5289 = ~n_5287 & ~n_5288;
assign n_5290 =  x_422 & ~n_1537;
assign n_5291 =  x_836 &  n_1537;
assign n_5292 = ~n_5290 & ~n_5291;
assign n_5293 =  x_422 & ~n_5292;
assign n_5294 = ~x_422 &  n_5292;
assign n_5295 = ~n_5293 & ~n_5294;
assign n_5296 =  x_421 & ~n_1537;
assign n_5297 =  x_835 &  n_1537;
assign n_5298 = ~n_5296 & ~n_5297;
assign n_5299 =  x_421 & ~n_5298;
assign n_5300 = ~x_421 &  n_5298;
assign n_5301 = ~n_5299 & ~n_5300;
assign n_5302 =  x_420 & ~n_1537;
assign n_5303 =  x_834 &  n_1537;
assign n_5304 = ~n_5302 & ~n_5303;
assign n_5305 =  x_420 & ~n_5304;
assign n_5306 = ~x_420 &  n_5304;
assign n_5307 = ~n_5305 & ~n_5306;
assign n_5308 =  x_419 & ~n_1537;
assign n_5309 =  x_833 &  n_1537;
assign n_5310 = ~n_5308 & ~n_5309;
assign n_5311 =  x_419 & ~n_5310;
assign n_5312 = ~x_419 &  n_5310;
assign n_5313 = ~n_5311 & ~n_5312;
assign n_5314 =  x_418 & ~n_1537;
assign n_5315 =  x_832 &  n_1537;
assign n_5316 = ~n_5314 & ~n_5315;
assign n_5317 =  x_418 & ~n_5316;
assign n_5318 = ~x_418 &  n_5316;
assign n_5319 = ~n_5317 & ~n_5318;
assign n_5320 =  x_417 & ~n_1537;
assign n_5321 =  x_831 &  n_1537;
assign n_5322 = ~n_5320 & ~n_5321;
assign n_5323 =  x_417 & ~n_5322;
assign n_5324 = ~x_417 &  n_5322;
assign n_5325 = ~n_5323 & ~n_5324;
assign n_5326 =  x_416 & ~n_1537;
assign n_5327 =  x_830 &  n_1537;
assign n_5328 = ~n_5326 & ~n_5327;
assign n_5329 =  x_416 & ~n_5328;
assign n_5330 = ~x_416 &  n_5328;
assign n_5331 = ~n_5329 & ~n_5330;
assign n_5332 =  x_415 & ~n_1537;
assign n_5333 =  x_829 &  n_1537;
assign n_5334 = ~n_5332 & ~n_5333;
assign n_5335 =  x_415 & ~n_5334;
assign n_5336 = ~x_415 &  n_5334;
assign n_5337 = ~n_5335 & ~n_5336;
assign n_5338 =  x_414 & ~n_1537;
assign n_5339 =  x_828 &  n_1537;
assign n_5340 = ~n_5338 & ~n_5339;
assign n_5341 =  x_414 & ~n_5340;
assign n_5342 = ~x_414 &  n_5340;
assign n_5343 = ~n_5341 & ~n_5342;
assign n_5344 =  x_413 & ~n_1537;
assign n_5345 =  x_827 &  n_1537;
assign n_5346 = ~n_5344 & ~n_5345;
assign n_5347 =  x_413 & ~n_5346;
assign n_5348 = ~x_413 &  n_5346;
assign n_5349 = ~n_5347 & ~n_5348;
assign n_5350 =  x_412 & ~n_1537;
assign n_5351 =  x_826 &  n_1537;
assign n_5352 = ~n_5350 & ~n_5351;
assign n_5353 =  x_412 & ~n_5352;
assign n_5354 = ~x_412 &  n_5352;
assign n_5355 = ~n_5353 & ~n_5354;
assign n_5356 =  x_411 & ~n_1537;
assign n_5357 =  x_825 &  n_1537;
assign n_5358 = ~n_5356 & ~n_5357;
assign n_5359 =  x_411 & ~n_5358;
assign n_5360 = ~x_411 &  n_5358;
assign n_5361 = ~n_5359 & ~n_5360;
assign n_5362 =  x_410 & ~n_1537;
assign n_5363 =  x_824 &  n_1537;
assign n_5364 = ~n_5362 & ~n_5363;
assign n_5365 =  x_410 & ~n_5364;
assign n_5366 = ~x_410 &  n_5364;
assign n_5367 = ~n_5365 & ~n_5366;
assign n_5368 =  x_409 & ~n_1537;
assign n_5369 =  x_823 &  n_1537;
assign n_5370 = ~n_5368 & ~n_5369;
assign n_5371 =  x_409 & ~n_5370;
assign n_5372 = ~x_409 &  n_5370;
assign n_5373 = ~n_5371 & ~n_5372;
assign n_5374 =  x_408 & ~n_1537;
assign n_5375 =  x_822 &  n_1537;
assign n_5376 = ~n_5374 & ~n_5375;
assign n_5377 =  x_408 & ~n_5376;
assign n_5378 = ~x_408 &  n_5376;
assign n_5379 = ~n_5377 & ~n_5378;
assign n_5380 =  x_407 & ~n_1537;
assign n_5381 =  x_821 &  n_1537;
assign n_5382 = ~n_5380 & ~n_5381;
assign n_5383 =  x_407 & ~n_5382;
assign n_5384 = ~x_407 &  n_5382;
assign n_5385 = ~n_5383 & ~n_5384;
assign n_5386 =  x_406 & ~n_1537;
assign n_5387 =  x_820 &  n_1537;
assign n_5388 = ~n_5386 & ~n_5387;
assign n_5389 =  x_406 & ~n_5388;
assign n_5390 = ~x_406 &  n_5388;
assign n_5391 = ~n_5389 & ~n_5390;
assign n_5392 =  x_405 & ~n_1537;
assign n_5393 =  x_819 &  n_1537;
assign n_5394 = ~n_5392 & ~n_5393;
assign n_5395 =  x_405 & ~n_5394;
assign n_5396 = ~x_405 &  n_5394;
assign n_5397 = ~n_5395 & ~n_5396;
assign n_5398 =  x_404 & ~n_1537;
assign n_5399 =  x_818 &  n_1537;
assign n_5400 = ~n_5398 & ~n_5399;
assign n_5401 =  x_404 & ~n_5400;
assign n_5402 = ~x_404 &  n_5400;
assign n_5403 = ~n_5401 & ~n_5402;
assign n_5404 =  x_403 & ~n_1537;
assign n_5405 =  x_817 &  n_1537;
assign n_5406 = ~n_5404 & ~n_5405;
assign n_5407 =  x_403 & ~n_5406;
assign n_5408 = ~x_403 &  n_5406;
assign n_5409 = ~n_5407 & ~n_5408;
assign n_5410 =  x_402 & ~n_1537;
assign n_5411 =  x_816 &  n_1537;
assign n_5412 = ~n_5410 & ~n_5411;
assign n_5413 =  x_402 & ~n_5412;
assign n_5414 = ~x_402 &  n_5412;
assign n_5415 = ~n_5413 & ~n_5414;
assign n_5416 =  x_401 & ~n_1537;
assign n_5417 =  x_815 &  n_1537;
assign n_5418 = ~n_5416 & ~n_5417;
assign n_5419 =  x_401 & ~n_5418;
assign n_5420 = ~x_401 &  n_5418;
assign n_5421 = ~n_5419 & ~n_5420;
assign n_5422 =  x_400 & ~n_1537;
assign n_5423 =  x_814 &  n_1537;
assign n_5424 = ~n_5422 & ~n_5423;
assign n_5425 =  x_400 & ~n_5424;
assign n_5426 = ~x_400 &  n_5424;
assign n_5427 = ~n_5425 & ~n_5426;
assign n_5428 =  x_399 & ~n_1537;
assign n_5429 =  x_813 &  n_1537;
assign n_5430 = ~n_5428 & ~n_5429;
assign n_5431 =  x_399 & ~n_5430;
assign n_5432 = ~x_399 &  n_5430;
assign n_5433 = ~n_5431 & ~n_5432;
assign n_5434 =  x_398 & ~n_1537;
assign n_5435 =  x_812 &  n_1537;
assign n_5436 = ~n_5434 & ~n_5435;
assign n_5437 =  x_398 & ~n_5436;
assign n_5438 = ~x_398 &  n_5436;
assign n_5439 = ~n_5437 & ~n_5438;
assign n_5440 =  x_397 & ~n_1537;
assign n_5441 =  x_811 &  n_1537;
assign n_5442 = ~n_5440 & ~n_5441;
assign n_5443 =  x_397 & ~n_5442;
assign n_5444 = ~x_397 &  n_5442;
assign n_5445 = ~n_5443 & ~n_5444;
assign n_5446 =  x_396 & ~n_1537;
assign n_5447 =  x_810 &  n_1537;
assign n_5448 = ~n_5446 & ~n_5447;
assign n_5449 =  x_396 & ~n_5448;
assign n_5450 = ~x_396 &  n_5448;
assign n_5451 = ~n_5449 & ~n_5450;
assign n_5452 =  x_395 & ~n_1537;
assign n_5453 =  x_809 &  n_1537;
assign n_5454 = ~n_5452 & ~n_5453;
assign n_5455 =  x_395 & ~n_5454;
assign n_5456 = ~x_395 &  n_5454;
assign n_5457 = ~n_5455 & ~n_5456;
assign n_5458 =  x_394 & ~n_1537;
assign n_5459 =  x_808 &  n_1537;
assign n_5460 = ~n_5458 & ~n_5459;
assign n_5461 =  x_394 & ~n_5460;
assign n_5462 = ~x_394 &  n_5460;
assign n_5463 = ~n_5461 & ~n_5462;
assign n_5464 =  x_393 & ~n_1537;
assign n_5465 =  x_393 &  n_5464;
assign n_5466 = ~x_393 & ~n_5464;
assign n_5467 = ~n_5465 & ~n_5466;
assign n_5468 =  n_990 &  n_1536;
assign n_5469 = ~n_3933 & ~n_5468;
assign n_5470 =  x_361 &  n_5469;
assign n_5471 =  x_870 &  n_5468;
assign n_5472 = ~n_2070 & ~n_5471;
assign n_5473 = ~n_5470 &  n_5472;
assign n_5474 =  x_361 & ~n_5473;
assign n_5475 = ~x_361 &  n_5473;
assign n_5476 = ~n_5474 & ~n_5475;
assign n_5477 =  x_869 &  n_5468;
assign n_5478 =  x_360 &  n_5469;
assign n_5479 = ~n_5477 & ~n_5478;
assign n_5480 =  x_360 & ~n_5479;
assign n_5481 = ~x_360 &  n_5479;
assign n_5482 = ~n_5480 & ~n_5481;
assign n_5483 =  x_868 &  n_5468;
assign n_5484 =  x_359 &  n_5469;
assign n_5485 = ~n_5483 & ~n_5484;
assign n_5486 =  x_359 & ~n_5485;
assign n_5487 = ~x_359 &  n_5485;
assign n_5488 = ~n_5486 & ~n_5487;
assign n_5489 =  x_867 &  n_5468;
assign n_5490 =  x_358 &  n_5469;
assign n_5491 = ~n_5489 & ~n_5490;
assign n_5492 =  x_358 & ~n_5491;
assign n_5493 = ~x_358 &  n_5491;
assign n_5494 = ~n_5492 & ~n_5493;
assign n_5495 =  x_866 &  n_5468;
assign n_5496 =  x_357 &  n_5469;
assign n_5497 = ~n_5495 & ~n_5496;
assign n_5498 =  x_357 & ~n_5497;
assign n_5499 = ~x_357 &  n_5497;
assign n_5500 = ~n_5498 & ~n_5499;
assign n_5501 =  x_865 &  n_5468;
assign n_5502 =  x_356 &  n_5469;
assign n_5503 = ~n_5501 & ~n_5502;
assign n_5504 =  x_356 & ~n_5503;
assign n_5505 = ~x_356 &  n_5503;
assign n_5506 = ~n_5504 & ~n_5505;
assign n_5507 =  x_864 &  n_5468;
assign n_5508 =  x_355 &  n_5469;
assign n_5509 = ~n_5507 & ~n_5508;
assign n_5510 =  x_355 & ~n_5509;
assign n_5511 = ~x_355 &  n_5509;
assign n_5512 = ~n_5510 & ~n_5511;
assign n_5513 =  x_863 &  n_5468;
assign n_5514 =  x_354 &  n_5469;
assign n_5515 = ~n_5513 & ~n_5514;
assign n_5516 =  x_354 & ~n_5515;
assign n_5517 = ~x_354 &  n_5515;
assign n_5518 = ~n_5516 & ~n_5517;
assign n_5519 =  x_862 &  n_5468;
assign n_5520 =  x_353 &  n_5469;
assign n_5521 = ~n_5519 & ~n_5520;
assign n_5522 =  x_353 & ~n_5521;
assign n_5523 = ~x_353 &  n_5521;
assign n_5524 = ~n_5522 & ~n_5523;
assign n_5525 =  x_861 &  n_5468;
assign n_5526 =  x_352 &  n_5469;
assign n_5527 = ~n_5525 & ~n_5526;
assign n_5528 =  x_352 & ~n_5527;
assign n_5529 = ~x_352 &  n_5527;
assign n_5530 = ~n_5528 & ~n_5529;
assign n_5531 =  x_351 &  n_5469;
assign n_5532 =  x_860 &  n_5468;
assign n_5533 = ~n_2070 & ~n_5532;
assign n_5534 = ~n_5531 &  n_5533;
assign n_5535 =  x_351 & ~n_5534;
assign n_5536 = ~x_351 &  n_5534;
assign n_5537 = ~n_5535 & ~n_5536;
assign n_5538 =  x_859 &  n_5468;
assign n_5539 =  x_350 &  n_5469;
assign n_5540 = ~n_5538 & ~n_5539;
assign n_5541 =  x_350 & ~n_5540;
assign n_5542 = ~x_350 &  n_5540;
assign n_5543 = ~n_5541 & ~n_5542;
assign n_5544 =  x_858 &  n_5468;
assign n_5545 =  x_349 &  n_5469;
assign n_5546 = ~n_5544 & ~n_5545;
assign n_5547 =  x_349 & ~n_5546;
assign n_5548 = ~x_349 &  n_5546;
assign n_5549 = ~n_5547 & ~n_5548;
assign n_5550 =  x_857 &  n_5468;
assign n_5551 =  x_348 &  n_5469;
assign n_5552 = ~n_5550 & ~n_5551;
assign n_5553 =  x_348 & ~n_5552;
assign n_5554 = ~x_348 &  n_5552;
assign n_5555 = ~n_5553 & ~n_5554;
assign n_5556 =  x_856 &  n_5468;
assign n_5557 =  x_347 &  n_5469;
assign n_5558 = ~n_5556 & ~n_5557;
assign n_5559 =  x_347 & ~n_5558;
assign n_5560 = ~x_347 &  n_5558;
assign n_5561 = ~n_5559 & ~n_5560;
assign n_5562 =  x_855 &  n_5468;
assign n_5563 =  x_346 &  n_5469;
assign n_5564 = ~n_5562 & ~n_5563;
assign n_5565 =  x_346 & ~n_5564;
assign n_5566 = ~x_346 &  n_5564;
assign n_5567 = ~n_5565 & ~n_5566;
assign n_5568 =  x_854 &  n_5468;
assign n_5569 =  x_345 &  n_5469;
assign n_5570 = ~n_5568 & ~n_5569;
assign n_5571 =  x_345 & ~n_5570;
assign n_5572 = ~x_345 &  n_5570;
assign n_5573 = ~n_5571 & ~n_5572;
assign n_5574 =  x_853 &  n_5468;
assign n_5575 =  x_344 &  n_5469;
assign n_5576 = ~n_5574 & ~n_5575;
assign n_5577 =  x_344 & ~n_5576;
assign n_5578 = ~x_344 &  n_5576;
assign n_5579 = ~n_5577 & ~n_5578;
assign n_5580 =  x_852 &  n_5468;
assign n_5581 =  x_343 &  n_5469;
assign n_5582 = ~n_5580 & ~n_5581;
assign n_5583 =  x_343 & ~n_5582;
assign n_5584 = ~x_343 &  n_5582;
assign n_5585 = ~n_5583 & ~n_5584;
assign n_5586 =  x_851 &  n_5468;
assign n_5587 =  x_342 &  n_5469;
assign n_5588 = ~n_5586 & ~n_5587;
assign n_5589 =  x_342 & ~n_5588;
assign n_5590 = ~x_342 &  n_5588;
assign n_5591 = ~n_5589 & ~n_5590;
assign n_5592 =  x_850 &  n_5468;
assign n_5593 =  x_341 &  n_5469;
assign n_5594 = ~n_5592 & ~n_5593;
assign n_5595 =  x_341 & ~n_5594;
assign n_5596 = ~x_341 &  n_5594;
assign n_5597 = ~n_5595 & ~n_5596;
assign n_5598 =  x_849 &  n_5468;
assign n_5599 =  x_340 &  n_5469;
assign n_5600 = ~n_5598 & ~n_5599;
assign n_5601 =  x_340 & ~n_5600;
assign n_5602 = ~x_340 &  n_5600;
assign n_5603 = ~n_5601 & ~n_5602;
assign n_5604 =  x_848 &  n_5468;
assign n_5605 =  x_339 &  n_5469;
assign n_5606 = ~n_5604 & ~n_5605;
assign n_5607 =  x_339 & ~n_5606;
assign n_5608 = ~x_339 &  n_5606;
assign n_5609 = ~n_5607 & ~n_5608;
assign n_5610 =  x_847 &  n_5468;
assign n_5611 =  x_338 &  n_5469;
assign n_5612 = ~n_5610 & ~n_5611;
assign n_5613 =  x_338 & ~n_5612;
assign n_5614 = ~x_338 &  n_5612;
assign n_5615 = ~n_5613 & ~n_5614;
assign n_5616 =  x_846 &  n_5468;
assign n_5617 =  x_337 &  n_5469;
assign n_5618 = ~n_5616 & ~n_5617;
assign n_5619 =  x_337 & ~n_5618;
assign n_5620 = ~x_337 &  n_5618;
assign n_5621 = ~n_5619 & ~n_5620;
assign n_5622 =  x_845 &  n_5468;
assign n_5623 =  x_336 &  n_5469;
assign n_5624 = ~n_5622 & ~n_5623;
assign n_5625 =  x_336 & ~n_5624;
assign n_5626 = ~x_336 &  n_5624;
assign n_5627 = ~n_5625 & ~n_5626;
assign n_5628 =  x_844 &  n_5468;
assign n_5629 =  x_335 &  n_5469;
assign n_5630 = ~n_5628 & ~n_5629;
assign n_5631 =  x_335 & ~n_5630;
assign n_5632 = ~x_335 &  n_5630;
assign n_5633 = ~n_5631 & ~n_5632;
assign n_5634 =  x_843 &  n_5468;
assign n_5635 =  x_334 &  n_5469;
assign n_5636 = ~n_5634 & ~n_5635;
assign n_5637 =  x_334 & ~n_5636;
assign n_5638 = ~x_334 &  n_5636;
assign n_5639 = ~n_5637 & ~n_5638;
assign n_5640 =  x_842 &  n_5468;
assign n_5641 =  x_333 &  n_5469;
assign n_5642 = ~n_5640 & ~n_5641;
assign n_5643 =  x_333 & ~n_5642;
assign n_5644 = ~x_333 &  n_5642;
assign n_5645 = ~n_5643 & ~n_5644;
assign n_5646 =  x_841 &  n_5468;
assign n_5647 =  x_332 &  n_5469;
assign n_5648 = ~n_5646 & ~n_5647;
assign n_5649 =  x_332 & ~n_5648;
assign n_5650 = ~x_332 &  n_5648;
assign n_5651 = ~n_5649 & ~n_5650;
assign n_5652 =  x_840 &  n_5468;
assign n_5653 =  x_331 &  n_5469;
assign n_5654 = ~n_5652 & ~n_5653;
assign n_5655 =  x_331 & ~n_5654;
assign n_5656 = ~x_331 &  n_5654;
assign n_5657 = ~n_5655 & ~n_5656;
assign n_5658 =  x_839 &  n_5468;
assign n_5659 =  x_330 &  n_5469;
assign n_5660 = ~n_5658 & ~n_5659;
assign n_5661 =  x_330 & ~n_5660;
assign n_5662 = ~x_330 &  n_5660;
assign n_5663 = ~n_5661 & ~n_5662;
assign n_5664 = ~n_1709 & ~n_1858;
assign n_5665 =  x_42 & ~n_5664;
assign n_5666 =  x_329 & ~n_5665;
assign n_5667 =  x_392 &  n_1859;
assign n_5668 =  x_966 &  n_1710;
assign n_5669 = ~n_5667 & ~n_5668;
assign n_5670 = ~n_5666 &  n_5669;
assign n_5671 =  x_329 & ~n_5670;
assign n_5672 = ~x_329 &  n_5670;
assign n_5673 = ~n_5671 & ~n_5672;
assign n_5674 =  x_328 & ~n_5665;
assign n_5675 =  x_391 &  n_1859;
assign n_5676 =  x_965 &  n_1710;
assign n_5677 = ~n_5675 & ~n_5676;
assign n_5678 = ~n_5674 &  n_5677;
assign n_5679 =  x_328 & ~n_5678;
assign n_5680 = ~x_328 &  n_5678;
assign n_5681 = ~n_5679 & ~n_5680;
assign n_5682 =  x_327 & ~n_5665;
assign n_5683 =  x_390 &  n_1859;
assign n_5684 =  x_964 &  n_1710;
assign n_5685 = ~n_5683 & ~n_5684;
assign n_5686 = ~n_5682 &  n_5685;
assign n_5687 =  x_327 & ~n_5686;
assign n_5688 = ~x_327 &  n_5686;
assign n_5689 = ~n_5687 & ~n_5688;
assign n_5690 =  x_326 & ~n_5665;
assign n_5691 =  x_389 &  n_1859;
assign n_5692 =  x_963 &  n_1710;
assign n_5693 = ~n_5691 & ~n_5692;
assign n_5694 = ~n_5690 &  n_5693;
assign n_5695 =  x_326 & ~n_5694;
assign n_5696 = ~x_326 &  n_5694;
assign n_5697 = ~n_5695 & ~n_5696;
assign n_5698 =  x_325 & ~n_5665;
assign n_5699 =  x_388 &  n_1859;
assign n_5700 =  x_962 &  n_1710;
assign n_5701 = ~n_5699 & ~n_5700;
assign n_5702 = ~n_5698 &  n_5701;
assign n_5703 =  x_325 & ~n_5702;
assign n_5704 = ~x_325 &  n_5702;
assign n_5705 = ~n_5703 & ~n_5704;
assign n_5706 =  x_324 & ~n_5665;
assign n_5707 =  x_387 &  n_1859;
assign n_5708 =  x_961 &  n_1710;
assign n_5709 = ~n_5707 & ~n_5708;
assign n_5710 = ~n_5706 &  n_5709;
assign n_5711 =  x_324 & ~n_5710;
assign n_5712 = ~x_324 &  n_5710;
assign n_5713 = ~n_5711 & ~n_5712;
assign n_5714 =  x_323 & ~n_5665;
assign n_5715 =  x_386 &  n_1859;
assign n_5716 =  x_960 &  n_1710;
assign n_5717 = ~n_5715 & ~n_5716;
assign n_5718 = ~n_5714 &  n_5717;
assign n_5719 =  x_323 & ~n_5718;
assign n_5720 = ~x_323 &  n_5718;
assign n_5721 = ~n_5719 & ~n_5720;
assign n_5722 =  x_322 & ~n_5665;
assign n_5723 =  x_385 &  n_1859;
assign n_5724 =  x_959 &  n_1710;
assign n_5725 = ~n_5723 & ~n_5724;
assign n_5726 = ~n_5722 &  n_5725;
assign n_5727 =  x_322 & ~n_5726;
assign n_5728 = ~x_322 &  n_5726;
assign n_5729 = ~n_5727 & ~n_5728;
assign n_5730 =  x_321 & ~n_5665;
assign n_5731 =  x_384 &  n_1859;
assign n_5732 =  x_958 &  n_1710;
assign n_5733 = ~n_5731 & ~n_5732;
assign n_5734 = ~n_5730 &  n_5733;
assign n_5735 =  x_321 & ~n_5734;
assign n_5736 = ~x_321 &  n_5734;
assign n_5737 = ~n_5735 & ~n_5736;
assign n_5738 =  x_320 & ~n_5665;
assign n_5739 =  x_383 &  n_1859;
assign n_5740 =  x_957 &  n_1710;
assign n_5741 = ~n_5739 & ~n_5740;
assign n_5742 = ~n_5738 &  n_5741;
assign n_5743 =  x_320 & ~n_5742;
assign n_5744 = ~x_320 &  n_5742;
assign n_5745 = ~n_5743 & ~n_5744;
assign n_5746 =  x_319 & ~n_5665;
assign n_5747 =  x_382 &  n_1859;
assign n_5748 =  x_956 &  n_1710;
assign n_5749 = ~n_5747 & ~n_5748;
assign n_5750 = ~n_5746 &  n_5749;
assign n_5751 =  x_319 & ~n_5750;
assign n_5752 = ~x_319 &  n_5750;
assign n_5753 = ~n_5751 & ~n_5752;
assign n_5754 =  x_318 & ~n_5665;
assign n_5755 =  x_381 &  n_1859;
assign n_5756 =  x_955 &  n_1710;
assign n_5757 = ~n_5755 & ~n_5756;
assign n_5758 = ~n_5754 &  n_5757;
assign n_5759 =  x_318 & ~n_5758;
assign n_5760 = ~x_318 &  n_5758;
assign n_5761 = ~n_5759 & ~n_5760;
assign n_5762 =  x_317 & ~n_5665;
assign n_5763 =  x_380 &  n_1859;
assign n_5764 =  x_954 &  n_1710;
assign n_5765 = ~n_5763 & ~n_5764;
assign n_5766 = ~n_5762 &  n_5765;
assign n_5767 =  x_317 & ~n_5766;
assign n_5768 = ~x_317 &  n_5766;
assign n_5769 = ~n_5767 & ~n_5768;
assign n_5770 =  x_316 & ~n_5665;
assign n_5771 =  x_379 &  n_1859;
assign n_5772 =  x_953 &  n_1710;
assign n_5773 = ~n_5771 & ~n_5772;
assign n_5774 = ~n_5770 &  n_5773;
assign n_5775 =  x_316 & ~n_5774;
assign n_5776 = ~x_316 &  n_5774;
assign n_5777 = ~n_5775 & ~n_5776;
assign n_5778 =  x_315 & ~n_5665;
assign n_5779 =  x_378 &  n_1859;
assign n_5780 =  x_952 &  n_1710;
assign n_5781 = ~n_5779 & ~n_5780;
assign n_5782 = ~n_5778 &  n_5781;
assign n_5783 =  x_315 & ~n_5782;
assign n_5784 = ~x_315 &  n_5782;
assign n_5785 = ~n_5783 & ~n_5784;
assign n_5786 =  x_314 & ~n_5665;
assign n_5787 =  x_377 &  n_1859;
assign n_5788 =  x_951 &  n_1710;
assign n_5789 = ~n_5787 & ~n_5788;
assign n_5790 = ~n_5786 &  n_5789;
assign n_5791 =  x_314 & ~n_5790;
assign n_5792 = ~x_314 &  n_5790;
assign n_5793 = ~n_5791 & ~n_5792;
assign n_5794 =  x_313 & ~n_5665;
assign n_5795 =  x_376 &  n_1859;
assign n_5796 =  x_950 &  n_1710;
assign n_5797 = ~n_5795 & ~n_5796;
assign n_5798 = ~n_5794 &  n_5797;
assign n_5799 =  x_313 & ~n_5798;
assign n_5800 = ~x_313 &  n_5798;
assign n_5801 = ~n_5799 & ~n_5800;
assign n_5802 =  x_312 & ~n_5665;
assign n_5803 =  x_375 &  n_1859;
assign n_5804 =  x_949 &  n_1710;
assign n_5805 = ~n_5803 & ~n_5804;
assign n_5806 = ~n_5802 &  n_5805;
assign n_5807 =  x_312 & ~n_5806;
assign n_5808 = ~x_312 &  n_5806;
assign n_5809 = ~n_5807 & ~n_5808;
assign n_5810 =  x_311 & ~n_5665;
assign n_5811 =  x_374 &  n_1859;
assign n_5812 =  x_948 &  n_1710;
assign n_5813 = ~n_5811 & ~n_5812;
assign n_5814 = ~n_5810 &  n_5813;
assign n_5815 =  x_311 & ~n_5814;
assign n_5816 = ~x_311 &  n_5814;
assign n_5817 = ~n_5815 & ~n_5816;
assign n_5818 =  x_310 & ~n_5665;
assign n_5819 =  x_373 &  n_1859;
assign n_5820 =  x_947 &  n_1710;
assign n_5821 = ~n_5819 & ~n_5820;
assign n_5822 = ~n_5818 &  n_5821;
assign n_5823 =  x_310 & ~n_5822;
assign n_5824 = ~x_310 &  n_5822;
assign n_5825 = ~n_5823 & ~n_5824;
assign n_5826 =  x_309 & ~n_5665;
assign n_5827 =  x_372 &  n_1859;
assign n_5828 =  x_946 &  n_1710;
assign n_5829 = ~n_5827 & ~n_5828;
assign n_5830 = ~n_5826 &  n_5829;
assign n_5831 =  x_309 & ~n_5830;
assign n_5832 = ~x_309 &  n_5830;
assign n_5833 = ~n_5831 & ~n_5832;
assign n_5834 =  x_308 & ~n_5665;
assign n_5835 =  x_371 &  n_1859;
assign n_5836 =  x_945 &  n_1710;
assign n_5837 = ~n_5835 & ~n_5836;
assign n_5838 = ~n_5834 &  n_5837;
assign n_5839 =  x_308 & ~n_5838;
assign n_5840 = ~x_308 &  n_5838;
assign n_5841 = ~n_5839 & ~n_5840;
assign n_5842 =  x_307 & ~n_5665;
assign n_5843 =  x_370 &  n_1859;
assign n_5844 =  x_944 &  n_1710;
assign n_5845 = ~n_5843 & ~n_5844;
assign n_5846 = ~n_5842 &  n_5845;
assign n_5847 =  x_307 & ~n_5846;
assign n_5848 = ~x_307 &  n_5846;
assign n_5849 = ~n_5847 & ~n_5848;
assign n_5850 =  x_306 & ~n_5665;
assign n_5851 =  x_369 &  n_1859;
assign n_5852 =  x_943 &  n_1710;
assign n_5853 = ~n_5851 & ~n_5852;
assign n_5854 = ~n_5850 &  n_5853;
assign n_5855 =  x_306 & ~n_5854;
assign n_5856 = ~x_306 &  n_5854;
assign n_5857 = ~n_5855 & ~n_5856;
assign n_5858 =  x_305 & ~n_5665;
assign n_5859 =  x_368 &  n_1859;
assign n_5860 =  x_942 &  n_1710;
assign n_5861 = ~n_5859 & ~n_5860;
assign n_5862 = ~n_5858 &  n_5861;
assign n_5863 =  x_305 & ~n_5862;
assign n_5864 = ~x_305 &  n_5862;
assign n_5865 = ~n_5863 & ~n_5864;
assign n_5866 =  x_304 & ~n_5665;
assign n_5867 =  x_367 &  n_1859;
assign n_5868 =  x_941 &  n_1710;
assign n_5869 = ~n_5867 & ~n_5868;
assign n_5870 = ~n_5866 &  n_5869;
assign n_5871 =  x_304 & ~n_5870;
assign n_5872 = ~x_304 &  n_5870;
assign n_5873 = ~n_5871 & ~n_5872;
assign n_5874 =  x_303 & ~n_5665;
assign n_5875 =  x_366 &  n_1859;
assign n_5876 =  x_940 &  n_1710;
assign n_5877 = ~n_5875 & ~n_5876;
assign n_5878 = ~n_5874 &  n_5877;
assign n_5879 =  x_303 & ~n_5878;
assign n_5880 = ~x_303 &  n_5878;
assign n_5881 = ~n_5879 & ~n_5880;
assign n_5882 =  x_302 & ~n_5665;
assign n_5883 =  x_365 &  n_1859;
assign n_5884 =  x_939 &  n_1710;
assign n_5885 = ~n_5883 & ~n_5884;
assign n_5886 = ~n_5882 &  n_5885;
assign n_5887 =  x_302 & ~n_5886;
assign n_5888 = ~x_302 &  n_5886;
assign n_5889 = ~n_5887 & ~n_5888;
assign n_5890 =  x_301 & ~n_5665;
assign n_5891 =  x_364 &  n_1859;
assign n_5892 =  x_938 &  n_1710;
assign n_5893 = ~n_5891 & ~n_5892;
assign n_5894 = ~n_5890 &  n_5893;
assign n_5895 =  x_301 & ~n_5894;
assign n_5896 = ~x_301 &  n_5894;
assign n_5897 = ~n_5895 & ~n_5896;
assign n_5898 =  x_300 & ~n_5665;
assign n_5899 =  x_363 &  n_1859;
assign n_5900 =  x_937 &  n_1710;
assign n_5901 = ~n_5899 & ~n_5900;
assign n_5902 = ~n_5898 &  n_5901;
assign n_5903 =  x_300 & ~n_5902;
assign n_5904 = ~x_300 &  n_5902;
assign n_5905 = ~n_5903 & ~n_5904;
assign n_5906 =  x_299 & ~n_5665;
assign n_5907 =  x_362 &  n_1859;
assign n_5908 =  x_936 &  n_1710;
assign n_5909 = ~n_5907 & ~n_5908;
assign n_5910 = ~n_5906 &  n_5909;
assign n_5911 =  x_299 & ~n_5910;
assign n_5912 = ~x_299 &  n_5910;
assign n_5913 = ~n_5911 & ~n_5912;
assign n_5914 =  x_935 &  n_1710;
assign n_5915 =  x_298 & ~n_5665;
assign n_5916 = ~n_5914 & ~n_5915;
assign n_5917 =  x_298 & ~n_5916;
assign n_5918 = ~x_298 &  n_5916;
assign n_5919 = ~n_5917 & ~n_5918;
assign n_5920 = ~n_2337 & ~n_3933;
assign n_5921 =  x_266 &  n_5920;
assign n_5922 =  x_870 &  n_2337;
assign n_5923 = ~n_2070 & ~n_5922;
assign n_5924 = ~n_5921 &  n_5923;
assign n_5925 =  x_266 & ~n_5924;
assign n_5926 = ~x_266 &  n_5924;
assign n_5927 = ~n_5925 & ~n_5926;
assign n_5928 =  x_265 &  n_5920;
assign n_5929 =  x_869 &  n_2337;
assign n_5930 = ~n_2070 & ~n_5929;
assign n_5931 = ~n_5928 &  n_5930;
assign n_5932 =  x_265 & ~n_5931;
assign n_5933 = ~x_265 &  n_5931;
assign n_5934 = ~n_5932 & ~n_5933;
assign n_5935 =  x_868 &  n_2337;
assign n_5936 =  x_264 &  n_5920;
assign n_5937 = ~n_5935 & ~n_5936;
assign n_5938 =  x_264 & ~n_5937;
assign n_5939 = ~x_264 &  n_5937;
assign n_5940 = ~n_5938 & ~n_5939;
assign n_5941 =  x_263 &  n_5920;
assign n_5942 =  x_867 &  n_2337;
assign n_5943 = ~n_2070 & ~n_5942;
assign n_5944 = ~n_5941 &  n_5943;
assign n_5945 =  x_263 & ~n_5944;
assign n_5946 = ~x_263 &  n_5944;
assign n_5947 = ~n_5945 & ~n_5946;
assign n_5948 =  x_866 &  n_2337;
assign n_5949 =  x_262 &  n_5920;
assign n_5950 = ~n_5948 & ~n_5949;
assign n_5951 =  x_262 & ~n_5950;
assign n_5952 = ~x_262 &  n_5950;
assign n_5953 = ~n_5951 & ~n_5952;
assign n_5954 =  x_865 &  n_2337;
assign n_5955 =  x_261 &  n_5920;
assign n_5956 = ~n_5954 & ~n_5955;
assign n_5957 =  x_261 & ~n_5956;
assign n_5958 = ~x_261 &  n_5956;
assign n_5959 = ~n_5957 & ~n_5958;
assign n_5960 =  x_864 &  n_2337;
assign n_5961 =  x_260 &  n_5920;
assign n_5962 = ~n_5960 & ~n_5961;
assign n_5963 =  x_260 & ~n_5962;
assign n_5964 = ~x_260 &  n_5962;
assign n_5965 = ~n_5963 & ~n_5964;
assign n_5966 =  x_863 &  n_2337;
assign n_5967 =  x_259 &  n_5920;
assign n_5968 = ~n_5966 & ~n_5967;
assign n_5969 =  x_259 & ~n_5968;
assign n_5970 = ~x_259 &  n_5968;
assign n_5971 = ~n_5969 & ~n_5970;
assign n_5972 =  x_862 &  n_2337;
assign n_5973 =  x_258 &  n_5920;
assign n_5974 = ~n_5972 & ~n_5973;
assign n_5975 =  x_258 & ~n_5974;
assign n_5976 = ~x_258 &  n_5974;
assign n_5977 = ~n_5975 & ~n_5976;
assign n_5978 =  x_861 &  n_2337;
assign n_5979 =  x_257 &  n_5920;
assign n_5980 = ~n_5978 & ~n_5979;
assign n_5981 =  x_257 & ~n_5980;
assign n_5982 = ~x_257 &  n_5980;
assign n_5983 = ~n_5981 & ~n_5982;
assign n_5984 =  x_256 &  n_5920;
assign n_5985 =  x_860 &  n_2337;
assign n_5986 = ~n_2070 & ~n_5985;
assign n_5987 = ~n_5984 &  n_5986;
assign n_5988 =  x_256 & ~n_5987;
assign n_5989 = ~x_256 &  n_5987;
assign n_5990 = ~n_5988 & ~n_5989;
assign n_5991 =  x_859 &  n_2337;
assign n_5992 =  x_255 &  n_5920;
assign n_5993 = ~n_5991 & ~n_5992;
assign n_5994 =  x_255 & ~n_5993;
assign n_5995 = ~x_255 &  n_5993;
assign n_5996 = ~n_5994 & ~n_5995;
assign n_5997 =  x_858 &  n_2337;
assign n_5998 =  x_254 &  n_5920;
assign n_5999 = ~n_5997 & ~n_5998;
assign n_6000 =  x_254 & ~n_5999;
assign n_6001 = ~x_254 &  n_5999;
assign n_6002 = ~n_6000 & ~n_6001;
assign n_6003 =  x_857 &  n_2337;
assign n_6004 =  x_253 &  n_5920;
assign n_6005 = ~n_6003 & ~n_6004;
assign n_6006 =  x_253 & ~n_6005;
assign n_6007 = ~x_253 &  n_6005;
assign n_6008 = ~n_6006 & ~n_6007;
assign n_6009 =  x_856 &  n_2337;
assign n_6010 =  x_252 &  n_5920;
assign n_6011 = ~n_6009 & ~n_6010;
assign n_6012 =  x_252 & ~n_6011;
assign n_6013 = ~x_252 &  n_6011;
assign n_6014 = ~n_6012 & ~n_6013;
assign n_6015 =  x_855 &  n_2337;
assign n_6016 =  x_251 &  n_5920;
assign n_6017 = ~n_6015 & ~n_6016;
assign n_6018 =  x_251 & ~n_6017;
assign n_6019 = ~x_251 &  n_6017;
assign n_6020 = ~n_6018 & ~n_6019;
assign n_6021 =  x_854 &  n_2337;
assign n_6022 =  x_250 &  n_5920;
assign n_6023 = ~n_6021 & ~n_6022;
assign n_6024 =  x_250 & ~n_6023;
assign n_6025 = ~x_250 &  n_6023;
assign n_6026 = ~n_6024 & ~n_6025;
assign n_6027 =  x_853 &  n_2337;
assign n_6028 =  x_249 &  n_5920;
assign n_6029 = ~n_6027 & ~n_6028;
assign n_6030 =  x_249 & ~n_6029;
assign n_6031 = ~x_249 &  n_6029;
assign n_6032 = ~n_6030 & ~n_6031;
assign n_6033 =  x_852 &  n_2337;
assign n_6034 =  x_248 &  n_5920;
assign n_6035 = ~n_6033 & ~n_6034;
assign n_6036 =  x_248 & ~n_6035;
assign n_6037 = ~x_248 &  n_6035;
assign n_6038 = ~n_6036 & ~n_6037;
assign n_6039 =  x_851 &  n_2337;
assign n_6040 =  x_247 &  n_5920;
assign n_6041 = ~n_6039 & ~n_6040;
assign n_6042 =  x_247 & ~n_6041;
assign n_6043 = ~x_247 &  n_6041;
assign n_6044 = ~n_6042 & ~n_6043;
assign n_6045 =  x_850 &  n_2337;
assign n_6046 =  x_246 &  n_5920;
assign n_6047 = ~n_6045 & ~n_6046;
assign n_6048 =  x_246 & ~n_6047;
assign n_6049 = ~x_246 &  n_6047;
assign n_6050 = ~n_6048 & ~n_6049;
assign n_6051 =  x_849 &  n_2337;
assign n_6052 =  x_245 &  n_5920;
assign n_6053 = ~n_6051 & ~n_6052;
assign n_6054 =  x_245 & ~n_6053;
assign n_6055 = ~x_245 &  n_6053;
assign n_6056 = ~n_6054 & ~n_6055;
assign n_6057 =  x_848 &  n_2337;
assign n_6058 =  x_244 &  n_5920;
assign n_6059 = ~n_6057 & ~n_6058;
assign n_6060 =  x_244 & ~n_6059;
assign n_6061 = ~x_244 &  n_6059;
assign n_6062 = ~n_6060 & ~n_6061;
assign n_6063 =  x_847 &  n_2337;
assign n_6064 =  x_243 &  n_5920;
assign n_6065 = ~n_6063 & ~n_6064;
assign n_6066 =  x_243 & ~n_6065;
assign n_6067 = ~x_243 &  n_6065;
assign n_6068 = ~n_6066 & ~n_6067;
assign n_6069 =  x_846 &  n_2337;
assign n_6070 =  x_242 &  n_5920;
assign n_6071 = ~n_6069 & ~n_6070;
assign n_6072 =  x_242 & ~n_6071;
assign n_6073 = ~x_242 &  n_6071;
assign n_6074 = ~n_6072 & ~n_6073;
assign n_6075 =  x_845 &  n_2337;
assign n_6076 =  x_241 &  n_5920;
assign n_6077 = ~n_6075 & ~n_6076;
assign n_6078 =  x_241 & ~n_6077;
assign n_6079 = ~x_241 &  n_6077;
assign n_6080 = ~n_6078 & ~n_6079;
assign n_6081 =  x_844 &  n_2337;
assign n_6082 =  x_240 &  n_5920;
assign n_6083 = ~n_6081 & ~n_6082;
assign n_6084 =  x_240 & ~n_6083;
assign n_6085 = ~x_240 &  n_6083;
assign n_6086 = ~n_6084 & ~n_6085;
assign n_6087 =  x_843 &  n_2337;
assign n_6088 =  x_239 &  n_5920;
assign n_6089 = ~n_6087 & ~n_6088;
assign n_6090 =  x_239 & ~n_6089;
assign n_6091 = ~x_239 &  n_6089;
assign n_6092 = ~n_6090 & ~n_6091;
assign n_6093 =  x_842 &  n_2337;
assign n_6094 =  x_238 &  n_5920;
assign n_6095 = ~n_6093 & ~n_6094;
assign n_6096 =  x_238 & ~n_6095;
assign n_6097 = ~x_238 &  n_6095;
assign n_6098 = ~n_6096 & ~n_6097;
assign n_6099 =  x_841 &  n_2337;
assign n_6100 =  x_237 &  n_5920;
assign n_6101 = ~n_6099 & ~n_6100;
assign n_6102 =  x_237 & ~n_6101;
assign n_6103 = ~x_237 &  n_6101;
assign n_6104 = ~n_6102 & ~n_6103;
assign n_6105 =  x_840 &  n_2337;
assign n_6106 =  x_236 &  n_5920;
assign n_6107 = ~n_6105 & ~n_6106;
assign n_6108 =  x_236 & ~n_6107;
assign n_6109 = ~x_236 &  n_6107;
assign n_6110 = ~n_6108 & ~n_6109;
assign n_6111 =  x_839 &  n_2337;
assign n_6112 =  x_235 &  n_5920;
assign n_6113 = ~n_6111 & ~n_6112;
assign n_6114 =  x_235 & ~n_6113;
assign n_6115 = ~x_235 &  n_6113;
assign n_6116 = ~n_6114 & ~n_6115;
assign n_6117 =  x_234 & ~n_1802;
assign n_6118 =  i_32 &  n_1802;
assign n_6119 = ~n_6117 & ~n_6118;
assign n_6120 =  x_234 & ~n_6119;
assign n_6121 = ~x_234 &  n_6119;
assign n_6122 = ~n_6120 & ~n_6121;
assign n_6123 =  x_233 & ~n_1802;
assign n_6124 =  i_31 &  n_1802;
assign n_6125 = ~n_6123 & ~n_6124;
assign n_6126 =  x_233 & ~n_6125;
assign n_6127 = ~x_233 &  n_6125;
assign n_6128 = ~n_6126 & ~n_6127;
assign n_6129 =  x_232 & ~n_1802;
assign n_6130 =  i_30 &  n_1802;
assign n_6131 = ~n_6129 & ~n_6130;
assign n_6132 =  x_232 & ~n_6131;
assign n_6133 = ~x_232 &  n_6131;
assign n_6134 = ~n_6132 & ~n_6133;
assign n_6135 =  x_231 & ~n_1802;
assign n_6136 =  i_29 &  n_1802;
assign n_6137 = ~n_6135 & ~n_6136;
assign n_6138 =  x_231 & ~n_6137;
assign n_6139 = ~x_231 &  n_6137;
assign n_6140 = ~n_6138 & ~n_6139;
assign n_6141 =  x_230 & ~n_1802;
assign n_6142 =  i_28 &  n_1802;
assign n_6143 = ~n_6141 & ~n_6142;
assign n_6144 =  x_230 & ~n_6143;
assign n_6145 = ~x_230 &  n_6143;
assign n_6146 = ~n_6144 & ~n_6145;
assign n_6147 =  x_229 & ~n_1802;
assign n_6148 =  i_27 &  n_1802;
assign n_6149 = ~n_6147 & ~n_6148;
assign n_6150 =  x_229 & ~n_6149;
assign n_6151 = ~x_229 &  n_6149;
assign n_6152 = ~n_6150 & ~n_6151;
assign n_6153 =  x_228 & ~n_1802;
assign n_6154 =  i_26 &  n_1802;
assign n_6155 = ~n_6153 & ~n_6154;
assign n_6156 =  x_228 & ~n_6155;
assign n_6157 = ~x_228 &  n_6155;
assign n_6158 = ~n_6156 & ~n_6157;
assign n_6159 =  x_227 & ~n_1802;
assign n_6160 =  i_25 &  n_1802;
assign n_6161 = ~n_6159 & ~n_6160;
assign n_6162 =  x_227 & ~n_6161;
assign n_6163 = ~x_227 &  n_6161;
assign n_6164 = ~n_6162 & ~n_6163;
assign n_6165 =  x_226 & ~n_1802;
assign n_6166 =  i_24 &  n_1802;
assign n_6167 = ~n_6165 & ~n_6166;
assign n_6168 =  x_226 & ~n_6167;
assign n_6169 = ~x_226 &  n_6167;
assign n_6170 = ~n_6168 & ~n_6169;
assign n_6171 =  x_225 & ~n_1802;
assign n_6172 =  i_23 &  n_1802;
assign n_6173 = ~n_6171 & ~n_6172;
assign n_6174 =  x_225 & ~n_6173;
assign n_6175 = ~x_225 &  n_6173;
assign n_6176 = ~n_6174 & ~n_6175;
assign n_6177 =  x_224 & ~n_1802;
assign n_6178 =  i_22 &  n_1802;
assign n_6179 = ~n_6177 & ~n_6178;
assign n_6180 =  x_224 & ~n_6179;
assign n_6181 = ~x_224 &  n_6179;
assign n_6182 = ~n_6180 & ~n_6181;
assign n_6183 =  x_223 & ~n_1802;
assign n_6184 =  i_21 &  n_1802;
assign n_6185 = ~n_6183 & ~n_6184;
assign n_6186 =  x_223 & ~n_6185;
assign n_6187 = ~x_223 &  n_6185;
assign n_6188 = ~n_6186 & ~n_6187;
assign n_6189 =  x_222 & ~n_1802;
assign n_6190 =  i_20 &  n_1802;
assign n_6191 = ~n_6189 & ~n_6190;
assign n_6192 =  x_222 & ~n_6191;
assign n_6193 = ~x_222 &  n_6191;
assign n_6194 = ~n_6192 & ~n_6193;
assign n_6195 =  x_221 & ~n_1802;
assign n_6196 =  i_19 &  n_1802;
assign n_6197 = ~n_6195 & ~n_6196;
assign n_6198 =  x_221 & ~n_6197;
assign n_6199 = ~x_221 &  n_6197;
assign n_6200 = ~n_6198 & ~n_6199;
assign n_6201 =  x_220 & ~n_1802;
assign n_6202 =  i_18 &  n_1802;
assign n_6203 = ~n_6201 & ~n_6202;
assign n_6204 =  x_220 & ~n_6203;
assign n_6205 = ~x_220 &  n_6203;
assign n_6206 = ~n_6204 & ~n_6205;
assign n_6207 =  x_219 & ~n_1802;
assign n_6208 =  i_17 &  n_1802;
assign n_6209 = ~n_6207 & ~n_6208;
assign n_6210 =  x_219 & ~n_6209;
assign n_6211 = ~x_219 &  n_6209;
assign n_6212 = ~n_6210 & ~n_6211;
assign n_6213 =  x_218 & ~n_1802;
assign n_6214 =  i_16 &  n_1802;
assign n_6215 = ~n_6213 & ~n_6214;
assign n_6216 =  x_218 & ~n_6215;
assign n_6217 = ~x_218 &  n_6215;
assign n_6218 = ~n_6216 & ~n_6217;
assign n_6219 =  x_217 & ~n_1802;
assign n_6220 =  i_15 &  n_1802;
assign n_6221 = ~n_6219 & ~n_6220;
assign n_6222 =  x_217 & ~n_6221;
assign n_6223 = ~x_217 &  n_6221;
assign n_6224 = ~n_6222 & ~n_6223;
assign n_6225 =  x_216 & ~n_1802;
assign n_6226 =  i_14 &  n_1802;
assign n_6227 = ~n_6225 & ~n_6226;
assign n_6228 =  x_216 & ~n_6227;
assign n_6229 = ~x_216 &  n_6227;
assign n_6230 = ~n_6228 & ~n_6229;
assign n_6231 =  x_215 & ~n_1802;
assign n_6232 =  i_13 &  n_1802;
assign n_6233 = ~n_6231 & ~n_6232;
assign n_6234 =  x_215 & ~n_6233;
assign n_6235 = ~x_215 &  n_6233;
assign n_6236 = ~n_6234 & ~n_6235;
assign n_6237 =  x_214 & ~n_1802;
assign n_6238 =  i_12 &  n_1802;
assign n_6239 = ~n_6237 & ~n_6238;
assign n_6240 =  x_214 & ~n_6239;
assign n_6241 = ~x_214 &  n_6239;
assign n_6242 = ~n_6240 & ~n_6241;
assign n_6243 =  x_213 & ~n_1802;
assign n_6244 =  i_11 &  n_1802;
assign n_6245 = ~n_6243 & ~n_6244;
assign n_6246 =  x_213 & ~n_6245;
assign n_6247 = ~x_213 &  n_6245;
assign n_6248 = ~n_6246 & ~n_6247;
assign n_6249 =  x_212 & ~n_1802;
assign n_6250 =  i_10 &  n_1802;
assign n_6251 = ~n_6249 & ~n_6250;
assign n_6252 =  x_212 & ~n_6251;
assign n_6253 = ~x_212 &  n_6251;
assign n_6254 = ~n_6252 & ~n_6253;
assign n_6255 =  x_211 & ~n_1802;
assign n_6256 =  i_9 &  n_1802;
assign n_6257 = ~n_6255 & ~n_6256;
assign n_6258 =  x_211 & ~n_6257;
assign n_6259 = ~x_211 &  n_6257;
assign n_6260 = ~n_6258 & ~n_6259;
assign n_6261 =  x_210 & ~n_1802;
assign n_6262 =  i_8 &  n_1802;
assign n_6263 = ~n_6261 & ~n_6262;
assign n_6264 =  x_210 & ~n_6263;
assign n_6265 = ~x_210 &  n_6263;
assign n_6266 = ~n_6264 & ~n_6265;
assign n_6267 =  x_209 & ~n_1802;
assign n_6268 =  i_7 &  n_1802;
assign n_6269 = ~n_6267 & ~n_6268;
assign n_6270 =  x_209 & ~n_6269;
assign n_6271 = ~x_209 &  n_6269;
assign n_6272 = ~n_6270 & ~n_6271;
assign n_6273 =  x_208 & ~n_1802;
assign n_6274 =  i_6 &  n_1802;
assign n_6275 = ~n_6273 & ~n_6274;
assign n_6276 =  x_208 & ~n_6275;
assign n_6277 = ~x_208 &  n_6275;
assign n_6278 = ~n_6276 & ~n_6277;
assign n_6279 =  x_207 & ~n_1802;
assign n_6280 =  i_5 &  n_1802;
assign n_6281 = ~n_6279 & ~n_6280;
assign n_6282 =  x_207 & ~n_6281;
assign n_6283 = ~x_207 &  n_6281;
assign n_6284 = ~n_6282 & ~n_6283;
assign n_6285 =  x_206 & ~n_1802;
assign n_6286 =  i_4 &  n_1802;
assign n_6287 = ~n_6285 & ~n_6286;
assign n_6288 =  x_206 & ~n_6287;
assign n_6289 = ~x_206 &  n_6287;
assign n_6290 = ~n_6288 & ~n_6289;
assign n_6291 =  x_205 & ~n_1802;
assign n_6292 =  i_3 &  n_1802;
assign n_6293 = ~n_6291 & ~n_6292;
assign n_6294 =  x_205 & ~n_6293;
assign n_6295 = ~x_205 &  n_6293;
assign n_6296 = ~n_6294 & ~n_6295;
assign n_6297 =  x_204 & ~n_1802;
assign n_6298 =  i_2 &  n_1802;
assign n_6299 = ~n_6297 & ~n_6298;
assign n_6300 =  x_204 & ~n_6299;
assign n_6301 = ~x_204 &  n_6299;
assign n_6302 = ~n_6300 & ~n_6301;
assign n_6303 =  x_203 & ~n_1802;
assign n_6304 =  i_1 &  n_1802;
assign n_6305 = ~n_6303 & ~n_6304;
assign n_6306 =  x_203 & ~n_6305;
assign n_6307 = ~x_203 &  n_6305;
assign n_6308 = ~n_6306 & ~n_6307;
assign n_6309 =  x_202 & ~n_1359;
assign n_6310 =  i_32 &  n_1359;
assign n_6311 = ~n_6309 & ~n_6310;
assign n_6312 =  x_202 & ~n_6311;
assign n_6313 = ~x_202 &  n_6311;
assign n_6314 = ~n_6312 & ~n_6313;
assign n_6315 =  x_201 & ~n_1359;
assign n_6316 =  i_31 &  n_1359;
assign n_6317 = ~n_6315 & ~n_6316;
assign n_6318 =  x_201 & ~n_6317;
assign n_6319 = ~x_201 &  n_6317;
assign n_6320 = ~n_6318 & ~n_6319;
assign n_6321 =  x_200 & ~n_1359;
assign n_6322 =  i_30 &  n_1359;
assign n_6323 = ~n_6321 & ~n_6322;
assign n_6324 =  x_200 & ~n_6323;
assign n_6325 = ~x_200 &  n_6323;
assign n_6326 = ~n_6324 & ~n_6325;
assign n_6327 =  x_199 & ~n_1359;
assign n_6328 =  i_29 &  n_1359;
assign n_6329 = ~n_6327 & ~n_6328;
assign n_6330 =  x_199 & ~n_6329;
assign n_6331 = ~x_199 &  n_6329;
assign n_6332 = ~n_6330 & ~n_6331;
assign n_6333 =  x_198 & ~n_1359;
assign n_6334 =  i_28 &  n_1359;
assign n_6335 = ~n_6333 & ~n_6334;
assign n_6336 =  x_198 & ~n_6335;
assign n_6337 = ~x_198 &  n_6335;
assign n_6338 = ~n_6336 & ~n_6337;
assign n_6339 =  x_197 & ~n_1359;
assign n_6340 =  i_27 &  n_1359;
assign n_6341 = ~n_6339 & ~n_6340;
assign n_6342 =  x_197 & ~n_6341;
assign n_6343 = ~x_197 &  n_6341;
assign n_6344 = ~n_6342 & ~n_6343;
assign n_6345 =  x_196 & ~n_1359;
assign n_6346 =  i_26 &  n_1359;
assign n_6347 = ~n_6345 & ~n_6346;
assign n_6348 =  x_196 & ~n_6347;
assign n_6349 = ~x_196 &  n_6347;
assign n_6350 = ~n_6348 & ~n_6349;
assign n_6351 =  x_195 & ~n_1359;
assign n_6352 =  i_25 &  n_1359;
assign n_6353 = ~n_6351 & ~n_6352;
assign n_6354 =  x_195 & ~n_6353;
assign n_6355 = ~x_195 &  n_6353;
assign n_6356 = ~n_6354 & ~n_6355;
assign n_6357 =  x_194 & ~n_1359;
assign n_6358 =  i_24 &  n_1359;
assign n_6359 = ~n_6357 & ~n_6358;
assign n_6360 =  x_194 & ~n_6359;
assign n_6361 = ~x_194 &  n_6359;
assign n_6362 = ~n_6360 & ~n_6361;
assign n_6363 =  x_193 & ~n_1359;
assign n_6364 =  i_23 &  n_1359;
assign n_6365 = ~n_6363 & ~n_6364;
assign n_6366 =  x_193 & ~n_6365;
assign n_6367 = ~x_193 &  n_6365;
assign n_6368 = ~n_6366 & ~n_6367;
assign n_6369 =  x_192 & ~n_1359;
assign n_6370 =  i_22 &  n_1359;
assign n_6371 = ~n_6369 & ~n_6370;
assign n_6372 =  x_192 & ~n_6371;
assign n_6373 = ~x_192 &  n_6371;
assign n_6374 = ~n_6372 & ~n_6373;
assign n_6375 =  x_191 & ~n_1359;
assign n_6376 =  i_21 &  n_1359;
assign n_6377 = ~n_6375 & ~n_6376;
assign n_6378 =  x_191 & ~n_6377;
assign n_6379 = ~x_191 &  n_6377;
assign n_6380 = ~n_6378 & ~n_6379;
assign n_6381 =  x_190 & ~n_1359;
assign n_6382 =  i_20 &  n_1359;
assign n_6383 = ~n_6381 & ~n_6382;
assign n_6384 =  x_190 & ~n_6383;
assign n_6385 = ~x_190 &  n_6383;
assign n_6386 = ~n_6384 & ~n_6385;
assign n_6387 =  x_189 & ~n_1359;
assign n_6388 =  i_19 &  n_1359;
assign n_6389 = ~n_6387 & ~n_6388;
assign n_6390 =  x_189 & ~n_6389;
assign n_6391 = ~x_189 &  n_6389;
assign n_6392 = ~n_6390 & ~n_6391;
assign n_6393 =  x_188 & ~n_1359;
assign n_6394 =  i_18 &  n_1359;
assign n_6395 = ~n_6393 & ~n_6394;
assign n_6396 =  x_188 & ~n_6395;
assign n_6397 = ~x_188 &  n_6395;
assign n_6398 = ~n_6396 & ~n_6397;
assign n_6399 =  x_187 & ~n_1359;
assign n_6400 =  i_17 &  n_1359;
assign n_6401 = ~n_6399 & ~n_6400;
assign n_6402 =  x_187 & ~n_6401;
assign n_6403 = ~x_187 &  n_6401;
assign n_6404 = ~n_6402 & ~n_6403;
assign n_6405 =  x_186 & ~n_1359;
assign n_6406 =  i_16 &  n_1359;
assign n_6407 = ~n_6405 & ~n_6406;
assign n_6408 =  x_186 & ~n_6407;
assign n_6409 = ~x_186 &  n_6407;
assign n_6410 = ~n_6408 & ~n_6409;
assign n_6411 =  x_185 & ~n_1359;
assign n_6412 =  i_15 &  n_1359;
assign n_6413 = ~n_6411 & ~n_6412;
assign n_6414 =  x_185 & ~n_6413;
assign n_6415 = ~x_185 &  n_6413;
assign n_6416 = ~n_6414 & ~n_6415;
assign n_6417 =  x_184 & ~n_1359;
assign n_6418 =  i_14 &  n_1359;
assign n_6419 = ~n_6417 & ~n_6418;
assign n_6420 =  x_184 & ~n_6419;
assign n_6421 = ~x_184 &  n_6419;
assign n_6422 = ~n_6420 & ~n_6421;
assign n_6423 =  x_183 & ~n_1359;
assign n_6424 =  i_13 &  n_1359;
assign n_6425 = ~n_6423 & ~n_6424;
assign n_6426 =  x_183 & ~n_6425;
assign n_6427 = ~x_183 &  n_6425;
assign n_6428 = ~n_6426 & ~n_6427;
assign n_6429 =  x_182 & ~n_1359;
assign n_6430 =  i_12 &  n_1359;
assign n_6431 = ~n_6429 & ~n_6430;
assign n_6432 =  x_182 & ~n_6431;
assign n_6433 = ~x_182 &  n_6431;
assign n_6434 = ~n_6432 & ~n_6433;
assign n_6435 =  x_181 & ~n_1359;
assign n_6436 =  i_11 &  n_1359;
assign n_6437 = ~n_6435 & ~n_6436;
assign n_6438 =  x_181 & ~n_6437;
assign n_6439 = ~x_181 &  n_6437;
assign n_6440 = ~n_6438 & ~n_6439;
assign n_6441 =  x_180 & ~n_1359;
assign n_6442 =  i_10 &  n_1359;
assign n_6443 = ~n_6441 & ~n_6442;
assign n_6444 =  x_180 & ~n_6443;
assign n_6445 = ~x_180 &  n_6443;
assign n_6446 = ~n_6444 & ~n_6445;
assign n_6447 =  x_179 & ~n_1359;
assign n_6448 =  i_9 &  n_1359;
assign n_6449 = ~n_6447 & ~n_6448;
assign n_6450 =  x_179 & ~n_6449;
assign n_6451 = ~x_179 &  n_6449;
assign n_6452 = ~n_6450 & ~n_6451;
assign n_6453 =  x_178 & ~n_1359;
assign n_6454 =  i_8 &  n_1359;
assign n_6455 = ~n_6453 & ~n_6454;
assign n_6456 =  x_178 & ~n_6455;
assign n_6457 = ~x_178 &  n_6455;
assign n_6458 = ~n_6456 & ~n_6457;
assign n_6459 =  x_177 & ~n_1359;
assign n_6460 =  i_7 &  n_1359;
assign n_6461 = ~n_6459 & ~n_6460;
assign n_6462 =  x_177 & ~n_6461;
assign n_6463 = ~x_177 &  n_6461;
assign n_6464 = ~n_6462 & ~n_6463;
assign n_6465 =  x_176 & ~n_1359;
assign n_6466 =  i_6 &  n_1359;
assign n_6467 = ~n_6465 & ~n_6466;
assign n_6468 =  x_176 & ~n_6467;
assign n_6469 = ~x_176 &  n_6467;
assign n_6470 = ~n_6468 & ~n_6469;
assign n_6471 =  x_175 & ~n_1359;
assign n_6472 =  i_5 &  n_1359;
assign n_6473 = ~n_6471 & ~n_6472;
assign n_6474 =  x_175 & ~n_6473;
assign n_6475 = ~x_175 &  n_6473;
assign n_6476 = ~n_6474 & ~n_6475;
assign n_6477 =  x_174 & ~n_1359;
assign n_6478 =  i_4 &  n_1359;
assign n_6479 = ~n_6477 & ~n_6478;
assign n_6480 =  x_174 & ~n_6479;
assign n_6481 = ~x_174 &  n_6479;
assign n_6482 = ~n_6480 & ~n_6481;
assign n_6483 =  x_173 & ~n_1359;
assign n_6484 =  i_3 &  n_1359;
assign n_6485 = ~n_6483 & ~n_6484;
assign n_6486 =  x_173 & ~n_6485;
assign n_6487 = ~x_173 &  n_6485;
assign n_6488 = ~n_6486 & ~n_6487;
assign n_6489 =  x_172 & ~n_1359;
assign n_6490 =  i_2 &  n_1359;
assign n_6491 = ~n_6489 & ~n_6490;
assign n_6492 =  x_172 & ~n_6491;
assign n_6493 = ~x_172 &  n_6491;
assign n_6494 = ~n_6492 & ~n_6493;
assign n_6495 =  x_171 & ~n_1359;
assign n_6496 =  i_1 &  n_1359;
assign n_6497 = ~n_6495 & ~n_6496;
assign n_6498 =  x_171 & ~n_6497;
assign n_6499 = ~x_171 &  n_6497;
assign n_6500 = ~n_6498 & ~n_6499;
assign n_6501 = ~x_40 &  n_891;
assign n_6502 = ~x_41 & ~n_814;
assign n_6503 = ~n_6501 &  n_6502;
assign n_6504 =  x_41 & ~n_1841;
assign n_6505 =  x_42 & ~n_6504;
assign n_6506 = ~n_6503 &  n_6505;
assign n_6507 =  x_170 & ~n_6506;
assign n_6508 =  x_934 &  n_2414;
assign n_6509 =  x_1062 &  n_1542;
assign n_6510 = ~n_6508 & ~n_6509;
assign n_6511 = ~n_6507 &  n_6510;
assign n_6512 =  x_170 & ~n_6511;
assign n_6513 = ~x_170 &  n_6511;
assign n_6514 = ~n_6512 & ~n_6513;
assign n_6515 =  x_169 & ~n_6506;
assign n_6516 =  x_933 &  n_2414;
assign n_6517 =  x_1061 &  n_1542;
assign n_6518 = ~n_6516 & ~n_6517;
assign n_6519 = ~n_6515 &  n_6518;
assign n_6520 =  x_169 & ~n_6519;
assign n_6521 = ~x_169 &  n_6519;
assign n_6522 = ~n_6520 & ~n_6521;
assign n_6523 =  x_168 & ~n_6506;
assign n_6524 =  x_932 &  n_2414;
assign n_6525 =  x_1060 &  n_1542;
assign n_6526 = ~n_6524 & ~n_6525;
assign n_6527 = ~n_6523 &  n_6526;
assign n_6528 =  x_168 & ~n_6527;
assign n_6529 = ~x_168 &  n_6527;
assign n_6530 = ~n_6528 & ~n_6529;
assign n_6531 =  x_167 & ~n_6506;
assign n_6532 =  x_931 &  n_2414;
assign n_6533 =  x_1059 &  n_1542;
assign n_6534 = ~n_6532 & ~n_6533;
assign n_6535 = ~n_6531 &  n_6534;
assign n_6536 =  x_167 & ~n_6535;
assign n_6537 = ~x_167 &  n_6535;
assign n_6538 = ~n_6536 & ~n_6537;
assign n_6539 =  x_166 & ~n_6506;
assign n_6540 =  x_930 &  n_2414;
assign n_6541 =  x_1058 &  n_1542;
assign n_6542 = ~n_6540 & ~n_6541;
assign n_6543 = ~n_6539 &  n_6542;
assign n_6544 =  x_166 & ~n_6543;
assign n_6545 = ~x_166 &  n_6543;
assign n_6546 = ~n_6544 & ~n_6545;
assign n_6547 =  x_165 & ~n_6506;
assign n_6548 =  x_929 &  n_2414;
assign n_6549 =  x_1057 &  n_1542;
assign n_6550 = ~n_6548 & ~n_6549;
assign n_6551 = ~n_6547 &  n_6550;
assign n_6552 =  x_165 & ~n_6551;
assign n_6553 = ~x_165 &  n_6551;
assign n_6554 = ~n_6552 & ~n_6553;
assign n_6555 =  x_164 & ~n_6506;
assign n_6556 =  x_928 &  n_2414;
assign n_6557 =  x_1056 &  n_1542;
assign n_6558 = ~n_6556 & ~n_6557;
assign n_6559 = ~n_6555 &  n_6558;
assign n_6560 =  x_164 & ~n_6559;
assign n_6561 = ~x_164 &  n_6559;
assign n_6562 = ~n_6560 & ~n_6561;
assign n_6563 =  x_163 & ~n_6506;
assign n_6564 =  x_927 &  n_2414;
assign n_6565 =  x_1055 &  n_1542;
assign n_6566 = ~n_6564 & ~n_6565;
assign n_6567 = ~n_6563 &  n_6566;
assign n_6568 =  x_163 & ~n_6567;
assign n_6569 = ~x_163 &  n_6567;
assign n_6570 = ~n_6568 & ~n_6569;
assign n_6571 =  x_162 & ~n_6506;
assign n_6572 =  x_926 &  n_2414;
assign n_6573 =  x_1054 &  n_1542;
assign n_6574 = ~n_6572 & ~n_6573;
assign n_6575 = ~n_6571 &  n_6574;
assign n_6576 =  x_162 & ~n_6575;
assign n_6577 = ~x_162 &  n_6575;
assign n_6578 = ~n_6576 & ~n_6577;
assign n_6579 =  x_161 & ~n_6506;
assign n_6580 =  x_925 &  n_2414;
assign n_6581 =  x_1053 &  n_1542;
assign n_6582 = ~n_6580 & ~n_6581;
assign n_6583 = ~n_6579 &  n_6582;
assign n_6584 =  x_161 & ~n_6583;
assign n_6585 = ~x_161 &  n_6583;
assign n_6586 = ~n_6584 & ~n_6585;
assign n_6587 =  x_160 & ~n_6506;
assign n_6588 =  x_924 &  n_2414;
assign n_6589 =  x_1052 &  n_1542;
assign n_6590 = ~n_6588 & ~n_6589;
assign n_6591 = ~n_6587 &  n_6590;
assign n_6592 =  x_160 & ~n_6591;
assign n_6593 = ~x_160 &  n_6591;
assign n_6594 = ~n_6592 & ~n_6593;
assign n_6595 =  x_159 & ~n_6506;
assign n_6596 =  x_923 &  n_2414;
assign n_6597 =  x_1051 &  n_1542;
assign n_6598 = ~n_6596 & ~n_6597;
assign n_6599 = ~n_6595 &  n_6598;
assign n_6600 =  x_159 & ~n_6599;
assign n_6601 = ~x_159 &  n_6599;
assign n_6602 = ~n_6600 & ~n_6601;
assign n_6603 =  x_158 & ~n_6506;
assign n_6604 =  x_922 &  n_2414;
assign n_6605 =  x_1050 &  n_1542;
assign n_6606 = ~n_6604 & ~n_6605;
assign n_6607 = ~n_6603 &  n_6606;
assign n_6608 =  x_158 & ~n_6607;
assign n_6609 = ~x_158 &  n_6607;
assign n_6610 = ~n_6608 & ~n_6609;
assign n_6611 =  x_157 & ~n_6506;
assign n_6612 =  x_921 &  n_2414;
assign n_6613 =  x_1049 &  n_1542;
assign n_6614 = ~n_6612 & ~n_6613;
assign n_6615 = ~n_6611 &  n_6614;
assign n_6616 =  x_157 & ~n_6615;
assign n_6617 = ~x_157 &  n_6615;
assign n_6618 = ~n_6616 & ~n_6617;
assign n_6619 =  x_156 & ~n_6506;
assign n_6620 =  x_920 &  n_2414;
assign n_6621 =  x_1048 &  n_1542;
assign n_6622 = ~n_6620 & ~n_6621;
assign n_6623 = ~n_6619 &  n_6622;
assign n_6624 =  x_156 & ~n_6623;
assign n_6625 = ~x_156 &  n_6623;
assign n_6626 = ~n_6624 & ~n_6625;
assign n_6627 =  x_155 & ~n_6506;
assign n_6628 =  x_919 &  n_2414;
assign n_6629 =  x_1047 &  n_1542;
assign n_6630 = ~n_6628 & ~n_6629;
assign n_6631 = ~n_6627 &  n_6630;
assign n_6632 =  x_155 & ~n_6631;
assign n_6633 = ~x_155 &  n_6631;
assign n_6634 = ~n_6632 & ~n_6633;
assign n_6635 =  x_154 & ~n_6506;
assign n_6636 =  x_918 &  n_2414;
assign n_6637 =  x_1046 &  n_1542;
assign n_6638 = ~n_6636 & ~n_6637;
assign n_6639 = ~n_6635 &  n_6638;
assign n_6640 =  x_154 & ~n_6639;
assign n_6641 = ~x_154 &  n_6639;
assign n_6642 = ~n_6640 & ~n_6641;
assign n_6643 =  x_153 & ~n_6506;
assign n_6644 =  x_917 &  n_2414;
assign n_6645 =  x_1045 &  n_1542;
assign n_6646 = ~n_6644 & ~n_6645;
assign n_6647 = ~n_6643 &  n_6646;
assign n_6648 =  x_153 & ~n_6647;
assign n_6649 = ~x_153 &  n_6647;
assign n_6650 = ~n_6648 & ~n_6649;
assign n_6651 =  x_152 & ~n_6506;
assign n_6652 =  x_916 &  n_2414;
assign n_6653 =  x_1044 &  n_1542;
assign n_6654 = ~n_6652 & ~n_6653;
assign n_6655 = ~n_6651 &  n_6654;
assign n_6656 =  x_152 & ~n_6655;
assign n_6657 = ~x_152 &  n_6655;
assign n_6658 = ~n_6656 & ~n_6657;
assign n_6659 =  x_151 & ~n_6506;
assign n_6660 =  x_915 &  n_2414;
assign n_6661 =  x_1043 &  n_1542;
assign n_6662 = ~n_6660 & ~n_6661;
assign n_6663 = ~n_6659 &  n_6662;
assign n_6664 =  x_151 & ~n_6663;
assign n_6665 = ~x_151 &  n_6663;
assign n_6666 = ~n_6664 & ~n_6665;
assign n_6667 =  x_150 & ~n_6506;
assign n_6668 =  x_914 &  n_2414;
assign n_6669 =  x_1042 &  n_1542;
assign n_6670 = ~n_6668 & ~n_6669;
assign n_6671 = ~n_6667 &  n_6670;
assign n_6672 =  x_150 & ~n_6671;
assign n_6673 = ~x_150 &  n_6671;
assign n_6674 = ~n_6672 & ~n_6673;
assign n_6675 =  x_149 & ~n_6506;
assign n_6676 =  x_913 &  n_2414;
assign n_6677 =  x_1041 &  n_1542;
assign n_6678 = ~n_6676 & ~n_6677;
assign n_6679 = ~n_6675 &  n_6678;
assign n_6680 =  x_149 & ~n_6679;
assign n_6681 = ~x_149 &  n_6679;
assign n_6682 = ~n_6680 & ~n_6681;
assign n_6683 =  x_148 & ~n_6506;
assign n_6684 =  x_912 &  n_2414;
assign n_6685 =  x_1040 &  n_1542;
assign n_6686 = ~n_6684 & ~n_6685;
assign n_6687 = ~n_6683 &  n_6686;
assign n_6688 =  x_148 & ~n_6687;
assign n_6689 = ~x_148 &  n_6687;
assign n_6690 = ~n_6688 & ~n_6689;
assign n_6691 =  x_147 & ~n_6506;
assign n_6692 =  x_911 &  n_2414;
assign n_6693 =  x_1039 &  n_1542;
assign n_6694 = ~n_6692 & ~n_6693;
assign n_6695 = ~n_6691 &  n_6694;
assign n_6696 =  x_147 & ~n_6695;
assign n_6697 = ~x_147 &  n_6695;
assign n_6698 = ~n_6696 & ~n_6697;
assign n_6699 =  x_146 & ~n_6506;
assign n_6700 =  x_910 &  n_2414;
assign n_6701 =  x_1038 &  n_1542;
assign n_6702 = ~n_6700 & ~n_6701;
assign n_6703 = ~n_6699 &  n_6702;
assign n_6704 =  x_146 & ~n_6703;
assign n_6705 = ~x_146 &  n_6703;
assign n_6706 = ~n_6704 & ~n_6705;
assign n_6707 =  x_145 & ~n_6506;
assign n_6708 =  x_909 &  n_2414;
assign n_6709 =  x_1037 &  n_1542;
assign n_6710 = ~n_6708 & ~n_6709;
assign n_6711 = ~n_6707 &  n_6710;
assign n_6712 =  x_145 & ~n_6711;
assign n_6713 = ~x_145 &  n_6711;
assign n_6714 = ~n_6712 & ~n_6713;
assign n_6715 =  x_144 & ~n_6506;
assign n_6716 =  x_908 &  n_2414;
assign n_6717 =  x_1036 &  n_1542;
assign n_6718 = ~n_6716 & ~n_6717;
assign n_6719 = ~n_6715 &  n_6718;
assign n_6720 =  x_144 & ~n_6719;
assign n_6721 = ~x_144 &  n_6719;
assign n_6722 = ~n_6720 & ~n_6721;
assign n_6723 =  x_143 & ~n_6506;
assign n_6724 =  x_907 &  n_2414;
assign n_6725 =  x_1035 &  n_1542;
assign n_6726 = ~n_6724 & ~n_6725;
assign n_6727 = ~n_6723 &  n_6726;
assign n_6728 =  x_143 & ~n_6727;
assign n_6729 = ~x_143 &  n_6727;
assign n_6730 = ~n_6728 & ~n_6729;
assign n_6731 =  x_142 & ~n_6506;
assign n_6732 =  x_906 &  n_2414;
assign n_6733 =  x_1034 &  n_1542;
assign n_6734 = ~n_6732 & ~n_6733;
assign n_6735 = ~n_6731 &  n_6734;
assign n_6736 =  x_142 & ~n_6735;
assign n_6737 = ~x_142 &  n_6735;
assign n_6738 = ~n_6736 & ~n_6737;
assign n_6739 =  x_141 & ~n_6506;
assign n_6740 =  x_905 &  n_2414;
assign n_6741 =  x_1033 &  n_1542;
assign n_6742 = ~n_6740 & ~n_6741;
assign n_6743 = ~n_6739 &  n_6742;
assign n_6744 =  x_141 & ~n_6743;
assign n_6745 = ~x_141 &  n_6743;
assign n_6746 = ~n_6744 & ~n_6745;
assign n_6747 =  x_140 & ~n_6506;
assign n_6748 =  x_904 &  n_2414;
assign n_6749 =  x_1032 &  n_1542;
assign n_6750 = ~n_6748 & ~n_6749;
assign n_6751 = ~n_6747 &  n_6750;
assign n_6752 =  x_140 & ~n_6751;
assign n_6753 = ~x_140 &  n_6751;
assign n_6754 = ~n_6752 & ~n_6753;
assign n_6755 =  x_139 & ~n_6506;
assign n_6756 =  x_903 &  n_2414;
assign n_6757 =  x_1031 &  n_1542;
assign n_6758 = ~n_6756 & ~n_6757;
assign n_6759 = ~n_6755 &  n_6758;
assign n_6760 =  x_139 & ~n_6759;
assign n_6761 = ~x_139 &  n_6759;
assign n_6762 = ~n_6760 & ~n_6761;
assign n_6763 =  x_138 & ~n_6506;
assign n_6764 =  x_1030 &  n_2414;
assign n_6765 =  x_74 &  n_1542;
assign n_6766 = ~n_6764 & ~n_6765;
assign n_6767 = ~n_6763 &  n_6766;
assign n_6768 =  x_138 & ~n_6767;
assign n_6769 = ~x_138 &  n_6767;
assign n_6770 = ~n_6768 & ~n_6769;
assign n_6771 =  x_137 & ~n_6506;
assign n_6772 =  x_1029 &  n_2414;
assign n_6773 =  x_73 &  n_1542;
assign n_6774 = ~n_6772 & ~n_6773;
assign n_6775 = ~n_6771 &  n_6774;
assign n_6776 =  x_137 & ~n_6775;
assign n_6777 = ~x_137 &  n_6775;
assign n_6778 = ~n_6776 & ~n_6777;
assign n_6779 =  x_136 & ~n_6506;
assign n_6780 =  x_1028 &  n_2414;
assign n_6781 =  x_72 &  n_1542;
assign n_6782 = ~n_6780 & ~n_6781;
assign n_6783 = ~n_6779 &  n_6782;
assign n_6784 =  x_136 & ~n_6783;
assign n_6785 = ~x_136 &  n_6783;
assign n_6786 = ~n_6784 & ~n_6785;
assign n_6787 =  x_135 & ~n_6506;
assign n_6788 =  x_1027 &  n_2414;
assign n_6789 =  x_71 &  n_1542;
assign n_6790 = ~n_6788 & ~n_6789;
assign n_6791 = ~n_6787 &  n_6790;
assign n_6792 =  x_135 & ~n_6791;
assign n_6793 = ~x_135 &  n_6791;
assign n_6794 = ~n_6792 & ~n_6793;
assign n_6795 =  x_134 & ~n_6506;
assign n_6796 =  x_1026 &  n_2414;
assign n_6797 =  x_70 &  n_1542;
assign n_6798 = ~n_6796 & ~n_6797;
assign n_6799 = ~n_6795 &  n_6798;
assign n_6800 =  x_134 & ~n_6799;
assign n_6801 = ~x_134 &  n_6799;
assign n_6802 = ~n_6800 & ~n_6801;
assign n_6803 =  x_133 & ~n_6506;
assign n_6804 =  x_1025 &  n_2414;
assign n_6805 =  x_69 &  n_1542;
assign n_6806 = ~n_6804 & ~n_6805;
assign n_6807 = ~n_6803 &  n_6806;
assign n_6808 =  x_133 & ~n_6807;
assign n_6809 = ~x_133 &  n_6807;
assign n_6810 = ~n_6808 & ~n_6809;
assign n_6811 =  x_132 & ~n_6506;
assign n_6812 =  x_1024 &  n_2414;
assign n_6813 =  x_68 &  n_1542;
assign n_6814 = ~n_6812 & ~n_6813;
assign n_6815 = ~n_6811 &  n_6814;
assign n_6816 =  x_132 & ~n_6815;
assign n_6817 = ~x_132 &  n_6815;
assign n_6818 = ~n_6816 & ~n_6817;
assign n_6819 =  x_131 & ~n_6506;
assign n_6820 =  x_1023 &  n_2414;
assign n_6821 =  x_67 &  n_1542;
assign n_6822 = ~n_6820 & ~n_6821;
assign n_6823 = ~n_6819 &  n_6822;
assign n_6824 =  x_131 & ~n_6823;
assign n_6825 = ~x_131 &  n_6823;
assign n_6826 = ~n_6824 & ~n_6825;
assign n_6827 =  x_130 & ~n_6506;
assign n_6828 =  x_1022 &  n_2414;
assign n_6829 =  x_66 &  n_1542;
assign n_6830 = ~n_6828 & ~n_6829;
assign n_6831 = ~n_6827 &  n_6830;
assign n_6832 =  x_130 & ~n_6831;
assign n_6833 = ~x_130 &  n_6831;
assign n_6834 = ~n_6832 & ~n_6833;
assign n_6835 =  x_129 & ~n_6506;
assign n_6836 =  x_1021 &  n_2414;
assign n_6837 =  x_65 &  n_1542;
assign n_6838 = ~n_6836 & ~n_6837;
assign n_6839 = ~n_6835 &  n_6838;
assign n_6840 =  x_129 & ~n_6839;
assign n_6841 = ~x_129 &  n_6839;
assign n_6842 = ~n_6840 & ~n_6841;
assign n_6843 =  x_128 & ~n_6506;
assign n_6844 =  x_1020 &  n_2414;
assign n_6845 =  x_64 &  n_1542;
assign n_6846 = ~n_6844 & ~n_6845;
assign n_6847 = ~n_6843 &  n_6846;
assign n_6848 =  x_128 & ~n_6847;
assign n_6849 = ~x_128 &  n_6847;
assign n_6850 = ~n_6848 & ~n_6849;
assign n_6851 =  x_127 & ~n_6506;
assign n_6852 =  x_1019 &  n_2414;
assign n_6853 =  x_63 &  n_1542;
assign n_6854 = ~n_6852 & ~n_6853;
assign n_6855 = ~n_6851 &  n_6854;
assign n_6856 =  x_127 & ~n_6855;
assign n_6857 = ~x_127 &  n_6855;
assign n_6858 = ~n_6856 & ~n_6857;
assign n_6859 =  x_126 & ~n_6506;
assign n_6860 =  x_1018 &  n_2414;
assign n_6861 =  x_62 &  n_1542;
assign n_6862 = ~n_6860 & ~n_6861;
assign n_6863 = ~n_6859 &  n_6862;
assign n_6864 =  x_126 & ~n_6863;
assign n_6865 = ~x_126 &  n_6863;
assign n_6866 = ~n_6864 & ~n_6865;
assign n_6867 =  x_125 & ~n_6506;
assign n_6868 =  x_1017 &  n_2414;
assign n_6869 =  x_61 &  n_1542;
assign n_6870 = ~n_6868 & ~n_6869;
assign n_6871 = ~n_6867 &  n_6870;
assign n_6872 =  x_125 & ~n_6871;
assign n_6873 = ~x_125 &  n_6871;
assign n_6874 = ~n_6872 & ~n_6873;
assign n_6875 =  x_124 & ~n_6506;
assign n_6876 =  x_1016 &  n_2414;
assign n_6877 =  x_60 &  n_1542;
assign n_6878 = ~n_6876 & ~n_6877;
assign n_6879 = ~n_6875 &  n_6878;
assign n_6880 =  x_124 & ~n_6879;
assign n_6881 = ~x_124 &  n_6879;
assign n_6882 = ~n_6880 & ~n_6881;
assign n_6883 =  x_123 & ~n_6506;
assign n_6884 =  x_1015 &  n_2414;
assign n_6885 =  x_59 &  n_1542;
assign n_6886 = ~n_6884 & ~n_6885;
assign n_6887 = ~n_6883 &  n_6886;
assign n_6888 =  x_123 & ~n_6887;
assign n_6889 = ~x_123 &  n_6887;
assign n_6890 = ~n_6888 & ~n_6889;
assign n_6891 =  x_122 & ~n_6506;
assign n_6892 =  x_1014 &  n_2414;
assign n_6893 =  x_58 &  n_1542;
assign n_6894 = ~n_6892 & ~n_6893;
assign n_6895 = ~n_6891 &  n_6894;
assign n_6896 =  x_122 & ~n_6895;
assign n_6897 = ~x_122 &  n_6895;
assign n_6898 = ~n_6896 & ~n_6897;
assign n_6899 =  x_121 & ~n_6506;
assign n_6900 =  x_1013 &  n_2414;
assign n_6901 =  x_57 &  n_1542;
assign n_6902 = ~n_6900 & ~n_6901;
assign n_6903 = ~n_6899 &  n_6902;
assign n_6904 =  x_121 & ~n_6903;
assign n_6905 = ~x_121 &  n_6903;
assign n_6906 = ~n_6904 & ~n_6905;
assign n_6907 =  x_120 & ~n_6506;
assign n_6908 =  x_1012 &  n_2414;
assign n_6909 =  x_56 &  n_1542;
assign n_6910 = ~n_6908 & ~n_6909;
assign n_6911 = ~n_6907 &  n_6910;
assign n_6912 =  x_120 & ~n_6911;
assign n_6913 = ~x_120 &  n_6911;
assign n_6914 = ~n_6912 & ~n_6913;
assign n_6915 =  x_119 & ~n_6506;
assign n_6916 =  x_1011 &  n_2414;
assign n_6917 =  x_55 &  n_1542;
assign n_6918 = ~n_6916 & ~n_6917;
assign n_6919 = ~n_6915 &  n_6918;
assign n_6920 =  x_119 & ~n_6919;
assign n_6921 = ~x_119 &  n_6919;
assign n_6922 = ~n_6920 & ~n_6921;
assign n_6923 =  x_118 & ~n_6506;
assign n_6924 =  x_1010 &  n_2414;
assign n_6925 =  x_54 &  n_1542;
assign n_6926 = ~n_6924 & ~n_6925;
assign n_6927 = ~n_6923 &  n_6926;
assign n_6928 =  x_118 & ~n_6927;
assign n_6929 = ~x_118 &  n_6927;
assign n_6930 = ~n_6928 & ~n_6929;
assign n_6931 =  x_117 & ~n_6506;
assign n_6932 =  x_1009 &  n_2414;
assign n_6933 =  x_53 &  n_1542;
assign n_6934 = ~n_6932 & ~n_6933;
assign n_6935 = ~n_6931 &  n_6934;
assign n_6936 =  x_117 & ~n_6935;
assign n_6937 = ~x_117 &  n_6935;
assign n_6938 = ~n_6936 & ~n_6937;
assign n_6939 =  x_116 & ~n_6506;
assign n_6940 =  x_1008 &  n_2414;
assign n_6941 =  x_52 &  n_1542;
assign n_6942 = ~n_6940 & ~n_6941;
assign n_6943 = ~n_6939 &  n_6942;
assign n_6944 =  x_116 & ~n_6943;
assign n_6945 = ~x_116 &  n_6943;
assign n_6946 = ~n_6944 & ~n_6945;
assign n_6947 =  x_115 & ~n_6506;
assign n_6948 =  x_1007 &  n_2414;
assign n_6949 =  x_51 &  n_1542;
assign n_6950 = ~n_6948 & ~n_6949;
assign n_6951 = ~n_6947 &  n_6950;
assign n_6952 =  x_115 & ~n_6951;
assign n_6953 = ~x_115 &  n_6951;
assign n_6954 = ~n_6952 & ~n_6953;
assign n_6955 =  x_114 & ~n_6506;
assign n_6956 =  x_1006 &  n_2414;
assign n_6957 =  x_50 &  n_1542;
assign n_6958 = ~n_6956 & ~n_6957;
assign n_6959 = ~n_6955 &  n_6958;
assign n_6960 =  x_114 & ~n_6959;
assign n_6961 = ~x_114 &  n_6959;
assign n_6962 = ~n_6960 & ~n_6961;
assign n_6963 =  x_113 & ~n_6506;
assign n_6964 =  x_1005 &  n_2414;
assign n_6965 =  x_49 &  n_1542;
assign n_6966 = ~n_6964 & ~n_6965;
assign n_6967 = ~n_6963 &  n_6966;
assign n_6968 =  x_113 & ~n_6967;
assign n_6969 = ~x_113 &  n_6967;
assign n_6970 = ~n_6968 & ~n_6969;
assign n_6971 =  x_112 & ~n_6506;
assign n_6972 =  x_1004 &  n_2414;
assign n_6973 =  x_48 &  n_1542;
assign n_6974 = ~n_6972 & ~n_6973;
assign n_6975 = ~n_6971 &  n_6974;
assign n_6976 =  x_112 & ~n_6975;
assign n_6977 = ~x_112 &  n_6975;
assign n_6978 = ~n_6976 & ~n_6977;
assign n_6979 =  x_111 & ~n_6506;
assign n_6980 =  x_1003 &  n_2414;
assign n_6981 =  x_47 &  n_1542;
assign n_6982 = ~n_6980 & ~n_6981;
assign n_6983 = ~n_6979 &  n_6982;
assign n_6984 =  x_111 & ~n_6983;
assign n_6985 = ~x_111 &  n_6983;
assign n_6986 = ~n_6984 & ~n_6985;
assign n_6987 =  x_110 & ~n_6506;
assign n_6988 =  x_1002 &  n_2414;
assign n_6989 =  x_46 &  n_1542;
assign n_6990 = ~n_6988 & ~n_6989;
assign n_6991 = ~n_6987 &  n_6990;
assign n_6992 =  x_110 & ~n_6991;
assign n_6993 = ~x_110 &  n_6991;
assign n_6994 = ~n_6992 & ~n_6993;
assign n_6995 =  x_109 & ~n_6506;
assign n_6996 =  x_1001 &  n_2414;
assign n_6997 =  x_45 &  n_1542;
assign n_6998 = ~n_6996 & ~n_6997;
assign n_6999 = ~n_6995 &  n_6998;
assign n_7000 =  x_109 & ~n_6999;
assign n_7001 = ~x_109 &  n_6999;
assign n_7002 = ~n_7000 & ~n_7001;
assign n_7003 =  x_108 & ~n_6506;
assign n_7004 =  x_1000 &  n_2414;
assign n_7005 =  x_44 &  n_1542;
assign n_7006 = ~n_7004 & ~n_7005;
assign n_7007 = ~n_7003 &  n_7006;
assign n_7008 =  x_108 & ~n_7007;
assign n_7009 = ~x_108 &  n_7007;
assign n_7010 = ~n_7008 & ~n_7009;
assign n_7011 =  x_107 & ~n_6506;
assign n_7012 =  x_999 &  n_2414;
assign n_7013 =  x_43 &  n_1542;
assign n_7014 = ~n_7012 & ~n_7013;
assign n_7015 = ~n_7011 &  n_7014;
assign n_7016 =  x_107 & ~n_7015;
assign n_7017 = ~x_107 &  n_7015;
assign n_7018 = ~n_7016 & ~n_7017;
assign n_7019 =  x_106 & ~n_1270;
assign n_7020 = ~n_7019 & ~n_2828;
assign n_7021 =  x_106 & ~n_7020;
assign n_7022 = ~x_106 &  n_7020;
assign n_7023 = ~n_7021 & ~n_7022;
assign n_7024 =  x_105 & ~n_1270;
assign n_7025 = ~n_7024 & ~n_2834;
assign n_7026 =  x_105 & ~n_7025;
assign n_7027 = ~x_105 &  n_7025;
assign n_7028 = ~n_7026 & ~n_7027;
assign n_7029 =  x_104 & ~n_1270;
assign n_7030 = ~n_7029 & ~n_2840;
assign n_7031 =  x_104 & ~n_7030;
assign n_7032 = ~x_104 &  n_7030;
assign n_7033 = ~n_7031 & ~n_7032;
assign n_7034 =  x_103 & ~n_1270;
assign n_7035 = ~n_7034 & ~n_2846;
assign n_7036 =  x_103 & ~n_7035;
assign n_7037 = ~x_103 &  n_7035;
assign n_7038 = ~n_7036 & ~n_7037;
assign n_7039 =  x_102 & ~n_1270;
assign n_7040 = ~n_7039 & ~n_2852;
assign n_7041 =  x_102 & ~n_7040;
assign n_7042 = ~x_102 &  n_7040;
assign n_7043 = ~n_7041 & ~n_7042;
assign n_7044 =  x_101 & ~n_1270;
assign n_7045 = ~n_7044 & ~n_2858;
assign n_7046 =  x_101 & ~n_7045;
assign n_7047 = ~x_101 &  n_7045;
assign n_7048 = ~n_7046 & ~n_7047;
assign n_7049 =  x_100 & ~n_1270;
assign n_7050 = ~n_7049 & ~n_2864;
assign n_7051 =  x_100 & ~n_7050;
assign n_7052 = ~x_100 &  n_7050;
assign n_7053 = ~n_7051 & ~n_7052;
assign n_7054 =  x_99 & ~n_1270;
assign n_7055 = ~n_7054 & ~n_2870;
assign n_7056 =  x_99 & ~n_7055;
assign n_7057 = ~x_99 &  n_7055;
assign n_7058 = ~n_7056 & ~n_7057;
assign n_7059 =  x_98 & ~n_1270;
assign n_7060 = ~n_7059 & ~n_2876;
assign n_7061 =  x_98 & ~n_7060;
assign n_7062 = ~x_98 &  n_7060;
assign n_7063 = ~n_7061 & ~n_7062;
assign n_7064 =  x_97 & ~n_1270;
assign n_7065 = ~n_7064 & ~n_2882;
assign n_7066 =  x_97 & ~n_7065;
assign n_7067 = ~x_97 &  n_7065;
assign n_7068 = ~n_7066 & ~n_7067;
assign n_7069 =  x_96 & ~n_1270;
assign n_7070 = ~n_7069 & ~n_2888;
assign n_7071 =  x_96 & ~n_7070;
assign n_7072 = ~x_96 &  n_7070;
assign n_7073 = ~n_7071 & ~n_7072;
assign n_7074 =  x_95 & ~n_1270;
assign n_7075 = ~n_7074 & ~n_2894;
assign n_7076 =  x_95 & ~n_7075;
assign n_7077 = ~x_95 &  n_7075;
assign n_7078 = ~n_7076 & ~n_7077;
assign n_7079 =  x_94 & ~n_1270;
assign n_7080 = ~n_7079 & ~n_2900;
assign n_7081 =  x_94 & ~n_7080;
assign n_7082 = ~x_94 &  n_7080;
assign n_7083 = ~n_7081 & ~n_7082;
assign n_7084 =  x_93 & ~n_1270;
assign n_7085 = ~n_7084 & ~n_2906;
assign n_7086 =  x_93 & ~n_7085;
assign n_7087 = ~x_93 &  n_7085;
assign n_7088 = ~n_7086 & ~n_7087;
assign n_7089 =  x_92 & ~n_1270;
assign n_7090 = ~n_7089 & ~n_2912;
assign n_7091 =  x_92 & ~n_7090;
assign n_7092 = ~x_92 &  n_7090;
assign n_7093 = ~n_7091 & ~n_7092;
assign n_7094 =  x_91 & ~n_1270;
assign n_7095 = ~n_7094 & ~n_2918;
assign n_7096 =  x_91 & ~n_7095;
assign n_7097 = ~x_91 &  n_7095;
assign n_7098 = ~n_7096 & ~n_7097;
assign n_7099 =  x_90 & ~n_1270;
assign n_7100 = ~n_7099 & ~n_2924;
assign n_7101 =  x_90 & ~n_7100;
assign n_7102 = ~x_90 &  n_7100;
assign n_7103 = ~n_7101 & ~n_7102;
assign n_7104 =  x_89 & ~n_1270;
assign n_7105 = ~n_7104 & ~n_2930;
assign n_7106 =  x_89 & ~n_7105;
assign n_7107 = ~x_89 &  n_7105;
assign n_7108 = ~n_7106 & ~n_7107;
assign n_7109 =  x_88 & ~n_1270;
assign n_7110 = ~n_7109 & ~n_2936;
assign n_7111 =  x_88 & ~n_7110;
assign n_7112 = ~x_88 &  n_7110;
assign n_7113 = ~n_7111 & ~n_7112;
assign n_7114 =  x_87 & ~n_1270;
assign n_7115 = ~n_7114 & ~n_2942;
assign n_7116 =  x_87 & ~n_7115;
assign n_7117 = ~x_87 &  n_7115;
assign n_7118 = ~n_7116 & ~n_7117;
assign n_7119 =  x_86 & ~n_1270;
assign n_7120 = ~n_7119 & ~n_2948;
assign n_7121 =  x_86 & ~n_7120;
assign n_7122 = ~x_86 &  n_7120;
assign n_7123 = ~n_7121 & ~n_7122;
assign n_7124 =  x_85 & ~n_1270;
assign n_7125 = ~n_7124 & ~n_2954;
assign n_7126 =  x_85 & ~n_7125;
assign n_7127 = ~x_85 &  n_7125;
assign n_7128 = ~n_7126 & ~n_7127;
assign n_7129 =  x_84 & ~n_1270;
assign n_7130 = ~n_7129 & ~n_2960;
assign n_7131 =  x_84 & ~n_7130;
assign n_7132 = ~x_84 &  n_7130;
assign n_7133 = ~n_7131 & ~n_7132;
assign n_7134 =  x_83 & ~n_1270;
assign n_7135 = ~n_7134 & ~n_2966;
assign n_7136 =  x_83 & ~n_7135;
assign n_7137 = ~x_83 &  n_7135;
assign n_7138 = ~n_7136 & ~n_7137;
assign n_7139 =  x_82 & ~n_1270;
assign n_7140 = ~n_7139 & ~n_2972;
assign n_7141 =  x_82 & ~n_7140;
assign n_7142 = ~x_82 &  n_7140;
assign n_7143 = ~n_7141 & ~n_7142;
assign n_7144 =  x_81 & ~n_1270;
assign n_7145 = ~n_7144 & ~n_2978;
assign n_7146 =  x_81 & ~n_7145;
assign n_7147 = ~x_81 &  n_7145;
assign n_7148 = ~n_7146 & ~n_7147;
assign n_7149 =  x_80 & ~n_1270;
assign n_7150 = ~n_7149 & ~n_2984;
assign n_7151 =  x_80 & ~n_7150;
assign n_7152 = ~x_80 &  n_7150;
assign n_7153 = ~n_7151 & ~n_7152;
assign n_7154 =  x_79 & ~n_1270;
assign n_7155 = ~n_7154 & ~n_2990;
assign n_7156 =  x_79 & ~n_7155;
assign n_7157 = ~x_79 &  n_7155;
assign n_7158 = ~n_7156 & ~n_7157;
assign n_7159 =  x_78 & ~n_1270;
assign n_7160 = ~n_7159 & ~n_2996;
assign n_7161 =  x_78 & ~n_7160;
assign n_7162 = ~x_78 &  n_7160;
assign n_7163 = ~n_7161 & ~n_7162;
assign n_7164 =  x_77 & ~n_1270;
assign n_7165 = ~n_7164 & ~n_3002;
assign n_7166 =  x_77 & ~n_7165;
assign n_7167 = ~x_77 &  n_7165;
assign n_7168 = ~n_7166 & ~n_7167;
assign n_7169 =  x_76 & ~n_1270;
assign n_7170 = ~n_7169 & ~n_3008;
assign n_7171 =  x_76 & ~n_7170;
assign n_7172 = ~x_76 &  n_7170;
assign n_7173 = ~n_7171 & ~n_7172;
assign n_7174 =  x_75 & ~n_1270;
assign n_7175 = ~n_7174 & ~n_3014;
assign n_7176 =  x_75 & ~n_7175;
assign n_7177 = ~x_75 &  n_7175;
assign n_7178 = ~n_7176 & ~n_7177;
assign n_7179 =  x_74 & ~n_9;
assign n_7180 =  x_266 &  n_9;
assign n_7181 = ~n_7179 & ~n_7180;
assign n_7182 =  x_74 & ~n_7181;
assign n_7183 = ~x_74 &  n_7181;
assign n_7184 = ~n_7182 & ~n_7183;
assign n_7185 =  x_73 & ~n_9;
assign n_7186 =  x_265 &  n_9;
assign n_7187 = ~n_7185 & ~n_7186;
assign n_7188 =  x_73 & ~n_7187;
assign n_7189 = ~x_73 &  n_7187;
assign n_7190 = ~n_7188 & ~n_7189;
assign n_7191 =  x_72 & ~n_9;
assign n_7192 =  x_264 &  n_9;
assign n_7193 = ~n_7191 & ~n_7192;
assign n_7194 =  x_72 & ~n_7193;
assign n_7195 = ~x_72 &  n_7193;
assign n_7196 = ~n_7194 & ~n_7195;
assign n_7197 =  x_71 & ~n_9;
assign n_7198 =  x_263 &  n_9;
assign n_7199 = ~n_7197 & ~n_7198;
assign n_7200 =  x_71 & ~n_7199;
assign n_7201 = ~x_71 &  n_7199;
assign n_7202 = ~n_7200 & ~n_7201;
assign n_7203 =  x_70 & ~n_9;
assign n_7204 =  x_262 &  n_9;
assign n_7205 = ~n_7203 & ~n_7204;
assign n_7206 =  x_70 & ~n_7205;
assign n_7207 = ~x_70 &  n_7205;
assign n_7208 = ~n_7206 & ~n_7207;
assign n_7209 =  x_69 & ~n_9;
assign n_7210 =  x_261 &  n_9;
assign n_7211 = ~n_7209 & ~n_7210;
assign n_7212 =  x_69 & ~n_7211;
assign n_7213 = ~x_69 &  n_7211;
assign n_7214 = ~n_7212 & ~n_7213;
assign n_7215 =  x_68 & ~n_9;
assign n_7216 =  x_260 &  n_9;
assign n_7217 = ~n_7215 & ~n_7216;
assign n_7218 =  x_68 & ~n_7217;
assign n_7219 = ~x_68 &  n_7217;
assign n_7220 = ~n_7218 & ~n_7219;
assign n_7221 =  x_67 & ~n_9;
assign n_7222 =  x_259 &  n_9;
assign n_7223 = ~n_7221 & ~n_7222;
assign n_7224 =  x_67 & ~n_7223;
assign n_7225 = ~x_67 &  n_7223;
assign n_7226 = ~n_7224 & ~n_7225;
assign n_7227 =  x_975 & ~n_1270;
assign n_7228 = ~n_2966 & ~n_7227;
assign n_7229 =  x_975 & ~n_7228;
assign n_7230 = ~x_975 &  n_7228;
assign n_7231 = ~n_7229 & ~n_7230;
assign n_7232 =  x_974 & ~n_1270;
assign n_7233 = ~n_2972 & ~n_7232;
assign n_7234 =  x_974 & ~n_7233;
assign n_7235 = ~x_974 &  n_7233;
assign n_7236 = ~n_7234 & ~n_7235;
assign n_7237 =  x_973 & ~n_1270;
assign n_7238 = ~n_2978 & ~n_7237;
assign n_7239 =  x_973 & ~n_7238;
assign n_7240 = ~x_973 &  n_7238;
assign n_7241 = ~n_7239 & ~n_7240;
assign n_7242 =  x_972 & ~n_1270;
assign n_7243 = ~n_2984 & ~n_7242;
assign n_7244 =  x_972 & ~n_7243;
assign n_7245 = ~x_972 &  n_7243;
assign n_7246 = ~n_7244 & ~n_7245;
assign n_7247 =  x_971 & ~n_1270;
assign n_7248 = ~n_2990 & ~n_7247;
assign n_7249 =  x_971 & ~n_7248;
assign n_7250 = ~x_971 &  n_7248;
assign n_7251 = ~n_7249 & ~n_7250;
assign n_7252 =  x_970 & ~n_1270;
assign n_7253 = ~n_2996 & ~n_7252;
assign n_7254 =  x_970 & ~n_7253;
assign n_7255 = ~x_970 &  n_7253;
assign n_7256 = ~n_7254 & ~n_7255;
assign n_7257 =  x_969 & ~n_1270;
assign n_7258 = ~n_3002 & ~n_7257;
assign n_7259 =  x_969 & ~n_7258;
assign n_7260 = ~x_969 &  n_7258;
assign n_7261 = ~n_7259 & ~n_7260;
assign n_7262 =  x_968 & ~n_1270;
assign n_7263 = ~n_3008 & ~n_7262;
assign n_7264 =  x_968 & ~n_7263;
assign n_7265 = ~x_968 &  n_7263;
assign n_7266 = ~n_7264 & ~n_7265;
assign n_7267 =  x_967 & ~n_1270;
assign n_7268 = ~n_3014 & ~n_7267;
assign n_7269 =  x_967 & ~n_7268;
assign n_7270 = ~x_967 &  n_7268;
assign n_7271 = ~n_7269 & ~n_7270;
assign n_7272 =  x_966 & ~n_6506;
assign n_7273 =  x_583 &  n_2414;
assign n_7274 =  x_456 &  n_1542;
assign n_7275 = ~n_7273 & ~n_7274;
assign n_7276 = ~n_7272 &  n_7275;
assign n_7277 =  x_966 & ~n_7276;
assign n_7278 = ~x_966 &  n_7276;
assign n_7279 = ~n_7277 & ~n_7278;
assign n_7280 =  x_965 & ~n_6506;
assign n_7281 =  x_582 &  n_2414;
assign n_7282 =  x_455 &  n_1542;
assign n_7283 = ~n_7281 & ~n_7282;
assign n_7284 = ~n_7280 &  n_7283;
assign n_7285 =  x_965 & ~n_7284;
assign n_7286 = ~x_965 &  n_7284;
assign n_7287 = ~n_7285 & ~n_7286;
assign n_7288 =  x_964 & ~n_6506;
assign n_7289 =  x_581 &  n_2414;
assign n_7290 =  x_454 &  n_1542;
assign n_7291 = ~n_7289 & ~n_7290;
assign n_7292 = ~n_7288 &  n_7291;
assign n_7293 =  x_964 & ~n_7292;
assign n_7294 = ~x_964 &  n_7292;
assign n_7295 = ~n_7293 & ~n_7294;
assign n_7296 =  x_963 & ~n_6506;
assign n_7297 =  x_580 &  n_2414;
assign n_7298 =  x_453 &  n_1542;
assign n_7299 = ~n_7297 & ~n_7298;
assign n_7300 = ~n_7296 &  n_7299;
assign n_7301 =  x_963 & ~n_7300;
assign n_7302 = ~x_963 &  n_7300;
assign n_7303 = ~n_7301 & ~n_7302;
assign n_7304 =  x_962 & ~n_6506;
assign n_7305 =  x_579 &  n_2414;
assign n_7306 =  x_452 &  n_1542;
assign n_7307 = ~n_7305 & ~n_7306;
assign n_7308 = ~n_7304 &  n_7307;
assign n_7309 =  x_962 & ~n_7308;
assign n_7310 = ~x_962 &  n_7308;
assign n_7311 = ~n_7309 & ~n_7310;
assign n_7312 =  x_961 & ~n_6506;
assign n_7313 =  x_578 &  n_2414;
assign n_7314 =  x_451 &  n_1542;
assign n_7315 = ~n_7313 & ~n_7314;
assign n_7316 = ~n_7312 &  n_7315;
assign n_7317 =  x_961 & ~n_7316;
assign n_7318 = ~x_961 &  n_7316;
assign n_7319 = ~n_7317 & ~n_7318;
assign n_7320 =  x_960 & ~n_6506;
assign n_7321 =  x_577 &  n_2414;
assign n_7322 =  x_450 &  n_1542;
assign n_7323 = ~n_7321 & ~n_7322;
assign n_7324 = ~n_7320 &  n_7323;
assign n_7325 =  x_960 & ~n_7324;
assign n_7326 = ~x_960 &  n_7324;
assign n_7327 = ~n_7325 & ~n_7326;
assign n_7328 =  x_959 & ~n_6506;
assign n_7329 =  x_576 &  n_2414;
assign n_7330 =  x_449 &  n_1542;
assign n_7331 = ~n_7329 & ~n_7330;
assign n_7332 = ~n_7328 &  n_7331;
assign n_7333 =  x_959 & ~n_7332;
assign n_7334 = ~x_959 &  n_7332;
assign n_7335 = ~n_7333 & ~n_7334;
assign n_7336 =  x_958 & ~n_6506;
assign n_7337 =  x_575 &  n_2414;
assign n_7338 =  x_448 &  n_1542;
assign n_7339 = ~n_7337 & ~n_7338;
assign n_7340 = ~n_7336 &  n_7339;
assign n_7341 =  x_958 & ~n_7340;
assign n_7342 = ~x_958 &  n_7340;
assign n_7343 = ~n_7341 & ~n_7342;
assign n_7344 =  x_957 & ~n_6506;
assign n_7345 =  x_574 &  n_2414;
assign n_7346 =  x_447 &  n_1542;
assign n_7347 = ~n_7345 & ~n_7346;
assign n_7348 = ~n_7344 &  n_7347;
assign n_7349 =  x_957 & ~n_7348;
assign n_7350 = ~x_957 &  n_7348;
assign n_7351 = ~n_7349 & ~n_7350;
assign n_7352 =  x_956 & ~n_6506;
assign n_7353 =  x_573 &  n_2414;
assign n_7354 =  x_446 &  n_1542;
assign n_7355 = ~n_7353 & ~n_7354;
assign n_7356 = ~n_7352 &  n_7355;
assign n_7357 =  x_956 & ~n_7356;
assign n_7358 = ~x_956 &  n_7356;
assign n_7359 = ~n_7357 & ~n_7358;
assign n_7360 =  x_955 & ~n_6506;
assign n_7361 =  x_572 &  n_2414;
assign n_7362 =  x_445 &  n_1542;
assign n_7363 = ~n_7361 & ~n_7362;
assign n_7364 = ~n_7360 &  n_7363;
assign n_7365 =  x_955 & ~n_7364;
assign n_7366 = ~x_955 &  n_7364;
assign n_7367 = ~n_7365 & ~n_7366;
assign n_7368 =  x_954 & ~n_6506;
assign n_7369 =  x_571 &  n_2414;
assign n_7370 =  x_444 &  n_1542;
assign n_7371 = ~n_7369 & ~n_7370;
assign n_7372 = ~n_7368 &  n_7371;
assign n_7373 =  x_954 & ~n_7372;
assign n_7374 = ~x_954 &  n_7372;
assign n_7375 = ~n_7373 & ~n_7374;
assign n_7376 =  x_953 & ~n_6506;
assign n_7377 =  x_570 &  n_2414;
assign n_7378 =  x_443 &  n_1542;
assign n_7379 = ~n_7377 & ~n_7378;
assign n_7380 = ~n_7376 &  n_7379;
assign n_7381 =  x_953 & ~n_7380;
assign n_7382 = ~x_953 &  n_7380;
assign n_7383 = ~n_7381 & ~n_7382;
assign n_7384 =  x_952 & ~n_6506;
assign n_7385 =  x_569 &  n_2414;
assign n_7386 =  x_442 &  n_1542;
assign n_7387 = ~n_7385 & ~n_7386;
assign n_7388 = ~n_7384 &  n_7387;
assign n_7389 =  x_952 & ~n_7388;
assign n_7390 = ~x_952 &  n_7388;
assign n_7391 = ~n_7389 & ~n_7390;
assign n_7392 =  x_951 & ~n_6506;
assign n_7393 =  x_568 &  n_2414;
assign n_7394 =  x_441 &  n_1542;
assign n_7395 = ~n_7393 & ~n_7394;
assign n_7396 = ~n_7392 &  n_7395;
assign n_7397 =  x_951 & ~n_7396;
assign n_7398 = ~x_951 &  n_7396;
assign n_7399 = ~n_7397 & ~n_7398;
assign n_7400 =  x_950 & ~n_6506;
assign n_7401 =  x_567 &  n_2414;
assign n_7402 =  x_440 &  n_1542;
assign n_7403 = ~n_7401 & ~n_7402;
assign n_7404 = ~n_7400 &  n_7403;
assign n_7405 =  x_950 & ~n_7404;
assign n_7406 = ~x_950 &  n_7404;
assign n_7407 = ~n_7405 & ~n_7406;
assign n_7408 =  x_949 & ~n_6506;
assign n_7409 =  x_566 &  n_2414;
assign n_7410 =  x_439 &  n_1542;
assign n_7411 = ~n_7409 & ~n_7410;
assign n_7412 = ~n_7408 &  n_7411;
assign n_7413 =  x_949 & ~n_7412;
assign n_7414 = ~x_949 &  n_7412;
assign n_7415 = ~n_7413 & ~n_7414;
assign n_7416 =  x_948 & ~n_6506;
assign n_7417 =  x_565 &  n_2414;
assign n_7418 =  x_438 &  n_1542;
assign n_7419 = ~n_7417 & ~n_7418;
assign n_7420 = ~n_7416 &  n_7419;
assign n_7421 =  x_948 & ~n_7420;
assign n_7422 = ~x_948 &  n_7420;
assign n_7423 = ~n_7421 & ~n_7422;
assign n_7424 =  x_947 & ~n_6506;
assign n_7425 =  x_564 &  n_2414;
assign n_7426 =  x_437 &  n_1542;
assign n_7427 = ~n_7425 & ~n_7426;
assign n_7428 = ~n_7424 &  n_7427;
assign n_7429 =  x_947 & ~n_7428;
assign n_7430 = ~x_947 &  n_7428;
assign n_7431 = ~n_7429 & ~n_7430;
assign n_7432 =  x_946 & ~n_6506;
assign n_7433 =  x_563 &  n_2414;
assign n_7434 =  x_436 &  n_1542;
assign n_7435 = ~n_7433 & ~n_7434;
assign n_7436 = ~n_7432 &  n_7435;
assign n_7437 =  x_946 & ~n_7436;
assign n_7438 = ~x_946 &  n_7436;
assign n_7439 = ~n_7437 & ~n_7438;
assign n_7440 =  x_945 & ~n_6506;
assign n_7441 =  x_562 &  n_2414;
assign n_7442 =  x_435 &  n_1542;
assign n_7443 = ~n_7441 & ~n_7442;
assign n_7444 = ~n_7440 &  n_7443;
assign n_7445 =  x_945 & ~n_7444;
assign n_7446 = ~x_945 &  n_7444;
assign n_7447 = ~n_7445 & ~n_7446;
assign n_7448 =  x_944 & ~n_6506;
assign n_7449 =  x_561 &  n_2414;
assign n_7450 =  x_434 &  n_1542;
assign n_7451 = ~n_7449 & ~n_7450;
assign n_7452 = ~n_7448 &  n_7451;
assign n_7453 =  x_944 & ~n_7452;
assign n_7454 = ~x_944 &  n_7452;
assign n_7455 = ~n_7453 & ~n_7454;
assign n_7456 =  x_943 & ~n_6506;
assign n_7457 =  x_560 &  n_2414;
assign n_7458 =  x_433 &  n_1542;
assign n_7459 = ~n_7457 & ~n_7458;
assign n_7460 = ~n_7456 &  n_7459;
assign n_7461 =  x_943 & ~n_7460;
assign n_7462 = ~x_943 &  n_7460;
assign n_7463 = ~n_7461 & ~n_7462;
assign n_7464 =  x_942 & ~n_6506;
assign n_7465 =  x_559 &  n_2414;
assign n_7466 =  x_432 &  n_1542;
assign n_7467 = ~n_7465 & ~n_7466;
assign n_7468 = ~n_7464 &  n_7467;
assign n_7469 =  x_942 & ~n_7468;
assign n_7470 = ~x_942 &  n_7468;
assign n_7471 = ~n_7469 & ~n_7470;
assign n_7472 =  x_941 & ~n_6506;
assign n_7473 =  x_558 &  n_2414;
assign n_7474 =  x_431 &  n_1542;
assign n_7475 = ~n_7473 & ~n_7474;
assign n_7476 = ~n_7472 &  n_7475;
assign n_7477 =  x_941 & ~n_7476;
assign n_7478 = ~x_941 &  n_7476;
assign n_7479 = ~n_7477 & ~n_7478;
assign n_7480 =  x_940 & ~n_6506;
assign n_7481 =  x_557 &  n_2414;
assign n_7482 =  x_430 &  n_1542;
assign n_7483 = ~n_7481 & ~n_7482;
assign n_7484 = ~n_7480 &  n_7483;
assign n_7485 =  x_940 & ~n_7484;
assign n_7486 = ~x_940 &  n_7484;
assign n_7487 = ~n_7485 & ~n_7486;
assign n_7488 =  x_939 & ~n_6506;
assign n_7489 =  x_556 &  n_2414;
assign n_7490 =  x_429 &  n_1542;
assign n_7491 = ~n_7489 & ~n_7490;
assign n_7492 = ~n_7488 &  n_7491;
assign n_7493 =  x_939 & ~n_7492;
assign n_7494 = ~x_939 &  n_7492;
assign n_7495 = ~n_7493 & ~n_7494;
assign n_7496 =  x_938 & ~n_6506;
assign n_7497 =  x_555 &  n_2414;
assign n_7498 =  x_428 &  n_1542;
assign n_7499 = ~n_7497 & ~n_7498;
assign n_7500 = ~n_7496 &  n_7499;
assign n_7501 =  x_938 & ~n_7500;
assign n_7502 = ~x_938 &  n_7500;
assign n_7503 = ~n_7501 & ~n_7502;
assign n_7504 =  x_937 & ~n_6506;
assign n_7505 =  x_554 &  n_2414;
assign n_7506 =  x_427 &  n_1542;
assign n_7507 = ~n_7505 & ~n_7506;
assign n_7508 = ~n_7504 &  n_7507;
assign n_7509 =  x_937 & ~n_7508;
assign n_7510 = ~x_937 &  n_7508;
assign n_7511 = ~n_7509 & ~n_7510;
assign n_7512 =  x_936 & ~n_6506;
assign n_7513 =  x_553 &  n_2414;
assign n_7514 =  x_426 &  n_1542;
assign n_7515 = ~n_7513 & ~n_7514;
assign n_7516 = ~n_7512 &  n_7515;
assign n_7517 =  x_936 & ~n_7516;
assign n_7518 = ~x_936 &  n_7516;
assign n_7519 = ~n_7517 & ~n_7518;
assign n_7520 =  x_935 & ~n_6506;
assign n_7521 =  x_552 &  n_2414;
assign n_7522 =  x_425 &  n_1542;
assign n_7523 = ~n_7521 & ~n_7522;
assign n_7524 = ~n_7520 &  n_7523;
assign n_7525 =  x_935 & ~n_7524;
assign n_7526 = ~x_935 &  n_7524;
assign n_7527 = ~n_7525 & ~n_7526;
assign n_7528 =  x_902 &  n_1964;
assign n_7529 = ~n_1964 & ~n_1398;
assign n_7530 =  x_934 &  n_7529;
assign n_7531 = ~n_7528 & ~n_7530;
assign n_7532 =  x_934 & ~n_7531;
assign n_7533 = ~x_934 &  n_7531;
assign n_7534 = ~n_7532 & ~n_7533;
assign n_7535 =  x_901 &  n_1964;
assign n_7536 =  x_933 &  n_7529;
assign n_7537 = ~n_7535 & ~n_7536;
assign n_7538 =  x_933 & ~n_7537;
assign n_7539 = ~x_933 &  n_7537;
assign n_7540 = ~n_7538 & ~n_7539;
assign n_7541 =  x_900 &  n_1964;
assign n_7542 =  x_932 &  n_7529;
assign n_7543 = ~n_7541 & ~n_7542;
assign n_7544 =  x_932 & ~n_7543;
assign n_7545 = ~x_932 &  n_7543;
assign n_7546 = ~n_7544 & ~n_7545;
assign n_7547 =  x_931 &  n_7529;
assign n_7548 =  x_42 & ~x_899;
assign n_7549 =  n_2156 & ~n_7548;
assign n_7550 = ~n_7547 & ~n_7549;
assign n_7551 =  x_931 & ~n_7550;
assign n_7552 = ~x_931 &  n_7550;
assign n_7553 = ~n_7551 & ~n_7552;
assign n_7554 =  x_930 &  n_7529;
assign n_7555 =  x_42 & ~x_898;
assign n_7556 =  n_2156 & ~n_7555;
assign n_7557 = ~n_7554 & ~n_7556;
assign n_7558 =  x_930 & ~n_7557;
assign n_7559 = ~x_930 &  n_7557;
assign n_7560 = ~n_7558 & ~n_7559;
assign n_7561 =  x_897 &  n_1964;
assign n_7562 =  x_929 &  n_7529;
assign n_7563 = ~n_7561 & ~n_7562;
assign n_7564 =  x_929 & ~n_7563;
assign n_7565 = ~x_929 &  n_7563;
assign n_7566 = ~n_7564 & ~n_7565;
assign n_7567 =  x_896 &  n_1964;
assign n_7568 =  x_928 &  n_7529;
assign n_7569 = ~n_7567 & ~n_7568;
assign n_7570 =  x_928 & ~n_7569;
assign n_7571 = ~x_928 &  n_7569;
assign n_7572 = ~n_7570 & ~n_7571;
assign n_7573 =  x_895 &  n_1964;
assign n_7574 =  x_927 &  n_7529;
assign n_7575 = ~n_7573 & ~n_7574;
assign n_7576 =  x_927 & ~n_7575;
assign n_7577 = ~x_927 &  n_7575;
assign n_7578 = ~n_7576 & ~n_7577;
assign n_7579 =  x_894 &  n_1964;
assign n_7580 =  x_926 &  n_7529;
assign n_7581 = ~n_7579 & ~n_7580;
assign n_7582 =  x_926 & ~n_7581;
assign n_7583 = ~x_926 &  n_7581;
assign n_7584 = ~n_7582 & ~n_7583;
assign n_7585 =  x_893 &  n_1964;
assign n_7586 =  x_925 &  n_7529;
assign n_7587 = ~n_7585 & ~n_7586;
assign n_7588 =  x_925 & ~n_7587;
assign n_7589 = ~x_925 &  n_7587;
assign n_7590 = ~n_7588 & ~n_7589;
assign n_7591 =  x_924 &  n_7529;
assign n_7592 =  x_42 & ~x_892;
assign n_7593 =  n_2156 & ~n_7592;
assign n_7594 = ~n_7591 & ~n_7593;
assign n_7595 =  x_924 & ~n_7594;
assign n_7596 = ~x_924 &  n_7594;
assign n_7597 = ~n_7595 & ~n_7596;
assign n_7598 =  x_891 &  n_1964;
assign n_7599 =  x_923 &  n_7529;
assign n_7600 = ~n_7598 & ~n_7599;
assign n_7601 =  x_923 & ~n_7600;
assign n_7602 = ~x_923 &  n_7600;
assign n_7603 = ~n_7601 & ~n_7602;
assign n_7604 =  x_890 &  n_1964;
assign n_7605 =  x_922 &  n_7529;
assign n_7606 = ~n_7604 & ~n_7605;
assign n_7607 =  x_922 & ~n_7606;
assign n_7608 = ~x_922 &  n_7606;
assign n_7609 = ~n_7607 & ~n_7608;
assign n_7610 =  x_889 &  n_1964;
assign n_7611 =  x_921 &  n_7529;
assign n_7612 = ~n_7610 & ~n_7611;
assign n_7613 =  x_921 & ~n_7612;
assign n_7614 = ~x_921 &  n_7612;
assign n_7615 = ~n_7613 & ~n_7614;
assign n_7616 =  x_888 &  n_1964;
assign n_7617 =  x_920 &  n_7529;
assign n_7618 = ~n_7616 & ~n_7617;
assign n_7619 =  x_920 & ~n_7618;
assign n_7620 = ~x_920 &  n_7618;
assign n_7621 = ~n_7619 & ~n_7620;
assign n_7622 =  x_887 &  n_1964;
assign n_7623 =  x_919 &  n_7529;
assign n_7624 = ~n_7622 & ~n_7623;
assign n_7625 =  x_919 & ~n_7624;
assign n_7626 = ~x_919 &  n_7624;
assign n_7627 = ~n_7625 & ~n_7626;
assign n_7628 =  x_886 &  n_1964;
assign n_7629 =  x_918 &  n_7529;
assign n_7630 = ~n_7628 & ~n_7629;
assign n_7631 =  x_918 & ~n_7630;
assign n_7632 = ~x_918 &  n_7630;
assign n_7633 = ~n_7631 & ~n_7632;
assign n_7634 =  x_885 &  n_1964;
assign n_7635 =  x_917 &  n_7529;
assign n_7636 = ~n_7634 & ~n_7635;
assign n_7637 =  x_917 & ~n_7636;
assign n_7638 = ~x_917 &  n_7636;
assign n_7639 = ~n_7637 & ~n_7638;
assign n_7640 =  x_884 &  n_1964;
assign n_7641 =  x_916 &  n_7529;
assign n_7642 = ~n_7640 & ~n_7641;
assign n_7643 =  x_916 & ~n_7642;
assign n_7644 = ~x_916 &  n_7642;
assign n_7645 = ~n_7643 & ~n_7644;
assign n_7646 =  x_883 &  n_1964;
assign n_7647 =  x_915 &  n_7529;
assign n_7648 = ~n_7646 & ~n_7647;
assign n_7649 =  x_915 & ~n_7648;
assign n_7650 = ~x_915 &  n_7648;
assign n_7651 = ~n_7649 & ~n_7650;
assign n_7652 =  x_882 &  n_1964;
assign n_7653 =  x_914 &  n_7529;
assign n_7654 = ~n_7652 & ~n_7653;
assign n_7655 =  x_914 & ~n_7654;
assign n_7656 = ~x_914 &  n_7654;
assign n_7657 = ~n_7655 & ~n_7656;
assign n_7658 =  x_881 &  n_1964;
assign n_7659 =  x_913 &  n_7529;
assign n_7660 = ~n_7658 & ~n_7659;
assign n_7661 =  x_913 & ~n_7660;
assign n_7662 = ~x_913 &  n_7660;
assign n_7663 = ~n_7661 & ~n_7662;
assign n_7664 =  x_880 &  n_1964;
assign n_7665 =  x_912 &  n_7529;
assign n_7666 = ~n_7664 & ~n_7665;
assign n_7667 =  x_912 & ~n_7666;
assign n_7668 = ~x_912 &  n_7666;
assign n_7669 = ~n_7667 & ~n_7668;
assign n_7670 =  x_879 &  n_1964;
assign n_7671 =  x_911 &  n_7529;
assign n_7672 = ~n_7670 & ~n_7671;
assign n_7673 =  x_911 & ~n_7672;
assign n_7674 = ~x_911 &  n_7672;
assign n_7675 = ~n_7673 & ~n_7674;
assign n_7676 =  x_878 &  n_1964;
assign n_7677 =  x_910 &  n_7529;
assign n_7678 = ~n_7676 & ~n_7677;
assign n_7679 =  x_910 & ~n_7678;
assign n_7680 = ~x_910 &  n_7678;
assign n_7681 = ~n_7679 & ~n_7680;
assign n_7682 =  x_877 &  n_1964;
assign n_7683 =  x_909 &  n_7529;
assign n_7684 = ~n_7682 & ~n_7683;
assign n_7685 =  x_909 & ~n_7684;
assign n_7686 = ~x_909 &  n_7684;
assign n_7687 = ~n_7685 & ~n_7686;
assign n_7688 =  x_876 &  n_1964;
assign n_7689 =  x_908 &  n_7529;
assign n_7690 = ~n_7688 & ~n_7689;
assign n_7691 =  x_908 & ~n_7690;
assign n_7692 = ~x_908 &  n_7690;
assign n_7693 = ~n_7691 & ~n_7692;
assign n_7694 =  x_875 &  n_1964;
assign n_7695 =  x_907 &  n_7529;
assign n_7696 = ~n_7694 & ~n_7695;
assign n_7697 =  x_907 & ~n_7696;
assign n_7698 = ~x_907 &  n_7696;
assign n_7699 = ~n_7697 & ~n_7698;
assign n_7700 =  x_874 &  n_1964;
assign n_7701 =  x_906 &  n_7529;
assign n_7702 = ~n_7700 & ~n_7701;
assign n_7703 =  x_906 & ~n_7702;
assign n_7704 = ~x_906 &  n_7702;
assign n_7705 = ~n_7703 & ~n_7704;
assign n_7706 =  x_873 &  n_1964;
assign n_7707 =  x_905 &  n_7529;
assign n_7708 = ~n_7706 & ~n_7707;
assign n_7709 =  x_905 & ~n_7708;
assign n_7710 = ~x_905 &  n_7708;
assign n_7711 = ~n_7709 & ~n_7710;
assign n_7712 =  x_872 &  n_1964;
assign n_7713 =  x_904 &  n_7529;
assign n_7714 = ~n_7712 & ~n_7713;
assign n_7715 =  x_904 & ~n_7714;
assign n_7716 = ~x_904 &  n_7714;
assign n_7717 = ~n_7715 & ~n_7716;
assign n_7718 =  x_871 &  n_1964;
assign n_7719 =  x_903 &  n_7529;
assign n_7720 = ~n_7718 & ~n_7719;
assign n_7721 =  x_903 & ~n_7720;
assign n_7722 = ~x_903 &  n_7720;
assign n_7723 = ~n_7721 & ~n_7722;
assign n_7724 = ~x_38 &  n_1667;
assign n_7725 =  x_902 & ~n_7724;
assign n_7726 =  x_902 &  n_7725;
assign n_7727 = ~x_902 & ~n_7725;
assign n_7728 = ~n_7726 & ~n_7727;
assign n_7729 =  x_901 & ~n_7724;
assign n_7730 =  x_901 &  n_7729;
assign n_7731 = ~x_901 & ~n_7729;
assign n_7732 = ~n_7730 & ~n_7731;
assign n_7733 =  x_900 & ~n_7724;
assign n_7734 =  x_900 &  n_7733;
assign n_7735 = ~x_900 & ~n_7733;
assign n_7736 = ~n_7734 & ~n_7735;
assign n_7737 = ~x_41 &  n_1842;
assign n_7738 =  x_899 &  n_7737;
assign n_7739 = ~x_899 & ~n_7737;
assign n_7740 = ~n_7738 & ~n_7739;
assign n_7741 = ~n_7724 & ~n_7740;
assign n_7742 =  x_899 & ~n_7741;
assign n_7743 = ~x_899 &  n_7741;
assign n_7744 = ~n_7742 & ~n_7743;
assign n_7745 = ~x_898 &  n_7738;
assign n_7746 =  x_898 & ~n_7738;
assign n_7747 = ~n_7724 & ~n_7746;
assign n_7748 = ~n_7745 &  n_7747;
assign n_7749 =  x_898 & ~n_7748;
assign n_7750 = ~x_898 &  n_7748;
assign n_7751 = ~n_7749 & ~n_7750;
assign n_7752 = ~n_7737 & ~n_7724;
assign n_7753 =  x_897 &  n_7752;
assign n_7754 =  x_898 &  x_899;
assign n_7755 =  x_897 &  n_7754;
assign n_7756 = ~x_897 & ~n_7754;
assign n_7757 = ~n_7755 & ~n_7756;
assign n_7758 =  n_7737 &  n_7757;
assign n_7759 = ~n_7753 & ~n_7758;
assign n_7760 =  x_897 & ~n_7759;
assign n_7761 = ~x_897 &  n_7759;
assign n_7762 = ~n_7760 & ~n_7761;
assign n_7763 =  x_896 &  n_7752;
assign n_7764 =  x_896 &  n_7755;
assign n_7765 = ~x_896 & ~n_7755;
assign n_7766 = ~n_7764 & ~n_7765;
assign n_7767 =  n_7737 &  n_7766;
assign n_7768 = ~n_7763 & ~n_7767;
assign n_7769 =  x_896 & ~n_7768;
assign n_7770 = ~x_896 &  n_7768;
assign n_7771 = ~n_7769 & ~n_7770;
assign n_7772 =  x_895 &  n_7752;
assign n_7773 =  x_895 &  n_7764;
assign n_7774 = ~x_895 & ~n_7764;
assign n_7775 = ~n_7773 & ~n_7774;
assign n_7776 =  n_7737 &  n_7775;
assign n_7777 = ~n_7772 & ~n_7776;
assign n_7778 =  x_895 & ~n_7777;
assign n_7779 = ~x_895 &  n_7777;
assign n_7780 = ~n_7778 & ~n_7779;
assign n_7781 =  x_894 &  n_7752;
assign n_7782 =  x_894 &  n_7773;
assign n_7783 = ~x_894 & ~n_7773;
assign n_7784 = ~n_7782 & ~n_7783;
assign n_7785 =  n_7737 &  n_7784;
assign n_7786 = ~n_7781 & ~n_7785;
assign n_7787 =  x_894 & ~n_7786;
assign n_7788 = ~x_894 &  n_7786;
assign n_7789 = ~n_7787 & ~n_7788;
assign n_7790 =  x_893 &  n_7752;
assign n_7791 =  x_893 &  n_7782;
assign n_7792 = ~x_893 & ~n_7782;
assign n_7793 = ~n_7791 & ~n_7792;
assign n_7794 =  n_7737 &  n_7793;
assign n_7795 = ~n_7790 & ~n_7794;
assign n_7796 =  x_893 & ~n_7795;
assign n_7797 = ~x_893 &  n_7795;
assign n_7798 = ~n_7796 & ~n_7797;
assign n_7799 =  n_7791 &  n_7737;
assign n_7800 =  x_892 & ~n_7799;
assign n_7801 = ~x_892 &  n_7799;
assign n_7802 = ~n_7724 & ~n_7801;
assign n_7803 = ~n_7800 &  n_7802;
assign n_7804 =  x_892 & ~n_7803;
assign n_7805 = ~x_892 &  n_7803;
assign n_7806 = ~n_7804 & ~n_7805;
assign n_7807 =  x_891 &  n_7752;
assign n_7808 =  x_892 &  n_7791;
assign n_7809 = ~x_891 & ~n_7808;
assign n_7810 =  x_891 &  n_7808;
assign n_7811 = ~n_7810 &  n_7737;
assign n_7812 = ~n_7809 &  n_7811;
assign n_7813 = ~n_7807 & ~n_7812;
assign n_7814 =  x_891 & ~n_7813;
assign n_7815 = ~x_891 &  n_7813;
assign n_7816 = ~n_7814 & ~n_7815;
assign n_7817 =  x_890 &  n_7752;
assign n_7818 = ~x_890 & ~n_7810;
assign n_7819 =  x_890 &  n_7810;
assign n_7820 = ~n_7819 &  n_7737;
assign n_7821 = ~n_7818 &  n_7820;
assign n_7822 = ~n_7817 & ~n_7821;
assign n_7823 =  x_890 & ~n_7822;
assign n_7824 = ~x_890 &  n_7822;
assign n_7825 = ~n_7823 & ~n_7824;
assign n_7826 =  x_889 &  n_7752;
assign n_7827 = ~x_889 & ~n_7819;
assign n_7828 =  x_889 &  n_7819;
assign n_7829 = ~n_7828 &  n_7737;
assign n_7830 = ~n_7827 &  n_7829;
assign n_7831 = ~n_7826 & ~n_7830;
assign n_7832 =  x_889 & ~n_7831;
assign n_7833 = ~x_889 &  n_7831;
assign n_7834 = ~n_7832 & ~n_7833;
assign n_7835 =  x_888 &  n_7752;
assign n_7836 = ~x_888 & ~n_7828;
assign n_7837 =  x_888 &  n_7828;
assign n_7838 = ~n_7837 &  n_7737;
assign n_7839 = ~n_7836 &  n_7838;
assign n_7840 = ~n_7835 & ~n_7839;
assign n_7841 =  x_888 & ~n_7840;
assign n_7842 = ~x_888 &  n_7840;
assign n_7843 = ~n_7841 & ~n_7842;
assign n_7844 =  x_887 &  n_7752;
assign n_7845 = ~x_887 & ~n_7837;
assign n_7846 =  x_887 &  n_7837;
assign n_7847 = ~n_7846 &  n_7737;
assign n_7848 = ~n_7845 &  n_7847;
assign n_7849 = ~n_7844 & ~n_7848;
assign n_7850 =  x_887 & ~n_7849;
assign n_7851 = ~x_887 &  n_7849;
assign n_7852 = ~n_7850 & ~n_7851;
assign n_7853 =  x_886 &  n_7752;
assign n_7854 = ~x_886 & ~n_7846;
assign n_7855 =  x_886 &  n_7846;
assign n_7856 = ~n_7855 &  n_7737;
assign n_7857 = ~n_7854 &  n_7856;
assign n_7858 = ~n_7853 & ~n_7857;
assign n_7859 =  x_886 & ~n_7858;
assign n_7860 = ~x_886 &  n_7858;
assign n_7861 = ~n_7859 & ~n_7860;
assign n_7862 =  x_885 &  n_7752;
assign n_7863 = ~x_885 & ~n_7855;
assign n_7864 =  x_885 &  n_7855;
assign n_7865 = ~n_7864 &  n_7737;
assign n_7866 = ~n_7863 &  n_7865;
assign n_7867 = ~n_7862 & ~n_7866;
assign n_7868 =  x_885 & ~n_7867;
assign n_7869 = ~x_885 &  n_7867;
assign n_7870 = ~n_7868 & ~n_7869;
assign n_7871 =  x_884 &  n_7752;
assign n_7872 = ~x_884 & ~n_7864;
assign n_7873 =  x_884 &  n_7864;
assign n_7874 = ~n_7873 &  n_7737;
assign n_7875 = ~n_7872 &  n_7874;
assign n_7876 = ~n_7871 & ~n_7875;
assign n_7877 =  x_884 & ~n_7876;
assign n_7878 = ~x_884 &  n_7876;
assign n_7879 = ~n_7877 & ~n_7878;
assign n_7880 =  x_883 &  n_7752;
assign n_7881 = ~x_883 & ~n_7873;
assign n_7882 =  x_883 &  n_7873;
assign n_7883 = ~n_7882 &  n_7737;
assign n_7884 = ~n_7881 &  n_7883;
assign n_7885 = ~n_7880 & ~n_7884;
assign n_7886 =  x_883 & ~n_7885;
assign n_7887 = ~x_883 &  n_7885;
assign n_7888 = ~n_7886 & ~n_7887;
assign n_7889 =  x_882 &  n_7752;
assign n_7890 = ~x_882 & ~n_7882;
assign n_7891 =  x_882 &  n_7882;
assign n_7892 = ~n_7891 &  n_7737;
assign n_7893 = ~n_7890 &  n_7892;
assign n_7894 = ~n_7889 & ~n_7893;
assign n_7895 =  x_882 & ~n_7894;
assign n_7896 = ~x_882 &  n_7894;
assign n_7897 = ~n_7895 & ~n_7896;
assign n_7898 =  x_881 &  n_7752;
assign n_7899 = ~x_881 & ~n_7891;
assign n_7900 =  x_881 &  n_7891;
assign n_7901 = ~n_7900 &  n_7737;
assign n_7902 = ~n_7899 &  n_7901;
assign n_7903 = ~n_7898 & ~n_7902;
assign n_7904 =  x_881 & ~n_7903;
assign n_7905 = ~x_881 &  n_7903;
assign n_7906 = ~n_7904 & ~n_7905;
assign n_7907 =  x_880 &  n_7752;
assign n_7908 = ~x_880 & ~n_7900;
assign n_7909 =  x_880 &  n_7900;
assign n_7910 = ~n_7909 &  n_7737;
assign n_7911 = ~n_7908 &  n_7910;
assign n_7912 = ~n_7907 & ~n_7911;
assign n_7913 =  x_880 & ~n_7912;
assign n_7914 = ~x_880 &  n_7912;
assign n_7915 = ~n_7913 & ~n_7914;
assign n_7916 =  x_879 &  n_7752;
assign n_7917 = ~x_879 & ~n_7909;
assign n_7918 =  x_879 &  n_7909;
assign n_7919 = ~n_7918 &  n_7737;
assign n_7920 = ~n_7917 &  n_7919;
assign n_7921 = ~n_7916 & ~n_7920;
assign n_7922 =  x_879 & ~n_7921;
assign n_7923 = ~x_879 &  n_7921;
assign n_7924 = ~n_7922 & ~n_7923;
assign n_7925 =  x_878 &  n_7752;
assign n_7926 = ~x_878 & ~n_7918;
assign n_7927 =  x_878 &  n_7918;
assign n_7928 = ~n_7927 &  n_7737;
assign n_7929 = ~n_7926 &  n_7928;
assign n_7930 = ~n_7925 & ~n_7929;
assign n_7931 =  x_878 & ~n_7930;
assign n_7932 = ~x_878 &  n_7930;
assign n_7933 = ~n_7931 & ~n_7932;
assign n_7934 =  x_877 &  n_7752;
assign n_7935 = ~x_877 & ~n_7927;
assign n_7936 =  x_877 &  n_7927;
assign n_7937 = ~n_7936 &  n_7737;
assign n_7938 = ~n_7935 &  n_7937;
assign n_7939 = ~n_7934 & ~n_7938;
assign n_7940 =  x_877 & ~n_7939;
assign n_7941 = ~x_877 &  n_7939;
assign n_7942 = ~n_7940 & ~n_7941;
assign n_7943 =  x_876 &  n_7752;
assign n_7944 = ~x_876 & ~n_7936;
assign n_7945 =  x_876 &  n_7936;
assign n_7946 = ~n_7945 &  n_7737;
assign n_7947 = ~n_7944 &  n_7946;
assign n_7948 = ~n_7943 & ~n_7947;
assign n_7949 =  x_876 & ~n_7948;
assign n_7950 = ~x_876 &  n_7948;
assign n_7951 = ~n_7949 & ~n_7950;
assign n_7952 =  x_875 &  n_7752;
assign n_7953 = ~x_875 & ~n_7945;
assign n_7954 =  x_875 &  n_7945;
assign n_7955 = ~n_7954 &  n_7737;
assign n_7956 = ~n_7953 &  n_7955;
assign n_7957 = ~n_7952 & ~n_7956;
assign n_7958 =  x_875 & ~n_7957;
assign n_7959 = ~x_875 &  n_7957;
assign n_7960 = ~n_7958 & ~n_7959;
assign n_7961 =  x_874 &  n_7752;
assign n_7962 = ~x_874 & ~n_7954;
assign n_7963 =  x_874 &  n_7954;
assign n_7964 = ~n_7963 &  n_7737;
assign n_7965 = ~n_7962 &  n_7964;
assign n_7966 = ~n_7961 & ~n_7965;
assign n_7967 =  x_874 & ~n_7966;
assign n_7968 = ~x_874 &  n_7966;
assign n_7969 = ~n_7967 & ~n_7968;
assign n_7970 =  x_873 &  n_7752;
assign n_7971 = ~x_873 & ~n_7963;
assign n_7972 =  x_873 &  n_7963;
assign n_7973 = ~n_7972 &  n_7737;
assign n_7974 = ~n_7971 &  n_7973;
assign n_7975 = ~n_7970 & ~n_7974;
assign n_7976 =  x_873 & ~n_7975;
assign n_7977 = ~x_873 &  n_7975;
assign n_7978 = ~n_7976 & ~n_7977;
assign n_7979 =  x_872 &  n_7972;
assign n_7980 = ~n_7979 &  n_7737;
assign n_7981 = ~n_7980 & ~n_7752;
assign n_7982 =  x_872 & ~n_7981;
assign n_7983 =  n_7972 &  n_7980;
assign n_7984 = ~n_7982 & ~n_7983;
assign n_7985 =  x_872 & ~n_7984;
assign n_7986 = ~x_872 &  n_7984;
assign n_7987 = ~n_7985 & ~n_7986;
assign n_7988 =  x_871 & ~n_7981;
assign n_7989 = ~x_871 &  n_7737;
assign n_7990 =  n_7979 &  n_7989;
assign n_7991 = ~n_7988 & ~n_7990;
assign n_7992 =  x_871 & ~n_7991;
assign n_7993 = ~x_871 &  n_7991;
assign n_7994 = ~n_7992 & ~n_7993;
assign n_7995 = ~x_870 & ~n_1665;
assign n_7996 =  x_870 & ~n_7995;
assign n_7997 = ~x_870 &  n_7995;
assign n_7998 = ~n_7996 & ~n_7997;
assign n_7999 =  x_869 & ~n_1665;
assign n_8000 =  x_869 &  n_7999;
assign n_8001 = ~x_869 & ~n_7999;
assign n_8002 = ~n_8000 & ~n_8001;
assign n_8003 =  x_868 & ~n_1665;
assign n_8004 =  x_868 &  n_8003;
assign n_8005 = ~x_868 & ~n_8003;
assign n_8006 = ~n_8004 & ~n_8005;
assign n_8007 = ~x_867 & ~n_1668;
assign n_8008 = ~n_1665 & ~n_1668;
assign n_8009 =  x_867 & ~n_8008;
assign n_8010 = ~n_8007 & ~n_8009;
assign n_8011 =  x_867 &  n_8010;
assign n_8012 = ~x_867 & ~n_8010;
assign n_8013 = ~n_8011 & ~n_8012;
assign n_8014 =  x_866 &  n_8008;
assign n_8015 =  x_866 &  x_867;
assign n_8016 = ~x_866 & ~x_867;
assign n_8017 = ~n_8015 & ~n_8016;
assign n_8018 =  n_1668 &  n_8017;
assign n_8019 = ~n_8014 & ~n_8018;
assign n_8020 =  x_866 & ~n_8019;
assign n_8021 = ~x_866 &  n_8019;
assign n_8022 = ~n_8020 & ~n_8021;
assign n_8023 =  x_865 &  n_8008;
assign n_8024 =  x_865 &  n_8015;
assign n_8025 = ~x_865 & ~n_8015;
assign n_8026 = ~n_8024 & ~n_8025;
assign n_8027 =  n_1668 &  n_8026;
assign n_8028 = ~n_8023 & ~n_8027;
assign n_8029 =  x_865 & ~n_8028;
assign n_8030 = ~x_865 &  n_8028;
assign n_8031 = ~n_8029 & ~n_8030;
assign n_8032 =  x_864 &  n_8008;
assign n_8033 =  x_864 &  n_8024;
assign n_8034 = ~x_864 & ~n_8024;
assign n_8035 = ~n_8033 & ~n_8034;
assign n_8036 =  n_1668 &  n_8035;
assign n_8037 = ~n_8032 & ~n_8036;
assign n_8038 =  x_864 & ~n_8037;
assign n_8039 = ~x_864 &  n_8037;
assign n_8040 = ~n_8038 & ~n_8039;
assign n_8041 =  x_863 &  n_8008;
assign n_8042 = ~x_863 & ~n_8033;
assign n_8043 =  x_863 &  n_8033;
assign n_8044 =  n_1668 & ~n_8043;
assign n_8045 = ~n_8042 &  n_8044;
assign n_8046 = ~n_8041 & ~n_8045;
assign n_8047 =  x_863 & ~n_8046;
assign n_8048 = ~x_863 &  n_8046;
assign n_8049 = ~n_8047 & ~n_8048;
assign n_8050 =  x_862 &  n_8043;
assign n_8051 =  n_1668 & ~n_8050;
assign n_8052 = ~n_8008 & ~n_8051;
assign n_8053 =  x_862 & ~n_8052;
assign n_8054 =  n_8043 &  n_8051;
assign n_8055 = ~n_8053 & ~n_8054;
assign n_8056 =  x_862 & ~n_8055;
assign n_8057 = ~x_862 &  n_8055;
assign n_8058 = ~n_8056 & ~n_8057;
assign n_8059 =  n_1668 &  n_8050;
assign n_8060 = ~x_861 & ~n_8059;
assign n_8061 =  x_861 &  n_8052;
assign n_8062 = ~n_8060 & ~n_8061;
assign n_8063 =  x_861 &  n_8062;
assign n_8064 = ~x_861 & ~n_8062;
assign n_8065 = ~n_8063 & ~n_8064;
assign n_8066 =  x_861 &  n_8059;
assign n_8067 =  x_860 & ~n_8066;
assign n_8068 = ~x_860 &  n_8066;
assign n_8069 = ~n_1665 & ~n_8068;
assign n_8070 = ~n_8067 &  n_8069;
assign n_8071 =  x_860 & ~n_8070;
assign n_8072 = ~x_860 &  n_8070;
assign n_8073 = ~n_8071 & ~n_8072;
assign n_8074 =  x_859 &  n_8008;
assign n_8075 =  x_860 &  x_861;
assign n_8076 =  n_8050 &  n_8075;
assign n_8077 = ~x_859 & ~n_8076;
assign n_8078 =  x_859 &  n_8076;
assign n_8079 =  n_1668 & ~n_8078;
assign n_8080 = ~n_8077 &  n_8079;
assign n_8081 = ~n_8074 & ~n_8080;
assign n_8082 =  x_859 & ~n_8081;
assign n_8083 = ~x_859 &  n_8081;
assign n_8084 = ~n_8082 & ~n_8083;
assign n_8085 =  x_858 &  n_8008;
assign n_8086 = ~x_858 & ~n_8078;
assign n_8087 =  x_858 &  n_8078;
assign n_8088 =  n_1668 & ~n_8087;
assign n_8089 = ~n_8086 &  n_8088;
assign n_8090 = ~n_8085 & ~n_8089;
assign n_8091 =  x_858 & ~n_8090;
assign n_8092 = ~x_858 &  n_8090;
assign n_8093 = ~n_8091 & ~n_8092;
assign n_8094 =  x_857 &  n_8008;
assign n_8095 = ~x_857 & ~n_8087;
assign n_8096 =  x_857 &  n_8087;
assign n_8097 =  n_1668 & ~n_8096;
assign n_8098 = ~n_8095 &  n_8097;
assign n_8099 = ~n_8094 & ~n_8098;
assign n_8100 =  x_857 & ~n_8099;
assign n_8101 = ~x_857 &  n_8099;
assign n_8102 = ~n_8100 & ~n_8101;
assign n_8103 =  x_856 &  n_8008;
assign n_8104 = ~x_856 & ~n_8096;
assign n_8105 =  x_856 &  n_8096;
assign n_8106 =  n_1668 & ~n_8105;
assign n_8107 = ~n_8104 &  n_8106;
assign n_8108 = ~n_8103 & ~n_8107;
assign n_8109 =  x_856 & ~n_8108;
assign n_8110 = ~x_856 &  n_8108;
assign n_8111 = ~n_8109 & ~n_8110;
assign n_8112 =  x_855 &  n_8008;
assign n_8113 = ~x_855 & ~n_8105;
assign n_8114 =  x_855 &  n_8105;
assign n_8115 =  n_1668 & ~n_8114;
assign n_8116 = ~n_8113 &  n_8115;
assign n_8117 = ~n_8112 & ~n_8116;
assign n_8118 =  x_855 & ~n_8117;
assign n_8119 = ~x_855 &  n_8117;
assign n_8120 = ~n_8118 & ~n_8119;
assign n_8121 =  x_854 &  n_8008;
assign n_8122 = ~x_854 & ~n_8114;
assign n_8123 =  x_854 &  n_8114;
assign n_8124 =  n_1668 & ~n_8123;
assign n_8125 = ~n_8122 &  n_8124;
assign n_8126 = ~n_8121 & ~n_8125;
assign n_8127 =  x_854 & ~n_8126;
assign n_8128 = ~x_854 &  n_8126;
assign n_8129 = ~n_8127 & ~n_8128;
assign n_8130 =  x_853 &  n_8008;
assign n_8131 = ~x_853 & ~n_8123;
assign n_8132 =  x_853 &  n_8123;
assign n_8133 =  n_1668 & ~n_8132;
assign n_8134 = ~n_8131 &  n_8133;
assign n_8135 = ~n_8130 & ~n_8134;
assign n_8136 =  x_853 & ~n_8135;
assign n_8137 = ~x_853 &  n_8135;
assign n_8138 = ~n_8136 & ~n_8137;
assign n_8139 =  x_852 &  n_8008;
assign n_8140 = ~x_852 & ~n_8132;
assign n_8141 =  x_852 &  n_8132;
assign n_8142 =  n_1668 & ~n_8141;
assign n_8143 = ~n_8140 &  n_8142;
assign n_8144 = ~n_8139 & ~n_8143;
assign n_8145 =  x_852 & ~n_8144;
assign n_8146 = ~x_852 &  n_8144;
assign n_8147 = ~n_8145 & ~n_8146;
assign n_8148 =  x_851 &  n_8008;
assign n_8149 = ~x_851 & ~n_8141;
assign n_8150 =  x_851 &  n_8141;
assign n_8151 =  n_1668 & ~n_8150;
assign n_8152 = ~n_8149 &  n_8151;
assign n_8153 = ~n_8148 & ~n_8152;
assign n_8154 =  x_851 & ~n_8153;
assign n_8155 = ~x_851 &  n_8153;
assign n_8156 = ~n_8154 & ~n_8155;
assign n_8157 =  x_850 &  n_8008;
assign n_8158 = ~x_850 & ~n_8150;
assign n_8159 =  x_850 &  n_8150;
assign n_8160 =  n_1668 & ~n_8159;
assign n_8161 = ~n_8158 &  n_8160;
assign n_8162 = ~n_8157 & ~n_8161;
assign n_8163 =  x_850 & ~n_8162;
assign n_8164 = ~x_850 &  n_8162;
assign n_8165 = ~n_8163 & ~n_8164;
assign n_8166 =  x_849 &  n_8008;
assign n_8167 = ~x_849 & ~n_8159;
assign n_8168 =  x_849 &  n_8159;
assign n_8169 =  n_1668 & ~n_8168;
assign n_8170 = ~n_8167 &  n_8169;
assign n_8171 = ~n_8166 & ~n_8170;
assign n_8172 =  x_849 & ~n_8171;
assign n_8173 = ~x_849 &  n_8171;
assign n_8174 = ~n_8172 & ~n_8173;
assign n_8175 =  x_848 &  n_8008;
assign n_8176 = ~x_848 & ~n_8168;
assign n_8177 =  x_848 &  n_8168;
assign n_8178 =  n_1668 & ~n_8177;
assign n_8179 = ~n_8176 &  n_8178;
assign n_8180 = ~n_8175 & ~n_8179;
assign n_8181 =  x_848 & ~n_8180;
assign n_8182 = ~x_848 &  n_8180;
assign n_8183 = ~n_8181 & ~n_8182;
assign n_8184 =  x_847 &  n_8008;
assign n_8185 = ~x_847 & ~n_8177;
assign n_8186 =  x_847 &  n_8177;
assign n_8187 =  n_1668 & ~n_8186;
assign n_8188 = ~n_8185 &  n_8187;
assign n_8189 = ~n_8184 & ~n_8188;
assign n_8190 =  x_847 & ~n_8189;
assign n_8191 = ~x_847 &  n_8189;
assign n_8192 = ~n_8190 & ~n_8191;
assign n_8193 =  x_846 &  n_8008;
assign n_8194 = ~x_846 & ~n_8186;
assign n_8195 =  x_846 &  n_8186;
assign n_8196 =  n_1668 & ~n_8195;
assign n_8197 = ~n_8194 &  n_8196;
assign n_8198 = ~n_8193 & ~n_8197;
assign n_8199 =  x_846 & ~n_8198;
assign n_8200 = ~x_846 &  n_8198;
assign n_8201 = ~n_8199 & ~n_8200;
assign n_8202 =  x_845 &  n_8008;
assign n_8203 = ~x_845 & ~n_8195;
assign n_8204 =  x_845 &  n_8195;
assign n_8205 =  n_1668 & ~n_8204;
assign n_8206 = ~n_8203 &  n_8205;
assign n_8207 = ~n_8202 & ~n_8206;
assign n_8208 =  x_845 & ~n_8207;
assign n_8209 = ~x_845 &  n_8207;
assign n_8210 = ~n_8208 & ~n_8209;
assign n_8211 =  x_844 &  n_8008;
assign n_8212 = ~x_844 & ~n_8204;
assign n_8213 =  x_844 &  n_8204;
assign n_8214 =  n_1668 & ~n_8213;
assign n_8215 = ~n_8212 &  n_8214;
assign n_8216 = ~n_8211 & ~n_8215;
assign n_8217 =  x_844 & ~n_8216;
assign n_8218 = ~x_844 &  n_8216;
assign n_8219 = ~n_8217 & ~n_8218;
assign n_8220 =  x_843 &  n_8008;
assign n_8221 = ~x_843 & ~n_8213;
assign n_8222 =  x_843 &  n_8213;
assign n_8223 =  n_1668 & ~n_8222;
assign n_8224 = ~n_8221 &  n_8223;
assign n_8225 = ~n_8220 & ~n_8224;
assign n_8226 =  x_843 & ~n_8225;
assign n_8227 = ~x_843 &  n_8225;
assign n_8228 = ~n_8226 & ~n_8227;
assign n_8229 =  x_842 &  n_8008;
assign n_8230 = ~x_842 & ~n_8222;
assign n_8231 =  x_842 &  n_8222;
assign n_8232 =  n_1668 & ~n_8231;
assign n_8233 = ~n_8230 &  n_8232;
assign n_8234 = ~n_8229 & ~n_8233;
assign n_8235 =  x_842 & ~n_8234;
assign n_8236 = ~x_842 &  n_8234;
assign n_8237 = ~n_8235 & ~n_8236;
assign n_8238 =  x_841 &  n_8008;
assign n_8239 = ~x_841 & ~n_8231;
assign n_8240 =  x_841 &  n_8231;
assign n_8241 =  n_1668 & ~n_8240;
assign n_8242 = ~n_8239 &  n_8241;
assign n_8243 = ~n_8238 & ~n_8242;
assign n_8244 =  x_841 & ~n_8243;
assign n_8245 = ~x_841 &  n_8243;
assign n_8246 = ~n_8244 & ~n_8245;
assign n_8247 =  x_840 &  n_8240;
assign n_8248 =  n_1668 & ~n_8247;
assign n_8249 = ~n_8248 & ~n_8008;
assign n_8250 =  x_840 & ~n_8249;
assign n_8251 =  n_8240 &  n_8248;
assign n_8252 = ~n_8250 & ~n_8251;
assign n_8253 =  x_840 & ~n_8252;
assign n_8254 = ~x_840 &  n_8252;
assign n_8255 = ~n_8253 & ~n_8254;
assign n_8256 =  x_839 & ~n_8249;
assign n_8257 = ~x_839 &  n_1668;
assign n_8258 =  n_8247 &  n_8257;
assign n_8259 = ~n_8256 & ~n_8258;
assign n_8260 =  x_839 & ~n_8259;
assign n_8261 = ~x_839 &  n_8259;
assign n_8262 = ~n_8260 & ~n_8261;
assign n_8263 = ~n_752 & ~n_812;
assign n_8264 =  n_828 &  n_816;
assign n_8265 = ~n_8263 &  n_8264;
assign n_8266 =  x_807 & ~n_8265;
assign n_8267 =  n_828 &  n_817;
assign n_8268 =  x_487 &  n_8267;
assign n_8269 =  x_424 &  n_1230;
assign n_8270 = ~n_8268 & ~n_8269;
assign n_8271 = ~n_8266 &  n_8270;
assign n_8272 =  x_807 & ~n_8271;
assign n_8273 = ~x_807 &  n_8271;
assign n_8274 = ~n_8272 & ~n_8273;
assign n_8275 =  x_806 & ~n_8265;
assign n_8276 =  x_486 &  n_8267;
assign n_8277 =  x_423 &  n_1230;
assign n_8278 = ~n_8276 & ~n_8277;
assign n_8279 = ~n_8275 &  n_8278;
assign n_8280 =  x_806 & ~n_8279;
assign n_8281 = ~x_806 &  n_8279;
assign n_8282 = ~n_8280 & ~n_8281;
assign n_8283 =  x_805 & ~n_8265;
assign n_8284 =  x_485 &  n_8267;
assign n_8285 =  x_422 &  n_1230;
assign n_8286 = ~n_8284 & ~n_8285;
assign n_8287 = ~n_8283 &  n_8286;
assign n_8288 =  x_805 & ~n_8287;
assign n_8289 = ~x_805 &  n_8287;
assign n_8290 = ~n_8288 & ~n_8289;
assign n_8291 =  x_804 & ~n_8265;
assign n_8292 =  x_484 &  n_8267;
assign n_8293 =  x_421 &  n_1230;
assign n_8294 = ~n_8292 & ~n_8293;
assign n_8295 = ~n_8291 &  n_8294;
assign n_8296 =  x_804 & ~n_8295;
assign n_8297 = ~x_804 &  n_8295;
assign n_8298 = ~n_8296 & ~n_8297;
assign n_8299 =  x_803 & ~n_8265;
assign n_8300 =  x_483 &  n_8267;
assign n_8301 =  x_420 &  n_1230;
assign n_8302 = ~n_8300 & ~n_8301;
assign n_8303 = ~n_8299 &  n_8302;
assign n_8304 =  x_803 & ~n_8303;
assign n_8305 = ~x_803 &  n_8303;
assign n_8306 = ~n_8304 & ~n_8305;
assign n_8307 =  x_802 & ~n_8265;
assign n_8308 =  x_482 &  n_8267;
assign n_8309 =  x_419 &  n_1230;
assign n_8310 = ~n_8308 & ~n_8309;
assign n_8311 = ~n_8307 &  n_8310;
assign n_8312 =  x_802 & ~n_8311;
assign n_8313 = ~x_802 &  n_8311;
assign n_8314 = ~n_8312 & ~n_8313;
assign n_8315 =  x_801 & ~n_8265;
assign n_8316 =  x_481 &  n_8267;
assign n_8317 =  x_418 &  n_1230;
assign n_8318 = ~n_8316 & ~n_8317;
assign n_8319 = ~n_8315 &  n_8318;
assign n_8320 =  x_801 & ~n_8319;
assign n_8321 = ~x_801 &  n_8319;
assign n_8322 = ~n_8320 & ~n_8321;
assign n_8323 =  x_800 & ~n_8265;
assign n_8324 =  x_480 &  n_8267;
assign n_8325 =  x_417 &  n_1230;
assign n_8326 = ~n_8324 & ~n_8325;
assign n_8327 = ~n_8323 &  n_8326;
assign n_8328 =  x_800 & ~n_8327;
assign n_8329 = ~x_800 &  n_8327;
assign n_8330 = ~n_8328 & ~n_8329;
assign n_8331 =  x_799 & ~n_8265;
assign n_8332 =  x_479 &  n_8267;
assign n_8333 =  x_416 &  n_1230;
assign n_8334 = ~n_8332 & ~n_8333;
assign n_8335 = ~n_8331 &  n_8334;
assign n_8336 =  x_799 & ~n_8335;
assign n_8337 = ~x_799 &  n_8335;
assign n_8338 = ~n_8336 & ~n_8337;
assign n_8339 =  x_798 & ~n_8265;
assign n_8340 =  x_478 &  n_8267;
assign n_8341 =  x_415 &  n_1230;
assign n_8342 = ~n_8340 & ~n_8341;
assign n_8343 = ~n_8339 &  n_8342;
assign n_8344 =  x_798 & ~n_8343;
assign n_8345 = ~x_798 &  n_8343;
assign n_8346 = ~n_8344 & ~n_8345;
assign n_8347 =  x_797 & ~n_8265;
assign n_8348 =  x_477 &  n_8267;
assign n_8349 =  x_414 &  n_1230;
assign n_8350 = ~n_8348 & ~n_8349;
assign n_8351 = ~n_8347 &  n_8350;
assign n_8352 =  x_797 & ~n_8351;
assign n_8353 = ~x_797 &  n_8351;
assign n_8354 = ~n_8352 & ~n_8353;
assign n_8355 =  x_796 & ~n_8265;
assign n_8356 =  x_476 &  n_8267;
assign n_8357 =  x_413 &  n_1230;
assign n_8358 = ~n_8356 & ~n_8357;
assign n_8359 = ~n_8355 &  n_8358;
assign n_8360 =  x_796 & ~n_8359;
assign n_8361 = ~x_796 &  n_8359;
assign n_8362 = ~n_8360 & ~n_8361;
assign n_8363 =  x_795 & ~n_8265;
assign n_8364 =  x_475 &  n_8267;
assign n_8365 =  x_412 &  n_1230;
assign n_8366 = ~n_8364 & ~n_8365;
assign n_8367 = ~n_8363 &  n_8366;
assign n_8368 =  x_795 & ~n_8367;
assign n_8369 = ~x_795 &  n_8367;
assign n_8370 = ~n_8368 & ~n_8369;
assign n_8371 =  x_794 & ~n_8265;
assign n_8372 =  x_474 &  n_8267;
assign n_8373 =  x_411 &  n_1230;
assign n_8374 = ~n_8372 & ~n_8373;
assign n_8375 = ~n_8371 &  n_8374;
assign n_8376 =  x_794 & ~n_8375;
assign n_8377 = ~x_794 &  n_8375;
assign n_8378 = ~n_8376 & ~n_8377;
assign n_8379 =  x_793 & ~n_8265;
assign n_8380 =  x_473 &  n_8267;
assign n_8381 =  x_410 &  n_1230;
assign n_8382 = ~n_8380 & ~n_8381;
assign n_8383 = ~n_8379 &  n_8382;
assign n_8384 =  x_793 & ~n_8383;
assign n_8385 = ~x_793 &  n_8383;
assign n_8386 = ~n_8384 & ~n_8385;
assign n_8387 =  x_792 & ~n_8265;
assign n_8388 =  x_472 &  n_8267;
assign n_8389 =  x_409 &  n_1230;
assign n_8390 = ~n_8388 & ~n_8389;
assign n_8391 = ~n_8387 &  n_8390;
assign n_8392 =  x_792 & ~n_8391;
assign n_8393 = ~x_792 &  n_8391;
assign n_8394 = ~n_8392 & ~n_8393;
assign n_8395 =  x_791 & ~n_8265;
assign n_8396 =  x_471 &  n_8267;
assign n_8397 =  x_408 &  n_1230;
assign n_8398 = ~n_8396 & ~n_8397;
assign n_8399 = ~n_8395 &  n_8398;
assign n_8400 =  x_791 & ~n_8399;
assign n_8401 = ~x_791 &  n_8399;
assign n_8402 = ~n_8400 & ~n_8401;
assign n_8403 =  x_790 & ~n_8265;
assign n_8404 =  x_470 &  n_8267;
assign n_8405 =  x_407 &  n_1230;
assign n_8406 = ~n_8404 & ~n_8405;
assign n_8407 = ~n_8403 &  n_8406;
assign n_8408 =  x_790 & ~n_8407;
assign n_8409 = ~x_790 &  n_8407;
assign n_8410 = ~n_8408 & ~n_8409;
assign n_8411 =  x_789 & ~n_8265;
assign n_8412 =  x_469 &  n_8267;
assign n_8413 =  x_406 &  n_1230;
assign n_8414 = ~n_8412 & ~n_8413;
assign n_8415 = ~n_8411 &  n_8414;
assign n_8416 =  x_789 & ~n_8415;
assign n_8417 = ~x_789 &  n_8415;
assign n_8418 = ~n_8416 & ~n_8417;
assign n_8419 =  x_788 & ~n_8265;
assign n_8420 =  x_468 &  n_8267;
assign n_8421 =  x_405 &  n_1230;
assign n_8422 = ~n_8420 & ~n_8421;
assign n_8423 = ~n_8419 &  n_8422;
assign n_8424 =  x_788 & ~n_8423;
assign n_8425 = ~x_788 &  n_8423;
assign n_8426 = ~n_8424 & ~n_8425;
assign n_8427 =  x_787 & ~n_8265;
assign n_8428 =  x_467 &  n_8267;
assign n_8429 =  x_404 &  n_1230;
assign n_8430 = ~n_8428 & ~n_8429;
assign n_8431 = ~n_8427 &  n_8430;
assign n_8432 =  x_787 & ~n_8431;
assign n_8433 = ~x_787 &  n_8431;
assign n_8434 = ~n_8432 & ~n_8433;
assign n_8435 =  x_786 & ~n_8265;
assign n_8436 =  x_466 &  n_8267;
assign n_8437 =  x_403 &  n_1230;
assign n_8438 = ~n_8436 & ~n_8437;
assign n_8439 = ~n_8435 &  n_8438;
assign n_8440 =  x_786 & ~n_8439;
assign n_8441 = ~x_786 &  n_8439;
assign n_8442 = ~n_8440 & ~n_8441;
assign n_8443 =  x_785 & ~n_8265;
assign n_8444 =  x_465 &  n_8267;
assign n_8445 =  x_402 &  n_1230;
assign n_8446 = ~n_8444 & ~n_8445;
assign n_8447 = ~n_8443 &  n_8446;
assign n_8448 =  x_785 & ~n_8447;
assign n_8449 = ~x_785 &  n_8447;
assign n_8450 = ~n_8448 & ~n_8449;
assign n_8451 =  x_784 & ~n_8265;
assign n_8452 =  x_464 &  n_8267;
assign n_8453 =  x_401 &  n_1230;
assign n_8454 = ~n_8452 & ~n_8453;
assign n_8455 = ~n_8451 &  n_8454;
assign n_8456 =  x_784 & ~n_8455;
assign n_8457 = ~x_784 &  n_8455;
assign n_8458 = ~n_8456 & ~n_8457;
assign n_8459 =  x_783 & ~n_8265;
assign n_8460 =  x_463 &  n_8267;
assign n_8461 =  x_400 &  n_1230;
assign n_8462 = ~n_8460 & ~n_8461;
assign n_8463 = ~n_8459 &  n_8462;
assign n_8464 =  x_783 & ~n_8463;
assign n_8465 = ~x_783 &  n_8463;
assign n_8466 = ~n_8464 & ~n_8465;
assign n_8467 =  x_782 & ~n_8265;
assign n_8468 =  x_462 &  n_8267;
assign n_8469 =  x_399 &  n_1230;
assign n_8470 = ~n_8468 & ~n_8469;
assign n_8471 = ~n_8467 &  n_8470;
assign n_8472 =  x_782 & ~n_8471;
assign n_8473 = ~x_782 &  n_8471;
assign n_8474 = ~n_8472 & ~n_8473;
assign n_8475 =  x_781 & ~n_8265;
assign n_8476 =  x_461 &  n_8267;
assign n_8477 =  x_398 &  n_1230;
assign n_8478 = ~n_8476 & ~n_8477;
assign n_8479 = ~n_8475 &  n_8478;
assign n_8480 =  x_781 & ~n_8479;
assign n_8481 = ~x_781 &  n_8479;
assign n_8482 = ~n_8480 & ~n_8481;
assign n_8483 =  x_780 & ~n_8265;
assign n_8484 =  x_460 &  n_8267;
assign n_8485 =  x_397 &  n_1230;
assign n_8486 = ~n_8484 & ~n_8485;
assign n_8487 = ~n_8483 &  n_8486;
assign n_8488 =  x_780 & ~n_8487;
assign n_8489 = ~x_780 &  n_8487;
assign n_8490 = ~n_8488 & ~n_8489;
assign n_8491 =  x_779 & ~n_8265;
assign n_8492 =  x_459 &  n_8267;
assign n_8493 =  x_396 &  n_1230;
assign n_8494 = ~n_8492 & ~n_8493;
assign n_8495 = ~n_8491 &  n_8494;
assign n_8496 =  x_779 & ~n_8495;
assign n_8497 = ~x_779 &  n_8495;
assign n_8498 = ~n_8496 & ~n_8497;
assign n_8499 =  x_778 & ~n_8265;
assign n_8500 =  x_458 &  n_8267;
assign n_8501 =  x_395 &  n_1230;
assign n_8502 = ~n_8500 & ~n_8501;
assign n_8503 = ~n_8499 &  n_8502;
assign n_8504 =  x_778 & ~n_8503;
assign n_8505 = ~x_778 &  n_8503;
assign n_8506 = ~n_8504 & ~n_8505;
assign n_8507 =  x_777 & ~n_8265;
assign n_8508 =  x_457 &  n_8267;
assign n_8509 =  x_394 &  n_1230;
assign n_8510 = ~n_8508 & ~n_8509;
assign n_8511 = ~n_8507 &  n_8510;
assign n_8512 =  x_777 & ~n_8511;
assign n_8513 = ~x_777 &  n_8511;
assign n_8514 = ~n_8512 & ~n_8513;
assign n_8515 =  x_393 &  n_1230;
assign n_8516 =  x_776 & ~n_8265;
assign n_8517 = ~n_8515 & ~n_8516;
assign n_8518 =  x_776 & ~n_8517;
assign n_8519 = ~x_776 &  n_8517;
assign n_8520 = ~n_8518 & ~n_8519;
assign n_8521 =  x_775 & ~n_1531;
assign n_8522 =  i_32 &  n_1531;
assign n_8523 = ~n_8521 & ~n_8522;
assign n_8524 =  x_775 & ~n_8523;
assign n_8525 = ~x_775 &  n_8523;
assign n_8526 = ~n_8524 & ~n_8525;
assign n_8527 =  x_774 & ~n_1531;
assign n_8528 =  i_31 &  n_1531;
assign n_8529 = ~n_8527 & ~n_8528;
assign n_8530 =  x_774 & ~n_8529;
assign n_8531 = ~x_774 &  n_8529;
assign n_8532 = ~n_8530 & ~n_8531;
assign n_8533 =  x_773 & ~n_1531;
assign n_8534 =  i_30 &  n_1531;
assign n_8535 = ~n_8533 & ~n_8534;
assign n_8536 =  x_773 & ~n_8535;
assign n_8537 = ~x_773 &  n_8535;
assign n_8538 = ~n_8536 & ~n_8537;
assign n_8539 =  x_772 & ~n_1531;
assign n_8540 =  i_29 &  n_1531;
assign n_8541 = ~n_8539 & ~n_8540;
assign n_8542 =  x_772 & ~n_8541;
assign n_8543 = ~x_772 &  n_8541;
assign n_8544 = ~n_8542 & ~n_8543;
assign n_8545 =  x_771 & ~n_1531;
assign n_8546 =  i_28 &  n_1531;
assign n_8547 = ~n_8545 & ~n_8546;
assign n_8548 =  x_771 & ~n_8547;
assign n_8549 = ~x_771 &  n_8547;
assign n_8550 = ~n_8548 & ~n_8549;
assign n_8551 =  x_770 & ~n_1531;
assign n_8552 =  i_27 &  n_1531;
assign n_8553 = ~n_8551 & ~n_8552;
assign n_8554 =  x_770 & ~n_8553;
assign n_8555 = ~x_770 &  n_8553;
assign n_8556 = ~n_8554 & ~n_8555;
assign n_8557 =  x_769 & ~n_1531;
assign n_8558 =  i_26 &  n_1531;
assign n_8559 = ~n_8557 & ~n_8558;
assign n_8560 =  x_769 & ~n_8559;
assign n_8561 = ~x_769 &  n_8559;
assign n_8562 = ~n_8560 & ~n_8561;
assign n_8563 =  x_768 & ~n_1531;
assign n_8564 =  i_25 &  n_1531;
assign n_8565 = ~n_8563 & ~n_8564;
assign n_8566 =  x_768 & ~n_8565;
assign n_8567 = ~x_768 &  n_8565;
assign n_8568 = ~n_8566 & ~n_8567;
assign n_8569 =  x_767 & ~n_1531;
assign n_8570 =  i_24 &  n_1531;
assign n_8571 = ~n_8569 & ~n_8570;
assign n_8572 =  x_767 & ~n_8571;
assign n_8573 = ~x_767 &  n_8571;
assign n_8574 = ~n_8572 & ~n_8573;
assign n_8575 =  x_766 & ~n_1531;
assign n_8576 =  i_23 &  n_1531;
assign n_8577 = ~n_8575 & ~n_8576;
assign n_8578 =  x_766 & ~n_8577;
assign n_8579 = ~x_766 &  n_8577;
assign n_8580 = ~n_8578 & ~n_8579;
assign n_8581 =  x_765 & ~n_1531;
assign n_8582 =  i_22 &  n_1531;
assign n_8583 = ~n_8581 & ~n_8582;
assign n_8584 =  x_765 & ~n_8583;
assign n_8585 = ~x_765 &  n_8583;
assign n_8586 = ~n_8584 & ~n_8585;
assign n_8587 =  x_764 & ~n_1531;
assign n_8588 =  i_21 &  n_1531;
assign n_8589 = ~n_8587 & ~n_8588;
assign n_8590 =  x_764 & ~n_8589;
assign n_8591 = ~x_764 &  n_8589;
assign n_8592 = ~n_8590 & ~n_8591;
assign n_8593 =  x_763 & ~n_1531;
assign n_8594 =  i_20 &  n_1531;
assign n_8595 = ~n_8593 & ~n_8594;
assign n_8596 =  x_763 & ~n_8595;
assign n_8597 = ~x_763 &  n_8595;
assign n_8598 = ~n_8596 & ~n_8597;
assign n_8599 =  x_762 & ~n_1531;
assign n_8600 =  i_19 &  n_1531;
assign n_8601 = ~n_8599 & ~n_8600;
assign n_8602 =  x_762 & ~n_8601;
assign n_8603 = ~x_762 &  n_8601;
assign n_8604 = ~n_8602 & ~n_8603;
assign n_8605 =  x_761 & ~n_1531;
assign n_8606 =  i_18 &  n_1531;
assign n_8607 = ~n_8605 & ~n_8606;
assign n_8608 =  x_761 & ~n_8607;
assign n_8609 = ~x_761 &  n_8607;
assign n_8610 = ~n_8608 & ~n_8609;
assign n_8611 =  x_760 & ~n_1531;
assign n_8612 =  i_17 &  n_1531;
assign n_8613 = ~n_8611 & ~n_8612;
assign n_8614 =  x_760 & ~n_8613;
assign n_8615 = ~x_760 &  n_8613;
assign n_8616 = ~n_8614 & ~n_8615;
assign n_8617 =  x_759 & ~n_1531;
assign n_8618 =  i_16 &  n_1531;
assign n_8619 = ~n_8617 & ~n_8618;
assign n_8620 =  x_759 & ~n_8619;
assign n_8621 = ~x_759 &  n_8619;
assign n_8622 = ~n_8620 & ~n_8621;
assign n_8623 =  x_758 & ~n_1531;
assign n_8624 =  i_15 &  n_1531;
assign n_8625 = ~n_8623 & ~n_8624;
assign n_8626 =  x_758 & ~n_8625;
assign n_8627 = ~x_758 &  n_8625;
assign n_8628 = ~n_8626 & ~n_8627;
assign n_8629 =  x_757 & ~n_1531;
assign n_8630 =  i_14 &  n_1531;
assign n_8631 = ~n_8629 & ~n_8630;
assign n_8632 =  x_757 & ~n_8631;
assign n_8633 = ~x_757 &  n_8631;
assign n_8634 = ~n_8632 & ~n_8633;
assign n_8635 =  x_756 & ~n_1531;
assign n_8636 =  i_13 &  n_1531;
assign n_8637 = ~n_8635 & ~n_8636;
assign n_8638 =  x_756 & ~n_8637;
assign n_8639 = ~x_756 &  n_8637;
assign n_8640 = ~n_8638 & ~n_8639;
assign n_8641 =  x_755 & ~n_1531;
assign n_8642 =  i_12 &  n_1531;
assign n_8643 = ~n_8641 & ~n_8642;
assign n_8644 =  x_755 & ~n_8643;
assign n_8645 = ~x_755 &  n_8643;
assign n_8646 = ~n_8644 & ~n_8645;
assign n_8647 =  x_754 & ~n_1531;
assign n_8648 =  i_11 &  n_1531;
assign n_8649 = ~n_8647 & ~n_8648;
assign n_8650 =  x_754 & ~n_8649;
assign n_8651 = ~x_754 &  n_8649;
assign n_8652 = ~n_8650 & ~n_8651;
assign n_8653 =  x_753 & ~n_1531;
assign n_8654 =  i_10 &  n_1531;
assign n_8655 = ~n_8653 & ~n_8654;
assign n_8656 =  x_753 & ~n_8655;
assign n_8657 = ~x_753 &  n_8655;
assign n_8658 = ~n_8656 & ~n_8657;
assign n_8659 =  x_752 & ~n_1531;
assign n_8660 =  i_9 &  n_1531;
assign n_8661 = ~n_8659 & ~n_8660;
assign n_8662 =  x_752 & ~n_8661;
assign n_8663 = ~x_752 &  n_8661;
assign n_8664 = ~n_8662 & ~n_8663;
assign n_8665 =  x_751 & ~n_1531;
assign n_8666 =  i_8 &  n_1531;
assign n_8667 = ~n_8665 & ~n_8666;
assign n_8668 =  x_751 & ~n_8667;
assign n_8669 = ~x_751 &  n_8667;
assign n_8670 = ~n_8668 & ~n_8669;
assign n_8671 =  x_750 & ~n_1531;
assign n_8672 =  i_7 &  n_1531;
assign n_8673 = ~n_8671 & ~n_8672;
assign n_8674 =  x_750 & ~n_8673;
assign n_8675 = ~x_750 &  n_8673;
assign n_8676 = ~n_8674 & ~n_8675;
assign n_8677 =  x_748 & ~n_1531;
assign n_8678 =  i_5 &  n_1531;
assign n_8679 = ~n_8677 & ~n_8678;
assign n_8680 =  x_748 & ~n_8679;
assign n_8681 = ~x_748 &  n_8679;
assign n_8682 = ~n_8680 & ~n_8681;
assign n_8683 =  x_749 & ~n_1531;
assign n_8684 =  i_6 &  n_1531;
assign n_8685 = ~n_8683 & ~n_8684;
assign n_8686 =  x_749 & ~n_8685;
assign n_8687 = ~x_749 &  n_8685;
assign n_8688 = ~n_8686 & ~n_8687;
assign n_8689 = ~n_8682 & ~n_8688;
assign n_8690 = ~n_8676 &  n_8689;
assign n_8691 = ~n_8670 &  n_8690;
assign n_8692 = ~n_8664 &  n_8691;
assign n_8693 = ~n_8658 &  n_8692;
assign n_8694 = ~n_8652 &  n_8693;
assign n_8695 = ~n_8646 &  n_8694;
assign n_8696 = ~n_8640 &  n_8695;
assign n_8697 = ~n_8634 &  n_8696;
assign n_8698 = ~n_8628 &  n_8697;
assign n_8699 = ~n_8622 &  n_8698;
assign n_8700 = ~n_8616 &  n_8699;
assign n_8701 = ~n_8610 &  n_8700;
assign n_8702 = ~n_8604 &  n_8701;
assign n_8703 = ~n_8598 &  n_8702;
assign n_8704 = ~n_8592 &  n_8703;
assign n_8705 = ~n_8586 &  n_8704;
assign n_8706 = ~n_8580 &  n_8705;
assign n_8707 = ~n_8574 &  n_8706;
assign n_8708 = ~n_8568 &  n_8707;
assign n_8709 = ~n_8562 &  n_8708;
assign n_8710 = ~n_8556 &  n_8709;
assign n_8711 = ~n_8550 &  n_8710;
assign n_8712 = ~n_8544 &  n_8711;
assign n_8713 = ~n_8538 &  n_8712;
assign n_8714 = ~n_8532 &  n_8713;
assign n_8715 = ~n_8526 &  n_8714;
assign n_8716 = ~n_8520 &  n_8715;
assign n_8717 = ~n_8514 &  n_8716;
assign n_8718 = ~n_8506 &  n_8717;
assign n_8719 = ~n_8498 &  n_8718;
assign n_8720 = ~n_8490 &  n_8719;
assign n_8721 = ~n_8482 &  n_8720;
assign n_8722 = ~n_8474 &  n_8721;
assign n_8723 = ~n_8466 &  n_8722;
assign n_8724 = ~n_8458 &  n_8723;
assign n_8725 = ~n_8450 &  n_8724;
assign n_8726 = ~n_8442 &  n_8725;
assign n_8727 = ~n_8434 &  n_8726;
assign n_8728 = ~n_8426 &  n_8727;
assign n_8729 = ~n_8418 &  n_8728;
assign n_8730 = ~n_8410 &  n_8729;
assign n_8731 = ~n_8402 &  n_8730;
assign n_8732 = ~n_8394 &  n_8731;
assign n_8733 = ~n_8386 &  n_8732;
assign n_8734 = ~n_8378 &  n_8733;
assign n_8735 = ~n_8370 &  n_8734;
assign n_8736 = ~n_8362 &  n_8735;
assign n_8737 = ~n_8354 &  n_8736;
assign n_8738 = ~n_8346 &  n_8737;
assign n_8739 = ~n_8338 &  n_8738;
assign n_8740 = ~n_8330 &  n_8739;
assign n_8741 = ~n_8322 &  n_8740;
assign n_8742 = ~n_8314 &  n_8741;
assign n_8743 = ~n_8306 &  n_8742;
assign n_8744 = ~n_8298 &  n_8743;
assign n_8745 = ~n_8290 &  n_8744;
assign n_8746 = ~n_8282 &  n_8745;
assign n_8747 = ~n_8274 &  n_8746;
assign n_8748 = ~n_8262 &  n_8747;
assign n_8749 = ~n_8255 &  n_8748;
assign n_8750 = ~n_8246 &  n_8749;
assign n_8751 = ~n_8237 &  n_8750;
assign n_8752 = ~n_8228 &  n_8751;
assign n_8753 = ~n_8219 &  n_8752;
assign n_8754 = ~n_8210 &  n_8753;
assign n_8755 = ~n_8201 &  n_8754;
assign n_8756 = ~n_8192 &  n_8755;
assign n_8757 = ~n_8183 &  n_8756;
assign n_8758 = ~n_8174 &  n_8757;
assign n_8759 = ~n_8165 &  n_8758;
assign n_8760 = ~n_8156 &  n_8759;
assign n_8761 = ~n_8147 &  n_8760;
assign n_8762 = ~n_8138 &  n_8761;
assign n_8763 = ~n_8129 &  n_8762;
assign n_8764 = ~n_8120 &  n_8763;
assign n_8765 = ~n_8111 &  n_8764;
assign n_8766 = ~n_8102 &  n_8765;
assign n_8767 = ~n_8093 &  n_8766;
assign n_8768 = ~n_8084 &  n_8767;
assign n_8769 = ~n_8073 &  n_8768;
assign n_8770 = ~n_8065 &  n_8769;
assign n_8771 = ~n_8058 &  n_8770;
assign n_8772 = ~n_8049 &  n_8771;
assign n_8773 = ~n_8040 &  n_8772;
assign n_8774 = ~n_8031 &  n_8773;
assign n_8775 = ~n_8022 &  n_8774;
assign n_8776 = ~n_8013 &  n_8775;
assign n_8777 = ~n_8006 &  n_8776;
assign n_8778 = ~n_8002 &  n_8777;
assign n_8779 = ~n_7998 &  n_8778;
assign n_8780 = ~n_7994 &  n_8779;
assign n_8781 = ~n_7987 &  n_8780;
assign n_8782 = ~n_7978 &  n_8781;
assign n_8783 = ~n_7969 &  n_8782;
assign n_8784 = ~n_7960 &  n_8783;
assign n_8785 = ~n_7951 &  n_8784;
assign n_8786 = ~n_7942 &  n_8785;
assign n_8787 = ~n_7933 &  n_8786;
assign n_8788 = ~n_7924 &  n_8787;
assign n_8789 = ~n_7915 &  n_8788;
assign n_8790 = ~n_7906 &  n_8789;
assign n_8791 = ~n_7897 &  n_8790;
assign n_8792 = ~n_7888 &  n_8791;
assign n_8793 = ~n_7879 &  n_8792;
assign n_8794 = ~n_7870 &  n_8793;
assign n_8795 = ~n_7861 &  n_8794;
assign n_8796 = ~n_7852 &  n_8795;
assign n_8797 = ~n_7843 &  n_8796;
assign n_8798 = ~n_7834 &  n_8797;
assign n_8799 = ~n_7825 &  n_8798;
assign n_8800 = ~n_7816 &  n_8799;
assign n_8801 = ~n_7806 &  n_8800;
assign n_8802 = ~n_7798 &  n_8801;
assign n_8803 = ~n_7789 &  n_8802;
assign n_8804 = ~n_7780 &  n_8803;
assign n_8805 = ~n_7771 &  n_8804;
assign n_8806 = ~n_7762 &  n_8805;
assign n_8807 = ~n_7751 &  n_8806;
assign n_8808 = ~n_7744 &  n_8807;
assign n_8809 = ~n_7736 &  n_8808;
assign n_8810 = ~n_7732 &  n_8809;
assign n_8811 = ~n_7728 &  n_8810;
assign n_8812 = ~n_7723 &  n_8811;
assign n_8813 = ~n_7717 &  n_8812;
assign n_8814 = ~n_7711 &  n_8813;
assign n_8815 = ~n_7705 &  n_8814;
assign n_8816 = ~n_7699 &  n_8815;
assign n_8817 = ~n_7693 &  n_8816;
assign n_8818 = ~n_7687 &  n_8817;
assign n_8819 = ~n_7681 &  n_8818;
assign n_8820 = ~n_7675 &  n_8819;
assign n_8821 = ~n_7669 &  n_8820;
assign n_8822 = ~n_7663 &  n_8821;
assign n_8823 = ~n_7657 &  n_8822;
assign n_8824 = ~n_7651 &  n_8823;
assign n_8825 = ~n_7645 &  n_8824;
assign n_8826 = ~n_7639 &  n_8825;
assign n_8827 = ~n_7633 &  n_8826;
assign n_8828 = ~n_7627 &  n_8827;
assign n_8829 = ~n_7621 &  n_8828;
assign n_8830 = ~n_7615 &  n_8829;
assign n_8831 = ~n_7609 &  n_8830;
assign n_8832 = ~n_7603 &  n_8831;
assign n_8833 = ~n_7597 &  n_8832;
assign n_8834 = ~n_7590 &  n_8833;
assign n_8835 = ~n_7584 &  n_8834;
assign n_8836 = ~n_7578 &  n_8835;
assign n_8837 = ~n_7572 &  n_8836;
assign n_8838 = ~n_7566 &  n_8837;
assign n_8839 = ~n_7560 &  n_8838;
assign n_8840 = ~n_7553 &  n_8839;
assign n_8841 = ~n_7546 &  n_8840;
assign n_8842 = ~n_7540 &  n_8841;
assign n_8843 = ~n_7534 &  n_8842;
assign n_8844 = ~n_7527 &  n_8843;
assign n_8845 = ~n_7519 &  n_8844;
assign n_8846 = ~n_7511 &  n_8845;
assign n_8847 = ~n_7503 &  n_8846;
assign n_8848 = ~n_7495 &  n_8847;
assign n_8849 = ~n_7487 &  n_8848;
assign n_8850 = ~n_7479 &  n_8849;
assign n_8851 = ~n_7471 &  n_8850;
assign n_8852 = ~n_7463 &  n_8851;
assign n_8853 = ~n_7455 &  n_8852;
assign n_8854 = ~n_7447 &  n_8853;
assign n_8855 = ~n_7439 &  n_8854;
assign n_8856 = ~n_7431 &  n_8855;
assign n_8857 = ~n_7423 &  n_8856;
assign n_8858 = ~n_7415 &  n_8857;
assign n_8859 = ~n_7407 &  n_8858;
assign n_8860 = ~n_7399 &  n_8859;
assign n_8861 = ~n_7391 &  n_8860;
assign n_8862 = ~n_7383 &  n_8861;
assign n_8863 = ~n_7375 &  n_8862;
assign n_8864 = ~n_7367 &  n_8863;
assign n_8865 = ~n_7359 &  n_8864;
assign n_8866 = ~n_7351 &  n_8865;
assign n_8867 = ~n_7343 &  n_8866;
assign n_8868 = ~n_7335 &  n_8867;
assign n_8869 = ~n_7327 &  n_8868;
assign n_8870 = ~n_7319 &  n_8869;
assign n_8871 = ~n_7311 &  n_8870;
assign n_8872 = ~n_7303 &  n_8871;
assign n_8873 = ~n_7295 &  n_8872;
assign n_8874 = ~n_7287 &  n_8873;
assign n_8875 = ~n_7279 &  n_8874;
assign n_8876 = ~n_7271 &  n_8875;
assign n_8877 = ~n_7266 &  n_8876;
assign n_8878 = ~n_7261 &  n_8877;
assign n_8879 = ~n_7256 &  n_8878;
assign n_8880 = ~n_7251 &  n_8879;
assign n_8881 = ~n_7246 &  n_8880;
assign n_8882 = ~n_7241 &  n_8881;
assign n_8883 = ~n_7236 &  n_8882;
assign n_8884 = ~n_7231 &  n_8883;
assign n_8885 = ~n_7226 &  n_8884;
assign n_8886 = ~n_7220 &  n_8885;
assign n_8887 = ~n_7214 &  n_8886;
assign n_8888 = ~n_7208 &  n_8887;
assign n_8889 = ~n_7202 &  n_8888;
assign n_8890 = ~n_7196 &  n_8889;
assign n_8891 = ~n_7190 &  n_8890;
assign n_8892 = ~n_7184 &  n_8891;
assign n_8893 = ~n_7178 &  n_8892;
assign n_8894 = ~n_7173 &  n_8893;
assign n_8895 = ~n_7168 &  n_8894;
assign n_8896 = ~n_7163 &  n_8895;
assign n_8897 = ~n_7158 &  n_8896;
assign n_8898 = ~n_7153 &  n_8897;
assign n_8899 = ~n_7148 &  n_8898;
assign n_8900 = ~n_7143 &  n_8899;
assign n_8901 = ~n_7138 &  n_8900;
assign n_8902 = ~n_7133 &  n_8901;
assign n_8903 = ~n_7128 &  n_8902;
assign n_8904 = ~n_7123 &  n_8903;
assign n_8905 = ~n_7118 &  n_8904;
assign n_8906 = ~n_7113 &  n_8905;
assign n_8907 = ~n_7108 &  n_8906;
assign n_8908 = ~n_7103 &  n_8907;
assign n_8909 = ~n_7098 &  n_8908;
assign n_8910 = ~n_7093 &  n_8909;
assign n_8911 = ~n_7088 &  n_8910;
assign n_8912 = ~n_7083 &  n_8911;
assign n_8913 = ~n_7078 &  n_8912;
assign n_8914 = ~n_7073 &  n_8913;
assign n_8915 = ~n_7068 &  n_8914;
assign n_8916 = ~n_7063 &  n_8915;
assign n_8917 = ~n_7058 &  n_8916;
assign n_8918 = ~n_7053 &  n_8917;
assign n_8919 = ~n_7048 &  n_8918;
assign n_8920 = ~n_7043 &  n_8919;
assign n_8921 = ~n_7038 &  n_8920;
assign n_8922 = ~n_7033 &  n_8921;
assign n_8923 = ~n_7028 &  n_8922;
assign n_8924 = ~n_7023 &  n_8923;
assign n_8925 = ~n_7018 &  n_8924;
assign n_8926 = ~n_7010 &  n_8925;
assign n_8927 = ~n_7002 &  n_8926;
assign n_8928 = ~n_6994 &  n_8927;
assign n_8929 = ~n_6986 &  n_8928;
assign n_8930 = ~n_6978 &  n_8929;
assign n_8931 = ~n_6970 &  n_8930;
assign n_8932 = ~n_6962 &  n_8931;
assign n_8933 = ~n_6954 &  n_8932;
assign n_8934 = ~n_6946 &  n_8933;
assign n_8935 = ~n_6938 &  n_8934;
assign n_8936 = ~n_6930 &  n_8935;
assign n_8937 = ~n_6922 &  n_8936;
assign n_8938 = ~n_6914 &  n_8937;
assign n_8939 = ~n_6906 &  n_8938;
assign n_8940 = ~n_6898 &  n_8939;
assign n_8941 = ~n_6890 &  n_8940;
assign n_8942 = ~n_6882 &  n_8941;
assign n_8943 = ~n_6874 &  n_8942;
assign n_8944 = ~n_6866 &  n_8943;
assign n_8945 = ~n_6858 &  n_8944;
assign n_8946 = ~n_6850 &  n_8945;
assign n_8947 = ~n_6842 &  n_8946;
assign n_8948 = ~n_6834 &  n_8947;
assign n_8949 = ~n_6826 &  n_8948;
assign n_8950 = ~n_6818 &  n_8949;
assign n_8951 = ~n_6810 &  n_8950;
assign n_8952 = ~n_6802 &  n_8951;
assign n_8953 = ~n_6794 &  n_8952;
assign n_8954 = ~n_6786 &  n_8953;
assign n_8955 = ~n_6778 &  n_8954;
assign n_8956 = ~n_6770 &  n_8955;
assign n_8957 = ~n_6762 &  n_8956;
assign n_8958 = ~n_6754 &  n_8957;
assign n_8959 = ~n_6746 &  n_8958;
assign n_8960 = ~n_6738 &  n_8959;
assign n_8961 = ~n_6730 &  n_8960;
assign n_8962 = ~n_6722 &  n_8961;
assign n_8963 = ~n_6714 &  n_8962;
assign n_8964 = ~n_6706 &  n_8963;
assign n_8965 = ~n_6698 &  n_8964;
assign n_8966 = ~n_6690 &  n_8965;
assign n_8967 = ~n_6682 &  n_8966;
assign n_8968 = ~n_6674 &  n_8967;
assign n_8969 = ~n_6666 &  n_8968;
assign n_8970 = ~n_6658 &  n_8969;
assign n_8971 = ~n_6650 &  n_8970;
assign n_8972 = ~n_6642 &  n_8971;
assign n_8973 = ~n_6634 &  n_8972;
assign n_8974 = ~n_6626 &  n_8973;
assign n_8975 = ~n_6618 &  n_8974;
assign n_8976 = ~n_6610 &  n_8975;
assign n_8977 = ~n_6602 &  n_8976;
assign n_8978 = ~n_6594 &  n_8977;
assign n_8979 = ~n_6586 &  n_8978;
assign n_8980 = ~n_6578 &  n_8979;
assign n_8981 = ~n_6570 &  n_8980;
assign n_8982 = ~n_6562 &  n_8981;
assign n_8983 = ~n_6554 &  n_8982;
assign n_8984 = ~n_6546 &  n_8983;
assign n_8985 = ~n_6538 &  n_8984;
assign n_8986 = ~n_6530 &  n_8985;
assign n_8987 = ~n_6522 &  n_8986;
assign n_8988 = ~n_6514 &  n_8987;
assign n_8989 = ~n_6500 &  n_8988;
assign n_8990 = ~n_6494 &  n_8989;
assign n_8991 = ~n_6488 &  n_8990;
assign n_8992 = ~n_6482 &  n_8991;
assign n_8993 = ~n_6476 &  n_8992;
assign n_8994 = ~n_6470 &  n_8993;
assign n_8995 = ~n_6464 &  n_8994;
assign n_8996 = ~n_6458 &  n_8995;
assign n_8997 = ~n_6452 &  n_8996;
assign n_8998 = ~n_6446 &  n_8997;
assign n_8999 = ~n_6440 &  n_8998;
assign n_9000 = ~n_6434 &  n_8999;
assign n_9001 = ~n_6428 &  n_9000;
assign n_9002 = ~n_6422 &  n_9001;
assign n_9003 = ~n_6416 &  n_9002;
assign n_9004 = ~n_6410 &  n_9003;
assign n_9005 = ~n_6404 &  n_9004;
assign n_9006 = ~n_6398 &  n_9005;
assign n_9007 = ~n_6392 &  n_9006;
assign n_9008 = ~n_6386 &  n_9007;
assign n_9009 = ~n_6380 &  n_9008;
assign n_9010 = ~n_6374 &  n_9009;
assign n_9011 = ~n_6368 &  n_9010;
assign n_9012 = ~n_6362 &  n_9011;
assign n_9013 = ~n_6356 &  n_9012;
assign n_9014 = ~n_6350 &  n_9013;
assign n_9015 = ~n_6344 &  n_9014;
assign n_9016 = ~n_6338 &  n_9015;
assign n_9017 = ~n_6332 &  n_9016;
assign n_9018 = ~n_6326 &  n_9017;
assign n_9019 = ~n_6320 &  n_9018;
assign n_9020 = ~n_6314 &  n_9019;
assign n_9021 = ~n_6308 &  n_9020;
assign n_9022 = ~n_6302 &  n_9021;
assign n_9023 = ~n_6296 &  n_9022;
assign n_9024 = ~n_6290 &  n_9023;
assign n_9025 = ~n_6284 &  n_9024;
assign n_9026 = ~n_6278 &  n_9025;
assign n_9027 = ~n_6272 &  n_9026;
assign n_9028 = ~n_6266 &  n_9027;
assign n_9029 = ~n_6260 &  n_9028;
assign n_9030 = ~n_6254 &  n_9029;
assign n_9031 = ~n_6248 &  n_9030;
assign n_9032 = ~n_6242 &  n_9031;
assign n_9033 = ~n_6236 &  n_9032;
assign n_9034 = ~n_6230 &  n_9033;
assign n_9035 = ~n_6224 &  n_9034;
assign n_9036 = ~n_6218 &  n_9035;
assign n_9037 = ~n_6212 &  n_9036;
assign n_9038 = ~n_6206 &  n_9037;
assign n_9039 = ~n_6200 &  n_9038;
assign n_9040 = ~n_6194 &  n_9039;
assign n_9041 = ~n_6188 &  n_9040;
assign n_9042 = ~n_6182 &  n_9041;
assign n_9043 = ~n_6176 &  n_9042;
assign n_9044 = ~n_6170 &  n_9043;
assign n_9045 = ~n_6164 &  n_9044;
assign n_9046 = ~n_6158 &  n_9045;
assign n_9047 = ~n_6152 &  n_9046;
assign n_9048 = ~n_6146 &  n_9047;
assign n_9049 = ~n_6140 &  n_9048;
assign n_9050 = ~n_6134 &  n_9049;
assign n_9051 = ~n_6128 &  n_9050;
assign n_9052 = ~n_6122 &  n_9051;
assign n_9053 = ~n_6116 &  n_9052;
assign n_9054 = ~n_6110 &  n_9053;
assign n_9055 = ~n_6104 &  n_9054;
assign n_9056 = ~n_6098 &  n_9055;
assign n_9057 = ~n_6092 &  n_9056;
assign n_9058 = ~n_6086 &  n_9057;
assign n_9059 = ~n_6080 &  n_9058;
assign n_9060 = ~n_6074 &  n_9059;
assign n_9061 = ~n_6068 &  n_9060;
assign n_9062 = ~n_6062 &  n_9061;
assign n_9063 = ~n_6056 &  n_9062;
assign n_9064 = ~n_6050 &  n_9063;
assign n_9065 = ~n_6044 &  n_9064;
assign n_9066 = ~n_6038 &  n_9065;
assign n_9067 = ~n_6032 &  n_9066;
assign n_9068 = ~n_6026 &  n_9067;
assign n_9069 = ~n_6020 &  n_9068;
assign n_9070 = ~n_6014 &  n_9069;
assign n_9071 = ~n_6008 &  n_9070;
assign n_9072 = ~n_6002 &  n_9071;
assign n_9073 = ~n_5996 &  n_9072;
assign n_9074 = ~n_5990 &  n_9073;
assign n_9075 = ~n_5983 &  n_9074;
assign n_9076 = ~n_5977 &  n_9075;
assign n_9077 = ~n_5971 &  n_9076;
assign n_9078 = ~n_5965 &  n_9077;
assign n_9079 = ~n_5959 &  n_9078;
assign n_9080 = ~n_5953 &  n_9079;
assign n_9081 = ~n_5947 &  n_9080;
assign n_9082 = ~n_5940 &  n_9081;
assign n_9083 = ~n_5934 &  n_9082;
assign n_9084 = ~n_5927 &  n_9083;
assign n_9085 = ~n_5919 &  n_9084;
assign n_9086 = ~n_5913 &  n_9085;
assign n_9087 = ~n_5905 &  n_9086;
assign n_9088 = ~n_5897 &  n_9087;
assign n_9089 = ~n_5889 &  n_9088;
assign n_9090 = ~n_5881 &  n_9089;
assign n_9091 = ~n_5873 &  n_9090;
assign n_9092 = ~n_5865 &  n_9091;
assign n_9093 = ~n_5857 &  n_9092;
assign n_9094 = ~n_5849 &  n_9093;
assign n_9095 = ~n_5841 &  n_9094;
assign n_9096 = ~n_5833 &  n_9095;
assign n_9097 = ~n_5825 &  n_9096;
assign n_9098 = ~n_5817 &  n_9097;
assign n_9099 = ~n_5809 &  n_9098;
assign n_9100 = ~n_5801 &  n_9099;
assign n_9101 = ~n_5793 &  n_9100;
assign n_9102 = ~n_5785 &  n_9101;
assign n_9103 = ~n_5777 &  n_9102;
assign n_9104 = ~n_5769 &  n_9103;
assign n_9105 = ~n_5761 &  n_9104;
assign n_9106 = ~n_5753 &  n_9105;
assign n_9107 = ~n_5745 &  n_9106;
assign n_9108 = ~n_5737 &  n_9107;
assign n_9109 = ~n_5729 &  n_9108;
assign n_9110 = ~n_5721 &  n_9109;
assign n_9111 = ~n_5713 &  n_9110;
assign n_9112 = ~n_5705 &  n_9111;
assign n_9113 = ~n_5697 &  n_9112;
assign n_9114 = ~n_5689 &  n_9113;
assign n_9115 = ~n_5681 &  n_9114;
assign n_9116 = ~n_5673 &  n_9115;
assign n_9117 = ~n_5663 &  n_9116;
assign n_9118 = ~n_5657 &  n_9117;
assign n_9119 = ~n_5651 &  n_9118;
assign n_9120 = ~n_5645 &  n_9119;
assign n_9121 = ~n_5639 &  n_9120;
assign n_9122 = ~n_5633 &  n_9121;
assign n_9123 = ~n_5627 &  n_9122;
assign n_9124 = ~n_5621 &  n_9123;
assign n_9125 = ~n_5615 &  n_9124;
assign n_9126 = ~n_5609 &  n_9125;
assign n_9127 = ~n_5603 &  n_9126;
assign n_9128 = ~n_5597 &  n_9127;
assign n_9129 = ~n_5591 &  n_9128;
assign n_9130 = ~n_5585 &  n_9129;
assign n_9131 = ~n_5579 &  n_9130;
assign n_9132 = ~n_5573 &  n_9131;
assign n_9133 = ~n_5567 &  n_9132;
assign n_9134 = ~n_5561 &  n_9133;
assign n_9135 = ~n_5555 &  n_9134;
assign n_9136 = ~n_5549 &  n_9135;
assign n_9137 = ~n_5543 &  n_9136;
assign n_9138 = ~n_5537 &  n_9137;
assign n_9139 = ~n_5530 &  n_9138;
assign n_9140 = ~n_5524 &  n_9139;
assign n_9141 = ~n_5518 &  n_9140;
assign n_9142 = ~n_5512 &  n_9141;
assign n_9143 = ~n_5506 &  n_9142;
assign n_9144 = ~n_5500 &  n_9143;
assign n_9145 = ~n_5494 &  n_9144;
assign n_9146 = ~n_5488 &  n_9145;
assign n_9147 = ~n_5482 &  n_9146;
assign n_9148 = ~n_5476 &  n_9147;
assign n_9149 = ~n_5467 &  n_9148;
assign n_9150 = ~n_5463 &  n_9149;
assign n_9151 = ~n_5457 &  n_9150;
assign n_9152 = ~n_5451 &  n_9151;
assign n_9153 = ~n_5445 &  n_9152;
assign n_9154 = ~n_5439 &  n_9153;
assign n_9155 = ~n_5433 &  n_9154;
assign n_9156 = ~n_5427 &  n_9155;
assign n_9157 = ~n_5421 &  n_9156;
assign n_9158 = ~n_5415 &  n_9157;
assign n_9159 = ~n_5409 &  n_9158;
assign n_9160 = ~n_5403 &  n_9159;
assign n_9161 = ~n_5397 &  n_9160;
assign n_9162 = ~n_5391 &  n_9161;
assign n_9163 = ~n_5385 &  n_9162;
assign n_9164 = ~n_5379 &  n_9163;
assign n_9165 = ~n_5373 &  n_9164;
assign n_9166 = ~n_5367 &  n_9165;
assign n_9167 = ~n_5361 &  n_9166;
assign n_9168 = ~n_5355 &  n_9167;
assign n_9169 = ~n_5349 &  n_9168;
assign n_9170 = ~n_5343 &  n_9169;
assign n_9171 = ~n_5337 &  n_9170;
assign n_9172 = ~n_5331 &  n_9171;
assign n_9173 = ~n_5325 &  n_9172;
assign n_9174 = ~n_5319 &  n_9173;
assign n_9175 = ~n_5313 &  n_9174;
assign n_9176 = ~n_5307 &  n_9175;
assign n_9177 = ~n_5301 &  n_9176;
assign n_9178 = ~n_5295 &  n_9177;
assign n_9179 = ~n_5289 &  n_9178;
assign n_9180 = ~n_5283 &  n_9179;
assign n_9181 = ~n_5277 &  n_9180;
assign n_9182 = ~n_5271 &  n_9181;
assign n_9183 = ~n_5265 &  n_9182;
assign n_9184 = ~n_5259 &  n_9183;
assign n_9185 = ~n_5253 &  n_9184;
assign n_9186 = ~n_5247 &  n_9185;
assign n_9187 = ~n_5241 &  n_9186;
assign n_9188 = ~n_5235 &  n_9187;
assign n_9189 = ~n_5229 &  n_9188;
assign n_9190 = ~n_5223 &  n_9189;
assign n_9191 = ~n_5217 &  n_9190;
assign n_9192 = ~n_5211 &  n_9191;
assign n_9193 = ~n_5205 &  n_9192;
assign n_9194 = ~n_5199 &  n_9193;
assign n_9195 = ~n_5193 &  n_9194;
assign n_9196 = ~n_5187 &  n_9195;
assign n_9197 = ~n_5181 &  n_9196;
assign n_9198 = ~n_5175 &  n_9197;
assign n_9199 = ~n_5169 &  n_9198;
assign n_9200 = ~n_5163 &  n_9199;
assign n_9201 = ~n_5157 &  n_9200;
assign n_9202 = ~n_5151 &  n_9201;
assign n_9203 = ~n_5145 &  n_9202;
assign n_9204 = ~n_5139 &  n_9203;
assign n_9205 = ~n_5133 &  n_9204;
assign n_9206 = ~n_5127 &  n_9205;
assign n_9207 = ~n_5121 &  n_9206;
assign n_9208 = ~n_5115 &  n_9207;
assign n_9209 = ~n_5109 &  n_9208;
assign n_9210 = ~n_5103 &  n_9209;
assign n_9211 = ~n_5097 &  n_9210;
assign n_9212 = ~n_5091 &  n_9211;
assign n_9213 = ~n_5085 &  n_9212;
assign n_9214 = ~n_5079 &  n_9213;
assign n_9215 = ~n_5073 &  n_9214;
assign n_9216 = ~n_5067 &  n_9215;
assign n_9217 = ~n_5061 &  n_9216;
assign n_9218 = ~n_5055 &  n_9217;
assign n_9219 = ~n_5049 &  n_9218;
assign n_9220 = ~n_5043 &  n_9219;
assign n_9221 = ~n_5037 &  n_9220;
assign n_9222 = ~n_5031 &  n_9221;
assign n_9223 = ~n_5025 &  n_9222;
assign n_9224 = ~n_5019 &  n_9223;
assign n_9225 = ~n_5013 &  n_9224;
assign n_9226 = ~n_5007 &  n_9225;
assign n_9227 = ~n_5001 &  n_9226;
assign n_9228 = ~n_4995 &  n_9227;
assign n_9229 = ~n_4989 &  n_9228;
assign n_9230 = ~n_4983 &  n_9229;
assign n_9231 = ~n_4977 &  n_9230;
assign n_9232 = ~n_4971 &  n_9231;
assign n_9233 = ~n_4965 &  n_9232;
assign n_9234 = ~n_4959 &  n_9233;
assign n_9235 = ~n_4953 &  n_9234;
assign n_9236 = ~n_4947 &  n_9235;
assign n_9237 = ~n_4941 &  n_9236;
assign n_9238 = ~n_4935 &  n_9237;
assign n_9239 = ~n_4929 &  n_9238;
assign n_9240 = ~n_4923 &  n_9239;
assign n_9241 = ~n_4917 &  n_9240;
assign n_9242 = ~n_4911 &  n_9241;
assign n_9243 = ~n_4905 &  n_9242;
assign n_9244 = ~n_4899 &  n_9243;
assign n_9245 = ~n_4892 &  n_9244;
assign n_9246 = ~n_4886 &  n_9245;
assign n_9247 = ~n_4880 &  n_9246;
assign n_9248 = ~n_4874 &  n_9247;
assign n_9249 = ~n_4868 &  n_9248;
assign n_9250 = ~n_4862 &  n_9249;
assign n_9251 = ~n_4856 &  n_9250;
assign n_9252 = ~n_4850 &  n_9251;
assign n_9253 = ~n_4844 &  n_9252;
assign n_9254 = ~n_4838 &  n_9253;
assign n_9255 = ~n_4832 &  n_9254;
assign n_9256 = ~n_4826 &  n_9255;
assign n_9257 = ~n_4820 &  n_9256;
assign n_9258 = ~n_4814 &  n_9257;
assign n_9259 = ~n_4808 &  n_9258;
assign n_9260 = ~n_4802 &  n_9259;
assign n_9261 = ~n_4796 &  n_9260;
assign n_9262 = ~n_4790 &  n_9261;
assign n_9263 = ~n_4784 &  n_9262;
assign n_9264 = ~n_4778 &  n_9263;
assign n_9265 = ~n_4772 &  n_9264;
assign n_9266 = ~n_4766 &  n_9265;
assign n_9267 = ~n_4760 &  n_9266;
assign n_9268 = ~n_4754 &  n_9267;
assign n_9269 = ~n_4748 &  n_9268;
assign n_9270 = ~n_4742 &  n_9269;
assign n_9271 = ~n_4736 &  n_9270;
assign n_9272 = ~n_4730 &  n_9271;
assign n_9273 = ~n_4724 &  n_9272;
assign n_9274 = ~n_4718 &  n_9273;
assign n_9275 = ~n_4712 &  n_9274;
assign n_9276 = ~n_4706 &  n_9275;
assign n_9277 = ~n_4700 &  n_9276;
assign n_9278 = ~n_4694 &  n_9277;
assign n_9279 = ~n_4688 &  n_9278;
assign n_9280 = ~n_4682 &  n_9279;
assign n_9281 = ~n_4676 &  n_9280;
assign n_9282 = ~n_4670 &  n_9281;
assign n_9283 = ~n_4664 &  n_9282;
assign n_9284 = ~n_4658 &  n_9283;
assign n_9285 = ~n_4652 &  n_9284;
assign n_9286 = ~n_4646 &  n_9285;
assign n_9287 = ~n_4640 &  n_9286;
assign n_9288 = ~n_4634 &  n_9287;
assign n_9289 = ~n_4628 &  n_9288;
assign n_9290 = ~n_4622 &  n_9289;
assign n_9291 = ~n_4616 &  n_9290;
assign n_9292 = ~n_4610 &  n_9291;
assign n_9293 = ~n_4604 &  n_9292;
assign n_9294 = ~n_4598 &  n_9293;
assign n_9295 = ~n_4592 &  n_9294;
assign n_9296 = ~n_4586 &  n_9295;
assign n_9297 = ~n_4580 &  n_9296;
assign n_9298 = ~n_4574 &  n_9297;
assign n_9299 = ~n_4568 &  n_9298;
assign n_9300 = ~n_4562 &  n_9299;
assign n_9301 = ~n_4556 &  n_9300;
assign n_9302 = ~n_4550 &  n_9301;
assign n_9303 = ~n_4544 &  n_9302;
assign n_9304 = ~n_4538 &  n_9303;
assign n_9305 = ~n_4532 &  n_9304;
assign n_9306 = ~n_4526 &  n_9305;
assign n_9307 = ~n_4520 &  n_9306;
assign n_9308 = ~n_4514 &  n_9307;
assign n_9309 = ~n_4508 &  n_9308;
assign n_9310 = ~n_4502 &  n_9309;
assign n_9311 = ~n_4496 &  n_9310;
assign n_9312 = ~n_4490 &  n_9311;
assign n_9313 = ~n_4484 &  n_9312;
assign n_9314 = ~n_4478 &  n_9313;
assign n_9315 = ~n_4472 &  n_9314;
assign n_9316 = ~n_4466 &  n_9315;
assign n_9317 = ~n_4460 &  n_9316;
assign n_9318 = ~n_4454 &  n_9317;
assign n_9319 = ~n_4448 &  n_9318;
assign n_9320 = ~n_4442 &  n_9319;
assign n_9321 = ~n_4436 &  n_9320;
assign n_9322 = ~n_4430 &  n_9321;
assign n_9323 = ~n_4424 &  n_9322;
assign n_9324 = ~n_4418 &  n_9323;
assign n_9325 = ~n_4412 &  n_9324;
assign n_9326 = ~n_4406 &  n_9325;
assign n_9327 = ~n_4400 &  n_9326;
assign n_9328 = ~n_4394 &  n_9327;
assign n_9329 = ~n_4388 &  n_9328;
assign n_9330 = ~n_4382 &  n_9329;
assign n_9331 = ~n_4376 &  n_9330;
assign n_9332 = ~n_4370 &  n_9331;
assign n_9333 = ~n_4364 &  n_9332;
assign n_9334 = ~n_4358 &  n_9333;
assign n_9335 = ~n_4352 &  n_9334;
assign n_9336 = ~n_4346 &  n_9335;
assign n_9337 = ~n_4340 &  n_9336;
assign n_9338 = ~n_4334 &  n_9337;
assign n_9339 = ~n_4328 &  n_9338;
assign n_9340 = ~n_4322 &  n_9339;
assign n_9341 = ~n_4316 &  n_9340;
assign n_9342 = ~n_4310 &  n_9341;
assign n_9343 = ~n_4304 &  n_9342;
assign n_9344 = ~n_4298 &  n_9343;
assign n_9345 = ~n_4292 &  n_9344;
assign n_9346 = ~n_4286 &  n_9345;
assign n_9347 = ~n_4280 &  n_9346;
assign n_9348 = ~n_4274 &  n_9347;
assign n_9349 = ~n_4268 &  n_9348;
assign n_9350 = ~n_4262 &  n_9349;
assign n_9351 = ~n_4256 &  n_9350;
assign n_9352 = ~n_4250 &  n_9351;
assign n_9353 = ~n_4244 &  n_9352;
assign n_9354 = ~n_4238 &  n_9353;
assign n_9355 = ~n_4232 &  n_9354;
assign n_9356 = ~n_4226 &  n_9355;
assign n_9357 = ~n_4220 &  n_9356;
assign n_9358 = ~n_4214 &  n_9357;
assign n_9359 = ~n_4208 &  n_9358;
assign n_9360 = ~n_4202 &  n_9359;
assign n_9361 = ~n_4196 &  n_9360;
assign n_9362 = ~n_4190 &  n_9361;
assign n_9363 = ~n_4184 &  n_9362;
assign n_9364 = ~n_4178 &  n_9363;
assign n_9365 = ~n_4172 &  n_9364;
assign n_9366 = ~n_4166 &  n_9365;
assign n_9367 = ~n_4160 &  n_9366;
assign n_9368 = ~n_4154 &  n_9367;
assign n_9369 = ~n_4148 &  n_9368;
assign n_9370 = ~n_4142 &  n_9369;
assign n_9371 = ~n_4136 &  n_9370;
assign n_9372 = ~n_4130 &  n_9371;
assign n_9373 = ~n_4124 &  n_9372;
assign n_9374 = ~n_4118 &  n_9373;
assign n_9375 = ~n_4112 &  n_9374;
assign n_9376 = ~n_4106 &  n_9375;
assign n_9377 = ~n_4100 &  n_9376;
assign n_9378 = ~n_4094 &  n_9377;
assign n_9379 = ~n_4088 &  n_9378;
assign n_9380 = ~n_4082 &  n_9379;
assign n_9381 = ~n_4076 &  n_9380;
assign n_9382 = ~n_4070 &  n_9381;
assign n_9383 = ~n_4064 &  n_9382;
assign n_9384 = ~n_4058 &  n_9383;
assign n_9385 = ~n_4052 &  n_9384;
assign n_9386 = ~n_4046 &  n_9385;
assign n_9387 = ~n_4040 &  n_9386;
assign n_9388 = ~n_4034 &  n_9387;
assign n_9389 = ~n_4028 &  n_9388;
assign n_9390 = ~n_4022 &  n_9389;
assign n_9391 = ~n_4016 &  n_9390;
assign n_9392 = ~n_4010 &  n_9391;
assign n_9393 = ~n_4004 &  n_9392;
assign n_9394 = ~n_3998 &  n_9393;
assign n_9395 = ~n_3992 &  n_9394;
assign n_9396 = ~n_3986 &  n_9395;
assign n_9397 = ~n_3980 &  n_9396;
assign n_9398 = ~n_3974 &  n_9397;
assign n_9399 = ~n_3968 &  n_9398;
assign n_9400 = ~n_3962 &  n_9399;
assign n_9401 = ~n_3956 &  n_9400;
assign n_9402 = ~n_3950 &  n_9401;
assign n_9403 = ~n_3944 &  n_9402;
assign n_9404 = ~n_3938 &  n_9403;
assign n_9405 = ~n_3930 &  n_9404;
assign n_9406 = ~n_3924 &  n_9405;
assign n_9407 = ~n_3918 &  n_9406;
assign n_9408 = ~n_3912 &  n_9407;
assign n_9409 = ~n_3906 &  n_9408;
assign n_9410 = ~n_3900 &  n_9409;
assign n_9411 = ~n_3894 &  n_9410;
assign n_9412 = ~n_3888 &  n_9411;
assign n_9413 = ~n_3882 &  n_9412;
assign n_9414 = ~n_3876 &  n_9413;
assign n_9415 = ~n_3870 &  n_9414;
assign n_9416 = ~n_3864 &  n_9415;
assign n_9417 = ~n_3858 &  n_9416;
assign n_9418 = ~n_3852 &  n_9417;
assign n_9419 = ~n_3846 &  n_9418;
assign n_9420 = ~n_3840 &  n_9419;
assign n_9421 = ~n_3834 &  n_9420;
assign n_9422 = ~n_3828 &  n_9421;
assign n_9423 = ~n_3822 &  n_9422;
assign n_9424 = ~n_3816 &  n_9423;
assign n_9425 = ~n_3810 &  n_9424;
assign n_9426 = ~n_3804 &  n_9425;
assign n_9427 = ~n_3798 &  n_9426;
assign n_9428 = ~n_3792 &  n_9427;
assign n_9429 = ~n_3786 &  n_9428;
assign n_9430 = ~n_3780 &  n_9429;
assign n_9431 = ~n_3774 &  n_9430;
assign n_9432 = ~n_3768 &  n_9431;
assign n_9433 = ~n_3762 &  n_9432;
assign n_9434 = ~n_3756 &  n_9433;
assign n_9435 = ~n_3750 &  n_9434;
assign n_9436 = ~n_3744 &  n_9435;
assign n_9437 = ~n_3738 &  n_9436;
assign n_9438 = ~n_3732 &  n_9437;
assign n_9439 = ~n_3726 &  n_9438;
assign n_9440 = ~n_3720 &  n_9439;
assign n_9441 = ~n_3714 &  n_9440;
assign n_9442 = ~n_3708 &  n_9441;
assign n_9443 = ~n_3702 &  n_9442;
assign n_9444 = ~n_3696 &  n_9443;
assign n_9445 = ~n_3690 &  n_9444;
assign n_9446 = ~n_3684 &  n_9445;
assign n_9447 = ~n_3678 &  n_9446;
assign n_9448 = ~n_3672 &  n_9447;
assign n_9449 = ~n_3666 &  n_9448;
assign n_9450 = ~n_3660 &  n_9449;
assign n_9451 = ~n_3654 &  n_9450;
assign n_9452 = ~n_3648 &  n_9451;
assign n_9453 = ~n_3642 &  n_9452;
assign n_9454 = ~n_3636 &  n_9453;
assign n_9455 = ~n_3630 &  n_9454;
assign n_9456 = ~n_3624 &  n_9455;
assign n_9457 = ~n_3618 &  n_9456;
assign n_9458 = ~n_3612 &  n_9457;
assign n_9459 = ~n_3606 &  n_9458;
assign n_9460 = ~n_3600 &  n_9459;
assign n_9461 = ~n_3594 &  n_9460;
assign n_9462 = ~n_3588 &  n_9461;
assign n_9463 = ~n_3582 &  n_9462;
assign n_9464 = ~n_3576 &  n_9463;
assign n_9465 = ~n_3570 &  n_9464;
assign n_9466 = ~n_3564 &  n_9465;
assign n_9467 = ~n_3558 &  n_9466;
assign n_9468 = ~n_3552 &  n_9467;
assign n_9469 = ~n_3546 &  n_9468;
assign n_9470 = ~n_3540 &  n_9469;
assign n_9471 = ~n_3534 &  n_9470;
assign n_9472 = ~n_3528 &  n_9471;
assign n_9473 = ~n_3522 &  n_9472;
assign n_9474 = ~n_3517 &  n_9473;
assign n_9475 = ~n_3512 &  n_9474;
assign n_9476 = ~n_3507 &  n_9475;
assign n_9477 = ~n_3502 &  n_9476;
assign n_9478 = ~n_3497 &  n_9477;
assign n_9479 = ~n_3492 &  n_9478;
assign n_9480 = ~n_3487 &  n_9479;
assign n_9481 = ~n_3482 &  n_9480;
assign n_9482 = ~n_3477 &  n_9481;
assign n_9483 = ~n_3472 &  n_9482;
assign n_9484 = ~n_3467 &  n_9483;
assign n_9485 = ~n_3462 &  n_9484;
assign n_9486 = ~n_3457 &  n_9485;
assign n_9487 = ~n_3452 &  n_9486;
assign n_9488 = ~n_3447 &  n_9487;
assign n_9489 = ~n_3442 &  n_9488;
assign n_9490 = ~n_3437 &  n_9489;
assign n_9491 = ~n_3432 &  n_9490;
assign n_9492 = ~n_3427 &  n_9491;
assign n_9493 = ~n_3422 &  n_9492;
assign n_9494 = ~n_3417 &  n_9493;
assign n_9495 = ~n_3412 &  n_9494;
assign n_9496 = ~n_3407 &  n_9495;
assign n_9497 = ~n_3401 &  n_9496;
assign n_9498 = ~n_3395 &  n_9497;
assign n_9499 = ~n_3389 &  n_9498;
assign n_9500 = ~n_3383 &  n_9499;
assign n_9501 = ~n_3377 &  n_9500;
assign n_9502 = ~n_3371 &  n_9501;
assign n_9503 = ~n_3365 &  n_9502;
assign n_9504 = ~n_3359 &  n_9503;
assign n_9505 = ~n_3353 &  n_9504;
assign n_9506 = ~n_3347 &  n_9505;
assign n_9507 = ~n_3341 &  n_9506;
assign n_9508 = ~n_3335 &  n_9507;
assign n_9509 = ~n_3329 &  n_9508;
assign n_9510 = ~n_3323 &  n_9509;
assign n_9511 = ~n_3317 &  n_9510;
assign n_9512 = ~n_3311 &  n_9511;
assign n_9513 = ~n_3305 &  n_9512;
assign n_9514 = ~n_3299 &  n_9513;
assign n_9515 = ~n_3293 &  n_9514;
assign n_9516 = ~n_3287 &  n_9515;
assign n_9517 = ~n_3281 &  n_9516;
assign n_9518 = ~n_3274 &  n_9517;
assign n_9519 = ~n_3268 &  n_9518;
assign n_9520 = ~n_3262 &  n_9519;
assign n_9521 = ~n_3256 &  n_9520;
assign n_9522 = ~n_3250 &  n_9521;
assign n_9523 = ~n_3243 &  n_9522;
assign n_9524 = ~n_3237 &  n_9523;
assign n_9525 = ~n_3231 &  n_9524;
assign n_9526 = ~n_3225 &  n_9525;
assign n_9527 = ~n_3218 &  n_9526;
assign n_9528 = ~n_3211 &  n_9527;
assign n_9529 = ~n_3205 &  n_9528;
assign n_9530 = ~n_3199 &  n_9529;
assign n_9531 = ~n_3193 &  n_9530;
assign n_9532 = ~n_3187 &  n_9531;
assign n_9533 = ~n_3181 &  n_9532;
assign n_9534 = ~n_3175 &  n_9533;
assign n_9535 = ~n_3169 &  n_9534;
assign n_9536 = ~n_3163 &  n_9535;
assign n_9537 = ~n_3157 &  n_9536;
assign n_9538 = ~n_3151 &  n_9537;
assign n_9539 = ~n_3145 &  n_9538;
assign n_9540 = ~n_3139 &  n_9539;
assign n_9541 = ~n_3133 &  n_9540;
assign n_9542 = ~n_3127 &  n_9541;
assign n_9543 = ~n_3121 &  n_9542;
assign n_9544 = ~n_3115 &  n_9543;
assign n_9545 = ~n_3109 &  n_9544;
assign n_9546 = ~n_3103 &  n_9545;
assign n_9547 = ~n_3097 &  n_9546;
assign n_9548 = ~n_3091 &  n_9547;
assign n_9549 = ~n_3085 &  n_9548;
assign n_9550 = ~n_3079 &  n_9549;
assign n_9551 = ~n_3073 &  n_9550;
assign n_9552 = ~n_3067 &  n_9551;
assign n_9553 = ~n_3061 &  n_9552;
assign n_9554 = ~n_3055 &  n_9553;
assign n_9555 = ~n_3049 &  n_9554;
assign n_9556 = ~n_3043 &  n_9555;
assign n_9557 = ~n_3037 &  n_9556;
assign n_9558 = ~n_3031 &  n_9557;
assign n_9559 = ~n_3025 &  n_9558;
assign n_9560 = ~n_3019 &  n_9559;
assign n_9561 = ~n_3013 &  n_9560;
assign n_9562 = ~n_3007 &  n_9561;
assign n_9563 = ~n_3001 &  n_9562;
assign n_9564 = ~n_2995 &  n_9563;
assign n_9565 = ~n_2989 &  n_9564;
assign n_9566 = ~n_2983 &  n_9565;
assign n_9567 = ~n_2977 &  n_9566;
assign n_9568 = ~n_2971 &  n_9567;
assign n_9569 = ~n_2965 &  n_9568;
assign n_9570 = ~n_2959 &  n_9569;
assign n_9571 = ~n_2953 &  n_9570;
assign n_9572 = ~n_2947 &  n_9571;
assign n_9573 = ~n_2941 &  n_9572;
assign n_9574 = ~n_2935 &  n_9573;
assign n_9575 = ~n_2929 &  n_9574;
assign n_9576 = ~n_2923 &  n_9575;
assign n_9577 = ~n_2917 &  n_9576;
assign n_9578 = ~n_2911 &  n_9577;
assign n_9579 = ~n_2905 &  n_9578;
assign n_9580 = ~n_2899 &  n_9579;
assign n_9581 = ~n_2893 &  n_9580;
assign n_9582 = ~n_2887 &  n_9581;
assign n_9583 = ~n_2881 &  n_9582;
assign n_9584 = ~n_2875 &  n_9583;
assign n_9585 = ~n_2869 &  n_9584;
assign n_9586 = ~n_2863 &  n_9585;
assign n_9587 = ~n_2857 &  n_9586;
assign n_9588 = ~n_2851 &  n_9587;
assign n_9589 = ~n_2845 &  n_9588;
assign n_9590 = ~n_2839 &  n_9589;
assign n_9591 = ~n_2833 &  n_9590;
assign n_9592 = ~n_2827 &  n_9591;
assign n_9593 = ~n_2823 &  n_9592;
assign n_9594 = ~n_2817 &  n_9593;
assign n_9595 = ~n_2811 &  n_9594;
assign n_9596 = ~n_2805 &  n_9595;
assign n_9597 = ~n_2799 &  n_9596;
assign n_9598 = ~n_2793 &  n_9597;
assign n_9599 = ~n_2787 &  n_9598;
assign n_9600 = ~n_2781 &  n_9599;
assign n_9601 = ~n_2775 &  n_9600;
assign n_9602 = ~n_2769 &  n_9601;
assign n_9603 = ~n_2763 &  n_9602;
assign n_9604 = ~n_2757 &  n_9603;
assign n_9605 = ~n_2751 &  n_9604;
assign n_9606 = ~n_2745 &  n_9605;
assign n_9607 = ~n_2739 &  n_9606;
assign n_9608 = ~n_2733 &  n_9607;
assign n_9609 = ~n_2727 &  n_9608;
assign n_9610 = ~n_2721 &  n_9609;
assign n_9611 = ~n_2715 &  n_9610;
assign n_9612 = ~n_2709 &  n_9611;
assign n_9613 = ~n_2703 &  n_9612;
assign n_9614 = ~n_2697 &  n_9613;
assign n_9615 = ~n_2691 &  n_9614;
assign n_9616 = ~n_2685 &  n_9615;
assign n_9617 = ~n_2679 &  n_9616;
assign n_9618 = ~n_2673 &  n_9617;
assign n_9619 = ~n_2667 &  n_9618;
assign n_9620 = ~n_2661 &  n_9619;
assign n_9621 = ~n_2655 &  n_9620;
assign n_9622 = ~n_2649 &  n_9621;
assign n_9623 = ~n_2643 &  n_9622;
assign n_9624 = ~n_2637 &  n_9623;
assign n_9625 = ~n_2580 &  n_9624;
assign n_9626 = ~n_2508 &  n_9625;
assign n_9627 = ~n_2443 &  n_9626;
assign n_9628 = ~n_2358 &  n_9627;
assign n_9629 = ~n_2267 &  n_9628;
assign n_9630 = ~n_2148 &  n_9629;
assign n_9631 = ~n_2021 &  n_9630;
assign n_9632 = ~n_1773 &  n_9631;
assign n_9633 = ~n_1456 &  n_9632;
assign n_9634 = ~n_153 &  n_9633;
assign n_9635 = ~n_147 &  n_9634;
assign n_9636 = ~n_141 &  n_9635;
assign n_9637 = ~n_135 &  n_9636;
assign n_9638 = ~n_129 &  n_9637;
assign n_9639 = ~n_123 &  n_9638;
assign n_9640 = ~n_117 &  n_9639;
assign n_9641 = ~n_111 &  n_9640;
assign n_9642 = ~n_105 &  n_9641;
assign n_9643 = ~n_99 &  n_9642;
assign n_9644 = ~n_93 &  n_9643;
assign n_9645 = ~n_87 &  n_9644;
assign n_9646 = ~n_81 &  n_9645;
assign n_9647 = ~n_75 &  n_9646;
assign n_9648 = ~n_69 &  n_9647;
assign n_9649 = ~n_63 &  n_9648;
assign n_9650 = ~n_57 &  n_9649;
assign n_9651 = ~n_51 &  n_9650;
assign n_9652 = ~n_45 &  n_9651;
assign n_9653 = ~n_39 &  n_9652;
assign n_9654 = ~n_33 &  n_9653;
assign n_9655 = ~n_27 &  n_9654;
assign n_9656 = ~n_21 &  n_9655;
assign n_9657 = ~n_15 &  n_9656;
assign o_1 = ~n_9657;
endmodule

