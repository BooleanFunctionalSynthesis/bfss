// Generated using findDep.cpp 
module query06_query42_1344n (v_1, v_2, v_3, v_4, v_5, v_6, v_7, v_8, v_9, v_10, v_11, v_12, v_13, v_14, v_15, v_16, v_17, v_18, v_19, v_20, v_21, v_22, v_23, v_24, v_25, v_27, v_28, v_29, v_30, v_31, v_32, v_33, v_34, v_35, v_36, v_37, v_38, v_39, v_40, v_41, v_42, v_43, v_44, v_45, v_46, v_47, v_48, v_49, v_50, v_51, v_52, v_53, v_54, v_55, v_56, v_57, v_58, v_59, v_60, v_61, v_62, v_63, v_64, v_65, v_66, v_67, v_68, v_69, v_70, v_71, v_72, v_73, v_74, v_75, v_76, v_77, v_78, v_79, v_80, v_81, v_82, v_83, v_84, v_85, v_86, v_87, v_88, v_89, v_90, v_91, v_92, v_93, v_94, v_95, v_96, v_100, v_101, v_102, v_103, v_104, v_105, v_106, v_107, v_108, v_109, v_110, v_111, v_112, v_113, v_117, v_120, v_121, v_122, v_126, v_127, v_128, v_131, v_132, v_26, v_97, v_98, v_99, v_114, v_115, v_116, v_118, v_119, v_123, v_124, v_125, v_129, v_130, v_133, v_134, v_135, v_136, v_137, v_138, v_139, v_140, v_141, v_142, v_143, v_144, v_145, v_146, v_147, v_148, v_149, v_150, v_151, v_152, v_153, v_154, v_155, v_156, v_157, v_158, v_159, v_160, v_161, v_162, v_163, v_164, v_165, v_166, v_167, v_168, v_169, v_170, v_171, v_172, v_173, v_174, v_175, v_176, v_177, v_178, v_179, v_180, v_181, v_182, v_183, v_184, v_185, v_186, v_187, v_188, v_189, v_190, v_191, v_192, v_193, v_194, v_195, v_196, v_197, v_198, v_199, v_200, v_201, v_202, v_203, v_204, v_205, v_206, v_207, v_208, v_209, v_210, v_211, v_212, v_213, v_214, v_215, v_216, v_217, v_218, v_219, v_220, v_221, v_222, v_223, v_224, v_225, v_226, v_227, v_228, v_229, v_230, v_231, v_232, v_233, v_234, v_235, v_236, v_237, v_238, v_239, v_240, v_241, v_242, v_243, v_244, v_245, v_246, v_247, v_248, v_249, v_250, v_251, v_252, v_253, v_254, v_255, v_256, v_257, v_258, v_259, v_260, v_261, v_262, v_263, v_264, v_265, v_266, v_267, v_268, v_269, v_270, v_271, v_272, v_273, v_274, v_275, v_276, v_277, v_278, v_279, v_280, v_281, v_282, v_283, v_284, v_285, v_286, v_287, v_288, v_289, v_290, v_291, v_292, v_293, v_294, v_295, v_296, v_297, v_298, v_299, v_300, v_301, v_302, v_303, v_304, v_305, v_306, v_307, v_308, v_309, v_310, v_311, v_312, v_313, v_314, v_315, v_316, v_317, v_318, v_319, v_320, v_321, v_322, v_323, v_324, v_325, v_326, v_327, v_328, v_329, v_330, v_331, v_332, v_333, v_334, v_335, v_336, v_337, v_338, v_339, v_340, v_341, v_342, v_343, v_344, v_345, v_346, v_347, v_348, v_349, v_350, v_351, v_352, v_353, v_354, v_355, v_356, v_357, v_358, v_359, v_360, v_361, v_362, v_363, v_364, v_365, v_366, v_367, v_368, v_369, v_370, v_371, v_372, v_373, v_374, v_375, v_376, v_377, v_378, v_379, v_380, v_381, v_382, v_383, v_384, v_385, v_386, v_387, v_388, v_389, v_390, v_391, v_392, v_393, v_394, v_395, v_396, v_397, v_398, v_399, v_400, v_401, v_402, v_403, v_404, v_405, v_406, v_407, v_408, v_409, v_410, v_411, v_412, v_413, v_414, v_415, v_416, v_417, v_418, v_419, v_420, v_421, v_422, v_423, v_424, v_425, v_426, v_427, v_428, v_429, v_430, v_431, v_432, v_433, v_434, v_435, v_436, v_437, v_438, v_439, v_440, v_441, v_442, v_443, v_444, v_445, v_446, v_447, v_448, v_449, v_450, v_451, v_452, v_453, v_454, v_455, v_456, v_457, v_458, v_459, v_460, v_461, v_462, v_463, v_464, v_465, v_466, v_467, v_468, v_469, v_470, v_471, v_472, v_473, v_474, v_475, v_476, v_477, v_478, v_479, v_480, v_481, v_482, v_483, v_484, v_485, v_486, v_487, v_488, v_489, v_490, v_491, v_492, v_493, v_494, v_495, v_496, v_497, v_498, v_499, v_500, v_501, v_502, v_503, v_504, v_505, v_506, v_507, v_508, v_509, v_510, v_511, v_512, v_513, v_514, v_515, v_516, v_517, v_518, v_519, v_520, v_521, v_522, v_523, v_524, v_525, v_526, v_527, v_528, v_529, v_530, v_531, v_532, v_533, v_534, v_535, v_536, v_537, v_538, v_539, v_540, v_541, v_542, v_543, v_544, v_545, v_546, v_547, v_548, v_549, v_550, v_551, v_552, v_553, v_554, v_555, v_556, v_557, v_558, v_559, v_560, v_561, v_562, v_563, v_564, v_565, v_566, v_567, v_568, v_569, v_570, v_571, v_572, v_573, v_574, v_575, v_576, v_577, v_578, v_579, v_580, v_581, v_582, v_583, v_584, v_585, v_586, v_587, v_588, v_589, v_590, v_591, v_592, v_593, v_594, v_595, v_596, v_597, v_598, v_599, v_600, v_601, v_602, v_603, v_604, v_605, v_606, v_607, v_608, v_609, v_610, v_611, v_612, v_613, v_614, v_615, v_616, v_617, v_618, v_619, v_620, v_621, v_622, v_623, v_624, v_625, v_626, v_627, v_628, v_629, v_630, v_631, v_632, v_633, v_634, v_635, v_636, v_637, v_638, v_639, v_640, v_641, v_642, v_643, v_644, v_645, v_646, v_647, v_648, v_649, v_650, v_651, v_652, v_653, v_654, v_655, v_656, v_657, v_658, v_659, v_660, v_661, v_662, v_663, v_664, v_665, v_666, v_667, v_668, v_669, v_670, v_671, v_672, v_673, v_674, v_675, v_676, v_677, v_678, v_679, v_680, v_681, v_682, v_683, v_684, v_685, v_686, v_687, v_688, v_689, v_690, v_691, v_692, v_693, v_694, v_695, v_696, v_697, v_698, v_699, v_700, v_701, v_702, v_703, v_704, v_705, v_706, v_707, v_708, v_709, v_710, v_711, v_712, v_713, v_714, v_715, v_716, v_717, v_718, v_719, v_720, v_721, v_722, v_723, v_724, v_725, v_726, v_727, v_728, v_729, v_730, v_731, v_732, v_733, v_734, v_735, v_736, v_737, v_738, v_739, v_740, v_741, v_742, v_743, v_744, v_745, v_746, v_747, v_748, v_749, v_750, v_751, v_752, v_753, v_754, v_755, v_756, v_757, v_758, v_759, v_760, v_761, v_762, v_763, v_764, v_765, v_766, v_767, v_768, v_769, v_770, v_771, v_772, v_773, v_774, v_775, v_776, v_777, v_778, v_779, v_780, v_781, v_782, v_783, v_784, v_785, v_786, v_787, v_788, v_789, v_790, v_791, v_792, v_793, v_794, v_795, v_796, v_797, v_798, v_799, v_800, v_801, v_802, v_803, v_804, v_805, v_806, v_807, v_808, v_809, v_810, v_811, v_812, v_813, v_814, v_815, v_816, v_817, v_818, v_819, v_820, v_821, v_822, v_823, v_824, v_825, v_826, v_827, v_828, v_829, v_830, v_831, v_832, v_833, v_834, v_835, v_836, v_837, v_838, v_839, v_840, v_841, v_842, v_843, v_844, v_845, v_846, v_847, v_848, v_849, v_850, v_851, v_852, v_853, v_854, v_855, v_856, v_857, v_858, v_859, v_860, v_861, v_862, v_863, v_864, v_865, v_866, v_867, v_868, v_869, v_870, v_871, v_872, v_873, v_874, v_875, v_876, v_877, v_878, v_879, v_880, v_881, v_882, v_883, v_884, v_885, v_886, v_887, v_888, v_889, v_890, v_891, v_892, v_893, v_894, v_895, v_896, v_897, v_898, v_899, v_900, v_901, v_902, v_903, v_904, v_905, v_906, v_907, v_908, v_909, v_910, v_911, v_912, v_913, v_914, v_915, v_916, v_917, v_918, v_919, v_920, v_921, v_922, v_923, v_924, v_925, v_926, v_927, v_928, v_929, v_930, v_931, v_932, v_933, v_934, v_935, v_936, v_937, v_938, v_939, v_940, v_941, v_942, v_943, v_944, v_945, v_946, v_947, v_948, v_949, v_950, v_951, v_952, v_953, v_954, v_955, v_956, v_957, v_958, v_959, v_960, v_961, v_962, v_963, v_964, v_965, v_966, v_967, v_968, v_969, v_970, v_971, v_972, v_973, v_974, v_975, v_976, v_977, v_978, v_979, v_980, v_981, v_982, v_983, v_984, v_985, v_986, v_987, v_988, v_989, v_990, v_991, v_992, v_993, v_994, v_995, v_996, v_997, v_998, v_999, v_1000, v_1001, v_1002, v_1003, v_1004, v_1005, v_1006, v_1007, v_1008, v_1009, v_1010, v_1011, v_1012, v_1013, v_1014, v_1015, v_1016, v_1017, v_1018, v_1019, v_1020, v_1021, v_1022, v_1023, v_1024, v_1025, v_1026, v_1027, v_1028, v_1029, v_1030, v_1031, v_1032, v_1033, v_1034, v_1035, v_1036, v_1037, v_1038, v_1039, v_1040, v_1041, v_1042, v_1043, v_1044, v_1045, v_1046, v_1047, v_1048, v_1049, v_1050, v_1051, v_1052, v_1053, v_1054, v_1055, v_1056, v_1057, v_1058, v_1059, v_1060, v_1061, v_1062, v_1063, v_1064, v_1065, v_1066, v_1067, v_1068, v_1069, v_1070, v_1071, v_1072, v_1073, v_1074, v_1075, v_1076, v_1077, v_1078, v_1079, v_1080, v_1081, v_1082, v_1083, v_1084, v_1085, v_1086, v_1087, v_1088, v_1089, v_1090, v_1091, v_1092, v_1093, v_1094, v_1095, v_1096, v_1097, v_1098, v_1099, v_1100, v_1101, v_1102, v_1103, v_1104, v_1105, v_1106, v_1107, v_1108, v_1109, v_1110, v_1111, v_1112, v_1113, v_1114, v_1115, v_1116, v_1117, v_1118, v_1119, v_1120, v_1121, v_1122, v_1123, v_1124, v_1125, v_1126, v_1127, v_1128, v_1129, v_1130, v_1131, v_1132, v_1133, v_1134, v_1135, v_1136, v_1137, v_1138, v_1139, v_1140, v_1141, v_1142, v_1143, v_1144, v_1145, v_1146, v_1147, v_1148, v_1149, v_1150, v_1151, v_1152, v_1153, v_1154, v_1155, v_1156, v_1157, v_1158, v_1159, v_1160, v_1161, v_1162, v_1163, v_1164, v_1165, v_1166, v_1167, v_1168, v_1169, v_1170, v_1171, v_1172, v_1173, v_1174, v_1175, v_1176, v_1177, v_1178, v_1179, v_1180, v_1181, v_1182, v_1183, v_1184, v_1185, v_1186, v_1187, v_1188, v_1189, v_1190, v_1191, v_1192, v_1193, v_1194, v_1195, v_1196, v_1197, v_1198, v_1199, v_1200, v_1201, v_1202, v_1203, v_1204, v_1205, v_1206, v_1207, v_1208, v_1209, v_1210, v_1211, v_1212, v_1213, v_1214, v_1215, v_1216, v_1217, v_1218, v_1219, v_1220, v_1221, v_1222, v_1223, v_1224, v_1225, v_1226, v_1227, v_1228, v_1229, v_1230, v_1231, v_1232, v_1233, v_1234, v_1235, v_1236, v_1237, v_1238, v_1239, v_1240, v_1241, v_1242, v_1243, v_1244, v_1245, v_1246, v_1247, v_1248, v_1249, v_1250, v_1251, v_1252, v_1253, v_1254, v_1255, v_1256, v_1257, v_1258, v_1259, v_1260, v_1261, v_1262, v_1263, v_1264, v_1265, v_1266, v_1267, v_1268, v_1269, v_1270, v_1271, v_1272, v_1273, v_1274, v_1275, v_1276, v_1277, v_1278, v_1279, v_1280, v_1281, v_1282, v_1283, v_1284, v_1285, v_1286, v_1287, v_1288, v_1289, v_1290, v_1291, v_1292, v_1293, v_1294, v_1295, v_1296, v_1297, v_1298, v_1299, v_1300, v_1301, v_1302, v_1303, v_1304, v_1305, v_1306, v_1307, v_1308, v_1309, v_1310, v_1311, v_1312, v_1313, v_1314, v_1315, v_1316, v_1317, v_1318, v_1319, v_1320, v_1321, v_1322, v_1323, v_1324, v_1325, v_1326, v_1327, v_1328, v_1329, v_1330, v_1331, v_1332, v_1333, v_1334, v_1335, v_1336, v_1337, v_1338, v_1339, v_1340, v_1341, v_1342, v_1343, v_1344, v_1345, v_1346, v_1347, v_1348, v_1349, v_1350, v_1351, v_1352, v_1353, v_1354, v_1355, v_1356, v_1357, v_1358, v_1359, v_1360, v_1361, v_1362, v_1363, v_1364, v_1365, v_1366, v_1367, v_1368, v_1369, v_1370, v_1371, v_1372, v_1373, v_1374, v_1375, v_1376, v_1377, v_1378, v_1379, v_1380, v_1381, v_1382, v_1383, v_1384, v_1385, v_1386, v_1387, v_1388, v_1389, v_1390, v_1391, v_1392, v_1393, v_1394, v_1395, v_1396, v_1397, v_1398, v_1399, v_1400, v_1401, v_1402, v_1403, v_1404, v_1405, v_1406, v_1407, v_1408, v_1409, v_1410, v_1411, v_1412, v_1413, v_1414, v_1415, v_1416, v_1417, v_1418, v_1419, v_1420, v_1421, v_1422, v_1423, v_1424, v_1425, v_1426, v_1427, v_1428, v_1429, v_1430, v_1431, v_1432, v_1433, v_1434, v_1435, v_1436, v_1437, v_1438, v_1439, v_1440, v_1441, v_1442, v_1443, v_1444, v_1445, v_1446, v_1447, v_1448, v_1449, v_1450, v_1451, v_1452, v_1453, v_1454, v_1455, v_1456, v_1457, v_1458, v_1459, v_1460, v_1461, v_1462, v_1463, v_1464, v_1465, v_1466, v_1467, v_1468, v_1469, v_1470, v_1471, v_1472, v_1473, v_1474, v_1475, v_1476, v_1477, v_1478, v_1479, v_1480, v_1481, v_1482, v_1483, v_1484, v_1485, v_1486, v_1487, v_1488, v_1489, v_1490, v_1491, v_1492, v_1493, v_1494, v_1495, v_1496, v_1497, v_1498, v_1499, v_1500, v_1501, v_1502, v_1503, v_1504, v_1505, v_1506, v_1507, v_1508, v_1509, v_1510, v_1511, v_1512, v_1513, v_1514, v_1515, v_1516, v_1517, v_1518, v_1519, v_1520, v_1521, v_1522, v_1523, v_1524, v_1525, v_1526, v_1527, v_1528, v_1529, v_1530, v_1531, v_1532, v_1533, v_1534, v_1535, v_1536, v_1537, v_1538, v_1539, v_1540, v_1541, v_1542, v_1543, v_1544, v_1545, v_1546, v_1547, v_1548, v_1549, v_1550, v_1551, v_1552, v_1553, v_1554, v_1555, v_1556, v_1557, v_1558, v_1559, v_1560, v_1561, v_1562, v_1563, v_1564, v_1565, v_1566, v_1567, v_1568, v_1569, v_1570, v_1571, v_1572, v_1573, v_1574, v_1575, v_1576, v_1577, v_1578, v_1579, v_1580, v_1581, v_1582, v_1583, v_1584, v_1585, v_1586, v_1587, v_1588, v_1589, v_1590, v_1591, v_1592, v_1593, v_1594, v_1595, v_1596, v_1597, v_1598, v_1599, v_1600, v_1601, v_1602, v_1603, v_1604, v_1605, v_1606, v_1607, v_1608, v_1609, v_1610, v_1611, v_1612, v_1613, v_1614, v_1615, v_1616, v_1617, v_1618, v_1619, v_1620, v_1621, v_1622, v_1623, v_1624, v_1625, v_1626, v_1627, v_1628, v_1629, v_1630, v_1631, v_1632, v_1633, v_1634, v_1635, v_1636, v_1637, v_1638, v_1639, v_1640, v_1641, v_1642, v_1643, v_1644, v_1645, v_1646, v_1647, v_1648, v_1649, v_1650, v_1651, v_1652, v_1653, v_1654, v_1655, v_1656, v_1657, v_1658, v_1659, v_1660, v_1661, v_1662, v_1663, v_1664, v_1665, v_1666, v_1667, v_1668, v_1669, v_1670, v_1671, v_1672, v_1673, v_1674, v_1675, v_1676, v_1677, v_1678, v_1679, v_1680, v_1681, v_1682, v_1683, v_1684, v_1685, v_1686, v_1687, v_1688, v_1689, v_1690, v_1691, v_1692, v_1693, v_1694, v_1695, v_1696, v_1697, v_1698, v_1699, v_1700, v_1701, v_1702, v_1703, v_1704, v_1705, v_1706, v_1707, v_1708, v_1709, v_1710, v_1711, v_1712, v_1713, v_1714, v_1715, v_1716, v_1717, v_1718, v_1719, v_1720, v_1721, v_1722, v_1723, v_1724, v_1725, v_1726, v_1727, v_1728, v_1729, v_1730, v_1731, v_1732, v_1733, v_1734, v_1735, v_1736, v_1737, v_1738, v_1739, v_1740, v_1741, v_1742, v_1743, v_1744, v_1745, v_1746, v_1747, v_1748, v_1749, v_1750, v_1751, v_1752, v_1753, v_1754, v_1755, v_1756, v_1757, v_1758, v_1759, v_1760, v_1761, v_1762, v_1763, v_1764, v_1765, v_1766, v_1767, v_1768, v_1769, v_1770, v_1771, v_1772, v_1773, v_1774, v_1775, v_1776, v_1777, v_1778, v_1779, v_1780, v_1781, v_1782, v_1783, v_1784, v_1785, v_1786, v_1787, v_1788, v_1789, v_1790, v_1791, v_1792, v_1793, v_1794, v_1795, v_1796, v_1797, v_1798, v_1799, v_1800, v_1801, v_1802, v_1803, v_1804, v_1805, v_1806, v_1807, v_1808, v_1809, v_1810, v_1811, v_1812, v_1813, v_1814, v_1815, v_1816, v_1817, v_1818, v_1819, v_1820, v_1821, v_1822, v_1823, v_1824, v_1825, v_1826, v_1827, v_1828, v_1829, v_1830, v_1831, v_1832, v_1833, v_1834, v_1835, v_1836, v_1837, v_1838, v_1839, v_1840, v_1841, v_1842, v_1843, v_1844, v_1845, v_1846, v_1847, v_1848, v_1849, v_1850, v_1851, v_1852, v_1853, v_1854, v_1855, v_1856, v_1857, v_1858, v_1859, v_1860, v_1861, v_1862, v_1863, v_1864, v_1865, v_1866, v_1867, v_1868, v_1869, v_1870, v_1871, v_1872, v_1873, v_1874, v_1875, v_1876, v_1877, v_1878, v_1879, v_1880, v_1881, v_1882, v_1883, v_1884, v_1885, v_1886, v_1887, v_1888, v_1889, v_1890, v_1891, v_1892, v_1893, v_1894, v_1895, v_1896, v_1897, v_1898, v_1899, v_1900, v_1901, v_1902, v_1903, v_1904, v_1905, v_1906, v_1907, v_1908, v_1909, v_1910, v_1911, v_1912, v_1913, v_1914, v_1915, v_1916, v_1917, v_1918, v_1919, v_1920, v_1921, v_1922, v_1923, v_1924, v_1925, v_1926, v_1927, v_1928, v_1929, v_1930, v_1931, v_1932, v_1933, v_1934, v_1935, v_1936, v_1937, v_1938, v_1939, v_1940, v_1941, v_1942, v_1943, v_1944, v_1945, v_1946, v_1947, v_1948, v_1949, v_1950, v_1951, v_1952, v_1953, v_1954, v_1955, v_1956, v_1957, v_1958, v_1959, v_1960, v_1961, v_1962, v_1963, v_1964, v_1965, v_1966, v_1967, v_1968, v_1969, v_1970, v_1971, v_1972, v_1973, v_1974, v_1975, v_1976, v_1977, v_1978, v_1979, v_1980, v_1981, v_1982, v_1983, v_1984, v_1985, v_1986, v_1987, v_1988, v_1989, v_1990, v_1991, v_1992, v_1993, v_1994, v_1995, v_1996, v_1997, v_1998, v_1999, v_2000, v_2001, v_2002, v_2003, v_2004, v_2005, v_2006, v_2007, v_2008, v_2009, v_2010, v_2011, v_2012, v_2013, v_2014, v_2015, v_2016, v_2017, v_2018, v_2019, v_2020, v_2021, v_2022, v_2023, v_2024, v_2025, v_2026, v_2027, v_2028, v_2029, v_2030, v_2031, v_2032, v_2033, v_2034, v_2035, v_2036, v_2037, v_2038, v_2039, v_2040, v_2041, v_2042, v_2043, v_2044, v_2045, v_2046, v_2047, v_2048, v_2049, v_2050, v_2051, v_2052, v_2053, v_2054, v_2055, v_2056, v_2057, v_2058, v_2059, v_2060, v_2061, v_2062, v_2063, v_2064, v_2065, v_2066, v_2067, v_2068, v_2069, v_2070, v_2071, v_2072, v_2073, v_2074, v_2075, v_2076, v_2077, v_2078, v_2079, v_2080, v_2081, v_2082, v_2083, v_2084, v_2085, v_2086, v_2087, v_2088, v_2089, v_2090, v_2091, v_2092, v_2093, v_2094, v_2095, v_2096, v_2097, v_2098, v_2099, v_2100, v_2101, v_2102, v_2103, v_2104, v_2105, v_2106, v_2107, v_2108, v_2109, v_2110, v_2111, v_2112, v_2113, v_2114, v_2115, v_2116, v_2117, v_2118, v_2119, v_2120, v_2121, v_2122, v_2123, v_2124, v_2125, v_2126, v_2127, v_2128, v_2129, v_2130, v_2131, v_2132, v_2133, v_2134, v_2135, v_2136, v_2137, v_2138, v_2139, v_2140, v_2141, v_2142, v_2143, v_2144, v_2145, v_2146, v_2147, v_2148, v_2149, v_2150, v_2151, v_2152, v_2153, v_2154, v_2155, v_2156, v_2157, v_2158, v_2159, v_2160, v_2161, v_2162, v_2163, v_2164, v_2165, v_2166, v_2167, v_2168, v_2169, v_2170, v_2171, v_2172, v_2173, v_2174, v_2175, v_2176, v_2177, v_2178, v_2179, v_2180, v_2181, v_2182, v_2183, v_2184, v_2185, v_2186, v_2187, v_2188, v_2189, v_2190, v_2191, v_2192, v_2193, v_2194, v_2195, v_2196, v_2197, v_2198, v_2199, v_2200, v_2201, v_2202, v_2203, v_2204, v_2205, v_2206, v_2207, v_2208, v_2209, v_2210, v_2211, v_2212, v_2213, v_2214, v_2215, v_2216, v_2217, v_2218, v_2219, v_2220, v_2221, v_2222, v_2223, v_2224, v_2225, v_2226, v_2227, v_2228, v_2229, v_2230, v_2231, v_2232, v_2233, v_2234, v_2235, v_2236, v_2237, v_2238, v_2239, v_2240, v_2241, v_2242, v_2243, v_2244, v_2245, v_2246, v_2247, v_2248, v_2249, v_2250, v_2251, v_2252, v_2253, v_2254, v_2255, v_2256, v_2257, v_2258, v_2259, v_2260, v_2261, v_2262, v_2263, v_2264, v_2265, v_2266, v_2267, v_2268, v_2269, v_2270, v_2271, v_2272, v_2273, v_2274, v_2275, v_2276, v_2277, v_2278, v_2279, v_2280, v_2281, v_2282, v_2283, v_2284, v_2285, v_2286, v_2287, v_2288, v_2289, v_2290, v_2291, v_2292, v_2293, v_2294, v_2295, v_2296, v_2297, v_2298, v_2299, v_2300, v_2301, v_2302, v_2303, v_2304, v_2305, v_2306, v_2307, v_2308, v_2309, v_2310, v_2311, v_2312, v_2313, v_2314, v_2315, v_2316, v_2317, v_2318, v_2319, v_2320, v_2321, v_2322, v_2323, v_2324, v_2325, v_2326, v_2327, v_2328, v_2329, v_2330, v_2331, v_2332, v_2333, v_2334, v_2335, v_2336, v_2337, v_2338, v_2339, v_2340, v_2341, v_2342, v_2343, v_2344, v_2345, v_2346, v_2347, v_2348, v_2349, v_2350, v_2351, v_2352, v_2353, v_2354, v_2355, v_2356, v_2357, v_2358, v_2359, v_2360, v_2361, v_2362, v_2363, v_2364, v_2365, v_2366, v_2367, v_2368, v_2369, v_2370, v_2371, v_2372, v_2373, v_2374, v_2375, v_2376, v_2377, v_2378, v_2379, v_2380, v_2381, v_2382, v_2383, v_2384, v_2385, v_2386, v_2387, v_2388, v_2389, v_2390, v_2391, v_2392, v_2393, v_2394, v_2395, v_2396, v_2397, v_2398, v_2399, v_2400, v_2401, v_2402, v_2403, v_2404, v_2405, v_2406, v_2407, v_2408, v_2409, v_2410, v_2411, v_2412, v_2413, v_2414, v_2415, v_2416, v_2417, v_2418, v_2419, v_2420, v_2421, v_2422, v_2423, v_2424, v_2425, v_2426, v_2427, v_2428, v_2429, v_2430, v_2431, v_2432, v_2433, v_2434, v_2435, v_2436, v_2437, v_2438, v_2439, v_2440, v_2441, v_2442, v_2443, v_2444, v_2445, v_2446, v_2447, v_2448, v_2449, v_2450, v_2451, v_2452, v_2453, v_2454, v_2455, v_2456, v_2457, v_2458, v_2459, v_2460, v_2461, v_2462, v_2463, v_2464, v_2465, v_2466, v_2467, v_2468, v_2469, v_2470, v_2471, v_2472, v_2473, v_2474, v_2475, v_2476, v_2477, v_2478, v_2479, v_2480, v_2481, v_2482, v_2483, v_2484, v_2485, v_2486, v_2487, v_2488, v_2489, v_2490, v_2491, v_2492, v_2493, v_2494, v_2495, v_2496, v_2497, v_2498, v_2499, v_2500, v_2501, v_2502, v_2503, v_2504, v_2505, v_2506, v_2507, v_2508, v_2509, v_2510, v_2511, v_2512, v_2513, v_2514, v_2515, v_2516, v_2517, v_2518, v_2519, v_2520, v_2521, v_2522, v_2523, v_2524, v_2525, v_2526, v_2527, v_2528, v_2529, v_2530, v_2531, v_2532, v_2533, v_2534, v_2535, v_2536, v_2537, v_2538, v_2539, v_2540, v_2541, v_2542, v_2543, v_2544, v_2545, v_2546, v_2547, v_2548, v_2549, v_2550, v_2551, v_2552, v_2553, v_2554, v_2555, v_2556, v_2557, v_2558, v_2559, v_2560, v_2561, v_2562, v_2563, v_2564, v_2565, v_2566, v_2567, v_2568, v_2569, v_2570, v_2571, v_2572, v_2573, v_2574, v_2575, v_2576, v_2577, v_2578, v_2579, v_2580, v_2581, v_2582, v_2583, v_2584, v_2585, v_2586, v_2587, v_2588, v_2589, v_2590, v_2591, v_2592, v_2593, v_2594, v_2595, v_2596, v_2597, v_2598, v_2599, v_2600, v_2601, v_2602, v_2603, v_2604, v_2605, v_2606, v_2607, v_2608, v_2609, v_2610, v_2611, v_2612, v_2613, v_2614, v_2615, v_2616, v_2617, v_2618, v_2619, v_2620, v_2621, v_2622, v_2623, v_2624, v_2625, v_2626, v_2627, v_2628, v_2629, v_2630, v_2631, v_2632, v_2633, v_2634, v_2635, v_2636, v_2637, v_2638, v_2639, v_2640, v_2641, v_2642, v_2643, v_2644, v_2645, v_2646, v_2647, v_2648, v_2649, v_2650, v_2651, v_2652, v_2653, v_2654, v_2655, v_2656, v_2657, v_2658, v_2659, v_2660, v_2661, v_2662, v_2663, v_2664, v_2665, v_2666, v_2667, v_2668, v_2669, v_2670, v_2671, v_2672, v_2673, v_2674, v_2675, v_2676, v_2677, v_2678, v_2679, v_2680, v_2681, v_2682, v_2683, v_2684, v_2685, v_2686, v_2687, v_2688, v_2689, v_2690, v_2691, v_2692, v_2693, v_2694, v_2695, v_2696, v_2697, v_2698, v_2699, v_2700, v_2701, v_2702, v_2703, v_2704, v_2705, v_2706, v_2707, v_2708, v_2709, v_2710, v_2711, v_2712, v_2713, v_2714, v_2715, v_2716, v_2717, v_2718, v_2719, v_2720, v_2721, v_2722, v_2723, v_2724, v_2725, v_2726, v_2727, v_2728, v_2729, v_2730, v_2731, v_2732, v_2733, v_2734, v_2735, v_2736, v_2737, v_2738, v_2739, v_2740, v_2741, v_2742, v_2743, v_2744, v_2745, v_2746, v_2747, v_2748, v_2749, v_2750, v_2751, v_2752, v_2753, v_2754, v_2755, v_2756, v_2757, v_2758, v_2759, v_2760, v_2761, v_2762, v_2763, v_2764, v_2765, v_2766, v_2767, v_2768, v_2769, v_2770, v_2771, v_2772, v_2773, v_2774, v_2775, v_2776, v_2777, v_2778, v_2779, v_2780, v_2781, v_2782, v_2783, v_2784, v_2785, v_2786, v_2787, v_2788, v_2789, v_2790, v_2791, v_2792, v_2793, v_2794, v_2795, v_2796, v_2797, v_2798, v_2799, v_2800, v_2801, v_2802, v_2803, v_2804, v_2805, v_2806, v_2807, v_2808, v_2809, v_2810, v_2811, v_2812, v_2813, v_2814, v_2815, v_2816, v_2817, v_2818, v_2819, v_2820, v_2821, v_2822, v_2823, v_2824, v_2825, v_2826, v_2827, v_2828, v_2829, v_2830, v_2831, v_2832, v_2833, v_2834, v_2835, v_2836, v_2837, v_2838, v_2839, v_2840, v_2841, v_2842, v_2843, v_2844, v_2845, v_2846, v_2847, v_2848, v_2849, v_2850, v_2851, v_2852, v_2853, v_2854, v_2855, v_2856, v_2857, v_2858, v_2859, v_2860, v_2861, v_2862, v_2863, v_2864, v_2865, v_2866, v_2867, v_2868, v_2869, v_2870, v_2871, v_2872, v_2873, v_2874, v_2875, v_2876, v_2877, v_2878, v_2879, v_2880, v_2881, v_2882, v_2883, v_2884, v_2885, v_2886, v_2887, v_2888, v_2889, v_2890, v_2891, v_2892, v_2893, v_2894, v_2895, v_2896, v_2897, v_2898, v_2899, v_2900, v_2901, v_2902, v_2903, v_2904, v_2905, v_2906, v_2907, v_2908, v_2909, v_2910, v_2911, v_2912, v_2913, v_2914, v_2915, v_2916, v_2917, v_2918, v_2919, v_2920, v_2921, v_2922, v_2923, v_2924, v_2925, v_2926, v_2927, v_2928, v_2929, v_2930, v_2931, v_2932, v_2933, v_2934, v_2935, v_2936, v_2937, v_2938, v_2939, v_2940, v_2941, v_2942, v_2943, v_2944, v_2945, v_2946, v_2947, v_2948, v_2949, v_2950, v_2951, v_2952, v_2953, v_2954, v_2955, v_2956, v_2957, v_2958, v_2959, v_2960, v_2961, v_2962, v_2963, v_2964, v_2965, v_2966, v_2967, v_2968, v_2969, v_2970, v_2971, v_2972, v_2973, v_2974, v_2975, v_2976, v_2977, v_2978, v_2979, v_2980, v_2981, v_2982, v_2983, v_2984, v_2985, v_2986, v_2987, v_2988, v_2989, v_2990, v_2991, v_2992, v_2993, v_2994, v_2995, v_2996, v_2997, v_2998, v_2999, v_3000, v_3001, v_3002, v_3003, v_3004, v_3005, v_3006, v_3007, v_3008, v_3009, v_3010, v_3011, v_3012, v_3013, v_3014, v_3015, v_3016, v_3017, v_3018, v_3019, v_3020, v_3021, v_3022, v_3023, v_3024, v_3025, v_3026, v_3027, v_3028, v_3029, v_3030, v_3031, v_3032, v_3033, v_3034, v_3035, v_3036, v_3037, v_3038, v_3039, v_3040, v_3041, v_3042, v_3043, v_3044, v_3045, v_3046, v_3047, v_3048, v_3049, v_3050, v_3051, v_3052, v_3053, v_3054, v_3055, v_3056, v_3057, v_3058, v_3059, v_3060, v_3061, v_3062, v_3063, v_3064, v_3065, v_3066, v_3067, v_3068, v_3069, v_3070, v_3071, v_3072, v_3073, v_3074, v_3075, v_3076, v_3077, v_3078, v_3079, v_3080, v_3081, v_3082, v_3083, v_3084, v_3085, v_3086, v_3087, v_3088, v_3089, v_3090, v_3091, v_3092, v_3093, v_3094, v_3095, v_3096, v_3097, v_3098, v_3099, v_3100, v_3101, v_3102, v_3103, v_3104, v_3105, v_3106, v_3107, v_3108, v_3109, v_3110, v_3111, v_3112, v_3113, v_3114, v_3115, v_3116, v_3117, v_3118, v_3119, v_3120, v_3121, v_3122, v_3123, v_3124, v_3125, v_3126, v_3127, v_3128, v_3129, v_3130, v_3131, v_3132, v_3133, v_3134, v_3135, v_3136, v_3137, v_3138, v_3139, v_3140, v_3141, v_3142, v_3143, v_3144, v_3145, v_3146, v_3147, v_3148, v_3149, v_3150, v_3151, v_3152, v_3153, v_3154, v_3155, v_3156, v_3157, v_3158, v_3159, v_3160, v_3161, v_3162, v_3163, v_3164, v_3165, v_3166, v_3167, v_3168, v_3169, v_3170, v_3171, v_3172, v_3173, v_3174, v_3175, v_3176, v_3177, v_3178, v_3179, v_3180, v_3181, v_3182, v_3183, v_3184, v_3185, v_3186, v_3187, v_3188, v_3189, v_3190, v_3191, v_3192, v_3193, v_3194, v_3195, v_3196, v_3197, v_3198, v_3199, v_3200, v_3201, v_3202, v_3203, v_3204, v_3205, v_3206, v_3207, v_3208, v_3209, v_3210, v_3211, v_3212, v_3213, v_3214, v_3215, v_3216, v_3217, v_3218, v_3219, v_3220, v_3221, v_3222, v_3223, v_3224, v_3225, v_3226, v_3227, v_3228, v_3229, v_3230, v_3231, v_3232, v_3233, v_3234, v_3235, v_3236, v_3237, v_3238, v_3239, v_3240, v_3241, v_3242, v_3243, v_3244, v_3245, v_3246, v_3247, v_3248, v_3249, v_3250, v_3251, v_3252, v_3253, v_3254, v_3255, v_3256, v_3257, v_3258, v_3259, v_3260, v_3261, v_3262, v_3263, v_3264, v_3265, v_3266, v_3267, v_3268, v_3269, v_3270, v_3271, v_3272, v_3273, v_3274, v_3275, v_3276, v_3277, v_3278, v_3279, v_3280, v_3281, v_3282, v_3283, v_3284, v_3285, v_3286, v_3287, v_3288, v_3289, v_3290, v_3291, v_3292, v_3293, v_3294, v_3295, v_3296, v_3297, v_3298, v_3299, v_3300, v_3301, v_3302, v_3303, v_3304, v_3305, v_3306, v_3307, v_3308, v_3309, v_3310, v_3311, v_3312, v_3313, v_3314, v_3315, v_3316, v_3317, v_3318, v_3319, v_3320, v_3321, v_3322, v_3323, v_3324, v_3325, v_3326, v_3327, v_3328, v_3329, v_3330, v_3331, v_3332, v_3333, v_3334, v_3335, v_3336, v_3337, v_3338, v_3339, v_3340, v_3341, v_3342, v_3343, v_3344, v_3345, v_3346, v_3347, v_3348, v_3349, v_3350, v_3351, v_3352, v_3353, v_3354, v_3355, v_3356, v_3357, v_3358, v_3359, v_3360, v_3361, v_3362, v_3363, v_3364, v_3365, v_3366, v_3367, v_3368, v_3369, v_3370, v_3371, v_3372, v_3373, v_3374, v_3375, v_3376, v_3377, v_3378, v_3379, v_3380, o_1);
input v_1;
input v_2;
input v_3;
input v_4;
input v_5;
input v_6;
input v_7;
input v_8;
input v_9;
input v_10;
input v_11;
input v_12;
input v_13;
input v_14;
input v_15;
input v_16;
input v_17;
input v_18;
input v_19;
input v_20;
input v_21;
input v_22;
input v_23;
input v_24;
input v_25;
input v_27;
input v_28;
input v_29;
input v_30;
input v_31;
input v_32;
input v_33;
input v_34;
input v_35;
input v_36;
input v_37;
input v_38;
input v_39;
input v_40;
input v_41;
input v_42;
input v_43;
input v_44;
input v_45;
input v_46;
input v_47;
input v_48;
input v_49;
input v_50;
input v_51;
input v_52;
input v_53;
input v_54;
input v_55;
input v_56;
input v_57;
input v_58;
input v_59;
input v_60;
input v_61;
input v_62;
input v_63;
input v_64;
input v_65;
input v_66;
input v_67;
input v_68;
input v_69;
input v_70;
input v_71;
input v_72;
input v_73;
input v_74;
input v_75;
input v_76;
input v_77;
input v_78;
input v_79;
input v_80;
input v_81;
input v_82;
input v_83;
input v_84;
input v_85;
input v_86;
input v_87;
input v_88;
input v_89;
input v_90;
input v_91;
input v_92;
input v_93;
input v_94;
input v_95;
input v_96;
input v_100;
input v_101;
input v_102;
input v_103;
input v_104;
input v_105;
input v_106;
input v_107;
input v_108;
input v_109;
input v_110;
input v_111;
input v_112;
input v_113;
input v_117;
input v_120;
input v_121;
input v_122;
input v_126;
input v_127;
input v_128;
input v_131;
input v_132;
input v_26;
input v_97;
input v_98;
input v_99;
input v_114;
input v_115;
input v_116;
input v_118;
input v_119;
input v_123;
input v_124;
input v_125;
input v_129;
input v_130;
input v_133;
input v_134;
input v_135;
input v_136;
input v_137;
input v_138;
input v_139;
input v_140;
input v_141;
input v_142;
input v_143;
input v_144;
input v_145;
input v_146;
input v_147;
input v_148;
input v_149;
input v_150;
input v_151;
input v_152;
input v_153;
input v_154;
input v_155;
input v_156;
input v_157;
input v_158;
input v_159;
input v_160;
input v_161;
input v_162;
input v_163;
input v_164;
input v_165;
input v_166;
input v_167;
input v_168;
input v_169;
input v_170;
input v_171;
input v_172;
input v_173;
input v_174;
input v_175;
input v_176;
input v_177;
input v_178;
input v_179;
input v_180;
input v_181;
input v_182;
input v_183;
input v_184;
input v_185;
input v_186;
input v_187;
input v_188;
input v_189;
input v_190;
input v_191;
input v_192;
input v_193;
input v_194;
input v_195;
input v_196;
input v_197;
input v_198;
input v_199;
input v_200;
input v_201;
input v_202;
input v_203;
input v_204;
input v_205;
input v_206;
input v_207;
input v_208;
input v_209;
input v_210;
input v_211;
input v_212;
input v_213;
input v_214;
input v_215;
input v_216;
input v_217;
input v_218;
input v_219;
input v_220;
input v_221;
input v_222;
input v_223;
input v_224;
input v_225;
input v_226;
input v_227;
input v_228;
input v_229;
input v_230;
input v_231;
input v_232;
input v_233;
input v_234;
input v_235;
input v_236;
input v_237;
input v_238;
input v_239;
input v_240;
input v_241;
input v_242;
input v_243;
input v_244;
input v_245;
input v_246;
input v_247;
input v_248;
input v_249;
input v_250;
input v_251;
input v_252;
input v_253;
input v_254;
input v_255;
input v_256;
input v_257;
input v_258;
input v_259;
input v_260;
input v_261;
input v_262;
input v_263;
input v_264;
input v_265;
input v_266;
input v_267;
input v_268;
input v_269;
input v_270;
input v_271;
input v_272;
input v_273;
input v_274;
input v_275;
input v_276;
input v_277;
input v_278;
input v_279;
input v_280;
input v_281;
input v_282;
input v_283;
input v_284;
input v_285;
input v_286;
input v_287;
input v_288;
input v_289;
input v_290;
input v_291;
input v_292;
input v_293;
input v_294;
input v_295;
input v_296;
input v_297;
input v_298;
input v_299;
input v_300;
input v_301;
input v_302;
input v_303;
input v_304;
input v_305;
input v_306;
input v_307;
input v_308;
input v_309;
input v_310;
input v_311;
input v_312;
input v_313;
input v_314;
input v_315;
input v_316;
input v_317;
input v_318;
input v_319;
input v_320;
input v_321;
input v_322;
input v_323;
input v_324;
input v_325;
input v_326;
input v_327;
input v_328;
input v_329;
input v_330;
input v_331;
input v_332;
input v_333;
input v_334;
input v_335;
input v_336;
input v_337;
input v_338;
input v_339;
input v_340;
input v_341;
input v_342;
input v_343;
input v_344;
input v_345;
input v_346;
input v_347;
input v_348;
input v_349;
input v_350;
input v_351;
input v_352;
input v_353;
input v_354;
input v_355;
input v_356;
input v_357;
input v_358;
input v_359;
input v_360;
input v_361;
input v_362;
input v_363;
input v_364;
input v_365;
input v_366;
input v_367;
input v_368;
input v_369;
input v_370;
input v_371;
input v_372;
input v_373;
input v_374;
input v_375;
input v_376;
input v_377;
input v_378;
input v_379;
input v_380;
input v_381;
input v_382;
input v_383;
input v_384;
input v_385;
input v_386;
input v_387;
input v_388;
input v_389;
input v_390;
input v_391;
input v_392;
input v_393;
input v_394;
input v_395;
input v_396;
input v_397;
input v_398;
input v_399;
input v_400;
input v_401;
input v_402;
input v_403;
input v_404;
input v_405;
input v_406;
input v_407;
input v_408;
input v_409;
input v_410;
input v_411;
input v_412;
input v_413;
input v_414;
input v_415;
input v_416;
input v_417;
input v_418;
input v_419;
input v_420;
input v_421;
input v_422;
input v_423;
input v_424;
input v_425;
input v_426;
input v_427;
input v_428;
input v_429;
input v_430;
input v_431;
input v_432;
input v_433;
input v_434;
input v_435;
input v_436;
input v_437;
input v_438;
input v_439;
input v_440;
input v_441;
input v_442;
input v_443;
input v_444;
input v_445;
input v_446;
input v_447;
input v_448;
input v_449;
input v_450;
input v_451;
input v_452;
input v_453;
input v_454;
input v_455;
input v_456;
input v_457;
input v_458;
input v_459;
input v_460;
input v_461;
input v_462;
input v_463;
input v_464;
input v_465;
input v_466;
input v_467;
input v_468;
input v_469;
input v_470;
input v_471;
input v_472;
input v_473;
input v_474;
input v_475;
input v_476;
input v_477;
input v_478;
input v_479;
input v_480;
input v_481;
input v_482;
input v_483;
input v_484;
input v_485;
input v_486;
input v_487;
input v_488;
input v_489;
input v_490;
input v_491;
input v_492;
input v_493;
input v_494;
input v_495;
input v_496;
input v_497;
input v_498;
input v_499;
input v_500;
input v_501;
input v_502;
input v_503;
input v_504;
input v_505;
input v_506;
input v_507;
input v_508;
input v_509;
input v_510;
input v_511;
input v_512;
input v_513;
input v_514;
input v_515;
input v_516;
input v_517;
input v_518;
input v_519;
input v_520;
input v_521;
input v_522;
input v_523;
input v_524;
input v_525;
input v_526;
input v_527;
input v_528;
input v_529;
input v_530;
input v_531;
input v_532;
input v_533;
input v_534;
input v_535;
input v_536;
input v_537;
input v_538;
input v_539;
input v_540;
input v_541;
input v_542;
input v_543;
input v_544;
input v_545;
input v_546;
input v_547;
input v_548;
input v_549;
input v_550;
input v_551;
input v_552;
input v_553;
input v_554;
input v_555;
input v_556;
input v_557;
input v_558;
input v_559;
input v_560;
input v_561;
input v_562;
input v_563;
input v_564;
input v_565;
input v_566;
input v_567;
input v_568;
input v_569;
input v_570;
input v_571;
input v_572;
input v_573;
input v_574;
input v_575;
input v_576;
input v_577;
input v_578;
input v_579;
input v_580;
input v_581;
input v_582;
input v_583;
input v_584;
input v_585;
input v_586;
input v_587;
input v_588;
input v_589;
input v_590;
input v_591;
input v_592;
input v_593;
input v_594;
input v_595;
input v_596;
input v_597;
input v_598;
input v_599;
input v_600;
input v_601;
input v_602;
input v_603;
input v_604;
input v_605;
input v_606;
input v_607;
input v_608;
input v_609;
input v_610;
input v_611;
input v_612;
input v_613;
input v_614;
input v_615;
input v_616;
input v_617;
input v_618;
input v_619;
input v_620;
input v_621;
input v_622;
input v_623;
input v_624;
input v_625;
input v_626;
input v_627;
input v_628;
input v_629;
input v_630;
input v_631;
input v_632;
input v_633;
input v_634;
input v_635;
input v_636;
input v_637;
input v_638;
input v_639;
input v_640;
input v_641;
input v_642;
input v_643;
input v_644;
input v_645;
input v_646;
input v_647;
input v_648;
input v_649;
input v_650;
input v_651;
input v_652;
input v_653;
input v_654;
input v_655;
input v_656;
input v_657;
input v_658;
input v_659;
input v_660;
input v_661;
input v_662;
input v_663;
input v_664;
input v_665;
input v_666;
input v_667;
input v_668;
input v_669;
input v_670;
input v_671;
input v_672;
input v_673;
input v_674;
input v_675;
input v_676;
input v_677;
input v_678;
input v_679;
input v_680;
input v_681;
input v_682;
input v_683;
input v_684;
input v_685;
input v_686;
input v_687;
input v_688;
input v_689;
input v_690;
input v_691;
input v_692;
input v_693;
input v_694;
input v_695;
input v_696;
input v_697;
input v_698;
input v_699;
input v_700;
input v_701;
input v_702;
input v_703;
input v_704;
input v_705;
input v_706;
input v_707;
input v_708;
input v_709;
input v_710;
input v_711;
input v_712;
input v_713;
input v_714;
input v_715;
input v_716;
input v_717;
input v_718;
input v_719;
input v_720;
input v_721;
input v_722;
input v_723;
input v_724;
input v_725;
input v_726;
input v_727;
input v_728;
input v_729;
input v_730;
input v_731;
input v_732;
input v_733;
input v_734;
input v_735;
input v_736;
input v_737;
input v_738;
input v_739;
input v_740;
input v_741;
input v_742;
input v_743;
input v_744;
input v_745;
input v_746;
input v_747;
input v_748;
input v_749;
input v_750;
input v_751;
input v_752;
input v_753;
input v_754;
input v_755;
input v_756;
input v_757;
input v_758;
input v_759;
input v_760;
input v_761;
input v_762;
input v_763;
input v_764;
input v_765;
input v_766;
input v_767;
input v_768;
input v_769;
input v_770;
input v_771;
input v_772;
input v_773;
input v_774;
input v_775;
input v_776;
input v_777;
input v_778;
input v_779;
input v_780;
input v_781;
input v_782;
input v_783;
input v_784;
input v_785;
input v_786;
input v_787;
input v_788;
input v_789;
input v_790;
input v_791;
input v_792;
input v_793;
input v_794;
input v_795;
input v_796;
input v_797;
input v_798;
input v_799;
input v_800;
input v_801;
input v_802;
input v_803;
input v_804;
input v_805;
input v_806;
input v_807;
input v_808;
input v_809;
input v_810;
input v_811;
input v_812;
input v_813;
input v_814;
input v_815;
input v_816;
input v_817;
input v_818;
input v_819;
input v_820;
input v_821;
input v_822;
input v_823;
input v_824;
input v_825;
input v_826;
input v_827;
input v_828;
input v_829;
input v_830;
input v_831;
input v_832;
input v_833;
input v_834;
input v_835;
input v_836;
input v_837;
input v_838;
input v_839;
input v_840;
input v_841;
input v_842;
input v_843;
input v_844;
input v_845;
input v_846;
input v_847;
input v_848;
input v_849;
input v_850;
input v_851;
input v_852;
input v_853;
input v_854;
input v_855;
input v_856;
input v_857;
input v_858;
input v_859;
input v_860;
input v_861;
input v_862;
input v_863;
input v_864;
input v_865;
input v_866;
input v_867;
input v_868;
input v_869;
input v_870;
input v_871;
input v_872;
input v_873;
input v_874;
input v_875;
input v_876;
input v_877;
input v_878;
input v_879;
input v_880;
input v_881;
input v_882;
input v_883;
input v_884;
input v_885;
input v_886;
input v_887;
input v_888;
input v_889;
input v_890;
input v_891;
input v_892;
input v_893;
input v_894;
input v_895;
input v_896;
input v_897;
input v_898;
input v_899;
input v_900;
input v_901;
input v_902;
input v_903;
input v_904;
input v_905;
input v_906;
input v_907;
input v_908;
input v_909;
input v_910;
input v_911;
input v_912;
input v_913;
input v_914;
input v_915;
input v_916;
input v_917;
input v_918;
input v_919;
input v_920;
input v_921;
input v_922;
input v_923;
input v_924;
input v_925;
input v_926;
input v_927;
input v_928;
input v_929;
input v_930;
input v_931;
input v_932;
input v_933;
input v_934;
input v_935;
input v_936;
input v_937;
input v_938;
input v_939;
input v_940;
input v_941;
input v_942;
input v_943;
input v_944;
input v_945;
input v_946;
input v_947;
input v_948;
input v_949;
input v_950;
input v_951;
input v_952;
input v_953;
input v_954;
input v_955;
input v_956;
input v_957;
input v_958;
input v_959;
input v_960;
input v_961;
input v_962;
input v_963;
input v_964;
input v_965;
input v_966;
input v_967;
input v_968;
input v_969;
input v_970;
input v_971;
input v_972;
input v_973;
input v_974;
input v_975;
input v_976;
input v_977;
input v_978;
input v_979;
input v_980;
input v_981;
input v_982;
input v_983;
input v_984;
input v_985;
input v_986;
input v_987;
input v_988;
input v_989;
input v_990;
input v_991;
input v_992;
input v_993;
input v_994;
input v_995;
input v_996;
input v_997;
input v_998;
input v_999;
input v_1000;
input v_1001;
input v_1002;
input v_1003;
input v_1004;
input v_1005;
input v_1006;
input v_1007;
input v_1008;
input v_1009;
input v_1010;
input v_1011;
input v_1012;
input v_1013;
input v_1014;
input v_1015;
input v_1016;
input v_1017;
input v_1018;
input v_1019;
input v_1020;
input v_1021;
input v_1022;
input v_1023;
input v_1024;
input v_1025;
input v_1026;
input v_1027;
input v_1028;
input v_1029;
input v_1030;
input v_1031;
input v_1032;
input v_1033;
input v_1034;
input v_1035;
input v_1036;
input v_1037;
input v_1038;
input v_1039;
input v_1040;
input v_1041;
input v_1042;
input v_1043;
input v_1044;
input v_1045;
input v_1046;
input v_1047;
input v_1048;
input v_1049;
input v_1050;
input v_1051;
input v_1052;
input v_1053;
input v_1054;
input v_1055;
input v_1056;
input v_1057;
input v_1058;
input v_1059;
input v_1060;
input v_1061;
input v_1062;
input v_1063;
input v_1064;
input v_1065;
input v_1066;
input v_1067;
input v_1068;
input v_1069;
input v_1070;
input v_1071;
input v_1072;
input v_1073;
input v_1074;
input v_1075;
input v_1076;
input v_1077;
input v_1078;
input v_1079;
input v_1080;
input v_1081;
input v_1082;
input v_1083;
input v_1084;
input v_1085;
input v_1086;
input v_1087;
input v_1088;
input v_1089;
input v_1090;
input v_1091;
input v_1092;
input v_1093;
input v_1094;
input v_1095;
input v_1096;
input v_1097;
input v_1098;
input v_1099;
input v_1100;
input v_1101;
input v_1102;
input v_1103;
input v_1104;
input v_1105;
input v_1106;
input v_1107;
input v_1108;
input v_1109;
input v_1110;
input v_1111;
input v_1112;
input v_1113;
input v_1114;
input v_1115;
input v_1116;
input v_1117;
input v_1118;
input v_1119;
input v_1120;
input v_1121;
input v_1122;
input v_1123;
input v_1124;
input v_1125;
input v_1126;
input v_1127;
input v_1128;
input v_1129;
input v_1130;
input v_1131;
input v_1132;
input v_1133;
input v_1134;
input v_1135;
input v_1136;
input v_1137;
input v_1138;
input v_1139;
input v_1140;
input v_1141;
input v_1142;
input v_1143;
input v_1144;
input v_1145;
input v_1146;
input v_1147;
input v_1148;
input v_1149;
input v_1150;
input v_1151;
input v_1152;
input v_1153;
input v_1154;
input v_1155;
input v_1156;
input v_1157;
input v_1158;
input v_1159;
input v_1160;
input v_1161;
input v_1162;
input v_1163;
input v_1164;
input v_1165;
input v_1166;
input v_1167;
input v_1168;
input v_1169;
input v_1170;
input v_1171;
input v_1172;
input v_1173;
input v_1174;
input v_1175;
input v_1176;
input v_1177;
input v_1178;
input v_1179;
input v_1180;
input v_1181;
input v_1182;
input v_1183;
input v_1184;
input v_1185;
input v_1186;
input v_1187;
input v_1188;
input v_1189;
input v_1190;
input v_1191;
input v_1192;
input v_1193;
input v_1194;
input v_1195;
input v_1196;
input v_1197;
input v_1198;
input v_1199;
input v_1200;
input v_1201;
input v_1202;
input v_1203;
input v_1204;
input v_1205;
input v_1206;
input v_1207;
input v_1208;
input v_1209;
input v_1210;
input v_1211;
input v_1212;
input v_1213;
input v_1214;
input v_1215;
input v_1216;
input v_1217;
input v_1218;
input v_1219;
input v_1220;
input v_1221;
input v_1222;
input v_1223;
input v_1224;
input v_1225;
input v_1226;
input v_1227;
input v_1228;
input v_1229;
input v_1230;
input v_1231;
input v_1232;
input v_1233;
input v_1234;
input v_1235;
input v_1236;
input v_1237;
input v_1238;
input v_1239;
input v_1240;
input v_1241;
input v_1242;
input v_1243;
input v_1244;
input v_1245;
input v_1246;
input v_1247;
input v_1248;
input v_1249;
input v_1250;
input v_1251;
input v_1252;
input v_1253;
input v_1254;
input v_1255;
input v_1256;
input v_1257;
input v_1258;
input v_1259;
input v_1260;
input v_1261;
input v_1262;
input v_1263;
input v_1264;
input v_1265;
input v_1266;
input v_1267;
input v_1268;
input v_1269;
input v_1270;
input v_1271;
input v_1272;
input v_1273;
input v_1274;
input v_1275;
input v_1276;
input v_1277;
input v_1278;
input v_1279;
input v_1280;
input v_1281;
input v_1282;
input v_1283;
input v_1284;
input v_1285;
input v_1286;
input v_1287;
input v_1288;
input v_1289;
input v_1290;
input v_1291;
input v_1292;
input v_1293;
input v_1294;
input v_1295;
input v_1296;
input v_1297;
input v_1298;
input v_1299;
input v_1300;
input v_1301;
input v_1302;
input v_1303;
input v_1304;
input v_1305;
input v_1306;
input v_1307;
input v_1308;
input v_1309;
input v_1310;
input v_1311;
input v_1312;
input v_1313;
input v_1314;
input v_1315;
input v_1316;
input v_1317;
input v_1318;
input v_1319;
input v_1320;
input v_1321;
input v_1322;
input v_1323;
input v_1324;
input v_1325;
input v_1326;
input v_1327;
input v_1328;
input v_1329;
input v_1330;
input v_1331;
input v_1332;
input v_1333;
input v_1334;
input v_1335;
input v_1336;
input v_1337;
input v_1338;
input v_1339;
input v_1340;
input v_1341;
input v_1342;
input v_1343;
input v_1344;
input v_1345;
input v_1346;
input v_1347;
input v_1348;
input v_1349;
input v_1350;
input v_1351;
input v_1352;
input v_1353;
input v_1354;
input v_1355;
input v_1356;
input v_1357;
input v_1358;
input v_1359;
input v_1360;
input v_1361;
input v_1362;
input v_1363;
input v_1364;
input v_1365;
input v_1366;
input v_1367;
input v_1368;
input v_1369;
input v_1370;
input v_1371;
input v_1372;
input v_1373;
input v_1374;
input v_1375;
input v_1376;
input v_1377;
input v_1378;
input v_1379;
input v_1380;
input v_1381;
input v_1382;
input v_1383;
input v_1384;
input v_1385;
input v_1386;
input v_1387;
input v_1388;
input v_1389;
input v_1390;
input v_1391;
input v_1392;
input v_1393;
input v_1394;
input v_1395;
input v_1396;
input v_1397;
input v_1398;
input v_1399;
input v_1400;
input v_1401;
input v_1402;
input v_1403;
input v_1404;
input v_1405;
input v_1406;
input v_1407;
input v_1408;
input v_1409;
input v_1410;
input v_1411;
input v_1412;
input v_1413;
input v_1414;
input v_1415;
input v_1416;
input v_1417;
input v_1418;
input v_1419;
input v_1420;
input v_1421;
input v_1422;
input v_1423;
input v_1424;
input v_1425;
input v_1426;
input v_1427;
input v_1428;
input v_1429;
input v_1430;
input v_1431;
input v_1432;
input v_1433;
input v_1434;
input v_1435;
input v_1436;
input v_1437;
input v_1438;
input v_1439;
input v_1440;
input v_1441;
input v_1442;
input v_1443;
input v_1444;
input v_1445;
input v_1446;
input v_1447;
input v_1448;
input v_1449;
input v_1450;
input v_1451;
input v_1452;
input v_1453;
input v_1454;
input v_1455;
input v_1456;
input v_1457;
input v_1458;
input v_1459;
input v_1460;
input v_1461;
input v_1462;
input v_1463;
input v_1464;
input v_1465;
input v_1466;
input v_1467;
input v_1468;
input v_1469;
input v_1470;
input v_1471;
input v_1472;
input v_1473;
input v_1474;
input v_1475;
input v_1476;
input v_1477;
input v_1478;
input v_1479;
input v_1480;
input v_1481;
input v_1482;
input v_1483;
input v_1484;
input v_1485;
input v_1486;
input v_1487;
input v_1488;
input v_1489;
input v_1490;
input v_1491;
input v_1492;
input v_1493;
input v_1494;
input v_1495;
input v_1496;
input v_1497;
input v_1498;
input v_1499;
input v_1500;
input v_1501;
input v_1502;
input v_1503;
input v_1504;
input v_1505;
input v_1506;
input v_1507;
input v_1508;
input v_1509;
input v_1510;
input v_1511;
input v_1512;
input v_1513;
input v_1514;
input v_1515;
input v_1516;
input v_1517;
input v_1518;
input v_1519;
input v_1520;
input v_1521;
input v_1522;
input v_1523;
input v_1524;
input v_1525;
input v_1526;
input v_1527;
input v_1528;
input v_1529;
input v_1530;
input v_1531;
input v_1532;
input v_1533;
input v_1534;
input v_1535;
input v_1536;
input v_1537;
input v_1538;
input v_1539;
input v_1540;
input v_1541;
input v_1542;
input v_1543;
input v_1544;
input v_1545;
input v_1546;
input v_1547;
input v_1548;
input v_1549;
input v_1550;
input v_1551;
input v_1552;
input v_1553;
input v_1554;
input v_1555;
input v_1556;
input v_1557;
input v_1558;
input v_1559;
input v_1560;
input v_1561;
input v_1562;
input v_1563;
input v_1564;
input v_1565;
input v_1566;
input v_1567;
input v_1568;
input v_1569;
input v_1570;
input v_1571;
input v_1572;
input v_1573;
input v_1574;
input v_1575;
input v_1576;
input v_1577;
input v_1578;
input v_1579;
input v_1580;
input v_1581;
input v_1582;
input v_1583;
input v_1584;
input v_1585;
input v_1586;
input v_1587;
input v_1588;
input v_1589;
input v_1590;
input v_1591;
input v_1592;
input v_1593;
input v_1594;
input v_1595;
input v_1596;
input v_1597;
input v_1598;
input v_1599;
input v_1600;
input v_1601;
input v_1602;
input v_1603;
input v_1604;
input v_1605;
input v_1606;
input v_1607;
input v_1608;
input v_1609;
input v_1610;
input v_1611;
input v_1612;
input v_1613;
input v_1614;
input v_1615;
input v_1616;
input v_1617;
input v_1618;
input v_1619;
input v_1620;
input v_1621;
input v_1622;
input v_1623;
input v_1624;
input v_1625;
input v_1626;
input v_1627;
input v_1628;
input v_1629;
input v_1630;
input v_1631;
input v_1632;
input v_1633;
input v_1634;
input v_1635;
input v_1636;
input v_1637;
input v_1638;
input v_1639;
input v_1640;
input v_1641;
input v_1642;
input v_1643;
input v_1644;
input v_1645;
input v_1646;
input v_1647;
input v_1648;
input v_1649;
input v_1650;
input v_1651;
input v_1652;
input v_1653;
input v_1654;
input v_1655;
input v_1656;
input v_1657;
input v_1658;
input v_1659;
input v_1660;
input v_1661;
input v_1662;
input v_1663;
input v_1664;
input v_1665;
input v_1666;
input v_1667;
input v_1668;
input v_1669;
input v_1670;
input v_1671;
input v_1672;
input v_1673;
input v_1674;
input v_1675;
input v_1676;
input v_1677;
input v_1678;
input v_1679;
input v_1680;
input v_1681;
input v_1682;
input v_1683;
input v_1684;
input v_1685;
input v_1686;
input v_1687;
input v_1688;
input v_1689;
input v_1690;
input v_1691;
input v_1692;
input v_1693;
input v_1694;
input v_1695;
input v_1696;
input v_1697;
input v_1698;
input v_1699;
input v_1700;
input v_1701;
input v_1702;
input v_1703;
input v_1704;
input v_1705;
input v_1706;
input v_1707;
input v_1708;
input v_1709;
input v_1710;
input v_1711;
input v_1712;
input v_1713;
input v_1714;
input v_1715;
input v_1716;
input v_1717;
input v_1718;
input v_1719;
input v_1720;
input v_1721;
input v_1722;
input v_1723;
input v_1724;
input v_1725;
input v_1726;
input v_1727;
input v_1728;
input v_1729;
input v_1730;
input v_1731;
input v_1732;
input v_1733;
input v_1734;
input v_1735;
input v_1736;
input v_1737;
input v_1738;
input v_1739;
input v_1740;
input v_1741;
input v_1742;
input v_1743;
input v_1744;
input v_1745;
input v_1746;
input v_1747;
input v_1748;
input v_1749;
input v_1750;
input v_1751;
input v_1752;
input v_1753;
input v_1754;
input v_1755;
input v_1756;
input v_1757;
input v_1758;
input v_1759;
input v_1760;
input v_1761;
input v_1762;
input v_1763;
input v_1764;
input v_1765;
input v_1766;
input v_1767;
input v_1768;
input v_1769;
input v_1770;
input v_1771;
input v_1772;
input v_1773;
input v_1774;
input v_1775;
input v_1776;
input v_1777;
input v_1778;
input v_1779;
input v_1780;
input v_1781;
input v_1782;
input v_1783;
input v_1784;
input v_1785;
input v_1786;
input v_1787;
input v_1788;
input v_1789;
input v_1790;
input v_1791;
input v_1792;
input v_1793;
input v_1794;
input v_1795;
input v_1796;
input v_1797;
input v_1798;
input v_1799;
input v_1800;
input v_1801;
input v_1802;
input v_1803;
input v_1804;
input v_1805;
input v_1806;
input v_1807;
input v_1808;
input v_1809;
input v_1810;
input v_1811;
input v_1812;
input v_1813;
input v_1814;
input v_1815;
input v_1816;
input v_1817;
input v_1818;
input v_1819;
input v_1820;
input v_1821;
input v_1822;
input v_1823;
input v_1824;
input v_1825;
input v_1826;
input v_1827;
input v_1828;
input v_1829;
input v_1830;
input v_1831;
input v_1832;
input v_1833;
input v_1834;
input v_1835;
input v_1836;
input v_1837;
input v_1838;
input v_1839;
input v_1840;
input v_1841;
input v_1842;
input v_1843;
input v_1844;
input v_1845;
input v_1846;
input v_1847;
input v_1848;
input v_1849;
input v_1850;
input v_1851;
input v_1852;
input v_1853;
input v_1854;
input v_1855;
input v_1856;
input v_1857;
input v_1858;
input v_1859;
input v_1860;
input v_1861;
input v_1862;
input v_1863;
input v_1864;
input v_1865;
input v_1866;
input v_1867;
input v_1868;
input v_1869;
input v_1870;
input v_1871;
input v_1872;
input v_1873;
input v_1874;
input v_1875;
input v_1876;
input v_1877;
input v_1878;
input v_1879;
input v_1880;
input v_1881;
input v_1882;
input v_1883;
input v_1884;
input v_1885;
input v_1886;
input v_1887;
input v_1888;
input v_1889;
input v_1890;
input v_1891;
input v_1892;
input v_1893;
input v_1894;
input v_1895;
input v_1896;
input v_1897;
input v_1898;
input v_1899;
input v_1900;
input v_1901;
input v_1902;
input v_1903;
input v_1904;
input v_1905;
input v_1906;
input v_1907;
input v_1908;
input v_1909;
input v_1910;
input v_1911;
input v_1912;
input v_1913;
input v_1914;
input v_1915;
input v_1916;
input v_1917;
input v_1918;
input v_1919;
input v_1920;
input v_1921;
input v_1922;
input v_1923;
input v_1924;
input v_1925;
input v_1926;
input v_1927;
input v_1928;
input v_1929;
input v_1930;
input v_1931;
input v_1932;
input v_1933;
input v_1934;
input v_1935;
input v_1936;
input v_1937;
input v_1938;
input v_1939;
input v_1940;
input v_1941;
input v_1942;
input v_1943;
input v_1944;
input v_1945;
input v_1946;
input v_1947;
input v_1948;
input v_1949;
input v_1950;
input v_1951;
input v_1952;
input v_1953;
input v_1954;
input v_1955;
input v_1956;
input v_1957;
input v_1958;
input v_1959;
input v_1960;
input v_1961;
input v_1962;
input v_1963;
input v_1964;
input v_1965;
input v_1966;
input v_1967;
input v_1968;
input v_1969;
input v_1970;
input v_1971;
input v_1972;
input v_1973;
input v_1974;
input v_1975;
input v_1976;
input v_1977;
input v_1978;
input v_1979;
input v_1980;
input v_1981;
input v_1982;
input v_1983;
input v_1984;
input v_1985;
input v_1986;
input v_1987;
input v_1988;
input v_1989;
input v_1990;
input v_1991;
input v_1992;
input v_1993;
input v_1994;
input v_1995;
input v_1996;
input v_1997;
input v_1998;
input v_1999;
input v_2000;
input v_2001;
input v_2002;
input v_2003;
input v_2004;
input v_2005;
input v_2006;
input v_2007;
input v_2008;
input v_2009;
input v_2010;
input v_2011;
input v_2012;
input v_2013;
input v_2014;
input v_2015;
input v_2016;
input v_2017;
input v_2018;
input v_2019;
input v_2020;
input v_2021;
input v_2022;
input v_2023;
input v_2024;
input v_2025;
input v_2026;
input v_2027;
input v_2028;
input v_2029;
input v_2030;
input v_2031;
input v_2032;
input v_2033;
input v_2034;
input v_2035;
input v_2036;
input v_2037;
input v_2038;
input v_2039;
input v_2040;
input v_2041;
input v_2042;
input v_2043;
input v_2044;
input v_2045;
input v_2046;
input v_2047;
input v_2048;
input v_2049;
input v_2050;
input v_2051;
input v_2052;
input v_2053;
input v_2054;
input v_2055;
input v_2056;
input v_2057;
input v_2058;
input v_2059;
input v_2060;
input v_2061;
input v_2062;
input v_2063;
input v_2064;
input v_2065;
input v_2066;
input v_2067;
input v_2068;
input v_2069;
input v_2070;
input v_2071;
input v_2072;
input v_2073;
input v_2074;
input v_2075;
input v_2076;
input v_2077;
input v_2078;
input v_2079;
input v_2080;
input v_2081;
input v_2082;
input v_2083;
input v_2084;
input v_2085;
input v_2086;
input v_2087;
input v_2088;
input v_2089;
input v_2090;
input v_2091;
input v_2092;
input v_2093;
input v_2094;
input v_2095;
input v_2096;
input v_2097;
input v_2098;
input v_2099;
input v_2100;
input v_2101;
input v_2102;
input v_2103;
input v_2104;
input v_2105;
input v_2106;
input v_2107;
input v_2108;
input v_2109;
input v_2110;
input v_2111;
input v_2112;
input v_2113;
input v_2114;
input v_2115;
input v_2116;
input v_2117;
input v_2118;
input v_2119;
input v_2120;
input v_2121;
input v_2122;
input v_2123;
input v_2124;
input v_2125;
input v_2126;
input v_2127;
input v_2128;
input v_2129;
input v_2130;
input v_2131;
input v_2132;
input v_2133;
input v_2134;
input v_2135;
input v_2136;
input v_2137;
input v_2138;
input v_2139;
input v_2140;
input v_2141;
input v_2142;
input v_2143;
input v_2144;
input v_2145;
input v_2146;
input v_2147;
input v_2148;
input v_2149;
input v_2150;
input v_2151;
input v_2152;
input v_2153;
input v_2154;
input v_2155;
input v_2156;
input v_2157;
input v_2158;
input v_2159;
input v_2160;
input v_2161;
input v_2162;
input v_2163;
input v_2164;
input v_2165;
input v_2166;
input v_2167;
input v_2168;
input v_2169;
input v_2170;
input v_2171;
input v_2172;
input v_2173;
input v_2174;
input v_2175;
input v_2176;
input v_2177;
input v_2178;
input v_2179;
input v_2180;
input v_2181;
input v_2182;
input v_2183;
input v_2184;
input v_2185;
input v_2186;
input v_2187;
input v_2188;
input v_2189;
input v_2190;
input v_2191;
input v_2192;
input v_2193;
input v_2194;
input v_2195;
input v_2196;
input v_2197;
input v_2198;
input v_2199;
input v_2200;
input v_2201;
input v_2202;
input v_2203;
input v_2204;
input v_2205;
input v_2206;
input v_2207;
input v_2208;
input v_2209;
input v_2210;
input v_2211;
input v_2212;
input v_2213;
input v_2214;
input v_2215;
input v_2216;
input v_2217;
input v_2218;
input v_2219;
input v_2220;
input v_2221;
input v_2222;
input v_2223;
input v_2224;
input v_2225;
input v_2226;
input v_2227;
input v_2228;
input v_2229;
input v_2230;
input v_2231;
input v_2232;
input v_2233;
input v_2234;
input v_2235;
input v_2236;
input v_2237;
input v_2238;
input v_2239;
input v_2240;
input v_2241;
input v_2242;
input v_2243;
input v_2244;
input v_2245;
input v_2246;
input v_2247;
input v_2248;
input v_2249;
input v_2250;
input v_2251;
input v_2252;
input v_2253;
input v_2254;
input v_2255;
input v_2256;
input v_2257;
input v_2258;
input v_2259;
input v_2260;
input v_2261;
input v_2262;
input v_2263;
input v_2264;
input v_2265;
input v_2266;
input v_2267;
input v_2268;
input v_2269;
input v_2270;
input v_2271;
input v_2272;
input v_2273;
input v_2274;
input v_2275;
input v_2276;
input v_2277;
input v_2278;
input v_2279;
input v_2280;
input v_2281;
input v_2282;
input v_2283;
input v_2284;
input v_2285;
input v_2286;
input v_2287;
input v_2288;
input v_2289;
input v_2290;
input v_2291;
input v_2292;
input v_2293;
input v_2294;
input v_2295;
input v_2296;
input v_2297;
input v_2298;
input v_2299;
input v_2300;
input v_2301;
input v_2302;
input v_2303;
input v_2304;
input v_2305;
input v_2306;
input v_2307;
input v_2308;
input v_2309;
input v_2310;
input v_2311;
input v_2312;
input v_2313;
input v_2314;
input v_2315;
input v_2316;
input v_2317;
input v_2318;
input v_2319;
input v_2320;
input v_2321;
input v_2322;
input v_2323;
input v_2324;
input v_2325;
input v_2326;
input v_2327;
input v_2328;
input v_2329;
input v_2330;
input v_2331;
input v_2332;
input v_2333;
input v_2334;
input v_2335;
input v_2336;
input v_2337;
input v_2338;
input v_2339;
input v_2340;
input v_2341;
input v_2342;
input v_2343;
input v_2344;
input v_2345;
input v_2346;
input v_2347;
input v_2348;
input v_2349;
input v_2350;
input v_2351;
input v_2352;
input v_2353;
input v_2354;
input v_2355;
input v_2356;
input v_2357;
input v_2358;
input v_2359;
input v_2360;
input v_2361;
input v_2362;
input v_2363;
input v_2364;
input v_2365;
input v_2366;
input v_2367;
input v_2368;
input v_2369;
input v_2370;
input v_2371;
input v_2372;
input v_2373;
input v_2374;
input v_2375;
input v_2376;
input v_2377;
input v_2378;
input v_2379;
input v_2380;
input v_2381;
input v_2382;
input v_2383;
input v_2384;
input v_2385;
input v_2386;
input v_2387;
input v_2388;
input v_2389;
input v_2390;
input v_2391;
input v_2392;
input v_2393;
input v_2394;
input v_2395;
input v_2396;
input v_2397;
input v_2398;
input v_2399;
input v_2400;
input v_2401;
input v_2402;
input v_2403;
input v_2404;
input v_2405;
input v_2406;
input v_2407;
input v_2408;
input v_2409;
input v_2410;
input v_2411;
input v_2412;
input v_2413;
input v_2414;
input v_2415;
input v_2416;
input v_2417;
input v_2418;
input v_2419;
input v_2420;
input v_2421;
input v_2422;
input v_2423;
input v_2424;
input v_2425;
input v_2426;
input v_2427;
input v_2428;
input v_2429;
input v_2430;
input v_2431;
input v_2432;
input v_2433;
input v_2434;
input v_2435;
input v_2436;
input v_2437;
input v_2438;
input v_2439;
input v_2440;
input v_2441;
input v_2442;
input v_2443;
input v_2444;
input v_2445;
input v_2446;
input v_2447;
input v_2448;
input v_2449;
input v_2450;
input v_2451;
input v_2452;
input v_2453;
input v_2454;
input v_2455;
input v_2456;
input v_2457;
input v_2458;
input v_2459;
input v_2460;
input v_2461;
input v_2462;
input v_2463;
input v_2464;
input v_2465;
input v_2466;
input v_2467;
input v_2468;
input v_2469;
input v_2470;
input v_2471;
input v_2472;
input v_2473;
input v_2474;
input v_2475;
input v_2476;
input v_2477;
input v_2478;
input v_2479;
input v_2480;
input v_2481;
input v_2482;
input v_2483;
input v_2484;
input v_2485;
input v_2486;
input v_2487;
input v_2488;
input v_2489;
input v_2490;
input v_2491;
input v_2492;
input v_2493;
input v_2494;
input v_2495;
input v_2496;
input v_2497;
input v_2498;
input v_2499;
input v_2500;
input v_2501;
input v_2502;
input v_2503;
input v_2504;
input v_2505;
input v_2506;
input v_2507;
input v_2508;
input v_2509;
input v_2510;
input v_2511;
input v_2512;
input v_2513;
input v_2514;
input v_2515;
input v_2516;
input v_2517;
input v_2518;
input v_2519;
input v_2520;
input v_2521;
input v_2522;
input v_2523;
input v_2524;
input v_2525;
input v_2526;
input v_2527;
input v_2528;
input v_2529;
input v_2530;
input v_2531;
input v_2532;
input v_2533;
input v_2534;
input v_2535;
input v_2536;
input v_2537;
input v_2538;
input v_2539;
input v_2540;
input v_2541;
input v_2542;
input v_2543;
input v_2544;
input v_2545;
input v_2546;
input v_2547;
input v_2548;
input v_2549;
input v_2550;
input v_2551;
input v_2552;
input v_2553;
input v_2554;
input v_2555;
input v_2556;
input v_2557;
input v_2558;
input v_2559;
input v_2560;
input v_2561;
input v_2562;
input v_2563;
input v_2564;
input v_2565;
input v_2566;
input v_2567;
input v_2568;
input v_2569;
input v_2570;
input v_2571;
input v_2572;
input v_2573;
input v_2574;
input v_2575;
input v_2576;
input v_2577;
input v_2578;
input v_2579;
input v_2580;
input v_2581;
input v_2582;
input v_2583;
input v_2584;
input v_2585;
input v_2586;
input v_2587;
input v_2588;
input v_2589;
input v_2590;
input v_2591;
input v_2592;
input v_2593;
input v_2594;
input v_2595;
input v_2596;
input v_2597;
input v_2598;
input v_2599;
input v_2600;
input v_2601;
input v_2602;
input v_2603;
input v_2604;
input v_2605;
input v_2606;
input v_2607;
input v_2608;
input v_2609;
input v_2610;
input v_2611;
input v_2612;
input v_2613;
input v_2614;
input v_2615;
input v_2616;
input v_2617;
input v_2618;
input v_2619;
input v_2620;
input v_2621;
input v_2622;
input v_2623;
input v_2624;
input v_2625;
input v_2626;
input v_2627;
input v_2628;
input v_2629;
input v_2630;
input v_2631;
input v_2632;
input v_2633;
input v_2634;
input v_2635;
input v_2636;
input v_2637;
input v_2638;
input v_2639;
input v_2640;
input v_2641;
input v_2642;
input v_2643;
input v_2644;
input v_2645;
input v_2646;
input v_2647;
input v_2648;
input v_2649;
input v_2650;
input v_2651;
input v_2652;
input v_2653;
input v_2654;
input v_2655;
input v_2656;
input v_2657;
input v_2658;
input v_2659;
input v_2660;
input v_2661;
input v_2662;
input v_2663;
input v_2664;
input v_2665;
input v_2666;
input v_2667;
input v_2668;
input v_2669;
input v_2670;
input v_2671;
input v_2672;
input v_2673;
input v_2674;
input v_2675;
input v_2676;
input v_2677;
input v_2678;
input v_2679;
input v_2680;
input v_2681;
input v_2682;
input v_2683;
input v_2684;
input v_2685;
input v_2686;
input v_2687;
input v_2688;
input v_2689;
input v_2690;
input v_2691;
input v_2692;
input v_2693;
input v_2694;
input v_2695;
input v_2696;
input v_2697;
input v_2698;
input v_2699;
input v_2700;
input v_2701;
input v_2702;
input v_2703;
input v_2704;
input v_2705;
input v_2706;
input v_2707;
input v_2708;
input v_2709;
input v_2710;
input v_2711;
input v_2712;
input v_2713;
input v_2714;
input v_2715;
input v_2716;
input v_2717;
input v_2718;
input v_2719;
input v_2720;
input v_2721;
input v_2722;
input v_2723;
input v_2724;
input v_2725;
input v_2726;
input v_2727;
input v_2728;
input v_2729;
input v_2730;
input v_2731;
input v_2732;
input v_2733;
input v_2734;
input v_2735;
input v_2736;
input v_2737;
input v_2738;
input v_2739;
input v_2740;
input v_2741;
input v_2742;
input v_2743;
input v_2744;
input v_2745;
input v_2746;
input v_2747;
input v_2748;
input v_2749;
input v_2750;
input v_2751;
input v_2752;
input v_2753;
input v_2754;
input v_2755;
input v_2756;
input v_2757;
input v_2758;
input v_2759;
input v_2760;
input v_2761;
input v_2762;
input v_2763;
input v_2764;
input v_2765;
input v_2766;
input v_2767;
input v_2768;
input v_2769;
input v_2770;
input v_2771;
input v_2772;
input v_2773;
input v_2774;
input v_2775;
input v_2776;
input v_2777;
input v_2778;
input v_2779;
input v_2780;
input v_2781;
input v_2782;
input v_2783;
input v_2784;
input v_2785;
input v_2786;
input v_2787;
input v_2788;
input v_2789;
input v_2790;
input v_2791;
input v_2792;
input v_2793;
input v_2794;
input v_2795;
input v_2796;
input v_2797;
input v_2798;
input v_2799;
input v_2800;
input v_2801;
input v_2802;
input v_2803;
input v_2804;
input v_2805;
input v_2806;
input v_2807;
input v_2808;
input v_2809;
input v_2810;
input v_2811;
input v_2812;
input v_2813;
input v_2814;
input v_2815;
input v_2816;
input v_2817;
input v_2818;
input v_2819;
input v_2820;
input v_2821;
input v_2822;
input v_2823;
input v_2824;
input v_2825;
input v_2826;
input v_2827;
input v_2828;
input v_2829;
input v_2830;
input v_2831;
input v_2832;
input v_2833;
input v_2834;
input v_2835;
input v_2836;
input v_2837;
input v_2838;
input v_2839;
input v_2840;
input v_2841;
input v_2842;
input v_2843;
input v_2844;
input v_2845;
input v_2846;
input v_2847;
input v_2848;
input v_2849;
input v_2850;
input v_2851;
input v_2852;
input v_2853;
input v_2854;
input v_2855;
input v_2856;
input v_2857;
input v_2858;
input v_2859;
input v_2860;
input v_2861;
input v_2862;
input v_2863;
input v_2864;
input v_2865;
input v_2866;
input v_2867;
input v_2868;
input v_2869;
input v_2870;
input v_2871;
input v_2872;
input v_2873;
input v_2874;
input v_2875;
input v_2876;
input v_2877;
input v_2878;
input v_2879;
input v_2880;
input v_2881;
input v_2882;
input v_2883;
input v_2884;
input v_2885;
input v_2886;
input v_2887;
input v_2888;
input v_2889;
input v_2890;
input v_2891;
input v_2892;
input v_2893;
input v_2894;
input v_2895;
input v_2896;
input v_2897;
input v_2898;
input v_2899;
input v_2900;
input v_2901;
input v_2902;
input v_2903;
input v_2904;
input v_2905;
input v_2906;
input v_2907;
input v_2908;
input v_2909;
input v_2910;
input v_2911;
input v_2912;
input v_2913;
input v_2914;
input v_2915;
input v_2916;
input v_2917;
input v_2918;
input v_2919;
input v_2920;
input v_2921;
input v_2922;
input v_2923;
input v_2924;
input v_2925;
input v_2926;
input v_2927;
input v_2928;
input v_2929;
input v_2930;
input v_2931;
input v_2932;
input v_2933;
input v_2934;
input v_2935;
input v_2936;
input v_2937;
input v_2938;
input v_2939;
input v_2940;
input v_2941;
input v_2942;
input v_2943;
input v_2944;
input v_2945;
input v_2946;
input v_2947;
input v_2948;
input v_2949;
input v_2950;
input v_2951;
input v_2952;
input v_2953;
input v_2954;
input v_2955;
input v_2956;
input v_2957;
input v_2958;
input v_2959;
input v_2960;
input v_2961;
input v_2962;
input v_2963;
input v_2964;
input v_2965;
input v_2966;
input v_2967;
input v_2968;
input v_2969;
input v_2970;
input v_2971;
input v_2972;
input v_2973;
input v_2974;
input v_2975;
input v_2976;
input v_2977;
input v_2978;
input v_2979;
input v_2980;
input v_2981;
input v_2982;
input v_2983;
input v_2984;
input v_2985;
input v_2986;
input v_2987;
input v_2988;
input v_2989;
input v_2990;
input v_2991;
input v_2992;
input v_2993;
input v_2994;
input v_2995;
input v_2996;
input v_2997;
input v_2998;
input v_2999;
input v_3000;
input v_3001;
input v_3002;
input v_3003;
input v_3004;
input v_3005;
input v_3006;
input v_3007;
input v_3008;
input v_3009;
input v_3010;
input v_3011;
input v_3012;
input v_3013;
input v_3014;
input v_3015;
input v_3016;
input v_3017;
input v_3018;
input v_3019;
input v_3020;
input v_3021;
input v_3022;
input v_3023;
input v_3024;
input v_3025;
input v_3026;
input v_3027;
input v_3028;
input v_3029;
input v_3030;
input v_3031;
input v_3032;
input v_3033;
input v_3034;
input v_3035;
input v_3036;
input v_3037;
input v_3038;
input v_3039;
input v_3040;
input v_3041;
input v_3042;
input v_3043;
input v_3044;
input v_3045;
input v_3046;
input v_3047;
input v_3048;
input v_3049;
input v_3050;
input v_3051;
input v_3052;
input v_3053;
input v_3054;
input v_3055;
input v_3056;
input v_3057;
input v_3058;
input v_3059;
input v_3060;
input v_3061;
input v_3062;
input v_3063;
input v_3064;
input v_3065;
input v_3066;
input v_3067;
input v_3068;
input v_3069;
input v_3070;
input v_3071;
input v_3072;
input v_3073;
input v_3074;
input v_3075;
input v_3076;
input v_3077;
input v_3078;
input v_3079;
input v_3080;
input v_3081;
input v_3082;
input v_3083;
input v_3084;
input v_3085;
input v_3086;
input v_3087;
input v_3088;
input v_3089;
input v_3090;
input v_3091;
input v_3092;
input v_3093;
input v_3094;
input v_3095;
input v_3096;
input v_3097;
input v_3098;
input v_3099;
input v_3100;
input v_3101;
input v_3102;
input v_3103;
input v_3104;
input v_3105;
input v_3106;
input v_3107;
input v_3108;
input v_3109;
input v_3110;
input v_3111;
input v_3112;
input v_3113;
input v_3114;
input v_3115;
input v_3116;
input v_3117;
input v_3118;
input v_3119;
input v_3120;
input v_3121;
input v_3122;
input v_3123;
input v_3124;
input v_3125;
input v_3126;
input v_3127;
input v_3128;
input v_3129;
input v_3130;
input v_3131;
input v_3132;
input v_3133;
input v_3134;
input v_3135;
input v_3136;
input v_3137;
input v_3138;
input v_3139;
input v_3140;
input v_3141;
input v_3142;
input v_3143;
input v_3144;
input v_3145;
input v_3146;
input v_3147;
input v_3148;
input v_3149;
input v_3150;
input v_3151;
input v_3152;
input v_3153;
input v_3154;
input v_3155;
input v_3156;
input v_3157;
input v_3158;
input v_3159;
input v_3160;
input v_3161;
input v_3162;
input v_3163;
input v_3164;
input v_3165;
input v_3166;
input v_3167;
input v_3168;
input v_3169;
input v_3170;
input v_3171;
input v_3172;
input v_3173;
input v_3174;
input v_3175;
input v_3176;
input v_3177;
input v_3178;
input v_3179;
input v_3180;
input v_3181;
input v_3182;
input v_3183;
input v_3184;
input v_3185;
input v_3186;
input v_3187;
input v_3188;
input v_3189;
input v_3190;
input v_3191;
input v_3192;
input v_3193;
input v_3194;
input v_3195;
input v_3196;
input v_3197;
input v_3198;
input v_3199;
input v_3200;
input v_3201;
input v_3202;
input v_3203;
input v_3204;
input v_3205;
input v_3206;
input v_3207;
input v_3208;
input v_3209;
input v_3210;
input v_3211;
input v_3212;
input v_3213;
input v_3214;
input v_3215;
input v_3216;
input v_3217;
input v_3218;
input v_3219;
input v_3220;
input v_3221;
input v_3222;
input v_3223;
input v_3224;
input v_3225;
input v_3226;
input v_3227;
input v_3228;
input v_3229;
input v_3230;
input v_3231;
input v_3232;
input v_3233;
input v_3234;
input v_3235;
input v_3236;
input v_3237;
input v_3238;
input v_3239;
input v_3240;
input v_3241;
input v_3242;
input v_3243;
input v_3244;
input v_3245;
input v_3246;
input v_3247;
input v_3248;
input v_3249;
input v_3250;
input v_3251;
input v_3252;
input v_3253;
input v_3254;
input v_3255;
input v_3256;
input v_3257;
input v_3258;
input v_3259;
input v_3260;
input v_3261;
input v_3262;
input v_3263;
input v_3264;
input v_3265;
input v_3266;
input v_3267;
input v_3268;
input v_3269;
input v_3270;
input v_3271;
input v_3272;
input v_3273;
input v_3274;
input v_3275;
input v_3276;
input v_3277;
input v_3278;
input v_3279;
input v_3280;
input v_3281;
input v_3282;
input v_3283;
input v_3284;
input v_3285;
input v_3286;
input v_3287;
input v_3288;
input v_3289;
input v_3290;
input v_3291;
input v_3292;
input v_3293;
input v_3294;
input v_3295;
input v_3296;
input v_3297;
input v_3298;
input v_3299;
input v_3300;
input v_3301;
input v_3302;
input v_3303;
input v_3304;
input v_3305;
input v_3306;
input v_3307;
input v_3308;
input v_3309;
input v_3310;
input v_3311;
input v_3312;
input v_3313;
input v_3314;
input v_3315;
input v_3316;
input v_3317;
input v_3318;
input v_3319;
input v_3320;
input v_3321;
input v_3322;
input v_3323;
input v_3324;
input v_3325;
input v_3326;
input v_3327;
input v_3328;
input v_3329;
input v_3330;
input v_3331;
input v_3332;
input v_3333;
input v_3334;
input v_3335;
input v_3336;
input v_3337;
input v_3338;
input v_3339;
input v_3340;
input v_3341;
input v_3342;
input v_3343;
input v_3344;
input v_3345;
input v_3346;
input v_3347;
input v_3348;
input v_3349;
input v_3350;
input v_3351;
input v_3352;
input v_3353;
input v_3354;
input v_3355;
input v_3356;
input v_3357;
input v_3358;
input v_3359;
input v_3360;
input v_3361;
input v_3362;
input v_3363;
input v_3364;
input v_3365;
input v_3366;
input v_3367;
input v_3368;
input v_3369;
input v_3370;
input v_3371;
input v_3372;
input v_3373;
input v_3374;
input v_3375;
input v_3376;
input v_3377;
input v_3378;
input v_3379;
input v_3380;
output o_1;
wire v_3381;
wire x_1;
wire x_2;
wire x_3;
wire x_4;
wire x_5;
wire x_6;
wire x_7;
wire x_8;
wire x_9;
wire x_10;
wire x_11;
wire x_12;
wire x_13;
wire x_14;
wire x_15;
wire x_16;
wire x_17;
wire x_18;
wire x_19;
wire x_20;
wire x_21;
wire x_22;
wire x_23;
wire x_24;
wire x_25;
wire x_26;
wire x_27;
wire x_28;
wire x_29;
wire x_30;
wire x_31;
wire x_32;
wire x_33;
wire x_34;
wire x_35;
wire x_36;
wire x_37;
wire x_38;
wire x_39;
wire x_40;
wire x_41;
wire x_42;
wire x_43;
wire x_44;
wire x_45;
wire x_46;
wire x_47;
wire x_48;
wire x_49;
wire x_50;
wire x_51;
wire x_52;
wire x_53;
wire x_54;
wire x_55;
wire x_56;
wire x_57;
wire x_58;
wire x_59;
wire x_60;
wire x_61;
wire x_62;
wire x_63;
wire x_64;
wire x_65;
wire x_66;
wire x_67;
wire x_68;
wire x_69;
wire x_70;
wire x_71;
wire x_72;
wire x_73;
wire x_74;
wire x_75;
wire x_76;
wire x_77;
wire x_78;
wire x_79;
wire x_80;
wire x_81;
wire x_82;
wire x_83;
wire x_84;
wire x_85;
wire x_86;
wire x_87;
wire x_88;
wire x_89;
wire x_90;
wire x_91;
wire x_92;
wire x_93;
wire x_94;
wire x_95;
wire x_96;
wire x_97;
wire x_98;
wire x_99;
wire x_100;
wire x_101;
wire x_102;
wire x_103;
wire x_104;
wire x_105;
wire x_106;
wire x_107;
wire x_108;
wire x_109;
wire x_110;
wire x_111;
wire x_112;
wire x_113;
wire x_114;
wire x_115;
wire x_116;
wire x_117;
wire x_118;
wire x_119;
wire x_120;
wire x_121;
wire x_122;
wire x_123;
wire x_124;
wire x_125;
wire x_126;
wire x_127;
wire x_128;
wire x_129;
wire x_130;
wire x_131;
wire x_132;
wire x_133;
wire x_134;
wire x_135;
wire x_136;
wire x_137;
wire x_138;
wire x_139;
wire x_140;
wire x_141;
wire x_142;
wire x_143;
wire x_144;
wire x_145;
wire x_146;
wire x_147;
wire x_148;
wire x_149;
wire x_150;
wire x_151;
wire x_152;
wire x_153;
wire x_154;
wire x_155;
wire x_156;
wire x_157;
wire x_158;
wire x_159;
wire x_160;
wire x_161;
wire x_162;
wire x_163;
wire x_164;
wire x_165;
wire x_166;
wire x_167;
wire x_168;
wire x_169;
wire x_170;
wire x_171;
wire x_172;
wire x_173;
wire x_174;
wire x_175;
wire x_176;
wire x_177;
wire x_178;
wire x_179;
wire x_180;
wire x_181;
wire x_182;
wire x_183;
wire x_184;
wire x_185;
wire x_186;
wire x_187;
wire x_188;
wire x_189;
wire x_190;
wire x_191;
wire x_192;
wire x_193;
wire x_194;
wire x_195;
wire x_196;
wire x_197;
wire x_198;
wire x_199;
wire x_200;
wire x_201;
wire x_202;
wire x_203;
wire x_204;
wire x_205;
wire x_206;
wire x_207;
wire x_208;
wire x_209;
wire x_210;
wire x_211;
wire x_212;
wire x_213;
wire x_214;
wire x_215;
wire x_216;
wire x_217;
wire x_218;
wire x_219;
wire x_220;
wire x_221;
wire x_222;
wire x_223;
wire x_224;
wire x_225;
wire x_226;
wire x_227;
wire x_228;
wire x_229;
wire x_230;
wire x_231;
wire x_232;
wire x_233;
wire x_234;
wire x_235;
wire x_236;
wire x_237;
wire x_238;
wire x_239;
wire x_240;
wire x_241;
wire x_242;
wire x_243;
wire x_244;
wire x_245;
wire x_246;
wire x_247;
wire x_248;
wire x_249;
wire x_250;
wire x_251;
wire x_252;
wire x_253;
wire x_254;
wire x_255;
wire x_256;
wire x_257;
wire x_258;
wire x_259;
wire x_260;
wire x_261;
wire x_262;
wire x_263;
wire x_264;
wire x_265;
wire x_266;
wire x_267;
wire x_268;
wire x_269;
wire x_270;
wire x_271;
wire x_272;
wire x_273;
wire x_274;
wire x_275;
wire x_276;
wire x_277;
wire x_278;
wire x_279;
wire x_280;
wire x_281;
wire x_282;
wire x_283;
wire x_284;
wire x_285;
wire x_286;
wire x_287;
wire x_288;
wire x_289;
wire x_290;
wire x_291;
wire x_292;
wire x_293;
wire x_294;
wire x_295;
wire x_296;
wire x_297;
wire x_298;
wire x_299;
wire x_300;
wire x_301;
wire x_302;
wire x_303;
wire x_304;
wire x_305;
wire x_306;
wire x_307;
wire x_308;
wire x_309;
wire x_310;
wire x_311;
wire x_312;
wire x_313;
wire x_314;
wire x_315;
wire x_316;
wire x_317;
wire x_318;
wire x_319;
wire x_320;
wire x_321;
wire x_322;
wire x_323;
wire x_324;
wire x_325;
wire x_326;
wire x_327;
wire x_328;
wire x_329;
wire x_330;
wire x_331;
wire x_332;
wire x_333;
wire x_334;
wire x_335;
wire x_336;
wire x_337;
wire x_338;
wire x_339;
wire x_340;
wire x_341;
wire x_342;
wire x_343;
wire x_344;
wire x_345;
wire x_346;
wire x_347;
wire x_348;
wire x_349;
wire x_350;
wire x_351;
wire x_352;
wire x_353;
wire x_354;
wire x_355;
wire x_356;
wire x_357;
wire x_358;
wire x_359;
wire x_360;
wire x_361;
wire x_362;
wire x_363;
wire x_364;
wire x_365;
wire x_366;
wire x_367;
wire x_368;
wire x_369;
wire x_370;
wire x_371;
wire x_372;
wire x_373;
wire x_374;
wire x_375;
wire x_376;
wire x_377;
wire x_378;
wire x_379;
wire x_380;
wire x_381;
wire x_382;
wire x_383;
wire x_384;
wire x_385;
wire x_386;
wire x_387;
wire x_388;
wire x_389;
wire x_390;
wire x_391;
wire x_392;
wire x_393;
wire x_394;
wire x_395;
wire x_396;
wire x_397;
wire x_398;
wire x_399;
wire x_400;
wire x_401;
wire x_402;
wire x_403;
wire x_404;
wire x_405;
wire x_406;
wire x_407;
wire x_408;
wire x_409;
wire x_410;
wire x_411;
wire x_412;
wire x_413;
wire x_414;
wire x_415;
wire x_416;
wire x_417;
wire x_418;
wire x_419;
wire x_420;
wire x_421;
wire x_422;
wire x_423;
wire x_424;
wire x_425;
wire x_426;
wire x_427;
wire x_428;
wire x_429;
wire x_430;
wire x_431;
wire x_432;
wire x_433;
wire x_434;
wire x_435;
wire x_436;
wire x_437;
wire x_438;
wire x_439;
wire x_440;
wire x_441;
wire x_442;
wire x_443;
wire x_444;
wire x_445;
wire x_446;
wire x_447;
wire x_448;
wire x_449;
wire x_450;
wire x_451;
wire x_452;
wire x_453;
wire x_454;
wire x_455;
wire x_456;
wire x_457;
wire x_458;
wire x_459;
wire x_460;
wire x_461;
wire x_462;
wire x_463;
wire x_464;
wire x_465;
wire x_466;
wire x_467;
wire x_468;
wire x_469;
wire x_470;
wire x_471;
wire x_472;
wire x_473;
wire x_474;
wire x_475;
wire x_476;
wire x_477;
wire x_478;
wire x_479;
wire x_480;
wire x_481;
wire x_482;
wire x_483;
wire x_484;
wire x_485;
wire x_486;
wire x_487;
wire x_488;
wire x_489;
wire x_490;
wire x_491;
wire x_492;
wire x_493;
wire x_494;
wire x_495;
wire x_496;
wire x_497;
wire x_498;
wire x_499;
wire x_500;
wire x_501;
wire x_502;
wire x_503;
wire x_504;
wire x_505;
wire x_506;
wire x_507;
wire x_508;
wire x_509;
wire x_510;
wire x_511;
wire x_512;
wire x_513;
wire x_514;
wire x_515;
wire x_516;
wire x_517;
wire x_518;
wire x_519;
wire x_520;
wire x_521;
wire x_522;
wire x_523;
wire x_524;
wire x_525;
wire x_526;
wire x_527;
wire x_528;
wire x_529;
wire x_530;
wire x_531;
wire x_532;
wire x_533;
wire x_534;
wire x_535;
wire x_536;
wire x_537;
wire x_538;
wire x_539;
wire x_540;
wire x_541;
wire x_542;
wire x_543;
wire x_544;
wire x_545;
wire x_546;
wire x_547;
wire x_548;
wire x_549;
wire x_550;
wire x_551;
wire x_552;
wire x_553;
wire x_554;
wire x_555;
wire x_556;
wire x_557;
wire x_558;
wire x_559;
wire x_560;
wire x_561;
wire x_562;
wire x_563;
wire x_564;
wire x_565;
wire x_566;
wire x_567;
wire x_568;
wire x_569;
wire x_570;
wire x_571;
wire x_572;
wire x_573;
wire x_574;
wire x_575;
wire x_576;
wire x_577;
wire x_578;
wire x_579;
wire x_580;
wire x_581;
wire x_582;
wire x_583;
wire x_584;
wire x_585;
wire x_586;
wire x_587;
wire x_588;
wire x_589;
wire x_590;
wire x_591;
wire x_592;
wire x_593;
wire x_594;
wire x_595;
wire x_596;
wire x_597;
wire x_598;
wire x_599;
wire x_600;
wire x_601;
wire x_602;
wire x_603;
wire x_604;
wire x_605;
wire x_606;
wire x_607;
wire x_608;
wire x_609;
wire x_610;
wire x_611;
wire x_612;
wire x_613;
wire x_614;
wire x_615;
wire x_616;
wire x_617;
wire x_618;
wire x_619;
wire x_620;
wire x_621;
wire x_622;
wire x_623;
wire x_624;
wire x_625;
wire x_626;
wire x_627;
wire x_628;
wire x_629;
wire x_630;
wire x_631;
wire x_632;
wire x_633;
wire x_634;
wire x_635;
wire x_636;
wire x_637;
wire x_638;
wire x_639;
wire x_640;
wire x_641;
wire x_642;
wire x_643;
wire x_644;
wire x_645;
wire x_646;
wire x_647;
wire x_648;
wire x_649;
wire x_650;
wire x_651;
wire x_652;
wire x_653;
wire x_654;
wire x_655;
wire x_656;
wire x_657;
wire x_658;
wire x_659;
wire x_660;
wire x_661;
wire x_662;
wire x_663;
wire x_664;
wire x_665;
wire x_666;
wire x_667;
wire x_668;
wire x_669;
wire x_670;
wire x_671;
wire x_672;
wire x_673;
wire x_674;
wire x_675;
wire x_676;
wire x_677;
wire x_678;
wire x_679;
wire x_680;
wire x_681;
wire x_682;
wire x_683;
wire x_684;
wire x_685;
wire x_686;
wire x_687;
wire x_688;
wire x_689;
wire x_690;
wire x_691;
wire x_692;
wire x_693;
wire x_694;
wire x_695;
wire x_696;
wire x_697;
wire x_698;
wire x_699;
wire x_700;
wire x_701;
wire x_702;
wire x_703;
wire x_704;
wire x_705;
wire x_706;
wire x_707;
wire x_708;
wire x_709;
wire x_710;
wire x_711;
wire x_712;
wire x_713;
wire x_714;
wire x_715;
wire x_716;
wire x_717;
wire x_718;
wire x_719;
wire x_720;
wire x_721;
wire x_722;
wire x_723;
wire x_724;
wire x_725;
wire x_726;
wire x_727;
wire x_728;
wire x_729;
wire x_730;
wire x_731;
wire x_732;
wire x_733;
wire x_734;
wire x_735;
wire x_736;
wire x_737;
wire x_738;
wire x_739;
wire x_740;
wire x_741;
wire x_742;
wire x_743;
wire x_744;
wire x_745;
wire x_746;
wire x_747;
wire x_748;
wire x_749;
wire x_750;
wire x_751;
wire x_752;
wire x_753;
wire x_754;
wire x_755;
wire x_756;
wire x_757;
wire x_758;
wire x_759;
wire x_760;
wire x_761;
wire x_762;
wire x_763;
wire x_764;
wire x_765;
wire x_766;
wire x_767;
wire x_768;
wire x_769;
wire x_770;
wire x_771;
wire x_772;
wire x_773;
wire x_774;
wire x_775;
wire x_776;
wire x_777;
wire x_778;
wire x_779;
wire x_780;
wire x_781;
wire x_782;
wire x_783;
wire x_784;
wire x_785;
wire x_786;
wire x_787;
wire x_788;
wire x_789;
wire x_790;
wire x_791;
wire x_792;
wire x_793;
wire x_794;
wire x_795;
wire x_796;
wire x_797;
wire x_798;
wire x_799;
wire x_800;
wire x_801;
wire x_802;
wire x_803;
wire x_804;
wire x_805;
wire x_806;
wire x_807;
wire x_808;
wire x_809;
wire x_810;
wire x_811;
wire x_812;
wire x_813;
wire x_814;
wire x_815;
wire x_816;
wire x_817;
wire x_818;
wire x_819;
wire x_820;
wire x_821;
wire x_822;
wire x_823;
wire x_824;
wire x_825;
wire x_826;
wire x_827;
wire x_828;
wire x_829;
wire x_830;
wire x_831;
wire x_832;
wire x_833;
wire x_834;
wire x_835;
wire x_836;
wire x_837;
wire x_838;
wire x_839;
wire x_840;
wire x_841;
wire x_842;
wire x_843;
wire x_844;
wire x_845;
wire x_846;
wire x_847;
wire x_848;
wire x_849;
wire x_850;
wire x_851;
wire x_852;
wire x_853;
wire x_854;
wire x_855;
wire x_856;
wire x_857;
wire x_858;
wire x_859;
wire x_860;
wire x_861;
wire x_862;
wire x_863;
wire x_864;
wire x_865;
wire x_866;
wire x_867;
wire x_868;
wire x_869;
wire x_870;
wire x_871;
wire x_872;
wire x_873;
wire x_874;
wire x_875;
wire x_876;
wire x_877;
wire x_878;
wire x_879;
wire x_880;
wire x_881;
wire x_882;
wire x_883;
wire x_884;
wire x_885;
wire x_886;
wire x_887;
wire x_888;
wire x_889;
wire x_890;
wire x_891;
wire x_892;
wire x_893;
wire x_894;
wire x_895;
wire x_896;
wire x_897;
wire x_898;
wire x_899;
wire x_900;
wire x_901;
wire x_902;
wire x_903;
wire x_904;
wire x_905;
wire x_906;
wire x_907;
wire x_908;
wire x_909;
wire x_910;
wire x_911;
wire x_912;
wire x_913;
wire x_914;
wire x_915;
wire x_916;
wire x_917;
wire x_918;
wire x_919;
wire x_920;
wire x_921;
wire x_922;
wire x_923;
wire x_924;
wire x_925;
wire x_926;
wire x_927;
wire x_928;
wire x_929;
wire x_930;
wire x_931;
wire x_932;
wire x_933;
wire x_934;
wire x_935;
wire x_936;
wire x_937;
wire x_938;
wire x_939;
wire x_940;
wire x_941;
wire x_942;
wire x_943;
wire x_944;
wire x_945;
wire x_946;
wire x_947;
wire x_948;
wire x_949;
wire x_950;
wire x_951;
wire x_952;
wire x_953;
wire x_954;
wire x_955;
wire x_956;
wire x_957;
wire x_958;
wire x_959;
wire x_960;
wire x_961;
wire x_962;
wire x_963;
wire x_964;
wire x_965;
wire x_966;
wire x_967;
wire x_968;
wire x_969;
wire x_970;
wire x_971;
wire x_972;
wire x_973;
wire x_974;
wire x_975;
wire x_976;
wire x_977;
wire x_978;
wire x_979;
wire x_980;
wire x_981;
wire x_982;
wire x_983;
wire x_984;
wire x_985;
wire x_986;
wire x_987;
wire x_988;
wire x_989;
wire x_990;
wire x_991;
wire x_992;
wire x_993;
wire x_994;
wire x_995;
wire x_996;
wire x_997;
wire x_998;
wire x_999;
wire x_1000;
wire x_1001;
wire x_1002;
wire x_1003;
wire x_1004;
wire x_1005;
wire x_1006;
wire x_1007;
wire x_1008;
wire x_1009;
wire x_1010;
wire x_1011;
wire x_1012;
wire x_1013;
wire x_1014;
wire x_1015;
wire x_1016;
wire x_1017;
wire x_1018;
wire x_1019;
wire x_1020;
wire x_1021;
wire x_1022;
wire x_1023;
wire x_1024;
wire x_1025;
wire x_1026;
wire x_1027;
wire x_1028;
wire x_1029;
wire x_1030;
wire x_1031;
wire x_1032;
wire x_1033;
wire x_1034;
wire x_1035;
wire x_1036;
wire x_1037;
wire x_1038;
wire x_1039;
wire x_1040;
wire x_1041;
wire x_1042;
wire x_1043;
wire x_1044;
wire x_1045;
wire x_1046;
wire x_1047;
wire x_1048;
wire x_1049;
wire x_1050;
wire x_1051;
wire x_1052;
wire x_1053;
wire x_1054;
wire x_1055;
wire x_1056;
wire x_1057;
wire x_1058;
wire x_1059;
wire x_1060;
wire x_1061;
wire x_1062;
wire x_1063;
wire x_1064;
wire x_1065;
wire x_1066;
wire x_1067;
wire x_1068;
wire x_1069;
wire x_1070;
wire x_1071;
wire x_1072;
wire x_1073;
wire x_1074;
wire x_1075;
wire x_1076;
wire x_1077;
wire x_1078;
wire x_1079;
wire x_1080;
wire x_1081;
wire x_1082;
wire x_1083;
wire x_1084;
wire x_1085;
wire x_1086;
wire x_1087;
wire x_1088;
wire x_1089;
wire x_1090;
wire x_1091;
wire x_1092;
wire x_1093;
wire x_1094;
wire x_1095;
wire x_1096;
wire x_1097;
wire x_1098;
wire x_1099;
wire x_1100;
wire x_1101;
wire x_1102;
wire x_1103;
wire x_1104;
wire x_1105;
wire x_1106;
wire x_1107;
wire x_1108;
wire x_1109;
wire x_1110;
wire x_1111;
wire x_1112;
wire x_1113;
wire x_1114;
wire x_1115;
wire x_1116;
wire x_1117;
wire x_1118;
wire x_1119;
wire x_1120;
wire x_1121;
wire x_1122;
wire x_1123;
wire x_1124;
wire x_1125;
wire x_1126;
wire x_1127;
wire x_1128;
wire x_1129;
wire x_1130;
wire x_1131;
wire x_1132;
wire x_1133;
wire x_1134;
wire x_1135;
wire x_1136;
wire x_1137;
wire x_1138;
wire x_1139;
wire x_1140;
wire x_1141;
wire x_1142;
wire x_1143;
wire x_1144;
wire x_1145;
wire x_1146;
wire x_1147;
wire x_1148;
wire x_1149;
wire x_1150;
wire x_1151;
wire x_1152;
wire x_1153;
wire x_1154;
wire x_1155;
wire x_1156;
wire x_1157;
wire x_1158;
wire x_1159;
wire x_1160;
wire x_1161;
wire x_1162;
wire x_1163;
wire x_1164;
wire x_1165;
wire x_1166;
wire x_1167;
wire x_1168;
wire x_1169;
wire x_1170;
wire x_1171;
wire x_1172;
wire x_1173;
wire x_1174;
wire x_1175;
wire x_1176;
wire x_1177;
wire x_1178;
wire x_1179;
wire x_1180;
wire x_1181;
wire x_1182;
wire x_1183;
wire x_1184;
wire x_1185;
wire x_1186;
wire x_1187;
wire x_1188;
wire x_1189;
wire x_1190;
wire x_1191;
wire x_1192;
wire x_1193;
wire x_1194;
wire x_1195;
wire x_1196;
wire x_1197;
wire x_1198;
wire x_1199;
wire x_1200;
wire x_1201;
wire x_1202;
wire x_1203;
wire x_1204;
wire x_1205;
wire x_1206;
wire x_1207;
wire x_1208;
wire x_1209;
wire x_1210;
wire x_1211;
wire x_1212;
wire x_1213;
wire x_1214;
wire x_1215;
wire x_1216;
wire x_1217;
wire x_1218;
wire x_1219;
wire x_1220;
wire x_1221;
wire x_1222;
wire x_1223;
wire x_1224;
wire x_1225;
wire x_1226;
wire x_1227;
wire x_1228;
wire x_1229;
wire x_1230;
wire x_1231;
wire x_1232;
wire x_1233;
wire x_1234;
wire x_1235;
wire x_1236;
wire x_1237;
wire x_1238;
wire x_1239;
wire x_1240;
wire x_1241;
wire x_1242;
wire x_1243;
wire x_1244;
wire x_1245;
wire x_1246;
wire x_1247;
wire x_1248;
wire x_1249;
wire x_1250;
wire x_1251;
wire x_1252;
wire x_1253;
wire x_1254;
wire x_1255;
wire x_1256;
wire x_1257;
wire x_1258;
wire x_1259;
wire x_1260;
wire x_1261;
wire x_1262;
wire x_1263;
wire x_1264;
wire x_1265;
wire x_1266;
wire x_1267;
wire x_1268;
wire x_1269;
wire x_1270;
wire x_1271;
wire x_1272;
wire x_1273;
wire x_1274;
wire x_1275;
wire x_1276;
wire x_1277;
wire x_1278;
wire x_1279;
wire x_1280;
wire x_1281;
wire x_1282;
wire x_1283;
wire x_1284;
wire x_1285;
wire x_1286;
wire x_1287;
wire x_1288;
wire x_1289;
wire x_1290;
wire x_1291;
wire x_1292;
wire x_1293;
wire x_1294;
wire x_1295;
wire x_1296;
wire x_1297;
wire x_1298;
wire x_1299;
wire x_1300;
wire x_1301;
wire x_1302;
wire x_1303;
wire x_1304;
wire x_1305;
wire x_1306;
wire x_1307;
wire x_1308;
wire x_1309;
wire x_1310;
wire x_1311;
wire x_1312;
wire x_1313;
wire x_1314;
wire x_1315;
wire x_1316;
wire x_1317;
wire x_1318;
wire x_1319;
wire x_1320;
wire x_1321;
wire x_1322;
wire x_1323;
wire x_1324;
wire x_1325;
wire x_1326;
wire x_1327;
wire x_1328;
wire x_1329;
wire x_1330;
wire x_1331;
wire x_1332;
wire x_1333;
wire x_1334;
wire x_1335;
wire x_1336;
wire x_1337;
wire x_1338;
wire x_1339;
wire x_1340;
wire x_1341;
wire x_1342;
wire x_1343;
wire x_1344;
wire x_1345;
wire x_1346;
wire x_1347;
wire x_1348;
wire x_1349;
wire x_1350;
wire x_1351;
wire x_1352;
wire x_1353;
wire x_1354;
wire x_1355;
wire x_1356;
wire x_1357;
wire x_1358;
wire x_1359;
wire x_1360;
wire x_1361;
wire x_1362;
wire x_1363;
wire x_1364;
wire x_1365;
wire x_1366;
wire x_1367;
wire x_1368;
wire x_1369;
wire x_1370;
wire x_1371;
wire x_1372;
wire x_1373;
wire x_1374;
wire x_1375;
wire x_1376;
wire x_1377;
wire x_1378;
wire x_1379;
wire x_1380;
wire x_1381;
wire x_1382;
wire x_1383;
wire x_1384;
wire x_1385;
wire x_1386;
wire x_1387;
wire x_1388;
wire x_1389;
wire x_1390;
wire x_1391;
wire x_1392;
wire x_1393;
wire x_1394;
wire x_1395;
wire x_1396;
wire x_1397;
wire x_1398;
wire x_1399;
wire x_1400;
wire x_1401;
wire x_1402;
wire x_1403;
wire x_1404;
wire x_1405;
wire x_1406;
wire x_1407;
wire x_1408;
wire x_1409;
wire x_1410;
wire x_1411;
wire x_1412;
wire x_1413;
wire x_1414;
wire x_1415;
wire x_1416;
wire x_1417;
wire x_1418;
wire x_1419;
wire x_1420;
wire x_1421;
wire x_1422;
wire x_1423;
wire x_1424;
wire x_1425;
wire x_1426;
wire x_1427;
wire x_1428;
wire x_1429;
wire x_1430;
wire x_1431;
wire x_1432;
wire x_1433;
wire x_1434;
wire x_1435;
wire x_1436;
wire x_1437;
wire x_1438;
wire x_1439;
wire x_1440;
wire x_1441;
wire x_1442;
wire x_1443;
wire x_1444;
wire x_1445;
wire x_1446;
wire x_1447;
wire x_1448;
wire x_1449;
wire x_1450;
wire x_1451;
wire x_1452;
wire x_1453;
wire x_1454;
wire x_1455;
wire x_1456;
wire x_1457;
wire x_1458;
wire x_1459;
wire x_1460;
wire x_1461;
wire x_1462;
wire x_1463;
wire x_1464;
wire x_1465;
wire x_1466;
wire x_1467;
wire x_1468;
wire x_1469;
wire x_1470;
wire x_1471;
wire x_1472;
wire x_1473;
wire x_1474;
wire x_1475;
wire x_1476;
wire x_1477;
wire x_1478;
wire x_1479;
wire x_1480;
wire x_1481;
wire x_1482;
wire x_1483;
wire x_1484;
wire x_1485;
wire x_1486;
wire x_1487;
wire x_1488;
wire x_1489;
wire x_1490;
wire x_1491;
wire x_1492;
wire x_1493;
wire x_1494;
wire x_1495;
wire x_1496;
wire x_1497;
wire x_1498;
wire x_1499;
wire x_1500;
wire x_1501;
wire x_1502;
wire x_1503;
wire x_1504;
wire x_1505;
wire x_1506;
wire x_1507;
wire x_1508;
wire x_1509;
wire x_1510;
wire x_1511;
wire x_1512;
wire x_1513;
wire x_1514;
wire x_1515;
wire x_1516;
wire x_1517;
wire x_1518;
wire x_1519;
wire x_1520;
wire x_1521;
wire x_1522;
wire x_1523;
wire x_1524;
wire x_1525;
wire x_1526;
wire x_1527;
wire x_1528;
wire x_1529;
wire x_1530;
wire x_1531;
wire x_1532;
wire x_1533;
wire x_1534;
wire x_1535;
wire x_1536;
wire x_1537;
wire x_1538;
wire x_1539;
wire x_1540;
wire x_1541;
wire x_1542;
wire x_1543;
wire x_1544;
wire x_1545;
wire x_1546;
wire x_1547;
wire x_1548;
wire x_1549;
wire x_1550;
wire x_1551;
wire x_1552;
wire x_1553;
wire x_1554;
wire x_1555;
wire x_1556;
wire x_1557;
wire x_1558;
wire x_1559;
wire x_1560;
wire x_1561;
wire x_1562;
wire x_1563;
wire x_1564;
wire x_1565;
wire x_1566;
wire x_1567;
wire x_1568;
wire x_1569;
wire x_1570;
wire x_1571;
wire x_1572;
wire x_1573;
wire x_1574;
wire x_1575;
wire x_1576;
wire x_1577;
wire x_1578;
wire x_1579;
wire x_1580;
wire x_1581;
wire x_1582;
wire x_1583;
wire x_1584;
wire x_1585;
wire x_1586;
wire x_1587;
wire x_1588;
wire x_1589;
wire x_1590;
wire x_1591;
wire x_1592;
wire x_1593;
wire x_1594;
wire x_1595;
wire x_1596;
wire x_1597;
wire x_1598;
wire x_1599;
wire x_1600;
wire x_1601;
wire x_1602;
wire x_1603;
wire x_1604;
wire x_1605;
wire x_1606;
wire x_1607;
wire x_1608;
wire x_1609;
wire x_1610;
wire x_1611;
wire x_1612;
wire x_1613;
wire x_1614;
wire x_1615;
wire x_1616;
wire x_1617;
wire x_1618;
wire x_1619;
wire x_1620;
wire x_1621;
wire x_1622;
wire x_1623;
wire x_1624;
wire x_1625;
wire x_1626;
wire x_1627;
wire x_1628;
wire x_1629;
wire x_1630;
wire x_1631;
wire x_1632;
wire x_1633;
wire x_1634;
wire x_1635;
wire x_1636;
wire x_1637;
wire x_1638;
wire x_1639;
wire x_1640;
wire x_1641;
wire x_1642;
wire x_1643;
wire x_1644;
wire x_1645;
wire x_1646;
wire x_1647;
wire x_1648;
wire x_1649;
wire x_1650;
wire x_1651;
wire x_1652;
wire x_1653;
wire x_1654;
wire x_1655;
wire x_1656;
wire x_1657;
wire x_1658;
wire x_1659;
wire x_1660;
wire x_1661;
wire x_1662;
wire x_1663;
wire x_1664;
wire x_1665;
wire x_1666;
wire x_1667;
wire x_1668;
wire x_1669;
wire x_1670;
wire x_1671;
wire x_1672;
wire x_1673;
wire x_1674;
wire x_1675;
wire x_1676;
wire x_1677;
wire x_1678;
wire x_1679;
wire x_1680;
wire x_1681;
wire x_1682;
wire x_1683;
wire x_1684;
wire x_1685;
wire x_1686;
wire x_1687;
wire x_1688;
wire x_1689;
wire x_1690;
wire x_1691;
wire x_1692;
wire x_1693;
wire x_1694;
wire x_1695;
wire x_1696;
wire x_1697;
wire x_1698;
wire x_1699;
wire x_1700;
wire x_1701;
wire x_1702;
wire x_1703;
wire x_1704;
wire x_1705;
wire x_1706;
wire x_1707;
wire x_1708;
wire x_1709;
wire x_1710;
wire x_1711;
wire x_1712;
wire x_1713;
wire x_1714;
wire x_1715;
wire x_1716;
wire x_1717;
wire x_1718;
wire x_1719;
wire x_1720;
wire x_1721;
wire x_1722;
wire x_1723;
wire x_1724;
wire x_1725;
wire x_1726;
wire x_1727;
wire x_1728;
wire x_1729;
wire x_1730;
wire x_1731;
wire x_1732;
wire x_1733;
wire x_1734;
wire x_1735;
wire x_1736;
wire x_1737;
wire x_1738;
wire x_1739;
wire x_1740;
wire x_1741;
wire x_1742;
wire x_1743;
wire x_1744;
wire x_1745;
wire x_1746;
wire x_1747;
wire x_1748;
wire x_1749;
wire x_1750;
wire x_1751;
wire x_1752;
wire x_1753;
wire x_1754;
wire x_1755;
wire x_1756;
wire x_1757;
wire x_1758;
wire x_1759;
wire x_1760;
wire x_1761;
wire x_1762;
wire x_1763;
wire x_1764;
wire x_1765;
wire x_1766;
wire x_1767;
wire x_1768;
wire x_1769;
wire x_1770;
wire x_1771;
wire x_1772;
wire x_1773;
wire x_1774;
wire x_1775;
wire x_1776;
wire x_1777;
wire x_1778;
wire x_1779;
wire x_1780;
wire x_1781;
wire x_1782;
wire x_1783;
wire x_1784;
wire x_1785;
wire x_1786;
wire x_1787;
wire x_1788;
wire x_1789;
wire x_1790;
wire x_1791;
wire x_1792;
wire x_1793;
wire x_1794;
wire x_1795;
wire x_1796;
wire x_1797;
wire x_1798;
wire x_1799;
wire x_1800;
wire x_1801;
wire x_1802;
wire x_1803;
wire x_1804;
wire x_1805;
wire x_1806;
wire x_1807;
wire x_1808;
wire x_1809;
wire x_1810;
wire x_1811;
wire x_1812;
wire x_1813;
wire x_1814;
wire x_1815;
wire x_1816;
wire x_1817;
wire x_1818;
wire x_1819;
wire x_1820;
wire x_1821;
wire x_1822;
wire x_1823;
wire x_1824;
wire x_1825;
wire x_1826;
wire x_1827;
wire x_1828;
wire x_1829;
wire x_1830;
wire x_1831;
wire x_1832;
wire x_1833;
wire x_1834;
wire x_1835;
wire x_1836;
wire x_1837;
wire x_1838;
wire x_1839;
wire x_1840;
wire x_1841;
wire x_1842;
wire x_1843;
wire x_1844;
wire x_1845;
wire x_1846;
wire x_1847;
wire x_1848;
wire x_1849;
wire x_1850;
wire x_1851;
wire x_1852;
wire x_1853;
wire x_1854;
wire x_1855;
wire x_1856;
wire x_1857;
wire x_1858;
wire x_1859;
wire x_1860;
wire x_1861;
wire x_1862;
wire x_1863;
wire x_1864;
wire x_1865;
wire x_1866;
wire x_1867;
wire x_1868;
wire x_1869;
wire x_1870;
wire x_1871;
wire x_1872;
wire x_1873;
wire x_1874;
wire x_1875;
wire x_1876;
wire x_1877;
wire x_1878;
wire x_1879;
wire x_1880;
wire x_1881;
wire x_1882;
wire x_1883;
wire x_1884;
wire x_1885;
wire x_1886;
wire x_1887;
wire x_1888;
wire x_1889;
wire x_1890;
wire x_1891;
wire x_1892;
wire x_1893;
wire x_1894;
wire x_1895;
wire x_1896;
wire x_1897;
wire x_1898;
wire x_1899;
wire x_1900;
wire x_1901;
wire x_1902;
wire x_1903;
wire x_1904;
wire x_1905;
wire x_1906;
wire x_1907;
wire x_1908;
wire x_1909;
wire x_1910;
wire x_1911;
wire x_1912;
wire x_1913;
wire x_1914;
wire x_1915;
wire x_1916;
wire x_1917;
wire x_1918;
wire x_1919;
wire x_1920;
wire x_1921;
wire x_1922;
wire x_1923;
wire x_1924;
wire x_1925;
wire x_1926;
wire x_1927;
wire x_1928;
wire x_1929;
wire x_1930;
wire x_1931;
wire x_1932;
wire x_1933;
wire x_1934;
wire x_1935;
wire x_1936;
wire x_1937;
wire x_1938;
wire x_1939;
wire x_1940;
wire x_1941;
wire x_1942;
wire x_1943;
wire x_1944;
wire x_1945;
wire x_1946;
wire x_1947;
wire x_1948;
wire x_1949;
wire x_1950;
wire x_1951;
wire x_1952;
wire x_1953;
wire x_1954;
wire x_1955;
wire x_1956;
wire x_1957;
wire x_1958;
wire x_1959;
wire x_1960;
wire x_1961;
wire x_1962;
wire x_1963;
wire x_1964;
wire x_1965;
wire x_1966;
wire x_1967;
wire x_1968;
wire x_1969;
wire x_1970;
wire x_1971;
wire x_1972;
wire x_1973;
wire x_1974;
wire x_1975;
wire x_1976;
wire x_1977;
wire x_1978;
wire x_1979;
wire x_1980;
wire x_1981;
wire x_1982;
wire x_1983;
wire x_1984;
wire x_1985;
wire x_1986;
wire x_1987;
wire x_1988;
wire x_1989;
wire x_1990;
wire x_1991;
wire x_1992;
wire x_1993;
wire x_1994;
wire x_1995;
wire x_1996;
wire x_1997;
wire x_1998;
wire x_1999;
wire x_2000;
wire x_2001;
wire x_2002;
wire x_2003;
wire x_2004;
wire x_2005;
wire x_2006;
wire x_2007;
wire x_2008;
wire x_2009;
wire x_2010;
wire x_2011;
wire x_2012;
wire x_2013;
wire x_2014;
wire x_2015;
wire x_2016;
wire x_2017;
wire x_2018;
wire x_2019;
wire x_2020;
wire x_2021;
wire x_2022;
wire x_2023;
wire x_2024;
wire x_2025;
wire x_2026;
wire x_2027;
wire x_2028;
wire x_2029;
wire x_2030;
wire x_2031;
wire x_2032;
wire x_2033;
wire x_2034;
wire x_2035;
wire x_2036;
wire x_2037;
wire x_2038;
wire x_2039;
wire x_2040;
wire x_2041;
wire x_2042;
wire x_2043;
wire x_2044;
wire x_2045;
wire x_2046;
wire x_2047;
wire x_2048;
wire x_2049;
wire x_2050;
wire x_2051;
wire x_2052;
wire x_2053;
wire x_2054;
wire x_2055;
wire x_2056;
wire x_2057;
wire x_2058;
wire x_2059;
wire x_2060;
wire x_2061;
wire x_2062;
wire x_2063;
wire x_2064;
wire x_2065;
wire x_2066;
wire x_2067;
wire x_2068;
wire x_2069;
wire x_2070;
wire x_2071;
wire x_2072;
wire x_2073;
wire x_2074;
wire x_2075;
wire x_2076;
wire x_2077;
wire x_2078;
wire x_2079;
wire x_2080;
wire x_2081;
wire x_2082;
wire x_2083;
wire x_2084;
wire x_2085;
wire x_2086;
wire x_2087;
wire x_2088;
wire x_2089;
wire x_2090;
wire x_2091;
wire x_2092;
wire x_2093;
wire x_2094;
wire x_2095;
wire x_2096;
wire x_2097;
wire x_2098;
wire x_2099;
wire x_2100;
wire x_2101;
wire x_2102;
wire x_2103;
wire x_2104;
wire x_2105;
wire x_2106;
wire x_2107;
wire x_2108;
wire x_2109;
wire x_2110;
wire x_2111;
wire x_2112;
wire x_2113;
wire x_2114;
wire x_2115;
wire x_2116;
wire x_2117;
wire x_2118;
wire x_2119;
wire x_2120;
wire x_2121;
wire x_2122;
wire x_2123;
wire x_2124;
wire x_2125;
wire x_2126;
wire x_2127;
wire x_2128;
wire x_2129;
wire x_2130;
wire x_2131;
wire x_2132;
wire x_2133;
wire x_2134;
wire x_2135;
wire x_2136;
wire x_2137;
wire x_2138;
wire x_2139;
wire x_2140;
wire x_2141;
wire x_2142;
wire x_2143;
wire x_2144;
wire x_2145;
wire x_2146;
wire x_2147;
wire x_2148;
wire x_2149;
wire x_2150;
wire x_2151;
wire x_2152;
wire x_2153;
wire x_2154;
wire x_2155;
wire x_2156;
wire x_2157;
wire x_2158;
wire x_2159;
wire x_2160;
wire x_2161;
wire x_2162;
wire x_2163;
wire x_2164;
wire x_2165;
wire x_2166;
wire x_2167;
wire x_2168;
wire x_2169;
wire x_2170;
wire x_2171;
wire x_2172;
wire x_2173;
wire x_2174;
wire x_2175;
wire x_2176;
wire x_2177;
wire x_2178;
wire x_2179;
wire x_2180;
wire x_2181;
wire x_2182;
wire x_2183;
wire x_2184;
wire x_2185;
wire x_2186;
wire x_2187;
wire x_2188;
wire x_2189;
wire x_2190;
wire x_2191;
wire x_2192;
wire x_2193;
wire x_2194;
wire x_2195;
wire x_2196;
wire x_2197;
wire x_2198;
wire x_2199;
wire x_2200;
wire x_2201;
wire x_2202;
wire x_2203;
wire x_2204;
wire x_2205;
wire x_2206;
wire x_2207;
wire x_2208;
wire x_2209;
wire x_2210;
wire x_2211;
wire x_2212;
wire x_2213;
wire x_2214;
wire x_2215;
wire x_2216;
wire x_2217;
wire x_2218;
wire x_2219;
wire x_2220;
wire x_2221;
wire x_2222;
wire x_2223;
wire x_2224;
wire x_2225;
wire x_2226;
wire x_2227;
wire x_2228;
wire x_2229;
wire x_2230;
wire x_2231;
wire x_2232;
wire x_2233;
wire x_2234;
wire x_2235;
wire x_2236;
wire x_2237;
wire x_2238;
wire x_2239;
wire x_2240;
wire x_2241;
wire x_2242;
wire x_2243;
wire x_2244;
wire x_2245;
wire x_2246;
wire x_2247;
wire x_2248;
wire x_2249;
wire x_2250;
wire x_2251;
wire x_2252;
wire x_2253;
wire x_2254;
wire x_2255;
wire x_2256;
wire x_2257;
wire x_2258;
wire x_2259;
wire x_2260;
wire x_2261;
wire x_2262;
wire x_2263;
wire x_2264;
wire x_2265;
wire x_2266;
wire x_2267;
wire x_2268;
wire x_2269;
wire x_2270;
wire x_2271;
wire x_2272;
wire x_2273;
wire x_2274;
wire x_2275;
wire x_2276;
wire x_2277;
wire x_2278;
wire x_2279;
wire x_2280;
wire x_2281;
wire x_2282;
wire x_2283;
wire x_2284;
wire x_2285;
wire x_2286;
wire x_2287;
wire x_2288;
wire x_2289;
wire x_2290;
wire x_2291;
wire x_2292;
wire x_2293;
wire x_2294;
wire x_2295;
wire x_2296;
wire x_2297;
wire x_2298;
wire x_2299;
wire x_2300;
wire x_2301;
wire x_2302;
wire x_2303;
wire x_2304;
wire x_2305;
wire x_2306;
wire x_2307;
wire x_2308;
wire x_2309;
wire x_2310;
wire x_2311;
wire x_2312;
wire x_2313;
wire x_2314;
wire x_2315;
wire x_2316;
wire x_2317;
wire x_2318;
wire x_2319;
wire x_2320;
wire x_2321;
wire x_2322;
wire x_2323;
wire x_2324;
wire x_2325;
wire x_2326;
wire x_2327;
wire x_2328;
wire x_2329;
wire x_2330;
wire x_2331;
wire x_2332;
wire x_2333;
wire x_2334;
wire x_2335;
wire x_2336;
wire x_2337;
wire x_2338;
wire x_2339;
wire x_2340;
wire x_2341;
wire x_2342;
wire x_2343;
wire x_2344;
wire x_2345;
wire x_2346;
wire x_2347;
wire x_2348;
wire x_2349;
wire x_2350;
wire x_2351;
wire x_2352;
wire x_2353;
wire x_2354;
wire x_2355;
wire x_2356;
wire x_2357;
wire x_2358;
wire x_2359;
wire x_2360;
wire x_2361;
wire x_2362;
wire x_2363;
wire x_2364;
wire x_2365;
wire x_2366;
wire x_2367;
wire x_2368;
wire x_2369;
wire x_2370;
wire x_2371;
wire x_2372;
wire x_2373;
wire x_2374;
wire x_2375;
wire x_2376;
wire x_2377;
wire x_2378;
wire x_2379;
wire x_2380;
wire x_2381;
wire x_2382;
wire x_2383;
wire x_2384;
wire x_2385;
wire x_2386;
wire x_2387;
wire x_2388;
wire x_2389;
wire x_2390;
wire x_2391;
wire x_2392;
wire x_2393;
wire x_2394;
wire x_2395;
wire x_2396;
wire x_2397;
wire x_2398;
wire x_2399;
wire x_2400;
wire x_2401;
wire x_2402;
wire x_2403;
wire x_2404;
wire x_2405;
wire x_2406;
wire x_2407;
wire x_2408;
wire x_2409;
wire x_2410;
wire x_2411;
wire x_2412;
wire x_2413;
wire x_2414;
wire x_2415;
wire x_2416;
wire x_2417;
wire x_2418;
wire x_2419;
wire x_2420;
wire x_2421;
wire x_2422;
wire x_2423;
wire x_2424;
wire x_2425;
wire x_2426;
wire x_2427;
wire x_2428;
wire x_2429;
wire x_2430;
wire x_2431;
wire x_2432;
wire x_2433;
wire x_2434;
wire x_2435;
wire x_2436;
wire x_2437;
wire x_2438;
wire x_2439;
wire x_2440;
wire x_2441;
wire x_2442;
wire x_2443;
wire x_2444;
wire x_2445;
wire x_2446;
wire x_2447;
wire x_2448;
wire x_2449;
wire x_2450;
wire x_2451;
wire x_2452;
wire x_2453;
wire x_2454;
wire x_2455;
wire x_2456;
wire x_2457;
wire x_2458;
wire x_2459;
wire x_2460;
wire x_2461;
wire x_2462;
wire x_2463;
wire x_2464;
wire x_2465;
wire x_2466;
wire x_2467;
wire x_2468;
wire x_2469;
wire x_2470;
wire x_2471;
wire x_2472;
wire x_2473;
wire x_2474;
wire x_2475;
wire x_2476;
wire x_2477;
wire x_2478;
wire x_2479;
wire x_2480;
wire x_2481;
wire x_2482;
wire x_2483;
wire x_2484;
wire x_2485;
wire x_2486;
wire x_2487;
wire x_2488;
wire x_2489;
wire x_2490;
wire x_2491;
wire x_2492;
wire x_2493;
wire x_2494;
wire x_2495;
wire x_2496;
wire x_2497;
wire x_2498;
wire x_2499;
wire x_2500;
wire x_2501;
wire x_2502;
wire x_2503;
wire x_2504;
wire x_2505;
wire x_2506;
wire x_2507;
wire x_2508;
wire x_2509;
wire x_2510;
wire x_2511;
wire x_2512;
wire x_2513;
wire x_2514;
wire x_2515;
wire x_2516;
wire x_2517;
wire x_2518;
wire x_2519;
wire x_2520;
wire x_2521;
wire x_2522;
wire x_2523;
wire x_2524;
wire x_2525;
wire x_2526;
wire x_2527;
wire x_2528;
wire x_2529;
wire x_2530;
wire x_2531;
wire x_2532;
wire x_2533;
wire x_2534;
wire x_2535;
wire x_2536;
wire x_2537;
wire x_2538;
wire x_2539;
wire x_2540;
wire x_2541;
wire x_2542;
wire x_2543;
wire x_2544;
wire x_2545;
wire x_2546;
wire x_2547;
wire x_2548;
wire x_2549;
wire x_2550;
wire x_2551;
wire x_2552;
wire x_2553;
wire x_2554;
wire x_2555;
wire x_2556;
wire x_2557;
wire x_2558;
wire x_2559;
wire x_2560;
wire x_2561;
wire x_2562;
wire x_2563;
wire x_2564;
wire x_2565;
wire x_2566;
wire x_2567;
wire x_2568;
wire x_2569;
wire x_2570;
wire x_2571;
wire x_2572;
wire x_2573;
wire x_2574;
wire x_2575;
wire x_2576;
wire x_2577;
wire x_2578;
wire x_2579;
wire x_2580;
wire x_2581;
wire x_2582;
wire x_2583;
wire x_2584;
wire x_2585;
wire x_2586;
wire x_2587;
wire x_2588;
wire x_2589;
wire x_2590;
wire x_2591;
wire x_2592;
wire x_2593;
wire x_2594;
wire x_2595;
wire x_2596;
wire x_2597;
wire x_2598;
wire x_2599;
wire x_2600;
wire x_2601;
wire x_2602;
wire x_2603;
wire x_2604;
wire x_2605;
wire x_2606;
wire x_2607;
wire x_2608;
wire x_2609;
wire x_2610;
wire x_2611;
wire x_2612;
wire x_2613;
wire x_2614;
wire x_2615;
wire x_2616;
wire x_2617;
wire x_2618;
wire x_2619;
wire x_2620;
wire x_2621;
wire x_2622;
wire x_2623;
wire x_2624;
wire x_2625;
wire x_2626;
wire x_2627;
wire x_2628;
wire x_2629;
wire x_2630;
wire x_2631;
wire x_2632;
wire x_2633;
wire x_2634;
wire x_2635;
wire x_2636;
wire x_2637;
wire x_2638;
wire x_2639;
wire x_2640;
wire x_2641;
wire x_2642;
wire x_2643;
wire x_2644;
wire x_2645;
wire x_2646;
wire x_2647;
wire x_2648;
wire x_2649;
wire x_2650;
wire x_2651;
wire x_2652;
wire x_2653;
wire x_2654;
wire x_2655;
wire x_2656;
wire x_2657;
wire x_2658;
wire x_2659;
wire x_2660;
wire x_2661;
wire x_2662;
wire x_2663;
wire x_2664;
wire x_2665;
wire x_2666;
wire x_2667;
wire x_2668;
wire x_2669;
wire x_2670;
wire x_2671;
wire x_2672;
wire x_2673;
wire x_2674;
wire x_2675;
wire x_2676;
wire x_2677;
wire x_2678;
wire x_2679;
wire x_2680;
wire x_2681;
wire x_2682;
wire x_2683;
wire x_2684;
wire x_2685;
wire x_2686;
wire x_2687;
wire x_2688;
wire x_2689;
wire x_2690;
wire x_2691;
wire x_2692;
wire x_2693;
wire x_2694;
wire x_2695;
wire x_2696;
wire x_2697;
wire x_2698;
wire x_2699;
wire x_2700;
wire x_2701;
wire x_2702;
wire x_2703;
wire x_2704;
wire x_2705;
wire x_2706;
wire x_2707;
wire x_2708;
wire x_2709;
wire x_2710;
wire x_2711;
wire x_2712;
wire x_2713;
wire x_2714;
wire x_2715;
wire x_2716;
wire x_2717;
wire x_2718;
wire x_2719;
wire x_2720;
wire x_2721;
wire x_2722;
wire x_2723;
wire x_2724;
wire x_2725;
wire x_2726;
wire x_2727;
wire x_2728;
wire x_2729;
wire x_2730;
wire x_2731;
wire x_2732;
wire x_2733;
wire x_2734;
wire x_2735;
wire x_2736;
wire x_2737;
wire x_2738;
wire x_2739;
wire x_2740;
wire x_2741;
wire x_2742;
wire x_2743;
wire x_2744;
wire x_2745;
wire x_2746;
wire x_2747;
wire x_2748;
wire x_2749;
wire x_2750;
wire x_2751;
wire x_2752;
wire x_2753;
wire x_2754;
wire x_2755;
wire x_2756;
wire x_2757;
wire x_2758;
wire x_2759;
wire x_2760;
wire x_2761;
wire x_2762;
wire x_2763;
wire x_2764;
wire x_2765;
wire x_2766;
wire x_2767;
wire x_2768;
wire x_2769;
wire x_2770;
wire x_2771;
wire x_2772;
wire x_2773;
wire x_2774;
wire x_2775;
wire x_2776;
wire x_2777;
wire x_2778;
wire x_2779;
wire x_2780;
wire x_2781;
wire x_2782;
wire x_2783;
wire x_2784;
wire x_2785;
wire x_2786;
wire x_2787;
wire x_2788;
wire x_2789;
wire x_2790;
wire x_2791;
wire x_2792;
wire x_2793;
wire x_2794;
wire x_2795;
wire x_2796;
wire x_2797;
wire x_2798;
wire x_2799;
wire x_2800;
wire x_2801;
wire x_2802;
wire x_2803;
wire x_2804;
wire x_2805;
wire x_2806;
wire x_2807;
wire x_2808;
wire x_2809;
wire x_2810;
wire x_2811;
wire x_2812;
wire x_2813;
wire x_2814;
wire x_2815;
wire x_2816;
wire x_2817;
wire x_2818;
wire x_2819;
wire x_2820;
wire x_2821;
wire x_2822;
wire x_2823;
wire x_2824;
wire x_2825;
wire x_2826;
wire x_2827;
wire x_2828;
wire x_2829;
wire x_2830;
wire x_2831;
wire x_2832;
wire x_2833;
wire x_2834;
wire x_2835;
wire x_2836;
wire x_2837;
wire x_2838;
wire x_2839;
wire x_2840;
wire x_2841;
wire x_2842;
wire x_2843;
wire x_2844;
wire x_2845;
wire x_2846;
wire x_2847;
wire x_2848;
wire x_2849;
wire x_2850;
wire x_2851;
wire x_2852;
wire x_2853;
wire x_2854;
wire x_2855;
wire x_2856;
wire x_2857;
wire x_2858;
wire x_2859;
wire x_2860;
wire x_2861;
wire x_2862;
wire x_2863;
wire x_2864;
wire x_2865;
wire x_2866;
wire x_2867;
wire x_2868;
wire x_2869;
wire x_2870;
wire x_2871;
wire x_2872;
wire x_2873;
wire x_2874;
wire x_2875;
wire x_2876;
wire x_2877;
wire x_2878;
wire x_2879;
wire x_2880;
wire x_2881;
wire x_2882;
wire x_2883;
wire x_2884;
wire x_2885;
wire x_2886;
wire x_2887;
wire x_2888;
wire x_2889;
wire x_2890;
wire x_2891;
wire x_2892;
wire x_2893;
wire x_2894;
wire x_2895;
wire x_2896;
wire x_2897;
wire x_2898;
wire x_2899;
wire x_2900;
wire x_2901;
wire x_2902;
wire x_2903;
wire x_2904;
wire x_2905;
wire x_2906;
wire x_2907;
wire x_2908;
wire x_2909;
wire x_2910;
wire x_2911;
wire x_2912;
wire x_2913;
wire x_2914;
wire x_2915;
wire x_2916;
wire x_2917;
wire x_2918;
wire x_2919;
wire x_2920;
wire x_2921;
wire x_2922;
wire x_2923;
wire x_2924;
wire x_2925;
wire x_2926;
wire x_2927;
wire x_2928;
wire x_2929;
wire x_2930;
wire x_2931;
wire x_2932;
wire x_2933;
wire x_2934;
wire x_2935;
wire x_2936;
wire x_2937;
wire x_2938;
wire x_2939;
wire x_2940;
wire x_2941;
wire x_2942;
wire x_2943;
wire x_2944;
wire x_2945;
wire x_2946;
wire x_2947;
wire x_2948;
wire x_2949;
wire x_2950;
wire x_2951;
wire x_2952;
wire x_2953;
wire x_2954;
wire x_2955;
wire x_2956;
wire x_2957;
wire x_2958;
wire x_2959;
wire x_2960;
wire x_2961;
wire x_2962;
wire x_2963;
wire x_2964;
wire x_2965;
wire x_2966;
wire x_2967;
wire x_2968;
wire x_2969;
wire x_2970;
wire x_2971;
wire x_2972;
wire x_2973;
wire x_2974;
wire x_2975;
wire x_2976;
wire x_2977;
wire x_2978;
wire x_2979;
wire x_2980;
wire x_2981;
wire x_2982;
wire x_2983;
wire x_2984;
wire x_2985;
wire x_2986;
wire x_2987;
wire x_2988;
wire x_2989;
wire x_2990;
wire x_2991;
wire x_2992;
wire x_2993;
wire x_2994;
wire x_2995;
wire x_2996;
wire x_2997;
wire x_2998;
wire x_2999;
wire x_3000;
wire x_3001;
wire x_3002;
wire x_3003;
wire x_3004;
wire x_3005;
wire x_3006;
wire x_3007;
wire x_3008;
wire x_3009;
wire x_3010;
wire x_3011;
wire x_3012;
wire x_3013;
wire x_3014;
wire x_3015;
wire x_3016;
wire x_3017;
wire x_3018;
wire x_3019;
wire x_3020;
wire x_3021;
wire x_3022;
wire x_3023;
wire x_3024;
wire x_3025;
wire x_3026;
wire x_3027;
wire x_3028;
wire x_3029;
wire x_3030;
wire x_3031;
wire x_3032;
wire x_3033;
wire x_3034;
wire x_3035;
wire x_3036;
wire x_3037;
wire x_3038;
wire x_3039;
wire x_3040;
wire x_3041;
wire x_3042;
wire x_3043;
wire x_3044;
wire x_3045;
wire x_3046;
wire x_3047;
wire x_3048;
wire x_3049;
wire x_3050;
wire x_3051;
wire x_3052;
wire x_3053;
wire x_3054;
wire x_3055;
wire x_3056;
wire x_3057;
wire x_3058;
wire x_3059;
wire x_3060;
wire x_3061;
wire x_3062;
wire x_3063;
wire x_3064;
wire x_3065;
wire x_3066;
wire x_3067;
wire x_3068;
wire x_3069;
wire x_3070;
wire x_3071;
wire x_3072;
wire x_3073;
wire x_3074;
wire x_3075;
wire x_3076;
wire x_3077;
wire x_3078;
wire x_3079;
wire x_3080;
wire x_3081;
wire x_3082;
wire x_3083;
wire x_3084;
wire x_3085;
wire x_3086;
wire x_3087;
wire x_3088;
wire x_3089;
wire x_3090;
wire x_3091;
wire x_3092;
wire x_3093;
wire x_3094;
wire x_3095;
wire x_3096;
wire x_3097;
wire x_3098;
wire x_3099;
wire x_3100;
wire x_3101;
wire x_3102;
wire x_3103;
wire x_3104;
wire x_3105;
wire x_3106;
wire x_3107;
wire x_3108;
wire x_3109;
wire x_3110;
wire x_3111;
wire x_3112;
wire x_3113;
wire x_3114;
wire x_3115;
wire x_3116;
wire x_3117;
wire x_3118;
wire x_3119;
wire x_3120;
wire x_3121;
wire x_3122;
wire x_3123;
wire x_3124;
wire x_3125;
wire x_3126;
wire x_3127;
wire x_3128;
wire x_3129;
wire x_3130;
wire x_3131;
wire x_3132;
wire x_3133;
wire x_3134;
wire x_3135;
wire x_3136;
wire x_3137;
wire x_3138;
wire x_3139;
wire x_3140;
wire x_3141;
wire x_3142;
wire x_3143;
wire x_3144;
wire x_3145;
wire x_3146;
wire x_3147;
wire x_3148;
wire x_3149;
wire x_3150;
wire x_3151;
wire x_3152;
wire x_3153;
wire x_3154;
wire x_3155;
wire x_3156;
wire x_3157;
wire x_3158;
wire x_3159;
wire x_3160;
wire x_3161;
wire x_3162;
wire x_3163;
wire x_3164;
wire x_3165;
wire x_3166;
wire x_3167;
wire x_3168;
wire x_3169;
wire x_3170;
wire x_3171;
wire x_3172;
wire x_3173;
wire x_3174;
wire x_3175;
wire x_3176;
wire x_3177;
wire x_3178;
wire x_3179;
wire x_3180;
wire x_3181;
wire x_3182;
wire x_3183;
wire x_3184;
wire x_3185;
wire x_3186;
wire x_3187;
wire x_3188;
wire x_3189;
wire x_3190;
wire x_3191;
wire x_3192;
wire x_3193;
wire x_3194;
wire x_3195;
wire x_3196;
wire x_3197;
wire x_3198;
wire x_3199;
wire x_3200;
wire x_3201;
wire x_3202;
wire x_3203;
wire x_3204;
wire x_3205;
wire x_3206;
wire x_3207;
wire x_3208;
wire x_3209;
wire x_3210;
wire x_3211;
wire x_3212;
wire x_3213;
wire x_3214;
wire x_3215;
wire x_3216;
wire x_3217;
wire x_3218;
wire x_3219;
wire x_3220;
wire x_3221;
wire x_3222;
wire x_3223;
wire x_3224;
wire x_3225;
wire x_3226;
wire x_3227;
wire x_3228;
wire x_3229;
wire x_3230;
wire x_3231;
wire x_3232;
wire x_3233;
wire x_3234;
wire x_3235;
wire x_3236;
wire x_3237;
wire x_3238;
wire x_3239;
wire x_3240;
wire x_3241;
wire x_3242;
wire x_3243;
wire x_3244;
wire x_3245;
wire x_3246;
wire x_3247;
wire x_3248;
wire x_3249;
wire x_3250;
wire x_3251;
wire x_3252;
wire x_3253;
wire x_3254;
wire x_3255;
wire x_3256;
wire x_3257;
wire x_3258;
wire x_3259;
wire x_3260;
wire x_3261;
wire x_3262;
wire x_3263;
wire x_3264;
wire x_3265;
wire x_3266;
wire x_3267;
wire x_3268;
wire x_3269;
wire x_3270;
wire x_3271;
wire x_3272;
wire x_3273;
wire x_3274;
wire x_3275;
wire x_3276;
wire x_3277;
wire x_3278;
wire x_3279;
wire x_3280;
wire x_3281;
wire x_3282;
wire x_3283;
wire x_3284;
wire x_3285;
wire x_3286;
wire x_3287;
wire x_3288;
wire x_3289;
wire x_3290;
wire x_3291;
wire x_3292;
wire x_3293;
wire x_3294;
wire x_3295;
wire x_3296;
wire x_3297;
wire x_3298;
wire x_3299;
wire x_3300;
wire x_3301;
wire x_3302;
wire x_3303;
wire x_3304;
wire x_3305;
wire x_3306;
wire x_3307;
wire x_3308;
wire x_3309;
wire x_3310;
wire x_3311;
wire x_3312;
wire x_3313;
wire x_3314;
wire x_3315;
wire x_3316;
wire x_3317;
wire x_3318;
wire x_3319;
wire x_3320;
wire x_3321;
wire x_3322;
wire x_3323;
wire x_3324;
wire x_3325;
wire x_3326;
wire x_3327;
wire x_3328;
wire x_3329;
wire x_3330;
wire x_3331;
wire x_3332;
wire x_3333;
wire x_3334;
wire x_3335;
wire x_3336;
wire x_3337;
wire x_3338;
wire x_3339;
wire x_3340;
wire x_3341;
wire x_3342;
wire x_3343;
wire x_3344;
wire x_3345;
wire x_3346;
wire x_3347;
wire x_3348;
wire x_3349;
wire x_3350;
wire x_3351;
wire x_3352;
wire x_3353;
wire x_3354;
wire x_3355;
wire x_3356;
wire x_3357;
wire x_3358;
wire x_3359;
wire x_3360;
wire x_3361;
wire x_3362;
wire x_3363;
wire x_3364;
wire x_3365;
wire x_3366;
wire x_3367;
wire x_3368;
wire x_3369;
wire x_3370;
wire x_3371;
wire x_3372;
wire x_3373;
wire x_3374;
wire x_3375;
wire x_3376;
wire x_3377;
wire x_3378;
wire x_3379;
wire x_3380;
wire x_3381;
wire x_3382;
wire x_3383;
wire x_3384;
wire x_3385;
wire x_3386;
wire x_3387;
wire x_3388;
wire x_3389;
wire x_3390;
wire x_3391;
wire x_3392;
wire x_3393;
wire x_3394;
wire x_3395;
wire x_3396;
wire x_3397;
wire x_3398;
wire x_3399;
wire x_3400;
wire x_3401;
wire x_3402;
wire x_3403;
wire x_3404;
wire x_3405;
wire x_3406;
wire x_3407;
wire x_3408;
wire x_3409;
wire x_3410;
wire x_3411;
wire x_3412;
wire x_3413;
wire x_3414;
wire x_3415;
wire x_3416;
wire x_3417;
wire x_3418;
wire x_3419;
wire x_3420;
wire x_3421;
wire x_3422;
wire x_3423;
wire x_3424;
wire x_3425;
wire x_3426;
wire x_3427;
wire x_3428;
wire x_3429;
wire x_3430;
wire x_3431;
wire x_3432;
wire x_3433;
wire x_3434;
wire x_3435;
wire x_3436;
wire x_3437;
wire x_3438;
wire x_3439;
wire x_3440;
wire x_3441;
wire x_3442;
wire x_3443;
wire x_3444;
wire x_3445;
wire x_3446;
wire x_3447;
wire x_3448;
wire x_3449;
wire x_3450;
wire x_3451;
wire x_3452;
wire x_3453;
wire x_3454;
wire x_3455;
wire x_3456;
wire x_3457;
wire x_3458;
wire x_3459;
wire x_3460;
wire x_3461;
wire x_3462;
wire x_3463;
wire x_3464;
wire x_3465;
wire x_3466;
wire x_3467;
wire x_3468;
wire x_3469;
wire x_3470;
wire x_3471;
wire x_3472;
wire x_3473;
wire x_3474;
wire x_3475;
wire x_3476;
wire x_3477;
wire x_3478;
wire x_3479;
wire x_3480;
wire x_3481;
wire x_3482;
wire x_3483;
wire x_3484;
wire x_3485;
wire x_3486;
wire x_3487;
wire x_3488;
wire x_3489;
wire x_3490;
wire x_3491;
wire x_3492;
wire x_3493;
wire x_3494;
wire x_3495;
wire x_3496;
wire x_3497;
wire x_3498;
wire x_3499;
wire x_3500;
wire x_3501;
wire x_3502;
wire x_3503;
wire x_3504;
wire x_3505;
wire x_3506;
wire x_3507;
wire x_3508;
wire x_3509;
wire x_3510;
wire x_3511;
wire x_3512;
wire x_3513;
wire x_3514;
wire x_3515;
wire x_3516;
wire x_3517;
wire x_3518;
wire x_3519;
wire x_3520;
wire x_3521;
wire x_3522;
wire x_3523;
wire x_3524;
wire x_3525;
wire x_3526;
wire x_3527;
wire x_3528;
wire x_3529;
wire x_3530;
wire x_3531;
wire x_3532;
wire x_3533;
wire x_3534;
wire x_3535;
wire x_3536;
wire x_3537;
wire x_3538;
wire x_3539;
wire x_3540;
wire x_3541;
wire x_3542;
wire x_3543;
wire x_3544;
wire x_3545;
wire x_3546;
wire x_3547;
wire x_3548;
wire x_3549;
wire x_3550;
wire x_3551;
wire x_3552;
wire x_3553;
wire x_3554;
wire x_3555;
wire x_3556;
wire x_3557;
wire x_3558;
wire x_3559;
wire x_3560;
wire x_3561;
wire x_3562;
wire x_3563;
wire x_3564;
wire x_3565;
wire x_3566;
wire x_3567;
wire x_3568;
wire x_3569;
wire x_3570;
wire x_3571;
wire x_3572;
wire x_3573;
wire x_3574;
wire x_3575;
wire x_3576;
wire x_3577;
wire x_3578;
wire x_3579;
wire x_3580;
wire x_3581;
wire x_3582;
wire x_3583;
wire x_3584;
wire x_3585;
wire x_3586;
wire x_3587;
wire x_3588;
wire x_3589;
wire x_3590;
wire x_3591;
wire x_3592;
wire x_3593;
wire x_3594;
wire x_3595;
wire x_3596;
wire x_3597;
wire x_3598;
wire x_3599;
wire x_3600;
wire x_3601;
wire x_3602;
wire x_3603;
wire x_3604;
wire x_3605;
wire x_3606;
wire x_3607;
wire x_3608;
wire x_3609;
wire x_3610;
wire x_3611;
wire x_3612;
wire x_3613;
wire x_3614;
wire x_3615;
wire x_3616;
wire x_3617;
wire x_3618;
wire x_3619;
wire x_3620;
wire x_3621;
wire x_3622;
wire x_3623;
wire x_3624;
wire x_3625;
wire x_3626;
wire x_3627;
wire x_3628;
wire x_3629;
wire x_3630;
wire x_3631;
wire x_3632;
wire x_3633;
wire x_3634;
wire x_3635;
wire x_3636;
wire x_3637;
wire x_3638;
wire x_3639;
wire x_3640;
wire x_3641;
wire x_3642;
wire x_3643;
wire x_3644;
wire x_3645;
wire x_3646;
wire x_3647;
wire x_3648;
wire x_3649;
wire x_3650;
wire x_3651;
wire x_3652;
wire x_3653;
wire x_3654;
wire x_3655;
wire x_3656;
wire x_3657;
wire x_3658;
wire x_3659;
wire x_3660;
wire x_3661;
wire x_3662;
wire x_3663;
wire x_3664;
wire x_3665;
wire x_3666;
wire x_3667;
wire x_3668;
wire x_3669;
wire x_3670;
wire x_3671;
wire x_3672;
wire x_3673;
wire x_3674;
wire x_3675;
wire x_3676;
wire x_3677;
wire x_3678;
wire x_3679;
wire x_3680;
wire x_3681;
wire x_3682;
wire x_3683;
wire x_3684;
wire x_3685;
wire x_3686;
wire x_3687;
wire x_3688;
wire x_3689;
wire x_3690;
wire x_3691;
wire x_3692;
wire x_3693;
wire x_3694;
wire x_3695;
wire x_3696;
wire x_3697;
wire x_3698;
wire x_3699;
wire x_3700;
wire x_3701;
wire x_3702;
wire x_3703;
wire x_3704;
wire x_3705;
wire x_3706;
wire x_3707;
wire x_3708;
wire x_3709;
wire x_3710;
wire x_3711;
wire x_3712;
wire x_3713;
wire x_3714;
wire x_3715;
wire x_3716;
wire x_3717;
wire x_3718;
wire x_3719;
wire x_3720;
wire x_3721;
wire x_3722;
wire x_3723;
wire x_3724;
wire x_3725;
wire x_3726;
wire x_3727;
wire x_3728;
wire x_3729;
wire x_3730;
wire x_3731;
wire x_3732;
wire x_3733;
wire x_3734;
wire x_3735;
wire x_3736;
wire x_3737;
wire x_3738;
wire x_3739;
wire x_3740;
wire x_3741;
wire x_3742;
wire x_3743;
wire x_3744;
wire x_3745;
wire x_3746;
wire x_3747;
wire x_3748;
wire x_3749;
wire x_3750;
wire x_3751;
wire x_3752;
wire x_3753;
wire x_3754;
wire x_3755;
wire x_3756;
wire x_3757;
wire x_3758;
wire x_3759;
wire x_3760;
wire x_3761;
wire x_3762;
wire x_3763;
wire x_3764;
wire x_3765;
wire x_3766;
wire x_3767;
wire x_3768;
wire x_3769;
wire x_3770;
wire x_3771;
wire x_3772;
wire x_3773;
wire x_3774;
wire x_3775;
wire x_3776;
wire x_3777;
wire x_3778;
wire x_3779;
wire x_3780;
wire x_3781;
wire x_3782;
wire x_3783;
wire x_3784;
wire x_3785;
wire x_3786;
wire x_3787;
wire x_3788;
wire x_3789;
wire x_3790;
wire x_3791;
wire x_3792;
wire x_3793;
wire x_3794;
wire x_3795;
wire x_3796;
wire x_3797;
wire x_3798;
wire x_3799;
wire x_3800;
wire x_3801;
wire x_3802;
wire x_3803;
wire x_3804;
wire x_3805;
wire x_3806;
wire x_3807;
wire x_3808;
wire x_3809;
wire x_3810;
wire x_3811;
wire x_3812;
wire x_3813;
wire x_3814;
wire x_3815;
wire x_3816;
wire x_3817;
wire x_3818;
wire x_3819;
wire x_3820;
wire x_3821;
wire x_3822;
wire x_3823;
wire x_3824;
wire x_3825;
wire x_3826;
wire x_3827;
wire x_3828;
wire x_3829;
wire x_3830;
wire x_3831;
wire x_3832;
wire x_3833;
wire x_3834;
wire x_3835;
wire x_3836;
wire x_3837;
wire x_3838;
wire x_3839;
wire x_3840;
wire x_3841;
wire x_3842;
wire x_3843;
wire x_3844;
wire x_3845;
wire x_3846;
wire x_3847;
wire x_3848;
wire x_3849;
wire x_3850;
wire x_3851;
wire x_3852;
wire x_3853;
wire x_3854;
wire x_3855;
wire x_3856;
wire x_3857;
wire x_3858;
wire x_3859;
wire x_3860;
wire x_3861;
wire x_3862;
wire x_3863;
wire x_3864;
wire x_3865;
wire x_3866;
wire x_3867;
wire x_3868;
wire x_3869;
wire x_3870;
wire x_3871;
wire x_3872;
wire x_3873;
wire x_3874;
wire x_3875;
wire x_3876;
wire x_3877;
wire x_3878;
wire x_3879;
wire x_3880;
wire x_3881;
wire x_3882;
wire x_3883;
wire x_3884;
wire x_3885;
wire x_3886;
wire x_3887;
wire x_3888;
wire x_3889;
wire x_3890;
wire x_3891;
wire x_3892;
wire x_3893;
wire x_3894;
wire x_3895;
wire x_3896;
wire x_3897;
wire x_3898;
wire x_3899;
wire x_3900;
wire x_3901;
wire x_3902;
wire x_3903;
wire x_3904;
wire x_3905;
wire x_3906;
wire x_3907;
wire x_3908;
wire x_3909;
wire x_3910;
wire x_3911;
wire x_3912;
wire x_3913;
wire x_3914;
wire x_3915;
wire x_3916;
wire x_3917;
wire x_3918;
wire x_3919;
wire x_3920;
wire x_3921;
wire x_3922;
wire x_3923;
wire x_3924;
wire x_3925;
wire x_3926;
wire x_3927;
wire x_3928;
wire x_3929;
wire x_3930;
wire x_3931;
wire x_3932;
wire x_3933;
wire x_3934;
wire x_3935;
wire x_3936;
wire x_3937;
wire x_3938;
wire x_3939;
wire x_3940;
wire x_3941;
wire x_3942;
wire x_3943;
wire x_3944;
wire x_3945;
wire x_3946;
wire x_3947;
wire x_3948;
wire x_3949;
wire x_3950;
wire x_3951;
wire x_3952;
wire x_3953;
wire x_3954;
wire x_3955;
wire x_3956;
wire x_3957;
wire x_3958;
wire x_3959;
wire x_3960;
wire x_3961;
wire x_3962;
wire x_3963;
wire x_3964;
wire x_3965;
wire x_3966;
wire x_3967;
wire x_3968;
wire x_3969;
wire x_3970;
wire x_3971;
wire x_3972;
wire x_3973;
wire x_3974;
wire x_3975;
wire x_3976;
wire x_3977;
wire x_3978;
wire x_3979;
wire x_3980;
wire x_3981;
wire x_3982;
wire x_3983;
wire x_3984;
wire x_3985;
wire x_3986;
wire x_3987;
wire x_3988;
wire x_3989;
wire x_3990;
wire x_3991;
wire x_3992;
wire x_3993;
wire x_3994;
wire x_3995;
wire x_3996;
wire x_3997;
wire x_3998;
wire x_3999;
wire x_4000;
wire x_4001;
wire x_4002;
wire x_4003;
wire x_4004;
wire x_4005;
wire x_4006;
wire x_4007;
wire x_4008;
wire x_4009;
wire x_4010;
wire x_4011;
wire x_4012;
wire x_4013;
wire x_4014;
wire x_4015;
wire x_4016;
wire x_4017;
wire x_4018;
wire x_4019;
wire x_4020;
wire x_4021;
wire x_4022;
wire x_4023;
wire x_4024;
wire x_4025;
wire x_4026;
wire x_4027;
wire x_4028;
wire x_4029;
wire x_4030;
wire x_4031;
wire x_4032;
wire x_4033;
wire x_4034;
wire x_4035;
wire x_4036;
wire x_4037;
wire x_4038;
wire x_4039;
wire x_4040;
wire x_4041;
wire x_4042;
wire x_4043;
wire x_4044;
wire x_4045;
wire x_4046;
wire x_4047;
wire x_4048;
wire x_4049;
wire x_4050;
wire x_4051;
wire x_4052;
wire x_4053;
wire x_4054;
wire x_4055;
wire x_4056;
wire x_4057;
wire x_4058;
wire x_4059;
wire x_4060;
wire x_4061;
wire x_4062;
wire x_4063;
wire x_4064;
wire x_4065;
wire x_4066;
wire x_4067;
wire x_4068;
wire x_4069;
wire x_4070;
wire x_4071;
wire x_4072;
wire x_4073;
wire x_4074;
wire x_4075;
wire x_4076;
wire x_4077;
wire x_4078;
wire x_4079;
wire x_4080;
wire x_4081;
wire x_4082;
wire x_4083;
wire x_4084;
wire x_4085;
wire x_4086;
wire x_4087;
wire x_4088;
wire x_4089;
wire x_4090;
wire x_4091;
wire x_4092;
wire x_4093;
wire x_4094;
wire x_4095;
wire x_4096;
wire x_4097;
wire x_4098;
wire x_4099;
wire x_4100;
wire x_4101;
wire x_4102;
wire x_4103;
wire x_4104;
wire x_4105;
wire x_4106;
wire x_4107;
wire x_4108;
wire x_4109;
wire x_4110;
wire x_4111;
wire x_4112;
wire x_4113;
wire x_4114;
wire x_4115;
wire x_4116;
wire x_4117;
wire x_4118;
wire x_4119;
wire x_4120;
wire x_4121;
wire x_4122;
wire x_4123;
wire x_4124;
wire x_4125;
wire x_4126;
wire x_4127;
wire x_4128;
wire x_4129;
wire x_4130;
wire x_4131;
wire x_4132;
wire x_4133;
wire x_4134;
wire x_4135;
wire x_4136;
wire x_4137;
wire x_4138;
wire x_4139;
wire x_4140;
wire x_4141;
wire x_4142;
wire x_4143;
wire x_4144;
wire x_4145;
wire x_4146;
wire x_4147;
wire x_4148;
wire x_4149;
wire x_4150;
wire x_4151;
wire x_4152;
wire x_4153;
wire x_4154;
wire x_4155;
wire x_4156;
wire x_4157;
wire x_4158;
wire x_4159;
wire x_4160;
wire x_4161;
wire x_4162;
wire x_4163;
wire x_4164;
wire x_4165;
wire x_4166;
wire x_4167;
wire x_4168;
wire x_4169;
wire x_4170;
wire x_4171;
wire x_4172;
wire x_4173;
wire x_4174;
wire x_4175;
wire x_4176;
wire x_4177;
wire x_4178;
wire x_4179;
wire x_4180;
wire x_4181;
wire x_4182;
wire x_4183;
wire x_4184;
wire x_4185;
wire x_4186;
wire x_4187;
wire x_4188;
wire x_4189;
wire x_4190;
wire x_4191;
wire x_4192;
wire x_4193;
wire x_4194;
wire x_4195;
wire x_4196;
wire x_4197;
wire x_4198;
wire x_4199;
wire x_4200;
wire x_4201;
wire x_4202;
wire x_4203;
wire x_4204;
wire x_4205;
wire x_4206;
wire x_4207;
wire x_4208;
wire x_4209;
wire x_4210;
wire x_4211;
wire x_4212;
wire x_4213;
wire x_4214;
wire x_4215;
wire x_4216;
wire x_4217;
wire x_4218;
wire x_4219;
wire x_4220;
wire x_4221;
wire x_4222;
wire x_4223;
wire x_4224;
wire x_4225;
wire x_4226;
wire x_4227;
wire x_4228;
wire x_4229;
wire x_4230;
wire x_4231;
wire x_4232;
wire x_4233;
wire x_4234;
wire x_4235;
wire x_4236;
wire x_4237;
wire x_4238;
wire x_4239;
wire x_4240;
wire x_4241;
wire x_4242;
wire x_4243;
wire x_4244;
wire x_4245;
wire x_4246;
wire x_4247;
wire x_4248;
wire x_4249;
wire x_4250;
wire x_4251;
wire x_4252;
wire x_4253;
wire x_4254;
wire x_4255;
wire x_4256;
wire x_4257;
wire x_4258;
wire x_4259;
wire x_4260;
wire x_4261;
wire x_4262;
wire x_4263;
wire x_4264;
wire x_4265;
wire x_4266;
wire x_4267;
wire x_4268;
wire x_4269;
wire x_4270;
wire x_4271;
wire x_4272;
wire x_4273;
wire x_4274;
wire x_4275;
wire x_4276;
wire x_4277;
wire x_4278;
wire x_4279;
wire x_4280;
wire x_4281;
wire x_4282;
wire x_4283;
wire x_4284;
wire x_4285;
wire x_4286;
wire x_4287;
wire x_4288;
wire x_4289;
wire x_4290;
wire x_4291;
wire x_4292;
wire x_4293;
wire x_4294;
wire x_4295;
wire x_4296;
wire x_4297;
wire x_4298;
wire x_4299;
wire x_4300;
wire x_4301;
wire x_4302;
wire x_4303;
wire x_4304;
wire x_4305;
wire x_4306;
wire x_4307;
wire x_4308;
wire x_4309;
wire x_4310;
wire x_4311;
wire x_4312;
wire x_4313;
wire x_4314;
wire x_4315;
wire x_4316;
wire x_4317;
wire x_4318;
wire x_4319;
wire x_4320;
wire x_4321;
wire x_4322;
wire x_4323;
wire x_4324;
wire x_4325;
wire x_4326;
wire x_4327;
wire x_4328;
wire x_4329;
wire x_4330;
wire x_4331;
wire x_4332;
wire x_4333;
wire x_4334;
wire x_4335;
wire x_4336;
wire x_4337;
wire x_4338;
wire x_4339;
wire x_4340;
wire x_4341;
wire x_4342;
wire x_4343;
wire x_4344;
wire x_4345;
wire x_4346;
wire x_4347;
wire x_4348;
wire x_4349;
wire x_4350;
wire x_4351;
wire x_4352;
wire x_4353;
wire x_4354;
wire x_4355;
wire x_4356;
wire x_4357;
wire x_4358;
wire x_4359;
wire x_4360;
wire x_4361;
wire x_4362;
wire x_4363;
wire x_4364;
wire x_4365;
wire x_4366;
wire x_4367;
wire x_4368;
wire x_4369;
wire x_4370;
wire x_4371;
wire x_4372;
wire x_4373;
wire x_4374;
wire x_4375;
wire x_4376;
wire x_4377;
wire x_4378;
wire x_4379;
wire x_4380;
wire x_4381;
wire x_4382;
wire x_4383;
wire x_4384;
wire x_4385;
wire x_4386;
wire x_4387;
wire x_4388;
wire x_4389;
wire x_4390;
wire x_4391;
wire x_4392;
wire x_4393;
wire x_4394;
wire x_4395;
wire x_4396;
wire x_4397;
wire x_4398;
wire x_4399;
wire x_4400;
wire x_4401;
wire x_4402;
wire x_4403;
wire x_4404;
wire x_4405;
wire x_4406;
wire x_4407;
wire x_4408;
wire x_4409;
wire x_4410;
wire x_4411;
wire x_4412;
wire x_4413;
wire x_4414;
wire x_4415;
wire x_4416;
wire x_4417;
wire x_4418;
wire x_4419;
wire x_4420;
wire x_4421;
wire x_4422;
wire x_4423;
wire x_4424;
wire x_4425;
wire x_4426;
wire x_4427;
wire x_4428;
wire x_4429;
wire x_4430;
wire x_4431;
wire x_4432;
wire x_4433;
wire x_4434;
wire x_4435;
wire x_4436;
wire x_4437;
wire x_4438;
wire x_4439;
wire x_4440;
wire x_4441;
wire x_4442;
wire x_4443;
wire x_4444;
wire x_4445;
wire x_4446;
wire x_4447;
wire x_4448;
wire x_4449;
wire x_4450;
wire x_4451;
wire x_4452;
wire x_4453;
wire x_4454;
wire x_4455;
wire x_4456;
wire x_4457;
wire x_4458;
wire x_4459;
wire x_4460;
wire x_4461;
wire x_4462;
wire x_4463;
wire x_4464;
wire x_4465;
wire x_4466;
wire x_4467;
wire x_4468;
wire x_4469;
wire x_4470;
wire x_4471;
wire x_4472;
wire x_4473;
wire x_4474;
wire x_4475;
wire x_4476;
wire x_4477;
wire x_4478;
wire x_4479;
wire x_4480;
wire x_4481;
wire x_4482;
wire x_4483;
wire x_4484;
wire x_4485;
wire x_4486;
wire x_4487;
wire x_4488;
wire x_4489;
wire x_4490;
wire x_4491;
wire x_4492;
wire x_4493;
wire x_4494;
wire x_4495;
wire x_4496;
wire x_4497;
wire x_4498;
wire x_4499;
wire x_4500;
wire x_4501;
wire x_4502;
wire x_4503;
wire x_4504;
wire x_4505;
wire x_4506;
wire x_4507;
wire x_4508;
wire x_4509;
wire x_4510;
wire x_4511;
wire x_4512;
wire x_4513;
wire x_4514;
wire x_4515;
wire x_4516;
wire x_4517;
wire x_4518;
wire x_4519;
wire x_4520;
wire x_4521;
wire x_4522;
wire x_4523;
wire x_4524;
wire x_4525;
wire x_4526;
wire x_4527;
wire x_4528;
wire x_4529;
wire x_4530;
wire x_4531;
wire x_4532;
wire x_4533;
wire x_4534;
wire x_4535;
wire x_4536;
wire x_4537;
wire x_4538;
wire x_4539;
wire x_4540;
wire x_4541;
wire x_4542;
wire x_4543;
wire x_4544;
wire x_4545;
wire x_4546;
wire x_4547;
wire x_4548;
wire x_4549;
wire x_4550;
wire x_4551;
wire x_4552;
wire x_4553;
wire x_4554;
wire x_4555;
wire x_4556;
wire x_4557;
wire x_4558;
wire x_4559;
wire x_4560;
wire x_4561;
wire x_4562;
wire x_4563;
wire x_4564;
wire x_4565;
wire x_4566;
wire x_4567;
wire x_4568;
wire x_4569;
wire x_4570;
wire x_4571;
wire x_4572;
wire x_4573;
wire x_4574;
wire x_4575;
wire x_4576;
wire x_4577;
wire x_4578;
wire x_4579;
wire x_4580;
wire x_4581;
wire x_4582;
wire x_4583;
wire x_4584;
wire x_4585;
wire x_4586;
wire x_4587;
wire x_4588;
wire x_4589;
wire x_4590;
wire x_4591;
wire x_4592;
wire x_4593;
wire x_4594;
wire x_4595;
wire x_4596;
wire x_4597;
wire x_4598;
wire x_4599;
wire x_4600;
wire x_4601;
wire x_4602;
wire x_4603;
wire x_4604;
wire x_4605;
wire x_4606;
wire x_4607;
wire x_4608;
wire x_4609;
wire x_4610;
wire x_4611;
wire x_4612;
wire x_4613;
wire x_4614;
wire x_4615;
wire x_4616;
wire x_4617;
wire x_4618;
wire x_4619;
wire x_4620;
wire x_4621;
wire x_4622;
wire x_4623;
wire x_4624;
wire x_4625;
wire x_4626;
wire x_4627;
wire x_4628;
wire x_4629;
wire x_4630;
wire x_4631;
wire x_4632;
wire x_4633;
wire x_4634;
wire x_4635;
wire x_4636;
wire x_4637;
wire x_4638;
wire x_4639;
wire x_4640;
wire x_4641;
wire x_4642;
wire x_4643;
wire x_4644;
wire x_4645;
wire x_4646;
wire x_4647;
wire x_4648;
wire x_4649;
wire x_4650;
wire x_4651;
wire x_4652;
wire x_4653;
wire x_4654;
wire x_4655;
wire x_4656;
wire x_4657;
wire x_4658;
wire x_4659;
wire x_4660;
wire x_4661;
wire x_4662;
wire x_4663;
wire x_4664;
wire x_4665;
wire x_4666;
wire x_4667;
wire x_4668;
wire x_4669;
wire x_4670;
wire x_4671;
wire x_4672;
wire x_4673;
wire x_4674;
wire x_4675;
wire x_4676;
wire x_4677;
wire x_4678;
wire x_4679;
wire x_4680;
wire x_4681;
wire x_4682;
wire x_4683;
wire x_4684;
wire x_4685;
wire x_4686;
wire x_4687;
wire x_4688;
wire x_4689;
wire x_4690;
wire x_4691;
wire x_4692;
wire x_4693;
wire x_4694;
wire x_4695;
wire x_4696;
wire x_4697;
wire x_4698;
wire x_4699;
wire x_4700;
wire x_4701;
wire x_4702;
wire x_4703;
wire x_4704;
wire x_4705;
wire x_4706;
wire x_4707;
wire x_4708;
wire x_4709;
wire x_4710;
wire x_4711;
wire x_4712;
wire x_4713;
wire x_4714;
wire x_4715;
wire x_4716;
wire x_4717;
wire x_4718;
wire x_4719;
wire x_4720;
wire x_4721;
wire x_4722;
wire x_4723;
wire x_4724;
wire x_4725;
wire x_4726;
wire x_4727;
wire x_4728;
wire x_4729;
wire x_4730;
wire x_4731;
wire x_4732;
wire x_4733;
wire x_4734;
wire x_4735;
wire x_4736;
wire x_4737;
wire x_4738;
wire x_4739;
wire x_4740;
wire x_4741;
wire x_4742;
wire x_4743;
wire x_4744;
wire x_4745;
wire x_4746;
wire x_4747;
wire x_4748;
wire x_4749;
wire x_4750;
wire x_4751;
wire x_4752;
wire x_4753;
wire x_4754;
wire x_4755;
wire x_4756;
wire x_4757;
wire x_4758;
wire x_4759;
wire x_4760;
wire x_4761;
wire x_4762;
wire x_4763;
wire x_4764;
wire x_4765;
wire x_4766;
wire x_4767;
wire x_4768;
wire x_4769;
wire x_4770;
wire x_4771;
wire x_4772;
wire x_4773;
wire x_4774;
wire x_4775;
wire x_4776;
wire x_4777;
wire x_4778;
wire x_4779;
wire x_4780;
wire x_4781;
wire x_4782;
wire x_4783;
wire x_4784;
wire x_4785;
wire x_4786;
wire x_4787;
wire x_4788;
wire x_4789;
wire x_4790;
wire x_4791;
wire x_4792;
wire x_4793;
wire x_4794;
wire x_4795;
wire x_4796;
wire x_4797;
wire x_4798;
wire x_4799;
wire x_4800;
wire x_4801;
wire x_4802;
wire x_4803;
wire x_4804;
wire x_4805;
wire x_4806;
wire x_4807;
wire x_4808;
wire x_4809;
wire x_4810;
wire x_4811;
wire x_4812;
wire x_4813;
wire x_4814;
wire x_4815;
wire x_4816;
wire x_4817;
wire x_4818;
wire x_4819;
wire x_4820;
wire x_4821;
wire x_4822;
wire x_4823;
wire x_4824;
wire x_4825;
wire x_4826;
wire x_4827;
wire x_4828;
wire x_4829;
wire x_4830;
wire x_4831;
wire x_4832;
wire x_4833;
wire x_4834;
wire x_4835;
wire x_4836;
wire x_4837;
wire x_4838;
wire x_4839;
wire x_4840;
wire x_4841;
wire x_4842;
wire x_4843;
wire x_4844;
wire x_4845;
wire x_4846;
wire x_4847;
wire x_4848;
wire x_4849;
wire x_4850;
wire x_4851;
wire x_4852;
wire x_4853;
wire x_4854;
wire x_4855;
wire x_4856;
wire x_4857;
wire x_4858;
wire x_4859;
wire x_4860;
wire x_4861;
wire x_4862;
wire x_4863;
wire x_4864;
wire x_4865;
wire x_4866;
wire x_4867;
wire x_4868;
wire x_4869;
wire x_4870;
wire x_4871;
wire x_4872;
wire x_4873;
wire x_4874;
wire x_4875;
wire x_4876;
wire x_4877;
wire x_4878;
wire x_4879;
wire x_4880;
wire x_4881;
wire x_4882;
wire x_4883;
wire x_4884;
wire x_4885;
wire x_4886;
wire x_4887;
wire x_4888;
wire x_4889;
wire x_4890;
wire x_4891;
wire x_4892;
wire x_4893;
wire x_4894;
wire x_4895;
wire x_4896;
wire x_4897;
wire x_4898;
wire x_4899;
wire x_4900;
wire x_4901;
wire x_4902;
wire x_4903;
wire x_4904;
wire x_4905;
wire x_4906;
wire x_4907;
wire x_4908;
wire x_4909;
wire x_4910;
wire x_4911;
wire x_4912;
wire x_4913;
wire x_4914;
wire x_4915;
wire x_4916;
wire x_4917;
wire x_4918;
wire x_4919;
wire x_4920;
wire x_4921;
wire x_4922;
wire x_4923;
wire x_4924;
wire x_4925;
wire x_4926;
wire x_4927;
wire x_4928;
wire x_4929;
wire x_4930;
wire x_4931;
wire x_4932;
wire x_4933;
wire x_4934;
wire x_4935;
wire x_4936;
wire x_4937;
wire x_4938;
wire x_4939;
wire x_4940;
wire x_4941;
wire x_4942;
wire x_4943;
wire x_4944;
wire x_4945;
wire x_4946;
wire x_4947;
wire x_4948;
wire x_4949;
wire x_4950;
wire x_4951;
wire x_4952;
wire x_4953;
wire x_4954;
wire x_4955;
wire x_4956;
wire x_4957;
wire x_4958;
wire x_4959;
wire x_4960;
wire x_4961;
wire x_4962;
wire x_4963;
wire x_4964;
wire x_4965;
wire x_4966;
wire x_4967;
wire x_4968;
wire x_4969;
wire x_4970;
wire x_4971;
wire x_4972;
wire x_4973;
wire x_4974;
wire x_4975;
wire x_4976;
wire x_4977;
wire x_4978;
wire x_4979;
wire x_4980;
wire x_4981;
wire x_4982;
wire x_4983;
wire x_4984;
wire x_4985;
wire x_4986;
wire x_4987;
wire x_4988;
wire x_4989;
wire x_4990;
wire x_4991;
wire x_4992;
wire x_4993;
wire x_4994;
wire x_4995;
wire x_4996;
wire x_4997;
wire x_4998;
wire x_4999;
wire x_5000;
wire x_5001;
wire x_5002;
wire x_5003;
wire x_5004;
wire x_5005;
wire x_5006;
wire x_5007;
wire x_5008;
wire x_5009;
wire x_5010;
wire x_5011;
wire x_5012;
wire x_5013;
wire x_5014;
wire x_5015;
wire x_5016;
wire x_5017;
wire x_5018;
wire x_5019;
wire x_5020;
wire x_5021;
wire x_5022;
wire x_5023;
wire x_5024;
wire x_5025;
wire x_5026;
wire x_5027;
wire x_5028;
wire x_5029;
wire x_5030;
wire x_5031;
wire x_5032;
wire x_5033;
wire x_5034;
wire x_5035;
wire x_5036;
wire x_5037;
wire x_5038;
wire x_5039;
wire x_5040;
wire x_5041;
wire x_5042;
wire x_5043;
wire x_5044;
wire x_5045;
wire x_5046;
wire x_5047;
wire x_5048;
wire x_5049;
wire x_5050;
wire x_5051;
wire x_5052;
wire x_5053;
wire x_5054;
wire x_5055;
wire x_5056;
wire x_5057;
wire x_5058;
wire x_5059;
wire x_5060;
wire x_5061;
wire x_5062;
wire x_5063;
wire x_5064;
wire x_5065;
wire x_5066;
wire x_5067;
wire x_5068;
wire x_5069;
wire x_5070;
wire x_5071;
wire x_5072;
wire x_5073;
wire x_5074;
wire x_5075;
wire x_5076;
wire x_5077;
wire x_5078;
wire x_5079;
wire x_5080;
wire x_5081;
wire x_5082;
wire x_5083;
wire x_5084;
wire x_5085;
wire x_5086;
wire x_5087;
wire x_5088;
wire x_5089;
wire x_5090;
wire x_5091;
wire x_5092;
wire x_5093;
wire x_5094;
wire x_5095;
wire x_5096;
wire x_5097;
wire x_5098;
wire x_5099;
wire x_5100;
wire x_5101;
wire x_5102;
wire x_5103;
wire x_5104;
wire x_5105;
wire x_5106;
wire x_5107;
wire x_5108;
wire x_5109;
wire x_5110;
wire x_5111;
wire x_5112;
wire x_5113;
wire x_5114;
wire x_5115;
wire x_5116;
wire x_5117;
wire x_5118;
wire x_5119;
wire x_5120;
wire x_5121;
wire x_5122;
wire x_5123;
wire x_5124;
wire x_5125;
wire x_5126;
wire x_5127;
wire x_5128;
wire x_5129;
wire x_5130;
wire x_5131;
wire x_5132;
wire x_5133;
wire x_5134;
wire x_5135;
wire x_5136;
wire x_5137;
wire x_5138;
wire x_5139;
wire x_5140;
wire x_5141;
wire x_5142;
wire x_5143;
wire x_5144;
wire x_5145;
wire x_5146;
wire x_5147;
wire x_5148;
wire x_5149;
wire x_5150;
wire x_5151;
wire x_5152;
wire x_5153;
wire x_5154;
wire x_5155;
wire x_5156;
wire x_5157;
wire x_5158;
wire x_5159;
wire x_5160;
wire x_5161;
wire x_5162;
wire x_5163;
wire x_5164;
wire x_5165;
wire x_5166;
wire x_5167;
wire x_5168;
wire x_5169;
wire x_5170;
wire x_5171;
wire x_5172;
wire x_5173;
wire x_5174;
wire x_5175;
wire x_5176;
wire x_5177;
wire x_5178;
wire x_5179;
wire x_5180;
wire x_5181;
wire x_5182;
wire x_5183;
wire x_5184;
wire x_5185;
wire x_5186;
wire x_5187;
wire x_5188;
wire x_5189;
wire x_5190;
wire x_5191;
wire x_5192;
wire x_5193;
wire x_5194;
wire x_5195;
wire x_5196;
wire x_5197;
wire x_5198;
wire x_5199;
wire x_5200;
wire x_5201;
wire x_5202;
wire x_5203;
wire x_5204;
wire x_5205;
wire x_5206;
wire x_5207;
wire x_5208;
wire x_5209;
wire x_5210;
wire x_5211;
wire x_5212;
wire x_5213;
wire x_5214;
wire x_5215;
wire x_5216;
wire x_5217;
wire x_5218;
wire x_5219;
wire x_5220;
wire x_5221;
wire x_5222;
wire x_5223;
wire x_5224;
wire x_5225;
wire x_5226;
wire x_5227;
wire x_5228;
wire x_5229;
wire x_5230;
wire x_5231;
wire x_5232;
wire x_5233;
wire x_5234;
wire x_5235;
wire x_5236;
wire x_5237;
wire x_5238;
wire x_5239;
wire x_5240;
wire x_5241;
wire x_5242;
wire x_5243;
wire x_5244;
wire x_5245;
wire x_5246;
wire x_5247;
wire x_5248;
wire x_5249;
wire x_5250;
wire x_5251;
wire x_5252;
wire x_5253;
wire x_5254;
wire x_5255;
wire x_5256;
wire x_5257;
wire x_5258;
wire x_5259;
wire x_5260;
wire x_5261;
wire x_5262;
wire x_5263;
wire x_5264;
wire x_5265;
wire x_5266;
wire x_5267;
wire x_5268;
wire x_5269;
wire x_5270;
wire x_5271;
wire x_5272;
wire x_5273;
wire x_5274;
wire x_5275;
wire x_5276;
wire x_5277;
wire x_5278;
wire x_5279;
wire x_5280;
wire x_5281;
wire x_5282;
wire x_5283;
wire x_5284;
wire x_5285;
wire x_5286;
wire x_5287;
wire x_5288;
wire x_5289;
wire x_5290;
wire x_5291;
wire x_5292;
wire x_5293;
wire x_5294;
wire x_5295;
wire x_5296;
wire x_5297;
wire x_5298;
wire x_5299;
wire x_5300;
wire x_5301;
wire x_5302;
wire x_5303;
wire x_5304;
wire x_5305;
wire x_5306;
wire x_5307;
wire x_5308;
wire x_5309;
wire x_5310;
wire x_5311;
wire x_5312;
wire x_5313;
wire x_5314;
wire x_5315;
wire x_5316;
wire x_5317;
wire x_5318;
wire x_5319;
wire x_5320;
wire x_5321;
wire x_5322;
wire x_5323;
wire x_5324;
wire x_5325;
wire x_5326;
wire x_5327;
wire x_5328;
wire x_5329;
wire x_5330;
wire x_5331;
wire x_5332;
wire x_5333;
wire x_5334;
wire x_5335;
wire x_5336;
wire x_5337;
wire x_5338;
wire x_5339;
wire x_5340;
wire x_5341;
wire x_5342;
wire x_5343;
wire x_5344;
wire x_5345;
wire x_5346;
wire x_5347;
wire x_5348;
wire x_5349;
wire x_5350;
wire x_5351;
wire x_5352;
wire x_5353;
wire x_5354;
wire x_5355;
wire x_5356;
wire x_5357;
wire x_5358;
wire x_5359;
wire x_5360;
wire x_5361;
wire x_5362;
wire x_5363;
wire x_5364;
wire x_5365;
wire x_5366;
wire x_5367;
wire x_5368;
wire x_5369;
wire x_5370;
wire x_5371;
wire x_5372;
wire x_5373;
wire x_5374;
wire x_5375;
wire x_5376;
wire x_5377;
wire x_5378;
wire x_5379;
wire x_5380;
wire x_5381;
wire x_5382;
wire x_5383;
wire x_5384;
wire x_5385;
wire x_5386;
wire x_5387;
wire x_5388;
wire x_5389;
wire x_5390;
wire x_5391;
wire x_5392;
wire x_5393;
wire x_5394;
wire x_5395;
wire x_5396;
wire x_5397;
wire x_5398;
wire x_5399;
wire x_5400;
wire x_5401;
wire x_5402;
wire x_5403;
wire x_5404;
wire x_5405;
wire x_5406;
wire x_5407;
wire x_5408;
wire x_5409;
wire x_5410;
wire x_5411;
wire x_5412;
wire x_5413;
wire x_5414;
wire x_5415;
wire x_5416;
wire x_5417;
wire x_5418;
wire x_5419;
wire x_5420;
wire x_5421;
wire x_5422;
wire x_5423;
wire x_5424;
wire x_5425;
wire x_5426;
wire x_5427;
wire x_5428;
wire x_5429;
wire x_5430;
wire x_5431;
wire x_5432;
wire x_5433;
wire x_5434;
wire x_5435;
wire x_5436;
wire x_5437;
wire x_5438;
wire x_5439;
wire x_5440;
wire x_5441;
wire x_5442;
wire x_5443;
wire x_5444;
wire x_5445;
wire x_5446;
wire x_5447;
wire x_5448;
wire x_5449;
wire x_5450;
wire x_5451;
wire x_5452;
wire x_5453;
wire x_5454;
wire x_5455;
wire x_5456;
wire x_5457;
wire x_5458;
wire x_5459;
wire x_5460;
wire x_5461;
wire x_5462;
wire x_5463;
wire x_5464;
wire x_5465;
wire x_5466;
wire x_5467;
wire x_5468;
wire x_5469;
wire x_5470;
wire x_5471;
wire x_5472;
wire x_5473;
wire x_5474;
wire x_5475;
wire x_5476;
wire x_5477;
wire x_5478;
wire x_5479;
wire x_5480;
wire x_5481;
wire x_5482;
wire x_5483;
wire x_5484;
wire x_5485;
wire x_5486;
wire x_5487;
wire x_5488;
wire x_5489;
wire x_5490;
wire x_5491;
wire x_5492;
wire x_5493;
wire x_5494;
wire x_5495;
wire x_5496;
wire x_5497;
wire x_5498;
wire x_5499;
wire x_5500;
wire x_5501;
wire x_5502;
wire x_5503;
wire x_5504;
wire x_5505;
wire x_5506;
wire x_5507;
wire x_5508;
wire x_5509;
wire x_5510;
wire x_5511;
wire x_5512;
wire x_5513;
wire x_5514;
wire x_5515;
wire x_5516;
wire x_5517;
wire x_5518;
wire x_5519;
wire x_5520;
wire x_5521;
wire x_5522;
wire x_5523;
wire x_5524;
wire x_5525;
wire x_5526;
wire x_5527;
wire x_5528;
wire x_5529;
wire x_5530;
wire x_5531;
wire x_5532;
wire x_5533;
wire x_5534;
wire x_5535;
wire x_5536;
wire x_5537;
wire x_5538;
wire x_5539;
wire x_5540;
wire x_5541;
wire x_5542;
wire x_5543;
wire x_5544;
wire x_5545;
wire x_5546;
wire x_5547;
wire x_5548;
wire x_5549;
wire x_5550;
wire x_5551;
wire x_5552;
wire x_5553;
wire x_5554;
wire x_5555;
wire x_5556;
wire x_5557;
wire x_5558;
wire x_5559;
wire x_5560;
wire x_5561;
wire x_5562;
wire x_5563;
wire x_5564;
wire x_5565;
wire x_5566;
wire x_5567;
wire x_5568;
wire x_5569;
wire x_5570;
wire x_5571;
wire x_5572;
wire x_5573;
wire x_5574;
wire x_5575;
wire x_5576;
wire x_5577;
wire x_5578;
wire x_5579;
wire x_5580;
wire x_5581;
wire x_5582;
wire x_5583;
wire x_5584;
wire x_5585;
wire x_5586;
wire x_5587;
wire x_5588;
wire x_5589;
wire x_5590;
wire x_5591;
wire x_5592;
wire x_5593;
wire x_5594;
wire x_5595;
wire x_5596;
wire x_5597;
wire x_5598;
wire x_5599;
wire x_5600;
wire x_5601;
wire x_5602;
wire x_5603;
wire x_5604;
wire x_5605;
wire x_5606;
wire x_5607;
wire x_5608;
wire x_5609;
wire x_5610;
wire x_5611;
wire x_5612;
wire x_5613;
wire x_5614;
wire x_5615;
wire x_5616;
wire x_5617;
wire x_5618;
wire x_5619;
wire x_5620;
wire x_5621;
wire x_5622;
wire x_5623;
wire x_5624;
wire x_5625;
wire x_5626;
wire x_5627;
wire x_5628;
wire x_5629;
wire x_5630;
wire x_5631;
wire x_5632;
wire x_5633;
wire x_5634;
wire x_5635;
wire x_5636;
wire x_5637;
wire x_5638;
wire x_5639;
wire x_5640;
wire x_5641;
wire x_5642;
wire x_5643;
wire x_5644;
wire x_5645;
wire x_5646;
wire x_5647;
wire x_5648;
wire x_5649;
wire x_5650;
wire x_5651;
wire x_5652;
wire x_5653;
wire x_5654;
wire x_5655;
wire x_5656;
wire x_5657;
wire x_5658;
wire x_5659;
wire x_5660;
wire x_5661;
wire x_5662;
wire x_5663;
wire x_5664;
wire x_5665;
wire x_5666;
wire x_5667;
wire x_5668;
wire x_5669;
wire x_5670;
wire x_5671;
wire x_5672;
wire x_5673;
wire x_5674;
wire x_5675;
wire x_5676;
wire x_5677;
wire x_5678;
wire x_5679;
wire x_5680;
wire x_5681;
wire x_5682;
wire x_5683;
wire x_5684;
wire x_5685;
wire x_5686;
wire x_5687;
wire x_5688;
wire x_5689;
wire x_5690;
wire x_5691;
wire x_5692;
wire x_5693;
wire x_5694;
wire x_5695;
wire x_5696;
wire x_5697;
wire x_5698;
wire x_5699;
wire x_5700;
wire x_5701;
wire x_5702;
wire x_5703;
wire x_5704;
wire x_5705;
wire x_5706;
wire x_5707;
wire x_5708;
wire x_5709;
wire x_5710;
wire x_5711;
wire x_5712;
wire x_5713;
wire x_5714;
wire x_5715;
wire x_5716;
wire x_5717;
wire x_5718;
wire x_5719;
wire x_5720;
wire x_5721;
wire x_5722;
wire x_5723;
wire x_5724;
wire x_5725;
wire x_5726;
wire x_5727;
wire x_5728;
wire x_5729;
wire x_5730;
wire x_5731;
wire x_5732;
wire x_5733;
wire x_5734;
wire x_5735;
wire x_5736;
wire x_5737;
wire x_5738;
wire x_5739;
wire x_5740;
wire x_5741;
wire x_5742;
wire x_5743;
wire x_5744;
wire x_5745;
wire x_5746;
wire x_5747;
wire x_5748;
wire x_5749;
wire x_5750;
wire x_5751;
wire x_5752;
wire x_5753;
wire x_5754;
wire x_5755;
wire x_5756;
wire x_5757;
wire x_5758;
wire x_5759;
wire x_5760;
wire x_5761;
wire x_5762;
wire x_5763;
wire x_5764;
wire x_5765;
wire x_5766;
wire x_5767;
wire x_5768;
wire x_5769;
wire x_5770;
wire x_5771;
wire x_5772;
wire x_5773;
wire x_5774;
wire x_5775;
wire x_5776;
wire x_5777;
wire x_5778;
wire x_5779;
wire x_5780;
wire x_5781;
wire x_5782;
wire x_5783;
wire x_5784;
wire x_5785;
wire x_5786;
wire x_5787;
wire x_5788;
wire x_5789;
wire x_5790;
wire x_5791;
wire x_5792;
wire x_5793;
wire x_5794;
wire x_5795;
wire x_5796;
wire x_5797;
wire x_5798;
wire x_5799;
wire x_5800;
wire x_5801;
wire x_5802;
wire x_5803;
wire x_5804;
wire x_5805;
wire x_5806;
wire x_5807;
wire x_5808;
wire x_5809;
wire x_5810;
wire x_5811;
wire x_5812;
wire x_5813;
wire x_5814;
wire x_5815;
wire x_5816;
wire x_5817;
wire x_5818;
wire x_5819;
wire x_5820;
wire x_5821;
wire x_5822;
wire x_5823;
wire x_5824;
wire x_5825;
wire x_5826;
wire x_5827;
wire x_5828;
wire x_5829;
wire x_5830;
wire x_5831;
wire x_5832;
wire x_5833;
wire x_5834;
wire x_5835;
wire x_5836;
wire x_5837;
wire x_5838;
wire x_5839;
wire x_5840;
wire x_5841;
wire x_5842;
wire x_5843;
wire x_5844;
wire x_5845;
wire x_5846;
wire x_5847;
wire x_5848;
wire x_5849;
wire x_5850;
wire x_5851;
wire x_5852;
wire x_5853;
wire x_5854;
wire x_5855;
wire x_5856;
wire x_5857;
wire x_5858;
wire x_5859;
wire x_5860;
wire x_5861;
wire x_5862;
wire x_5863;
wire x_5864;
wire x_5865;
wire x_5866;
wire x_5867;
wire x_5868;
wire x_5869;
wire x_5870;
wire x_5871;
wire x_5872;
wire x_5873;
wire x_5874;
wire x_5875;
wire x_5876;
wire x_5877;
wire x_5878;
wire x_5879;
wire x_5880;
wire x_5881;
wire x_5882;
wire x_5883;
wire x_5884;
wire x_5885;
wire x_5886;
wire x_5887;
wire x_5888;
wire x_5889;
wire x_5890;
wire x_5891;
wire x_5892;
wire x_5893;
wire x_5894;
wire x_5895;
wire x_5896;
wire x_5897;
wire x_5898;
wire x_5899;
wire x_5900;
wire x_5901;
wire x_5902;
wire x_5903;
wire x_5904;
wire x_5905;
wire x_5906;
wire x_5907;
wire x_5908;
wire x_5909;
wire x_5910;
wire x_5911;
wire x_5912;
wire x_5913;
wire x_5914;
wire x_5915;
wire x_5916;
wire x_5917;
wire x_5918;
wire x_5919;
wire x_5920;
wire x_5921;
wire x_5922;
wire x_5923;
wire x_5924;
wire x_5925;
wire x_5926;
wire x_5927;
wire x_5928;
wire x_5929;
wire x_5930;
wire x_5931;
wire x_5932;
wire x_5933;
wire x_5934;
wire x_5935;
wire x_5936;
wire x_5937;
wire x_5938;
wire x_5939;
wire x_5940;
wire x_5941;
wire x_5942;
wire x_5943;
wire x_5944;
wire x_5945;
wire x_5946;
wire x_5947;
wire x_5948;
wire x_5949;
wire x_5950;
wire x_5951;
wire x_5952;
wire x_5953;
wire x_5954;
wire x_5955;
wire x_5956;
wire x_5957;
wire x_5958;
wire x_5959;
wire x_5960;
wire x_5961;
wire x_5962;
wire x_5963;
wire x_5964;
wire x_5965;
wire x_5966;
wire x_5967;
wire x_5968;
wire x_5969;
wire x_5970;
wire x_5971;
wire x_5972;
wire x_5973;
wire x_5974;
wire x_5975;
wire x_5976;
wire x_5977;
wire x_5978;
wire x_5979;
wire x_5980;
wire x_5981;
wire x_5982;
wire x_5983;
wire x_5984;
wire x_5985;
wire x_5986;
wire x_5987;
wire x_5988;
wire x_5989;
wire x_5990;
wire x_5991;
wire x_5992;
wire x_5993;
wire x_5994;
wire x_5995;
wire x_5996;
wire x_5997;
wire x_5998;
wire x_5999;
wire x_6000;
wire x_6001;
wire x_6002;
wire x_6003;
wire x_6004;
wire x_6005;
wire x_6006;
wire x_6007;
wire x_6008;
wire x_6009;
wire x_6010;
wire x_6011;
wire x_6012;
wire x_6013;
wire x_6014;
wire x_6015;
wire x_6016;
wire x_6017;
wire x_6018;
wire x_6019;
wire x_6020;
wire x_6021;
wire x_6022;
wire x_6023;
wire x_6024;
wire x_6025;
wire x_6026;
wire x_6027;
wire x_6028;
wire x_6029;
wire x_6030;
wire x_6031;
wire x_6032;
wire x_6033;
wire x_6034;
wire x_6035;
wire x_6036;
wire x_6037;
wire x_6038;
wire x_6039;
wire x_6040;
wire x_6041;
wire x_6042;
wire x_6043;
wire x_6044;
wire x_6045;
wire x_6046;
wire x_6047;
wire x_6048;
wire x_6049;
wire x_6050;
wire x_6051;
wire x_6052;
wire x_6053;
wire x_6054;
wire x_6055;
wire x_6056;
wire x_6057;
wire x_6058;
wire x_6059;
wire x_6060;
wire x_6061;
wire x_6062;
wire x_6063;
wire x_6064;
wire x_6065;
wire x_6066;
wire x_6067;
wire x_6068;
wire x_6069;
wire x_6070;
wire x_6071;
wire x_6072;
wire x_6073;
wire x_6074;
wire x_6075;
wire x_6076;
wire x_6077;
wire x_6078;
wire x_6079;
wire x_6080;
wire x_6081;
wire x_6082;
wire x_6083;
wire x_6084;
wire x_6085;
wire x_6086;
wire x_6087;
wire x_6088;
wire x_6089;
wire x_6090;
wire x_6091;
wire x_6092;
wire x_6093;
wire x_6094;
wire x_6095;
wire x_6096;
wire x_6097;
wire x_6098;
wire x_6099;
wire x_6100;
wire x_6101;
wire x_6102;
wire x_6103;
wire x_6104;
wire x_6105;
wire x_6106;
wire x_6107;
wire x_6108;
wire x_6109;
wire x_6110;
wire x_6111;
wire x_6112;
wire x_6113;
wire x_6114;
wire x_6115;
wire x_6116;
wire x_6117;
wire x_6118;
wire x_6119;
wire x_6120;
wire x_6121;
wire x_6122;
wire x_6123;
wire x_6124;
wire x_6125;
wire x_6126;
wire x_6127;
wire x_6128;
wire x_6129;
wire x_6130;
wire x_6131;
wire x_6132;
wire x_6133;
wire x_6134;
wire x_6135;
wire x_6136;
wire x_6137;
wire x_6138;
wire x_6139;
wire x_6140;
wire x_6141;
wire x_6142;
wire x_6143;
wire x_6144;
wire x_6145;
wire x_6146;
wire x_6147;
wire x_6148;
wire x_6149;
wire x_6150;
wire x_6151;
wire x_6152;
wire x_6153;
wire x_6154;
wire x_6155;
wire x_6156;
wire x_6157;
wire x_6158;
wire x_6159;
wire x_6160;
wire x_6161;
wire x_6162;
wire x_6163;
wire x_6164;
wire x_6165;
wire x_6166;
wire x_6167;
wire x_6168;
wire x_6169;
wire x_6170;
wire x_6171;
wire x_6172;
wire x_6173;
wire x_6174;
wire x_6175;
wire x_6176;
wire x_6177;
wire x_6178;
wire x_6179;
wire x_6180;
wire x_6181;
wire x_6182;
wire x_6183;
wire x_6184;
wire x_6185;
wire x_6186;
wire x_6187;
wire x_6188;
wire x_6189;
wire x_6190;
wire x_6191;
wire x_6192;
wire x_6193;
wire x_6194;
wire x_6195;
wire x_6196;
wire x_6197;
wire x_6198;
wire x_6199;
wire x_6200;
wire x_6201;
wire x_6202;
wire x_6203;
wire x_6204;
wire x_6205;
wire x_6206;
wire x_6207;
wire x_6208;
wire x_6209;
wire x_6210;
wire x_6211;
wire x_6212;
wire x_6213;
wire x_6214;
wire x_6215;
wire x_6216;
wire x_6217;
wire x_6218;
wire x_6219;
wire x_6220;
wire x_6221;
wire x_6222;
wire x_6223;
wire x_6224;
wire x_6225;
wire x_6226;
wire x_6227;
wire x_6228;
wire x_6229;
wire x_6230;
wire x_6231;
wire x_6232;
wire x_6233;
wire x_6234;
wire x_6235;
wire x_6236;
wire x_6237;
wire x_6238;
wire x_6239;
wire x_6240;
wire x_6241;
wire x_6242;
wire x_6243;
wire x_6244;
wire x_6245;
wire x_6246;
wire x_6247;
wire x_6248;
wire x_6249;
wire x_6250;
wire x_6251;
wire x_6252;
wire x_6253;
wire x_6254;
wire x_6255;
wire x_6256;
wire x_6257;
wire x_6258;
wire x_6259;
wire x_6260;
wire x_6261;
wire x_6262;
wire x_6263;
wire x_6264;
wire x_6265;
wire x_6266;
wire x_6267;
wire x_6268;
wire x_6269;
wire x_6270;
wire x_6271;
wire x_6272;
wire x_6273;
wire x_6274;
wire x_6275;
wire x_6276;
wire x_6277;
wire x_6278;
wire x_6279;
wire x_6280;
wire x_6281;
wire x_6282;
wire x_6283;
wire x_6284;
wire x_6285;
wire x_6286;
wire x_6287;
wire x_6288;
wire x_6289;
wire x_6290;
wire x_6291;
wire x_6292;
wire x_6293;
wire x_6294;
wire x_6295;
wire x_6296;
wire x_6297;
wire x_6298;
wire x_6299;
wire x_6300;
wire x_6301;
wire x_6302;
wire x_6303;
wire x_6304;
wire x_6305;
wire x_6306;
wire x_6307;
wire x_6308;
wire x_6309;
wire x_6310;
wire x_6311;
wire x_6312;
wire x_6313;
wire x_6314;
wire x_6315;
wire x_6316;
wire x_6317;
wire x_6318;
wire x_6319;
wire x_6320;
wire x_6321;
wire x_6322;
wire x_6323;
wire x_6324;
wire x_6325;
wire x_6326;
wire x_6327;
wire x_6328;
wire x_6329;
wire x_6330;
wire x_6331;
wire x_6332;
wire x_6333;
wire x_6334;
wire x_6335;
wire x_6336;
wire x_6337;
wire x_6338;
wire x_6339;
wire x_6340;
wire x_6341;
wire x_6342;
wire x_6343;
wire x_6344;
wire x_6345;
wire x_6346;
wire x_6347;
wire x_6348;
wire x_6349;
wire x_6350;
wire x_6351;
wire x_6352;
wire x_6353;
wire x_6354;
wire x_6355;
wire x_6356;
wire x_6357;
wire x_6358;
wire x_6359;
wire x_6360;
wire x_6361;
wire x_6362;
wire x_6363;
wire x_6364;
wire x_6365;
wire x_6366;
wire x_6367;
wire x_6368;
wire x_6369;
wire x_6370;
wire x_6371;
wire x_6372;
wire x_6373;
wire x_6374;
wire x_6375;
wire x_6376;
wire x_6377;
wire x_6378;
wire x_6379;
wire x_6380;
wire x_6381;
wire x_6382;
wire x_6383;
wire x_6384;
wire x_6385;
wire x_6386;
wire x_6387;
wire x_6388;
wire x_6389;
wire x_6390;
wire x_6391;
wire x_6392;
wire x_6393;
wire x_6394;
wire x_6395;
wire x_6396;
wire x_6397;
wire x_6398;
wire x_6399;
wire x_6400;
wire x_6401;
wire x_6402;
wire x_6403;
wire x_6404;
wire x_6405;
wire x_6406;
wire x_6407;
wire x_6408;
wire x_6409;
wire x_6410;
wire x_6411;
wire x_6412;
wire x_6413;
wire x_6414;
wire x_6415;
wire x_6416;
wire x_6417;
wire x_6418;
wire x_6419;
wire x_6420;
wire x_6421;
wire x_6422;
wire x_6423;
wire x_6424;
wire x_6425;
wire x_6426;
wire x_6427;
wire x_6428;
wire x_6429;
wire x_6430;
wire x_6431;
wire x_6432;
wire x_6433;
wire x_6434;
wire x_6435;
wire x_6436;
wire x_6437;
wire x_6438;
wire x_6439;
wire x_6440;
wire x_6441;
wire x_6442;
wire x_6443;
wire x_6444;
wire x_6445;
wire x_6446;
wire x_6447;
wire x_6448;
wire x_6449;
wire x_6450;
wire x_6451;
wire x_6452;
wire x_6453;
wire x_6454;
wire x_6455;
wire x_6456;
wire x_6457;
wire x_6458;
wire x_6459;
wire x_6460;
wire x_6461;
wire x_6462;
wire x_6463;
wire x_6464;
wire x_6465;
wire x_6466;
wire x_6467;
wire x_6468;
wire x_6469;
wire x_6470;
wire x_6471;
wire x_6472;
wire x_6473;
wire x_6474;
wire x_6475;
wire x_6476;
wire x_6477;
wire x_6478;
wire x_6479;
wire x_6480;
wire x_6481;
wire x_6482;
wire x_6483;
wire x_6484;
wire x_6485;
wire x_6486;
wire x_6487;
wire x_6488;
wire x_6489;
wire x_6490;
wire x_6491;
wire x_6492;
wire x_6493;
wire x_6494;
wire x_6495;
wire x_6496;
wire x_6497;
wire x_6498;
wire x_6499;
wire x_6500;
wire x_6501;
wire x_6502;
wire x_6503;
wire x_6504;
wire x_6505;
wire x_6506;
wire x_6507;
wire x_6508;
wire x_6509;
wire x_6510;
wire x_6511;
wire x_6512;
wire x_6513;
wire x_6514;
wire x_6515;
wire x_6516;
wire x_6517;
wire x_6518;
wire x_6519;
wire x_6520;
wire x_6521;
wire x_6522;
wire x_6523;
wire x_6524;
wire x_6525;
wire x_6526;
wire x_6527;
wire x_6528;
wire x_6529;
wire x_6530;
wire x_6531;
wire x_6532;
wire x_6533;
wire x_6534;
wire x_6535;
wire x_6536;
wire x_6537;
wire x_6538;
wire x_6539;
wire x_6540;
wire x_6541;
wire x_6542;
wire x_6543;
wire x_6544;
wire x_6545;
wire x_6546;
wire x_6547;
wire x_6548;
wire x_6549;
wire x_6550;
wire x_6551;
wire x_6552;
wire x_6553;
wire x_6554;
wire x_6555;
wire x_6556;
wire x_6557;
wire x_6558;
wire x_6559;
wire x_6560;
wire x_6561;
wire x_6562;
wire x_6563;
wire x_6564;
wire x_6565;
wire x_6566;
wire x_6567;
wire x_6568;
wire x_6569;
wire x_6570;
wire x_6571;
wire x_6572;
wire x_6573;
wire x_6574;
wire x_6575;
wire x_6576;
wire x_6577;
wire x_6578;
wire x_6579;
wire x_6580;
wire x_6581;
wire x_6582;
wire x_6583;
wire x_6584;
wire x_6585;
wire x_6586;
wire x_6587;
wire x_6588;
wire x_6589;
wire x_6590;
wire x_6591;
wire x_6592;
wire x_6593;
wire x_6594;
wire x_6595;
wire x_6596;
wire x_6597;
wire x_6598;
wire x_6599;
wire x_6600;
wire x_6601;
wire x_6602;
wire x_6603;
wire x_6604;
wire x_6605;
wire x_6606;
wire x_6607;
wire x_6608;
wire x_6609;
wire x_6610;
wire x_6611;
wire x_6612;
wire x_6613;
wire x_6614;
wire x_6615;
wire x_6616;
wire x_6617;
wire x_6618;
wire x_6619;
wire x_6620;
wire x_6621;
wire x_6622;
wire x_6623;
wire x_6624;
wire x_6625;
wire x_6626;
wire x_6627;
wire x_6628;
wire x_6629;
wire x_6630;
wire x_6631;
wire x_6632;
wire x_6633;
wire x_6634;
wire x_6635;
wire x_6636;
wire x_6637;
wire x_6638;
wire x_6639;
wire x_6640;
wire x_6641;
wire x_6642;
wire x_6643;
wire x_6644;
wire x_6645;
wire x_6646;
wire x_6647;
wire x_6648;
wire x_6649;
wire x_6650;
wire x_6651;
wire x_6652;
wire x_6653;
wire x_6654;
wire x_6655;
wire x_6656;
wire x_6657;
wire x_6658;
wire x_6659;
wire x_6660;
wire x_6661;
wire x_6662;
wire x_6663;
wire x_6664;
wire x_6665;
wire x_6666;
wire x_6667;
wire x_6668;
wire x_6669;
wire x_6670;
wire x_6671;
wire x_6672;
wire x_6673;
wire x_6674;
wire x_6675;
wire x_6676;
wire x_6677;
wire x_6678;
wire x_6679;
wire x_6680;
wire x_6681;
wire x_6682;
wire x_6683;
wire x_6684;
wire x_6685;
wire x_6686;
wire x_6687;
wire x_6688;
wire x_6689;
wire x_6690;
wire x_6691;
wire x_6692;
wire x_6693;
wire x_6694;
wire x_6695;
wire x_6696;
wire x_6697;
wire x_6698;
wire x_6699;
wire x_6700;
wire x_6701;
wire x_6702;
wire x_6703;
wire x_6704;
wire x_6705;
wire x_6706;
wire x_6707;
wire x_6708;
wire x_6709;
wire x_6710;
wire x_6711;
wire x_6712;
wire x_6713;
wire x_6714;
wire x_6715;
wire x_6716;
wire x_6717;
wire x_6718;
wire x_6719;
wire x_6720;
wire x_6721;
wire x_6722;
wire x_6723;
wire x_6724;
wire x_6725;
wire x_6726;
wire x_6727;
wire x_6728;
wire x_6729;
wire x_6730;
wire x_6731;
wire x_6732;
wire x_6733;
wire x_6734;
wire x_6735;
wire x_6736;
wire x_6737;
wire x_6738;
wire x_6739;
wire x_6740;
wire x_6741;
wire x_6742;
wire x_6743;
wire x_6744;
wire x_6745;
wire x_6746;
wire x_6747;
wire x_6748;
wire x_6749;
wire x_6750;
wire x_6751;
wire x_6752;
wire x_6753;
wire x_6754;
wire x_6755;
wire x_6756;
wire x_6757;
wire x_6758;
wire x_6759;
wire x_6760;
wire x_6761;
wire x_6762;
wire x_6763;
wire x_6764;
wire x_6765;
wire x_6766;
wire x_6767;
wire x_6768;
wire x_6769;
wire x_6770;
wire x_6771;
wire x_6772;
wire x_6773;
wire x_6774;
wire x_6775;
wire x_6776;
wire x_6777;
wire x_6778;
wire x_6779;
wire x_6780;
wire x_6781;
wire x_6782;
wire x_6783;
wire x_6784;
wire x_6785;
wire x_6786;
wire x_6787;
wire x_6788;
wire x_6789;
wire x_6790;
wire x_6791;
wire x_6792;
wire x_6793;
wire x_6794;
wire x_6795;
wire x_6796;
wire x_6797;
wire x_6798;
wire x_6799;
wire x_6800;
wire x_6801;
wire x_6802;
wire x_6803;
wire x_6804;
wire x_6805;
wire x_6806;
wire x_6807;
wire x_6808;
wire x_6809;
wire x_6810;
wire x_6811;
wire x_6812;
wire x_6813;
wire x_6814;
wire x_6815;
wire x_6816;
wire x_6817;
wire x_6818;
wire x_6819;
wire x_6820;
wire x_6821;
wire x_6822;
wire x_6823;
wire x_6824;
wire x_6825;
wire x_6826;
wire x_6827;
wire x_6828;
wire x_6829;
wire x_6830;
wire x_6831;
wire x_6832;
wire x_6833;
wire x_6834;
wire x_6835;
wire x_6836;
wire x_6837;
wire x_6838;
wire x_6839;
wire x_6840;
wire x_6841;
wire x_6842;
wire x_6843;
wire x_6844;
wire x_6845;
wire x_6846;
wire x_6847;
wire x_6848;
wire x_6849;
wire x_6850;
wire x_6851;
wire x_6852;
wire x_6853;
wire x_6854;
wire x_6855;
wire x_6856;
wire x_6857;
wire x_6858;
wire x_6859;
wire x_6860;
wire x_6861;
wire x_6862;
wire x_6863;
wire x_6864;
wire x_6865;
wire x_6866;
wire x_6867;
wire x_6868;
wire x_6869;
wire x_6870;
wire x_6871;
wire x_6872;
wire x_6873;
wire x_6874;
wire x_6875;
wire x_6876;
wire x_6877;
wire x_6878;
wire x_6879;
wire x_6880;
wire x_6881;
wire x_6882;
wire x_6883;
wire x_6884;
wire x_6885;
wire x_6886;
wire x_6887;
wire x_6888;
wire x_6889;
wire x_6890;
wire x_6891;
wire x_6892;
wire x_6893;
wire x_6894;
wire x_6895;
wire x_6896;
wire x_6897;
wire x_6898;
wire x_6899;
wire x_6900;
wire x_6901;
wire x_6902;
wire x_6903;
wire x_6904;
wire x_6905;
wire x_6906;
wire x_6907;
wire x_6908;
wire x_6909;
wire x_6910;
wire x_6911;
wire x_6912;
wire x_6913;
wire x_6914;
wire x_6915;
wire x_6916;
wire x_6917;
wire x_6918;
wire x_6919;
wire x_6920;
wire x_6921;
wire x_6922;
wire x_6923;
wire x_6924;
wire x_6925;
wire x_6926;
wire x_6927;
wire x_6928;
wire x_6929;
wire x_6930;
wire x_6931;
wire x_6932;
wire x_6933;
wire x_6934;
wire x_6935;
wire x_6936;
wire x_6937;
wire x_6938;
wire x_6939;
wire x_6940;
wire x_6941;
wire x_6942;
wire x_6943;
wire x_6944;
wire x_6945;
wire x_6946;
wire x_6947;
wire x_6948;
wire x_6949;
wire x_6950;
wire x_6951;
wire x_6952;
wire x_6953;
wire x_6954;
wire x_6955;
wire x_6956;
wire x_6957;
wire x_6958;
wire x_6959;
wire x_6960;
wire x_6961;
wire x_6962;
wire x_6963;
wire x_6964;
wire x_6965;
wire x_6966;
wire x_6967;
wire x_6968;
wire x_6969;
wire x_6970;
wire x_6971;
wire x_6972;
wire x_6973;
wire x_6974;
wire x_6975;
wire x_6976;
wire x_6977;
wire x_6978;
wire x_6979;
wire x_6980;
wire x_6981;
wire x_6982;
wire x_6983;
wire x_6984;
wire x_6985;
wire x_6986;
wire x_6987;
wire x_6988;
wire x_6989;
wire x_6990;
wire x_6991;
wire x_6992;
wire x_6993;
wire x_6994;
wire x_6995;
wire x_6996;
wire x_6997;
wire x_6998;
wire x_6999;
wire x_7000;
wire x_7001;
wire x_7002;
wire x_7003;
wire x_7004;
wire x_7005;
wire x_7006;
wire x_7007;
wire x_7008;
wire x_7009;
wire x_7010;
wire x_7011;
wire x_7012;
wire x_7013;
wire x_7014;
wire x_7015;
wire x_7016;
wire x_7017;
wire x_7018;
wire x_7019;
wire x_7020;
wire x_7021;
wire x_7022;
wire x_7023;
wire x_7024;
wire x_7025;
wire x_7026;
wire x_7027;
wire x_7028;
wire x_7029;
wire x_7030;
wire x_7031;
wire x_7032;
wire x_7033;
wire x_7034;
wire x_7035;
wire x_7036;
wire x_7037;
wire x_7038;
wire x_7039;
wire x_7040;
wire x_7041;
wire x_7042;
wire x_7043;
wire x_7044;
wire x_7045;
wire x_7046;
wire x_7047;
wire x_7048;
wire x_7049;
wire x_7050;
wire x_7051;
wire x_7052;
wire x_7053;
wire x_7054;
wire x_7055;
wire x_7056;
wire x_7057;
wire x_7058;
wire x_7059;
wire x_7060;
wire x_7061;
wire x_7062;
wire x_7063;
wire x_7064;
wire x_7065;
wire x_7066;
wire x_7067;
wire x_7068;
wire x_7069;
wire x_7070;
wire x_7071;
wire x_7072;
wire x_7073;
wire x_7074;
wire x_7075;
wire x_7076;
wire x_7077;
wire x_7078;
wire x_7079;
wire x_7080;
wire x_7081;
wire x_7082;
wire x_7083;
wire x_7084;
wire x_7085;
wire x_7086;
wire x_7087;
wire x_7088;
wire x_7089;
wire x_7090;
wire x_7091;
wire x_7092;
wire x_7093;
wire x_7094;
wire x_7095;
wire x_7096;
wire x_7097;
wire x_7098;
wire x_7099;
wire x_7100;
wire x_7101;
wire x_7102;
wire x_7103;
wire x_7104;
wire x_7105;
wire x_7106;
wire x_7107;
wire x_7108;
wire x_7109;
wire x_7110;
wire x_7111;
wire x_7112;
wire x_7113;
wire x_7114;
wire x_7115;
wire x_7116;
wire x_7117;
wire x_7118;
wire x_7119;
wire x_7120;
wire x_7121;
wire x_7122;
wire x_7123;
wire x_7124;
wire x_7125;
wire x_7126;
wire x_7127;
wire x_7128;
wire x_7129;
wire x_7130;
wire x_7131;
wire x_7132;
wire x_7133;
wire x_7134;
wire x_7135;
wire x_7136;
wire x_7137;
wire x_7138;
wire x_7139;
wire x_7140;
wire x_7141;
wire x_7142;
wire x_7143;
wire x_7144;
wire x_7145;
wire x_7146;
wire x_7147;
wire x_7148;
wire x_7149;
wire x_7150;
wire x_7151;
wire x_7152;
wire x_7153;
wire x_7154;
wire x_7155;
wire x_7156;
wire x_7157;
wire x_7158;
wire x_7159;
wire x_7160;
wire x_7161;
wire x_7162;
wire x_7163;
wire x_7164;
wire x_7165;
wire x_7166;
wire x_7167;
wire x_7168;
wire x_7169;
wire x_7170;
wire x_7171;
wire x_7172;
wire x_7173;
wire x_7174;
wire x_7175;
wire x_7176;
wire x_7177;
wire x_7178;
wire x_7179;
wire x_7180;
wire x_7181;
wire x_7182;
wire x_7183;
wire x_7184;
wire x_7185;
wire x_7186;
wire x_7187;
wire x_7188;
wire x_7189;
wire x_7190;
wire x_7191;
wire x_7192;
wire x_7193;
wire x_7194;
wire x_7195;
wire x_7196;
wire x_7197;
wire x_7198;
wire x_7199;
wire x_7200;
wire x_7201;
wire x_7202;
wire x_7203;
wire x_7204;
wire x_7205;
wire x_7206;
wire x_7207;
wire x_7208;
wire x_7209;
wire x_7210;
wire x_7211;
wire x_7212;
wire x_7213;
wire x_7214;
wire x_7215;
wire x_7216;
wire x_7217;
wire x_7218;
wire x_7219;
wire x_7220;
wire x_7221;
wire x_7222;
wire x_7223;
wire x_7224;
wire x_7225;
wire x_7226;
wire x_7227;
wire x_7228;
wire x_7229;
wire x_7230;
wire x_7231;
wire x_7232;
wire x_7233;
wire x_7234;
wire x_7235;
wire x_7236;
wire x_7237;
wire x_7238;
wire x_7239;
wire x_7240;
wire x_7241;
wire x_7242;
wire x_7243;
wire x_7244;
wire x_7245;
wire x_7246;
wire x_7247;
wire x_7248;
wire x_7249;
wire x_7250;
wire x_7251;
wire x_7252;
wire x_7253;
wire x_7254;
wire x_7255;
wire x_7256;
wire x_7257;
wire x_7258;
wire x_7259;
wire x_7260;
wire x_7261;
wire x_7262;
wire x_7263;
wire x_7264;
wire x_7265;
wire x_7266;
wire x_7267;
wire x_7268;
wire x_7269;
wire x_7270;
wire x_7271;
wire x_7272;
wire x_7273;
wire x_7274;
wire x_7275;
wire x_7276;
wire x_7277;
wire x_7278;
wire x_7279;
wire x_7280;
wire x_7281;
wire x_7282;
wire x_7283;
wire x_7284;
wire x_7285;
wire x_7286;
wire x_7287;
wire x_7288;
wire x_7289;
wire x_7290;
wire x_7291;
wire x_7292;
wire x_7293;
wire x_7294;
wire x_7295;
wire x_7296;
wire x_7297;
wire x_7298;
wire x_7299;
wire x_7300;
wire x_7301;
wire x_7302;
wire x_7303;
wire x_7304;
wire x_7305;
wire x_7306;
wire x_7307;
wire x_7308;
wire x_7309;
wire x_7310;
wire x_7311;
wire x_7312;
wire x_7313;
wire x_7314;
wire x_7315;
wire x_7316;
wire x_7317;
wire x_7318;
wire x_7319;
wire x_7320;
wire x_7321;
wire x_7322;
wire x_7323;
wire x_7324;
wire x_7325;
wire x_7326;
wire x_7327;
wire x_7328;
wire x_7329;
wire x_7330;
wire x_7331;
wire x_7332;
wire x_7333;
wire x_7334;
wire x_7335;
wire x_7336;
wire x_7337;
wire x_7338;
wire x_7339;
wire x_7340;
wire x_7341;
wire x_7342;
wire x_7343;
wire x_7344;
wire x_7345;
wire x_7346;
wire x_7347;
wire x_7348;
wire x_7349;
wire x_7350;
wire x_7351;
wire x_7352;
wire x_7353;
wire x_7354;
wire x_7355;
wire x_7356;
wire x_7357;
wire x_7358;
wire x_7359;
wire x_7360;
wire x_7361;
wire x_7362;
wire x_7363;
wire x_7364;
wire x_7365;
wire x_7366;
wire x_7367;
wire x_7368;
wire x_7369;
wire x_7370;
wire x_7371;
wire x_7372;
wire x_7373;
wire x_7374;
wire x_7375;
wire x_7376;
wire x_7377;
wire x_7378;
wire x_7379;
wire x_7380;
wire x_7381;
wire x_7382;
wire x_7383;
wire x_7384;
wire x_7385;
wire x_7386;
wire x_7387;
wire x_7388;
wire x_7389;
wire x_7390;
wire x_7391;
wire x_7392;
wire x_7393;
wire x_7394;
wire x_7395;
wire x_7396;
wire x_7397;
wire x_7398;
wire x_7399;
wire x_7400;
wire x_7401;
wire x_7402;
wire x_7403;
wire x_7404;
wire x_7405;
wire x_7406;
wire x_7407;
wire x_7408;
wire x_7409;
wire x_7410;
wire x_7411;
wire x_7412;
wire x_7413;
wire x_7414;
wire x_7415;
wire x_7416;
wire x_7417;
wire x_7418;
wire x_7419;
wire x_7420;
wire x_7421;
wire x_7422;
wire x_7423;
wire x_7424;
wire x_7425;
wire x_7426;
wire x_7427;
wire x_7428;
wire x_7429;
wire x_7430;
wire x_7431;
wire x_7432;
wire x_7433;
wire x_7434;
wire x_7435;
wire x_7436;
wire x_7437;
wire x_7438;
wire x_7439;
wire x_7440;
wire x_7441;
wire x_7442;
wire x_7443;
wire x_7444;
wire x_7445;
wire x_7446;
wire x_7447;
wire x_7448;
wire x_7449;
wire x_7450;
wire x_7451;
wire x_7452;
wire x_7453;
wire x_7454;
wire x_7455;
wire x_7456;
wire x_7457;
wire x_7458;
wire x_7459;
wire x_7460;
wire x_7461;
wire x_7462;
wire x_7463;
wire x_7464;
wire x_7465;
wire x_7466;
wire x_7467;
wire x_7468;
wire x_7469;
wire x_7470;
wire x_7471;
wire x_7472;
wire x_7473;
wire x_7474;
wire x_7475;
wire x_7476;
wire x_7477;
wire x_7478;
wire x_7479;
wire x_7480;
wire x_7481;
wire x_7482;
wire x_7483;
wire x_7484;
wire x_7485;
wire x_7486;
wire x_7487;
wire x_7488;
wire x_7489;
wire x_7490;
wire x_7491;
wire x_7492;
wire x_7493;
wire x_7494;
wire x_7495;
wire x_7496;
wire x_7497;
wire x_7498;
wire x_7499;
wire x_7500;
wire x_7501;
wire x_7502;
wire x_7503;
wire x_7504;
wire x_7505;
wire x_7506;
wire x_7507;
wire x_7508;
wire x_7509;
wire x_7510;
wire x_7511;
wire x_7512;
wire x_7513;
wire x_7514;
wire x_7515;
wire x_7516;
wire x_7517;
wire x_7518;
wire x_7519;
wire x_7520;
wire x_7521;
wire x_7522;
wire x_7523;
wire x_7524;
wire x_7525;
wire x_7526;
wire x_7527;
wire x_7528;
wire x_7529;
wire x_7530;
wire x_7531;
wire x_7532;
wire x_7533;
wire x_7534;
wire x_7535;
wire x_7536;
wire x_7537;
wire x_7538;
wire x_7539;
wire x_7540;
wire x_7541;
wire x_7542;
wire x_7543;
wire x_7544;
wire x_7545;
wire x_7546;
wire x_7547;
wire x_7548;
wire x_7549;
wire x_7550;
wire x_7551;
wire x_7552;
wire x_7553;
wire x_7554;
wire x_7555;
wire x_7556;
wire x_7557;
wire x_7558;
wire x_7559;
wire x_7560;
wire x_7561;
wire x_7562;
wire x_7563;
wire x_7564;
wire x_7565;
wire x_7566;
wire x_7567;
wire x_7568;
wire x_7569;
wire x_7570;
wire x_7571;
wire x_7572;
wire x_7573;
wire x_7574;
wire x_7575;
wire x_7576;
wire x_7577;
wire x_7578;
wire x_7579;
wire x_7580;
wire x_7581;
wire x_7582;
wire x_7583;
wire x_7584;
wire x_7585;
wire x_7586;
wire x_7587;
wire x_7588;
wire x_7589;
wire x_7590;
wire x_7591;
wire x_7592;
wire x_7593;
wire x_7594;
wire x_7595;
wire x_7596;
wire x_7597;
wire x_7598;
wire x_7599;
wire x_7600;
wire x_7601;
wire x_7602;
wire x_7603;
wire x_7604;
wire x_7605;
wire x_7606;
wire x_7607;
wire x_7608;
wire x_7609;
wire x_7610;
wire x_7611;
wire x_7612;
wire x_7613;
wire x_7614;
wire x_7615;
wire x_7616;
wire x_7617;
wire x_7618;
wire x_7619;
wire x_7620;
wire x_7621;
wire x_7622;
wire x_7623;
wire x_7624;
wire x_7625;
wire x_7626;
wire x_7627;
wire x_7628;
wire x_7629;
wire x_7630;
wire x_7631;
wire x_7632;
wire x_7633;
wire x_7634;
wire x_7635;
wire x_7636;
wire x_7637;
wire x_7638;
wire x_7639;
wire x_7640;
wire x_7641;
wire x_7642;
wire x_7643;
wire x_7644;
wire x_7645;
wire x_7646;
wire x_7647;
wire x_7648;
wire x_7649;
wire x_7650;
wire x_7651;
wire x_7652;
wire x_7653;
wire x_7654;
wire x_7655;
wire x_7656;
wire x_7657;
wire x_7658;
wire x_7659;
wire x_7660;
wire x_7661;
wire x_7662;
wire x_7663;
wire x_7664;
wire x_7665;
wire x_7666;
wire x_7667;
wire x_7668;
wire x_7669;
wire x_7670;
wire x_7671;
wire x_7672;
wire x_7673;
wire x_7674;
wire x_7675;
wire x_7676;
wire x_7677;
wire x_7678;
wire x_7679;
wire x_7680;
wire x_7681;
wire x_7682;
wire x_7683;
wire x_7684;
wire x_7685;
wire x_7686;
wire x_7687;
wire x_7688;
wire x_7689;
wire x_7690;
wire x_7691;
wire x_7692;
wire x_7693;
wire x_7694;
wire x_7695;
wire x_7696;
wire x_7697;
wire x_7698;
wire x_7699;
wire x_7700;
wire x_7701;
wire x_7702;
wire x_7703;
wire x_7704;
wire x_7705;
wire x_7706;
wire x_7707;
wire x_7708;
wire x_7709;
wire x_7710;
wire x_7711;
wire x_7712;
wire x_7713;
wire x_7714;
wire x_7715;
wire x_7716;
wire x_7717;
wire x_7718;
wire x_7719;
wire x_7720;
wire x_7721;
wire x_7722;
wire x_7723;
wire x_7724;
wire x_7725;
wire x_7726;
wire x_7727;
wire x_7728;
wire x_7729;
wire x_7730;
wire x_7731;
wire x_7732;
wire x_7733;
wire x_7734;
wire x_7735;
wire x_7736;
wire x_7737;
wire x_7738;
wire x_7739;
wire x_7740;
wire x_7741;
wire x_7742;
wire x_7743;
wire x_7744;
wire x_7745;
wire x_7746;
wire x_7747;
wire x_7748;
wire x_7749;
wire x_7750;
wire x_7751;
wire x_7752;
wire x_7753;
wire x_7754;
wire x_7755;
wire x_7756;
wire x_7757;
wire x_7758;
wire x_7759;
wire x_7760;
wire x_7761;
wire x_7762;
wire x_7763;
wire x_7764;
wire x_7765;
wire x_7766;
wire x_7767;
wire x_7768;
wire x_7769;
wire x_7770;
wire x_7771;
wire x_7772;
wire x_7773;
wire x_7774;
wire x_7775;
wire x_7776;
wire x_7777;
wire x_7778;
wire x_7779;
wire x_7780;
wire x_7781;
wire x_7782;
wire x_7783;
wire x_7784;
wire x_7785;
wire x_7786;
wire x_7787;
wire x_7788;
wire x_7789;
wire x_7790;
wire x_7791;
wire x_7792;
wire x_7793;
wire x_7794;
wire x_7795;
wire x_7796;
wire x_7797;
wire x_7798;
wire x_7799;
wire x_7800;
wire x_7801;
wire x_7802;
wire x_7803;
wire x_7804;
wire x_7805;
wire x_7806;
wire x_7807;
wire x_7808;
wire x_7809;
wire x_7810;
wire x_7811;
wire x_7812;
wire x_7813;
wire x_7814;
wire x_7815;
wire x_7816;
wire x_7817;
wire x_7818;
wire x_7819;
wire x_7820;
wire x_7821;
wire x_7822;
wire x_7823;
wire x_7824;
wire x_7825;
wire x_7826;
wire x_7827;
wire x_7828;
wire x_7829;
wire x_7830;
wire x_7831;
wire x_7832;
wire x_7833;
wire x_7834;
wire x_7835;
wire x_7836;
wire x_7837;
wire x_7838;
wire x_7839;
wire x_7840;
wire x_7841;
wire x_7842;
wire x_7843;
wire x_7844;
wire x_7845;
wire x_7846;
wire x_7847;
wire x_7848;
wire x_7849;
wire x_7850;
wire x_7851;
wire x_7852;
wire x_7853;
wire x_7854;
wire x_7855;
wire x_7856;
wire x_7857;
wire x_7858;
wire x_7859;
wire x_7860;
wire x_7861;
wire x_7862;
wire x_7863;
wire x_7864;
wire x_7865;
wire x_7866;
wire x_7867;
wire x_7868;
wire x_7869;
wire x_7870;
wire x_7871;
wire x_7872;
wire x_7873;
wire x_7874;
wire x_7875;
wire x_7876;
wire x_7877;
wire x_7878;
wire x_7879;
wire x_7880;
wire x_7881;
wire x_7882;
wire x_7883;
wire x_7884;
wire x_7885;
wire x_7886;
wire x_7887;
wire x_7888;
wire x_7889;
wire x_7890;
wire x_7891;
wire x_7892;
wire x_7893;
wire x_7894;
wire x_7895;
wire x_7896;
wire x_7897;
wire x_7898;
wire x_7899;
wire x_7900;
wire x_7901;
wire x_7902;
wire x_7903;
wire x_7904;
wire x_7905;
wire x_7906;
wire x_7907;
wire x_7908;
wire x_7909;
wire x_7910;
wire x_7911;
wire x_7912;
wire x_7913;
wire x_7914;
wire x_7915;
wire x_7916;
wire x_7917;
wire x_7918;
wire x_7919;
wire x_7920;
wire x_7921;
wire x_7922;
wire x_7923;
wire x_7924;
wire x_7925;
wire x_7926;
wire x_7927;
wire x_7928;
wire x_7929;
wire x_7930;
wire x_7931;
wire x_7932;
wire x_7933;
wire x_7934;
wire x_7935;
wire x_7936;
wire x_7937;
wire x_7938;
wire x_7939;
wire x_7940;
wire x_7941;
wire x_7942;
wire x_7943;
wire x_7944;
wire x_7945;
wire x_7946;
wire x_7947;
wire x_7948;
wire x_7949;
wire x_7950;
wire x_7951;
wire x_7952;
wire x_7953;
wire x_7954;
wire x_7955;
wire x_7956;
wire x_7957;
wire x_7958;
wire x_7959;
wire x_7960;
wire x_7961;
wire x_7962;
wire x_7963;
wire x_7964;
wire x_7965;
wire x_7966;
wire x_7967;
wire x_7968;
wire x_7969;
wire x_7970;
wire x_7971;
wire x_7972;
wire x_7973;
wire x_7974;
wire x_7975;
wire x_7976;
wire x_7977;
wire x_7978;
wire x_7979;
wire x_7980;
wire x_7981;
wire x_7982;
wire x_7983;
wire x_7984;
wire x_7985;
wire x_7986;
wire x_7987;
wire x_7988;
wire x_7989;
wire x_7990;
wire x_7991;
wire x_7992;
wire x_7993;
wire x_7994;
wire x_7995;
wire x_7996;
wire x_7997;
wire x_7998;
wire x_7999;
wire x_8000;
wire x_8001;
wire x_8002;
wire x_8003;
wire x_8004;
wire x_8005;
wire x_8006;
wire x_8007;
wire x_8008;
wire x_8009;
wire x_8010;
wire x_8011;
wire x_8012;
wire x_8013;
wire x_8014;
wire x_8015;
wire x_8016;
wire x_8017;
wire x_8018;
wire x_8019;
wire x_8020;
wire x_8021;
wire x_8022;
wire x_8023;
wire x_8024;
wire x_8025;
wire x_8026;
wire x_8027;
wire x_8028;
wire x_8029;
wire x_8030;
wire x_8031;
wire x_8032;
wire x_8033;
wire x_8034;
wire x_8035;
wire x_8036;
wire x_8037;
wire x_8038;
wire x_8039;
wire x_8040;
wire x_8041;
wire x_8042;
wire x_8043;
wire x_8044;
wire x_8045;
wire x_8046;
wire x_8047;
wire x_8048;
wire x_8049;
wire x_8050;
wire x_8051;
wire x_8052;
wire x_8053;
wire x_8054;
wire x_8055;
wire x_8056;
wire x_8057;
wire x_8058;
wire x_8059;
wire x_8060;
wire x_8061;
wire x_8062;
wire x_8063;
wire x_8064;
wire x_8065;
wire x_8066;
wire x_8067;
wire x_8068;
wire x_8069;
wire x_8070;
wire x_8071;
wire x_8072;
wire x_8073;
wire x_8074;
wire x_8075;
wire x_8076;
wire x_8077;
wire x_8078;
wire x_8079;
wire x_8080;
wire x_8081;
wire x_8082;
wire x_8083;
wire x_8084;
wire x_8085;
wire x_8086;
wire x_8087;
wire x_8088;
wire x_8089;
wire x_8090;
wire x_8091;
wire x_8092;
wire x_8093;
wire x_8094;
wire x_8095;
wire x_8096;
wire x_8097;
wire x_8098;
wire x_8099;
wire x_8100;
wire x_8101;
wire x_8102;
wire x_8103;
wire x_8104;
wire x_8105;
wire x_8106;
wire x_8107;
wire x_8108;
wire x_8109;
wire x_8110;
wire x_8111;
wire x_8112;
wire x_8113;
wire x_8114;
wire x_8115;
wire x_8116;
wire x_8117;
wire x_8118;
wire x_8119;
wire x_8120;
wire x_8121;
wire x_8122;
wire x_8123;
wire x_8124;
wire x_8125;
wire x_8126;
wire x_8127;
wire x_8128;
wire x_8129;
wire x_8130;
wire x_8131;
wire x_8132;
wire x_8133;
wire x_8134;
wire x_8135;
wire x_8136;
wire x_8137;
wire x_8138;
wire x_8139;
wire x_8140;
wire x_8141;
wire x_8142;
wire x_8143;
wire x_8144;
wire x_8145;
wire x_8146;
wire x_8147;
wire x_8148;
wire x_8149;
wire x_8150;
wire x_8151;
wire x_8152;
wire x_8153;
wire x_8154;
wire x_8155;
wire x_8156;
wire x_8157;
wire x_8158;
wire x_8159;
wire x_8160;
wire x_8161;
wire x_8162;
wire x_8163;
wire x_8164;
wire x_8165;
wire x_8166;
wire x_8167;
wire x_8168;
wire x_8169;
wire x_8170;
wire x_8171;
wire x_8172;
wire x_8173;
wire x_8174;
wire x_8175;
wire x_8176;
wire x_8177;
wire x_8178;
wire x_8179;
wire x_8180;
wire x_8181;
wire x_8182;
wire x_8183;
wire x_8184;
wire x_8185;
wire x_8186;
wire x_8187;
wire x_8188;
wire x_8189;
wire x_8190;
wire x_8191;
wire x_8192;
wire x_8193;
wire x_8194;
wire x_8195;
wire x_8196;
wire x_8197;
wire x_8198;
wire x_8199;
wire x_8200;
wire x_8201;
wire x_8202;
wire x_8203;
wire x_8204;
wire x_8205;
wire x_8206;
wire x_8207;
wire x_8208;
wire x_8209;
wire x_8210;
wire x_8211;
wire x_8212;
wire x_8213;
wire x_8214;
wire x_8215;
wire x_8216;
wire x_8217;
wire x_8218;
wire x_8219;
wire x_8220;
wire x_8221;
wire x_8222;
wire x_8223;
wire x_8224;
wire x_8225;
wire x_8226;
wire x_8227;
wire x_8228;
wire x_8229;
wire x_8230;
wire x_8231;
wire x_8232;
wire x_8233;
wire x_8234;
wire x_8235;
wire x_8236;
wire x_8237;
wire x_8238;
wire x_8239;
wire x_8240;
wire x_8241;
wire x_8242;
wire x_8243;
wire x_8244;
wire x_8245;
wire x_8246;
wire x_8247;
wire x_8248;
wire x_8249;
wire x_8250;
wire x_8251;
wire x_8252;
wire x_8253;
wire x_8254;
wire x_8255;
wire x_8256;
wire x_8257;
wire x_8258;
wire x_8259;
wire x_8260;
wire x_8261;
wire x_8262;
wire x_8263;
wire x_8264;
wire x_8265;
wire x_8266;
wire x_8267;
wire x_8268;
wire x_8269;
wire x_8270;
wire x_8271;
wire x_8272;
wire x_8273;
wire x_8274;
wire x_8275;
wire x_8276;
wire x_8277;
wire x_8278;
wire x_8279;
wire x_8280;
wire x_8281;
wire x_8282;
wire x_8283;
wire x_8284;
wire x_8285;
wire x_8286;
wire x_8287;
wire x_8288;
wire x_8289;
wire x_8290;
wire x_8291;
wire x_8292;
wire x_8293;
wire x_8294;
wire x_8295;
wire x_8296;
wire x_8297;
wire x_8298;
wire x_8299;
wire x_8300;
wire x_8301;
wire x_8302;
wire x_8303;
wire x_8304;
wire x_8305;
wire x_8306;
wire x_8307;
wire x_8308;
wire x_8309;
wire x_8310;
wire x_8311;
wire x_8312;
wire x_8313;
wire x_8314;
wire x_8315;
wire x_8316;
wire x_8317;
wire x_8318;
wire x_8319;
wire x_8320;
wire x_8321;
wire x_8322;
wire x_8323;
wire x_8324;
wire x_8325;
wire x_8326;
wire x_8327;
wire x_8328;
wire x_8329;
wire x_8330;
wire x_8331;
wire x_8332;
wire x_8333;
wire x_8334;
wire x_8335;
wire x_8336;
wire x_8337;
wire x_8338;
wire x_8339;
wire x_8340;
wire x_8341;
wire x_8342;
wire x_8343;
wire x_8344;
wire x_8345;
wire x_8346;
wire x_8347;
wire x_8348;
wire x_8349;
wire x_8350;
wire x_8351;
wire x_8352;
wire x_8353;
wire x_8354;
wire x_8355;
wire x_8356;
wire x_8357;
wire x_8358;
wire x_8359;
wire x_8360;
wire x_8361;
wire x_8362;
wire x_8363;
wire x_8364;
wire x_8365;
wire x_8366;
wire x_8367;
wire x_8368;
wire x_8369;
wire x_8370;
wire x_8371;
wire x_8372;
wire x_8373;
wire x_8374;
wire x_8375;
wire x_8376;
wire x_8377;
wire x_8378;
wire x_8379;
wire x_8380;
wire x_8381;
wire x_8382;
wire x_8383;
wire x_8384;
wire x_8385;
wire x_8386;
wire x_8387;
wire x_8388;
wire x_8389;
wire x_8390;
wire x_8391;
wire x_8392;
wire x_8393;
wire x_8394;
wire x_8395;
wire x_8396;
wire x_8397;
wire x_8398;
wire x_8399;
wire x_8400;
wire x_8401;
wire x_8402;
wire x_8403;
wire x_8404;
wire x_8405;
wire x_8406;
wire x_8407;
wire x_8408;
wire x_8409;
wire x_8410;
wire x_8411;
wire x_8412;
wire x_8413;
wire x_8414;
wire x_8415;
wire x_8416;
wire x_8417;
wire x_8418;
wire x_8419;
wire x_8420;
wire x_8421;
wire x_8422;
wire x_8423;
wire x_8424;
wire x_8425;
wire x_8426;
wire x_8427;
wire x_8428;
wire x_8429;
wire x_8430;
wire x_8431;
wire x_8432;
wire x_8433;
wire x_8434;
wire x_8435;
wire x_8436;
wire x_8437;
wire x_8438;
wire x_8439;
wire x_8440;
wire x_8441;
wire x_8442;
wire x_8443;
wire x_8444;
wire x_8445;
wire x_8446;
wire x_8447;
wire x_8448;
wire x_8449;
wire x_8450;
wire x_8451;
wire x_8452;
wire x_8453;
wire x_8454;
wire x_8455;
wire x_8456;
wire x_8457;
wire x_8458;
wire x_8459;
wire x_8460;
wire x_8461;
wire x_8462;
wire x_8463;
wire x_8464;
wire x_8465;
wire x_8466;
wire x_8467;
wire x_8468;
wire x_8469;
wire x_8470;
wire x_8471;
wire x_8472;
wire x_8473;
wire x_8474;
wire x_8475;
wire x_8476;
wire x_8477;
wire x_8478;
wire x_8479;
wire x_8480;
wire x_8481;
wire x_8482;
wire x_8483;
wire x_8484;
wire x_8485;
wire x_8486;
wire x_8487;
wire x_8488;
wire x_8489;
wire x_8490;
wire x_8491;
wire x_8492;
wire x_8493;
wire x_8494;
wire x_8495;
wire x_8496;
wire x_8497;
wire x_8498;
wire x_8499;
wire x_8500;
wire x_8501;
wire x_8502;
wire x_8503;
wire x_8504;
wire x_8505;
wire x_8506;
wire x_8507;
wire x_8508;
wire x_8509;
wire x_8510;
wire x_8511;
wire x_8512;
wire x_8513;
wire x_8514;
wire x_8515;
wire x_8516;
wire x_8517;
wire x_8518;
wire x_8519;
wire x_8520;
wire x_8521;
wire x_8522;
wire x_8523;
wire x_8524;
wire x_8525;
wire x_8526;
wire x_8527;
wire x_8528;
wire x_8529;
wire x_8530;
wire x_8531;
wire x_8532;
wire x_8533;
wire x_8534;
wire x_8535;
wire x_8536;
wire x_8537;
wire x_8538;
wire x_8539;
wire x_8540;
wire x_8541;
wire x_8542;
wire x_8543;
wire x_8544;
wire x_8545;
wire x_8546;
wire x_8547;
wire x_8548;
wire x_8549;
wire x_8550;
wire x_8551;
wire x_8552;
wire x_8553;
wire x_8554;
wire x_8555;
wire x_8556;
wire x_8557;
wire x_8558;
wire x_8559;
wire x_8560;
wire x_8561;
wire x_8562;
wire x_8563;
wire x_8564;
wire x_8565;
wire x_8566;
wire x_8567;
wire x_8568;
wire x_8569;
wire x_8570;
wire x_8571;
wire x_8572;
wire x_8573;
wire x_8574;
wire x_8575;
wire x_8576;
wire x_8577;
wire x_8578;
wire x_8579;
wire x_8580;
wire x_8581;
wire x_8582;
wire x_8583;
wire x_8584;
wire x_8585;
wire x_8586;
wire x_8587;
wire x_8588;
wire x_8589;
wire x_8590;
wire x_8591;
wire x_8592;
wire x_8593;
wire x_8594;
wire x_8595;
wire x_8596;
wire x_8597;
wire x_8598;
wire x_8599;
wire x_8600;
wire x_8601;
wire x_8602;
wire x_8603;
wire x_8604;
wire x_8605;
wire x_8606;
wire x_8607;
wire x_8608;
wire x_8609;
wire x_8610;
wire x_8611;
wire x_8612;
wire x_8613;
wire x_8614;
wire x_8615;
wire x_8616;
wire x_8617;
wire x_8618;
wire x_8619;
wire x_8620;
wire x_8621;
wire x_8622;
wire x_8623;
wire x_8624;
wire x_8625;
wire x_8626;
wire x_8627;
wire x_8628;
wire x_8629;
wire x_8630;
wire x_8631;
wire x_8632;
wire x_8633;
wire x_8634;
wire x_8635;
wire x_8636;
wire x_8637;
wire x_8638;
wire x_8639;
wire x_8640;
wire x_8641;
wire x_8642;
wire x_8643;
wire x_8644;
wire x_8645;
wire x_8646;
wire x_8647;
wire x_8648;
wire x_8649;
wire x_8650;
wire x_8651;
wire x_8652;
wire x_8653;
wire x_8654;
wire x_8655;
wire x_8656;
wire x_8657;
wire x_8658;
wire x_8659;
wire x_8660;
wire x_8661;
wire x_8662;
wire x_8663;
wire x_8664;
wire x_8665;
wire x_8666;
wire x_8667;
wire x_8668;
wire x_8669;
wire x_8670;
wire x_8671;
wire x_8672;
wire x_8673;
wire x_8674;
wire x_8675;
wire x_8676;
wire x_8677;
wire x_8678;
wire x_8679;
wire x_8680;
wire x_8681;
wire x_8682;
wire x_8683;
wire x_8684;
wire x_8685;
wire x_8686;
wire x_8687;
wire x_8688;
wire x_8689;
wire x_8690;
wire x_8691;
wire x_8692;
wire x_8693;
wire x_8694;
wire x_8695;
wire x_8696;
wire x_8697;
wire x_8698;
wire x_8699;
wire x_8700;
wire x_8701;
wire x_8702;
wire x_8703;
wire x_8704;
wire x_8705;
wire x_8706;
wire x_8707;
wire x_8708;
wire x_8709;
wire x_8710;
wire x_8711;
wire x_8712;
wire x_8713;
wire x_8714;
wire x_8715;
wire x_8716;
wire x_8717;
wire x_8718;
wire x_8719;
wire x_8720;
wire x_8721;
wire x_8722;
wire x_8723;
wire x_8724;
wire x_8725;
wire x_8726;
wire x_8727;
wire x_8728;
wire x_8729;
wire x_8730;
wire x_8731;
wire x_8732;
wire x_8733;
wire x_8734;
wire x_8735;
wire x_8736;
wire x_8737;
wire x_8738;
wire x_8739;
wire x_8740;
wire x_8741;
wire x_8742;
wire x_8743;
wire x_8744;
wire x_8745;
wire x_8746;
wire x_8747;
wire x_8748;
wire x_8749;
wire x_8750;
wire x_8751;
wire x_8752;
wire x_8753;
wire x_8754;
wire x_8755;
wire x_8756;
wire x_8757;
wire x_8758;
wire x_8759;
wire x_8760;
wire x_8761;
wire x_8762;
wire x_8763;
wire x_8764;
wire x_8765;
wire x_8766;
wire x_8767;
wire x_8768;
wire x_8769;
wire x_8770;
wire x_8771;
wire x_8772;
wire x_8773;
wire x_8774;
wire x_8775;
wire x_8776;
wire x_8777;
wire x_8778;
wire x_8779;
wire x_8780;
wire x_8781;
wire x_8782;
wire x_8783;
wire x_8784;
wire x_8785;
wire x_8786;
wire x_8787;
wire x_8788;
wire x_8789;
wire x_8790;
wire x_8791;
wire x_8792;
wire x_8793;
wire x_8794;
wire x_8795;
wire x_8796;
wire x_8797;
wire x_8798;
wire x_8799;
wire x_8800;
wire x_8801;
wire x_8802;
wire x_8803;
wire x_8804;
wire x_8805;
wire x_8806;
wire x_8807;
wire x_8808;
wire x_8809;
wire x_8810;
wire x_8811;
wire x_8812;
wire x_8813;
wire x_8814;
wire x_8815;
wire x_8816;
wire x_8817;
wire x_8818;
wire x_8819;
wire x_8820;
wire x_8821;
wire x_8822;
wire x_8823;
wire x_8824;
wire x_8825;
wire x_8826;
wire x_8827;
wire x_8828;
wire x_8829;
wire x_8830;
wire x_8831;
wire x_8832;
wire x_8833;
wire x_8834;
wire x_8835;
wire x_8836;
wire x_8837;
wire x_8838;
wire x_8839;
wire x_8840;
wire x_8841;
wire x_8842;
wire x_8843;
wire x_8844;
wire x_8845;
wire x_8846;
wire x_8847;
wire x_8848;
wire x_8849;
wire x_8850;
wire x_8851;
wire x_8852;
wire x_8853;
wire x_8854;
wire x_8855;
wire x_8856;
wire x_8857;
wire x_8858;
wire x_8859;
wire x_8860;
wire x_8861;
wire x_8862;
wire x_8863;
wire x_8864;
wire x_8865;
wire x_8866;
wire x_8867;
wire x_8868;
wire x_8869;
wire x_8870;
wire x_8871;
wire x_8872;
wire x_8873;
wire x_8874;
wire x_8875;
wire x_8876;
wire x_8877;
wire x_8878;
wire x_8879;
wire x_8880;
wire x_8881;
wire x_8882;
wire x_8883;
wire x_8884;
wire x_8885;
wire x_8886;
wire x_8887;
wire x_8888;
wire x_8889;
wire x_8890;
wire x_8891;
wire x_8892;
wire x_8893;
wire x_8894;
wire x_8895;
wire x_8896;
wire x_8897;
wire x_8898;
wire x_8899;
wire x_8900;
wire x_8901;
wire x_8902;
wire x_8903;
wire x_8904;
wire x_8905;
wire x_8906;
wire x_8907;
wire x_8908;
wire x_8909;
wire x_8910;
wire x_8911;
wire x_8912;
wire x_8913;
wire x_8914;
wire x_8915;
wire x_8916;
wire x_8917;
wire x_8918;
wire x_8919;
wire x_8920;
wire x_8921;
wire x_8922;
wire x_8923;
wire x_8924;
wire x_8925;
wire x_8926;
wire x_8927;
wire x_8928;
wire x_8929;
wire x_8930;
wire x_8931;
wire x_8932;
wire x_8933;
wire x_8934;
wire x_8935;
wire x_8936;
wire x_8937;
wire x_8938;
wire x_8939;
wire x_8940;
wire x_8941;
wire x_8942;
wire x_8943;
wire x_8944;
wire x_8945;
wire x_8946;
wire x_8947;
wire x_8948;
wire x_8949;
wire x_8950;
wire x_8951;
wire x_8952;
wire x_8953;
wire x_8954;
wire x_8955;
wire x_8956;
wire x_8957;
wire x_8958;
wire x_8959;
wire x_8960;
wire x_8961;
wire x_8962;
wire x_8963;
wire x_8964;
wire x_8965;
wire x_8966;
wire x_8967;
wire x_8968;
wire x_8969;
wire x_8970;
wire x_8971;
wire x_8972;
wire x_8973;
wire x_8974;
wire x_8975;
wire x_8976;
wire x_8977;
wire x_8978;
wire x_8979;
wire x_8980;
wire x_8981;
wire x_8982;
wire x_8983;
wire x_8984;
wire x_8985;
wire x_8986;
wire x_8987;
wire x_8988;
wire x_8989;
wire x_8990;
wire x_8991;
wire x_8992;
wire x_8993;
wire x_8994;
wire x_8995;
wire x_8996;
wire x_8997;
wire x_8998;
wire x_8999;
wire x_9000;
wire x_9001;
wire x_9002;
wire x_9003;
wire x_9004;
wire x_9005;
wire x_9006;
wire x_9007;
wire x_9008;
wire x_9009;
wire x_9010;
wire x_9011;
wire x_9012;
wire x_9013;
wire x_9014;
wire x_9015;
wire x_9016;
wire x_9017;
wire x_9018;
wire x_9019;
wire x_9020;
wire x_9021;
wire x_9022;
wire x_9023;
wire x_9024;
wire x_9025;
wire x_9026;
wire x_9027;
wire x_9028;
wire x_9029;
wire x_9030;
wire x_9031;
wire x_9032;
wire x_9033;
wire x_9034;
wire x_9035;
wire x_9036;
wire x_9037;
wire x_9038;
wire x_9039;
wire x_9040;
wire x_9041;
wire x_9042;
wire x_9043;
wire x_9044;
wire x_9045;
wire x_9046;
wire x_9047;
wire x_9048;
wire x_9049;
wire x_9050;
wire x_9051;
wire x_9052;
wire x_9053;
wire x_9054;
wire x_9055;
wire x_9056;
wire x_9057;
wire x_9058;
wire x_9059;
wire x_9060;
wire x_9061;
wire x_9062;
wire x_9063;
wire x_9064;
wire x_9065;
wire x_9066;
wire x_9067;
wire x_9068;
wire x_9069;
wire x_9070;
wire x_9071;
wire x_9072;
wire x_9073;
wire x_9074;
wire x_9075;
wire x_9076;
wire x_9077;
wire x_9078;
wire x_9079;
wire x_9080;
wire x_9081;
wire x_9082;
wire x_9083;
wire x_9084;
wire x_9085;
wire x_9086;
wire x_9087;
wire x_9088;
wire x_9089;
wire x_9090;
wire x_9091;
wire x_9092;
wire x_9093;
wire x_9094;
wire x_9095;
wire x_9096;
wire x_9097;
wire x_9098;
wire x_9099;
wire x_9100;
wire x_9101;
wire x_9102;
wire x_9103;
wire x_9104;
wire x_9105;
wire x_9106;
wire x_9107;
wire x_9108;
wire x_9109;
wire x_9110;
wire x_9111;
wire x_9112;
wire x_9113;
wire x_9114;
wire x_9115;
wire x_9116;
wire x_9117;
wire x_9118;
wire x_9119;
wire x_9120;
wire x_9121;
wire x_9122;
wire x_9123;
wire x_9124;
wire x_9125;
wire x_9126;
wire x_9127;
wire x_9128;
wire x_9129;
wire x_9130;
wire x_9131;
wire x_9132;
wire x_9133;
wire x_9134;
wire x_9135;
wire x_9136;
wire x_9137;
wire x_9138;
wire x_9139;
wire x_9140;
wire x_9141;
wire x_9142;
wire x_9143;
wire x_9144;
wire x_9145;
wire x_9146;
wire x_9147;
wire x_9148;
wire x_9149;
wire x_9150;
wire x_9151;
wire x_9152;
wire x_9153;
wire x_9154;
wire x_9155;
wire x_9156;
wire x_9157;
wire x_9158;
wire x_9159;
wire x_9160;
wire x_9161;
wire x_9162;
wire x_9163;
wire x_9164;
wire x_9165;
wire x_9166;
wire x_9167;
wire x_9168;
wire x_9169;
wire x_9170;
wire x_9171;
wire x_9172;
wire x_9173;
wire x_9174;
wire x_9175;
wire x_9176;
wire x_9177;
wire x_9178;
wire x_9179;
wire x_9180;
wire x_9181;
wire x_9182;
wire x_9183;
wire x_9184;
wire x_9185;
wire x_9186;
wire x_9187;
wire x_9188;
wire x_9189;
wire x_9190;
wire x_9191;
wire x_9192;
wire x_9193;
wire x_9194;
wire x_9195;
wire x_9196;
wire x_9197;
wire x_9198;
wire x_9199;
wire x_9200;
wire x_9201;
wire x_9202;
wire x_9203;
wire x_9204;
wire x_9205;
wire x_9206;
wire x_9207;
wire x_9208;
wire x_9209;
wire x_9210;
wire x_9211;
wire x_9212;
wire x_9213;
wire x_9214;
wire x_9215;
wire x_9216;
wire x_9217;
wire x_9218;
wire x_9219;
wire x_9220;
wire x_9221;
wire x_9222;
wire x_9223;
wire x_9224;
wire x_9225;
wire x_9226;
wire x_9227;
wire x_9228;
wire x_9229;
wire x_9230;
wire x_9231;
wire x_9232;
wire x_9233;
wire x_9234;
wire x_9235;
wire x_9236;
wire x_9237;
wire x_9238;
wire x_9239;
wire x_9240;
wire x_9241;
wire x_9242;
wire x_9243;
wire x_9244;
wire x_9245;
wire x_9246;
wire x_9247;
wire x_9248;
wire x_9249;
wire x_9250;
wire x_9251;
wire x_9252;
wire x_9253;
wire x_9254;
wire x_9255;
wire x_9256;
wire x_9257;
wire x_9258;
wire x_9259;
wire x_9260;
wire x_9261;
wire x_9262;
wire x_9263;
wire x_9264;
wire x_9265;
wire x_9266;
wire x_9267;
wire x_9268;
wire x_9269;
wire x_9270;
wire x_9271;
wire x_9272;
wire x_9273;
wire x_9274;
wire x_9275;
wire x_9276;
wire x_9277;
wire x_9278;
wire x_9279;
wire x_9280;
wire x_9281;
wire x_9282;
wire x_9283;
wire x_9284;
wire x_9285;
wire x_9286;
wire x_9287;
wire x_9288;
wire x_9289;
wire x_9290;
wire x_9291;
wire x_9292;
wire x_9293;
wire x_9294;
wire x_9295;
wire x_9296;
wire x_9297;
wire x_9298;
wire x_9299;
wire x_9300;
wire x_9301;
wire x_9302;
wire x_9303;
wire x_9304;
wire x_9305;
wire x_9306;
wire x_9307;
wire x_9308;
wire x_9309;
wire x_9310;
wire x_9311;
wire x_9312;
wire x_9313;
wire x_9314;
wire x_9315;
wire x_9316;
wire x_9317;
wire x_9318;
wire x_9319;
wire x_9320;
wire x_9321;
wire x_9322;
wire x_9323;
wire x_9324;
wire x_9325;
wire x_9326;
wire x_9327;
wire x_9328;
wire x_9329;
wire x_9330;
wire x_9331;
wire x_9332;
wire x_9333;
wire x_9334;
wire x_9335;
wire x_9336;
wire x_9337;
wire x_9338;
wire x_9339;
wire x_9340;
wire x_9341;
wire x_9342;
wire x_9343;
wire x_9344;
wire x_9345;
wire x_9346;
wire x_9347;
wire x_9348;
wire x_9349;
wire x_9350;
wire x_9351;
wire x_9352;
wire x_9353;
wire x_9354;
wire x_9355;
wire x_9356;
wire x_9357;
wire x_9358;
wire x_9359;
wire x_9360;
wire x_9361;
wire x_9362;
wire x_9363;
wire x_9364;
wire x_9365;
wire x_9366;
wire x_9367;
wire x_9368;
wire x_9369;
wire x_9370;
wire x_9371;
wire x_9372;
wire x_9373;
wire x_9374;
wire x_9375;
wire x_9376;
wire x_9377;
wire x_9378;
wire x_9379;
wire x_9380;
wire x_9381;
wire x_9382;
wire x_9383;
wire x_9384;
wire x_9385;
wire x_9386;
wire x_9387;
wire x_9388;
wire x_9389;
wire x_9390;
wire x_9391;
wire x_9392;
wire x_9393;
wire x_9394;
wire x_9395;
wire x_9396;
wire x_9397;
wire x_9398;
wire x_9399;
wire x_9400;
wire x_9401;
wire x_9402;
wire x_9403;
wire x_9404;
wire x_9405;
wire x_9406;
wire x_9407;
wire x_9408;
wire x_9409;
wire x_9410;
wire x_9411;
wire x_9412;
wire x_9413;
wire x_9414;
wire x_9415;
wire x_9416;
wire x_9417;
wire x_9418;
wire x_9419;
wire x_9420;
wire x_9421;
wire x_9422;
wire x_9423;
wire x_9424;
wire x_9425;
wire x_9426;
wire x_9427;
wire x_9428;
wire x_9429;
wire x_9430;
wire x_9431;
wire x_9432;
wire x_9433;
wire x_9434;
wire x_9435;
wire x_9436;
wire x_9437;
wire x_9438;
wire x_9439;
wire x_9440;
wire x_9441;
wire x_9442;
wire x_9443;
wire x_9444;
wire x_9445;
wire x_9446;
wire x_9447;
wire x_9448;
wire x_9449;
wire x_9450;
wire x_9451;
wire x_9452;
wire x_9453;
wire x_9454;
wire x_9455;
wire x_9456;
wire x_9457;
wire x_9458;
wire x_9459;
wire x_9460;
wire x_9461;
wire x_9462;
wire x_9463;
wire x_9464;
wire x_9465;
wire x_9466;
wire x_9467;
wire x_9468;
wire x_9469;
wire x_9470;
wire x_9471;
wire x_9472;
wire x_9473;
wire x_9474;
wire x_9475;
wire x_9476;
wire x_9477;
wire x_9478;
wire x_9479;
wire x_9480;
wire x_9481;
wire x_9482;
wire x_9483;
wire x_9484;
wire x_9485;
wire x_9486;
wire x_9487;
wire x_9488;
wire x_9489;
wire x_9490;
wire x_9491;
wire x_9492;
wire x_9493;
wire x_9494;
wire x_9495;
wire x_9496;
wire x_9497;
wire x_9498;
wire x_9499;
wire x_9500;
wire x_9501;
wire x_9502;
wire x_9503;
wire x_9504;
wire x_9505;
wire x_9506;
wire x_9507;
wire x_9508;
wire x_9509;
wire x_9510;
wire x_9511;
wire x_9512;
wire x_9513;
wire x_9514;
wire x_9515;
wire x_9516;
wire x_9517;
wire x_9518;
wire x_9519;
wire x_9520;
wire x_9521;
wire x_9522;
wire x_9523;
wire x_9524;
wire x_9525;
wire x_9526;
wire x_9527;
wire x_9528;
wire x_9529;
wire x_9530;
wire x_9531;
wire x_9532;
wire x_9533;
wire x_9534;
wire x_9535;
wire x_9536;
wire x_9537;
wire x_9538;
wire x_9539;
wire x_9540;
wire x_9541;
wire x_9542;
wire x_9543;
wire x_9544;
wire x_9545;
wire x_9546;
wire x_9547;
wire x_9548;
wire x_9549;
wire x_9550;
wire x_9551;
wire x_9552;
wire x_9553;
wire x_9554;
wire x_9555;
wire x_9556;
wire x_9557;
wire x_9558;
wire x_9559;
wire x_9560;
wire x_9561;
wire x_9562;
wire x_9563;
wire x_9564;
wire x_9565;
wire x_9566;
wire x_9567;
wire x_9568;
wire x_9569;
wire x_9570;
wire x_9571;
wire x_9572;
wire x_9573;
wire x_9574;
wire x_9575;
wire x_9576;
wire x_9577;
wire x_9578;
wire x_9579;
wire x_9580;
wire x_9581;
wire x_9582;
wire x_9583;
wire x_9584;
wire x_9585;
wire x_9586;
wire x_9587;
wire x_9588;
wire x_9589;
wire x_9590;
wire x_9591;
wire x_9592;
wire x_9593;
wire x_9594;
wire x_9595;
wire x_9596;
wire x_9597;
wire x_9598;
wire x_9599;
wire x_9600;
wire x_9601;
wire x_9602;
wire x_9603;
wire x_9604;
wire x_9605;
wire x_9606;
wire x_9607;
wire x_9608;
wire x_9609;
wire x_9610;
wire x_9611;
wire x_9612;
wire x_9613;
wire x_9614;
wire x_9615;
wire x_9616;
wire x_9617;
wire x_9618;
wire x_9619;
wire x_9620;
wire x_9621;
wire x_9622;
wire x_9623;
wire x_9624;
wire x_9625;
wire x_9626;
wire x_9627;
wire x_9628;
wire x_9629;
wire x_9630;
wire x_9631;
wire x_9632;
wire x_9633;
wire x_9634;
wire x_9635;
wire x_9636;
wire x_9637;
wire x_9638;
wire x_9639;
wire x_9640;
wire x_9641;
wire x_9642;
wire x_9643;
wire x_9644;
wire x_9645;
wire x_9646;
wire x_9647;
wire x_9648;
wire x_9649;
wire x_9650;
wire x_9651;
wire x_9652;
wire x_9653;
wire x_9654;
wire x_9655;
wire x_9656;
wire x_9657;
wire x_9658;
wire x_9659;
wire x_9660;
wire x_9661;
wire x_9662;
wire x_9663;
wire x_9664;
wire x_9665;
wire x_9666;
wire x_9667;
wire x_9668;
wire x_9669;
wire x_9670;
wire x_9671;
wire x_9672;
wire x_9673;
wire x_9674;
wire x_9675;
wire x_9676;
wire x_9677;
wire x_9678;
wire x_9679;
wire x_9680;
wire x_9681;
wire x_9682;
wire x_9683;
wire x_9684;
wire x_9685;
wire x_9686;
wire x_9687;
wire x_9688;
wire x_9689;
wire x_9690;
wire x_9691;
wire x_9692;
wire x_9693;
wire x_9694;
wire x_9695;
wire x_9696;
wire x_9697;
wire x_9698;
wire x_9699;
wire x_9700;
wire x_9701;
wire x_9702;
wire x_9703;
wire x_9704;
wire x_9705;
wire x_9706;
wire x_9707;
wire x_9708;
wire x_9709;
wire x_9710;
wire x_9711;
wire x_9712;
wire x_9713;
wire x_9714;
wire x_9715;
wire x_9716;
wire x_9717;
wire x_9718;
wire x_9719;
wire x_9720;
wire x_9721;
wire x_9722;
wire x_9723;
wire x_9724;
wire x_9725;
wire x_9726;
wire x_9727;
wire x_9728;
wire x_9729;
wire x_9730;
wire x_9731;
wire x_9732;
wire x_9733;
wire x_9734;
wire x_9735;
wire x_9736;
wire x_9737;
wire x_9738;
wire x_9739;
wire x_9740;
wire x_9741;
wire x_9742;
wire x_9743;
wire x_9744;
wire x_9745;
wire x_9746;
wire x_9747;
wire x_9748;
wire x_9749;
wire x_9750;
wire x_9751;
wire x_9752;
wire x_9753;
wire x_9754;
wire x_9755;
wire x_9756;
wire x_9757;
wire x_9758;
wire x_9759;
wire x_9760;
wire x_9761;
wire x_9762;
wire x_9763;
wire x_9764;
wire x_9765;
wire x_9766;
wire x_9767;
wire x_9768;
wire x_9769;
wire x_9770;
wire x_9771;
wire x_9772;
wire x_9773;
wire x_9774;
wire x_9775;
wire x_9776;
wire x_9777;
wire x_9778;
wire x_9779;
wire x_9780;
wire x_9781;
wire x_9782;
wire x_9783;
wire x_9784;
wire x_9785;
wire x_9786;
wire x_9787;
wire x_9788;
wire x_9789;
wire x_9790;
wire x_9791;
wire x_9792;
wire x_9793;
wire x_9794;
wire x_9795;
wire x_9796;
wire x_9797;
wire x_9798;
wire x_9799;
wire x_9800;
wire x_9801;
wire x_9802;
wire x_9803;
wire x_9804;
wire x_9805;
wire x_9806;
wire x_9807;
wire x_9808;
wire x_9809;
wire x_9810;
wire x_9811;
wire x_9812;
wire x_9813;
wire x_9814;
wire x_9815;
wire x_9816;
wire x_9817;
wire x_9818;
wire x_9819;
wire x_9820;
wire x_9821;
wire x_9822;
wire x_9823;
wire x_9824;
wire x_9825;
wire x_9826;
wire x_9827;
wire x_9828;
wire x_9829;
wire x_9830;
wire x_9831;
wire x_9832;
wire x_9833;
wire x_9834;
wire x_9835;
wire x_9836;
wire x_9837;
wire x_9838;
wire x_9839;
wire x_9840;
wire x_9841;
wire x_9842;
wire x_9843;
wire x_9844;
wire x_9845;
wire x_9846;
wire x_9847;
wire x_9848;
wire x_9849;
wire x_9850;
wire x_9851;
wire x_9852;
wire x_9853;
wire x_9854;
wire x_9855;
wire x_9856;
wire x_9857;
wire x_9858;
wire x_9859;
wire x_9860;
wire x_9861;
wire x_9862;
wire x_9863;
wire x_9864;
wire x_9865;
wire x_9866;
wire x_9867;
wire x_9868;
wire x_9869;
wire x_9870;
wire x_9871;
wire x_9872;
wire x_9873;
wire x_9874;
wire x_9875;
wire x_9876;
wire x_9877;
wire x_9878;
wire x_9879;
wire x_9880;
wire x_9881;
wire x_9882;
wire x_9883;
wire x_9884;
wire x_9885;
wire x_9886;
wire x_9887;
wire x_9888;
wire x_9889;
wire x_9890;
wire x_9891;
wire x_9892;
wire x_9893;
wire x_9894;
wire x_9895;
wire x_9896;
wire x_9897;
wire x_9898;
wire x_9899;
wire x_9900;
wire x_9901;
wire x_9902;
wire x_9903;
wire x_9904;
wire x_9905;
wire x_9906;
wire x_9907;
wire x_9908;
wire x_9909;
wire x_9910;
wire x_9911;
wire x_9912;
wire x_9913;
wire x_9914;
wire x_9915;
wire x_9916;
wire x_9917;
wire x_9918;
wire x_9919;
wire x_9920;
wire x_9921;
wire x_9922;
wire x_9923;
wire x_9924;
wire x_9925;
wire x_9926;
wire x_9927;
wire x_9928;
wire x_9929;
wire x_9930;
wire x_9931;
wire x_9932;
wire x_9933;
wire x_9934;
wire x_9935;
wire x_9936;
wire x_9937;
wire x_9938;
wire x_9939;
wire x_9940;
wire x_9941;
wire x_9942;
wire x_9943;
wire x_9944;
wire x_9945;
wire x_9946;
wire x_9947;
wire x_9948;
wire x_9949;
wire x_9950;
wire x_9951;
wire x_9952;
wire x_9953;
wire x_9954;
wire x_9955;
wire x_9956;
wire x_9957;
wire x_9958;
wire x_9959;
wire x_9960;
wire x_9961;
wire x_9962;
wire x_9963;
wire x_9964;
wire x_9965;
wire x_9966;
wire x_9967;
wire x_9968;
wire x_9969;
wire x_9970;
wire x_9971;
wire x_9972;
wire x_9973;
wire x_9974;
wire x_9975;
wire x_9976;
wire x_9977;
wire x_9978;
wire x_9979;
wire x_9980;
wire x_9981;
wire x_9982;
wire x_9983;
wire x_9984;
wire x_9985;
wire x_9986;
wire x_9987;
wire x_9988;
wire x_9989;
wire x_9990;
wire x_9991;
wire x_9992;
wire x_9993;
wire x_9994;
wire x_9995;
wire x_9996;
wire x_9997;
wire x_9998;
wire x_9999;
wire x_10000;
wire x_10001;
wire x_10002;
wire x_10003;
wire x_10004;
wire x_10005;
wire x_10006;
wire x_10007;
wire x_10008;
wire x_10009;
wire x_10010;
wire x_10011;
wire x_10012;
wire x_10013;
wire x_10014;
wire x_10015;
wire x_10016;
wire x_10017;
wire x_10018;
wire x_10019;
wire x_10020;
wire x_10021;
wire x_10022;
wire x_10023;
wire x_10024;
wire x_10025;
wire x_10026;
wire x_10027;
wire x_10028;
wire x_10029;
wire x_10030;
wire x_10031;
wire x_10032;
wire x_10033;
wire x_10034;
wire x_10035;
wire x_10036;
wire x_10037;
wire x_10038;
wire x_10039;
wire x_10040;
wire x_10041;
wire x_10042;
wire x_10043;
wire x_10044;
wire x_10045;
wire x_10046;
wire x_10047;
wire x_10048;
wire x_10049;
wire x_10050;
wire x_10051;
wire x_10052;
wire x_10053;
wire x_10054;
wire x_10055;
wire x_10056;
wire x_10057;
wire x_10058;
wire x_10059;
wire x_10060;
wire x_10061;
wire x_10062;
wire x_10063;
wire x_10064;
wire x_10065;
wire x_10066;
wire x_10067;
wire x_10068;
wire x_10069;
wire x_10070;
wire x_10071;
wire x_10072;
wire x_10073;
wire x_10074;
wire x_10075;
wire x_10076;
wire x_10077;
wire x_10078;
wire x_10079;
wire x_10080;
wire x_10081;
wire x_10082;
wire x_10083;
wire x_10084;
wire x_10085;
wire x_10086;
wire x_10087;
wire x_10088;
wire x_10089;
wire x_10090;
wire x_10091;
wire x_10092;
wire x_10093;
wire x_10094;
wire x_10095;
wire x_10096;
wire x_10097;
wire x_10098;
wire x_10099;
wire x_10100;
wire x_10101;
wire x_10102;
wire x_10103;
wire x_10104;
wire x_10105;
wire x_10106;
wire x_10107;
wire x_10108;
wire x_10109;
wire x_10110;
wire x_10111;
wire x_10112;
wire x_10113;
wire x_10114;
wire x_10115;
wire x_10116;
wire x_10117;
wire x_10118;
wire x_10119;
wire x_10120;
wire x_10121;
wire x_10122;
wire x_10123;
wire x_10124;
wire x_10125;
wire x_10126;
wire x_10127;
wire x_10128;
wire x_10129;
wire x_10130;
wire x_10131;
wire x_10132;
wire x_10133;
wire x_10134;
wire x_10135;
wire x_10136;
wire x_10137;
wire x_10138;
wire x_10139;
wire x_10140;
wire x_10141;
wire x_10142;
wire x_10143;
wire x_10144;
wire x_10145;
wire x_10146;
wire x_10147;
wire x_10148;
wire x_10149;
wire x_10150;
wire x_10151;
wire x_10152;
wire x_10153;
wire x_10154;
wire x_10155;
wire x_10156;
wire x_10157;
wire x_10158;
wire x_10159;
wire x_10160;
wire x_10161;
wire x_10162;
wire x_10163;
wire x_10164;
wire x_10165;
wire x_10166;
wire x_10167;
wire x_10168;
wire x_10169;
wire x_10170;
wire x_10171;
wire x_10172;
wire x_10173;
wire x_10174;
wire x_10175;
wire x_10176;
wire x_10177;
wire x_10178;
wire x_10179;
wire x_10180;
wire x_10181;
wire x_10182;
wire x_10183;
wire x_10184;
wire x_10185;
wire x_10186;
wire x_10187;
wire x_10188;
wire x_10189;
wire x_10190;
wire x_10191;
wire x_10192;
wire x_10193;
wire x_10194;
wire x_10195;
wire x_10196;
wire x_10197;
wire x_10198;
wire x_10199;
wire x_10200;
wire x_10201;
wire x_10202;
wire x_10203;
wire x_10204;
wire x_10205;
wire x_10206;
wire x_10207;
wire x_10208;
wire x_10209;
wire x_10210;
wire x_10211;
wire x_10212;
wire x_10213;
wire x_10214;
wire x_10215;
wire x_10216;
wire x_10217;
wire x_10218;
wire x_10219;
wire x_10220;
wire x_10221;
wire x_10222;
wire x_10223;
wire x_10224;
wire x_10225;
wire x_10226;
wire x_10227;
wire x_10228;
wire x_10229;
wire x_10230;
wire x_10231;
wire x_10232;
wire x_10233;
wire x_10234;
wire x_10235;
wire x_10236;
wire x_10237;
wire x_10238;
wire x_10239;
wire x_10240;
wire x_10241;
wire x_10242;
wire x_10243;
wire x_10244;
wire x_10245;
wire x_10246;
wire x_10247;
wire x_10248;
wire x_10249;
wire x_10250;
wire x_10251;
wire x_10252;
wire x_10253;
wire x_10254;
wire x_10255;
wire x_10256;
wire x_10257;
wire x_10258;
wire x_10259;
wire x_10260;
wire x_10261;
wire x_10262;
wire x_10263;
wire x_10264;
wire x_10265;
wire x_10266;
wire x_10267;
wire x_10268;
wire x_10269;
wire x_10270;
wire x_10271;
wire x_10272;
wire x_10273;
wire x_10274;
wire x_10275;
wire x_10276;
wire x_10277;
wire x_10278;
wire x_10279;
wire x_10280;
wire x_10281;
wire x_10282;
wire x_10283;
wire x_10284;
wire x_10285;
wire x_10286;
wire x_10287;
wire x_10288;
wire x_10289;
wire x_10290;
wire x_10291;
wire x_10292;
wire x_10293;
wire x_10294;
wire x_10295;
wire x_10296;
wire x_10297;
wire x_10298;
wire x_10299;
wire x_10300;
wire x_10301;
wire x_10302;
wire x_10303;
wire x_10304;
wire x_10305;
wire x_10306;
wire x_10307;
wire x_10308;
wire x_10309;
wire x_10310;
wire x_10311;
wire x_10312;
wire x_10313;
wire x_10314;
wire x_10315;
wire x_10316;
wire x_10317;
wire x_10318;
wire x_10319;
wire x_10320;
wire x_10321;
wire x_10322;
wire x_10323;
wire x_10324;
wire x_10325;
wire x_10326;
wire x_10327;
wire x_10328;
wire x_10329;
wire x_10330;
wire x_10331;
wire x_10332;
wire x_10333;
wire x_10334;
wire x_10335;
wire x_10336;
wire x_10337;
wire x_10338;
wire x_10339;
wire x_10340;
wire x_10341;
wire x_10342;
wire x_10343;
wire x_10344;
wire x_10345;
wire x_10346;
wire x_10347;
wire x_10348;
wire x_10349;
wire x_10350;
wire x_10351;
wire x_10352;
wire x_10353;
wire x_10354;
wire x_10355;
wire x_10356;
wire x_10357;
wire x_10358;
wire x_10359;
wire x_10360;
wire x_10361;
wire x_10362;
wire x_10363;
wire x_10364;
wire x_10365;
wire x_10366;
wire x_10367;
wire x_10368;
wire x_10369;
wire x_10370;
wire x_10371;
wire x_10372;
wire x_10373;
wire x_10374;
wire x_10375;
wire x_10376;
wire x_10377;
wire x_10378;
wire x_10379;
wire x_10380;
wire x_10381;
wire x_10382;
wire x_10383;
wire x_10384;
wire x_10385;
wire x_10386;
wire x_10387;
wire x_10388;
wire x_10389;
wire x_10390;
wire x_10391;
wire x_10392;
wire x_10393;
wire x_10394;
wire x_10395;
wire x_10396;
wire x_10397;
wire x_10398;
wire x_10399;
wire x_10400;
wire x_10401;
wire x_10402;
wire x_10403;
wire x_10404;
wire x_10405;
wire x_10406;
wire x_10407;
wire x_10408;
wire x_10409;
wire x_10410;
wire x_10411;
wire x_10412;
wire x_10413;
wire x_10414;
wire x_10415;
wire x_10416;
wire x_10417;
wire x_10418;
wire x_10419;
wire x_10420;
wire x_10421;
wire x_10422;
wire x_10423;
wire x_10424;
wire x_10425;
wire x_10426;
wire x_10427;
wire x_10428;
wire x_10429;
wire x_10430;
wire x_10431;
wire x_10432;
wire x_10433;
wire x_10434;
wire x_10435;
wire x_10436;
wire x_10437;
wire x_10438;
wire x_10439;
wire x_10440;
wire x_10441;
wire x_10442;
wire x_10443;
wire x_10444;
wire x_10445;
wire x_10446;
wire x_10447;
wire x_10448;
wire x_10449;
wire x_10450;
wire x_10451;
wire x_10452;
wire x_10453;
wire x_10454;
wire x_10455;
wire x_10456;
wire x_10457;
wire x_10458;
wire x_10459;
wire x_10460;
wire x_10461;
wire x_10462;
wire x_10463;
wire x_10464;
wire x_10465;
wire x_10466;
wire x_10467;
wire x_10468;
wire x_10469;
wire x_10470;
wire x_10471;
wire x_10472;
wire x_10473;
wire x_10474;
wire x_10475;
wire x_10476;
wire x_10477;
wire x_10478;
wire x_10479;
wire x_10480;
wire x_10481;
wire x_10482;
wire x_10483;
wire x_10484;
wire x_10485;
wire x_10486;
wire x_10487;
wire x_10488;
wire x_10489;
wire x_10490;
wire x_10491;
wire x_10492;
wire x_10493;
wire x_10494;
wire x_10495;
wire x_10496;
wire x_10497;
wire x_10498;
wire x_10499;
wire x_10500;
wire x_10501;
wire x_10502;
wire x_10503;
wire x_10504;
wire x_10505;
wire x_10506;
wire x_10507;
wire x_10508;
wire x_10509;
wire x_10510;
wire x_10511;
wire x_10512;
wire x_10513;
wire x_10514;
wire x_10515;
wire x_10516;
wire x_10517;
wire x_10518;
wire x_10519;
wire x_10520;
wire x_10521;
wire x_10522;
wire x_10523;
wire x_10524;
wire x_10525;
wire x_10526;
wire x_10527;
wire x_10528;
wire x_10529;
wire x_10530;
wire x_10531;
wire x_10532;
wire x_10533;
wire x_10534;
wire x_10535;
wire x_10536;
wire x_10537;
wire x_10538;
wire x_10539;
wire x_10540;
wire x_10541;
wire x_10542;
wire x_10543;
wire x_10544;
wire x_10545;
wire x_10546;
wire x_10547;
wire x_10548;
wire x_10549;
wire x_10550;
wire x_10551;
wire x_10552;
wire x_10553;
wire x_10554;
wire x_10555;
wire x_10556;
wire x_10557;
wire x_10558;
wire x_10559;
wire x_10560;
wire x_10561;
wire x_10562;
wire x_10563;
wire x_10564;
wire x_10565;
wire x_10566;
wire x_10567;
wire x_10568;
wire x_10569;
wire x_10570;
wire x_10571;
wire x_10572;
wire x_10573;
wire x_10574;
wire x_10575;
wire x_10576;
wire x_10577;
wire x_10578;
wire x_10579;
wire x_10580;
wire x_10581;
wire x_10582;
wire x_10583;
wire x_10584;
wire x_10585;
wire x_10586;
wire x_10587;
wire x_10588;
wire x_10589;
wire x_10590;
wire x_10591;
wire x_10592;
wire x_10593;
wire x_10594;
wire x_10595;
wire x_10596;
wire x_10597;
wire x_10598;
wire x_10599;
wire x_10600;
wire x_10601;
wire x_10602;
wire x_10603;
wire x_10604;
wire x_10605;
wire x_10606;
wire x_10607;
wire x_10608;
wire x_10609;
wire x_10610;
wire x_10611;
wire x_10612;
wire x_10613;
wire x_10614;
wire x_10615;
wire x_10616;
wire x_10617;
wire x_10618;
wire x_10619;
wire x_10620;
wire x_10621;
wire x_10622;
wire x_10623;
wire x_10624;
wire x_10625;
wire x_10626;
wire x_10627;
wire x_10628;
wire x_10629;
wire x_10630;
wire x_10631;
wire x_10632;
wire x_10633;
wire x_10634;
wire x_10635;
wire x_10636;
wire x_10637;
wire x_10638;
wire x_10639;
wire x_10640;
wire x_10641;
wire x_10642;
wire x_10643;
wire x_10644;
wire x_10645;
wire x_10646;
wire x_10647;
wire x_10648;
wire x_10649;
wire x_10650;
wire x_10651;
wire x_10652;
wire x_10653;
wire x_10654;
wire x_10655;
wire x_10656;
wire x_10657;
wire x_10658;
wire x_10659;
wire x_10660;
wire x_10661;
wire x_10662;
wire x_10663;
wire x_10664;
wire x_10665;
wire x_10666;
wire x_10667;
wire x_10668;
wire x_10669;
wire x_10670;
wire x_10671;
wire x_10672;
wire x_10673;
wire x_10674;
wire x_10675;
wire x_10676;
wire x_10677;
wire x_10678;
wire x_10679;
wire x_10680;
wire x_10681;
wire x_10682;
wire x_10683;
wire x_10684;
wire x_10685;
wire x_10686;
wire x_10687;
wire x_10688;
wire x_10689;
wire x_10690;
wire x_10691;
wire x_10692;
wire x_10693;
wire x_10694;
wire x_10695;
wire x_10696;
wire x_10697;
wire x_10698;
wire x_10699;
wire x_10700;
wire x_10701;
wire x_10702;
wire x_10703;
wire x_10704;
wire x_10705;
wire x_10706;
wire x_10707;
wire x_10708;
wire x_10709;
wire x_10710;
wire x_10711;
wire x_10712;
wire x_10713;
wire x_10714;
wire x_10715;
wire x_10716;
wire x_10717;
wire x_10718;
wire x_10719;
wire x_10720;
wire x_10721;
wire x_10722;
wire x_10723;
wire x_10724;
wire x_10725;
wire x_10726;
wire x_10727;
wire x_10728;
wire x_10729;
wire x_10730;
wire x_10731;
wire x_10732;
wire x_10733;
wire x_10734;
wire x_10735;
wire x_10736;
wire x_10737;
wire x_10738;
wire x_10739;
wire x_10740;
wire x_10741;
wire x_10742;
wire x_10743;
wire x_10744;
wire x_10745;
wire x_10746;
wire x_10747;
wire x_10748;
wire x_10749;
wire x_10750;
wire x_10751;
wire x_10752;
wire x_10753;
wire x_10754;
wire x_10755;
wire x_10756;
wire x_10757;
wire x_10758;
wire x_10759;
wire x_10760;
wire x_10761;
wire x_10762;
wire x_10763;
wire x_10764;
wire x_10765;
wire x_10766;
wire x_10767;
wire x_10768;
wire x_10769;
wire x_10770;
wire x_10771;
wire x_10772;
wire x_10773;
wire x_10774;
wire x_10775;
wire x_10776;
wire x_10777;
wire x_10778;
wire x_10779;
wire x_10780;
wire x_10781;
wire x_10782;
wire x_10783;
wire x_10784;
wire x_10785;
wire x_10786;
wire x_10787;
wire x_10788;
wire x_10789;
wire x_10790;
wire x_10791;
wire x_10792;
wire x_10793;
wire x_10794;
wire x_10795;
wire x_10796;
wire x_10797;
wire x_10798;
wire x_10799;
wire x_10800;
wire x_10801;
wire x_10802;
wire x_10803;
wire x_10804;
wire x_10805;
wire x_10806;
wire x_10807;
wire x_10808;
wire x_10809;
wire x_10810;
wire x_10811;
wire x_10812;
wire x_10813;
wire x_10814;
wire x_10815;
wire x_10816;
wire x_10817;
wire x_10818;
wire x_10819;
wire x_10820;
wire x_10821;
wire x_10822;
wire x_10823;
wire x_10824;
wire x_10825;
wire x_10826;
wire x_10827;
wire x_10828;
wire x_10829;
wire x_10830;
wire x_10831;
wire x_10832;
wire x_10833;
wire x_10834;
wire x_10835;
wire x_10836;
wire x_10837;
wire x_10838;
wire x_10839;
wire x_10840;
wire x_10841;
wire x_10842;
wire x_10843;
wire x_10844;
wire x_10845;
wire x_10846;
wire x_10847;
wire x_10848;
wire x_10849;
wire x_10850;
wire x_10851;
wire x_10852;
wire x_10853;
wire x_10854;
wire x_10855;
wire x_10856;
wire x_10857;
wire x_10858;
wire x_10859;
wire x_10860;
wire x_10861;
wire x_10862;
wire x_10863;
wire x_10864;
wire x_10865;
wire x_10866;
wire x_10867;
wire x_10868;
wire x_10869;
wire x_10870;
wire x_10871;
wire x_10872;
wire x_10873;
wire x_10874;
wire x_10875;
wire x_10876;
wire x_10877;
wire x_10878;
wire x_10879;
wire x_10880;
wire x_10881;
wire x_10882;
wire x_10883;
wire x_10884;
wire x_10885;
wire x_10886;
wire x_10887;
wire x_10888;
wire x_10889;
wire x_10890;
wire x_10891;
wire x_10892;
wire x_10893;
wire x_10894;
wire x_10895;
wire x_10896;
wire x_10897;
wire x_10898;
wire x_10899;
wire x_10900;
wire x_10901;
wire x_10902;
wire x_10903;
wire x_10904;
wire x_10905;
wire x_10906;
wire x_10907;
wire x_10908;
wire x_10909;
wire x_10910;
wire x_10911;
wire x_10912;
wire x_10913;
wire x_10914;
wire x_10915;
wire x_10916;
wire x_10917;
wire x_10918;
wire x_10919;
wire x_10920;
wire x_10921;
wire x_10922;
wire x_10923;
wire x_10924;
wire x_10925;
wire x_10926;
wire x_10927;
wire x_10928;
wire x_10929;
wire x_10930;
wire x_10931;
wire x_10932;
wire x_10933;
wire x_10934;
wire x_10935;
wire x_10936;
wire x_10937;
wire x_10938;
wire x_10939;
wire x_10940;
wire x_10941;
wire x_10942;
wire x_10943;
wire x_10944;
wire x_10945;
wire x_10946;
wire x_10947;
wire x_10948;
wire x_10949;
wire x_10950;
wire x_10951;
wire x_10952;
wire x_10953;
wire x_10954;
wire x_10955;
wire x_10956;
wire x_10957;
wire x_10958;
wire x_10959;
wire x_10960;
wire x_10961;
wire x_10962;
wire x_10963;
wire x_10964;
wire x_10965;
wire x_10966;
wire x_10967;
wire x_10968;
wire x_10969;
wire x_10970;
wire x_10971;
wire x_10972;
wire x_10973;
wire x_10974;
wire x_10975;
wire x_10976;
wire x_10977;
wire x_10978;
wire x_10979;
wire x_10980;
wire x_10981;
wire x_10982;
wire x_10983;
wire x_10984;
wire x_10985;
wire x_10986;
wire x_10987;
wire x_10988;
wire x_10989;
wire x_10990;
wire x_10991;
wire x_10992;
wire x_10993;
wire x_10994;
wire x_10995;
wire x_10996;
wire x_10997;
wire x_10998;
wire x_10999;
wire x_11000;
wire x_11001;
wire x_11002;
wire x_11003;
wire x_11004;
wire x_11005;
wire x_11006;
wire x_11007;
wire x_11008;
wire x_11009;
wire x_11010;
wire x_11011;
wire x_11012;
wire x_11013;
wire x_11014;
wire x_11015;
wire x_11016;
wire x_11017;
wire x_11018;
wire x_11019;
wire x_11020;
wire x_11021;
wire x_11022;
wire x_11023;
wire x_11024;
wire x_11025;
wire x_11026;
wire x_11027;
wire x_11028;
wire x_11029;
wire x_11030;
wire x_11031;
wire x_11032;
wire x_11033;
wire x_11034;
wire x_11035;
wire x_11036;
wire x_11037;
wire x_11038;
wire x_11039;
wire x_11040;
wire x_11041;
wire x_11042;
wire x_11043;
wire x_11044;
wire x_11045;
wire x_11046;
wire x_11047;
wire x_11048;
wire x_11049;
wire x_11050;
wire x_11051;
wire x_11052;
wire x_11053;
wire x_11054;
wire x_11055;
wire x_11056;
wire x_11057;
wire x_11058;
wire x_11059;
wire x_11060;
wire x_11061;
wire x_11062;
wire x_11063;
wire x_11064;
wire x_11065;
wire x_11066;
wire x_11067;
wire x_11068;
wire x_11069;
wire x_11070;
wire x_11071;
wire x_11072;
wire x_11073;
wire x_11074;
wire x_11075;
wire x_11076;
wire x_11077;
wire x_11078;
wire x_11079;
wire x_11080;
wire x_11081;
wire x_11082;
wire x_11083;
wire x_11084;
wire x_11085;
wire x_11086;
wire x_11087;
wire x_11088;
wire x_11089;
wire x_11090;
wire x_11091;
wire x_11092;
wire x_11093;
wire x_11094;
wire x_11095;
wire x_11096;
wire x_11097;
wire x_11098;
wire x_11099;
wire x_11100;
wire x_11101;
wire x_11102;
wire x_11103;
wire x_11104;
wire x_11105;
wire x_11106;
wire x_11107;
wire x_11108;
wire x_11109;
wire x_11110;
wire x_11111;
wire x_11112;
wire x_11113;
wire x_11114;
wire x_11115;
wire x_11116;
wire x_11117;
wire x_11118;
wire x_11119;
wire x_11120;
wire x_11121;
wire x_11122;
wire x_11123;
wire x_11124;
wire x_11125;
wire x_11126;
wire x_11127;
wire x_11128;
wire x_11129;
wire x_11130;
wire x_11131;
wire x_11132;
wire x_11133;
wire x_11134;
wire x_11135;
wire x_11136;
wire x_11137;
wire x_11138;
wire x_11139;
wire x_11140;
wire x_11141;
wire x_11142;
wire x_11143;
wire x_11144;
wire x_11145;
wire x_11146;
wire x_11147;
wire x_11148;
wire x_11149;
wire x_11150;
wire x_11151;
wire x_11152;
wire x_11153;
wire x_11154;
wire x_11155;
wire x_11156;
wire x_11157;
wire x_11158;
wire x_11159;
wire x_11160;
wire x_11161;
wire x_11162;
wire x_11163;
wire x_11164;
wire x_11165;
wire x_11166;
wire x_11167;
wire x_11168;
wire x_11169;
wire x_11170;
wire x_11171;
wire x_11172;
wire x_11173;
wire x_11174;
wire x_11175;
wire x_11176;
wire x_11177;
wire x_11178;
wire x_11179;
wire x_11180;
wire x_11181;
wire x_11182;
wire x_11183;
wire x_11184;
wire x_11185;
wire x_11186;
wire x_11187;
wire x_11188;
wire x_11189;
wire x_11190;
wire x_11191;
wire x_11192;
wire x_11193;
wire x_11194;
wire x_11195;
wire x_11196;
wire x_11197;
wire x_11198;
wire x_11199;
wire x_11200;
wire x_11201;
wire x_11202;
wire x_11203;
wire x_11204;
wire x_11205;
wire x_11206;
wire x_11207;
wire x_11208;
wire x_11209;
wire x_11210;
wire x_11211;
wire x_11212;
wire x_11213;
wire x_11214;
wire x_11215;
wire x_11216;
wire x_11217;
wire x_11218;
wire x_11219;
wire x_11220;
wire x_11221;
wire x_11222;
wire x_11223;
wire x_11224;
wire x_11225;
wire x_11226;
wire x_11227;
wire x_11228;
wire x_11229;
wire x_11230;
wire x_11231;
wire x_11232;
wire x_11233;
wire x_11234;
wire x_11235;
wire x_11236;
wire x_11237;
wire x_11238;
wire x_11239;
wire x_11240;
wire x_11241;
wire x_11242;
wire x_11243;
wire x_11244;
wire x_11245;
wire x_11246;
wire x_11247;
wire x_11248;
wire x_11249;
wire x_11250;
wire x_11251;
wire x_11252;
wire x_11253;
wire x_11254;
wire x_11255;
wire x_11256;
wire x_11257;
wire x_11258;
wire x_11259;
wire x_11260;
wire x_11261;
wire x_11262;
wire x_11263;
wire x_11264;
wire x_11265;
wire x_11266;
wire x_11267;
wire x_11268;
wire x_11269;
wire x_11270;
wire x_11271;
wire x_11272;
wire x_11273;
wire x_11274;
wire x_11275;
wire x_11276;
wire x_11277;
wire x_11278;
wire x_11279;
wire x_11280;
wire x_11281;
wire x_11282;
wire x_11283;
wire x_11284;
wire x_11285;
wire x_11286;
wire x_11287;
wire x_11288;
wire x_11289;
wire x_11290;
wire x_11291;
wire x_11292;
wire x_11293;
wire x_11294;
wire x_11295;
wire x_11296;
wire x_11297;
wire x_11298;
wire x_11299;
wire x_11300;
wire x_11301;
wire x_11302;
wire x_11303;
wire x_11304;
wire x_11305;
wire x_11306;
wire x_11307;
wire x_11308;
wire x_11309;
wire x_11310;
wire x_11311;
wire x_11312;
wire x_11313;
wire x_11314;
wire x_11315;
wire x_11316;
wire x_11317;
wire x_11318;
wire x_11319;
wire x_11320;
wire x_11321;
wire x_11322;
wire x_11323;
wire x_11324;
wire x_11325;
wire x_11326;
wire x_11327;
wire x_11328;
wire x_11329;
wire x_11330;
wire x_11331;
wire x_11332;
wire x_11333;
wire x_11334;
wire x_11335;
wire x_11336;
wire x_11337;
wire x_11338;
wire x_11339;
wire x_11340;
wire x_11341;
wire x_11342;
wire x_11343;
wire x_11344;
wire x_11345;
wire x_11346;
wire x_11347;
wire x_11348;
wire x_11349;
wire x_11350;
wire x_11351;
wire x_11352;
wire x_11353;
wire x_11354;
wire x_11355;
wire x_11356;
wire x_11357;
wire x_11358;
wire x_11359;
wire x_11360;
wire x_11361;
wire x_11362;
wire x_11363;
wire x_11364;
wire x_11365;
wire x_11366;
wire x_11367;
wire x_11368;
wire x_11369;
wire x_11370;
wire x_11371;
wire x_11372;
wire x_11373;
wire x_11374;
wire x_11375;
wire x_11376;
wire x_11377;
wire x_11378;
wire x_11379;
wire x_11380;
wire x_11381;
wire x_11382;
wire x_11383;
wire x_11384;
wire x_11385;
wire x_11386;
wire x_11387;
wire x_11388;
wire x_11389;
wire x_11390;
wire x_11391;
wire x_11392;
wire x_11393;
wire x_11394;
wire x_11395;
wire x_11396;
wire x_11397;
wire x_11398;
wire x_11399;
wire x_11400;
wire x_11401;
wire x_11402;
wire x_11403;
wire x_11404;
wire x_11405;
wire x_11406;
wire x_11407;
wire x_11408;
wire x_11409;
wire x_11410;
wire x_11411;
wire x_11412;
wire x_11413;
wire x_11414;
wire x_11415;
wire x_11416;
wire x_11417;
wire x_11418;
wire x_11419;
wire x_11420;
wire x_11421;
wire x_11422;
wire x_11423;
wire x_11424;
wire x_11425;
wire x_11426;
wire x_11427;
wire x_11428;
wire x_11429;
wire x_11430;
wire x_11431;
wire x_11432;
wire x_11433;
wire x_11434;
wire x_11435;
wire x_11436;
wire x_11437;
wire x_11438;
wire x_11439;
wire x_11440;
wire x_11441;
wire x_11442;
wire x_11443;
wire x_11444;
wire x_11445;
wire x_11446;
wire x_11447;
wire x_11448;
wire x_11449;
wire x_11450;
wire x_11451;
wire x_11452;
wire x_11453;
wire x_11454;
wire x_11455;
wire x_11456;
wire x_11457;
wire x_11458;
wire x_11459;
wire x_11460;
wire x_11461;
wire x_11462;
wire x_11463;
wire x_11464;
wire x_11465;
wire x_11466;
wire x_11467;
wire x_11468;
wire x_11469;
wire x_11470;
wire x_11471;
wire x_11472;
wire x_11473;
wire x_11474;
wire x_11475;
wire x_11476;
wire x_11477;
wire x_11478;
wire x_11479;
wire x_11480;
wire x_11481;
wire x_11482;
wire x_11483;
wire x_11484;
wire x_11485;
wire x_11486;
wire x_11487;
wire x_11488;
wire x_11489;
wire x_11490;
wire x_11491;
wire x_11492;
wire x_11493;
wire x_11494;
wire x_11495;
wire x_11496;
wire x_11497;
wire x_11498;
wire x_11499;
wire x_11500;
wire x_11501;
wire x_11502;
wire x_11503;
wire x_11504;
wire x_11505;
wire x_11506;
wire x_11507;
wire x_11508;
wire x_11509;
wire x_11510;
wire x_11511;
wire x_11512;
wire x_11513;
wire x_11514;
wire x_11515;
wire x_11516;
wire x_11517;
wire x_11518;
wire x_11519;
wire x_11520;
wire x_11521;
wire x_11522;
wire x_11523;
wire x_11524;
wire x_11525;
wire x_11526;
wire x_11527;
wire x_11528;
wire x_11529;
wire x_11530;
wire x_11531;
wire x_11532;
wire x_11533;
wire x_11534;
wire x_11535;
wire x_11536;
wire x_11537;
wire x_11538;
wire x_11539;
wire x_11540;
wire x_11541;
wire x_11542;
wire x_11543;
wire x_11544;
wire x_11545;
wire x_11546;
wire x_11547;
wire x_11548;
wire x_11549;
wire x_11550;
wire x_11551;
wire x_11552;
wire x_11553;
wire x_11554;
wire x_11555;
wire x_11556;
wire x_11557;
wire x_11558;
wire x_11559;
wire x_11560;
wire x_11561;
wire x_11562;
wire x_11563;
wire x_11564;
wire x_11565;
wire x_11566;
wire x_11567;
wire x_11568;
wire x_11569;
wire x_11570;
wire x_11571;
wire x_11572;
wire x_11573;
wire x_11574;
wire x_11575;
wire x_11576;
wire x_11577;
wire x_11578;
wire x_11579;
wire x_11580;
wire x_11581;
wire x_11582;
wire x_11583;
wire x_11584;
wire x_11585;
wire x_11586;
wire x_11587;
wire x_11588;
wire x_11589;
wire x_11590;
wire x_11591;
wire x_11592;
wire x_11593;
wire x_11594;
wire x_11595;
wire x_11596;
wire x_11597;
wire x_11598;
wire x_11599;
wire x_11600;
wire x_11601;
wire x_11602;
wire x_11603;
wire x_11604;
wire x_11605;
wire x_11606;
wire x_11607;
wire x_11608;
wire x_11609;
wire x_11610;
wire x_11611;
wire x_11612;
wire x_11613;
wire x_11614;
wire x_11615;
wire x_11616;
wire x_11617;
wire x_11618;
wire x_11619;
wire x_11620;
wire x_11621;
wire x_11622;
wire x_11623;
wire x_11624;
wire x_11625;
wire x_11626;
wire x_11627;
wire x_11628;
wire x_11629;
wire x_11630;
wire x_11631;
wire x_11632;
wire x_11633;
wire x_11634;
wire x_11635;
wire x_11636;
wire x_11637;
wire x_11638;
wire x_11639;
wire x_11640;
wire x_11641;
wire x_11642;
wire x_11643;
wire x_11644;
wire x_11645;
wire x_11646;
wire x_11647;
wire x_11648;
wire x_11649;
wire x_11650;
wire x_11651;
wire x_11652;
wire x_11653;
wire x_11654;
wire x_11655;
wire x_11656;
wire x_11657;
wire x_11658;
wire x_11659;
wire x_11660;
wire x_11661;
wire x_11662;
wire x_11663;
wire x_11664;
wire x_11665;
wire x_11666;
wire x_11667;
wire x_11668;
wire x_11669;
wire x_11670;
wire x_11671;
wire x_11672;
wire x_11673;
wire x_11674;
wire x_11675;
wire x_11676;
wire x_11677;
wire x_11678;
wire x_11679;
wire x_11680;
wire x_11681;
wire x_11682;
wire x_11683;
wire x_11684;
wire x_11685;
wire x_11686;
wire x_11687;
wire x_11688;
wire x_11689;
wire x_11690;
wire x_11691;
wire x_11692;
wire x_11693;
wire x_11694;
wire x_11695;
wire x_11696;
wire x_11697;
wire x_11698;
wire x_11699;
wire x_11700;
wire x_11701;
wire x_11702;
wire x_11703;
wire x_11704;
wire x_11705;
wire x_11706;
wire x_11707;
wire x_11708;
wire x_11709;
wire x_11710;
wire x_11711;
wire x_11712;
wire x_11713;
wire x_11714;
wire x_11715;
wire x_11716;
wire x_11717;
wire x_11718;
wire x_11719;
wire x_11720;
wire x_11721;
wire x_11722;
wire x_11723;
wire x_11724;
wire x_11725;
wire x_11726;
wire x_11727;
wire x_11728;
wire x_11729;
wire x_11730;
wire x_11731;
wire x_11732;
wire x_11733;
wire x_11734;
wire x_11735;
wire x_11736;
wire x_11737;
wire x_11738;
wire x_11739;
wire x_11740;
wire x_11741;
wire x_11742;
wire x_11743;
wire x_11744;
wire x_11745;
wire x_11746;
wire x_11747;
wire x_11748;
wire x_11749;
wire x_11750;
wire x_11751;
wire x_11752;
wire x_11753;
wire x_11754;
wire x_11755;
wire x_11756;
wire x_11757;
wire x_11758;
wire x_11759;
wire x_11760;
wire x_11761;
wire x_11762;
wire x_11763;
wire x_11764;
wire x_11765;
wire x_11766;
wire x_11767;
wire x_11768;
wire x_11769;
wire x_11770;
wire x_11771;
wire x_11772;
wire x_11773;
wire x_11774;
wire x_11775;
wire x_11776;
wire x_11777;
wire x_11778;
wire x_11779;
wire x_11780;
wire x_11781;
wire x_11782;
wire x_11783;
wire x_11784;
wire x_11785;
wire x_11786;
wire x_11787;
wire x_11788;
wire x_11789;
wire x_11790;
wire x_11791;
wire x_11792;
wire x_11793;
wire x_11794;
wire x_11795;
wire x_11796;
wire x_11797;
wire x_11798;
wire x_11799;
wire x_11800;
wire x_11801;
wire x_11802;
wire x_11803;
wire x_11804;
wire x_11805;
wire x_11806;
wire x_11807;
wire x_11808;
wire x_11809;
wire x_11810;
wire x_11811;
wire x_11812;
wire x_11813;
wire x_11814;
wire x_11815;
wire x_11816;
wire x_11817;
wire x_11818;
wire x_11819;
wire x_11820;
wire x_11821;
wire x_11822;
wire x_11823;
wire x_11824;
wire x_11825;
wire x_11826;
wire x_11827;
wire x_11828;
wire x_11829;
wire x_11830;
wire x_11831;
wire x_11832;
wire x_11833;
wire x_11834;
wire x_11835;
wire x_11836;
wire x_11837;
wire x_11838;
wire x_11839;
wire x_11840;
wire x_11841;
wire x_11842;
wire x_11843;
wire x_11844;
wire x_11845;
wire x_11846;
wire x_11847;
wire x_11848;
wire x_11849;
wire x_11850;
wire x_11851;
wire x_11852;
wire x_11853;
wire x_11854;
wire x_11855;
wire x_11856;
wire x_11857;
wire x_11858;
wire x_11859;
wire x_11860;
wire x_11861;
wire x_11862;
wire x_11863;
wire x_11864;
wire x_11865;
wire x_11866;
wire x_11867;
wire x_11868;
wire x_11869;
wire x_11870;
wire x_11871;
wire x_11872;
wire x_11873;
wire x_11874;
wire x_11875;
wire x_11876;
wire x_11877;
wire x_11878;
wire x_11879;
wire x_11880;
wire x_11881;
wire x_11882;
wire x_11883;
wire x_11884;
wire x_11885;
wire x_11886;
wire x_11887;
wire x_11888;
wire x_11889;
wire x_11890;
wire x_11891;
wire x_11892;
wire x_11893;
wire x_11894;
wire x_11895;
wire x_11896;
wire x_11897;
wire x_11898;
wire x_11899;
wire x_11900;
wire x_11901;
wire x_11902;
wire x_11903;
wire x_11904;
wire x_11905;
wire x_11906;
wire x_11907;
wire x_11908;
wire x_11909;
wire x_11910;
wire x_11911;
wire x_11912;
wire x_11913;
wire x_11914;
wire x_11915;
wire x_11916;
wire x_11917;
wire x_11918;
wire x_11919;
wire x_11920;
wire x_11921;
wire x_11922;
wire x_11923;
wire x_11924;
wire x_11925;
wire x_11926;
wire x_11927;
wire x_11928;
wire x_11929;
wire x_11930;
wire x_11931;
wire x_11932;
wire x_11933;
wire x_11934;
wire x_11935;
wire x_11936;
wire x_11937;
wire x_11938;
wire x_11939;
wire x_11940;
wire x_11941;
wire x_11942;
wire x_11943;
wire x_11944;
wire x_11945;
wire x_11946;
wire x_11947;
wire x_11948;
wire x_11949;
wire x_11950;
wire x_11951;
wire x_11952;
wire x_11953;
wire x_11954;
wire x_11955;
wire x_11956;
wire x_11957;
wire x_11958;
wire x_11959;
wire x_11960;
wire x_11961;
wire x_11962;
wire x_11963;
wire x_11964;
wire x_11965;
wire x_11966;
wire x_11967;
wire x_11968;
wire x_11969;
wire x_11970;
wire x_11971;
wire x_11972;
wire x_11973;
wire x_11974;
wire x_11975;
wire x_11976;
wire x_11977;
wire x_11978;
wire x_11979;
wire x_11980;
wire x_11981;
wire x_11982;
wire x_11983;
wire x_11984;
wire x_11985;
wire x_11986;
wire x_11987;
wire x_11988;
wire x_11989;
wire x_11990;
wire x_11991;
wire x_11992;
wire x_11993;
wire x_11994;
wire x_11995;
wire x_11996;
wire x_11997;
wire x_11998;
wire x_11999;
wire x_12000;
wire x_12001;
wire x_12002;
wire x_12003;
wire x_12004;
wire x_12005;
wire x_12006;
wire x_12007;
wire x_12008;
wire x_12009;
wire x_12010;
wire x_12011;
wire x_12012;
wire x_12013;
wire x_12014;
wire x_12015;
wire x_12016;
wire x_12017;
wire x_12018;
wire x_12019;
wire x_12020;
wire x_12021;
wire x_12022;
wire x_12023;
wire x_12024;
wire x_12025;
wire x_12026;
wire x_12027;
wire x_12028;
wire x_12029;
wire x_12030;
wire x_12031;
wire x_12032;
wire x_12033;
wire x_12034;
wire x_12035;
wire x_12036;
wire x_12037;
wire x_12038;
wire x_12039;
wire x_12040;
wire x_12041;
wire x_12042;
wire x_12043;
wire x_12044;
wire x_12045;
wire x_12046;
wire x_12047;
wire x_12048;
wire x_12049;
wire x_12050;
wire x_12051;
wire x_12052;
wire x_12053;
wire x_12054;
wire x_12055;
wire x_12056;
wire x_12057;
wire x_12058;
wire x_12059;
wire x_12060;
wire x_12061;
wire x_12062;
wire x_12063;
wire x_12064;
wire x_12065;
wire x_12066;
wire x_12067;
wire x_12068;
wire x_12069;
wire x_12070;
wire x_12071;
wire x_12072;
wire x_12073;
wire x_12074;
wire x_12075;
wire x_12076;
wire x_12077;
wire x_12078;
wire x_12079;
wire x_12080;
wire x_12081;
wire x_12082;
wire x_12083;
wire x_12084;
wire x_12085;
wire x_12086;
wire x_12087;
wire x_12088;
wire x_12089;
wire x_12090;
wire x_12091;
wire x_12092;
wire x_12093;
wire x_12094;
wire x_12095;
wire x_12096;
wire x_12097;
wire x_12098;
wire x_12099;
wire x_12100;
wire x_12101;
wire x_12102;
wire x_12103;
wire x_12104;
wire x_12105;
wire x_12106;
wire x_12107;
wire x_12108;
wire x_12109;
wire x_12110;
wire x_12111;
wire x_12112;
wire x_12113;
wire x_12114;
wire x_12115;
wire x_12116;
wire x_12117;
wire x_12118;
wire x_12119;
wire x_12120;
wire x_12121;
wire x_12122;
wire x_12123;
wire x_12124;
wire x_12125;
wire x_12126;
wire x_12127;
wire x_12128;
wire x_12129;
wire x_12130;
wire x_12131;
wire x_12132;
wire x_12133;
wire x_12134;
wire x_12135;
wire x_12136;
wire x_12137;
wire x_12138;
wire x_12139;
wire x_12140;
wire x_12141;
wire x_12142;
wire x_12143;
wire x_12144;
wire x_12145;
wire x_12146;
wire x_12147;
wire x_12148;
wire x_12149;
wire x_12150;
wire x_12151;
wire x_12152;
wire x_12153;
wire x_12154;
wire x_12155;
wire x_12156;
wire x_12157;
wire x_12158;
wire x_12159;
wire x_12160;
wire x_12161;
wire x_12162;
wire x_12163;
wire x_12164;
wire x_12165;
wire x_12166;
wire x_12167;
wire x_12168;
wire x_12169;
wire x_12170;
wire x_12171;
wire x_12172;
wire x_12173;
wire x_12174;
wire x_12175;
wire x_12176;
wire x_12177;
wire x_12178;
wire x_12179;
wire x_12180;
wire x_12181;
wire x_12182;
wire x_12183;
wire x_12184;
wire x_12185;
wire x_12186;
wire x_12187;
wire x_12188;
wire x_12189;
wire x_12190;
wire x_12191;
wire x_12192;
wire x_12193;
wire x_12194;
wire x_12195;
wire x_12196;
wire x_12197;
wire x_12198;
wire x_12199;
wire x_12200;
wire x_12201;
wire x_12202;
wire x_12203;
wire x_12204;
wire x_12205;
wire x_12206;
wire x_12207;
wire x_12208;
wire x_12209;
wire x_12210;
wire x_12211;
wire x_12212;
wire x_12213;
wire x_12214;
wire x_12215;
wire x_12216;
wire x_12217;
wire x_12218;
wire x_12219;
wire x_12220;
wire x_12221;
wire x_12222;
wire x_12223;
wire x_12224;
wire x_12225;
wire x_12226;
wire x_12227;
wire x_12228;
wire x_12229;
wire x_12230;
wire x_12231;
wire x_12232;
wire x_12233;
wire x_12234;
wire x_12235;
wire x_12236;
wire x_12237;
wire x_12238;
wire x_12239;
wire x_12240;
wire x_12241;
wire x_12242;
wire x_12243;
wire x_12244;
wire x_12245;
wire x_12246;
wire x_12247;
wire x_12248;
wire x_12249;
wire x_12250;
wire x_12251;
wire x_12252;
wire x_12253;
wire x_12254;
wire x_12255;
wire x_12256;
wire x_12257;
wire x_12258;
wire x_12259;
wire x_12260;
wire x_12261;
wire x_12262;
wire x_12263;
wire x_12264;
wire x_12265;
wire x_12266;
wire x_12267;
wire x_12268;
wire x_12269;
wire x_12270;
wire x_12271;
wire x_12272;
wire x_12273;
wire x_12274;
wire x_12275;
wire x_12276;
wire x_12277;
wire x_12278;
wire x_12279;
wire x_12280;
wire x_12281;
wire x_12282;
wire x_12283;
wire x_12284;
wire x_12285;
wire x_12286;
wire x_12287;
wire x_12288;
wire x_12289;
wire x_12290;
wire x_12291;
wire x_12292;
wire x_12293;
wire x_12294;
wire x_12295;
wire x_12296;
wire x_12297;
wire x_12298;
wire x_12299;
wire x_12300;
wire x_12301;
wire x_12302;
wire x_12303;
wire x_12304;
wire x_12305;
wire x_12306;
wire x_12307;
wire x_12308;
wire x_12309;
wire x_12310;
wire x_12311;
wire x_12312;
wire x_12313;
wire x_12314;
wire x_12315;
wire x_12316;
wire x_12317;
wire x_12318;
wire x_12319;
wire x_12320;
wire x_12321;
wire x_12322;
wire x_12323;
wire x_12324;
wire x_12325;
wire x_12326;
wire x_12327;
wire x_12328;
wire x_12329;
wire x_12330;
wire x_12331;
wire x_12332;
wire x_12333;
wire x_12334;
wire x_12335;
wire x_12336;
wire x_12337;
wire x_12338;
wire x_12339;
wire x_12340;
wire x_12341;
wire x_12342;
wire x_12343;
wire x_12344;
wire x_12345;
wire x_12346;
wire x_12347;
wire x_12348;
wire x_12349;
wire x_12350;
wire x_12351;
wire x_12352;
wire x_12353;
wire x_12354;
wire x_12355;
wire x_12356;
wire x_12357;
wire x_12358;
wire x_12359;
wire x_12360;
wire x_12361;
wire x_12362;
wire x_12363;
wire x_12364;
wire x_12365;
wire x_12366;
wire x_12367;
wire x_12368;
wire x_12369;
wire x_12370;
wire x_12371;
wire x_12372;
wire x_12373;
wire x_12374;
wire x_12375;
wire x_12376;
wire x_12377;
wire x_12378;
wire x_12379;
wire x_12380;
wire x_12381;
wire x_12382;
wire x_12383;
wire x_12384;
wire x_12385;
wire x_12386;
wire x_12387;
wire x_12388;
wire x_12389;
wire x_12390;
wire x_12391;
wire x_12392;
wire x_12393;
wire x_12394;
wire x_12395;
wire x_12396;
wire x_12397;
wire x_12398;
wire x_12399;
wire x_12400;
wire x_12401;
wire x_12402;
wire x_12403;
wire x_12404;
wire x_12405;
wire x_12406;
wire x_12407;
wire x_12408;
wire x_12409;
wire x_12410;
wire x_12411;
wire x_12412;
wire x_12413;
wire x_12414;
wire x_12415;
wire x_12416;
wire x_12417;
wire x_12418;
wire x_12419;
wire x_12420;
wire x_12421;
wire x_12422;
wire x_12423;
wire x_12424;
wire x_12425;
wire x_12426;
wire x_12427;
wire x_12428;
wire x_12429;
wire x_12430;
wire x_12431;
wire x_12432;
wire x_12433;
wire x_12434;
wire x_12435;
wire x_12436;
wire x_12437;
wire x_12438;
wire x_12439;
wire x_12440;
wire x_12441;
wire x_12442;
wire x_12443;
wire x_12444;
wire x_12445;
wire x_12446;
wire x_12447;
wire x_12448;
wire x_12449;
wire x_12450;
wire x_12451;
wire x_12452;
wire x_12453;
wire x_12454;
wire x_12455;
wire x_12456;
wire x_12457;
wire x_12458;
wire x_12459;
wire x_12460;
wire x_12461;
wire x_12462;
wire x_12463;
wire x_12464;
wire x_12465;
wire x_12466;
wire x_12467;
wire x_12468;
wire x_12469;
wire x_12470;
wire x_12471;
wire x_12472;
wire x_12473;
wire x_12474;
wire x_12475;
wire x_12476;
wire x_12477;
wire x_12478;
wire x_12479;
wire x_12480;
wire x_12481;
wire x_12482;
wire x_12483;
wire x_12484;
wire x_12485;
wire x_12486;
wire x_12487;
wire x_12488;
wire x_12489;
wire x_12490;
wire x_12491;
wire x_12492;
wire x_12493;
wire x_12494;
wire x_12495;
wire x_12496;
wire x_12497;
wire x_12498;
wire x_12499;
wire x_12500;
wire x_12501;
wire x_12502;
wire x_12503;
wire x_12504;
wire x_12505;
wire x_12506;
wire x_12507;
wire x_12508;
wire x_12509;
wire x_12510;
wire x_12511;
wire x_12512;
wire x_12513;
wire x_12514;
wire x_12515;
wire x_12516;
wire x_12517;
wire x_12518;
wire x_12519;
wire x_12520;
wire x_12521;
wire x_12522;
wire x_12523;
wire x_12524;
wire x_12525;
wire x_12526;
wire x_12527;
wire x_12528;
wire x_12529;
wire x_12530;
wire x_12531;
wire x_12532;
wire x_12533;
wire x_12534;
wire x_12535;
wire x_12536;
wire x_12537;
wire x_12538;
wire x_12539;
wire x_12540;
wire x_12541;
wire x_12542;
wire x_12543;
wire x_12544;
wire x_12545;
wire x_12546;
wire x_12547;
wire x_12548;
wire x_12549;
wire x_12550;
wire x_12551;
wire x_12552;
wire x_12553;
wire x_12554;
wire x_12555;
wire x_12556;
wire x_12557;
wire x_12558;
wire x_12559;
wire x_12560;
wire x_12561;
wire x_12562;
wire x_12563;
wire x_12564;
wire x_12565;
wire x_12566;
wire x_12567;
wire x_12568;
wire x_12569;
wire x_12570;
wire x_12571;
wire x_12572;
wire x_12573;
wire x_12574;
wire x_12575;
wire x_12576;
wire x_12577;
wire x_12578;
wire x_12579;
wire x_12580;
wire x_12581;
wire x_12582;
wire x_12583;
wire x_12584;
wire x_12585;
wire x_12586;
wire x_12587;
wire x_12588;
wire x_12589;
wire x_12590;
wire x_12591;
wire x_12592;
wire x_12593;
wire x_12594;
wire x_12595;
wire x_12596;
wire x_12597;
wire x_12598;
wire x_12599;
wire x_12600;
wire x_12601;
wire x_12602;
wire x_12603;
wire x_12604;
wire x_12605;
wire x_12606;
wire x_12607;
wire x_12608;
wire x_12609;
wire x_12610;
wire x_12611;
wire x_12612;
wire x_12613;
wire x_12614;
wire x_12615;
wire x_12616;
wire x_12617;
wire x_12618;
wire x_12619;
wire x_12620;
wire x_12621;
wire x_12622;
wire x_12623;
wire x_12624;
wire x_12625;
wire x_12626;
wire x_12627;
wire x_12628;
wire x_12629;
wire x_12630;
wire x_12631;
wire x_12632;
wire x_12633;
wire x_12634;
wire x_12635;
wire x_12636;
wire x_12637;
wire x_12638;
wire x_12639;
wire x_12640;
wire x_12641;
wire x_12642;
wire x_12643;
wire x_12644;
wire x_12645;
wire x_12646;
wire x_12647;
wire x_12648;
wire x_12649;
wire x_12650;
wire x_12651;
wire x_12652;
wire x_12653;
wire x_12654;
wire x_12655;
wire x_12656;
wire x_12657;
wire x_12658;
wire x_12659;
wire x_12660;
wire x_12661;
wire x_12662;
wire x_12663;
wire x_12664;
wire x_12665;
wire x_12666;
wire x_12667;
wire x_12668;
wire x_12669;
wire x_12670;
wire x_12671;
wire x_12672;
wire x_12673;
wire x_12674;
wire x_12675;
wire x_12676;
wire x_12677;
wire x_12678;
wire x_12679;
wire x_12680;
wire x_12681;
wire x_12682;
wire x_12683;
wire x_12684;
wire x_12685;
wire x_12686;
wire x_12687;
wire x_12688;
wire x_12689;
wire x_12690;
wire x_12691;
wire x_12692;
wire x_12693;
wire x_12694;
wire x_12695;
wire x_12696;
wire x_12697;
wire x_12698;
wire x_12699;
wire x_12700;
wire x_12701;
wire x_12702;
wire x_12703;
wire x_12704;
wire x_12705;
wire x_12706;
wire x_12707;
wire x_12708;
wire x_12709;
wire x_12710;
wire x_12711;
wire x_12712;
wire x_12713;
wire x_12714;
wire x_12715;
wire x_12716;
wire x_12717;
wire x_12718;
wire x_12719;
wire x_12720;
wire x_12721;
wire x_12722;
wire x_12723;
wire x_12724;
wire x_12725;
wire x_12726;
wire x_12727;
wire x_12728;
wire x_12729;
wire x_12730;
wire x_12731;
wire x_12732;
wire x_12733;
wire x_12734;
wire x_12735;
wire x_12736;
wire x_12737;
wire x_12738;
wire x_12739;
wire x_12740;
wire x_12741;
wire x_12742;
wire x_12743;
wire x_12744;
wire x_12745;
wire x_12746;
wire x_12747;
wire x_12748;
wire x_12749;
wire x_12750;
wire x_12751;
wire x_12752;
wire x_12753;
wire x_12754;
wire x_12755;
wire x_12756;
wire x_12757;
wire x_12758;
wire x_12759;
wire x_12760;
wire x_12761;
wire x_12762;
wire x_12763;
wire x_12764;
wire x_12765;
wire x_12766;
wire x_12767;
wire x_12768;
wire x_12769;
wire x_12770;
wire x_12771;
wire x_12772;
wire x_12773;
wire x_12774;
wire x_12775;
wire x_12776;
wire x_12777;
wire x_12778;
wire x_12779;
wire x_12780;
wire x_12781;
wire x_12782;
wire x_12783;
wire x_12784;
wire x_12785;
wire x_12786;
wire x_12787;
wire x_12788;
wire x_12789;
wire x_12790;
wire x_12791;
wire x_12792;
wire x_12793;
wire x_12794;
wire x_12795;
wire x_12796;
wire x_12797;
wire x_12798;
wire x_12799;
wire x_12800;
wire x_12801;
wire x_12802;
wire x_12803;
wire x_12804;
wire x_12805;
wire x_12806;
wire x_12807;
wire x_12808;
wire x_12809;
wire x_12810;
wire x_12811;
wire x_12812;
wire x_12813;
wire x_12814;
wire x_12815;
wire x_12816;
wire x_12817;
wire x_12818;
wire x_12819;
wire x_12820;
wire x_12821;
wire x_12822;
wire x_12823;
wire x_12824;
wire x_12825;
wire x_12826;
wire x_12827;
wire x_12828;
wire x_12829;
wire x_12830;
wire x_12831;
wire x_12832;
wire x_12833;
wire x_12834;
wire x_12835;
wire x_12836;
wire x_12837;
wire x_12838;
wire x_12839;
wire x_12840;
wire x_12841;
wire x_12842;
wire x_12843;
wire x_12844;
wire x_12845;
wire x_12846;
wire x_12847;
wire x_12848;
wire x_12849;
wire x_12850;
wire x_12851;
wire x_12852;
wire x_12853;
wire x_12854;
wire x_12855;
wire x_12856;
wire x_12857;
wire x_12858;
wire x_12859;
wire x_12860;
wire x_12861;
wire x_12862;
wire x_12863;
wire x_12864;
wire x_12865;
wire x_12866;
wire x_12867;
wire x_12868;
wire x_12869;
wire x_12870;
wire x_12871;
wire x_12872;
wire x_12873;
wire x_12874;
wire x_12875;
wire x_12876;
wire x_12877;
wire x_12878;
wire x_12879;
wire x_12880;
wire x_12881;
wire x_12882;
wire x_12883;
wire x_12884;
wire x_12885;
wire x_12886;
wire x_12887;
wire x_12888;
wire x_12889;
wire x_12890;
wire x_12891;
wire x_12892;
wire x_12893;
wire x_12894;
wire x_12895;
wire x_12896;
wire x_12897;
wire x_12898;
wire x_12899;
wire x_12900;
wire x_12901;
wire x_12902;
wire x_12903;
wire x_12904;
wire x_12905;
wire x_12906;
wire x_12907;
wire x_12908;
wire x_12909;
wire x_12910;
wire x_12911;
wire x_12912;
wire x_12913;
wire x_12914;
wire x_12915;
wire x_12916;
wire x_12917;
wire x_12918;
wire x_12919;
wire x_12920;
wire x_12921;
wire x_12922;
wire x_12923;
wire x_12924;
wire x_12925;
wire x_12926;
wire x_12927;
wire x_12928;
wire x_12929;
wire x_12930;
wire x_12931;
wire x_12932;
wire x_12933;
wire x_12934;
wire x_12935;
wire x_12936;
wire x_12937;
wire x_12938;
wire x_12939;
wire x_12940;
wire x_12941;
wire x_12942;
wire x_12943;
wire x_12944;
wire x_12945;
wire x_12946;
wire x_12947;
wire x_12948;
wire x_12949;
wire x_12950;
wire x_12951;
wire x_12952;
wire x_12953;
wire x_12954;
wire x_12955;
wire x_12956;
wire x_12957;
wire x_12958;
wire x_12959;
wire x_12960;
wire x_12961;
wire x_12962;
wire x_12963;
wire x_12964;
wire x_12965;
wire x_12966;
wire x_12967;
wire x_12968;
wire x_12969;
wire x_12970;
wire x_12971;
wire x_12972;
wire x_12973;
wire x_12974;
wire x_12975;
wire x_12976;
wire x_12977;
wire x_12978;
wire x_12979;
wire x_12980;
wire x_12981;
wire x_12982;
wire x_12983;
wire x_12984;
wire x_12985;
wire x_12986;
wire x_12987;
wire x_12988;
wire x_12989;
wire x_12990;
wire x_12991;
wire x_12992;
wire x_12993;
wire x_12994;
wire x_12995;
wire x_12996;
wire x_12997;
wire x_12998;
wire x_12999;
wire x_13000;
wire x_13001;
wire x_13002;
wire x_13003;
wire x_13004;
wire x_13005;
wire x_13006;
wire x_13007;
wire x_13008;
wire x_13009;
wire x_13010;
wire x_13011;
wire x_13012;
wire x_13013;
wire x_13014;
wire x_13015;
wire x_13016;
wire x_13017;
wire x_13018;
wire x_13019;
wire x_13020;
wire x_13021;
wire x_13022;
wire x_13023;
wire x_13024;
wire x_13025;
wire x_13026;
wire x_13027;
wire x_13028;
wire x_13029;
wire x_13030;
wire x_13031;
wire x_13032;
wire x_13033;
wire x_13034;
wire x_13035;
wire x_13036;
wire x_13037;
wire x_13038;
wire x_13039;
wire x_13040;
wire x_13041;
wire x_13042;
wire x_13043;
wire x_13044;
wire x_13045;
wire x_13046;
wire x_13047;
wire x_13048;
wire x_13049;
wire x_13050;
wire x_13051;
wire x_13052;
wire x_13053;
wire x_13054;
wire x_13055;
wire x_13056;
wire x_13057;
wire x_13058;
wire x_13059;
wire x_13060;
wire x_13061;
wire x_13062;
wire x_13063;
wire x_13064;
wire x_13065;
wire x_13066;
wire x_13067;
wire x_13068;
wire x_13069;
wire x_13070;
wire x_13071;
wire x_13072;
wire x_13073;
wire x_13074;
wire x_13075;
wire x_13076;
wire x_13077;
wire x_13078;
wire x_13079;
wire x_13080;
wire x_13081;
wire x_13082;
wire x_13083;
wire x_13084;
wire x_13085;
wire x_13086;
wire x_13087;
wire x_13088;
wire x_13089;
wire x_13090;
wire x_13091;
wire x_13092;
wire x_13093;
wire x_13094;
wire x_13095;
wire x_13096;
wire x_13097;
wire x_13098;
wire x_13099;
wire x_13100;
wire x_13101;
wire x_13102;
wire x_13103;
wire x_13104;
wire x_13105;
wire x_13106;
wire x_13107;
wire x_13108;
wire x_13109;
wire x_13110;
wire x_13111;
wire x_13112;
wire x_13113;
wire x_13114;
wire x_13115;
wire x_13116;
wire x_13117;
wire x_13118;
wire x_13119;
wire x_13120;
wire x_13121;
wire x_13122;
wire x_13123;
wire x_13124;
wire x_13125;
wire x_13126;
wire x_13127;
wire x_13128;
wire x_13129;
wire x_13130;
wire x_13131;
wire x_13132;
wire x_13133;
wire x_13134;
wire x_13135;
wire x_13136;
wire x_13137;
wire x_13138;
wire x_13139;
wire x_13140;
wire x_13141;
wire x_13142;
wire x_13143;
wire x_13144;
wire x_13145;
wire x_13146;
wire x_13147;
wire x_13148;
wire x_13149;
wire x_13150;
wire x_13151;
wire x_13152;
wire x_13153;
wire x_13154;
wire x_13155;
wire x_13156;
wire x_13157;
wire x_13158;
wire x_13159;
wire x_13160;
wire x_13161;
wire x_13162;
wire x_13163;
wire x_13164;
wire x_13165;
wire x_13166;
wire x_13167;
wire x_13168;
wire x_13169;
wire x_13170;
wire x_13171;
wire x_13172;
wire x_13173;
wire x_13174;
wire x_13175;
wire x_13176;
wire x_13177;
wire x_13178;
wire x_13179;
wire x_13180;
wire x_13181;
wire x_13182;
wire x_13183;
wire x_13184;
wire x_13185;
wire x_13186;
wire x_13187;
wire x_13188;
wire x_13189;
wire x_13190;
wire x_13191;
wire x_13192;
wire x_13193;
wire x_13194;
wire x_13195;
wire x_13196;
wire x_13197;
wire x_13198;
wire x_13199;
wire x_13200;
wire x_13201;
wire x_13202;
wire x_13203;
wire x_13204;
wire x_13205;
wire x_13206;
wire x_13207;
wire x_13208;
wire x_13209;
wire x_13210;
wire x_13211;
wire x_13212;
wire x_13213;
wire x_13214;
wire x_13215;
wire x_13216;
wire x_13217;
wire x_13218;
wire x_13219;
wire x_13220;
wire x_13221;
wire x_13222;
wire x_13223;
wire x_13224;
wire x_13225;
wire x_13226;
wire x_13227;
wire x_13228;
wire x_13229;
wire x_13230;
wire x_13231;
wire x_13232;
wire x_13233;
wire x_13234;
wire x_13235;
wire x_13236;
wire x_13237;
wire x_13238;
wire x_13239;
wire x_13240;
wire x_13241;
wire x_13242;
wire x_13243;
wire x_13244;
wire x_13245;
wire x_13246;
wire x_13247;
wire x_13248;
wire x_13249;
wire x_13250;
wire x_13251;
wire x_13252;
wire x_13253;
wire x_13254;
wire x_13255;
wire x_13256;
wire x_13257;
wire x_13258;
wire x_13259;
wire x_13260;
wire x_13261;
wire x_13262;
wire x_13263;
wire x_13264;
wire x_13265;
wire x_13266;
wire x_13267;
wire x_13268;
wire x_13269;
wire x_13270;
wire x_13271;
wire x_13272;
wire x_13273;
wire x_13274;
wire x_13275;
wire x_13276;
wire x_13277;
wire x_13278;
wire x_13279;
wire x_13280;
wire x_13281;
wire x_13282;
wire x_13283;
wire x_13284;
wire x_13285;
wire x_13286;
wire x_13287;
wire x_13288;
wire x_13289;
wire x_13290;
wire x_13291;
wire x_13292;
wire x_13293;
wire x_13294;
wire x_13295;
wire x_13296;
wire x_13297;
wire x_13298;
wire x_13299;
wire x_13300;
wire x_13301;
wire x_13302;
wire x_13303;
wire x_13304;
wire x_13305;
wire x_13306;
wire x_13307;
wire x_13308;
wire x_13309;
wire x_13310;
wire x_13311;
wire x_13312;
wire x_13313;
wire x_13314;
wire x_13315;
wire x_13316;
wire x_13317;
wire x_13318;
wire x_13319;
wire x_13320;
wire x_13321;
wire x_13322;
wire x_13323;
wire x_13324;
wire x_13325;
wire x_13326;
wire x_13327;
wire x_13328;
wire x_13329;
wire x_13330;
wire x_13331;
wire x_13332;
wire x_13333;
wire x_13334;
wire x_13335;
wire x_13336;
wire x_13337;
wire x_13338;
wire x_13339;
wire x_13340;
wire x_13341;
wire x_13342;
wire x_13343;
wire x_13344;
wire x_13345;
wire x_13346;
wire x_13347;
wire x_13348;
wire x_13349;
wire x_13350;
wire x_13351;
wire x_13352;
wire x_13353;
wire x_13354;
wire x_13355;
wire x_13356;
wire x_13357;
wire x_13358;
wire x_13359;
wire x_13360;
wire x_13361;
wire x_13362;
wire x_13363;
wire x_13364;
wire x_13365;
wire x_13366;
wire x_13367;
wire x_13368;
wire x_13369;
wire x_13370;
wire x_13371;
wire x_13372;
wire x_13373;
wire x_13374;
wire x_13375;
wire x_13376;
wire x_13377;
wire x_13378;
wire x_13379;
wire x_13380;
wire x_13381;
wire x_13382;
wire x_13383;
wire x_13384;
wire x_13385;
wire x_13386;
wire x_13387;
wire x_13388;
wire x_13389;
wire x_13390;
wire x_13391;
wire x_13392;
wire x_13393;
wire x_13394;
wire x_13395;
wire x_13396;
wire x_13397;
wire x_13398;
wire x_13399;
wire x_13400;
wire x_13401;
wire x_13402;
wire x_13403;
wire x_13404;
wire x_13405;
wire x_13406;
wire x_13407;
wire x_13408;
wire x_13409;
wire x_13410;
wire x_13411;
wire x_13412;
wire x_13413;
wire x_13414;
wire x_13415;
wire x_13416;
wire x_13417;
wire x_13418;
wire x_13419;
wire x_13420;
wire x_13421;
wire x_13422;
wire x_13423;
wire x_13424;
wire x_13425;
wire x_13426;
wire x_13427;
wire x_13428;
wire x_13429;
wire x_13430;
wire x_13431;
wire x_13432;
wire x_13433;
wire x_13434;
wire x_13435;
wire x_13436;
wire x_13437;
wire x_13438;
wire x_13439;
wire x_13440;
wire x_13441;
wire x_13442;
wire x_13443;
wire x_13444;
wire x_13445;
wire x_13446;
wire x_13447;
wire x_13448;
wire x_13449;
wire x_13450;
wire x_13451;
wire x_13452;
wire x_13453;
wire x_13454;
wire x_13455;
wire x_13456;
wire x_13457;
wire x_13458;
wire x_13459;
wire x_13460;
wire x_13461;
wire x_13462;
wire x_13463;
wire x_13464;
wire x_13465;
wire x_13466;
wire x_13467;
wire x_13468;
wire x_13469;
wire x_13470;
wire x_13471;
wire x_13472;
wire x_13473;
wire x_13474;
wire x_13475;
wire x_13476;
wire x_13477;
wire x_13478;
wire x_13479;
wire x_13480;
wire x_13481;
wire x_13482;
wire x_13483;
wire x_13484;
wire x_13485;
wire x_13486;
wire x_13487;
wire x_13488;
wire x_13489;
wire x_13490;
wire x_13491;
wire x_13492;
wire x_13493;
wire x_13494;
wire x_13495;
wire x_13496;
wire x_13497;
wire x_13498;
wire x_13499;
wire x_13500;
wire x_13501;
wire x_13502;
wire x_13503;
wire x_13504;
wire x_13505;
wire x_13506;
wire x_13507;
wire x_13508;
wire x_13509;
wire x_13510;
wire x_13511;
wire x_13512;
wire x_13513;
wire x_13514;
wire x_13515;
wire x_13516;
wire x_13517;
wire x_13518;
wire x_13519;
wire x_13520;
wire x_13521;
wire x_13522;
wire x_13523;
wire x_13524;
wire x_13525;
wire x_13526;
wire x_13527;
wire x_13528;
wire x_13529;
wire x_13530;
wire x_13531;
wire x_13532;
wire x_13533;
wire x_13534;
wire x_13535;
wire x_13536;
wire x_13537;
wire x_13538;
wire x_13539;
wire x_13540;
wire x_13541;
wire x_13542;
wire x_13543;
wire x_13544;
wire x_13545;
wire x_13546;
wire x_13547;
wire x_13548;
wire x_13549;
wire x_13550;
wire x_13551;
wire x_13552;
wire x_13553;
wire x_13554;
wire x_13555;
wire x_13556;
wire x_13557;
wire x_13558;
wire x_13559;
wire x_13560;
wire x_13561;
wire x_13562;
wire x_13563;
wire x_13564;
wire x_13565;
wire x_13566;
wire x_13567;
wire x_13568;
wire x_13569;
wire x_13570;
wire x_13571;
wire x_13572;
wire x_13573;
wire x_13574;
wire x_13575;
wire x_13576;
wire x_13577;
wire x_13578;
wire x_13579;
wire x_13580;
wire x_13581;
wire x_13582;
wire x_13583;
wire x_13584;
wire x_13585;
wire x_13586;
wire x_13587;
wire x_13588;
wire x_13589;
wire x_13590;
wire x_13591;
wire x_13592;
wire x_13593;
wire x_13594;
wire x_13595;
wire x_13596;
wire x_13597;
wire x_13598;
wire x_13599;
wire x_13600;
wire x_13601;
wire x_13602;
wire x_13603;
wire x_13604;
wire x_13605;
wire x_13606;
wire x_13607;
wire x_13608;
wire x_13609;
wire x_13610;
wire x_13611;
wire x_13612;
wire x_13613;
wire x_13614;
wire x_13615;
wire x_13616;
wire x_13617;
wire x_13618;
wire x_13619;
wire x_13620;
wire x_13621;
wire x_13622;
wire x_13623;
wire x_13624;
wire x_13625;
wire x_13626;
wire x_13627;
wire x_13628;
wire x_13629;
wire x_13630;
wire x_13631;
wire x_13632;
wire x_13633;
wire x_13634;
wire x_13635;
wire x_13636;
wire x_13637;
wire x_13638;
wire x_13639;
wire x_13640;
wire x_13641;
wire x_13642;
wire x_13643;
wire x_13644;
wire x_13645;
wire x_13646;
wire x_13647;
wire x_13648;
wire x_13649;
wire x_13650;
wire x_13651;
wire x_13652;
wire x_13653;
wire x_13654;
wire x_13655;
wire x_13656;
wire x_13657;
wire x_13658;
wire x_13659;
wire x_13660;
wire x_13661;
wire x_13662;
wire x_13663;
wire x_13664;
wire x_13665;
wire x_13666;
wire x_13667;
wire x_13668;
wire x_13669;
wire x_13670;
wire x_13671;
wire x_13672;
wire x_13673;
wire x_13674;
wire x_13675;
wire x_13676;
wire x_13677;
wire x_13678;
wire x_13679;
wire x_13680;
wire x_13681;
wire x_13682;
wire x_13683;
wire x_13684;
wire x_13685;
wire x_13686;
wire x_13687;
wire x_13688;
wire x_13689;
wire x_13690;
wire x_13691;
wire x_13692;
wire x_13693;
wire x_13694;
wire x_13695;
wire x_13696;
wire x_13697;
wire x_13698;
wire x_13699;
wire x_13700;
wire x_13701;
wire x_13702;
wire x_13703;
wire x_13704;
wire x_13705;
wire x_13706;
wire x_13707;
wire x_13708;
wire x_13709;
wire x_13710;
wire x_13711;
wire x_13712;
wire x_13713;
wire x_13714;
wire x_13715;
wire x_13716;
wire x_13717;
wire x_13718;
wire x_13719;
wire x_13720;
wire x_13721;
wire x_13722;
wire x_13723;
wire x_13724;
wire x_13725;
wire x_13726;
wire x_13727;
wire x_13728;
wire x_13729;
wire x_13730;
wire x_13731;
wire x_13732;
wire x_13733;
wire x_13734;
wire x_13735;
wire x_13736;
wire x_13737;
wire x_13738;
wire x_13739;
wire x_13740;
wire x_13741;
wire x_13742;
wire x_13743;
wire x_13744;
wire x_13745;
wire x_13746;
wire x_13747;
wire x_13748;
wire x_13749;
wire x_13750;
wire x_13751;
wire x_13752;
wire x_13753;
wire x_13754;
wire x_13755;
wire x_13756;
wire x_13757;
wire x_13758;
wire x_13759;
wire x_13760;
wire x_13761;
wire x_13762;
wire x_13763;
wire x_13764;
wire x_13765;
wire x_13766;
wire x_13767;
wire x_13768;
wire x_13769;
wire x_13770;
wire x_13771;
wire x_13772;
wire x_13773;
wire x_13774;
wire x_13775;
wire x_13776;
wire x_13777;
wire x_13778;
wire x_13779;
wire x_13780;
wire x_13781;
wire x_13782;
wire x_13783;
wire x_13784;
wire x_13785;
wire x_13786;
wire x_13787;
wire x_13788;
wire x_13789;
wire x_13790;
wire x_13791;
wire x_13792;
wire x_13793;
wire x_13794;
wire x_13795;
wire x_13796;
wire x_13797;
wire x_13798;
wire x_13799;
wire x_13800;
wire x_13801;
wire x_13802;
wire x_13803;
wire x_13804;
wire x_13805;
wire x_13806;
wire x_13807;
wire x_13808;
wire x_13809;
wire x_13810;
wire x_13811;
wire x_13812;
wire x_13813;
wire x_13814;
wire x_13815;
wire x_13816;
wire x_13817;
wire x_13818;
wire x_13819;
wire x_13820;
wire x_13821;
wire x_13822;
wire x_13823;
wire x_13824;
wire x_13825;
wire x_13826;
wire x_13827;
wire x_13828;
wire x_13829;
wire x_13830;
wire x_13831;
wire x_13832;
wire x_13833;
wire x_13834;
wire x_13835;
wire x_13836;
wire x_13837;
wire x_13838;
wire x_13839;
wire x_13840;
wire x_13841;
wire x_13842;
wire x_13843;
wire x_13844;
wire x_13845;
wire x_13846;
wire x_13847;
wire x_13848;
wire x_13849;
wire x_13850;
wire x_13851;
wire x_13852;
wire x_13853;
wire x_13854;
wire x_13855;
wire x_13856;
wire x_13857;
wire x_13858;
wire x_13859;
wire x_13860;
wire x_13861;
wire x_13862;
wire x_13863;
wire x_13864;
wire x_13865;
wire x_13866;
wire x_13867;
wire x_13868;
wire x_13869;
wire x_13870;
wire x_13871;
wire x_13872;
wire x_13873;
wire x_13874;
wire x_13875;
wire x_13876;
wire x_13877;
wire x_13878;
wire x_13879;
wire x_13880;
wire x_13881;
wire x_13882;
wire x_13883;
wire x_13884;
wire x_13885;
wire x_13886;
wire x_13887;
wire x_13888;
wire x_13889;
wire x_13890;
wire x_13891;
wire x_13892;
wire x_13893;
wire x_13894;
wire x_13895;
wire x_13896;
wire x_13897;
wire x_13898;
wire x_13899;
wire x_13900;
wire x_13901;
wire x_13902;
wire x_13903;
wire x_13904;
wire x_13905;
wire x_13906;
wire x_13907;
wire x_13908;
wire x_13909;
wire x_13910;
wire x_13911;
wire x_13912;
wire x_13913;
wire x_13914;
wire x_13915;
wire x_13916;
wire x_13917;
wire x_13918;
wire x_13919;
wire x_13920;
wire x_13921;
wire x_13922;
wire x_13923;
wire x_13924;
wire x_13925;
wire x_13926;
wire x_13927;
wire x_13928;
wire x_13929;
wire x_13930;
wire x_13931;
wire x_13932;
wire x_13933;
wire x_13934;
wire x_13935;
wire x_13936;
wire x_13937;
wire x_13938;
wire x_13939;
wire x_13940;
wire x_13941;
wire x_13942;
wire x_13943;
wire x_13944;
wire x_13945;
wire x_13946;
wire x_13947;
wire x_13948;
wire x_13949;
wire x_13950;
wire x_13951;
wire x_13952;
wire x_13953;
wire x_13954;
wire x_13955;
wire x_13956;
wire x_13957;
wire x_13958;
wire x_13959;
wire x_13960;
wire x_13961;
wire x_13962;
wire x_13963;
wire x_13964;
wire x_13965;
wire x_13966;
wire x_13967;
wire x_13968;
wire x_13969;
wire x_13970;
wire x_13971;
wire x_13972;
wire x_13973;
wire x_13974;
wire x_13975;
wire x_13976;
wire x_13977;
wire x_13978;
wire x_13979;
wire x_13980;
wire x_13981;
wire x_13982;
wire x_13983;
wire x_13984;
wire x_13985;
wire x_13986;
wire x_13987;
wire x_13988;
wire x_13989;
wire x_13990;
wire x_13991;
wire x_13992;
wire x_13993;
wire x_13994;
wire x_13995;
wire x_13996;
wire x_13997;
wire x_13998;
wire x_13999;
wire x_14000;
wire x_14001;
wire x_14002;
wire x_14003;
wire x_14004;
wire x_14005;
wire x_14006;
wire x_14007;
wire x_14008;
wire x_14009;
wire x_14010;
wire x_14011;
wire x_14012;
wire x_14013;
wire x_14014;
wire x_14015;
wire x_14016;
wire x_14017;
wire x_14018;
wire x_14019;
wire x_14020;
wire x_14021;
wire x_14022;
wire x_14023;
wire x_14024;
wire x_14025;
wire x_14026;
wire x_14027;
wire x_14028;
wire x_14029;
wire x_14030;
wire x_14031;
wire x_14032;
wire x_14033;
wire x_14034;
wire x_14035;
wire x_14036;
wire x_14037;
wire x_14038;
wire x_14039;
wire x_14040;
wire x_14041;
wire x_14042;
wire x_14043;
wire x_14044;
wire x_14045;
wire x_14046;
wire x_14047;
wire x_14048;
wire x_14049;
wire x_14050;
wire x_14051;
wire x_14052;
wire x_14053;
wire x_14054;
wire x_14055;
wire x_14056;
wire x_14057;
wire x_14058;
wire x_14059;
wire x_14060;
wire x_14061;
wire x_14062;
wire x_14063;
wire x_14064;
wire x_14065;
wire x_14066;
wire x_14067;
wire x_14068;
wire x_14069;
wire x_14070;
wire x_14071;
wire x_14072;
wire x_14073;
wire x_14074;
wire x_14075;
wire x_14076;
wire x_14077;
wire x_14078;
wire x_14079;
wire x_14080;
wire x_14081;
wire x_14082;
wire x_14083;
wire x_14084;
wire x_14085;
wire x_14086;
wire x_14087;
wire x_14088;
wire x_14089;
wire x_14090;
wire x_14091;
wire x_14092;
wire x_14093;
wire x_14094;
wire x_14095;
wire x_14096;
wire x_14097;
wire x_14098;
wire x_14099;
wire x_14100;
wire x_14101;
wire x_14102;
wire x_14103;
wire x_14104;
wire x_14105;
wire x_14106;
wire x_14107;
wire x_14108;
wire x_14109;
wire x_14110;
wire x_14111;
wire x_14112;
wire x_14113;
wire x_14114;
wire x_14115;
wire x_14116;
wire x_14117;
wire x_14118;
wire x_14119;
wire x_14120;
wire x_14121;
wire x_14122;
wire x_14123;
wire x_14124;
wire x_14125;
wire x_14126;
wire x_14127;
wire x_14128;
wire x_14129;
wire x_14130;
wire x_14131;
wire x_14132;
wire x_14133;
wire x_14134;
wire x_14135;
wire x_14136;
wire x_14137;
wire x_14138;
wire x_14139;
wire x_14140;
wire x_14141;
wire x_14142;
wire x_14143;
wire x_14144;
wire x_14145;
wire x_14146;
wire x_14147;
wire x_14148;
wire x_14149;
wire x_14150;
wire x_14151;
wire x_14152;
wire x_14153;
wire x_14154;
wire x_14155;
wire x_14156;
wire x_14157;
wire x_14158;
wire x_14159;
wire x_14160;
wire x_14161;
wire x_14162;
wire x_14163;
wire x_14164;
wire x_14165;
wire x_14166;
wire x_14167;
wire x_14168;
wire x_14169;
wire x_14170;
wire x_14171;
wire x_14172;
wire x_14173;
wire x_14174;
wire x_14175;
wire x_14176;
wire x_14177;
wire x_14178;
wire x_14179;
wire x_14180;
wire x_14181;
wire x_14182;
wire x_14183;
wire x_14184;
wire x_14185;
wire x_14186;
wire x_14187;
wire x_14188;
wire x_14189;
wire x_14190;
wire x_14191;
wire x_14192;
wire x_14193;
wire x_14194;
wire x_14195;
wire x_14196;
wire x_14197;
wire x_14198;
wire x_14199;
wire x_14200;
wire x_14201;
wire x_14202;
wire x_14203;
wire x_14204;
wire x_14205;
wire x_14206;
wire x_14207;
wire x_14208;
wire x_14209;
wire x_14210;
wire x_14211;
wire x_14212;
wire x_14213;
wire x_14214;
wire x_14215;
wire x_14216;
wire x_14217;
wire x_14218;
wire x_14219;
wire x_14220;
wire x_14221;
wire x_14222;
wire x_14223;
wire x_14224;
wire x_14225;
wire x_14226;
wire x_14227;
wire x_14228;
wire x_14229;
wire x_14230;
wire x_14231;
wire x_14232;
wire x_14233;
wire x_14234;
wire x_14235;
wire x_14236;
wire x_14237;
wire x_14238;
wire x_14239;
wire x_14240;
wire x_14241;
wire x_14242;
wire x_14243;
wire x_14244;
wire x_14245;
wire x_14246;
wire x_14247;
wire x_14248;
wire x_14249;
wire x_14250;
wire x_14251;
wire x_14252;
wire x_14253;
wire x_14254;
wire x_14255;
wire x_14256;
wire x_14257;
wire x_14258;
wire x_14259;
wire x_14260;
wire x_14261;
wire x_14262;
wire x_14263;
wire x_14264;
wire x_14265;
wire x_14266;
wire x_14267;
wire x_14268;
wire x_14269;
wire x_14270;
wire x_14271;
wire x_14272;
wire x_14273;
wire x_14274;
wire x_14275;
wire x_14276;
wire x_14277;
wire x_14278;
wire x_14279;
wire x_14280;
wire x_14281;
wire x_14282;
wire x_14283;
wire x_14284;
wire x_14285;
wire x_14286;
wire x_14287;
wire x_14288;
wire x_14289;
wire x_14290;
wire x_14291;
wire x_14292;
wire x_14293;
wire x_14294;
wire x_14295;
wire x_14296;
wire x_14297;
wire x_14298;
wire x_14299;
wire x_14300;
wire x_14301;
wire x_14302;
wire x_14303;
wire x_14304;
wire x_14305;
wire x_14306;
wire x_14307;
wire x_14308;
wire x_14309;
wire x_14310;
wire x_14311;
wire x_14312;
wire x_14313;
wire x_14314;
wire x_14315;
wire x_14316;
wire x_14317;
wire x_14318;
wire x_14319;
wire x_14320;
wire x_14321;
wire x_14322;
wire x_14323;
wire x_14324;
wire x_14325;
wire x_14326;
wire x_14327;
wire x_14328;
wire x_14329;
wire x_14330;
wire x_14331;
wire x_14332;
wire x_14333;
wire x_14334;
wire x_14335;
wire x_14336;
wire x_14337;
wire x_14338;
wire x_14339;
wire x_14340;
wire x_14341;
wire x_14342;
wire x_14343;
wire x_14344;
wire x_14345;
wire x_14346;
wire x_14347;
wire x_14348;
wire x_14349;
wire x_14350;
wire x_14351;
wire x_14352;
wire x_14353;
wire x_14354;
wire x_14355;
wire x_14356;
wire x_14357;
wire x_14358;
wire x_14359;
wire x_14360;
wire x_14361;
wire x_14362;
wire x_14363;
wire x_14364;
wire x_14365;
wire x_14366;
wire x_14367;
wire x_14368;
wire x_14369;
wire x_14370;
wire x_14371;
wire x_14372;
wire x_14373;
wire x_14374;
wire x_14375;
wire x_14376;
wire x_14377;
wire x_14378;
wire x_14379;
wire x_14380;
wire x_14381;
wire x_14382;
wire x_14383;
wire x_14384;
wire x_14385;
wire x_14386;
wire x_14387;
wire x_14388;
wire x_14389;
wire x_14390;
wire x_14391;
wire x_14392;
wire x_14393;
wire x_14394;
wire x_14395;
wire x_14396;
wire x_14397;
wire x_14398;
wire x_14399;
wire x_14400;
wire x_14401;
wire x_14402;
wire x_14403;
wire x_14404;
wire x_14405;
wire x_14406;
wire x_14407;
wire x_14408;
wire x_14409;
wire x_14410;
wire x_14411;
wire x_14412;
wire x_14413;
wire x_14414;
wire x_14415;
wire x_14416;
wire x_14417;
wire x_14418;
wire x_14419;
wire x_14420;
wire x_14421;
wire x_14422;
wire x_14423;
wire x_14424;
wire x_14425;
wire x_14426;
wire x_14427;
wire x_14428;
wire x_14429;
wire x_14430;
wire x_14431;
wire x_14432;
wire x_14433;
wire x_14434;
wire x_14435;
wire x_14436;
wire x_14437;
wire x_14438;
wire x_14439;
wire x_14440;
wire x_14441;
wire x_14442;
wire x_14443;
wire x_14444;
wire x_14445;
wire x_14446;
wire x_14447;
wire x_14448;
wire x_14449;
wire x_14450;
wire x_14451;
wire x_14452;
wire x_14453;
wire x_14454;
wire x_14455;
wire x_14456;
wire x_14457;
wire x_14458;
wire x_14459;
wire x_14460;
wire x_14461;
wire x_14462;
wire x_14463;
wire x_14464;
wire x_14465;
wire x_14466;
wire x_14467;
wire x_14468;
wire x_14469;
wire x_14470;
wire x_14471;
wire x_14472;
wire x_14473;
wire x_14474;
wire x_14475;
wire x_14476;
wire x_14477;
wire x_14478;
wire x_14479;
wire x_14480;
wire x_14481;
wire x_14482;
wire x_14483;
wire x_14484;
wire x_14485;
wire x_14486;
wire x_14487;
wire x_14488;
wire x_14489;
wire x_14490;
wire x_14491;
wire x_14492;
wire x_14493;
wire x_14494;
wire x_14495;
wire x_14496;
wire x_14497;
wire x_14498;
wire x_14499;
wire x_14500;
wire x_14501;
wire x_14502;
wire x_14503;
wire x_14504;
wire x_14505;
wire x_14506;
wire x_14507;
wire x_14508;
wire x_14509;
wire x_14510;
wire x_14511;
wire x_14512;
wire x_14513;
wire x_14514;
wire x_14515;
wire x_14516;
wire x_14517;
wire x_14518;
wire x_14519;
wire x_14520;
wire x_14521;
wire x_14522;
wire x_14523;
wire x_14524;
wire x_14525;
wire x_14526;
wire x_14527;
wire x_14528;
wire x_14529;
wire x_14530;
wire x_14531;
wire x_14532;
wire x_14533;
wire x_14534;
wire x_14535;
wire x_14536;
wire x_14537;
wire x_14538;
wire x_14539;
wire x_14540;
wire x_14541;
wire x_14542;
wire x_14543;
wire x_14544;
wire x_14545;
wire x_14546;
wire x_14547;
wire x_14548;
wire x_14549;
wire x_14550;
wire x_14551;
wire x_14552;
wire x_14553;
wire x_14554;
wire x_14555;
wire x_14556;
wire x_14557;
wire x_14558;
wire x_14559;
wire x_14560;
wire x_14561;
wire x_14562;
wire x_14563;
wire x_14564;
wire x_14565;
wire x_14566;
wire x_14567;
wire x_14568;
wire x_14569;
wire x_14570;
wire x_14571;
wire x_14572;
wire x_14573;
wire x_14574;
wire x_14575;
wire x_14576;
wire x_14577;
wire x_14578;
wire x_14579;
wire x_14580;
wire x_14581;
wire x_14582;
wire x_14583;
wire x_14584;
wire x_14585;
wire x_14586;
wire x_14587;
wire x_14588;
wire x_14589;
wire x_14590;
wire x_14591;
wire x_14592;
wire x_14593;
wire x_14594;
wire x_14595;
wire x_14596;
wire x_14597;
wire x_14598;
wire x_14599;
wire x_14600;
wire x_14601;
wire x_14602;
wire x_14603;
wire x_14604;
wire x_14605;
wire x_14606;
wire x_14607;
wire x_14608;
wire x_14609;
wire x_14610;
wire x_14611;
wire x_14612;
wire x_14613;
wire x_14614;
wire x_14615;
wire x_14616;
wire x_14617;
wire x_14618;
wire x_14619;
wire x_14620;
wire x_14621;
wire x_14622;
wire x_14623;
wire x_14624;
wire x_14625;
wire x_14626;
wire x_14627;
wire x_14628;
wire x_14629;
wire x_14630;
wire x_14631;
wire x_14632;
wire x_14633;
wire x_14634;
wire x_14635;
wire x_14636;
wire x_14637;
wire x_14638;
wire x_14639;
wire x_14640;
wire x_14641;
wire x_14642;
wire x_14643;
wire x_14644;
wire x_14645;
wire x_14646;
wire x_14647;
wire x_14648;
wire x_14649;
wire x_14650;
wire x_14651;
wire x_14652;
wire x_14653;
wire x_14654;
wire x_14655;
wire x_14656;
wire x_14657;
wire x_14658;
wire x_14659;
wire x_14660;
wire x_14661;
wire x_14662;
wire x_14663;
wire x_14664;
wire x_14665;
wire x_14666;
wire x_14667;
wire x_14668;
wire x_14669;
wire x_14670;
wire x_14671;
wire x_14672;
wire x_14673;
wire x_14674;
wire x_14675;
wire x_14676;
wire x_14677;
wire x_14678;
wire x_14679;
wire x_14680;
wire x_14681;
wire x_14682;
wire x_14683;
wire x_14684;
wire x_14685;
wire x_14686;
wire x_14687;
wire x_14688;
wire x_14689;
wire x_14690;
wire x_14691;
wire x_14692;
wire x_14693;
wire x_14694;
wire x_14695;
wire x_14696;
wire x_14697;
wire x_14698;
wire x_14699;
wire x_14700;
wire x_14701;
wire x_14702;
wire x_14703;
wire x_14704;
wire x_14705;
wire x_14706;
wire x_14707;
wire x_14708;
wire x_14709;
wire x_14710;
wire x_14711;
wire x_14712;
wire x_14713;
wire x_14714;
wire x_14715;
wire x_14716;
wire x_14717;
wire x_14718;
wire x_14719;
wire x_14720;
wire x_14721;
wire x_14722;
wire x_14723;
wire x_14724;
wire x_14725;
wire x_14726;
wire x_14727;
wire x_14728;
wire x_14729;
wire x_14730;
wire x_14731;
wire x_14732;
wire x_14733;
wire x_14734;
wire x_14735;
wire x_14736;
wire x_14737;
wire x_14738;
wire x_14739;
wire x_14740;
wire x_14741;
wire x_14742;
wire x_14743;
wire x_14744;
wire x_14745;
wire x_14746;
wire x_14747;
wire x_14748;
wire x_14749;
wire x_14750;
wire x_14751;
wire x_14752;
wire x_14753;
wire x_14754;
wire x_14755;
wire x_14756;
wire x_14757;
wire x_14758;
wire x_14759;
wire x_14760;
wire x_14761;
wire x_14762;
wire x_14763;
wire x_14764;
wire x_14765;
wire x_14766;
wire x_14767;
wire x_14768;
wire x_14769;
wire x_14770;
wire x_14771;
wire x_14772;
wire x_14773;
wire x_14774;
wire x_14775;
wire x_14776;
wire x_14777;
wire x_14778;
wire x_14779;
wire x_14780;
wire x_14781;
wire x_14782;
wire x_14783;
wire x_14784;
wire x_14785;
wire x_14786;
wire x_14787;
wire x_14788;
wire x_14789;
wire x_14790;
wire x_14791;
wire x_14792;
wire x_14793;
wire x_14794;
wire x_14795;
wire x_14796;
wire x_14797;
wire x_14798;
wire x_14799;
wire x_14800;
wire x_14801;
wire x_14802;
wire x_14803;
wire x_14804;
wire x_14805;
wire x_14806;
wire x_14807;
wire x_14808;
wire x_14809;
wire x_14810;
wire x_14811;
wire x_14812;
wire x_14813;
wire x_14814;
wire x_14815;
wire x_14816;
wire x_14817;
wire x_14818;
wire x_14819;
wire x_14820;
wire x_14821;
wire x_14822;
wire x_14823;
wire x_14824;
wire x_14825;
wire x_14826;
wire x_14827;
wire x_14828;
wire x_14829;
wire x_14830;
wire x_14831;
wire x_14832;
wire x_14833;
wire x_14834;
wire x_14835;
wire x_14836;
wire x_14837;
wire x_14838;
wire x_14839;
wire x_14840;
wire x_14841;
wire x_14842;
wire x_14843;
wire x_14844;
wire x_14845;
wire x_14846;
wire x_14847;
wire x_14848;
wire x_14849;
wire x_14850;
wire x_14851;
wire x_14852;
wire x_14853;
wire x_14854;
wire x_14855;
wire x_14856;
wire x_14857;
wire x_14858;
wire x_14859;
wire x_14860;
wire x_14861;
wire x_14862;
wire x_14863;
wire x_14864;
wire x_14865;
wire x_14866;
wire x_14867;
wire x_14868;
wire x_14869;
wire x_14870;
wire x_14871;
wire x_14872;
wire x_14873;
wire x_14874;
wire x_14875;
wire x_14876;
wire x_14877;
wire x_14878;
wire x_14879;
wire x_14880;
wire x_14881;
wire x_14882;
wire x_14883;
wire x_14884;
wire x_14885;
wire x_14886;
wire x_14887;
wire x_14888;
wire x_14889;
wire x_14890;
wire x_14891;
wire x_14892;
wire x_14893;
wire x_14894;
wire x_14895;
wire x_14896;
wire x_14897;
wire x_14898;
wire x_14899;
wire x_14900;
wire x_14901;
wire x_14902;
wire x_14903;
wire x_14904;
wire x_14905;
wire x_14906;
wire x_14907;
wire x_14908;
wire x_14909;
wire x_14910;
wire x_14911;
wire x_14912;
wire x_14913;
wire x_14914;
wire x_14915;
wire x_14916;
wire x_14917;
wire x_14918;
wire x_14919;
wire x_14920;
wire x_14921;
wire x_14922;
wire x_14923;
wire x_14924;
wire x_14925;
wire x_14926;
wire x_14927;
wire x_14928;
wire x_14929;
wire x_14930;
wire x_14931;
wire x_14932;
wire x_14933;
wire x_14934;
wire x_14935;
wire x_14936;
wire x_14937;
wire x_14938;
wire x_14939;
wire x_14940;
wire x_14941;
wire x_14942;
wire x_14943;
wire x_14944;
wire x_14945;
wire x_14946;
wire x_14947;
wire x_14948;
wire x_14949;
wire x_14950;
wire x_14951;
wire x_14952;
wire x_14953;
wire x_14954;
wire x_14955;
wire x_14956;
wire x_14957;
wire x_14958;
wire x_14959;
wire x_14960;
wire x_14961;
wire x_14962;
wire x_14963;
wire x_14964;
wire x_14965;
wire x_14966;
wire x_14967;
wire x_14968;
wire x_14969;
wire x_14970;
wire x_14971;
wire x_14972;
wire x_14973;
wire x_14974;
wire x_14975;
wire x_14976;
wire x_14977;
wire x_14978;
wire x_14979;
wire x_14980;
wire x_14981;
wire x_14982;
wire x_14983;
wire x_14984;
wire x_14985;
wire x_14986;
wire x_14987;
wire x_14988;
wire x_14989;
wire x_14990;
wire x_14991;
wire x_14992;
wire x_14993;
wire x_14994;
wire x_14995;
wire x_14996;
wire x_14997;
wire x_14998;
wire x_14999;
wire x_15000;
wire x_15001;
wire x_15002;
wire x_15003;
wire x_15004;
wire x_15005;
wire x_15006;
wire x_15007;
wire x_15008;
wire x_15009;
wire x_15010;
wire x_15011;
wire x_15012;
wire x_15013;
wire x_15014;
wire x_15015;
wire x_15016;
wire x_15017;
wire x_15018;
wire x_15019;
wire x_15020;
wire x_15021;
wire x_15022;
wire x_15023;
wire x_15024;
wire x_15025;
wire x_15026;
wire x_15027;
wire x_15028;
wire x_15029;
wire x_15030;
wire x_15031;
wire x_15032;
wire x_15033;
wire x_15034;
wire x_15035;
wire x_15036;
wire x_15037;
wire x_15038;
wire x_15039;
wire x_15040;
wire x_15041;
wire x_15042;
wire x_15043;
wire x_15044;
wire x_15045;
wire x_15046;
wire x_15047;
wire x_15048;
wire x_15049;
wire x_15050;
wire x_15051;
wire x_15052;
wire x_15053;
wire x_15054;
wire x_15055;
wire x_15056;
wire x_15057;
wire x_15058;
wire x_15059;
wire x_15060;
wire x_15061;
wire x_15062;
wire x_15063;
wire x_15064;
wire x_15065;
wire x_15066;
wire x_15067;
wire x_15068;
wire x_15069;
wire x_15070;
wire x_15071;
wire x_15072;
wire x_15073;
wire x_15074;
wire x_15075;
wire x_15076;
wire x_15077;
wire x_15078;
wire x_15079;
wire x_15080;
wire x_15081;
wire x_15082;
wire x_15083;
wire x_15084;
wire x_15085;
wire x_15086;
wire x_15087;
wire x_15088;
wire x_15089;
wire x_15090;
wire x_15091;
wire x_15092;
wire x_15093;
wire x_15094;
wire x_15095;
wire x_15096;
wire x_15097;
wire x_15098;
wire x_15099;
wire x_15100;
wire x_15101;
wire x_15102;
wire x_15103;
wire x_15104;
wire x_15105;
wire x_15106;
wire x_15107;
wire x_15108;
wire x_15109;
wire x_15110;
wire x_15111;
wire x_15112;
wire x_15113;
wire x_15114;
wire x_15115;
wire x_15116;
wire x_15117;
wire x_15118;
wire x_15119;
wire x_15120;
wire x_15121;
wire x_15122;
wire x_15123;
wire x_15124;
wire x_15125;
wire x_15126;
wire x_15127;
wire x_15128;
wire x_15129;
wire x_15130;
wire x_15131;
wire x_15132;
wire x_15133;
wire x_15134;
wire x_15135;
wire x_15136;
wire x_15137;
wire x_15138;
wire x_15139;
wire x_15140;
wire x_15141;
wire x_15142;
wire x_15143;
wire x_15144;
wire x_15145;
wire x_15146;
wire x_15147;
wire x_15148;
wire x_15149;
wire x_15150;
wire x_15151;
wire x_15152;
wire x_15153;
wire x_15154;
wire x_15155;
wire x_15156;
wire x_15157;
wire x_15158;
wire x_15159;
wire x_15160;
wire x_15161;
wire x_15162;
wire x_15163;
wire x_15164;
wire x_15165;
wire x_15166;
wire x_15167;
wire x_15168;
wire x_15169;
wire x_15170;
wire x_15171;
wire x_15172;
wire x_15173;
wire x_15174;
wire x_15175;
wire x_15176;
wire x_15177;
wire x_15178;
wire x_15179;
wire x_15180;
wire x_15181;
wire x_15182;
wire x_15183;
wire x_15184;
wire x_15185;
wire x_15186;
wire x_15187;
wire x_15188;
wire x_15189;
wire x_15190;
wire x_15191;
wire x_15192;
wire x_15193;
wire x_15194;
wire x_15195;
wire x_15196;
wire x_15197;
wire x_15198;
wire x_15199;
wire x_15200;
wire x_15201;
wire x_15202;
wire x_15203;
wire x_15204;
wire x_15205;
wire x_15206;
wire x_15207;
wire x_15208;
wire x_15209;
wire x_15210;
wire x_15211;
wire x_15212;
wire x_15213;
wire x_15214;
wire x_15215;
wire x_15216;
wire x_15217;
wire x_15218;
wire x_15219;
wire x_15220;
wire x_15221;
wire x_15222;
wire x_15223;
wire x_15224;
wire x_15225;
wire x_15226;
wire x_15227;
wire x_15228;
wire x_15229;
wire x_15230;
wire x_15231;
wire x_15232;
wire x_15233;
wire x_15234;
wire x_15235;
wire x_15236;
wire x_15237;
wire x_15238;
wire x_15239;
wire x_15240;
wire x_15241;
wire x_15242;
wire x_15243;
wire x_15244;
wire x_15245;
wire x_15246;
wire x_15247;
wire x_15248;
wire x_15249;
wire x_15250;
wire x_15251;
wire x_15252;
wire x_15253;
wire x_15254;
wire x_15255;
wire x_15256;
wire x_15257;
wire x_15258;
wire x_15259;
wire x_15260;
wire x_15261;
wire x_15262;
wire x_15263;
wire x_15264;
wire x_15265;
wire x_15266;
wire x_15267;
wire x_15268;
wire x_15269;
wire x_15270;
wire x_15271;
wire x_15272;
wire x_15273;
wire x_15274;
wire x_15275;
wire x_15276;
wire x_15277;
wire x_15278;
wire x_15279;
wire x_15280;
wire x_15281;
wire x_15282;
wire x_15283;
wire x_15284;
wire x_15285;
wire x_15286;
wire x_15287;
wire x_15288;
wire x_15289;
wire x_15290;
wire x_15291;
wire x_15292;
wire x_15293;
wire x_15294;
wire x_15295;
wire x_15296;
wire x_15297;
wire x_15298;
wire x_15299;
wire x_15300;
wire x_15301;
wire x_15302;
wire x_15303;
wire x_15304;
wire x_15305;
wire x_15306;
wire x_15307;
wire x_15308;
wire x_15309;
wire x_15310;
wire x_15311;
wire x_15312;
wire x_15313;
wire x_15314;
wire x_15315;
wire x_15316;
wire x_15317;
wire x_15318;
wire x_15319;
wire x_15320;
wire x_15321;
wire x_15322;
wire x_15323;
wire x_15324;
wire x_15325;
wire x_15326;
wire x_15327;
wire x_15328;
wire x_15329;
wire x_15330;
wire x_15331;
wire x_15332;
wire x_15333;
wire x_15334;
wire x_15335;
wire x_15336;
wire x_15337;
wire x_15338;
wire x_15339;
wire x_15340;
wire x_15341;
wire x_15342;
wire x_15343;
wire x_15344;
wire x_15345;
wire x_15346;
wire x_15347;
wire x_15348;
wire x_15349;
wire x_15350;
wire x_15351;
wire x_15352;
wire x_15353;
wire x_15354;
wire x_15355;
wire x_15356;
wire x_15357;
wire x_15358;
wire x_15359;
wire x_15360;
wire x_15361;
wire x_15362;
wire x_15363;
wire x_15364;
wire x_15365;
wire x_15366;
wire x_15367;
wire x_15368;
wire x_15369;
wire x_15370;
wire x_15371;
wire x_15372;
wire x_15373;
wire x_15374;
wire x_15375;
wire x_15376;
wire x_15377;
wire x_15378;
wire x_15379;
wire x_15380;
wire x_15381;
wire x_15382;
wire x_15383;
wire x_15384;
wire x_15385;
wire x_15386;
wire x_15387;
wire x_15388;
wire x_15389;
wire x_15390;
wire x_15391;
wire x_15392;
wire x_15393;
wire x_15394;
wire x_15395;
wire x_15396;
wire x_15397;
wire x_15398;
wire x_15399;
wire x_15400;
wire x_15401;
wire x_15402;
wire x_15403;
wire x_15404;
wire x_15405;
wire x_15406;
wire x_15407;
wire x_15408;
wire x_15409;
wire x_15410;
wire x_15411;
wire x_15412;
wire x_15413;
wire x_15414;
wire x_15415;
wire x_15416;
wire x_15417;
wire x_15418;
wire x_15419;
wire x_15420;
wire x_15421;
wire x_15422;
wire x_15423;
wire x_15424;
wire x_15425;
wire x_15426;
wire x_15427;
wire x_15428;
wire x_15429;
wire x_15430;
wire x_15431;
wire x_15432;
wire x_15433;
wire x_15434;
wire x_15435;
wire x_15436;
wire x_15437;
wire x_15438;
wire x_15439;
wire x_15440;
wire x_15441;
wire x_15442;
wire x_15443;
wire x_15444;
wire x_15445;
wire x_15446;
wire x_15447;
wire x_15448;
wire x_15449;
wire x_15450;
wire x_15451;
wire x_15452;
wire x_15453;
wire x_15454;
wire x_15455;
wire x_15456;
wire x_15457;
wire x_15458;
wire x_15459;
wire x_15460;
wire x_15461;
wire x_15462;
wire x_15463;
wire x_15464;
wire x_15465;
wire x_15466;
wire x_15467;
wire x_15468;
wire x_15469;
wire x_15470;
wire x_15471;
wire x_15472;
wire x_15473;
wire x_15474;
wire x_15475;
wire x_15476;
wire x_15477;
wire x_15478;
wire x_15479;
wire x_15480;
wire x_15481;
wire x_15482;
wire x_15483;
wire x_15484;
wire x_15485;
wire x_15486;
wire x_15487;
wire x_15488;
wire x_15489;
wire x_15490;
wire x_15491;
wire x_15492;
wire x_15493;
wire x_15494;
wire x_15495;
wire x_15496;
wire x_15497;
wire x_15498;
wire x_15499;
wire x_15500;
wire x_15501;
wire x_15502;
wire x_15503;
wire x_15504;
wire x_15505;
wire x_15506;
wire x_15507;
wire x_15508;
wire x_15509;
wire x_15510;
wire x_15511;
wire x_15512;
wire x_15513;
wire x_15514;
wire x_15515;
wire x_15516;
wire x_15517;
wire x_15518;
wire x_15519;
wire x_15520;
wire x_15521;
wire x_15522;
wire x_15523;
wire x_15524;
wire x_15525;
wire x_15526;
wire x_15527;
wire x_15528;
wire x_15529;
wire x_15530;
wire x_15531;
wire x_15532;
wire x_15533;
wire x_15534;
wire x_15535;
wire x_15536;
wire x_15537;
wire x_15538;
wire x_15539;
wire x_15540;
wire x_15541;
wire x_15542;
wire x_15543;
wire x_15544;
wire x_15545;
wire x_15546;
wire x_15547;
wire x_15548;
wire x_15549;
wire x_15550;
wire x_15551;
wire x_15552;
wire x_15553;
wire x_15554;
wire x_15555;
wire x_15556;
wire x_15557;
wire x_15558;
wire x_15559;
wire x_15560;
wire x_15561;
wire x_15562;
wire x_15563;
wire x_15564;
wire x_15565;
wire x_15566;
wire x_15567;
wire x_15568;
wire x_15569;
wire x_15570;
wire x_15571;
wire x_15572;
wire x_15573;
wire x_15574;
wire x_15575;
wire x_15576;
wire x_15577;
wire x_15578;
wire x_15579;
wire x_15580;
wire x_15581;
wire x_15582;
wire x_15583;
wire x_15584;
wire x_15585;
wire x_15586;
wire x_15587;
wire x_15588;
wire x_15589;
wire x_15590;
wire x_15591;
wire x_15592;
wire x_15593;
wire x_15594;
wire x_15595;
wire x_15596;
wire x_15597;
wire x_15598;
wire x_15599;
wire x_15600;
wire x_15601;
wire x_15602;
wire x_15603;
wire x_15604;
wire x_15605;
wire x_15606;
wire x_15607;
wire x_15608;
wire x_15609;
wire x_15610;
wire x_15611;
wire x_15612;
wire x_15613;
wire x_15614;
wire x_15615;
wire x_15616;
wire x_15617;
wire x_15618;
wire x_15619;
wire x_15620;
wire x_15621;
wire x_15622;
wire x_15623;
wire x_15624;
wire x_15625;
wire x_15626;
wire x_15627;
wire x_15628;
wire x_15629;
wire x_15630;
wire x_15631;
wire x_15632;
wire x_15633;
wire x_15634;
wire x_15635;
wire x_15636;
wire x_15637;
wire x_15638;
wire x_15639;
wire x_15640;
wire x_15641;
wire x_15642;
wire x_15643;
wire x_15644;
wire x_15645;
wire x_15646;
wire x_15647;
wire x_15648;
wire x_15649;
wire x_15650;
wire x_15651;
wire x_15652;
wire x_15653;
wire x_15654;
wire x_15655;
wire x_15656;
wire x_15657;
wire x_15658;
wire x_15659;
wire x_15660;
wire x_15661;
wire x_15662;
wire x_15663;
wire x_15664;
wire x_15665;
wire x_15666;
wire x_15667;
wire x_15668;
wire x_15669;
wire x_15670;
wire x_15671;
wire x_15672;
wire x_15673;
wire x_15674;
wire x_15675;
wire x_15676;
wire x_15677;
wire x_15678;
wire x_15679;
wire x_15680;
wire x_15681;
wire x_15682;
wire x_15683;
wire x_15684;
wire x_15685;
wire x_15686;
wire x_15687;
wire x_15688;
wire x_15689;
wire x_15690;
wire x_15691;
wire x_15692;
wire x_15693;
wire x_15694;
wire x_15695;
wire x_15696;
wire x_15697;
wire x_15698;
wire x_15699;
wire x_15700;
wire x_15701;
wire x_15702;
wire x_15703;
wire x_15704;
wire x_15705;
wire x_15706;
wire x_15707;
wire x_15708;
wire x_15709;
wire x_15710;
wire x_15711;
wire x_15712;
wire x_15713;
wire x_15714;
wire x_15715;
wire x_15716;
wire x_15717;
wire x_15718;
wire x_15719;
wire x_15720;
wire x_15721;
wire x_15722;
wire x_15723;
wire x_15724;
wire x_15725;
wire x_15726;
wire x_15727;
wire x_15728;
wire x_15729;
wire x_15730;
wire x_15731;
wire x_15732;
wire x_15733;
wire x_15734;
wire x_15735;
wire x_15736;
wire x_15737;
wire x_15738;
wire x_15739;
wire x_15740;
wire x_15741;
wire x_15742;
wire x_15743;
wire x_15744;
wire x_15745;
wire x_15746;
wire x_15747;
wire x_15748;
wire x_15749;
wire x_15750;
wire x_15751;
wire x_15752;
wire x_15753;
wire x_15754;
wire x_15755;
wire x_15756;
wire x_15757;
wire x_15758;
wire x_15759;
wire x_15760;
wire x_15761;
wire x_15762;
wire x_15763;
wire x_15764;
wire x_15765;
wire x_15766;
wire x_15767;
wire x_15768;
wire x_15769;
wire x_15770;
wire x_15771;
wire x_15772;
wire x_15773;
wire x_15774;
wire x_15775;
wire x_15776;
wire x_15777;
wire x_15778;
wire x_15779;
wire x_15780;
wire x_15781;
wire x_15782;
wire x_15783;
wire x_15784;
wire x_15785;
wire x_15786;
wire x_15787;
wire x_15788;
wire x_15789;
wire x_15790;
wire x_15791;
wire x_15792;
wire x_15793;
wire x_15794;
wire x_15795;
wire x_15796;
wire x_15797;
wire x_15798;
wire x_15799;
wire x_15800;
wire x_15801;
wire x_15802;
wire x_15803;
wire x_15804;
wire x_15805;
wire x_15806;
wire x_15807;
wire x_15808;
wire x_15809;
wire x_15810;
wire x_15811;
wire x_15812;
wire x_15813;
wire x_15814;
wire x_15815;
wire x_15816;
wire x_15817;
wire x_15818;
wire x_15819;
wire x_15820;
wire x_15821;
wire x_15822;
wire x_15823;
wire x_15824;
wire x_15825;
wire x_15826;
wire x_15827;
wire x_15828;
wire x_15829;
wire x_15830;
wire x_15831;
wire x_15832;
wire x_15833;
wire x_15834;
wire x_15835;
wire x_15836;
wire x_15837;
wire x_15838;
wire x_15839;
wire x_15840;
wire x_15841;
wire x_15842;
wire x_15843;
wire x_15844;
wire x_15845;
wire x_15846;
wire x_15847;
wire x_15848;
wire x_15849;
wire x_15850;
wire x_15851;
wire x_15852;
wire x_15853;
wire x_15854;
wire x_15855;
wire x_15856;
wire x_15857;
wire x_15858;
wire x_15859;
wire x_15860;
wire x_15861;
wire x_15862;
wire x_15863;
wire x_15864;
wire x_15865;
wire x_15866;
wire x_15867;
wire x_15868;
wire x_15869;
wire x_15870;
wire x_15871;
wire x_15872;
wire x_15873;
wire x_15874;
wire x_15875;
wire x_15876;
wire x_15877;
wire x_15878;
wire x_15879;
wire x_15880;
wire x_15881;
wire x_15882;
wire x_15883;
wire x_15884;
wire x_15885;
wire x_15886;
wire x_15887;
wire x_15888;
wire x_15889;
wire x_15890;
wire x_15891;
wire x_15892;
wire x_15893;
wire x_15894;
wire x_15895;
wire x_15896;
wire x_15897;
wire x_15898;
wire x_15899;
wire x_15900;
wire x_15901;
wire x_15902;
wire x_15903;
wire x_15904;
wire x_15905;
wire x_15906;
wire x_15907;
wire x_15908;
wire x_15909;
wire x_15910;
wire x_15911;
wire x_15912;
wire x_15913;
wire x_15914;
wire x_15915;
wire x_15916;
wire x_15917;
wire x_15918;
wire x_15919;
wire x_15920;
wire x_15921;
wire x_15922;
wire x_15923;
wire x_15924;
wire x_15925;
wire x_15926;
wire x_15927;
wire x_15928;
wire x_15929;
wire x_15930;
wire x_15931;
wire x_15932;
wire x_15933;
wire x_15934;
wire x_15935;
wire x_15936;
wire x_15937;
wire x_15938;
wire x_15939;
wire x_15940;
wire x_15941;
wire x_15942;
wire x_15943;
wire x_15944;
wire x_15945;
wire x_15946;
wire x_15947;
wire x_15948;
wire x_15949;
wire x_15950;
wire x_15951;
wire x_15952;
wire x_15953;
wire x_15954;
wire x_15955;
wire x_15956;
wire x_15957;
wire x_15958;
wire x_15959;
wire x_15960;
wire x_15961;
wire x_15962;
wire x_15963;
wire x_15964;
wire x_15965;
wire x_15966;
wire x_15967;
wire x_15968;
wire x_15969;
wire x_15970;
wire x_15971;
wire x_15972;
wire x_15973;
wire x_15974;
wire x_15975;
wire x_15976;
wire x_15977;
wire x_15978;
wire x_15979;
wire x_15980;
wire x_15981;
wire x_15982;
wire x_15983;
wire x_15984;
wire x_15985;
wire x_15986;
wire x_15987;
wire x_15988;
wire x_15989;
wire x_15990;
wire x_15991;
wire x_15992;
wire x_15993;
wire x_15994;
wire x_15995;
wire x_15996;
wire x_15997;
wire x_15998;
wire x_15999;
wire x_16000;
wire x_16001;
wire x_16002;
wire x_16003;
wire x_16004;
wire x_16005;
wire x_16006;
wire x_16007;
wire x_16008;
wire x_16009;
wire x_16010;
wire x_16011;
wire x_16012;
wire x_16013;
wire x_16014;
wire x_16015;
wire x_16016;
wire x_16017;
wire x_16018;
wire x_16019;
wire x_16020;
wire x_16021;
wire x_16022;
wire x_16023;
wire x_16024;
wire x_16025;
wire x_16026;
wire x_16027;
wire x_16028;
wire x_16029;
wire x_16030;
wire x_16031;
wire x_16032;
wire x_16033;
wire x_16034;
wire x_16035;
wire x_16036;
wire x_16037;
wire x_16038;
wire x_16039;
wire x_16040;
wire x_16041;
wire x_16042;
wire x_16043;
wire x_16044;
wire x_16045;
wire x_16046;
wire x_16047;
wire x_16048;
wire x_16049;
wire x_16050;
wire x_16051;
wire x_16052;
wire x_16053;
wire x_16054;
wire x_16055;
wire x_16056;
wire x_16057;
wire x_16058;
wire x_16059;
wire x_16060;
wire x_16061;
wire x_16062;
wire x_16063;
wire x_16064;
wire x_16065;
wire x_16066;
wire x_16067;
wire x_16068;
wire x_16069;
wire x_16070;
wire x_16071;
wire x_16072;
wire x_16073;
wire x_16074;
wire x_16075;
wire x_16076;
wire x_16077;
wire x_16078;
wire x_16079;
wire x_16080;
wire x_16081;
wire x_16082;
wire x_16083;
wire x_16084;
wire x_16085;
wire x_16086;
wire x_16087;
wire x_16088;
wire x_16089;
wire x_16090;
wire x_16091;
wire x_16092;
wire x_16093;
wire x_16094;
wire x_16095;
wire x_16096;
wire x_16097;
wire x_16098;
wire x_16099;
wire x_16100;
wire x_16101;
wire x_16102;
wire x_16103;
wire x_16104;
wire x_16105;
wire x_16106;
wire x_16107;
wire x_16108;
wire x_16109;
wire x_16110;
wire x_16111;
wire x_16112;
wire x_16113;
wire x_16114;
wire x_16115;
wire x_16116;
wire x_16117;
wire x_16118;
wire x_16119;
wire x_16120;
wire x_16121;
wire x_16122;
wire x_16123;
wire x_16124;
wire x_16125;
wire x_16126;
wire x_16127;
wire x_16128;
wire x_16129;
wire x_16130;
wire x_16131;
wire x_16132;
wire x_16133;
wire x_16134;
wire x_16135;
wire x_16136;
wire x_16137;
wire x_16138;
wire x_16139;
wire x_16140;
wire x_16141;
wire x_16142;
wire x_16143;
wire x_16144;
wire x_16145;
wire x_16146;
wire x_16147;
wire x_16148;
wire x_16149;
wire x_16150;
wire x_16151;
wire x_16152;
wire x_16153;
wire x_16154;
wire x_16155;
wire x_16156;
wire x_16157;
wire x_16158;
wire x_16159;
wire x_16160;
wire x_16161;
wire x_16162;
wire x_16163;
wire x_16164;
wire x_16165;
wire x_16166;
wire x_16167;
wire x_16168;
wire x_16169;
wire x_16170;
wire x_16171;
wire x_16172;
wire x_16173;
wire x_16174;
wire x_16175;
wire x_16176;
wire x_16177;
wire x_16178;
wire x_16179;
wire x_16180;
wire x_16181;
wire x_16182;
wire x_16183;
wire x_16184;
wire x_16185;
wire x_16186;
wire x_16187;
wire x_16188;
wire x_16189;
wire x_16190;
wire x_16191;
wire x_16192;
wire x_16193;
wire x_16194;
wire x_16195;
wire x_16196;
wire x_16197;
wire x_16198;
wire x_16199;
wire x_16200;
wire x_16201;
wire x_16202;
wire x_16203;
wire x_16204;
wire x_16205;
wire x_16206;
wire x_16207;
wire x_16208;
wire x_16209;
wire x_16210;
wire x_16211;
wire x_16212;
wire x_16213;
wire x_16214;
wire x_16215;
wire x_16216;
wire x_16217;
wire x_16218;
wire x_16219;
wire x_16220;
wire x_16221;
wire x_16222;
wire x_16223;
wire x_16224;
wire x_16225;
wire x_16226;
wire x_16227;
wire x_16228;
wire x_16229;
wire x_16230;
wire x_16231;
wire x_16232;
wire x_16233;
wire x_16234;
wire x_16235;
wire x_16236;
wire x_16237;
wire x_16238;
wire x_16239;
wire x_16240;
wire x_16241;
wire x_16242;
wire x_16243;
wire x_16244;
wire x_16245;
wire x_16246;
wire x_16247;
wire x_16248;
wire x_16249;
wire x_16250;
wire x_16251;
wire x_16252;
wire x_16253;
wire x_16254;
wire x_16255;
wire x_16256;
wire x_16257;
wire x_16258;
wire x_16259;
wire x_16260;
wire x_16261;
wire x_16262;
wire x_16263;
wire x_16264;
wire x_16265;
wire x_16266;
wire x_16267;
wire x_16268;
wire x_16269;
wire x_16270;
wire x_16271;
wire x_16272;
wire x_16273;
wire x_16274;
wire x_16275;
wire x_16276;
wire x_16277;
wire x_16278;
wire x_16279;
wire x_16280;
wire x_16281;
wire x_16282;
wire x_16283;
wire x_16284;
wire x_16285;
wire x_16286;
wire x_16287;
wire x_16288;
wire x_16289;
wire x_16290;
wire x_16291;
wire x_16292;
wire x_16293;
wire x_16294;
wire x_16295;
wire x_16296;
wire x_16297;
wire x_16298;
wire x_16299;
wire x_16300;
wire x_16301;
wire x_16302;
wire x_16303;
wire x_16304;
wire x_16305;
wire x_16306;
wire x_16307;
wire x_16308;
wire x_16309;
wire x_16310;
wire x_16311;
wire x_16312;
wire x_16313;
wire x_16314;
wire x_16315;
wire x_16316;
wire x_16317;
wire x_16318;
wire x_16319;
wire x_16320;
wire x_16321;
wire x_16322;
wire x_16323;
wire x_16324;
wire x_16325;
wire x_16326;
wire x_16327;
wire x_16328;
wire x_16329;
wire x_16330;
wire x_16331;
wire x_16332;
wire x_16333;
wire x_16334;
wire x_16335;
wire x_16336;
wire x_16337;
wire x_16338;
wire x_16339;
wire x_16340;
wire x_16341;
wire x_16342;
wire x_16343;
wire x_16344;
wire x_16345;
wire x_16346;
wire x_16347;
wire x_16348;
wire x_16349;
wire x_16350;
wire x_16351;
wire x_16352;
wire x_16353;
wire x_16354;
wire x_16355;
wire x_16356;
wire x_16357;
wire x_16358;
wire x_16359;
wire x_16360;
wire x_16361;
wire x_16362;
wire x_16363;
wire x_16364;
wire x_16365;
wire x_16366;
wire x_16367;
wire x_16368;
wire x_16369;
wire x_16370;
wire x_16371;
wire x_16372;
wire x_16373;
wire x_16374;
wire x_16375;
wire x_16376;
wire x_16377;
wire x_16378;
wire x_16379;
wire x_16380;
wire x_16381;
wire x_16382;
wire x_16383;
wire x_16384;
wire x_16385;
wire x_16386;
wire x_16387;
wire x_16388;
wire x_16389;
wire x_16390;
wire x_16391;
wire x_16392;
wire x_16393;
wire x_16394;
wire x_16395;
wire x_16396;
wire x_16397;
wire x_16398;
wire x_16399;
wire x_16400;
wire x_16401;
wire x_16402;
wire x_16403;
wire x_16404;
wire x_16405;
wire x_16406;
wire x_16407;
wire x_16408;
wire x_16409;
wire x_16410;
wire x_16411;
wire x_16412;
wire x_16413;
wire x_16414;
wire x_16415;
wire x_16416;
wire x_16417;
wire x_16418;
wire x_16419;
wire x_16420;
wire x_16421;
wire x_16422;
wire x_16423;
wire x_16424;
wire x_16425;
wire x_16426;
wire x_16427;
wire x_16428;
wire x_16429;
wire x_16430;
wire x_16431;
wire x_16432;
wire x_16433;
wire x_16434;
wire x_16435;
wire x_16436;
wire x_16437;
wire x_16438;
wire x_16439;
wire x_16440;
wire x_16441;
wire x_16442;
wire x_16443;
wire x_16444;
wire x_16445;
wire x_16446;
wire x_16447;
wire x_16448;
wire x_16449;
wire x_16450;
wire x_16451;
wire x_16452;
wire x_16453;
wire x_16454;
wire x_16455;
wire x_16456;
wire x_16457;
wire x_16458;
wire x_16459;
wire x_16460;
wire x_16461;
wire x_16462;
wire x_16463;
wire x_16464;
wire x_16465;
wire x_16466;
wire x_16467;
wire x_16468;
wire x_16469;
wire x_16470;
wire x_16471;
wire x_16472;
wire x_16473;
wire x_16474;
wire x_16475;
wire x_16476;
wire x_16477;
wire x_16478;
wire x_16479;
wire x_16480;
wire x_16481;
wire x_16482;
wire x_16483;
wire x_16484;
wire x_16485;
wire x_16486;
wire x_16487;
wire x_16488;
wire x_16489;
wire x_16490;
wire x_16491;
wire x_16492;
wire x_16493;
wire x_16494;
wire x_16495;
wire x_16496;
wire x_16497;
wire x_16498;
wire x_16499;
wire x_16500;
wire x_16501;
wire x_16502;
wire x_16503;
wire x_16504;
wire x_16505;
wire x_16506;
wire x_16507;
wire x_16508;
wire x_16509;
wire x_16510;
wire x_16511;
wire x_16512;
wire x_16513;
wire x_16514;
wire x_16515;
wire x_16516;
wire x_16517;
wire x_16518;
wire x_16519;
wire x_16520;
wire x_16521;
wire x_16522;
wire x_16523;
wire x_16524;
wire x_16525;
wire x_16526;
wire x_16527;
wire x_16528;
wire x_16529;
wire x_16530;
wire x_16531;
wire x_16532;
wire x_16533;
wire x_16534;
wire x_16535;
wire x_16536;
wire x_16537;
wire x_16538;
wire x_16539;
wire x_16540;
wire x_16541;
wire x_16542;
wire x_16543;
wire x_16544;
wire x_16545;
wire x_16546;
wire x_16547;
wire x_16548;
wire x_16549;
wire x_16550;
wire x_16551;
wire x_16552;
wire x_16553;
wire x_16554;
wire x_16555;
wire x_16556;
wire x_16557;
wire x_16558;
wire x_16559;
wire x_16560;
wire x_16561;
wire x_16562;
wire x_16563;
wire x_16564;
wire x_16565;
wire x_16566;
wire x_16567;
wire x_16568;
wire x_16569;
wire x_16570;
wire x_16571;
wire x_16572;
wire x_16573;
wire x_16574;
wire x_16575;
wire x_16576;
wire x_16577;
wire x_16578;
wire x_16579;
wire x_16580;
wire x_16581;
wire x_16582;
wire x_16583;
wire x_16584;
wire x_16585;
wire x_16586;
wire x_16587;
wire x_16588;
wire x_16589;
wire x_16590;
wire x_16591;
wire x_16592;
wire x_16593;
wire x_16594;
wire x_16595;
wire x_16596;
wire x_16597;
wire x_16598;
wire x_16599;
wire x_16600;
wire x_16601;
wire x_16602;
wire x_16603;
wire x_16604;
wire x_16605;
wire x_16606;
wire x_16607;
wire x_16608;
wire x_16609;
wire x_16610;
wire x_16611;
wire x_16612;
wire x_16613;
wire x_16614;
wire x_16615;
wire x_16616;
wire x_16617;
wire x_16618;
wire x_16619;
wire x_16620;
wire x_16621;
wire x_16622;
wire x_16623;
wire x_16624;
wire x_16625;
wire x_16626;
wire x_16627;
wire x_16628;
wire x_16629;
wire x_16630;
wire x_16631;
wire x_16632;
wire x_16633;
wire x_16634;
wire x_16635;
wire x_16636;
wire x_16637;
wire x_16638;
wire x_16639;
wire x_16640;
wire x_16641;
wire x_16642;
wire x_16643;
wire x_16644;
wire x_16645;
wire x_16646;
wire x_16647;
wire x_16648;
wire x_16649;
wire x_16650;
wire x_16651;
wire x_16652;
wire x_16653;
wire x_16654;
wire x_16655;
wire x_16656;
wire x_16657;
wire x_16658;
wire x_16659;
wire x_16660;
wire x_16661;
wire x_16662;
wire x_16663;
wire x_16664;
wire x_16665;
wire x_16666;
wire x_16667;
wire x_16668;
wire x_16669;
wire x_16670;
wire x_16671;
wire x_16672;
wire x_16673;
wire x_16674;
wire x_16675;
wire x_16676;
wire x_16677;
wire x_16678;
wire x_16679;
wire x_16680;
wire x_16681;
wire x_16682;
wire x_16683;
wire x_16684;
wire x_16685;
wire x_16686;
wire x_16687;
wire x_16688;
wire x_16689;
wire x_16690;
wire x_16691;
wire x_16692;
wire x_16693;
wire x_16694;
wire x_16695;
wire x_16696;
wire x_16697;
wire x_16698;
wire x_16699;
wire x_16700;
wire x_16701;
wire x_16702;
wire x_16703;
wire x_16704;
wire x_16705;
wire x_16706;
wire x_16707;
wire x_16708;
wire x_16709;
wire x_16710;
wire x_16711;
wire x_16712;
wire x_16713;
wire x_16714;
wire x_16715;
wire x_16716;
wire x_16717;
wire x_16718;
wire x_16719;
wire x_16720;
wire x_16721;
wire x_16722;
wire x_16723;
wire x_16724;
wire x_16725;
wire x_16726;
wire x_16727;
wire x_16728;
wire x_16729;
wire x_16730;
wire x_16731;
wire x_16732;
wire x_16733;
wire x_16734;
wire x_16735;
wire x_16736;
wire x_16737;
wire x_16738;
wire x_16739;
wire x_16740;
wire x_16741;
wire x_16742;
wire x_16743;
wire x_16744;
wire x_16745;
wire x_16746;
wire x_16747;
wire x_16748;
wire x_16749;
wire x_16750;
wire x_16751;
wire x_16752;
wire x_16753;
wire x_16754;
wire x_16755;
wire x_16756;
wire x_16757;
wire x_16758;
wire x_16759;
wire x_16760;
wire x_16761;
wire x_16762;
wire x_16763;
wire x_16764;
wire x_16765;
wire x_16766;
wire x_16767;
wire x_16768;
wire x_16769;
wire x_16770;
wire x_16771;
wire x_16772;
wire x_16773;
wire x_16774;
wire x_16775;
wire x_16776;
wire x_16777;
wire x_16778;
wire x_16779;
wire x_16780;
wire x_16781;
wire x_16782;
wire x_16783;
wire x_16784;
wire x_16785;
wire x_16786;
wire x_16787;
wire x_16788;
wire x_16789;
wire x_16790;
wire x_16791;
wire x_16792;
wire x_16793;
wire x_16794;
wire x_16795;
wire x_16796;
wire x_16797;
wire x_16798;
wire x_16799;
wire x_16800;
wire x_16801;
wire x_16802;
wire x_16803;
wire x_16804;
wire x_16805;
wire x_16806;
wire x_16807;
wire x_16808;
wire x_16809;
wire x_16810;
wire x_16811;
wire x_16812;
wire x_16813;
wire x_16814;
wire x_16815;
wire x_16816;
wire x_16817;
wire x_16818;
wire x_16819;
wire x_16820;
wire x_16821;
wire x_16822;
wire x_16823;
wire x_16824;
wire x_16825;
wire x_16826;
wire x_16827;
wire x_16828;
wire x_16829;
wire x_16830;
wire x_16831;
wire x_16832;
wire x_16833;
wire x_16834;
wire x_16835;
wire x_16836;
wire x_16837;
wire x_16838;
wire x_16839;
wire x_16840;
wire x_16841;
wire x_16842;
wire x_16843;
wire x_16844;
wire x_16845;
wire x_16846;
wire x_16847;
wire x_16848;
wire x_16849;
wire x_16850;
wire x_16851;
wire x_16852;
wire x_16853;
wire x_16854;
wire x_16855;
wire x_16856;
wire x_16857;
wire x_16858;
wire x_16859;
wire x_16860;
wire x_16861;
wire x_16862;
wire x_16863;
wire x_16864;
wire x_16865;
wire x_16866;
wire x_16867;
wire x_16868;
wire x_16869;
wire x_16870;
wire x_16871;
wire x_16872;
wire x_16873;
wire x_16874;
wire x_16875;
wire x_16876;
wire x_16877;
wire x_16878;
wire x_16879;
wire x_16880;
wire x_16881;
wire x_16882;
wire x_16883;
wire x_16884;
wire x_16885;
wire x_16886;
wire x_16887;
wire x_16888;
wire x_16889;
wire x_16890;
wire x_16891;
wire x_16892;
wire x_16893;
wire x_16894;
wire x_16895;
wire x_16896;
wire x_16897;
wire x_16898;
wire x_16899;
wire x_16900;
wire x_16901;
wire x_16902;
wire x_16903;
wire x_16904;
wire x_16905;
wire x_16906;
wire x_16907;
wire x_16908;
wire x_16909;
wire x_16910;
wire x_16911;
wire x_16912;
wire x_16913;
wire x_16914;
wire x_16915;
wire x_16916;
wire x_16917;
wire x_16918;
wire x_16919;
wire x_16920;
wire x_16921;
wire x_16922;
wire x_16923;
wire x_16924;
wire x_16925;
wire x_16926;
wire x_16927;
wire x_16928;
wire x_16929;
wire x_16930;
wire x_16931;
wire x_16932;
wire x_16933;
wire x_16934;
wire x_16935;
wire x_16936;
wire x_16937;
wire x_16938;
wire x_16939;
wire x_16940;
wire x_16941;
wire x_16942;
wire x_16943;
wire x_16944;
wire x_16945;
wire x_16946;
wire x_16947;
wire x_16948;
wire x_16949;
wire x_16950;
wire x_16951;
wire x_16952;
wire x_16953;
wire x_16954;
wire x_16955;
wire x_16956;
wire x_16957;
wire x_16958;
wire x_16959;
wire x_16960;
wire x_16961;
wire x_16962;
wire x_16963;
wire x_16964;
wire x_16965;
wire x_16966;
wire x_16967;
wire x_16968;
wire x_16969;
wire x_16970;
wire x_16971;
wire x_16972;
wire x_16973;
wire x_16974;
wire x_16975;
wire x_16976;
wire x_16977;
wire x_16978;
wire x_16979;
wire x_16980;
wire x_16981;
wire x_16982;
wire x_16983;
wire x_16984;
wire x_16985;
wire x_16986;
wire x_16987;
wire x_16988;
wire x_16989;
wire x_16990;
wire x_16991;
wire x_16992;
wire x_16993;
wire x_16994;
wire x_16995;
wire x_16996;
wire x_16997;
wire x_16998;
wire x_16999;
wire x_17000;
wire x_17001;
wire x_17002;
wire x_17003;
wire x_17004;
wire x_17005;
wire x_17006;
wire x_17007;
wire x_17008;
wire x_17009;
wire x_17010;
wire x_17011;
wire x_17012;
wire x_17013;
wire x_17014;
wire x_17015;
wire x_17016;
wire x_17017;
wire x_17018;
wire x_17019;
wire x_17020;
wire x_17021;
wire x_17022;
wire x_17023;
wire x_17024;
wire x_17025;
wire x_17026;
wire x_17027;
wire x_17028;
wire x_17029;
wire x_17030;
wire x_17031;
wire x_17032;
wire x_17033;
wire x_17034;
wire x_17035;
wire x_17036;
wire x_17037;
wire x_17038;
wire x_17039;
wire x_17040;
wire x_17041;
wire x_17042;
wire x_17043;
wire x_17044;
wire x_17045;
wire x_17046;
wire x_17047;
wire x_17048;
wire x_17049;
wire x_17050;
wire x_17051;
wire x_17052;
wire x_17053;
wire x_17054;
wire x_17055;
wire x_17056;
wire x_17057;
wire x_17058;
wire x_17059;
wire x_17060;
wire x_17061;
wire x_17062;
wire x_17063;
wire x_17064;
wire x_17065;
wire x_17066;
wire x_17067;
wire x_17068;
wire x_17069;
wire x_17070;
wire x_17071;
wire x_17072;
wire x_17073;
wire x_17074;
wire x_17075;
wire x_17076;
wire x_17077;
wire x_17078;
wire x_17079;
wire x_17080;
wire x_17081;
wire x_17082;
wire x_17083;
wire x_17084;
wire x_17085;
wire x_17086;
wire x_17087;
wire x_17088;
wire x_17089;
wire x_17090;
wire x_17091;
wire x_17092;
wire x_17093;
wire x_17094;
wire x_17095;
wire x_17096;
wire x_17097;
wire x_17098;
wire x_17099;
wire x_17100;
wire x_17101;
wire x_17102;
wire x_17103;
wire x_17104;
wire x_17105;
wire x_17106;
wire x_17107;
wire x_17108;
wire x_17109;
wire x_17110;
wire x_17111;
wire x_17112;
wire x_17113;
wire x_17114;
wire x_17115;
wire x_17116;
wire x_17117;
wire x_17118;
wire x_17119;
wire x_17120;
wire x_17121;
wire x_17122;
wire x_17123;
wire x_17124;
wire x_17125;
wire x_17126;
wire x_17127;
wire x_17128;
wire x_17129;
wire x_17130;
wire x_17131;
wire x_17132;
wire x_17133;
wire x_17134;
wire x_17135;
wire x_17136;
wire x_17137;
wire x_17138;
wire x_17139;
wire x_17140;
wire x_17141;
wire x_17142;
wire x_17143;
wire x_17144;
wire x_17145;
wire x_17146;
wire x_17147;
wire x_17148;
wire x_17149;
wire x_17150;
wire x_17151;
wire x_17152;
wire x_17153;
wire x_17154;
wire x_17155;
wire x_17156;
wire x_17157;
wire x_17158;
wire x_17159;
wire x_17160;
wire x_17161;
wire x_17162;
wire x_17163;
wire x_17164;
wire x_17165;
wire x_17166;
wire x_17167;
wire x_17168;
wire x_17169;
wire x_17170;
wire x_17171;
wire x_17172;
wire x_17173;
wire x_17174;
wire x_17175;
wire x_17176;
wire x_17177;
wire x_17178;
wire x_17179;
wire x_17180;
wire x_17181;
wire x_17182;
wire x_17183;
wire x_17184;
wire x_17185;
wire x_17186;
wire x_17187;
wire x_17188;
wire x_17189;
wire x_17190;
wire x_17191;
wire x_17192;
wire x_17193;
wire x_17194;
wire x_17195;
wire x_17196;
wire x_17197;
wire x_17198;
wire x_17199;
wire x_17200;
wire x_17201;
wire x_17202;
wire x_17203;
wire x_17204;
wire x_17205;
wire x_17206;
wire x_17207;
wire x_17208;
wire x_17209;
wire x_17210;
wire x_17211;
wire x_17212;
wire x_17213;
wire x_17214;
wire x_17215;
wire x_17216;
wire x_17217;
wire x_17218;
wire x_17219;
wire x_17220;
wire x_17221;
wire x_17222;
wire x_17223;
wire x_17224;
wire x_17225;
wire x_17226;
wire x_17227;
wire x_17228;
wire x_17229;
wire x_17230;
wire x_17231;
wire x_17232;
wire x_17233;
wire x_17234;
wire x_17235;
wire x_17236;
wire x_17237;
wire x_17238;
wire x_17239;
wire x_17240;
wire x_17241;
wire x_17242;
wire x_17243;
wire x_17244;
wire x_17245;
wire x_17246;
wire x_17247;
wire x_17248;
wire x_17249;
wire x_17250;
wire x_17251;
wire x_17252;
wire x_17253;
wire x_17254;
wire x_17255;
wire x_17256;
wire x_17257;
wire x_17258;
wire x_17259;
wire x_17260;
wire x_17261;
wire x_17262;
wire x_17263;
wire x_17264;
wire x_17265;
wire x_17266;
wire x_17267;
wire x_17268;
wire x_17269;
wire x_17270;
wire x_17271;
wire x_17272;
wire x_17273;
wire x_17274;
wire x_17275;
wire x_17276;
wire x_17277;
wire x_17278;
wire x_17279;
wire x_17280;
wire x_17281;
wire x_17282;
wire x_17283;
wire x_17284;
wire x_17285;
wire x_17286;
wire x_17287;
wire x_17288;
wire x_17289;
wire x_17290;
wire x_17291;
wire x_17292;
wire x_17293;
wire x_17294;
wire x_17295;
wire x_17296;
wire x_17297;
wire x_17298;
wire x_17299;
wire x_17300;
wire x_17301;
wire x_17302;
wire x_17303;
wire x_17304;
wire x_17305;
wire x_17306;
wire x_17307;
wire x_17308;
wire x_17309;
wire x_17310;
wire x_17311;
wire x_17312;
wire x_17313;
wire x_17314;
wire x_17315;
wire x_17316;
wire x_17317;
wire x_17318;
wire x_17319;
wire x_17320;
wire x_17321;
wire x_17322;
wire x_17323;
wire x_17324;
wire x_17325;
wire x_17326;
wire x_17327;
wire x_17328;
wire x_17329;
wire x_17330;
wire x_17331;
wire x_17332;
wire x_17333;
wire x_17334;
wire x_17335;
wire x_17336;
wire x_17337;
wire x_17338;
wire x_17339;
wire x_17340;
wire x_17341;
wire x_17342;
wire x_17343;
wire x_17344;
wire x_17345;
wire x_17346;
wire x_17347;
wire x_17348;
wire x_17349;
wire x_17350;
wire x_17351;
wire x_17352;
wire x_17353;
wire x_17354;
wire x_17355;
wire x_17356;
wire x_17357;
wire x_17358;
wire x_17359;
wire x_17360;
wire x_17361;
wire x_17362;
wire x_17363;
wire x_17364;
wire x_17365;
wire x_17366;
wire x_17367;
wire x_17368;
wire x_17369;
wire x_17370;
wire x_17371;
wire x_17372;
wire x_17373;
wire x_17374;
wire x_17375;
wire x_17376;
wire x_17377;
wire x_17378;
wire x_17379;
wire x_17380;
wire x_17381;
wire x_17382;
wire x_17383;
wire x_17384;
wire x_17385;
wire x_17386;
wire x_17387;
wire x_17388;
wire x_17389;
wire x_17390;
wire x_17391;
wire x_17392;
wire x_17393;
wire x_17394;
wire x_17395;
wire x_17396;
wire x_17397;
wire x_17398;
wire x_17399;
wire x_17400;
wire x_17401;
wire x_17402;
wire x_17403;
wire x_17404;
wire x_17405;
wire x_17406;
wire x_17407;
wire x_17408;
wire x_17409;
wire x_17410;
wire x_17411;
wire x_17412;
wire x_17413;
wire x_17414;
wire x_17415;
wire x_17416;
wire x_17417;
wire x_17418;
wire x_17419;
wire x_17420;
wire x_17421;
wire x_17422;
wire x_17423;
wire x_17424;
wire x_17425;
wire x_17426;
wire x_17427;
wire x_17428;
wire x_17429;
wire x_17430;
wire x_17431;
wire x_17432;
wire x_17433;
wire x_17434;
wire x_17435;
wire x_17436;
wire x_17437;
wire x_17438;
wire x_17439;
wire x_17440;
wire x_17441;
wire x_17442;
wire x_17443;
wire x_17444;
wire x_17445;
wire x_17446;
wire x_17447;
wire x_17448;
wire x_17449;
wire x_17450;
wire x_17451;
wire x_17452;
wire x_17453;
wire x_17454;
wire x_17455;
wire x_17456;
wire x_17457;
wire x_17458;
wire x_17459;
wire x_17460;
wire x_17461;
wire x_17462;
wire x_17463;
wire x_17464;
wire x_17465;
wire x_17466;
wire x_17467;
wire x_17468;
wire x_17469;
wire x_17470;
wire x_17471;
wire x_17472;
wire x_17473;
wire x_17474;
wire x_17475;
wire x_17476;
wire x_17477;
wire x_17478;
wire x_17479;
wire x_17480;
wire x_17481;
wire x_17482;
wire x_17483;
wire x_17484;
wire x_17485;
wire x_17486;
wire x_17487;
wire x_17488;
wire x_17489;
wire x_17490;
wire x_17491;
wire x_17492;
wire x_17493;
wire x_17494;
wire x_17495;
wire x_17496;
wire x_17497;
wire x_17498;
wire x_17499;
wire x_17500;
wire x_17501;
wire x_17502;
wire x_17503;
wire x_17504;
wire x_17505;
wire x_17506;
wire x_17507;
wire x_17508;
wire x_17509;
wire x_17510;
wire x_17511;
wire x_17512;
wire x_17513;
wire x_17514;
wire x_17515;
wire x_17516;
wire x_17517;
wire x_17518;
wire x_17519;
wire x_17520;
wire x_17521;
wire x_17522;
wire x_17523;
wire x_17524;
wire x_17525;
wire x_17526;
wire x_17527;
wire x_17528;
wire x_17529;
wire x_17530;
wire x_17531;
wire x_17532;
wire x_17533;
wire x_17534;
wire x_17535;
wire x_17536;
wire x_17537;
wire x_17538;
wire x_17539;
wire x_17540;
wire x_17541;
wire x_17542;
wire x_17543;
wire x_17544;
wire x_17545;
wire x_17546;
wire x_17547;
wire x_17548;
wire x_17549;
wire x_17550;
wire x_17551;
wire x_17552;
wire x_17553;
wire x_17554;
wire x_17555;
wire x_17556;
wire x_17557;
wire x_17558;
wire x_17559;
wire x_17560;
wire x_17561;
wire x_17562;
wire x_17563;
wire x_17564;
wire x_17565;
wire x_17566;
wire x_17567;
wire x_17568;
wire x_17569;
wire x_17570;
wire x_17571;
wire x_17572;
wire x_17573;
wire x_17574;
wire x_17575;
wire x_17576;
wire x_17577;
wire x_17578;
wire x_17579;
wire x_17580;
wire x_17581;
wire x_17582;
wire x_17583;
wire x_17584;
wire x_17585;
wire x_17586;
wire x_17587;
wire x_17588;
wire x_17589;
wire x_17590;
wire x_17591;
wire x_17592;
wire x_17593;
wire x_17594;
wire x_17595;
wire x_17596;
wire x_17597;
wire x_17598;
wire x_17599;
wire x_17600;
wire x_17601;
wire x_17602;
wire x_17603;
wire x_17604;
wire x_17605;
wire x_17606;
wire x_17607;
wire x_17608;
wire x_17609;
wire x_17610;
wire x_17611;
wire x_17612;
wire x_17613;
wire x_17614;
wire x_17615;
wire x_17616;
wire x_17617;
wire x_17618;
wire x_17619;
wire x_17620;
wire x_17621;
wire x_17622;
wire x_17623;
wire x_17624;
wire x_17625;
wire x_17626;
wire x_17627;
wire x_17628;
wire x_17629;
wire x_17630;
wire x_17631;
wire x_17632;
wire x_17633;
wire x_17634;
wire x_17635;
wire x_17636;
wire x_17637;
wire x_17638;
wire x_17639;
wire x_17640;
wire x_17641;
wire x_17642;
wire x_17643;
wire x_17644;
wire x_17645;
wire x_17646;
wire x_17647;
wire x_17648;
wire x_17649;
wire x_17650;
wire x_17651;
wire x_17652;
wire x_17653;
wire x_17654;
wire x_17655;
wire x_17656;
wire x_17657;
wire x_17658;
wire x_17659;
wire x_17660;
wire x_17661;
wire x_17662;
wire x_17663;
wire x_17664;
wire x_17665;
wire x_17666;
wire x_17667;
wire x_17668;
wire x_17669;
wire x_17670;
wire x_17671;
wire x_17672;
wire x_17673;
wire x_17674;
wire x_17675;
wire x_17676;
wire x_17677;
wire x_17678;
wire x_17679;
wire x_17680;
wire x_17681;
wire x_17682;
wire x_17683;
wire x_17684;
wire x_17685;
wire x_17686;
wire x_17687;
wire x_17688;
wire x_17689;
wire x_17690;
wire x_17691;
wire x_17692;
wire x_17693;
wire x_17694;
wire x_17695;
wire x_17696;
wire x_17697;
wire x_17698;
wire x_17699;
wire x_17700;
wire x_17701;
wire x_17702;
wire x_17703;
wire x_17704;
wire x_17705;
wire x_17706;
wire x_17707;
wire x_17708;
wire x_17709;
wire x_17710;
wire x_17711;
wire x_17712;
wire x_17713;
wire x_17714;
wire x_17715;
wire x_17716;
wire x_17717;
wire x_17718;
wire x_17719;
wire x_17720;
wire x_17721;
wire x_17722;
wire x_17723;
wire x_17724;
wire x_17725;
wire x_17726;
wire x_17727;
wire x_17728;
wire x_17729;
wire x_17730;
wire x_17731;
wire x_17732;
wire x_17733;
wire x_17734;
wire x_17735;
wire x_17736;
wire x_17737;
wire x_17738;
wire x_17739;
wire x_17740;
wire x_17741;
wire x_17742;
wire x_17743;
wire x_17744;
wire x_17745;
wire x_17746;
wire x_17747;
wire x_17748;
wire x_17749;
wire x_17750;
wire x_17751;
wire x_17752;
wire x_17753;
wire x_17754;
wire x_17755;
wire x_17756;
wire x_17757;
wire x_17758;
wire x_17759;
wire x_17760;
wire x_17761;
wire x_17762;
wire x_17763;
wire x_17764;
wire x_17765;
wire x_17766;
wire x_17767;
wire x_17768;
wire x_17769;
wire x_17770;
wire x_17771;
wire x_17772;
wire x_17773;
wire x_17774;
wire x_17775;
wire x_17776;
wire x_17777;
wire x_17778;
wire x_17779;
wire x_17780;
wire x_17781;
wire x_17782;
wire x_17783;
wire x_17784;
wire x_17785;
wire x_17786;
wire x_17787;
wire x_17788;
wire x_17789;
wire x_17790;
wire x_17791;
wire x_17792;
wire x_17793;
wire x_17794;
wire x_17795;
wire x_17796;
wire x_17797;
wire x_17798;
wire x_17799;
wire x_17800;
wire x_17801;
wire x_17802;
wire x_17803;
wire x_17804;
wire x_17805;
wire x_17806;
wire x_17807;
wire x_17808;
wire x_17809;
wire x_17810;
wire x_17811;
wire x_17812;
wire x_17813;
wire x_17814;
wire x_17815;
wire x_17816;
wire x_17817;
wire x_17818;
wire x_17819;
wire x_17820;
wire x_17821;
wire x_17822;
wire x_17823;
wire x_17824;
wire x_17825;
wire x_17826;
wire x_17827;
wire x_17828;
wire x_17829;
wire x_17830;
wire x_17831;
wire x_17832;
wire x_17833;
wire x_17834;
wire x_17835;
wire x_17836;
wire x_17837;
wire x_17838;
wire x_17839;
wire x_17840;
wire x_17841;
wire x_17842;
wire x_17843;
wire x_17844;
wire x_17845;
wire x_17846;
wire x_17847;
wire x_17848;
wire x_17849;
wire x_17850;
wire x_17851;
wire x_17852;
wire x_17853;
wire x_17854;
wire x_17855;
wire x_17856;
wire x_17857;
wire x_17858;
wire x_17859;
wire x_17860;
wire x_17861;
wire x_17862;
wire x_17863;
wire x_17864;
wire x_17865;
wire x_17866;
wire x_17867;
wire x_17868;
wire x_17869;
wire x_17870;
wire x_17871;
wire x_17872;
wire x_17873;
wire x_17874;
wire x_17875;
wire x_17876;
wire x_17877;
wire x_17878;
wire x_17879;
wire x_17880;
wire x_17881;
wire x_17882;
wire x_17883;
wire x_17884;
wire x_17885;
wire x_17886;
wire x_17887;
wire x_17888;
wire x_17889;
wire x_17890;
wire x_17891;
wire x_17892;
wire x_17893;
wire x_17894;
wire x_17895;
wire x_17896;
wire x_17897;
wire x_17898;
wire x_17899;
wire x_17900;
wire x_17901;
wire x_17902;
wire x_17903;
wire x_17904;
wire x_17905;
wire x_17906;
wire x_17907;
wire x_17908;
wire x_17909;
wire x_17910;
wire x_17911;
wire x_17912;
wire x_17913;
wire x_17914;
wire x_17915;
wire x_17916;
wire x_17917;
wire x_17918;
wire x_17919;
wire x_17920;
wire x_17921;
wire x_17922;
wire x_17923;
wire x_17924;
wire x_17925;
wire x_17926;
wire x_17927;
wire x_17928;
wire x_17929;
wire x_17930;
wire x_17931;
wire x_17932;
wire x_17933;
wire x_17934;
wire x_17935;
wire x_17936;
wire x_17937;
wire x_17938;
wire x_17939;
wire x_17940;
wire x_17941;
wire x_17942;
wire x_17943;
wire x_17944;
wire x_17945;
wire x_17946;
wire x_17947;
wire x_17948;
wire x_17949;
wire x_17950;
wire x_17951;
wire x_17952;
wire x_17953;
wire x_17954;
wire x_17955;
wire x_17956;
wire x_17957;
wire x_17958;
wire x_17959;
wire x_17960;
wire x_17961;
wire x_17962;
wire x_17963;
wire x_17964;
wire x_17965;
wire x_17966;
wire x_17967;
wire x_17968;
wire x_17969;
wire x_17970;
wire x_17971;
wire x_17972;
wire x_17973;
wire x_17974;
wire x_17975;
wire x_17976;
wire x_17977;
wire x_17978;
wire x_17979;
wire x_17980;
wire x_17981;
wire x_17982;
wire x_17983;
wire x_17984;
wire x_17985;
wire x_17986;
wire x_17987;
wire x_17988;
wire x_17989;
wire x_17990;
wire x_17991;
wire x_17992;
wire x_17993;
wire x_17994;
wire x_17995;
wire x_17996;
wire x_17997;
wire x_17998;
wire x_17999;
wire x_18000;
wire x_18001;
wire x_18002;
wire x_18003;
wire x_18004;
wire x_18005;
wire x_18006;
wire x_18007;
wire x_18008;
wire x_18009;
wire x_18010;
wire x_18011;
wire x_18012;
wire x_18013;
wire x_18014;
wire x_18015;
wire x_18016;
wire x_18017;
wire x_18018;
wire x_18019;
wire x_18020;
wire x_18021;
wire x_18022;
wire x_18023;
wire x_18024;
wire x_18025;
wire x_18026;
wire x_18027;
wire x_18028;
wire x_18029;
wire x_18030;
wire x_18031;
wire x_18032;
wire x_18033;
wire x_18034;
wire x_18035;
wire x_18036;
wire x_18037;
wire x_18038;
wire x_18039;
wire x_18040;
wire x_18041;
wire x_18042;
wire x_18043;
wire x_18044;
wire x_18045;
wire x_18046;
wire x_18047;
wire x_18048;
wire x_18049;
wire x_18050;
wire x_18051;
wire x_18052;
wire x_18053;
wire x_18054;
wire x_18055;
wire x_18056;
wire x_18057;
wire x_18058;
wire x_18059;
wire x_18060;
wire x_18061;
wire x_18062;
wire x_18063;
wire x_18064;
wire x_18065;
wire x_18066;
wire x_18067;
wire x_18068;
wire x_18069;
wire x_18070;
wire x_18071;
wire x_18072;
wire x_18073;
wire x_18074;
wire x_18075;
wire x_18076;
wire x_18077;
wire x_18078;
wire x_18079;
wire x_18080;
wire x_18081;
wire x_18082;
wire x_18083;
wire x_18084;
wire x_18085;
wire x_18086;
wire x_18087;
wire x_18088;
wire x_18089;
wire x_18090;
wire x_18091;
wire x_18092;
wire x_18093;
wire x_18094;
wire x_18095;
wire x_18096;
wire x_18097;
wire x_18098;
wire x_18099;
wire x_18100;
wire x_18101;
wire x_18102;
wire x_18103;
wire x_18104;
wire x_18105;
wire x_18106;
wire x_18107;
wire x_18108;
wire x_18109;
wire x_18110;
wire x_18111;
wire x_18112;
wire x_18113;
wire x_18114;
wire x_18115;
wire x_18116;
wire x_18117;
wire x_18118;
wire x_18119;
wire x_18120;
wire x_18121;
wire x_18122;
wire x_18123;
wire x_18124;
wire x_18125;
wire x_18126;
wire x_18127;
wire x_18128;
wire x_18129;
wire x_18130;
wire x_18131;
wire x_18132;
wire x_18133;
wire x_18134;
wire x_18135;
wire x_18136;
wire x_18137;
wire x_18138;
wire x_18139;
wire x_18140;
wire x_18141;
wire x_18142;
wire x_18143;
wire x_18144;
wire x_18145;
wire x_18146;
wire x_18147;
wire x_18148;
wire x_18149;
wire x_18150;
wire x_18151;
wire x_18152;
wire x_18153;
wire x_18154;
wire x_18155;
wire x_18156;
wire x_18157;
wire x_18158;
wire x_18159;
wire x_18160;
wire x_18161;
wire x_18162;
wire x_18163;
wire x_18164;
wire x_18165;
wire x_18166;
wire x_18167;
wire x_18168;
wire x_18169;
wire x_18170;
wire x_18171;
wire x_18172;
wire x_18173;
wire x_18174;
wire x_18175;
wire x_18176;
wire x_18177;
wire x_18178;
wire x_18179;
wire x_18180;
wire x_18181;
wire x_18182;
wire x_18183;
wire x_18184;
wire x_18185;
wire x_18186;
wire x_18187;
wire x_18188;
wire x_18189;
wire x_18190;
wire x_18191;
wire x_18192;
wire x_18193;
wire x_18194;
wire x_18195;
wire x_18196;
wire x_18197;
wire x_18198;
wire x_18199;
wire x_18200;
wire x_18201;
wire x_18202;
wire x_18203;
wire x_18204;
wire x_18205;
wire x_18206;
wire x_18207;
wire x_18208;
wire x_18209;
wire x_18210;
wire x_18211;
wire x_18212;
wire x_18213;
wire x_18214;
wire x_18215;
wire x_18216;
wire x_18217;
wire x_18218;
wire x_18219;
wire x_18220;
wire x_18221;
wire x_18222;
wire x_18223;
wire x_18224;
wire x_18225;
wire x_18226;
wire x_18227;
wire x_18228;
wire x_18229;
wire x_18230;
wire x_18231;
wire x_18232;
wire x_18233;
wire x_18234;
wire x_18235;
wire x_18236;
wire x_18237;
wire x_18238;
wire x_18239;
wire x_18240;
wire x_18241;
wire x_18242;
wire x_18243;
wire x_18244;
wire x_18245;
wire x_18246;
wire x_18247;
wire x_18248;
wire x_18249;
wire x_18250;
wire x_18251;
wire x_18252;
wire x_18253;
wire x_18254;
wire x_18255;
wire x_18256;
wire x_18257;
wire x_18258;
wire x_18259;
wire x_18260;
wire x_18261;
wire x_18262;
wire x_18263;
wire x_18264;
wire x_18265;
wire x_18266;
wire x_18267;
wire x_18268;
wire x_18269;
wire x_18270;
wire x_18271;
wire x_18272;
wire x_18273;
wire x_18274;
wire x_18275;
wire x_18276;
wire x_18277;
wire x_18278;
wire x_18279;
wire x_18280;
wire x_18281;
wire x_18282;
wire x_18283;
wire x_18284;
wire x_18285;
wire x_18286;
wire x_18287;
wire x_18288;
wire x_18289;
wire x_18290;
wire x_18291;
wire x_18292;
wire x_18293;
wire x_18294;
wire x_18295;
wire x_18296;
wire x_18297;
wire x_18298;
wire x_18299;
wire x_18300;
wire x_18301;
wire x_18302;
wire x_18303;
wire x_18304;
wire x_18305;
wire x_18306;
wire x_18307;
wire x_18308;
wire x_18309;
wire x_18310;
wire x_18311;
wire x_18312;
wire x_18313;
wire x_18314;
wire x_18315;
wire x_18316;
wire x_18317;
wire x_18318;
wire x_18319;
wire x_18320;
wire x_18321;
wire x_18322;
wire x_18323;
wire x_18324;
wire x_18325;
wire x_18326;
wire x_18327;
wire x_18328;
wire x_18329;
wire x_18330;
wire x_18331;
wire x_18332;
wire x_18333;
wire x_18334;
wire x_18335;
wire x_18336;
wire x_18337;
wire x_18338;
wire x_18339;
wire x_18340;
wire x_18341;
wire x_18342;
wire x_18343;
wire x_18344;
wire x_18345;
wire x_18346;
wire x_18347;
wire x_18348;
wire x_18349;
wire x_18350;
wire x_18351;
wire x_18352;
wire x_18353;
wire x_18354;
wire x_18355;
wire x_18356;
wire x_18357;
wire x_18358;
wire x_18359;
wire x_18360;
wire x_18361;
wire x_18362;
wire x_18363;
wire x_18364;
wire x_18365;
wire x_18366;
wire x_18367;
wire x_18368;
wire x_18369;
wire x_18370;
wire x_18371;
wire x_18372;
wire x_18373;
wire x_18374;
wire x_18375;
wire x_18376;
wire x_18377;
wire x_18378;
wire x_18379;
wire x_18380;
wire x_18381;
wire x_18382;
wire x_18383;
wire x_18384;
wire x_18385;
wire x_18386;
wire x_18387;
wire x_18388;
wire x_18389;
wire x_18390;
wire x_18391;
wire x_18392;
wire x_18393;
wire x_18394;
wire x_18395;
wire x_18396;
wire x_18397;
wire x_18398;
wire x_18399;
wire x_18400;
wire x_18401;
wire x_18402;
wire x_18403;
wire x_18404;
wire x_18405;
wire x_18406;
wire x_18407;
wire x_18408;
wire x_18409;
wire x_18410;
wire x_18411;
wire x_18412;
wire x_18413;
wire x_18414;
wire x_18415;
wire x_18416;
wire x_18417;
wire x_18418;
wire x_18419;
wire x_18420;
wire x_18421;
wire x_18422;
wire x_18423;
wire x_18424;
wire x_18425;
wire x_18426;
wire x_18427;
wire x_18428;
wire x_18429;
wire x_18430;
wire x_18431;
wire x_18432;
wire x_18433;
wire x_18434;
wire x_18435;
wire x_18436;
wire x_18437;
wire x_18438;
wire x_18439;
wire x_18440;
wire x_18441;
wire x_18442;
wire x_18443;
wire x_18444;
wire x_18445;
wire x_18446;
wire x_18447;
wire x_18448;
wire x_18449;
wire x_18450;
wire x_18451;
wire x_18452;
wire x_18453;
wire x_18454;
wire x_18455;
wire x_18456;
wire x_18457;
wire x_18458;
wire x_18459;
wire x_18460;
wire x_18461;
wire x_18462;
wire x_18463;
wire x_18464;
wire x_18465;
wire x_18466;
wire x_18467;
wire x_18468;
wire x_18469;
wire x_18470;
wire x_18471;
wire x_18472;
wire x_18473;
wire x_18474;
wire x_18475;
wire x_18476;
wire x_18477;
wire x_18478;
wire x_18479;
wire x_18480;
wire x_18481;
wire x_18482;
wire x_18483;
wire x_18484;
wire x_18485;
wire x_18486;
wire x_18487;
wire x_18488;
wire x_18489;
wire x_18490;
wire x_18491;
wire x_18492;
wire x_18493;
wire x_18494;
wire x_18495;
wire x_18496;
wire x_18497;
wire x_18498;
wire x_18499;
wire x_18500;
wire x_18501;
wire x_18502;
wire x_18503;
wire x_18504;
wire x_18505;
wire x_18506;
wire x_18507;
wire x_18508;
wire x_18509;
wire x_18510;
wire x_18511;
wire x_18512;
wire x_18513;
wire x_18514;
wire x_18515;
wire x_18516;
wire x_18517;
wire x_18518;
wire x_18519;
wire x_18520;
wire x_18521;
wire x_18522;
wire x_18523;
wire x_18524;
wire x_18525;
wire x_18526;
wire x_18527;
wire x_18528;
wire x_18529;
wire x_18530;
wire x_18531;
wire x_18532;
wire x_18533;
wire x_18534;
wire x_18535;
wire x_18536;
wire x_18537;
wire x_18538;
wire x_18539;
wire x_18540;
wire x_18541;
wire x_18542;
wire x_18543;
wire x_18544;
wire x_18545;
wire x_18546;
wire x_18547;
wire x_18548;
wire x_18549;
wire x_18550;
wire x_18551;
wire x_18552;
wire x_18553;
wire x_18554;
wire x_18555;
wire x_18556;
wire x_18557;
wire x_18558;
wire x_18559;
wire x_18560;
wire x_18561;
wire x_18562;
wire x_18563;
wire x_18564;
wire x_18565;
wire x_18566;
wire x_18567;
wire x_18568;
wire x_18569;
wire x_18570;
wire x_18571;
wire x_18572;
wire x_18573;
wire x_18574;
wire x_18575;
wire x_18576;
wire x_18577;
wire x_18578;
wire x_18579;
wire x_18580;
wire x_18581;
wire x_18582;
wire x_18583;
wire x_18584;
wire x_18585;
wire x_18586;
wire x_18587;
wire x_18588;
wire x_18589;
wire x_18590;
wire x_18591;
wire x_18592;
wire x_18593;
wire x_18594;
wire x_18595;
wire x_18596;
wire x_18597;
wire x_18598;
wire x_18599;
wire x_18600;
wire x_18601;
wire x_18602;
wire x_18603;
wire x_18604;
wire x_18605;
wire x_18606;
wire x_18607;
wire x_18608;
wire x_18609;
wire x_18610;
wire x_18611;
wire x_18612;
wire x_18613;
wire x_18614;
wire x_18615;
wire x_18616;
wire x_18617;
wire x_18618;
wire x_18619;
wire x_18620;
wire x_18621;
wire x_18622;
wire x_18623;
wire x_18624;
wire x_18625;
wire x_18626;
wire x_18627;
wire x_18628;
wire x_18629;
wire x_18630;
wire x_18631;
wire x_18632;
wire x_18633;
wire x_18634;
wire x_18635;
wire x_18636;
wire x_18637;
wire x_18638;
wire x_18639;
wire x_18640;
wire x_18641;
wire x_18642;
wire x_18643;
wire x_18644;
wire x_18645;
wire x_18646;
wire x_18647;
wire x_18648;
wire x_18649;
wire x_18650;
wire x_18651;
wire x_18652;
wire x_18653;
wire x_18654;
wire x_18655;
wire x_18656;
wire x_18657;
wire x_18658;
wire x_18659;
wire x_18660;
wire x_18661;
wire x_18662;
wire x_18663;
wire x_18664;
wire x_18665;
wire x_18666;
wire x_18667;
wire x_18668;
wire x_18669;
wire x_18670;
wire x_18671;
wire x_18672;
wire x_18673;
wire x_18674;
wire x_18675;
wire x_18676;
wire x_18677;
wire x_18678;
wire x_18679;
wire x_18680;
wire x_18681;
wire x_18682;
wire x_18683;
wire x_18684;
wire x_18685;
wire x_18686;
wire x_18687;
wire x_18688;
wire x_18689;
wire x_18690;
wire x_18691;
wire x_18692;
wire x_18693;
wire x_18694;
wire x_18695;
wire x_18696;
wire x_18697;
wire x_18698;
wire x_18699;
wire x_18700;
wire x_18701;
wire x_18702;
wire x_18703;
wire x_18704;
wire x_18705;
wire x_18706;
wire x_18707;
wire x_18708;
wire x_18709;
wire x_18710;
wire x_18711;
wire x_18712;
wire x_18713;
wire x_18714;
wire x_18715;
wire x_18716;
wire x_18717;
wire x_18718;
wire x_18719;
wire x_18720;
wire x_18721;
wire x_18722;
wire x_18723;
wire x_18724;
wire x_18725;
wire x_18726;
wire x_18727;
wire x_18728;
wire x_18729;
wire x_18730;
wire x_18731;
wire x_18732;
wire x_18733;
wire x_18734;
wire x_18735;
wire x_18736;
wire x_18737;
wire x_18738;
wire x_18739;
wire x_18740;
wire x_18741;
wire x_18742;
wire x_18743;
wire x_18744;
wire x_18745;
wire x_18746;
wire x_18747;
wire x_18748;
wire x_18749;
wire x_18750;
wire x_18751;
wire x_18752;
wire x_18753;
wire x_18754;
wire x_18755;
wire x_18756;
wire x_18757;
wire x_18758;
wire x_18759;
wire x_18760;
wire x_18761;
wire x_18762;
wire x_18763;
wire x_18764;
wire x_18765;
wire x_18766;
wire x_18767;
wire x_18768;
wire x_18769;
wire x_18770;
wire x_18771;
wire x_18772;
wire x_18773;
wire x_18774;
wire x_18775;
wire x_18776;
wire x_18777;
wire x_18778;
wire x_18779;
wire x_18780;
wire x_18781;
wire x_18782;
wire x_18783;
wire x_18784;
wire x_18785;
wire x_18786;
wire x_18787;
wire x_18788;
wire x_18789;
wire x_18790;
wire x_18791;
wire x_18792;
wire x_18793;
wire x_18794;
wire x_18795;
wire x_18796;
wire x_18797;
wire x_18798;
wire x_18799;
wire x_18800;
wire x_18801;
wire x_18802;
wire x_18803;
wire x_18804;
wire x_18805;
wire x_18806;
wire x_18807;
wire x_18808;
wire x_18809;
wire x_18810;
wire x_18811;
wire x_18812;
wire x_18813;
wire x_18814;
wire x_18815;
wire x_18816;
wire x_18817;
wire x_18818;
wire x_18819;
wire x_18820;
wire x_18821;
wire x_18822;
wire x_18823;
wire x_18824;
wire x_18825;
wire x_18826;
wire x_18827;
wire x_18828;
wire x_18829;
wire x_18830;
wire x_18831;
wire x_18832;
wire x_18833;
wire x_18834;
wire x_18835;
wire x_18836;
wire x_18837;
wire x_18838;
wire x_18839;
wire x_18840;
wire x_18841;
wire x_18842;
wire x_18843;
wire x_18844;
wire x_18845;
wire x_18846;
wire x_18847;
wire x_18848;
wire x_18849;
wire x_18850;
wire x_18851;
wire x_18852;
wire x_18853;
wire x_18854;
wire x_18855;
wire x_18856;
wire x_18857;
wire x_18858;
wire x_18859;
wire x_18860;
wire x_18861;
wire x_18862;
wire x_18863;
wire x_18864;
wire x_18865;
wire x_18866;
wire x_18867;
wire x_18868;
wire x_18869;
wire x_18870;
wire x_18871;
wire x_18872;
wire x_18873;
wire x_18874;
wire x_18875;
wire x_18876;
wire x_18877;
wire x_18878;
wire x_18879;
wire x_18880;
wire x_18881;
wire x_18882;
wire x_18883;
wire x_18884;
wire x_18885;
wire x_18886;
wire x_18887;
wire x_18888;
wire x_18889;
wire x_18890;
wire x_18891;
wire x_18892;
wire x_18893;
wire x_18894;
wire x_18895;
wire x_18896;
wire x_18897;
wire x_18898;
wire x_18899;
wire x_18900;
wire x_18901;
wire x_18902;
wire x_18903;
wire x_18904;
wire x_18905;
wire x_18906;
wire x_18907;
wire x_18908;
wire x_18909;
wire x_18910;
wire x_18911;
wire x_18912;
wire x_18913;
wire x_18914;
wire x_18915;
wire x_18916;
wire x_18917;
wire x_18918;
wire x_18919;
wire x_18920;
wire x_18921;
wire x_18922;
wire x_18923;
wire x_18924;
wire x_18925;
wire x_18926;
wire x_18927;
wire x_18928;
wire x_18929;
wire x_18930;
wire x_18931;
wire x_18932;
wire x_18933;
wire x_18934;
wire x_18935;
wire x_18936;
wire x_18937;
wire x_18938;
wire x_18939;
wire x_18940;
wire x_18941;
wire x_18942;
wire x_18943;
wire x_18944;
wire x_18945;
wire x_18946;
wire x_18947;
wire x_18948;
wire x_18949;
wire x_18950;
wire x_18951;
wire x_18952;
wire x_18953;
wire x_18954;
wire x_18955;
wire x_18956;
wire x_18957;
wire x_18958;
wire x_18959;
wire x_18960;
wire x_18961;
wire x_18962;
wire x_18963;
wire x_18964;
wire x_18965;
wire x_18966;
wire x_18967;
wire x_18968;
wire x_18969;
wire x_18970;
wire x_18971;
wire x_18972;
wire x_18973;
wire x_18974;
wire x_18975;
wire x_18976;
wire x_18977;
wire x_18978;
wire x_18979;
wire x_18980;
wire x_18981;
wire x_18982;
wire x_18983;
wire x_18984;
wire x_18985;
wire x_18986;
wire x_18987;
wire x_18988;
wire x_18989;
wire x_18990;
wire x_18991;
wire x_18992;
wire x_18993;
wire x_18994;
wire x_18995;
wire x_18996;
wire x_18997;
wire x_18998;
wire x_18999;
wire x_19000;
wire x_19001;
wire x_19002;
wire x_19003;
wire x_19004;
wire x_19005;
wire x_19006;
wire x_19007;
wire x_19008;
wire x_19009;
wire x_19010;
wire x_19011;
wire x_19012;
wire x_19013;
wire x_19014;
wire x_19015;
wire x_19016;
wire x_19017;
wire x_19018;
wire x_19019;
wire x_19020;
wire x_19021;
wire x_19022;
wire x_19023;
wire x_19024;
wire x_19025;
wire x_19026;
wire x_19027;
wire x_19028;
wire x_19029;
wire x_19030;
wire x_19031;
wire x_19032;
wire x_19033;
wire x_19034;
wire x_19035;
wire x_19036;
wire x_19037;
wire x_19038;
wire x_19039;
wire x_19040;
wire x_19041;
wire x_19042;
wire x_19043;
wire x_19044;
wire x_19045;
wire x_19046;
wire x_19047;
wire x_19048;
wire x_19049;
wire x_19050;
wire x_19051;
wire x_19052;
wire x_19053;
wire x_19054;
wire x_19055;
wire x_19056;
wire x_19057;
wire x_19058;
wire x_19059;
wire x_19060;
wire x_19061;
wire x_19062;
wire x_19063;
wire x_19064;
wire x_19065;
wire x_19066;
wire x_19067;
wire x_19068;
wire x_19069;
wire x_19070;
wire x_19071;
wire x_19072;
wire x_19073;
wire x_19074;
wire x_19075;
wire x_19076;
wire x_19077;
wire x_19078;
wire x_19079;
wire x_19080;
wire x_19081;
wire x_19082;
wire x_19083;
wire x_19084;
wire x_19085;
wire x_19086;
wire x_19087;
wire x_19088;
wire x_19089;
wire x_19090;
wire x_19091;
wire x_19092;
wire x_19093;
wire x_19094;
wire x_19095;
wire x_19096;
wire x_19097;
wire x_19098;
wire x_19099;
wire x_19100;
wire x_19101;
wire x_19102;
wire x_19103;
wire x_19104;
wire x_19105;
wire x_19106;
wire x_19107;
wire x_19108;
wire x_19109;
wire x_19110;
wire x_19111;
wire x_19112;
wire x_19113;
wire x_19114;
wire x_19115;
wire x_19116;
wire x_19117;
wire x_19118;
wire x_19119;
wire x_19120;
wire x_19121;
wire x_19122;
wire x_19123;
wire x_19124;
wire x_19125;
wire x_19126;
wire x_19127;
wire x_19128;
wire x_19129;
wire x_19130;
wire x_19131;
wire x_19132;
wire x_19133;
wire x_19134;
wire x_19135;
wire x_19136;
wire x_19137;
wire x_19138;
wire x_19139;
wire x_19140;
wire x_19141;
wire x_19142;
wire x_19143;
wire x_19144;
wire x_19145;
wire x_19146;
wire x_19147;
wire x_19148;
wire x_19149;
wire x_19150;
wire x_19151;
wire x_19152;
wire x_19153;
wire x_19154;
wire x_19155;
wire x_19156;
wire x_19157;
wire x_19158;
wire x_19159;
wire x_19160;
wire x_19161;
wire x_19162;
wire x_19163;
wire x_19164;
wire x_19165;
wire x_19166;
wire x_19167;
wire x_19168;
wire x_19169;
wire x_19170;
wire x_19171;
wire x_19172;
wire x_19173;
wire x_19174;
wire x_19175;
wire x_19176;
wire x_19177;
wire x_19178;
wire x_19179;
wire x_19180;
wire x_19181;
wire x_19182;
wire x_19183;
wire x_19184;
wire x_19185;
wire x_19186;
wire x_19187;
wire x_19188;
wire x_19189;
wire x_19190;
wire x_19191;
wire x_19192;
wire x_19193;
wire x_19194;
wire x_19195;
wire x_19196;
wire x_19197;
wire x_19198;
wire x_19199;
wire x_19200;
wire x_19201;
wire x_19202;
wire x_19203;
wire x_19204;
wire x_19205;
wire x_19206;
wire x_19207;
wire x_19208;
wire x_19209;
wire x_19210;
wire x_19211;
wire x_19212;
wire x_19213;
wire x_19214;
wire x_19215;
wire x_19216;
wire x_19217;
wire x_19218;
wire x_19219;
wire x_19220;
wire x_19221;
wire x_19222;
wire x_19223;
wire x_19224;
wire x_19225;
wire x_19226;
wire x_19227;
wire x_19228;
wire x_19229;
wire x_19230;
wire x_19231;
wire x_19232;
wire x_19233;
wire x_19234;
wire x_19235;
wire x_19236;
wire x_19237;
wire x_19238;
wire x_19239;
wire x_19240;
wire x_19241;
wire x_19242;
wire x_19243;
wire x_19244;
wire x_19245;
wire x_19246;
wire x_19247;
wire x_19248;
wire x_19249;
wire x_19250;
wire x_19251;
wire x_19252;
wire x_19253;
wire x_19254;
wire x_19255;
wire x_19256;
wire x_19257;
wire x_19258;
wire x_19259;
wire x_19260;
wire x_19261;
wire x_19262;
wire x_19263;
wire x_19264;
wire x_19265;
wire x_19266;
wire x_19267;
wire x_19268;
wire x_19269;
wire x_19270;
wire x_19271;
wire x_19272;
wire x_19273;
wire x_19274;
wire x_19275;
wire x_19276;
wire x_19277;
wire x_19278;
wire x_19279;
wire x_19280;
wire x_19281;
wire x_19282;
wire x_19283;
wire x_19284;
wire x_19285;
wire x_19286;
wire x_19287;
wire x_19288;
wire x_19289;
wire x_19290;
wire x_19291;
wire x_19292;
wire x_19293;
wire x_19294;
wire x_19295;
wire x_19296;
wire x_19297;
wire x_19298;
wire x_19299;
wire x_19300;
wire x_19301;
wire x_19302;
wire x_19303;
wire x_19304;
wire x_19305;
wire x_19306;
wire x_19307;
wire x_19308;
wire x_19309;
wire x_19310;
wire x_19311;
wire x_19312;
wire x_19313;
wire x_19314;
wire x_19315;
wire x_19316;
wire x_19317;
wire x_19318;
wire x_19319;
wire x_19320;
wire x_19321;
wire x_19322;
wire x_19323;
wire x_19324;
wire x_19325;
wire x_19326;
wire x_19327;
wire x_19328;
wire x_19329;
wire x_19330;
wire x_19331;
wire x_19332;
wire x_19333;
wire x_19334;
wire x_19335;
wire x_19336;
wire x_19337;
wire x_19338;
wire x_19339;
wire x_19340;
wire x_19341;
wire x_19342;
wire x_19343;
wire x_19344;
wire x_19345;
wire x_19346;
wire x_19347;
wire x_19348;
wire x_19349;
wire x_19350;
wire x_19351;
wire x_19352;
wire x_19353;
wire x_19354;
wire x_19355;
wire x_19356;
wire x_19357;
wire x_19358;
wire x_19359;
wire x_19360;
wire x_19361;
wire x_19362;
wire x_19363;
wire x_19364;
wire x_19365;
wire x_19366;
wire x_19367;
wire x_19368;
wire x_19369;
wire x_19370;
wire x_19371;
wire x_19372;
wire x_19373;
wire x_19374;
wire x_19375;
wire x_19376;
wire x_19377;
wire x_19378;
wire x_19379;
wire x_19380;
wire x_19381;
wire x_19382;
wire x_19383;
wire x_19384;
wire x_19385;
wire x_19386;
wire x_19387;
wire x_19388;
wire x_19389;
wire x_19390;
wire x_19391;
wire x_19392;
wire x_19393;
wire x_19394;
wire x_19395;
wire x_19396;
wire x_19397;
wire x_19398;
wire x_19399;
wire x_19400;
wire x_19401;
wire x_19402;
wire x_19403;
wire x_19404;
wire x_19405;
wire x_19406;
wire x_19407;
wire x_19408;
wire x_19409;
wire x_19410;
wire x_19411;
wire x_19412;
wire x_19413;
wire x_19414;
wire x_19415;
wire x_19416;
wire x_19417;
wire x_19418;
wire x_19419;
wire x_19420;
wire x_19421;
wire x_19422;
wire x_19423;
wire x_19424;
wire x_19425;
wire x_19426;
wire x_19427;
wire x_19428;
wire x_19429;
wire x_19430;
wire x_19431;
wire x_19432;
wire x_19433;
wire x_19434;
wire x_19435;
wire x_19436;
wire x_19437;
wire x_19438;
wire x_19439;
wire x_19440;
wire x_19441;
wire x_19442;
wire x_19443;
wire x_19444;
wire x_19445;
wire x_19446;
wire x_19447;
wire x_19448;
wire x_19449;
wire x_19450;
wire x_19451;
wire x_19452;
wire x_19453;
wire x_19454;
wire x_19455;
wire x_19456;
wire x_19457;
wire x_19458;
wire x_19459;
wire x_19460;
wire x_19461;
wire x_19462;
wire x_19463;
wire x_19464;
wire x_19465;
wire x_19466;
wire x_19467;
wire x_19468;
wire x_19469;
wire x_19470;
wire x_19471;
wire x_19472;
wire x_19473;
wire x_19474;
wire x_19475;
wire x_19476;
wire x_19477;
wire x_19478;
wire x_19479;
wire x_19480;
wire x_19481;
wire x_19482;
wire x_19483;
wire x_19484;
wire x_19485;
wire x_19486;
wire x_19487;
wire x_19488;
wire x_19489;
wire x_19490;
wire x_19491;
wire x_19492;
wire x_19493;
wire x_19494;
wire x_19495;
wire x_19496;
wire x_19497;
wire x_19498;
wire x_19499;
wire x_19500;
wire x_19501;
wire x_19502;
wire x_19503;
wire x_19504;
wire x_19505;
wire x_19506;
wire x_19507;
wire x_19508;
wire x_19509;
wire x_19510;
wire x_19511;
wire x_19512;
wire x_19513;
wire x_19514;
wire x_19515;
wire x_19516;
wire x_19517;
wire x_19518;
wire x_19519;
wire x_19520;
wire x_19521;
wire x_19522;
wire x_19523;
wire x_19524;
wire x_19525;
wire x_19526;
wire x_19527;
wire x_19528;
wire x_19529;
wire x_19530;
wire x_19531;
wire x_19532;
wire x_19533;
wire x_19534;
wire x_19535;
wire x_19536;
wire x_19537;
wire x_19538;
wire x_19539;
wire x_19540;
wire x_19541;
wire x_19542;
wire x_19543;
wire x_19544;
wire x_19545;
wire x_19546;
wire x_19547;
wire x_19548;
wire x_19549;
wire x_19550;
wire x_19551;
wire x_19552;
wire x_19553;
wire x_19554;
wire x_19555;
wire x_19556;
wire x_19557;
wire x_19558;
wire x_19559;
wire x_19560;
wire x_19561;
wire x_19562;
wire x_19563;
wire x_19564;
wire x_19565;
wire x_19566;
wire x_19567;
wire x_19568;
wire x_19569;
wire x_19570;
wire x_19571;
wire x_19572;
wire x_19573;
wire x_19574;
wire x_19575;
wire x_19576;
wire x_19577;
wire x_19578;
wire x_19579;
wire x_19580;
wire x_19581;
wire x_19582;
wire x_19583;
wire x_19584;
wire x_19585;
wire x_19586;
wire x_19587;
wire x_19588;
wire x_19589;
wire x_19590;
wire x_19591;
wire x_19592;
wire x_19593;
wire x_19594;
wire x_19595;
wire x_19596;
wire x_19597;
wire x_19598;
wire x_19599;
wire x_19600;
wire x_19601;
wire x_19602;
wire x_19603;
wire x_19604;
wire x_19605;
wire x_19606;
wire x_19607;
wire x_19608;
wire x_19609;
wire x_19610;
wire x_19611;
wire x_19612;
wire x_19613;
wire x_19614;
wire x_19615;
wire x_19616;
wire x_19617;
wire x_19618;
wire x_19619;
wire x_19620;
wire x_19621;
wire x_19622;
wire x_19623;
wire x_19624;
wire x_19625;
wire x_19626;
wire x_19627;
wire x_19628;
wire x_19629;
wire x_19630;
wire x_19631;
wire x_19632;
wire x_19633;
wire x_19634;
wire x_19635;
wire x_19636;
wire x_19637;
wire x_19638;
wire x_19639;
wire x_19640;
wire x_19641;
wire x_19642;
wire x_19643;
wire x_19644;
wire x_19645;
wire x_19646;
wire x_19647;
wire x_19648;
wire x_19649;
wire x_19650;
wire x_19651;
wire x_19652;
wire x_19653;
wire x_19654;
wire x_19655;
wire x_19656;
wire x_19657;
wire x_19658;
wire x_19659;
wire x_19660;
wire x_19661;
wire x_19662;
wire x_19663;
wire x_19664;
wire x_19665;
wire x_19666;
wire x_19667;
wire x_19668;
wire x_19669;
wire x_19670;
wire x_19671;
wire x_19672;
wire x_19673;
wire x_19674;
wire x_19675;
wire x_19676;
wire x_19677;
wire x_19678;
wire x_19679;
wire x_19680;
wire x_19681;
wire x_19682;
wire x_19683;
wire x_19684;
wire x_19685;
wire x_19686;
wire x_19687;
wire x_19688;
wire x_19689;
wire x_19690;
wire x_19691;
wire x_19692;
wire x_19693;
wire x_19694;
wire x_19695;
wire x_19696;
wire x_19697;
wire x_19698;
wire x_19699;
wire x_19700;
wire x_19701;
wire x_19702;
wire x_19703;
wire x_19704;
wire x_19705;
wire x_19706;
wire x_19707;
wire x_19708;
wire x_19709;
wire x_19710;
wire x_19711;
wire x_19712;
wire x_19713;
wire x_19714;
wire x_19715;
wire x_19716;
wire x_19717;
wire x_19718;
wire x_19719;
wire x_19720;
wire x_19721;
wire x_19722;
wire x_19723;
wire x_19724;
wire x_19725;
wire x_19726;
wire x_19727;
wire x_19728;
wire x_19729;
wire x_19730;
wire x_19731;
wire x_19732;
wire x_19733;
wire x_19734;
wire x_19735;
wire x_19736;
wire x_19737;
wire x_19738;
wire x_19739;
wire x_19740;
wire x_19741;
wire x_19742;
wire x_19743;
wire x_19744;
wire x_19745;
wire x_19746;
wire x_19747;
wire x_19748;
wire x_19749;
wire x_19750;
wire x_19751;
wire x_19752;
wire x_19753;
wire x_19754;
wire x_19755;
wire x_19756;
wire x_19757;
wire x_19758;
wire x_19759;
wire x_19760;
wire x_19761;
wire x_19762;
wire x_19763;
wire x_19764;
wire x_19765;
wire x_19766;
wire x_19767;
wire x_19768;
wire x_19769;
wire x_19770;
wire x_19771;
wire x_19772;
wire x_19773;
wire x_19774;
wire x_19775;
wire x_19776;
wire x_19777;
wire x_19778;
wire x_19779;
wire x_19780;
wire x_19781;
wire x_19782;
wire x_19783;
wire x_19784;
wire x_19785;
wire x_19786;
wire x_19787;
wire x_19788;
wire x_19789;
wire x_19790;
wire x_19791;
wire x_19792;
wire x_19793;
wire x_19794;
wire x_19795;
wire x_19796;
wire x_19797;
wire x_19798;
wire x_19799;
wire x_19800;
wire x_19801;
wire x_19802;
wire x_19803;
wire x_19804;
wire x_19805;
wire x_19806;
wire x_19807;
wire x_19808;
wire x_19809;
wire x_19810;
wire x_19811;
wire x_19812;
wire x_19813;
wire x_19814;
wire x_19815;
wire x_19816;
wire x_19817;
wire x_19818;
wire x_19819;
wire x_19820;
wire x_19821;
wire x_19822;
wire x_19823;
wire x_19824;
wire x_19825;
wire x_19826;
wire x_19827;
wire x_19828;
wire x_19829;
wire x_19830;
wire x_19831;
wire x_19832;
wire x_19833;
wire x_19834;
wire x_19835;
wire x_19836;
wire x_19837;
wire x_19838;
wire x_19839;
wire x_19840;
wire x_19841;
wire x_19842;
wire x_19843;
wire x_19844;
wire x_19845;
wire x_19846;
wire x_19847;
wire x_19848;
wire x_19849;
wire x_19850;
wire x_19851;
wire x_19852;
wire x_19853;
wire x_19854;
wire x_19855;
wire x_19856;
wire x_19857;
wire x_19858;
wire x_19859;
wire x_19860;
wire x_19861;
wire x_19862;
wire x_19863;
wire x_19864;
wire x_19865;
wire x_19866;
wire x_19867;
wire x_19868;
wire x_19869;
wire x_19870;
wire x_19871;
wire x_19872;
wire x_19873;
wire x_19874;
wire x_19875;
wire x_19876;
wire x_19877;
wire x_19878;
wire x_19879;
wire x_19880;
wire x_19881;
wire x_19882;
wire x_19883;
wire x_19884;
wire x_19885;
wire x_19886;
wire x_19887;
wire x_19888;
wire x_19889;
wire x_19890;
wire x_19891;
wire x_19892;
wire x_19893;
wire x_19894;
wire x_19895;
wire x_19896;
wire x_19897;
wire x_19898;
wire x_19899;
wire x_19900;
wire x_19901;
wire x_19902;
wire x_19903;
wire x_19904;
wire x_19905;
wire x_19906;
wire x_19907;
wire x_19908;
wire x_19909;
wire x_19910;
wire x_19911;
wire x_19912;
wire x_19913;
wire x_19914;
wire x_19915;
wire x_19916;
wire x_19917;
wire x_19918;
wire x_19919;
wire x_19920;
wire x_19921;
wire x_19922;
wire x_19923;
wire x_19924;
wire x_19925;
wire x_19926;
wire x_19927;
wire x_19928;
wire x_19929;
wire x_19930;
wire x_19931;
wire x_19932;
wire x_19933;
wire x_19934;
wire x_19935;
wire x_19936;
wire x_19937;
wire x_19938;
wire x_19939;
wire x_19940;
wire x_19941;
wire x_19942;
wire x_19943;
wire x_19944;
wire x_19945;
wire x_19946;
wire x_19947;
wire x_19948;
wire x_19949;
wire x_19950;
wire x_19951;
wire x_19952;
wire x_19953;
wire x_19954;
wire x_19955;
wire x_19956;
wire x_19957;
wire x_19958;
wire x_19959;
wire x_19960;
wire x_19961;
wire x_19962;
wire x_19963;
wire x_19964;
wire x_19965;
wire x_19966;
wire x_19967;
wire x_19968;
wire x_19969;
wire x_19970;
wire x_19971;
wire x_19972;
wire x_19973;
wire x_19974;
wire x_19975;
wire x_19976;
wire x_19977;
wire x_19978;
wire x_19979;
wire x_19980;
wire x_19981;
wire x_19982;
wire x_19983;
wire x_19984;
wire x_19985;
wire x_19986;
wire x_19987;
wire x_19988;
wire x_19989;
wire x_19990;
wire x_19991;
wire x_19992;
wire x_19993;
wire x_19994;
wire x_19995;
wire x_19996;
wire x_19997;
wire x_19998;
wire x_19999;
wire x_20000;
wire x_20001;
wire x_20002;
wire x_20003;
wire x_20004;
wire x_20005;
wire x_20006;
wire x_20007;
wire x_20008;
wire x_20009;
wire x_20010;
wire x_20011;
wire x_20012;
wire x_20013;
wire x_20014;
wire x_20015;
wire x_20016;
wire x_20017;
wire x_20018;
wire x_20019;
wire x_20020;
wire x_20021;
wire x_20022;
wire x_20023;
wire x_20024;
wire x_20025;
wire x_20026;
wire x_20027;
wire x_20028;
wire x_20029;
wire x_20030;
wire x_20031;
wire x_20032;
wire x_20033;
wire x_20034;
wire x_20035;
wire x_20036;
wire x_20037;
wire x_20038;
wire x_20039;
wire x_20040;
wire x_20041;
wire x_20042;
wire x_20043;
wire x_20044;
wire x_20045;
wire x_20046;
wire x_20047;
wire x_20048;
wire x_20049;
wire x_20050;
wire x_20051;
wire x_20052;
wire x_20053;
wire x_20054;
wire x_20055;
wire x_20056;
wire x_20057;
wire x_20058;
wire x_20059;
wire x_20060;
wire x_20061;
wire x_20062;
wire x_20063;
wire x_20064;
wire x_20065;
wire x_20066;
wire x_20067;
wire x_20068;
wire x_20069;
wire x_20070;
wire x_20071;
wire x_20072;
wire x_20073;
wire x_20074;
wire x_20075;
wire x_20076;
wire x_20077;
wire x_20078;
wire x_20079;
wire x_20080;
wire x_20081;
wire x_20082;
wire x_20083;
wire x_20084;
wire x_20085;
wire x_20086;
wire x_20087;
wire x_20088;
wire x_20089;
wire x_20090;
wire x_20091;
wire x_20092;
wire x_20093;
wire x_20094;
wire x_20095;
wire x_20096;
wire x_20097;
wire x_20098;
wire x_20099;
wire x_20100;
wire x_20101;
wire x_20102;
wire x_20103;
wire x_20104;
wire x_20105;
wire x_20106;
wire x_20107;
wire x_20108;
wire x_20109;
wire x_20110;
wire x_20111;
wire x_20112;
wire x_20113;
wire x_20114;
wire x_20115;
wire x_20116;
wire x_20117;
wire x_20118;
wire x_20119;
wire x_20120;
wire x_20121;
wire x_20122;
wire x_20123;
wire x_20124;
wire x_20125;
wire x_20126;
wire x_20127;
wire x_20128;
wire x_20129;
wire x_20130;
wire x_20131;
wire x_20132;
wire x_20133;
wire x_20134;
wire x_20135;
wire x_20136;
wire x_20137;
wire x_20138;
wire x_20139;
wire x_20140;
wire x_20141;
wire x_20142;
wire x_20143;
wire x_20144;
wire x_20145;
wire x_20146;
wire x_20147;
wire x_20148;
wire x_20149;
wire x_20150;
wire x_20151;
wire x_20152;
wire x_20153;
wire x_20154;
wire x_20155;
wire x_20156;
wire x_20157;
wire x_20158;
wire x_20159;
wire x_20160;
wire x_20161;
wire x_20162;
wire x_20163;
wire x_20164;
wire x_20165;
wire x_20166;
wire x_20167;
wire x_20168;
wire x_20169;
wire x_20170;
wire x_20171;
wire x_20172;
wire x_20173;
wire x_20174;
wire x_20175;
wire x_20176;
wire x_20177;
wire x_20178;
wire x_20179;
wire x_20180;
wire x_20181;
wire x_20182;
wire x_20183;
wire x_20184;
wire x_20185;
wire x_20186;
wire x_20187;
wire x_20188;
wire x_20189;
wire x_20190;
wire x_20191;
wire x_20192;
wire x_20193;
wire x_20194;
wire x_20195;
wire x_20196;
wire x_20197;
wire x_20198;
wire x_20199;
wire x_20200;
wire x_20201;
wire x_20202;
wire x_20203;
wire x_20204;
wire x_20205;
wire x_20206;
wire x_20207;
wire x_20208;
wire x_20209;
wire x_20210;
wire x_20211;
wire x_20212;
wire x_20213;
wire x_20214;
wire x_20215;
wire x_20216;
wire x_20217;
wire x_20218;
wire x_20219;
wire x_20220;
wire x_20221;
wire x_20222;
wire x_20223;
wire x_20224;
wire x_20225;
wire x_20226;
wire x_20227;
wire x_20228;
wire x_20229;
wire x_20230;
wire x_20231;
wire x_20232;
wire x_20233;
wire x_20234;
wire x_20235;
wire x_20236;
wire x_20237;
wire x_20238;
wire x_20239;
wire x_20240;
wire x_20241;
wire x_20242;
wire x_20243;
wire x_20244;
wire x_20245;
wire x_20246;
wire x_20247;
wire x_20248;
wire x_20249;
wire x_20250;
wire x_20251;
wire x_20252;
wire x_20253;
wire x_20254;
wire x_20255;
wire x_20256;
wire x_20257;
wire x_20258;
wire x_20259;
wire x_20260;
wire x_20261;
wire x_20262;
wire x_20263;
wire x_20264;
wire x_20265;
wire x_20266;
wire x_20267;
wire x_20268;
wire x_20269;
wire x_20270;
wire x_20271;
wire x_20272;
wire x_20273;
wire x_20274;
wire x_20275;
wire x_20276;
wire x_20277;
wire x_20278;
wire x_20279;
wire x_20280;
wire x_20281;
wire x_20282;
wire x_20283;
wire x_20284;
wire x_20285;
wire x_20286;
wire x_20287;
wire x_20288;
wire x_20289;
wire x_20290;
wire x_20291;
wire x_20292;
wire x_20293;
wire x_20294;
wire x_20295;
wire x_20296;
wire x_20297;
wire x_20298;
wire x_20299;
wire x_20300;
wire x_20301;
wire x_20302;
wire x_20303;
wire x_20304;
wire x_20305;
wire x_20306;
wire x_20307;
wire x_20308;
wire x_20309;
wire x_20310;
wire x_20311;
wire x_20312;
wire x_20313;
wire x_20314;
wire x_20315;
wire x_20316;
wire x_20317;
wire x_20318;
wire x_20319;
wire x_20320;
wire x_20321;
wire x_20322;
wire x_20323;
wire x_20324;
wire x_20325;
wire x_20326;
wire x_20327;
wire x_20328;
wire x_20329;
wire x_20330;
wire x_20331;
wire x_20332;
wire x_20333;
wire x_20334;
wire x_20335;
wire x_20336;
wire x_20337;
wire x_20338;
wire x_20339;
wire x_20340;
wire x_20341;
wire x_20342;
wire x_20343;
wire x_20344;
wire x_20345;
wire x_20346;
wire x_20347;
wire x_20348;
wire x_20349;
wire x_20350;
wire x_20351;
wire x_20352;
wire x_20353;
wire x_20354;
wire x_20355;
wire x_20356;
wire x_20357;
wire x_20358;
wire x_20359;
wire x_20360;
wire x_20361;
wire x_20362;
wire x_20363;
wire x_20364;
wire x_20365;
wire x_20366;
wire x_20367;
wire x_20368;
wire x_20369;
wire x_20370;
wire x_20371;
wire x_20372;
wire x_20373;
wire x_20374;
wire x_20375;
wire x_20376;
wire x_20377;
wire x_20378;
wire x_20379;
wire x_20380;
wire x_20381;
wire x_20382;
wire x_20383;
wire x_20384;
wire x_20385;
wire x_20386;
wire x_20387;
wire x_20388;
wire x_20389;
wire x_20390;
wire x_20391;
wire x_20392;
wire x_20393;
wire x_20394;
wire x_20395;
wire x_20396;
wire x_20397;
wire x_20398;
wire x_20399;
wire x_20400;
wire x_20401;
wire x_20402;
wire x_20403;
wire x_20404;
wire x_20405;
wire x_20406;
wire x_20407;
wire x_20408;
wire x_20409;
wire x_20410;
wire x_20411;
wire x_20412;
wire x_20413;
wire x_20414;
wire x_20415;
wire x_20416;
wire x_20417;
wire x_20418;
wire x_20419;
wire x_20420;
wire x_20421;
wire x_20422;
wire x_20423;
wire x_20424;
wire x_20425;
wire x_20426;
wire x_20427;
wire x_20428;
wire x_20429;
wire x_20430;
wire x_20431;
wire x_20432;
wire x_20433;
wire x_20434;
wire x_20435;
wire x_20436;
wire x_20437;
wire x_20438;
wire x_20439;
wire x_20440;
wire x_20441;
wire x_20442;
wire x_20443;
wire x_20444;
wire x_20445;
wire x_20446;
wire x_20447;
wire x_20448;
wire x_20449;
wire x_20450;
wire x_20451;
wire x_20452;
wire x_20453;
wire x_20454;
wire x_20455;
wire x_20456;
wire x_20457;
wire x_20458;
wire x_20459;
wire x_20460;
wire x_20461;
wire x_20462;
wire x_20463;
wire x_20464;
wire x_20465;
wire x_20466;
wire x_20467;
wire x_20468;
wire x_20469;
wire x_20470;
wire x_20471;
wire x_20472;
wire x_20473;
wire x_20474;
wire x_20475;
wire x_20476;
wire x_20477;
wire x_20478;
wire x_20479;
wire x_20480;
wire x_20481;
wire x_20482;
wire x_20483;
wire x_20484;
wire x_20485;
wire x_20486;
wire x_20487;
wire x_20488;
wire x_20489;
wire x_20490;
wire x_20491;
wire x_20492;
wire x_20493;
wire x_20494;
wire x_20495;
wire x_20496;
wire x_20497;
wire x_20498;
wire x_20499;
wire x_20500;
wire x_20501;
wire x_20502;
wire x_20503;
wire x_20504;
wire x_20505;
wire x_20506;
wire x_20507;
wire x_20508;
wire x_20509;
wire x_20510;
wire x_20511;
wire x_20512;
wire x_20513;
wire x_20514;
wire x_20515;
wire x_20516;
wire x_20517;
wire x_20518;
wire x_20519;
wire x_20520;
wire x_20521;
wire x_20522;
wire x_20523;
wire x_20524;
wire x_20525;
wire x_20526;
wire x_20527;
wire x_20528;
wire x_20529;
wire x_20530;
wire x_20531;
wire x_20532;
wire x_20533;
wire x_20534;
wire x_20535;
wire x_20536;
wire x_20537;
wire x_20538;
wire x_20539;
wire x_20540;
wire x_20541;
wire x_20542;
wire x_20543;
wire x_20544;
wire x_20545;
wire x_20546;
wire x_20547;
wire x_20548;
wire x_20549;
wire x_20550;
wire x_20551;
wire x_20552;
wire x_20553;
wire x_20554;
wire x_20555;
wire x_20556;
wire x_20557;
wire x_20558;
wire x_20559;
wire x_20560;
wire x_20561;
wire x_20562;
wire x_20563;
wire x_20564;
wire x_20565;
wire x_20566;
wire x_20567;
wire x_20568;
wire x_20569;
wire x_20570;
wire x_20571;
wire x_20572;
wire x_20573;
wire x_20574;
wire x_20575;
wire x_20576;
wire x_20577;
wire x_20578;
wire x_20579;
wire x_20580;
wire x_20581;
wire x_20582;
wire x_20583;
wire x_20584;
wire x_20585;
wire x_20586;
wire x_20587;
wire x_20588;
wire x_20589;
wire x_20590;
wire x_20591;
wire x_20592;
wire x_20593;
wire x_20594;
wire x_20595;
wire x_20596;
wire x_20597;
wire x_20598;
wire x_20599;
wire x_20600;
wire x_20601;
wire x_20602;
wire x_20603;
wire x_20604;
wire x_20605;
wire x_20606;
wire x_20607;
wire x_20608;
wire x_20609;
wire x_20610;
wire x_20611;
wire x_20612;
wire x_20613;
wire x_20614;
wire x_20615;
wire x_20616;
wire x_20617;
wire x_20618;
wire x_20619;
wire x_20620;
wire x_20621;
wire x_20622;
wire x_20623;
wire x_20624;
wire x_20625;
wire x_20626;
wire x_20627;
wire x_20628;
wire x_20629;
wire x_20630;
wire x_20631;
wire x_20632;
wire x_20633;
wire x_20634;
wire x_20635;
wire x_20636;
wire x_20637;
wire x_20638;
wire x_20639;
wire x_20640;
wire x_20641;
wire x_20642;
wire x_20643;
wire x_20644;
wire x_20645;
wire x_20646;
wire x_20647;
wire x_20648;
wire x_20649;
wire x_20650;
wire x_20651;
wire x_20652;
wire x_20653;
wire x_20654;
wire x_20655;
wire x_20656;
wire x_20657;
wire x_20658;
wire x_20659;
wire x_20660;
wire x_20661;
wire x_20662;
wire x_20663;
wire x_20664;
wire x_20665;
wire x_20666;
wire x_20667;
wire x_20668;
wire x_20669;
wire x_20670;
wire x_20671;
wire x_20672;
wire x_20673;
wire x_20674;
wire x_20675;
wire x_20676;
wire x_20677;
wire x_20678;
wire x_20679;
wire x_20680;
wire x_20681;
wire x_20682;
wire x_20683;
wire x_20684;
wire x_20685;
wire x_20686;
wire x_20687;
wire x_20688;
wire x_20689;
wire x_20690;
wire x_20691;
wire x_20692;
wire x_20693;
wire x_20694;
wire x_20695;
wire x_20696;
wire x_20697;
wire x_20698;
wire x_20699;
wire x_20700;
wire x_20701;
wire x_20702;
wire x_20703;
wire x_20704;
wire x_20705;
wire x_20706;
wire x_20707;
wire x_20708;
wire x_20709;
wire x_20710;
wire x_20711;
wire x_20712;
wire x_20713;
wire x_20714;
wire x_20715;
wire x_20716;
wire x_20717;
wire x_20718;
wire x_20719;
wire x_20720;
wire x_20721;
wire x_20722;
wire x_20723;
wire x_20724;
wire x_20725;
wire x_20726;
wire x_20727;
wire x_20728;
wire x_20729;
wire x_20730;
wire x_20731;
wire x_20732;
wire x_20733;
wire x_20734;
wire x_20735;
wire x_20736;
wire x_20737;
wire x_20738;
wire x_20739;
wire x_20740;
wire x_20741;
wire x_20742;
wire x_20743;
wire x_20744;
wire x_20745;
wire x_20746;
wire x_20747;
wire x_20748;
wire x_20749;
wire x_20750;
wire x_20751;
wire x_20752;
wire x_20753;
wire x_20754;
wire x_20755;
wire x_20756;
wire x_20757;
wire x_20758;
wire x_20759;
wire x_20760;
wire x_20761;
wire x_20762;
wire x_20763;
wire x_20764;
wire x_20765;
wire x_20766;
wire x_20767;
wire x_20768;
wire x_20769;
wire x_20770;
wire x_20771;
wire x_20772;
wire x_20773;
wire x_20774;
wire x_20775;
wire x_20776;
wire x_20777;
wire x_20778;
wire x_20779;
wire x_20780;
wire x_20781;
wire x_20782;
wire x_20783;
wire x_20784;
wire x_20785;
wire x_20786;
wire x_20787;
wire x_20788;
wire x_20789;
wire x_20790;
wire x_20791;
wire x_20792;
wire x_20793;
wire x_20794;
wire x_20795;
wire x_20796;
wire x_20797;
wire x_20798;
wire x_20799;
wire x_20800;
wire x_20801;
wire x_20802;
wire x_20803;
wire x_20804;
wire x_20805;
wire x_20806;
wire x_20807;
wire x_20808;
wire x_20809;
wire x_20810;
wire x_20811;
wire x_20812;
wire x_20813;
wire x_20814;
wire x_20815;
wire x_20816;
wire x_20817;
wire x_20818;
wire x_20819;
wire x_20820;
wire x_20821;
wire x_20822;
wire x_20823;
wire x_20824;
wire x_20825;
wire x_20826;
wire x_20827;
wire x_20828;
wire x_20829;
wire x_20830;
wire x_20831;
wire x_20832;
wire x_20833;
wire x_20834;
wire x_20835;
wire x_20836;
wire x_20837;
wire x_20838;
wire x_20839;
wire x_20840;
wire x_20841;
wire x_20842;
wire x_20843;
wire x_20844;
wire x_20845;
wire x_20846;
wire x_20847;
wire x_20848;
wire x_20849;
wire x_20850;
wire x_20851;
wire x_20852;
wire x_20853;
wire x_20854;
wire x_20855;
wire x_20856;
wire x_20857;
wire x_20858;
wire x_20859;
wire x_20860;
wire x_20861;
wire x_20862;
wire x_20863;
wire x_20864;
wire x_20865;
wire x_20866;
wire x_20867;
wire x_20868;
wire x_20869;
wire x_20870;
wire x_20871;
wire x_20872;
wire x_20873;
wire x_20874;
wire x_20875;
wire x_20876;
wire x_20877;
wire x_20878;
wire x_20879;
wire x_20880;
wire x_20881;
wire x_20882;
wire x_20883;
wire x_20884;
wire x_20885;
wire x_20886;
wire x_20887;
wire x_20888;
wire x_20889;
wire x_20890;
wire x_20891;
wire x_20892;
wire x_20893;
wire x_20894;
wire x_20895;
wire x_20896;
wire x_20897;
wire x_20898;
wire x_20899;
wire x_20900;
wire x_20901;
wire x_20902;
wire x_20903;
wire x_20904;
wire x_20905;
wire x_20906;
wire x_20907;
wire x_20908;
wire x_20909;
wire x_20910;
wire x_20911;
wire x_20912;
wire x_20913;
wire x_20914;
wire x_20915;
wire x_20916;
wire x_20917;
wire x_20918;
wire x_20919;
wire x_20920;
wire x_20921;
wire x_20922;
wire x_20923;
wire x_20924;
wire x_20925;
wire x_20926;
wire x_20927;
wire x_20928;
wire x_20929;
wire x_20930;
wire x_20931;
wire x_20932;
wire x_20933;
wire x_20934;
wire x_20935;
wire x_20936;
wire x_20937;
wire x_20938;
wire x_20939;
wire x_20940;
wire x_20941;
wire x_20942;
wire x_20943;
wire x_20944;
wire x_20945;
wire x_20946;
wire x_20947;
wire x_20948;
wire x_20949;
wire x_20950;
wire x_20951;
wire x_20952;
wire x_20953;
wire x_20954;
wire x_20955;
wire x_20956;
wire x_20957;
wire x_20958;
wire x_20959;
wire x_20960;
wire x_20961;
wire x_20962;
wire x_20963;
wire x_20964;
wire x_20965;
wire x_20966;
wire x_20967;
wire x_20968;
wire x_20969;
wire x_20970;
wire x_20971;
wire x_20972;
wire x_20973;
wire x_20974;
wire x_20975;
wire x_20976;
wire x_20977;
wire x_20978;
wire x_20979;
wire x_20980;
wire x_20981;
wire x_20982;
wire x_20983;
wire x_20984;
wire x_20985;
wire x_20986;
wire x_20987;
wire x_20988;
wire x_20989;
wire x_20990;
wire x_20991;
wire x_20992;
wire x_20993;
wire x_20994;
wire x_20995;
wire x_20996;
wire x_20997;
wire x_20998;
wire x_20999;
wire x_21000;
wire x_21001;
wire x_21002;
wire x_21003;
wire x_21004;
wire x_21005;
wire x_21006;
wire x_21007;
wire x_21008;
wire x_21009;
wire x_21010;
wire x_21011;
wire x_21012;
wire x_21013;
wire x_21014;
wire x_21015;
wire x_21016;
wire x_21017;
wire x_21018;
wire x_21019;
wire x_21020;
wire x_21021;
wire x_21022;
wire x_21023;
wire x_21024;
wire x_21025;
wire x_21026;
wire x_21027;
wire x_21028;
wire x_21029;
wire x_21030;
wire x_21031;
wire x_21032;
wire x_21033;
wire x_21034;
wire x_21035;
wire x_21036;
wire x_21037;
wire x_21038;
wire x_21039;
wire x_21040;
wire x_21041;
wire x_21042;
wire x_21043;
wire x_21044;
wire x_21045;
wire x_21046;
wire x_21047;
wire x_21048;
wire x_21049;
wire x_21050;
wire x_21051;
wire x_21052;
wire x_21053;
wire x_21054;
wire x_21055;
wire x_21056;
wire x_21057;
wire x_21058;
wire x_21059;
wire x_21060;
wire x_21061;
wire x_21062;
wire x_21063;
wire x_21064;
wire x_21065;
wire x_21066;
wire x_21067;
wire x_21068;
wire x_21069;
wire x_21070;
wire x_21071;
wire x_21072;
wire x_21073;
wire x_21074;
wire x_21075;
wire x_21076;
wire x_21077;
wire x_21078;
wire x_21079;
wire x_21080;
wire x_21081;
wire x_21082;
wire x_21083;
wire x_21084;
wire x_21085;
wire x_21086;
wire x_21087;
wire x_21088;
wire x_21089;
wire x_21090;
wire x_21091;
wire x_21092;
wire x_21093;
wire x_21094;
wire x_21095;
wire x_21096;
wire x_21097;
wire x_21098;
wire x_21099;
wire x_21100;
wire x_21101;
wire x_21102;
wire x_21103;
wire x_21104;
wire x_21105;
wire x_21106;
wire x_21107;
wire x_21108;
wire x_21109;
wire x_21110;
wire x_21111;
wire x_21112;
wire x_21113;
wire x_21114;
wire x_21115;
wire x_21116;
wire x_21117;
wire x_21118;
wire x_21119;
wire x_21120;
wire x_21121;
wire x_21122;
wire x_21123;
wire x_21124;
wire x_21125;
wire x_21126;
wire x_21127;
wire x_21128;
wire x_21129;
wire x_21130;
wire x_21131;
wire x_21132;
wire x_21133;
wire x_21134;
wire x_21135;
wire x_21136;
wire x_21137;
wire x_21138;
wire x_21139;
wire x_21140;
wire x_21141;
wire x_21142;
wire x_21143;
wire x_21144;
wire x_21145;
wire x_21146;
wire x_21147;
wire x_21148;
wire x_21149;
wire x_21150;
wire x_21151;
wire x_21152;
wire x_21153;
wire x_21154;
wire x_21155;
wire x_21156;
wire x_21157;
wire x_21158;
wire x_21159;
wire x_21160;
wire x_21161;
wire x_21162;
wire x_21163;
wire x_21164;
wire x_21165;
wire x_21166;
wire x_21167;
wire x_21168;
wire x_21169;
wire x_21170;
wire x_21171;
wire x_21172;
wire x_21173;
wire x_21174;
wire x_21175;
wire x_21176;
wire x_21177;
wire x_21178;
wire x_21179;
wire x_21180;
wire x_21181;
wire x_21182;
wire x_21183;
wire x_21184;
wire x_21185;
wire x_21186;
wire x_21187;
wire x_21188;
wire x_21189;
wire x_21190;
wire x_21191;
wire x_21192;
wire x_21193;
wire x_21194;
wire x_21195;
wire x_21196;
wire x_21197;
wire x_21198;
wire x_21199;
wire x_21200;
wire x_21201;
wire x_21202;
wire x_21203;
wire x_21204;
wire x_21205;
wire x_21206;
wire x_21207;
wire x_21208;
wire x_21209;
wire x_21210;
wire x_21211;
wire x_21212;
wire x_21213;
wire x_21214;
wire x_21215;
wire x_21216;
wire x_21217;
wire x_21218;
wire x_21219;
wire x_21220;
wire x_21221;
wire x_21222;
wire x_21223;
wire x_21224;
wire x_21225;
wire x_21226;
wire x_21227;
wire x_21228;
wire x_21229;
wire x_21230;
wire x_21231;
wire x_21232;
wire x_21233;
wire x_21234;
wire x_21235;
wire x_21236;
wire x_21237;
wire x_21238;
wire x_21239;
wire x_21240;
wire x_21241;
wire x_21242;
wire x_21243;
wire x_21244;
wire x_21245;
wire x_21246;
wire x_21247;
wire x_21248;
wire x_21249;
wire x_21250;
wire x_21251;
wire x_21252;
wire x_21253;
wire x_21254;
wire x_21255;
wire x_21256;
wire x_21257;
wire x_21258;
wire x_21259;
wire x_21260;
wire x_21261;
wire x_21262;
wire x_21263;
wire x_21264;
wire x_21265;
wire x_21266;
wire x_21267;
wire x_21268;
wire x_21269;
wire x_21270;
wire x_21271;
wire x_21272;
wire x_21273;
wire x_21274;
wire x_21275;
wire x_21276;
wire x_21277;
wire x_21278;
wire x_21279;
wire x_21280;
wire x_21281;
wire x_21282;
wire x_21283;
wire x_21284;
wire x_21285;
wire x_21286;
wire x_21287;
wire x_21288;
wire x_21289;
wire x_21290;
wire x_21291;
wire x_21292;
wire x_21293;
wire x_21294;
wire x_21295;
wire x_21296;
wire x_21297;
wire x_21298;
wire x_21299;
wire x_21300;
wire x_21301;
wire x_21302;
wire x_21303;
wire x_21304;
wire x_21305;
wire x_21306;
wire x_21307;
wire x_21308;
wire x_21309;
wire x_21310;
wire x_21311;
wire x_21312;
wire x_21313;
wire x_21314;
wire x_21315;
wire x_21316;
wire x_21317;
wire x_21318;
wire x_21319;
wire x_21320;
wire x_21321;
wire x_21322;
wire x_21323;
wire x_21324;
wire x_21325;
wire x_21326;
wire x_21327;
wire x_21328;
wire x_21329;
wire x_21330;
wire x_21331;
wire x_21332;
wire x_21333;
wire x_21334;
wire x_21335;
wire x_21336;
wire x_21337;
wire x_21338;
wire x_21339;
wire x_21340;
wire x_21341;
wire x_21342;
wire x_21343;
wire x_21344;
wire x_21345;
wire x_21346;
wire x_21347;
wire x_21348;
wire x_21349;
wire x_21350;
wire x_21351;
wire x_21352;
wire x_21353;
wire x_21354;
wire x_21355;
wire x_21356;
wire x_21357;
wire x_21358;
wire x_21359;
wire x_21360;
wire x_21361;
wire x_21362;
wire x_21363;
wire x_21364;
wire x_21365;
wire x_21366;
wire x_21367;
wire x_21368;
wire x_21369;
wire x_21370;
wire x_21371;
wire x_21372;
wire x_21373;
wire x_21374;
wire x_21375;
wire x_21376;
wire x_21377;
wire x_21378;
wire x_21379;
wire x_21380;
wire x_21381;
wire x_21382;
wire x_21383;
wire x_21384;
wire x_21385;
wire x_21386;
wire x_21387;
wire x_21388;
wire x_21389;
wire x_21390;
wire x_21391;
wire x_21392;
wire x_21393;
wire x_21394;
wire x_21395;
wire x_21396;
wire x_21397;
wire x_21398;
wire x_21399;
wire x_21400;
wire x_21401;
wire x_21402;
wire x_21403;
wire x_21404;
wire x_21405;
wire x_21406;
wire x_21407;
wire x_21408;
wire x_21409;
wire x_21410;
wire x_21411;
wire x_21412;
wire x_21413;
wire x_21414;
wire x_21415;
wire x_21416;
wire x_21417;
wire x_21418;
wire x_21419;
wire x_21420;
wire x_21421;
wire x_21422;
wire x_21423;
wire x_21424;
wire x_21425;
wire x_21426;
wire x_21427;
wire x_21428;
wire x_21429;
wire x_21430;
wire x_21431;
wire x_21432;
wire x_21433;
wire x_21434;
wire x_21435;
wire x_21436;
wire x_21437;
wire x_21438;
wire x_21439;
wire x_21440;
wire x_21441;
wire x_21442;
wire x_21443;
wire x_21444;
wire x_21445;
wire x_21446;
wire x_21447;
wire x_21448;
wire x_21449;
wire x_21450;
wire x_21451;
wire x_21452;
wire x_21453;
wire x_21454;
wire x_21455;
wire x_21456;
wire x_21457;
wire x_21458;
wire x_21459;
wire x_21460;
wire x_21461;
wire x_21462;
wire x_21463;
wire x_21464;
wire x_21465;
wire x_21466;
wire x_21467;
wire x_21468;
wire x_21469;
wire x_21470;
wire x_21471;
wire x_21472;
wire x_21473;
wire x_21474;
wire x_21475;
wire x_21476;
wire x_21477;
wire x_21478;
wire x_21479;
wire x_21480;
wire x_21481;
wire x_21482;
wire x_21483;
wire x_21484;
wire x_21485;
wire x_21486;
wire x_21487;
wire x_21488;
wire x_21489;
wire x_21490;
wire x_21491;
wire x_21492;
wire x_21493;
wire x_21494;
wire x_21495;
wire x_21496;
wire x_21497;
wire x_21498;
wire x_21499;
wire x_21500;
wire x_21501;
wire x_21502;
wire x_21503;
wire x_21504;
wire x_21505;
wire x_21506;
wire x_21507;
wire x_21508;
wire x_21509;
wire x_21510;
wire x_21511;
wire x_21512;
wire x_21513;
wire x_21514;
wire x_21515;
wire x_21516;
wire x_21517;
wire x_21518;
wire x_21519;
wire x_21520;
wire x_21521;
wire x_21522;
wire x_21523;
wire x_21524;
wire x_21525;
wire x_21526;
wire x_21527;
wire x_21528;
wire x_21529;
wire x_21530;
wire x_21531;
wire x_21532;
wire x_21533;
wire x_21534;
wire x_21535;
wire x_21536;
wire x_21537;
wire x_21538;
wire x_21539;
wire x_21540;
wire x_21541;
wire x_21542;
wire x_21543;
wire x_21544;
wire x_21545;
wire x_21546;
wire x_21547;
wire x_21548;
wire x_21549;
wire x_21550;
wire x_21551;
wire x_21552;
wire x_21553;
wire x_21554;
wire x_21555;
wire x_21556;
wire x_21557;
wire x_21558;
wire x_21559;
wire x_21560;
wire x_21561;
wire x_21562;
wire x_21563;
wire x_21564;
wire x_21565;
wire x_21566;
wire x_21567;
wire x_21568;
wire x_21569;
wire x_21570;
wire x_21571;
wire x_21572;
wire x_21573;
wire x_21574;
wire x_21575;
wire x_21576;
wire x_21577;
wire x_21578;
wire x_21579;
wire x_21580;
wire x_21581;
wire x_21582;
wire x_21583;
wire x_21584;
wire x_21585;
wire x_21586;
wire x_21587;
wire x_21588;
wire x_21589;
wire x_21590;
wire x_21591;
wire x_21592;
wire x_21593;
wire x_21594;
wire x_21595;
wire x_21596;
wire x_21597;
wire x_21598;
wire x_21599;
wire x_21600;
wire x_21601;
wire x_21602;
wire x_21603;
wire x_21604;
wire x_21605;
wire x_21606;
wire x_21607;
wire x_21608;
wire x_21609;
wire x_21610;
wire x_21611;
wire x_21612;
wire x_21613;
wire x_21614;
wire x_21615;
wire x_21616;
wire x_21617;
wire x_21618;
wire x_21619;
wire x_21620;
wire x_21621;
wire x_21622;
wire x_21623;
wire x_21624;
wire x_21625;
wire x_21626;
wire x_21627;
wire x_21628;
wire x_21629;
wire x_21630;
wire x_21631;
wire x_21632;
wire x_21633;
wire x_21634;
wire x_21635;
wire x_21636;
wire x_21637;
wire x_21638;
wire x_21639;
wire x_21640;
wire x_21641;
wire x_21642;
wire x_21643;
wire x_21644;
wire x_21645;
wire x_21646;
wire x_21647;
wire x_21648;
wire x_21649;
wire x_21650;
wire x_21651;
wire x_21652;
wire x_21653;
wire x_21654;
wire x_21655;
wire x_21656;
wire x_21657;
wire x_21658;
wire x_21659;
wire x_21660;
wire x_21661;
wire x_21662;
wire x_21663;
wire x_21664;
wire x_21665;
wire x_21666;
wire x_21667;
wire x_21668;
wire x_21669;
wire x_21670;
wire x_21671;
wire x_21672;
wire x_21673;
wire x_21674;
wire x_21675;
wire x_21676;
wire x_21677;
wire x_21678;
wire x_21679;
wire x_21680;
wire x_21681;
wire x_21682;
wire x_21683;
wire x_21684;
wire x_21685;
wire x_21686;
wire x_21687;
wire x_21688;
wire x_21689;
wire x_21690;
wire x_21691;
wire x_21692;
wire x_21693;
wire x_21694;
wire x_21695;
wire x_21696;
wire x_21697;
wire x_21698;
wire x_21699;
wire x_21700;
wire x_21701;
wire x_21702;
wire x_21703;
wire x_21704;
wire x_21705;
wire x_21706;
wire x_21707;
wire x_21708;
wire x_21709;
wire x_21710;
wire x_21711;
wire x_21712;
wire x_21713;
wire x_21714;
wire x_21715;
wire x_21716;
wire x_21717;
wire x_21718;
wire x_21719;
wire x_21720;
wire x_21721;
wire x_21722;
wire x_21723;
wire x_21724;
wire x_21725;
wire x_21726;
wire x_21727;
wire x_21728;
wire x_21729;
wire x_21730;
wire x_21731;
wire x_21732;
wire x_21733;
wire x_21734;
wire x_21735;
wire x_21736;
wire x_21737;
wire x_21738;
wire x_21739;
wire x_21740;
wire x_21741;
wire x_21742;
wire x_21743;
wire x_21744;
wire x_21745;
wire x_21746;
wire x_21747;
wire x_21748;
wire x_21749;
wire x_21750;
wire x_21751;
wire x_21752;
wire x_21753;
wire x_21754;
wire x_21755;
wire x_21756;
wire x_21757;
wire x_21758;
wire x_21759;
wire x_21760;
wire x_21761;
wire x_21762;
wire x_21763;
wire x_21764;
wire x_21765;
wire x_21766;
wire x_21767;
wire x_21768;
wire x_21769;
wire x_21770;
wire x_21771;
wire x_21772;
wire x_21773;
wire x_21774;
wire x_21775;
wire x_21776;
wire x_21777;
wire x_21778;
wire x_21779;
wire x_21780;
wire x_21781;
wire x_21782;
wire x_21783;
wire x_21784;
wire x_21785;
wire x_21786;
wire x_21787;
wire x_21788;
wire x_21789;
wire x_21790;
wire x_21791;
wire x_21792;
wire x_21793;
wire x_21794;
wire x_21795;
wire x_21796;
wire x_21797;
wire x_21798;
wire x_21799;
wire x_21800;
wire x_21801;
wire x_21802;
wire x_21803;
wire x_21804;
wire x_21805;
wire x_21806;
wire x_21807;
wire x_21808;
wire x_21809;
wire x_21810;
wire x_21811;
wire x_21812;
wire x_21813;
wire x_21814;
wire x_21815;
wire x_21816;
wire x_21817;
wire x_21818;
wire x_21819;
wire x_21820;
wire x_21821;
wire x_21822;
wire x_21823;
wire x_21824;
wire x_21825;
wire x_21826;
wire x_21827;
wire x_21828;
wire x_21829;
wire x_21830;
wire x_21831;
wire x_21832;
wire x_21833;
wire x_21834;
wire x_21835;
wire x_21836;
wire x_21837;
wire x_21838;
wire x_21839;
wire x_21840;
wire x_21841;
wire x_21842;
wire x_21843;
wire x_21844;
wire x_21845;
wire x_21846;
wire x_21847;
wire x_21848;
wire x_21849;
wire x_21850;
wire x_21851;
wire x_21852;
wire x_21853;
wire x_21854;
wire x_21855;
wire x_21856;
wire x_21857;
wire x_21858;
wire x_21859;
wire x_21860;
wire x_21861;
wire x_21862;
wire x_21863;
wire x_21864;
wire x_21865;
wire x_21866;
wire x_21867;
wire x_21868;
wire x_21869;
wire x_21870;
wire x_21871;
wire x_21872;
wire x_21873;
wire x_21874;
wire x_21875;
wire x_21876;
wire x_21877;
wire x_21878;
wire x_21879;
wire x_21880;
wire x_21881;
wire x_21882;
wire x_21883;
wire x_21884;
wire x_21885;
wire x_21886;
wire x_21887;
wire x_21888;
wire x_21889;
wire x_21890;
wire x_21891;
wire x_21892;
wire x_21893;
wire x_21894;
wire x_21895;
wire x_21896;
wire x_21897;
wire x_21898;
wire x_21899;
wire x_21900;
wire x_21901;
wire x_21902;
wire x_21903;
wire x_21904;
wire x_21905;
wire x_21906;
wire x_21907;
wire x_21908;
wire x_21909;
wire x_21910;
wire x_21911;
wire x_21912;
wire x_21913;
wire x_21914;
wire x_21915;
wire x_21916;
wire x_21917;
wire x_21918;
wire x_21919;
wire x_21920;
wire x_21921;
wire x_21922;
wire x_21923;
wire x_21924;
wire x_21925;
wire x_21926;
wire x_21927;
wire x_21928;
wire x_21929;
wire x_21930;
wire x_21931;
wire x_21932;
wire x_21933;
wire x_21934;
wire x_21935;
wire x_21936;
wire x_21937;
wire x_21938;
wire x_21939;
wire x_21940;
wire x_21941;
wire x_21942;
wire x_21943;
wire x_21944;
wire x_21945;
wire x_21946;
wire x_21947;
wire x_21948;
wire x_21949;
wire x_21950;
wire x_21951;
wire x_21952;
wire x_21953;
wire x_21954;
wire x_21955;
wire x_21956;
wire x_21957;
wire x_21958;
wire x_21959;
wire x_21960;
wire x_21961;
wire x_21962;
wire x_21963;
wire x_21964;
wire x_21965;
wire x_21966;
wire x_21967;
wire x_21968;
wire x_21969;
wire x_21970;
wire x_21971;
wire x_21972;
wire x_21973;
wire x_21974;
wire x_21975;
wire x_21976;
wire x_21977;
wire x_21978;
wire x_21979;
wire x_21980;
wire x_21981;
wire x_21982;
wire x_21983;
wire x_21984;
wire x_21985;
wire x_21986;
wire x_21987;
wire x_21988;
wire x_21989;
wire x_21990;
wire x_21991;
wire x_21992;
wire x_21993;
wire x_21994;
wire x_21995;
wire x_21996;
wire x_21997;
wire x_21998;
wire x_21999;
wire x_22000;
wire x_22001;
wire x_22002;
wire x_22003;
wire x_22004;
wire x_22005;
wire x_22006;
wire x_22007;
wire x_22008;
wire x_22009;
wire x_22010;
wire x_22011;
wire x_22012;
wire x_22013;
wire x_22014;
wire x_22015;
wire x_22016;
wire x_22017;
wire x_22018;
wire x_22019;
wire x_22020;
wire x_22021;
wire x_22022;
wire x_22023;
wire x_22024;
wire x_22025;
wire x_22026;
wire x_22027;
wire x_22028;
wire x_22029;
wire x_22030;
wire x_22031;
wire x_22032;
wire x_22033;
wire x_22034;
wire x_22035;
wire x_22036;
wire x_22037;
wire x_22038;
wire x_22039;
wire x_22040;
wire x_22041;
wire x_22042;
wire x_22043;
wire x_22044;
wire x_22045;
wire x_22046;
wire x_22047;
wire x_22048;
wire x_22049;
wire x_22050;
wire x_22051;
wire x_22052;
wire x_22053;
wire x_22054;
wire x_22055;
wire x_22056;
wire x_22057;
wire x_22058;
wire x_22059;
wire x_22060;
wire x_22061;
wire x_22062;
wire x_22063;
wire x_22064;
wire x_22065;
wire x_22066;
wire x_22067;
wire x_22068;
wire x_22069;
wire x_22070;
wire x_22071;
wire x_22072;
wire x_22073;
wire x_22074;
wire x_22075;
wire x_22076;
wire x_22077;
wire x_22078;
wire x_22079;
wire x_22080;
wire x_22081;
wire x_22082;
wire x_22083;
wire x_22084;
wire x_22085;
wire x_22086;
wire x_22087;
wire x_22088;
wire x_22089;
wire x_22090;
wire x_22091;
wire x_22092;
wire x_22093;
wire x_22094;
wire x_22095;
wire x_22096;
wire x_22097;
wire x_22098;
wire x_22099;
wire x_22100;
wire x_22101;
wire x_22102;
wire x_22103;
wire x_22104;
wire x_22105;
wire x_22106;
wire x_22107;
wire x_22108;
wire x_22109;
wire x_22110;
wire x_22111;
wire x_22112;
wire x_22113;
wire x_22114;
wire x_22115;
wire x_22116;
wire x_22117;
wire x_22118;
wire x_22119;
wire x_22120;
wire x_22121;
wire x_22122;
wire x_22123;
wire x_22124;
wire x_22125;
wire x_22126;
wire x_22127;
wire x_22128;
wire x_22129;
wire x_22130;
wire x_22131;
wire x_22132;
wire x_22133;
wire x_22134;
wire x_22135;
wire x_22136;
wire x_22137;
wire x_22138;
wire x_22139;
wire x_22140;
wire x_22141;
wire x_22142;
wire x_22143;
wire x_22144;
wire x_22145;
wire x_22146;
wire x_22147;
wire x_22148;
wire x_22149;
wire x_22150;
wire x_22151;
wire x_22152;
wire x_22153;
wire x_22154;
wire x_22155;
wire x_22156;
wire x_22157;
wire x_22158;
wire x_22159;
wire x_22160;
wire x_22161;
wire x_22162;
wire x_22163;
wire x_22164;
wire x_22165;
wire x_22166;
wire x_22167;
wire x_22168;
wire x_22169;
wire x_22170;
wire x_22171;
wire x_22172;
wire x_22173;
wire x_22174;
wire x_22175;
wire x_22176;
wire x_22177;
wire x_22178;
wire x_22179;
wire x_22180;
wire x_22181;
wire x_22182;
wire x_22183;
wire x_22184;
wire x_22185;
wire x_22186;
wire x_22187;
wire x_22188;
wire x_22189;
wire x_22190;
wire x_22191;
wire x_22192;
wire x_22193;
wire x_22194;
wire x_22195;
wire x_22196;
wire x_22197;
wire x_22198;
wire x_22199;
wire x_22200;
wire x_22201;
wire x_22202;
wire x_22203;
wire x_22204;
wire x_22205;
wire x_22206;
wire x_22207;
wire x_22208;
wire x_22209;
wire x_22210;
wire x_22211;
wire x_22212;
wire x_22213;
wire x_22214;
wire x_22215;
wire x_22216;
wire x_22217;
wire x_22218;
wire x_22219;
wire x_22220;
wire x_22221;
wire x_22222;
wire x_22223;
wire x_22224;
wire x_22225;
wire x_22226;
wire x_22227;
wire x_22228;
wire x_22229;
wire x_22230;
wire x_22231;
wire x_22232;
wire x_22233;
wire x_22234;
wire x_22235;
wire x_22236;
wire x_22237;
wire x_22238;
wire x_22239;
wire x_22240;
wire x_22241;
wire x_22242;
wire x_22243;
wire x_22244;
wire x_22245;
wire x_22246;
wire x_22247;
wire x_22248;
wire x_22249;
wire x_22250;
wire x_22251;
wire x_22252;
wire x_22253;
wire x_22254;
wire x_22255;
wire x_22256;
wire x_22257;
wire x_22258;
wire x_22259;
wire x_22260;
wire x_22261;
wire x_22262;
wire x_22263;
wire x_22264;
wire x_22265;
wire x_22266;
wire x_22267;
wire x_22268;
wire x_22269;
wire x_22270;
wire x_22271;
wire x_22272;
wire x_22273;
wire x_22274;
wire x_22275;
wire x_22276;
wire x_22277;
wire x_22278;
wire x_22279;
wire x_22280;
wire x_22281;
wire x_22282;
wire x_22283;
wire x_22284;
wire x_22285;
wire x_22286;
wire x_22287;
wire x_22288;
wire x_22289;
wire x_22290;
wire x_22291;
wire x_22292;
wire x_22293;
wire x_22294;
wire x_22295;
wire x_22296;
wire x_22297;
wire x_22298;
wire x_22299;
wire x_22300;
wire x_22301;
wire x_22302;
wire x_22303;
wire x_22304;
wire x_22305;
wire x_22306;
wire x_22307;
wire x_22308;
wire x_22309;
wire x_22310;
wire x_22311;
wire x_22312;
wire x_22313;
wire x_22314;
wire x_22315;
wire x_22316;
wire x_22317;
wire x_22318;
wire x_22319;
wire x_22320;
wire x_22321;
wire x_22322;
wire x_22323;
wire x_22324;
wire x_22325;
wire x_22326;
wire x_22327;
wire x_22328;
wire x_22329;
wire x_22330;
wire x_22331;
wire x_22332;
wire x_22333;
wire x_22334;
wire x_22335;
wire x_22336;
wire x_22337;
wire x_22338;
wire x_22339;
wire x_22340;
wire x_22341;
wire x_22342;
wire x_22343;
wire x_22344;
wire x_22345;
wire x_22346;
wire x_22347;
wire x_22348;
wire x_22349;
wire x_22350;
wire x_22351;
wire x_22352;
wire x_22353;
wire x_22354;
wire x_22355;
wire x_22356;
wire x_22357;
wire x_22358;
wire x_22359;
wire x_22360;
wire x_22361;
wire x_22362;
wire x_22363;
wire x_22364;
wire x_22365;
wire x_22366;
wire x_22367;
wire x_22368;
wire x_22369;
wire x_22370;
wire x_22371;
wire x_22372;
wire x_22373;
wire x_22374;
wire x_22375;
wire x_22376;
wire x_22377;
wire x_22378;
wire x_22379;
wire x_22380;
wire x_22381;
wire x_22382;
wire x_22383;
wire x_22384;
wire x_22385;
wire x_22386;
wire x_22387;
wire x_22388;
wire x_22389;
wire x_22390;
wire x_22391;
wire x_22392;
wire x_22393;
wire x_22394;
wire x_22395;
wire x_22396;
wire x_22397;
wire x_22398;
wire x_22399;
wire x_22400;
wire x_22401;
wire x_22402;
wire x_22403;
wire x_22404;
wire x_22405;
wire x_22406;
wire x_22407;
wire x_22408;
wire x_22409;
wire x_22410;
wire x_22411;
wire x_22412;
wire x_22413;
wire x_22414;
wire x_22415;
wire x_22416;
wire x_22417;
wire x_22418;
wire x_22419;
wire x_22420;
wire x_22421;
wire x_22422;
wire x_22423;
wire x_22424;
wire x_22425;
wire x_22426;
wire x_22427;
wire x_22428;
wire x_22429;
wire x_22430;
wire x_22431;
wire x_22432;
wire x_22433;
wire x_22434;
wire x_22435;
wire x_22436;
wire x_22437;
wire x_22438;
wire x_22439;
wire x_22440;
wire x_22441;
wire x_22442;
wire x_22443;
wire x_22444;
wire x_22445;
wire x_22446;
wire x_22447;
wire x_22448;
wire x_22449;
wire x_22450;
wire x_22451;
wire x_22452;
wire x_22453;
wire x_22454;
wire x_22455;
wire x_22456;
wire x_22457;
wire x_22458;
wire x_22459;
wire x_22460;
wire x_22461;
wire x_22462;
wire x_22463;
wire x_22464;
wire x_22465;
wire x_22466;
wire x_22467;
wire x_22468;
wire x_22469;
wire x_22470;
wire x_22471;
wire x_22472;
wire x_22473;
wire x_22474;
wire x_22475;
wire x_22476;
wire x_22477;
wire x_22478;
wire x_22479;
wire x_22480;
wire x_22481;
wire x_22482;
wire x_22483;
wire x_22484;
wire x_22485;
wire x_22486;
wire x_22487;
wire x_22488;
wire x_22489;
wire x_22490;
wire x_22491;
wire x_22492;
wire x_22493;
wire x_22494;
wire x_22495;
wire x_22496;
wire x_22497;
assign v_3381 = 0;
assign x_1 = ~v_3380 | ~v_2730 | ~v_2066 | ~v_1382;
assign x_2 = v_3380 | ~v_3136;
assign x_3 = v_3380 | ~v_3185;
assign x_4 = v_3380 | ~v_3210;
assign x_5 = v_3380 | ~v_3221;
assign x_6 = v_3380 | ~v_3256;
assign x_7 = v_3380 | ~v_3275;
assign x_8 = v_3380 | ~v_3284;
assign x_9 = v_3380 | ~v_3293;
assign x_10 = v_3380 | ~v_3302;
assign x_11 = v_3380 | ~v_3311;
assign x_12 = v_3380 | ~v_3320;
assign x_13 = v_3380 | ~v_3337;
assign x_14 = v_3380 | ~v_3346;
assign x_15 = v_3380 | ~v_3355;
assign x_16 = v_3380 | ~v_3364;
assign x_17 = v_3380 | ~v_3379;
assign x_18 = v_5 | v_4 | v_6 | v_3 | v_2 | v_1 | ~v_1041 | ~v_1040 | ~v_3378 | v_3379;
assign x_19 = v_3378 | ~v_3371;
assign x_20 = v_3378 | ~v_3377;
assign x_21 = v_26 | ~v_3376 | ~v_1037 | ~v_1819 | ~v_2483 | ~v_3253 | ~v_3272 | ~v_3334 | v_3377;
assign x_22 = v_3376 | ~v_3375;
assign x_23 = v_3376 | ~v_698;
assign x_24 = v_3376 | ~v_699;
assign x_25 = v_3376 | ~v_700;
assign x_26 = v_3376 | ~v_701;
assign x_27 = ~v_3374 | ~v_3373 | ~v_3372 | v_3375;
assign x_28 = v_3374 | ~v_1372;
assign x_29 = v_3374 | ~v_2986;
assign x_30 = v_3374 | ~v_2987;
assign x_31 = v_3374 | ~v_2988;
assign x_32 = v_3374 | ~v_2959;
assign x_33 = v_3374 | ~v_2960;
assign x_34 = v_3374 | ~v_2961;
assign x_35 = v_3374 | ~v_2962;
assign x_36 = v_3374 | ~v_763;
assign x_37 = v_3374 | ~v_764;
assign x_38 = v_3374 | ~v_726;
assign x_39 = v_3374 | ~v_1373;
assign x_40 = v_3374 | ~v_2963;
assign x_41 = v_3374 | ~v_731;
assign x_42 = v_3374 | ~v_2964;
assign x_43 = v_3374 | ~v_2993;
assign x_44 = v_3374 | ~v_1374;
assign x_45 = v_3374 | ~v_1375;
assign x_46 = v_3374 | ~v_76;
assign x_47 = v_3374 | ~v_75;
assign x_48 = v_3374 | ~v_74;
assign x_49 = v_3374 | ~v_73;
assign x_50 = v_3374 | ~v_72;
assign x_51 = v_3374 | ~v_71;
assign x_52 = v_3374 | ~v_70;
assign x_53 = v_3374 | ~v_69;
assign x_54 = v_3374 | ~v_68;
assign x_55 = v_3373 | ~v_1367;
assign x_56 = v_3373 | ~v_1368;
assign x_57 = v_3373 | ~v_2977;
assign x_58 = v_3373 | ~v_2978;
assign x_59 = v_3373 | ~v_2948;
assign x_60 = v_3373 | ~v_2949;
assign x_61 = v_3373 | ~v_2950;
assign x_62 = v_3373 | ~v_750;
assign x_63 = v_3373 | ~v_714;
assign x_64 = v_3373 | ~v_2951;
assign x_65 = v_3373 | ~v_2952;
assign x_66 = v_3373 | ~v_2979;
assign x_67 = v_3373 | ~v_2984;
assign x_68 = v_3373 | ~v_757;
assign x_69 = v_3373 | ~v_1369;
assign x_70 = v_3373 | ~v_721;
assign x_71 = v_3373 | ~v_1370;
assign x_72 = v_3373 | ~v_2954;
assign x_73 = v_3373 | ~v_51;
assign x_74 = v_3373 | ~v_50;
assign x_75 = v_3373 | ~v_49;
assign x_76 = v_3373 | ~v_48;
assign x_77 = v_3373 | ~v_47;
assign x_78 = v_3373 | ~v_46;
assign x_79 = v_3373 | ~v_45;
assign x_80 = v_3373 | ~v_44;
assign x_81 = v_3373 | ~v_43;
assign x_82 = v_3372 | ~v_1362;
assign x_83 = v_3372 | ~v_2968;
assign x_84 = v_3372 | ~v_2969;
assign x_85 = v_3372 | ~v_2970;
assign x_86 = v_3372 | ~v_2938;
assign x_87 = v_3372 | ~v_2939;
assign x_88 = v_3372 | ~v_2940;
assign x_89 = v_3372 | ~v_2941;
assign x_90 = v_3372 | ~v_739;
assign x_91 = v_3372 | ~v_705;
assign x_92 = v_3372 | ~v_706;
assign x_93 = v_3372 | ~v_2971;
assign x_94 = v_3372 | ~v_2942;
assign x_95 = v_3372 | ~v_1363;
assign x_96 = v_3372 | ~v_746;
assign x_97 = v_3372 | ~v_1364;
assign x_98 = v_3372 | ~v_1365;
assign x_99 = v_3372 | ~v_2943;
assign x_100 = v_3372 | ~v_25;
assign x_101 = v_3372 | ~v_24;
assign x_102 = v_3372 | ~v_23;
assign x_103 = v_3372 | ~v_22;
assign x_104 = v_3372 | ~v_21;
assign x_105 = v_3372 | ~v_20;
assign x_106 = v_3372 | ~v_19;
assign x_107 = v_3372 | ~v_18;
assign x_108 = v_3372 | ~v_17;
assign x_109 = ~v_2932 | ~v_3370 | v_3371;
assign x_110 = v_3370 | ~v_3326;
assign x_111 = v_3370 | ~v_3263;
assign x_112 = v_3370 | ~v_3236;
assign x_113 = v_3370 | ~v_3369;
assign x_114 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_3368 | v_3369;
assign x_115 = v_3368 | ~v_3365;
assign x_116 = v_3368 | ~v_3366;
assign x_117 = v_3368 | ~v_3367;
assign x_118 = v_76 | v_69 | v_68 | v_75 | v_74 | v_73 | v_72 | v_71 | v_70 | ~v_1356 | ~v_1355 | ~v_2790 | ~v_2761 | ~v_278 | ~v_2760 | ~v_1354 | ~v_273 | ~v_311 | ~v_310 | ~v_2759 | ~v_2758 | ~v_2757 | ~v_2756 | ~v_2785 | ~v_2784 | ~v_2783 | ~v_1353 | v_3367;
assign x_119 = v_50 | v_51 | v_49 | v_48 | v_46 | v_45 | v_43 | ~v_2751 | v_47 | v_44 | ~v_1351 | ~v_268 | ~v_1350 | ~v_304 | ~v_2781 | ~v_2776 | ~v_2749 | ~v_2748 | ~v_261 | ~v_297 | ~v_2747 | ~v_2746 | ~v_2745 | ~v_2775 | ~v_2774 | ~v_1349 | ~v_1348 | v_3366;
assign x_120 = v_25 | v_24 | v_23 | v_22 | v_21 | v_20 | v_19 | v_18 | v_17 | ~v_2740 | ~v_1346 | ~v_1345 | ~v_293 | ~v_1344 | ~v_2739 | ~v_2768 | ~v_253 | ~v_252 | ~v_286 | ~v_2738 | ~v_2737 | ~v_2736 | ~v_2735 | ~v_2767 | ~v_2766 | ~v_2765 | ~v_1343 | v_3365;
assign x_121 = v_9 | v_5 | v_4 | v_10 | v_3 | v_2 | v_1 | ~v_1041 | ~v_1040 | ~v_3363 | v_3364;
assign x_122 = v_3363 | ~v_3359;
assign x_123 = v_3363 | ~v_3362;
assign x_124 = v_26 | ~v_3110 | ~v_1037 | ~v_1819 | ~v_2483 | ~v_3109 | ~v_3108 | ~v_3107 | ~v_3102 | ~v_3361 | ~v_3360 | v_3362;
assign x_125 = v_3361 | ~v_3198;
assign x_126 = v_3361 | ~v_3130;
assign x_127 = v_3360 | ~v_3179;
assign x_128 = v_3360 | ~v_3216;
assign x_129 = ~v_2932 | ~v_3358 | v_3359;
assign x_130 = v_3358 | ~v_3356;
assign x_131 = v_3358 | ~v_3357;
assign x_132 = v_3358 | ~v_2899;
assign x_133 = v_3358 | ~v_2904;
assign x_134 = v_3358 | ~v_2905;
assign x_135 = v_3358 | ~v_2906;
assign x_136 = v_3358 | ~v_2907;
assign x_137 = ~v_2927 | ~v_3186 | v_3357;
assign x_138 = ~v_3211 | ~v_3155 | v_3356;
assign x_139 = v_9 | v_5 | v_6 | v_10 | v_3 | v_2 | v_1 | ~v_1041 | ~v_1040 | ~v_3354 | v_3355;
assign x_140 = v_3354 | ~v_3350;
assign x_141 = v_3354 | ~v_3353;
assign x_142 = v_26 | ~v_1037 | ~v_1819 | ~v_2483 | ~v_3129 | ~v_3128 | ~v_3123 | ~v_3118 | ~v_3117 | ~v_3352 | ~v_3351 | v_3353;
assign x_143 = v_3352 | ~v_3247;
assign x_144 = v_3352 | ~v_3216;
assign x_145 = v_3351 | ~v_3251;
assign x_146 = v_3351 | ~v_3111;
assign x_147 = ~v_2932 | ~v_3349 | v_3350;
assign x_148 = v_3349 | ~v_3347;
assign x_149 = v_3349 | ~v_3348;
assign x_150 = v_3349 | ~v_2914;
assign x_151 = v_3349 | ~v_2915;
assign x_152 = v_3349 | ~v_2920;
assign x_153 = v_3349 | ~v_2925;
assign x_154 = v_3349 | ~v_2926;
assign x_155 = ~v_3211 | ~v_3230 | v_3348;
assign x_156 = ~v_2908 | ~v_3234 | v_3347;
assign x_157 = v_9 | v_7 | v_5 | v_6 | v_8 | v_10 | v_2 | v_1 | ~v_1041 | ~v_1040 | ~v_3345 | v_3346;
assign x_158 = v_3345 | ~v_3341;
assign x_159 = v_3345 | ~v_3344;
assign x_160 = v_26 | ~v_1037 | ~v_1819 | ~v_2483 | ~v_3126 | ~v_3125 | ~v_3124 | ~v_3250 | ~v_3249 | ~v_3343 | ~v_3342 | v_3344;
assign x_161 = v_3343 | ~v_3073;
assign x_162 = v_3343 | ~v_3247;
assign x_163 = v_3342 | ~v_3202;
assign x_164 = v_3342 | ~v_3130;
assign x_165 = ~v_2932 | ~v_3340 | v_3341;
assign x_166 = v_3340 | ~v_3338;
assign x_167 = v_3340 | ~v_3339;
assign x_168 = v_3340 | ~v_3232;
assign x_169 = v_3340 | ~v_3233;
assign x_170 = v_3340 | ~v_2921;
assign x_171 = v_3340 | ~v_2922;
assign x_172 = v_3340 | ~v_2923;
assign x_173 = ~v_3230 | ~v_2870 | v_3339;
assign x_174 = ~v_2927 | ~v_3190 | v_3338;
assign x_175 = v_9 | v_7 | v_5 | v_4 | v_8 | v_10 | v_2 | v_1 | ~v_1041 | ~v_1040 | ~v_3336 | v_3337;
assign x_176 = v_3336 | ~v_3328;
assign x_177 = v_3336 | ~v_3335;
assign x_178 = v_26 | ~v_1037 | ~v_1819 | ~v_2483 | ~v_3334 | ~v_3252 | ~v_3271 | ~v_3333 | v_3335;
assign x_179 = v_3334 | ~v_3111;
assign x_180 = v_3334 | ~v_3202;
assign x_181 = v_3333 | ~v_3332;
assign x_182 = v_3333 | ~v_698;
assign x_183 = v_3333 | ~v_699;
assign x_184 = v_3333 | ~v_700;
assign x_185 = v_3333 | ~v_701;
assign x_186 = ~v_3331 | ~v_3330 | ~v_3329 | v_3332;
assign x_187 = v_3331 | ~v_682;
assign x_188 = v_3331 | ~v_683;
assign x_189 = v_3331 | ~v_906;
assign x_190 = v_3331 | ~v_907;
assign x_191 = v_3331 | ~v_3023;
assign x_192 = v_3331 | ~v_3024;
assign x_193 = v_3331 | ~v_3007;
assign x_194 = v_3331 | ~v_3025;
assign x_195 = v_3331 | ~v_2959;
assign x_196 = v_3331 | ~v_2962;
assign x_197 = v_3331 | ~v_3008;
assign x_198 = v_3331 | ~v_3009;
assign x_199 = v_3331 | ~v_1323;
assign x_200 = v_3331 | ~v_1324;
assign x_201 = v_3331 | ~v_1325;
assign x_202 = v_3331 | ~v_3010;
assign x_203 = v_3331 | ~v_3026;
assign x_204 = v_3331 | ~v_1326;
assign x_205 = v_3331 | ~v_113;
assign x_206 = v_3331 | ~v_112;
assign x_207 = v_3331 | ~v_106;
assign x_208 = v_3331 | ~v_105;
assign x_209 = v_3331 | ~v_76;
assign x_210 = v_3331 | ~v_75;
assign x_211 = v_3331 | ~v_74;
assign x_212 = v_3331 | ~v_73;
assign x_213 = v_3331 | ~v_69;
assign x_214 = v_3330 | ~v_2948;
assign x_215 = v_3330 | ~v_1318;
assign x_216 = v_3330 | ~v_2951;
assign x_217 = v_3330 | ~v_3002;
assign x_218 = v_3330 | ~v_3018;
assign x_219 = v_3330 | ~v_1319;
assign x_220 = v_3330 | ~v_3019;
assign x_221 = v_3330 | ~v_900;
assign x_222 = v_3330 | ~v_3003;
assign x_223 = v_3330 | ~v_3004;
assign x_224 = v_3330 | ~v_3020;
assign x_225 = v_3330 | ~v_677;
assign x_226 = v_3330 | ~v_3021;
assign x_227 = v_3330 | ~v_902;
assign x_228 = v_3330 | ~v_1320;
assign x_229 = v_3330 | ~v_678;
assign x_230 = v_3330 | ~v_1321;
assign x_231 = v_3330 | ~v_3005;
assign x_232 = v_3330 | ~v_111;
assign x_233 = v_3330 | ~v_110;
assign x_234 = v_3330 | ~v_102;
assign x_235 = v_3330 | ~v_101;
assign x_236 = v_3330 | ~v_51;
assign x_237 = v_3330 | ~v_50;
assign x_238 = v_3330 | ~v_49;
assign x_239 = v_3330 | ~v_48;
assign x_240 = v_3330 | ~v_44;
assign x_241 = v_3329 | ~v_646;
assign x_242 = v_3329 | ~v_885;
assign x_243 = v_3329 | ~v_3013;
assign x_244 = v_3329 | ~v_2997;
assign x_245 = v_3329 | ~v_2998;
assign x_246 = v_3329 | ~v_3014;
assign x_247 = v_3329 | ~v_2939;
assign x_248 = v_3329 | ~v_1313;
assign x_249 = v_3329 | ~v_1314;
assign x_250 = v_3329 | ~v_3015;
assign x_251 = v_3329 | ~v_1315;
assign x_252 = v_3329 | ~v_661;
assign x_253 = v_3329 | ~v_890;
assign x_254 = v_3329 | ~v_2999;
assign x_255 = v_3329 | ~v_3000;
assign x_256 = v_3329 | ~v_1316;
assign x_257 = v_3329 | ~v_3016;
assign x_258 = v_3329 | ~v_109;
assign x_259 = v_3329 | ~v_108;
assign x_260 = v_3329 | ~v_95;
assign x_261 = v_3329 | ~v_94;
assign x_262 = v_3329 | ~v_2943;
assign x_263 = v_3329 | ~v_25;
assign x_264 = v_3329 | ~v_24;
assign x_265 = v_3329 | ~v_23;
assign x_266 = v_3329 | ~v_22;
assign x_267 = v_3329 | ~v_18;
assign x_268 = ~v_2932 | ~v_3327 | v_3328;
assign x_269 = v_3327 | ~v_3325;
assign x_270 = v_3327 | ~v_3262;
assign x_271 = v_3327 | ~v_3235;
assign x_272 = v_3327 | ~v_3326;
assign x_273 = ~v_3190 | ~v_2908 | v_3326;
assign x_274 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_3324 | v_3325;
assign x_275 = v_3324 | ~v_3321;
assign x_276 = v_3324 | ~v_3322;
assign x_277 = v_3324 | ~v_3323;
assign x_278 = v_76 | v_69 | v_75 | v_74 | v_73 | v_106 | v_105 | v_113 | v_112 | ~v_1306 | ~v_2823 | ~v_2807 | ~v_1305 | ~v_1304 | ~v_1303 | ~v_2806 | ~v_2805 | ~v_2759 | ~v_2756 | ~v_2822 | ~v_2804 | ~v_2821 | ~v_2820 | ~v_454 | ~v_453 | ~v_230 | ~v_229 | v_3323;
assign x_279 = v_50 | v_51 | v_49 | v_48 | v_44 | v_101 | ~v_2802 | v_102 | v_111 | v_110 | ~v_1301 | ~v_225 | ~v_1300 | ~v_449 | ~v_2818 | ~v_224 | ~v_2817 | ~v_2801 | ~v_2800 | ~v_447 | ~v_2816 | ~v_1299 | ~v_2815 | ~v_2799 | ~v_2748 | ~v_1298 | ~v_2745 | v_3322;
assign x_280 = v_25 | v_24 | v_23 | v_22 | v_18 | ~v_2740 | ~v_2813 | v_95 | v_94 | v_108 | v_109 | ~v_1296 | ~v_2797 | ~v_2796 | ~v_437 | ~v_208 | ~v_1295 | ~v_2812 | ~v_1294 | ~v_1293 | ~v_2736 | ~v_2811 | ~v_2795 | ~v_2794 | ~v_2810 | ~v_432 | ~v_193 | v_3321;
assign x_281 = v_7 | v_5 | v_4 | v_6 | v_8 | v_2 | v_1 | ~v_1041 | ~v_1040 | ~v_3319 | v_3320;
assign x_282 = v_3319 | ~v_3315;
assign x_283 = v_3319 | ~v_3318;
assign x_284 = v_26 | ~v_1037 | ~v_1819 | ~v_2483 | ~v_3170 | ~v_3169 | ~v_3168 | ~v_3201 | ~v_3199 | ~v_3317 | ~v_3316 | v_3318;
assign x_285 = v_3317 | ~v_3251;
assign x_286 = v_3317 | ~v_3174;
assign x_287 = v_3316 | ~v_3073;
assign x_288 = v_3316 | ~v_3206;
assign x_289 = ~v_2932 | ~v_3314 | v_3315;
assign x_290 = v_3314 | ~v_3312;
assign x_291 = v_3314 | ~v_3313;
assign x_292 = v_3314 | ~v_3187;
assign x_293 = v_3314 | ~v_3189;
assign x_294 = v_3314 | ~v_3144;
assign x_295 = v_3314 | ~v_3145;
assign x_296 = v_3314 | ~v_3146;
assign x_297 = ~v_3150 | ~v_3234 | v_3313;
assign x_298 = ~v_3194 | ~v_2870 | v_3312;
assign x_299 = v_9 | v_7 | v_4 | v_6 | v_8 | v_10 | v_2 | v_1 | ~v_1041 | ~v_1040 | ~v_3310 | v_3311;
assign x_300 = v_3310 | ~v_3306;
assign x_301 = v_3310 | ~v_3309;
assign x_302 = v_26 | ~v_1037 | ~v_1819 | ~v_2483 | ~v_3072 | ~v_3071 | ~v_3070 | ~v_3069 | ~v_3052 | ~v_3308 | ~v_3307 | v_3309;
assign x_303 = v_3308 | ~v_3116;
assign x_304 = v_3308 | ~v_3251;
assign x_305 = v_3307 | ~v_3202;
assign x_306 = v_3307 | ~v_3216;
assign x_307 = ~v_2932 | ~v_3305 | v_3306;
assign x_308 = v_3305 | ~v_3303;
assign x_309 = v_3305 | ~v_3304;
assign x_310 = v_3305 | ~v_2849;
assign x_311 = v_3305 | ~v_2866;
assign x_312 = v_3305 | ~v_2867;
assign x_313 = v_3305 | ~v_2868;
assign x_314 = v_3305 | ~v_2869;
assign x_315 = ~v_3234 | ~v_2913 | v_3304;
assign x_316 = ~v_3211 | ~v_3190 | v_3303;
assign x_317 = v_9 | v_7 | v_5 | v_6 | v_8 | v_10 | v_3 | v_1 | ~v_1041 | ~v_1040 | ~v_3301 | v_3302;
assign x_318 = v_3301 | ~v_3297;
assign x_319 = v_3301 | ~v_3300;
assign x_320 = v_26 | ~v_1037 | ~v_1819 | ~v_2483 | ~v_3121 | ~v_3120 | ~v_3119 | ~v_3246 | ~v_3245 | ~v_3299 | ~v_3298 | v_3300;
assign x_321 = v_3299 | ~v_3251;
assign x_322 = v_3299 | ~v_3179;
assign x_323 = v_3298 | ~v_3206;
assign x_324 = v_3298 | ~v_3130;
assign x_325 = ~v_2932 | ~v_3296 | v_3297;
assign x_326 = v_3296 | ~v_3294;
assign x_327 = v_3296 | ~v_3295;
assign x_328 = v_3296 | ~v_3228;
assign x_329 = v_3296 | ~v_3229;
assign x_330 = v_3296 | ~v_2916;
assign x_331 = v_3296 | ~v_2917;
assign x_332 = v_3296 | ~v_2918;
assign x_333 = ~v_3155 | ~v_3234 | v_3295;
assign x_334 = ~v_2927 | ~v_3194 | v_3294;
assign x_335 = v_9 | v_7 | v_5 | v_4 | v_8 | v_10 | v_3 | v_1 | ~v_1041 | ~v_1040 | ~v_3292 | v_3293;
assign x_336 = v_3292 | ~v_3288;
assign x_337 = v_3292 | ~v_3291;
assign x_338 = v_26 | ~v_1037 | ~v_1819 | ~v_2483 | ~v_3100 | ~v_3095 | ~v_3090 | ~v_3178 | ~v_3176 | ~v_3290 | ~v_3289 | v_3291;
assign x_339 = v_3290 | ~v_3247;
assign x_340 = v_3290 | ~v_3198;
assign x_341 = v_3289 | ~v_3111;
assign x_342 = v_3289 | ~v_3206;
assign x_343 = ~v_2932 | ~v_3287 | v_3288;
assign x_344 = v_3287 | ~v_3285;
assign x_345 = v_3287 | ~v_3286;
assign x_346 = v_3287 | ~v_3152;
assign x_347 = v_3287 | ~v_3154;
assign x_348 = v_3287 | ~v_2887;
assign x_349 = v_3287 | ~v_2892;
assign x_350 = v_3287 | ~v_2897;
assign x_351 = ~v_3186 | ~v_3230 | v_3286;
assign x_352 = ~v_3194 | ~v_2908 | v_3285;
assign x_353 = v_7 | v_5 | v_4 | v_6 | v_8 | v_3 | v_1 | ~v_1041 | ~v_1040 | ~v_3283 | v_3284;
assign x_354 = v_3283 | ~v_3279;
assign x_355 = v_3283 | ~v_3282;
assign x_356 = v_26 | ~v_1037 | ~v_1819 | ~v_2483 | ~v_3163 | ~v_3162 | ~v_3161 | ~v_3205 | ~v_3204 | ~v_3281 | ~v_3280 | v_3282;
assign x_357 = v_3281 | ~v_3247;
assign x_358 = v_3281 | ~v_3174;
assign x_359 = v_3280 | ~v_3179;
assign x_360 = v_3280 | ~v_3202;
assign x_361 = ~v_2932 | ~v_3278 | v_3279;
assign x_362 = v_3278 | ~v_3276;
assign x_363 = v_3278 | ~v_3277;
assign x_364 = v_3278 | ~v_3192;
assign x_365 = v_3278 | ~v_3193;
assign x_366 = v_3278 | ~v_3137;
assign x_367 = v_3278 | ~v_3138;
assign x_368 = v_3278 | ~v_3139;
assign x_369 = ~v_3150 | ~v_3230 | v_3277;
assign x_370 = ~v_3190 | ~v_3155 | v_3276;
assign x_371 = v_9 | v_7 | v_4 | v_6 | v_8 | v_10 | v_3 | v_1 | ~v_1041 | ~v_1040 | ~v_3274 | v_3275;
assign x_372 = v_3274 | ~v_3265;
assign x_373 = v_3274 | ~v_3273;
assign x_374 = v_26 | ~v_1037 | ~v_1819 | ~v_2483 | ~v_3272 | ~v_3271 | ~v_3248 | ~v_3270 | v_3273;
assign x_375 = v_3272 | ~v_3216;
assign x_376 = v_3272 | ~v_3206;
assign x_377 = v_3271 | ~v_3073;
assign x_378 = v_3271 | ~v_3179;
assign x_379 = v_3270 | ~v_3269;
assign x_380 = v_3270 | ~v_698;
assign x_381 = v_3270 | ~v_699;
assign x_382 = v_3270 | ~v_700;
assign x_383 = v_3270 | ~v_701;
assign x_384 = ~v_3268 | ~v_3267 | ~v_3266 | v_3269;
assign x_385 = v_3268 | ~v_1218;
assign x_386 = v_3268 | ~v_1219;
assign x_387 = v_3268 | ~v_2956;
assign x_388 = v_3268 | ~v_814;
assign x_389 = v_3268 | ~v_2957;
assign x_390 = v_3268 | ~v_815;
assign x_391 = v_3268 | ~v_2958;
assign x_392 = v_3268 | ~v_2959;
assign x_393 = v_3268 | ~v_2962;
assign x_394 = v_3268 | ~v_632;
assign x_395 = v_3268 | ~v_633;
assign x_396 = v_3268 | ~v_1220;
assign x_397 = v_3268 | ~v_1221;
assign x_398 = v_3268 | ~v_3084;
assign x_399 = v_3268 | ~v_3085;
assign x_400 = v_3268 | ~v_3086;
assign x_401 = v_3268 | ~v_3087;
assign x_402 = v_3268 | ~v_2965;
assign x_403 = v_3268 | ~v_113;
assign x_404 = v_3268 | ~v_112;
assign x_405 = v_3268 | ~v_106;
assign x_406 = v_3268 | ~v_105;
assign x_407 = v_3268 | ~v_76;
assign x_408 = v_3268 | ~v_75;
assign x_409 = v_3268 | ~v_74;
assign x_410 = v_3268 | ~v_73;
assign x_411 = v_3268 | ~v_69;
assign x_412 = v_3267 | ~v_1213;
assign x_413 = v_3267 | ~v_1214;
assign x_414 = v_3267 | ~v_2945;
assign x_415 = v_3267 | ~v_803;
assign x_416 = v_3267 | ~v_2946;
assign x_417 = v_3267 | ~v_804;
assign x_418 = v_3267 | ~v_2947;
assign x_419 = v_3267 | ~v_2948;
assign x_420 = v_3267 | ~v_2951;
assign x_421 = v_3267 | ~v_613;
assign x_422 = v_3267 | ~v_614;
assign x_423 = v_3267 | ~v_1215;
assign x_424 = v_3267 | ~v_1216;
assign x_425 = v_3267 | ~v_3079;
assign x_426 = v_3267 | ~v_3080;
assign x_427 = v_3267 | ~v_3081;
assign x_428 = v_3267 | ~v_3082;
assign x_429 = v_3267 | ~v_2953;
assign x_430 = v_3267 | ~v_111;
assign x_431 = v_3267 | ~v_110;
assign x_432 = v_3267 | ~v_102;
assign x_433 = v_3267 | ~v_101;
assign x_434 = v_3267 | ~v_51;
assign x_435 = v_3267 | ~v_50;
assign x_436 = v_3267 | ~v_49;
assign x_437 = v_3267 | ~v_48;
assign x_438 = v_3267 | ~v_44;
assign x_439 = v_3266 | ~v_1208;
assign x_440 = v_3266 | ~v_1209;
assign x_441 = v_3266 | ~v_2934;
assign x_442 = v_3266 | ~v_792;
assign x_443 = v_3266 | ~v_2935;
assign x_444 = v_3266 | ~v_793;
assign x_445 = v_3266 | ~v_2936;
assign x_446 = v_3266 | ~v_2937;
assign x_447 = v_3266 | ~v_2939;
assign x_448 = v_3266 | ~v_594;
assign x_449 = v_3266 | ~v_595;
assign x_450 = v_3266 | ~v_1210;
assign x_451 = v_3266 | ~v_1211;
assign x_452 = v_3266 | ~v_3074;
assign x_453 = v_3266 | ~v_3075;
assign x_454 = v_3266 | ~v_3076;
assign x_455 = v_3266 | ~v_3077;
assign x_456 = v_3266 | ~v_109;
assign x_457 = v_3266 | ~v_108;
assign x_458 = v_3266 | ~v_95;
assign x_459 = v_3266 | ~v_94;
assign x_460 = v_3266 | ~v_2943;
assign x_461 = v_3266 | ~v_25;
assign x_462 = v_3266 | ~v_24;
assign x_463 = v_3266 | ~v_23;
assign x_464 = v_3266 | ~v_22;
assign x_465 = v_3266 | ~v_18;
assign x_466 = ~v_2932 | ~v_3264 | v_3265;
assign x_467 = v_3264 | ~v_3261;
assign x_468 = v_3264 | ~v_3231;
assign x_469 = v_3264 | ~v_3262;
assign x_470 = v_3264 | ~v_3263;
assign x_471 = ~v_3194 | ~v_3211 | v_3263;
assign x_472 = ~v_3155 | ~v_2870 | v_3262;
assign x_473 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_3260 | v_3261;
assign x_474 = v_3260 | ~v_3257;
assign x_475 = v_3260 | ~v_3258;
assign x_476 = v_3260 | ~v_3259;
assign x_477 = v_76 | v_69 | v_75 | v_74 | v_73 | v_106 | v_105 | v_113 | v_112 | ~v_2762 | ~v_2884 | ~v_2883 | ~v_2882 | ~v_2881 | ~v_1200 | ~v_1199 | ~v_180 | ~v_179 | ~v_2759 | ~v_2756 | ~v_2755 | ~v_362 | ~v_2754 | ~v_361 | ~v_2753 | ~v_1198 | ~v_1197 | v_3259;
assign x_478 = v_50 | v_51 | v_49 | v_48 | v_44 | v_101 | v_102 | v_111 | v_110 | ~v_2750 | ~v_2879 | ~v_2878 | ~v_2877 | ~v_2876 | ~v_1195 | ~v_1194 | ~v_161 | ~v_160 | ~v_2748 | ~v_2745 | ~v_2744 | ~v_351 | ~v_2743 | ~v_350 | ~v_2742 | ~v_1193 | ~v_1192 | v_3258;
assign x_479 = v_25 | v_24 | v_23 | v_22 | v_18 | ~v_2740 | v_95 | v_94 | v_108 | v_109 | ~v_2874 | ~v_2873 | ~v_2872 | ~v_2871 | ~v_1190 | ~v_1189 | ~v_142 | ~v_141 | ~v_2736 | ~v_2734 | ~v_2733 | ~v_340 | ~v_2732 | ~v_339 | ~v_2731 | ~v_1188 | ~v_1187 | v_3257;
assign x_480 = v_9 | v_7 | v_5 | v_6 | v_8 | v_10 | v_3 | v_2 | ~v_1041 | ~v_1040 | ~v_3255 | v_3256;
assign x_481 = v_3255 | ~v_3238;
assign x_482 = v_3255 | ~v_3254;
assign x_483 = v_26 | ~v_1037 | ~v_1819 | ~v_2483 | ~v_3253 | ~v_3252 | ~v_3248 | ~v_3243 | v_3254;
assign x_484 = v_3253 | ~v_3130;
assign x_485 = v_3253 | ~v_3174;
assign x_486 = v_3252 | ~v_3251;
assign x_487 = v_3252 | ~v_3198;
assign x_488 = ~v_3126 | ~v_3125 | ~v_3124 | ~v_3250 | ~v_3249 | v_3251;
assign x_489 = v_3250 | ~v_3122;
assign x_490 = v_3250 | ~v_3028;
assign x_491 = v_3250 | ~v_698;
assign x_492 = v_3250 | ~v_699;
assign x_493 = v_3250 | ~v_700;
assign x_494 = v_3250 | ~v_701;
assign x_495 = v_3249 | ~v_3244;
assign x_496 = v_3249 | ~v_3068;
assign x_497 = v_3249 | ~v_698;
assign x_498 = v_3249 | ~v_699;
assign x_499 = v_3249 | ~v_700;
assign x_500 = v_3249 | ~v_701;
assign x_501 = v_3248 | ~v_3116;
assign x_502 = v_3248 | ~v_3247;
assign x_503 = ~v_3121 | ~v_3120 | ~v_3119 | ~v_3246 | ~v_3245 | v_3247;
assign x_504 = v_3246 | ~v_3127;
assign x_505 = v_3246 | ~v_3099;
assign x_506 = v_3246 | ~v_698;
assign x_507 = v_3246 | ~v_699;
assign x_508 = v_3246 | ~v_700;
assign x_509 = v_3246 | ~v_701;
assign x_510 = v_3245 | ~v_3244;
assign x_511 = v_3245 | ~v_3094;
assign x_512 = v_3245 | ~v_698;
assign x_513 = v_3245 | ~v_699;
assign x_514 = v_3245 | ~v_700;
assign x_515 = v_3245 | ~v_701;
assign x_516 = ~v_3129 | ~v_3118 | ~v_3117 | v_3244;
assign x_517 = v_3243 | ~v_3242;
assign x_518 = v_3243 | ~v_698;
assign x_519 = v_3243 | ~v_699;
assign x_520 = v_3243 | ~v_700;
assign x_521 = v_3243 | ~v_701;
assign x_522 = ~v_3241 | ~v_3240 | ~v_3239 | v_3242;
assign x_523 = v_3241 | ~v_1167;
assign x_524 = v_3241 | ~v_1168;
assign x_525 = v_3241 | ~v_2959;
assign x_526 = v_3241 | ~v_2962;
assign x_527 = v_3241 | ~v_634;
assign x_528 = v_3241 | ~v_635;
assign x_529 = v_3241 | ~v_1169;
assign x_530 = v_3241 | ~v_1170;
assign x_531 = v_3241 | ~v_3046;
assign x_532 = v_3241 | ~v_3047;
assign x_533 = v_3241 | ~v_2989;
assign x_534 = v_3241 | ~v_2990;
assign x_535 = v_3241 | ~v_3048;
assign x_536 = v_3241 | ~v_3049;
assign x_537 = v_3241 | ~v_2991;
assign x_538 = v_3241 | ~v_2992;
assign x_539 = v_3241 | ~v_688;
assign x_540 = v_3241 | ~v_689;
assign x_541 = v_3241 | ~v_132;
assign x_542 = v_3241 | ~v_127;
assign x_543 = v_3241 | ~v_113;
assign x_544 = v_3241 | ~v_112;
assign x_545 = v_3241 | ~v_106;
assign x_546 = v_3241 | ~v_105;
assign x_547 = v_3241 | ~v_76;
assign x_548 = v_3241 | ~v_75;
assign x_549 = v_3241 | ~v_69;
assign x_550 = v_3240 | ~v_2948;
assign x_551 = v_3240 | ~v_2951;
assign x_552 = v_3240 | ~v_615;
assign x_553 = v_3240 | ~v_616;
assign x_554 = v_3240 | ~v_1162;
assign x_555 = v_3240 | ~v_1163;
assign x_556 = v_3240 | ~v_3041;
assign x_557 = v_3240 | ~v_3042;
assign x_558 = v_3240 | ~v_2980;
assign x_559 = v_3240 | ~v_2981;
assign x_560 = v_3240 | ~v_3043;
assign x_561 = v_3240 | ~v_3044;
assign x_562 = v_3240 | ~v_2982;
assign x_563 = v_3240 | ~v_2983;
assign x_564 = v_3240 | ~v_669;
assign x_565 = v_3240 | ~v_670;
assign x_566 = v_3240 | ~v_1164;
assign x_567 = v_3240 | ~v_1165;
assign x_568 = v_3240 | ~v_131;
assign x_569 = v_3240 | ~v_126;
assign x_570 = v_3240 | ~v_111;
assign x_571 = v_3240 | ~v_110;
assign x_572 = v_3240 | ~v_102;
assign x_573 = v_3240 | ~v_101;
assign x_574 = v_3240 | ~v_51;
assign x_575 = v_3240 | ~v_50;
assign x_576 = v_3240 | ~v_44;
assign x_577 = v_3239 | ~v_2939;
assign x_578 = v_3239 | ~v_596;
assign x_579 = v_3239 | ~v_597;
assign x_580 = v_3239 | ~v_1157;
assign x_581 = v_3239 | ~v_1158;
assign x_582 = v_3239 | ~v_3036;
assign x_583 = v_3239 | ~v_3037;
assign x_584 = v_3239 | ~v_2972;
assign x_585 = v_3239 | ~v_2973;
assign x_586 = v_3239 | ~v_3038;
assign x_587 = v_3239 | ~v_3039;
assign x_588 = v_3239 | ~v_2974;
assign x_589 = v_3239 | ~v_2975;
assign x_590 = v_3239 | ~v_653;
assign x_591 = v_3239 | ~v_654;
assign x_592 = v_3239 | ~v_1159;
assign x_593 = v_3239 | ~v_1160;
assign x_594 = v_3239 | ~v_128;
assign x_595 = v_3239 | ~v_122;
assign x_596 = v_3239 | ~v_109;
assign x_597 = v_3239 | ~v_108;
assign x_598 = v_3239 | ~v_95;
assign x_599 = v_3239 | ~v_94;
assign x_600 = v_3239 | ~v_2943;
assign x_601 = v_3239 | ~v_25;
assign x_602 = v_3239 | ~v_24;
assign x_603 = v_3239 | ~v_18;
assign x_604 = ~v_2932 | ~v_3237 | v_3238;
assign x_605 = v_3237 | ~v_3226;
assign x_606 = v_3237 | ~v_3231;
assign x_607 = v_3237 | ~v_3235;
assign x_608 = v_3237 | ~v_3236;
assign x_609 = ~v_3150 | ~v_2927 | v_3236;
assign x_610 = ~v_3186 | ~v_3234 | v_3235;
assign x_611 = v_3234 | ~v_3232;
assign x_612 = v_3234 | ~v_3233;
assign x_613 = v_3234 | ~v_2921;
assign x_614 = v_3234 | ~v_2922;
assign x_615 = v_3234 | ~v_2923;
assign x_616 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2825 | ~v_2919 | v_3233;
assign x_617 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2865 | ~v_3227 | v_3232;
assign x_618 = ~v_3230 | ~v_2913 | v_3231;
assign x_619 = v_3230 | ~v_3228;
assign x_620 = v_3230 | ~v_3229;
assign x_621 = v_3230 | ~v_2916;
assign x_622 = v_3230 | ~v_2917;
assign x_623 = v_3230 | ~v_2918;
assign x_624 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2896 | ~v_2924 | v_3229;
assign x_625 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2891 | ~v_3227 | v_3228;
assign x_626 = v_3227 | ~v_2914;
assign x_627 = v_3227 | ~v_2915;
assign x_628 = v_3227 | ~v_2926;
assign x_629 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_3225 | v_3226;
assign x_630 = v_3225 | ~v_3222;
assign x_631 = v_3225 | ~v_3223;
assign x_632 = v_3225 | ~v_3224;
assign x_633 = v_76 | v_69 | v_75 | v_106 | v_105 | v_132 | v_127 | v_113 | v_112 | ~v_236 | ~v_235 | ~v_2789 | ~v_2788 | ~v_2846 | ~v_2845 | ~v_2787 | ~v_2786 | ~v_2844 | ~v_2843 | ~v_1141 | ~v_1140 | ~v_182 | ~v_181 | ~v_2759 | ~v_2756 | ~v_1139 | ~v_1138 | v_3224;
assign x_634 = v_50 | v_51 | v_44 | v_101 | v_102 | v_111 | v_110 | v_131 | v_126 | ~v_1136 | ~v_1135 | ~v_217 | ~v_216 | ~v_2780 | ~v_2779 | ~v_2841 | ~v_2840 | ~v_2778 | ~v_2777 | ~v_2839 | ~v_2838 | ~v_1134 | ~v_1133 | ~v_163 | ~v_162 | ~v_2748 | ~v_2745 | v_3223;
assign x_635 = v_25 | v_24 | v_18 | ~v_2740 | v_95 | v_94 | v_108 | v_109 | v_128 | v_122 | ~v_1131 | ~v_1130 | ~v_201 | ~v_200 | ~v_2772 | ~v_2771 | ~v_2836 | ~v_2835 | ~v_2770 | ~v_2769 | ~v_2834 | ~v_2833 | ~v_1129 | ~v_1128 | ~v_144 | ~v_143 | ~v_2736 | v_3222;
assign x_636 = v_9 | v_7 | v_4 | v_6 | v_8 | v_10 | v_3 | v_2 | ~v_1041 | ~v_1040 | ~v_3220 | v_3221;
assign x_637 = v_3220 | ~v_3215;
assign x_638 = v_3220 | ~v_3219;
assign x_639 = v_26 | ~v_1037 | ~v_1819 | ~v_2483 | ~v_3034 | ~v_3029 | ~v_2996 | ~v_3115 | ~v_3113 | ~v_3218 | ~v_3217 | v_3219;
assign x_640 = v_3218 | ~v_3073;
assign x_641 = v_3218 | ~v_3198;
assign x_642 = v_3217 | ~v_3216;
assign x_643 = v_3217 | ~v_3174;
assign x_644 = ~v_3063 | ~v_3133 | ~v_3062 | ~v_3057 | ~v_3132 | v_3216;
assign x_645 = ~v_2932 | ~v_3214 | v_3215;
assign x_646 = v_3214 | ~v_3212;
assign x_647 = v_3214 | ~v_3213;
assign x_648 = v_3214 | ~v_2910;
assign x_649 = v_3214 | ~v_2912;
assign x_650 = v_3214 | ~v_2793;
assign x_651 = v_3214 | ~v_2826;
assign x_652 = v_3214 | ~v_2831;
assign x_653 = ~v_3186 | ~v_2870 | v_3213;
assign x_654 = ~v_3150 | ~v_3211 | v_3212;
assign x_655 = v_3211 | ~v_2929;
assign x_656 = v_3211 | ~v_2854;
assign x_657 = v_3211 | ~v_2859;
assign x_658 = v_3211 | ~v_2930;
assign x_659 = v_3211 | ~v_2860;
assign x_660 = v_7 | v_5 | v_4 | v_6 | v_8 | v_3 | v_2 | ~v_1041 | ~v_1040 | ~v_3209 | v_3210;
assign x_661 = v_3209 | ~v_3197;
assign x_662 = v_3209 | ~v_3208;
assign x_663 = v_26 | ~v_1037 | ~v_1819 | ~v_2483 | ~v_3173 | ~v_3172 | ~v_3167 | ~v_3166 | ~v_3165 | ~v_3207 | ~v_3203 | v_3208;
assign x_664 = v_3207 | ~v_3116;
assign x_665 = v_3207 | ~v_3206;
assign x_666 = ~v_3163 | ~v_3162 | ~v_3161 | ~v_3205 | ~v_3204 | v_3206;
assign x_667 = v_3205 | ~v_3099;
assign x_668 = v_3205 | ~v_3171;
assign x_669 = v_3205 | ~v_698;
assign x_670 = v_3205 | ~v_699;
assign x_671 = v_3205 | ~v_700;
assign x_672 = v_3205 | ~v_701;
assign x_673 = v_3204 | ~v_3089;
assign x_674 = v_3204 | ~v_3200;
assign x_675 = v_3204 | ~v_698;
assign x_676 = v_3204 | ~v_699;
assign x_677 = v_3204 | ~v_700;
assign x_678 = v_3204 | ~v_701;
assign x_679 = v_3203 | ~v_3198;
assign x_680 = v_3203 | ~v_3202;
assign x_681 = ~v_3170 | ~v_3169 | ~v_3168 | ~v_3201 | ~v_3199 | v_3202;
assign x_682 = v_3201 | ~v_3200;
assign x_683 = v_3201 | ~v_3051;
assign x_684 = v_3201 | ~v_698;
assign x_685 = v_3201 | ~v_699;
assign x_686 = v_3201 | ~v_700;
assign x_687 = v_3201 | ~v_701;
assign x_688 = ~v_3173 | ~v_3167 | ~v_3166 | v_3200;
assign x_689 = v_3199 | ~v_3164;
assign x_690 = v_3199 | ~v_3028;
assign x_691 = v_3199 | ~v_698;
assign x_692 = v_3199 | ~v_699;
assign x_693 = v_3199 | ~v_700;
assign x_694 = v_3199 | ~v_701;
assign x_695 = ~v_3105 | ~v_3104 | ~v_3103 | ~v_3182 | ~v_3181 | v_3198;
assign x_696 = ~v_2932 | ~v_3196 | v_3197;
assign x_697 = v_3196 | ~v_3191;
assign x_698 = v_3196 | ~v_3195;
assign x_699 = v_3196 | ~v_3141;
assign x_700 = v_3196 | ~v_3142;
assign x_701 = v_3196 | ~v_3143;
assign x_702 = v_3196 | ~v_3148;
assign x_703 = v_3196 | ~v_3149;
assign x_704 = ~v_3194 | ~v_2913 | v_3195;
assign x_705 = v_3194 | ~v_3192;
assign x_706 = v_3194 | ~v_3193;
assign x_707 = v_3194 | ~v_3137;
assign x_708 = v_3194 | ~v_3138;
assign x_709 = v_3194 | ~v_3139;
assign x_710 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_3147 | ~v_2896 | v_3193;
assign x_711 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_3188 | ~v_2886 | v_3192;
assign x_712 = ~v_3190 | ~v_3186 | v_3191;
assign x_713 = v_3190 | ~v_3187;
assign x_714 = v_3190 | ~v_3189;
assign x_715 = v_3190 | ~v_3144;
assign x_716 = v_3190 | ~v_3145;
assign x_717 = v_3190 | ~v_3146;
assign x_718 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2848 | ~v_3188 | v_3189;
assign x_719 = v_3188 | ~v_3142;
assign x_720 = v_3188 | ~v_3143;
assign x_721 = v_3188 | ~v_3149;
assign x_722 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2825 | ~v_3140 | v_3187;
assign x_723 = v_3186 | ~v_3157;
assign x_724 = v_3186 | ~v_3158;
assign x_725 = v_3186 | ~v_2900;
assign x_726 = v_3186 | ~v_2901;
assign x_727 = v_3186 | ~v_2902;
assign x_728 = v_9 | v_7 | v_5 | v_4 | v_8 | v_10 | v_3 | v_2 | ~v_1041 | ~v_1040 | ~v_3184 | v_3185;
assign x_729 = v_3184 | ~v_3160;
assign x_730 = v_3184 | ~v_3183;
assign x_731 = v_26 | ~v_1037 | ~v_1819 | ~v_2483 | ~v_3105 | ~v_3104 | ~v_3103 | ~v_3182 | ~v_3181 | ~v_3180 | ~v_3175 | v_3183;
assign x_732 = v_3182 | ~v_3177;
assign x_733 = v_3182 | ~v_2995;
assign x_734 = v_3182 | ~v_698;
assign x_735 = v_3182 | ~v_699;
assign x_736 = v_3182 | ~v_700;
assign x_737 = v_3182 | ~v_701;
assign x_738 = v_3181 | ~v_3101;
assign x_739 = v_3181 | ~v_3033;
assign x_740 = v_3181 | ~v_698;
assign x_741 = v_3181 | ~v_699;
assign x_742 = v_3181 | ~v_700;
assign x_743 = v_3181 | ~v_701;
assign x_744 = v_3180 | ~v_3116;
assign x_745 = v_3180 | ~v_3179;
assign x_746 = ~v_3100 | ~v_3095 | ~v_3090 | ~v_3178 | ~v_3176 | v_3179;
assign x_747 = v_3178 | ~v_3177;
assign x_748 = v_3178 | ~v_3094;
assign x_749 = v_3178 | ~v_698;
assign x_750 = v_3178 | ~v_699;
assign x_751 = v_3178 | ~v_700;
assign x_752 = v_3178 | ~v_701;
assign x_753 = ~v_3110 | ~v_3109 | ~v_3108 | v_3177;
assign x_754 = v_3176 | ~v_3106;
assign x_755 = v_3176 | ~v_3089;
assign x_756 = v_3176 | ~v_698;
assign x_757 = v_3176 | ~v_699;
assign x_758 = v_3176 | ~v_700;
assign x_759 = v_3176 | ~v_701;
assign x_760 = v_3175 | ~v_3111;
assign x_761 = v_3175 | ~v_3174;
assign x_762 = ~v_3173 | ~v_3172 | ~v_3167 | ~v_3166 | ~v_3165 | v_3174;
assign x_763 = v_3173 | ~v_2995;
assign x_764 = v_3173 | ~v_698;
assign x_765 = v_3173 | ~v_699;
assign x_766 = v_3173 | ~v_700;
assign x_767 = v_3173 | ~v_701;
assign x_768 = v_3172 | ~v_3012;
assign x_769 = v_3172 | ~v_3171;
assign x_770 = v_3172 | ~v_698;
assign x_771 = v_3172 | ~v_699;
assign x_772 = v_3172 | ~v_700;
assign x_773 = v_3172 | ~v_701;
assign x_774 = ~v_3170 | ~v_3169 | ~v_3168 | v_3171;
assign x_775 = v_3170 | ~v_3068;
assign x_776 = v_3170 | ~v_698;
assign x_777 = v_3170 | ~v_699;
assign x_778 = v_3170 | ~v_700;
assign x_779 = v_3170 | ~v_701;
assign x_780 = v_3169 | ~v_3094;
assign x_781 = v_3169 | ~v_3028;
assign x_782 = v_3169 | ~v_698;
assign x_783 = v_3169 | ~v_699;
assign x_784 = v_3169 | ~v_700;
assign x_785 = v_3169 | ~v_701;
assign x_786 = v_3168 | ~v_3051;
assign x_787 = v_3168 | ~v_2995;
assign x_788 = v_3168 | ~v_698;
assign x_789 = v_3168 | ~v_699;
assign x_790 = v_3168 | ~v_700;
assign x_791 = v_3168 | ~v_701;
assign x_792 = v_3167 | ~v_3012;
assign x_793 = v_3167 | ~v_3068;
assign x_794 = v_3167 | ~v_698;
assign x_795 = v_3167 | ~v_699;
assign x_796 = v_3167 | ~v_700;
assign x_797 = v_3167 | ~v_701;
assign x_798 = v_3166 | ~v_3033;
assign x_799 = v_3166 | ~v_3094;
assign x_800 = v_3166 | ~v_698;
assign x_801 = v_3166 | ~v_699;
assign x_802 = v_3166 | ~v_700;
assign x_803 = v_3166 | ~v_701;
assign x_804 = v_3165 | ~v_3164;
assign x_805 = v_3165 | ~v_3033;
assign x_806 = v_3165 | ~v_698;
assign x_807 = v_3165 | ~v_699;
assign x_808 = v_3165 | ~v_700;
assign x_809 = v_3165 | ~v_701;
assign x_810 = ~v_3163 | ~v_3162 | ~v_3161 | v_3164;
assign x_811 = v_3163 | ~v_3094;
assign x_812 = v_3163 | ~v_698;
assign x_813 = v_3163 | ~v_699;
assign x_814 = v_3163 | ~v_700;
assign x_815 = v_3163 | ~v_701;
assign x_816 = v_3162 | ~v_3099;
assign x_817 = v_3162 | ~v_3068;
assign x_818 = v_3162 | ~v_698;
assign x_819 = v_3162 | ~v_699;
assign x_820 = v_3162 | ~v_700;
assign x_821 = v_3162 | ~v_701;
assign x_822 = v_3161 | ~v_3089;
assign x_823 = v_3161 | ~v_2995;
assign x_824 = v_3161 | ~v_698;
assign x_825 = v_3161 | ~v_699;
assign x_826 = v_3161 | ~v_700;
assign x_827 = v_3161 | ~v_701;
assign x_828 = ~v_2932 | ~v_3159 | v_3160;
assign x_829 = v_3159 | ~v_3151;
assign x_830 = v_3159 | ~v_3156;
assign x_831 = v_3159 | ~v_3157;
assign x_832 = v_3159 | ~v_3158;
assign x_833 = v_3159 | ~v_2900;
assign x_834 = v_3159 | ~v_2901;
assign x_835 = v_3159 | ~v_2902;
assign x_836 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2792 | ~v_3153 | v_3158;
assign x_837 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2830 | ~v_2898 | v_3157;
assign x_838 = ~v_3155 | ~v_2913 | v_3156;
assign x_839 = v_3155 | ~v_3152;
assign x_840 = v_3155 | ~v_3154;
assign x_841 = v_3155 | ~v_2887;
assign x_842 = v_3155 | ~v_2892;
assign x_843 = v_3155 | ~v_2897;
assign x_844 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2891 | ~v_3153 | v_3154;
assign x_845 = v_3153 | ~v_2905;
assign x_846 = v_3153 | ~v_2906;
assign x_847 = v_3153 | ~v_2907;
assign x_848 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2886 | ~v_2903 | v_3152;
assign x_849 = ~v_3150 | ~v_2908 | v_3151;
assign x_850 = v_3150 | ~v_3141;
assign x_851 = v_3150 | ~v_3142;
assign x_852 = v_3150 | ~v_3143;
assign x_853 = v_3150 | ~v_3148;
assign x_854 = v_3150 | ~v_3149;
assign x_855 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2792 | v_3149;
assign x_856 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_3147 | ~v_2809 | v_3148;
assign x_857 = v_3147 | ~v_3144;
assign x_858 = v_3147 | ~v_3145;
assign x_859 = v_3147 | ~v_3146;
assign x_860 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2865 | v_3146;
assign x_861 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2825 | ~v_2891 | v_3145;
assign x_862 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2792 | ~v_2848 | v_3144;
assign x_863 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2865 | ~v_2809 | v_3143;
assign x_864 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2891 | ~v_2830 | v_3142;
assign x_865 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2830 | ~v_3140 | v_3141;
assign x_866 = v_3140 | ~v_3137;
assign x_867 = v_3140 | ~v_3138;
assign x_868 = v_3140 | ~v_3139;
assign x_869 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2891 | v_3139;
assign x_870 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2865 | ~v_2896 | v_3138;
assign x_871 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2792 | ~v_2886 | v_3137;
assign x_872 = v_9 | v_4 | v_6 | v_10 | v_3 | v_2 | v_1 | ~v_1041 | ~v_1040 | ~v_3135 | v_3136;
assign x_873 = v_3135 | ~v_2933;
assign x_874 = v_3135 | ~v_3134;
assign x_875 = v_26 | ~v_1037 | ~v_1819 | ~v_2483 | ~v_3063 | ~v_3133 | ~v_3062 | ~v_3057 | ~v_3132 | ~v_3131 | ~v_3112 | v_3134;
assign x_876 = v_3133 | ~v_3114;
assign x_877 = v_3133 | ~v_3061;
assign x_878 = v_3133 | ~v_698;
assign x_879 = v_3133 | ~v_699;
assign x_880 = v_3133 | ~v_700;
assign x_881 = v_3133 | ~v_701;
assign x_882 = v_3132 | ~v_3035;
assign x_883 = v_3132 | ~v_3056;
assign x_884 = v_3132 | ~v_698;
assign x_885 = v_3132 | ~v_699;
assign x_886 = v_3132 | ~v_700;
assign x_887 = v_3132 | ~v_701;
assign x_888 = v_3131 | ~v_3116;
assign x_889 = v_3131 | ~v_3130;
assign x_890 = ~v_3129 | ~v_3128 | ~v_3123 | ~v_3118 | ~v_3117 | v_3130;
assign x_891 = v_3129 | ~v_3056;
assign x_892 = v_3129 | ~v_698;
assign x_893 = v_3129 | ~v_699;
assign x_894 = v_3129 | ~v_700;
assign x_895 = v_3129 | ~v_701;
assign x_896 = v_3128 | ~v_3127;
assign x_897 = v_3128 | ~v_3061;
assign x_898 = v_3128 | ~v_698;
assign x_899 = v_3128 | ~v_699;
assign x_900 = v_3128 | ~v_700;
assign x_901 = v_3128 | ~v_701;
assign x_902 = ~v_3126 | ~v_3125 | ~v_3124 | v_3127;
assign x_903 = v_3126 | ~v_3051;
assign x_904 = v_3126 | ~v_698;
assign x_905 = v_3126 | ~v_699;
assign x_906 = v_3126 | ~v_700;
assign x_907 = v_3126 | ~v_701;
assign x_908 = v_3125 | ~v_3056;
assign x_909 = v_3125 | ~v_3068;
assign x_910 = v_3125 | ~v_698;
assign x_911 = v_3125 | ~v_699;
assign x_912 = v_3125 | ~v_700;
assign x_913 = v_3125 | ~v_701;
assign x_914 = v_3124 | ~v_3089;
assign x_915 = v_3124 | ~v_3028;
assign x_916 = v_3124 | ~v_698;
assign x_917 = v_3124 | ~v_699;
assign x_918 = v_3124 | ~v_700;
assign x_919 = v_3124 | ~v_701;
assign x_920 = v_3123 | ~v_2967;
assign x_921 = v_3123 | ~v_3122;
assign x_922 = v_3123 | ~v_698;
assign x_923 = v_3123 | ~v_699;
assign x_924 = v_3123 | ~v_700;
assign x_925 = v_3123 | ~v_701;
assign x_926 = ~v_3121 | ~v_3120 | ~v_3119 | v_3122;
assign x_927 = v_3121 | ~v_3089;
assign x_928 = v_3121 | ~v_698;
assign x_929 = v_3121 | ~v_699;
assign x_930 = v_3121 | ~v_700;
assign x_931 = v_3121 | ~v_701;
assign x_932 = v_3120 | ~v_3056;
assign x_933 = v_3120 | ~v_3094;
assign x_934 = v_3120 | ~v_698;
assign x_935 = v_3120 | ~v_699;
assign x_936 = v_3120 | ~v_700;
assign x_937 = v_3120 | ~v_701;
assign x_938 = v_3119 | ~v_3099;
assign x_939 = v_3119 | ~v_3051;
assign x_940 = v_3119 | ~v_698;
assign x_941 = v_3119 | ~v_699;
assign x_942 = v_3119 | ~v_700;
assign x_943 = v_3119 | ~v_701;
assign x_944 = v_3118 | ~v_3051;
assign x_945 = v_3118 | ~v_3061;
assign x_946 = v_3118 | ~v_698;
assign x_947 = v_3118 | ~v_699;
assign x_948 = v_3118 | ~v_700;
assign x_949 = v_3118 | ~v_701;
assign x_950 = v_3117 | ~v_2967;
assign x_951 = v_3117 | ~v_3089;
assign x_952 = v_3117 | ~v_698;
assign x_953 = v_3117 | ~v_699;
assign x_954 = v_3117 | ~v_700;
assign x_955 = v_3117 | ~v_701;
assign x_956 = ~v_3034 | ~v_3029 | ~v_2996 | ~v_3115 | ~v_3113 | v_3116;
assign x_957 = v_3115 | ~v_3114;
assign x_958 = v_3115 | ~v_3012;
assign x_959 = v_3115 | ~v_698;
assign x_960 = v_3115 | ~v_699;
assign x_961 = v_3115 | ~v_700;
assign x_962 = v_3115 | ~v_701;
assign x_963 = ~v_3072 | ~v_3071 | ~v_3070 | v_3114;
assign x_964 = v_3113 | ~v_3064;
assign x_965 = v_3113 | ~v_2995;
assign x_966 = v_3113 | ~v_698;
assign x_967 = v_3113 | ~v_699;
assign x_968 = v_3113 | ~v_700;
assign x_969 = v_3113 | ~v_701;
assign x_970 = v_3112 | ~v_3073;
assign x_971 = v_3112 | ~v_3111;
assign x_972 = ~v_3110 | ~v_3109 | ~v_3108 | ~v_3107 | ~v_3102 | v_3111;
assign x_973 = v_3110 | ~v_3061;
assign x_974 = v_3110 | ~v_698;
assign x_975 = v_3110 | ~v_699;
assign x_976 = v_3110 | ~v_700;
assign x_977 = v_3110 | ~v_701;
assign x_978 = v_3109 | ~v_3056;
assign x_979 = v_3109 | ~v_3012;
assign x_980 = v_3109 | ~v_698;
assign x_981 = v_3109 | ~v_699;
assign x_982 = v_3109 | ~v_700;
assign x_983 = v_3109 | ~v_701;
assign x_984 = v_3108 | ~v_2967;
assign x_985 = v_3108 | ~v_3099;
assign x_986 = v_3108 | ~v_698;
assign x_987 = v_3108 | ~v_699;
assign x_988 = v_3108 | ~v_700;
assign x_989 = v_3108 | ~v_701;
assign x_990 = v_3107 | ~v_3106;
assign x_991 = v_3107 | ~v_3056;
assign x_992 = v_3107 | ~v_698;
assign x_993 = v_3107 | ~v_699;
assign x_994 = v_3107 | ~v_700;
assign x_995 = v_3107 | ~v_701;
assign x_996 = ~v_3105 | ~v_3104 | ~v_3103 | v_3106;
assign x_997 = v_3105 | ~v_3012;
assign x_998 = v_3105 | ~v_698;
assign x_999 = v_3105 | ~v_699;
assign x_1000 = v_3105 | ~v_700;
assign x_1001 = v_3105 | ~v_701;
assign x_1002 = v_3104 | ~v_2995;
assign x_1003 = v_3104 | ~v_3061;
assign x_1004 = v_3104 | ~v_698;
assign x_1005 = v_3104 | ~v_699;
assign x_1006 = v_3104 | ~v_700;
assign x_1007 = v_3104 | ~v_701;
assign x_1008 = v_3103 | ~v_3099;
assign x_1009 = v_3103 | ~v_3033;
assign x_1010 = v_3103 | ~v_698;
assign x_1011 = v_3103 | ~v_699;
assign x_1012 = v_3103 | ~v_700;
assign x_1013 = v_3103 | ~v_701;
assign x_1014 = v_3102 | ~v_3101;
assign x_1015 = v_3102 | ~v_2967;
assign x_1016 = v_3102 | ~v_698;
assign x_1017 = v_3102 | ~v_699;
assign x_1018 = v_3102 | ~v_700;
assign x_1019 = v_3102 | ~v_701;
assign x_1020 = ~v_3100 | ~v_3095 | ~v_3090 | v_3101;
assign x_1021 = v_3100 | ~v_3099;
assign x_1022 = v_3100 | ~v_698;
assign x_1023 = v_3100 | ~v_699;
assign x_1024 = v_3100 | ~v_700;
assign x_1025 = v_3100 | ~v_701;
assign x_1026 = ~v_3098 | ~v_3097 | ~v_3096 | v_3099;
assign x_1027 = v_3098 | ~v_782;
assign x_1028 = v_3098 | ~v_783;
assign x_1029 = v_3098 | ~v_682;
assign x_1030 = v_3098 | ~v_683;
assign x_1031 = v_3098 | ~v_3007;
assign x_1032 = v_3098 | ~v_2959;
assign x_1033 = v_3098 | ~v_2962;
assign x_1034 = v_3098 | ~v_3008;
assign x_1035 = v_3098 | ~v_3009;
assign x_1036 = v_3098 | ~v_632;
assign x_1037 = v_3098 | ~v_633;
assign x_1038 = v_3098 | ~v_784;
assign x_1039 = v_3098 | ~v_785;
assign x_1040 = v_3098 | ~v_3084;
assign x_1041 = v_3098 | ~v_3085;
assign x_1042 = v_3098 | ~v_3086;
assign x_1043 = v_3098 | ~v_3087;
assign x_1044 = v_3098 | ~v_3010;
assign x_1045 = v_3098 | ~v_121;
assign x_1046 = v_3098 | ~v_113;
assign x_1047 = v_3098 | ~v_112;
assign x_1048 = v_3098 | ~v_106;
assign x_1049 = v_3098 | ~v_105;
assign x_1050 = v_3098 | ~v_104;
assign x_1051 = v_3098 | ~v_75;
assign x_1052 = v_3098 | ~v_74;
assign x_1053 = v_3098 | ~v_73;
assign x_1054 = v_3097 | ~v_777;
assign x_1055 = v_3097 | ~v_778;
assign x_1056 = v_3097 | ~v_2948;
assign x_1057 = v_3097 | ~v_2951;
assign x_1058 = v_3097 | ~v_613;
assign x_1059 = v_3097 | ~v_614;
assign x_1060 = v_3097 | ~v_779;
assign x_1061 = v_3097 | ~v_780;
assign x_1062 = v_3097 | ~v_3079;
assign x_1063 = v_3097 | ~v_3080;
assign x_1064 = v_3097 | ~v_3081;
assign x_1065 = v_3097 | ~v_3002;
assign x_1066 = v_3097 | ~v_3003;
assign x_1067 = v_3097 | ~v_3004;
assign x_1068 = v_3097 | ~v_677;
assign x_1069 = v_3097 | ~v_678;
assign x_1070 = v_3097 | ~v_3082;
assign x_1071 = v_3097 | ~v_120;
assign x_1072 = v_3097 | ~v_3005;
assign x_1073 = v_3097 | ~v_111;
assign x_1074 = v_3097 | ~v_110;
assign x_1075 = v_3097 | ~v_102;
assign x_1076 = v_3097 | ~v_101;
assign x_1077 = v_3097 | ~v_100;
assign x_1078 = v_3097 | ~v_50;
assign x_1079 = v_3097 | ~v_49;
assign x_1080 = v_3097 | ~v_48;
assign x_1081 = v_3096 | ~v_772;
assign x_1082 = v_3096 | ~v_773;
assign x_1083 = v_3096 | ~v_646;
assign x_1084 = v_3096 | ~v_2997;
assign x_1085 = v_3096 | ~v_2998;
assign x_1086 = v_3096 | ~v_2939;
assign x_1087 = v_3096 | ~v_594;
assign x_1088 = v_3096 | ~v_595;
assign x_1089 = v_3096 | ~v_774;
assign x_1090 = v_3096 | ~v_775;
assign x_1091 = v_3096 | ~v_3074;
assign x_1092 = v_3096 | ~v_3075;
assign x_1093 = v_3096 | ~v_3076;
assign x_1094 = v_3096 | ~v_3077;
assign x_1095 = v_3096 | ~v_661;
assign x_1096 = v_3096 | ~v_2999;
assign x_1097 = v_3096 | ~v_3000;
assign x_1098 = v_3096 | ~v_117;
assign x_1099 = v_3096 | ~v_109;
assign x_1100 = v_3096 | ~v_108;
assign x_1101 = v_3096 | ~v_95;
assign x_1102 = v_3096 | ~v_94;
assign x_1103 = v_3096 | ~v_93;
assign x_1104 = v_3096 | ~v_2943;
assign x_1105 = v_3096 | ~v_24;
assign x_1106 = v_3096 | ~v_23;
assign x_1107 = v_3096 | ~v_22;
assign x_1108 = v_3095 | ~v_3094;
assign x_1109 = v_3095 | ~v_3061;
assign x_1110 = v_3095 | ~v_698;
assign x_1111 = v_3095 | ~v_699;
assign x_1112 = v_3095 | ~v_700;
assign x_1113 = v_3095 | ~v_701;
assign x_1114 = ~v_3093 | ~v_3092 | ~v_3091 | v_3094;
assign x_1115 = v_3093 | ~v_761;
assign x_1116 = v_3093 | ~v_762;
assign x_1117 = v_3093 | ~v_2986;
assign x_1118 = v_3093 | ~v_2987;
assign x_1119 = v_3093 | ~v_2988;
assign x_1120 = v_3093 | ~v_2959;
assign x_1121 = v_3093 | ~v_2962;
assign x_1122 = v_3093 | ~v_763;
assign x_1123 = v_3093 | ~v_764;
assign x_1124 = v_3093 | ~v_765;
assign x_1125 = v_3093 | ~v_766;
assign x_1126 = v_3093 | ~v_632;
assign x_1127 = v_3093 | ~v_633;
assign x_1128 = v_3093 | ~v_3084;
assign x_1129 = v_3093 | ~v_3085;
assign x_1130 = v_3093 | ~v_3086;
assign x_1131 = v_3093 | ~v_3087;
assign x_1132 = v_3093 | ~v_2993;
assign x_1133 = v_3093 | ~v_113;
assign x_1134 = v_3093 | ~v_112;
assign x_1135 = v_3093 | ~v_104;
assign x_1136 = v_3093 | ~v_76;
assign x_1137 = v_3093 | ~v_75;
assign x_1138 = v_3093 | ~v_74;
assign x_1139 = v_3093 | ~v_73;
assign x_1140 = v_3093 | ~v_72;
assign x_1141 = v_3093 | ~v_70;
assign x_1142 = v_3092 | ~v_2977;
assign x_1143 = v_3092 | ~v_2978;
assign x_1144 = v_3092 | ~v_2948;
assign x_1145 = v_3092 | ~v_750;
assign x_1146 = v_3092 | ~v_2951;
assign x_1147 = v_3092 | ~v_2979;
assign x_1148 = v_3092 | ~v_751;
assign x_1149 = v_3092 | ~v_752;
assign x_1150 = v_3092 | ~v_613;
assign x_1151 = v_3092 | ~v_614;
assign x_1152 = v_3092 | ~v_3079;
assign x_1153 = v_3092 | ~v_3080;
assign x_1154 = v_3092 | ~v_3081;
assign x_1155 = v_3092 | ~v_753;
assign x_1156 = v_3092 | ~v_754;
assign x_1157 = v_3092 | ~v_2984;
assign x_1158 = v_3092 | ~v_757;
assign x_1159 = v_3092 | ~v_3082;
assign x_1160 = v_3092 | ~v_111;
assign x_1161 = v_3092 | ~v_110;
assign x_1162 = v_3092 | ~v_100;
assign x_1163 = v_3092 | ~v_51;
assign x_1164 = v_3092 | ~v_50;
assign x_1165 = v_3092 | ~v_49;
assign x_1166 = v_3092 | ~v_48;
assign x_1167 = v_3092 | ~v_47;
assign x_1168 = v_3092 | ~v_45;
assign x_1169 = v_3091 | ~v_2968;
assign x_1170 = v_3091 | ~v_2969;
assign x_1171 = v_3091 | ~v_2970;
assign x_1172 = v_3091 | ~v_2939;
assign x_1173 = v_3091 | ~v_739;
assign x_1174 = v_3091 | ~v_2971;
assign x_1175 = v_3091 | ~v_740;
assign x_1176 = v_3091 | ~v_741;
assign x_1177 = v_3091 | ~v_594;
assign x_1178 = v_3091 | ~v_595;
assign x_1179 = v_3091 | ~v_3074;
assign x_1180 = v_3091 | ~v_3075;
assign x_1181 = v_3091 | ~v_3076;
assign x_1182 = v_3091 | ~v_3077;
assign x_1183 = v_3091 | ~v_742;
assign x_1184 = v_3091 | ~v_743;
assign x_1185 = v_3091 | ~v_746;
assign x_1186 = v_3091 | ~v_109;
assign x_1187 = v_3091 | ~v_108;
assign x_1188 = v_3091 | ~v_93;
assign x_1189 = v_3091 | ~v_2943;
assign x_1190 = v_3091 | ~v_25;
assign x_1191 = v_3091 | ~v_24;
assign x_1192 = v_3091 | ~v_23;
assign x_1193 = v_3091 | ~v_22;
assign x_1194 = v_3091 | ~v_21;
assign x_1195 = v_3091 | ~v_19;
assign x_1196 = v_3090 | ~v_3089;
assign x_1197 = v_3090 | ~v_3012;
assign x_1198 = v_3090 | ~v_698;
assign x_1199 = v_3090 | ~v_699;
assign x_1200 = v_3090 | ~v_700;
assign x_1201 = v_3090 | ~v_701;
assign x_1202 = ~v_3088 | ~v_3083 | ~v_3078 | v_3089;
assign x_1203 = v_3088 | ~v_630;
assign x_1204 = v_3088 | ~v_631;
assign x_1205 = v_3088 | ~v_2959;
assign x_1206 = v_3088 | ~v_2962;
assign x_1207 = v_3088 | ~v_632;
assign x_1208 = v_3088 | ~v_633;
assign x_1209 = v_3088 | ~v_634;
assign x_1210 = v_3088 | ~v_635;
assign x_1211 = v_3088 | ~v_636;
assign x_1212 = v_3088 | ~v_637;
assign x_1213 = v_3088 | ~v_3046;
assign x_1214 = v_3088 | ~v_3047;
assign x_1215 = v_3088 | ~v_3048;
assign x_1216 = v_3088 | ~v_3049;
assign x_1217 = v_3088 | ~v_3084;
assign x_1218 = v_3088 | ~v_3085;
assign x_1219 = v_3088 | ~v_3086;
assign x_1220 = v_3088 | ~v_3087;
assign x_1221 = v_3088 | ~v_127;
assign x_1222 = v_3088 | ~v_113;
assign x_1223 = v_3088 | ~v_112;
assign x_1224 = v_3088 | ~v_107;
assign x_1225 = v_3088 | ~v_106;
assign x_1226 = v_3088 | ~v_105;
assign x_1227 = v_3088 | ~v_104;
assign x_1228 = v_3088 | ~v_76;
assign x_1229 = v_3088 | ~v_73;
assign x_1230 = ~v_86 | ~v_114 | v_3087;
assign x_1231 = ~v_78 | v_114 | v_3086;
assign x_1232 = ~v_88 | ~v_115 | v_3085;
assign x_1233 = ~v_80 | v_115 | v_3084;
assign x_1234 = v_3083 | ~v_611;
assign x_1235 = v_3083 | ~v_612;
assign x_1236 = v_3083 | ~v_2948;
assign x_1237 = v_3083 | ~v_2951;
assign x_1238 = v_3083 | ~v_613;
assign x_1239 = v_3083 | ~v_614;
assign x_1240 = v_3083 | ~v_615;
assign x_1241 = v_3083 | ~v_616;
assign x_1242 = v_3083 | ~v_617;
assign x_1243 = v_3083 | ~v_618;
assign x_1244 = v_3083 | ~v_3041;
assign x_1245 = v_3083 | ~v_3042;
assign x_1246 = v_3083 | ~v_3043;
assign x_1247 = v_3083 | ~v_3044;
assign x_1248 = v_3083 | ~v_3079;
assign x_1249 = v_3083 | ~v_3080;
assign x_1250 = v_3083 | ~v_3081;
assign x_1251 = v_3083 | ~v_3082;
assign x_1252 = v_3083 | ~v_126;
assign x_1253 = v_3083 | ~v_111;
assign x_1254 = v_3083 | ~v_110;
assign x_1255 = v_3083 | ~v_103;
assign x_1256 = v_3083 | ~v_102;
assign x_1257 = v_3083 | ~v_101;
assign x_1258 = v_3083 | ~v_100;
assign x_1259 = v_3083 | ~v_51;
assign x_1260 = v_3083 | ~v_48;
assign x_1261 = ~v_61 | ~v_114 | v_3082;
assign x_1262 = ~v_53 | v_114 | v_3081;
assign x_1263 = ~v_63 | ~v_115 | v_3080;
assign x_1264 = ~v_55 | v_115 | v_3079;
assign x_1265 = v_3078 | ~v_592;
assign x_1266 = v_3078 | ~v_593;
assign x_1267 = v_3078 | ~v_2939;
assign x_1268 = v_3078 | ~v_594;
assign x_1269 = v_3078 | ~v_595;
assign x_1270 = v_3078 | ~v_596;
assign x_1271 = v_3078 | ~v_597;
assign x_1272 = v_3078 | ~v_598;
assign x_1273 = v_3078 | ~v_599;
assign x_1274 = v_3078 | ~v_3036;
assign x_1275 = v_3078 | ~v_3037;
assign x_1276 = v_3078 | ~v_3038;
assign x_1277 = v_3078 | ~v_3039;
assign x_1278 = v_3078 | ~v_3074;
assign x_1279 = v_3078 | ~v_3075;
assign x_1280 = v_3078 | ~v_3076;
assign x_1281 = v_3078 | ~v_3077;
assign x_1282 = v_3078 | ~v_122;
assign x_1283 = v_3078 | ~v_109;
assign x_1284 = v_3078 | ~v_108;
assign x_1285 = v_3078 | ~v_96;
assign x_1286 = v_3078 | ~v_95;
assign x_1287 = v_3078 | ~v_94;
assign x_1288 = v_3078 | ~v_93;
assign x_1289 = v_3078 | ~v_2943;
assign x_1290 = v_3078 | ~v_25;
assign x_1291 = v_3078 | ~v_22;
assign x_1292 = ~v_36 | ~v_114 | v_3077;
assign x_1293 = ~v_28 | v_114 | v_3076;
assign x_1294 = ~v_38 | ~v_115 | v_3075;
assign x_1295 = ~v_30 | v_115 | v_3074;
assign x_1296 = ~v_3072 | ~v_3071 | ~v_3070 | ~v_3069 | ~v_3052 | v_3073;
assign x_1297 = v_3072 | ~v_3028;
assign x_1298 = v_3072 | ~v_698;
assign x_1299 = v_3072 | ~v_699;
assign x_1300 = v_3072 | ~v_700;
assign x_1301 = v_3072 | ~v_701;
assign x_1302 = v_3071 | ~v_2967;
assign x_1303 = v_3071 | ~v_3068;
assign x_1304 = v_3071 | ~v_698;
assign x_1305 = v_3071 | ~v_699;
assign x_1306 = v_3071 | ~v_700;
assign x_1307 = v_3071 | ~v_701;
assign x_1308 = v_3070 | ~v_3033;
assign x_1309 = v_3070 | ~v_3051;
assign x_1310 = v_3070 | ~v_698;
assign x_1311 = v_3070 | ~v_699;
assign x_1312 = v_3070 | ~v_700;
assign x_1313 = v_3070 | ~v_701;
assign x_1314 = v_3069 | ~v_3064;
assign x_1315 = v_3069 | ~v_3068;
assign x_1316 = v_3069 | ~v_698;
assign x_1317 = v_3069 | ~v_699;
assign x_1318 = v_3069 | ~v_700;
assign x_1319 = v_3069 | ~v_701;
assign x_1320 = ~v_3067 | ~v_3066 | ~v_3065 | v_3068;
assign x_1321 = v_3067 | ~v_906;
assign x_1322 = v_3067 | ~v_907;
assign x_1323 = v_3067 | ~v_3023;
assign x_1324 = v_3067 | ~v_3024;
assign x_1325 = v_3067 | ~v_3025;
assign x_1326 = v_3067 | ~v_2986;
assign x_1327 = v_3067 | ~v_2987;
assign x_1328 = v_3067 | ~v_2988;
assign x_1329 = v_3067 | ~v_2959;
assign x_1330 = v_3067 | ~v_2962;
assign x_1331 = v_3067 | ~v_908;
assign x_1332 = v_3067 | ~v_909;
assign x_1333 = v_3067 | ~v_910;
assign x_1334 = v_3067 | ~v_763;
assign x_1335 = v_3067 | ~v_764;
assign x_1336 = v_3067 | ~v_3026;
assign x_1337 = v_3067 | ~v_2993;
assign x_1338 = v_3067 | ~v_914;
assign x_1339 = v_3067 | ~v_121;
assign x_1340 = v_3067 | ~v_113;
assign x_1341 = v_3067 | ~v_112;
assign x_1342 = v_3067 | ~v_104;
assign x_1343 = v_3067 | ~v_75;
assign x_1344 = v_3067 | ~v_74;
assign x_1345 = v_3067 | ~v_73;
assign x_1346 = v_3067 | ~v_72;
assign x_1347 = v_3067 | ~v_70;
assign x_1348 = v_3066 | ~v_2977;
assign x_1349 = v_3066 | ~v_2978;
assign x_1350 = v_3066 | ~v_2948;
assign x_1351 = v_3066 | ~v_896;
assign x_1352 = v_3066 | ~v_750;
assign x_1353 = v_3066 | ~v_2951;
assign x_1354 = v_3066 | ~v_2979;
assign x_1355 = v_3066 | ~v_3018;
assign x_1356 = v_3066 | ~v_897;
assign x_1357 = v_3066 | ~v_3019;
assign x_1358 = v_3066 | ~v_2984;
assign x_1359 = v_3066 | ~v_757;
assign x_1360 = v_3066 | ~v_900;
assign x_1361 = v_3066 | ~v_3020;
assign x_1362 = v_3066 | ~v_3021;
assign x_1363 = v_3066 | ~v_901;
assign x_1364 = v_3066 | ~v_902;
assign x_1365 = v_3066 | ~v_903;
assign x_1366 = v_3066 | ~v_120;
assign x_1367 = v_3066 | ~v_111;
assign x_1368 = v_3066 | ~v_110;
assign x_1369 = v_3066 | ~v_100;
assign x_1370 = v_3066 | ~v_50;
assign x_1371 = v_3066 | ~v_49;
assign x_1372 = v_3066 | ~v_48;
assign x_1373 = v_3066 | ~v_47;
assign x_1374 = v_3066 | ~v_45;
assign x_1375 = v_3065 | ~v_885;
assign x_1376 = v_3065 | ~v_3013;
assign x_1377 = v_3065 | ~v_3014;
assign x_1378 = v_3065 | ~v_2968;
assign x_1379 = v_3065 | ~v_2969;
assign x_1380 = v_3065 | ~v_2970;
assign x_1381 = v_3065 | ~v_2939;
assign x_1382 = v_3065 | ~v_886;
assign x_1383 = v_3065 | ~v_887;
assign x_1384 = v_3065 | ~v_739;
assign x_1385 = v_3065 | ~v_2971;
assign x_1386 = v_3065 | ~v_3015;
assign x_1387 = v_3065 | ~v_746;
assign x_1388 = v_3065 | ~v_890;
assign x_1389 = v_3065 | ~v_891;
assign x_1390 = v_3065 | ~v_892;
assign x_1391 = v_3065 | ~v_117;
assign x_1392 = v_3065 | ~v_3016;
assign x_1393 = v_3065 | ~v_109;
assign x_1394 = v_3065 | ~v_108;
assign x_1395 = v_3065 | ~v_93;
assign x_1396 = v_3065 | ~v_2943;
assign x_1397 = v_3065 | ~v_24;
assign x_1398 = v_3065 | ~v_23;
assign x_1399 = v_3065 | ~v_22;
assign x_1400 = v_3065 | ~v_21;
assign x_1401 = v_3065 | ~v_19;
assign x_1402 = ~v_3063 | ~v_3062 | ~v_3057 | v_3064;
assign x_1403 = v_3063 | ~v_2967;
assign x_1404 = v_3063 | ~v_698;
assign x_1405 = v_3063 | ~v_699;
assign x_1406 = v_3063 | ~v_700;
assign x_1407 = v_3063 | ~v_701;
assign x_1408 = v_3062 | ~v_3028;
assign x_1409 = v_3062 | ~v_3061;
assign x_1410 = v_3062 | ~v_698;
assign x_1411 = v_3062 | ~v_699;
assign x_1412 = v_3062 | ~v_700;
assign x_1413 = v_3062 | ~v_701;
assign x_1414 = ~v_3060 | ~v_3059 | ~v_3058 | v_3061;
assign x_1415 = v_3060 | ~v_682;
assign x_1416 = v_3060 | ~v_683;
assign x_1417 = v_3060 | ~v_3007;
assign x_1418 = v_3060 | ~v_2959;
assign x_1419 = v_3060 | ~v_2960;
assign x_1420 = v_3060 | ~v_2961;
assign x_1421 = v_3060 | ~v_2962;
assign x_1422 = v_3060 | ~v_3008;
assign x_1423 = v_3060 | ~v_3009;
assign x_1424 = v_3060 | ~v_725;
assign x_1425 = v_3060 | ~v_726;
assign x_1426 = v_3060 | ~v_727;
assign x_1427 = v_3060 | ~v_728;
assign x_1428 = v_3060 | ~v_3010;
assign x_1429 = v_3060 | ~v_2963;
assign x_1430 = v_3060 | ~v_731;
assign x_1431 = v_3060 | ~v_2964;
assign x_1432 = v_3060 | ~v_734;
assign x_1433 = v_3060 | ~v_107;
assign x_1434 = v_3060 | ~v_106;
assign x_1435 = v_3060 | ~v_105;
assign x_1436 = v_3060 | ~v_104;
assign x_1437 = v_3060 | ~v_76;
assign x_1438 = v_3060 | ~v_74;
assign x_1439 = v_3060 | ~v_73;
assign x_1440 = v_3060 | ~v_71;
assign x_1441 = v_3060 | ~v_68;
assign x_1442 = v_3059 | ~v_2948;
assign x_1443 = v_3059 | ~v_2949;
assign x_1444 = v_3059 | ~v_2950;
assign x_1445 = v_3059 | ~v_714;
assign x_1446 = v_3059 | ~v_715;
assign x_1447 = v_3059 | ~v_2951;
assign x_1448 = v_3059 | ~v_2952;
assign x_1449 = v_3059 | ~v_3002;
assign x_1450 = v_3059 | ~v_718;
assign x_1451 = v_3059 | ~v_721;
assign x_1452 = v_3059 | ~v_3003;
assign x_1453 = v_3059 | ~v_3004;
assign x_1454 = v_3059 | ~v_677;
assign x_1455 = v_3059 | ~v_722;
assign x_1456 = v_3059 | ~v_678;
assign x_1457 = v_3059 | ~v_723;
assign x_1458 = v_3059 | ~v_3005;
assign x_1459 = v_3059 | ~v_103;
assign x_1460 = v_3059 | ~v_102;
assign x_1461 = v_3059 | ~v_101;
assign x_1462 = v_3059 | ~v_100;
assign x_1463 = v_3059 | ~v_2954;
assign x_1464 = v_3059 | ~v_51;
assign x_1465 = v_3059 | ~v_49;
assign x_1466 = v_3059 | ~v_48;
assign x_1467 = v_3059 | ~v_46;
assign x_1468 = v_3059 | ~v_43;
assign x_1469 = v_3058 | ~v_646;
assign x_1470 = v_3058 | ~v_2997;
assign x_1471 = v_3058 | ~v_2998;
assign x_1472 = v_3058 | ~v_2938;
assign x_1473 = v_3058 | ~v_2939;
assign x_1474 = v_3058 | ~v_2940;
assign x_1475 = v_3058 | ~v_2941;
assign x_1476 = v_3058 | ~v_703;
assign x_1477 = v_3058 | ~v_704;
assign x_1478 = v_3058 | ~v_705;
assign x_1479 = v_3058 | ~v_706;
assign x_1480 = v_3058 | ~v_2942;
assign x_1481 = v_3058 | ~v_661;
assign x_1482 = v_3058 | ~v_711;
assign x_1483 = v_3058 | ~v_2999;
assign x_1484 = v_3058 | ~v_3000;
assign x_1485 = v_3058 | ~v_712;
assign x_1486 = v_3058 | ~v_96;
assign x_1487 = v_3058 | ~v_95;
assign x_1488 = v_3058 | ~v_94;
assign x_1489 = v_3058 | ~v_93;
assign x_1490 = v_3058 | ~v_2943;
assign x_1491 = v_3058 | ~v_25;
assign x_1492 = v_3058 | ~v_23;
assign x_1493 = v_3058 | ~v_22;
assign x_1494 = v_3058 | ~v_20;
assign x_1495 = v_3058 | ~v_17;
assign x_1496 = v_3057 | ~v_3056;
assign x_1497 = v_3057 | ~v_3033;
assign x_1498 = v_3057 | ~v_698;
assign x_1499 = v_3057 | ~v_699;
assign x_1500 = v_3057 | ~v_700;
assign x_1501 = v_3057 | ~v_701;
assign x_1502 = ~v_3055 | ~v_3054 | ~v_3053 | v_3056;
assign x_1503 = v_3055 | ~v_852;
assign x_1504 = v_3055 | ~v_853;
assign x_1505 = v_3055 | ~v_2959;
assign x_1506 = v_3055 | ~v_2960;
assign x_1507 = v_3055 | ~v_2961;
assign x_1508 = v_3055 | ~v_2962;
assign x_1509 = v_3055 | ~v_726;
assign x_1510 = v_3055 | ~v_634;
assign x_1511 = v_3055 | ~v_635;
assign x_1512 = v_3055 | ~v_854;
assign x_1513 = v_3055 | ~v_855;
assign x_1514 = v_3055 | ~v_3046;
assign x_1515 = v_3055 | ~v_3047;
assign x_1516 = v_3055 | ~v_3048;
assign x_1517 = v_3055 | ~v_3049;
assign x_1518 = v_3055 | ~v_2963;
assign x_1519 = v_3055 | ~v_731;
assign x_1520 = v_3055 | ~v_2964;
assign x_1521 = v_3055 | ~v_127;
assign x_1522 = v_3055 | ~v_106;
assign x_1523 = v_3055 | ~v_105;
assign x_1524 = v_3055 | ~v_104;
assign x_1525 = v_3055 | ~v_76;
assign x_1526 = v_3055 | ~v_75;
assign x_1527 = v_3055 | ~v_73;
assign x_1528 = v_3055 | ~v_71;
assign x_1529 = v_3055 | ~v_68;
assign x_1530 = v_3054 | ~v_847;
assign x_1531 = v_3054 | ~v_848;
assign x_1532 = v_3054 | ~v_2948;
assign x_1533 = v_3054 | ~v_2949;
assign x_1534 = v_3054 | ~v_2950;
assign x_1535 = v_3054 | ~v_714;
assign x_1536 = v_3054 | ~v_2951;
assign x_1537 = v_3054 | ~v_2952;
assign x_1538 = v_3054 | ~v_615;
assign x_1539 = v_3054 | ~v_616;
assign x_1540 = v_3054 | ~v_849;
assign x_1541 = v_3054 | ~v_850;
assign x_1542 = v_3054 | ~v_3041;
assign x_1543 = v_3054 | ~v_3042;
assign x_1544 = v_3054 | ~v_3043;
assign x_1545 = v_3054 | ~v_3044;
assign x_1546 = v_3054 | ~v_721;
assign x_1547 = v_3054 | ~v_126;
assign x_1548 = v_3054 | ~v_102;
assign x_1549 = v_3054 | ~v_101;
assign x_1550 = v_3054 | ~v_100;
assign x_1551 = v_3054 | ~v_2954;
assign x_1552 = v_3054 | ~v_51;
assign x_1553 = v_3054 | ~v_50;
assign x_1554 = v_3054 | ~v_48;
assign x_1555 = v_3054 | ~v_46;
assign x_1556 = v_3054 | ~v_43;
assign x_1557 = v_3053 | ~v_842;
assign x_1558 = v_3053 | ~v_843;
assign x_1559 = v_3053 | ~v_2938;
assign x_1560 = v_3053 | ~v_2939;
assign x_1561 = v_3053 | ~v_2940;
assign x_1562 = v_3053 | ~v_2941;
assign x_1563 = v_3053 | ~v_705;
assign x_1564 = v_3053 | ~v_706;
assign x_1565 = v_3053 | ~v_2942;
assign x_1566 = v_3053 | ~v_596;
assign x_1567 = v_3053 | ~v_597;
assign x_1568 = v_3053 | ~v_844;
assign x_1569 = v_3053 | ~v_845;
assign x_1570 = v_3053 | ~v_3036;
assign x_1571 = v_3053 | ~v_3037;
assign x_1572 = v_3053 | ~v_3038;
assign x_1573 = v_3053 | ~v_3039;
assign x_1574 = v_3053 | ~v_122;
assign x_1575 = v_3053 | ~v_95;
assign x_1576 = v_3053 | ~v_94;
assign x_1577 = v_3053 | ~v_93;
assign x_1578 = v_3053 | ~v_2943;
assign x_1579 = v_3053 | ~v_25;
assign x_1580 = v_3053 | ~v_24;
assign x_1581 = v_3053 | ~v_22;
assign x_1582 = v_3053 | ~v_20;
assign x_1583 = v_3053 | ~v_17;
assign x_1584 = v_3052 | ~v_3035;
assign x_1585 = v_3052 | ~v_3051;
assign x_1586 = v_3052 | ~v_698;
assign x_1587 = v_3052 | ~v_699;
assign x_1588 = v_3052 | ~v_700;
assign x_1589 = v_3052 | ~v_701;
assign x_1590 = ~v_3050 | ~v_3045 | ~v_3040 | v_3051;
assign x_1591 = v_3050 | ~v_951;
assign x_1592 = v_3050 | ~v_952;
assign x_1593 = v_3050 | ~v_906;
assign x_1594 = v_3050 | ~v_907;
assign x_1595 = v_3050 | ~v_3023;
assign x_1596 = v_3050 | ~v_3024;
assign x_1597 = v_3050 | ~v_3025;
assign x_1598 = v_3050 | ~v_2959;
assign x_1599 = v_3050 | ~v_2962;
assign x_1600 = v_3050 | ~v_953;
assign x_1601 = v_3050 | ~v_954;
assign x_1602 = v_3050 | ~v_634;
assign x_1603 = v_3050 | ~v_635;
assign x_1604 = v_3050 | ~v_3046;
assign x_1605 = v_3050 | ~v_3047;
assign x_1606 = v_3050 | ~v_3048;
assign x_1607 = v_3050 | ~v_3049;
assign x_1608 = v_3050 | ~v_3026;
assign x_1609 = v_3050 | ~v_127;
assign x_1610 = v_3050 | ~v_113;
assign x_1611 = v_3050 | ~v_112;
assign x_1612 = v_3050 | ~v_106;
assign x_1613 = v_3050 | ~v_105;
assign x_1614 = v_3050 | ~v_104;
assign x_1615 = v_3050 | ~v_76;
assign x_1616 = v_3050 | ~v_75;
assign x_1617 = v_3050 | ~v_73;
assign x_1618 = ~v_87 | ~v_123 | v_3049;
assign x_1619 = ~v_79 | v_123 | v_3048;
assign x_1620 = ~v_90 | ~v_124 | v_3047;
assign x_1621 = ~v_82 | v_124 | v_3046;
assign x_1622 = v_3045 | ~v_946;
assign x_1623 = v_3045 | ~v_947;
assign x_1624 = v_3045 | ~v_2948;
assign x_1625 = v_3045 | ~v_2951;
assign x_1626 = v_3045 | ~v_948;
assign x_1627 = v_3045 | ~v_949;
assign x_1628 = v_3045 | ~v_615;
assign x_1629 = v_3045 | ~v_616;
assign x_1630 = v_3045 | ~v_3041;
assign x_1631 = v_3045 | ~v_3042;
assign x_1632 = v_3045 | ~v_3043;
assign x_1633 = v_3045 | ~v_3044;
assign x_1634 = v_3045 | ~v_3018;
assign x_1635 = v_3045 | ~v_3019;
assign x_1636 = v_3045 | ~v_900;
assign x_1637 = v_3045 | ~v_3020;
assign x_1638 = v_3045 | ~v_3021;
assign x_1639 = v_3045 | ~v_902;
assign x_1640 = v_3045 | ~v_126;
assign x_1641 = v_3045 | ~v_111;
assign x_1642 = v_3045 | ~v_110;
assign x_1643 = v_3045 | ~v_102;
assign x_1644 = v_3045 | ~v_101;
assign x_1645 = v_3045 | ~v_100;
assign x_1646 = v_3045 | ~v_51;
assign x_1647 = v_3045 | ~v_50;
assign x_1648 = v_3045 | ~v_48;
assign x_1649 = ~v_62 | ~v_123 | v_3044;
assign x_1650 = ~v_54 | v_123 | v_3043;
assign x_1651 = ~v_65 | ~v_124 | v_3042;
assign x_1652 = ~v_57 | v_124 | v_3041;
assign x_1653 = v_3040 | ~v_941;
assign x_1654 = v_3040 | ~v_942;
assign x_1655 = v_3040 | ~v_885;
assign x_1656 = v_3040 | ~v_3013;
assign x_1657 = v_3040 | ~v_3014;
assign x_1658 = v_3040 | ~v_2939;
assign x_1659 = v_3040 | ~v_943;
assign x_1660 = v_3040 | ~v_944;
assign x_1661 = v_3040 | ~v_596;
assign x_1662 = v_3040 | ~v_597;
assign x_1663 = v_3040 | ~v_3036;
assign x_1664 = v_3040 | ~v_3037;
assign x_1665 = v_3040 | ~v_3038;
assign x_1666 = v_3040 | ~v_3039;
assign x_1667 = v_3040 | ~v_3015;
assign x_1668 = v_3040 | ~v_890;
assign x_1669 = v_3040 | ~v_122;
assign x_1670 = v_3040 | ~v_3016;
assign x_1671 = v_3040 | ~v_109;
assign x_1672 = v_3040 | ~v_108;
assign x_1673 = v_3040 | ~v_95;
assign x_1674 = v_3040 | ~v_94;
assign x_1675 = v_3040 | ~v_93;
assign x_1676 = v_3040 | ~v_2943;
assign x_1677 = v_3040 | ~v_25;
assign x_1678 = v_3040 | ~v_24;
assign x_1679 = v_3040 | ~v_22;
assign x_1680 = ~v_37 | ~v_123 | v_3039;
assign x_1681 = ~v_29 | v_123 | v_3038;
assign x_1682 = ~v_40 | ~v_124 | v_3037;
assign x_1683 = ~v_32 | v_124 | v_3036;
assign x_1684 = ~v_3034 | ~v_3029 | ~v_2996 | v_3035;
assign x_1685 = v_3034 | ~v_3033;
assign x_1686 = v_3034 | ~v_698;
assign x_1687 = v_3034 | ~v_699;
assign x_1688 = v_3034 | ~v_700;
assign x_1689 = v_3034 | ~v_701;
assign x_1690 = ~v_3032 | ~v_3031 | ~v_3030 | v_3033;
assign x_1691 = v_3032 | ~v_812;
assign x_1692 = v_3032 | ~v_813;
assign x_1693 = v_3032 | ~v_2956;
assign x_1694 = v_3032 | ~v_814;
assign x_1695 = v_3032 | ~v_2957;
assign x_1696 = v_3032 | ~v_815;
assign x_1697 = v_3032 | ~v_2958;
assign x_1698 = v_3032 | ~v_2959;
assign x_1699 = v_3032 | ~v_2962;
assign x_1700 = v_3032 | ~v_816;
assign x_1701 = v_3032 | ~v_817;
assign x_1702 = v_3032 | ~v_2989;
assign x_1703 = v_3032 | ~v_2990;
assign x_1704 = v_3032 | ~v_2991;
assign x_1705 = v_3032 | ~v_2992;
assign x_1706 = v_3032 | ~v_688;
assign x_1707 = v_3032 | ~v_689;
assign x_1708 = v_3032 | ~v_2965;
assign x_1709 = v_3032 | ~v_132;
assign x_1710 = v_3032 | ~v_121;
assign x_1711 = v_3032 | ~v_113;
assign x_1712 = v_3032 | ~v_112;
assign x_1713 = v_3032 | ~v_106;
assign x_1714 = v_3032 | ~v_105;
assign x_1715 = v_3032 | ~v_104;
assign x_1716 = v_3032 | ~v_75;
assign x_1717 = v_3032 | ~v_74;
assign x_1718 = v_3031 | ~v_801;
assign x_1719 = v_3031 | ~v_802;
assign x_1720 = v_3031 | ~v_2945;
assign x_1721 = v_3031 | ~v_803;
assign x_1722 = v_3031 | ~v_2946;
assign x_1723 = v_3031 | ~v_804;
assign x_1724 = v_3031 | ~v_2947;
assign x_1725 = v_3031 | ~v_2948;
assign x_1726 = v_3031 | ~v_2951;
assign x_1727 = v_3031 | ~v_805;
assign x_1728 = v_3031 | ~v_806;
assign x_1729 = v_3031 | ~v_2980;
assign x_1730 = v_3031 | ~v_2981;
assign x_1731 = v_3031 | ~v_2982;
assign x_1732 = v_3031 | ~v_2983;
assign x_1733 = v_3031 | ~v_669;
assign x_1734 = v_3031 | ~v_670;
assign x_1735 = v_3031 | ~v_2953;
assign x_1736 = v_3031 | ~v_131;
assign x_1737 = v_3031 | ~v_120;
assign x_1738 = v_3031 | ~v_111;
assign x_1739 = v_3031 | ~v_110;
assign x_1740 = v_3031 | ~v_102;
assign x_1741 = v_3031 | ~v_101;
assign x_1742 = v_3031 | ~v_100;
assign x_1743 = v_3031 | ~v_50;
assign x_1744 = v_3031 | ~v_49;
assign x_1745 = v_3030 | ~v_790;
assign x_1746 = v_3030 | ~v_791;
assign x_1747 = v_3030 | ~v_2934;
assign x_1748 = v_3030 | ~v_792;
assign x_1749 = v_3030 | ~v_2935;
assign x_1750 = v_3030 | ~v_793;
assign x_1751 = v_3030 | ~v_2936;
assign x_1752 = v_3030 | ~v_2937;
assign x_1753 = v_3030 | ~v_2939;
assign x_1754 = v_3030 | ~v_794;
assign x_1755 = v_3030 | ~v_795;
assign x_1756 = v_3030 | ~v_2972;
assign x_1757 = v_3030 | ~v_2973;
assign x_1758 = v_3030 | ~v_2974;
assign x_1759 = v_3030 | ~v_2975;
assign x_1760 = v_3030 | ~v_653;
assign x_1761 = v_3030 | ~v_654;
assign x_1762 = v_3030 | ~v_128;
assign x_1763 = v_3030 | ~v_117;
assign x_1764 = v_3030 | ~v_109;
assign x_1765 = v_3030 | ~v_108;
assign x_1766 = v_3030 | ~v_95;
assign x_1767 = v_3030 | ~v_94;
assign x_1768 = v_3030 | ~v_93;
assign x_1769 = v_3030 | ~v_2943;
assign x_1770 = v_3030 | ~v_24;
assign x_1771 = v_3030 | ~v_23;
assign x_1772 = v_3029 | ~v_3012;
assign x_1773 = v_3029 | ~v_3028;
assign x_1774 = v_3029 | ~v_698;
assign x_1775 = v_3029 | ~v_699;
assign x_1776 = v_3029 | ~v_700;
assign x_1777 = v_3029 | ~v_701;
assign x_1778 = ~v_3027 | ~v_3022 | ~v_3017 | v_3028;
assign x_1779 = v_3027 | ~v_2956;
assign x_1780 = v_3027 | ~v_814;
assign x_1781 = v_3027 | ~v_2957;
assign x_1782 = v_3027 | ~v_815;
assign x_1783 = v_3027 | ~v_2958;
assign x_1784 = v_3027 | ~v_930;
assign x_1785 = v_3027 | ~v_931;
assign x_1786 = v_3027 | ~v_932;
assign x_1787 = v_3027 | ~v_933;
assign x_1788 = v_3027 | ~v_906;
assign x_1789 = v_3027 | ~v_907;
assign x_1790 = v_3027 | ~v_3023;
assign x_1791 = v_3027 | ~v_3024;
assign x_1792 = v_3027 | ~v_3025;
assign x_1793 = v_3027 | ~v_2959;
assign x_1794 = v_3027 | ~v_2962;
assign x_1795 = v_3027 | ~v_3026;
assign x_1796 = v_3027 | ~v_2965;
assign x_1797 = v_3027 | ~v_113;
assign x_1798 = v_3027 | ~v_112;
assign x_1799 = v_3027 | ~v_107;
assign x_1800 = v_3027 | ~v_106;
assign x_1801 = v_3027 | ~v_105;
assign x_1802 = v_3027 | ~v_104;
assign x_1803 = v_3027 | ~v_76;
assign x_1804 = v_3027 | ~v_74;
assign x_1805 = v_3027 | ~v_73;
assign x_1806 = ~v_80 | v_98 | v_3026;
assign x_1807 = ~v_88 | ~v_98 | v_3025;
assign x_1808 = ~v_86 | ~v_97 | v_3024;
assign x_1809 = ~v_78 | v_97 | v_3023;
assign x_1810 = v_3022 | ~v_2945;
assign x_1811 = v_3022 | ~v_803;
assign x_1812 = v_3022 | ~v_2946;
assign x_1813 = v_3022 | ~v_804;
assign x_1814 = v_3022 | ~v_2947;
assign x_1815 = v_3022 | ~v_925;
assign x_1816 = v_3022 | ~v_926;
assign x_1817 = v_3022 | ~v_2948;
assign x_1818 = v_3022 | ~v_2951;
assign x_1819 = v_3022 | ~v_927;
assign x_1820 = v_3022 | ~v_928;
assign x_1821 = v_3022 | ~v_3018;
assign x_1822 = v_3022 | ~v_3019;
assign x_1823 = v_3022 | ~v_900;
assign x_1824 = v_3022 | ~v_3020;
assign x_1825 = v_3022 | ~v_3021;
assign x_1826 = v_3022 | ~v_902;
assign x_1827 = v_3022 | ~v_2953;
assign x_1828 = v_3022 | ~v_111;
assign x_1829 = v_3022 | ~v_110;
assign x_1830 = v_3022 | ~v_103;
assign x_1831 = v_3022 | ~v_102;
assign x_1832 = v_3022 | ~v_101;
assign x_1833 = v_3022 | ~v_100;
assign x_1834 = v_3022 | ~v_51;
assign x_1835 = v_3022 | ~v_49;
assign x_1836 = v_3022 | ~v_48;
assign x_1837 = ~v_55 | v_98 | v_3021;
assign x_1838 = ~v_63 | ~v_98 | v_3020;
assign x_1839 = ~v_53 | v_97 | v_3019;
assign x_1840 = ~v_61 | ~v_97 | v_3018;
assign x_1841 = v_3017 | ~v_2934;
assign x_1842 = v_3017 | ~v_792;
assign x_1843 = v_3017 | ~v_2935;
assign x_1844 = v_3017 | ~v_793;
assign x_1845 = v_3017 | ~v_2936;
assign x_1846 = v_3017 | ~v_2937;
assign x_1847 = v_3017 | ~v_920;
assign x_1848 = v_3017 | ~v_921;
assign x_1849 = v_3017 | ~v_885;
assign x_1850 = v_3017 | ~v_3013;
assign x_1851 = v_3017 | ~v_3014;
assign x_1852 = v_3017 | ~v_2939;
assign x_1853 = v_3017 | ~v_922;
assign x_1854 = v_3017 | ~v_3015;
assign x_1855 = v_3017 | ~v_890;
assign x_1856 = v_3017 | ~v_923;
assign x_1857 = v_3017 | ~v_3016;
assign x_1858 = v_3017 | ~v_109;
assign x_1859 = v_3017 | ~v_108;
assign x_1860 = v_3017 | ~v_96;
assign x_1861 = v_3017 | ~v_95;
assign x_1862 = v_3017 | ~v_94;
assign x_1863 = v_3017 | ~v_93;
assign x_1864 = v_3017 | ~v_2943;
assign x_1865 = v_3017 | ~v_25;
assign x_1866 = v_3017 | ~v_23;
assign x_1867 = v_3017 | ~v_22;
assign x_1868 = ~v_30 | v_98 | v_3016;
assign x_1869 = ~v_36 | ~v_97 | v_3015;
assign x_1870 = ~v_38 | ~v_98 | v_3014;
assign x_1871 = ~v_28 | v_97 | v_3013;
assign x_1872 = ~v_3011 | ~v_3006 | ~v_3001 | v_3012;
assign x_1873 = v_3011 | ~v_680;
assign x_1874 = v_3011 | ~v_681;
assign x_1875 = v_3011 | ~v_682;
assign x_1876 = v_3011 | ~v_683;
assign x_1877 = v_3011 | ~v_3007;
assign x_1878 = v_3011 | ~v_2959;
assign x_1879 = v_3011 | ~v_2962;
assign x_1880 = v_3011 | ~v_3008;
assign x_1881 = v_3011 | ~v_3009;
assign x_1882 = v_3011 | ~v_686;
assign x_1883 = v_3011 | ~v_687;
assign x_1884 = v_3011 | ~v_2989;
assign x_1885 = v_3011 | ~v_2990;
assign x_1886 = v_3011 | ~v_2991;
assign x_1887 = v_3011 | ~v_2992;
assign x_1888 = v_3011 | ~v_688;
assign x_1889 = v_3011 | ~v_689;
assign x_1890 = v_3011 | ~v_3010;
assign x_1891 = v_3011 | ~v_132;
assign x_1892 = v_3011 | ~v_113;
assign x_1893 = v_3011 | ~v_112;
assign x_1894 = v_3011 | ~v_106;
assign x_1895 = v_3011 | ~v_105;
assign x_1896 = v_3011 | ~v_104;
assign x_1897 = v_3011 | ~v_76;
assign x_1898 = v_3011 | ~v_75;
assign x_1899 = v_3011 | ~v_74;
assign x_1900 = ~v_79 | v_97 | v_3010;
assign x_1901 = ~v_90 | ~v_98 | v_3009;
assign x_1902 = ~v_82 | v_98 | v_3008;
assign x_1903 = ~v_87 | ~v_97 | v_3007;
assign x_1904 = v_3006 | ~v_2948;
assign x_1905 = v_3006 | ~v_2951;
assign x_1906 = v_3006 | ~v_665;
assign x_1907 = v_3006 | ~v_666;
assign x_1908 = v_3006 | ~v_2980;
assign x_1909 = v_3006 | ~v_2981;
assign x_1910 = v_3006 | ~v_2982;
assign x_1911 = v_3006 | ~v_2983;
assign x_1912 = v_3006 | ~v_667;
assign x_1913 = v_3006 | ~v_668;
assign x_1914 = v_3006 | ~v_669;
assign x_1915 = v_3006 | ~v_670;
assign x_1916 = v_3006 | ~v_3002;
assign x_1917 = v_3006 | ~v_3003;
assign x_1918 = v_3006 | ~v_3004;
assign x_1919 = v_3006 | ~v_677;
assign x_1920 = v_3006 | ~v_678;
assign x_1921 = v_3006 | ~v_131;
assign x_1922 = v_3006 | ~v_3005;
assign x_1923 = v_3006 | ~v_111;
assign x_1924 = v_3006 | ~v_110;
assign x_1925 = v_3006 | ~v_102;
assign x_1926 = v_3006 | ~v_101;
assign x_1927 = v_3006 | ~v_100;
assign x_1928 = v_3006 | ~v_51;
assign x_1929 = v_3006 | ~v_50;
assign x_1930 = v_3006 | ~v_49;
assign x_1931 = ~v_57 | v_98 | v_3005;
assign x_1932 = ~v_65 | ~v_98 | v_3004;
assign x_1933 = ~v_54 | v_97 | v_3003;
assign x_1934 = ~v_62 | ~v_97 | v_3002;
assign x_1935 = v_3001 | ~v_646;
assign x_1936 = v_3001 | ~v_2997;
assign x_1937 = v_3001 | ~v_2998;
assign x_1938 = v_3001 | ~v_2939;
assign x_1939 = v_3001 | ~v_649;
assign x_1940 = v_3001 | ~v_650;
assign x_1941 = v_3001 | ~v_2972;
assign x_1942 = v_3001 | ~v_2973;
assign x_1943 = v_3001 | ~v_2974;
assign x_1944 = v_3001 | ~v_2975;
assign x_1945 = v_3001 | ~v_651;
assign x_1946 = v_3001 | ~v_652;
assign x_1947 = v_3001 | ~v_653;
assign x_1948 = v_3001 | ~v_654;
assign x_1949 = v_3001 | ~v_661;
assign x_1950 = v_3001 | ~v_2999;
assign x_1951 = v_3001 | ~v_3000;
assign x_1952 = v_3001 | ~v_128;
assign x_1953 = v_3001 | ~v_109;
assign x_1954 = v_3001 | ~v_108;
assign x_1955 = v_3001 | ~v_95;
assign x_1956 = v_3001 | ~v_94;
assign x_1957 = v_3001 | ~v_93;
assign x_1958 = v_3001 | ~v_2943;
assign x_1959 = v_3001 | ~v_25;
assign x_1960 = v_3001 | ~v_24;
assign x_1961 = v_3001 | ~v_23;
assign x_1962 = ~v_32 | v_98 | v_3000;
assign x_1963 = ~v_40 | ~v_98 | v_2999;
assign x_1964 = ~v_37 | ~v_97 | v_2998;
assign x_1965 = ~v_29 | v_97 | v_2997;
assign x_1966 = v_2996 | ~v_2967;
assign x_1967 = v_2996 | ~v_2995;
assign x_1968 = v_2996 | ~v_698;
assign x_1969 = v_2996 | ~v_699;
assign x_1970 = v_2996 | ~v_700;
assign x_1971 = v_2996 | ~v_701;
assign x_1972 = ~v_2994 | ~v_2985 | ~v_2976 | v_2995;
assign x_1973 = v_2994 | ~v_871;
assign x_1974 = v_2994 | ~v_872;
assign x_1975 = v_2994 | ~v_873;
assign x_1976 = v_2994 | ~v_874;
assign x_1977 = v_2994 | ~v_2986;
assign x_1978 = v_2994 | ~v_2987;
assign x_1979 = v_2994 | ~v_2988;
assign x_1980 = v_2994 | ~v_2959;
assign x_1981 = v_2994 | ~v_2962;
assign x_1982 = v_2994 | ~v_763;
assign x_1983 = v_2994 | ~v_764;
assign x_1984 = v_2994 | ~v_2989;
assign x_1985 = v_2994 | ~v_2990;
assign x_1986 = v_2994 | ~v_2991;
assign x_1987 = v_2994 | ~v_2992;
assign x_1988 = v_2994 | ~v_688;
assign x_1989 = v_2994 | ~v_689;
assign x_1990 = v_2994 | ~v_2993;
assign x_1991 = v_2994 | ~v_132;
assign x_1992 = v_2994 | ~v_113;
assign x_1993 = v_2994 | ~v_112;
assign x_1994 = v_2994 | ~v_104;
assign x_1995 = v_2994 | ~v_76;
assign x_1996 = v_2994 | ~v_75;
assign x_1997 = v_2994 | ~v_74;
assign x_1998 = v_2994 | ~v_72;
assign x_1999 = v_2994 | ~v_70;
assign x_2000 = ~v_26 | ~v_87 | v_2993;
assign x_2001 = ~v_88 | ~v_124 | v_2992;
assign x_2002 = ~v_80 | v_124 | v_2991;
assign x_2003 = ~v_86 | ~v_123 | v_2990;
assign x_2004 = ~v_78 | v_123 | v_2989;
assign x_2005 = ~v_26 | ~v_90 | v_2988;
assign x_2006 = v_26 | ~v_82 | v_2987;
assign x_2007 = v_26 | ~v_79 | v_2986;
assign x_2008 = v_2985 | ~v_866;
assign x_2009 = v_2985 | ~v_867;
assign x_2010 = v_2985 | ~v_2977;
assign x_2011 = v_2985 | ~v_2978;
assign x_2012 = v_2985 | ~v_2948;
assign x_2013 = v_2985 | ~v_750;
assign x_2014 = v_2985 | ~v_2951;
assign x_2015 = v_2985 | ~v_2979;
assign x_2016 = v_2985 | ~v_2980;
assign x_2017 = v_2985 | ~v_2981;
assign x_2018 = v_2985 | ~v_2982;
assign x_2019 = v_2985 | ~v_2983;
assign x_2020 = v_2985 | ~v_868;
assign x_2021 = v_2985 | ~v_669;
assign x_2022 = v_2985 | ~v_670;
assign x_2023 = v_2985 | ~v_869;
assign x_2024 = v_2985 | ~v_2984;
assign x_2025 = v_2985 | ~v_757;
assign x_2026 = v_2985 | ~v_131;
assign x_2027 = v_2985 | ~v_111;
assign x_2028 = v_2985 | ~v_110;
assign x_2029 = v_2985 | ~v_100;
assign x_2030 = v_2985 | ~v_51;
assign x_2031 = v_2985 | ~v_50;
assign x_2032 = v_2985 | ~v_49;
assign x_2033 = v_2985 | ~v_47;
assign x_2034 = v_2985 | ~v_45;
assign x_2035 = ~v_26 | ~v_62 | v_2984;
assign x_2036 = ~v_63 | ~v_124 | v_2983;
assign x_2037 = ~v_55 | v_124 | v_2982;
assign x_2038 = ~v_61 | ~v_123 | v_2981;
assign x_2039 = ~v_53 | v_123 | v_2980;
assign x_2040 = v_26 | ~v_54 | v_2979;
assign x_2041 = ~v_26 | ~v_65 | v_2978;
assign x_2042 = v_26 | ~v_57 | v_2977;
assign x_2043 = v_2976 | ~v_861;
assign x_2044 = v_2976 | ~v_862;
assign x_2045 = v_2976 | ~v_2968;
assign x_2046 = v_2976 | ~v_2969;
assign x_2047 = v_2976 | ~v_2970;
assign x_2048 = v_2976 | ~v_2939;
assign x_2049 = v_2976 | ~v_739;
assign x_2050 = v_2976 | ~v_2971;
assign x_2051 = v_2976 | ~v_2972;
assign x_2052 = v_2976 | ~v_2973;
assign x_2053 = v_2976 | ~v_2974;
assign x_2054 = v_2976 | ~v_2975;
assign x_2055 = v_2976 | ~v_653;
assign x_2056 = v_2976 | ~v_654;
assign x_2057 = v_2976 | ~v_863;
assign x_2058 = v_2976 | ~v_864;
assign x_2059 = v_2976 | ~v_746;
assign x_2060 = v_2976 | ~v_128;
assign x_2061 = v_2976 | ~v_109;
assign x_2062 = v_2976 | ~v_108;
assign x_2063 = v_2976 | ~v_93;
assign x_2064 = v_2976 | ~v_2943;
assign x_2065 = v_2976 | ~v_25;
assign x_2066 = v_2976 | ~v_24;
assign x_2067 = v_2976 | ~v_23;
assign x_2068 = v_2976 | ~v_21;
assign x_2069 = v_2976 | ~v_19;
assign x_2070 = ~v_38 | ~v_124 | v_2975;
assign x_2071 = ~v_30 | v_124 | v_2974;
assign x_2072 = ~v_36 | ~v_123 | v_2973;
assign x_2073 = ~v_28 | v_123 | v_2972;
assign x_2074 = ~v_26 | ~v_40 | v_2971;
assign x_2075 = ~v_26 | ~v_37 | v_2970;
assign x_2076 = ~v_32 | v_26 | v_2969;
assign x_2077 = ~v_29 | v_26 | v_2968;
assign x_2078 = ~v_2966 | ~v_2955 | ~v_2944 | v_2967;
assign x_2079 = v_2966 | ~v_835;
assign x_2080 = v_2966 | ~v_836;
assign x_2081 = v_2966 | ~v_2956;
assign x_2082 = v_2966 | ~v_814;
assign x_2083 = v_2966 | ~v_2957;
assign x_2084 = v_2966 | ~v_815;
assign x_2085 = v_2966 | ~v_2958;
assign x_2086 = v_2966 | ~v_837;
assign x_2087 = v_2966 | ~v_838;
assign x_2088 = v_2966 | ~v_2959;
assign x_2089 = v_2966 | ~v_2960;
assign x_2090 = v_2966 | ~v_2961;
assign x_2091 = v_2966 | ~v_2962;
assign x_2092 = v_2966 | ~v_726;
assign x_2093 = v_2966 | ~v_2963;
assign x_2094 = v_2966 | ~v_731;
assign x_2095 = v_2966 | ~v_2964;
assign x_2096 = v_2966 | ~v_2965;
assign x_2097 = v_2966 | ~v_106;
assign x_2098 = v_2966 | ~v_105;
assign x_2099 = v_2966 | ~v_104;
assign x_2100 = v_2966 | ~v_76;
assign x_2101 = v_2966 | ~v_75;
assign x_2102 = v_2966 | ~v_74;
assign x_2103 = v_2966 | ~v_73;
assign x_2104 = v_2966 | ~v_71;
assign x_2105 = v_2966 | ~v_68;
assign x_2106 = ~v_87 | ~v_114 | v_2965;
assign x_2107 = ~v_26 | ~v_88 | v_2964;
assign x_2108 = ~v_26 | ~v_86 | v_2963;
assign x_2109 = ~v_26 | ~v_85 | v_2962;
assign x_2110 = v_26 | ~v_80 | v_2961;
assign x_2111 = v_26 | ~v_78 | v_2960;
assign x_2112 = v_26 | ~v_77 | v_2959;
assign x_2113 = ~v_79 | v_114 | v_2958;
assign x_2114 = ~v_90 | ~v_115 | v_2957;
assign x_2115 = ~v_82 | v_115 | v_2956;
assign x_2116 = v_2955 | ~v_830;
assign x_2117 = v_2955 | ~v_831;
assign x_2118 = v_2955 | ~v_2945;
assign x_2119 = v_2955 | ~v_803;
assign x_2120 = v_2955 | ~v_2946;
assign x_2121 = v_2955 | ~v_804;
assign x_2122 = v_2955 | ~v_2947;
assign x_2123 = v_2955 | ~v_2948;
assign x_2124 = v_2955 | ~v_2949;
assign x_2125 = v_2955 | ~v_2950;
assign x_2126 = v_2955 | ~v_714;
assign x_2127 = v_2955 | ~v_2951;
assign x_2128 = v_2955 | ~v_2952;
assign x_2129 = v_2955 | ~v_832;
assign x_2130 = v_2955 | ~v_833;
assign x_2131 = v_2955 | ~v_721;
assign x_2132 = v_2955 | ~v_2953;
assign x_2133 = v_2955 | ~v_102;
assign x_2134 = v_2955 | ~v_101;
assign x_2135 = v_2955 | ~v_100;
assign x_2136 = v_2955 | ~v_2954;
assign x_2137 = v_2955 | ~v_51;
assign x_2138 = v_2955 | ~v_50;
assign x_2139 = v_2955 | ~v_49;
assign x_2140 = v_2955 | ~v_48;
assign x_2141 = v_2955 | ~v_46;
assign x_2142 = v_2955 | ~v_43;
assign x_2143 = ~v_26 | ~v_61 | v_2954;
assign x_2144 = ~v_62 | ~v_114 | v_2953;
assign x_2145 = ~v_26 | ~v_63 | v_2952;
assign x_2146 = ~v_26 | ~v_60 | v_2951;
assign x_2147 = v_26 | ~v_55 | v_2950;
assign x_2148 = v_26 | ~v_53 | v_2949;
assign x_2149 = v_26 | ~v_52 | v_2948;
assign x_2150 = ~v_54 | v_114 | v_2947;
assign x_2151 = ~v_65 | ~v_115 | v_2946;
assign x_2152 = ~v_57 | v_115 | v_2945;
assign x_2153 = v_2944 | ~v_825;
assign x_2154 = v_2944 | ~v_826;
assign x_2155 = v_2944 | ~v_2934;
assign x_2156 = v_2944 | ~v_792;
assign x_2157 = v_2944 | ~v_2935;
assign x_2158 = v_2944 | ~v_793;
assign x_2159 = v_2944 | ~v_2936;
assign x_2160 = v_2944 | ~v_2937;
assign x_2161 = v_2944 | ~v_2938;
assign x_2162 = v_2944 | ~v_2939;
assign x_2163 = v_2944 | ~v_2940;
assign x_2164 = v_2944 | ~v_2941;
assign x_2165 = v_2944 | ~v_705;
assign x_2166 = v_2944 | ~v_706;
assign x_2167 = v_2944 | ~v_2942;
assign x_2168 = v_2944 | ~v_827;
assign x_2169 = v_2944 | ~v_828;
assign x_2170 = v_2944 | ~v_95;
assign x_2171 = v_2944 | ~v_94;
assign x_2172 = v_2944 | ~v_93;
assign x_2173 = v_2944 | ~v_2943;
assign x_2174 = v_2944 | ~v_25;
assign x_2175 = v_2944 | ~v_24;
assign x_2176 = v_2944 | ~v_23;
assign x_2177 = v_2944 | ~v_22;
assign x_2178 = v_2944 | ~v_20;
assign x_2179 = v_2944 | ~v_17;
assign x_2180 = ~v_27 | v_26 | v_2943;
assign x_2181 = ~v_28 | v_26 | v_2942;
assign x_2182 = ~v_26 | ~v_38 | v_2941;
assign x_2183 = ~v_26 | ~v_36 | v_2940;
assign x_2184 = ~v_26 | ~v_35 | v_2939;
assign x_2185 = ~v_30 | v_26 | v_2938;
assign x_2186 = ~v_37 | ~v_114 | v_2937;
assign x_2187 = ~v_29 | v_114 | v_2936;
assign x_2188 = ~v_40 | ~v_115 | v_2935;
assign x_2189 = ~v_32 | v_115 | v_2934;
assign x_2190 = ~v_2932 | ~v_2931 | v_2933;
assign x_2191 = v_2932 | ~v_2274;
assign x_2192 = v_2932 | ~v_1600;
assign x_2193 = v_2932 | ~v_585;
assign x_2194 = v_2932 | ~v_26;
assign x_2195 = v_2931 | ~v_2909;
assign x_2196 = v_2931 | ~v_2928;
assign x_2197 = v_2931 | ~v_2929;
assign x_2198 = v_2931 | ~v_2854;
assign x_2199 = v_2931 | ~v_2859;
assign x_2200 = v_2931 | ~v_2930;
assign x_2201 = v_2931 | ~v_2860;
assign x_2202 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2858 | ~v_2911 | v_2930;
assign x_2203 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2853 | ~v_2832 | v_2929;
assign x_2204 = ~v_2927 | ~v_2913 | v_2928;
assign x_2205 = v_2927 | ~v_2914;
assign x_2206 = v_2927 | ~v_2915;
assign x_2207 = v_2927 | ~v_2920;
assign x_2208 = v_2927 | ~v_2925;
assign x_2209 = v_2927 | ~v_2926;
assign x_2210 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2853 | v_2926;
assign x_2211 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2858 | ~v_2924 | v_2925;
assign x_2212 = v_2924 | ~v_2921;
assign x_2213 = v_2924 | ~v_2922;
assign x_2214 = v_2924 | ~v_2923;
assign x_2215 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2848 | v_2923;
assign x_2216 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2865 | ~v_2853 | v_2922;
assign x_2217 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2825 | ~v_2886 | v_2921;
assign x_2218 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2919 | ~v_2764 | v_2920;
assign x_2219 = v_2919 | ~v_2916;
assign x_2220 = v_2919 | ~v_2917;
assign x_2221 = v_2919 | ~v_2918;
assign x_2222 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2886 | v_2918;
assign x_2223 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2891 | ~v_2853 | v_2917;
assign x_2224 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2848 | ~v_2896 | v_2916;
assign x_2225 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2858 | ~v_2848 | v_2915;
assign x_2226 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2886 | ~v_2764 | v_2914;
assign x_2227 = v_2913 | ~v_2910;
assign x_2228 = v_2913 | ~v_2912;
assign x_2229 = v_2913 | ~v_2793;
assign x_2230 = v_2913 | ~v_2826;
assign x_2231 = v_2913 | ~v_2831;
assign x_2232 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2809 | ~v_2911 | v_2912;
assign x_2233 = v_2911 | ~v_2867;
assign x_2234 = v_2911 | ~v_2868;
assign x_2235 = v_2911 | ~v_2869;
assign x_2236 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2792 | ~v_2861 | v_2910;
assign x_2237 = ~v_2908 | ~v_2870 | v_2909;
assign x_2238 = v_2908 | ~v_2899;
assign x_2239 = v_2908 | ~v_2904;
assign x_2240 = v_2908 | ~v_2905;
assign x_2241 = v_2908 | ~v_2906;
assign x_2242 = v_2908 | ~v_2907;
assign x_2243 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2858 | v_2907;
assign x_2244 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2809 | ~v_2853 | v_2906;
assign x_2245 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2896 | ~v_2764 | v_2905;
assign x_2246 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2853 | ~v_2903 | v_2904;
assign x_2247 = v_2903 | ~v_2900;
assign x_2248 = v_2903 | ~v_2901;
assign x_2249 = v_2903 | ~v_2902;
assign x_2250 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2809 | v_2902;
assign x_2251 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2858 | ~v_2792 | v_2901;
assign x_2252 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2830 | ~v_2896 | v_2900;
assign x_2253 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2764 | ~v_2898 | v_2899;
assign x_2254 = v_2898 | ~v_2887;
assign x_2255 = v_2898 | ~v_2892;
assign x_2256 = v_2898 | ~v_2897;
assign x_2257 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2896 | v_2897;
assign x_2258 = v_2896 | ~v_2893;
assign x_2259 = v_2896 | ~v_2894;
assign x_2260 = v_2896 | ~v_2895;
assign x_2261 = v_75 | v_74 | v_73 | v_106 | v_105 | v_104 | v_113 | v_112 | v_121 | ~v_2807 | ~v_2884 | ~v_2883 | ~v_2882 | ~v_2881 | ~v_332 | ~v_331 | ~v_180 | ~v_179 | ~v_2806 | ~v_2805 | ~v_2759 | ~v_2756 | ~v_2804 | ~v_230 | ~v_229 | ~v_330 | ~v_329 | v_2895;
assign x_2262 = v_50 | v_49 | v_48 | v_101 | v_100 | ~v_2802 | v_102 | v_111 | v_110 | v_120 | ~v_2879 | ~v_225 | ~v_224 | ~v_2801 | ~v_2800 | ~v_2799 | ~v_2878 | ~v_2877 | ~v_2876 | ~v_327 | ~v_326 | ~v_161 | ~v_160 | ~v_2748 | ~v_2745 | ~v_325 | ~v_324 | v_2894;
assign x_2263 = v_24 | v_23 | v_22 | ~v_2740 | v_95 | v_94 | v_93 | v_108 | v_109 | v_117 | ~v_2797 | ~v_2796 | ~v_208 | ~v_2874 | ~v_2873 | ~v_2872 | ~v_2871 | ~v_322 | ~v_321 | ~v_142 | ~v_141 | ~v_2736 | ~v_2795 | ~v_2794 | ~v_193 | ~v_320 | ~v_319 | v_2893;
assign x_2264 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2858 | ~v_2891 | v_2892;
assign x_2265 = v_2891 | ~v_2888;
assign x_2266 = v_2891 | ~v_2889;
assign x_2267 = v_2891 | ~v_2890;
assign x_2268 = v_76 | v_75 | v_74 | v_73 | v_72 | v_70 | v_104 | v_113 | v_112 | ~v_2790 | ~v_2884 | ~v_2883 | ~v_2882 | ~v_2881 | ~v_180 | ~v_179 | ~v_313 | ~v_312 | ~v_311 | ~v_310 | ~v_2759 | ~v_2756 | ~v_2785 | ~v_2784 | ~v_2783 | ~v_309 | ~v_308 | v_2890;
assign x_2269 = v_50 | v_51 | v_49 | v_48 | v_45 | v_47 | v_100 | v_111 | v_110 | ~v_2879 | ~v_304 | ~v_2781 | ~v_301 | ~v_300 | ~v_2878 | ~v_2877 | ~v_2876 | ~v_161 | ~v_160 | ~v_299 | ~v_298 | ~v_2776 | ~v_2748 | ~v_297 | ~v_2745 | ~v_2775 | ~v_2774 | v_2889;
assign x_2270 = v_25 | v_24 | v_23 | v_22 | v_21 | v_19 | ~v_2740 | v_93 | v_108 | v_109 | ~v_293 | ~v_290 | ~v_289 | ~v_2874 | ~v_2873 | ~v_2872 | ~v_2871 | ~v_142 | ~v_141 | ~v_288 | ~v_287 | ~v_2768 | ~v_286 | ~v_2736 | ~v_2767 | ~v_2766 | ~v_2765 | v_2888;
assign x_2271 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2809 | ~v_2886 | v_2887;
assign x_2272 = v_2886 | ~v_2875;
assign x_2273 = v_2886 | ~v_2880;
assign x_2274 = v_2886 | ~v_2885;
assign x_2275 = v_76 | v_73 | v_107 | v_106 | v_105 | v_104 | v_127 | v_113 | v_112 | ~v_2884 | ~v_2883 | ~v_2882 | ~v_2881 | ~v_2846 | ~v_2845 | ~v_2844 | ~v_2843 | ~v_184 | ~v_183 | ~v_182 | ~v_181 | ~v_180 | ~v_179 | ~v_2759 | ~v_2756 | ~v_178 | ~v_177 | v_2885;
assign x_2276 = v_2884 | v_114;
assign x_2277 = v_2884 | v_86;
assign x_2278 = v_2883 | ~v_114;
assign x_2279 = v_2883 | v_78;
assign x_2280 = v_2882 | v_115;
assign x_2281 = v_2882 | v_88;
assign x_2282 = v_2881 | ~v_115;
assign x_2283 = v_2881 | v_80;
assign x_2284 = v_51 | v_48 | v_103 | v_101 | v_100 | v_102 | v_111 | v_110 | v_126 | ~v_2879 | ~v_2878 | ~v_2877 | ~v_2876 | ~v_2841 | ~v_2840 | ~v_2839 | ~v_2838 | ~v_165 | ~v_164 | ~v_163 | ~v_162 | ~v_161 | ~v_160 | ~v_2748 | ~v_2745 | ~v_159 | ~v_158 | v_2880;
assign x_2285 = v_2879 | v_114;
assign x_2286 = v_2879 | v_61;
assign x_2287 = v_2878 | ~v_114;
assign x_2288 = v_2878 | v_53;
assign x_2289 = v_2877 | v_115;
assign x_2290 = v_2877 | v_63;
assign x_2291 = v_2876 | ~v_115;
assign x_2292 = v_2876 | v_55;
assign x_2293 = v_25 | v_22 | ~v_2740 | v_96 | v_95 | v_94 | v_93 | v_108 | v_109 | v_122 | ~v_2874 | ~v_2873 | ~v_2872 | ~v_2871 | ~v_2836 | ~v_2835 | ~v_2834 | ~v_2833 | ~v_146 | ~v_145 | ~v_144 | ~v_143 | ~v_142 | ~v_141 | ~v_2736 | ~v_140 | ~v_139 | v_2875;
assign x_2294 = v_2874 | v_114;
assign x_2295 = v_2874 | v_36;
assign x_2296 = v_2873 | ~v_114;
assign x_2297 = v_2873 | v_28;
assign x_2298 = v_2872 | v_115;
assign x_2299 = v_2872 | v_38;
assign x_2300 = v_2871 | ~v_115;
assign x_2301 = v_2871 | v_30;
assign x_2302 = v_2870 | ~v_2849;
assign x_2303 = v_2870 | ~v_2866;
assign x_2304 = v_2870 | ~v_2867;
assign x_2305 = v_2870 | ~v_2868;
assign x_2306 = v_2870 | ~v_2869;
assign x_2307 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2825 | v_2869;
assign x_2308 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2865 | ~v_2764 | v_2868;
assign x_2309 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2848 | ~v_2830 | v_2867;
assign x_2310 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2865 | ~v_2861 | v_2866;
assign x_2311 = v_2865 | ~v_2862;
assign x_2312 = v_2865 | ~v_2863;
assign x_2313 = v_2865 | ~v_2864;
assign x_2314 = v_75 | v_74 | v_73 | v_72 | v_70 | v_104 | v_113 | v_112 | v_121 | ~v_461 | ~v_2790 | ~v_2823 | ~v_311 | ~v_310 | ~v_457 | ~v_456 | ~v_455 | ~v_2759 | ~v_2756 | ~v_2785 | ~v_2784 | ~v_2783 | ~v_2822 | ~v_2821 | ~v_2820 | ~v_454 | ~v_453 | v_2864;
assign x_2315 = v_50 | v_49 | v_48 | v_45 | v_47 | v_100 | v_111 | v_110 | v_120 | ~v_450 | ~v_449 | ~v_448 | ~v_2818 | ~v_2817 | ~v_447 | ~v_304 | ~v_2781 | ~v_2816 | ~v_444 | ~v_2815 | ~v_2776 | ~v_2748 | ~v_297 | ~v_443 | ~v_2745 | ~v_2775 | ~v_2774 | v_2863;
assign x_2316 = v_24 | v_23 | v_22 | v_21 | v_19 | ~v_2740 | ~v_2813 | v_93 | v_108 | v_109 | v_117 | ~v_439 | ~v_438 | ~v_437 | ~v_293 | ~v_2812 | ~v_2768 | ~v_286 | ~v_434 | ~v_433 | ~v_2736 | ~v_2767 | ~v_2766 | ~v_2765 | ~v_2811 | ~v_2810 | ~v_432 | v_2862;
assign x_2317 = v_2861 | ~v_2854;
assign x_2318 = v_2861 | ~v_2859;
assign x_2319 = v_2861 | ~v_2860;
assign x_2320 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2764 | v_2860;
assign x_2321 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2858 | ~v_2825 | v_2859;
assign x_2322 = v_2858 | ~v_2855;
assign x_2323 = v_2858 | ~v_2856;
assign x_2324 = v_2858 | ~v_2857;
assign x_2325 = v_76 | v_68 | v_74 | v_73 | v_71 | v_107 | v_106 | v_105 | v_104 | ~v_281 | ~v_2761 | ~v_278 | ~v_2760 | ~v_2807 | ~v_275 | ~v_274 | ~v_273 | ~v_272 | ~v_2806 | ~v_2805 | ~v_2759 | ~v_2758 | ~v_2757 | ~v_2756 | ~v_2804 | ~v_230 | ~v_229 | v_2857;
assign x_2326 = v_51 | v_49 | v_48 | v_46 | v_43 | ~v_2751 | v_103 | v_101 | v_100 | ~v_2802 | v_102 | ~v_270 | ~v_225 | ~v_269 | ~v_224 | ~v_2801 | ~v_2800 | ~v_268 | ~v_265 | ~v_2799 | ~v_2749 | ~v_2748 | ~v_262 | ~v_261 | ~v_2747 | ~v_2746 | ~v_2745 | v_2856;
assign x_2327 = v_25 | v_23 | v_22 | v_20 | v_17 | ~v_2740 | v_96 | v_95 | v_94 | v_93 | ~v_259 | ~v_2797 | ~v_2796 | ~v_258 | ~v_208 | ~v_2739 | ~v_253 | ~v_252 | ~v_251 | ~v_250 | ~v_2738 | ~v_2737 | ~v_2736 | ~v_2735 | ~v_2795 | ~v_2794 | ~v_193 | v_2855;
assign x_2328 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2830 | ~v_2853 | v_2854;
assign x_2329 = v_2853 | ~v_2850;
assign x_2330 = v_2853 | ~v_2851;
assign x_2331 = v_2853 | ~v_2852;
assign x_2332 = v_76 | v_68 | v_75 | v_73 | v_71 | v_106 | v_105 | v_104 | v_127 | ~v_2761 | ~v_278 | ~v_2760 | ~v_2846 | ~v_2845 | ~v_2844 | ~v_2843 | ~v_402 | ~v_401 | ~v_182 | ~v_181 | ~v_273 | ~v_2759 | ~v_2758 | ~v_2757 | ~v_2756 | ~v_400 | ~v_399 | v_2852;
assign x_2333 = v_50 | v_51 | v_48 | v_46 | v_43 | ~v_2751 | v_101 | v_100 | v_102 | v_126 | ~v_268 | ~v_2841 | ~v_2840 | ~v_2839 | ~v_2838 | ~v_397 | ~v_396 | ~v_163 | ~v_162 | ~v_2749 | ~v_2748 | ~v_261 | ~v_2747 | ~v_2746 | ~v_2745 | ~v_395 | ~v_394 | v_2851;
assign x_2334 = v_25 | v_24 | v_22 | v_20 | v_17 | ~v_2740 | v_95 | v_94 | v_93 | v_122 | ~v_2836 | ~v_2835 | ~v_2834 | ~v_2833 | ~v_392 | ~v_391 | ~v_144 | ~v_143 | ~v_2739 | ~v_253 | ~v_252 | ~v_2738 | ~v_2737 | ~v_2736 | ~v_2735 | ~v_390 | ~v_389 | v_2850;
assign x_2335 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2848 | ~v_2832 | v_2849;
assign x_2336 = v_2848 | ~v_2837;
assign x_2337 = v_2848 | ~v_2842;
assign x_2338 = v_2848 | ~v_2847;
assign x_2339 = v_76 | v_75 | v_73 | v_106 | v_105 | v_104 | v_127 | v_113 | v_112 | ~v_2823 | ~v_2846 | ~v_2845 | ~v_2844 | ~v_2843 | ~v_182 | ~v_181 | ~v_501 | ~v_500 | ~v_2759 | ~v_2756 | ~v_2822 | ~v_2821 | ~v_2820 | ~v_454 | ~v_453 | ~v_499 | ~v_498 | v_2847;
assign x_2340 = v_2846 | v_123;
assign x_2341 = v_2846 | v_87;
assign x_2342 = v_2845 | ~v_123;
assign x_2343 = v_2845 | v_79;
assign x_2344 = v_2844 | v_124;
assign x_2345 = v_2844 | v_90;
assign x_2346 = v_2843 | ~v_124;
assign x_2347 = v_2843 | v_82;
assign x_2348 = v_50 | v_51 | v_48 | v_101 | v_100 | v_102 | v_111 | v_110 | v_126 | ~v_449 | ~v_2818 | ~v_2817 | ~v_447 | ~v_2816 | ~v_2815 | ~v_2841 | ~v_2840 | ~v_2839 | ~v_2838 | ~v_163 | ~v_162 | ~v_496 | ~v_495 | ~v_2748 | ~v_2745 | ~v_494 | ~v_493 | v_2842;
assign x_2349 = v_2841 | v_123;
assign x_2350 = v_2841 | v_62;
assign x_2351 = v_2840 | ~v_123;
assign x_2352 = v_2840 | v_54;
assign x_2353 = v_2839 | v_124;
assign x_2354 = v_2839 | v_65;
assign x_2355 = v_2838 | ~v_124;
assign x_2356 = v_2838 | v_57;
assign x_2357 = v_25 | v_24 | v_22 | ~v_2740 | ~v_2813 | v_95 | v_94 | v_93 | v_108 | v_109 | v_122 | ~v_437 | ~v_2812 | ~v_2836 | ~v_2835 | ~v_2834 | ~v_2833 | ~v_144 | ~v_143 | ~v_491 | ~v_490 | ~v_2736 | ~v_2811 | ~v_2810 | ~v_432 | ~v_489 | ~v_488 | v_2837;
assign x_2358 = v_2836 | v_123;
assign x_2359 = v_2836 | v_37;
assign x_2360 = v_2835 | ~v_123;
assign x_2361 = v_2835 | v_29;
assign x_2362 = v_2834 | v_124;
assign x_2363 = v_2834 | v_40;
assign x_2364 = v_2833 | ~v_124;
assign x_2365 = v_2833 | v_32;
assign x_2366 = v_2832 | ~v_2793;
assign x_2367 = v_2832 | ~v_2826;
assign x_2368 = v_2832 | ~v_2831;
assign x_2369 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2830 | v_2831;
assign x_2370 = v_2830 | ~v_2827;
assign x_2371 = v_2830 | ~v_2828;
assign x_2372 = v_2830 | ~v_2829;
assign x_2373 = v_75 | v_74 | v_106 | v_105 | v_104 | v_132 | v_113 | v_112 | v_121 | ~v_2762 | ~v_236 | ~v_235 | ~v_2789 | ~v_2788 | ~v_2787 | ~v_2786 | ~v_364 | ~v_363 | ~v_2759 | ~v_2756 | ~v_2755 | ~v_362 | ~v_2754 | ~v_361 | ~v_2753 | ~v_360 | ~v_359 | v_2829;
assign x_2374 = v_50 | v_49 | v_101 | v_100 | v_102 | v_111 | v_110 | v_131 | ~v_2750 | v_120 | ~v_217 | ~v_216 | ~v_2780 | ~v_2779 | ~v_2778 | ~v_2777 | ~v_353 | ~v_352 | ~v_2748 | ~v_2745 | ~v_2744 | ~v_351 | ~v_2743 | ~v_350 | ~v_2742 | ~v_349 | ~v_348 | v_2828;
assign x_2375 = v_24 | v_23 | ~v_2740 | v_95 | v_94 | v_93 | v_108 | v_109 | v_128 | v_117 | ~v_201 | ~v_200 | ~v_2772 | ~v_2771 | ~v_2770 | ~v_2769 | ~v_342 | ~v_341 | ~v_2736 | ~v_2734 | ~v_2733 | ~v_340 | ~v_2732 | ~v_339 | ~v_2731 | ~v_338 | ~v_337 | v_2827;
assign x_2376 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2825 | ~v_2809 | v_2826;
assign x_2377 = v_2825 | ~v_2814;
assign x_2378 = v_2825 | ~v_2819;
assign x_2379 = v_2825 | ~v_2824;
assign x_2380 = v_76 | v_74 | v_73 | v_107 | v_106 | v_105 | v_104 | v_113 | v_112 | ~v_2762 | ~v_2823 | ~v_2759 | ~v_2756 | ~v_2822 | ~v_2821 | ~v_2820 | ~v_454 | ~v_453 | ~v_480 | ~v_479 | ~v_478 | ~v_477 | ~v_2755 | ~v_362 | ~v_2754 | ~v_361 | ~v_2753 | v_2824;
assign x_2381 = v_2823 | ~v_98;
assign x_2382 = v_2823 | v_80;
assign x_2383 = v_2822 | v_88;
assign x_2384 = v_2822 | v_98;
assign x_2385 = v_2821 | v_97;
assign x_2386 = v_2821 | v_86;
assign x_2387 = v_2820 | ~v_97;
assign x_2388 = v_2820 | v_78;
assign x_2389 = v_51 | v_49 | v_48 | v_103 | v_101 | v_100 | v_102 | v_111 | v_110 | ~v_2750 | ~v_449 | ~v_2818 | ~v_2817 | ~v_447 | ~v_2816 | ~v_2815 | ~v_475 | ~v_474 | ~v_2748 | ~v_2745 | ~v_473 | ~v_472 | ~v_2744 | ~v_351 | ~v_2743 | ~v_350 | ~v_2742 | v_2819;
assign x_2390 = v_2818 | ~v_98;
assign x_2391 = v_2818 | v_55;
assign x_2392 = v_2817 | v_98;
assign x_2393 = v_2817 | v_63;
assign x_2394 = v_2816 | ~v_97;
assign x_2395 = v_2816 | v_53;
assign x_2396 = v_2815 | v_97;
assign x_2397 = v_2815 | v_61;
assign x_2398 = v_25 | v_23 | v_22 | ~v_2740 | ~v_2813 | v_96 | v_95 | v_94 | v_93 | v_108 | v_109 | ~v_470 | ~v_437 | ~v_2812 | ~v_469 | ~v_2736 | ~v_2811 | ~v_2810 | ~v_432 | ~v_468 | ~v_467 | ~v_2734 | ~v_2733 | ~v_340 | ~v_2732 | ~v_339 | ~v_2731 | v_2814;
assign x_2399 = v_2813 | ~v_98;
assign x_2400 = v_2813 | v_30;
assign x_2401 = v_2812 | v_97;
assign x_2402 = v_2812 | v_36;
assign x_2403 = v_2811 | v_98;
assign x_2404 = v_2811 | v_38;
assign x_2405 = v_2810 | ~v_97;
assign x_2406 = v_2810 | v_28;
assign x_2407 = v_2809 | ~v_2798;
assign x_2408 = v_2809 | ~v_2803;
assign x_2409 = v_2809 | ~v_2808;
assign x_2410 = v_76 | v_75 | v_74 | v_106 | v_105 | v_104 | v_132 | v_113 | v_112 | ~v_2807 | ~v_236 | ~v_235 | ~v_2789 | ~v_2788 | ~v_2787 | ~v_2786 | ~v_234 | ~v_233 | ~v_2806 | ~v_2805 | ~v_2759 | ~v_2756 | ~v_2804 | ~v_230 | ~v_229 | ~v_228 | ~v_227 | v_2808;
assign x_2411 = v_2807 | ~v_97;
assign x_2412 = v_2807 | v_79;
assign x_2413 = v_2806 | v_90;
assign x_2414 = v_2806 | v_98;
assign x_2415 = v_2805 | ~v_98;
assign x_2416 = v_2805 | v_82;
assign x_2417 = v_2804 | v_97;
assign x_2418 = v_2804 | v_87;
assign x_2419 = v_50 | v_51 | v_49 | v_101 | v_100 | ~v_2802 | v_102 | v_111 | v_110 | v_131 | ~v_225 | ~v_224 | ~v_2801 | ~v_2800 | ~v_2799 | ~v_217 | ~v_216 | ~v_215 | ~v_214 | ~v_2780 | ~v_2779 | ~v_2778 | ~v_2777 | ~v_213 | ~v_212 | ~v_2748 | ~v_2745 | v_2803;
assign x_2420 = v_2802 | ~v_98;
assign x_2421 = v_2802 | v_57;
assign x_2422 = v_2801 | v_98;
assign x_2423 = v_2801 | v_65;
assign x_2424 = v_2800 | ~v_97;
assign x_2425 = v_2800 | v_54;
assign x_2426 = v_2799 | v_97;
assign x_2427 = v_2799 | v_62;
assign x_2428 = v_25 | v_24 | v_23 | ~v_2740 | v_95 | v_94 | v_93 | v_108 | v_109 | v_128 | ~v_2797 | ~v_2796 | ~v_208 | ~v_201 | ~v_200 | ~v_199 | ~v_198 | ~v_2772 | ~v_2771 | ~v_2770 | ~v_2769 | ~v_197 | ~v_196 | ~v_2736 | ~v_2795 | ~v_2794 | ~v_193 | v_2798;
assign x_2429 = v_2797 | ~v_98;
assign x_2430 = v_2797 | v_32;
assign x_2431 = v_2796 | v_98;
assign x_2432 = v_2796 | v_40;
assign x_2433 = v_2795 | v_97;
assign x_2434 = v_2795 | v_37;
assign x_2435 = v_2794 | ~v_97;
assign x_2436 = v_2794 | v_29;
assign x_2437 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2792 | ~v_2764 | v_2793;
assign x_2438 = v_2792 | ~v_2773;
assign x_2439 = v_2792 | ~v_2782;
assign x_2440 = v_2792 | ~v_2791;
assign x_2441 = v_76 | v_75 | v_74 | v_72 | v_70 | v_104 | v_132 | v_113 | v_112 | ~v_2790 | ~v_236 | ~v_235 | ~v_2789 | ~v_2788 | ~v_2787 | ~v_2786 | ~v_311 | ~v_310 | ~v_2759 | ~v_2756 | ~v_2785 | ~v_2784 | ~v_2783 | ~v_421 | ~v_420 | ~v_419 | ~v_418 | v_2791;
assign x_2442 = v_2790 | v_87;
assign x_2443 = v_2790 | v_26;
assign x_2444 = v_2789 | v_124;
assign x_2445 = v_2789 | v_88;
assign x_2446 = v_2788 | ~v_124;
assign x_2447 = v_2788 | v_80;
assign x_2448 = v_2787 | v_123;
assign x_2449 = v_2787 | v_86;
assign x_2450 = v_2786 | ~v_123;
assign x_2451 = v_2786 | v_78;
assign x_2452 = v_2785 | v_90;
assign x_2453 = v_2785 | v_26;
assign x_2454 = v_2784 | v_82;
assign x_2455 = v_2784 | ~v_26;
assign x_2456 = v_2783 | v_79;
assign x_2457 = v_2783 | ~v_26;
assign x_2458 = v_50 | v_51 | v_49 | v_45 | v_47 | v_100 | v_111 | v_110 | v_131 | ~v_304 | ~v_2781 | ~v_416 | ~v_217 | ~v_216 | ~v_415 | ~v_2780 | ~v_2779 | ~v_2778 | ~v_2777 | ~v_2776 | ~v_2748 | ~v_297 | ~v_2745 | ~v_2775 | ~v_2774 | ~v_414 | ~v_413 | v_2782;
assign x_2459 = v_2781 | v_62;
assign x_2460 = v_2781 | v_26;
assign x_2461 = v_2780 | v_124;
assign x_2462 = v_2780 | v_63;
assign x_2463 = v_2779 | ~v_124;
assign x_2464 = v_2779 | v_55;
assign x_2465 = v_2778 | v_123;
assign x_2466 = v_2778 | v_61;
assign x_2467 = v_2777 | ~v_123;
assign x_2468 = v_2777 | v_53;
assign x_2469 = v_2776 | v_54;
assign x_2470 = v_2776 | ~v_26;
assign x_2471 = v_2775 | v_65;
assign x_2472 = v_2775 | v_26;
assign x_2473 = v_2774 | v_57;
assign x_2474 = v_2774 | ~v_26;
assign x_2475 = v_25 | v_24 | v_23 | v_21 | v_19 | ~v_2740 | v_93 | v_108 | v_109 | v_128 | ~v_293 | ~v_411 | ~v_410 | ~v_201 | ~v_200 | ~v_2772 | ~v_2771 | ~v_2770 | ~v_2769 | ~v_2768 | ~v_286 | ~v_2736 | ~v_2767 | ~v_2766 | ~v_2765 | ~v_409 | ~v_408 | v_2773;
assign x_2476 = v_2772 | v_124;
assign x_2477 = v_2772 | v_38;
assign x_2478 = v_2771 | ~v_124;
assign x_2479 = v_2771 | v_30;
assign x_2480 = v_2770 | v_123;
assign x_2481 = v_2770 | v_36;
assign x_2482 = v_2769 | ~v_123;
assign x_2483 = v_2769 | v_28;
assign x_2484 = v_2768 | v_40;
assign x_2485 = v_2768 | v_26;
assign x_2486 = v_2767 | v_37;
assign x_2487 = v_2767 | v_26;
assign x_2488 = v_2766 | v_32;
assign x_2489 = v_2766 | ~v_26;
assign x_2490 = v_2765 | v_29;
assign x_2491 = v_2765 | ~v_26;
assign x_2492 = v_2764 | ~v_2741;
assign x_2493 = v_2764 | ~v_2752;
assign x_2494 = v_2764 | ~v_2763;
assign x_2495 = v_76 | v_68 | v_75 | v_74 | v_73 | v_71 | v_106 | v_105 | v_104 | ~v_2762 | ~v_2761 | ~v_278 | ~v_2760 | ~v_273 | ~v_2759 | ~v_2758 | ~v_2757 | ~v_2756 | ~v_385 | ~v_384 | ~v_2755 | ~v_362 | ~v_2754 | ~v_361 | ~v_2753 | ~v_383 | ~v_382 | v_2763;
assign x_2496 = v_2762 | v_114;
assign x_2497 = v_2762 | v_87;
assign x_2498 = v_2761 | v_88;
assign x_2499 = v_2761 | v_26;
assign x_2500 = v_2760 | v_86;
assign x_2501 = v_2760 | v_26;
assign x_2502 = v_2759 | v_85;
assign x_2503 = v_2759 | v_26;
assign x_2504 = v_2758 | v_80;
assign x_2505 = v_2758 | ~v_26;
assign x_2506 = v_2757 | v_78;
assign x_2507 = v_2757 | ~v_26;
assign x_2508 = v_2756 | v_77;
assign x_2509 = v_2756 | ~v_26;
assign x_2510 = v_2755 | ~v_114;
assign x_2511 = v_2755 | v_79;
assign x_2512 = v_2754 | v_115;
assign x_2513 = v_2754 | v_90;
assign x_2514 = v_2753 | ~v_115;
assign x_2515 = v_2753 | v_82;
assign x_2516 = v_50 | v_51 | v_49 | v_48 | v_46 | v_43 | ~v_2751 | v_101 | v_100 | v_102 | ~v_2750 | ~v_268 | ~v_380 | ~v_379 | ~v_2749 | ~v_2748 | ~v_261 | ~v_2747 | ~v_2746 | ~v_2745 | ~v_2744 | ~v_351 | ~v_2743 | ~v_350 | ~v_2742 | ~v_378 | ~v_377 | v_2752;
assign x_2517 = v_2751 | v_61;
assign x_2518 = v_2751 | v_26;
assign x_2519 = v_2750 | v_114;
assign x_2520 = v_2750 | v_62;
assign x_2521 = v_2749 | v_63;
assign x_2522 = v_2749 | v_26;
assign x_2523 = v_2748 | v_60;
assign x_2524 = v_2748 | v_26;
assign x_2525 = v_2747 | v_55;
assign x_2526 = v_2747 | ~v_26;
assign x_2527 = v_2746 | v_53;
assign x_2528 = v_2746 | ~v_26;
assign x_2529 = v_2745 | v_52;
assign x_2530 = v_2745 | ~v_26;
assign x_2531 = v_2744 | ~v_114;
assign x_2532 = v_2744 | v_54;
assign x_2533 = v_2743 | v_115;
assign x_2534 = v_2743 | v_65;
assign x_2535 = v_2742 | ~v_115;
assign x_2536 = v_2742 | v_57;
assign x_2537 = v_25 | v_24 | v_23 | v_22 | v_20 | v_17 | ~v_2740 | v_95 | v_94 | v_93 | ~v_375 | ~v_374 | ~v_2739 | ~v_253 | ~v_252 | ~v_2738 | ~v_2737 | ~v_2736 | ~v_2735 | ~v_2734 | ~v_2733 | ~v_340 | ~v_2732 | ~v_339 | ~v_2731 | ~v_373 | ~v_372 | v_2741;
assign x_2538 = v_2740 | v_27;
assign x_2539 = v_2740 | ~v_26;
assign x_2540 = v_2739 | v_28;
assign x_2541 = v_2739 | ~v_26;
assign x_2542 = v_2738 | v_38;
assign x_2543 = v_2738 | v_26;
assign x_2544 = v_2737 | v_36;
assign x_2545 = v_2737 | v_26;
assign x_2546 = v_2736 | v_35;
assign x_2547 = v_2736 | v_26;
assign x_2548 = v_2735 | v_30;
assign x_2549 = v_2735 | ~v_26;
assign x_2550 = v_2734 | v_114;
assign x_2551 = v_2734 | v_37;
assign x_2552 = v_2733 | ~v_114;
assign x_2553 = v_2733 | v_29;
assign x_2554 = v_2732 | v_115;
assign x_2555 = v_2732 | v_40;
assign x_2556 = v_2731 | ~v_115;
assign x_2557 = v_2731 | v_32;
assign x_2558 = v_2730 | ~v_2486;
assign x_2559 = v_2730 | ~v_2535;
assign x_2560 = v_2730 | ~v_2560;
assign x_2561 = v_2730 | ~v_2571;
assign x_2562 = v_2730 | ~v_2606;
assign x_2563 = v_2730 | ~v_2625;
assign x_2564 = v_2730 | ~v_2634;
assign x_2565 = v_2730 | ~v_2643;
assign x_2566 = v_2730 | ~v_2652;
assign x_2567 = v_2730 | ~v_2661;
assign x_2568 = v_2730 | ~v_2670;
assign x_2569 = v_2730 | ~v_2687;
assign x_2570 = v_2730 | ~v_2696;
assign x_2571 = v_2730 | ~v_2705;
assign x_2572 = v_2730 | ~v_2714;
assign x_2573 = v_2730 | ~v_2729;
assign x_2574 = v_9 | v_7 | v_5 | v_4 | v_6 | v_3 | v_2 | v_1 | ~v_1041 | ~v_1040 | ~v_2728 | v_2729;
assign x_2575 = v_2728 | ~v_2721;
assign x_2576 = v_2728 | ~v_2727;
assign x_2577 = v_99 | ~v_2483 | ~v_1022 | ~v_1811 | ~v_2603 | ~v_2622 | ~v_2684 | ~v_2726 | v_2727;
assign x_2578 = v_2726 | ~v_2725;
assign x_2579 = v_2726 | ~v_698;
assign x_2580 = v_2726 | ~v_699;
assign x_2581 = v_2726 | ~v_700;
assign x_2582 = v_2726 | ~v_701;
assign x_2583 = ~v_2724 | ~v_2723 | ~v_2722 | v_2725;
assign x_2584 = v_2724 | ~v_1372;
assign x_2585 = v_2724 | ~v_2301;
assign x_2586 = v_2724 | ~v_2302;
assign x_2587 = v_2724 | ~v_763;
assign x_2588 = v_2724 | ~v_764;
assign x_2589 = v_2724 | ~v_2329;
assign x_2590 = v_2724 | ~v_2330;
assign x_2591 = v_2724 | ~v_726;
assign x_2592 = v_2724 | ~v_2303;
assign x_2593 = v_2724 | ~v_2304;
assign x_2594 = v_2724 | ~v_1373;
assign x_2595 = v_2724 | ~v_2305;
assign x_2596 = v_2724 | ~v_2333;
assign x_2597 = v_2724 | ~v_731;
assign x_2598 = v_2724 | ~v_1374;
assign x_2599 = v_2724 | ~v_2307;
assign x_2600 = v_2724 | ~v_2336;
assign x_2601 = v_2724 | ~v_1375;
assign x_2602 = v_2724 | ~v_112;
assign x_2603 = v_2724 | ~v_105;
assign x_2604 = v_2724 | ~v_76;
assign x_2605 = v_2724 | ~v_75;
assign x_2606 = v_2724 | ~v_74;
assign x_2607 = v_2724 | ~v_73;
assign x_2608 = v_2724 | ~v_72;
assign x_2609 = v_2724 | ~v_71;
assign x_2610 = v_2724 | ~v_69;
assign x_2611 = v_2723 | ~v_1367;
assign x_2612 = v_2723 | ~v_1368;
assign x_2613 = v_2723 | ~v_2290;
assign x_2614 = v_2723 | ~v_2291;
assign x_2615 = v_2723 | ~v_750;
assign x_2616 = v_2723 | ~v_714;
assign x_2617 = v_2723 | ~v_2322;
assign x_2618 = v_2723 | ~v_2292;
assign x_2619 = v_2723 | ~v_2323;
assign x_2620 = v_2723 | ~v_2293;
assign x_2621 = v_2723 | ~v_757;
assign x_2622 = v_2723 | ~v_1369;
assign x_2623 = v_2723 | ~v_721;
assign x_2624 = v_2723 | ~v_2295;
assign x_2625 = v_2723 | ~v_2326;
assign x_2626 = v_2723 | ~v_2327;
assign x_2627 = v_2723 | ~v_2296;
assign x_2628 = v_2723 | ~v_110;
assign x_2629 = v_2723 | ~v_101;
assign x_2630 = v_2723 | ~v_1370;
assign x_2631 = v_2723 | ~v_51;
assign x_2632 = v_2723 | ~v_50;
assign x_2633 = v_2723 | ~v_49;
assign x_2634 = v_2723 | ~v_48;
assign x_2635 = v_2723 | ~v_47;
assign x_2636 = v_2723 | ~v_46;
assign x_2637 = v_2723 | ~v_44;
assign x_2638 = v_2722 | ~v_1362;
assign x_2639 = v_2722 | ~v_2279;
assign x_2640 = v_2722 | ~v_739;
assign x_2641 = v_2722 | ~v_2311;
assign x_2642 = v_2722 | ~v_2280;
assign x_2643 = v_2722 | ~v_2281;
assign x_2644 = v_2722 | ~v_705;
assign x_2645 = v_2722 | ~v_706;
assign x_2646 = v_2722 | ~v_1363;
assign x_2647 = v_2722 | ~v_2282;
assign x_2648 = v_2722 | ~v_2283;
assign x_2649 = v_2722 | ~v_746;
assign x_2650 = v_2722 | ~v_1364;
assign x_2651 = v_2722 | ~v_2316;
assign x_2652 = v_2722 | ~v_2317;
assign x_2653 = v_2722 | ~v_1365;
assign x_2654 = v_2722 | ~v_2286;
assign x_2655 = v_2722 | ~v_2318;
assign x_2656 = v_2722 | ~v_108;
assign x_2657 = v_2722 | ~v_94;
assign x_2658 = v_2722 | ~v_25;
assign x_2659 = v_2722 | ~v_24;
assign x_2660 = v_2722 | ~v_23;
assign x_2661 = v_2722 | ~v_22;
assign x_2662 = v_2722 | ~v_21;
assign x_2663 = v_2722 | ~v_20;
assign x_2664 = v_2722 | ~v_18;
assign x_2665 = ~v_2275 | ~v_2720 | v_2721;
assign x_2666 = v_2720 | ~v_2719;
assign x_2667 = v_2720 | ~v_2676;
assign x_2668 = v_2720 | ~v_2613;
assign x_2669 = v_2720 | ~v_2586;
assign x_2670 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2718 | v_2719;
assign x_2671 = v_2718 | ~v_2715;
assign x_2672 = v_2718 | ~v_2716;
assign x_2673 = v_2718 | ~v_2717;
assign x_2674 = v_76 | v_69 | v_75 | v_74 | v_73 | v_72 | v_71 | v_105 | ~v_1356 | v_112 | ~v_2126 | ~v_2097 | ~v_1355 | ~v_278 | ~v_2123 | ~v_2095 | ~v_1354 | ~v_2094 | ~v_2093 | ~v_273 | ~v_2120 | ~v_2119 | ~v_311 | ~v_310 | ~v_2092 | ~v_2091 | ~v_1353 | v_2717;
assign x_2675 = v_50 | v_51 | v_49 | v_48 | v_46 | v_47 | v_44 | ~v_1351 | v_101 | v_110 | ~v_2086 | ~v_2117 | ~v_2116 | ~v_2085 | ~v_268 | ~v_1350 | ~v_304 | ~v_2083 | ~v_2113 | ~v_2082 | ~v_2112 | ~v_261 | ~v_297 | ~v_2081 | ~v_2080 | ~v_1349 | ~v_1348 | v_2716;
assign x_2676 = v_25 | v_24 | v_23 | v_22 | v_21 | v_20 | v_18 | ~v_2108 | v_94 | ~v_2076 | v_108 | ~v_1346 | ~v_2107 | ~v_2106 | ~v_1345 | ~v_293 | ~v_2073 | ~v_2072 | ~v_1344 | ~v_253 | ~v_252 | ~v_2071 | ~v_2070 | ~v_2101 | ~v_286 | ~v_2069 | ~v_1343 | v_2715;
assign x_2677 = v_7 | v_5 | v_4 | v_10 | v_3 | v_2 | v_1 | ~v_1041 | ~v_1040 | ~v_2713 | v_2714;
assign x_2678 = v_2713 | ~v_2709;
assign x_2679 = v_2713 | ~v_2712;
assign x_2680 = v_99 | ~v_2483 | ~v_1022 | ~v_1811 | ~v_2453 | ~v_2452 | ~v_2451 | ~v_2450 | ~v_2445 | ~v_2711 | ~v_2710 | v_2712;
assign x_2681 = v_2711 | ~v_2548;
assign x_2682 = v_2711 | ~v_2473;
assign x_2683 = v_2710 | ~v_2529;
assign x_2684 = v_2710 | ~v_2566;
assign x_2685 = ~v_2275 | ~v_2708 | v_2709;
assign x_2686 = v_2708 | ~v_2706;
assign x_2687 = v_2708 | ~v_2707;
assign x_2688 = v_2708 | ~v_2235;
assign x_2689 = v_2708 | ~v_2240;
assign x_2690 = v_2708 | ~v_2241;
assign x_2691 = v_2708 | ~v_2242;
assign x_2692 = v_2708 | ~v_2243;
assign x_2693 = ~v_2263 | ~v_2536 | v_2707;
assign x_2694 = ~v_2561 | ~v_2505 | v_2706;
assign x_2695 = v_9 | v_7 | v_5 | v_6 | v_10 | v_3 | v_2 | v_1 | ~v_1041 | ~v_1040 | ~v_2704 | v_2705;
assign x_2696 = v_2704 | ~v_2700;
assign x_2697 = v_2704 | ~v_2703;
assign x_2698 = v_99 | ~v_2483 | ~v_1022 | ~v_1811 | ~v_2472 | ~v_2471 | ~v_2466 | ~v_2461 | ~v_2460 | ~v_2702 | ~v_2701 | v_2703;
assign x_2699 = v_2702 | ~v_2597;
assign x_2700 = v_2702 | ~v_2566;
assign x_2701 = v_2701 | ~v_2601;
assign x_2702 = v_2701 | ~v_2454;
assign x_2703 = ~v_2275 | ~v_2699 | v_2700;
assign x_2704 = v_2699 | ~v_2697;
assign x_2705 = v_2699 | ~v_2698;
assign x_2706 = v_2699 | ~v_2250;
assign x_2707 = v_2699 | ~v_2251;
assign x_2708 = v_2699 | ~v_2256;
assign x_2709 = v_2699 | ~v_2261;
assign x_2710 = v_2699 | ~v_2262;
assign x_2711 = ~v_2561 | ~v_2580 | v_2698;
assign x_2712 = ~v_2244 | ~v_2584 | v_2697;
assign x_2713 = v_9 | v_5 | v_6 | v_8 | v_10 | v_2 | v_1 | ~v_1041 | ~v_1040 | ~v_2695 | v_2696;
assign x_2714 = v_2695 | ~v_2691;
assign x_2715 = v_2695 | ~v_2694;
assign x_2716 = v_99 | ~v_2483 | ~v_1022 | ~v_1811 | ~v_2469 | ~v_2468 | ~v_2467 | ~v_2600 | ~v_2599 | ~v_2693 | ~v_2692 | v_2694;
assign x_2717 = v_2693 | ~v_2416;
assign x_2718 = v_2693 | ~v_2597;
assign x_2719 = v_2692 | ~v_2552;
assign x_2720 = v_2692 | ~v_2473;
assign x_2721 = ~v_2275 | ~v_2690 | v_2691;
assign x_2722 = v_2690 | ~v_2688;
assign x_2723 = v_2690 | ~v_2689;
assign x_2724 = v_2690 | ~v_2582;
assign x_2725 = v_2690 | ~v_2583;
assign x_2726 = v_2690 | ~v_2257;
assign x_2727 = v_2690 | ~v_2258;
assign x_2728 = v_2690 | ~v_2259;
assign x_2729 = ~v_2580 | ~v_2206 | v_2689;
assign x_2730 = ~v_2263 | ~v_2540 | v_2688;
assign x_2731 = v_5 | v_4 | v_8 | v_10 | v_2 | v_1 | ~v_1041 | ~v_1040 | ~v_2686 | v_2687;
assign x_2732 = v_2686 | ~v_2678;
assign x_2733 = v_2686 | ~v_2685;
assign x_2734 = v_99 | ~v_2483 | ~v_1022 | ~v_1811 | ~v_2684 | ~v_2602 | ~v_2621 | ~v_2683 | v_2685;
assign x_2735 = v_2684 | ~v_2454;
assign x_2736 = v_2684 | ~v_2552;
assign x_2737 = v_2683 | ~v_2682;
assign x_2738 = v_2683 | ~v_698;
assign x_2739 = v_2683 | ~v_699;
assign x_2740 = v_2683 | ~v_700;
assign x_2741 = v_2683 | ~v_701;
assign x_2742 = ~v_2681 | ~v_2680 | ~v_2679 | v_2682;
assign x_2743 = v_2681 | ~v_682;
assign x_2744 = v_2681 | ~v_683;
assign x_2745 = v_2681 | ~v_906;
assign x_2746 = v_2681 | ~v_907;
assign x_2747 = v_2681 | ~v_2301;
assign x_2748 = v_2681 | ~v_2302;
assign x_2749 = v_2681 | ~v_2350;
assign x_2750 = v_2681 | ~v_2366;
assign x_2751 = v_2681 | ~v_2367;
assign x_2752 = v_2681 | ~v_2351;
assign x_2753 = v_2681 | ~v_2352;
assign x_2754 = v_2681 | ~v_1323;
assign x_2755 = v_2681 | ~v_1324;
assign x_2756 = v_2681 | ~v_1325;
assign x_2757 = v_2681 | ~v_2368;
assign x_2758 = v_2681 | ~v_2353;
assign x_2759 = v_2681 | ~v_1326;
assign x_2760 = v_2681 | ~v_2369;
assign x_2761 = v_2681 | ~v_113;
assign x_2762 = v_2681 | ~v_106;
assign x_2763 = v_2681 | ~v_76;
assign x_2764 = v_2681 | ~v_75;
assign x_2765 = v_2681 | ~v_74;
assign x_2766 = v_2681 | ~v_73;
assign x_2767 = v_2681 | ~v_70;
assign x_2768 = v_2681 | ~v_69;
assign x_2769 = v_2681 | ~v_68;
assign x_2770 = v_2680 | ~v_2290;
assign x_2771 = v_2680 | ~v_2291;
assign x_2772 = v_2680 | ~v_1318;
assign x_2773 = v_2680 | ~v_2345;
assign x_2774 = v_2680 | ~v_2346;
assign x_2775 = v_2680 | ~v_2361;
assign x_2776 = v_2680 | ~v_1319;
assign x_2777 = v_2680 | ~v_2362;
assign x_2778 = v_2680 | ~v_900;
assign x_2779 = v_2680 | ~v_2347;
assign x_2780 = v_2680 | ~v_2348;
assign x_2781 = v_2680 | ~v_2363;
assign x_2782 = v_2680 | ~v_677;
assign x_2783 = v_2680 | ~v_2364;
assign x_2784 = v_2680 | ~v_902;
assign x_2785 = v_2680 | ~v_1320;
assign x_2786 = v_2680 | ~v_678;
assign x_2787 = v_2680 | ~v_1321;
assign x_2788 = v_2680 | ~v_111;
assign x_2789 = v_2680 | ~v_102;
assign x_2790 = v_2680 | ~v_51;
assign x_2791 = v_2680 | ~v_50;
assign x_2792 = v_2680 | ~v_49;
assign x_2793 = v_2680 | ~v_48;
assign x_2794 = v_2680 | ~v_45;
assign x_2795 = v_2680 | ~v_44;
assign x_2796 = v_2680 | ~v_43;
assign x_2797 = v_2679 | ~v_646;
assign x_2798 = v_2679 | ~v_885;
assign x_2799 = v_2679 | ~v_2279;
assign x_2800 = v_2679 | ~v_2340;
assign x_2801 = v_2679 | ~v_2341;
assign x_2802 = v_2679 | ~v_2356;
assign x_2803 = v_2679 | ~v_2357;
assign x_2804 = v_2679 | ~v_2358;
assign x_2805 = v_2679 | ~v_1313;
assign x_2806 = v_2679 | ~v_1314;
assign x_2807 = v_2679 | ~v_2359;
assign x_2808 = v_2679 | ~v_2282;
assign x_2809 = v_2679 | ~v_1315;
assign x_2810 = v_2679 | ~v_661;
assign x_2811 = v_2679 | ~v_890;
assign x_2812 = v_2679 | ~v_2342;
assign x_2813 = v_2679 | ~v_2343;
assign x_2814 = v_2679 | ~v_1316;
assign x_2815 = v_2679 | ~v_109;
assign x_2816 = v_2679 | ~v_95;
assign x_2817 = v_2679 | ~v_25;
assign x_2818 = v_2679 | ~v_24;
assign x_2819 = v_2679 | ~v_23;
assign x_2820 = v_2679 | ~v_22;
assign x_2821 = v_2679 | ~v_19;
assign x_2822 = v_2679 | ~v_18;
assign x_2823 = v_2679 | ~v_17;
assign x_2824 = ~v_2275 | ~v_2677 | v_2678;
assign x_2825 = v_2677 | ~v_2675;
assign x_2826 = v_2677 | ~v_2612;
assign x_2827 = v_2677 | ~v_2585;
assign x_2828 = v_2677 | ~v_2676;
assign x_2829 = ~v_2540 | ~v_2244 | v_2676;
assign x_2830 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2674 | v_2675;
assign x_2831 = v_2674 | ~v_2671;
assign x_2832 = v_2674 | ~v_2672;
assign x_2833 = v_2674 | ~v_2673;
assign x_2834 = v_76 | v_69 | v_68 | v_75 | v_74 | v_73 | v_70 | v_106 | v_113 | ~v_2159 | ~v_1306 | ~v_2143 | ~v_2158 | ~v_1305 | ~v_1304 | ~v_1303 | ~v_2142 | ~v_2141 | ~v_2157 | ~v_2156 | ~v_2140 | ~v_2092 | ~v_2091 | ~v_454 | ~v_453 | ~v_230 | ~v_229 | v_2673;
assign x_2835 = v_50 | v_51 | v_49 | v_48 | v_45 | v_43 | v_44 | v_102 | v_111 | ~v_1301 | ~v_225 | ~v_1300 | ~v_449 | ~v_2154 | ~v_224 | ~v_2153 | ~v_2138 | ~v_2137 | ~v_447 | ~v_2152 | ~v_1299 | ~v_2151 | ~v_2136 | ~v_2135 | ~v_1298 | ~v_2081 | ~v_2080 | v_2672;
assign x_2836 = v_25 | v_24 | v_23 | v_22 | v_19 | v_18 | v_17 | v_95 | v_109 | ~v_1296 | ~v_2133 | ~v_2132 | ~v_437 | ~v_208 | ~v_1295 | ~v_2073 | ~v_2149 | ~v_1294 | ~v_1293 | ~v_2148 | ~v_2147 | ~v_2146 | ~v_2131 | ~v_2130 | ~v_2069 | ~v_432 | ~v_193 | v_2671;
assign x_2837 = v_9 | v_5 | v_4 | v_6 | v_8 | v_2 | v_1 | ~v_1041 | ~v_1040 | ~v_2669 | v_2670;
assign x_2838 = v_2669 | ~v_2665;
assign x_2839 = v_2669 | ~v_2668;
assign x_2840 = v_99 | ~v_2483 | ~v_1022 | ~v_1811 | ~v_2520 | ~v_2519 | ~v_2518 | ~v_2551 | ~v_2549 | ~v_2667 | ~v_2666 | v_2668;
assign x_2841 = v_2667 | ~v_2601;
assign x_2842 = v_2667 | ~v_2524;
assign x_2843 = v_2666 | ~v_2416;
assign x_2844 = v_2666 | ~v_2556;
assign x_2845 = ~v_2275 | ~v_2664 | v_2665;
assign x_2846 = v_2664 | ~v_2662;
assign x_2847 = v_2664 | ~v_2663;
assign x_2848 = v_2664 | ~v_2537;
assign x_2849 = v_2664 | ~v_2539;
assign x_2850 = v_2664 | ~v_2494;
assign x_2851 = v_2664 | ~v_2495;
assign x_2852 = v_2664 | ~v_2496;
assign x_2853 = ~v_2500 | ~v_2584 | v_2663;
assign x_2854 = ~v_2544 | ~v_2206 | v_2662;
assign x_2855 = v_9 | v_4 | v_6 | v_8 | v_10 | v_2 | v_1 | ~v_1041 | ~v_1040 | ~v_2660 | v_2661;
assign x_2856 = v_2660 | ~v_2656;
assign x_2857 = v_2660 | ~v_2659;
assign x_2858 = v_99 | ~v_2483 | ~v_1022 | ~v_1811 | ~v_2415 | ~v_2414 | ~v_2413 | ~v_2412 | ~v_2395 | ~v_2658 | ~v_2657 | v_2659;
assign x_2859 = v_2658 | ~v_2459;
assign x_2860 = v_2658 | ~v_2601;
assign x_2861 = v_2657 | ~v_2552;
assign x_2862 = v_2657 | ~v_2566;
assign x_2863 = ~v_2275 | ~v_2655 | v_2656;
assign x_2864 = v_2655 | ~v_2653;
assign x_2865 = v_2655 | ~v_2654;
assign x_2866 = v_2655 | ~v_2185;
assign x_2867 = v_2655 | ~v_2202;
assign x_2868 = v_2655 | ~v_2203;
assign x_2869 = v_2655 | ~v_2204;
assign x_2870 = v_2655 | ~v_2205;
assign x_2871 = ~v_2584 | ~v_2249 | v_2654;
assign x_2872 = ~v_2561 | ~v_2540 | v_2653;
assign x_2873 = v_9 | v_7 | v_5 | v_6 | v_8 | v_10 | v_3 | v_1 | ~v_1041 | ~v_1040 | ~v_2651 | v_2652;
assign x_2874 = v_2651 | ~v_2647;
assign x_2875 = v_2651 | ~v_2650;
assign x_2876 = v_99 | ~v_2483 | ~v_1022 | ~v_1811 | ~v_2464 | ~v_2463 | ~v_2462 | ~v_2596 | ~v_2595 | ~v_2649 | ~v_2648 | v_2650;
assign x_2877 = v_2649 | ~v_2601;
assign x_2878 = v_2649 | ~v_2529;
assign x_2879 = v_2648 | ~v_2556;
assign x_2880 = v_2648 | ~v_2473;
assign x_2881 = ~v_2275 | ~v_2646 | v_2647;
assign x_2882 = v_2646 | ~v_2644;
assign x_2883 = v_2646 | ~v_2645;
assign x_2884 = v_2646 | ~v_2578;
assign x_2885 = v_2646 | ~v_2579;
assign x_2886 = v_2646 | ~v_2252;
assign x_2887 = v_2646 | ~v_2253;
assign x_2888 = v_2646 | ~v_2254;
assign x_2889 = ~v_2505 | ~v_2584 | v_2645;
assign x_2890 = ~v_2263 | ~v_2544 | v_2644;
assign x_2891 = v_7 | v_5 | v_4 | v_8 | v_10 | v_3 | v_1 | ~v_1041 | ~v_1040 | ~v_2642 | v_2643;
assign x_2892 = v_2642 | ~v_2638;
assign x_2893 = v_2642 | ~v_2641;
assign x_2894 = v_99 | ~v_2483 | ~v_1022 | ~v_1811 | ~v_2443 | ~v_2438 | ~v_2433 | ~v_2528 | ~v_2526 | ~v_2640 | ~v_2639 | v_2641;
assign x_2895 = v_2640 | ~v_2597;
assign x_2896 = v_2640 | ~v_2548;
assign x_2897 = v_2639 | ~v_2454;
assign x_2898 = v_2639 | ~v_2556;
assign x_2899 = ~v_2275 | ~v_2637 | v_2638;
assign x_2900 = v_2637 | ~v_2635;
assign x_2901 = v_2637 | ~v_2636;
assign x_2902 = v_2637 | ~v_2502;
assign x_2903 = v_2637 | ~v_2504;
assign x_2904 = v_2637 | ~v_2223;
assign x_2905 = v_2637 | ~v_2228;
assign x_2906 = v_2637 | ~v_2233;
assign x_2907 = ~v_2536 | ~v_2580 | v_2636;
assign x_2908 = ~v_2544 | ~v_2244 | v_2635;
assign x_2909 = v_9 | v_7 | v_5 | v_4 | v_6 | v_8 | v_3 | v_1 | ~v_1041 | ~v_1040 | ~v_2633 | v_2634;
assign x_2910 = v_2633 | ~v_2629;
assign x_2911 = v_2633 | ~v_2632;
assign x_2912 = v_99 | ~v_2483 | ~v_1022 | ~v_1811 | ~v_2513 | ~v_2512 | ~v_2511 | ~v_2555 | ~v_2554 | ~v_2631 | ~v_2630 | v_2632;
assign x_2913 = v_2631 | ~v_2597;
assign x_2914 = v_2631 | ~v_2524;
assign x_2915 = v_2630 | ~v_2529;
assign x_2916 = v_2630 | ~v_2552;
assign x_2917 = ~v_2275 | ~v_2628 | v_2629;
assign x_2918 = v_2628 | ~v_2626;
assign x_2919 = v_2628 | ~v_2627;
assign x_2920 = v_2628 | ~v_2542;
assign x_2921 = v_2628 | ~v_2543;
assign x_2922 = v_2628 | ~v_2487;
assign x_2923 = v_2628 | ~v_2488;
assign x_2924 = v_2628 | ~v_2489;
assign x_2925 = ~v_2500 | ~v_2580 | v_2627;
assign x_2926 = ~v_2540 | ~v_2505 | v_2626;
assign x_2927 = v_9 | v_7 | v_4 | v_6 | v_8 | v_10 | v_3 | v_1 | ~v_1041 | ~v_1040 | ~v_2624 | v_2625;
assign x_2928 = v_2624 | ~v_2615;
assign x_2929 = v_2624 | ~v_2623;
assign x_2930 = v_99 | ~v_2483 | ~v_1022 | ~v_1811 | ~v_2622 | ~v_2621 | ~v_2598 | ~v_2620 | v_2623;
assign x_2931 = v_2622 | ~v_2566;
assign x_2932 = v_2622 | ~v_2556;
assign x_2933 = v_2621 | ~v_2416;
assign x_2934 = v_2621 | ~v_2529;
assign x_2935 = v_2620 | ~v_2619;
assign x_2936 = v_2620 | ~v_698;
assign x_2937 = v_2620 | ~v_699;
assign x_2938 = v_2620 | ~v_700;
assign x_2939 = v_2620 | ~v_701;
assign x_2940 = ~v_2618 | ~v_2617 | ~v_2616 | v_2619;
assign x_2941 = v_2618 | ~v_1218;
assign x_2942 = v_2618 | ~v_1219;
assign x_2943 = v_2618 | ~v_814;
assign x_2944 = v_2618 | ~v_815;
assign x_2945 = v_2618 | ~v_2299;
assign x_2946 = v_2618 | ~v_2300;
assign x_2947 = v_2618 | ~v_2427;
assign x_2948 = v_2618 | ~v_2428;
assign x_2949 = v_2618 | ~v_2301;
assign x_2950 = v_2618 | ~v_2302;
assign x_2951 = v_2618 | ~v_632;
assign x_2952 = v_2618 | ~v_633;
assign x_2953 = v_2618 | ~v_1220;
assign x_2954 = v_2618 | ~v_1221;
assign x_2955 = v_2618 | ~v_2429;
assign x_2956 = v_2618 | ~v_2430;
assign x_2957 = v_2618 | ~v_2306;
assign x_2958 = v_2618 | ~v_2308;
assign x_2959 = v_2618 | ~v_113;
assign x_2960 = v_2618 | ~v_112;
assign x_2961 = v_2618 | ~v_106;
assign x_2962 = v_2618 | ~v_105;
assign x_2963 = v_2618 | ~v_76;
assign x_2964 = v_2618 | ~v_75;
assign x_2965 = v_2618 | ~v_74;
assign x_2966 = v_2618 | ~v_73;
assign x_2967 = v_2618 | ~v_69;
assign x_2968 = v_2617 | ~v_1213;
assign x_2969 = v_2617 | ~v_1214;
assign x_2970 = v_2617 | ~v_803;
assign x_2971 = v_2617 | ~v_804;
assign x_2972 = v_2617 | ~v_2288;
assign x_2973 = v_2617 | ~v_2289;
assign x_2974 = v_2617 | ~v_2422;
assign x_2975 = v_2617 | ~v_2423;
assign x_2976 = v_2617 | ~v_2290;
assign x_2977 = v_2617 | ~v_2291;
assign x_2978 = v_2617 | ~v_613;
assign x_2979 = v_2617 | ~v_614;
assign x_2980 = v_2617 | ~v_1215;
assign x_2981 = v_2617 | ~v_1216;
assign x_2982 = v_2617 | ~v_2424;
assign x_2983 = v_2617 | ~v_2294;
assign x_2984 = v_2617 | ~v_2425;
assign x_2985 = v_2617 | ~v_2297;
assign x_2986 = v_2617 | ~v_111;
assign x_2987 = v_2617 | ~v_110;
assign x_2988 = v_2617 | ~v_102;
assign x_2989 = v_2617 | ~v_101;
assign x_2990 = v_2617 | ~v_51;
assign x_2991 = v_2617 | ~v_50;
assign x_2992 = v_2617 | ~v_49;
assign x_2993 = v_2617 | ~v_48;
assign x_2994 = v_2617 | ~v_44;
assign x_2995 = v_2616 | ~v_1208;
assign x_2996 = v_2616 | ~v_1209;
assign x_2997 = v_2616 | ~v_792;
assign x_2998 = v_2616 | ~v_793;
assign x_2999 = v_2616 | ~v_2277;
assign x_3000 = v_2616 | ~v_2278;
assign x_3001 = v_2616 | ~v_2417;
assign x_3002 = v_2616 | ~v_2418;
assign x_3003 = v_2616 | ~v_2279;
assign x_3004 = v_2616 | ~v_594;
assign x_3005 = v_2616 | ~v_595;
assign x_3006 = v_2616 | ~v_1210;
assign x_3007 = v_2616 | ~v_1211;
assign x_3008 = v_2616 | ~v_2282;
assign x_3009 = v_2616 | ~v_2419;
assign x_3010 = v_2616 | ~v_2420;
assign x_3011 = v_2616 | ~v_2284;
assign x_3012 = v_2616 | ~v_2285;
assign x_3013 = v_2616 | ~v_109;
assign x_3014 = v_2616 | ~v_108;
assign x_3015 = v_2616 | ~v_95;
assign x_3016 = v_2616 | ~v_94;
assign x_3017 = v_2616 | ~v_25;
assign x_3018 = v_2616 | ~v_24;
assign x_3019 = v_2616 | ~v_23;
assign x_3020 = v_2616 | ~v_22;
assign x_3021 = v_2616 | ~v_18;
assign x_3022 = ~v_2275 | ~v_2614 | v_2615;
assign x_3023 = v_2614 | ~v_2611;
assign x_3024 = v_2614 | ~v_2581;
assign x_3025 = v_2614 | ~v_2612;
assign x_3026 = v_2614 | ~v_2613;
assign x_3027 = ~v_2544 | ~v_2561 | v_2613;
assign x_3028 = ~v_2505 | ~v_2206 | v_2612;
assign x_3029 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2610 | v_2611;
assign x_3030 = v_2610 | ~v_2607;
assign x_3031 = v_2610 | ~v_2608;
assign x_3032 = v_2610 | ~v_2609;
assign x_3033 = v_76 | v_69 | v_75 | v_74 | v_73 | v_106 | v_105 | v_113 | v_112 | ~v_2098 | ~v_2096 | ~v_2220 | ~v_2219 | ~v_1200 | ~v_1199 | ~v_180 | ~v_179 | ~v_2092 | ~v_2091 | ~v_2218 | ~v_2217 | ~v_2090 | ~v_2089 | ~v_362 | ~v_361 | ~v_1198 | ~v_1197 | v_2609;
assign x_3034 = v_50 | v_51 | v_49 | v_48 | v_44 | v_101 | v_102 | v_111 | v_110 | ~v_2087 | ~v_2215 | ~v_2084 | ~v_2214 | ~v_1195 | ~v_1194 | ~v_161 | ~v_160 | ~v_2081 | ~v_2080 | ~v_2213 | ~v_2212 | ~v_2079 | ~v_2078 | ~v_351 | ~v_350 | ~v_1193 | ~v_1192 | v_2608;
assign x_3035 = v_25 | v_24 | v_23 | v_22 | v_18 | v_95 | v_94 | v_108 | v_109 | ~v_2075 | ~v_2074 | ~v_2210 | ~v_2209 | ~v_2073 | ~v_1190 | ~v_1189 | ~v_142 | ~v_141 | ~v_2069 | ~v_2208 | ~v_2207 | ~v_2068 | ~v_2067 | ~v_340 | ~v_339 | ~v_1188 | ~v_1187 | v_2607;
assign x_3036 = v_9 | v_7 | v_5 | v_6 | v_8 | v_10 | v_3 | v_2 | ~v_1041 | ~v_1040 | ~v_2605 | v_2606;
assign x_3037 = v_2605 | ~v_2588;
assign x_3038 = v_2605 | ~v_2604;
assign x_3039 = v_99 | ~v_2483 | ~v_1022 | ~v_1811 | ~v_2603 | ~v_2602 | ~v_2598 | ~v_2593 | v_2604;
assign x_3040 = v_2603 | ~v_2473;
assign x_3041 = v_2603 | ~v_2524;
assign x_3042 = v_2602 | ~v_2601;
assign x_3043 = v_2602 | ~v_2548;
assign x_3044 = ~v_2469 | ~v_2468 | ~v_2467 | ~v_2600 | ~v_2599 | v_2601;
assign x_3045 = v_2600 | ~v_2465;
assign x_3046 = v_2600 | ~v_2371;
assign x_3047 = v_2600 | ~v_698;
assign x_3048 = v_2600 | ~v_699;
assign x_3049 = v_2600 | ~v_700;
assign x_3050 = v_2600 | ~v_701;
assign x_3051 = v_2599 | ~v_2594;
assign x_3052 = v_2599 | ~v_2411;
assign x_3053 = v_2599 | ~v_698;
assign x_3054 = v_2599 | ~v_699;
assign x_3055 = v_2599 | ~v_700;
assign x_3056 = v_2599 | ~v_701;
assign x_3057 = v_2598 | ~v_2459;
assign x_3058 = v_2598 | ~v_2597;
assign x_3059 = ~v_2464 | ~v_2463 | ~v_2462 | ~v_2596 | ~v_2595 | v_2597;
assign x_3060 = v_2596 | ~v_2470;
assign x_3061 = v_2596 | ~v_2442;
assign x_3062 = v_2596 | ~v_698;
assign x_3063 = v_2596 | ~v_699;
assign x_3064 = v_2596 | ~v_700;
assign x_3065 = v_2596 | ~v_701;
assign x_3066 = v_2595 | ~v_2594;
assign x_3067 = v_2595 | ~v_2437;
assign x_3068 = v_2595 | ~v_698;
assign x_3069 = v_2595 | ~v_699;
assign x_3070 = v_2595 | ~v_700;
assign x_3071 = v_2595 | ~v_701;
assign x_3072 = ~v_2472 | ~v_2461 | ~v_2460 | v_2594;
assign x_3073 = v_2593 | ~v_2592;
assign x_3074 = v_2593 | ~v_698;
assign x_3075 = v_2593 | ~v_699;
assign x_3076 = v_2593 | ~v_700;
assign x_3077 = v_2593 | ~v_701;
assign x_3078 = ~v_2591 | ~v_2590 | ~v_2589 | v_2592;
assign x_3079 = v_2591 | ~v_1167;
assign x_3080 = v_2591 | ~v_1168;
assign x_3081 = v_2591 | ~v_2301;
assign x_3082 = v_2591 | ~v_2302;
assign x_3083 = v_2591 | ~v_2389;
assign x_3084 = v_2591 | ~v_2390;
assign x_3085 = v_2591 | ~v_634;
assign x_3086 = v_2591 | ~v_635;
assign x_3087 = v_2591 | ~v_1169;
assign x_3088 = v_2591 | ~v_1170;
assign x_3089 = v_2591 | ~v_2331;
assign x_3090 = v_2591 | ~v_2332;
assign x_3091 = v_2591 | ~v_688;
assign x_3092 = v_2591 | ~v_689;
assign x_3093 = v_2591 | ~v_2334;
assign x_3094 = v_2591 | ~v_2335;
assign x_3095 = v_2591 | ~v_2391;
assign x_3096 = v_2591 | ~v_2392;
assign x_3097 = v_2591 | ~v_132;
assign x_3098 = v_2591 | ~v_127;
assign x_3099 = v_2591 | ~v_113;
assign x_3100 = v_2591 | ~v_112;
assign x_3101 = v_2591 | ~v_106;
assign x_3102 = v_2591 | ~v_105;
assign x_3103 = v_2591 | ~v_76;
assign x_3104 = v_2591 | ~v_75;
assign x_3105 = v_2591 | ~v_69;
assign x_3106 = v_2590 | ~v_2290;
assign x_3107 = v_2590 | ~v_2291;
assign x_3108 = v_2590 | ~v_2384;
assign x_3109 = v_2590 | ~v_2385;
assign x_3110 = v_2590 | ~v_615;
assign x_3111 = v_2590 | ~v_616;
assign x_3112 = v_2590 | ~v_1162;
assign x_3113 = v_2590 | ~v_1163;
assign x_3114 = v_2590 | ~v_2320;
assign x_3115 = v_2590 | ~v_2321;
assign x_3116 = v_2590 | ~v_669;
assign x_3117 = v_2590 | ~v_670;
assign x_3118 = v_2590 | ~v_1164;
assign x_3119 = v_2590 | ~v_1165;
assign x_3120 = v_2590 | ~v_2324;
assign x_3121 = v_2590 | ~v_2325;
assign x_3122 = v_2590 | ~v_2386;
assign x_3123 = v_2590 | ~v_2387;
assign x_3124 = v_2590 | ~v_131;
assign x_3125 = v_2590 | ~v_126;
assign x_3126 = v_2590 | ~v_111;
assign x_3127 = v_2590 | ~v_110;
assign x_3128 = v_2590 | ~v_102;
assign x_3129 = v_2590 | ~v_101;
assign x_3130 = v_2590 | ~v_51;
assign x_3131 = v_2590 | ~v_50;
assign x_3132 = v_2590 | ~v_44;
assign x_3133 = v_2589 | ~v_2279;
assign x_3134 = v_2589 | ~v_2379;
assign x_3135 = v_2589 | ~v_2380;
assign x_3136 = v_2589 | ~v_596;
assign x_3137 = v_2589 | ~v_597;
assign x_3138 = v_2589 | ~v_1157;
assign x_3139 = v_2589 | ~v_1158;
assign x_3140 = v_2589 | ~v_2312;
assign x_3141 = v_2589 | ~v_2313;
assign x_3142 = v_2589 | ~v_653;
assign x_3143 = v_2589 | ~v_654;
assign x_3144 = v_2589 | ~v_1159;
assign x_3145 = v_2589 | ~v_1160;
assign x_3146 = v_2589 | ~v_2282;
assign x_3147 = v_2589 | ~v_2314;
assign x_3148 = v_2589 | ~v_2315;
assign x_3149 = v_2589 | ~v_2381;
assign x_3150 = v_2589 | ~v_2382;
assign x_3151 = v_2589 | ~v_128;
assign x_3152 = v_2589 | ~v_122;
assign x_3153 = v_2589 | ~v_109;
assign x_3154 = v_2589 | ~v_108;
assign x_3155 = v_2589 | ~v_95;
assign x_3156 = v_2589 | ~v_94;
assign x_3157 = v_2589 | ~v_25;
assign x_3158 = v_2589 | ~v_24;
assign x_3159 = v_2589 | ~v_18;
assign x_3160 = ~v_2275 | ~v_2587 | v_2588;
assign x_3161 = v_2587 | ~v_2576;
assign x_3162 = v_2587 | ~v_2581;
assign x_3163 = v_2587 | ~v_2585;
assign x_3164 = v_2587 | ~v_2586;
assign x_3165 = ~v_2500 | ~v_2263 | v_2586;
assign x_3166 = ~v_2536 | ~v_2584 | v_2585;
assign x_3167 = v_2584 | ~v_2582;
assign x_3168 = v_2584 | ~v_2583;
assign x_3169 = v_2584 | ~v_2257;
assign x_3170 = v_2584 | ~v_2258;
assign x_3171 = v_2584 | ~v_2259;
assign x_3172 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2161 | ~v_2255 | v_2583;
assign x_3173 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2201 | ~v_2577 | v_2582;
assign x_3174 = ~v_2580 | ~v_2249 | v_2581;
assign x_3175 = v_2580 | ~v_2578;
assign x_3176 = v_2580 | ~v_2579;
assign x_3177 = v_2580 | ~v_2252;
assign x_3178 = v_2580 | ~v_2253;
assign x_3179 = v_2580 | ~v_2254;
assign x_3180 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2232 | ~v_2260 | v_2579;
assign x_3181 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2227 | ~v_2577 | v_2578;
assign x_3182 = v_2577 | ~v_2250;
assign x_3183 = v_2577 | ~v_2251;
assign x_3184 = v_2577 | ~v_2262;
assign x_3185 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2575 | v_2576;
assign x_3186 = v_2575 | ~v_2572;
assign x_3187 = v_2575 | ~v_2573;
assign x_3188 = v_2575 | ~v_2574;
assign x_3189 = v_76 | v_69 | v_75 | v_106 | v_105 | v_132 | v_127 | v_113 | v_112 | ~v_2182 | ~v_2181 | ~v_2125 | ~v_2124 | ~v_236 | ~v_235 | ~v_2122 | ~v_2121 | ~v_1141 | ~v_1140 | ~v_182 | ~v_181 | ~v_2180 | ~v_2179 | ~v_2092 | ~v_2091 | ~v_1139 | ~v_1138 | v_2574;
assign x_3190 = v_50 | v_51 | v_44 | v_101 | v_102 | v_111 | v_110 | v_131 | v_126 | ~v_2177 | ~v_2176 | ~v_2115 | ~v_2114 | ~v_1136 | ~v_1135 | ~v_217 | ~v_216 | ~v_2111 | ~v_2110 | ~v_1134 | ~v_1133 | ~v_163 | ~v_162 | ~v_2175 | ~v_2174 | ~v_2081 | ~v_2080 | v_2573;
assign x_3191 = v_25 | v_24 | v_18 | v_95 | v_94 | v_108 | v_109 | v_128 | v_122 | ~v_2172 | ~v_2171 | ~v_2105 | ~v_2104 | ~v_2073 | ~v_1131 | ~v_1130 | ~v_201 | ~v_200 | ~v_2103 | ~v_2102 | ~v_1129 | ~v_1128 | ~v_144 | ~v_143 | ~v_2170 | ~v_2169 | ~v_2069 | v_2572;
assign x_3192 = v_9 | v_7 | v_4 | v_6 | v_8 | v_10 | v_3 | v_2 | ~v_1041 | ~v_1040 | ~v_2570 | v_2571;
assign x_3193 = v_2570 | ~v_2565;
assign x_3194 = v_2570 | ~v_2569;
assign x_3195 = v_99 | ~v_2483 | ~v_1022 | ~v_1811 | ~v_2377 | ~v_2372 | ~v_2339 | ~v_2458 | ~v_2456 | ~v_2568 | ~v_2567 | v_2569;
assign x_3196 = v_2568 | ~v_2416;
assign x_3197 = v_2568 | ~v_2548;
assign x_3198 = v_2567 | ~v_2566;
assign x_3199 = v_2567 | ~v_2524;
assign x_3200 = ~v_2406 | ~v_2476 | ~v_2405 | ~v_2400 | ~v_2475 | v_2566;
assign x_3201 = ~v_2275 | ~v_2564 | v_2565;
assign x_3202 = v_2564 | ~v_2562;
assign x_3203 = v_2564 | ~v_2563;
assign x_3204 = v_2564 | ~v_2246;
assign x_3205 = v_2564 | ~v_2248;
assign x_3206 = v_2564 | ~v_2129;
assign x_3207 = v_2564 | ~v_2162;
assign x_3208 = v_2564 | ~v_2167;
assign x_3209 = ~v_2536 | ~v_2206 | v_2563;
assign x_3210 = ~v_2500 | ~v_2561 | v_2562;
assign x_3211 = v_2561 | ~v_2265;
assign x_3212 = v_2561 | ~v_2190;
assign x_3213 = v_2561 | ~v_2195;
assign x_3214 = v_2561 | ~v_2266;
assign x_3215 = v_2561 | ~v_2196;
assign x_3216 = v_9 | v_7 | v_5 | v_4 | v_6 | v_8 | v_3 | v_2 | ~v_1041 | ~v_1040 | ~v_2559 | v_2560;
assign x_3217 = v_2559 | ~v_2547;
assign x_3218 = v_2559 | ~v_2558;
assign x_3219 = v_99 | ~v_2483 | ~v_1022 | ~v_1811 | ~v_2523 | ~v_2522 | ~v_2517 | ~v_2516 | ~v_2515 | ~v_2557 | ~v_2553 | v_2558;
assign x_3220 = v_2557 | ~v_2459;
assign x_3221 = v_2557 | ~v_2556;
assign x_3222 = ~v_2513 | ~v_2512 | ~v_2511 | ~v_2555 | ~v_2554 | v_2556;
assign x_3223 = v_2555 | ~v_2442;
assign x_3224 = v_2555 | ~v_2521;
assign x_3225 = v_2555 | ~v_698;
assign x_3226 = v_2555 | ~v_699;
assign x_3227 = v_2555 | ~v_700;
assign x_3228 = v_2555 | ~v_701;
assign x_3229 = v_2554 | ~v_2432;
assign x_3230 = v_2554 | ~v_2550;
assign x_3231 = v_2554 | ~v_698;
assign x_3232 = v_2554 | ~v_699;
assign x_3233 = v_2554 | ~v_700;
assign x_3234 = v_2554 | ~v_701;
assign x_3235 = v_2553 | ~v_2548;
assign x_3236 = v_2553 | ~v_2552;
assign x_3237 = ~v_2520 | ~v_2519 | ~v_2518 | ~v_2551 | ~v_2549 | v_2552;
assign x_3238 = v_2551 | ~v_2550;
assign x_3239 = v_2551 | ~v_2394;
assign x_3240 = v_2551 | ~v_698;
assign x_3241 = v_2551 | ~v_699;
assign x_3242 = v_2551 | ~v_700;
assign x_3243 = v_2551 | ~v_701;
assign x_3244 = ~v_2523 | ~v_2517 | ~v_2516 | v_2550;
assign x_3245 = v_2549 | ~v_2514;
assign x_3246 = v_2549 | ~v_2371;
assign x_3247 = v_2549 | ~v_698;
assign x_3248 = v_2549 | ~v_699;
assign x_3249 = v_2549 | ~v_700;
assign x_3250 = v_2549 | ~v_701;
assign x_3251 = ~v_2448 | ~v_2447 | ~v_2446 | ~v_2532 | ~v_2531 | v_2548;
assign x_3252 = ~v_2275 | ~v_2546 | v_2547;
assign x_3253 = v_2546 | ~v_2541;
assign x_3254 = v_2546 | ~v_2545;
assign x_3255 = v_2546 | ~v_2491;
assign x_3256 = v_2546 | ~v_2492;
assign x_3257 = v_2546 | ~v_2493;
assign x_3258 = v_2546 | ~v_2498;
assign x_3259 = v_2546 | ~v_2499;
assign x_3260 = ~v_2544 | ~v_2249 | v_2545;
assign x_3261 = v_2544 | ~v_2542;
assign x_3262 = v_2544 | ~v_2543;
assign x_3263 = v_2544 | ~v_2487;
assign x_3264 = v_2544 | ~v_2488;
assign x_3265 = v_2544 | ~v_2489;
assign x_3266 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2497 | ~v_2232 | v_2543;
assign x_3267 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2538 | ~v_2222 | v_2542;
assign x_3268 = ~v_2540 | ~v_2536 | v_2541;
assign x_3269 = v_2540 | ~v_2537;
assign x_3270 = v_2540 | ~v_2539;
assign x_3271 = v_2540 | ~v_2494;
assign x_3272 = v_2540 | ~v_2495;
assign x_3273 = v_2540 | ~v_2496;
assign x_3274 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2184 | ~v_2538 | v_2539;
assign x_3275 = v_2538 | ~v_2492;
assign x_3276 = v_2538 | ~v_2493;
assign x_3277 = v_2538 | ~v_2499;
assign x_3278 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2161 | ~v_2490 | v_2537;
assign x_3279 = v_2536 | ~v_2507;
assign x_3280 = v_2536 | ~v_2508;
assign x_3281 = v_2536 | ~v_2236;
assign x_3282 = v_2536 | ~v_2237;
assign x_3283 = v_2536 | ~v_2238;
assign x_3284 = v_7 | v_5 | v_4 | v_8 | v_10 | v_3 | v_2 | ~v_1041 | ~v_1040 | ~v_2534 | v_2535;
assign x_3285 = v_2534 | ~v_2510;
assign x_3286 = v_2534 | ~v_2533;
assign x_3287 = v_99 | ~v_2483 | ~v_1022 | ~v_1811 | ~v_2448 | ~v_2447 | ~v_2446 | ~v_2532 | ~v_2531 | ~v_2530 | ~v_2525 | v_2533;
assign x_3288 = v_2532 | ~v_2527;
assign x_3289 = v_2532 | ~v_2338;
assign x_3290 = v_2532 | ~v_698;
assign x_3291 = v_2532 | ~v_699;
assign x_3292 = v_2532 | ~v_700;
assign x_3293 = v_2532 | ~v_701;
assign x_3294 = v_2531 | ~v_2444;
assign x_3295 = v_2531 | ~v_2376;
assign x_3296 = v_2531 | ~v_698;
assign x_3297 = v_2531 | ~v_699;
assign x_3298 = v_2531 | ~v_700;
assign x_3299 = v_2531 | ~v_701;
assign x_3300 = v_2530 | ~v_2459;
assign x_3301 = v_2530 | ~v_2529;
assign x_3302 = ~v_2443 | ~v_2438 | ~v_2433 | ~v_2528 | ~v_2526 | v_2529;
assign x_3303 = v_2528 | ~v_2527;
assign x_3304 = v_2528 | ~v_2437;
assign x_3305 = v_2528 | ~v_698;
assign x_3306 = v_2528 | ~v_699;
assign x_3307 = v_2528 | ~v_700;
assign x_3308 = v_2528 | ~v_701;
assign x_3309 = ~v_2453 | ~v_2452 | ~v_2451 | v_2527;
assign x_3310 = v_2526 | ~v_2449;
assign x_3311 = v_2526 | ~v_2432;
assign x_3312 = v_2526 | ~v_698;
assign x_3313 = v_2526 | ~v_699;
assign x_3314 = v_2526 | ~v_700;
assign x_3315 = v_2526 | ~v_701;
assign x_3316 = v_2525 | ~v_2454;
assign x_3317 = v_2525 | ~v_2524;
assign x_3318 = ~v_2523 | ~v_2522 | ~v_2517 | ~v_2516 | ~v_2515 | v_2524;
assign x_3319 = v_2523 | ~v_2338;
assign x_3320 = v_2523 | ~v_698;
assign x_3321 = v_2523 | ~v_699;
assign x_3322 = v_2523 | ~v_700;
assign x_3323 = v_2523 | ~v_701;
assign x_3324 = v_2522 | ~v_2355;
assign x_3325 = v_2522 | ~v_2521;
assign x_3326 = v_2522 | ~v_698;
assign x_3327 = v_2522 | ~v_699;
assign x_3328 = v_2522 | ~v_700;
assign x_3329 = v_2522 | ~v_701;
assign x_3330 = ~v_2520 | ~v_2519 | ~v_2518 | v_2521;
assign x_3331 = v_2520 | ~v_2411;
assign x_3332 = v_2520 | ~v_698;
assign x_3333 = v_2520 | ~v_699;
assign x_3334 = v_2520 | ~v_700;
assign x_3335 = v_2520 | ~v_701;
assign x_3336 = v_2519 | ~v_2437;
assign x_3337 = v_2519 | ~v_2371;
assign x_3338 = v_2519 | ~v_698;
assign x_3339 = v_2519 | ~v_699;
assign x_3340 = v_2519 | ~v_700;
assign x_3341 = v_2519 | ~v_701;
assign x_3342 = v_2518 | ~v_2394;
assign x_3343 = v_2518 | ~v_2338;
assign x_3344 = v_2518 | ~v_698;
assign x_3345 = v_2518 | ~v_699;
assign x_3346 = v_2518 | ~v_700;
assign x_3347 = v_2518 | ~v_701;
assign x_3348 = v_2517 | ~v_2355;
assign x_3349 = v_2517 | ~v_2411;
assign x_3350 = v_2517 | ~v_698;
assign x_3351 = v_2517 | ~v_699;
assign x_3352 = v_2517 | ~v_700;
assign x_3353 = v_2517 | ~v_701;
assign x_3354 = v_2516 | ~v_2376;
assign x_3355 = v_2516 | ~v_2437;
assign x_3356 = v_2516 | ~v_698;
assign x_3357 = v_2516 | ~v_699;
assign x_3358 = v_2516 | ~v_700;
assign x_3359 = v_2516 | ~v_701;
assign x_3360 = v_2515 | ~v_2514;
assign x_3361 = v_2515 | ~v_2376;
assign x_3362 = v_2515 | ~v_698;
assign x_3363 = v_2515 | ~v_699;
assign x_3364 = v_2515 | ~v_700;
assign x_3365 = v_2515 | ~v_701;
assign x_3366 = ~v_2513 | ~v_2512 | ~v_2511 | v_2514;
assign x_3367 = v_2513 | ~v_2437;
assign x_3368 = v_2513 | ~v_698;
assign x_3369 = v_2513 | ~v_699;
assign x_3370 = v_2513 | ~v_700;
assign x_3371 = v_2513 | ~v_701;
assign x_3372 = v_2512 | ~v_2442;
assign x_3373 = v_2512 | ~v_2411;
assign x_3374 = v_2512 | ~v_698;
assign x_3375 = v_2512 | ~v_699;
assign x_3376 = v_2512 | ~v_700;
assign x_3377 = v_2512 | ~v_701;
assign x_3378 = v_2511 | ~v_2432;
assign x_3379 = v_2511 | ~v_2338;
assign x_3380 = v_2511 | ~v_698;
assign x_3381 = v_2511 | ~v_699;
assign x_3382 = v_2511 | ~v_700;
assign x_3383 = v_2511 | ~v_701;
assign x_3384 = ~v_2275 | ~v_2509 | v_2510;
assign x_3385 = v_2509 | ~v_2501;
assign x_3386 = v_2509 | ~v_2506;
assign x_3387 = v_2509 | ~v_2507;
assign x_3388 = v_2509 | ~v_2508;
assign x_3389 = v_2509 | ~v_2236;
assign x_3390 = v_2509 | ~v_2237;
assign x_3391 = v_2509 | ~v_2238;
assign x_3392 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2128 | ~v_2503 | v_2508;
assign x_3393 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2166 | ~v_2234 | v_2507;
assign x_3394 = ~v_2505 | ~v_2249 | v_2506;
assign x_3395 = v_2505 | ~v_2502;
assign x_3396 = v_2505 | ~v_2504;
assign x_3397 = v_2505 | ~v_2223;
assign x_3398 = v_2505 | ~v_2228;
assign x_3399 = v_2505 | ~v_2233;
assign x_3400 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2227 | ~v_2503 | v_2504;
assign x_3401 = v_2503 | ~v_2241;
assign x_3402 = v_2503 | ~v_2242;
assign x_3403 = v_2503 | ~v_2243;
assign x_3404 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2222 | ~v_2239 | v_2502;
assign x_3405 = ~v_2500 | ~v_2244 | v_2501;
assign x_3406 = v_2500 | ~v_2491;
assign x_3407 = v_2500 | ~v_2492;
assign x_3408 = v_2500 | ~v_2493;
assign x_3409 = v_2500 | ~v_2498;
assign x_3410 = v_2500 | ~v_2499;
assign x_3411 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2128 | v_2499;
assign x_3412 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2497 | ~v_2145 | v_2498;
assign x_3413 = v_2497 | ~v_2494;
assign x_3414 = v_2497 | ~v_2495;
assign x_3415 = v_2497 | ~v_2496;
assign x_3416 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2201 | v_2496;
assign x_3417 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2161 | ~v_2227 | v_2495;
assign x_3418 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2128 | ~v_2184 | v_2494;
assign x_3419 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2201 | ~v_2145 | v_2493;
assign x_3420 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2227 | ~v_2166 | v_2492;
assign x_3421 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2166 | ~v_2490 | v_2491;
assign x_3422 = v_2490 | ~v_2487;
assign x_3423 = v_2490 | ~v_2488;
assign x_3424 = v_2490 | ~v_2489;
assign x_3425 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2227 | v_2489;
assign x_3426 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2201 | ~v_2232 | v_2488;
assign x_3427 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2128 | ~v_2222 | v_2487;
assign x_3428 = v_9 | v_7 | v_4 | v_6 | v_10 | v_3 | v_2 | v_1 | ~v_1041 | ~v_1040 | ~v_2485 | v_2486;
assign x_3429 = v_2485 | ~v_2276;
assign x_3430 = v_2485 | ~v_2484;
assign x_3431 = v_99 | ~v_2483 | ~v_1022 | ~v_1811 | ~v_2406 | ~v_2476 | ~v_2405 | ~v_2400 | ~v_2475 | ~v_2474 | ~v_2455 | v_2484;
assign x_3432 = v_2483 | ~v_2479;
assign x_3433 = v_2483 | ~v_2482;
assign x_3434 = v_98 | ~v_1033 | ~v_1032 | ~v_2481 | ~v_2480 | v_2482;
assign x_3435 = v_2481 | ~v_1030;
assign x_3436 = v_2481 | v_119;
assign x_3437 = v_2480 | ~v_1815;
assign x_3438 = v_2480 | v_130;
assign x_3439 = v_97 | ~v_1012 | ~v_1011 | ~v_2478 | ~v_2477 | v_2479;
assign x_3440 = v_2478 | ~v_1017;
assign x_3441 = v_2478 | v_114;
assign x_3442 = v_2477 | ~v_1807;
assign x_3443 = v_2477 | v_123;
assign x_3444 = v_2476 | ~v_2457;
assign x_3445 = v_2476 | ~v_2404;
assign x_3446 = v_2476 | ~v_698;
assign x_3447 = v_2476 | ~v_699;
assign x_3448 = v_2476 | ~v_700;
assign x_3449 = v_2476 | ~v_701;
assign x_3450 = v_2475 | ~v_2378;
assign x_3451 = v_2475 | ~v_2399;
assign x_3452 = v_2475 | ~v_698;
assign x_3453 = v_2475 | ~v_699;
assign x_3454 = v_2475 | ~v_700;
assign x_3455 = v_2475 | ~v_701;
assign x_3456 = v_2474 | ~v_2459;
assign x_3457 = v_2474 | ~v_2473;
assign x_3458 = ~v_2472 | ~v_2471 | ~v_2466 | ~v_2461 | ~v_2460 | v_2473;
assign x_3459 = v_2472 | ~v_2399;
assign x_3460 = v_2472 | ~v_698;
assign x_3461 = v_2472 | ~v_699;
assign x_3462 = v_2472 | ~v_700;
assign x_3463 = v_2472 | ~v_701;
assign x_3464 = v_2471 | ~v_2404;
assign x_3465 = v_2471 | ~v_2470;
assign x_3466 = v_2471 | ~v_698;
assign x_3467 = v_2471 | ~v_699;
assign x_3468 = v_2471 | ~v_700;
assign x_3469 = v_2471 | ~v_701;
assign x_3470 = ~v_2469 | ~v_2468 | ~v_2467 | v_2470;
assign x_3471 = v_2469 | ~v_2394;
assign x_3472 = v_2469 | ~v_698;
assign x_3473 = v_2469 | ~v_699;
assign x_3474 = v_2469 | ~v_700;
assign x_3475 = v_2469 | ~v_701;
assign x_3476 = v_2468 | ~v_2399;
assign x_3477 = v_2468 | ~v_2411;
assign x_3478 = v_2468 | ~v_698;
assign x_3479 = v_2468 | ~v_699;
assign x_3480 = v_2468 | ~v_700;
assign x_3481 = v_2468 | ~v_701;
assign x_3482 = v_2467 | ~v_2432;
assign x_3483 = v_2467 | ~v_2371;
assign x_3484 = v_2467 | ~v_698;
assign x_3485 = v_2467 | ~v_699;
assign x_3486 = v_2467 | ~v_700;
assign x_3487 = v_2467 | ~v_701;
assign x_3488 = v_2466 | ~v_2310;
assign x_3489 = v_2466 | ~v_2465;
assign x_3490 = v_2466 | ~v_698;
assign x_3491 = v_2466 | ~v_699;
assign x_3492 = v_2466 | ~v_700;
assign x_3493 = v_2466 | ~v_701;
assign x_3494 = ~v_2464 | ~v_2463 | ~v_2462 | v_2465;
assign x_3495 = v_2464 | ~v_2432;
assign x_3496 = v_2464 | ~v_698;
assign x_3497 = v_2464 | ~v_699;
assign x_3498 = v_2464 | ~v_700;
assign x_3499 = v_2464 | ~v_701;
assign x_3500 = v_2463 | ~v_2399;
assign x_3501 = v_2463 | ~v_2437;
assign x_3502 = v_2463 | ~v_698;
assign x_3503 = v_2463 | ~v_699;
assign x_3504 = v_2463 | ~v_700;
assign x_3505 = v_2463 | ~v_701;
assign x_3506 = v_2462 | ~v_2442;
assign x_3507 = v_2462 | ~v_2394;
assign x_3508 = v_2462 | ~v_698;
assign x_3509 = v_2462 | ~v_699;
assign x_3510 = v_2462 | ~v_700;
assign x_3511 = v_2462 | ~v_701;
assign x_3512 = v_2461 | ~v_2404;
assign x_3513 = v_2461 | ~v_2394;
assign x_3514 = v_2461 | ~v_698;
assign x_3515 = v_2461 | ~v_699;
assign x_3516 = v_2461 | ~v_700;
assign x_3517 = v_2461 | ~v_701;
assign x_3518 = v_2460 | ~v_2310;
assign x_3519 = v_2460 | ~v_2432;
assign x_3520 = v_2460 | ~v_698;
assign x_3521 = v_2460 | ~v_699;
assign x_3522 = v_2460 | ~v_700;
assign x_3523 = v_2460 | ~v_701;
assign x_3524 = ~v_2377 | ~v_2372 | ~v_2339 | ~v_2458 | ~v_2456 | v_2459;
assign x_3525 = v_2458 | ~v_2457;
assign x_3526 = v_2458 | ~v_2355;
assign x_3527 = v_2458 | ~v_698;
assign x_3528 = v_2458 | ~v_699;
assign x_3529 = v_2458 | ~v_700;
assign x_3530 = v_2458 | ~v_701;
assign x_3531 = ~v_2415 | ~v_2414 | ~v_2413 | v_2457;
assign x_3532 = v_2456 | ~v_2407;
assign x_3533 = v_2456 | ~v_2338;
assign x_3534 = v_2456 | ~v_698;
assign x_3535 = v_2456 | ~v_699;
assign x_3536 = v_2456 | ~v_700;
assign x_3537 = v_2456 | ~v_701;
assign x_3538 = v_2455 | ~v_2416;
assign x_3539 = v_2455 | ~v_2454;
assign x_3540 = ~v_2453 | ~v_2452 | ~v_2451 | ~v_2450 | ~v_2445 | v_2454;
assign x_3541 = v_2453 | ~v_2404;
assign x_3542 = v_2453 | ~v_698;
assign x_3543 = v_2453 | ~v_699;
assign x_3544 = v_2453 | ~v_700;
assign x_3545 = v_2453 | ~v_701;
assign x_3546 = v_2452 | ~v_2399;
assign x_3547 = v_2452 | ~v_2355;
assign x_3548 = v_2452 | ~v_698;
assign x_3549 = v_2452 | ~v_699;
assign x_3550 = v_2452 | ~v_700;
assign x_3551 = v_2452 | ~v_701;
assign x_3552 = v_2451 | ~v_2310;
assign x_3553 = v_2451 | ~v_2442;
assign x_3554 = v_2451 | ~v_698;
assign x_3555 = v_2451 | ~v_699;
assign x_3556 = v_2451 | ~v_700;
assign x_3557 = v_2451 | ~v_701;
assign x_3558 = v_2450 | ~v_2449;
assign x_3559 = v_2450 | ~v_2399;
assign x_3560 = v_2450 | ~v_698;
assign x_3561 = v_2450 | ~v_699;
assign x_3562 = v_2450 | ~v_700;
assign x_3563 = v_2450 | ~v_701;
assign x_3564 = ~v_2448 | ~v_2447 | ~v_2446 | v_2449;
assign x_3565 = v_2448 | ~v_2355;
assign x_3566 = v_2448 | ~v_698;
assign x_3567 = v_2448 | ~v_699;
assign x_3568 = v_2448 | ~v_700;
assign x_3569 = v_2448 | ~v_701;
assign x_3570 = v_2447 | ~v_2404;
assign x_3571 = v_2447 | ~v_2338;
assign x_3572 = v_2447 | ~v_698;
assign x_3573 = v_2447 | ~v_699;
assign x_3574 = v_2447 | ~v_700;
assign x_3575 = v_2447 | ~v_701;
assign x_3576 = v_2446 | ~v_2442;
assign x_3577 = v_2446 | ~v_2376;
assign x_3578 = v_2446 | ~v_698;
assign x_3579 = v_2446 | ~v_699;
assign x_3580 = v_2446 | ~v_700;
assign x_3581 = v_2446 | ~v_701;
assign x_3582 = v_2445 | ~v_2444;
assign x_3583 = v_2445 | ~v_2310;
assign x_3584 = v_2445 | ~v_698;
assign x_3585 = v_2445 | ~v_699;
assign x_3586 = v_2445 | ~v_700;
assign x_3587 = v_2445 | ~v_701;
assign x_3588 = ~v_2443 | ~v_2438 | ~v_2433 | v_2444;
assign x_3589 = v_2443 | ~v_2442;
assign x_3590 = v_2443 | ~v_698;
assign x_3591 = v_2443 | ~v_699;
assign x_3592 = v_2443 | ~v_700;
assign x_3593 = v_2443 | ~v_701;
assign x_3594 = ~v_2441 | ~v_2440 | ~v_2439 | v_2442;
assign x_3595 = v_2441 | ~v_2427;
assign x_3596 = v_2441 | ~v_2428;
assign x_3597 = v_2441 | ~v_782;
assign x_3598 = v_2441 | ~v_783;
assign x_3599 = v_2441 | ~v_682;
assign x_3600 = v_2441 | ~v_683;
assign x_3601 = v_2441 | ~v_2301;
assign x_3602 = v_2441 | ~v_2302;
assign x_3603 = v_2441 | ~v_2350;
assign x_3604 = v_2441 | ~v_2351;
assign x_3605 = v_2441 | ~v_2352;
assign x_3606 = v_2441 | ~v_632;
assign x_3607 = v_2441 | ~v_633;
assign x_3608 = v_2441 | ~v_784;
assign x_3609 = v_2441 | ~v_785;
assign x_3610 = v_2441 | ~v_2353;
assign x_3611 = v_2441 | ~v_2429;
assign x_3612 = v_2441 | ~v_2430;
assign x_3613 = v_2441 | ~v_121;
assign x_3614 = v_2441 | ~v_113;
assign x_3615 = v_2441 | ~v_112;
assign x_3616 = v_2441 | ~v_106;
assign x_3617 = v_2441 | ~v_104;
assign x_3618 = v_2441 | ~v_75;
assign x_3619 = v_2441 | ~v_74;
assign x_3620 = v_2441 | ~v_73;
assign x_3621 = v_2441 | ~v_70;
assign x_3622 = v_2440 | ~v_2422;
assign x_3623 = v_2440 | ~v_2423;
assign x_3624 = v_2440 | ~v_777;
assign x_3625 = v_2440 | ~v_778;
assign x_3626 = v_2440 | ~v_2290;
assign x_3627 = v_2440 | ~v_2291;
assign x_3628 = v_2440 | ~v_613;
assign x_3629 = v_2440 | ~v_614;
assign x_3630 = v_2440 | ~v_779;
assign x_3631 = v_2440 | ~v_780;
assign x_3632 = v_2440 | ~v_2345;
assign x_3633 = v_2440 | ~v_2346;
assign x_3634 = v_2440 | ~v_2424;
assign x_3635 = v_2440 | ~v_2347;
assign x_3636 = v_2440 | ~v_2348;
assign x_3637 = v_2440 | ~v_677;
assign x_3638 = v_2440 | ~v_678;
assign x_3639 = v_2440 | ~v_2425;
assign x_3640 = v_2440 | ~v_120;
assign x_3641 = v_2440 | ~v_111;
assign x_3642 = v_2440 | ~v_110;
assign x_3643 = v_2440 | ~v_102;
assign x_3644 = v_2440 | ~v_100;
assign x_3645 = v_2440 | ~v_50;
assign x_3646 = v_2440 | ~v_49;
assign x_3647 = v_2440 | ~v_48;
assign x_3648 = v_2440 | ~v_45;
assign x_3649 = v_2439 | ~v_2417;
assign x_3650 = v_2439 | ~v_2418;
assign x_3651 = v_2439 | ~v_772;
assign x_3652 = v_2439 | ~v_773;
assign x_3653 = v_2439 | ~v_646;
assign x_3654 = v_2439 | ~v_2279;
assign x_3655 = v_2439 | ~v_2340;
assign x_3656 = v_2439 | ~v_2341;
assign x_3657 = v_2439 | ~v_594;
assign x_3658 = v_2439 | ~v_595;
assign x_3659 = v_2439 | ~v_774;
assign x_3660 = v_2439 | ~v_775;
assign x_3661 = v_2439 | ~v_2282;
assign x_3662 = v_2439 | ~v_2419;
assign x_3663 = v_2439 | ~v_2420;
assign x_3664 = v_2439 | ~v_661;
assign x_3665 = v_2439 | ~v_2342;
assign x_3666 = v_2439 | ~v_2343;
assign x_3667 = v_2439 | ~v_117;
assign x_3668 = v_2439 | ~v_109;
assign x_3669 = v_2439 | ~v_108;
assign x_3670 = v_2439 | ~v_95;
assign x_3671 = v_2439 | ~v_93;
assign x_3672 = v_2439 | ~v_24;
assign x_3673 = v_2439 | ~v_23;
assign x_3674 = v_2439 | ~v_22;
assign x_3675 = v_2439 | ~v_19;
assign x_3676 = v_2438 | ~v_2404;
assign x_3677 = v_2438 | ~v_2437;
assign x_3678 = v_2438 | ~v_698;
assign x_3679 = v_2438 | ~v_699;
assign x_3680 = v_2438 | ~v_700;
assign x_3681 = v_2438 | ~v_701;
assign x_3682 = ~v_2436 | ~v_2435 | ~v_2434 | v_2437;
assign x_3683 = v_2436 | ~v_761;
assign x_3684 = v_2436 | ~v_762;
assign x_3685 = v_2436 | ~v_2427;
assign x_3686 = v_2436 | ~v_2428;
assign x_3687 = v_2436 | ~v_2301;
assign x_3688 = v_2436 | ~v_2302;
assign x_3689 = v_2436 | ~v_763;
assign x_3690 = v_2436 | ~v_764;
assign x_3691 = v_2436 | ~v_2329;
assign x_3692 = v_2436 | ~v_2330;
assign x_3693 = v_2436 | ~v_765;
assign x_3694 = v_2436 | ~v_766;
assign x_3695 = v_2436 | ~v_632;
assign x_3696 = v_2436 | ~v_633;
assign x_3697 = v_2436 | ~v_2333;
assign x_3698 = v_2436 | ~v_2429;
assign x_3699 = v_2436 | ~v_2430;
assign x_3700 = v_2436 | ~v_2336;
assign x_3701 = v_2436 | ~v_113;
assign x_3702 = v_2436 | ~v_112;
assign x_3703 = v_2436 | ~v_105;
assign x_3704 = v_2436 | ~v_104;
assign x_3705 = v_2436 | ~v_76;
assign x_3706 = v_2436 | ~v_75;
assign x_3707 = v_2436 | ~v_74;
assign x_3708 = v_2436 | ~v_73;
assign x_3709 = v_2436 | ~v_72;
assign x_3710 = v_2435 | ~v_2422;
assign x_3711 = v_2435 | ~v_2423;
assign x_3712 = v_2435 | ~v_2290;
assign x_3713 = v_2435 | ~v_2291;
assign x_3714 = v_2435 | ~v_750;
assign x_3715 = v_2435 | ~v_751;
assign x_3716 = v_2435 | ~v_752;
assign x_3717 = v_2435 | ~v_613;
assign x_3718 = v_2435 | ~v_614;
assign x_3719 = v_2435 | ~v_753;
assign x_3720 = v_2435 | ~v_754;
assign x_3721 = v_2435 | ~v_2322;
assign x_3722 = v_2435 | ~v_2323;
assign x_3723 = v_2435 | ~v_2424;
assign x_3724 = v_2435 | ~v_757;
assign x_3725 = v_2435 | ~v_2326;
assign x_3726 = v_2435 | ~v_2327;
assign x_3727 = v_2435 | ~v_2425;
assign x_3728 = v_2435 | ~v_111;
assign x_3729 = v_2435 | ~v_110;
assign x_3730 = v_2435 | ~v_101;
assign x_3731 = v_2435 | ~v_100;
assign x_3732 = v_2435 | ~v_51;
assign x_3733 = v_2435 | ~v_50;
assign x_3734 = v_2435 | ~v_49;
assign x_3735 = v_2435 | ~v_48;
assign x_3736 = v_2435 | ~v_47;
assign x_3737 = v_2434 | ~v_2417;
assign x_3738 = v_2434 | ~v_2418;
assign x_3739 = v_2434 | ~v_2279;
assign x_3740 = v_2434 | ~v_739;
assign x_3741 = v_2434 | ~v_2311;
assign x_3742 = v_2434 | ~v_740;
assign x_3743 = v_2434 | ~v_741;
assign x_3744 = v_2434 | ~v_594;
assign x_3745 = v_2434 | ~v_595;
assign x_3746 = v_2434 | ~v_742;
assign x_3747 = v_2434 | ~v_743;
assign x_3748 = v_2434 | ~v_2282;
assign x_3749 = v_2434 | ~v_2419;
assign x_3750 = v_2434 | ~v_2420;
assign x_3751 = v_2434 | ~v_746;
assign x_3752 = v_2434 | ~v_2316;
assign x_3753 = v_2434 | ~v_2317;
assign x_3754 = v_2434 | ~v_2318;
assign x_3755 = v_2434 | ~v_109;
assign x_3756 = v_2434 | ~v_108;
assign x_3757 = v_2434 | ~v_94;
assign x_3758 = v_2434 | ~v_93;
assign x_3759 = v_2434 | ~v_25;
assign x_3760 = v_2434 | ~v_24;
assign x_3761 = v_2434 | ~v_23;
assign x_3762 = v_2434 | ~v_22;
assign x_3763 = v_2434 | ~v_21;
assign x_3764 = v_2433 | ~v_2432;
assign x_3765 = v_2433 | ~v_2355;
assign x_3766 = v_2433 | ~v_698;
assign x_3767 = v_2433 | ~v_699;
assign x_3768 = v_2433 | ~v_700;
assign x_3769 = v_2433 | ~v_701;
assign x_3770 = ~v_2431 | ~v_2426 | ~v_2421 | v_2432;
assign x_3771 = v_2431 | ~v_630;
assign x_3772 = v_2431 | ~v_631;
assign x_3773 = v_2431 | ~v_2427;
assign x_3774 = v_2431 | ~v_2428;
assign x_3775 = v_2431 | ~v_2301;
assign x_3776 = v_2431 | ~v_2302;
assign x_3777 = v_2431 | ~v_632;
assign x_3778 = v_2431 | ~v_633;
assign x_3779 = v_2431 | ~v_2389;
assign x_3780 = v_2431 | ~v_2390;
assign x_3781 = v_2431 | ~v_634;
assign x_3782 = v_2431 | ~v_635;
assign x_3783 = v_2431 | ~v_636;
assign x_3784 = v_2431 | ~v_637;
assign x_3785 = v_2431 | ~v_2429;
assign x_3786 = v_2431 | ~v_2430;
assign x_3787 = v_2431 | ~v_2391;
assign x_3788 = v_2431 | ~v_2392;
assign x_3789 = v_2431 | ~v_127;
assign x_3790 = v_2431 | ~v_113;
assign x_3791 = v_2431 | ~v_112;
assign x_3792 = v_2431 | ~v_107;
assign x_3793 = v_2431 | ~v_106;
assign x_3794 = v_2431 | ~v_105;
assign x_3795 = v_2431 | ~v_104;
assign x_3796 = v_2431 | ~v_76;
assign x_3797 = v_2431 | ~v_73;
assign x_3798 = ~v_86 | ~v_119 | v_2430;
assign x_3799 = ~v_78 | v_119 | v_2429;
assign x_3800 = ~v_88 | ~v_118 | v_2428;
assign x_3801 = ~v_80 | v_118 | v_2427;
assign x_3802 = v_2426 | ~v_611;
assign x_3803 = v_2426 | ~v_612;
assign x_3804 = v_2426 | ~v_2422;
assign x_3805 = v_2426 | ~v_2423;
assign x_3806 = v_2426 | ~v_2290;
assign x_3807 = v_2426 | ~v_2291;
assign x_3808 = v_2426 | ~v_613;
assign x_3809 = v_2426 | ~v_614;
assign x_3810 = v_2426 | ~v_2384;
assign x_3811 = v_2426 | ~v_2385;
assign x_3812 = v_2426 | ~v_615;
assign x_3813 = v_2426 | ~v_616;
assign x_3814 = v_2426 | ~v_617;
assign x_3815 = v_2426 | ~v_618;
assign x_3816 = v_2426 | ~v_2424;
assign x_3817 = v_2426 | ~v_2386;
assign x_3818 = v_2426 | ~v_2387;
assign x_3819 = v_2426 | ~v_2425;
assign x_3820 = v_2426 | ~v_126;
assign x_3821 = v_2426 | ~v_111;
assign x_3822 = v_2426 | ~v_110;
assign x_3823 = v_2426 | ~v_103;
assign x_3824 = v_2426 | ~v_102;
assign x_3825 = v_2426 | ~v_101;
assign x_3826 = v_2426 | ~v_100;
assign x_3827 = v_2426 | ~v_51;
assign x_3828 = v_2426 | ~v_48;
assign x_3829 = ~v_61 | ~v_119 | v_2425;
assign x_3830 = ~v_53 | v_119 | v_2424;
assign x_3831 = ~v_63 | ~v_118 | v_2423;
assign x_3832 = ~v_55 | v_118 | v_2422;
assign x_3833 = v_2421 | ~v_592;
assign x_3834 = v_2421 | ~v_593;
assign x_3835 = v_2421 | ~v_2417;
assign x_3836 = v_2421 | ~v_2418;
assign x_3837 = v_2421 | ~v_2279;
assign x_3838 = v_2421 | ~v_594;
assign x_3839 = v_2421 | ~v_595;
assign x_3840 = v_2421 | ~v_2379;
assign x_3841 = v_2421 | ~v_2380;
assign x_3842 = v_2421 | ~v_596;
assign x_3843 = v_2421 | ~v_597;
assign x_3844 = v_2421 | ~v_598;
assign x_3845 = v_2421 | ~v_599;
assign x_3846 = v_2421 | ~v_2282;
assign x_3847 = v_2421 | ~v_2419;
assign x_3848 = v_2421 | ~v_2420;
assign x_3849 = v_2421 | ~v_2381;
assign x_3850 = v_2421 | ~v_2382;
assign x_3851 = v_2421 | ~v_122;
assign x_3852 = v_2421 | ~v_109;
assign x_3853 = v_2421 | ~v_108;
assign x_3854 = v_2421 | ~v_96;
assign x_3855 = v_2421 | ~v_95;
assign x_3856 = v_2421 | ~v_94;
assign x_3857 = v_2421 | ~v_93;
assign x_3858 = v_2421 | ~v_25;
assign x_3859 = v_2421 | ~v_22;
assign x_3860 = ~v_36 | ~v_119 | v_2420;
assign x_3861 = ~v_28 | v_119 | v_2419;
assign x_3862 = ~v_38 | ~v_118 | v_2418;
assign x_3863 = ~v_30 | v_118 | v_2417;
assign x_3864 = ~v_2415 | ~v_2414 | ~v_2413 | ~v_2412 | ~v_2395 | v_2416;
assign x_3865 = v_2415 | ~v_2371;
assign x_3866 = v_2415 | ~v_698;
assign x_3867 = v_2415 | ~v_699;
assign x_3868 = v_2415 | ~v_700;
assign x_3869 = v_2415 | ~v_701;
assign x_3870 = v_2414 | ~v_2310;
assign x_3871 = v_2414 | ~v_2411;
assign x_3872 = v_2414 | ~v_698;
assign x_3873 = v_2414 | ~v_699;
assign x_3874 = v_2414 | ~v_700;
assign x_3875 = v_2414 | ~v_701;
assign x_3876 = v_2413 | ~v_2376;
assign x_3877 = v_2413 | ~v_2394;
assign x_3878 = v_2413 | ~v_698;
assign x_3879 = v_2413 | ~v_699;
assign x_3880 = v_2413 | ~v_700;
assign x_3881 = v_2413 | ~v_701;
assign x_3882 = v_2412 | ~v_2407;
assign x_3883 = v_2412 | ~v_2411;
assign x_3884 = v_2412 | ~v_698;
assign x_3885 = v_2412 | ~v_699;
assign x_3886 = v_2412 | ~v_700;
assign x_3887 = v_2412 | ~v_701;
assign x_3888 = ~v_2410 | ~v_2409 | ~v_2408 | v_2411;
assign x_3889 = v_2410 | ~v_906;
assign x_3890 = v_2410 | ~v_907;
assign x_3891 = v_2410 | ~v_2301;
assign x_3892 = v_2410 | ~v_2302;
assign x_3893 = v_2410 | ~v_2366;
assign x_3894 = v_2410 | ~v_2367;
assign x_3895 = v_2410 | ~v_908;
assign x_3896 = v_2410 | ~v_909;
assign x_3897 = v_2410 | ~v_910;
assign x_3898 = v_2410 | ~v_763;
assign x_3899 = v_2410 | ~v_764;
assign x_3900 = v_2410 | ~v_2329;
assign x_3901 = v_2410 | ~v_2330;
assign x_3902 = v_2410 | ~v_2368;
assign x_3903 = v_2410 | ~v_2333;
assign x_3904 = v_2410 | ~v_2369;
assign x_3905 = v_2410 | ~v_914;
assign x_3906 = v_2410 | ~v_2336;
assign x_3907 = v_2410 | ~v_121;
assign x_3908 = v_2410 | ~v_113;
assign x_3909 = v_2410 | ~v_105;
assign x_3910 = v_2410 | ~v_104;
assign x_3911 = v_2410 | ~v_75;
assign x_3912 = v_2410 | ~v_74;
assign x_3913 = v_2410 | ~v_73;
assign x_3914 = v_2410 | ~v_72;
assign x_3915 = v_2410 | ~v_68;
assign x_3916 = v_2409 | ~v_2290;
assign x_3917 = v_2409 | ~v_2291;
assign x_3918 = v_2409 | ~v_896;
assign x_3919 = v_2409 | ~v_750;
assign x_3920 = v_2409 | ~v_2322;
assign x_3921 = v_2409 | ~v_2323;
assign x_3922 = v_2409 | ~v_2361;
assign x_3923 = v_2409 | ~v_2362;
assign x_3924 = v_2409 | ~v_897;
assign x_3925 = v_2409 | ~v_757;
assign x_3926 = v_2409 | ~v_900;
assign x_3927 = v_2409 | ~v_2363;
assign x_3928 = v_2409 | ~v_2326;
assign x_3929 = v_2409 | ~v_2327;
assign x_3930 = v_2409 | ~v_901;
assign x_3931 = v_2409 | ~v_2364;
assign x_3932 = v_2409 | ~v_902;
assign x_3933 = v_2409 | ~v_903;
assign x_3934 = v_2409 | ~v_120;
assign x_3935 = v_2409 | ~v_111;
assign x_3936 = v_2409 | ~v_101;
assign x_3937 = v_2409 | ~v_100;
assign x_3938 = v_2409 | ~v_50;
assign x_3939 = v_2409 | ~v_49;
assign x_3940 = v_2409 | ~v_48;
assign x_3941 = v_2409 | ~v_47;
assign x_3942 = v_2409 | ~v_43;
assign x_3943 = v_2408 | ~v_885;
assign x_3944 = v_2408 | ~v_2279;
assign x_3945 = v_2408 | ~v_2356;
assign x_3946 = v_2408 | ~v_2357;
assign x_3947 = v_2408 | ~v_2358;
assign x_3948 = v_2408 | ~v_886;
assign x_3949 = v_2408 | ~v_887;
assign x_3950 = v_2408 | ~v_739;
assign x_3951 = v_2408 | ~v_2311;
assign x_3952 = v_2408 | ~v_2359;
assign x_3953 = v_2408 | ~v_2282;
assign x_3954 = v_2408 | ~v_746;
assign x_3955 = v_2408 | ~v_890;
assign x_3956 = v_2408 | ~v_2316;
assign x_3957 = v_2408 | ~v_891;
assign x_3958 = v_2408 | ~v_2317;
assign x_3959 = v_2408 | ~v_892;
assign x_3960 = v_2408 | ~v_117;
assign x_3961 = v_2408 | ~v_2318;
assign x_3962 = v_2408 | ~v_109;
assign x_3963 = v_2408 | ~v_94;
assign x_3964 = v_2408 | ~v_93;
assign x_3965 = v_2408 | ~v_24;
assign x_3966 = v_2408 | ~v_23;
assign x_3967 = v_2408 | ~v_22;
assign x_3968 = v_2408 | ~v_21;
assign x_3969 = v_2408 | ~v_17;
assign x_3970 = ~v_2406 | ~v_2405 | ~v_2400 | v_2407;
assign x_3971 = v_2406 | ~v_2310;
assign x_3972 = v_2406 | ~v_698;
assign x_3973 = v_2406 | ~v_699;
assign x_3974 = v_2406 | ~v_700;
assign x_3975 = v_2406 | ~v_701;
assign x_3976 = v_2405 | ~v_2404;
assign x_3977 = v_2405 | ~v_2371;
assign x_3978 = v_2405 | ~v_698;
assign x_3979 = v_2405 | ~v_699;
assign x_3980 = v_2405 | ~v_700;
assign x_3981 = v_2405 | ~v_701;
assign x_3982 = ~v_2403 | ~v_2402 | ~v_2401 | v_2404;
assign x_3983 = v_2403 | ~v_682;
assign x_3984 = v_2403 | ~v_683;
assign x_3985 = v_2403 | ~v_2301;
assign x_3986 = v_2403 | ~v_2302;
assign x_3987 = v_2403 | ~v_2350;
assign x_3988 = v_2403 | ~v_2351;
assign x_3989 = v_2403 | ~v_2352;
assign x_3990 = v_2403 | ~v_725;
assign x_3991 = v_2403 | ~v_726;
assign x_3992 = v_2403 | ~v_727;
assign x_3993 = v_2403 | ~v_728;
assign x_3994 = v_2403 | ~v_2303;
assign x_3995 = v_2403 | ~v_2304;
assign x_3996 = v_2403 | ~v_2305;
assign x_3997 = v_2403 | ~v_2353;
assign x_3998 = v_2403 | ~v_731;
assign x_3999 = v_2403 | ~v_734;
assign x_4000 = v_2403 | ~v_2307;
assign x_4001 = v_2403 | ~v_112;
assign x_4002 = v_2403 | ~v_107;
assign x_4003 = v_2403 | ~v_106;
assign x_4004 = v_2403 | ~v_104;
assign x_4005 = v_2403 | ~v_76;
assign x_4006 = v_2403 | ~v_74;
assign x_4007 = v_2403 | ~v_73;
assign x_4008 = v_2403 | ~v_71;
assign x_4009 = v_2403 | ~v_70;
assign x_4010 = v_2402 | ~v_2290;
assign x_4011 = v_2402 | ~v_2291;
assign x_4012 = v_2402 | ~v_714;
assign x_4013 = v_2402 | ~v_715;
assign x_4014 = v_2402 | ~v_2345;
assign x_4015 = v_2402 | ~v_2292;
assign x_4016 = v_2402 | ~v_2346;
assign x_4017 = v_2402 | ~v_718;
assign x_4018 = v_2402 | ~v_2293;
assign x_4019 = v_2402 | ~v_721;
assign x_4020 = v_2402 | ~v_2347;
assign x_4021 = v_2402 | ~v_2348;
assign x_4022 = v_2402 | ~v_2295;
assign x_4023 = v_2402 | ~v_677;
assign x_4024 = v_2402 | ~v_722;
assign x_4025 = v_2402 | ~v_678;
assign x_4026 = v_2402 | ~v_2296;
assign x_4027 = v_2402 | ~v_723;
assign x_4028 = v_2402 | ~v_110;
assign x_4029 = v_2402 | ~v_103;
assign x_4030 = v_2402 | ~v_102;
assign x_4031 = v_2402 | ~v_100;
assign x_4032 = v_2402 | ~v_51;
assign x_4033 = v_2402 | ~v_49;
assign x_4034 = v_2402 | ~v_48;
assign x_4035 = v_2402 | ~v_46;
assign x_4036 = v_2402 | ~v_45;
assign x_4037 = v_2401 | ~v_646;
assign x_4038 = v_2401 | ~v_2279;
assign x_4039 = v_2401 | ~v_2340;
assign x_4040 = v_2401 | ~v_2341;
assign x_4041 = v_2401 | ~v_703;
assign x_4042 = v_2401 | ~v_704;
assign x_4043 = v_2401 | ~v_2280;
assign x_4044 = v_2401 | ~v_2281;
assign x_4045 = v_2401 | ~v_705;
assign x_4046 = v_2401 | ~v_706;
assign x_4047 = v_2401 | ~v_2282;
assign x_4048 = v_2401 | ~v_2283;
assign x_4049 = v_2401 | ~v_661;
assign x_4050 = v_2401 | ~v_2342;
assign x_4051 = v_2401 | ~v_711;
assign x_4052 = v_2401 | ~v_712;
assign x_4053 = v_2401 | ~v_2343;
assign x_4054 = v_2401 | ~v_2286;
assign x_4055 = v_2401 | ~v_108;
assign x_4056 = v_2401 | ~v_96;
assign x_4057 = v_2401 | ~v_95;
assign x_4058 = v_2401 | ~v_93;
assign x_4059 = v_2401 | ~v_25;
assign x_4060 = v_2401 | ~v_23;
assign x_4061 = v_2401 | ~v_22;
assign x_4062 = v_2401 | ~v_20;
assign x_4063 = v_2401 | ~v_19;
assign x_4064 = v_2400 | ~v_2399;
assign x_4065 = v_2400 | ~v_2376;
assign x_4066 = v_2400 | ~v_698;
assign x_4067 = v_2400 | ~v_699;
assign x_4068 = v_2400 | ~v_700;
assign x_4069 = v_2400 | ~v_701;
assign x_4070 = ~v_2398 | ~v_2397 | ~v_2396 | v_2399;
assign x_4071 = v_2398 | ~v_852;
assign x_4072 = v_2398 | ~v_853;
assign x_4073 = v_2398 | ~v_2301;
assign x_4074 = v_2398 | ~v_2302;
assign x_4075 = v_2398 | ~v_726;
assign x_4076 = v_2398 | ~v_2303;
assign x_4077 = v_2398 | ~v_2304;
assign x_4078 = v_2398 | ~v_2389;
assign x_4079 = v_2398 | ~v_2390;
assign x_4080 = v_2398 | ~v_634;
assign x_4081 = v_2398 | ~v_635;
assign x_4082 = v_2398 | ~v_854;
assign x_4083 = v_2398 | ~v_855;
assign x_4084 = v_2398 | ~v_2305;
assign x_4085 = v_2398 | ~v_731;
assign x_4086 = v_2398 | ~v_2391;
assign x_4087 = v_2398 | ~v_2392;
assign x_4088 = v_2398 | ~v_2307;
assign x_4089 = v_2398 | ~v_127;
assign x_4090 = v_2398 | ~v_112;
assign x_4091 = v_2398 | ~v_106;
assign x_4092 = v_2398 | ~v_105;
assign x_4093 = v_2398 | ~v_104;
assign x_4094 = v_2398 | ~v_76;
assign x_4095 = v_2398 | ~v_75;
assign x_4096 = v_2398 | ~v_73;
assign x_4097 = v_2398 | ~v_71;
assign x_4098 = v_2397 | ~v_847;
assign x_4099 = v_2397 | ~v_848;
assign x_4100 = v_2397 | ~v_2290;
assign x_4101 = v_2397 | ~v_2291;
assign x_4102 = v_2397 | ~v_714;
assign x_4103 = v_2397 | ~v_2384;
assign x_4104 = v_2397 | ~v_2385;
assign x_4105 = v_2397 | ~v_615;
assign x_4106 = v_2397 | ~v_616;
assign x_4107 = v_2397 | ~v_849;
assign x_4108 = v_2397 | ~v_850;
assign x_4109 = v_2397 | ~v_2292;
assign x_4110 = v_2397 | ~v_2293;
assign x_4111 = v_2397 | ~v_2386;
assign x_4112 = v_2397 | ~v_2387;
assign x_4113 = v_2397 | ~v_721;
assign x_4114 = v_2397 | ~v_2295;
assign x_4115 = v_2397 | ~v_2296;
assign x_4116 = v_2397 | ~v_126;
assign x_4117 = v_2397 | ~v_110;
assign x_4118 = v_2397 | ~v_102;
assign x_4119 = v_2397 | ~v_101;
assign x_4120 = v_2397 | ~v_100;
assign x_4121 = v_2397 | ~v_51;
assign x_4122 = v_2397 | ~v_50;
assign x_4123 = v_2397 | ~v_48;
assign x_4124 = v_2397 | ~v_46;
assign x_4125 = v_2396 | ~v_842;
assign x_4126 = v_2396 | ~v_843;
assign x_4127 = v_2396 | ~v_2279;
assign x_4128 = v_2396 | ~v_2280;
assign x_4129 = v_2396 | ~v_2281;
assign x_4130 = v_2396 | ~v_705;
assign x_4131 = v_2396 | ~v_706;
assign x_4132 = v_2396 | ~v_2379;
assign x_4133 = v_2396 | ~v_2380;
assign x_4134 = v_2396 | ~v_596;
assign x_4135 = v_2396 | ~v_597;
assign x_4136 = v_2396 | ~v_844;
assign x_4137 = v_2396 | ~v_845;
assign x_4138 = v_2396 | ~v_2282;
assign x_4139 = v_2396 | ~v_2283;
assign x_4140 = v_2396 | ~v_2381;
assign x_4141 = v_2396 | ~v_2382;
assign x_4142 = v_2396 | ~v_122;
assign x_4143 = v_2396 | ~v_2286;
assign x_4144 = v_2396 | ~v_108;
assign x_4145 = v_2396 | ~v_95;
assign x_4146 = v_2396 | ~v_94;
assign x_4147 = v_2396 | ~v_93;
assign x_4148 = v_2396 | ~v_25;
assign x_4149 = v_2396 | ~v_24;
assign x_4150 = v_2396 | ~v_22;
assign x_4151 = v_2396 | ~v_20;
assign x_4152 = v_2395 | ~v_2378;
assign x_4153 = v_2395 | ~v_2394;
assign x_4154 = v_2395 | ~v_698;
assign x_4155 = v_2395 | ~v_699;
assign x_4156 = v_2395 | ~v_700;
assign x_4157 = v_2395 | ~v_701;
assign x_4158 = ~v_2393 | ~v_2388 | ~v_2383 | v_2394;
assign x_4159 = v_2393 | ~v_951;
assign x_4160 = v_2393 | ~v_952;
assign x_4161 = v_2393 | ~v_906;
assign x_4162 = v_2393 | ~v_907;
assign x_4163 = v_2393 | ~v_2301;
assign x_4164 = v_2393 | ~v_2302;
assign x_4165 = v_2393 | ~v_2366;
assign x_4166 = v_2393 | ~v_2367;
assign x_4167 = v_2393 | ~v_953;
assign x_4168 = v_2393 | ~v_954;
assign x_4169 = v_2393 | ~v_2389;
assign x_4170 = v_2393 | ~v_2390;
assign x_4171 = v_2393 | ~v_634;
assign x_4172 = v_2393 | ~v_635;
assign x_4173 = v_2393 | ~v_2368;
assign x_4174 = v_2393 | ~v_2391;
assign x_4175 = v_2393 | ~v_2392;
assign x_4176 = v_2393 | ~v_2369;
assign x_4177 = v_2393 | ~v_127;
assign x_4178 = v_2393 | ~v_113;
assign x_4179 = v_2393 | ~v_106;
assign x_4180 = v_2393 | ~v_105;
assign x_4181 = v_2393 | ~v_104;
assign x_4182 = v_2393 | ~v_76;
assign x_4183 = v_2393 | ~v_75;
assign x_4184 = v_2393 | ~v_73;
assign x_4185 = v_2393 | ~v_68;
assign x_4186 = ~v_87 | ~v_130 | v_2392;
assign x_4187 = ~v_79 | v_130 | v_2391;
assign x_4188 = ~v_90 | ~v_129 | v_2390;
assign x_4189 = ~v_82 | v_129 | v_2389;
assign x_4190 = v_2388 | ~v_946;
assign x_4191 = v_2388 | ~v_947;
assign x_4192 = v_2388 | ~v_2290;
assign x_4193 = v_2388 | ~v_2291;
assign x_4194 = v_2388 | ~v_948;
assign x_4195 = v_2388 | ~v_949;
assign x_4196 = v_2388 | ~v_2384;
assign x_4197 = v_2388 | ~v_2385;
assign x_4198 = v_2388 | ~v_615;
assign x_4199 = v_2388 | ~v_616;
assign x_4200 = v_2388 | ~v_2361;
assign x_4201 = v_2388 | ~v_2362;
assign x_4202 = v_2388 | ~v_2386;
assign x_4203 = v_2388 | ~v_2387;
assign x_4204 = v_2388 | ~v_900;
assign x_4205 = v_2388 | ~v_2363;
assign x_4206 = v_2388 | ~v_2364;
assign x_4207 = v_2388 | ~v_902;
assign x_4208 = v_2388 | ~v_126;
assign x_4209 = v_2388 | ~v_111;
assign x_4210 = v_2388 | ~v_102;
assign x_4211 = v_2388 | ~v_101;
assign x_4212 = v_2388 | ~v_100;
assign x_4213 = v_2388 | ~v_51;
assign x_4214 = v_2388 | ~v_50;
assign x_4215 = v_2388 | ~v_48;
assign x_4216 = v_2388 | ~v_43;
assign x_4217 = ~v_62 | ~v_130 | v_2387;
assign x_4218 = ~v_54 | v_130 | v_2386;
assign x_4219 = ~v_65 | ~v_129 | v_2385;
assign x_4220 = ~v_57 | v_129 | v_2384;
assign x_4221 = v_2383 | ~v_941;
assign x_4222 = v_2383 | ~v_942;
assign x_4223 = v_2383 | ~v_885;
assign x_4224 = v_2383 | ~v_2279;
assign x_4225 = v_2383 | ~v_2356;
assign x_4226 = v_2383 | ~v_2357;
assign x_4227 = v_2383 | ~v_2358;
assign x_4228 = v_2383 | ~v_943;
assign x_4229 = v_2383 | ~v_944;
assign x_4230 = v_2383 | ~v_2379;
assign x_4231 = v_2383 | ~v_2380;
assign x_4232 = v_2383 | ~v_596;
assign x_4233 = v_2383 | ~v_597;
assign x_4234 = v_2383 | ~v_2359;
assign x_4235 = v_2383 | ~v_2282;
assign x_4236 = v_2383 | ~v_2381;
assign x_4237 = v_2383 | ~v_2382;
assign x_4238 = v_2383 | ~v_890;
assign x_4239 = v_2383 | ~v_122;
assign x_4240 = v_2383 | ~v_109;
assign x_4241 = v_2383 | ~v_95;
assign x_4242 = v_2383 | ~v_94;
assign x_4243 = v_2383 | ~v_93;
assign x_4244 = v_2383 | ~v_25;
assign x_4245 = v_2383 | ~v_24;
assign x_4246 = v_2383 | ~v_22;
assign x_4247 = v_2383 | ~v_17;
assign x_4248 = ~v_37 | ~v_130 | v_2382;
assign x_4249 = ~v_29 | v_130 | v_2381;
assign x_4250 = ~v_40 | ~v_129 | v_2380;
assign x_4251 = ~v_32 | v_129 | v_2379;
assign x_4252 = ~v_2377 | ~v_2372 | ~v_2339 | v_2378;
assign x_4253 = v_2377 | ~v_2376;
assign x_4254 = v_2377 | ~v_698;
assign x_4255 = v_2377 | ~v_699;
assign x_4256 = v_2377 | ~v_700;
assign x_4257 = v_2377 | ~v_701;
assign x_4258 = ~v_2375 | ~v_2374 | ~v_2373 | v_2376;
assign x_4259 = v_2375 | ~v_812;
assign x_4260 = v_2375 | ~v_813;
assign x_4261 = v_2375 | ~v_814;
assign x_4262 = v_2375 | ~v_815;
assign x_4263 = v_2375 | ~v_2299;
assign x_4264 = v_2375 | ~v_2300;
assign x_4265 = v_2375 | ~v_2301;
assign x_4266 = v_2375 | ~v_2302;
assign x_4267 = v_2375 | ~v_816;
assign x_4268 = v_2375 | ~v_817;
assign x_4269 = v_2375 | ~v_2331;
assign x_4270 = v_2375 | ~v_2332;
assign x_4271 = v_2375 | ~v_688;
assign x_4272 = v_2375 | ~v_689;
assign x_4273 = v_2375 | ~v_2334;
assign x_4274 = v_2375 | ~v_2335;
assign x_4275 = v_2375 | ~v_2306;
assign x_4276 = v_2375 | ~v_2308;
assign x_4277 = v_2375 | ~v_132;
assign x_4278 = v_2375 | ~v_121;
assign x_4279 = v_2375 | ~v_113;
assign x_4280 = v_2375 | ~v_112;
assign x_4281 = v_2375 | ~v_106;
assign x_4282 = v_2375 | ~v_105;
assign x_4283 = v_2375 | ~v_104;
assign x_4284 = v_2375 | ~v_75;
assign x_4285 = v_2375 | ~v_74;
assign x_4286 = v_2374 | ~v_801;
assign x_4287 = v_2374 | ~v_802;
assign x_4288 = v_2374 | ~v_803;
assign x_4289 = v_2374 | ~v_804;
assign x_4290 = v_2374 | ~v_2288;
assign x_4291 = v_2374 | ~v_2289;
assign x_4292 = v_2374 | ~v_2290;
assign x_4293 = v_2374 | ~v_2291;
assign x_4294 = v_2374 | ~v_805;
assign x_4295 = v_2374 | ~v_806;
assign x_4296 = v_2374 | ~v_2320;
assign x_4297 = v_2374 | ~v_2321;
assign x_4298 = v_2374 | ~v_669;
assign x_4299 = v_2374 | ~v_670;
assign x_4300 = v_2374 | ~v_2324;
assign x_4301 = v_2374 | ~v_2325;
assign x_4302 = v_2374 | ~v_2294;
assign x_4303 = v_2374 | ~v_2297;
assign x_4304 = v_2374 | ~v_131;
assign x_4305 = v_2374 | ~v_120;
assign x_4306 = v_2374 | ~v_111;
assign x_4307 = v_2374 | ~v_110;
assign x_4308 = v_2374 | ~v_102;
assign x_4309 = v_2374 | ~v_101;
assign x_4310 = v_2374 | ~v_100;
assign x_4311 = v_2374 | ~v_50;
assign x_4312 = v_2374 | ~v_49;
assign x_4313 = v_2373 | ~v_790;
assign x_4314 = v_2373 | ~v_791;
assign x_4315 = v_2373 | ~v_792;
assign x_4316 = v_2373 | ~v_793;
assign x_4317 = v_2373 | ~v_2277;
assign x_4318 = v_2373 | ~v_2278;
assign x_4319 = v_2373 | ~v_2279;
assign x_4320 = v_2373 | ~v_794;
assign x_4321 = v_2373 | ~v_795;
assign x_4322 = v_2373 | ~v_2312;
assign x_4323 = v_2373 | ~v_2313;
assign x_4324 = v_2373 | ~v_653;
assign x_4325 = v_2373 | ~v_654;
assign x_4326 = v_2373 | ~v_2282;
assign x_4327 = v_2373 | ~v_2314;
assign x_4328 = v_2373 | ~v_2315;
assign x_4329 = v_2373 | ~v_2284;
assign x_4330 = v_2373 | ~v_2285;
assign x_4331 = v_2373 | ~v_128;
assign x_4332 = v_2373 | ~v_117;
assign x_4333 = v_2373 | ~v_109;
assign x_4334 = v_2373 | ~v_108;
assign x_4335 = v_2373 | ~v_95;
assign x_4336 = v_2373 | ~v_94;
assign x_4337 = v_2373 | ~v_93;
assign x_4338 = v_2373 | ~v_24;
assign x_4339 = v_2373 | ~v_23;
assign x_4340 = v_2372 | ~v_2355;
assign x_4341 = v_2372 | ~v_2371;
assign x_4342 = v_2372 | ~v_698;
assign x_4343 = v_2372 | ~v_699;
assign x_4344 = v_2372 | ~v_700;
assign x_4345 = v_2372 | ~v_701;
assign x_4346 = ~v_2370 | ~v_2365 | ~v_2360 | v_2371;
assign x_4347 = v_2370 | ~v_814;
assign x_4348 = v_2370 | ~v_815;
assign x_4349 = v_2370 | ~v_2299;
assign x_4350 = v_2370 | ~v_2300;
assign x_4351 = v_2370 | ~v_930;
assign x_4352 = v_2370 | ~v_931;
assign x_4353 = v_2370 | ~v_932;
assign x_4354 = v_2370 | ~v_933;
assign x_4355 = v_2370 | ~v_906;
assign x_4356 = v_2370 | ~v_907;
assign x_4357 = v_2370 | ~v_2301;
assign x_4358 = v_2370 | ~v_2302;
assign x_4359 = v_2370 | ~v_2366;
assign x_4360 = v_2370 | ~v_2367;
assign x_4361 = v_2370 | ~v_2368;
assign x_4362 = v_2370 | ~v_2306;
assign x_4363 = v_2370 | ~v_2369;
assign x_4364 = v_2370 | ~v_2308;
assign x_4365 = v_2370 | ~v_113;
assign x_4366 = v_2370 | ~v_107;
assign x_4367 = v_2370 | ~v_106;
assign x_4368 = v_2370 | ~v_105;
assign x_4369 = v_2370 | ~v_104;
assign x_4370 = v_2370 | ~v_76;
assign x_4371 = v_2370 | ~v_74;
assign x_4372 = v_2370 | ~v_73;
assign x_4373 = v_2370 | ~v_68;
assign x_4374 = ~v_88 | ~v_99 | v_2369;
assign x_4375 = ~v_80 | v_99 | v_2368;
assign x_4376 = ~v_86 | ~v_99 | v_2367;
assign x_4377 = ~v_78 | v_99 | v_2366;
assign x_4378 = v_2365 | ~v_803;
assign x_4379 = v_2365 | ~v_804;
assign x_4380 = v_2365 | ~v_2288;
assign x_4381 = v_2365 | ~v_2289;
assign x_4382 = v_2365 | ~v_925;
assign x_4383 = v_2365 | ~v_926;
assign x_4384 = v_2365 | ~v_2290;
assign x_4385 = v_2365 | ~v_2291;
assign x_4386 = v_2365 | ~v_927;
assign x_4387 = v_2365 | ~v_928;
assign x_4388 = v_2365 | ~v_2361;
assign x_4389 = v_2365 | ~v_2362;
assign x_4390 = v_2365 | ~v_2294;
assign x_4391 = v_2365 | ~v_900;
assign x_4392 = v_2365 | ~v_2363;
assign x_4393 = v_2365 | ~v_2364;
assign x_4394 = v_2365 | ~v_902;
assign x_4395 = v_2365 | ~v_2297;
assign x_4396 = v_2365 | ~v_111;
assign x_4397 = v_2365 | ~v_103;
assign x_4398 = v_2365 | ~v_102;
assign x_4399 = v_2365 | ~v_101;
assign x_4400 = v_2365 | ~v_100;
assign x_4401 = v_2365 | ~v_51;
assign x_4402 = v_2365 | ~v_49;
assign x_4403 = v_2365 | ~v_48;
assign x_4404 = v_2365 | ~v_43;
assign x_4405 = ~v_55 | v_99 | v_2364;
assign x_4406 = ~v_63 | ~v_99 | v_2363;
assign x_4407 = ~v_53 | v_99 | v_2362;
assign x_4408 = ~v_61 | ~v_99 | v_2361;
assign x_4409 = v_2360 | ~v_792;
assign x_4410 = v_2360 | ~v_793;
assign x_4411 = v_2360 | ~v_2277;
assign x_4412 = v_2360 | ~v_2278;
assign x_4413 = v_2360 | ~v_920;
assign x_4414 = v_2360 | ~v_921;
assign x_4415 = v_2360 | ~v_885;
assign x_4416 = v_2360 | ~v_2279;
assign x_4417 = v_2360 | ~v_2356;
assign x_4418 = v_2360 | ~v_2357;
assign x_4419 = v_2360 | ~v_2358;
assign x_4420 = v_2360 | ~v_922;
assign x_4421 = v_2360 | ~v_2359;
assign x_4422 = v_2360 | ~v_2282;
assign x_4423 = v_2360 | ~v_2284;
assign x_4424 = v_2360 | ~v_2285;
assign x_4425 = v_2360 | ~v_890;
assign x_4426 = v_2360 | ~v_923;
assign x_4427 = v_2360 | ~v_109;
assign x_4428 = v_2360 | ~v_96;
assign x_4429 = v_2360 | ~v_95;
assign x_4430 = v_2360 | ~v_94;
assign x_4431 = v_2360 | ~v_93;
assign x_4432 = v_2360 | ~v_25;
assign x_4433 = v_2360 | ~v_23;
assign x_4434 = v_2360 | ~v_22;
assign x_4435 = v_2360 | ~v_17;
assign x_4436 = ~v_36 | ~v_99 | v_2359;
assign x_4437 = ~v_38 | ~v_99 | v_2358;
assign x_4438 = ~v_30 | v_99 | v_2357;
assign x_4439 = ~v_28 | v_99 | v_2356;
assign x_4440 = ~v_2354 | ~v_2349 | ~v_2344 | v_2355;
assign x_4441 = v_2354 | ~v_680;
assign x_4442 = v_2354 | ~v_681;
assign x_4443 = v_2354 | ~v_682;
assign x_4444 = v_2354 | ~v_683;
assign x_4445 = v_2354 | ~v_2301;
assign x_4446 = v_2354 | ~v_2302;
assign x_4447 = v_2354 | ~v_2350;
assign x_4448 = v_2354 | ~v_2351;
assign x_4449 = v_2354 | ~v_2352;
assign x_4450 = v_2354 | ~v_686;
assign x_4451 = v_2354 | ~v_687;
assign x_4452 = v_2354 | ~v_2331;
assign x_4453 = v_2354 | ~v_2332;
assign x_4454 = v_2354 | ~v_688;
assign x_4455 = v_2354 | ~v_689;
assign x_4456 = v_2354 | ~v_2353;
assign x_4457 = v_2354 | ~v_2334;
assign x_4458 = v_2354 | ~v_2335;
assign x_4459 = v_2354 | ~v_132;
assign x_4460 = v_2354 | ~v_113;
assign x_4461 = v_2354 | ~v_112;
assign x_4462 = v_2354 | ~v_106;
assign x_4463 = v_2354 | ~v_104;
assign x_4464 = v_2354 | ~v_76;
assign x_4465 = v_2354 | ~v_75;
assign x_4466 = v_2354 | ~v_74;
assign x_4467 = v_2354 | ~v_70;
assign x_4468 = ~v_79 | v_99 | v_2353;
assign x_4469 = ~v_90 | ~v_99 | v_2352;
assign x_4470 = ~v_82 | v_99 | v_2351;
assign x_4471 = ~v_87 | ~v_99 | v_2350;
assign x_4472 = v_2349 | ~v_2290;
assign x_4473 = v_2349 | ~v_2291;
assign x_4474 = v_2349 | ~v_665;
assign x_4475 = v_2349 | ~v_666;
assign x_4476 = v_2349 | ~v_2320;
assign x_4477 = v_2349 | ~v_2321;
assign x_4478 = v_2349 | ~v_667;
assign x_4479 = v_2349 | ~v_668;
assign x_4480 = v_2349 | ~v_669;
assign x_4481 = v_2349 | ~v_670;
assign x_4482 = v_2349 | ~v_2345;
assign x_4483 = v_2349 | ~v_2346;
assign x_4484 = v_2349 | ~v_2324;
assign x_4485 = v_2349 | ~v_2325;
assign x_4486 = v_2349 | ~v_2347;
assign x_4487 = v_2349 | ~v_2348;
assign x_4488 = v_2349 | ~v_677;
assign x_4489 = v_2349 | ~v_678;
assign x_4490 = v_2349 | ~v_131;
assign x_4491 = v_2349 | ~v_111;
assign x_4492 = v_2349 | ~v_110;
assign x_4493 = v_2349 | ~v_102;
assign x_4494 = v_2349 | ~v_100;
assign x_4495 = v_2349 | ~v_51;
assign x_4496 = v_2349 | ~v_50;
assign x_4497 = v_2349 | ~v_49;
assign x_4498 = v_2349 | ~v_45;
assign x_4499 = ~v_54 | v_99 | v_2348;
assign x_4500 = ~v_65 | ~v_99 | v_2347;
assign x_4501 = ~v_57 | v_99 | v_2346;
assign x_4502 = ~v_62 | ~v_99 | v_2345;
assign x_4503 = v_2344 | ~v_646;
assign x_4504 = v_2344 | ~v_2279;
assign x_4505 = v_2344 | ~v_2340;
assign x_4506 = v_2344 | ~v_2341;
assign x_4507 = v_2344 | ~v_649;
assign x_4508 = v_2344 | ~v_650;
assign x_4509 = v_2344 | ~v_2312;
assign x_4510 = v_2344 | ~v_2313;
assign x_4511 = v_2344 | ~v_651;
assign x_4512 = v_2344 | ~v_652;
assign x_4513 = v_2344 | ~v_653;
assign x_4514 = v_2344 | ~v_654;
assign x_4515 = v_2344 | ~v_2282;
assign x_4516 = v_2344 | ~v_2314;
assign x_4517 = v_2344 | ~v_2315;
assign x_4518 = v_2344 | ~v_661;
assign x_4519 = v_2344 | ~v_2342;
assign x_4520 = v_2344 | ~v_2343;
assign x_4521 = v_2344 | ~v_128;
assign x_4522 = v_2344 | ~v_109;
assign x_4523 = v_2344 | ~v_108;
assign x_4524 = v_2344 | ~v_95;
assign x_4525 = v_2344 | ~v_93;
assign x_4526 = v_2344 | ~v_25;
assign x_4527 = v_2344 | ~v_24;
assign x_4528 = v_2344 | ~v_23;
assign x_4529 = v_2344 | ~v_19;
assign x_4530 = ~v_32 | v_99 | v_2343;
assign x_4531 = ~v_40 | ~v_99 | v_2342;
assign x_4532 = ~v_37 | ~v_99 | v_2341;
assign x_4533 = ~v_29 | v_99 | v_2340;
assign x_4534 = v_2339 | ~v_2310;
assign x_4535 = v_2339 | ~v_2338;
assign x_4536 = v_2339 | ~v_698;
assign x_4537 = v_2339 | ~v_699;
assign x_4538 = v_2339 | ~v_700;
assign x_4539 = v_2339 | ~v_701;
assign x_4540 = ~v_2337 | ~v_2328 | ~v_2319 | v_2338;
assign x_4541 = v_2337 | ~v_871;
assign x_4542 = v_2337 | ~v_872;
assign x_4543 = v_2337 | ~v_873;
assign x_4544 = v_2337 | ~v_874;
assign x_4545 = v_2337 | ~v_2301;
assign x_4546 = v_2337 | ~v_2302;
assign x_4547 = v_2337 | ~v_763;
assign x_4548 = v_2337 | ~v_764;
assign x_4549 = v_2337 | ~v_2329;
assign x_4550 = v_2337 | ~v_2330;
assign x_4551 = v_2337 | ~v_2331;
assign x_4552 = v_2337 | ~v_2332;
assign x_4553 = v_2337 | ~v_688;
assign x_4554 = v_2337 | ~v_689;
assign x_4555 = v_2337 | ~v_2333;
assign x_4556 = v_2337 | ~v_2334;
assign x_4557 = v_2337 | ~v_2335;
assign x_4558 = v_2337 | ~v_2336;
assign x_4559 = v_2337 | ~v_132;
assign x_4560 = v_2337 | ~v_113;
assign x_4561 = v_2337 | ~v_112;
assign x_4562 = v_2337 | ~v_105;
assign x_4563 = v_2337 | ~v_104;
assign x_4564 = v_2337 | ~v_76;
assign x_4565 = v_2337 | ~v_75;
assign x_4566 = v_2337 | ~v_74;
assign x_4567 = v_2337 | ~v_72;
assign x_4568 = ~v_87 | ~v_98 | v_2336;
assign x_4569 = ~v_86 | ~v_130 | v_2335;
assign x_4570 = ~v_78 | v_130 | v_2334;
assign x_4571 = ~v_79 | v_98 | v_2333;
assign x_4572 = ~v_88 | ~v_129 | v_2332;
assign x_4573 = ~v_80 | v_129 | v_2331;
assign x_4574 = ~v_90 | ~v_97 | v_2330;
assign x_4575 = ~v_82 | v_97 | v_2329;
assign x_4576 = v_2328 | ~v_866;
assign x_4577 = v_2328 | ~v_867;
assign x_4578 = v_2328 | ~v_2290;
assign x_4579 = v_2328 | ~v_2291;
assign x_4580 = v_2328 | ~v_750;
assign x_4581 = v_2328 | ~v_2320;
assign x_4582 = v_2328 | ~v_2321;
assign x_4583 = v_2328 | ~v_868;
assign x_4584 = v_2328 | ~v_669;
assign x_4585 = v_2328 | ~v_670;
assign x_4586 = v_2328 | ~v_869;
assign x_4587 = v_2328 | ~v_2322;
assign x_4588 = v_2328 | ~v_2323;
assign x_4589 = v_2328 | ~v_2324;
assign x_4590 = v_2328 | ~v_2325;
assign x_4591 = v_2328 | ~v_757;
assign x_4592 = v_2328 | ~v_2326;
assign x_4593 = v_2328 | ~v_2327;
assign x_4594 = v_2328 | ~v_131;
assign x_4595 = v_2328 | ~v_111;
assign x_4596 = v_2328 | ~v_110;
assign x_4597 = v_2328 | ~v_101;
assign x_4598 = v_2328 | ~v_100;
assign x_4599 = v_2328 | ~v_51;
assign x_4600 = v_2328 | ~v_50;
assign x_4601 = v_2328 | ~v_49;
assign x_4602 = v_2328 | ~v_47;
assign x_4603 = ~v_65 | ~v_97 | v_2327;
assign x_4604 = ~v_54 | v_98 | v_2326;
assign x_4605 = ~v_61 | ~v_130 | v_2325;
assign x_4606 = ~v_53 | v_130 | v_2324;
assign x_4607 = ~v_62 | ~v_98 | v_2323;
assign x_4608 = ~v_57 | v_97 | v_2322;
assign x_4609 = ~v_63 | ~v_129 | v_2321;
assign x_4610 = ~v_55 | v_129 | v_2320;
assign x_4611 = v_2319 | ~v_861;
assign x_4612 = v_2319 | ~v_862;
assign x_4613 = v_2319 | ~v_2279;
assign x_4614 = v_2319 | ~v_739;
assign x_4615 = v_2319 | ~v_2311;
assign x_4616 = v_2319 | ~v_2312;
assign x_4617 = v_2319 | ~v_2313;
assign x_4618 = v_2319 | ~v_653;
assign x_4619 = v_2319 | ~v_654;
assign x_4620 = v_2319 | ~v_863;
assign x_4621 = v_2319 | ~v_864;
assign x_4622 = v_2319 | ~v_2282;
assign x_4623 = v_2319 | ~v_2314;
assign x_4624 = v_2319 | ~v_2315;
assign x_4625 = v_2319 | ~v_746;
assign x_4626 = v_2319 | ~v_2316;
assign x_4627 = v_2319 | ~v_2317;
assign x_4628 = v_2319 | ~v_128;
assign x_4629 = v_2319 | ~v_2318;
assign x_4630 = v_2319 | ~v_109;
assign x_4631 = v_2319 | ~v_108;
assign x_4632 = v_2319 | ~v_94;
assign x_4633 = v_2319 | ~v_93;
assign x_4634 = v_2319 | ~v_25;
assign x_4635 = v_2319 | ~v_24;
assign x_4636 = v_2319 | ~v_23;
assign x_4637 = v_2319 | ~v_21;
assign x_4638 = ~v_29 | v_98 | v_2318;
assign x_4639 = ~v_32 | v_97 | v_2317;
assign x_4640 = ~v_40 | ~v_97 | v_2316;
assign x_4641 = ~v_36 | ~v_130 | v_2315;
assign x_4642 = ~v_28 | v_130 | v_2314;
assign x_4643 = ~v_38 | ~v_129 | v_2313;
assign x_4644 = ~v_30 | v_129 | v_2312;
assign x_4645 = ~v_37 | ~v_98 | v_2311;
assign x_4646 = ~v_2309 | ~v_2298 | ~v_2287 | v_2310;
assign x_4647 = v_2309 | ~v_835;
assign x_4648 = v_2309 | ~v_836;
assign x_4649 = v_2309 | ~v_814;
assign x_4650 = v_2309 | ~v_815;
assign x_4651 = v_2309 | ~v_2299;
assign x_4652 = v_2309 | ~v_2300;
assign x_4653 = v_2309 | ~v_837;
assign x_4654 = v_2309 | ~v_838;
assign x_4655 = v_2309 | ~v_2301;
assign x_4656 = v_2309 | ~v_2302;
assign x_4657 = v_2309 | ~v_726;
assign x_4658 = v_2309 | ~v_2303;
assign x_4659 = v_2309 | ~v_2304;
assign x_4660 = v_2309 | ~v_2305;
assign x_4661 = v_2309 | ~v_731;
assign x_4662 = v_2309 | ~v_2306;
assign x_4663 = v_2309 | ~v_2307;
assign x_4664 = v_2309 | ~v_2308;
assign x_4665 = v_2309 | ~v_112;
assign x_4666 = v_2309 | ~v_106;
assign x_4667 = v_2309 | ~v_105;
assign x_4668 = v_2309 | ~v_104;
assign x_4669 = v_2309 | ~v_76;
assign x_4670 = v_2309 | ~v_75;
assign x_4671 = v_2309 | ~v_74;
assign x_4672 = v_2309 | ~v_73;
assign x_4673 = v_2309 | ~v_71;
assign x_4674 = ~v_87 | ~v_119 | v_2308;
assign x_4675 = ~v_88 | ~v_97 | v_2307;
assign x_4676 = ~v_79 | v_119 | v_2306;
assign x_4677 = ~v_80 | v_97 | v_2305;
assign x_4678 = ~v_86 | ~v_98 | v_2304;
assign x_4679 = ~v_78 | v_98 | v_2303;
assign x_4680 = ~v_85 | ~v_99 | v_2302;
assign x_4681 = ~v_77 | v_99 | v_2301;
assign x_4682 = ~v_90 | ~v_118 | v_2300;
assign x_4683 = ~v_82 | v_118 | v_2299;
assign x_4684 = v_2298 | ~v_830;
assign x_4685 = v_2298 | ~v_831;
assign x_4686 = v_2298 | ~v_803;
assign x_4687 = v_2298 | ~v_804;
assign x_4688 = v_2298 | ~v_2288;
assign x_4689 = v_2298 | ~v_2289;
assign x_4690 = v_2298 | ~v_2290;
assign x_4691 = v_2298 | ~v_2291;
assign x_4692 = v_2298 | ~v_714;
assign x_4693 = v_2298 | ~v_832;
assign x_4694 = v_2298 | ~v_833;
assign x_4695 = v_2298 | ~v_2292;
assign x_4696 = v_2298 | ~v_2293;
assign x_4697 = v_2298 | ~v_2294;
assign x_4698 = v_2298 | ~v_721;
assign x_4699 = v_2298 | ~v_2295;
assign x_4700 = v_2298 | ~v_2296;
assign x_4701 = v_2298 | ~v_2297;
assign x_4702 = v_2298 | ~v_110;
assign x_4703 = v_2298 | ~v_102;
assign x_4704 = v_2298 | ~v_101;
assign x_4705 = v_2298 | ~v_100;
assign x_4706 = v_2298 | ~v_51;
assign x_4707 = v_2298 | ~v_50;
assign x_4708 = v_2298 | ~v_49;
assign x_4709 = v_2298 | ~v_48;
assign x_4710 = v_2298 | ~v_46;
assign x_4711 = ~v_62 | ~v_119 | v_2297;
assign x_4712 = ~v_55 | v_97 | v_2296;
assign x_4713 = ~v_63 | ~v_97 | v_2295;
assign x_4714 = ~v_54 | v_119 | v_2294;
assign x_4715 = ~v_53 | v_98 | v_2293;
assign x_4716 = ~v_61 | ~v_98 | v_2292;
assign x_4717 = ~v_60 | ~v_99 | v_2291;
assign x_4718 = ~v_52 | v_99 | v_2290;
assign x_4719 = ~v_65 | ~v_118 | v_2289;
assign x_4720 = ~v_57 | v_118 | v_2288;
assign x_4721 = v_2287 | ~v_825;
assign x_4722 = v_2287 | ~v_826;
assign x_4723 = v_2287 | ~v_792;
assign x_4724 = v_2287 | ~v_793;
assign x_4725 = v_2287 | ~v_2277;
assign x_4726 = v_2287 | ~v_2278;
assign x_4727 = v_2287 | ~v_2279;
assign x_4728 = v_2287 | ~v_2280;
assign x_4729 = v_2287 | ~v_2281;
assign x_4730 = v_2287 | ~v_705;
assign x_4731 = v_2287 | ~v_706;
assign x_4732 = v_2287 | ~v_827;
assign x_4733 = v_2287 | ~v_2282;
assign x_4734 = v_2287 | ~v_2283;
assign x_4735 = v_2287 | ~v_2284;
assign x_4736 = v_2287 | ~v_2285;
assign x_4737 = v_2287 | ~v_828;
assign x_4738 = v_2287 | ~v_2286;
assign x_4739 = v_2287 | ~v_108;
assign x_4740 = v_2287 | ~v_95;
assign x_4741 = v_2287 | ~v_94;
assign x_4742 = v_2287 | ~v_93;
assign x_4743 = v_2287 | ~v_25;
assign x_4744 = v_2287 | ~v_24;
assign x_4745 = v_2287 | ~v_23;
assign x_4746 = v_2287 | ~v_22;
assign x_4747 = v_2287 | ~v_20;
assign x_4748 = ~v_28 | v_98 | v_2286;
assign x_4749 = ~v_37 | ~v_119 | v_2285;
assign x_4750 = ~v_29 | v_119 | v_2284;
assign x_4751 = ~v_36 | ~v_98 | v_2283;
assign x_4752 = ~v_35 | ~v_99 | v_2282;
assign x_4753 = ~v_38 | ~v_97 | v_2281;
assign x_4754 = ~v_30 | v_97 | v_2280;
assign x_4755 = ~v_27 | v_99 | v_2279;
assign x_4756 = ~v_40 | ~v_118 | v_2278;
assign x_4757 = ~v_32 | v_118 | v_2277;
assign x_4758 = ~v_2275 | ~v_2267 | v_2276;
assign x_4759 = v_2275 | ~v_1592;
assign x_4760 = v_2275 | ~v_570;
assign x_4761 = v_2275 | ~v_2274;
assign x_4762 = v_2275 | ~v_99;
assign x_4763 = ~v_2273 | ~v_2270 | v_2274;
assign x_4764 = v_2273 | ~v_2271;
assign x_4765 = v_2273 | ~v_2272;
assign x_4766 = v_2273 | ~v_580;
assign x_4767 = v_2273 | ~v_581;
assign x_4768 = v_2273 | ~v_98;
assign x_4769 = ~v_119 | ~v_578 | v_2272;
assign x_4770 = ~v_130 | ~v_1596 | v_2271;
assign x_4771 = v_2270 | ~v_2268;
assign x_4772 = v_2270 | ~v_2269;
assign x_4773 = v_2270 | ~v_559;
assign x_4774 = v_2270 | ~v_560;
assign x_4775 = v_2270 | ~v_97;
assign x_4776 = ~v_114 | ~v_565 | v_2269;
assign x_4777 = ~v_123 | ~v_1588 | v_2268;
assign x_4778 = v_2267 | ~v_2245;
assign x_4779 = v_2267 | ~v_2264;
assign x_4780 = v_2267 | ~v_2265;
assign x_4781 = v_2267 | ~v_2190;
assign x_4782 = v_2267 | ~v_2195;
assign x_4783 = v_2267 | ~v_2266;
assign x_4784 = v_2267 | ~v_2196;
assign x_4785 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2194 | ~v_2247 | v_2266;
assign x_4786 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2189 | ~v_2168 | v_2265;
assign x_4787 = ~v_2263 | ~v_2249 | v_2264;
assign x_4788 = v_2263 | ~v_2250;
assign x_4789 = v_2263 | ~v_2251;
assign x_4790 = v_2263 | ~v_2256;
assign x_4791 = v_2263 | ~v_2261;
assign x_4792 = v_2263 | ~v_2262;
assign x_4793 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2189 | v_2262;
assign x_4794 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2260 | ~v_2194 | v_2261;
assign x_4795 = v_2260 | ~v_2257;
assign x_4796 = v_2260 | ~v_2258;
assign x_4797 = v_2260 | ~v_2259;
assign x_4798 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2184 | v_2259;
assign x_4799 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2201 | ~v_2189 | v_2258;
assign x_4800 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2161 | ~v_2222 | v_2257;
assign x_4801 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2255 | ~v_2100 | v_2256;
assign x_4802 = v_2255 | ~v_2252;
assign x_4803 = v_2255 | ~v_2253;
assign x_4804 = v_2255 | ~v_2254;
assign x_4805 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2222 | v_2254;
assign x_4806 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2227 | ~v_2189 | v_2253;
assign x_4807 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2184 | ~v_2232 | v_2252;
assign x_4808 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2184 | ~v_2194 | v_2251;
assign x_4809 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2222 | ~v_2100 | v_2250;
assign x_4810 = v_2249 | ~v_2246;
assign x_4811 = v_2249 | ~v_2248;
assign x_4812 = v_2249 | ~v_2129;
assign x_4813 = v_2249 | ~v_2162;
assign x_4814 = v_2249 | ~v_2167;
assign x_4815 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2145 | ~v_2247 | v_2248;
assign x_4816 = v_2247 | ~v_2203;
assign x_4817 = v_2247 | ~v_2204;
assign x_4818 = v_2247 | ~v_2205;
assign x_4819 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2128 | ~v_2197 | v_2246;
assign x_4820 = ~v_2244 | ~v_2206 | v_2245;
assign x_4821 = v_2244 | ~v_2235;
assign x_4822 = v_2244 | ~v_2240;
assign x_4823 = v_2244 | ~v_2241;
assign x_4824 = v_2244 | ~v_2242;
assign x_4825 = v_2244 | ~v_2243;
assign x_4826 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2194 | v_2243;
assign x_4827 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2145 | ~v_2189 | v_2242;
assign x_4828 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2232 | ~v_2100 | v_2241;
assign x_4829 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2189 | ~v_2239 | v_2240;
assign x_4830 = v_2239 | ~v_2236;
assign x_4831 = v_2239 | ~v_2237;
assign x_4832 = v_2239 | ~v_2238;
assign x_4833 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2145 | v_2238;
assign x_4834 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2128 | ~v_2194 | v_2237;
assign x_4835 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2166 | ~v_2232 | v_2236;
assign x_4836 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2100 | ~v_2234 | v_2235;
assign x_4837 = v_2234 | ~v_2223;
assign x_4838 = v_2234 | ~v_2228;
assign x_4839 = v_2234 | ~v_2233;
assign x_4840 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2232 | v_2233;
assign x_4841 = v_2232 | ~v_2229;
assign x_4842 = v_2232 | ~v_2230;
assign x_4843 = v_2232 | ~v_2231;
assign x_4844 = v_75 | v_74 | v_73 | v_70 | v_106 | v_104 | v_113 | v_112 | v_121 | ~v_2220 | ~v_2219 | ~v_2143 | ~v_332 | ~v_331 | ~v_180 | ~v_179 | ~v_2142 | ~v_2141 | ~v_2140 | ~v_2092 | ~v_2091 | ~v_230 | ~v_229 | ~v_330 | ~v_329 | ~v_2218 | ~v_2217 | v_2231;
assign x_4845 = v_50 | v_49 | v_48 | v_45 | v_100 | v_102 | v_111 | v_110 | v_120 | ~v_2215 | ~v_225 | ~v_224 | ~v_2138 | ~v_2137 | ~v_2214 | ~v_2136 | ~v_2135 | ~v_327 | ~v_326 | ~v_161 | ~v_160 | ~v_2081 | ~v_2080 | ~v_325 | ~v_324 | ~v_2213 | ~v_2212 | v_2230;
assign x_4846 = v_24 | v_23 | v_22 | v_19 | v_95 | v_93 | v_108 | v_109 | v_117 | ~v_2133 | ~v_2132 | ~v_208 | ~v_2210 | ~v_2209 | ~v_2073 | ~v_322 | ~v_321 | ~v_142 | ~v_141 | ~v_2131 | ~v_2130 | ~v_2069 | ~v_193 | ~v_320 | ~v_319 | ~v_2208 | ~v_2207 | v_2229;
assign x_4847 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2227 | ~v_2194 | v_2228;
assign x_4848 = v_2227 | ~v_2224;
assign x_4849 = v_2227 | ~v_2225;
assign x_4850 = v_2227 | ~v_2226;
assign x_4851 = v_76 | v_75 | v_74 | v_73 | v_72 | v_105 | v_104 | v_113 | v_112 | ~v_2126 | ~v_2220 | ~v_2219 | ~v_2123 | ~v_180 | ~v_179 | ~v_313 | ~v_312 | ~v_2120 | ~v_2119 | ~v_311 | ~v_310 | ~v_2092 | ~v_2091 | ~v_2218 | ~v_2217 | ~v_309 | ~v_308 | v_2226;
assign x_4852 = v_50 | v_51 | v_49 | v_48 | v_47 | v_101 | v_100 | v_111 | v_110 | ~v_2215 | ~v_2117 | ~v_2116 | ~v_304 | ~v_2214 | ~v_2113 | ~v_2112 | ~v_301 | ~v_300 | ~v_161 | ~v_160 | ~v_299 | ~v_298 | ~v_297 | ~v_2081 | ~v_2080 | ~v_2213 | ~v_2212 | v_2225;
assign x_4853 = v_25 | v_24 | v_23 | v_22 | v_21 | ~v_2108 | v_94 | v_93 | v_108 | v_109 | ~v_2107 | ~v_2106 | ~v_293 | ~v_2210 | ~v_2209 | ~v_2073 | ~v_290 | ~v_289 | ~v_142 | ~v_141 | ~v_288 | ~v_287 | ~v_2101 | ~v_286 | ~v_2069 | ~v_2208 | ~v_2207 | v_2224;
assign x_4854 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2145 | ~v_2222 | v_2223;
assign x_4855 = v_2222 | ~v_2211;
assign x_4856 = v_2222 | ~v_2216;
assign x_4857 = v_2222 | ~v_2221;
assign x_4858 = v_76 | v_73 | v_107 | v_106 | v_105 | v_104 | v_127 | v_113 | v_112 | ~v_2182 | ~v_2181 | ~v_2220 | ~v_2219 | ~v_184 | ~v_183 | ~v_182 | ~v_181 | ~v_2180 | ~v_2179 | ~v_180 | ~v_179 | ~v_2092 | ~v_2091 | ~v_2218 | ~v_2217 | ~v_178 | ~v_177 | v_2221;
assign x_4859 = v_2220 | v_119;
assign x_4860 = v_2220 | v_86;
assign x_4861 = v_2219 | ~v_119;
assign x_4862 = v_2219 | v_78;
assign x_4863 = v_2218 | v_118;
assign x_4864 = v_2218 | v_88;
assign x_4865 = v_2217 | ~v_118;
assign x_4866 = v_2217 | v_80;
assign x_4867 = v_51 | v_48 | v_103 | v_101 | v_100 | v_102 | v_111 | v_110 | v_126 | ~v_2215 | ~v_2177 | ~v_2176 | ~v_2214 | ~v_165 | ~v_164 | ~v_163 | ~v_162 | ~v_2175 | ~v_2174 | ~v_161 | ~v_160 | ~v_2081 | ~v_2080 | ~v_2213 | ~v_2212 | ~v_159 | ~v_158 | v_2216;
assign x_4868 = v_2215 | v_119;
assign x_4869 = v_2215 | v_61;
assign x_4870 = v_2214 | ~v_119;
assign x_4871 = v_2214 | v_53;
assign x_4872 = v_2213 | v_118;
assign x_4873 = v_2213 | v_63;
assign x_4874 = v_2212 | ~v_118;
assign x_4875 = v_2212 | v_55;
assign x_4876 = v_25 | v_22 | v_96 | v_95 | v_94 | v_93 | v_108 | v_109 | v_122 | ~v_2172 | ~v_2171 | ~v_2210 | ~v_2209 | ~v_2073 | ~v_146 | ~v_145 | ~v_144 | ~v_143 | ~v_2170 | ~v_2169 | ~v_142 | ~v_141 | ~v_2069 | ~v_2208 | ~v_2207 | ~v_140 | ~v_139 | v_2211;
assign x_4877 = v_2210 | v_119;
assign x_4878 = v_2210 | v_36;
assign x_4879 = v_2209 | ~v_119;
assign x_4880 = v_2209 | v_28;
assign x_4881 = v_2208 | v_118;
assign x_4882 = v_2208 | v_38;
assign x_4883 = v_2207 | ~v_118;
assign x_4884 = v_2207 | v_30;
assign x_4885 = v_2206 | ~v_2185;
assign x_4886 = v_2206 | ~v_2202;
assign x_4887 = v_2206 | ~v_2203;
assign x_4888 = v_2206 | ~v_2204;
assign x_4889 = v_2206 | ~v_2205;
assign x_4890 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2161 | v_2205;
assign x_4891 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2201 | ~v_2100 | v_2204;
assign x_4892 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2184 | ~v_2166 | v_2203;
assign x_4893 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2201 | ~v_2197 | v_2202;
assign x_4894 = v_2201 | ~v_2198;
assign x_4895 = v_2201 | ~v_2199;
assign x_4896 = v_2201 | ~v_2200;
assign x_4897 = v_68 | v_75 | v_74 | v_73 | v_72 | v_105 | v_104 | v_113 | v_121 | ~v_2126 | ~v_2159 | ~v_461 | ~v_2123 | ~v_2158 | ~v_2120 | ~v_2119 | ~v_311 | ~v_310 | ~v_457 | ~v_456 | ~v_455 | ~v_2157 | ~v_2156 | ~v_2092 | ~v_2091 | ~v_454 | ~v_453 | v_2200;
assign x_4898 = v_50 | v_49 | v_48 | v_43 | v_47 | v_101 | v_100 | v_111 | v_120 | ~v_450 | ~v_449 | ~v_2154 | ~v_448 | ~v_2117 | ~v_2116 | ~v_2153 | ~v_447 | ~v_304 | ~v_2152 | ~v_444 | ~v_2151 | ~v_2113 | ~v_2112 | ~v_297 | ~v_443 | ~v_2081 | ~v_2080 | v_2199;
assign x_4899 = v_24 | v_23 | v_22 | v_21 | v_17 | ~v_2108 | v_94 | v_93 | v_109 | v_117 | ~v_439 | ~v_2107 | ~v_438 | ~v_2106 | ~v_437 | ~v_293 | ~v_2073 | ~v_2149 | ~v_2101 | ~v_286 | ~v_434 | ~v_433 | ~v_2148 | ~v_2147 | ~v_2146 | ~v_2069 | ~v_432 | v_2198;
assign x_4900 = v_2197 | ~v_2190;
assign x_4901 = v_2197 | ~v_2195;
assign x_4902 = v_2197 | ~v_2196;
assign x_4903 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2100 | v_2196;
assign x_4904 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2161 | ~v_2194 | v_2195;
assign x_4905 = v_2194 | ~v_2191;
assign x_4906 = v_2194 | ~v_2192;
assign x_4907 = v_2194 | ~v_2193;
assign x_4908 = v_76 | v_74 | v_73 | v_71 | v_70 | v_107 | v_106 | v_104 | v_112 | ~v_2097 | ~v_281 | ~v_278 | ~v_2143 | ~v_2095 | ~v_2094 | ~v_2093 | ~v_275 | ~v_274 | ~v_273 | ~v_272 | ~v_2142 | ~v_2141 | ~v_2140 | ~v_2092 | ~v_2091 | ~v_230 | ~v_229 | v_2193;
assign x_4909 = v_51 | v_49 | v_48 | v_46 | v_45 | v_103 | v_100 | v_102 | v_110 | ~v_270 | ~v_2086 | ~v_225 | ~v_269 | ~v_224 | ~v_2085 | ~v_2138 | ~v_2137 | ~v_268 | ~v_2083 | ~v_265 | ~v_2136 | ~v_2082 | ~v_2135 | ~v_262 | ~v_261 | ~v_2081 | ~v_2080 | v_2192;
assign x_4910 = v_25 | v_23 | v_22 | v_20 | v_19 | v_96 | v_95 | ~v_2076 | v_93 | v_108 | ~v_2133 | ~v_259 | ~v_258 | ~v_2132 | ~v_208 | ~v_2073 | ~v_2072 | ~v_253 | ~v_252 | ~v_2071 | ~v_2070 | ~v_251 | ~v_250 | ~v_2131 | ~v_2130 | ~v_2069 | ~v_193 | v_2191;
assign x_4911 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2166 | ~v_2189 | v_2190;
assign x_4912 = v_2189 | ~v_2186;
assign x_4913 = v_2189 | ~v_2187;
assign x_4914 = v_2189 | ~v_2188;
assign x_4915 = v_76 | v_75 | v_73 | v_71 | v_106 | v_105 | v_104 | v_127 | v_112 | ~v_2097 | ~v_2182 | ~v_2181 | ~v_278 | ~v_2095 | ~v_402 | ~v_401 | ~v_182 | ~v_181 | ~v_2180 | ~v_2179 | ~v_2094 | ~v_2093 | ~v_273 | ~v_2092 | ~v_2091 | ~v_400 | ~v_399 | v_2188;
assign x_4916 = v_50 | v_51 | v_48 | v_46 | v_101 | v_100 | v_102 | v_110 | v_126 | ~v_2086 | ~v_2085 | ~v_268 | ~v_2177 | ~v_2176 | ~v_2083 | ~v_2082 | ~v_397 | ~v_396 | ~v_163 | ~v_162 | ~v_2175 | ~v_2174 | ~v_261 | ~v_2081 | ~v_2080 | ~v_395 | ~v_394 | v_2187;
assign x_4917 = v_25 | v_24 | v_22 | v_20 | v_95 | v_94 | ~v_2076 | v_93 | v_108 | v_122 | ~v_2172 | ~v_2171 | ~v_2073 | ~v_2072 | ~v_392 | ~v_391 | ~v_144 | ~v_143 | ~v_2170 | ~v_2169 | ~v_253 | ~v_252 | ~v_2071 | ~v_2070 | ~v_2069 | ~v_390 | ~v_389 | v_2186;
assign x_4918 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2184 | ~v_2168 | v_2185;
assign x_4919 = v_2184 | ~v_2173;
assign x_4920 = v_2184 | ~v_2178;
assign x_4921 = v_2184 | ~v_2183;
assign x_4922 = v_76 | v_68 | v_75 | v_73 | v_106 | v_105 | v_104 | v_127 | v_113 | ~v_2159 | ~v_2182 | ~v_2181 | ~v_2158 | ~v_182 | ~v_181 | ~v_2180 | ~v_2179 | ~v_501 | ~v_500 | ~v_2157 | ~v_2156 | ~v_2092 | ~v_2091 | ~v_454 | ~v_453 | ~v_499 | ~v_498 | v_2183;
assign x_4923 = v_2182 | v_130;
assign x_4924 = v_2182 | v_87;
assign x_4925 = v_2181 | ~v_130;
assign x_4926 = v_2181 | v_79;
assign x_4927 = v_2180 | v_129;
assign x_4928 = v_2180 | v_90;
assign x_4929 = v_2179 | ~v_129;
assign x_4930 = v_2179 | v_82;
assign x_4931 = v_50 | v_51 | v_48 | v_43 | v_101 | v_100 | v_102 | v_111 | v_126 | ~v_449 | ~v_2154 | ~v_2153 | ~v_447 | ~v_2177 | ~v_2176 | ~v_2152 | ~v_2151 | ~v_163 | ~v_162 | ~v_2175 | ~v_2174 | ~v_496 | ~v_495 | ~v_2081 | ~v_2080 | ~v_494 | ~v_493 | v_2178;
assign x_4932 = v_2177 | v_130;
assign x_4933 = v_2177 | v_62;
assign x_4934 = v_2176 | ~v_130;
assign x_4935 = v_2176 | v_54;
assign x_4936 = v_2175 | v_129;
assign x_4937 = v_2175 | v_65;
assign x_4938 = v_2174 | ~v_129;
assign x_4939 = v_2174 | v_57;
assign x_4940 = v_25 | v_24 | v_22 | v_17 | v_95 | v_94 | v_93 | v_109 | v_122 | ~v_437 | ~v_2172 | ~v_2171 | ~v_2073 | ~v_2149 | ~v_144 | ~v_143 | ~v_2170 | ~v_2169 | ~v_491 | ~v_490 | ~v_2148 | ~v_2147 | ~v_2146 | ~v_2069 | ~v_432 | ~v_489 | ~v_488 | v_2173;
assign x_4941 = v_2172 | v_130;
assign x_4942 = v_2172 | v_37;
assign x_4943 = v_2171 | ~v_130;
assign x_4944 = v_2171 | v_29;
assign x_4945 = v_2170 | v_129;
assign x_4946 = v_2170 | v_40;
assign x_4947 = v_2169 | ~v_129;
assign x_4948 = v_2169 | v_32;
assign x_4949 = v_2168 | ~v_2129;
assign x_4950 = v_2168 | ~v_2162;
assign x_4951 = v_2168 | ~v_2167;
assign x_4952 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2166 | v_2167;
assign x_4953 = v_2166 | ~v_2163;
assign x_4954 = v_2166 | ~v_2164;
assign x_4955 = v_2166 | ~v_2165;
assign x_4956 = v_75 | v_74 | v_106 | v_105 | v_104 | v_132 | v_113 | v_112 | v_121 | ~v_2098 | ~v_2096 | ~v_2125 | ~v_2124 | ~v_236 | ~v_235 | ~v_2122 | ~v_2121 | ~v_364 | ~v_363 | ~v_2092 | ~v_2091 | ~v_2090 | ~v_2089 | ~v_362 | ~v_361 | ~v_360 | ~v_359 | v_2165;
assign x_4957 = v_50 | v_49 | v_101 | v_100 | v_102 | v_111 | v_110 | v_131 | v_120 | ~v_2087 | ~v_2084 | ~v_2115 | ~v_2114 | ~v_217 | ~v_216 | ~v_2111 | ~v_2110 | ~v_353 | ~v_352 | ~v_2081 | ~v_2080 | ~v_2079 | ~v_2078 | ~v_351 | ~v_350 | ~v_349 | ~v_348 | v_2164;
assign x_4958 = v_24 | v_23 | v_95 | v_94 | v_93 | v_108 | v_109 | v_128 | v_117 | ~v_2075 | ~v_2074 | ~v_2105 | ~v_2104 | ~v_2073 | ~v_201 | ~v_200 | ~v_2103 | ~v_2102 | ~v_342 | ~v_341 | ~v_2069 | ~v_2068 | ~v_2067 | ~v_340 | ~v_339 | ~v_338 | ~v_337 | v_2163;
assign x_4959 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2161 | ~v_2145 | v_2162;
assign x_4960 = v_2161 | ~v_2150;
assign x_4961 = v_2161 | ~v_2155;
assign x_4962 = v_2161 | ~v_2160;
assign x_4963 = v_76 | v_68 | v_74 | v_73 | v_107 | v_106 | v_105 | v_104 | v_113 | ~v_2098 | ~v_2159 | ~v_2096 | ~v_2158 | ~v_2157 | ~v_2156 | ~v_2092 | ~v_2091 | ~v_454 | ~v_453 | ~v_480 | ~v_479 | ~v_478 | ~v_477 | ~v_2090 | ~v_2089 | ~v_362 | ~v_361 | v_2160;
assign x_4964 = v_2159 | v_99;
assign x_4965 = v_2159 | v_88;
assign x_4966 = v_2158 | ~v_99;
assign x_4967 = v_2158 | v_80;
assign x_4968 = v_2157 | v_99;
assign x_4969 = v_2157 | v_86;
assign x_4970 = v_2156 | ~v_99;
assign x_4971 = v_2156 | v_78;
assign x_4972 = v_51 | v_49 | v_48 | v_43 | v_103 | v_101 | v_100 | v_102 | v_111 | ~v_2087 | ~v_449 | ~v_2154 | ~v_2153 | ~v_447 | ~v_2084 | ~v_2152 | ~v_2151 | ~v_475 | ~v_474 | ~v_2081 | ~v_2080 | ~v_473 | ~v_472 | ~v_2079 | ~v_2078 | ~v_351 | ~v_350 | v_2155;
assign x_4973 = v_2154 | ~v_99;
assign x_4974 = v_2154 | v_55;
assign x_4975 = v_2153 | v_99;
assign x_4976 = v_2153 | v_63;
assign x_4977 = v_2152 | ~v_99;
assign x_4978 = v_2152 | v_53;
assign x_4979 = v_2151 | v_99;
assign x_4980 = v_2151 | v_61;
assign x_4981 = v_25 | v_23 | v_22 | v_17 | v_96 | v_95 | v_94 | v_93 | v_109 | ~v_470 | ~v_437 | ~v_2075 | ~v_2074 | ~v_2073 | ~v_2149 | ~v_469 | ~v_2148 | ~v_2147 | ~v_2146 | ~v_2069 | ~v_432 | ~v_468 | ~v_467 | ~v_2068 | ~v_2067 | ~v_340 | ~v_339 | v_2150;
assign x_4982 = v_2149 | v_99;
assign x_4983 = v_2149 | v_36;
assign x_4984 = v_2148 | v_99;
assign x_4985 = v_2148 | v_38;
assign x_4986 = v_2147 | ~v_99;
assign x_4987 = v_2147 | v_30;
assign x_4988 = v_2146 | ~v_99;
assign x_4989 = v_2146 | v_28;
assign x_4990 = v_2145 | ~v_2134;
assign x_4991 = v_2145 | ~v_2139;
assign x_4992 = v_2145 | ~v_2144;
assign x_4993 = v_76 | v_75 | v_74 | v_70 | v_106 | v_104 | v_132 | v_113 | v_112 | ~v_2125 | ~v_2124 | ~v_2143 | ~v_236 | ~v_235 | ~v_2122 | ~v_2121 | ~v_234 | ~v_233 | ~v_2142 | ~v_2141 | ~v_2140 | ~v_2092 | ~v_2091 | ~v_230 | ~v_229 | ~v_228 | ~v_227 | v_2144;
assign x_4994 = v_2143 | ~v_99;
assign x_4995 = v_2143 | v_79;
assign x_4996 = v_2142 | v_99;
assign x_4997 = v_2142 | v_90;
assign x_4998 = v_2141 | ~v_99;
assign x_4999 = v_2141 | v_82;
assign x_5000 = v_2140 | v_99;
assign x_5001 = v_2140 | v_87;
assign x_5002 = v_50 | v_51 | v_49 | v_45 | v_100 | v_102 | v_111 | v_110 | v_131 | ~v_225 | ~v_224 | ~v_2138 | ~v_2137 | ~v_2115 | ~v_2114 | ~v_2136 | ~v_2135 | ~v_217 | ~v_216 | ~v_215 | ~v_214 | ~v_2111 | ~v_2110 | ~v_213 | ~v_212 | ~v_2081 | ~v_2080 | v_2139;
assign x_5003 = v_2138 | ~v_99;
assign x_5004 = v_2138 | v_54;
assign x_5005 = v_2137 | v_99;
assign x_5006 = v_2137 | v_65;
assign x_5007 = v_2136 | ~v_99;
assign x_5008 = v_2136 | v_57;
assign x_5009 = v_2135 | v_99;
assign x_5010 = v_2135 | v_62;
assign x_5011 = v_25 | v_24 | v_23 | v_19 | v_95 | v_93 | v_108 | v_109 | v_128 | ~v_2133 | ~v_2132 | ~v_208 | ~v_2105 | ~v_2104 | ~v_2073 | ~v_201 | ~v_200 | ~v_199 | ~v_198 | ~v_2103 | ~v_2102 | ~v_197 | ~v_196 | ~v_2131 | ~v_2130 | ~v_2069 | ~v_193 | v_2134;
assign x_5012 = v_2133 | ~v_99;
assign x_5013 = v_2133 | v_32;
assign x_5014 = v_2132 | v_99;
assign x_5015 = v_2132 | v_40;
assign x_5016 = v_2131 | v_99;
assign x_5017 = v_2131 | v_37;
assign x_5018 = v_2130 | ~v_99;
assign x_5019 = v_2130 | v_29;
assign x_5020 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2128 | ~v_2100 | v_2129;
assign x_5021 = v_2128 | ~v_2109;
assign x_5022 = v_2128 | ~v_2118;
assign x_5023 = v_2128 | ~v_2127;
assign x_5024 = v_76 | v_75 | v_74 | v_72 | v_105 | v_104 | v_132 | v_113 | v_112 | ~v_2126 | ~v_2125 | ~v_2124 | ~v_2123 | ~v_236 | ~v_235 | ~v_2122 | ~v_2121 | ~v_2120 | ~v_2119 | ~v_311 | ~v_310 | ~v_2092 | ~v_2091 | ~v_421 | ~v_420 | ~v_419 | ~v_418 | v_2127;
assign x_5025 = v_2126 | v_87;
assign x_5026 = v_2126 | v_98;
assign x_5027 = v_2125 | v_130;
assign x_5028 = v_2125 | v_86;
assign x_5029 = v_2124 | ~v_130;
assign x_5030 = v_2124 | v_78;
assign x_5031 = v_2123 | ~v_98;
assign x_5032 = v_2123 | v_79;
assign x_5033 = v_2122 | v_129;
assign x_5034 = v_2122 | v_88;
assign x_5035 = v_2121 | ~v_129;
assign x_5036 = v_2121 | v_80;
assign x_5037 = v_2120 | v_97;
assign x_5038 = v_2120 | v_90;
assign x_5039 = v_2119 | ~v_97;
assign x_5040 = v_2119 | v_82;
assign x_5041 = v_50 | v_51 | v_49 | v_47 | v_101 | v_100 | v_111 | v_110 | v_131 | ~v_2117 | ~v_2116 | ~v_304 | ~v_2115 | ~v_2114 | ~v_2113 | ~v_2112 | ~v_416 | ~v_217 | ~v_216 | ~v_415 | ~v_2111 | ~v_2110 | ~v_297 | ~v_2081 | ~v_2080 | ~v_414 | ~v_413 | v_2118;
assign x_5042 = v_2117 | v_97;
assign x_5043 = v_2117 | v_65;
assign x_5044 = v_2116 | ~v_98;
assign x_5045 = v_2116 | v_54;
assign x_5046 = v_2115 | v_130;
assign x_5047 = v_2115 | v_61;
assign x_5048 = v_2114 | ~v_130;
assign x_5049 = v_2114 | v_53;
assign x_5050 = v_2113 | v_98;
assign x_5051 = v_2113 | v_62;
assign x_5052 = v_2112 | ~v_97;
assign x_5053 = v_2112 | v_57;
assign x_5054 = v_2111 | v_129;
assign x_5055 = v_2111 | v_63;
assign x_5056 = v_2110 | ~v_129;
assign x_5057 = v_2110 | v_55;
assign x_5058 = v_25 | v_24 | v_23 | v_21 | ~v_2108 | v_94 | v_93 | v_108 | v_109 | v_128 | ~v_2107 | ~v_2106 | ~v_293 | ~v_2105 | ~v_2104 | ~v_2073 | ~v_411 | ~v_410 | ~v_201 | ~v_200 | ~v_2103 | ~v_2102 | ~v_2101 | ~v_286 | ~v_2069 | ~v_409 | ~v_408 | v_2109;
assign x_5059 = v_2108 | ~v_98;
assign x_5060 = v_2108 | v_29;
assign x_5061 = v_2107 | ~v_97;
assign x_5062 = v_2107 | v_32;
assign x_5063 = v_2106 | v_97;
assign x_5064 = v_2106 | v_40;
assign x_5065 = v_2105 | v_130;
assign x_5066 = v_2105 | v_36;
assign x_5067 = v_2104 | ~v_130;
assign x_5068 = v_2104 | v_28;
assign x_5069 = v_2103 | v_129;
assign x_5070 = v_2103 | v_38;
assign x_5071 = v_2102 | ~v_129;
assign x_5072 = v_2102 | v_30;
assign x_5073 = v_2101 | v_98;
assign x_5074 = v_2101 | v_37;
assign x_5075 = v_2100 | ~v_2077;
assign x_5076 = v_2100 | ~v_2088;
assign x_5077 = v_2100 | ~v_2099;
assign x_5078 = v_76 | v_75 | v_74 | v_73 | v_71 | v_106 | v_105 | v_104 | v_112 | ~v_2098 | ~v_2097 | ~v_2096 | ~v_278 | ~v_2095 | ~v_2094 | ~v_2093 | ~v_273 | ~v_2092 | ~v_2091 | ~v_385 | ~v_384 | ~v_2090 | ~v_2089 | ~v_362 | ~v_361 | ~v_383 | ~v_382 | v_2099;
assign x_5079 = v_2098 | v_119;
assign x_5080 = v_2098 | v_87;
assign x_5081 = v_2097 | v_97;
assign x_5082 = v_2097 | v_88;
assign x_5083 = v_2096 | ~v_119;
assign x_5084 = v_2096 | v_79;
assign x_5085 = v_2095 | ~v_97;
assign x_5086 = v_2095 | v_80;
assign x_5087 = v_2094 | v_98;
assign x_5088 = v_2094 | v_86;
assign x_5089 = v_2093 | ~v_98;
assign x_5090 = v_2093 | v_78;
assign x_5091 = v_2092 | v_99;
assign x_5092 = v_2092 | v_85;
assign x_5093 = v_2091 | ~v_99;
assign x_5094 = v_2091 | v_77;
assign x_5095 = v_2090 | v_118;
assign x_5096 = v_2090 | v_90;
assign x_5097 = v_2089 | ~v_118;
assign x_5098 = v_2089 | v_82;
assign x_5099 = v_50 | v_51 | v_49 | v_48 | v_46 | v_101 | v_100 | v_102 | v_110 | ~v_2087 | ~v_2086 | ~v_2085 | ~v_268 | ~v_2084 | ~v_2083 | ~v_2082 | ~v_380 | ~v_379 | ~v_261 | ~v_2081 | ~v_2080 | ~v_2079 | ~v_2078 | ~v_351 | ~v_350 | ~v_378 | ~v_377 | v_2088;
assign x_5100 = v_2087 | v_119;
assign x_5101 = v_2087 | v_62;
assign x_5102 = v_2086 | ~v_97;
assign x_5103 = v_2086 | v_55;
assign x_5104 = v_2085 | v_97;
assign x_5105 = v_2085 | v_63;
assign x_5106 = v_2084 | ~v_119;
assign x_5107 = v_2084 | v_54;
assign x_5108 = v_2083 | ~v_98;
assign x_5109 = v_2083 | v_53;
assign x_5110 = v_2082 | v_98;
assign x_5111 = v_2082 | v_61;
assign x_5112 = v_2081 | v_99;
assign x_5113 = v_2081 | v_60;
assign x_5114 = v_2080 | ~v_99;
assign x_5115 = v_2080 | v_52;
assign x_5116 = v_2079 | v_118;
assign x_5117 = v_2079 | v_65;
assign x_5118 = v_2078 | ~v_118;
assign x_5119 = v_2078 | v_57;
assign x_5120 = v_25 | v_24 | v_23 | v_22 | v_20 | v_95 | v_94 | ~v_2076 | v_93 | v_108 | ~v_375 | ~v_2075 | ~v_2074 | ~v_2073 | ~v_2072 | ~v_374 | ~v_253 | ~v_252 | ~v_2071 | ~v_2070 | ~v_2069 | ~v_2068 | ~v_2067 | ~v_340 | ~v_339 | ~v_373 | ~v_372 | v_2077;
assign x_5121 = v_2076 | ~v_98;
assign x_5122 = v_2076 | v_28;
assign x_5123 = v_2075 | v_119;
assign x_5124 = v_2075 | v_37;
assign x_5125 = v_2074 | ~v_119;
assign x_5126 = v_2074 | v_29;
assign x_5127 = v_2073 | v_99;
assign x_5128 = v_2073 | v_35;
assign x_5129 = v_2072 | v_98;
assign x_5130 = v_2072 | v_36;
assign x_5131 = v_2071 | v_97;
assign x_5132 = v_2071 | v_38;
assign x_5133 = v_2070 | ~v_97;
assign x_5134 = v_2070 | v_30;
assign x_5135 = v_2069 | ~v_99;
assign x_5136 = v_2069 | v_27;
assign x_5137 = v_2068 | v_118;
assign x_5138 = v_2068 | v_40;
assign x_5139 = v_2067 | ~v_118;
assign x_5140 = v_2067 | v_32;
assign x_5141 = v_2066 | ~v_1822;
assign x_5142 = v_2066 | ~v_1887;
assign x_5143 = v_2066 | ~v_1910;
assign x_5144 = v_2066 | ~v_1933;
assign x_5145 = v_2066 | ~v_1942;
assign x_5146 = v_2066 | ~v_1961;
assign x_5147 = v_2066 | ~v_1978;
assign x_5148 = v_2066 | ~v_1987;
assign x_5149 = v_2066 | ~v_1996;
assign x_5150 = v_2066 | ~v_2005;
assign x_5151 = v_2066 | ~v_2014;
assign x_5152 = v_2066 | ~v_2023;
assign x_5153 = v_2066 | ~v_2032;
assign x_5154 = v_2066 | ~v_2041;
assign x_5155 = v_2066 | ~v_2050;
assign x_5156 = v_2066 | ~v_2065;
assign x_5157 = v_9 | v_7 | v_5 | v_4 | v_6 | v_3 | v_2 | v_1 | ~v_1041 | ~v_1040 | ~v_2064 | v_2065;
assign x_5158 = v_2064 | ~v_2057;
assign x_5159 = v_2064 | ~v_2063;
assign x_5160 = v_116 | ~v_1819 | ~v_1811 | ~v_1006 | ~v_1958 | ~v_1975 | ~v_1884 | ~v_2062 | v_2063;
assign x_5161 = v_2062 | ~v_2061;
assign x_5162 = v_2062 | ~v_698;
assign x_5163 = v_2062 | ~v_699;
assign x_5164 = v_2062 | ~v_700;
assign x_5165 = v_2062 | ~v_701;
assign x_5166 = ~v_2060 | ~v_2059 | ~v_2058 | v_2061;
assign x_5167 = v_2060 | ~v_1675;
assign x_5168 = v_2060 | ~v_1676;
assign x_5169 = v_2060 | ~v_1372;
assign x_5170 = v_2060 | ~v_1625;
assign x_5171 = v_2060 | ~v_1626;
assign x_5172 = v_2060 | ~v_763;
assign x_5173 = v_2060 | ~v_764;
assign x_5174 = v_2060 | ~v_726;
assign x_5175 = v_2060 | ~v_1373;
assign x_5176 = v_2060 | ~v_1677;
assign x_5177 = v_2060 | ~v_1678;
assign x_5178 = v_2060 | ~v_1754;
assign x_5179 = v_2060 | ~v_1755;
assign x_5180 = v_2060 | ~v_1756;
assign x_5181 = v_2060 | ~v_731;
assign x_5182 = v_2060 | ~v_1374;
assign x_5183 = v_2060 | ~v_1757;
assign x_5184 = v_2060 | ~v_1375;
assign x_5185 = v_2060 | ~v_112;
assign x_5186 = v_2060 | ~v_105;
assign x_5187 = v_2060 | ~v_76;
assign x_5188 = v_2060 | ~v_75;
assign x_5189 = v_2060 | ~v_74;
assign x_5190 = v_2060 | ~v_73;
assign x_5191 = v_2060 | ~v_72;
assign x_5192 = v_2060 | ~v_71;
assign x_5193 = v_2060 | ~v_69;
assign x_5194 = v_2059 | ~v_1670;
assign x_5195 = v_2059 | ~v_1671;
assign x_5196 = v_2059 | ~v_1367;
assign x_5197 = v_2059 | ~v_1368;
assign x_5198 = v_2059 | ~v_1614;
assign x_5199 = v_2059 | ~v_1615;
assign x_5200 = v_2059 | ~v_750;
assign x_5201 = v_2059 | ~v_714;
assign x_5202 = v_2059 | ~v_1672;
assign x_5203 = v_2059 | ~v_1673;
assign x_5204 = v_2059 | ~v_1749;
assign x_5205 = v_2059 | ~v_1750;
assign x_5206 = v_2059 | ~v_1751;
assign x_5207 = v_2059 | ~v_1752;
assign x_5208 = v_2059 | ~v_757;
assign x_5209 = v_2059 | ~v_1369;
assign x_5210 = v_2059 | ~v_721;
assign x_5211 = v_2059 | ~v_110;
assign x_5212 = v_2059 | ~v_101;
assign x_5213 = v_2059 | ~v_1370;
assign x_5214 = v_2059 | ~v_51;
assign x_5215 = v_2059 | ~v_50;
assign x_5216 = v_2059 | ~v_49;
assign x_5217 = v_2059 | ~v_48;
assign x_5218 = v_2059 | ~v_47;
assign x_5219 = v_2059 | ~v_46;
assign x_5220 = v_2059 | ~v_44;
assign x_5221 = v_2058 | ~v_1665;
assign x_5222 = v_2058 | ~v_1666;
assign x_5223 = v_2058 | ~v_1362;
assign x_5224 = v_2058 | ~v_1603;
assign x_5225 = v_2058 | ~v_1604;
assign x_5226 = v_2058 | ~v_739;
assign x_5227 = v_2058 | ~v_705;
assign x_5228 = v_2058 | ~v_706;
assign x_5229 = v_2058 | ~v_1667;
assign x_5230 = v_2058 | ~v_1744;
assign x_5231 = v_2058 | ~v_1745;
assign x_5232 = v_2058 | ~v_1746;
assign x_5233 = v_2058 | ~v_1363;
assign x_5234 = v_2058 | ~v_746;
assign x_5235 = v_2058 | ~v_1364;
assign x_5236 = v_2058 | ~v_1365;
assign x_5237 = v_2058 | ~v_1668;
assign x_5238 = v_2058 | ~v_1747;
assign x_5239 = v_2058 | ~v_108;
assign x_5240 = v_2058 | ~v_94;
assign x_5241 = v_2058 | ~v_25;
assign x_5242 = v_2058 | ~v_24;
assign x_5243 = v_2058 | ~v_23;
assign x_5244 = v_2058 | ~v_22;
assign x_5245 = v_2058 | ~v_21;
assign x_5246 = v_2058 | ~v_20;
assign x_5247 = v_2058 | ~v_18;
assign x_5248 = ~v_1601 | ~v_2056 | v_2057;
assign x_5249 = v_2056 | ~v_2055;
assign x_5250 = v_2056 | ~v_1852;
assign x_5251 = v_2056 | ~v_1967;
assign x_5252 = v_2056 | ~v_1949;
assign x_5253 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_2054 | v_2055;
assign x_5254 = v_2054 | ~v_2051;
assign x_5255 = v_2054 | ~v_2052;
assign x_5256 = v_2054 | ~v_2053;
assign x_5257 = v_76 | v_69 | v_75 | v_74 | v_73 | v_72 | v_71 | v_105 | ~v_1356 | v_112 | ~v_1537 | ~v_1355 | ~v_278 | ~v_1536 | ~v_1535 | ~v_1534 | ~v_1458 | ~v_1457 | ~v_1354 | ~v_273 | ~v_311 | ~v_310 | ~v_1406 | ~v_1405 | ~v_1353 | ~v_1456 | ~v_1455 | v_2053;
assign x_5258 = v_50 | v_51 | v_49 | v_48 | v_46 | v_47 | v_44 | ~v_1351 | v_101 | v_110 | ~v_268 | ~v_1350 | ~v_304 | ~v_1532 | ~v_1531 | ~v_1530 | ~v_1529 | ~v_1453 | ~v_1452 | ~v_261 | ~v_297 | ~v_1395 | ~v_1394 | ~v_1349 | ~v_1348 | ~v_1451 | ~v_1450 | v_2052;
assign x_5259 = v_25 | v_24 | v_23 | v_22 | v_21 | v_20 | v_18 | v_94 | v_108 | ~v_1527 | ~v_1448 | ~v_1346 | ~v_1345 | ~v_293 | ~v_1344 | ~v_1526 | ~v_1525 | ~v_1524 | ~v_1447 | ~v_253 | ~v_252 | ~v_286 | ~v_1384 | ~v_1383 | ~v_1343 | ~v_1446 | ~v_1445 | v_2051;
assign x_5260 = v_9 | v_7 | v_5 | v_4 | v_10 | v_3 | v_2 | v_1 | ~v_1041 | ~v_1040 | ~v_2049 | v_2050;
assign x_5261 = v_2049 | ~v_2045;
assign x_5262 = v_2049 | ~v_2048;
assign x_5263 = v_116 | ~v_1819 | ~v_1811 | ~v_1006 | ~v_1867 | ~v_1882 | ~v_1866 | ~v_1865 | ~v_1881 | ~v_2047 | ~v_2046 | v_2048;
assign x_5264 = v_2047 | ~v_1873;
assign x_5265 = v_2047 | ~v_1925;
assign x_5266 = v_2046 | ~v_1879;
assign x_5267 = v_2046 | ~v_1780;
assign x_5268 = ~v_1601 | ~v_2044 | v_2045;
assign x_5269 = v_2044 | ~v_2042;
assign x_5270 = v_2044 | ~v_2043;
assign x_5271 = v_2044 | ~v_1849;
assign x_5272 = v_2044 | ~v_1833;
assign x_5273 = v_2044 | ~v_1834;
assign x_5274 = v_2044 | ~v_1850;
assign x_5275 = v_2044 | ~v_1835;
assign x_5276 = ~v_1914 | ~v_1841 | v_2043;
assign x_5277 = ~v_1560 | ~v_1847 | v_2042;
assign x_5278 = v_7 | v_4 | v_6 | v_8 | v_10 | v_3 | v_2 | ~v_1041 | ~v_1040 | ~v_2040 | v_2041;
assign x_5279 = v_2040 | ~v_2036;
assign x_5280 = v_2040 | ~v_2039;
assign x_5281 = v_116 | ~v_1819 | ~v_1811 | ~v_1006 | ~v_1776 | ~v_1775 | ~v_1774 | ~v_1798 | ~v_1796 | ~v_2038 | ~v_2037 | v_2039;
assign x_5282 = v_2038 | ~v_1875;
assign x_5283 = v_2038 | ~v_1873;
assign x_5284 = v_2037 | ~v_1780;
assign x_5285 = v_2037 | ~v_1906;
assign x_5286 = ~v_1601 | ~v_2035 | v_2036;
assign x_5287 = v_2035 | ~v_2033;
assign x_5288 = v_2035 | ~v_2034;
assign x_5289 = v_2035 | ~v_1576;
assign x_5290 = v_2035 | ~v_1578;
assign x_5291 = v_2035 | ~v_1554;
assign x_5292 = v_2035 | ~v_1555;
assign x_5293 = v_2035 | ~v_1556;
assign x_5294 = ~v_1841 | ~v_1843 | v_2034;
assign x_5295 = ~v_1895 | ~v_1560 | v_2033;
assign x_5296 = v_9 | v_7 | v_5 | v_4 | v_6 | v_8 | v_3 | v_2 | ~v_1041 | ~v_1040 | ~v_2031 | v_2032;
assign x_5297 = v_2031 | ~v_2027;
assign x_5298 = v_2031 | ~v_2030;
assign x_5299 = v_116 | ~v_1819 | ~v_1811 | ~v_1006 | ~v_1736 | ~v_1735 | ~v_1730 | ~v_1905 | ~v_1904 | ~v_2029 | ~v_2028 | v_2030;
assign x_5300 = v_2029 | ~v_1799;
assign x_5301 = v_2029 | ~v_1902;
assign x_5302 = v_2028 | ~v_1873;
assign x_5303 = v_2028 | ~v_1742;
assign x_5304 = ~v_1601 | ~v_2026 | v_2027;
assign x_5305 = v_2026 | ~v_2024;
assign x_5306 = v_2026 | ~v_2025;
assign x_5307 = v_2026 | ~v_1893;
assign x_5308 = v_2026 | ~v_1894;
assign x_5309 = v_2026 | ~v_1510;
assign x_5310 = v_2026 | ~v_1515;
assign x_5311 = v_2026 | ~v_1516;
assign x_5312 = ~v_1891 | ~v_1579 | v_2025;
assign x_5313 = ~v_1522 | ~v_1841 | v_2024;
assign x_5314 = v_9 | v_7 | v_5 | v_4 | v_8 | v_10 | v_3 | v_2 | ~v_1041 | ~v_1040 | ~v_2022 | v_2023;
assign x_5315 = v_2022 | ~v_2018;
assign x_5316 = v_2022 | ~v_2021;
assign x_5317 = v_116 | ~v_1819 | ~v_1811 | ~v_1006 | ~v_1872 | ~v_1871 | ~v_1870 | ~v_1869 | ~v_1864 | ~v_2020 | ~v_2019 | v_2021;
assign x_5318 = v_2020 | ~v_1799;
assign x_5319 = v_2020 | ~v_1879;
assign x_5320 = v_2019 | ~v_1883;
assign x_5321 = v_2019 | ~v_1906;
assign x_5322 = ~v_1601 | ~v_2017 | v_2018;
assign x_5323 = v_2017 | ~v_2015;
assign x_5324 = v_2017 | ~v_2016;
assign x_5325 = v_2017 | ~v_1832;
assign x_5326 = v_2017 | ~v_1837;
assign x_5327 = v_2017 | ~v_1838;
assign x_5328 = v_2017 | ~v_1839;
assign x_5329 = v_2017 | ~v_1840;
assign x_5330 = ~v_1847 | ~v_1579 | v_2016;
assign x_5331 = ~v_1895 | ~v_1851 | v_2015;
assign x_5332 = v_7 | v_4 | v_6 | v_10 | v_3 | v_2 | v_1 | ~v_1041 | ~v_1040 | ~v_2013 | v_2014;
assign x_5333 = v_2013 | ~v_2009;
assign x_5334 = v_2013 | ~v_2012;
assign x_5335 = v_116 | ~v_1819 | ~v_1811 | ~v_1006 | ~v_1779 | ~v_1778 | ~v_1773 | ~v_1768 | ~v_1767 | ~v_2011 | ~v_2010 | v_2012;
assign x_5336 = v_2011 | ~v_1799;
assign x_5337 = v_2011 | ~v_1925;
assign x_5338 = v_2010 | ~v_1875;
assign x_5339 = v_2010 | ~v_1883;
assign x_5340 = ~v_1601 | ~v_2008 | v_2009;
assign x_5341 = v_2008 | ~v_2006;
assign x_5342 = v_2008 | ~v_2007;
assign x_5343 = v_2008 | ~v_1547;
assign x_5344 = v_2008 | ~v_1548;
assign x_5345 = v_2008 | ~v_1553;
assign x_5346 = v_2008 | ~v_1558;
assign x_5347 = v_2008 | ~v_1559;
assign x_5348 = ~v_1914 | ~v_1579 | v_2007;
assign x_5349 = ~v_1851 | ~v_1843 | v_2006;
assign x_5350 = v_9 | v_5 | v_6 | v_8 | v_10 | v_3 | v_1 | ~v_1041 | ~v_1040 | ~v_2004 | v_2005;
assign x_5351 = v_2004 | ~v_2000;
assign x_5352 = v_2004 | ~v_2003;
assign x_5353 = v_116 | ~v_1819 | ~v_1811 | ~v_1006 | ~v_1789 | ~v_1788 | ~v_1787 | ~v_1928 | ~v_1927 | ~v_2002 | ~v_2001 | v_2003;
assign x_5354 = v_2002 | ~v_1795;
assign x_5355 = v_2002 | ~v_1879;
assign x_5356 = v_2001 | ~v_1902;
assign x_5357 = v_2001 | ~v_1925;
assign x_5358 = ~v_1601 | ~v_1999 | v_2000;
assign x_5359 = v_1999 | ~v_1997;
assign x_5360 = v_1999 | ~v_1998;
assign x_5361 = v_1999 | ~v_1916;
assign x_5362 = v_1999 | ~v_1917;
assign x_5363 = v_1999 | ~v_1567;
assign x_5364 = v_1999 | ~v_1568;
assign x_5365 = v_1999 | ~v_1569;
assign x_5366 = ~v_1847 | ~v_1575 | v_1998;
assign x_5367 = ~v_1914 | ~v_1891 | v_1997;
assign x_5368 = v_9 | v_5 | v_4 | v_6 | v_8 | v_3 | v_1 | ~v_1041 | ~v_1040 | ~v_1995 | v_1996;
assign x_5369 = v_1995 | ~v_1991;
assign x_5370 = v_1995 | ~v_1994;
assign x_5371 = v_116 | ~v_1819 | ~v_1811 | ~v_1006 | ~v_1719 | ~v_1714 | ~v_1681 | ~v_1901 | ~v_1900 | ~v_1993 | ~v_1992 | v_1994;
assign x_5372 = v_1993 | ~v_1929;
assign x_5373 = v_1993 | ~v_1906;
assign x_5374 = v_1992 | ~v_1879;
assign x_5375 = v_1992 | ~v_1742;
assign x_5376 = ~v_1601 | ~v_1990 | v_1991;
assign x_5377 = v_1990 | ~v_1988;
assign x_5378 = v_1990 | ~v_1989;
assign x_5379 = v_1990 | ~v_1889;
assign x_5380 = v_1990 | ~v_1890;
assign x_5381 = v_1990 | ~v_1461;
assign x_5382 = v_1990 | ~v_1494;
assign x_5383 = v_1990 | ~v_1499;
assign x_5384 = ~v_1895 | ~v_1918 | v_1989;
assign x_5385 = ~v_1522 | ~v_1847 | v_1988;
assign x_5386 = v_9 | v_5 | v_4 | v_8 | v_10 | v_3 | v_1 | ~v_1041 | ~v_1040 | ~v_1986 | v_1987;
assign x_5387 = v_1986 | ~v_1982;
assign x_5388 = v_1986 | ~v_1985;
assign x_5389 = v_116 | ~v_1819 | ~v_1811 | ~v_1006 | ~v_1862 | ~v_1861 | ~v_1860 | ~v_1878 | ~v_1877 | ~v_1984 | ~v_1983 | v_1985;
assign x_5390 = v_1984 | ~v_1929;
assign x_5391 = v_1984 | ~v_1873;
assign x_5392 = v_1983 | ~v_1883;
assign x_5393 = v_1983 | ~v_1902;
assign x_5394 = ~v_1601 | ~v_1981 | v_1982;
assign x_5395 = v_1981 | ~v_1979;
assign x_5396 = v_1981 | ~v_1980;
assign x_5397 = v_1981 | ~v_1845;
assign x_5398 = v_1981 | ~v_1846;
assign x_5399 = v_1981 | ~v_1828;
assign x_5400 = v_1981 | ~v_1829;
assign x_5401 = v_1981 | ~v_1830;
assign x_5402 = ~v_1841 | ~v_1918 | v_1980;
assign x_5403 = ~v_1891 | ~v_1851 | v_1979;
assign x_5404 = v_4 | v_6 | v_8 | v_10 | v_3 | v_1 | ~v_1041 | ~v_1040 | ~v_1977 | v_1978;
assign x_5405 = v_1977 | ~v_1969;
assign x_5406 = v_1977 | ~v_1976;
assign x_5407 = v_116 | ~v_1819 | ~v_1811 | ~v_1006 | ~v_1975 | ~v_1957 | ~v_1880 | ~v_1974 | v_1976;
assign x_5408 = v_1975 | ~v_1780;
assign x_5409 = v_1975 | ~v_1902;
assign x_5410 = v_1974 | ~v_1973;
assign x_5411 = v_1974 | ~v_698;
assign x_5412 = v_1974 | ~v_699;
assign x_5413 = v_1974 | ~v_700;
assign x_5414 = v_1974 | ~v_701;
assign x_5415 = ~v_1972 | ~v_1971 | ~v_1970 | v_1973;
assign x_5416 = v_1972 | ~v_1655;
assign x_5417 = v_1972 | ~v_1656;
assign x_5418 = v_1972 | ~v_1218;
assign x_5419 = v_1972 | ~v_1219;
assign x_5420 = v_1972 | ~v_814;
assign x_5421 = v_1972 | ~v_815;
assign x_5422 = v_1972 | ~v_1625;
assign x_5423 = v_1972 | ~v_1626;
assign x_5424 = v_1972 | ~v_632;
assign x_5425 = v_1972 | ~v_633;
assign x_5426 = v_1972 | ~v_1629;
assign x_5427 = v_1972 | ~v_1630;
assign x_5428 = v_1972 | ~v_1220;
assign x_5429 = v_1972 | ~v_1221;
assign x_5430 = v_1972 | ~v_1661;
assign x_5431 = v_1972 | ~v_1662;
assign x_5432 = v_1972 | ~v_1632;
assign x_5433 = v_1972 | ~v_1633;
assign x_5434 = v_1972 | ~v_113;
assign x_5435 = v_1972 | ~v_106;
assign x_5436 = v_1972 | ~v_76;
assign x_5437 = v_1972 | ~v_75;
assign x_5438 = v_1972 | ~v_74;
assign x_5439 = v_1972 | ~v_73;
assign x_5440 = v_1972 | ~v_70;
assign x_5441 = v_1972 | ~v_69;
assign x_5442 = v_1972 | ~v_68;
assign x_5443 = v_1971 | ~v_1646;
assign x_5444 = v_1971 | ~v_1647;
assign x_5445 = v_1971 | ~v_1213;
assign x_5446 = v_1971 | ~v_1214;
assign x_5447 = v_1971 | ~v_803;
assign x_5448 = v_1971 | ~v_804;
assign x_5449 = v_1971 | ~v_1614;
assign x_5450 = v_1971 | ~v_1615;
assign x_5451 = v_1971 | ~v_613;
assign x_5452 = v_1971 | ~v_614;
assign x_5453 = v_1971 | ~v_1618;
assign x_5454 = v_1971 | ~v_1619;
assign x_5455 = v_1971 | ~v_1215;
assign x_5456 = v_1971 | ~v_1216;
assign x_5457 = v_1971 | ~v_1652;
assign x_5458 = v_1971 | ~v_1653;
assign x_5459 = v_1971 | ~v_1622;
assign x_5460 = v_1971 | ~v_1623;
assign x_5461 = v_1971 | ~v_111;
assign x_5462 = v_1971 | ~v_102;
assign x_5463 = v_1971 | ~v_51;
assign x_5464 = v_1971 | ~v_50;
assign x_5465 = v_1971 | ~v_49;
assign x_5466 = v_1971 | ~v_48;
assign x_5467 = v_1971 | ~v_45;
assign x_5468 = v_1971 | ~v_44;
assign x_5469 = v_1971 | ~v_43;
assign x_5470 = v_1970 | ~v_1637;
assign x_5471 = v_1970 | ~v_1638;
assign x_5472 = v_1970 | ~v_1208;
assign x_5473 = v_1970 | ~v_1209;
assign x_5474 = v_1970 | ~v_792;
assign x_5475 = v_1970 | ~v_793;
assign x_5476 = v_1970 | ~v_1603;
assign x_5477 = v_1970 | ~v_1604;
assign x_5478 = v_1970 | ~v_594;
assign x_5479 = v_1970 | ~v_595;
assign x_5480 = v_1970 | ~v_1607;
assign x_5481 = v_1970 | ~v_1608;
assign x_5482 = v_1970 | ~v_1210;
assign x_5483 = v_1970 | ~v_1211;
assign x_5484 = v_1970 | ~v_1642;
assign x_5485 = v_1970 | ~v_1643;
assign x_5486 = v_1970 | ~v_1610;
assign x_5487 = v_1970 | ~v_1611;
assign x_5488 = v_1970 | ~v_109;
assign x_5489 = v_1970 | ~v_95;
assign x_5490 = v_1970 | ~v_25;
assign x_5491 = v_1970 | ~v_24;
assign x_5492 = v_1970 | ~v_23;
assign x_5493 = v_1970 | ~v_22;
assign x_5494 = v_1970 | ~v_19;
assign x_5495 = v_1970 | ~v_18;
assign x_5496 = v_1970 | ~v_17;
assign x_5497 = ~v_1601 | ~v_1968 | v_1969;
assign x_5498 = v_1968 | ~v_1966;
assign x_5499 = v_1968 | ~v_1848;
assign x_5500 = v_1968 | ~v_1948;
assign x_5501 = v_1968 | ~v_1967;
assign x_5502 = ~v_1891 | ~v_1560 | v_1967;
assign x_5503 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1965 | v_1966;
assign x_5504 = v_1965 | ~v_1962;
assign x_5505 = v_1965 | ~v_1963;
assign x_5506 = v_1965 | ~v_1964;
assign x_5507 = v_76 | v_69 | v_68 | v_75 | v_74 | v_73 | v_70 | v_106 | v_113 | ~v_1413 | ~v_1412 | ~v_1442 | ~v_1441 | ~v_1200 | ~v_1199 | ~v_1410 | ~v_1409 | ~v_180 | ~v_179 | ~v_1406 | ~v_1405 | ~v_362 | ~v_361 | ~v_1198 | ~v_1197 | ~v_1436 | ~v_1435 | v_1964;
assign x_5508 = v_50 | v_51 | v_49 | v_48 | v_45 | v_43 | v_44 | v_102 | v_111 | ~v_1403 | ~v_1402 | ~v_1433 | ~v_1432 | ~v_1195 | ~v_1194 | ~v_1399 | ~v_1398 | ~v_161 | ~v_160 | ~v_1395 | ~v_1394 | ~v_351 | ~v_350 | ~v_1193 | ~v_1192 | ~v_1427 | ~v_1426 | v_1963;
assign x_5509 = v_25 | v_24 | v_23 | v_22 | v_19 | v_18 | v_17 | v_95 | v_109 | ~v_1391 | ~v_1390 | ~v_1423 | ~v_1422 | ~v_1190 | ~v_1189 | ~v_1388 | ~v_1387 | ~v_142 | ~v_141 | ~v_1384 | ~v_1383 | ~v_340 | ~v_339 | ~v_1188 | ~v_1187 | ~v_1418 | ~v_1417 | v_1962;
assign x_5510 = v_9 | v_7 | v_5 | v_6 | v_8 | v_10 | v_3 | v_2 | ~v_1041 | ~v_1040 | ~v_1960 | v_1961;
assign x_5511 = v_1960 | ~v_1951;
assign x_5512 = v_1960 | ~v_1959;
assign x_5513 = v_116 | ~v_1819 | ~v_1811 | ~v_1006 | ~v_1958 | ~v_1957 | ~v_1874 | ~v_1956 | v_1959;
assign x_5514 = v_1958 | ~v_1925;
assign x_5515 = v_1958 | ~v_1906;
assign x_5516 = v_1957 | ~v_1929;
assign x_5517 = v_1957 | ~v_1799;
assign x_5518 = v_1956 | ~v_1955;
assign x_5519 = v_1956 | ~v_698;
assign x_5520 = v_1956 | ~v_699;
assign x_5521 = v_1956 | ~v_700;
assign x_5522 = v_1956 | ~v_701;
assign x_5523 = ~v_1954 | ~v_1953 | ~v_1952 | v_1955;
assign x_5524 = v_1954 | ~v_1708;
assign x_5525 = v_1954 | ~v_1167;
assign x_5526 = v_1954 | ~v_1168;
assign x_5527 = v_1954 | ~v_1625;
assign x_5528 = v_1954 | ~v_1626;
assign x_5529 = v_1954 | ~v_634;
assign x_5530 = v_1954 | ~v_635;
assign x_5531 = v_1954 | ~v_1692;
assign x_5532 = v_1954 | ~v_1693;
assign x_5533 = v_1954 | ~v_1169;
assign x_5534 = v_1954 | ~v_1170;
assign x_5535 = v_1954 | ~v_688;
assign x_5536 = v_1954 | ~v_689;
assign x_5537 = v_1954 | ~v_1709;
assign x_5538 = v_1954 | ~v_1710;
assign x_5539 = v_1954 | ~v_1694;
assign x_5540 = v_1954 | ~v_1695;
assign x_5541 = v_1954 | ~v_1711;
assign x_5542 = v_1954 | ~v_132;
assign x_5543 = v_1954 | ~v_127;
assign x_5544 = v_1954 | ~v_113;
assign x_5545 = v_1954 | ~v_112;
assign x_5546 = v_1954 | ~v_106;
assign x_5547 = v_1954 | ~v_105;
assign x_5548 = v_1954 | ~v_76;
assign x_5549 = v_1954 | ~v_75;
assign x_5550 = v_1954 | ~v_69;
assign x_5551 = v_1953 | ~v_1703;
assign x_5552 = v_1953 | ~v_1704;
assign x_5553 = v_1953 | ~v_1614;
assign x_5554 = v_1953 | ~v_1615;
assign x_5555 = v_1953 | ~v_615;
assign x_5556 = v_1953 | ~v_616;
assign x_5557 = v_1953 | ~v_1687;
assign x_5558 = v_1953 | ~v_1688;
assign x_5559 = v_1953 | ~v_1162;
assign x_5560 = v_1953 | ~v_1163;
assign x_5561 = v_1953 | ~v_669;
assign x_5562 = v_1953 | ~v_670;
assign x_5563 = v_1953 | ~v_1164;
assign x_5564 = v_1953 | ~v_1165;
assign x_5565 = v_1953 | ~v_1705;
assign x_5566 = v_1953 | ~v_1706;
assign x_5567 = v_1953 | ~v_1689;
assign x_5568 = v_1953 | ~v_1690;
assign x_5569 = v_1953 | ~v_131;
assign x_5570 = v_1953 | ~v_126;
assign x_5571 = v_1953 | ~v_111;
assign x_5572 = v_1953 | ~v_110;
assign x_5573 = v_1953 | ~v_102;
assign x_5574 = v_1953 | ~v_101;
assign x_5575 = v_1953 | ~v_51;
assign x_5576 = v_1953 | ~v_50;
assign x_5577 = v_1953 | ~v_44;
assign x_5578 = v_1952 | ~v_1698;
assign x_5579 = v_1952 | ~v_1699;
assign x_5580 = v_1952 | ~v_1603;
assign x_5581 = v_1952 | ~v_1604;
assign x_5582 = v_1952 | ~v_596;
assign x_5583 = v_1952 | ~v_597;
assign x_5584 = v_1952 | ~v_1682;
assign x_5585 = v_1952 | ~v_1683;
assign x_5586 = v_1952 | ~v_1157;
assign x_5587 = v_1952 | ~v_1158;
assign x_5588 = v_1952 | ~v_653;
assign x_5589 = v_1952 | ~v_654;
assign x_5590 = v_1952 | ~v_1159;
assign x_5591 = v_1952 | ~v_1160;
assign x_5592 = v_1952 | ~v_1700;
assign x_5593 = v_1952 | ~v_1701;
assign x_5594 = v_1952 | ~v_1684;
assign x_5595 = v_1952 | ~v_1685;
assign x_5596 = v_1952 | ~v_128;
assign x_5597 = v_1952 | ~v_122;
assign x_5598 = v_1952 | ~v_109;
assign x_5599 = v_1952 | ~v_108;
assign x_5600 = v_1952 | ~v_95;
assign x_5601 = v_1952 | ~v_94;
assign x_5602 = v_1952 | ~v_25;
assign x_5603 = v_1952 | ~v_24;
assign x_5604 = v_1952 | ~v_18;
assign x_5605 = ~v_1601 | ~v_1950 | v_1951;
assign x_5606 = v_1950 | ~v_1947;
assign x_5607 = v_1950 | ~v_1842;
assign x_5608 = v_1950 | ~v_1948;
assign x_5609 = v_1950 | ~v_1949;
assign x_5610 = ~v_1895 | ~v_1914 | v_1949;
assign x_5611 = ~v_1579 | ~v_1918 | v_1948;
assign x_5612 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1946 | v_1947;
assign x_5613 = v_1946 | ~v_1943;
assign x_5614 = v_1946 | ~v_1944;
assign x_5615 = v_1946 | ~v_1945;
assign x_5616 = v_76 | v_69 | v_75 | v_106 | v_105 | v_132 | v_127 | v_113 | v_112 | ~v_1491 | ~v_1475 | ~v_1474 | ~v_1490 | ~v_1489 | ~v_236 | ~v_235 | ~v_1141 | ~v_1140 | ~v_1473 | ~v_1472 | ~v_182 | ~v_181 | ~v_1406 | ~v_1405 | ~v_1139 | ~v_1138 | ~v_1488 | v_1945;
assign x_5617 = v_50 | v_51 | v_44 | v_101 | v_102 | v_111 | v_110 | v_131 | v_126 | ~v_1470 | ~v_1469 | ~v_1486 | ~v_1485 | ~v_1136 | ~v_1135 | ~v_217 | ~v_216 | ~v_1134 | ~v_1133 | ~v_1468 | ~v_1467 | ~v_163 | ~v_162 | ~v_1395 | ~v_1394 | ~v_1484 | ~v_1483 | v_1944;
assign x_5618 = v_25 | v_24 | v_18 | v_95 | v_94 | v_108 | v_109 | v_128 | v_122 | ~v_1465 | ~v_1464 | ~v_1481 | ~v_1480 | ~v_1131 | ~v_1130 | ~v_201 | ~v_200 | ~v_1129 | ~v_1128 | ~v_1463 | ~v_1462 | ~v_144 | ~v_143 | ~v_1384 | ~v_1383 | ~v_1479 | ~v_1478 | v_1943;
assign x_5619 = v_9 | v_7 | v_5 | v_6 | v_10 | v_3 | v_2 | v_1 | ~v_1041 | ~v_1040 | ~v_1941 | v_1942;
assign x_5620 = v_1941 | ~v_1937;
assign x_5621 = v_1941 | ~v_1940;
assign x_5622 = v_116 | ~v_1819 | ~v_1811 | ~v_1006 | ~v_1784 | ~v_1924 | ~v_1922 | ~v_1783 | ~v_1782 | ~v_1939 | ~v_1938 | v_1940;
assign x_5623 = v_1939 | ~v_1929;
assign x_5624 = v_1939 | ~v_1780;
assign x_5625 = v_1938 | ~v_1795;
assign x_5626 = v_1938 | ~v_1883;
assign x_5627 = ~v_1601 | ~v_1936 | v_1937;
assign x_5628 = v_1936 | ~v_1934;
assign x_5629 = v_1936 | ~v_1935;
assign x_5630 = v_1936 | ~v_1562;
assign x_5631 = v_1936 | ~v_1563;
assign x_5632 = v_1936 | ~v_1911;
assign x_5633 = v_1936 | ~v_1913;
assign x_5634 = v_1936 | ~v_1564;
assign x_5635 = ~v_1560 | ~v_1918 | v_1935;
assign x_5636 = ~v_1851 | ~v_1575 | v_1934;
assign x_5637 = v_9 | v_7 | v_5 | v_6 | v_8 | v_10 | v_2 | v_1 | ~v_1041 | ~v_1040 | ~v_1932 | v_1933;
assign x_5638 = v_1932 | ~v_1921;
assign x_5639 = v_1932 | ~v_1931;
assign x_5640 = v_116 | ~v_1819 | ~v_1811 | ~v_1006 | ~v_1794 | ~v_1793 | ~v_1792 | ~v_1791 | ~v_1786 | ~v_1930 | ~v_1926 | v_1931;
assign x_5641 = v_1930 | ~v_1929;
assign x_5642 = v_1930 | ~v_1875;
assign x_5643 = ~v_1789 | ~v_1788 | ~v_1787 | ~v_1928 | ~v_1927 | v_1929;
assign x_5644 = v_1928 | ~v_1923;
assign x_5645 = v_1928 | ~v_1664;
assign x_5646 = v_1928 | ~v_698;
assign x_5647 = v_1928 | ~v_699;
assign x_5648 = v_1928 | ~v_700;
assign x_5649 = v_1928 | ~v_701;
assign x_5650 = v_1927 | ~v_1785;
assign x_5651 = v_1927 | ~v_1718;
assign x_5652 = v_1927 | ~v_698;
assign x_5653 = v_1927 | ~v_699;
assign x_5654 = v_1927 | ~v_700;
assign x_5655 = v_1927 | ~v_701;
assign x_5656 = v_1926 | ~v_1742;
assign x_5657 = v_1926 | ~v_1925;
assign x_5658 = ~v_1784 | ~v_1924 | ~v_1922 | ~v_1783 | ~v_1782 | v_1925;
assign x_5659 = v_1924 | ~v_1766;
assign x_5660 = v_1924 | ~v_1923;
assign x_5661 = v_1924 | ~v_698;
assign x_5662 = v_1924 | ~v_699;
assign x_5663 = v_1924 | ~v_700;
assign x_5664 = v_1924 | ~v_701;
assign x_5665 = ~v_1794 | ~v_1793 | ~v_1792 | v_1923;
assign x_5666 = v_1922 | ~v_1759;
assign x_5667 = v_1922 | ~v_1790;
assign x_5668 = v_1922 | ~v_698;
assign x_5669 = v_1922 | ~v_699;
assign x_5670 = v_1922 | ~v_700;
assign x_5671 = v_1922 | ~v_701;
assign x_5672 = ~v_1601 | ~v_1920 | v_1921;
assign x_5673 = v_1920 | ~v_1915;
assign x_5674 = v_1920 | ~v_1919;
assign x_5675 = v_1920 | ~v_1566;
assign x_5676 = v_1920 | ~v_1571;
assign x_5677 = v_1920 | ~v_1572;
assign x_5678 = v_1920 | ~v_1573;
assign x_5679 = v_1920 | ~v_1574;
assign x_5680 = ~v_1843 | ~v_1918 | v_1919;
assign x_5681 = v_1918 | ~v_1916;
assign x_5682 = v_1918 | ~v_1917;
assign x_5683 = v_1918 | ~v_1567;
assign x_5684 = v_1918 | ~v_1568;
assign x_5685 = v_1918 | ~v_1569;
assign x_5686 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1444 | ~v_1912 | v_1917;
assign x_5687 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1498 | ~v_1565 | v_1916;
assign x_5688 = ~v_1914 | ~v_1522 | v_1915;
assign x_5689 = v_1914 | ~v_1562;
assign x_5690 = v_1914 | ~v_1563;
assign x_5691 = v_1914 | ~v_1911;
assign x_5692 = v_1914 | ~v_1913;
assign x_5693 = v_1914 | ~v_1564;
assign x_5694 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1912 | ~v_1546 | v_1913;
assign x_5695 = v_1912 | ~v_1572;
assign x_5696 = v_1912 | ~v_1573;
assign x_5697 = v_1912 | ~v_1574;
assign x_5698 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1570 | ~v_1539 | v_1911;
assign x_5699 = v_9 | v_7 | v_5 | v_4 | v_6 | v_8 | v_2 | v_1 | ~v_1041 | ~v_1040 | ~v_1909 | v_1910;
assign x_5700 = v_1909 | ~v_1898;
assign x_5701 = v_1909 | ~v_1908;
assign x_5702 = v_116 | ~v_1819 | ~v_1811 | ~v_1006 | ~v_1741 | ~v_1740 | ~v_1739 | ~v_1738 | ~v_1721 | ~v_1907 | ~v_1903 | v_1908;
assign x_5703 = v_1907 | ~v_1795;
assign x_5704 = v_1907 | ~v_1906;
assign x_5705 = ~v_1736 | ~v_1735 | ~v_1730 | ~v_1905 | ~v_1904 | v_1906;
assign x_5706 = v_1905 | ~v_1720;
assign x_5707 = v_1905 | ~v_1734;
assign x_5708 = v_1905 | ~v_698;
assign x_5709 = v_1905 | ~v_699;
assign x_5710 = v_1905 | ~v_700;
assign x_5711 = v_1905 | ~v_701;
assign x_5712 = v_1904 | ~v_1899;
assign x_5713 = v_1904 | ~v_1729;
assign x_5714 = v_1904 | ~v_698;
assign x_5715 = v_1904 | ~v_699;
assign x_5716 = v_1904 | ~v_700;
assign x_5717 = v_1904 | ~v_701;
assign x_5718 = v_1903 | ~v_1875;
assign x_5719 = v_1903 | ~v_1902;
assign x_5720 = ~v_1719 | ~v_1714 | ~v_1681 | ~v_1901 | ~v_1900 | v_1902;
assign x_5721 = v_1901 | ~v_1697;
assign x_5722 = v_1901 | ~v_1737;
assign x_5723 = v_1901 | ~v_698;
assign x_5724 = v_1901 | ~v_699;
assign x_5725 = v_1901 | ~v_700;
assign x_5726 = v_1901 | ~v_701;
assign x_5727 = v_1900 | ~v_1899;
assign x_5728 = v_1900 | ~v_1664;
assign x_5729 = v_1900 | ~v_698;
assign x_5730 = v_1900 | ~v_699;
assign x_5731 = v_1900 | ~v_700;
assign x_5732 = v_1900 | ~v_701;
assign x_5733 = ~v_1741 | ~v_1740 | ~v_1739 | v_1899;
assign x_5734 = ~v_1601 | ~v_1897 | v_1898;
assign x_5735 = v_1897 | ~v_1892;
assign x_5736 = v_1897 | ~v_1896;
assign x_5737 = v_1897 | ~v_1501;
assign x_5738 = v_1897 | ~v_1518;
assign x_5739 = v_1897 | ~v_1519;
assign x_5740 = v_1897 | ~v_1520;
assign x_5741 = v_1897 | ~v_1521;
assign x_5742 = ~v_1895 | ~v_1575 | v_1896;
assign x_5743 = v_1895 | ~v_1893;
assign x_5744 = v_1895 | ~v_1894;
assign x_5745 = v_1895 | ~v_1510;
assign x_5746 = v_1895 | ~v_1515;
assign x_5747 = v_1895 | ~v_1516;
assign x_5748 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1514 | ~v_1500 | v_1894;
assign x_5749 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1509 | ~v_1888 | v_1893;
assign x_5750 = ~v_1891 | ~v_1843 | v_1892;
assign x_5751 = v_1891 | ~v_1889;
assign x_5752 = v_1891 | ~v_1890;
assign x_5753 = v_1891 | ~v_1461;
assign x_5754 = v_1891 | ~v_1494;
assign x_5755 = v_1891 | ~v_1499;
assign x_5756 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1517 | ~v_1477 | v_1890;
assign x_5757 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1444 | ~v_1888 | v_1889;
assign x_5758 = v_1888 | ~v_1519;
assign x_5759 = v_1888 | ~v_1520;
assign x_5760 = v_1888 | ~v_1521;
assign x_5761 = v_9 | v_7 | v_5 | v_4 | v_8 | v_10 | v_2 | v_1 | ~v_1041 | ~v_1040 | ~v_1886 | v_1887;
assign x_5762 = v_1886 | ~v_1854;
assign x_5763 = v_1886 | ~v_1885;
assign x_5764 = v_116 | ~v_1819 | ~v_1811 | ~v_1006 | ~v_1884 | ~v_1880 | ~v_1874 | ~v_1859 | v_1885;
assign x_5765 = v_1884 | ~v_1883;
assign x_5766 = v_1884 | ~v_1742;
assign x_5767 = ~v_1867 | ~v_1882 | ~v_1866 | ~v_1865 | ~v_1881 | v_1883;
assign x_5768 = v_1882 | ~v_1876;
assign x_5769 = v_1882 | ~v_1772;
assign x_5770 = v_1882 | ~v_698;
assign x_5771 = v_1882 | ~v_699;
assign x_5772 = v_1882 | ~v_700;
assign x_5773 = v_1882 | ~v_701;
assign x_5774 = v_1881 | ~v_1863;
assign x_5775 = v_1881 | ~v_1759;
assign x_5776 = v_1881 | ~v_698;
assign x_5777 = v_1881 | ~v_699;
assign x_5778 = v_1881 | ~v_700;
assign x_5779 = v_1881 | ~v_701;
assign x_5780 = v_1880 | ~v_1875;
assign x_5781 = v_1880 | ~v_1879;
assign x_5782 = ~v_1862 | ~v_1861 | ~v_1860 | ~v_1878 | ~v_1877 | v_1879;
assign x_5783 = v_1878 | ~v_1868;
assign x_5784 = v_1878 | ~v_1718;
assign x_5785 = v_1878 | ~v_698;
assign x_5786 = v_1878 | ~v_699;
assign x_5787 = v_1878 | ~v_700;
assign x_5788 = v_1878 | ~v_701;
assign x_5789 = v_1877 | ~v_1876;
assign x_5790 = v_1877 | ~v_1697;
assign x_5791 = v_1877 | ~v_698;
assign x_5792 = v_1877 | ~v_699;
assign x_5793 = v_1877 | ~v_700;
assign x_5794 = v_1877 | ~v_701;
assign x_5795 = ~v_1872 | ~v_1871 | ~v_1870 | v_1876;
assign x_5796 = ~v_1761 | ~v_1760 | ~v_1743 | ~v_1802 | ~v_1801 | v_1875;
assign x_5797 = v_1874 | ~v_1795;
assign x_5798 = v_1874 | ~v_1873;
assign x_5799 = ~v_1872 | ~v_1871 | ~v_1870 | ~v_1869 | ~v_1864 | v_1873;
assign x_5800 = v_1872 | ~v_1729;
assign x_5801 = v_1872 | ~v_698;
assign x_5802 = v_1872 | ~v_699;
assign x_5803 = v_1872 | ~v_700;
assign x_5804 = v_1872 | ~v_701;
assign x_5805 = v_1871 | ~v_1766;
assign x_5806 = v_1871 | ~v_1713;
assign x_5807 = v_1871 | ~v_698;
assign x_5808 = v_1871 | ~v_699;
assign x_5809 = v_1871 | ~v_700;
assign x_5810 = v_1871 | ~v_701;
assign x_5811 = v_1870 | ~v_1664;
assign x_5812 = v_1870 | ~v_1734;
assign x_5813 = v_1870 | ~v_698;
assign x_5814 = v_1870 | ~v_699;
assign x_5815 = v_1870 | ~v_700;
assign x_5816 = v_1870 | ~v_701;
assign x_5817 = v_1869 | ~v_1868;
assign x_5818 = v_1869 | ~v_1713;
assign x_5819 = v_1869 | ~v_698;
assign x_5820 = v_1869 | ~v_699;
assign x_5821 = v_1869 | ~v_700;
assign x_5822 = v_1869 | ~v_701;
assign x_5823 = ~v_1867 | ~v_1866 | ~v_1865 | v_1868;
assign x_5824 = v_1867 | ~v_1766;
assign x_5825 = v_1867 | ~v_698;
assign x_5826 = v_1867 | ~v_699;
assign x_5827 = v_1867 | ~v_700;
assign x_5828 = v_1867 | ~v_701;
assign x_5829 = v_1866 | ~v_1772;
assign x_5830 = v_1866 | ~v_1729;
assign x_5831 = v_1866 | ~v_698;
assign x_5832 = v_1866 | ~v_699;
assign x_5833 = v_1866 | ~v_700;
assign x_5834 = v_1866 | ~v_701;
assign x_5835 = v_1865 | ~v_1759;
assign x_5836 = v_1865 | ~v_1664;
assign x_5837 = v_1865 | ~v_698;
assign x_5838 = v_1865 | ~v_699;
assign x_5839 = v_1865 | ~v_700;
assign x_5840 = v_1865 | ~v_701;
assign x_5841 = v_1864 | ~v_1863;
assign x_5842 = v_1864 | ~v_1734;
assign x_5843 = v_1864 | ~v_698;
assign x_5844 = v_1864 | ~v_699;
assign x_5845 = v_1864 | ~v_700;
assign x_5846 = v_1864 | ~v_701;
assign x_5847 = ~v_1862 | ~v_1861 | ~v_1860 | v_1863;
assign x_5848 = v_1862 | ~v_1664;
assign x_5849 = v_1862 | ~v_698;
assign x_5850 = v_1862 | ~v_699;
assign x_5851 = v_1862 | ~v_700;
assign x_5852 = v_1862 | ~v_701;
assign x_5853 = v_1861 | ~v_1766;
assign x_5854 = v_1861 | ~v_1718;
assign x_5855 = v_1861 | ~v_698;
assign x_5856 = v_1861 | ~v_699;
assign x_5857 = v_1861 | ~v_700;
assign x_5858 = v_1861 | ~v_701;
assign x_5859 = v_1860 | ~v_1697;
assign x_5860 = v_1860 | ~v_1729;
assign x_5861 = v_1860 | ~v_698;
assign x_5862 = v_1860 | ~v_699;
assign x_5863 = v_1860 | ~v_700;
assign x_5864 = v_1860 | ~v_701;
assign x_5865 = v_1859 | ~v_1858;
assign x_5866 = v_1859 | ~v_698;
assign x_5867 = v_1859 | ~v_699;
assign x_5868 = v_1859 | ~v_700;
assign x_5869 = v_1859 | ~v_701;
assign x_5870 = ~v_1857 | ~v_1856 | ~v_1855 | v_1858;
assign x_5871 = v_1857 | ~v_1657;
assign x_5872 = v_1857 | ~v_682;
assign x_5873 = v_1857 | ~v_683;
assign x_5874 = v_1857 | ~v_906;
assign x_5875 = v_1857 | ~v_907;
assign x_5876 = v_1857 | ~v_1625;
assign x_5877 = v_1857 | ~v_1626;
assign x_5878 = v_1857 | ~v_1627;
assign x_5879 = v_1857 | ~v_1628;
assign x_5880 = v_1857 | ~v_1658;
assign x_5881 = v_1857 | ~v_1323;
assign x_5882 = v_1857 | ~v_1324;
assign x_5883 = v_1857 | ~v_1325;
assign x_5884 = v_1857 | ~v_1659;
assign x_5885 = v_1857 | ~v_1660;
assign x_5886 = v_1857 | ~v_1631;
assign x_5887 = v_1857 | ~v_1326;
assign x_5888 = v_1857 | ~v_1634;
assign x_5889 = v_1857 | ~v_113;
assign x_5890 = v_1857 | ~v_112;
assign x_5891 = v_1857 | ~v_106;
assign x_5892 = v_1857 | ~v_105;
assign x_5893 = v_1857 | ~v_76;
assign x_5894 = v_1857 | ~v_75;
assign x_5895 = v_1857 | ~v_74;
assign x_5896 = v_1857 | ~v_73;
assign x_5897 = v_1857 | ~v_69;
assign x_5898 = v_1856 | ~v_1648;
assign x_5899 = v_1856 | ~v_1649;
assign x_5900 = v_1856 | ~v_1614;
assign x_5901 = v_1856 | ~v_1615;
assign x_5902 = v_1856 | ~v_1616;
assign x_5903 = v_1856 | ~v_1617;
assign x_5904 = v_1856 | ~v_1318;
assign x_5905 = v_1856 | ~v_1650;
assign x_5906 = v_1856 | ~v_1651;
assign x_5907 = v_1856 | ~v_1620;
assign x_5908 = v_1856 | ~v_1621;
assign x_5909 = v_1856 | ~v_1319;
assign x_5910 = v_1856 | ~v_900;
assign x_5911 = v_1856 | ~v_677;
assign x_5912 = v_1856 | ~v_902;
assign x_5913 = v_1856 | ~v_1320;
assign x_5914 = v_1856 | ~v_678;
assign x_5915 = v_1856 | ~v_1321;
assign x_5916 = v_1856 | ~v_111;
assign x_5917 = v_1856 | ~v_110;
assign x_5918 = v_1856 | ~v_102;
assign x_5919 = v_1856 | ~v_101;
assign x_5920 = v_1856 | ~v_51;
assign x_5921 = v_1856 | ~v_50;
assign x_5922 = v_1856 | ~v_49;
assign x_5923 = v_1856 | ~v_48;
assign x_5924 = v_1856 | ~v_44;
assign x_5925 = v_1855 | ~v_1639;
assign x_5926 = v_1855 | ~v_1640;
assign x_5927 = v_1855 | ~v_646;
assign x_5928 = v_1855 | ~v_885;
assign x_5929 = v_1855 | ~v_1603;
assign x_5930 = v_1855 | ~v_1604;
assign x_5931 = v_1855 | ~v_1605;
assign x_5932 = v_1855 | ~v_1606;
assign x_5933 = v_1855 | ~v_1313;
assign x_5934 = v_1855 | ~v_1314;
assign x_5935 = v_1855 | ~v_1641;
assign x_5936 = v_1855 | ~v_1609;
assign x_5937 = v_1855 | ~v_1315;
assign x_5938 = v_1855 | ~v_661;
assign x_5939 = v_1855 | ~v_890;
assign x_5940 = v_1855 | ~v_1316;
assign x_5941 = v_1855 | ~v_1644;
assign x_5942 = v_1855 | ~v_1612;
assign x_5943 = v_1855 | ~v_109;
assign x_5944 = v_1855 | ~v_108;
assign x_5945 = v_1855 | ~v_95;
assign x_5946 = v_1855 | ~v_94;
assign x_5947 = v_1855 | ~v_25;
assign x_5948 = v_1855 | ~v_24;
assign x_5949 = v_1855 | ~v_23;
assign x_5950 = v_1855 | ~v_22;
assign x_5951 = v_1855 | ~v_18;
assign x_5952 = ~v_1601 | ~v_1853 | v_1854;
assign x_5953 = v_1853 | ~v_1827;
assign x_5954 = v_1853 | ~v_1842;
assign x_5955 = v_1853 | ~v_1848;
assign x_5956 = v_1853 | ~v_1852;
assign x_5957 = ~v_1522 | ~v_1851 | v_1852;
assign x_5958 = v_1851 | ~v_1849;
assign x_5959 = v_1851 | ~v_1833;
assign x_5960 = v_1851 | ~v_1834;
assign x_5961 = v_1851 | ~v_1850;
assign x_5962 = v_1851 | ~v_1835;
assign x_5963 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1552 | ~v_1844 | v_1850;
assign x_5964 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1539 | ~v_1831 | v_1849;
assign x_5965 = ~v_1847 | ~v_1843 | v_1848;
assign x_5966 = v_1847 | ~v_1845;
assign x_5967 = v_1847 | ~v_1846;
assign x_5968 = v_1847 | ~v_1828;
assign x_5969 = v_1847 | ~v_1829;
assign x_5970 = v_1847 | ~v_1830;
assign x_5971 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1498 | ~v_1836 | v_1846;
assign x_5972 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1477 | ~v_1844 | v_1845;
assign x_5973 = v_1844 | ~v_1838;
assign x_5974 = v_1844 | ~v_1839;
assign x_5975 = v_1844 | ~v_1840;
assign x_5976 = v_1843 | ~v_1581;
assign x_5977 = v_1843 | ~v_1582;
assign x_5978 = v_1843 | ~v_1523;
assign x_5979 = v_1843 | ~v_1540;
assign x_5980 = v_1843 | ~v_1541;
assign x_5981 = ~v_1841 | ~v_1575 | v_1842;
assign x_5982 = v_1841 | ~v_1832;
assign x_5983 = v_1841 | ~v_1837;
assign x_5984 = v_1841 | ~v_1838;
assign x_5985 = v_1841 | ~v_1839;
assign x_5986 = v_1841 | ~v_1840;
assign x_5987 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1509 | v_1840;
assign x_5988 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1493 | ~v_1546 | v_1839;
assign x_5989 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1514 | ~v_1444 | v_1838;
assign x_5990 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1493 | ~v_1836 | v_1837;
assign x_5991 = v_1836 | ~v_1833;
assign x_5992 = v_1836 | ~v_1834;
assign x_5993 = v_1836 | ~v_1835;
assign x_5994 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1546 | v_1835;
assign x_5995 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1509 | ~v_1552 | v_1834;
assign x_5996 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1444 | ~v_1539 | v_1833;
assign x_5997 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1514 | ~v_1831 | v_1832;
assign x_5998 = v_1831 | ~v_1828;
assign x_5999 = v_1831 | ~v_1829;
assign x_6000 = v_1831 | ~v_1830;
assign x_6001 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1444 | v_1830;
assign x_6002 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1498 | ~v_1546 | v_1829;
assign x_6003 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1509 | ~v_1477 | v_1828;
assign x_6004 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1826 | v_1827;
assign x_6005 = v_1826 | ~v_1823;
assign x_6006 = v_1826 | ~v_1824;
assign x_6007 = v_1826 | ~v_1825;
assign x_6008 = v_76 | v_69 | v_75 | v_74 | v_73 | v_106 | v_105 | v_113 | v_112 | ~v_1414 | ~v_1306 | ~v_1411 | ~v_1440 | ~v_1439 | ~v_1305 | ~v_1304 | ~v_1303 | ~v_1438 | ~v_1408 | ~v_1407 | ~v_1406 | ~v_1405 | ~v_454 | ~v_453 | ~v_230 | ~v_229 | ~v_1437 | v_1825;
assign x_6009 = v_50 | v_51 | v_49 | v_48 | v_44 | v_101 | v_102 | v_111 | v_110 | ~v_1301 | ~v_225 | ~v_1300 | ~v_449 | ~v_224 | ~v_447 | ~v_1299 | ~v_1401 | ~v_1400 | ~v_1431 | ~v_1430 | ~v_1298 | ~v_1397 | ~v_1396 | ~v_1395 | ~v_1394 | ~v_1429 | ~v_1428 | v_1824;
assign x_6010 = v_25 | v_24 | v_23 | v_22 | v_18 | v_95 | v_94 | v_108 | v_109 | ~v_1392 | ~v_1424 | ~v_1296 | ~v_437 | ~v_208 | ~v_1295 | ~v_1389 | ~v_1421 | ~v_1294 | ~v_1293 | ~v_1386 | ~v_1385 | ~v_1384 | ~v_1383 | ~v_432 | ~v_193 | ~v_1420 | ~v_1419 | v_1823;
assign x_6011 = v_7 | v_4 | v_6 | v_8 | v_10 | v_2 | v_1 | ~v_1041 | ~v_1040 | ~v_1821 | v_1822;
assign x_6012 = v_1821 | ~v_1602;
assign x_6013 = v_1821 | ~v_1820;
assign x_6014 = v_116 | ~v_1819 | ~v_1811 | ~v_1006 | ~v_1761 | ~v_1760 | ~v_1743 | ~v_1802 | ~v_1801 | ~v_1800 | ~v_1781 | v_1820;
assign x_6015 = v_1819 | ~v_1814;
assign x_6016 = v_1819 | ~v_1818;
assign x_6017 = v_115 | ~v_1029 | ~v_1028 | ~v_1817 | ~v_1816 | v_1818;
assign x_6018 = v_1817 | ~v_1034;
assign x_6019 = v_1817 | v_118;
assign x_6020 = v_1816 | ~v_1815;
assign x_6021 = v_1816 | v_133;
assign x_6022 = v_124 | ~v_1027 | ~v_1026 | v_1815;
assign x_6023 = v_114 | ~v_1000 | ~v_999 | ~v_1813 | ~v_1812 | v_1814;
assign x_6024 = v_1813 | ~v_997;
assign x_6025 = v_1813 | v_97;
assign x_6026 = v_1812 | ~v_1803;
assign x_6027 = v_1812 | v_123;
assign x_6028 = v_1811 | ~v_1806;
assign x_6029 = v_1811 | ~v_1810;
assign x_6030 = v_118 | ~v_1016 | ~v_1015 | ~v_1809 | ~v_1808 | v_1810;
assign x_6031 = v_1809 | ~v_1013;
assign x_6032 = v_1809 | v_115;
assign x_6033 = v_1808 | ~v_1807;
assign x_6034 = v_1808 | v_133;
assign x_6035 = v_129 | ~v_1020 | ~v_1019 | v_1807;
assign x_6036 = v_119 | ~v_996 | ~v_995 | ~v_1805 | ~v_1804 | v_1806;
assign x_6037 = v_1805 | ~v_1001;
assign x_6038 = v_1805 | v_98;
assign x_6039 = v_1804 | ~v_1803;
assign x_6040 = v_1804 | v_130;
assign x_6041 = v_134 | ~v_1004 | ~v_1003 | v_1803;
assign x_6042 = v_1802 | ~v_1777;
assign x_6043 = v_1802 | ~v_1725;
assign x_6044 = v_1802 | ~v_698;
assign x_6045 = v_1802 | ~v_699;
assign x_6046 = v_1802 | ~v_700;
assign x_6047 = v_1802 | ~v_701;
assign x_6048 = v_1801 | ~v_1797;
assign x_6049 = v_1801 | ~v_1680;
assign x_6050 = v_1801 | ~v_698;
assign x_6051 = v_1801 | ~v_699;
assign x_6052 = v_1801 | ~v_700;
assign x_6053 = v_1801 | ~v_701;
assign x_6054 = v_1800 | ~v_1795;
assign x_6055 = v_1800 | ~v_1799;
assign x_6056 = ~v_1776 | ~v_1775 | ~v_1774 | ~v_1798 | ~v_1796 | v_1799;
assign x_6057 = v_1798 | ~v_1797;
assign x_6058 = v_1798 | ~v_1713;
assign x_6059 = v_1798 | ~v_698;
assign x_6060 = v_1798 | ~v_699;
assign x_6061 = v_1798 | ~v_700;
assign x_6062 = v_1798 | ~v_701;
assign x_6063 = ~v_1779 | ~v_1773 | ~v_1768 | v_1797;
assign x_6064 = v_1796 | ~v_1762;
assign x_6065 = v_1796 | ~v_1729;
assign x_6066 = v_1796 | ~v_698;
assign x_6067 = v_1796 | ~v_699;
assign x_6068 = v_1796 | ~v_700;
assign x_6069 = v_1796 | ~v_701;
assign x_6070 = ~v_1794 | ~v_1793 | ~v_1792 | ~v_1791 | ~v_1786 | v_1795;
assign x_6071 = v_1794 | ~v_1725;
assign x_6072 = v_1794 | ~v_698;
assign x_6073 = v_1794 | ~v_699;
assign x_6074 = v_1794 | ~v_700;
assign x_6075 = v_1794 | ~v_701;
assign x_6076 = v_1793 | ~v_1772;
assign x_6077 = v_1793 | ~v_1680;
assign x_6078 = v_1793 | ~v_698;
assign x_6079 = v_1793 | ~v_699;
assign x_6080 = v_1793 | ~v_700;
assign x_6081 = v_1793 | ~v_701;
assign x_6082 = v_1792 | ~v_1636;
assign x_6083 = v_1792 | ~v_1697;
assign x_6084 = v_1792 | ~v_698;
assign x_6085 = v_1792 | ~v_699;
assign x_6086 = v_1792 | ~v_700;
assign x_6087 = v_1792 | ~v_701;
assign x_6088 = v_1791 | ~v_1790;
assign x_6089 = v_1791 | ~v_1636;
assign x_6090 = v_1791 | ~v_698;
assign x_6091 = v_1791 | ~v_699;
assign x_6092 = v_1791 | ~v_700;
assign x_6093 = v_1791 | ~v_701;
assign x_6094 = ~v_1789 | ~v_1788 | ~v_1787 | v_1790;
assign x_6095 = v_1789 | ~v_1697;
assign x_6096 = v_1789 | ~v_698;
assign x_6097 = v_1789 | ~v_699;
assign x_6098 = v_1789 | ~v_700;
assign x_6099 = v_1789 | ~v_701;
assign x_6100 = v_1788 | ~v_1772;
assign x_6101 = v_1788 | ~v_1718;
assign x_6102 = v_1788 | ~v_698;
assign x_6103 = v_1788 | ~v_699;
assign x_6104 = v_1788 | ~v_700;
assign x_6105 = v_1788 | ~v_701;
assign x_6106 = v_1787 | ~v_1725;
assign x_6107 = v_1787 | ~v_1664;
assign x_6108 = v_1787 | ~v_698;
assign x_6109 = v_1787 | ~v_699;
assign x_6110 = v_1787 | ~v_700;
assign x_6111 = v_1787 | ~v_701;
assign x_6112 = v_1786 | ~v_1785;
assign x_6113 = v_1786 | ~v_1680;
assign x_6114 = v_1786 | ~v_698;
assign x_6115 = v_1786 | ~v_699;
assign x_6116 = v_1786 | ~v_700;
assign x_6117 = v_1786 | ~v_701;
assign x_6118 = ~v_1784 | ~v_1783 | ~v_1782 | v_1785;
assign x_6119 = v_1784 | ~v_1772;
assign x_6120 = v_1784 | ~v_698;
assign x_6121 = v_1784 | ~v_699;
assign x_6122 = v_1784 | ~v_700;
assign x_6123 = v_1784 | ~v_701;
assign x_6124 = v_1783 | ~v_1759;
assign x_6125 = v_1783 | ~v_1697;
assign x_6126 = v_1783 | ~v_698;
assign x_6127 = v_1783 | ~v_699;
assign x_6128 = v_1783 | ~v_700;
assign x_6129 = v_1783 | ~v_701;
assign x_6130 = v_1782 | ~v_1766;
assign x_6131 = v_1782 | ~v_1725;
assign x_6132 = v_1782 | ~v_698;
assign x_6133 = v_1782 | ~v_699;
assign x_6134 = v_1782 | ~v_700;
assign x_6135 = v_1782 | ~v_701;
assign x_6136 = v_1781 | ~v_1742;
assign x_6137 = v_1781 | ~v_1780;
assign x_6138 = ~v_1779 | ~v_1778 | ~v_1773 | ~v_1768 | ~v_1767 | v_1780;
assign x_6139 = v_1779 | ~v_1759;
assign x_6140 = v_1779 | ~v_698;
assign x_6141 = v_1779 | ~v_699;
assign x_6142 = v_1779 | ~v_700;
assign x_6143 = v_1779 | ~v_701;
assign x_6144 = v_1778 | ~v_1777;
assign x_6145 = v_1778 | ~v_1772;
assign x_6146 = v_1778 | ~v_698;
assign x_6147 = v_1778 | ~v_699;
assign x_6148 = v_1778 | ~v_700;
assign x_6149 = v_1778 | ~v_701;
assign x_6150 = ~v_1776 | ~v_1775 | ~v_1774 | v_1777;
assign x_6151 = v_1776 | ~v_1734;
assign x_6152 = v_1776 | ~v_698;
assign x_6153 = v_1776 | ~v_699;
assign x_6154 = v_1776 | ~v_700;
assign x_6155 = v_1776 | ~v_701;
assign x_6156 = v_1775 | ~v_1759;
assign x_6157 = v_1775 | ~v_1713;
assign x_6158 = v_1775 | ~v_698;
assign x_6159 = v_1775 | ~v_699;
assign x_6160 = v_1775 | ~v_700;
assign x_6161 = v_1775 | ~v_701;
assign x_6162 = v_1774 | ~v_1636;
assign x_6163 = v_1774 | ~v_1729;
assign x_6164 = v_1774 | ~v_698;
assign x_6165 = v_1774 | ~v_699;
assign x_6166 = v_1774 | ~v_700;
assign x_6167 = v_1774 | ~v_701;
assign x_6168 = v_1773 | ~v_1772;
assign x_6169 = v_1773 | ~v_1734;
assign x_6170 = v_1773 | ~v_698;
assign x_6171 = v_1773 | ~v_699;
assign x_6172 = v_1773 | ~v_700;
assign x_6173 = v_1773 | ~v_701;
assign x_6174 = ~v_1771 | ~v_1770 | ~v_1769 | v_1772;
assign x_6175 = v_1771 | ~v_852;
assign x_6176 = v_1771 | ~v_853;
assign x_6177 = v_1771 | ~v_1625;
assign x_6178 = v_1771 | ~v_1626;
assign x_6179 = v_1771 | ~v_726;
assign x_6180 = v_1771 | ~v_634;
assign x_6181 = v_1771 | ~v_635;
assign x_6182 = v_1771 | ~v_1692;
assign x_6183 = v_1771 | ~v_1693;
assign x_6184 = v_1771 | ~v_854;
assign x_6185 = v_1771 | ~v_855;
assign x_6186 = v_1771 | ~v_1754;
assign x_6187 = v_1771 | ~v_1755;
assign x_6188 = v_1771 | ~v_1756;
assign x_6189 = v_1771 | ~v_731;
assign x_6190 = v_1771 | ~v_1694;
assign x_6191 = v_1771 | ~v_1695;
assign x_6192 = v_1771 | ~v_1757;
assign x_6193 = v_1771 | ~v_127;
assign x_6194 = v_1771 | ~v_112;
assign x_6195 = v_1771 | ~v_106;
assign x_6196 = v_1771 | ~v_105;
assign x_6197 = v_1771 | ~v_104;
assign x_6198 = v_1771 | ~v_76;
assign x_6199 = v_1771 | ~v_75;
assign x_6200 = v_1771 | ~v_73;
assign x_6201 = v_1771 | ~v_71;
assign x_6202 = v_1770 | ~v_847;
assign x_6203 = v_1770 | ~v_848;
assign x_6204 = v_1770 | ~v_1614;
assign x_6205 = v_1770 | ~v_1615;
assign x_6206 = v_1770 | ~v_714;
assign x_6207 = v_1770 | ~v_615;
assign x_6208 = v_1770 | ~v_616;
assign x_6209 = v_1770 | ~v_1687;
assign x_6210 = v_1770 | ~v_1688;
assign x_6211 = v_1770 | ~v_849;
assign x_6212 = v_1770 | ~v_850;
assign x_6213 = v_1770 | ~v_1749;
assign x_6214 = v_1770 | ~v_1750;
assign x_6215 = v_1770 | ~v_1751;
assign x_6216 = v_1770 | ~v_1752;
assign x_6217 = v_1770 | ~v_1689;
assign x_6218 = v_1770 | ~v_1690;
assign x_6219 = v_1770 | ~v_721;
assign x_6220 = v_1770 | ~v_126;
assign x_6221 = v_1770 | ~v_110;
assign x_6222 = v_1770 | ~v_102;
assign x_6223 = v_1770 | ~v_101;
assign x_6224 = v_1770 | ~v_100;
assign x_6225 = v_1770 | ~v_51;
assign x_6226 = v_1770 | ~v_50;
assign x_6227 = v_1770 | ~v_48;
assign x_6228 = v_1770 | ~v_46;
assign x_6229 = v_1769 | ~v_842;
assign x_6230 = v_1769 | ~v_843;
assign x_6231 = v_1769 | ~v_1603;
assign x_6232 = v_1769 | ~v_1604;
assign x_6233 = v_1769 | ~v_705;
assign x_6234 = v_1769 | ~v_706;
assign x_6235 = v_1769 | ~v_596;
assign x_6236 = v_1769 | ~v_597;
assign x_6237 = v_1769 | ~v_1682;
assign x_6238 = v_1769 | ~v_1683;
assign x_6239 = v_1769 | ~v_844;
assign x_6240 = v_1769 | ~v_845;
assign x_6241 = v_1769 | ~v_1744;
assign x_6242 = v_1769 | ~v_1745;
assign x_6243 = v_1769 | ~v_1746;
assign x_6244 = v_1769 | ~v_1684;
assign x_6245 = v_1769 | ~v_1685;
assign x_6246 = v_1769 | ~v_1747;
assign x_6247 = v_1769 | ~v_122;
assign x_6248 = v_1769 | ~v_108;
assign x_6249 = v_1769 | ~v_95;
assign x_6250 = v_1769 | ~v_94;
assign x_6251 = v_1769 | ~v_93;
assign x_6252 = v_1769 | ~v_25;
assign x_6253 = v_1769 | ~v_24;
assign x_6254 = v_1769 | ~v_22;
assign x_6255 = v_1769 | ~v_20;
assign x_6256 = v_1768 | ~v_1766;
assign x_6257 = v_1768 | ~v_1636;
assign x_6258 = v_1768 | ~v_698;
assign x_6259 = v_1768 | ~v_699;
assign x_6260 = v_1768 | ~v_700;
assign x_6261 = v_1768 | ~v_701;
assign x_6262 = v_1767 | ~v_1762;
assign x_6263 = v_1767 | ~v_1766;
assign x_6264 = v_1767 | ~v_698;
assign x_6265 = v_1767 | ~v_699;
assign x_6266 = v_1767 | ~v_700;
assign x_6267 = v_1767 | ~v_701;
assign x_6268 = ~v_1765 | ~v_1764 | ~v_1763 | v_1766;
assign x_6269 = v_1765 | ~v_1657;
assign x_6270 = v_1765 | ~v_682;
assign x_6271 = v_1765 | ~v_683;
assign x_6272 = v_1765 | ~v_1625;
assign x_6273 = v_1765 | ~v_1626;
assign x_6274 = v_1765 | ~v_1658;
assign x_6275 = v_1765 | ~v_725;
assign x_6276 = v_1765 | ~v_726;
assign x_6277 = v_1765 | ~v_727;
assign x_6278 = v_1765 | ~v_728;
assign x_6279 = v_1765 | ~v_1659;
assign x_6280 = v_1765 | ~v_1660;
assign x_6281 = v_1765 | ~v_1754;
assign x_6282 = v_1765 | ~v_1755;
assign x_6283 = v_1765 | ~v_1756;
assign x_6284 = v_1765 | ~v_731;
assign x_6285 = v_1765 | ~v_734;
assign x_6286 = v_1765 | ~v_1757;
assign x_6287 = v_1765 | ~v_112;
assign x_6288 = v_1765 | ~v_107;
assign x_6289 = v_1765 | ~v_106;
assign x_6290 = v_1765 | ~v_105;
assign x_6291 = v_1765 | ~v_104;
assign x_6292 = v_1765 | ~v_76;
assign x_6293 = v_1765 | ~v_74;
assign x_6294 = v_1765 | ~v_73;
assign x_6295 = v_1765 | ~v_71;
assign x_6296 = v_1764 | ~v_1648;
assign x_6297 = v_1764 | ~v_1649;
assign x_6298 = v_1764 | ~v_1614;
assign x_6299 = v_1764 | ~v_1615;
assign x_6300 = v_1764 | ~v_714;
assign x_6301 = v_1764 | ~v_715;
assign x_6302 = v_1764 | ~v_1650;
assign x_6303 = v_1764 | ~v_1651;
assign x_6304 = v_1764 | ~v_1749;
assign x_6305 = v_1764 | ~v_1750;
assign x_6306 = v_1764 | ~v_1751;
assign x_6307 = v_1764 | ~v_1752;
assign x_6308 = v_1764 | ~v_718;
assign x_6309 = v_1764 | ~v_721;
assign x_6310 = v_1764 | ~v_677;
assign x_6311 = v_1764 | ~v_722;
assign x_6312 = v_1764 | ~v_678;
assign x_6313 = v_1764 | ~v_723;
assign x_6314 = v_1764 | ~v_110;
assign x_6315 = v_1764 | ~v_103;
assign x_6316 = v_1764 | ~v_102;
assign x_6317 = v_1764 | ~v_101;
assign x_6318 = v_1764 | ~v_100;
assign x_6319 = v_1764 | ~v_51;
assign x_6320 = v_1764 | ~v_49;
assign x_6321 = v_1764 | ~v_48;
assign x_6322 = v_1764 | ~v_46;
assign x_6323 = v_1763 | ~v_1639;
assign x_6324 = v_1763 | ~v_1640;
assign x_6325 = v_1763 | ~v_646;
assign x_6326 = v_1763 | ~v_1603;
assign x_6327 = v_1763 | ~v_1604;
assign x_6328 = v_1763 | ~v_703;
assign x_6329 = v_1763 | ~v_704;
assign x_6330 = v_1763 | ~v_705;
assign x_6331 = v_1763 | ~v_706;
assign x_6332 = v_1763 | ~v_1641;
assign x_6333 = v_1763 | ~v_1744;
assign x_6334 = v_1763 | ~v_1745;
assign x_6335 = v_1763 | ~v_1746;
assign x_6336 = v_1763 | ~v_661;
assign x_6337 = v_1763 | ~v_711;
assign x_6338 = v_1763 | ~v_712;
assign x_6339 = v_1763 | ~v_1644;
assign x_6340 = v_1763 | ~v_1747;
assign x_6341 = v_1763 | ~v_108;
assign x_6342 = v_1763 | ~v_96;
assign x_6343 = v_1763 | ~v_95;
assign x_6344 = v_1763 | ~v_94;
assign x_6345 = v_1763 | ~v_93;
assign x_6346 = v_1763 | ~v_25;
assign x_6347 = v_1763 | ~v_23;
assign x_6348 = v_1763 | ~v_22;
assign x_6349 = v_1763 | ~v_20;
assign x_6350 = ~v_1761 | ~v_1760 | ~v_1743 | v_1762;
assign x_6351 = v_1761 | ~v_1636;
assign x_6352 = v_1761 | ~v_698;
assign x_6353 = v_1761 | ~v_699;
assign x_6354 = v_1761 | ~v_700;
assign x_6355 = v_1761 | ~v_701;
assign x_6356 = v_1760 | ~v_1759;
assign x_6357 = v_1760 | ~v_1680;
assign x_6358 = v_1760 | ~v_698;
assign x_6359 = v_1760 | ~v_699;
assign x_6360 = v_1760 | ~v_700;
assign x_6361 = v_1760 | ~v_701;
assign x_6362 = ~v_1758 | ~v_1753 | ~v_1748 | v_1759;
assign x_6363 = v_1758 | ~v_835;
assign x_6364 = v_1758 | ~v_836;
assign x_6365 = v_1758 | ~v_814;
assign x_6366 = v_1758 | ~v_815;
assign x_6367 = v_1758 | ~v_837;
assign x_6368 = v_1758 | ~v_838;
assign x_6369 = v_1758 | ~v_1625;
assign x_6370 = v_1758 | ~v_1626;
assign x_6371 = v_1758 | ~v_726;
assign x_6372 = v_1758 | ~v_1629;
assign x_6373 = v_1758 | ~v_1630;
assign x_6374 = v_1758 | ~v_1754;
assign x_6375 = v_1758 | ~v_1755;
assign x_6376 = v_1758 | ~v_1756;
assign x_6377 = v_1758 | ~v_731;
assign x_6378 = v_1758 | ~v_1632;
assign x_6379 = v_1758 | ~v_1633;
assign x_6380 = v_1758 | ~v_1757;
assign x_6381 = v_1758 | ~v_112;
assign x_6382 = v_1758 | ~v_106;
assign x_6383 = v_1758 | ~v_104;
assign x_6384 = v_1758 | ~v_76;
assign x_6385 = v_1758 | ~v_75;
assign x_6386 = v_1758 | ~v_74;
assign x_6387 = v_1758 | ~v_73;
assign x_6388 = v_1758 | ~v_71;
assign x_6389 = v_1758 | ~v_70;
assign x_6390 = ~v_88 | ~v_114 | v_1757;
assign x_6391 = ~v_80 | v_114 | v_1756;
assign x_6392 = ~v_86 | ~v_115 | v_1755;
assign x_6393 = ~v_78 | v_115 | v_1754;
assign x_6394 = v_1753 | ~v_830;
assign x_6395 = v_1753 | ~v_831;
assign x_6396 = v_1753 | ~v_803;
assign x_6397 = v_1753 | ~v_804;
assign x_6398 = v_1753 | ~v_1614;
assign x_6399 = v_1753 | ~v_1615;
assign x_6400 = v_1753 | ~v_714;
assign x_6401 = v_1753 | ~v_1618;
assign x_6402 = v_1753 | ~v_1619;
assign x_6403 = v_1753 | ~v_1749;
assign x_6404 = v_1753 | ~v_1750;
assign x_6405 = v_1753 | ~v_1751;
assign x_6406 = v_1753 | ~v_1752;
assign x_6407 = v_1753 | ~v_832;
assign x_6408 = v_1753 | ~v_833;
assign x_6409 = v_1753 | ~v_1622;
assign x_6410 = v_1753 | ~v_1623;
assign x_6411 = v_1753 | ~v_721;
assign x_6412 = v_1753 | ~v_110;
assign x_6413 = v_1753 | ~v_102;
assign x_6414 = v_1753 | ~v_100;
assign x_6415 = v_1753 | ~v_51;
assign x_6416 = v_1753 | ~v_50;
assign x_6417 = v_1753 | ~v_49;
assign x_6418 = v_1753 | ~v_48;
assign x_6419 = v_1753 | ~v_46;
assign x_6420 = v_1753 | ~v_45;
assign x_6421 = ~v_63 | ~v_114 | v_1752;
assign x_6422 = ~v_55 | v_114 | v_1751;
assign x_6423 = ~v_61 | ~v_115 | v_1750;
assign x_6424 = ~v_53 | v_115 | v_1749;
assign x_6425 = v_1748 | ~v_825;
assign x_6426 = v_1748 | ~v_826;
assign x_6427 = v_1748 | ~v_792;
assign x_6428 = v_1748 | ~v_793;
assign x_6429 = v_1748 | ~v_1603;
assign x_6430 = v_1748 | ~v_1604;
assign x_6431 = v_1748 | ~v_705;
assign x_6432 = v_1748 | ~v_706;
assign x_6433 = v_1748 | ~v_1607;
assign x_6434 = v_1748 | ~v_1608;
assign x_6435 = v_1748 | ~v_1744;
assign x_6436 = v_1748 | ~v_1745;
assign x_6437 = v_1748 | ~v_1746;
assign x_6438 = v_1748 | ~v_827;
assign x_6439 = v_1748 | ~v_1610;
assign x_6440 = v_1748 | ~v_1611;
assign x_6441 = v_1748 | ~v_1747;
assign x_6442 = v_1748 | ~v_828;
assign x_6443 = v_1748 | ~v_108;
assign x_6444 = v_1748 | ~v_95;
assign x_6445 = v_1748 | ~v_93;
assign x_6446 = v_1748 | ~v_25;
assign x_6447 = v_1748 | ~v_24;
assign x_6448 = v_1748 | ~v_23;
assign x_6449 = v_1748 | ~v_22;
assign x_6450 = v_1748 | ~v_20;
assign x_6451 = v_1748 | ~v_19;
assign x_6452 = ~v_38 | ~v_114 | v_1747;
assign x_6453 = ~v_30 | v_114 | v_1746;
assign x_6454 = ~v_36 | ~v_115 | v_1745;
assign x_6455 = ~v_28 | v_115 | v_1744;
assign x_6456 = v_1743 | ~v_1725;
assign x_6457 = v_1743 | ~v_1734;
assign x_6458 = v_1743 | ~v_698;
assign x_6459 = v_1743 | ~v_699;
assign x_6460 = v_1743 | ~v_700;
assign x_6461 = v_1743 | ~v_701;
assign x_6462 = ~v_1741 | ~v_1740 | ~v_1739 | ~v_1738 | ~v_1721 | v_1742;
assign x_6463 = v_1741 | ~v_1680;
assign x_6464 = v_1741 | ~v_698;
assign x_6465 = v_1741 | ~v_699;
assign x_6466 = v_1741 | ~v_700;
assign x_6467 = v_1741 | ~v_701;
assign x_6468 = v_1740 | ~v_1636;
assign x_6469 = v_1740 | ~v_1718;
assign x_6470 = v_1740 | ~v_698;
assign x_6471 = v_1740 | ~v_699;
assign x_6472 = v_1740 | ~v_700;
assign x_6473 = v_1740 | ~v_701;
assign x_6474 = v_1739 | ~v_1725;
assign x_6475 = v_1739 | ~v_1713;
assign x_6476 = v_1739 | ~v_698;
assign x_6477 = v_1739 | ~v_699;
assign x_6478 = v_1739 | ~v_700;
assign x_6479 = v_1739 | ~v_701;
assign x_6480 = v_1738 | ~v_1725;
assign x_6481 = v_1738 | ~v_1737;
assign x_6482 = v_1738 | ~v_698;
assign x_6483 = v_1738 | ~v_699;
assign x_6484 = v_1738 | ~v_700;
assign x_6485 = v_1738 | ~v_701;
assign x_6486 = ~v_1736 | ~v_1735 | ~v_1730 | v_1737;
assign x_6487 = v_1736 | ~v_1713;
assign x_6488 = v_1736 | ~v_698;
assign x_6489 = v_1736 | ~v_699;
assign x_6490 = v_1736 | ~v_700;
assign x_6491 = v_1736 | ~v_701;
assign x_6492 = v_1735 | ~v_1718;
assign x_6493 = v_1735 | ~v_1734;
assign x_6494 = v_1735 | ~v_698;
assign x_6495 = v_1735 | ~v_699;
assign x_6496 = v_1735 | ~v_700;
assign x_6497 = v_1735 | ~v_701;
assign x_6498 = ~v_1733 | ~v_1732 | ~v_1731 | v_1734;
assign x_6499 = v_1733 | ~v_1708;
assign x_6500 = v_1733 | ~v_812;
assign x_6501 = v_1733 | ~v_813;
assign x_6502 = v_1733 | ~v_814;
assign x_6503 = v_1733 | ~v_815;
assign x_6504 = v_1733 | ~v_1625;
assign x_6505 = v_1733 | ~v_1626;
assign x_6506 = v_1733 | ~v_1629;
assign x_6507 = v_1733 | ~v_1630;
assign x_6508 = v_1733 | ~v_816;
assign x_6509 = v_1733 | ~v_817;
assign x_6510 = v_1733 | ~v_688;
assign x_6511 = v_1733 | ~v_689;
assign x_6512 = v_1733 | ~v_1709;
assign x_6513 = v_1733 | ~v_1710;
assign x_6514 = v_1733 | ~v_1632;
assign x_6515 = v_1733 | ~v_1633;
assign x_6516 = v_1733 | ~v_1711;
assign x_6517 = v_1733 | ~v_132;
assign x_6518 = v_1733 | ~v_121;
assign x_6519 = v_1733 | ~v_113;
assign x_6520 = v_1733 | ~v_112;
assign x_6521 = v_1733 | ~v_106;
assign x_6522 = v_1733 | ~v_104;
assign x_6523 = v_1733 | ~v_75;
assign x_6524 = v_1733 | ~v_74;
assign x_6525 = v_1733 | ~v_70;
assign x_6526 = v_1732 | ~v_1703;
assign x_6527 = v_1732 | ~v_1704;
assign x_6528 = v_1732 | ~v_801;
assign x_6529 = v_1732 | ~v_802;
assign x_6530 = v_1732 | ~v_803;
assign x_6531 = v_1732 | ~v_804;
assign x_6532 = v_1732 | ~v_1614;
assign x_6533 = v_1732 | ~v_1615;
assign x_6534 = v_1732 | ~v_1618;
assign x_6535 = v_1732 | ~v_1619;
assign x_6536 = v_1732 | ~v_805;
assign x_6537 = v_1732 | ~v_806;
assign x_6538 = v_1732 | ~v_669;
assign x_6539 = v_1732 | ~v_670;
assign x_6540 = v_1732 | ~v_1705;
assign x_6541 = v_1732 | ~v_1706;
assign x_6542 = v_1732 | ~v_1622;
assign x_6543 = v_1732 | ~v_1623;
assign x_6544 = v_1732 | ~v_131;
assign x_6545 = v_1732 | ~v_120;
assign x_6546 = v_1732 | ~v_111;
assign x_6547 = v_1732 | ~v_110;
assign x_6548 = v_1732 | ~v_102;
assign x_6549 = v_1732 | ~v_100;
assign x_6550 = v_1732 | ~v_50;
assign x_6551 = v_1732 | ~v_49;
assign x_6552 = v_1732 | ~v_45;
assign x_6553 = v_1731 | ~v_1698;
assign x_6554 = v_1731 | ~v_1699;
assign x_6555 = v_1731 | ~v_790;
assign x_6556 = v_1731 | ~v_791;
assign x_6557 = v_1731 | ~v_792;
assign x_6558 = v_1731 | ~v_793;
assign x_6559 = v_1731 | ~v_1603;
assign x_6560 = v_1731 | ~v_1604;
assign x_6561 = v_1731 | ~v_1607;
assign x_6562 = v_1731 | ~v_1608;
assign x_6563 = v_1731 | ~v_794;
assign x_6564 = v_1731 | ~v_795;
assign x_6565 = v_1731 | ~v_653;
assign x_6566 = v_1731 | ~v_654;
assign x_6567 = v_1731 | ~v_1700;
assign x_6568 = v_1731 | ~v_1701;
assign x_6569 = v_1731 | ~v_1610;
assign x_6570 = v_1731 | ~v_1611;
assign x_6571 = v_1731 | ~v_128;
assign x_6572 = v_1731 | ~v_117;
assign x_6573 = v_1731 | ~v_109;
assign x_6574 = v_1731 | ~v_108;
assign x_6575 = v_1731 | ~v_95;
assign x_6576 = v_1731 | ~v_93;
assign x_6577 = v_1731 | ~v_24;
assign x_6578 = v_1731 | ~v_23;
assign x_6579 = v_1731 | ~v_19;
assign x_6580 = v_1730 | ~v_1729;
assign x_6581 = v_1730 | ~v_1680;
assign x_6582 = v_1730 | ~v_698;
assign x_6583 = v_1730 | ~v_699;
assign x_6584 = v_1730 | ~v_700;
assign x_6585 = v_1730 | ~v_701;
assign x_6586 = ~v_1728 | ~v_1727 | ~v_1726 | v_1729;
assign x_6587 = v_1728 | ~v_1708;
assign x_6588 = v_1728 | ~v_680;
assign x_6589 = v_1728 | ~v_681;
assign x_6590 = v_1728 | ~v_1657;
assign x_6591 = v_1728 | ~v_682;
assign x_6592 = v_1728 | ~v_683;
assign x_6593 = v_1728 | ~v_1625;
assign x_6594 = v_1728 | ~v_1626;
assign x_6595 = v_1728 | ~v_1658;
assign x_6596 = v_1728 | ~v_686;
assign x_6597 = v_1728 | ~v_687;
assign x_6598 = v_1728 | ~v_1659;
assign x_6599 = v_1728 | ~v_1660;
assign x_6600 = v_1728 | ~v_688;
assign x_6601 = v_1728 | ~v_689;
assign x_6602 = v_1728 | ~v_1709;
assign x_6603 = v_1728 | ~v_1710;
assign x_6604 = v_1728 | ~v_1711;
assign x_6605 = v_1728 | ~v_132;
assign x_6606 = v_1728 | ~v_113;
assign x_6607 = v_1728 | ~v_112;
assign x_6608 = v_1728 | ~v_106;
assign x_6609 = v_1728 | ~v_105;
assign x_6610 = v_1728 | ~v_104;
assign x_6611 = v_1728 | ~v_76;
assign x_6612 = v_1728 | ~v_75;
assign x_6613 = v_1728 | ~v_74;
assign x_6614 = v_1727 | ~v_1703;
assign x_6615 = v_1727 | ~v_1704;
assign x_6616 = v_1727 | ~v_1648;
assign x_6617 = v_1727 | ~v_1649;
assign x_6618 = v_1727 | ~v_1614;
assign x_6619 = v_1727 | ~v_1615;
assign x_6620 = v_1727 | ~v_665;
assign x_6621 = v_1727 | ~v_666;
assign x_6622 = v_1727 | ~v_1650;
assign x_6623 = v_1727 | ~v_1651;
assign x_6624 = v_1727 | ~v_667;
assign x_6625 = v_1727 | ~v_668;
assign x_6626 = v_1727 | ~v_669;
assign x_6627 = v_1727 | ~v_670;
assign x_6628 = v_1727 | ~v_1705;
assign x_6629 = v_1727 | ~v_1706;
assign x_6630 = v_1727 | ~v_677;
assign x_6631 = v_1727 | ~v_678;
assign x_6632 = v_1727 | ~v_131;
assign x_6633 = v_1727 | ~v_111;
assign x_6634 = v_1727 | ~v_110;
assign x_6635 = v_1727 | ~v_102;
assign x_6636 = v_1727 | ~v_101;
assign x_6637 = v_1727 | ~v_100;
assign x_6638 = v_1727 | ~v_51;
assign x_6639 = v_1727 | ~v_50;
assign x_6640 = v_1727 | ~v_49;
assign x_6641 = v_1726 | ~v_1698;
assign x_6642 = v_1726 | ~v_1699;
assign x_6643 = v_1726 | ~v_1639;
assign x_6644 = v_1726 | ~v_1640;
assign x_6645 = v_1726 | ~v_646;
assign x_6646 = v_1726 | ~v_1603;
assign x_6647 = v_1726 | ~v_1604;
assign x_6648 = v_1726 | ~v_649;
assign x_6649 = v_1726 | ~v_650;
assign x_6650 = v_1726 | ~v_1641;
assign x_6651 = v_1726 | ~v_651;
assign x_6652 = v_1726 | ~v_652;
assign x_6653 = v_1726 | ~v_653;
assign x_6654 = v_1726 | ~v_654;
assign x_6655 = v_1726 | ~v_1700;
assign x_6656 = v_1726 | ~v_1701;
assign x_6657 = v_1726 | ~v_661;
assign x_6658 = v_1726 | ~v_1644;
assign x_6659 = v_1726 | ~v_128;
assign x_6660 = v_1726 | ~v_109;
assign x_6661 = v_1726 | ~v_108;
assign x_6662 = v_1726 | ~v_95;
assign x_6663 = v_1726 | ~v_94;
assign x_6664 = v_1726 | ~v_93;
assign x_6665 = v_1726 | ~v_25;
assign x_6666 = v_1726 | ~v_24;
assign x_6667 = v_1726 | ~v_23;
assign x_6668 = ~v_1724 | ~v_1723 | ~v_1722 | v_1725;
assign x_6669 = v_1724 | ~v_951;
assign x_6670 = v_1724 | ~v_952;
assign x_6671 = v_1724 | ~v_906;
assign x_6672 = v_1724 | ~v_907;
assign x_6673 = v_1724 | ~v_1625;
assign x_6674 = v_1724 | ~v_1626;
assign x_6675 = v_1724 | ~v_1627;
assign x_6676 = v_1724 | ~v_1628;
assign x_6677 = v_1724 | ~v_953;
assign x_6678 = v_1724 | ~v_954;
assign x_6679 = v_1724 | ~v_634;
assign x_6680 = v_1724 | ~v_635;
assign x_6681 = v_1724 | ~v_1692;
assign x_6682 = v_1724 | ~v_1693;
assign x_6683 = v_1724 | ~v_1631;
assign x_6684 = v_1724 | ~v_1694;
assign x_6685 = v_1724 | ~v_1695;
assign x_6686 = v_1724 | ~v_1634;
assign x_6687 = v_1724 | ~v_127;
assign x_6688 = v_1724 | ~v_113;
assign x_6689 = v_1724 | ~v_112;
assign x_6690 = v_1724 | ~v_106;
assign x_6691 = v_1724 | ~v_105;
assign x_6692 = v_1724 | ~v_104;
assign x_6693 = v_1724 | ~v_76;
assign x_6694 = v_1724 | ~v_75;
assign x_6695 = v_1724 | ~v_73;
assign x_6696 = v_1723 | ~v_946;
assign x_6697 = v_1723 | ~v_947;
assign x_6698 = v_1723 | ~v_1614;
assign x_6699 = v_1723 | ~v_1615;
assign x_6700 = v_1723 | ~v_1616;
assign x_6701 = v_1723 | ~v_1617;
assign x_6702 = v_1723 | ~v_948;
assign x_6703 = v_1723 | ~v_949;
assign x_6704 = v_1723 | ~v_615;
assign x_6705 = v_1723 | ~v_616;
assign x_6706 = v_1723 | ~v_1687;
assign x_6707 = v_1723 | ~v_1688;
assign x_6708 = v_1723 | ~v_1620;
assign x_6709 = v_1723 | ~v_1621;
assign x_6710 = v_1723 | ~v_1689;
assign x_6711 = v_1723 | ~v_1690;
assign x_6712 = v_1723 | ~v_900;
assign x_6713 = v_1723 | ~v_902;
assign x_6714 = v_1723 | ~v_126;
assign x_6715 = v_1723 | ~v_111;
assign x_6716 = v_1723 | ~v_110;
assign x_6717 = v_1723 | ~v_102;
assign x_6718 = v_1723 | ~v_101;
assign x_6719 = v_1723 | ~v_100;
assign x_6720 = v_1723 | ~v_51;
assign x_6721 = v_1723 | ~v_50;
assign x_6722 = v_1723 | ~v_48;
assign x_6723 = v_1722 | ~v_941;
assign x_6724 = v_1722 | ~v_942;
assign x_6725 = v_1722 | ~v_885;
assign x_6726 = v_1722 | ~v_1603;
assign x_6727 = v_1722 | ~v_1604;
assign x_6728 = v_1722 | ~v_1605;
assign x_6729 = v_1722 | ~v_1606;
assign x_6730 = v_1722 | ~v_943;
assign x_6731 = v_1722 | ~v_944;
assign x_6732 = v_1722 | ~v_596;
assign x_6733 = v_1722 | ~v_597;
assign x_6734 = v_1722 | ~v_1682;
assign x_6735 = v_1722 | ~v_1683;
assign x_6736 = v_1722 | ~v_1609;
assign x_6737 = v_1722 | ~v_1684;
assign x_6738 = v_1722 | ~v_1685;
assign x_6739 = v_1722 | ~v_890;
assign x_6740 = v_1722 | ~v_1612;
assign x_6741 = v_1722 | ~v_122;
assign x_6742 = v_1722 | ~v_109;
assign x_6743 = v_1722 | ~v_108;
assign x_6744 = v_1722 | ~v_95;
assign x_6745 = v_1722 | ~v_94;
assign x_6746 = v_1722 | ~v_93;
assign x_6747 = v_1722 | ~v_25;
assign x_6748 = v_1722 | ~v_24;
assign x_6749 = v_1722 | ~v_22;
assign x_6750 = v_1721 | ~v_1636;
assign x_6751 = v_1721 | ~v_1720;
assign x_6752 = v_1721 | ~v_698;
assign x_6753 = v_1721 | ~v_699;
assign x_6754 = v_1721 | ~v_700;
assign x_6755 = v_1721 | ~v_701;
assign x_6756 = ~v_1719 | ~v_1714 | ~v_1681 | v_1720;
assign x_6757 = v_1719 | ~v_1718;
assign x_6758 = v_1719 | ~v_698;
assign x_6759 = v_1719 | ~v_699;
assign x_6760 = v_1719 | ~v_700;
assign x_6761 = v_1719 | ~v_701;
assign x_6762 = ~v_1717 | ~v_1716 | ~v_1715 | v_1718;
assign x_6763 = v_1717 | ~v_1655;
assign x_6764 = v_1717 | ~v_1656;
assign x_6765 = v_1717 | ~v_1675;
assign x_6766 = v_1717 | ~v_1676;
assign x_6767 = v_1717 | ~v_761;
assign x_6768 = v_1717 | ~v_762;
assign x_6769 = v_1717 | ~v_1625;
assign x_6770 = v_1717 | ~v_1626;
assign x_6771 = v_1717 | ~v_763;
assign x_6772 = v_1717 | ~v_764;
assign x_6773 = v_1717 | ~v_765;
assign x_6774 = v_1717 | ~v_766;
assign x_6775 = v_1717 | ~v_1677;
assign x_6776 = v_1717 | ~v_1678;
assign x_6777 = v_1717 | ~v_632;
assign x_6778 = v_1717 | ~v_633;
assign x_6779 = v_1717 | ~v_1661;
assign x_6780 = v_1717 | ~v_1662;
assign x_6781 = v_1717 | ~v_113;
assign x_6782 = v_1717 | ~v_105;
assign x_6783 = v_1717 | ~v_104;
assign x_6784 = v_1717 | ~v_76;
assign x_6785 = v_1717 | ~v_75;
assign x_6786 = v_1717 | ~v_74;
assign x_6787 = v_1717 | ~v_73;
assign x_6788 = v_1717 | ~v_72;
assign x_6789 = v_1717 | ~v_68;
assign x_6790 = v_1716 | ~v_1646;
assign x_6791 = v_1716 | ~v_1647;
assign x_6792 = v_1716 | ~v_1670;
assign x_6793 = v_1716 | ~v_1671;
assign x_6794 = v_1716 | ~v_1614;
assign x_6795 = v_1716 | ~v_1615;
assign x_6796 = v_1716 | ~v_750;
assign x_6797 = v_1716 | ~v_751;
assign x_6798 = v_1716 | ~v_752;
assign x_6799 = v_1716 | ~v_1672;
assign x_6800 = v_1716 | ~v_1673;
assign x_6801 = v_1716 | ~v_613;
assign x_6802 = v_1716 | ~v_614;
assign x_6803 = v_1716 | ~v_753;
assign x_6804 = v_1716 | ~v_754;
assign x_6805 = v_1716 | ~v_1652;
assign x_6806 = v_1716 | ~v_1653;
assign x_6807 = v_1716 | ~v_757;
assign x_6808 = v_1716 | ~v_111;
assign x_6809 = v_1716 | ~v_101;
assign x_6810 = v_1716 | ~v_100;
assign x_6811 = v_1716 | ~v_51;
assign x_6812 = v_1716 | ~v_50;
assign x_6813 = v_1716 | ~v_49;
assign x_6814 = v_1716 | ~v_48;
assign x_6815 = v_1716 | ~v_47;
assign x_6816 = v_1716 | ~v_43;
assign x_6817 = v_1715 | ~v_1637;
assign x_6818 = v_1715 | ~v_1638;
assign x_6819 = v_1715 | ~v_1665;
assign x_6820 = v_1715 | ~v_1666;
assign x_6821 = v_1715 | ~v_1603;
assign x_6822 = v_1715 | ~v_1604;
assign x_6823 = v_1715 | ~v_739;
assign x_6824 = v_1715 | ~v_740;
assign x_6825 = v_1715 | ~v_741;
assign x_6826 = v_1715 | ~v_1667;
assign x_6827 = v_1715 | ~v_594;
assign x_6828 = v_1715 | ~v_595;
assign x_6829 = v_1715 | ~v_742;
assign x_6830 = v_1715 | ~v_743;
assign x_6831 = v_1715 | ~v_1642;
assign x_6832 = v_1715 | ~v_1643;
assign x_6833 = v_1715 | ~v_746;
assign x_6834 = v_1715 | ~v_1668;
assign x_6835 = v_1715 | ~v_109;
assign x_6836 = v_1715 | ~v_94;
assign x_6837 = v_1715 | ~v_93;
assign x_6838 = v_1715 | ~v_25;
assign x_6839 = v_1715 | ~v_24;
assign x_6840 = v_1715 | ~v_23;
assign x_6841 = v_1715 | ~v_22;
assign x_6842 = v_1715 | ~v_21;
assign x_6843 = v_1715 | ~v_17;
assign x_6844 = v_1714 | ~v_1697;
assign x_6845 = v_1714 | ~v_1713;
assign x_6846 = v_1714 | ~v_698;
assign x_6847 = v_1714 | ~v_699;
assign x_6848 = v_1714 | ~v_700;
assign x_6849 = v_1714 | ~v_701;
assign x_6850 = ~v_1712 | ~v_1707 | ~v_1702 | v_1713;
assign x_6851 = v_1712 | ~v_1675;
assign x_6852 = v_1712 | ~v_1676;
assign x_6853 = v_1712 | ~v_1708;
assign x_6854 = v_1712 | ~v_871;
assign x_6855 = v_1712 | ~v_872;
assign x_6856 = v_1712 | ~v_873;
assign x_6857 = v_1712 | ~v_874;
assign x_6858 = v_1712 | ~v_1625;
assign x_6859 = v_1712 | ~v_1626;
assign x_6860 = v_1712 | ~v_763;
assign x_6861 = v_1712 | ~v_764;
assign x_6862 = v_1712 | ~v_1677;
assign x_6863 = v_1712 | ~v_1678;
assign x_6864 = v_1712 | ~v_688;
assign x_6865 = v_1712 | ~v_689;
assign x_6866 = v_1712 | ~v_1709;
assign x_6867 = v_1712 | ~v_1710;
assign x_6868 = v_1712 | ~v_1711;
assign x_6869 = v_1712 | ~v_132;
assign x_6870 = v_1712 | ~v_113;
assign x_6871 = v_1712 | ~v_112;
assign x_6872 = v_1712 | ~v_105;
assign x_6873 = v_1712 | ~v_104;
assign x_6874 = v_1712 | ~v_76;
assign x_6875 = v_1712 | ~v_75;
assign x_6876 = v_1712 | ~v_74;
assign x_6877 = v_1712 | ~v_72;
assign x_6878 = ~v_88 | ~v_134 | v_1711;
assign x_6879 = ~v_86 | ~v_133 | v_1710;
assign x_6880 = ~v_78 | v_133 | v_1709;
assign x_6881 = ~v_80 | v_134 | v_1708;
assign x_6882 = v_1707 | ~v_1670;
assign x_6883 = v_1707 | ~v_1671;
assign x_6884 = v_1707 | ~v_1703;
assign x_6885 = v_1707 | ~v_1704;
assign x_6886 = v_1707 | ~v_866;
assign x_6887 = v_1707 | ~v_867;
assign x_6888 = v_1707 | ~v_1614;
assign x_6889 = v_1707 | ~v_1615;
assign x_6890 = v_1707 | ~v_750;
assign x_6891 = v_1707 | ~v_1672;
assign x_6892 = v_1707 | ~v_1673;
assign x_6893 = v_1707 | ~v_868;
assign x_6894 = v_1707 | ~v_669;
assign x_6895 = v_1707 | ~v_670;
assign x_6896 = v_1707 | ~v_869;
assign x_6897 = v_1707 | ~v_1705;
assign x_6898 = v_1707 | ~v_1706;
assign x_6899 = v_1707 | ~v_757;
assign x_6900 = v_1707 | ~v_131;
assign x_6901 = v_1707 | ~v_111;
assign x_6902 = v_1707 | ~v_110;
assign x_6903 = v_1707 | ~v_101;
assign x_6904 = v_1707 | ~v_100;
assign x_6905 = v_1707 | ~v_51;
assign x_6906 = v_1707 | ~v_50;
assign x_6907 = v_1707 | ~v_49;
assign x_6908 = v_1707 | ~v_47;
assign x_6909 = ~v_61 | ~v_133 | v_1706;
assign x_6910 = ~v_53 | v_133 | v_1705;
assign x_6911 = ~v_63 | ~v_134 | v_1704;
assign x_6912 = ~v_55 | v_134 | v_1703;
assign x_6913 = v_1702 | ~v_1665;
assign x_6914 = v_1702 | ~v_1666;
assign x_6915 = v_1702 | ~v_1698;
assign x_6916 = v_1702 | ~v_1699;
assign x_6917 = v_1702 | ~v_861;
assign x_6918 = v_1702 | ~v_862;
assign x_6919 = v_1702 | ~v_1603;
assign x_6920 = v_1702 | ~v_1604;
assign x_6921 = v_1702 | ~v_739;
assign x_6922 = v_1702 | ~v_1667;
assign x_6923 = v_1702 | ~v_653;
assign x_6924 = v_1702 | ~v_654;
assign x_6925 = v_1702 | ~v_863;
assign x_6926 = v_1702 | ~v_864;
assign x_6927 = v_1702 | ~v_1700;
assign x_6928 = v_1702 | ~v_1701;
assign x_6929 = v_1702 | ~v_746;
assign x_6930 = v_1702 | ~v_1668;
assign x_6931 = v_1702 | ~v_128;
assign x_6932 = v_1702 | ~v_109;
assign x_6933 = v_1702 | ~v_108;
assign x_6934 = v_1702 | ~v_94;
assign x_6935 = v_1702 | ~v_93;
assign x_6936 = v_1702 | ~v_25;
assign x_6937 = v_1702 | ~v_24;
assign x_6938 = v_1702 | ~v_23;
assign x_6939 = v_1702 | ~v_21;
assign x_6940 = ~v_36 | ~v_133 | v_1701;
assign x_6941 = ~v_28 | v_133 | v_1700;
assign x_6942 = ~v_38 | ~v_134 | v_1699;
assign x_6943 = ~v_30 | v_134 | v_1698;
assign x_6944 = ~v_1696 | ~v_1691 | ~v_1686 | v_1697;
assign x_6945 = v_1696 | ~v_1655;
assign x_6946 = v_1696 | ~v_1656;
assign x_6947 = v_1696 | ~v_630;
assign x_6948 = v_1696 | ~v_631;
assign x_6949 = v_1696 | ~v_1625;
assign x_6950 = v_1696 | ~v_1626;
assign x_6951 = v_1696 | ~v_632;
assign x_6952 = v_1696 | ~v_633;
assign x_6953 = v_1696 | ~v_634;
assign x_6954 = v_1696 | ~v_635;
assign x_6955 = v_1696 | ~v_1692;
assign x_6956 = v_1696 | ~v_1693;
assign x_6957 = v_1696 | ~v_636;
assign x_6958 = v_1696 | ~v_637;
assign x_6959 = v_1696 | ~v_1661;
assign x_6960 = v_1696 | ~v_1662;
assign x_6961 = v_1696 | ~v_1694;
assign x_6962 = v_1696 | ~v_1695;
assign x_6963 = v_1696 | ~v_127;
assign x_6964 = v_1696 | ~v_113;
assign x_6965 = v_1696 | ~v_107;
assign x_6966 = v_1696 | ~v_106;
assign x_6967 = v_1696 | ~v_105;
assign x_6968 = v_1696 | ~v_104;
assign x_6969 = v_1696 | ~v_76;
assign x_6970 = v_1696 | ~v_73;
assign x_6971 = v_1696 | ~v_68;
assign x_6972 = ~v_87 | ~v_133 | v_1695;
assign x_6973 = ~v_79 | v_133 | v_1694;
assign x_6974 = ~v_90 | ~v_134 | v_1693;
assign x_6975 = ~v_82 | v_134 | v_1692;
assign x_6976 = v_1691 | ~v_1646;
assign x_6977 = v_1691 | ~v_1647;
assign x_6978 = v_1691 | ~v_611;
assign x_6979 = v_1691 | ~v_612;
assign x_6980 = v_1691 | ~v_1614;
assign x_6981 = v_1691 | ~v_1615;
assign x_6982 = v_1691 | ~v_613;
assign x_6983 = v_1691 | ~v_614;
assign x_6984 = v_1691 | ~v_615;
assign x_6985 = v_1691 | ~v_616;
assign x_6986 = v_1691 | ~v_1687;
assign x_6987 = v_1691 | ~v_1688;
assign x_6988 = v_1691 | ~v_617;
assign x_6989 = v_1691 | ~v_618;
assign x_6990 = v_1691 | ~v_1652;
assign x_6991 = v_1691 | ~v_1653;
assign x_6992 = v_1691 | ~v_1689;
assign x_6993 = v_1691 | ~v_1690;
assign x_6994 = v_1691 | ~v_126;
assign x_6995 = v_1691 | ~v_111;
assign x_6996 = v_1691 | ~v_103;
assign x_6997 = v_1691 | ~v_102;
assign x_6998 = v_1691 | ~v_101;
assign x_6999 = v_1691 | ~v_100;
assign x_7000 = v_1691 | ~v_51;
assign x_7001 = v_1691 | ~v_48;
assign x_7002 = v_1691 | ~v_43;
assign x_7003 = ~v_62 | ~v_133 | v_1690;
assign x_7004 = ~v_54 | v_133 | v_1689;
assign x_7005 = ~v_65 | ~v_134 | v_1688;
assign x_7006 = ~v_57 | v_134 | v_1687;
assign x_7007 = v_1686 | ~v_1637;
assign x_7008 = v_1686 | ~v_1638;
assign x_7009 = v_1686 | ~v_592;
assign x_7010 = v_1686 | ~v_593;
assign x_7011 = v_1686 | ~v_1603;
assign x_7012 = v_1686 | ~v_1604;
assign x_7013 = v_1686 | ~v_594;
assign x_7014 = v_1686 | ~v_595;
assign x_7015 = v_1686 | ~v_596;
assign x_7016 = v_1686 | ~v_597;
assign x_7017 = v_1686 | ~v_1682;
assign x_7018 = v_1686 | ~v_1683;
assign x_7019 = v_1686 | ~v_598;
assign x_7020 = v_1686 | ~v_599;
assign x_7021 = v_1686 | ~v_1642;
assign x_7022 = v_1686 | ~v_1643;
assign x_7023 = v_1686 | ~v_1684;
assign x_7024 = v_1686 | ~v_1685;
assign x_7025 = v_1686 | ~v_122;
assign x_7026 = v_1686 | ~v_109;
assign x_7027 = v_1686 | ~v_96;
assign x_7028 = v_1686 | ~v_95;
assign x_7029 = v_1686 | ~v_94;
assign x_7030 = v_1686 | ~v_93;
assign x_7031 = v_1686 | ~v_25;
assign x_7032 = v_1686 | ~v_22;
assign x_7033 = v_1686 | ~v_17;
assign x_7034 = ~v_37 | ~v_133 | v_1685;
assign x_7035 = ~v_29 | v_133 | v_1684;
assign x_7036 = ~v_40 | ~v_134 | v_1683;
assign x_7037 = ~v_32 | v_134 | v_1682;
assign x_7038 = v_1681 | ~v_1664;
assign x_7039 = v_1681 | ~v_1680;
assign x_7040 = v_1681 | ~v_698;
assign x_7041 = v_1681 | ~v_699;
assign x_7042 = v_1681 | ~v_700;
assign x_7043 = v_1681 | ~v_701;
assign x_7044 = ~v_1679 | ~v_1674 | ~v_1669 | v_1680;
assign x_7045 = v_1679 | ~v_1675;
assign x_7046 = v_1679 | ~v_1676;
assign x_7047 = v_1679 | ~v_906;
assign x_7048 = v_1679 | ~v_907;
assign x_7049 = v_1679 | ~v_1625;
assign x_7050 = v_1679 | ~v_1626;
assign x_7051 = v_1679 | ~v_1627;
assign x_7052 = v_1679 | ~v_1628;
assign x_7053 = v_1679 | ~v_908;
assign x_7054 = v_1679 | ~v_909;
assign x_7055 = v_1679 | ~v_910;
assign x_7056 = v_1679 | ~v_763;
assign x_7057 = v_1679 | ~v_764;
assign x_7058 = v_1679 | ~v_1677;
assign x_7059 = v_1679 | ~v_1678;
assign x_7060 = v_1679 | ~v_1631;
assign x_7061 = v_1679 | ~v_914;
assign x_7062 = v_1679 | ~v_1634;
assign x_7063 = v_1679 | ~v_121;
assign x_7064 = v_1679 | ~v_113;
assign x_7065 = v_1679 | ~v_112;
assign x_7066 = v_1679 | ~v_105;
assign x_7067 = v_1679 | ~v_104;
assign x_7068 = v_1679 | ~v_75;
assign x_7069 = v_1679 | ~v_74;
assign x_7070 = v_1679 | ~v_73;
assign x_7071 = v_1679 | ~v_72;
assign x_7072 = ~v_90 | ~v_114 | v_1678;
assign x_7073 = ~v_82 | v_114 | v_1677;
assign x_7074 = ~v_87 | ~v_115 | v_1676;
assign x_7075 = ~v_79 | v_115 | v_1675;
assign x_7076 = v_1674 | ~v_1670;
assign x_7077 = v_1674 | ~v_1671;
assign x_7078 = v_1674 | ~v_1614;
assign x_7079 = v_1674 | ~v_1615;
assign x_7080 = v_1674 | ~v_1616;
assign x_7081 = v_1674 | ~v_1617;
assign x_7082 = v_1674 | ~v_896;
assign x_7083 = v_1674 | ~v_750;
assign x_7084 = v_1674 | ~v_1672;
assign x_7085 = v_1674 | ~v_1673;
assign x_7086 = v_1674 | ~v_1620;
assign x_7087 = v_1674 | ~v_1621;
assign x_7088 = v_1674 | ~v_897;
assign x_7089 = v_1674 | ~v_757;
assign x_7090 = v_1674 | ~v_900;
assign x_7091 = v_1674 | ~v_901;
assign x_7092 = v_1674 | ~v_902;
assign x_7093 = v_1674 | ~v_903;
assign x_7094 = v_1674 | ~v_120;
assign x_7095 = v_1674 | ~v_111;
assign x_7096 = v_1674 | ~v_110;
assign x_7097 = v_1674 | ~v_101;
assign x_7098 = v_1674 | ~v_100;
assign x_7099 = v_1674 | ~v_50;
assign x_7100 = v_1674 | ~v_49;
assign x_7101 = v_1674 | ~v_48;
assign x_7102 = v_1674 | ~v_47;
assign x_7103 = ~v_65 | ~v_114 | v_1673;
assign x_7104 = ~v_57 | v_114 | v_1672;
assign x_7105 = ~v_62 | ~v_115 | v_1671;
assign x_7106 = ~v_54 | v_115 | v_1670;
assign x_7107 = v_1669 | ~v_1665;
assign x_7108 = v_1669 | ~v_1666;
assign x_7109 = v_1669 | ~v_885;
assign x_7110 = v_1669 | ~v_1603;
assign x_7111 = v_1669 | ~v_1604;
assign x_7112 = v_1669 | ~v_1605;
assign x_7113 = v_1669 | ~v_1606;
assign x_7114 = v_1669 | ~v_886;
assign x_7115 = v_1669 | ~v_887;
assign x_7116 = v_1669 | ~v_739;
assign x_7117 = v_1669 | ~v_1667;
assign x_7118 = v_1669 | ~v_1609;
assign x_7119 = v_1669 | ~v_746;
assign x_7120 = v_1669 | ~v_890;
assign x_7121 = v_1669 | ~v_891;
assign x_7122 = v_1669 | ~v_892;
assign x_7123 = v_1669 | ~v_1612;
assign x_7124 = v_1669 | ~v_1668;
assign x_7125 = v_1669 | ~v_117;
assign x_7126 = v_1669 | ~v_109;
assign x_7127 = v_1669 | ~v_108;
assign x_7128 = v_1669 | ~v_94;
assign x_7129 = v_1669 | ~v_93;
assign x_7130 = v_1669 | ~v_24;
assign x_7131 = v_1669 | ~v_23;
assign x_7132 = v_1669 | ~v_22;
assign x_7133 = v_1669 | ~v_21;
assign x_7134 = ~v_32 | v_114 | v_1668;
assign x_7135 = ~v_40 | ~v_114 | v_1667;
assign x_7136 = ~v_37 | ~v_115 | v_1666;
assign x_7137 = ~v_29 | v_115 | v_1665;
assign x_7138 = ~v_1663 | ~v_1654 | ~v_1645 | v_1664;
assign x_7139 = v_1663 | ~v_1655;
assign x_7140 = v_1663 | ~v_1656;
assign x_7141 = v_1663 | ~v_1657;
assign x_7142 = v_1663 | ~v_782;
assign x_7143 = v_1663 | ~v_783;
assign x_7144 = v_1663 | ~v_682;
assign x_7145 = v_1663 | ~v_683;
assign x_7146 = v_1663 | ~v_1625;
assign x_7147 = v_1663 | ~v_1626;
assign x_7148 = v_1663 | ~v_1658;
assign x_7149 = v_1663 | ~v_632;
assign x_7150 = v_1663 | ~v_633;
assign x_7151 = v_1663 | ~v_784;
assign x_7152 = v_1663 | ~v_785;
assign x_7153 = v_1663 | ~v_1659;
assign x_7154 = v_1663 | ~v_1660;
assign x_7155 = v_1663 | ~v_1661;
assign x_7156 = v_1663 | ~v_1662;
assign x_7157 = v_1663 | ~v_121;
assign x_7158 = v_1663 | ~v_113;
assign x_7159 = v_1663 | ~v_106;
assign x_7160 = v_1663 | ~v_105;
assign x_7161 = v_1663 | ~v_104;
assign x_7162 = v_1663 | ~v_75;
assign x_7163 = v_1663 | ~v_74;
assign x_7164 = v_1663 | ~v_73;
assign x_7165 = v_1663 | ~v_68;
assign x_7166 = ~v_86 | ~v_116 | v_1662;
assign x_7167 = ~v_78 | v_116 | v_1661;
assign x_7168 = ~v_90 | ~v_119 | v_1660;
assign x_7169 = ~v_82 | v_119 | v_1659;
assign x_7170 = ~v_87 | ~v_118 | v_1658;
assign x_7171 = ~v_79 | v_118 | v_1657;
assign x_7172 = ~v_88 | ~v_116 | v_1656;
assign x_7173 = ~v_80 | v_116 | v_1655;
assign x_7174 = v_1654 | ~v_1646;
assign x_7175 = v_1654 | ~v_1647;
assign x_7176 = v_1654 | ~v_1648;
assign x_7177 = v_1654 | ~v_1649;
assign x_7178 = v_1654 | ~v_777;
assign x_7179 = v_1654 | ~v_778;
assign x_7180 = v_1654 | ~v_1614;
assign x_7181 = v_1654 | ~v_1615;
assign x_7182 = v_1654 | ~v_613;
assign x_7183 = v_1654 | ~v_614;
assign x_7184 = v_1654 | ~v_779;
assign x_7185 = v_1654 | ~v_780;
assign x_7186 = v_1654 | ~v_1650;
assign x_7187 = v_1654 | ~v_1651;
assign x_7188 = v_1654 | ~v_1652;
assign x_7189 = v_1654 | ~v_1653;
assign x_7190 = v_1654 | ~v_677;
assign x_7191 = v_1654 | ~v_678;
assign x_7192 = v_1654 | ~v_120;
assign x_7193 = v_1654 | ~v_111;
assign x_7194 = v_1654 | ~v_102;
assign x_7195 = v_1654 | ~v_101;
assign x_7196 = v_1654 | ~v_100;
assign x_7197 = v_1654 | ~v_50;
assign x_7198 = v_1654 | ~v_49;
assign x_7199 = v_1654 | ~v_48;
assign x_7200 = v_1654 | ~v_43;
assign x_7201 = ~v_61 | ~v_116 | v_1653;
assign x_7202 = ~v_53 | v_116 | v_1652;
assign x_7203 = ~v_65 | ~v_119 | v_1651;
assign x_7204 = ~v_57 | v_119 | v_1650;
assign x_7205 = ~v_62 | ~v_118 | v_1649;
assign x_7206 = ~v_54 | v_118 | v_1648;
assign x_7207 = ~v_63 | ~v_116 | v_1647;
assign x_7208 = ~v_55 | v_116 | v_1646;
assign x_7209 = v_1645 | ~v_1637;
assign x_7210 = v_1645 | ~v_1638;
assign x_7211 = v_1645 | ~v_1639;
assign x_7212 = v_1645 | ~v_1640;
assign x_7213 = v_1645 | ~v_772;
assign x_7214 = v_1645 | ~v_773;
assign x_7215 = v_1645 | ~v_646;
assign x_7216 = v_1645 | ~v_1603;
assign x_7217 = v_1645 | ~v_1604;
assign x_7218 = v_1645 | ~v_594;
assign x_7219 = v_1645 | ~v_595;
assign x_7220 = v_1645 | ~v_774;
assign x_7221 = v_1645 | ~v_775;
assign x_7222 = v_1645 | ~v_1641;
assign x_7223 = v_1645 | ~v_1642;
assign x_7224 = v_1645 | ~v_1643;
assign x_7225 = v_1645 | ~v_661;
assign x_7226 = v_1645 | ~v_1644;
assign x_7227 = v_1645 | ~v_117;
assign x_7228 = v_1645 | ~v_109;
assign x_7229 = v_1645 | ~v_95;
assign x_7230 = v_1645 | ~v_94;
assign x_7231 = v_1645 | ~v_93;
assign x_7232 = v_1645 | ~v_24;
assign x_7233 = v_1645 | ~v_23;
assign x_7234 = v_1645 | ~v_22;
assign x_7235 = v_1645 | ~v_17;
assign x_7236 = ~v_32 | v_119 | v_1644;
assign x_7237 = ~v_36 | ~v_116 | v_1643;
assign x_7238 = ~v_28 | v_116 | v_1642;
assign x_7239 = ~v_40 | ~v_119 | v_1641;
assign x_7240 = ~v_37 | ~v_118 | v_1640;
assign x_7241 = ~v_29 | v_118 | v_1639;
assign x_7242 = ~v_38 | ~v_116 | v_1638;
assign x_7243 = ~v_30 | v_116 | v_1637;
assign x_7244 = ~v_1635 | ~v_1624 | ~v_1613 | v_1636;
assign x_7245 = v_1635 | ~v_814;
assign x_7246 = v_1635 | ~v_815;
assign x_7247 = v_1635 | ~v_930;
assign x_7248 = v_1635 | ~v_931;
assign x_7249 = v_1635 | ~v_932;
assign x_7250 = v_1635 | ~v_933;
assign x_7251 = v_1635 | ~v_906;
assign x_7252 = v_1635 | ~v_907;
assign x_7253 = v_1635 | ~v_1625;
assign x_7254 = v_1635 | ~v_1626;
assign x_7255 = v_1635 | ~v_1627;
assign x_7256 = v_1635 | ~v_1628;
assign x_7257 = v_1635 | ~v_1629;
assign x_7258 = v_1635 | ~v_1630;
assign x_7259 = v_1635 | ~v_1631;
assign x_7260 = v_1635 | ~v_1632;
assign x_7261 = v_1635 | ~v_1633;
assign x_7262 = v_1635 | ~v_1634;
assign x_7263 = v_1635 | ~v_113;
assign x_7264 = v_1635 | ~v_112;
assign x_7265 = v_1635 | ~v_107;
assign x_7266 = v_1635 | ~v_106;
assign x_7267 = v_1635 | ~v_104;
assign x_7268 = v_1635 | ~v_76;
assign x_7269 = v_1635 | ~v_74;
assign x_7270 = v_1635 | ~v_73;
assign x_7271 = v_1635 | ~v_70;
assign x_7272 = ~v_88 | ~v_119 | v_1634;
assign x_7273 = ~v_87 | ~v_116 | v_1633;
assign x_7274 = ~v_79 | v_116 | v_1632;
assign x_7275 = ~v_80 | v_119 | v_1631;
assign x_7276 = ~v_90 | ~v_116 | v_1630;
assign x_7277 = ~v_82 | v_116 | v_1629;
assign x_7278 = ~v_86 | ~v_118 | v_1628;
assign x_7279 = ~v_78 | v_118 | v_1627;
assign x_7280 = ~v_85 | ~v_116 | v_1626;
assign x_7281 = ~v_77 | v_116 | v_1625;
assign x_7282 = v_1624 | ~v_803;
assign x_7283 = v_1624 | ~v_804;
assign x_7284 = v_1624 | ~v_925;
assign x_7285 = v_1624 | ~v_926;
assign x_7286 = v_1624 | ~v_1614;
assign x_7287 = v_1624 | ~v_1615;
assign x_7288 = v_1624 | ~v_1616;
assign x_7289 = v_1624 | ~v_1617;
assign x_7290 = v_1624 | ~v_1618;
assign x_7291 = v_1624 | ~v_1619;
assign x_7292 = v_1624 | ~v_927;
assign x_7293 = v_1624 | ~v_928;
assign x_7294 = v_1624 | ~v_1620;
assign x_7295 = v_1624 | ~v_1621;
assign x_7296 = v_1624 | ~v_1622;
assign x_7297 = v_1624 | ~v_1623;
assign x_7298 = v_1624 | ~v_900;
assign x_7299 = v_1624 | ~v_902;
assign x_7300 = v_1624 | ~v_111;
assign x_7301 = v_1624 | ~v_110;
assign x_7302 = v_1624 | ~v_103;
assign x_7303 = v_1624 | ~v_102;
assign x_7304 = v_1624 | ~v_100;
assign x_7305 = v_1624 | ~v_51;
assign x_7306 = v_1624 | ~v_49;
assign x_7307 = v_1624 | ~v_48;
assign x_7308 = v_1624 | ~v_45;
assign x_7309 = ~v_62 | ~v_116 | v_1623;
assign x_7310 = ~v_54 | v_116 | v_1622;
assign x_7311 = ~v_63 | ~v_119 | v_1621;
assign x_7312 = ~v_55 | v_119 | v_1620;
assign x_7313 = ~v_65 | ~v_116 | v_1619;
assign x_7314 = ~v_57 | v_116 | v_1618;
assign x_7315 = ~v_61 | ~v_118 | v_1617;
assign x_7316 = ~v_53 | v_118 | v_1616;
assign x_7317 = ~v_60 | ~v_116 | v_1615;
assign x_7318 = ~v_52 | v_116 | v_1614;
assign x_7319 = v_1613 | ~v_792;
assign x_7320 = v_1613 | ~v_793;
assign x_7321 = v_1613 | ~v_920;
assign x_7322 = v_1613 | ~v_921;
assign x_7323 = v_1613 | ~v_885;
assign x_7324 = v_1613 | ~v_1603;
assign x_7325 = v_1613 | ~v_1604;
assign x_7326 = v_1613 | ~v_1605;
assign x_7327 = v_1613 | ~v_1606;
assign x_7328 = v_1613 | ~v_1607;
assign x_7329 = v_1613 | ~v_1608;
assign x_7330 = v_1613 | ~v_922;
assign x_7331 = v_1613 | ~v_1609;
assign x_7332 = v_1613 | ~v_1610;
assign x_7333 = v_1613 | ~v_1611;
assign x_7334 = v_1613 | ~v_890;
assign x_7335 = v_1613 | ~v_1612;
assign x_7336 = v_1613 | ~v_923;
assign x_7337 = v_1613 | ~v_109;
assign x_7338 = v_1613 | ~v_108;
assign x_7339 = v_1613 | ~v_96;
assign x_7340 = v_1613 | ~v_95;
assign x_7341 = v_1613 | ~v_93;
assign x_7342 = v_1613 | ~v_25;
assign x_7343 = v_1613 | ~v_23;
assign x_7344 = v_1613 | ~v_22;
assign x_7345 = v_1613 | ~v_19;
assign x_7346 = ~v_38 | ~v_119 | v_1612;
assign x_7347 = ~v_37 | ~v_116 | v_1611;
assign x_7348 = ~v_29 | v_116 | v_1610;
assign x_7349 = ~v_30 | v_119 | v_1609;
assign x_7350 = ~v_40 | ~v_116 | v_1608;
assign x_7351 = ~v_32 | v_116 | v_1607;
assign x_7352 = ~v_36 | ~v_118 | v_1606;
assign x_7353 = ~v_28 | v_118 | v_1605;
assign x_7354 = ~v_35 | ~v_116 | v_1604;
assign x_7355 = ~v_27 | v_116 | v_1603;
assign x_7356 = ~v_1601 | ~v_1583 | v_1602;
assign x_7357 = v_1601 | ~v_554;
assign x_7358 = v_1601 | ~v_1592;
assign x_7359 = v_1601 | ~v_1600;
assign x_7360 = v_1601 | ~v_116;
assign x_7361 = ~v_1599 | ~v_1595 | v_1600;
assign x_7362 = v_1599 | ~v_1597;
assign x_7363 = v_1599 | ~v_1598;
assign x_7364 = v_1599 | ~v_576;
assign x_7365 = v_1599 | ~v_577;
assign x_7366 = v_1599 | ~v_115;
assign x_7367 = ~v_118 | ~v_582 | v_1598;
assign x_7368 = ~v_133 | ~v_1596 | v_1597;
assign x_7369 = v_1596 | ~v_574;
assign x_7370 = v_1596 | ~v_575;
assign x_7371 = v_1596 | ~v_124;
assign x_7372 = v_1595 | ~v_1593;
assign x_7373 = v_1595 | ~v_1594;
assign x_7374 = v_1595 | ~v_547;
assign x_7375 = v_1595 | ~v_548;
assign x_7376 = v_1595 | ~v_114;
assign x_7377 = ~v_97 | ~v_545 | v_1594;
assign x_7378 = ~v_123 | ~v_1584 | v_1593;
assign x_7379 = ~v_1591 | ~v_1587 | v_1592;
assign x_7380 = v_1591 | ~v_1589;
assign x_7381 = v_1591 | ~v_1590;
assign x_7382 = v_1591 | ~v_563;
assign x_7383 = v_1591 | ~v_564;
assign x_7384 = v_1591 | ~v_118;
assign x_7385 = ~v_115 | ~v_561 | v_1590;
assign x_7386 = ~v_133 | ~v_1588 | v_1589;
assign x_7387 = v_1588 | ~v_567;
assign x_7388 = v_1588 | ~v_568;
assign x_7389 = v_1588 | ~v_129;
assign x_7390 = v_1587 | ~v_1585;
assign x_7391 = v_1587 | ~v_1586;
assign x_7392 = v_1587 | ~v_543;
assign x_7393 = v_1587 | ~v_544;
assign x_7394 = v_1587 | ~v_119;
assign x_7395 = ~v_98 | ~v_549 | v_1586;
assign x_7396 = ~v_130 | ~v_1584 | v_1585;
assign x_7397 = v_1584 | ~v_551;
assign x_7398 = v_1584 | ~v_552;
assign x_7399 = v_1584 | ~v_134;
assign x_7400 = v_1583 | ~v_1561;
assign x_7401 = v_1583 | ~v_1580;
assign x_7402 = v_1583 | ~v_1581;
assign x_7403 = v_1583 | ~v_1582;
assign x_7404 = v_1583 | ~v_1523;
assign x_7405 = v_1583 | ~v_1540;
assign x_7406 = v_1583 | ~v_1541;
assign x_7407 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1505 | ~v_1557 | v_1582;
assign x_7408 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1460 | ~v_1577 | v_1581;
assign x_7409 = ~v_1579 | ~v_1575 | v_1580;
assign x_7410 = v_1579 | ~v_1576;
assign x_7411 = v_1579 | ~v_1578;
assign x_7412 = v_1579 | ~v_1554;
assign x_7413 = v_1579 | ~v_1555;
assign x_7414 = v_1579 | ~v_1556;
assign x_7415 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1493 | ~v_1577 | v_1578;
assign x_7416 = v_1577 | ~v_1548;
assign x_7417 = v_1577 | ~v_1553;
assign x_7418 = v_1577 | ~v_1559;
assign x_7419 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1509 | ~v_1542 | v_1576;
assign x_7420 = v_1575 | ~v_1566;
assign x_7421 = v_1575 | ~v_1571;
assign x_7422 = v_1575 | ~v_1572;
assign x_7423 = v_1575 | ~v_1573;
assign x_7424 = v_1575 | ~v_1574;
assign x_7425 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1505 | v_1574;
assign x_7426 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1460 | ~v_1552 | v_1573;
assign x_7427 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1477 | ~v_1416 | v_1572;
assign x_7428 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1416 | ~v_1570 | v_1571;
assign x_7429 = v_1570 | ~v_1567;
assign x_7430 = v_1570 | ~v_1568;
assign x_7431 = v_1570 | ~v_1569;
assign x_7432 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1477 | v_1569;
assign x_7433 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1498 | ~v_1552 | v_1568;
assign x_7434 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1444 | ~v_1505 | v_1567;
assign x_7435 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1460 | ~v_1565 | v_1566;
assign x_7436 = v_1565 | ~v_1562;
assign x_7437 = v_1565 | ~v_1563;
assign x_7438 = v_1565 | ~v_1564;
assign x_7439 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1552 | v_1564;
assign x_7440 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1477 | ~v_1539 | v_1563;
assign x_7441 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1505 | ~v_1546 | v_1562;
assign x_7442 = ~v_1560 | ~v_1522 | v_1561;
assign x_7443 = v_1560 | ~v_1547;
assign x_7444 = v_1560 | ~v_1548;
assign x_7445 = v_1560 | ~v_1553;
assign x_7446 = v_1560 | ~v_1558;
assign x_7447 = v_1560 | ~v_1559;
assign x_7448 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1539 | v_1559;
assign x_7449 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1552 | ~v_1557 | v_1558;
assign x_7450 = v_1557 | ~v_1554;
assign x_7451 = v_1557 | ~v_1555;
assign x_7452 = v_1557 | ~v_1556;
assign x_7453 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1514 | v_1556;
assign x_7454 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1493 | ~v_1539 | v_1555;
assign x_7455 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1509 | ~v_1416 | v_1554;
assign x_7456 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1514 | ~v_1552 | v_1553;
assign x_7457 = v_1552 | ~v_1549;
assign x_7458 = v_1552 | ~v_1550;
assign x_7459 = v_1552 | ~v_1551;
assign x_7460 = v_76 | v_75 | v_73 | v_71 | v_106 | v_105 | v_104 | v_127 | v_112 | ~v_1537 | ~v_1475 | ~v_1474 | ~v_278 | ~v_1536 | ~v_1535 | ~v_1534 | ~v_402 | ~v_401 | ~v_1473 | ~v_1472 | ~v_182 | ~v_181 | ~v_273 | ~v_1406 | ~v_1405 | ~v_400 | ~v_399 | v_1551;
assign x_7461 = v_50 | v_51 | v_48 | v_46 | v_101 | v_100 | v_102 | v_110 | v_126 | ~v_268 | ~v_1470 | ~v_1469 | ~v_1532 | ~v_1531 | ~v_1530 | ~v_1529 | ~v_397 | ~v_396 | ~v_1468 | ~v_1467 | ~v_163 | ~v_162 | ~v_261 | ~v_1395 | ~v_1394 | ~v_395 | ~v_394 | v_1550;
assign x_7462 = v_25 | v_24 | v_22 | v_20 | v_95 | v_94 | v_93 | v_108 | v_122 | ~v_1527 | ~v_1465 | ~v_1464 | ~v_1526 | ~v_1525 | ~v_1524 | ~v_392 | ~v_391 | ~v_1463 | ~v_1462 | ~v_144 | ~v_143 | ~v_253 | ~v_252 | ~v_1384 | ~v_1383 | ~v_390 | ~v_389 | v_1549;
assign x_7463 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1416 | ~v_1546 | v_1548;
assign x_7464 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1546 | ~v_1542 | v_1547;
assign x_7465 = v_1546 | ~v_1543;
assign x_7466 = v_1546 | ~v_1544;
assign x_7467 = v_1546 | ~v_1545;
assign x_7468 = v_76 | v_74 | v_73 | v_71 | v_107 | v_106 | v_105 | v_104 | v_112 | ~v_1537 | ~v_281 | ~v_278 | ~v_1536 | ~v_1535 | ~v_1534 | ~v_1440 | ~v_1439 | ~v_275 | ~v_274 | ~v_273 | ~v_272 | ~v_1438 | ~v_1406 | ~v_1405 | ~v_230 | ~v_229 | ~v_1437 | v_1545;
assign x_7469 = v_51 | v_49 | v_48 | v_46 | v_103 | v_101 | v_100 | v_102 | v_110 | ~v_270 | ~v_225 | ~v_269 | ~v_224 | ~v_268 | ~v_265 | ~v_1532 | ~v_1531 | ~v_1530 | ~v_1529 | ~v_1431 | ~v_1430 | ~v_262 | ~v_261 | ~v_1395 | ~v_1394 | ~v_1429 | ~v_1428 | v_1544;
assign x_7470 = v_25 | v_23 | v_22 | v_20 | v_96 | v_95 | v_94 | v_93 | v_108 | ~v_1527 | ~v_1424 | ~v_259 | ~v_258 | ~v_208 | ~v_1526 | ~v_1525 | ~v_1524 | ~v_1421 | ~v_253 | ~v_252 | ~v_251 | ~v_250 | ~v_1384 | ~v_1383 | ~v_193 | ~v_1420 | ~v_1419 | v_1543;
assign x_7471 = v_1542 | ~v_1523;
assign x_7472 = v_1542 | ~v_1540;
assign x_7473 = v_1542 | ~v_1541;
assign x_7474 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1416 | v_1541;
assign x_7475 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1460 | ~v_1539 | v_1540;
assign x_7476 = v_1539 | ~v_1528;
assign x_7477 = v_1539 | ~v_1533;
assign x_7478 = v_1539 | ~v_1538;
assign x_7479 = v_76 | v_75 | v_74 | v_73 | v_71 | v_70 | v_106 | v_104 | v_112 | ~v_1537 | ~v_1413 | ~v_1412 | ~v_278 | ~v_1536 | ~v_1535 | ~v_1534 | ~v_1410 | ~v_1409 | ~v_273 | ~v_1406 | ~v_1405 | ~v_385 | ~v_384 | ~v_362 | ~v_361 | ~v_383 | ~v_382 | v_1538;
assign x_7480 = v_1537 | v_114;
assign x_7481 = v_1537 | v_88;
assign x_7482 = v_1536 | ~v_114;
assign x_7483 = v_1536 | v_80;
assign x_7484 = v_1535 | v_115;
assign x_7485 = v_1535 | v_86;
assign x_7486 = v_1534 | ~v_115;
assign x_7487 = v_1534 | v_78;
assign x_7488 = v_50 | v_51 | v_49 | v_48 | v_46 | v_45 | v_100 | v_102 | v_110 | ~v_268 | ~v_1403 | ~v_1402 | ~v_380 | ~v_379 | ~v_1532 | ~v_1531 | ~v_1530 | ~v_1529 | ~v_1399 | ~v_1398 | ~v_261 | ~v_1395 | ~v_1394 | ~v_351 | ~v_350 | ~v_378 | ~v_377 | v_1533;
assign x_7489 = v_1532 | v_114;
assign x_7490 = v_1532 | v_63;
assign x_7491 = v_1531 | ~v_114;
assign x_7492 = v_1531 | v_55;
assign x_7493 = v_1530 | v_115;
assign x_7494 = v_1530 | v_61;
assign x_7495 = v_1529 | ~v_115;
assign x_7496 = v_1529 | v_53;
assign x_7497 = v_25 | v_24 | v_23 | v_22 | v_20 | v_19 | v_95 | v_93 | v_108 | ~v_375 | ~v_1527 | ~v_1391 | ~v_1390 | ~v_374 | ~v_1526 | ~v_1525 | ~v_1524 | ~v_1388 | ~v_1387 | ~v_253 | ~v_252 | ~v_1384 | ~v_1383 | ~v_340 | ~v_339 | ~v_373 | ~v_372 | v_1528;
assign x_7498 = v_1527 | v_114;
assign x_7499 = v_1527 | v_38;
assign x_7500 = v_1526 | ~v_114;
assign x_7501 = v_1526 | v_30;
assign x_7502 = v_1525 | v_115;
assign x_7503 = v_1525 | v_36;
assign x_7504 = v_1524 | ~v_115;
assign x_7505 = v_1524 | v_28;
assign x_7506 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1514 | ~v_1505 | v_1523;
assign x_7507 = v_1522 | ~v_1501;
assign x_7508 = v_1522 | ~v_1518;
assign x_7509 = v_1522 | ~v_1519;
assign x_7510 = v_1522 | ~v_1520;
assign x_7511 = v_1522 | ~v_1521;
assign x_7512 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1460 | v_1521;
assign x_7513 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1498 | ~v_1416 | v_1520;
assign x_7514 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1493 | ~v_1505 | v_1519;
assign x_7515 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1517 | ~v_1505 | v_1518;
assign x_7516 = v_1517 | ~v_1510;
assign x_7517 = v_1517 | ~v_1515;
assign x_7518 = v_1517 | ~v_1516;
assign x_7519 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1493 | v_1516;
assign x_7520 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1514 | ~v_1498 | v_1515;
assign x_7521 = v_1514 | ~v_1511;
assign x_7522 = v_1514 | ~v_1512;
assign x_7523 = v_1514 | ~v_1513;
assign x_7524 = v_75 | v_74 | v_70 | v_106 | v_104 | v_132 | v_113 | v_112 | v_121 | ~v_1491 | ~v_1413 | ~v_1412 | ~v_1490 | ~v_1489 | ~v_236 | ~v_235 | ~v_364 | ~v_363 | ~v_1410 | ~v_1409 | ~v_1406 | ~v_1405 | ~v_362 | ~v_361 | ~v_360 | ~v_359 | ~v_1488 | v_1513;
assign x_7525 = v_50 | v_49 | v_45 | v_100 | v_102 | v_111 | v_110 | v_131 | v_120 | ~v_1403 | ~v_1402 | ~v_1486 | ~v_1485 | ~v_217 | ~v_216 | ~v_353 | ~v_352 | ~v_1399 | ~v_1398 | ~v_1395 | ~v_1394 | ~v_351 | ~v_350 | ~v_349 | ~v_348 | ~v_1484 | ~v_1483 | v_1512;
assign x_7526 = v_24 | v_23 | v_19 | v_95 | v_93 | v_108 | v_109 | v_128 | v_117 | ~v_1391 | ~v_1390 | ~v_1481 | ~v_1480 | ~v_201 | ~v_200 | ~v_342 | ~v_341 | ~v_1388 | ~v_1387 | ~v_1384 | ~v_1383 | ~v_340 | ~v_339 | ~v_338 | ~v_337 | ~v_1479 | ~v_1478 | v_1511;
assign x_7527 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1460 | ~v_1509 | v_1510;
assign x_7528 = v_1509 | ~v_1506;
assign x_7529 = v_1509 | ~v_1507;
assign x_7530 = v_1509 | ~v_1508;
assign x_7531 = v_76 | v_75 | v_74 | v_106 | v_105 | v_104 | v_132 | v_113 | v_112 | ~v_1491 | ~v_1490 | ~v_1489 | ~v_236 | ~v_235 | ~v_1440 | ~v_1439 | ~v_234 | ~v_233 | ~v_1438 | ~v_1406 | ~v_1405 | ~v_230 | ~v_229 | ~v_1437 | ~v_228 | ~v_227 | ~v_1488 | v_1508;
assign x_7532 = v_50 | v_51 | v_49 | v_101 | v_100 | v_102 | v_111 | v_110 | v_131 | ~v_225 | ~v_224 | ~v_1486 | ~v_1485 | ~v_217 | ~v_216 | ~v_215 | ~v_214 | ~v_1431 | ~v_1430 | ~v_213 | ~v_212 | ~v_1395 | ~v_1394 | ~v_1429 | ~v_1428 | ~v_1484 | ~v_1483 | v_1507;
assign x_7533 = v_25 | v_24 | v_23 | v_95 | v_94 | v_93 | v_108 | v_109 | v_128 | ~v_1424 | ~v_208 | ~v_1481 | ~v_1480 | ~v_201 | ~v_200 | ~v_199 | ~v_198 | ~v_1421 | ~v_197 | ~v_196 | ~v_1384 | ~v_1383 | ~v_193 | ~v_1420 | ~v_1419 | ~v_1479 | ~v_1478 | v_1506;
assign x_7534 = v_1505 | ~v_1502;
assign x_7535 = v_1505 | ~v_1503;
assign x_7536 = v_1505 | ~v_1504;
assign x_7537 = v_76 | v_75 | v_73 | v_106 | v_105 | v_104 | v_127 | v_113 | v_112 | ~v_1414 | ~v_1475 | ~v_1474 | ~v_1411 | ~v_1473 | ~v_1472 | ~v_182 | ~v_181 | ~v_501 | ~v_500 | ~v_1408 | ~v_1407 | ~v_1406 | ~v_1405 | ~v_454 | ~v_453 | ~v_499 | ~v_498 | v_1504;
assign x_7538 = v_50 | v_51 | v_48 | v_101 | v_100 | v_102 | v_111 | v_110 | v_126 | ~v_449 | ~v_447 | ~v_1470 | ~v_1469 | ~v_1401 | ~v_1400 | ~v_1468 | ~v_1467 | ~v_163 | ~v_162 | ~v_496 | ~v_495 | ~v_1397 | ~v_1396 | ~v_1395 | ~v_1394 | ~v_494 | ~v_493 | v_1503;
assign x_7539 = v_25 | v_24 | v_22 | v_95 | v_94 | v_93 | v_108 | v_109 | v_122 | ~v_1392 | ~v_437 | ~v_1465 | ~v_1464 | ~v_1389 | ~v_1463 | ~v_1462 | ~v_144 | ~v_143 | ~v_491 | ~v_490 | ~v_1386 | ~v_1385 | ~v_1384 | ~v_1383 | ~v_432 | ~v_489 | ~v_488 | v_1502;
assign x_7540 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1500 | ~v_1416 | v_1501;
assign x_7541 = v_1500 | ~v_1461;
assign x_7542 = v_1500 | ~v_1494;
assign x_7543 = v_1500 | ~v_1499;
assign x_7544 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1498 | v_1499;
assign x_7545 = v_1498 | ~v_1495;
assign x_7546 = v_1498 | ~v_1496;
assign x_7547 = v_1498 | ~v_1497;
assign x_7548 = v_76 | v_68 | v_75 | v_74 | v_73 | v_72 | v_105 | v_104 | v_113 | ~v_1442 | ~v_1441 | ~v_180 | ~v_179 | ~v_1458 | ~v_1457 | ~v_313 | ~v_312 | ~v_311 | ~v_310 | ~v_1406 | ~v_1405 | ~v_309 | ~v_308 | ~v_1456 | ~v_1455 | ~v_1436 | ~v_1435 | v_1497;
assign x_7549 = v_50 | v_51 | v_49 | v_48 | v_43 | v_47 | v_101 | v_100 | v_111 | ~v_304 | ~v_1433 | ~v_1432 | ~v_301 | ~v_300 | ~v_161 | ~v_160 | ~v_1453 | ~v_1452 | ~v_299 | ~v_298 | ~v_297 | ~v_1395 | ~v_1394 | ~v_1451 | ~v_1450 | ~v_1427 | ~v_1426 | v_1496;
assign x_7550 = v_25 | v_24 | v_23 | v_22 | v_21 | v_17 | v_94 | v_93 | v_109 | ~v_1448 | ~v_293 | ~v_1423 | ~v_1422 | ~v_290 | ~v_289 | ~v_142 | ~v_141 | ~v_1447 | ~v_288 | ~v_287 | ~v_286 | ~v_1384 | ~v_1383 | ~v_1446 | ~v_1445 | ~v_1418 | ~v_1417 | v_1495;
assign x_7551 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1493 | ~v_1477 | v_1494;
assign x_7552 = v_1493 | ~v_1482;
assign x_7553 = v_1493 | ~v_1487;
assign x_7554 = v_1493 | ~v_1492;
assign x_7555 = v_76 | v_75 | v_74 | v_72 | v_105 | v_104 | v_132 | v_113 | v_112 | ~v_1491 | ~v_1490 | ~v_1489 | ~v_236 | ~v_235 | ~v_1458 | ~v_1457 | ~v_311 | ~v_310 | ~v_1406 | ~v_1405 | ~v_421 | ~v_420 | ~v_419 | ~v_418 | ~v_1488 | ~v_1456 | ~v_1455 | v_1492;
assign x_7556 = v_1491 | v_134;
assign x_7557 = v_1491 | v_88;
assign x_7558 = v_1490 | v_133;
assign x_7559 = v_1490 | v_86;
assign x_7560 = v_1489 | ~v_133;
assign x_7561 = v_1489 | v_78;
assign x_7562 = v_1488 | ~v_134;
assign x_7563 = v_1488 | v_80;
assign x_7564 = v_50 | v_51 | v_49 | v_47 | v_101 | v_100 | v_111 | v_110 | v_131 | ~v_304 | ~v_1486 | ~v_1485 | ~v_416 | ~v_217 | ~v_216 | ~v_415 | ~v_1453 | ~v_1452 | ~v_297 | ~v_1395 | ~v_1394 | ~v_414 | ~v_413 | ~v_1484 | ~v_1483 | ~v_1451 | ~v_1450 | v_1487;
assign x_7565 = v_1486 | v_133;
assign x_7566 = v_1486 | v_61;
assign x_7567 = v_1485 | ~v_133;
assign x_7568 = v_1485 | v_53;
assign x_7569 = v_1484 | v_134;
assign x_7570 = v_1484 | v_63;
assign x_7571 = v_1483 | ~v_134;
assign x_7572 = v_1483 | v_55;
assign x_7573 = v_25 | v_24 | v_23 | v_21 | v_94 | v_93 | v_108 | v_109 | v_128 | ~v_1448 | ~v_293 | ~v_1481 | ~v_1480 | ~v_411 | ~v_410 | ~v_201 | ~v_200 | ~v_1447 | ~v_286 | ~v_1384 | ~v_1383 | ~v_409 | ~v_408 | ~v_1479 | ~v_1478 | ~v_1446 | ~v_1445 | v_1482;
assign x_7574 = v_1481 | v_133;
assign x_7575 = v_1481 | v_36;
assign x_7576 = v_1480 | ~v_133;
assign x_7577 = v_1480 | v_28;
assign x_7578 = v_1479 | v_134;
assign x_7579 = v_1479 | v_38;
assign x_7580 = v_1478 | ~v_134;
assign x_7581 = v_1478 | v_30;
assign x_7582 = v_1477 | ~v_1466;
assign x_7583 = v_1477 | ~v_1471;
assign x_7584 = v_1477 | ~v_1476;
assign x_7585 = v_76 | v_68 | v_73 | v_107 | v_106 | v_105 | v_104 | v_127 | v_113 | ~v_1475 | ~v_1474 | ~v_1442 | ~v_1441 | ~v_184 | ~v_183 | ~v_1473 | ~v_1472 | ~v_182 | ~v_181 | ~v_180 | ~v_179 | ~v_1406 | ~v_1405 | ~v_178 | ~v_177 | ~v_1436 | ~v_1435 | v_1476;
assign x_7586 = v_1475 | v_133;
assign x_7587 = v_1475 | v_87;
assign x_7588 = v_1474 | ~v_133;
assign x_7589 = v_1474 | v_79;
assign x_7590 = v_1473 | v_134;
assign x_7591 = v_1473 | v_90;
assign x_7592 = v_1472 | ~v_134;
assign x_7593 = v_1472 | v_82;
assign x_7594 = v_51 | v_48 | v_43 | v_103 | v_101 | v_100 | v_102 | v_111 | v_126 | ~v_1470 | ~v_1469 | ~v_1433 | ~v_1432 | ~v_165 | ~v_164 | ~v_1468 | ~v_1467 | ~v_163 | ~v_162 | ~v_161 | ~v_160 | ~v_1395 | ~v_1394 | ~v_159 | ~v_158 | ~v_1427 | ~v_1426 | v_1471;
assign x_7595 = v_1470 | v_133;
assign x_7596 = v_1470 | v_62;
assign x_7597 = v_1469 | ~v_133;
assign x_7598 = v_1469 | v_54;
assign x_7599 = v_1468 | v_134;
assign x_7600 = v_1468 | v_65;
assign x_7601 = v_1467 | ~v_134;
assign x_7602 = v_1467 | v_57;
assign x_7603 = v_25 | v_22 | v_17 | v_96 | v_95 | v_94 | v_93 | v_109 | v_122 | ~v_1465 | ~v_1464 | ~v_1423 | ~v_1422 | ~v_146 | ~v_145 | ~v_1463 | ~v_1462 | ~v_144 | ~v_143 | ~v_142 | ~v_141 | ~v_1384 | ~v_1383 | ~v_140 | ~v_139 | ~v_1418 | ~v_1417 | v_1466;
assign x_7604 = v_1465 | v_133;
assign x_7605 = v_1465 | v_37;
assign x_7606 = v_1464 | ~v_133;
assign x_7607 = v_1464 | v_29;
assign x_7608 = v_1463 | v_134;
assign x_7609 = v_1463 | v_40;
assign x_7610 = v_1462 | ~v_134;
assign x_7611 = v_1462 | v_32;
assign x_7612 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1460 | ~v_1444 | v_1461;
assign x_7613 = v_1460 | ~v_1449;
assign x_7614 = v_1460 | ~v_1454;
assign x_7615 = v_1460 | ~v_1459;
assign x_7616 = v_75 | v_74 | v_73 | v_72 | v_105 | v_104 | v_113 | v_112 | ~v_1414 | v_121 | ~v_461 | ~v_1411 | ~v_1458 | ~v_1457 | ~v_311 | ~v_310 | ~v_457 | ~v_456 | ~v_455 | ~v_1408 | ~v_1407 | ~v_1406 | ~v_1405 | ~v_454 | ~v_453 | ~v_1456 | ~v_1455 | v_1459;
assign x_7617 = v_1458 | v_114;
assign x_7618 = v_1458 | v_90;
assign x_7619 = v_1457 | ~v_114;
assign x_7620 = v_1457 | v_82;
assign x_7621 = v_1456 | v_115;
assign x_7622 = v_1456 | v_87;
assign x_7623 = v_1455 | ~v_115;
assign x_7624 = v_1455 | v_79;
assign x_7625 = v_50 | v_49 | v_48 | v_47 | v_101 | v_100 | v_111 | v_110 | v_120 | ~v_450 | ~v_449 | ~v_448 | ~v_447 | ~v_304 | ~v_444 | ~v_1401 | ~v_1400 | ~v_1453 | ~v_1452 | ~v_297 | ~v_443 | ~v_1397 | ~v_1396 | ~v_1395 | ~v_1394 | ~v_1451 | ~v_1450 | v_1454;
assign x_7626 = v_1453 | v_114;
assign x_7627 = v_1453 | v_65;
assign x_7628 = v_1452 | ~v_114;
assign x_7629 = v_1452 | v_57;
assign x_7630 = v_1451 | v_115;
assign x_7631 = v_1451 | v_62;
assign x_7632 = v_1450 | ~v_115;
assign x_7633 = v_1450 | v_54;
assign x_7634 = v_24 | v_23 | v_22 | v_21 | v_94 | v_93 | v_108 | v_109 | v_117 | ~v_1448 | ~v_1392 | ~v_439 | ~v_438 | ~v_437 | ~v_293 | ~v_1389 | ~v_1447 | ~v_286 | ~v_434 | ~v_433 | ~v_1386 | ~v_1385 | ~v_1384 | ~v_1383 | ~v_432 | ~v_1446 | ~v_1445 | v_1449;
assign x_7635 = v_1448 | ~v_114;
assign x_7636 = v_1448 | v_32;
assign x_7637 = v_1447 | v_114;
assign x_7638 = v_1447 | v_40;
assign x_7639 = v_1446 | v_115;
assign x_7640 = v_1446 | v_37;
assign x_7641 = v_1445 | ~v_115;
assign x_7642 = v_1445 | v_29;
assign x_7643 = v_1444 | ~v_1425;
assign x_7644 = v_1444 | ~v_1434;
assign x_7645 = v_1444 | ~v_1443;
assign x_7646 = v_68 | v_75 | v_74 | v_73 | v_106 | v_105 | v_104 | v_113 | v_121 | ~v_1442 | ~v_1441 | ~v_1440 | ~v_1439 | ~v_332 | ~v_331 | ~v_180 | ~v_179 | ~v_1438 | ~v_1406 | ~v_1405 | ~v_230 | ~v_229 | ~v_330 | ~v_329 | ~v_1437 | ~v_1436 | ~v_1435 | v_1443;
assign x_7647 = v_1442 | v_116;
assign x_7648 = v_1442 | v_86;
assign x_7649 = v_1441 | ~v_116;
assign x_7650 = v_1441 | v_78;
assign x_7651 = v_1440 | v_119;
assign x_7652 = v_1440 | v_90;
assign x_7653 = v_1439 | ~v_119;
assign x_7654 = v_1439 | v_82;
assign x_7655 = v_1438 | v_118;
assign x_7656 = v_1438 | v_87;
assign x_7657 = v_1437 | ~v_118;
assign x_7658 = v_1437 | v_79;
assign x_7659 = v_1436 | v_116;
assign x_7660 = v_1436 | v_88;
assign x_7661 = v_1435 | ~v_116;
assign x_7662 = v_1435 | v_80;
assign x_7663 = v_50 | v_49 | v_48 | v_43 | v_101 | v_100 | v_102 | v_111 | v_120 | ~v_225 | ~v_224 | ~v_1433 | ~v_1432 | ~v_1431 | ~v_1430 | ~v_327 | ~v_326 | ~v_161 | ~v_160 | ~v_1395 | ~v_1394 | ~v_325 | ~v_324 | ~v_1429 | ~v_1428 | ~v_1427 | ~v_1426 | v_1434;
assign x_7664 = v_1433 | v_116;
assign x_7665 = v_1433 | v_61;
assign x_7666 = v_1432 | ~v_116;
assign x_7667 = v_1432 | v_53;
assign x_7668 = v_1431 | v_119;
assign x_7669 = v_1431 | v_65;
assign x_7670 = v_1430 | ~v_119;
assign x_7671 = v_1430 | v_57;
assign x_7672 = v_1429 | v_118;
assign x_7673 = v_1429 | v_62;
assign x_7674 = v_1428 | ~v_118;
assign x_7675 = v_1428 | v_54;
assign x_7676 = v_1427 | v_116;
assign x_7677 = v_1427 | v_63;
assign x_7678 = v_1426 | ~v_116;
assign x_7679 = v_1426 | v_55;
assign x_7680 = v_24 | v_23 | v_22 | v_17 | v_95 | v_94 | v_93 | v_109 | v_117 | ~v_1424 | ~v_208 | ~v_1423 | ~v_1422 | ~v_1421 | ~v_322 | ~v_321 | ~v_142 | ~v_141 | ~v_1384 | ~v_1383 | ~v_193 | ~v_320 | ~v_319 | ~v_1420 | ~v_1419 | ~v_1418 | ~v_1417 | v_1425;
assign x_7681 = v_1424 | ~v_119;
assign x_7682 = v_1424 | v_32;
assign x_7683 = v_1423 | v_116;
assign x_7684 = v_1423 | v_36;
assign x_7685 = v_1422 | ~v_116;
assign x_7686 = v_1422 | v_28;
assign x_7687 = v_1421 | v_119;
assign x_7688 = v_1421 | v_40;
assign x_7689 = v_1420 | v_118;
assign x_7690 = v_1420 | v_37;
assign x_7691 = v_1419 | ~v_118;
assign x_7692 = v_1419 | v_29;
assign x_7693 = v_1418 | v_116;
assign x_7694 = v_1418 | v_38;
assign x_7695 = v_1417 | ~v_116;
assign x_7696 = v_1417 | v_30;
assign x_7697 = v_1416 | ~v_1393;
assign x_7698 = v_1416 | ~v_1404;
assign x_7699 = v_1416 | ~v_1415;
assign x_7700 = v_76 | v_74 | v_73 | v_70 | v_107 | v_106 | v_104 | v_113 | v_112 | ~v_1414 | ~v_1413 | ~v_1412 | ~v_1411 | ~v_1410 | ~v_1409 | ~v_1408 | ~v_1407 | ~v_1406 | ~v_1405 | ~v_454 | ~v_453 | ~v_480 | ~v_479 | ~v_478 | ~v_477 | ~v_362 | ~v_361 | v_1415;
assign x_7701 = v_1414 | v_119;
assign x_7702 = v_1414 | v_88;
assign x_7703 = v_1413 | v_116;
assign x_7704 = v_1413 | v_87;
assign x_7705 = v_1412 | ~v_116;
assign x_7706 = v_1412 | v_79;
assign x_7707 = v_1411 | ~v_119;
assign x_7708 = v_1411 | v_80;
assign x_7709 = v_1410 | v_116;
assign x_7710 = v_1410 | v_90;
assign x_7711 = v_1409 | ~v_116;
assign x_7712 = v_1409 | v_82;
assign x_7713 = v_1408 | v_118;
assign x_7714 = v_1408 | v_86;
assign x_7715 = v_1407 | ~v_118;
assign x_7716 = v_1407 | v_78;
assign x_7717 = v_1406 | v_116;
assign x_7718 = v_1406 | v_85;
assign x_7719 = v_1405 | ~v_116;
assign x_7720 = v_1405 | v_77;
assign x_7721 = v_51 | v_49 | v_48 | v_45 | v_103 | v_100 | v_102 | v_111 | v_110 | ~v_449 | ~v_447 | ~v_1403 | ~v_1402 | ~v_1401 | ~v_1400 | ~v_475 | ~v_474 | ~v_1399 | ~v_1398 | ~v_1397 | ~v_1396 | ~v_1395 | ~v_1394 | ~v_473 | ~v_472 | ~v_351 | ~v_350 | v_1404;
assign x_7722 = v_1403 | v_116;
assign x_7723 = v_1403 | v_62;
assign x_7724 = v_1402 | ~v_116;
assign x_7725 = v_1402 | v_54;
assign x_7726 = v_1401 | v_119;
assign x_7727 = v_1401 | v_63;
assign x_7728 = v_1400 | ~v_119;
assign x_7729 = v_1400 | v_55;
assign x_7730 = v_1399 | v_116;
assign x_7731 = v_1399 | v_65;
assign x_7732 = v_1398 | ~v_116;
assign x_7733 = v_1398 | v_57;
assign x_7734 = v_1397 | v_118;
assign x_7735 = v_1397 | v_61;
assign x_7736 = v_1396 | ~v_118;
assign x_7737 = v_1396 | v_53;
assign x_7738 = v_1395 | v_116;
assign x_7739 = v_1395 | v_60;
assign x_7740 = v_1394 | ~v_116;
assign x_7741 = v_1394 | v_52;
assign x_7742 = v_25 | v_23 | v_22 | v_19 | v_96 | v_95 | v_93 | v_108 | v_109 | ~v_470 | ~v_1392 | ~v_437 | ~v_1391 | ~v_1390 | ~v_1389 | ~v_469 | ~v_1388 | ~v_1387 | ~v_1386 | ~v_1385 | ~v_1384 | ~v_1383 | ~v_432 | ~v_468 | ~v_467 | ~v_340 | ~v_339 | v_1393;
assign x_7743 = v_1392 | v_119;
assign x_7744 = v_1392 | v_38;
assign x_7745 = v_1391 | v_116;
assign x_7746 = v_1391 | v_37;
assign x_7747 = v_1390 | ~v_116;
assign x_7748 = v_1390 | v_29;
assign x_7749 = v_1389 | ~v_119;
assign x_7750 = v_1389 | v_30;
assign x_7751 = v_1388 | v_116;
assign x_7752 = v_1388 | v_40;
assign x_7753 = v_1387 | ~v_116;
assign x_7754 = v_1387 | v_32;
assign x_7755 = v_1386 | v_118;
assign x_7756 = v_1386 | v_36;
assign x_7757 = v_1385 | ~v_118;
assign x_7758 = v_1385 | v_28;
assign x_7759 = v_1384 | v_116;
assign x_7760 = v_1384 | v_35;
assign x_7761 = v_1383 | ~v_116;
assign x_7762 = v_1383 | v_27;
assign x_7763 = v_1382 | ~v_1042;
assign x_7764 = v_1382 | ~v_1067;
assign x_7765 = v_1382 | ~v_1116;
assign x_7766 = v_1382 | ~v_1127;
assign x_7767 = v_1382 | ~v_1186;
assign x_7768 = v_1382 | ~v_1229;
assign x_7769 = v_1382 | ~v_1238;
assign x_7770 = v_1382 | ~v_1247;
assign x_7771 = v_1382 | ~v_1256;
assign x_7772 = v_1382 | ~v_1265;
assign x_7773 = v_1382 | ~v_1274;
assign x_7774 = v_1382 | ~v_1283;
assign x_7775 = v_1382 | ~v_1292;
assign x_7776 = v_1382 | ~v_1333;
assign x_7777 = v_1382 | ~v_1342;
assign x_7778 = v_1382 | ~v_1381;
assign x_7779 = v_9 | v_7 | v_5 | v_4 | v_6 | v_3 | v_2 | v_1 | ~v_1041 | ~v_1040 | ~v_1380 | v_1381;
assign x_7780 = v_1380 | ~v_1361;
assign x_7781 = v_1380 | ~v_1379;
assign x_7782 = v_125 | ~v_1037 | ~v_1022 | ~v_1006 | ~v_1183 | ~v_1226 | ~v_1330 | ~v_1378 | v_1379;
assign x_7783 = v_1378 | ~v_1377;
assign x_7784 = v_1378 | ~v_698;
assign x_7785 = v_1378 | ~v_699;
assign x_7786 = v_1378 | ~v_700;
assign x_7787 = v_1378 | ~v_701;
assign x_7788 = ~v_1376 | ~v_1371 | ~v_1366 | v_1377;
assign x_7789 = v_1376 | ~v_759;
assign x_7790 = v_1376 | ~v_760;
assign x_7791 = v_1376 | ~v_1372;
assign x_7792 = v_1376 | ~v_763;
assign x_7793 = v_1376 | ~v_764;
assign x_7794 = v_1376 | ~v_726;
assign x_7795 = v_1376 | ~v_1373;
assign x_7796 = v_1376 | ~v_729;
assign x_7797 = v_1376 | ~v_730;
assign x_7798 = v_1376 | ~v_731;
assign x_7799 = v_1376 | ~v_732;
assign x_7800 = v_1376 | ~v_733;
assign x_7801 = v_1376 | ~v_767;
assign x_7802 = v_1376 | ~v_768;
assign x_7803 = v_1376 | ~v_642;
assign x_7804 = v_1376 | ~v_643;
assign x_7805 = v_1376 | ~v_1374;
assign x_7806 = v_1376 | ~v_1375;
assign x_7807 = v_1376 | ~v_112;
assign x_7808 = v_1376 | ~v_105;
assign x_7809 = v_1376 | ~v_76;
assign x_7810 = v_1376 | ~v_75;
assign x_7811 = v_1376 | ~v_74;
assign x_7812 = v_1376 | ~v_73;
assign x_7813 = v_1376 | ~v_72;
assign x_7814 = v_1376 | ~v_71;
assign x_7815 = v_1376 | ~v_69;
assign x_7816 = ~v_26 | ~v_91 | v_1375;
assign x_7817 = ~v_16 | ~v_26 | v_1374;
assign x_7818 = ~v_13 | v_26 | v_1373;
assign x_7819 = v_26 | ~v_83 | v_1372;
assign x_7820 = v_1371 | ~v_748;
assign x_7821 = v_1371 | ~v_749;
assign x_7822 = v_1371 | ~v_1367;
assign x_7823 = v_1371 | ~v_1368;
assign x_7824 = v_1371 | ~v_750;
assign x_7825 = v_1371 | ~v_714;
assign x_7826 = v_1371 | ~v_716;
assign x_7827 = v_1371 | ~v_717;
assign x_7828 = v_1371 | ~v_719;
assign x_7829 = v_1371 | ~v_720;
assign x_7830 = v_1371 | ~v_755;
assign x_7831 = v_1371 | ~v_756;
assign x_7832 = v_1371 | ~v_623;
assign x_7833 = v_1371 | ~v_624;
assign x_7834 = v_1371 | ~v_757;
assign x_7835 = v_1371 | ~v_1369;
assign x_7836 = v_1371 | ~v_721;
assign x_7837 = v_1371 | ~v_110;
assign x_7838 = v_1371 | ~v_101;
assign x_7839 = v_1371 | ~v_1370;
assign x_7840 = v_1371 | ~v_51;
assign x_7841 = v_1371 | ~v_50;
assign x_7842 = v_1371 | ~v_49;
assign x_7843 = v_1371 | ~v_48;
assign x_7844 = v_1371 | ~v_47;
assign x_7845 = v_1371 | ~v_46;
assign x_7846 = v_1371 | ~v_44;
assign x_7847 = ~v_26 | ~v_66 | v_1370;
assign x_7848 = ~v_14 | ~v_26 | v_1369;
assign x_7849 = v_26 | ~v_58 | v_1368;
assign x_7850 = ~v_12 | v_26 | v_1367;
assign x_7851 = v_1366 | ~v_737;
assign x_7852 = v_1366 | ~v_738;
assign x_7853 = v_1366 | ~v_1362;
assign x_7854 = v_1366 | ~v_739;
assign x_7855 = v_1366 | ~v_705;
assign x_7856 = v_1366 | ~v_706;
assign x_7857 = v_1366 | ~v_707;
assign x_7858 = v_1366 | ~v_708;
assign x_7859 = v_1366 | ~v_1363;
assign x_7860 = v_1366 | ~v_709;
assign x_7861 = v_1366 | ~v_710;
assign x_7862 = v_1366 | ~v_744;
assign x_7863 = v_1366 | ~v_745;
assign x_7864 = v_1366 | ~v_604;
assign x_7865 = v_1366 | ~v_605;
assign x_7866 = v_1366 | ~v_746;
assign x_7867 = v_1366 | ~v_1364;
assign x_7868 = v_1366 | ~v_1365;
assign x_7869 = v_1366 | ~v_108;
assign x_7870 = v_1366 | ~v_94;
assign x_7871 = v_1366 | ~v_25;
assign x_7872 = v_1366 | ~v_24;
assign x_7873 = v_1366 | ~v_23;
assign x_7874 = v_1366 | ~v_22;
assign x_7875 = v_1366 | ~v_21;
assign x_7876 = v_1366 | ~v_20;
assign x_7877 = v_1366 | ~v_18;
assign x_7878 = ~v_15 | ~v_26 | v_1365;
assign x_7879 = ~v_11 | v_26 | v_1364;
assign x_7880 = ~v_26 | ~v_41 | v_1363;
assign x_7881 = ~v_33 | v_26 | v_1362;
assign x_7882 = ~v_586 | ~v_1360 | v_1361;
assign x_7883 = v_1360 | ~v_1359;
assign x_7884 = v_1360 | ~v_1310;
assign x_7885 = v_1360 | ~v_1205;
assign x_7886 = v_1360 | ~v_1154;
assign x_7887 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1358 | v_1359;
assign x_7888 = v_1358 | ~v_1347;
assign x_7889 = v_1358 | ~v_1352;
assign x_7890 = v_1358 | ~v_1357;
assign x_7891 = v_76 | v_69 | v_75 | v_74 | v_73 | v_72 | v_71 | v_105 | ~v_1356 | v_112 | ~v_1355 | ~v_190 | ~v_189 | ~v_315 | ~v_314 | ~v_280 | ~v_279 | ~v_278 | ~v_277 | ~v_276 | ~v_1354 | ~v_273 | ~v_311 | ~v_310 | ~v_1353 | ~v_307 | ~v_306 | v_1357;
assign x_7892 = v_1356 | v_91;
assign x_7893 = v_1356 | v_26;
assign x_7894 = v_1355 | v_26;
assign x_7895 = v_1355 | v_16;
assign x_7896 = v_1354 | v_13;
assign x_7897 = v_1354 | ~v_26;
assign x_7898 = v_1353 | v_83;
assign x_7899 = v_1353 | ~v_26;
assign x_7900 = v_50 | v_51 | v_49 | v_48 | v_46 | v_47 | v_44 | ~v_1351 | v_101 | v_110 | ~v_268 | ~v_1350 | ~v_304 | ~v_171 | ~v_170 | ~v_303 | ~v_302 | ~v_267 | ~v_266 | ~v_264 | ~v_263 | ~v_261 | ~v_297 | ~v_1349 | ~v_1348 | ~v_296 | ~v_295 | v_1352;
assign x_7901 = v_1351 | v_66;
assign x_7902 = v_1351 | v_26;
assign x_7903 = v_1350 | v_26;
assign x_7904 = v_1350 | v_14;
assign x_7905 = v_1349 | v_58;
assign x_7906 = v_1349 | ~v_26;
assign x_7907 = v_1348 | v_12;
assign x_7908 = v_1348 | ~v_26;
assign x_7909 = v_25 | v_24 | v_23 | v_22 | v_21 | v_20 | v_18 | v_94 | v_108 | ~v_1346 | ~v_1345 | ~v_293 | ~v_152 | ~v_151 | ~v_292 | ~v_291 | ~v_257 | ~v_256 | ~v_1344 | ~v_255 | ~v_254 | ~v_253 | ~v_252 | ~v_286 | ~v_1343 | ~v_285 | ~v_284 | v_1347;
assign x_7910 = v_1346 | v_26;
assign x_7911 = v_1346 | v_15;
assign x_7912 = v_1345 | v_11;
assign x_7913 = v_1345 | ~v_26;
assign x_7914 = v_1344 | v_41;
assign x_7915 = v_1344 | v_26;
assign x_7916 = v_1343 | v_33;
assign x_7917 = v_1343 | ~v_26;
assign x_7918 = v_7 | v_5 | v_6 | v_8 | v_10 | v_2 | v_1 | ~v_1041 | ~v_1040 | ~v_1341 | v_1342;
assign x_7919 = v_1341 | ~v_1337;
assign x_7920 = v_1341 | ~v_1340;
assign x_7921 = v_125 | ~v_1037 | ~v_1022 | ~v_1006 | ~v_1106 | ~v_1105 | ~v_1104 | ~v_1180 | ~v_1179 | ~v_1339 | ~v_1338 | v_1340;
assign x_7922 = v_1339 | ~v_1095;
assign x_7923 = v_1339 | ~v_1177;
assign x_7924 = v_1338 | ~v_961;
assign x_7925 = v_1338 | ~v_1110;
assign x_7926 = ~v_586 | ~v_1336 | v_1337;
assign x_7927 = v_1336 | ~v_1334;
assign x_7928 = v_1336 | ~v_1335;
assign x_7929 = v_1336 | ~v_1150;
assign x_7930 = v_1336 | ~v_1151;
assign x_7931 = v_1336 | ~v_1080;
assign x_7932 = v_1336 | ~v_1081;
assign x_7933 = v_1336 | ~v_1082;
assign x_7934 = ~v_1148 | ~v_1071 | v_1335;
assign x_7935 = ~v_1086 | ~v_508 | v_1334;
assign x_7936 = v_9 | v_7 | v_5 | v_4 | v_8 | v_10 | v_2 | v_1 | ~v_1041 | ~v_1040 | ~v_1332 | v_1333;
assign x_7937 = v_1332 | ~v_1312;
assign x_7938 = v_1332 | ~v_1331;
assign x_7939 = v_125 | ~v_1037 | ~v_1022 | ~v_1006 | ~v_1330 | ~v_1182 | ~v_1225 | ~v_1329 | v_1331;
assign x_7940 = v_1330 | ~v_1058;
assign x_7941 = v_1330 | ~v_961;
assign x_7942 = v_1329 | ~v_1328;
assign x_7943 = v_1329 | ~v_698;
assign x_7944 = v_1329 | ~v_699;
assign x_7945 = v_1329 | ~v_700;
assign x_7946 = v_1329 | ~v_701;
assign x_7947 = ~v_1327 | ~v_1322 | ~v_1317 | v_1328;
assign x_7948 = v_1327 | ~v_905;
assign x_7949 = v_1327 | ~v_682;
assign x_7950 = v_1327 | ~v_683;
assign x_7951 = v_1327 | ~v_906;
assign x_7952 = v_1327 | ~v_907;
assign x_7953 = v_1327 | ~v_1323;
assign x_7954 = v_1327 | ~v_1324;
assign x_7955 = v_1327 | ~v_1325;
assign x_7956 = v_1327 | ~v_684;
assign x_7957 = v_1327 | ~v_685;
assign x_7958 = v_1327 | ~v_911;
assign x_7959 = v_1327 | ~v_912;
assign x_7960 = v_1327 | ~v_692;
assign x_7961 = v_1327 | ~v_693;
assign x_7962 = v_1327 | ~v_642;
assign x_7963 = v_1327 | ~v_643;
assign x_7964 = v_1327 | ~v_913;
assign x_7965 = v_1327 | ~v_1326;
assign x_7966 = v_1327 | ~v_113;
assign x_7967 = v_1327 | ~v_112;
assign x_7968 = v_1327 | ~v_106;
assign x_7969 = v_1327 | ~v_105;
assign x_7970 = v_1327 | ~v_76;
assign x_7971 = v_1327 | ~v_75;
assign x_7972 = v_1327 | ~v_74;
assign x_7973 = v_1327 | ~v_73;
assign x_7974 = v_1327 | ~v_69;
assign x_7975 = ~v_13 | v_99 | v_1326;
assign x_7976 = ~v_91 | ~v_99 | v_1325;
assign x_7977 = ~v_83 | v_99 | v_1324;
assign x_7978 = ~v_16 | ~v_99 | v_1323;
assign x_7979 = v_1322 | ~v_894;
assign x_7980 = v_1322 | ~v_895;
assign x_7981 = v_1322 | ~v_1318;
assign x_7982 = v_1322 | ~v_663;
assign x_7983 = v_1322 | ~v_664;
assign x_7984 = v_1322 | ~v_1319;
assign x_7985 = v_1322 | ~v_898;
assign x_7986 = v_1322 | ~v_899;
assign x_7987 = v_1322 | ~v_673;
assign x_7988 = v_1322 | ~v_674;
assign x_7989 = v_1322 | ~v_623;
assign x_7990 = v_1322 | ~v_624;
assign x_7991 = v_1322 | ~v_900;
assign x_7992 = v_1322 | ~v_677;
assign x_7993 = v_1322 | ~v_902;
assign x_7994 = v_1322 | ~v_1320;
assign x_7995 = v_1322 | ~v_678;
assign x_7996 = v_1322 | ~v_1321;
assign x_7997 = v_1322 | ~v_111;
assign x_7998 = v_1322 | ~v_110;
assign x_7999 = v_1322 | ~v_102;
assign x_8000 = v_1322 | ~v_101;
assign x_8001 = v_1322 | ~v_51;
assign x_8002 = v_1322 | ~v_50;
assign x_8003 = v_1322 | ~v_49;
assign x_8004 = v_1322 | ~v_48;
assign x_8005 = v_1322 | ~v_44;
assign x_8006 = ~v_12 | v_99 | v_1321;
assign x_8007 = ~v_58 | v_99 | v_1320;
assign x_8008 = ~v_14 | ~v_99 | v_1319;
assign x_8009 = ~v_66 | ~v_99 | v_1318;
assign x_8010 = v_1317 | ~v_883;
assign x_8011 = v_1317 | ~v_884;
assign x_8012 = v_1317 | ~v_646;
assign x_8013 = v_1317 | ~v_885;
assign x_8014 = v_1317 | ~v_1313;
assign x_8015 = v_1317 | ~v_1314;
assign x_8016 = v_1317 | ~v_647;
assign x_8017 = v_1317 | ~v_648;
assign x_8018 = v_1317 | ~v_888;
assign x_8019 = v_1317 | ~v_889;
assign x_8020 = v_1317 | ~v_657;
assign x_8021 = v_1317 | ~v_658;
assign x_8022 = v_1317 | ~v_604;
assign x_8023 = v_1317 | ~v_605;
assign x_8024 = v_1317 | ~v_1315;
assign x_8025 = v_1317 | ~v_661;
assign x_8026 = v_1317 | ~v_890;
assign x_8027 = v_1317 | ~v_1316;
assign x_8028 = v_1317 | ~v_109;
assign x_8029 = v_1317 | ~v_108;
assign x_8030 = v_1317 | ~v_95;
assign x_8031 = v_1317 | ~v_94;
assign x_8032 = v_1317 | ~v_25;
assign x_8033 = v_1317 | ~v_24;
assign x_8034 = v_1317 | ~v_23;
assign x_8035 = v_1317 | ~v_22;
assign x_8036 = v_1317 | ~v_18;
assign x_8037 = ~v_41 | ~v_99 | v_1316;
assign x_8038 = ~v_33 | v_99 | v_1315;
assign x_8039 = ~v_15 | ~v_99 | v_1314;
assign x_8040 = ~v_11 | v_99 | v_1313;
assign x_8041 = ~v_586 | ~v_1311 | v_1312;
assign x_8042 = v_1311 | ~v_1309;
assign x_8043 = v_1311 | ~v_1204;
assign x_8044 = v_1311 | ~v_1153;
assign x_8045 = v_1311 | ~v_1310;
assign x_8046 = ~v_508 | ~v_1046 | v_1310;
assign x_8047 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1308 | v_1309;
assign x_8048 = v_1308 | ~v_1297;
assign x_8049 = v_1308 | ~v_1302;
assign x_8050 = v_1308 | ~v_1307;
assign x_8051 = v_76 | v_69 | v_75 | v_74 | v_73 | v_106 | v_105 | v_113 | v_112 | ~v_1306 | ~v_460 | ~v_190 | ~v_189 | ~v_240 | ~v_239 | ~v_459 | ~v_458 | ~v_232 | ~v_231 | ~v_1305 | ~v_1304 | ~v_1303 | ~v_454 | ~v_453 | ~v_230 | ~v_229 | ~v_452 | v_1307;
assign x_8052 = v_1306 | ~v_99;
assign x_8053 = v_1306 | v_13;
assign x_8054 = v_1305 | v_99;
assign x_8055 = v_1305 | v_91;
assign x_8056 = v_1304 | ~v_99;
assign x_8057 = v_1304 | v_83;
assign x_8058 = v_1303 | v_99;
assign x_8059 = v_1303 | v_16;
assign x_8060 = v_50 | v_51 | v_49 | v_48 | v_44 | v_101 | v_102 | v_111 | v_110 | ~v_1301 | ~v_225 | ~v_1300 | ~v_449 | ~v_224 | ~v_447 | ~v_171 | ~v_170 | ~v_221 | ~v_220 | ~v_446 | ~v_445 | ~v_1299 | ~v_211 | ~v_210 | ~v_1298 | ~v_442 | ~v_441 | v_1302;
assign x_8061 = v_1301 | ~v_99;
assign x_8062 = v_1301 | v_12;
assign x_8063 = v_1300 | ~v_99;
assign x_8064 = v_1300 | v_58;
assign x_8065 = v_1299 | v_99;
assign x_8066 = v_1299 | v_14;
assign x_8067 = v_1298 | v_99;
assign x_8068 = v_1298 | v_66;
assign x_8069 = v_25 | v_24 | v_23 | v_22 | v_18 | v_95 | v_94 | v_108 | v_109 | ~v_1296 | ~v_437 | ~v_208 | ~v_1295 | ~v_152 | ~v_151 | ~v_205 | ~v_204 | ~v_436 | ~v_435 | ~v_195 | ~v_194 | ~v_1294 | ~v_1293 | ~v_432 | ~v_193 | ~v_431 | ~v_430 | v_1297;
assign x_8070 = v_1296 | v_99;
assign x_8071 = v_1296 | v_41;
assign x_8072 = v_1295 | ~v_99;
assign x_8073 = v_1295 | v_33;
assign x_8074 = v_1294 | v_99;
assign x_8075 = v_1294 | v_15;
assign x_8076 = v_1293 | ~v_99;
assign x_8077 = v_1293 | v_11;
assign x_8078 = v_9 | v_7 | v_5 | v_4 | v_6 | v_8 | v_2 | v_1 | ~v_1041 | ~v_1040 | ~v_1291 | v_1292;
assign x_8079 = v_1291 | ~v_1287;
assign x_8080 = v_1291 | ~v_1290;
assign x_8081 = v_125 | ~v_1037 | ~v_1022 | ~v_1006 | ~v_960 | ~v_959 | ~v_958 | ~v_957 | ~v_936 | ~v_1289 | ~v_1288 | v_1290;
assign x_8082 = v_1289 | ~v_1181;
assign x_8083 = v_1289 | ~v_1059;
assign x_8084 = v_1288 | ~v_1095;
assign x_8085 = v_1288 | ~v_980;
assign x_8086 = ~v_586 | ~v_1286 | v_1287;
assign x_8087 = v_1286 | ~v_1284;
assign x_8088 = v_1286 | ~v_1285;
assign x_8089 = v_1286 | ~v_483;
assign x_8090 = v_1286 | ~v_504;
assign x_8091 = v_1286 | ~v_505;
assign x_8092 = v_1286 | ~v_506;
assign x_8093 = v_1286 | ~v_507;
assign x_8094 = ~v_1047 | ~v_1152 | v_1285;
assign x_8095 = ~v_527 | ~v_1071 | v_1284;
assign x_8096 = v_9 | v_7 | v_4 | v_6 | v_8 | v_10 | v_2 | v_1 | ~v_1041 | ~v_1040 | ~v_1282 | v_1283;
assign x_8097 = v_1282 | ~v_1278;
assign x_8098 = v_1282 | ~v_1281;
assign x_8099 = v_125 | ~v_1037 | ~v_1022 | ~v_1006 | ~v_970 | ~v_969 | ~v_968 | ~v_1094 | ~v_1093 | ~v_1280 | ~v_1279 | v_1281;
assign x_8100 = v_1280 | ~v_976;
assign x_8101 = v_1280 | ~v_1181;
assign x_8102 = v_1279 | ~v_961;
assign x_8103 = v_1279 | ~v_1122;
assign x_8104 = ~v_586 | ~v_1277 | v_1278;
assign x_8105 = v_1277 | ~v_1275;
assign x_8106 = v_1277 | ~v_1276;
assign x_8107 = v_1277 | ~v_1069;
assign x_8108 = v_1277 | ~v_1070;
assign x_8109 = v_1277 | ~v_515;
assign x_8110 = v_1277 | ~v_516;
assign x_8111 = v_1277 | ~v_517;
assign x_8112 = ~v_1152 | ~v_523 | v_1276;
assign x_8113 = ~v_1117 | ~v_508 | v_1275;
assign x_8114 = v_9 | v_7 | v_5 | v_4 | v_10 | v_3 | v_2 | v_1 | ~v_1041 | ~v_1040 | ~v_1273 | v_1274;
assign x_8115 = v_1273 | ~v_1269;
assign x_8116 = v_1273 | ~v_1272;
assign x_8117 = v_125 | ~v_1037 | ~v_1022 | ~v_1006 | ~v_859 | ~v_858 | ~v_841 | ~v_1057 | ~v_1055 | ~v_1271 | ~v_1270 | v_1272;
assign x_8118 = v_1271 | ~v_881;
assign x_8119 = v_1271 | ~v_1110;
assign x_8120 = v_1270 | ~v_1063;
assign x_8121 = v_1270 | ~v_1122;
assign x_8122 = ~v_586 | ~v_1268 | v_1269;
assign x_8123 = v_1268 | ~v_1266;
assign x_8124 = v_1268 | ~v_1267;
assign x_8125 = v_1268 | ~v_1043;
assign x_8126 = v_1268 | ~v_1045;
assign x_8127 = v_1268 | ~v_388;
assign x_8128 = v_1268 | ~v_405;
assign x_8129 = v_1268 | ~v_406;
assign x_8130 = ~v_1086 | ~v_428 | v_1267;
assign x_8131 = ~v_1117 | ~v_1051 | v_1266;
assign x_8132 = v_7 | v_5 | v_6 | v_10 | v_3 | v_2 | v_1 | ~v_1041 | ~v_1040 | ~v_1264 | v_1265;
assign x_8133 = v_1264 | ~v_1260;
assign x_8134 = v_1264 | ~v_1263;
assign x_8135 = v_125 | ~v_1037 | ~v_1022 | ~v_1006 | ~v_1109 | ~v_1108 | ~v_1103 | ~v_1102 | ~v_1101 | ~v_1262 | ~v_1261 | v_1263;
assign x_8136 = v_1262 | ~v_1177;
assign x_8137 = v_1262 | ~v_1122;
assign x_8138 = v_1261 | ~v_1181;
assign x_8139 = v_1261 | ~v_1058;
assign x_8140 = ~v_586 | ~v_1259 | v_1260;
assign x_8141 = v_1259 | ~v_1257;
assign x_8142 = v_1259 | ~v_1258;
assign x_8143 = v_1259 | ~v_1077;
assign x_8144 = v_1259 | ~v_1078;
assign x_8145 = v_1259 | ~v_1079;
assign x_8146 = v_1259 | ~v_1084;
assign x_8147 = v_1259 | ~v_1085;
assign x_8148 = ~v_1117 | ~v_1148 | v_1258;
assign x_8149 = ~v_1046 | ~v_1152 | v_1257;
assign x_8150 = v_7 | v_5 | v_6 | v_8 | v_10 | v_3 | v_1 | ~v_1041 | ~v_1040 | ~v_1255 | v_1256;
assign x_8151 = v_1255 | ~v_1251;
assign x_8152 = v_1255 | ~v_1254;
assign x_8153 = v_125 | ~v_1037 | ~v_1022 | ~v_1006 | ~v_1099 | ~v_1098 | ~v_1097 | ~v_1176 | ~v_1175 | ~v_1253 | ~v_1252 | v_1254;
assign x_8154 = v_1253 | ~v_1063;
assign x_8155 = v_1253 | ~v_1181;
assign x_8156 = v_1252 | ~v_980;
assign x_8157 = v_1252 | ~v_1110;
assign x_8158 = ~v_586 | ~v_1250 | v_1251;
assign x_8159 = v_1250 | ~v_1248;
assign x_8160 = v_1250 | ~v_1249;
assign x_8161 = v_1250 | ~v_1146;
assign x_8162 = v_1250 | ~v_1147;
assign x_8163 = v_1250 | ~v_1073;
assign x_8164 = v_1250 | ~v_1074;
assign x_8165 = v_1250 | ~v_1075;
assign x_8166 = ~v_1152 | ~v_1051 | v_1249;
assign x_8167 = ~v_1086 | ~v_527 | v_1248;
assign x_8168 = v_9 | v_7 | v_5 | v_4 | v_8 | v_10 | v_3 | v_1 | ~v_1041 | ~v_1040 | ~v_1246 | v_1247;
assign x_8169 = v_1246 | ~v_1242;
assign x_8170 = v_1246 | ~v_1245;
assign x_8171 = v_125 | ~v_1037 | ~v_1022 | ~v_1006 | ~v_788 | ~v_771 | ~v_702 | ~v_1062 | ~v_1061 | ~v_1244 | ~v_1243 | v_1245;
assign x_8172 = v_1244 | ~v_881;
assign x_8173 = v_1244 | ~v_1177;
assign x_8174 = v_1243 | ~v_1058;
assign x_8175 = v_1243 | ~v_980;
assign x_8176 = ~v_586 | ~v_1241 | v_1242;
assign x_8177 = v_1241 | ~v_1239;
assign x_8178 = v_1241 | ~v_1240;
assign x_8179 = v_1241 | ~v_1049;
assign x_8180 = v_1241 | ~v_1050;
assign x_8181 = v_1241 | ~v_249;
assign x_8182 = v_1241 | ~v_318;
assign x_8183 = v_1241 | ~v_335;
assign x_8184 = ~v_1148 | ~v_428 | v_1240;
assign x_8185 = ~v_527 | ~v_1046 | v_1239;
assign x_8186 = v_9 | v_7 | v_5 | v_4 | v_6 | v_8 | v_3 | v_1 | ~v_1041 | ~v_1040 | ~v_1237 | v_1238;
assign x_8187 = v_1237 | ~v_1233;
assign x_8188 = v_1237 | ~v_1236;
assign x_8189 = v_125 | ~v_1037 | ~v_1022 | ~v_1006 | ~v_918 | ~v_917 | ~v_882 | ~v_979 | ~v_977 | ~v_1235 | ~v_1234 | v_1236;
assign x_8190 = v_1235 | ~v_1177;
assign x_8191 = v_1235 | ~v_1059;
assign x_8192 = v_1234 | ~v_1063;
assign x_8193 = v_1234 | ~v_961;
assign x_8194 = ~v_586 | ~v_1232 | v_1233;
assign x_8195 = v_1232 | ~v_1230;
assign x_8196 = v_1232 | ~v_1231;
assign x_8197 = v_1232 | ~v_524;
assign x_8198 = v_1232 | ~v_526;
assign x_8199 = v_1232 | ~v_429;
assign x_8200 = v_1232 | ~v_464;
assign x_8201 = v_1232 | ~v_465;
assign x_8202 = ~v_1047 | ~v_1148 | v_1231;
assign x_8203 = ~v_508 | ~v_1051 | v_1230;
assign x_8204 = v_9 | v_7 | v_4 | v_6 | v_8 | v_10 | v_3 | v_1 | ~v_1041 | ~v_1040 | ~v_1228 | v_1229;
assign x_8205 = v_1228 | ~v_1207;
assign x_8206 = v_1228 | ~v_1227;
assign x_8207 = v_125 | ~v_1037 | ~v_1022 | ~v_1006 | ~v_1226 | ~v_1225 | ~v_1178 | ~v_1224 | v_1227;
assign x_8208 = v_1226 | ~v_1122;
assign x_8209 = v_1226 | ~v_980;
assign x_8210 = v_1225 | ~v_1063;
assign x_8211 = v_1225 | ~v_1095;
assign x_8212 = v_1224 | ~v_1223;
assign x_8213 = v_1224 | ~v_698;
assign x_8214 = v_1224 | ~v_699;
assign x_8215 = v_1224 | ~v_700;
assign x_8216 = v_1224 | ~v_701;
assign x_8217 = ~v_1222 | ~v_1217 | ~v_1212 | v_1223;
assign x_8218 = v_1222 | ~v_628;
assign x_8219 = v_1222 | ~v_629;
assign x_8220 = v_1222 | ~v_1218;
assign x_8221 = v_1222 | ~v_1219;
assign x_8222 = v_1222 | ~v_814;
assign x_8223 = v_1222 | ~v_815;
assign x_8224 = v_1222 | ~v_632;
assign x_8225 = v_1222 | ~v_633;
assign x_8226 = v_1222 | ~v_1220;
assign x_8227 = v_1222 | ~v_1221;
assign x_8228 = v_1222 | ~v_818;
assign x_8229 = v_1222 | ~v_819;
assign x_8230 = v_1222 | ~v_640;
assign x_8231 = v_1222 | ~v_641;
assign x_8232 = v_1222 | ~v_820;
assign x_8233 = v_1222 | ~v_642;
assign x_8234 = v_1222 | ~v_643;
assign x_8235 = v_1222 | ~v_821;
assign x_8236 = v_1222 | ~v_113;
assign x_8237 = v_1222 | ~v_112;
assign x_8238 = v_1222 | ~v_106;
assign x_8239 = v_1222 | ~v_105;
assign x_8240 = v_1222 | ~v_76;
assign x_8241 = v_1222 | ~v_75;
assign x_8242 = v_1222 | ~v_74;
assign x_8243 = v_1222 | ~v_73;
assign x_8244 = v_1222 | ~v_69;
assign x_8245 = ~v_91 | ~v_116 | v_1221;
assign x_8246 = ~v_83 | v_116 | v_1220;
assign x_8247 = ~v_16 | ~v_116 | v_1219;
assign x_8248 = ~v_13 | v_116 | v_1218;
assign x_8249 = v_1217 | ~v_609;
assign x_8250 = v_1217 | ~v_610;
assign x_8251 = v_1217 | ~v_1213;
assign x_8252 = v_1217 | ~v_1214;
assign x_8253 = v_1217 | ~v_803;
assign x_8254 = v_1217 | ~v_804;
assign x_8255 = v_1217 | ~v_613;
assign x_8256 = v_1217 | ~v_614;
assign x_8257 = v_1217 | ~v_1215;
assign x_8258 = v_1217 | ~v_1216;
assign x_8259 = v_1217 | ~v_807;
assign x_8260 = v_1217 | ~v_808;
assign x_8261 = v_1217 | ~v_621;
assign x_8262 = v_1217 | ~v_622;
assign x_8263 = v_1217 | ~v_809;
assign x_8264 = v_1217 | ~v_810;
assign x_8265 = v_1217 | ~v_623;
assign x_8266 = v_1217 | ~v_624;
assign x_8267 = v_1217 | ~v_111;
assign x_8268 = v_1217 | ~v_110;
assign x_8269 = v_1217 | ~v_102;
assign x_8270 = v_1217 | ~v_101;
assign x_8271 = v_1217 | ~v_51;
assign x_8272 = v_1217 | ~v_50;
assign x_8273 = v_1217 | ~v_49;
assign x_8274 = v_1217 | ~v_48;
assign x_8275 = v_1217 | ~v_44;
assign x_8276 = ~v_66 | ~v_116 | v_1216;
assign x_8277 = ~v_58 | v_116 | v_1215;
assign x_8278 = ~v_14 | ~v_116 | v_1214;
assign x_8279 = ~v_12 | v_116 | v_1213;
assign x_8280 = v_1212 | ~v_590;
assign x_8281 = v_1212 | ~v_591;
assign x_8282 = v_1212 | ~v_1208;
assign x_8283 = v_1212 | ~v_1209;
assign x_8284 = v_1212 | ~v_792;
assign x_8285 = v_1212 | ~v_793;
assign x_8286 = v_1212 | ~v_594;
assign x_8287 = v_1212 | ~v_595;
assign x_8288 = v_1212 | ~v_1210;
assign x_8289 = v_1212 | ~v_1211;
assign x_8290 = v_1212 | ~v_796;
assign x_8291 = v_1212 | ~v_797;
assign x_8292 = v_1212 | ~v_602;
assign x_8293 = v_1212 | ~v_603;
assign x_8294 = v_1212 | ~v_798;
assign x_8295 = v_1212 | ~v_799;
assign x_8296 = v_1212 | ~v_604;
assign x_8297 = v_1212 | ~v_605;
assign x_8298 = v_1212 | ~v_109;
assign x_8299 = v_1212 | ~v_108;
assign x_8300 = v_1212 | ~v_95;
assign x_8301 = v_1212 | ~v_94;
assign x_8302 = v_1212 | ~v_25;
assign x_8303 = v_1212 | ~v_24;
assign x_8304 = v_1212 | ~v_23;
assign x_8305 = v_1212 | ~v_22;
assign x_8306 = v_1212 | ~v_18;
assign x_8307 = ~v_41 | ~v_116 | v_1211;
assign x_8308 = ~v_33 | v_116 | v_1210;
assign x_8309 = ~v_15 | ~v_116 | v_1209;
assign x_8310 = ~v_11 | v_116 | v_1208;
assign x_8311 = ~v_586 | ~v_1206 | v_1207;
assign x_8312 = v_1206 | ~v_1203;
assign x_8313 = v_1206 | ~v_1149;
assign x_8314 = v_1206 | ~v_1204;
assign x_8315 = v_1206 | ~v_1205;
assign x_8316 = ~v_527 | ~v_1117 | v_1205;
assign x_8317 = ~v_1071 | ~v_1051 | v_1204;
assign x_8318 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1202 | v_1203;
assign x_8319 = v_1202 | ~v_1191;
assign x_8320 = v_1202 | ~v_1196;
assign x_8321 = v_1202 | ~v_1201;
assign x_8322 = v_76 | v_69 | v_75 | v_74 | v_73 | v_106 | v_105 | v_113 | v_112 | ~v_368 | ~v_190 | ~v_189 | ~v_367 | ~v_188 | ~v_187 | ~v_366 | ~v_365 | ~v_1200 | ~v_1199 | ~v_180 | ~v_179 | ~v_362 | ~v_361 | ~v_1198 | ~v_1197 | ~v_176 | ~v_175 | v_1201;
assign x_8323 = v_1200 | v_116;
assign x_8324 = v_1200 | v_91;
assign x_8325 = v_1199 | ~v_116;
assign x_8326 = v_1199 | v_83;
assign x_8327 = v_1198 | v_116;
assign x_8328 = v_1198 | v_16;
assign x_8329 = v_1197 | ~v_116;
assign x_8330 = v_1197 | v_13;
assign x_8331 = v_50 | v_51 | v_49 | v_48 | v_44 | v_101 | v_102 | v_111 | v_110 | ~v_171 | ~v_170 | ~v_357 | ~v_356 | ~v_169 | ~v_168 | ~v_355 | ~v_354 | ~v_1195 | ~v_1194 | ~v_161 | ~v_160 | ~v_351 | ~v_350 | ~v_1193 | ~v_1192 | ~v_157 | ~v_156 | v_1196;
assign x_8332 = v_1195 | v_116;
assign x_8333 = v_1195 | v_66;
assign x_8334 = v_1194 | ~v_116;
assign x_8335 = v_1194 | v_58;
assign x_8336 = v_1193 | v_116;
assign x_8337 = v_1193 | v_14;
assign x_8338 = v_1192 | ~v_116;
assign x_8339 = v_1192 | v_12;
assign x_8340 = v_25 | v_24 | v_23 | v_22 | v_18 | v_95 | v_94 | v_108 | v_109 | ~v_152 | ~v_151 | ~v_346 | ~v_345 | ~v_150 | ~v_149 | ~v_344 | ~v_343 | ~v_1190 | ~v_1189 | ~v_142 | ~v_141 | ~v_340 | ~v_339 | ~v_1188 | ~v_1187 | ~v_138 | ~v_137 | v_1191;
assign x_8341 = v_1190 | v_116;
assign x_8342 = v_1190 | v_41;
assign x_8343 = v_1189 | ~v_116;
assign x_8344 = v_1189 | v_33;
assign x_8345 = v_1188 | v_116;
assign x_8346 = v_1188 | v_15;
assign x_8347 = v_1187 | ~v_116;
assign x_8348 = v_1187 | v_11;
assign x_8349 = v_5 | v_6 | v_8 | v_10 | v_3 | v_2 | ~v_1041 | ~v_1040 | ~v_1185 | v_1186;
assign x_8350 = v_1185 | ~v_1156;
assign x_8351 = v_1185 | ~v_1184;
assign x_8352 = v_125 | ~v_1037 | ~v_1022 | ~v_1006 | ~v_1183 | ~v_1182 | ~v_1178 | ~v_1173 | v_1184;
assign x_8353 = v_1183 | ~v_1110;
assign x_8354 = v_1183 | ~v_1059;
assign x_8355 = v_1182 | ~v_881;
assign x_8356 = v_1182 | ~v_1181;
assign x_8357 = ~v_1106 | ~v_1105 | ~v_1104 | ~v_1180 | ~v_1179 | v_1181;
assign x_8358 = v_1180 | ~v_1174;
assign x_8359 = v_1180 | ~v_916;
assign x_8360 = v_1180 | ~v_698;
assign x_8361 = v_1180 | ~v_699;
assign x_8362 = v_1180 | ~v_700;
assign x_8363 = v_1180 | ~v_701;
assign x_8364 = v_1179 | ~v_1100;
assign x_8365 = v_1179 | ~v_935;
assign x_8366 = v_1179 | ~v_698;
assign x_8367 = v_1179 | ~v_699;
assign x_8368 = v_1179 | ~v_700;
assign x_8369 = v_1179 | ~v_701;
assign x_8370 = v_1178 | ~v_976;
assign x_8371 = v_1178 | ~v_1177;
assign x_8372 = ~v_1099 | ~v_1098 | ~v_1097 | ~v_1176 | ~v_1175 | v_1177;
assign x_8373 = v_1176 | ~v_1107;
assign x_8374 = v_1176 | ~v_787;
assign x_8375 = v_1176 | ~v_698;
assign x_8376 = v_1176 | ~v_699;
assign x_8377 = v_1176 | ~v_700;
assign x_8378 = v_1176 | ~v_701;
assign x_8379 = v_1175 | ~v_1174;
assign x_8380 = v_1175 | ~v_770;
assign x_8381 = v_1175 | ~v_698;
assign x_8382 = v_1175 | ~v_699;
assign x_8383 = v_1175 | ~v_700;
assign x_8384 = v_1175 | ~v_701;
assign x_8385 = ~v_1109 | ~v_1103 | ~v_1102 | v_1174;
assign x_8386 = v_1173 | ~v_1172;
assign x_8387 = v_1173 | ~v_698;
assign x_8388 = v_1173 | ~v_699;
assign x_8389 = v_1173 | ~v_700;
assign x_8390 = v_1173 | ~v_701;
assign x_8391 = ~v_1171 | ~v_1166 | ~v_1161 | v_1172;
assign x_8392 = v_1171 | ~v_626;
assign x_8393 = v_1171 | ~v_627;
assign x_8394 = v_1171 | ~v_1167;
assign x_8395 = v_1171 | ~v_1168;
assign x_8396 = v_1171 | ~v_634;
assign x_8397 = v_1171 | ~v_635;
assign x_8398 = v_1171 | ~v_1169;
assign x_8399 = v_1171 | ~v_1170;
assign x_8400 = v_1171 | ~v_638;
assign x_8401 = v_1171 | ~v_639;
assign x_8402 = v_1171 | ~v_688;
assign x_8403 = v_1171 | ~v_689;
assign x_8404 = v_1171 | ~v_690;
assign x_8405 = v_1171 | ~v_691;
assign x_8406 = v_1171 | ~v_694;
assign x_8407 = v_1171 | ~v_695;
assign x_8408 = v_1171 | ~v_642;
assign x_8409 = v_1171 | ~v_643;
assign x_8410 = v_1171 | ~v_132;
assign x_8411 = v_1171 | ~v_127;
assign x_8412 = v_1171 | ~v_113;
assign x_8413 = v_1171 | ~v_106;
assign x_8414 = v_1171 | ~v_76;
assign x_8415 = v_1171 | ~v_75;
assign x_8416 = v_1171 | ~v_70;
assign x_8417 = v_1171 | ~v_69;
assign x_8418 = v_1171 | ~v_68;
assign x_8419 = ~v_91 | ~v_125 | v_1170;
assign x_8420 = ~v_83 | v_125 | v_1169;
assign x_8421 = ~v_16 | ~v_125 | v_1168;
assign x_8422 = ~v_13 | v_125 | v_1167;
assign x_8423 = v_1166 | ~v_607;
assign x_8424 = v_1166 | ~v_608;
assign x_8425 = v_1166 | ~v_615;
assign x_8426 = v_1166 | ~v_616;
assign x_8427 = v_1166 | ~v_1162;
assign x_8428 = v_1166 | ~v_1163;
assign x_8429 = v_1166 | ~v_619;
assign x_8430 = v_1166 | ~v_620;
assign x_8431 = v_1166 | ~v_669;
assign x_8432 = v_1166 | ~v_670;
assign x_8433 = v_1166 | ~v_1164;
assign x_8434 = v_1166 | ~v_1165;
assign x_8435 = v_1166 | ~v_671;
assign x_8436 = v_1166 | ~v_672;
assign x_8437 = v_1166 | ~v_675;
assign x_8438 = v_1166 | ~v_676;
assign x_8439 = v_1166 | ~v_623;
assign x_8440 = v_1166 | ~v_624;
assign x_8441 = v_1166 | ~v_131;
assign x_8442 = v_1166 | ~v_126;
assign x_8443 = v_1166 | ~v_111;
assign x_8444 = v_1166 | ~v_102;
assign x_8445 = v_1166 | ~v_51;
assign x_8446 = v_1166 | ~v_50;
assign x_8447 = v_1166 | ~v_45;
assign x_8448 = v_1166 | ~v_44;
assign x_8449 = v_1166 | ~v_43;
assign x_8450 = ~v_12 | v_125 | v_1165;
assign x_8451 = ~v_14 | ~v_125 | v_1164;
assign x_8452 = ~v_66 | ~v_125 | v_1163;
assign x_8453 = ~v_58 | v_125 | v_1162;
assign x_8454 = v_1161 | ~v_588;
assign x_8455 = v_1161 | ~v_589;
assign x_8456 = v_1161 | ~v_596;
assign x_8457 = v_1161 | ~v_597;
assign x_8458 = v_1161 | ~v_1157;
assign x_8459 = v_1161 | ~v_1158;
assign x_8460 = v_1161 | ~v_600;
assign x_8461 = v_1161 | ~v_601;
assign x_8462 = v_1161 | ~v_653;
assign x_8463 = v_1161 | ~v_654;
assign x_8464 = v_1161 | ~v_1159;
assign x_8465 = v_1161 | ~v_1160;
assign x_8466 = v_1161 | ~v_655;
assign x_8467 = v_1161 | ~v_656;
assign x_8468 = v_1161 | ~v_659;
assign x_8469 = v_1161 | ~v_660;
assign x_8470 = v_1161 | ~v_604;
assign x_8471 = v_1161 | ~v_605;
assign x_8472 = v_1161 | ~v_128;
assign x_8473 = v_1161 | ~v_122;
assign x_8474 = v_1161 | ~v_109;
assign x_8475 = v_1161 | ~v_95;
assign x_8476 = v_1161 | ~v_25;
assign x_8477 = v_1161 | ~v_24;
assign x_8478 = v_1161 | ~v_19;
assign x_8479 = v_1161 | ~v_18;
assign x_8480 = v_1161 | ~v_17;
assign x_8481 = ~v_15 | ~v_125 | v_1160;
assign x_8482 = ~v_11 | v_125 | v_1159;
assign x_8483 = ~v_41 | ~v_125 | v_1158;
assign x_8484 = ~v_33 | v_125 | v_1157;
assign x_8485 = ~v_586 | ~v_1155 | v_1156;
assign x_8486 = v_1155 | ~v_1144;
assign x_8487 = v_1155 | ~v_1149;
assign x_8488 = v_1155 | ~v_1153;
assign x_8489 = v_1155 | ~v_1154;
assign x_8490 = ~v_1047 | ~v_1086 | v_1154;
assign x_8491 = ~v_1152 | ~v_428 | v_1153;
assign x_8492 = v_1152 | ~v_1150;
assign x_8493 = v_1152 | ~v_1151;
assign x_8494 = v_1152 | ~v_1080;
assign x_8495 = v_1152 | ~v_1081;
assign x_8496 = v_1152 | ~v_1082;
assign x_8497 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_463 | ~v_1145 | v_1151;
assign x_8498 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_482 | ~v_1076 | v_1150;
assign x_8499 = ~v_1148 | ~v_523 | v_1149;
assign x_8500 = v_1148 | ~v_1146;
assign x_8501 = v_1148 | ~v_1147;
assign x_8502 = v_1148 | ~v_1073;
assign x_8503 = v_1148 | ~v_1074;
assign x_8504 = v_1148 | ~v_1075;
assign x_8505 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_334 | ~v_1083 | v_1147;
assign x_8506 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_317 | ~v_1145 | v_1146;
assign x_8507 = v_1145 | ~v_1078;
assign x_8508 = v_1145 | ~v_1079;
assign x_8509 = v_1145 | ~v_1085;
assign x_8510 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1143 | v_1144;
assign x_8511 = v_1143 | ~v_1132;
assign x_8512 = v_1143 | ~v_1137;
assign x_8513 = v_1143 | ~v_1142;
assign x_8514 = v_76 | v_69 | v_68 | v_75 | v_70 | v_106 | v_132 | v_127 | v_113 | ~v_190 | ~v_189 | ~v_242 | ~v_241 | ~v_238 | ~v_237 | ~v_236 | ~v_235 | ~v_186 | ~v_185 | ~v_1141 | ~v_1140 | ~v_182 | ~v_181 | ~v_1139 | ~v_1138 | ~v_174 | ~v_173 | v_1142;
assign x_8515 = v_1141 | v_125;
assign x_8516 = v_1141 | v_91;
assign x_8517 = v_1140 | ~v_125;
assign x_8518 = v_1140 | v_83;
assign x_8519 = v_1139 | v_125;
assign x_8520 = v_1139 | v_16;
assign x_8521 = v_1138 | ~v_125;
assign x_8522 = v_1138 | v_13;
assign x_8523 = v_50 | v_51 | v_45 | v_43 | v_44 | v_102 | v_111 | v_131 | v_126 | ~v_171 | ~v_170 | ~v_223 | ~v_222 | ~v_219 | ~v_218 | ~v_1136 | ~v_1135 | ~v_217 | ~v_216 | ~v_167 | ~v_166 | ~v_1134 | ~v_1133 | ~v_163 | ~v_162 | ~v_155 | ~v_154 | v_1137;
assign x_8524 = v_1136 | ~v_125;
assign x_8525 = v_1136 | v_12;
assign x_8526 = v_1135 | v_125;
assign x_8527 = v_1135 | v_14;
assign x_8528 = v_1134 | v_125;
assign x_8529 = v_1134 | v_66;
assign x_8530 = v_1133 | ~v_125;
assign x_8531 = v_1133 | v_58;
assign x_8532 = v_25 | v_24 | v_19 | v_18 | v_17 | v_95 | v_109 | v_128 | v_122 | ~v_152 | ~v_151 | ~v_207 | ~v_206 | ~v_203 | ~v_202 | ~v_1131 | ~v_1130 | ~v_201 | ~v_200 | ~v_148 | ~v_147 | ~v_1129 | ~v_1128 | ~v_144 | ~v_143 | ~v_136 | ~v_135 | v_1132;
assign x_8533 = v_1131 | v_125;
assign x_8534 = v_1131 | v_15;
assign x_8535 = v_1130 | ~v_125;
assign x_8536 = v_1130 | v_11;
assign x_8537 = v_1129 | v_125;
assign x_8538 = v_1129 | v_41;
assign x_8539 = v_1128 | ~v_125;
assign x_8540 = v_1128 | v_33;
assign x_8541 = v_9 | v_4 | v_6 | v_8 | v_10 | v_3 | v_2 | ~v_1041 | ~v_1040 | ~v_1126 | v_1127;
assign x_8542 = v_1126 | ~v_1121;
assign x_8543 = v_1126 | ~v_1125;
assign x_8544 = v_125 | ~v_1037 | ~v_1022 | ~v_1006 | ~v_975 | ~v_974 | ~v_973 | ~v_972 | ~v_967 | ~v_1124 | ~v_1123 | v_1125;
assign x_8545 = v_1124 | ~v_881;
assign x_8546 = v_1124 | ~v_1095;
assign x_8547 = v_1123 | ~v_1122;
assign x_8548 = v_1123 | ~v_1059;
assign x_8549 = ~v_965 | ~v_1113 | ~v_964 | ~v_963 | ~v_1112 | v_1122;
assign x_8550 = ~v_586 | ~v_1120 | v_1121;
assign x_8551 = v_1120 | ~v_1118;
assign x_8552 = v_1120 | ~v_1119;
assign x_8553 = v_1120 | ~v_514;
assign x_8554 = v_1120 | ~v_519;
assign x_8555 = v_1120 | ~v_520;
assign x_8556 = v_1120 | ~v_521;
assign x_8557 = v_1120 | ~v_522;
assign x_8558 = ~v_1071 | ~v_428 | v_1119;
assign x_8559 = ~v_1047 | ~v_1117 | v_1118;
assign x_8560 = v_1117 | ~v_1088;
assign x_8561 = v_1117 | ~v_510;
assign x_8562 = v_1117 | ~v_511;
assign x_8563 = v_1117 | ~v_1089;
assign x_8564 = v_1117 | ~v_512;
assign x_8565 = v_9 | v_7 | v_4 | v_6 | v_10 | v_3 | v_2 | v_1 | ~v_1041 | ~v_1040 | ~v_1115 | v_1116;
assign x_8566 = v_1115 | ~v_1091;
assign x_8567 = v_1115 | ~v_1114;
assign x_8568 = v_125 | ~v_1037 | ~v_1022 | ~v_1006 | ~v_965 | ~v_1113 | ~v_964 | ~v_963 | ~v_1112 | ~v_1111 | ~v_1096 | v_1114;
assign x_8569 = v_1113 | ~v_971;
assign x_8570 = v_1113 | ~v_736;
assign x_8571 = v_1113 | ~v_698;
assign x_8572 = v_1113 | ~v_699;
assign x_8573 = v_1113 | ~v_700;
assign x_8574 = v_1113 | ~v_701;
assign x_8575 = v_1112 | ~v_1092;
assign x_8576 = v_1112 | ~v_857;
assign x_8577 = v_1112 | ~v_698;
assign x_8578 = v_1112 | ~v_699;
assign x_8579 = v_1112 | ~v_700;
assign x_8580 = v_1112 | ~v_701;
assign x_8581 = v_1111 | ~v_976;
assign x_8582 = v_1111 | ~v_1110;
assign x_8583 = ~v_1109 | ~v_1108 | ~v_1103 | ~v_1102 | ~v_1101 | v_1110;
assign x_8584 = v_1109 | ~v_857;
assign x_8585 = v_1109 | ~v_698;
assign x_8586 = v_1109 | ~v_699;
assign x_8587 = v_1109 | ~v_700;
assign x_8588 = v_1109 | ~v_701;
assign x_8589 = v_1108 | ~v_736;
assign x_8590 = v_1108 | ~v_1107;
assign x_8591 = v_1108 | ~v_698;
assign x_8592 = v_1108 | ~v_699;
assign x_8593 = v_1108 | ~v_700;
assign x_8594 = v_1108 | ~v_701;
assign x_8595 = ~v_1106 | ~v_1105 | ~v_1104 | v_1107;
assign x_8596 = v_1106 | ~v_956;
assign x_8597 = v_1106 | ~v_698;
assign x_8598 = v_1106 | ~v_699;
assign x_8599 = v_1106 | ~v_700;
assign x_8600 = v_1106 | ~v_701;
assign x_8601 = v_1105 | ~v_645;
assign x_8602 = v_1105 | ~v_935;
assign x_8603 = v_1105 | ~v_698;
assign x_8604 = v_1105 | ~v_699;
assign x_8605 = v_1105 | ~v_700;
assign x_8606 = v_1105 | ~v_701;
assign x_8607 = v_1104 | ~v_857;
assign x_8608 = v_1104 | ~v_916;
assign x_8609 = v_1104 | ~v_698;
assign x_8610 = v_1104 | ~v_699;
assign x_8611 = v_1104 | ~v_700;
assign x_8612 = v_1104 | ~v_701;
assign x_8613 = v_1103 | ~v_736;
assign x_8614 = v_1103 | ~v_956;
assign x_8615 = v_1103 | ~v_698;
assign x_8616 = v_1103 | ~v_699;
assign x_8617 = v_1103 | ~v_700;
assign x_8618 = v_1103 | ~v_701;
assign x_8619 = v_1102 | ~v_840;
assign x_8620 = v_1102 | ~v_645;
assign x_8621 = v_1102 | ~v_698;
assign x_8622 = v_1102 | ~v_699;
assign x_8623 = v_1102 | ~v_700;
assign x_8624 = v_1102 | ~v_701;
assign x_8625 = v_1101 | ~v_1100;
assign x_8626 = v_1101 | ~v_840;
assign x_8627 = v_1101 | ~v_698;
assign x_8628 = v_1101 | ~v_699;
assign x_8629 = v_1101 | ~v_700;
assign x_8630 = v_1101 | ~v_701;
assign x_8631 = ~v_1099 | ~v_1098 | ~v_1097 | v_1100;
assign x_8632 = v_1099 | ~v_645;
assign x_8633 = v_1099 | ~v_698;
assign x_8634 = v_1099 | ~v_699;
assign x_8635 = v_1099 | ~v_700;
assign x_8636 = v_1099 | ~v_701;
assign x_8637 = v_1098 | ~v_787;
assign x_8638 = v_1098 | ~v_956;
assign x_8639 = v_1098 | ~v_698;
assign x_8640 = v_1098 | ~v_699;
assign x_8641 = v_1098 | ~v_700;
assign x_8642 = v_1098 | ~v_701;
assign x_8643 = v_1097 | ~v_857;
assign x_8644 = v_1097 | ~v_770;
assign x_8645 = v_1097 | ~v_698;
assign x_8646 = v_1097 | ~v_699;
assign x_8647 = v_1097 | ~v_700;
assign x_8648 = v_1097 | ~v_701;
assign x_8649 = v_1096 | ~v_1095;
assign x_8650 = v_1096 | ~v_1058;
assign x_8651 = ~v_970 | ~v_969 | ~v_968 | ~v_1094 | ~v_1093 | v_1095;
assign x_8652 = v_1094 | ~v_966;
assign x_8653 = v_1094 | ~v_916;
assign x_8654 = v_1094 | ~v_698;
assign x_8655 = v_1094 | ~v_699;
assign x_8656 = v_1094 | ~v_700;
assign x_8657 = v_1094 | ~v_701;
assign x_8658 = v_1093 | ~v_1092;
assign x_8659 = v_1093 | ~v_956;
assign x_8660 = v_1093 | ~v_698;
assign x_8661 = v_1093 | ~v_699;
assign x_8662 = v_1093 | ~v_700;
assign x_8663 = v_1093 | ~v_701;
assign x_8664 = ~v_975 | ~v_974 | ~v_973 | v_1092;
assign x_8665 = ~v_586 | ~v_1090 | v_1091;
assign x_8666 = v_1090 | ~v_1072;
assign x_8667 = v_1090 | ~v_1087;
assign x_8668 = v_1090 | ~v_1088;
assign x_8669 = v_1090 | ~v_510;
assign x_8670 = v_1090 | ~v_511;
assign x_8671 = v_1090 | ~v_1089;
assign x_8672 = v_1090 | ~v_512;
assign x_8673 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_283 | ~v_518 | v_1089;
assign x_8674 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_404 | ~v_1068 | v_1088;
assign x_8675 = ~v_1086 | ~v_523 | v_1087;
assign x_8676 = v_1086 | ~v_1077;
assign x_8677 = v_1086 | ~v_1078;
assign x_8678 = v_1086 | ~v_1079;
assign x_8679 = v_1086 | ~v_1084;
assign x_8680 = v_1086 | ~v_1085;
assign x_8681 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_404 | v_1085;
assign x_8682 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_1083 | ~v_283 | v_1084;
assign x_8683 = v_1083 | ~v_1080;
assign x_8684 = v_1083 | ~v_1081;
assign x_8685 = v_1083 | ~v_1082;
assign x_8686 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_503 | v_1082;
assign x_8687 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_482 | ~v_192 | v_1081;
assign x_8688 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_463 | ~v_404 | v_1080;
assign x_8689 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_503 | ~v_283 | v_1079;
assign x_8690 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_192 | ~v_387 | v_1078;
assign x_8691 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_387 | ~v_1076 | v_1077;
assign x_8692 = v_1076 | ~v_1073;
assign x_8693 = v_1076 | ~v_1074;
assign x_8694 = v_1076 | ~v_1075;
assign x_8695 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_192 | v_1075;
assign x_8696 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_503 | ~v_334 | v_1074;
assign x_8697 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_317 | ~v_404 | v_1073;
assign x_8698 = ~v_1046 | ~v_1071 | v_1072;
assign x_8699 = v_1071 | ~v_1069;
assign x_8700 = v_1071 | ~v_1070;
assign x_8701 = v_1071 | ~v_515;
assign x_8702 = v_1071 | ~v_516;
assign x_8703 = v_1071 | ~v_517;
assign x_8704 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_463 | ~v_513 | v_1070;
assign x_8705 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_503 | ~v_1068 | v_1069;
assign x_8706 = v_1068 | ~v_520;
assign x_8707 = v_1068 | ~v_521;
assign x_8708 = v_1068 | ~v_522;
assign x_8709 = v_9 | v_5 | v_4 | v_8 | v_10 | v_3 | v_2 | ~v_1041 | ~v_1040 | ~v_1066 | v_1067;
assign x_8710 = v_1066 | ~v_1054;
assign x_8711 = v_1066 | ~v_1065;
assign x_8712 = v_125 | ~v_1037 | ~v_1022 | ~v_1006 | ~v_880 | ~v_879 | ~v_878 | ~v_877 | ~v_824 | ~v_1064 | ~v_1060 | v_1065;
assign x_8713 = v_1064 | ~v_976;
assign x_8714 = v_1064 | ~v_1063;
assign x_8715 = ~v_788 | ~v_771 | ~v_702 | ~v_1062 | ~v_1061 | v_1063;
assign x_8716 = v_1062 | ~v_860;
assign x_8717 = v_1062 | ~v_770;
assign x_8718 = v_1062 | ~v_698;
assign x_8719 = v_1062 | ~v_699;
assign x_8720 = v_1062 | ~v_700;
assign x_8721 = v_1062 | ~v_701;
assign x_8722 = v_1061 | ~v_1056;
assign x_8723 = v_1061 | ~v_645;
assign x_8724 = v_1061 | ~v_698;
assign x_8725 = v_1061 | ~v_699;
assign x_8726 = v_1061 | ~v_700;
assign x_8727 = v_1061 | ~v_701;
assign x_8728 = v_1060 | ~v_1058;
assign x_8729 = v_1060 | ~v_1059;
assign x_8730 = ~v_939 | ~v_983 | ~v_938 | ~v_937 | ~v_982 | v_1059;
assign x_8731 = ~v_859 | ~v_858 | ~v_841 | ~v_1057 | ~v_1055 | v_1058;
assign x_8732 = v_1057 | ~v_1056;
assign x_8733 = v_1057 | ~v_857;
assign x_8734 = v_1057 | ~v_698;
assign x_8735 = v_1057 | ~v_699;
assign x_8736 = v_1057 | ~v_700;
assign x_8737 = v_1057 | ~v_701;
assign x_8738 = ~v_880 | ~v_879 | ~v_878 | v_1056;
assign x_8739 = v_1055 | ~v_789;
assign x_8740 = v_1055 | ~v_840;
assign x_8741 = v_1055 | ~v_698;
assign x_8742 = v_1055 | ~v_699;
assign x_8743 = v_1055 | ~v_700;
assign x_8744 = v_1055 | ~v_701;
assign x_8745 = ~v_586 | ~v_1053 | v_1054;
assign x_8746 = v_1053 | ~v_1048;
assign x_8747 = v_1053 | ~v_1052;
assign x_8748 = v_1053 | ~v_371;
assign x_8749 = v_1053 | ~v_424;
assign x_8750 = v_1053 | ~v_425;
assign x_8751 = v_1053 | ~v_426;
assign x_8752 = v_1053 | ~v_427;
assign x_8753 = ~v_1051 | ~v_523 | v_1052;
assign x_8754 = v_1051 | ~v_1049;
assign x_8755 = v_1051 | ~v_1050;
assign x_8756 = v_1051 | ~v_249;
assign x_8757 = v_1051 | ~v_318;
assign x_8758 = v_1051 | ~v_335;
assign x_8759 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_317 | ~v_407 | v_1050;
assign x_8760 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_192 | ~v_1044 | v_1049;
assign x_8761 = ~v_1047 | ~v_1046 | v_1048;
assign x_8762 = v_1047 | ~v_529;
assign x_8763 = v_1047 | ~v_484;
assign x_8764 = v_1047 | ~v_485;
assign x_8765 = v_1047 | ~v_530;
assign x_8766 = v_1047 | ~v_486;
assign x_8767 = v_1046 | ~v_1043;
assign x_8768 = v_1046 | ~v_1045;
assign x_8769 = v_1046 | ~v_388;
assign x_8770 = v_1046 | ~v_405;
assign x_8771 = v_1046 | ~v_406;
assign x_8772 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_404 | ~v_1044 | v_1045;
assign x_8773 = v_1044 | ~v_425;
assign x_8774 = v_1044 | ~v_426;
assign x_8775 = v_1044 | ~v_427;
assign x_8776 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_387 | ~v_336 | v_1043;
assign x_8777 = v_9 | v_5 | v_4 | v_6 | v_8 | v_3 | v_2 | ~v_1041 | ~v_1040 | ~v_1039 | v_1042;
assign x_8778 = v_1041 | ~v_8;
assign x_8779 = v_1041 | ~v_7;
assign x_8780 = v_1041 | ~v_3;
assign x_8781 = v_1041 | ~v_2;
assign x_8782 = v_1041 | ~v_1;
assign x_8783 = v_1040 | ~v_10;
assign x_8784 = v_1040 | ~v_9;
assign x_8785 = v_1040 | ~v_6;
assign x_8786 = v_1040 | ~v_5;
assign x_8787 = v_1040 | ~v_4;
assign x_8788 = v_1039 | ~v_587;
assign x_8789 = v_1039 | ~v_1038;
assign x_8790 = v_125 | ~v_1037 | ~v_1022 | ~v_1006 | ~v_939 | ~v_983 | ~v_938 | ~v_937 | ~v_982 | ~v_981 | ~v_962 | v_1038;
assign x_8791 = v_1037 | ~v_1025;
assign x_8792 = v_1037 | ~v_1036;
assign x_8793 = v_124 | ~v_1035 | ~v_1031 | ~v_1027 | ~v_1026 | v_1036;
assign x_8794 = v_1035 | ~v_1034;
assign x_8795 = v_1035 | v_129;
assign x_8796 = v_98 | ~v_1033 | ~v_1032 | v_1034;
assign x_8797 = v_1033 | v_115;
assign x_8798 = v_1033 | v_119;
assign x_8799 = v_1032 | v_124;
assign x_8800 = v_1032 | v_130;
assign x_8801 = v_1031 | ~v_1030;
assign x_8802 = v_1031 | v_134;
assign x_8803 = v_115 | ~v_1029 | ~v_1028 | v_1030;
assign x_8804 = v_1029 | v_118;
assign x_8805 = v_1029 | v_98;
assign x_8806 = v_1028 | v_124;
assign x_8807 = v_1028 | v_133;
assign x_8808 = v_1027 | v_129;
assign x_8809 = v_1027 | v_98;
assign x_8810 = v_1026 | v_115;
assign x_8811 = v_1026 | v_134;
assign x_8812 = v_123 | ~v_1024 | ~v_989 | ~v_988 | ~v_1023 | v_1025;
assign x_8813 = v_1024 | ~v_1008;
assign x_8814 = v_1024 | v_114;
assign x_8815 = v_1023 | ~v_986;
assign x_8816 = v_1023 | v_97;
assign x_8817 = v_1022 | ~v_1010;
assign x_8818 = v_1022 | ~v_1021;
assign x_8819 = v_129 | ~v_1020 | ~v_1019 | ~v_1018 | ~v_1014 | v_1021;
assign x_8820 = v_1020 | v_124;
assign x_8821 = v_1020 | v_97;
assign x_8822 = v_1019 | v_118;
assign x_8823 = v_1019 | v_134;
assign x_8824 = v_1018 | ~v_1017;
assign x_8825 = v_1018 | v_134;
assign x_8826 = v_118 | ~v_1016 | ~v_1015 | v_1017;
assign x_8827 = v_1016 | v_115;
assign x_8828 = v_1016 | v_97;
assign x_8829 = v_1015 | v_129;
assign x_8830 = v_1015 | v_133;
assign x_8831 = v_1014 | ~v_1013;
assign x_8832 = v_1014 | v_124;
assign x_8833 = v_97 | ~v_1012 | ~v_1011 | v_1013;
assign x_8834 = v_1012 | v_118;
assign x_8835 = v_1012 | v_114;
assign x_8836 = v_1011 | v_123;
assign x_8837 = v_1011 | v_129;
assign x_8838 = v_130 | ~v_985 | ~v_984 | ~v_1009 | ~v_1007 | v_1010;
assign x_8839 = v_1009 | ~v_1008;
assign x_8840 = v_1009 | v_119;
assign x_8841 = v_133 | ~v_993 | ~v_992 | v_1008;
assign x_8842 = v_1007 | ~v_990;
assign x_8843 = v_1007 | v_98;
assign x_8844 = v_1006 | ~v_994;
assign x_8845 = v_1006 | ~v_1005;
assign x_8846 = v_134 | ~v_1004 | ~v_1003 | ~v_1002 | ~v_998 | v_1005;
assign x_8847 = v_1004 | v_124;
assign x_8848 = v_1004 | v_114;
assign x_8849 = v_1003 | v_129;
assign x_8850 = v_1003 | v_119;
assign x_8851 = v_1002 | ~v_1001;
assign x_8852 = v_1002 | v_124;
assign x_8853 = v_114 | ~v_1000 | ~v_999 | v_1001;
assign x_8854 = v_1000 | v_119;
assign x_8855 = v_1000 | v_97;
assign x_8856 = v_999 | v_123;
assign x_8857 = v_999 | v_134;
assign x_8858 = v_998 | ~v_997;
assign x_8859 = v_998 | v_129;
assign x_8860 = v_119 | ~v_996 | ~v_995 | v_997;
assign x_8861 = v_996 | v_114;
assign x_8862 = v_996 | v_98;
assign x_8863 = v_995 | v_134;
assign x_8864 = v_995 | v_130;
assign x_8865 = v_133 | ~v_993 | ~v_992 | ~v_991 | ~v_987 | v_994;
assign x_8866 = v_993 | v_123;
assign x_8867 = v_993 | v_115;
assign x_8868 = v_992 | v_118;
assign x_8869 = v_992 | v_130;
assign x_8870 = v_991 | ~v_990;
assign x_8871 = v_991 | v_115;
assign x_8872 = v_123 | ~v_989 | ~v_988 | v_990;
assign x_8873 = v_989 | v_130;
assign x_8874 = v_989 | v_97;
assign x_8875 = v_988 | v_133;
assign x_8876 = v_988 | v_114;
assign x_8877 = v_987 | ~v_986;
assign x_8878 = v_987 | v_118;
assign x_8879 = v_130 | ~v_985 | ~v_984 | v_986;
assign x_8880 = v_985 | v_123;
assign x_8881 = v_985 | v_98;
assign x_8882 = v_984 | v_133;
assign x_8883 = v_984 | v_119;
assign x_8884 = v_983 | ~v_697;
assign x_8885 = v_983 | ~v_978;
assign x_8886 = v_983 | ~v_698;
assign x_8887 = v_983 | ~v_699;
assign x_8888 = v_983 | ~v_700;
assign x_8889 = v_983 | ~v_701;
assign x_8890 = v_982 | ~v_919;
assign x_8891 = v_982 | ~v_823;
assign x_8892 = v_982 | ~v_698;
assign x_8893 = v_982 | ~v_699;
assign x_8894 = v_982 | ~v_700;
assign x_8895 = v_982 | ~v_701;
assign x_8896 = v_981 | ~v_976;
assign x_8897 = v_981 | ~v_980;
assign x_8898 = ~v_918 | ~v_917 | ~v_882 | ~v_979 | ~v_977 | v_980;
assign x_8899 = v_979 | ~v_787;
assign x_8900 = v_979 | ~v_978;
assign x_8901 = v_979 | ~v_698;
assign x_8902 = v_979 | ~v_699;
assign x_8903 = v_979 | ~v_700;
assign x_8904 = v_979 | ~v_701;
assign x_8905 = ~v_960 | ~v_959 | ~v_958 | v_978;
assign x_8906 = v_977 | ~v_645;
assign x_8907 = v_977 | ~v_940;
assign x_8908 = v_977 | ~v_698;
assign x_8909 = v_977 | ~v_699;
assign x_8910 = v_977 | ~v_700;
assign x_8911 = v_977 | ~v_701;
assign x_8912 = ~v_975 | ~v_974 | ~v_973 | ~v_972 | ~v_967 | v_976;
assign x_8913 = v_975 | ~v_823;
assign x_8914 = v_975 | ~v_698;
assign x_8915 = v_975 | ~v_699;
assign x_8916 = v_975 | ~v_700;
assign x_8917 = v_975 | ~v_701;
assign x_8918 = v_974 | ~v_697;
assign x_8919 = v_974 | ~v_935;
assign x_8920 = v_974 | ~v_698;
assign x_8921 = v_974 | ~v_699;
assign x_8922 = v_974 | ~v_700;
assign x_8923 = v_974 | ~v_701;
assign x_8924 = v_973 | ~v_840;
assign x_8925 = v_973 | ~v_876;
assign x_8926 = v_973 | ~v_698;
assign x_8927 = v_973 | ~v_699;
assign x_8928 = v_973 | ~v_700;
assign x_8929 = v_973 | ~v_701;
assign x_8930 = v_972 | ~v_971;
assign x_8931 = v_972 | ~v_697;
assign x_8932 = v_972 | ~v_698;
assign x_8933 = v_972 | ~v_699;
assign x_8934 = v_972 | ~v_700;
assign x_8935 = v_972 | ~v_701;
assign x_8936 = ~v_970 | ~v_969 | ~v_968 | v_971;
assign x_8937 = v_970 | ~v_935;
assign x_8938 = v_970 | ~v_698;
assign x_8939 = v_970 | ~v_699;
assign x_8940 = v_970 | ~v_700;
assign x_8941 = v_970 | ~v_701;
assign x_8942 = v_969 | ~v_840;
assign x_8943 = v_969 | ~v_916;
assign x_8944 = v_969 | ~v_698;
assign x_8945 = v_969 | ~v_699;
assign x_8946 = v_969 | ~v_700;
assign x_8947 = v_969 | ~v_701;
assign x_8948 = v_968 | ~v_823;
assign x_8949 = v_968 | ~v_956;
assign x_8950 = v_968 | ~v_698;
assign x_8951 = v_968 | ~v_699;
assign x_8952 = v_968 | ~v_700;
assign x_8953 = v_968 | ~v_701;
assign x_8954 = v_967 | ~v_966;
assign x_8955 = v_967 | ~v_876;
assign x_8956 = v_967 | ~v_698;
assign x_8957 = v_967 | ~v_699;
assign x_8958 = v_967 | ~v_700;
assign x_8959 = v_967 | ~v_701;
assign x_8960 = ~v_965 | ~v_964 | ~v_963 | v_966;
assign x_8961 = v_965 | ~v_840;
assign x_8962 = v_965 | ~v_698;
assign x_8963 = v_965 | ~v_699;
assign x_8964 = v_965 | ~v_700;
assign x_8965 = v_965 | ~v_701;
assign x_8966 = v_964 | ~v_736;
assign x_8967 = v_964 | ~v_935;
assign x_8968 = v_964 | ~v_698;
assign x_8969 = v_964 | ~v_699;
assign x_8970 = v_964 | ~v_700;
assign x_8971 = v_964 | ~v_701;
assign x_8972 = v_963 | ~v_857;
assign x_8973 = v_963 | ~v_823;
assign x_8974 = v_963 | ~v_698;
assign x_8975 = v_963 | ~v_699;
assign x_8976 = v_963 | ~v_700;
assign x_8977 = v_963 | ~v_701;
assign x_8978 = v_962 | ~v_881;
assign x_8979 = v_962 | ~v_961;
assign x_8980 = ~v_960 | ~v_959 | ~v_958 | ~v_957 | ~v_936 | v_961;
assign x_8981 = v_960 | ~v_770;
assign x_8982 = v_960 | ~v_935;
assign x_8983 = v_960 | ~v_698;
assign x_8984 = v_960 | ~v_699;
assign x_8985 = v_960 | ~v_700;
assign x_8986 = v_960 | ~v_701;
assign x_8987 = v_959 | ~v_916;
assign x_8988 = v_959 | ~v_698;
assign x_8989 = v_959 | ~v_699;
assign x_8990 = v_959 | ~v_700;
assign x_8991 = v_959 | ~v_701;
assign x_8992 = v_958 | ~v_956;
assign x_8993 = v_958 | ~v_876;
assign x_8994 = v_958 | ~v_698;
assign x_8995 = v_958 | ~v_699;
assign x_8996 = v_958 | ~v_700;
assign x_8997 = v_958 | ~v_701;
assign x_8998 = v_957 | ~v_940;
assign x_8999 = v_957 | ~v_956;
assign x_9000 = v_957 | ~v_698;
assign x_9001 = v_957 | ~v_699;
assign x_9002 = v_957 | ~v_700;
assign x_9003 = v_957 | ~v_701;
assign x_9004 = ~v_955 | ~v_950 | ~v_945 | v_956;
assign x_9005 = v_955 | ~v_626;
assign x_9006 = v_955 | ~v_627;
assign x_9007 = v_955 | ~v_905;
assign x_9008 = v_955 | ~v_951;
assign x_9009 = v_955 | ~v_952;
assign x_9010 = v_955 | ~v_906;
assign x_9011 = v_955 | ~v_907;
assign x_9012 = v_955 | ~v_953;
assign x_9013 = v_955 | ~v_954;
assign x_9014 = v_955 | ~v_634;
assign x_9015 = v_955 | ~v_635;
assign x_9016 = v_955 | ~v_638;
assign x_9017 = v_955 | ~v_639;
assign x_9018 = v_955 | ~v_911;
assign x_9019 = v_955 | ~v_912;
assign x_9020 = v_955 | ~v_642;
assign x_9021 = v_955 | ~v_643;
assign x_9022 = v_955 | ~v_913;
assign x_9023 = v_955 | ~v_127;
assign x_9024 = v_955 | ~v_113;
assign x_9025 = v_955 | ~v_112;
assign x_9026 = v_955 | ~v_106;
assign x_9027 = v_955 | ~v_104;
assign x_9028 = v_955 | ~v_76;
assign x_9029 = v_955 | ~v_75;
assign x_9030 = v_955 | ~v_73;
assign x_9031 = v_955 | ~v_70;
assign x_9032 = ~v_91 | ~v_129 | v_954;
assign x_9033 = ~v_83 | v_129 | v_953;
assign x_9034 = ~v_16 | ~v_130 | v_952;
assign x_9035 = ~v_13 | v_130 | v_951;
assign x_9036 = v_950 | ~v_607;
assign x_9037 = v_950 | ~v_608;
assign x_9038 = v_950 | ~v_894;
assign x_9039 = v_950 | ~v_895;
assign x_9040 = v_950 | ~v_946;
assign x_9041 = v_950 | ~v_947;
assign x_9042 = v_950 | ~v_948;
assign x_9043 = v_950 | ~v_949;
assign x_9044 = v_950 | ~v_615;
assign x_9045 = v_950 | ~v_616;
assign x_9046 = v_950 | ~v_619;
assign x_9047 = v_950 | ~v_620;
assign x_9048 = v_950 | ~v_898;
assign x_9049 = v_950 | ~v_899;
assign x_9050 = v_950 | ~v_623;
assign x_9051 = v_950 | ~v_624;
assign x_9052 = v_950 | ~v_900;
assign x_9053 = v_950 | ~v_902;
assign x_9054 = v_950 | ~v_126;
assign x_9055 = v_950 | ~v_111;
assign x_9056 = v_950 | ~v_110;
assign x_9057 = v_950 | ~v_102;
assign x_9058 = v_950 | ~v_100;
assign x_9059 = v_950 | ~v_51;
assign x_9060 = v_950 | ~v_50;
assign x_9061 = v_950 | ~v_48;
assign x_9062 = v_950 | ~v_45;
assign x_9063 = ~v_66 | ~v_129 | v_949;
assign x_9064 = ~v_58 | v_129 | v_948;
assign x_9065 = ~v_14 | ~v_130 | v_947;
assign x_9066 = ~v_12 | v_130 | v_946;
assign x_9067 = v_945 | ~v_588;
assign x_9068 = v_945 | ~v_589;
assign x_9069 = v_945 | ~v_883;
assign x_9070 = v_945 | ~v_884;
assign x_9071 = v_945 | ~v_941;
assign x_9072 = v_945 | ~v_942;
assign x_9073 = v_945 | ~v_885;
assign x_9074 = v_945 | ~v_943;
assign x_9075 = v_945 | ~v_944;
assign x_9076 = v_945 | ~v_596;
assign x_9077 = v_945 | ~v_597;
assign x_9078 = v_945 | ~v_600;
assign x_9079 = v_945 | ~v_601;
assign x_9080 = v_945 | ~v_888;
assign x_9081 = v_945 | ~v_889;
assign x_9082 = v_945 | ~v_604;
assign x_9083 = v_945 | ~v_605;
assign x_9084 = v_945 | ~v_890;
assign x_9085 = v_945 | ~v_122;
assign x_9086 = v_945 | ~v_109;
assign x_9087 = v_945 | ~v_108;
assign x_9088 = v_945 | ~v_95;
assign x_9089 = v_945 | ~v_93;
assign x_9090 = v_945 | ~v_25;
assign x_9091 = v_945 | ~v_24;
assign x_9092 = v_945 | ~v_22;
assign x_9093 = v_945 | ~v_19;
assign x_9094 = ~v_41 | ~v_129 | v_944;
assign x_9095 = ~v_33 | v_129 | v_943;
assign x_9096 = ~v_15 | ~v_130 | v_942;
assign x_9097 = ~v_11 | v_130 | v_941;
assign x_9098 = ~v_939 | ~v_938 | ~v_937 | v_940;
assign x_9099 = v_939 | ~v_876;
assign x_9100 = v_939 | ~v_698;
assign x_9101 = v_939 | ~v_699;
assign x_9102 = v_939 | ~v_700;
assign x_9103 = v_939 | ~v_701;
assign x_9104 = v_938 | ~v_697;
assign x_9105 = v_938 | ~v_916;
assign x_9106 = v_938 | ~v_698;
assign x_9107 = v_938 | ~v_699;
assign x_9108 = v_938 | ~v_700;
assign x_9109 = v_938 | ~v_701;
assign x_9110 = v_937 | ~v_823;
assign x_9111 = v_937 | ~v_770;
assign x_9112 = v_937 | ~v_698;
assign x_9113 = v_937 | ~v_699;
assign x_9114 = v_937 | ~v_700;
assign x_9115 = v_937 | ~v_701;
assign x_9116 = v_936 | ~v_919;
assign x_9117 = v_936 | ~v_935;
assign x_9118 = v_936 | ~v_698;
assign x_9119 = v_936 | ~v_699;
assign x_9120 = v_936 | ~v_700;
assign x_9121 = v_936 | ~v_701;
assign x_9122 = ~v_934 | ~v_929 | ~v_924 | v_935;
assign x_9123 = v_934 | ~v_905;
assign x_9124 = v_934 | ~v_814;
assign x_9125 = v_934 | ~v_815;
assign x_9126 = v_934 | ~v_930;
assign x_9127 = v_934 | ~v_931;
assign x_9128 = v_934 | ~v_932;
assign x_9129 = v_934 | ~v_933;
assign x_9130 = v_934 | ~v_906;
assign x_9131 = v_934 | ~v_907;
assign x_9132 = v_934 | ~v_818;
assign x_9133 = v_934 | ~v_819;
assign x_9134 = v_934 | ~v_911;
assign x_9135 = v_934 | ~v_912;
assign x_9136 = v_934 | ~v_820;
assign x_9137 = v_934 | ~v_642;
assign x_9138 = v_934 | ~v_643;
assign x_9139 = v_934 | ~v_821;
assign x_9140 = v_934 | ~v_913;
assign x_9141 = v_934 | ~v_113;
assign x_9142 = v_934 | ~v_112;
assign x_9143 = v_934 | ~v_107;
assign x_9144 = v_934 | ~v_106;
assign x_9145 = v_934 | ~v_105;
assign x_9146 = v_934 | ~v_104;
assign x_9147 = v_934 | ~v_76;
assign x_9148 = v_934 | ~v_74;
assign x_9149 = v_934 | ~v_73;
assign x_9150 = ~v_91 | ~v_118 | v_933;
assign x_9151 = ~v_83 | v_118 | v_932;
assign x_9152 = ~v_16 | ~v_119 | v_931;
assign x_9153 = ~v_13 | v_119 | v_930;
assign x_9154 = v_929 | ~v_894;
assign x_9155 = v_929 | ~v_895;
assign x_9156 = v_929 | ~v_803;
assign x_9157 = v_929 | ~v_804;
assign x_9158 = v_929 | ~v_925;
assign x_9159 = v_929 | ~v_926;
assign x_9160 = v_929 | ~v_807;
assign x_9161 = v_929 | ~v_808;
assign x_9162 = v_929 | ~v_927;
assign x_9163 = v_929 | ~v_928;
assign x_9164 = v_929 | ~v_898;
assign x_9165 = v_929 | ~v_899;
assign x_9166 = v_929 | ~v_809;
assign x_9167 = v_929 | ~v_810;
assign x_9168 = v_929 | ~v_623;
assign x_9169 = v_929 | ~v_624;
assign x_9170 = v_929 | ~v_900;
assign x_9171 = v_929 | ~v_902;
assign x_9172 = v_929 | ~v_111;
assign x_9173 = v_929 | ~v_110;
assign x_9174 = v_929 | ~v_103;
assign x_9175 = v_929 | ~v_102;
assign x_9176 = v_929 | ~v_101;
assign x_9177 = v_929 | ~v_100;
assign x_9178 = v_929 | ~v_51;
assign x_9179 = v_929 | ~v_49;
assign x_9180 = v_929 | ~v_48;
assign x_9181 = ~v_12 | v_119 | v_928;
assign x_9182 = ~v_14 | ~v_119 | v_927;
assign x_9183 = ~v_66 | ~v_118 | v_926;
assign x_9184 = ~v_58 | v_118 | v_925;
assign x_9185 = v_924 | ~v_883;
assign x_9186 = v_924 | ~v_884;
assign x_9187 = v_924 | ~v_792;
assign x_9188 = v_924 | ~v_793;
assign x_9189 = v_924 | ~v_920;
assign x_9190 = v_924 | ~v_921;
assign x_9191 = v_924 | ~v_885;
assign x_9192 = v_924 | ~v_796;
assign x_9193 = v_924 | ~v_797;
assign x_9194 = v_924 | ~v_922;
assign x_9195 = v_924 | ~v_888;
assign x_9196 = v_924 | ~v_889;
assign x_9197 = v_924 | ~v_798;
assign x_9198 = v_924 | ~v_799;
assign x_9199 = v_924 | ~v_604;
assign x_9200 = v_924 | ~v_605;
assign x_9201 = v_924 | ~v_890;
assign x_9202 = v_924 | ~v_923;
assign x_9203 = v_924 | ~v_109;
assign x_9204 = v_924 | ~v_108;
assign x_9205 = v_924 | ~v_96;
assign x_9206 = v_924 | ~v_95;
assign x_9207 = v_924 | ~v_94;
assign x_9208 = v_924 | ~v_93;
assign x_9209 = v_924 | ~v_25;
assign x_9210 = v_924 | ~v_23;
assign x_9211 = v_924 | ~v_22;
assign x_9212 = ~v_11 | v_119 | v_923;
assign x_9213 = ~v_15 | ~v_119 | v_922;
assign x_9214 = ~v_41 | ~v_118 | v_921;
assign x_9215 = ~v_33 | v_118 | v_920;
assign x_9216 = ~v_918 | ~v_917 | ~v_882 | v_919;
assign x_9217 = v_918 | ~v_770;
assign x_9218 = v_918 | ~v_698;
assign x_9219 = v_918 | ~v_699;
assign x_9220 = v_918 | ~v_700;
assign x_9221 = v_918 | ~v_701;
assign x_9222 = v_917 | ~v_787;
assign x_9223 = v_917 | ~v_916;
assign x_9224 = v_917 | ~v_698;
assign x_9225 = v_917 | ~v_699;
assign x_9226 = v_917 | ~v_700;
assign x_9227 = v_917 | ~v_701;
assign x_9228 = ~v_915 | ~v_904 | ~v_893 | v_916;
assign x_9229 = v_915 | ~v_905;
assign x_9230 = v_915 | ~v_759;
assign x_9231 = v_915 | ~v_760;
assign x_9232 = v_915 | ~v_906;
assign x_9233 = v_915 | ~v_907;
assign x_9234 = v_915 | ~v_908;
assign x_9235 = v_915 | ~v_909;
assign x_9236 = v_915 | ~v_910;
assign x_9237 = v_915 | ~v_763;
assign x_9238 = v_915 | ~v_764;
assign x_9239 = v_915 | ~v_911;
assign x_9240 = v_915 | ~v_912;
assign x_9241 = v_915 | ~v_767;
assign x_9242 = v_915 | ~v_768;
assign x_9243 = v_915 | ~v_642;
assign x_9244 = v_915 | ~v_643;
assign x_9245 = v_915 | ~v_913;
assign x_9246 = v_915 | ~v_914;
assign x_9247 = v_915 | ~v_121;
assign x_9248 = v_915 | ~v_113;
assign x_9249 = v_915 | ~v_112;
assign x_9250 = v_915 | ~v_105;
assign x_9251 = v_915 | ~v_104;
assign x_9252 = v_915 | ~v_75;
assign x_9253 = v_915 | ~v_74;
assign x_9254 = v_915 | ~v_73;
assign x_9255 = v_915 | ~v_72;
assign x_9256 = ~v_13 | v_98 | v_914;
assign x_9257 = ~v_88 | ~v_130 | v_913;
assign x_9258 = ~v_86 | ~v_129 | v_912;
assign x_9259 = ~v_78 | v_129 | v_911;
assign x_9260 = ~v_16 | ~v_98 | v_910;
assign x_9261 = ~v_91 | ~v_97 | v_909;
assign x_9262 = ~v_83 | v_97 | v_908;
assign x_9263 = ~v_89 | ~v_99 | v_907;
assign x_9264 = ~v_81 | v_99 | v_906;
assign x_9265 = ~v_80 | v_130 | v_905;
assign x_9266 = v_904 | ~v_894;
assign x_9267 = v_904 | ~v_895;
assign x_9268 = v_904 | ~v_748;
assign x_9269 = v_904 | ~v_749;
assign x_9270 = v_904 | ~v_896;
assign x_9271 = v_904 | ~v_750;
assign x_9272 = v_904 | ~v_897;
assign x_9273 = v_904 | ~v_898;
assign x_9274 = v_904 | ~v_899;
assign x_9275 = v_904 | ~v_755;
assign x_9276 = v_904 | ~v_756;
assign x_9277 = v_904 | ~v_623;
assign x_9278 = v_904 | ~v_624;
assign x_9279 = v_904 | ~v_757;
assign x_9280 = v_904 | ~v_900;
assign x_9281 = v_904 | ~v_901;
assign x_9282 = v_904 | ~v_902;
assign x_9283 = v_904 | ~v_903;
assign x_9284 = v_904 | ~v_120;
assign x_9285 = v_904 | ~v_111;
assign x_9286 = v_904 | ~v_110;
assign x_9287 = v_904 | ~v_101;
assign x_9288 = v_904 | ~v_100;
assign x_9289 = v_904 | ~v_50;
assign x_9290 = v_904 | ~v_49;
assign x_9291 = v_904 | ~v_48;
assign x_9292 = v_904 | ~v_47;
assign x_9293 = ~v_58 | v_97 | v_903;
assign x_9294 = ~v_64 | ~v_99 | v_902;
assign x_9295 = ~v_12 | v_98 | v_901;
assign x_9296 = ~v_56 | v_99 | v_900;
assign x_9297 = ~v_61 | ~v_129 | v_899;
assign x_9298 = ~v_53 | v_129 | v_898;
assign x_9299 = ~v_14 | ~v_98 | v_897;
assign x_9300 = ~v_66 | ~v_97 | v_896;
assign x_9301 = ~v_63 | ~v_130 | v_895;
assign x_9302 = ~v_55 | v_130 | v_894;
assign x_9303 = v_893 | ~v_883;
assign x_9304 = v_893 | ~v_884;
assign x_9305 = v_893 | ~v_737;
assign x_9306 = v_893 | ~v_738;
assign x_9307 = v_893 | ~v_885;
assign x_9308 = v_893 | ~v_886;
assign x_9309 = v_893 | ~v_887;
assign x_9310 = v_893 | ~v_739;
assign x_9311 = v_893 | ~v_888;
assign x_9312 = v_893 | ~v_889;
assign x_9313 = v_893 | ~v_744;
assign x_9314 = v_893 | ~v_745;
assign x_9315 = v_893 | ~v_604;
assign x_9316 = v_893 | ~v_605;
assign x_9317 = v_893 | ~v_746;
assign x_9318 = v_893 | ~v_890;
assign x_9319 = v_893 | ~v_891;
assign x_9320 = v_893 | ~v_892;
assign x_9321 = v_893 | ~v_117;
assign x_9322 = v_893 | ~v_109;
assign x_9323 = v_893 | ~v_108;
assign x_9324 = v_893 | ~v_94;
assign x_9325 = v_893 | ~v_93;
assign x_9326 = v_893 | ~v_24;
assign x_9327 = v_893 | ~v_23;
assign x_9328 = v_893 | ~v_22;
assign x_9329 = v_893 | ~v_21;
assign x_9330 = ~v_41 | ~v_97 | v_892;
assign x_9331 = ~v_33 | v_97 | v_891;
assign x_9332 = ~v_31 | v_99 | v_890;
assign x_9333 = ~v_36 | ~v_129 | v_889;
assign x_9334 = ~v_28 | v_129 | v_888;
assign x_9335 = ~v_15 | ~v_98 | v_887;
assign x_9336 = ~v_11 | v_98 | v_886;
assign x_9337 = ~v_39 | ~v_99 | v_885;
assign x_9338 = ~v_38 | ~v_130 | v_884;
assign x_9339 = ~v_30 | v_130 | v_883;
assign x_9340 = v_882 | ~v_645;
assign x_9341 = v_882 | ~v_876;
assign x_9342 = v_882 | ~v_698;
assign x_9343 = v_882 | ~v_699;
assign x_9344 = v_882 | ~v_700;
assign x_9345 = v_882 | ~v_701;
assign x_9346 = ~v_880 | ~v_879 | ~v_878 | ~v_877 | ~v_824 | v_881;
assign x_9347 = v_880 | ~v_697;
assign x_9348 = v_880 | ~v_698;
assign x_9349 = v_880 | ~v_699;
assign x_9350 = v_880 | ~v_700;
assign x_9351 = v_880 | ~v_701;
assign x_9352 = v_879 | ~v_736;
assign x_9353 = v_879 | ~v_876;
assign x_9354 = v_879 | ~v_698;
assign x_9355 = v_879 | ~v_699;
assign x_9356 = v_879 | ~v_700;
assign x_9357 = v_879 | ~v_701;
assign x_9358 = v_878 | ~v_787;
assign x_9359 = v_878 | ~v_823;
assign x_9360 = v_878 | ~v_698;
assign x_9361 = v_878 | ~v_699;
assign x_9362 = v_878 | ~v_700;
assign x_9363 = v_878 | ~v_701;
assign x_9364 = v_877 | ~v_860;
assign x_9365 = v_877 | ~v_876;
assign x_9366 = v_877 | ~v_698;
assign x_9367 = v_877 | ~v_699;
assign x_9368 = v_877 | ~v_700;
assign x_9369 = v_877 | ~v_701;
assign x_9370 = ~v_875 | ~v_870 | ~v_865 | v_876;
assign x_9371 = v_875 | ~v_759;
assign x_9372 = v_875 | ~v_760;
assign x_9373 = v_875 | ~v_871;
assign x_9374 = v_875 | ~v_872;
assign x_9375 = v_875 | ~v_873;
assign x_9376 = v_875 | ~v_874;
assign x_9377 = v_875 | ~v_763;
assign x_9378 = v_875 | ~v_764;
assign x_9379 = v_875 | ~v_688;
assign x_9380 = v_875 | ~v_689;
assign x_9381 = v_875 | ~v_690;
assign x_9382 = v_875 | ~v_691;
assign x_9383 = v_875 | ~v_767;
assign x_9384 = v_875 | ~v_768;
assign x_9385 = v_875 | ~v_694;
assign x_9386 = v_875 | ~v_695;
assign x_9387 = v_875 | ~v_642;
assign x_9388 = v_875 | ~v_643;
assign x_9389 = v_875 | ~v_132;
assign x_9390 = v_875 | ~v_113;
assign x_9391 = v_875 | ~v_105;
assign x_9392 = v_875 | ~v_104;
assign x_9393 = v_875 | ~v_76;
assign x_9394 = v_875 | ~v_75;
assign x_9395 = v_875 | ~v_74;
assign x_9396 = v_875 | ~v_72;
assign x_9397 = v_875 | ~v_68;
assign x_9398 = ~v_91 | ~v_123 | v_874;
assign x_9399 = ~v_83 | v_123 | v_873;
assign x_9400 = ~v_16 | ~v_124 | v_872;
assign x_9401 = ~v_13 | v_124 | v_871;
assign x_9402 = v_870 | ~v_748;
assign x_9403 = v_870 | ~v_749;
assign x_9404 = v_870 | ~v_866;
assign x_9405 = v_870 | ~v_867;
assign x_9406 = v_870 | ~v_750;
assign x_9407 = v_870 | ~v_868;
assign x_9408 = v_870 | ~v_669;
assign x_9409 = v_870 | ~v_670;
assign x_9410 = v_870 | ~v_869;
assign x_9411 = v_870 | ~v_671;
assign x_9412 = v_870 | ~v_672;
assign x_9413 = v_870 | ~v_755;
assign x_9414 = v_870 | ~v_756;
assign x_9415 = v_870 | ~v_675;
assign x_9416 = v_870 | ~v_676;
assign x_9417 = v_870 | ~v_623;
assign x_9418 = v_870 | ~v_624;
assign x_9419 = v_870 | ~v_757;
assign x_9420 = v_870 | ~v_131;
assign x_9421 = v_870 | ~v_111;
assign x_9422 = v_870 | ~v_101;
assign x_9423 = v_870 | ~v_100;
assign x_9424 = v_870 | ~v_51;
assign x_9425 = v_870 | ~v_50;
assign x_9426 = v_870 | ~v_49;
assign x_9427 = v_870 | ~v_47;
assign x_9428 = v_870 | ~v_43;
assign x_9429 = ~v_12 | v_124 | v_869;
assign x_9430 = ~v_14 | ~v_124 | v_868;
assign x_9431 = ~v_66 | ~v_123 | v_867;
assign x_9432 = ~v_58 | v_123 | v_866;
assign x_9433 = v_865 | ~v_737;
assign x_9434 = v_865 | ~v_738;
assign x_9435 = v_865 | ~v_861;
assign x_9436 = v_865 | ~v_862;
assign x_9437 = v_865 | ~v_739;
assign x_9438 = v_865 | ~v_653;
assign x_9439 = v_865 | ~v_654;
assign x_9440 = v_865 | ~v_863;
assign x_9441 = v_865 | ~v_864;
assign x_9442 = v_865 | ~v_655;
assign x_9443 = v_865 | ~v_656;
assign x_9444 = v_865 | ~v_744;
assign x_9445 = v_865 | ~v_745;
assign x_9446 = v_865 | ~v_659;
assign x_9447 = v_865 | ~v_660;
assign x_9448 = v_865 | ~v_604;
assign x_9449 = v_865 | ~v_605;
assign x_9450 = v_865 | ~v_746;
assign x_9451 = v_865 | ~v_128;
assign x_9452 = v_865 | ~v_109;
assign x_9453 = v_865 | ~v_94;
assign x_9454 = v_865 | ~v_93;
assign x_9455 = v_865 | ~v_25;
assign x_9456 = v_865 | ~v_24;
assign x_9457 = v_865 | ~v_23;
assign x_9458 = v_865 | ~v_21;
assign x_9459 = v_865 | ~v_17;
assign x_9460 = ~v_15 | ~v_124 | v_864;
assign x_9461 = ~v_11 | v_124 | v_863;
assign x_9462 = ~v_41 | ~v_123 | v_862;
assign x_9463 = ~v_33 | v_123 | v_861;
assign x_9464 = ~v_859 | ~v_858 | ~v_841 | v_860;
assign x_9465 = v_859 | ~v_736;
assign x_9466 = v_859 | ~v_698;
assign x_9467 = v_859 | ~v_699;
assign x_9468 = v_859 | ~v_700;
assign x_9469 = v_859 | ~v_701;
assign x_9470 = v_858 | ~v_857;
assign x_9471 = v_858 | ~v_697;
assign x_9472 = v_858 | ~v_698;
assign x_9473 = v_858 | ~v_699;
assign x_9474 = v_858 | ~v_700;
assign x_9475 = v_858 | ~v_701;
assign x_9476 = ~v_856 | ~v_851 | ~v_846 | v_857;
assign x_9477 = v_856 | ~v_626;
assign x_9478 = v_856 | ~v_627;
assign x_9479 = v_856 | ~v_852;
assign x_9480 = v_856 | ~v_853;
assign x_9481 = v_856 | ~v_726;
assign x_9482 = v_856 | ~v_634;
assign x_9483 = v_856 | ~v_635;
assign x_9484 = v_856 | ~v_854;
assign x_9485 = v_856 | ~v_855;
assign x_9486 = v_856 | ~v_638;
assign x_9487 = v_856 | ~v_639;
assign x_9488 = v_856 | ~v_729;
assign x_9489 = v_856 | ~v_730;
assign x_9490 = v_856 | ~v_731;
assign x_9491 = v_856 | ~v_732;
assign x_9492 = v_856 | ~v_733;
assign x_9493 = v_856 | ~v_642;
assign x_9494 = v_856 | ~v_643;
assign x_9495 = v_856 | ~v_127;
assign x_9496 = v_856 | ~v_112;
assign x_9497 = v_856 | ~v_106;
assign x_9498 = v_856 | ~v_104;
assign x_9499 = v_856 | ~v_76;
assign x_9500 = v_856 | ~v_75;
assign x_9501 = v_856 | ~v_73;
assign x_9502 = v_856 | ~v_71;
assign x_9503 = v_856 | ~v_70;
assign x_9504 = ~v_91 | ~v_124 | v_855;
assign x_9505 = ~v_83 | v_124 | v_854;
assign x_9506 = ~v_16 | ~v_123 | v_853;
assign x_9507 = ~v_13 | v_123 | v_852;
assign x_9508 = v_851 | ~v_607;
assign x_9509 = v_851 | ~v_608;
assign x_9510 = v_851 | ~v_847;
assign x_9511 = v_851 | ~v_848;
assign x_9512 = v_851 | ~v_714;
assign x_9513 = v_851 | ~v_615;
assign x_9514 = v_851 | ~v_616;
assign x_9515 = v_851 | ~v_849;
assign x_9516 = v_851 | ~v_850;
assign x_9517 = v_851 | ~v_619;
assign x_9518 = v_851 | ~v_620;
assign x_9519 = v_851 | ~v_716;
assign x_9520 = v_851 | ~v_717;
assign x_9521 = v_851 | ~v_719;
assign x_9522 = v_851 | ~v_720;
assign x_9523 = v_851 | ~v_623;
assign x_9524 = v_851 | ~v_624;
assign x_9525 = v_851 | ~v_721;
assign x_9526 = v_851 | ~v_126;
assign x_9527 = v_851 | ~v_110;
assign x_9528 = v_851 | ~v_102;
assign x_9529 = v_851 | ~v_100;
assign x_9530 = v_851 | ~v_51;
assign x_9531 = v_851 | ~v_50;
assign x_9532 = v_851 | ~v_48;
assign x_9533 = v_851 | ~v_46;
assign x_9534 = v_851 | ~v_45;
assign x_9535 = ~v_66 | ~v_124 | v_850;
assign x_9536 = ~v_58 | v_124 | v_849;
assign x_9537 = ~v_14 | ~v_123 | v_848;
assign x_9538 = ~v_12 | v_123 | v_847;
assign x_9539 = v_846 | ~v_588;
assign x_9540 = v_846 | ~v_589;
assign x_9541 = v_846 | ~v_842;
assign x_9542 = v_846 | ~v_843;
assign x_9543 = v_846 | ~v_705;
assign x_9544 = v_846 | ~v_706;
assign x_9545 = v_846 | ~v_596;
assign x_9546 = v_846 | ~v_597;
assign x_9547 = v_846 | ~v_844;
assign x_9548 = v_846 | ~v_845;
assign x_9549 = v_846 | ~v_600;
assign x_9550 = v_846 | ~v_601;
assign x_9551 = v_846 | ~v_707;
assign x_9552 = v_846 | ~v_708;
assign x_9553 = v_846 | ~v_709;
assign x_9554 = v_846 | ~v_710;
assign x_9555 = v_846 | ~v_604;
assign x_9556 = v_846 | ~v_605;
assign x_9557 = v_846 | ~v_122;
assign x_9558 = v_846 | ~v_108;
assign x_9559 = v_846 | ~v_95;
assign x_9560 = v_846 | ~v_93;
assign x_9561 = v_846 | ~v_25;
assign x_9562 = v_846 | ~v_24;
assign x_9563 = v_846 | ~v_22;
assign x_9564 = v_846 | ~v_20;
assign x_9565 = v_846 | ~v_19;
assign x_9566 = ~v_41 | ~v_124 | v_845;
assign x_9567 = ~v_33 | v_124 | v_844;
assign x_9568 = ~v_15 | ~v_123 | v_843;
assign x_9569 = ~v_11 | v_123 | v_842;
assign x_9570 = v_841 | ~v_840;
assign x_9571 = v_841 | ~v_787;
assign x_9572 = v_841 | ~v_698;
assign x_9573 = v_841 | ~v_699;
assign x_9574 = v_841 | ~v_700;
assign x_9575 = v_841 | ~v_701;
assign x_9576 = ~v_839 | ~v_834 | ~v_829 | v_840;
assign x_9577 = v_839 | ~v_835;
assign x_9578 = v_839 | ~v_836;
assign x_9579 = v_839 | ~v_814;
assign x_9580 = v_839 | ~v_815;
assign x_9581 = v_839 | ~v_837;
assign x_9582 = v_839 | ~v_838;
assign x_9583 = v_839 | ~v_726;
assign x_9584 = v_839 | ~v_818;
assign x_9585 = v_839 | ~v_819;
assign x_9586 = v_839 | ~v_729;
assign x_9587 = v_839 | ~v_730;
assign x_9588 = v_839 | ~v_731;
assign x_9589 = v_839 | ~v_732;
assign x_9590 = v_839 | ~v_733;
assign x_9591 = v_839 | ~v_820;
assign x_9592 = v_839 | ~v_642;
assign x_9593 = v_839 | ~v_643;
assign x_9594 = v_839 | ~v_821;
assign x_9595 = v_839 | ~v_112;
assign x_9596 = v_839 | ~v_106;
assign x_9597 = v_839 | ~v_105;
assign x_9598 = v_839 | ~v_104;
assign x_9599 = v_839 | ~v_76;
assign x_9600 = v_839 | ~v_75;
assign x_9601 = v_839 | ~v_74;
assign x_9602 = v_839 | ~v_73;
assign x_9603 = v_839 | ~v_71;
assign x_9604 = ~v_16 | ~v_114 | v_838;
assign x_9605 = ~v_13 | v_114 | v_837;
assign x_9606 = ~v_91 | ~v_115 | v_836;
assign x_9607 = ~v_83 | v_115 | v_835;
assign x_9608 = v_834 | ~v_830;
assign x_9609 = v_834 | ~v_831;
assign x_9610 = v_834 | ~v_803;
assign x_9611 = v_834 | ~v_804;
assign x_9612 = v_834 | ~v_714;
assign x_9613 = v_834 | ~v_807;
assign x_9614 = v_834 | ~v_808;
assign x_9615 = v_834 | ~v_716;
assign x_9616 = v_834 | ~v_717;
assign x_9617 = v_834 | ~v_832;
assign x_9618 = v_834 | ~v_833;
assign x_9619 = v_834 | ~v_719;
assign x_9620 = v_834 | ~v_720;
assign x_9621 = v_834 | ~v_809;
assign x_9622 = v_834 | ~v_810;
assign x_9623 = v_834 | ~v_623;
assign x_9624 = v_834 | ~v_624;
assign x_9625 = v_834 | ~v_721;
assign x_9626 = v_834 | ~v_110;
assign x_9627 = v_834 | ~v_102;
assign x_9628 = v_834 | ~v_101;
assign x_9629 = v_834 | ~v_100;
assign x_9630 = v_834 | ~v_51;
assign x_9631 = v_834 | ~v_50;
assign x_9632 = v_834 | ~v_49;
assign x_9633 = v_834 | ~v_48;
assign x_9634 = v_834 | ~v_46;
assign x_9635 = ~v_12 | v_114 | v_833;
assign x_9636 = ~v_14 | ~v_114 | v_832;
assign x_9637 = ~v_66 | ~v_115 | v_831;
assign x_9638 = ~v_58 | v_115 | v_830;
assign x_9639 = v_829 | ~v_825;
assign x_9640 = v_829 | ~v_826;
assign x_9641 = v_829 | ~v_792;
assign x_9642 = v_829 | ~v_793;
assign x_9643 = v_829 | ~v_705;
assign x_9644 = v_829 | ~v_706;
assign x_9645 = v_829 | ~v_796;
assign x_9646 = v_829 | ~v_797;
assign x_9647 = v_829 | ~v_707;
assign x_9648 = v_829 | ~v_708;
assign x_9649 = v_829 | ~v_827;
assign x_9650 = v_829 | ~v_709;
assign x_9651 = v_829 | ~v_710;
assign x_9652 = v_829 | ~v_798;
assign x_9653 = v_829 | ~v_799;
assign x_9654 = v_829 | ~v_604;
assign x_9655 = v_829 | ~v_605;
assign x_9656 = v_829 | ~v_828;
assign x_9657 = v_829 | ~v_108;
assign x_9658 = v_829 | ~v_95;
assign x_9659 = v_829 | ~v_94;
assign x_9660 = v_829 | ~v_93;
assign x_9661 = v_829 | ~v_25;
assign x_9662 = v_829 | ~v_24;
assign x_9663 = v_829 | ~v_23;
assign x_9664 = v_829 | ~v_22;
assign x_9665 = v_829 | ~v_20;
assign x_9666 = ~v_11 | v_114 | v_828;
assign x_9667 = ~v_15 | ~v_114 | v_827;
assign x_9668 = ~v_41 | ~v_115 | v_826;
assign x_9669 = ~v_33 | v_115 | v_825;
assign x_9670 = v_824 | ~v_789;
assign x_9671 = v_824 | ~v_823;
assign x_9672 = v_824 | ~v_698;
assign x_9673 = v_824 | ~v_699;
assign x_9674 = v_824 | ~v_700;
assign x_9675 = v_824 | ~v_701;
assign x_9676 = ~v_822 | ~v_811 | ~v_800 | v_823;
assign x_9677 = v_822 | ~v_812;
assign x_9678 = v_822 | ~v_813;
assign x_9679 = v_822 | ~v_814;
assign x_9680 = v_822 | ~v_815;
assign x_9681 = v_822 | ~v_816;
assign x_9682 = v_822 | ~v_817;
assign x_9683 = v_822 | ~v_818;
assign x_9684 = v_822 | ~v_819;
assign x_9685 = v_822 | ~v_688;
assign x_9686 = v_822 | ~v_689;
assign x_9687 = v_822 | ~v_690;
assign x_9688 = v_822 | ~v_691;
assign x_9689 = v_822 | ~v_820;
assign x_9690 = v_822 | ~v_694;
assign x_9691 = v_822 | ~v_695;
assign x_9692 = v_822 | ~v_642;
assign x_9693 = v_822 | ~v_643;
assign x_9694 = v_822 | ~v_821;
assign x_9695 = v_822 | ~v_132;
assign x_9696 = v_822 | ~v_121;
assign x_9697 = v_822 | ~v_113;
assign x_9698 = v_822 | ~v_106;
assign x_9699 = v_822 | ~v_105;
assign x_9700 = v_822 | ~v_104;
assign x_9701 = v_822 | ~v_75;
assign x_9702 = v_822 | ~v_74;
assign x_9703 = v_822 | ~v_68;
assign x_9704 = ~v_87 | ~v_134 | v_821;
assign x_9705 = ~v_79 | v_134 | v_820;
assign x_9706 = ~v_90 | ~v_133 | v_819;
assign x_9707 = ~v_82 | v_133 | v_818;
assign x_9708 = ~v_91 | ~v_133 | v_817;
assign x_9709 = ~v_83 | v_133 | v_816;
assign x_9710 = ~v_92 | ~v_116 | v_815;
assign x_9711 = ~v_84 | v_116 | v_814;
assign x_9712 = ~v_16 | ~v_134 | v_813;
assign x_9713 = ~v_13 | v_134 | v_812;
assign x_9714 = v_811 | ~v_801;
assign x_9715 = v_811 | ~v_802;
assign x_9716 = v_811 | ~v_803;
assign x_9717 = v_811 | ~v_804;
assign x_9718 = v_811 | ~v_805;
assign x_9719 = v_811 | ~v_806;
assign x_9720 = v_811 | ~v_807;
assign x_9721 = v_811 | ~v_808;
assign x_9722 = v_811 | ~v_669;
assign x_9723 = v_811 | ~v_670;
assign x_9724 = v_811 | ~v_671;
assign x_9725 = v_811 | ~v_672;
assign x_9726 = v_811 | ~v_809;
assign x_9727 = v_811 | ~v_810;
assign x_9728 = v_811 | ~v_675;
assign x_9729 = v_811 | ~v_676;
assign x_9730 = v_811 | ~v_623;
assign x_9731 = v_811 | ~v_624;
assign x_9732 = v_811 | ~v_131;
assign x_9733 = v_811 | ~v_120;
assign x_9734 = v_811 | ~v_111;
assign x_9735 = v_811 | ~v_102;
assign x_9736 = v_811 | ~v_101;
assign x_9737 = v_811 | ~v_100;
assign x_9738 = v_811 | ~v_50;
assign x_9739 = v_811 | ~v_49;
assign x_9740 = v_811 | ~v_43;
assign x_9741 = ~v_62 | ~v_134 | v_810;
assign x_9742 = ~v_54 | v_134 | v_809;
assign x_9743 = ~v_65 | ~v_133 | v_808;
assign x_9744 = ~v_57 | v_133 | v_807;
assign x_9745 = ~v_66 | ~v_133 | v_806;
assign x_9746 = ~v_58 | v_133 | v_805;
assign x_9747 = ~v_67 | ~v_116 | v_804;
assign x_9748 = ~v_59 | v_116 | v_803;
assign x_9749 = ~v_14 | ~v_134 | v_802;
assign x_9750 = ~v_12 | v_134 | v_801;
assign x_9751 = v_800 | ~v_790;
assign x_9752 = v_800 | ~v_791;
assign x_9753 = v_800 | ~v_792;
assign x_9754 = v_800 | ~v_793;
assign x_9755 = v_800 | ~v_794;
assign x_9756 = v_800 | ~v_795;
assign x_9757 = v_800 | ~v_796;
assign x_9758 = v_800 | ~v_797;
assign x_9759 = v_800 | ~v_653;
assign x_9760 = v_800 | ~v_654;
assign x_9761 = v_800 | ~v_655;
assign x_9762 = v_800 | ~v_656;
assign x_9763 = v_800 | ~v_798;
assign x_9764 = v_800 | ~v_799;
assign x_9765 = v_800 | ~v_659;
assign x_9766 = v_800 | ~v_660;
assign x_9767 = v_800 | ~v_604;
assign x_9768 = v_800 | ~v_605;
assign x_9769 = v_800 | ~v_128;
assign x_9770 = v_800 | ~v_117;
assign x_9771 = v_800 | ~v_109;
assign x_9772 = v_800 | ~v_95;
assign x_9773 = v_800 | ~v_94;
assign x_9774 = v_800 | ~v_93;
assign x_9775 = v_800 | ~v_24;
assign x_9776 = v_800 | ~v_23;
assign x_9777 = v_800 | ~v_17;
assign x_9778 = ~v_37 | ~v_134 | v_799;
assign x_9779 = ~v_29 | v_134 | v_798;
assign x_9780 = ~v_40 | ~v_133 | v_797;
assign x_9781 = ~v_32 | v_133 | v_796;
assign x_9782 = ~v_41 | ~v_133 | v_795;
assign x_9783 = ~v_33 | v_133 | v_794;
assign x_9784 = ~v_42 | ~v_116 | v_793;
assign x_9785 = ~v_34 | v_116 | v_792;
assign x_9786 = ~v_15 | ~v_134 | v_791;
assign x_9787 = ~v_11 | v_134 | v_790;
assign x_9788 = ~v_788 | ~v_771 | ~v_702 | v_789;
assign x_9789 = v_788 | ~v_787;
assign x_9790 = v_788 | ~v_698;
assign x_9791 = v_788 | ~v_699;
assign x_9792 = v_788 | ~v_700;
assign x_9793 = v_788 | ~v_701;
assign x_9794 = ~v_786 | ~v_781 | ~v_776 | v_787;
assign x_9795 = v_786 | ~v_628;
assign x_9796 = v_786 | ~v_629;
assign x_9797 = v_786 | ~v_782;
assign x_9798 = v_786 | ~v_783;
assign x_9799 = v_786 | ~v_682;
assign x_9800 = v_786 | ~v_683;
assign x_9801 = v_786 | ~v_684;
assign x_9802 = v_786 | ~v_685;
assign x_9803 = v_786 | ~v_632;
assign x_9804 = v_786 | ~v_633;
assign x_9805 = v_786 | ~v_784;
assign x_9806 = v_786 | ~v_785;
assign x_9807 = v_786 | ~v_640;
assign x_9808 = v_786 | ~v_641;
assign x_9809 = v_786 | ~v_692;
assign x_9810 = v_786 | ~v_693;
assign x_9811 = v_786 | ~v_642;
assign x_9812 = v_786 | ~v_643;
assign x_9813 = v_786 | ~v_121;
assign x_9814 = v_786 | ~v_113;
assign x_9815 = v_786 | ~v_112;
assign x_9816 = v_786 | ~v_106;
assign x_9817 = v_786 | ~v_105;
assign x_9818 = v_786 | ~v_104;
assign x_9819 = v_786 | ~v_75;
assign x_9820 = v_786 | ~v_74;
assign x_9821 = v_786 | ~v_73;
assign x_9822 = ~v_91 | ~v_119 | v_785;
assign x_9823 = ~v_83 | v_119 | v_784;
assign x_9824 = ~v_16 | ~v_118 | v_783;
assign x_9825 = ~v_13 | v_118 | v_782;
assign x_9826 = v_781 | ~v_609;
assign x_9827 = v_781 | ~v_610;
assign x_9828 = v_781 | ~v_777;
assign x_9829 = v_781 | ~v_778;
assign x_9830 = v_781 | ~v_663;
assign x_9831 = v_781 | ~v_664;
assign x_9832 = v_781 | ~v_613;
assign x_9833 = v_781 | ~v_614;
assign x_9834 = v_781 | ~v_779;
assign x_9835 = v_781 | ~v_780;
assign x_9836 = v_781 | ~v_621;
assign x_9837 = v_781 | ~v_622;
assign x_9838 = v_781 | ~v_673;
assign x_9839 = v_781 | ~v_674;
assign x_9840 = v_781 | ~v_623;
assign x_9841 = v_781 | ~v_624;
assign x_9842 = v_781 | ~v_677;
assign x_9843 = v_781 | ~v_678;
assign x_9844 = v_781 | ~v_120;
assign x_9845 = v_781 | ~v_111;
assign x_9846 = v_781 | ~v_110;
assign x_9847 = v_781 | ~v_102;
assign x_9848 = v_781 | ~v_101;
assign x_9849 = v_781 | ~v_100;
assign x_9850 = v_781 | ~v_50;
assign x_9851 = v_781 | ~v_49;
assign x_9852 = v_781 | ~v_48;
assign x_9853 = ~v_66 | ~v_119 | v_780;
assign x_9854 = ~v_58 | v_119 | v_779;
assign x_9855 = ~v_14 | ~v_118 | v_778;
assign x_9856 = ~v_12 | v_118 | v_777;
assign x_9857 = v_776 | ~v_590;
assign x_9858 = v_776 | ~v_591;
assign x_9859 = v_776 | ~v_772;
assign x_9860 = v_776 | ~v_773;
assign x_9861 = v_776 | ~v_646;
assign x_9862 = v_776 | ~v_647;
assign x_9863 = v_776 | ~v_648;
assign x_9864 = v_776 | ~v_594;
assign x_9865 = v_776 | ~v_595;
assign x_9866 = v_776 | ~v_774;
assign x_9867 = v_776 | ~v_775;
assign x_9868 = v_776 | ~v_602;
assign x_9869 = v_776 | ~v_603;
assign x_9870 = v_776 | ~v_657;
assign x_9871 = v_776 | ~v_658;
assign x_9872 = v_776 | ~v_604;
assign x_9873 = v_776 | ~v_605;
assign x_9874 = v_776 | ~v_661;
assign x_9875 = v_776 | ~v_117;
assign x_9876 = v_776 | ~v_109;
assign x_9877 = v_776 | ~v_108;
assign x_9878 = v_776 | ~v_95;
assign x_9879 = v_776 | ~v_94;
assign x_9880 = v_776 | ~v_93;
assign x_9881 = v_776 | ~v_24;
assign x_9882 = v_776 | ~v_23;
assign x_9883 = v_776 | ~v_22;
assign x_9884 = ~v_41 | ~v_119 | v_775;
assign x_9885 = ~v_33 | v_119 | v_774;
assign x_9886 = ~v_15 | ~v_118 | v_773;
assign x_9887 = ~v_11 | v_118 | v_772;
assign x_9888 = v_771 | ~v_736;
assign x_9889 = v_771 | ~v_770;
assign x_9890 = v_771 | ~v_698;
assign x_9891 = v_771 | ~v_699;
assign x_9892 = v_771 | ~v_700;
assign x_9893 = v_771 | ~v_701;
assign x_9894 = ~v_769 | ~v_758 | ~v_747 | v_770;
assign x_9895 = v_769 | ~v_628;
assign x_9896 = v_769 | ~v_629;
assign x_9897 = v_769 | ~v_759;
assign x_9898 = v_769 | ~v_760;
assign x_9899 = v_769 | ~v_761;
assign x_9900 = v_769 | ~v_762;
assign x_9901 = v_769 | ~v_763;
assign x_9902 = v_769 | ~v_764;
assign x_9903 = v_769 | ~v_765;
assign x_9904 = v_769 | ~v_766;
assign x_9905 = v_769 | ~v_632;
assign x_9906 = v_769 | ~v_633;
assign x_9907 = v_769 | ~v_640;
assign x_9908 = v_769 | ~v_641;
assign x_9909 = v_769 | ~v_767;
assign x_9910 = v_769 | ~v_768;
assign x_9911 = v_769 | ~v_642;
assign x_9912 = v_769 | ~v_643;
assign x_9913 = v_769 | ~v_113;
assign x_9914 = v_769 | ~v_112;
assign x_9915 = v_769 | ~v_105;
assign x_9916 = v_769 | ~v_104;
assign x_9917 = v_769 | ~v_76;
assign x_9918 = v_769 | ~v_75;
assign x_9919 = v_769 | ~v_74;
assign x_9920 = v_769 | ~v_73;
assign x_9921 = v_769 | ~v_72;
assign x_9922 = ~v_87 | ~v_124 | v_768;
assign x_9923 = ~v_79 | v_124 | v_767;
assign x_9924 = ~v_91 | ~v_114 | v_766;
assign x_9925 = ~v_83 | v_114 | v_765;
assign x_9926 = ~v_26 | ~v_92 | v_764;
assign x_9927 = v_26 | ~v_84 | v_763;
assign x_9928 = ~v_16 | ~v_115 | v_762;
assign x_9929 = ~v_13 | v_115 | v_761;
assign x_9930 = ~v_90 | ~v_123 | v_760;
assign x_9931 = ~v_82 | v_123 | v_759;
assign x_9932 = v_758 | ~v_609;
assign x_9933 = v_758 | ~v_610;
assign x_9934 = v_758 | ~v_748;
assign x_9935 = v_758 | ~v_749;
assign x_9936 = v_758 | ~v_750;
assign x_9937 = v_758 | ~v_751;
assign x_9938 = v_758 | ~v_752;
assign x_9939 = v_758 | ~v_613;
assign x_9940 = v_758 | ~v_614;
assign x_9941 = v_758 | ~v_753;
assign x_9942 = v_758 | ~v_754;
assign x_9943 = v_758 | ~v_621;
assign x_9944 = v_758 | ~v_622;
assign x_9945 = v_758 | ~v_755;
assign x_9946 = v_758 | ~v_756;
assign x_9947 = v_758 | ~v_623;
assign x_9948 = v_758 | ~v_624;
assign x_9949 = v_758 | ~v_757;
assign x_9950 = v_758 | ~v_111;
assign x_9951 = v_758 | ~v_110;
assign x_9952 = v_758 | ~v_101;
assign x_9953 = v_758 | ~v_100;
assign x_9954 = v_758 | ~v_51;
assign x_9955 = v_758 | ~v_50;
assign x_9956 = v_758 | ~v_49;
assign x_9957 = v_758 | ~v_48;
assign x_9958 = v_758 | ~v_47;
assign x_9959 = ~v_26 | ~v_67 | v_757;
assign x_9960 = ~v_62 | ~v_124 | v_756;
assign x_9961 = ~v_54 | v_124 | v_755;
assign x_9962 = ~v_12 | v_115 | v_754;
assign x_9963 = ~v_14 | ~v_115 | v_753;
assign x_9964 = ~v_66 | ~v_114 | v_752;
assign x_9965 = ~v_58 | v_114 | v_751;
assign x_9966 = v_26 | ~v_59 | v_750;
assign x_9967 = ~v_65 | ~v_123 | v_749;
assign x_9968 = ~v_57 | v_123 | v_748;
assign x_9969 = v_747 | ~v_590;
assign x_9970 = v_747 | ~v_591;
assign x_9971 = v_747 | ~v_737;
assign x_9972 = v_747 | ~v_738;
assign x_9973 = v_747 | ~v_739;
assign x_9974 = v_747 | ~v_740;
assign x_9975 = v_747 | ~v_741;
assign x_9976 = v_747 | ~v_594;
assign x_9977 = v_747 | ~v_595;
assign x_9978 = v_747 | ~v_742;
assign x_9979 = v_747 | ~v_743;
assign x_9980 = v_747 | ~v_602;
assign x_9981 = v_747 | ~v_603;
assign x_9982 = v_747 | ~v_744;
assign x_9983 = v_747 | ~v_745;
assign x_9984 = v_747 | ~v_604;
assign x_9985 = v_747 | ~v_605;
assign x_9986 = v_747 | ~v_746;
assign x_9987 = v_747 | ~v_109;
assign x_9988 = v_747 | ~v_108;
assign x_9989 = v_747 | ~v_94;
assign x_9990 = v_747 | ~v_93;
assign x_9991 = v_747 | ~v_25;
assign x_9992 = v_747 | ~v_24;
assign x_9993 = v_747 | ~v_23;
assign x_9994 = v_747 | ~v_22;
assign x_9995 = v_747 | ~v_21;
assign x_9996 = ~v_26 | ~v_42 | v_746;
assign x_9997 = ~v_37 | ~v_124 | v_745;
assign x_9998 = ~v_29 | v_124 | v_744;
assign x_9999 = ~v_15 | ~v_115 | v_743;
assign x_10000 = ~v_11 | v_115 | v_742;
assign x_10001 = ~v_41 | ~v_114 | v_741;
assign x_10002 = ~v_33 | v_114 | v_740;
assign x_10003 = ~v_34 | v_26 | v_739;
assign x_10004 = ~v_40 | ~v_123 | v_738;
assign x_10005 = ~v_32 | v_123 | v_737;
assign x_10006 = ~v_735 | ~v_724 | ~v_713 | v_736;
assign x_10007 = v_735 | ~v_682;
assign x_10008 = v_735 | ~v_683;
assign x_10009 = v_735 | ~v_725;
assign x_10010 = v_735 | ~v_726;
assign x_10011 = v_735 | ~v_727;
assign x_10012 = v_735 | ~v_728;
assign x_10013 = v_735 | ~v_684;
assign x_10014 = v_735 | ~v_685;
assign x_10015 = v_735 | ~v_729;
assign x_10016 = v_735 | ~v_730;
assign x_10017 = v_735 | ~v_731;
assign x_10018 = v_735 | ~v_732;
assign x_10019 = v_735 | ~v_733;
assign x_10020 = v_735 | ~v_692;
assign x_10021 = v_735 | ~v_693;
assign x_10022 = v_735 | ~v_642;
assign x_10023 = v_735 | ~v_643;
assign x_10024 = v_735 | ~v_734;
assign x_10025 = v_735 | ~v_112;
assign x_10026 = v_735 | ~v_107;
assign x_10027 = v_735 | ~v_106;
assign x_10028 = v_735 | ~v_105;
assign x_10029 = v_735 | ~v_104;
assign x_10030 = v_735 | ~v_76;
assign x_10031 = v_735 | ~v_74;
assign x_10032 = v_735 | ~v_73;
assign x_10033 = v_735 | ~v_71;
assign x_10034 = ~v_13 | v_97 | v_734;
assign x_10035 = ~v_86 | ~v_124 | v_733;
assign x_10036 = ~v_78 | v_124 | v_732;
assign x_10037 = ~v_26 | ~v_89 | v_731;
assign x_10038 = ~v_88 | ~v_123 | v_730;
assign x_10039 = ~v_80 | v_123 | v_729;
assign x_10040 = ~v_91 | ~v_98 | v_728;
assign x_10041 = ~v_83 | v_98 | v_727;
assign x_10042 = v_26 | ~v_81 | v_726;
assign x_10043 = ~v_16 | ~v_97 | v_725;
assign x_10044 = v_724 | ~v_714;
assign x_10045 = v_724 | ~v_715;
assign x_10046 = v_724 | ~v_663;
assign x_10047 = v_724 | ~v_664;
assign x_10048 = v_724 | ~v_716;
assign x_10049 = v_724 | ~v_717;
assign x_10050 = v_724 | ~v_718;
assign x_10051 = v_724 | ~v_719;
assign x_10052 = v_724 | ~v_720;
assign x_10053 = v_724 | ~v_673;
assign x_10054 = v_724 | ~v_674;
assign x_10055 = v_724 | ~v_623;
assign x_10056 = v_724 | ~v_624;
assign x_10057 = v_724 | ~v_721;
assign x_10058 = v_724 | ~v_677;
assign x_10059 = v_724 | ~v_722;
assign x_10060 = v_724 | ~v_678;
assign x_10061 = v_724 | ~v_723;
assign x_10062 = v_724 | ~v_110;
assign x_10063 = v_724 | ~v_103;
assign x_10064 = v_724 | ~v_102;
assign x_10065 = v_724 | ~v_101;
assign x_10066 = v_724 | ~v_100;
assign x_10067 = v_724 | ~v_51;
assign x_10068 = v_724 | ~v_49;
assign x_10069 = v_724 | ~v_48;
assign x_10070 = v_724 | ~v_46;
assign x_10071 = ~v_12 | v_97 | v_723;
assign x_10072 = ~v_58 | v_98 | v_722;
assign x_10073 = ~v_26 | ~v_64 | v_721;
assign x_10074 = ~v_61 | ~v_124 | v_720;
assign x_10075 = ~v_53 | v_124 | v_719;
assign x_10076 = ~v_14 | ~v_97 | v_718;
assign x_10077 = ~v_63 | ~v_123 | v_717;
assign x_10078 = ~v_55 | v_123 | v_716;
assign x_10079 = ~v_66 | ~v_98 | v_715;
assign x_10080 = v_26 | ~v_56 | v_714;
assign x_10081 = v_713 | ~v_646;
assign x_10082 = v_713 | ~v_703;
assign x_10083 = v_713 | ~v_704;
assign x_10084 = v_713 | ~v_705;
assign x_10085 = v_713 | ~v_706;
assign x_10086 = v_713 | ~v_647;
assign x_10087 = v_713 | ~v_648;
assign x_10088 = v_713 | ~v_707;
assign x_10089 = v_713 | ~v_708;
assign x_10090 = v_713 | ~v_709;
assign x_10091 = v_713 | ~v_710;
assign x_10092 = v_713 | ~v_657;
assign x_10093 = v_713 | ~v_658;
assign x_10094 = v_713 | ~v_604;
assign x_10095 = v_713 | ~v_605;
assign x_10096 = v_713 | ~v_661;
assign x_10097 = v_713 | ~v_711;
assign x_10098 = v_713 | ~v_712;
assign x_10099 = v_713 | ~v_108;
assign x_10100 = v_713 | ~v_96;
assign x_10101 = v_713 | ~v_95;
assign x_10102 = v_713 | ~v_94;
assign x_10103 = v_713 | ~v_93;
assign x_10104 = v_713 | ~v_25;
assign x_10105 = v_713 | ~v_23;
assign x_10106 = v_713 | ~v_22;
assign x_10107 = v_713 | ~v_20;
assign x_10108 = ~v_41 | ~v_98 | v_712;
assign x_10109 = ~v_33 | v_98 | v_711;
assign x_10110 = ~v_36 | ~v_124 | v_710;
assign x_10111 = ~v_28 | v_124 | v_709;
assign x_10112 = ~v_38 | ~v_123 | v_708;
assign x_10113 = ~v_30 | v_123 | v_707;
assign x_10114 = ~v_26 | ~v_39 | v_706;
assign x_10115 = ~v_31 | v_26 | v_705;
assign x_10116 = ~v_15 | ~v_97 | v_704;
assign x_10117 = ~v_11 | v_97 | v_703;
assign x_10118 = v_702 | ~v_645;
assign x_10119 = v_702 | ~v_697;
assign x_10120 = v_702 | ~v_698;
assign x_10121 = v_702 | ~v_699;
assign x_10122 = v_702 | ~v_700;
assign x_10123 = v_702 | ~v_701;
assign x_10124 = ~v_12 | v_11 | v_701;
assign x_10125 = ~v_13 | v_12 | v_700;
assign x_10126 = ~v_15 | v_14 | v_699;
assign x_10127 = ~v_14 | v_16 | v_698;
assign x_10128 = ~v_696 | ~v_679 | ~v_662 | v_697;
assign x_10129 = v_696 | ~v_680;
assign x_10130 = v_696 | ~v_681;
assign x_10131 = v_696 | ~v_682;
assign x_10132 = v_696 | ~v_683;
assign x_10133 = v_696 | ~v_684;
assign x_10134 = v_696 | ~v_685;
assign x_10135 = v_696 | ~v_686;
assign x_10136 = v_696 | ~v_687;
assign x_10137 = v_696 | ~v_688;
assign x_10138 = v_696 | ~v_689;
assign x_10139 = v_696 | ~v_690;
assign x_10140 = v_696 | ~v_691;
assign x_10141 = v_696 | ~v_692;
assign x_10142 = v_696 | ~v_693;
assign x_10143 = v_696 | ~v_694;
assign x_10144 = v_696 | ~v_695;
assign x_10145 = v_696 | ~v_642;
assign x_10146 = v_696 | ~v_643;
assign x_10147 = v_696 | ~v_132;
assign x_10148 = v_696 | ~v_113;
assign x_10149 = v_696 | ~v_106;
assign x_10150 = v_696 | ~v_105;
assign x_10151 = v_696 | ~v_104;
assign x_10152 = v_696 | ~v_76;
assign x_10153 = v_696 | ~v_75;
assign x_10154 = v_696 | ~v_74;
assign x_10155 = v_696 | ~v_68;
assign x_10156 = ~v_88 | ~v_125 | v_695;
assign x_10157 = ~v_80 | v_125 | v_694;
assign x_10158 = ~v_87 | ~v_129 | v_693;
assign x_10159 = ~v_79 | v_129 | v_692;
assign x_10160 = ~v_86 | ~v_125 | v_691;
assign x_10161 = ~v_78 | v_125 | v_690;
assign x_10162 = ~v_89 | ~v_125 | v_689;
assign x_10163 = ~v_81 | v_125 | v_688;
assign x_10164 = ~v_91 | ~v_130 | v_687;
assign x_10165 = ~v_83 | v_130 | v_686;
assign x_10166 = ~v_90 | ~v_130 | v_685;
assign x_10167 = ~v_82 | v_130 | v_684;
assign x_10168 = ~v_92 | ~v_99 | v_683;
assign x_10169 = ~v_84 | v_99 | v_682;
assign x_10170 = ~v_16 | ~v_129 | v_681;
assign x_10171 = ~v_13 | v_129 | v_680;
assign x_10172 = v_679 | ~v_663;
assign x_10173 = v_679 | ~v_664;
assign x_10174 = v_679 | ~v_665;
assign x_10175 = v_679 | ~v_666;
assign x_10176 = v_679 | ~v_667;
assign x_10177 = v_679 | ~v_668;
assign x_10178 = v_679 | ~v_669;
assign x_10179 = v_679 | ~v_670;
assign x_10180 = v_679 | ~v_671;
assign x_10181 = v_679 | ~v_672;
assign x_10182 = v_679 | ~v_673;
assign x_10183 = v_679 | ~v_674;
assign x_10184 = v_679 | ~v_675;
assign x_10185 = v_679 | ~v_676;
assign x_10186 = v_679 | ~v_623;
assign x_10187 = v_679 | ~v_624;
assign x_10188 = v_679 | ~v_677;
assign x_10189 = v_679 | ~v_678;
assign x_10190 = v_679 | ~v_131;
assign x_10191 = v_679 | ~v_111;
assign x_10192 = v_679 | ~v_102;
assign x_10193 = v_679 | ~v_101;
assign x_10194 = v_679 | ~v_100;
assign x_10195 = v_679 | ~v_51;
assign x_10196 = v_679 | ~v_50;
assign x_10197 = v_679 | ~v_49;
assign x_10198 = v_679 | ~v_43;
assign x_10199 = ~v_67 | ~v_99 | v_678;
assign x_10200 = ~v_59 | v_99 | v_677;
assign x_10201 = ~v_63 | ~v_125 | v_676;
assign x_10202 = ~v_55 | v_125 | v_675;
assign x_10203 = ~v_62 | ~v_129 | v_674;
assign x_10204 = ~v_54 | v_129 | v_673;
assign x_10205 = ~v_61 | ~v_125 | v_672;
assign x_10206 = ~v_53 | v_125 | v_671;
assign x_10207 = ~v_64 | ~v_125 | v_670;
assign x_10208 = ~v_56 | v_125 | v_669;
assign x_10209 = ~v_12 | v_129 | v_668;
assign x_10210 = ~v_14 | ~v_129 | v_667;
assign x_10211 = ~v_66 | ~v_130 | v_666;
assign x_10212 = ~v_58 | v_130 | v_665;
assign x_10213 = ~v_65 | ~v_130 | v_664;
assign x_10214 = ~v_57 | v_130 | v_663;
assign x_10215 = v_662 | ~v_646;
assign x_10216 = v_662 | ~v_647;
assign x_10217 = v_662 | ~v_648;
assign x_10218 = v_662 | ~v_649;
assign x_10219 = v_662 | ~v_650;
assign x_10220 = v_662 | ~v_651;
assign x_10221 = v_662 | ~v_652;
assign x_10222 = v_662 | ~v_653;
assign x_10223 = v_662 | ~v_654;
assign x_10224 = v_662 | ~v_655;
assign x_10225 = v_662 | ~v_656;
assign x_10226 = v_662 | ~v_657;
assign x_10227 = v_662 | ~v_658;
assign x_10228 = v_662 | ~v_659;
assign x_10229 = v_662 | ~v_660;
assign x_10230 = v_662 | ~v_604;
assign x_10231 = v_662 | ~v_605;
assign x_10232 = v_662 | ~v_661;
assign x_10233 = v_662 | ~v_128;
assign x_10234 = v_662 | ~v_109;
assign x_10235 = v_662 | ~v_95;
assign x_10236 = v_662 | ~v_94;
assign x_10237 = v_662 | ~v_93;
assign x_10238 = v_662 | ~v_25;
assign x_10239 = v_662 | ~v_24;
assign x_10240 = v_662 | ~v_23;
assign x_10241 = v_662 | ~v_17;
assign x_10242 = ~v_42 | ~v_99 | v_661;
assign x_10243 = ~v_38 | ~v_125 | v_660;
assign x_10244 = ~v_30 | v_125 | v_659;
assign x_10245 = ~v_37 | ~v_129 | v_658;
assign x_10246 = ~v_29 | v_129 | v_657;
assign x_10247 = ~v_36 | ~v_125 | v_656;
assign x_10248 = ~v_28 | v_125 | v_655;
assign x_10249 = ~v_39 | ~v_125 | v_654;
assign x_10250 = ~v_31 | v_125 | v_653;
assign x_10251 = ~v_15 | ~v_129 | v_652;
assign x_10252 = ~v_11 | v_129 | v_651;
assign x_10253 = ~v_41 | ~v_130 | v_650;
assign x_10254 = ~v_33 | v_130 | v_649;
assign x_10255 = ~v_40 | ~v_130 | v_648;
assign x_10256 = ~v_32 | v_130 | v_647;
assign x_10257 = ~v_34 | v_99 | v_646;
assign x_10258 = ~v_644 | ~v_625 | ~v_606 | v_645;
assign x_10259 = v_644 | ~v_626;
assign x_10260 = v_644 | ~v_627;
assign x_10261 = v_644 | ~v_628;
assign x_10262 = v_644 | ~v_629;
assign x_10263 = v_644 | ~v_630;
assign x_10264 = v_644 | ~v_631;
assign x_10265 = v_644 | ~v_632;
assign x_10266 = v_644 | ~v_633;
assign x_10267 = v_644 | ~v_634;
assign x_10268 = v_644 | ~v_635;
assign x_10269 = v_644 | ~v_636;
assign x_10270 = v_644 | ~v_637;
assign x_10271 = v_644 | ~v_638;
assign x_10272 = v_644 | ~v_639;
assign x_10273 = v_644 | ~v_640;
assign x_10274 = v_644 | ~v_641;
assign x_10275 = v_644 | ~v_642;
assign x_10276 = v_644 | ~v_643;
assign x_10277 = v_644 | ~v_127;
assign x_10278 = v_644 | ~v_113;
assign x_10279 = v_644 | ~v_112;
assign x_10280 = v_644 | ~v_107;
assign x_10281 = v_644 | ~v_106;
assign x_10282 = v_644 | ~v_104;
assign x_10283 = v_644 | ~v_76;
assign x_10284 = v_644 | ~v_73;
assign x_10285 = v_644 | ~v_70;
assign x_10286 = ~v_85 | ~v_125 | v_643;
assign x_10287 = ~v_77 | v_125 | v_642;
assign x_10288 = ~v_86 | ~v_134 | v_641;
assign x_10289 = ~v_78 | v_134 | v_640;
assign x_10290 = ~v_90 | ~v_125 | v_639;
assign x_10291 = ~v_82 | v_125 | v_638;
assign x_10292 = ~v_91 | ~v_134 | v_637;
assign x_10293 = ~v_83 | v_134 | v_636;
assign x_10294 = ~v_92 | ~v_125 | v_635;
assign x_10295 = ~v_84 | v_125 | v_634;
assign x_10296 = ~v_89 | ~v_116 | v_633;
assign x_10297 = ~v_81 | v_116 | v_632;
assign x_10298 = ~v_16 | ~v_133 | v_631;
assign x_10299 = ~v_13 | v_133 | v_630;
assign x_10300 = ~v_88 | ~v_133 | v_629;
assign x_10301 = ~v_80 | v_133 | v_628;
assign x_10302 = ~v_87 | ~v_125 | v_627;
assign x_10303 = ~v_79 | v_125 | v_626;
assign x_10304 = v_625 | ~v_607;
assign x_10305 = v_625 | ~v_608;
assign x_10306 = v_625 | ~v_609;
assign x_10307 = v_625 | ~v_610;
assign x_10308 = v_625 | ~v_611;
assign x_10309 = v_625 | ~v_612;
assign x_10310 = v_625 | ~v_613;
assign x_10311 = v_625 | ~v_614;
assign x_10312 = v_625 | ~v_615;
assign x_10313 = v_625 | ~v_616;
assign x_10314 = v_625 | ~v_617;
assign x_10315 = v_625 | ~v_618;
assign x_10316 = v_625 | ~v_619;
assign x_10317 = v_625 | ~v_620;
assign x_10318 = v_625 | ~v_621;
assign x_10319 = v_625 | ~v_622;
assign x_10320 = v_625 | ~v_623;
assign x_10321 = v_625 | ~v_624;
assign x_10322 = v_625 | ~v_126;
assign x_10323 = v_625 | ~v_111;
assign x_10324 = v_625 | ~v_110;
assign x_10325 = v_625 | ~v_103;
assign x_10326 = v_625 | ~v_102;
assign x_10327 = v_625 | ~v_100;
assign x_10328 = v_625 | ~v_51;
assign x_10329 = v_625 | ~v_48;
assign x_10330 = v_625 | ~v_45;
assign x_10331 = ~v_60 | ~v_125 | v_624;
assign x_10332 = ~v_52 | v_125 | v_623;
assign x_10333 = ~v_61 | ~v_134 | v_622;
assign x_10334 = ~v_53 | v_134 | v_621;
assign x_10335 = ~v_65 | ~v_125 | v_620;
assign x_10336 = ~v_57 | v_125 | v_619;
assign x_10337 = ~v_66 | ~v_134 | v_618;
assign x_10338 = ~v_58 | v_134 | v_617;
assign x_10339 = ~v_67 | ~v_125 | v_616;
assign x_10340 = ~v_59 | v_125 | v_615;
assign x_10341 = ~v_64 | ~v_116 | v_614;
assign x_10342 = ~v_56 | v_116 | v_613;
assign x_10343 = ~v_14 | ~v_133 | v_612;
assign x_10344 = ~v_12 | v_133 | v_611;
assign x_10345 = ~v_63 | ~v_133 | v_610;
assign x_10346 = ~v_55 | v_133 | v_609;
assign x_10347 = ~v_62 | ~v_125 | v_608;
assign x_10348 = ~v_54 | v_125 | v_607;
assign x_10349 = v_606 | ~v_588;
assign x_10350 = v_606 | ~v_589;
assign x_10351 = v_606 | ~v_590;
assign x_10352 = v_606 | ~v_591;
assign x_10353 = v_606 | ~v_592;
assign x_10354 = v_606 | ~v_593;
assign x_10355 = v_606 | ~v_594;
assign x_10356 = v_606 | ~v_595;
assign x_10357 = v_606 | ~v_596;
assign x_10358 = v_606 | ~v_597;
assign x_10359 = v_606 | ~v_598;
assign x_10360 = v_606 | ~v_599;
assign x_10361 = v_606 | ~v_600;
assign x_10362 = v_606 | ~v_601;
assign x_10363 = v_606 | ~v_602;
assign x_10364 = v_606 | ~v_603;
assign x_10365 = v_606 | ~v_604;
assign x_10366 = v_606 | ~v_605;
assign x_10367 = v_606 | ~v_122;
assign x_10368 = v_606 | ~v_109;
assign x_10369 = v_606 | ~v_108;
assign x_10370 = v_606 | ~v_96;
assign x_10371 = v_606 | ~v_95;
assign x_10372 = v_606 | ~v_93;
assign x_10373 = v_606 | ~v_25;
assign x_10374 = v_606 | ~v_22;
assign x_10375 = v_606 | ~v_19;
assign x_10376 = ~v_35 | ~v_125 | v_605;
assign x_10377 = ~v_27 | v_125 | v_604;
assign x_10378 = ~v_36 | ~v_134 | v_603;
assign x_10379 = ~v_28 | v_134 | v_602;
assign x_10380 = ~v_40 | ~v_125 | v_601;
assign x_10381 = ~v_32 | v_125 | v_600;
assign x_10382 = ~v_41 | ~v_134 | v_599;
assign x_10383 = ~v_33 | v_134 | v_598;
assign x_10384 = ~v_42 | ~v_125 | v_597;
assign x_10385 = ~v_34 | v_125 | v_596;
assign x_10386 = ~v_39 | ~v_116 | v_595;
assign x_10387 = ~v_31 | v_116 | v_594;
assign x_10388 = ~v_15 | ~v_133 | v_593;
assign x_10389 = ~v_11 | v_133 | v_592;
assign x_10390 = ~v_38 | ~v_133 | v_591;
assign x_10391 = ~v_30 | v_133 | v_590;
assign x_10392 = ~v_37 | ~v_125 | v_589;
assign x_10393 = ~v_29 | v_125 | v_588;
assign x_10394 = ~v_586 | ~v_531 | v_587;
assign x_10395 = v_586 | ~v_554;
assign x_10396 = v_586 | ~v_570;
assign x_10397 = v_586 | ~v_585;
assign x_10398 = v_586 | ~v_125;
assign x_10399 = ~v_584 | ~v_573 | v_585;
assign x_10400 = v_584 | ~v_574;
assign x_10401 = v_584 | ~v_575;
assign x_10402 = v_584 | ~v_579;
assign x_10403 = v_584 | ~v_583;
assign x_10404 = v_584 | ~v_124;
assign x_10405 = ~v_129 | ~v_582 | v_583;
assign x_10406 = v_582 | ~v_580;
assign x_10407 = v_582 | ~v_581;
assign x_10408 = v_582 | ~v_98;
assign x_10409 = ~v_115 | ~v_119 | v_581;
assign x_10410 = ~v_124 | ~v_130 | v_580;
assign x_10411 = ~v_134 | ~v_578 | v_579;
assign x_10412 = v_578 | ~v_576;
assign x_10413 = v_578 | ~v_577;
assign x_10414 = v_578 | ~v_115;
assign x_10415 = ~v_98 | ~v_118 | v_577;
assign x_10416 = ~v_124 | ~v_133 | v_576;
assign x_10417 = ~v_98 | ~v_129 | v_575;
assign x_10418 = ~v_115 | ~v_134 | v_574;
assign x_10419 = v_573 | ~v_571;
assign x_10420 = v_573 | ~v_536;
assign x_10421 = v_573 | ~v_537;
assign x_10422 = v_573 | ~v_572;
assign x_10423 = v_573 | ~v_123;
assign x_10424 = ~v_114 | ~v_556 | v_572;
assign x_10425 = ~v_97 | ~v_534 | v_571;
assign x_10426 = ~v_569 | ~v_558 | v_570;
assign x_10427 = v_569 | ~v_562;
assign x_10428 = v_569 | ~v_566;
assign x_10429 = v_569 | ~v_567;
assign x_10430 = v_569 | ~v_568;
assign x_10431 = v_569 | ~v_129;
assign x_10432 = ~v_97 | ~v_124 | v_568;
assign x_10433 = ~v_118 | ~v_134 | v_567;
assign x_10434 = ~v_134 | ~v_565 | v_566;
assign x_10435 = v_565 | ~v_563;
assign x_10436 = v_565 | ~v_564;
assign x_10437 = v_565 | ~v_118;
assign x_10438 = ~v_97 | ~v_115 | v_564;
assign x_10439 = ~v_129 | ~v_133 | v_563;
assign x_10440 = ~v_124 | ~v_561 | v_562;
assign x_10441 = v_561 | ~v_559;
assign x_10442 = v_561 | ~v_560;
assign x_10443 = v_561 | ~v_97;
assign x_10444 = ~v_114 | ~v_118 | v_560;
assign x_10445 = ~v_123 | ~v_129 | v_559;
assign x_10446 = v_558 | ~v_555;
assign x_10447 = v_558 | ~v_557;
assign x_10448 = v_558 | ~v_532;
assign x_10449 = v_558 | ~v_533;
assign x_10450 = v_558 | ~v_130;
assign x_10451 = ~v_119 | ~v_556 | v_557;
assign x_10452 = v_556 | ~v_540;
assign x_10453 = v_556 | ~v_541;
assign x_10454 = v_556 | ~v_133;
assign x_10455 = ~v_98 | ~v_538 | v_555;
assign x_10456 = ~v_553 | ~v_542 | v_554;
assign x_10457 = v_553 | ~v_546;
assign x_10458 = v_553 | ~v_550;
assign x_10459 = v_553 | ~v_551;
assign x_10460 = v_553 | ~v_552;
assign x_10461 = v_553 | ~v_134;
assign x_10462 = ~v_114 | ~v_124 | v_552;
assign x_10463 = ~v_119 | ~v_129 | v_551;
assign x_10464 = ~v_124 | ~v_549 | v_550;
assign x_10465 = v_549 | ~v_547;
assign x_10466 = v_549 | ~v_548;
assign x_10467 = v_549 | ~v_114;
assign x_10468 = ~v_97 | ~v_119 | v_548;
assign x_10469 = ~v_123 | ~v_134 | v_547;
assign x_10470 = ~v_129 | ~v_545 | v_546;
assign x_10471 = v_545 | ~v_543;
assign x_10472 = v_545 | ~v_544;
assign x_10473 = v_545 | ~v_119;
assign x_10474 = ~v_98 | ~v_114 | v_544;
assign x_10475 = ~v_130 | ~v_134 | v_543;
assign x_10476 = v_542 | ~v_535;
assign x_10477 = v_542 | ~v_539;
assign x_10478 = v_542 | ~v_540;
assign x_10479 = v_542 | ~v_541;
assign x_10480 = v_542 | ~v_133;
assign x_10481 = ~v_115 | ~v_123 | v_541;
assign x_10482 = ~v_118 | ~v_130 | v_540;
assign x_10483 = ~v_115 | ~v_538 | v_539;
assign x_10484 = v_538 | ~v_536;
assign x_10485 = v_538 | ~v_537;
assign x_10486 = v_538 | ~v_123;
assign x_10487 = ~v_97 | ~v_130 | v_537;
assign x_10488 = ~v_114 | ~v_133 | v_536;
assign x_10489 = ~v_118 | ~v_534 | v_535;
assign x_10490 = v_534 | ~v_532;
assign x_10491 = v_534 | ~v_533;
assign x_10492 = v_534 | ~v_130;
assign x_10493 = ~v_98 | ~v_123 | v_533;
assign x_10494 = ~v_119 | ~v_133 | v_532;
assign x_10495 = v_531 | ~v_509;
assign x_10496 = v_531 | ~v_528;
assign x_10497 = v_531 | ~v_529;
assign x_10498 = v_531 | ~v_484;
assign x_10499 = v_531 | ~v_485;
assign x_10500 = v_531 | ~v_530;
assign x_10501 = v_531 | ~v_486;
assign x_10502 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_525 | ~v_244 | v_530;
assign x_10503 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_370 | ~v_466 | v_529;
assign x_10504 = ~v_527 | ~v_523 | v_528;
assign x_10505 = v_527 | ~v_524;
assign x_10506 = v_527 | ~v_526;
assign x_10507 = v_527 | ~v_429;
assign x_10508 = v_527 | ~v_464;
assign x_10509 = v_527 | ~v_465;
assign x_10510 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_525 | ~v_334 | v_526;
assign x_10511 = v_525 | ~v_505;
assign x_10512 = v_525 | ~v_506;
assign x_10513 = v_525 | ~v_507;
assign x_10514 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_487 | ~v_192 | v_524;
assign x_10515 = v_523 | ~v_514;
assign x_10516 = v_523 | ~v_519;
assign x_10517 = v_523 | ~v_520;
assign x_10518 = v_523 | ~v_521;
assign x_10519 = v_523 | ~v_522;
assign x_10520 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_370 | v_522;
assign x_10521 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_482 | ~v_244 | v_521;
assign x_10522 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_423 | ~v_387 | v_520;
assign x_10523 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_244 | ~v_518 | v_519;
assign x_10524 = v_518 | ~v_515;
assign x_10525 = v_518 | ~v_516;
assign x_10526 = v_518 | ~v_517;
assign x_10527 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_482 | v_517;
assign x_10528 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_463 | ~v_387 | v_516;
assign x_10529 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_503 | ~v_370 | v_515;
assign x_10530 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_423 | ~v_513 | v_514;
assign x_10531 = v_513 | ~v_510;
assign x_10532 = v_513 | ~v_511;
assign x_10533 = v_513 | ~v_512;
assign x_10534 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_387 | v_512;
assign x_10535 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_482 | ~v_283 | v_511;
assign x_10536 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_370 | ~v_404 | v_510;
assign x_10537 = ~v_508 | ~v_428 | v_509;
assign x_10538 = v_508 | ~v_483;
assign x_10539 = v_508 | ~v_504;
assign x_10540 = v_508 | ~v_505;
assign x_10541 = v_508 | ~v_506;
assign x_10542 = v_508 | ~v_507;
assign x_10543 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_482 | ~v_317 | v_507;
assign x_10544 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_463 | v_506;
assign x_10545 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_423 | ~v_503 | v_505;
assign x_10546 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_503 | ~v_487 | v_504;
assign x_10547 = v_503 | ~v_492;
assign x_10548 = v_503 | ~v_497;
assign x_10549 = v_503 | ~v_502;
assign x_10550 = v_76 | v_75 | v_73 | v_70 | v_106 | v_104 | v_127 | v_113 | v_112 | ~v_460 | ~v_190 | ~v_189 | ~v_459 | ~v_458 | ~v_186 | ~v_185 | ~v_182 | ~v_181 | ~v_501 | ~v_500 | ~v_454 | ~v_453 | ~v_499 | ~v_498 | ~v_452 | ~v_174 | ~v_173 | v_502;
assign x_10551 = v_501 | v_129;
assign x_10552 = v_501 | v_91;
assign x_10553 = v_500 | ~v_129;
assign x_10554 = v_500 | v_83;
assign x_10555 = v_499 | v_130;
assign x_10556 = v_499 | v_16;
assign x_10557 = v_498 | ~v_130;
assign x_10558 = v_498 | v_13;
assign x_10559 = v_50 | v_51 | v_48 | v_45 | v_100 | v_102 | v_111 | v_110 | v_126 | ~v_449 | ~v_447 | ~v_171 | ~v_170 | ~v_446 | ~v_445 | ~v_167 | ~v_166 | ~v_163 | ~v_162 | ~v_496 | ~v_495 | ~v_494 | ~v_493 | ~v_442 | ~v_441 | ~v_155 | ~v_154 | v_497;
assign x_10560 = v_496 | v_129;
assign x_10561 = v_496 | v_66;
assign x_10562 = v_495 | ~v_129;
assign x_10563 = v_495 | v_58;
assign x_10564 = v_494 | v_130;
assign x_10565 = v_494 | v_14;
assign x_10566 = v_493 | ~v_130;
assign x_10567 = v_493 | v_12;
assign x_10568 = v_25 | v_24 | v_22 | v_19 | v_95 | v_93 | v_108 | v_109 | v_122 | ~v_437 | ~v_152 | ~v_151 | ~v_436 | ~v_435 | ~v_148 | ~v_147 | ~v_144 | ~v_143 | ~v_491 | ~v_490 | ~v_432 | ~v_489 | ~v_488 | ~v_431 | ~v_430 | ~v_136 | ~v_135 | v_492;
assign x_10569 = v_491 | v_129;
assign x_10570 = v_491 | v_41;
assign x_10571 = v_490 | ~v_129;
assign x_10572 = v_490 | v_33;
assign x_10573 = v_489 | v_130;
assign x_10574 = v_489 | v_15;
assign x_10575 = v_488 | ~v_130;
assign x_10576 = v_488 | v_11;
assign x_10577 = v_487 | ~v_484;
assign x_10578 = v_487 | ~v_485;
assign x_10579 = v_487 | ~v_486;
assign x_10580 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_423 | v_486;
assign x_10581 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_463 | ~v_244 | v_485;
assign x_10582 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_317 | ~v_370 | v_484;
assign x_10583 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_482 | ~v_466 | v_483;
assign x_10584 = v_482 | ~v_471;
assign x_10585 = v_482 | ~v_476;
assign x_10586 = v_482 | ~v_481;
assign x_10587 = v_76 | v_74 | v_73 | v_107 | v_106 | v_105 | v_104 | v_113 | v_112 | ~v_460 | ~v_368 | ~v_190 | ~v_189 | ~v_367 | ~v_459 | ~v_458 | ~v_366 | ~v_365 | ~v_454 | ~v_453 | ~v_480 | ~v_479 | ~v_478 | ~v_477 | ~v_362 | ~v_361 | ~v_452 | v_481;
assign x_10588 = v_480 | v_118;
assign x_10589 = v_480 | v_91;
assign x_10590 = v_479 | ~v_118;
assign x_10591 = v_479 | v_83;
assign x_10592 = v_478 | v_119;
assign x_10593 = v_478 | v_16;
assign x_10594 = v_477 | ~v_119;
assign x_10595 = v_477 | v_13;
assign x_10596 = v_51 | v_49 | v_48 | v_103 | v_101 | v_100 | v_102 | v_111 | v_110 | ~v_449 | ~v_447 | ~v_171 | ~v_170 | ~v_357 | ~v_356 | ~v_446 | ~v_445 | ~v_475 | ~v_474 | ~v_355 | ~v_354 | ~v_473 | ~v_472 | ~v_351 | ~v_350 | ~v_442 | ~v_441 | v_476;
assign x_10597 = v_475 | ~v_119;
assign x_10598 = v_475 | v_12;
assign x_10599 = v_474 | v_119;
assign x_10600 = v_474 | v_14;
assign x_10601 = v_473 | v_118;
assign x_10602 = v_473 | v_66;
assign x_10603 = v_472 | ~v_118;
assign x_10604 = v_472 | v_58;
assign x_10605 = v_25 | v_23 | v_22 | v_96 | v_95 | v_94 | v_93 | v_108 | v_109 | ~v_470 | ~v_437 | ~v_152 | ~v_151 | ~v_346 | ~v_345 | ~v_436 | ~v_435 | ~v_469 | ~v_344 | ~v_343 | ~v_432 | ~v_468 | ~v_467 | ~v_340 | ~v_339 | ~v_431 | ~v_430 | v_471;
assign x_10606 = v_470 | ~v_119;
assign x_10607 = v_470 | v_11;
assign x_10608 = v_469 | v_119;
assign x_10609 = v_469 | v_15;
assign x_10610 = v_468 | v_118;
assign x_10611 = v_468 | v_41;
assign x_10612 = v_467 | ~v_118;
assign x_10613 = v_467 | v_33;
assign x_10614 = v_466 | ~v_429;
assign x_10615 = v_466 | ~v_464;
assign x_10616 = v_466 | ~v_465;
assign x_10617 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_317 | v_465;
assign x_10618 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_463 | ~v_334 | v_464;
assign x_10619 = v_463 | ~v_440;
assign x_10620 = v_463 | ~v_451;
assign x_10621 = v_463 | ~v_462;
assign x_10622 = v_75 | v_74 | v_73 | v_72 | v_105 | v_104 | v_113 | v_112 | v_121 | ~v_461 | ~v_460 | ~v_190 | ~v_189 | ~v_315 | ~v_314 | ~v_459 | ~v_458 | ~v_311 | ~v_310 | ~v_457 | ~v_456 | ~v_455 | ~v_454 | ~v_453 | ~v_307 | ~v_306 | ~v_452 | v_462;
assign x_10623 = v_461 | ~v_98;
assign x_10624 = v_461 | v_13;
assign x_10625 = v_460 | v_130;
assign x_10626 = v_460 | v_88;
assign x_10627 = v_459 | v_129;
assign x_10628 = v_459 | v_86;
assign x_10629 = v_458 | ~v_129;
assign x_10630 = v_458 | v_78;
assign x_10631 = v_457 | v_98;
assign x_10632 = v_457 | v_16;
assign x_10633 = v_456 | v_97;
assign x_10634 = v_456 | v_91;
assign x_10635 = v_455 | ~v_97;
assign x_10636 = v_455 | v_83;
assign x_10637 = v_454 | v_99;
assign x_10638 = v_454 | v_89;
assign x_10639 = v_453 | ~v_99;
assign x_10640 = v_453 | v_81;
assign x_10641 = v_452 | ~v_130;
assign x_10642 = v_452 | v_80;
assign x_10643 = v_50 | v_49 | v_48 | v_47 | v_101 | v_100 | v_111 | v_110 | v_120 | ~v_450 | ~v_449 | ~v_448 | ~v_447 | ~v_304 | ~v_171 | ~v_170 | ~v_303 | ~v_302 | ~v_446 | ~v_445 | ~v_444 | ~v_297 | ~v_443 | ~v_296 | ~v_295 | ~v_442 | ~v_441 | v_451;
assign x_10644 = v_450 | ~v_97;
assign x_10645 = v_450 | v_58;
assign x_10646 = v_449 | v_99;
assign x_10647 = v_449 | v_64;
assign x_10648 = v_448 | ~v_98;
assign x_10649 = v_448 | v_12;
assign x_10650 = v_447 | ~v_99;
assign x_10651 = v_447 | v_56;
assign x_10652 = v_446 | v_129;
assign x_10653 = v_446 | v_61;
assign x_10654 = v_445 | ~v_129;
assign x_10655 = v_445 | v_53;
assign x_10656 = v_444 | v_98;
assign x_10657 = v_444 | v_14;
assign x_10658 = v_443 | v_97;
assign x_10659 = v_443 | v_66;
assign x_10660 = v_442 | v_130;
assign x_10661 = v_442 | v_63;
assign x_10662 = v_441 | ~v_130;
assign x_10663 = v_441 | v_55;
assign x_10664 = v_24 | v_23 | v_22 | v_21 | v_94 | v_93 | v_108 | v_109 | v_117 | ~v_439 | ~v_438 | ~v_437 | ~v_293 | ~v_152 | ~v_151 | ~v_292 | ~v_291 | ~v_436 | ~v_435 | ~v_286 | ~v_434 | ~v_433 | ~v_432 | ~v_285 | ~v_284 | ~v_431 | ~v_430 | v_440;
assign x_10665 = v_439 | v_97;
assign x_10666 = v_439 | v_41;
assign x_10667 = v_438 | ~v_97;
assign x_10668 = v_438 | v_33;
assign x_10669 = v_437 | ~v_99;
assign x_10670 = v_437 | v_31;
assign x_10671 = v_436 | v_129;
assign x_10672 = v_436 | v_36;
assign x_10673 = v_435 | ~v_129;
assign x_10674 = v_435 | v_28;
assign x_10675 = v_434 | v_98;
assign x_10676 = v_434 | v_15;
assign x_10677 = v_433 | ~v_98;
assign x_10678 = v_433 | v_11;
assign x_10679 = v_432 | v_99;
assign x_10680 = v_432 | v_39;
assign x_10681 = v_431 | v_130;
assign x_10682 = v_431 | v_38;
assign x_10683 = v_430 | ~v_130;
assign x_10684 = v_430 | v_30;
assign x_10685 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_423 | ~v_192 | v_429;
assign x_10686 = v_428 | ~v_371;
assign x_10687 = v_428 | ~v_424;
assign x_10688 = v_428 | ~v_425;
assign x_10689 = v_428 | ~v_426;
assign x_10690 = v_428 | ~v_427;
assign x_10691 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_244 | v_427;
assign x_10692 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_423 | ~v_283 | v_426;
assign x_10693 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_370 | ~v_334 | v_425;
assign x_10694 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_423 | ~v_407 | v_424;
assign x_10695 = v_423 | ~v_412;
assign x_10696 = v_423 | ~v_417;
assign x_10697 = v_423 | ~v_422;
assign x_10698 = v_76 | v_68 | v_75 | v_74 | v_72 | v_105 | v_104 | v_132 | v_113 | ~v_190 | ~v_189 | ~v_242 | ~v_241 | ~v_315 | ~v_314 | ~v_238 | ~v_237 | ~v_236 | ~v_235 | ~v_311 | ~v_310 | ~v_421 | ~v_420 | ~v_419 | ~v_418 | ~v_307 | ~v_306 | v_422;
assign x_10699 = v_421 | v_123;
assign x_10700 = v_421 | v_91;
assign x_10701 = v_420 | ~v_123;
assign x_10702 = v_420 | v_83;
assign x_10703 = v_419 | v_124;
assign x_10704 = v_419 | v_16;
assign x_10705 = v_418 | ~v_124;
assign x_10706 = v_418 | v_13;
assign x_10707 = v_50 | v_51 | v_49 | v_43 | v_47 | v_101 | v_100 | v_111 | v_131 | ~v_304 | ~v_171 | ~v_170 | ~v_223 | ~v_222 | ~v_303 | ~v_302 | ~v_219 | ~v_218 | ~v_416 | ~v_217 | ~v_216 | ~v_415 | ~v_297 | ~v_414 | ~v_413 | ~v_296 | ~v_295 | v_417;
assign x_10708 = v_416 | ~v_124;
assign x_10709 = v_416 | v_12;
assign x_10710 = v_415 | v_124;
assign x_10711 = v_415 | v_14;
assign x_10712 = v_414 | v_123;
assign x_10713 = v_414 | v_66;
assign x_10714 = v_413 | ~v_123;
assign x_10715 = v_413 | v_58;
assign x_10716 = v_25 | v_24 | v_23 | v_21 | v_17 | v_94 | v_93 | v_109 | v_128 | ~v_293 | ~v_152 | ~v_151 | ~v_207 | ~v_206 | ~v_292 | ~v_291 | ~v_203 | ~v_202 | ~v_411 | ~v_410 | ~v_201 | ~v_200 | ~v_286 | ~v_409 | ~v_408 | ~v_285 | ~v_284 | v_412;
assign x_10717 = v_411 | v_124;
assign x_10718 = v_411 | v_15;
assign x_10719 = v_410 | ~v_124;
assign x_10720 = v_410 | v_11;
assign x_10721 = v_409 | v_123;
assign x_10722 = v_409 | v_41;
assign x_10723 = v_408 | ~v_123;
assign x_10724 = v_408 | v_33;
assign x_10725 = v_407 | ~v_388;
assign x_10726 = v_407 | ~v_405;
assign x_10727 = v_407 | ~v_406;
assign x_10728 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_283 | v_406;
assign x_10729 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_244 | ~v_404 | v_405;
assign x_10730 = v_404 | ~v_393;
assign x_10731 = v_404 | ~v_398;
assign x_10732 = v_404 | ~v_403;
assign x_10733 = v_76 | v_75 | v_73 | v_71 | v_70 | v_106 | v_104 | v_127 | v_112 | ~v_190 | ~v_189 | ~v_280 | ~v_279 | ~v_278 | ~v_277 | ~v_276 | ~v_186 | ~v_185 | ~v_402 | ~v_401 | ~v_182 | ~v_181 | ~v_273 | ~v_400 | ~v_399 | ~v_174 | ~v_173 | v_403;
assign x_10734 = v_402 | v_124;
assign x_10735 = v_402 | v_91;
assign x_10736 = v_401 | ~v_124;
assign x_10737 = v_401 | v_83;
assign x_10738 = v_400 | v_123;
assign x_10739 = v_400 | v_16;
assign x_10740 = v_399 | ~v_123;
assign x_10741 = v_399 | v_13;
assign x_10742 = v_50 | v_51 | v_48 | v_46 | v_45 | v_100 | v_102 | v_110 | v_126 | ~v_268 | ~v_171 | ~v_170 | ~v_267 | ~v_266 | ~v_264 | ~v_263 | ~v_167 | ~v_166 | ~v_397 | ~v_396 | ~v_163 | ~v_162 | ~v_261 | ~v_395 | ~v_394 | ~v_155 | ~v_154 | v_398;
assign x_10743 = v_397 | v_124;
assign x_10744 = v_397 | v_66;
assign x_10745 = v_396 | ~v_124;
assign x_10746 = v_396 | v_58;
assign x_10747 = v_395 | v_123;
assign x_10748 = v_395 | v_14;
assign x_10749 = v_394 | ~v_123;
assign x_10750 = v_394 | v_12;
assign x_10751 = v_25 | v_24 | v_22 | v_20 | v_19 | v_95 | v_93 | v_108 | v_122 | ~v_152 | ~v_151 | ~v_257 | ~v_256 | ~v_255 | ~v_254 | ~v_148 | ~v_147 | ~v_392 | ~v_391 | ~v_144 | ~v_143 | ~v_253 | ~v_252 | ~v_390 | ~v_389 | ~v_136 | ~v_135 | v_393;
assign x_10752 = v_392 | v_124;
assign x_10753 = v_392 | v_41;
assign x_10754 = v_391 | ~v_124;
assign x_10755 = v_391 | v_33;
assign x_10756 = v_390 | v_123;
assign x_10757 = v_390 | v_15;
assign x_10758 = v_389 | ~v_123;
assign x_10759 = v_389 | v_11;
assign x_10760 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_334 | ~v_387 | v_388;
assign x_10761 = v_387 | ~v_376;
assign x_10762 = v_387 | ~v_381;
assign x_10763 = v_387 | ~v_386;
assign x_10764 = v_76 | v_75 | v_74 | v_73 | v_71 | v_106 | v_105 | v_104 | v_112 | ~v_368 | ~v_190 | ~v_189 | ~v_367 | ~v_280 | ~v_279 | ~v_278 | ~v_277 | ~v_276 | ~v_366 | ~v_365 | ~v_273 | ~v_385 | ~v_384 | ~v_362 | ~v_361 | ~v_383 | ~v_382 | v_386;
assign x_10765 = v_385 | v_114;
assign x_10766 = v_385 | v_16;
assign x_10767 = v_384 | ~v_114;
assign x_10768 = v_384 | v_13;
assign x_10769 = v_383 | v_115;
assign x_10770 = v_383 | v_91;
assign x_10771 = v_382 | ~v_115;
assign x_10772 = v_382 | v_83;
assign x_10773 = v_50 | v_51 | v_49 | v_48 | v_46 | v_101 | v_100 | v_102 | v_110 | ~v_268 | ~v_171 | ~v_170 | ~v_357 | ~v_356 | ~v_267 | ~v_266 | ~v_380 | ~v_379 | ~v_264 | ~v_263 | ~v_355 | ~v_354 | ~v_261 | ~v_351 | ~v_350 | ~v_378 | ~v_377 | v_381;
assign x_10774 = v_380 | ~v_114;
assign x_10775 = v_380 | v_12;
assign x_10776 = v_379 | v_114;
assign x_10777 = v_379 | v_14;
assign x_10778 = v_378 | v_115;
assign x_10779 = v_378 | v_66;
assign x_10780 = v_377 | ~v_115;
assign x_10781 = v_377 | v_58;
assign x_10782 = v_25 | v_24 | v_23 | v_22 | v_20 | v_95 | v_94 | v_93 | v_108 | ~v_375 | ~v_152 | ~v_151 | ~v_346 | ~v_345 | ~v_257 | ~v_256 | ~v_374 | ~v_255 | ~v_254 | ~v_344 | ~v_343 | ~v_253 | ~v_252 | ~v_340 | ~v_339 | ~v_373 | ~v_372 | v_376;
assign x_10783 = v_375 | ~v_114;
assign x_10784 = v_375 | v_11;
assign x_10785 = v_374 | v_114;
assign x_10786 = v_374 | v_15;
assign x_10787 = v_373 | v_115;
assign x_10788 = v_373 | v_41;
assign x_10789 = v_372 | ~v_115;
assign x_10790 = v_372 | v_33;
assign x_10791 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_370 | ~v_336 | v_371;
assign x_10792 = v_370 | ~v_347;
assign x_10793 = v_370 | ~v_358;
assign x_10794 = v_370 | ~v_369;
assign x_10795 = v_68 | v_75 | v_74 | v_106 | v_105 | v_104 | v_132 | v_113 | v_121 | ~v_368 | ~v_190 | ~v_189 | ~v_242 | ~v_241 | ~v_367 | ~v_238 | ~v_237 | ~v_236 | ~v_235 | ~v_366 | ~v_365 | ~v_364 | ~v_363 | ~v_362 | ~v_361 | ~v_360 | ~v_359 | v_369;
assign x_10796 = v_368 | v_134;
assign x_10797 = v_368 | v_87;
assign x_10798 = v_367 | ~v_134;
assign x_10799 = v_367 | v_79;
assign x_10800 = v_366 | v_133;
assign x_10801 = v_366 | v_90;
assign x_10802 = v_365 | ~v_133;
assign x_10803 = v_365 | v_82;
assign x_10804 = v_364 | v_133;
assign x_10805 = v_364 | v_91;
assign x_10806 = v_363 | ~v_133;
assign x_10807 = v_363 | v_83;
assign x_10808 = v_362 | v_116;
assign x_10809 = v_362 | v_92;
assign x_10810 = v_361 | ~v_116;
assign x_10811 = v_361 | v_84;
assign x_10812 = v_360 | v_134;
assign x_10813 = v_360 | v_16;
assign x_10814 = v_359 | ~v_134;
assign x_10815 = v_359 | v_13;
assign x_10816 = v_50 | v_49 | v_43 | v_101 | v_100 | v_102 | v_111 | v_131 | v_120 | ~v_171 | ~v_170 | ~v_223 | ~v_222 | ~v_357 | ~v_356 | ~v_219 | ~v_218 | ~v_217 | ~v_216 | ~v_355 | ~v_354 | ~v_353 | ~v_352 | ~v_351 | ~v_350 | ~v_349 | ~v_348 | v_358;
assign x_10817 = v_357 | v_134;
assign x_10818 = v_357 | v_62;
assign x_10819 = v_356 | ~v_134;
assign x_10820 = v_356 | v_54;
assign x_10821 = v_355 | v_133;
assign x_10822 = v_355 | v_65;
assign x_10823 = v_354 | ~v_133;
assign x_10824 = v_354 | v_57;
assign x_10825 = v_353 | v_133;
assign x_10826 = v_353 | v_66;
assign x_10827 = v_352 | ~v_133;
assign x_10828 = v_352 | v_58;
assign x_10829 = v_351 | v_116;
assign x_10830 = v_351 | v_67;
assign x_10831 = v_350 | ~v_116;
assign x_10832 = v_350 | v_59;
assign x_10833 = v_349 | v_134;
assign x_10834 = v_349 | v_14;
assign x_10835 = v_348 | ~v_134;
assign x_10836 = v_348 | v_12;
assign x_10837 = v_24 | v_23 | v_17 | v_95 | v_94 | v_93 | v_109 | v_128 | v_117 | ~v_152 | ~v_151 | ~v_207 | ~v_206 | ~v_346 | ~v_345 | ~v_203 | ~v_202 | ~v_201 | ~v_200 | ~v_344 | ~v_343 | ~v_342 | ~v_341 | ~v_340 | ~v_339 | ~v_338 | ~v_337 | v_347;
assign x_10838 = v_346 | v_134;
assign x_10839 = v_346 | v_37;
assign x_10840 = v_345 | ~v_134;
assign x_10841 = v_345 | v_29;
assign x_10842 = v_344 | v_133;
assign x_10843 = v_344 | v_40;
assign x_10844 = v_343 | ~v_133;
assign x_10845 = v_343 | v_32;
assign x_10846 = v_342 | v_133;
assign x_10847 = v_342 | v_41;
assign x_10848 = v_341 | ~v_133;
assign x_10849 = v_341 | v_33;
assign x_10850 = v_340 | v_116;
assign x_10851 = v_340 | v_42;
assign x_10852 = v_339 | ~v_116;
assign x_10853 = v_339 | v_34;
assign x_10854 = v_338 | v_134;
assign x_10855 = v_338 | v_15;
assign x_10856 = v_337 | ~v_134;
assign x_10857 = v_337 | v_11;
assign x_10858 = v_336 | ~v_249;
assign x_10859 = v_336 | ~v_318;
assign x_10860 = v_336 | ~v_335;
assign x_10861 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_334 | v_335;
assign x_10862 = v_334 | ~v_323;
assign x_10863 = v_334 | ~v_328;
assign x_10864 = v_334 | ~v_333;
assign x_10865 = v_75 | v_74 | v_73 | v_106 | v_105 | v_104 | v_113 | v_112 | v_121 | ~v_190 | ~v_189 | ~v_240 | ~v_239 | ~v_188 | ~v_187 | ~v_332 | ~v_331 | ~v_180 | ~v_179 | ~v_232 | ~v_231 | ~v_230 | ~v_229 | ~v_330 | ~v_329 | ~v_176 | ~v_175 | v_333;
assign x_10866 = v_332 | v_119;
assign x_10867 = v_332 | v_91;
assign x_10868 = v_331 | ~v_119;
assign x_10869 = v_331 | v_83;
assign x_10870 = v_330 | v_118;
assign x_10871 = v_330 | v_16;
assign x_10872 = v_329 | ~v_118;
assign x_10873 = v_329 | v_13;
assign x_10874 = v_50 | v_49 | v_48 | v_101 | v_100 | v_102 | v_111 | v_110 | v_120 | ~v_225 | ~v_224 | ~v_171 | ~v_170 | ~v_221 | ~v_220 | ~v_169 | ~v_168 | ~v_327 | ~v_326 | ~v_161 | ~v_160 | ~v_211 | ~v_210 | ~v_325 | ~v_324 | ~v_157 | ~v_156 | v_328;
assign x_10875 = v_327 | v_119;
assign x_10876 = v_327 | v_66;
assign x_10877 = v_326 | ~v_119;
assign x_10878 = v_326 | v_58;
assign x_10879 = v_325 | v_118;
assign x_10880 = v_325 | v_14;
assign x_10881 = v_324 | ~v_118;
assign x_10882 = v_324 | v_12;
assign x_10883 = v_24 | v_23 | v_22 | v_95 | v_94 | v_93 | v_108 | v_109 | v_117 | ~v_208 | ~v_152 | ~v_151 | ~v_205 | ~v_204 | ~v_150 | ~v_149 | ~v_322 | ~v_321 | ~v_142 | ~v_141 | ~v_195 | ~v_194 | ~v_193 | ~v_320 | ~v_319 | ~v_138 | ~v_137 | v_323;
assign x_10884 = v_322 | v_119;
assign x_10885 = v_322 | v_41;
assign x_10886 = v_321 | ~v_119;
assign x_10887 = v_321 | v_33;
assign x_10888 = v_320 | v_118;
assign x_10889 = v_320 | v_15;
assign x_10890 = v_319 | ~v_118;
assign x_10891 = v_319 | v_11;
assign x_10892 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_317 | ~v_283 | v_318;
assign x_10893 = v_317 | ~v_294;
assign x_10894 = v_317 | ~v_305;
assign x_10895 = v_317 | ~v_316;
assign x_10896 = v_76 | v_75 | v_74 | v_73 | v_72 | v_105 | v_104 | v_113 | v_112 | ~v_190 | ~v_189 | ~v_315 | ~v_314 | ~v_188 | ~v_187 | ~v_180 | ~v_179 | ~v_313 | ~v_312 | ~v_311 | ~v_310 | ~v_309 | ~v_308 | ~v_307 | ~v_306 | ~v_176 | ~v_175 | v_316;
assign x_10897 = v_315 | v_124;
assign x_10898 = v_315 | v_87;
assign x_10899 = v_314 | ~v_124;
assign x_10900 = v_314 | v_79;
assign x_10901 = v_313 | v_114;
assign x_10902 = v_313 | v_91;
assign x_10903 = v_312 | ~v_114;
assign x_10904 = v_312 | v_83;
assign x_10905 = v_311 | v_92;
assign x_10906 = v_311 | v_26;
assign x_10907 = v_310 | v_84;
assign x_10908 = v_310 | ~v_26;
assign x_10909 = v_309 | v_115;
assign x_10910 = v_309 | v_16;
assign x_10911 = v_308 | ~v_115;
assign x_10912 = v_308 | v_13;
assign x_10913 = v_307 | v_123;
assign x_10914 = v_307 | v_90;
assign x_10915 = v_306 | ~v_123;
assign x_10916 = v_306 | v_82;
assign x_10917 = v_50 | v_51 | v_49 | v_48 | v_47 | v_101 | v_100 | v_111 | v_110 | ~v_304 | ~v_171 | ~v_170 | ~v_303 | ~v_302 | ~v_169 | ~v_168 | ~v_301 | ~v_300 | ~v_161 | ~v_160 | ~v_299 | ~v_298 | ~v_297 | ~v_296 | ~v_295 | ~v_157 | ~v_156 | v_305;
assign x_10918 = v_304 | v_67;
assign x_10919 = v_304 | v_26;
assign x_10920 = v_303 | v_124;
assign x_10921 = v_303 | v_62;
assign x_10922 = v_302 | ~v_124;
assign x_10923 = v_302 | v_54;
assign x_10924 = v_301 | ~v_115;
assign x_10925 = v_301 | v_12;
assign x_10926 = v_300 | v_115;
assign x_10927 = v_300 | v_14;
assign x_10928 = v_299 | v_114;
assign x_10929 = v_299 | v_66;
assign x_10930 = v_298 | ~v_114;
assign x_10931 = v_298 | v_58;
assign x_10932 = v_297 | v_59;
assign x_10933 = v_297 | ~v_26;
assign x_10934 = v_296 | v_123;
assign x_10935 = v_296 | v_65;
assign x_10936 = v_295 | ~v_123;
assign x_10937 = v_295 | v_57;
assign x_10938 = v_25 | v_24 | v_23 | v_22 | v_21 | v_94 | v_93 | v_108 | v_109 | ~v_293 | ~v_152 | ~v_151 | ~v_292 | ~v_291 | ~v_150 | ~v_149 | ~v_290 | ~v_289 | ~v_142 | ~v_141 | ~v_288 | ~v_287 | ~v_286 | ~v_285 | ~v_284 | ~v_138 | ~v_137 | v_294;
assign x_10939 = v_293 | v_42;
assign x_10940 = v_293 | v_26;
assign x_10941 = v_292 | v_124;
assign x_10942 = v_292 | v_37;
assign x_10943 = v_291 | ~v_124;
assign x_10944 = v_291 | v_29;
assign x_10945 = v_290 | v_115;
assign x_10946 = v_290 | v_15;
assign x_10947 = v_289 | ~v_115;
assign x_10948 = v_289 | v_11;
assign x_10949 = v_288 | v_114;
assign x_10950 = v_288 | v_41;
assign x_10951 = v_287 | ~v_114;
assign x_10952 = v_287 | v_33;
assign x_10953 = v_286 | v_34;
assign x_10954 = v_286 | ~v_26;
assign x_10955 = v_285 | v_123;
assign x_10956 = v_285 | v_40;
assign x_10957 = v_284 | ~v_123;
assign x_10958 = v_284 | v_32;
assign x_10959 = v_283 | ~v_260;
assign x_10960 = v_283 | ~v_271;
assign x_10961 = v_283 | ~v_282;
assign x_10962 = v_76 | v_74 | v_73 | v_71 | v_107 | v_106 | v_105 | v_104 | v_112 | ~v_281 | ~v_190 | ~v_189 | ~v_240 | ~v_239 | ~v_280 | ~v_279 | ~v_278 | ~v_277 | ~v_276 | ~v_232 | ~v_231 | ~v_275 | ~v_274 | ~v_273 | ~v_272 | ~v_230 | ~v_229 | v_282;
assign x_10963 = v_281 | ~v_97;
assign x_10964 = v_281 | v_13;
assign x_10965 = v_280 | v_124;
assign x_10966 = v_280 | v_86;
assign x_10967 = v_279 | ~v_124;
assign x_10968 = v_279 | v_78;
assign x_10969 = v_278 | v_89;
assign x_10970 = v_278 | v_26;
assign x_10971 = v_277 | v_123;
assign x_10972 = v_277 | v_88;
assign x_10973 = v_276 | ~v_123;
assign x_10974 = v_276 | v_80;
assign x_10975 = v_275 | v_91;
assign x_10976 = v_275 | v_98;
assign x_10977 = v_274 | ~v_98;
assign x_10978 = v_274 | v_83;
assign x_10979 = v_273 | v_81;
assign x_10980 = v_273 | ~v_26;
assign x_10981 = v_272 | v_97;
assign x_10982 = v_272 | v_16;
assign x_10983 = v_51 | v_49 | v_48 | v_46 | v_103 | v_101 | v_100 | v_102 | v_110 | ~v_270 | ~v_225 | ~v_269 | ~v_224 | ~v_268 | ~v_171 | ~v_170 | ~v_221 | ~v_220 | ~v_267 | ~v_266 | ~v_265 | ~v_264 | ~v_263 | ~v_211 | ~v_210 | ~v_262 | ~v_261 | v_271;
assign x_10984 = v_270 | ~v_97;
assign x_10985 = v_270 | v_12;
assign x_10986 = v_269 | ~v_98;
assign x_10987 = v_269 | v_58;
assign x_10988 = v_268 | v_64;
assign x_10989 = v_268 | v_26;
assign x_10990 = v_267 | v_124;
assign x_10991 = v_267 | v_61;
assign x_10992 = v_266 | ~v_124;
assign x_10993 = v_266 | v_53;
assign x_10994 = v_265 | v_97;
assign x_10995 = v_265 | v_14;
assign x_10996 = v_264 | v_123;
assign x_10997 = v_264 | v_63;
assign x_10998 = v_263 | ~v_123;
assign x_10999 = v_263 | v_55;
assign x_11000 = v_262 | v_98;
assign x_11001 = v_262 | v_66;
assign x_11002 = v_261 | v_56;
assign x_11003 = v_261 | ~v_26;
assign x_11004 = v_25 | v_23 | v_22 | v_20 | v_96 | v_95 | v_94 | v_93 | v_108 | ~v_259 | ~v_258 | ~v_208 | ~v_152 | ~v_151 | ~v_205 | ~v_204 | ~v_257 | ~v_256 | ~v_255 | ~v_254 | ~v_195 | ~v_194 | ~v_253 | ~v_252 | ~v_251 | ~v_250 | ~v_193 | v_260;
assign x_11005 = v_259 | v_98;
assign x_11006 = v_259 | v_41;
assign x_11007 = v_258 | ~v_98;
assign x_11008 = v_258 | v_33;
assign x_11009 = v_257 | v_124;
assign x_11010 = v_257 | v_36;
assign x_11011 = v_256 | ~v_124;
assign x_11012 = v_256 | v_28;
assign x_11013 = v_255 | v_123;
assign x_11014 = v_255 | v_38;
assign x_11015 = v_254 | ~v_123;
assign x_11016 = v_254 | v_30;
assign x_11017 = v_253 | v_39;
assign x_11018 = v_253 | v_26;
assign x_11019 = v_252 | v_31;
assign x_11020 = v_252 | ~v_26;
assign x_11021 = v_251 | v_97;
assign x_11022 = v_251 | v_15;
assign x_11023 = v_250 | ~v_97;
assign x_11024 = v_250 | v_11;
assign x_11025 = ~v_248 | ~v_247 | ~v_246 | ~v_245 | ~v_244 | ~v_192 | v_249;
assign x_11026 = v_248 | v_12;
assign x_11027 = v_248 | ~v_11;
assign x_11028 = v_247 | v_13;
assign x_11029 = v_247 | ~v_12;
assign x_11030 = v_246 | v_15;
assign x_11031 = v_246 | ~v_14;
assign x_11032 = v_245 | v_14;
assign x_11033 = v_245 | ~v_16;
assign x_11034 = v_244 | ~v_209;
assign x_11035 = v_244 | ~v_226;
assign x_11036 = v_244 | ~v_243;
assign x_11037 = v_76 | v_68 | v_75 | v_74 | v_106 | v_105 | v_104 | v_132 | v_113 | ~v_190 | ~v_189 | ~v_242 | ~v_241 | ~v_240 | ~v_239 | ~v_238 | ~v_237 | ~v_236 | ~v_235 | ~v_234 | ~v_233 | ~v_232 | ~v_231 | ~v_230 | ~v_229 | ~v_228 | ~v_227 | v_243;
assign x_11038 = v_242 | v_125;
assign x_11039 = v_242 | v_88;
assign x_11040 = v_241 | ~v_125;
assign x_11041 = v_241 | v_80;
assign x_11042 = v_240 | v_129;
assign x_11043 = v_240 | v_87;
assign x_11044 = v_239 | ~v_129;
assign x_11045 = v_239 | v_79;
assign x_11046 = v_238 | v_125;
assign x_11047 = v_238 | v_86;
assign x_11048 = v_237 | ~v_125;
assign x_11049 = v_237 | v_78;
assign x_11050 = v_236 | v_125;
assign x_11051 = v_236 | v_89;
assign x_11052 = v_235 | ~v_125;
assign x_11053 = v_235 | v_81;
assign x_11054 = v_234 | v_130;
assign x_11055 = v_234 | v_91;
assign x_11056 = v_233 | ~v_130;
assign x_11057 = v_233 | v_83;
assign x_11058 = v_232 | v_130;
assign x_11059 = v_232 | v_90;
assign x_11060 = v_231 | ~v_130;
assign x_11061 = v_231 | v_82;
assign x_11062 = v_230 | v_92;
assign x_11063 = v_230 | v_99;
assign x_11064 = v_229 | ~v_99;
assign x_11065 = v_229 | v_84;
assign x_11066 = v_228 | v_129;
assign x_11067 = v_228 | v_16;
assign x_11068 = v_227 | ~v_129;
assign x_11069 = v_227 | v_13;
assign x_11070 = v_50 | v_51 | v_49 | v_43 | v_101 | v_100 | v_102 | v_111 | v_131 | ~v_225 | ~v_224 | ~v_171 | ~v_170 | ~v_223 | ~v_222 | ~v_221 | ~v_220 | ~v_219 | ~v_218 | ~v_217 | ~v_216 | ~v_215 | ~v_214 | ~v_213 | ~v_212 | ~v_211 | ~v_210 | v_226;
assign x_11071 = v_225 | v_99;
assign x_11072 = v_225 | v_67;
assign x_11073 = v_224 | ~v_99;
assign x_11074 = v_224 | v_59;
assign x_11075 = v_223 | v_125;
assign x_11076 = v_223 | v_63;
assign x_11077 = v_222 | ~v_125;
assign x_11078 = v_222 | v_55;
assign x_11079 = v_221 | v_129;
assign x_11080 = v_221 | v_62;
assign x_11081 = v_220 | ~v_129;
assign x_11082 = v_220 | v_54;
assign x_11083 = v_219 | v_125;
assign x_11084 = v_219 | v_61;
assign x_11085 = v_218 | ~v_125;
assign x_11086 = v_218 | v_53;
assign x_11087 = v_217 | v_125;
assign x_11088 = v_217 | v_64;
assign x_11089 = v_216 | ~v_125;
assign x_11090 = v_216 | v_56;
assign x_11091 = v_215 | ~v_129;
assign x_11092 = v_215 | v_12;
assign x_11093 = v_214 | v_129;
assign x_11094 = v_214 | v_14;
assign x_11095 = v_213 | v_130;
assign x_11096 = v_213 | v_66;
assign x_11097 = v_212 | ~v_130;
assign x_11098 = v_212 | v_58;
assign x_11099 = v_211 | v_130;
assign x_11100 = v_211 | v_65;
assign x_11101 = v_210 | ~v_130;
assign x_11102 = v_210 | v_57;
assign x_11103 = v_25 | v_24 | v_23 | v_17 | v_95 | v_94 | v_93 | v_109 | v_128 | ~v_208 | ~v_152 | ~v_151 | ~v_207 | ~v_206 | ~v_205 | ~v_204 | ~v_203 | ~v_202 | ~v_201 | ~v_200 | ~v_199 | ~v_198 | ~v_197 | ~v_196 | ~v_195 | ~v_194 | ~v_193 | v_209;
assign x_11104 = v_208 | v_99;
assign x_11105 = v_208 | v_42;
assign x_11106 = v_207 | v_125;
assign x_11107 = v_207 | v_38;
assign x_11108 = v_206 | ~v_125;
assign x_11109 = v_206 | v_30;
assign x_11110 = v_205 | v_129;
assign x_11111 = v_205 | v_37;
assign x_11112 = v_204 | ~v_129;
assign x_11113 = v_204 | v_29;
assign x_11114 = v_203 | v_125;
assign x_11115 = v_203 | v_36;
assign x_11116 = v_202 | ~v_125;
assign x_11117 = v_202 | v_28;
assign x_11118 = v_201 | v_125;
assign x_11119 = v_201 | v_39;
assign x_11120 = v_200 | ~v_125;
assign x_11121 = v_200 | v_31;
assign x_11122 = v_199 | v_129;
assign x_11123 = v_199 | v_15;
assign x_11124 = v_198 | ~v_129;
assign x_11125 = v_198 | v_11;
assign x_11126 = v_197 | v_130;
assign x_11127 = v_197 | v_41;
assign x_11128 = v_196 | ~v_130;
assign x_11129 = v_196 | v_33;
assign x_11130 = v_195 | v_130;
assign x_11131 = v_195 | v_40;
assign x_11132 = v_194 | ~v_130;
assign x_11133 = v_194 | v_32;
assign x_11134 = v_193 | ~v_99;
assign x_11135 = v_193 | v_34;
assign x_11136 = v_192 | ~v_153;
assign x_11137 = v_192 | ~v_172;
assign x_11138 = v_192 | ~v_191;
assign x_11139 = v_76 | v_73 | v_70 | v_107 | v_106 | v_104 | v_127 | v_113 | v_112 | ~v_190 | ~v_189 | ~v_188 | ~v_187 | ~v_186 | ~v_185 | ~v_184 | ~v_183 | ~v_182 | ~v_181 | ~v_180 | ~v_179 | ~v_178 | ~v_177 | ~v_176 | ~v_175 | ~v_174 | ~v_173 | v_191;
assign x_11140 = v_190 | v_125;
assign x_11141 = v_190 | v_85;
assign x_11142 = v_189 | ~v_125;
assign x_11143 = v_189 | v_77;
assign x_11144 = v_188 | v_134;
assign x_11145 = v_188 | v_86;
assign x_11146 = v_187 | ~v_134;
assign x_11147 = v_187 | v_78;
assign x_11148 = v_186 | v_125;
assign x_11149 = v_186 | v_90;
assign x_11150 = v_185 | ~v_125;
assign x_11151 = v_185 | v_82;
assign x_11152 = v_184 | v_134;
assign x_11153 = v_184 | v_91;
assign x_11154 = v_183 | ~v_134;
assign x_11155 = v_183 | v_83;
assign x_11156 = v_182 | v_125;
assign x_11157 = v_182 | v_92;
assign x_11158 = v_181 | ~v_125;
assign x_11159 = v_181 | v_84;
assign x_11160 = v_180 | v_116;
assign x_11161 = v_180 | v_89;
assign x_11162 = v_179 | ~v_116;
assign x_11163 = v_179 | v_81;
assign x_11164 = v_178 | v_133;
assign x_11165 = v_178 | v_16;
assign x_11166 = v_177 | ~v_133;
assign x_11167 = v_177 | v_13;
assign x_11168 = v_176 | v_133;
assign x_11169 = v_176 | v_88;
assign x_11170 = v_175 | ~v_133;
assign x_11171 = v_175 | v_80;
assign x_11172 = v_174 | v_125;
assign x_11173 = v_174 | v_87;
assign x_11174 = v_173 | ~v_125;
assign x_11175 = v_173 | v_79;
assign x_11176 = v_51 | v_48 | v_45 | v_103 | v_100 | v_102 | v_111 | v_110 | v_126 | ~v_171 | ~v_170 | ~v_169 | ~v_168 | ~v_167 | ~v_166 | ~v_165 | ~v_164 | ~v_163 | ~v_162 | ~v_161 | ~v_160 | ~v_159 | ~v_158 | ~v_157 | ~v_156 | ~v_155 | ~v_154 | v_172;
assign x_11177 = v_171 | v_125;
assign x_11178 = v_171 | v_60;
assign x_11179 = v_170 | ~v_125;
assign x_11180 = v_170 | v_52;
assign x_11181 = v_169 | v_134;
assign x_11182 = v_169 | v_61;
assign x_11183 = v_168 | ~v_134;
assign x_11184 = v_168 | v_53;
assign x_11185 = v_167 | v_125;
assign x_11186 = v_167 | v_65;
assign x_11187 = v_166 | ~v_125;
assign x_11188 = v_166 | v_57;
assign x_11189 = v_165 | v_134;
assign x_11190 = v_165 | v_66;
assign x_11191 = v_164 | ~v_134;
assign x_11192 = v_164 | v_58;
assign x_11193 = v_163 | v_125;
assign x_11194 = v_163 | v_67;
assign x_11195 = v_162 | ~v_125;
assign x_11196 = v_162 | v_59;
assign x_11197 = v_161 | v_116;
assign x_11198 = v_161 | v_64;
assign x_11199 = v_160 | ~v_116;
assign x_11200 = v_160 | v_56;
assign x_11201 = v_159 | v_133;
assign x_11202 = v_159 | v_14;
assign x_11203 = v_158 | ~v_133;
assign x_11204 = v_158 | v_12;
assign x_11205 = v_157 | v_133;
assign x_11206 = v_157 | v_63;
assign x_11207 = v_156 | ~v_133;
assign x_11208 = v_156 | v_55;
assign x_11209 = v_155 | v_125;
assign x_11210 = v_155 | v_62;
assign x_11211 = v_154 | ~v_125;
assign x_11212 = v_154 | v_54;
assign x_11213 = v_25 | v_22 | v_19 | v_96 | v_95 | v_93 | v_108 | v_109 | v_122 | ~v_152 | ~v_151 | ~v_150 | ~v_149 | ~v_148 | ~v_147 | ~v_146 | ~v_145 | ~v_144 | ~v_143 | ~v_142 | ~v_141 | ~v_140 | ~v_139 | ~v_138 | ~v_137 | ~v_136 | ~v_135 | v_153;
assign x_11214 = v_152 | v_125;
assign x_11215 = v_152 | v_35;
assign x_11216 = v_151 | ~v_125;
assign x_11217 = v_151 | v_27;
assign x_11218 = v_150 | v_134;
assign x_11219 = v_150 | v_36;
assign x_11220 = v_149 | ~v_134;
assign x_11221 = v_149 | v_28;
assign x_11222 = v_148 | v_125;
assign x_11223 = v_148 | v_40;
assign x_11224 = v_147 | ~v_125;
assign x_11225 = v_147 | v_32;
assign x_11226 = v_146 | v_134;
assign x_11227 = v_146 | v_41;
assign x_11228 = v_145 | ~v_134;
assign x_11229 = v_145 | v_33;
assign x_11230 = v_144 | v_125;
assign x_11231 = v_144 | v_42;
assign x_11232 = v_143 | ~v_125;
assign x_11233 = v_143 | v_34;
assign x_11234 = v_142 | v_116;
assign x_11235 = v_142 | v_39;
assign x_11236 = v_141 | ~v_116;
assign x_11237 = v_141 | v_31;
assign x_11238 = v_140 | v_133;
assign x_11239 = v_140 | v_15;
assign x_11240 = v_139 | ~v_133;
assign x_11241 = v_139 | v_11;
assign x_11242 = v_138 | v_133;
assign x_11243 = v_138 | v_38;
assign x_11244 = v_137 | ~v_133;
assign x_11245 = v_137 | v_30;
assign x_11246 = v_136 | v_125;
assign x_11247 = v_136 | v_37;
assign x_11248 = v_135 | ~v_125;
assign x_11249 = v_135 | v_29;
assign x_11250 = x_1 & x_2;
assign x_11251 = x_4 & x_5;
assign x_11252 = x_3 & x_11251;
assign x_11253 = x_11250 & x_11252;
assign x_11254 = x_6 & x_7;
assign x_11255 = x_9 & x_10;
assign x_11256 = x_8 & x_11255;
assign x_11257 = x_11254 & x_11256;
assign x_11258 = x_11253 & x_11257;
assign x_11259 = x_11 & x_12;
assign x_11260 = x_14 & x_15;
assign x_11261 = x_13 & x_11260;
assign x_11262 = x_11259 & x_11261;
assign x_11263 = x_17 & x_18;
assign x_11264 = x_16 & x_11263;
assign x_11265 = x_20 & x_21;
assign x_11266 = x_19 & x_11265;
assign x_11267 = x_11264 & x_11266;
assign x_11268 = x_11262 & x_11267;
assign x_11269 = x_11258 & x_11268;
assign x_11270 = x_22 & x_23;
assign x_11271 = x_25 & x_26;
assign x_11272 = x_24 & x_11271;
assign x_11273 = x_11270 & x_11272;
assign x_11274 = x_28 & x_29;
assign x_11275 = x_27 & x_11274;
assign x_11276 = x_31 & x_32;
assign x_11277 = x_30 & x_11276;
assign x_11278 = x_11275 & x_11277;
assign x_11279 = x_11273 & x_11278;
assign x_11280 = x_33 & x_34;
assign x_11281 = x_36 & x_37;
assign x_11282 = x_35 & x_11281;
assign x_11283 = x_11280 & x_11282;
assign x_11284 = x_39 & x_40;
assign x_11285 = x_38 & x_11284;
assign x_11286 = x_42 & x_43;
assign x_11287 = x_41 & x_11286;
assign x_11288 = x_11285 & x_11287;
assign x_11289 = x_11283 & x_11288;
assign x_11290 = x_11279 & x_11289;
assign x_11291 = x_11269 & x_11290;
assign x_11292 = x_44 & x_45;
assign x_11293 = x_47 & x_48;
assign x_11294 = x_46 & x_11293;
assign x_11295 = x_11292 & x_11294;
assign x_11296 = x_50 & x_51;
assign x_11297 = x_49 & x_11296;
assign x_11298 = x_53 & x_54;
assign x_11299 = x_52 & x_11298;
assign x_11300 = x_11297 & x_11299;
assign x_11301 = x_11295 & x_11300;
assign x_11302 = x_55 & x_56;
assign x_11303 = x_58 & x_59;
assign x_11304 = x_57 & x_11303;
assign x_11305 = x_11302 & x_11304;
assign x_11306 = x_61 & x_62;
assign x_11307 = x_60 & x_11306;
assign x_11308 = x_64 & x_65;
assign x_11309 = x_63 & x_11308;
assign x_11310 = x_11307 & x_11309;
assign x_11311 = x_11305 & x_11310;
assign x_11312 = x_11301 & x_11311;
assign x_11313 = x_66 & x_67;
assign x_11314 = x_69 & x_70;
assign x_11315 = x_68 & x_11314;
assign x_11316 = x_11313 & x_11315;
assign x_11317 = x_72 & x_73;
assign x_11318 = x_71 & x_11317;
assign x_11319 = x_75 & x_76;
assign x_11320 = x_74 & x_11319;
assign x_11321 = x_11318 & x_11320;
assign x_11322 = x_11316 & x_11321;
assign x_11323 = x_77 & x_78;
assign x_11324 = x_80 & x_81;
assign x_11325 = x_79 & x_11324;
assign x_11326 = x_11323 & x_11325;
assign x_11327 = x_83 & x_84;
assign x_11328 = x_82 & x_11327;
assign x_11329 = x_86 & x_87;
assign x_11330 = x_85 & x_11329;
assign x_11331 = x_11328 & x_11330;
assign x_11332 = x_11326 & x_11331;
assign x_11333 = x_11322 & x_11332;
assign x_11334 = x_11312 & x_11333;
assign x_11335 = x_11291 & x_11334;
assign x_11336 = x_88 & x_89;
assign x_11337 = x_91 & x_92;
assign x_11338 = x_90 & x_11337;
assign x_11339 = x_11336 & x_11338;
assign x_11340 = x_94 & x_95;
assign x_11341 = x_93 & x_11340;
assign x_11342 = x_97 & x_98;
assign x_11343 = x_96 & x_11342;
assign x_11344 = x_11341 & x_11343;
assign x_11345 = x_11339 & x_11344;
assign x_11346 = x_99 & x_100;
assign x_11347 = x_102 & x_103;
assign x_11348 = x_101 & x_11347;
assign x_11349 = x_11346 & x_11348;
assign x_11350 = x_105 & x_106;
assign x_11351 = x_104 & x_11350;
assign x_11352 = x_108 & x_109;
assign x_11353 = x_107 & x_11352;
assign x_11354 = x_11351 & x_11353;
assign x_11355 = x_11349 & x_11354;
assign x_11356 = x_11345 & x_11355;
assign x_11357 = x_110 & x_111;
assign x_11358 = x_113 & x_114;
assign x_11359 = x_112 & x_11358;
assign x_11360 = x_11357 & x_11359;
assign x_11361 = x_116 & x_117;
assign x_11362 = x_115 & x_11361;
assign x_11363 = x_119 & x_120;
assign x_11364 = x_118 & x_11363;
assign x_11365 = x_11362 & x_11364;
assign x_11366 = x_11360 & x_11365;
assign x_11367 = x_121 & x_122;
assign x_11368 = x_124 & x_125;
assign x_11369 = x_123 & x_11368;
assign x_11370 = x_11367 & x_11369;
assign x_11371 = x_127 & x_128;
assign x_11372 = x_126 & x_11371;
assign x_11373 = x_130 & x_131;
assign x_11374 = x_129 & x_11373;
assign x_11375 = x_11372 & x_11374;
assign x_11376 = x_11370 & x_11375;
assign x_11377 = x_11366 & x_11376;
assign x_11378 = x_11356 & x_11377;
assign x_11379 = x_132 & x_133;
assign x_11380 = x_135 & x_136;
assign x_11381 = x_134 & x_11380;
assign x_11382 = x_11379 & x_11381;
assign x_11383 = x_138 & x_139;
assign x_11384 = x_137 & x_11383;
assign x_11385 = x_141 & x_142;
assign x_11386 = x_140 & x_11385;
assign x_11387 = x_11384 & x_11386;
assign x_11388 = x_11382 & x_11387;
assign x_11389 = x_143 & x_144;
assign x_11390 = x_146 & x_147;
assign x_11391 = x_145 & x_11390;
assign x_11392 = x_11389 & x_11391;
assign x_11393 = x_149 & x_150;
assign x_11394 = x_148 & x_11393;
assign x_11395 = x_152 & x_153;
assign x_11396 = x_151 & x_11395;
assign x_11397 = x_11394 & x_11396;
assign x_11398 = x_11392 & x_11397;
assign x_11399 = x_11388 & x_11398;
assign x_11400 = x_154 & x_155;
assign x_11401 = x_157 & x_158;
assign x_11402 = x_156 & x_11401;
assign x_11403 = x_11400 & x_11402;
assign x_11404 = x_160 & x_161;
assign x_11405 = x_159 & x_11404;
assign x_11406 = x_163 & x_164;
assign x_11407 = x_162 & x_11406;
assign x_11408 = x_11405 & x_11407;
assign x_11409 = x_11403 & x_11408;
assign x_11410 = x_165 & x_166;
assign x_11411 = x_168 & x_169;
assign x_11412 = x_167 & x_11411;
assign x_11413 = x_11410 & x_11412;
assign x_11414 = x_171 & x_172;
assign x_11415 = x_170 & x_11414;
assign x_11416 = x_174 & x_175;
assign x_11417 = x_173 & x_11416;
assign x_11418 = x_11415 & x_11417;
assign x_11419 = x_11413 & x_11418;
assign x_11420 = x_11409 & x_11419;
assign x_11421 = x_11399 & x_11420;
assign x_11422 = x_11378 & x_11421;
assign x_11423 = x_11335 & x_11422;
assign x_11424 = x_176 & x_177;
assign x_11425 = x_179 & x_180;
assign x_11426 = x_178 & x_11425;
assign x_11427 = x_11424 & x_11426;
assign x_11428 = x_182 & x_183;
assign x_11429 = x_181 & x_11428;
assign x_11430 = x_185 & x_186;
assign x_11431 = x_184 & x_11430;
assign x_11432 = x_11429 & x_11431;
assign x_11433 = x_11427 & x_11432;
assign x_11434 = x_187 & x_188;
assign x_11435 = x_190 & x_191;
assign x_11436 = x_189 & x_11435;
assign x_11437 = x_11434 & x_11436;
assign x_11438 = x_193 & x_194;
assign x_11439 = x_192 & x_11438;
assign x_11440 = x_196 & x_197;
assign x_11441 = x_195 & x_11440;
assign x_11442 = x_11439 & x_11441;
assign x_11443 = x_11437 & x_11442;
assign x_11444 = x_11433 & x_11443;
assign x_11445 = x_198 & x_199;
assign x_11446 = x_201 & x_202;
assign x_11447 = x_200 & x_11446;
assign x_11448 = x_11445 & x_11447;
assign x_11449 = x_204 & x_205;
assign x_11450 = x_203 & x_11449;
assign x_11451 = x_207 & x_208;
assign x_11452 = x_206 & x_11451;
assign x_11453 = x_11450 & x_11452;
assign x_11454 = x_11448 & x_11453;
assign x_11455 = x_209 & x_210;
assign x_11456 = x_212 & x_213;
assign x_11457 = x_211 & x_11456;
assign x_11458 = x_11455 & x_11457;
assign x_11459 = x_215 & x_216;
assign x_11460 = x_214 & x_11459;
assign x_11461 = x_218 & x_219;
assign x_11462 = x_217 & x_11461;
assign x_11463 = x_11460 & x_11462;
assign x_11464 = x_11458 & x_11463;
assign x_11465 = x_11454 & x_11464;
assign x_11466 = x_11444 & x_11465;
assign x_11467 = x_220 & x_221;
assign x_11468 = x_223 & x_224;
assign x_11469 = x_222 & x_11468;
assign x_11470 = x_11467 & x_11469;
assign x_11471 = x_226 & x_227;
assign x_11472 = x_225 & x_11471;
assign x_11473 = x_229 & x_230;
assign x_11474 = x_228 & x_11473;
assign x_11475 = x_11472 & x_11474;
assign x_11476 = x_11470 & x_11475;
assign x_11477 = x_231 & x_232;
assign x_11478 = x_234 & x_235;
assign x_11479 = x_233 & x_11478;
assign x_11480 = x_11477 & x_11479;
assign x_11481 = x_237 & x_238;
assign x_11482 = x_236 & x_11481;
assign x_11483 = x_240 & x_241;
assign x_11484 = x_239 & x_11483;
assign x_11485 = x_11482 & x_11484;
assign x_11486 = x_11480 & x_11485;
assign x_11487 = x_11476 & x_11486;
assign x_11488 = x_242 & x_243;
assign x_11489 = x_245 & x_246;
assign x_11490 = x_244 & x_11489;
assign x_11491 = x_11488 & x_11490;
assign x_11492 = x_248 & x_249;
assign x_11493 = x_247 & x_11492;
assign x_11494 = x_251 & x_252;
assign x_11495 = x_250 & x_11494;
assign x_11496 = x_11493 & x_11495;
assign x_11497 = x_11491 & x_11496;
assign x_11498 = x_253 & x_254;
assign x_11499 = x_256 & x_257;
assign x_11500 = x_255 & x_11499;
assign x_11501 = x_11498 & x_11500;
assign x_11502 = x_259 & x_260;
assign x_11503 = x_258 & x_11502;
assign x_11504 = x_262 & x_263;
assign x_11505 = x_261 & x_11504;
assign x_11506 = x_11503 & x_11505;
assign x_11507 = x_11501 & x_11506;
assign x_11508 = x_11497 & x_11507;
assign x_11509 = x_11487 & x_11508;
assign x_11510 = x_11466 & x_11509;
assign x_11511 = x_264 & x_265;
assign x_11512 = x_267 & x_268;
assign x_11513 = x_266 & x_11512;
assign x_11514 = x_11511 & x_11513;
assign x_11515 = x_270 & x_271;
assign x_11516 = x_269 & x_11515;
assign x_11517 = x_273 & x_274;
assign x_11518 = x_272 & x_11517;
assign x_11519 = x_11516 & x_11518;
assign x_11520 = x_11514 & x_11519;
assign x_11521 = x_275 & x_276;
assign x_11522 = x_278 & x_279;
assign x_11523 = x_277 & x_11522;
assign x_11524 = x_11521 & x_11523;
assign x_11525 = x_281 & x_282;
assign x_11526 = x_280 & x_11525;
assign x_11527 = x_284 & x_285;
assign x_11528 = x_283 & x_11527;
assign x_11529 = x_11526 & x_11528;
assign x_11530 = x_11524 & x_11529;
assign x_11531 = x_11520 & x_11530;
assign x_11532 = x_286 & x_287;
assign x_11533 = x_289 & x_290;
assign x_11534 = x_288 & x_11533;
assign x_11535 = x_11532 & x_11534;
assign x_11536 = x_292 & x_293;
assign x_11537 = x_291 & x_11536;
assign x_11538 = x_295 & x_296;
assign x_11539 = x_294 & x_11538;
assign x_11540 = x_11537 & x_11539;
assign x_11541 = x_11535 & x_11540;
assign x_11542 = x_297 & x_298;
assign x_11543 = x_300 & x_301;
assign x_11544 = x_299 & x_11543;
assign x_11545 = x_11542 & x_11544;
assign x_11546 = x_303 & x_304;
assign x_11547 = x_302 & x_11546;
assign x_11548 = x_306 & x_307;
assign x_11549 = x_305 & x_11548;
assign x_11550 = x_11547 & x_11549;
assign x_11551 = x_11545 & x_11550;
assign x_11552 = x_11541 & x_11551;
assign x_11553 = x_11531 & x_11552;
assign x_11554 = x_308 & x_309;
assign x_11555 = x_311 & x_312;
assign x_11556 = x_310 & x_11555;
assign x_11557 = x_11554 & x_11556;
assign x_11558 = x_314 & x_315;
assign x_11559 = x_313 & x_11558;
assign x_11560 = x_317 & x_318;
assign x_11561 = x_316 & x_11560;
assign x_11562 = x_11559 & x_11561;
assign x_11563 = x_11557 & x_11562;
assign x_11564 = x_319 & x_320;
assign x_11565 = x_322 & x_323;
assign x_11566 = x_321 & x_11565;
assign x_11567 = x_11564 & x_11566;
assign x_11568 = x_325 & x_326;
assign x_11569 = x_324 & x_11568;
assign x_11570 = x_328 & x_329;
assign x_11571 = x_327 & x_11570;
assign x_11572 = x_11569 & x_11571;
assign x_11573 = x_11567 & x_11572;
assign x_11574 = x_11563 & x_11573;
assign x_11575 = x_330 & x_331;
assign x_11576 = x_333 & x_334;
assign x_11577 = x_332 & x_11576;
assign x_11578 = x_11575 & x_11577;
assign x_11579 = x_336 & x_337;
assign x_11580 = x_335 & x_11579;
assign x_11581 = x_339 & x_340;
assign x_11582 = x_338 & x_11581;
assign x_11583 = x_11580 & x_11582;
assign x_11584 = x_11578 & x_11583;
assign x_11585 = x_341 & x_342;
assign x_11586 = x_344 & x_345;
assign x_11587 = x_343 & x_11586;
assign x_11588 = x_11585 & x_11587;
assign x_11589 = x_347 & x_348;
assign x_11590 = x_346 & x_11589;
assign x_11591 = x_350 & x_351;
assign x_11592 = x_349 & x_11591;
assign x_11593 = x_11590 & x_11592;
assign x_11594 = x_11588 & x_11593;
assign x_11595 = x_11584 & x_11594;
assign x_11596 = x_11574 & x_11595;
assign x_11597 = x_11553 & x_11596;
assign x_11598 = x_11510 & x_11597;
assign x_11599 = x_11423 & x_11598;
assign x_11600 = x_352 & x_353;
assign x_11601 = x_355 & x_356;
assign x_11602 = x_354 & x_11601;
assign x_11603 = x_11600 & x_11602;
assign x_11604 = x_358 & x_359;
assign x_11605 = x_357 & x_11604;
assign x_11606 = x_361 & x_362;
assign x_11607 = x_360 & x_11606;
assign x_11608 = x_11605 & x_11607;
assign x_11609 = x_11603 & x_11608;
assign x_11610 = x_363 & x_364;
assign x_11611 = x_366 & x_367;
assign x_11612 = x_365 & x_11611;
assign x_11613 = x_11610 & x_11612;
assign x_11614 = x_369 & x_370;
assign x_11615 = x_368 & x_11614;
assign x_11616 = x_372 & x_373;
assign x_11617 = x_371 & x_11616;
assign x_11618 = x_11615 & x_11617;
assign x_11619 = x_11613 & x_11618;
assign x_11620 = x_11609 & x_11619;
assign x_11621 = x_374 & x_375;
assign x_11622 = x_377 & x_378;
assign x_11623 = x_376 & x_11622;
assign x_11624 = x_11621 & x_11623;
assign x_11625 = x_380 & x_381;
assign x_11626 = x_379 & x_11625;
assign x_11627 = x_383 & x_384;
assign x_11628 = x_382 & x_11627;
assign x_11629 = x_11626 & x_11628;
assign x_11630 = x_11624 & x_11629;
assign x_11631 = x_385 & x_386;
assign x_11632 = x_388 & x_389;
assign x_11633 = x_387 & x_11632;
assign x_11634 = x_11631 & x_11633;
assign x_11635 = x_391 & x_392;
assign x_11636 = x_390 & x_11635;
assign x_11637 = x_394 & x_395;
assign x_11638 = x_393 & x_11637;
assign x_11639 = x_11636 & x_11638;
assign x_11640 = x_11634 & x_11639;
assign x_11641 = x_11630 & x_11640;
assign x_11642 = x_11620 & x_11641;
assign x_11643 = x_396 & x_397;
assign x_11644 = x_399 & x_400;
assign x_11645 = x_398 & x_11644;
assign x_11646 = x_11643 & x_11645;
assign x_11647 = x_402 & x_403;
assign x_11648 = x_401 & x_11647;
assign x_11649 = x_405 & x_406;
assign x_11650 = x_404 & x_11649;
assign x_11651 = x_11648 & x_11650;
assign x_11652 = x_11646 & x_11651;
assign x_11653 = x_407 & x_408;
assign x_11654 = x_410 & x_411;
assign x_11655 = x_409 & x_11654;
assign x_11656 = x_11653 & x_11655;
assign x_11657 = x_413 & x_414;
assign x_11658 = x_412 & x_11657;
assign x_11659 = x_416 & x_417;
assign x_11660 = x_415 & x_11659;
assign x_11661 = x_11658 & x_11660;
assign x_11662 = x_11656 & x_11661;
assign x_11663 = x_11652 & x_11662;
assign x_11664 = x_418 & x_419;
assign x_11665 = x_421 & x_422;
assign x_11666 = x_420 & x_11665;
assign x_11667 = x_11664 & x_11666;
assign x_11668 = x_424 & x_425;
assign x_11669 = x_423 & x_11668;
assign x_11670 = x_427 & x_428;
assign x_11671 = x_426 & x_11670;
assign x_11672 = x_11669 & x_11671;
assign x_11673 = x_11667 & x_11672;
assign x_11674 = x_429 & x_430;
assign x_11675 = x_432 & x_433;
assign x_11676 = x_431 & x_11675;
assign x_11677 = x_11674 & x_11676;
assign x_11678 = x_435 & x_436;
assign x_11679 = x_434 & x_11678;
assign x_11680 = x_438 & x_439;
assign x_11681 = x_437 & x_11680;
assign x_11682 = x_11679 & x_11681;
assign x_11683 = x_11677 & x_11682;
assign x_11684 = x_11673 & x_11683;
assign x_11685 = x_11663 & x_11684;
assign x_11686 = x_11642 & x_11685;
assign x_11687 = x_440 & x_441;
assign x_11688 = x_443 & x_444;
assign x_11689 = x_442 & x_11688;
assign x_11690 = x_11687 & x_11689;
assign x_11691 = x_446 & x_447;
assign x_11692 = x_445 & x_11691;
assign x_11693 = x_449 & x_450;
assign x_11694 = x_448 & x_11693;
assign x_11695 = x_11692 & x_11694;
assign x_11696 = x_11690 & x_11695;
assign x_11697 = x_451 & x_452;
assign x_11698 = x_454 & x_455;
assign x_11699 = x_453 & x_11698;
assign x_11700 = x_11697 & x_11699;
assign x_11701 = x_457 & x_458;
assign x_11702 = x_456 & x_11701;
assign x_11703 = x_460 & x_461;
assign x_11704 = x_459 & x_11703;
assign x_11705 = x_11702 & x_11704;
assign x_11706 = x_11700 & x_11705;
assign x_11707 = x_11696 & x_11706;
assign x_11708 = x_462 & x_463;
assign x_11709 = x_465 & x_466;
assign x_11710 = x_464 & x_11709;
assign x_11711 = x_11708 & x_11710;
assign x_11712 = x_468 & x_469;
assign x_11713 = x_467 & x_11712;
assign x_11714 = x_471 & x_472;
assign x_11715 = x_470 & x_11714;
assign x_11716 = x_11713 & x_11715;
assign x_11717 = x_11711 & x_11716;
assign x_11718 = x_473 & x_474;
assign x_11719 = x_476 & x_477;
assign x_11720 = x_475 & x_11719;
assign x_11721 = x_11718 & x_11720;
assign x_11722 = x_479 & x_480;
assign x_11723 = x_478 & x_11722;
assign x_11724 = x_482 & x_483;
assign x_11725 = x_481 & x_11724;
assign x_11726 = x_11723 & x_11725;
assign x_11727 = x_11721 & x_11726;
assign x_11728 = x_11717 & x_11727;
assign x_11729 = x_11707 & x_11728;
assign x_11730 = x_484 & x_485;
assign x_11731 = x_487 & x_488;
assign x_11732 = x_486 & x_11731;
assign x_11733 = x_11730 & x_11732;
assign x_11734 = x_490 & x_491;
assign x_11735 = x_489 & x_11734;
assign x_11736 = x_493 & x_494;
assign x_11737 = x_492 & x_11736;
assign x_11738 = x_11735 & x_11737;
assign x_11739 = x_11733 & x_11738;
assign x_11740 = x_495 & x_496;
assign x_11741 = x_498 & x_499;
assign x_11742 = x_497 & x_11741;
assign x_11743 = x_11740 & x_11742;
assign x_11744 = x_501 & x_502;
assign x_11745 = x_500 & x_11744;
assign x_11746 = x_504 & x_505;
assign x_11747 = x_503 & x_11746;
assign x_11748 = x_11745 & x_11747;
assign x_11749 = x_11743 & x_11748;
assign x_11750 = x_11739 & x_11749;
assign x_11751 = x_506 & x_507;
assign x_11752 = x_509 & x_510;
assign x_11753 = x_508 & x_11752;
assign x_11754 = x_11751 & x_11753;
assign x_11755 = x_512 & x_513;
assign x_11756 = x_511 & x_11755;
assign x_11757 = x_515 & x_516;
assign x_11758 = x_514 & x_11757;
assign x_11759 = x_11756 & x_11758;
assign x_11760 = x_11754 & x_11759;
assign x_11761 = x_517 & x_518;
assign x_11762 = x_520 & x_521;
assign x_11763 = x_519 & x_11762;
assign x_11764 = x_11761 & x_11763;
assign x_11765 = x_523 & x_524;
assign x_11766 = x_522 & x_11765;
assign x_11767 = x_526 & x_527;
assign x_11768 = x_525 & x_11767;
assign x_11769 = x_11766 & x_11768;
assign x_11770 = x_11764 & x_11769;
assign x_11771 = x_11760 & x_11770;
assign x_11772 = x_11750 & x_11771;
assign x_11773 = x_11729 & x_11772;
assign x_11774 = x_11686 & x_11773;
assign x_11775 = x_528 & x_529;
assign x_11776 = x_531 & x_532;
assign x_11777 = x_530 & x_11776;
assign x_11778 = x_11775 & x_11777;
assign x_11779 = x_534 & x_535;
assign x_11780 = x_533 & x_11779;
assign x_11781 = x_537 & x_538;
assign x_11782 = x_536 & x_11781;
assign x_11783 = x_11780 & x_11782;
assign x_11784 = x_11778 & x_11783;
assign x_11785 = x_539 & x_540;
assign x_11786 = x_542 & x_543;
assign x_11787 = x_541 & x_11786;
assign x_11788 = x_11785 & x_11787;
assign x_11789 = x_545 & x_546;
assign x_11790 = x_544 & x_11789;
assign x_11791 = x_548 & x_549;
assign x_11792 = x_547 & x_11791;
assign x_11793 = x_11790 & x_11792;
assign x_11794 = x_11788 & x_11793;
assign x_11795 = x_11784 & x_11794;
assign x_11796 = x_550 & x_551;
assign x_11797 = x_553 & x_554;
assign x_11798 = x_552 & x_11797;
assign x_11799 = x_11796 & x_11798;
assign x_11800 = x_556 & x_557;
assign x_11801 = x_555 & x_11800;
assign x_11802 = x_559 & x_560;
assign x_11803 = x_558 & x_11802;
assign x_11804 = x_11801 & x_11803;
assign x_11805 = x_11799 & x_11804;
assign x_11806 = x_561 & x_562;
assign x_11807 = x_564 & x_565;
assign x_11808 = x_563 & x_11807;
assign x_11809 = x_11806 & x_11808;
assign x_11810 = x_567 & x_568;
assign x_11811 = x_566 & x_11810;
assign x_11812 = x_570 & x_571;
assign x_11813 = x_569 & x_11812;
assign x_11814 = x_11811 & x_11813;
assign x_11815 = x_11809 & x_11814;
assign x_11816 = x_11805 & x_11815;
assign x_11817 = x_11795 & x_11816;
assign x_11818 = x_572 & x_573;
assign x_11819 = x_575 & x_576;
assign x_11820 = x_574 & x_11819;
assign x_11821 = x_11818 & x_11820;
assign x_11822 = x_578 & x_579;
assign x_11823 = x_577 & x_11822;
assign x_11824 = x_581 & x_582;
assign x_11825 = x_580 & x_11824;
assign x_11826 = x_11823 & x_11825;
assign x_11827 = x_11821 & x_11826;
assign x_11828 = x_583 & x_584;
assign x_11829 = x_586 & x_587;
assign x_11830 = x_585 & x_11829;
assign x_11831 = x_11828 & x_11830;
assign x_11832 = x_589 & x_590;
assign x_11833 = x_588 & x_11832;
assign x_11834 = x_592 & x_593;
assign x_11835 = x_591 & x_11834;
assign x_11836 = x_11833 & x_11835;
assign x_11837 = x_11831 & x_11836;
assign x_11838 = x_11827 & x_11837;
assign x_11839 = x_594 & x_595;
assign x_11840 = x_597 & x_598;
assign x_11841 = x_596 & x_11840;
assign x_11842 = x_11839 & x_11841;
assign x_11843 = x_600 & x_601;
assign x_11844 = x_599 & x_11843;
assign x_11845 = x_603 & x_604;
assign x_11846 = x_602 & x_11845;
assign x_11847 = x_11844 & x_11846;
assign x_11848 = x_11842 & x_11847;
assign x_11849 = x_605 & x_606;
assign x_11850 = x_608 & x_609;
assign x_11851 = x_607 & x_11850;
assign x_11852 = x_11849 & x_11851;
assign x_11853 = x_611 & x_612;
assign x_11854 = x_610 & x_11853;
assign x_11855 = x_614 & x_615;
assign x_11856 = x_613 & x_11855;
assign x_11857 = x_11854 & x_11856;
assign x_11858 = x_11852 & x_11857;
assign x_11859 = x_11848 & x_11858;
assign x_11860 = x_11838 & x_11859;
assign x_11861 = x_11817 & x_11860;
assign x_11862 = x_616 & x_617;
assign x_11863 = x_619 & x_620;
assign x_11864 = x_618 & x_11863;
assign x_11865 = x_11862 & x_11864;
assign x_11866 = x_622 & x_623;
assign x_11867 = x_621 & x_11866;
assign x_11868 = x_625 & x_626;
assign x_11869 = x_624 & x_11868;
assign x_11870 = x_11867 & x_11869;
assign x_11871 = x_11865 & x_11870;
assign x_11872 = x_627 & x_628;
assign x_11873 = x_630 & x_631;
assign x_11874 = x_629 & x_11873;
assign x_11875 = x_11872 & x_11874;
assign x_11876 = x_633 & x_634;
assign x_11877 = x_632 & x_11876;
assign x_11878 = x_636 & x_637;
assign x_11879 = x_635 & x_11878;
assign x_11880 = x_11877 & x_11879;
assign x_11881 = x_11875 & x_11880;
assign x_11882 = x_11871 & x_11881;
assign x_11883 = x_638 & x_639;
assign x_11884 = x_641 & x_642;
assign x_11885 = x_640 & x_11884;
assign x_11886 = x_11883 & x_11885;
assign x_11887 = x_644 & x_645;
assign x_11888 = x_643 & x_11887;
assign x_11889 = x_647 & x_648;
assign x_11890 = x_646 & x_11889;
assign x_11891 = x_11888 & x_11890;
assign x_11892 = x_11886 & x_11891;
assign x_11893 = x_649 & x_650;
assign x_11894 = x_652 & x_653;
assign x_11895 = x_651 & x_11894;
assign x_11896 = x_11893 & x_11895;
assign x_11897 = x_655 & x_656;
assign x_11898 = x_654 & x_11897;
assign x_11899 = x_658 & x_659;
assign x_11900 = x_657 & x_11899;
assign x_11901 = x_11898 & x_11900;
assign x_11902 = x_11896 & x_11901;
assign x_11903 = x_11892 & x_11902;
assign x_11904 = x_11882 & x_11903;
assign x_11905 = x_660 & x_661;
assign x_11906 = x_663 & x_664;
assign x_11907 = x_662 & x_11906;
assign x_11908 = x_11905 & x_11907;
assign x_11909 = x_666 & x_667;
assign x_11910 = x_665 & x_11909;
assign x_11911 = x_669 & x_670;
assign x_11912 = x_668 & x_11911;
assign x_11913 = x_11910 & x_11912;
assign x_11914 = x_11908 & x_11913;
assign x_11915 = x_671 & x_672;
assign x_11916 = x_674 & x_675;
assign x_11917 = x_673 & x_11916;
assign x_11918 = x_11915 & x_11917;
assign x_11919 = x_677 & x_678;
assign x_11920 = x_676 & x_11919;
assign x_11921 = x_680 & x_681;
assign x_11922 = x_679 & x_11921;
assign x_11923 = x_11920 & x_11922;
assign x_11924 = x_11918 & x_11923;
assign x_11925 = x_11914 & x_11924;
assign x_11926 = x_682 & x_683;
assign x_11927 = x_685 & x_686;
assign x_11928 = x_684 & x_11927;
assign x_11929 = x_11926 & x_11928;
assign x_11930 = x_688 & x_689;
assign x_11931 = x_687 & x_11930;
assign x_11932 = x_691 & x_692;
assign x_11933 = x_690 & x_11932;
assign x_11934 = x_11931 & x_11933;
assign x_11935 = x_11929 & x_11934;
assign x_11936 = x_693 & x_694;
assign x_11937 = x_696 & x_697;
assign x_11938 = x_695 & x_11937;
assign x_11939 = x_11936 & x_11938;
assign x_11940 = x_699 & x_700;
assign x_11941 = x_698 & x_11940;
assign x_11942 = x_702 & x_703;
assign x_11943 = x_701 & x_11942;
assign x_11944 = x_11941 & x_11943;
assign x_11945 = x_11939 & x_11944;
assign x_11946 = x_11935 & x_11945;
assign x_11947 = x_11925 & x_11946;
assign x_11948 = x_11904 & x_11947;
assign x_11949 = x_11861 & x_11948;
assign x_11950 = x_11774 & x_11949;
assign x_11951 = x_11599 & x_11950;
assign x_11952 = x_704 & x_705;
assign x_11953 = x_707 & x_708;
assign x_11954 = x_706 & x_11953;
assign x_11955 = x_11952 & x_11954;
assign x_11956 = x_709 & x_710;
assign x_11957 = x_712 & x_713;
assign x_11958 = x_711 & x_11957;
assign x_11959 = x_11956 & x_11958;
assign x_11960 = x_11955 & x_11959;
assign x_11961 = x_714 & x_715;
assign x_11962 = x_717 & x_718;
assign x_11963 = x_716 & x_11962;
assign x_11964 = x_11961 & x_11963;
assign x_11965 = x_720 & x_721;
assign x_11966 = x_719 & x_11965;
assign x_11967 = x_723 & x_724;
assign x_11968 = x_722 & x_11967;
assign x_11969 = x_11966 & x_11968;
assign x_11970 = x_11964 & x_11969;
assign x_11971 = x_11960 & x_11970;
assign x_11972 = x_725 & x_726;
assign x_11973 = x_728 & x_729;
assign x_11974 = x_727 & x_11973;
assign x_11975 = x_11972 & x_11974;
assign x_11976 = x_731 & x_732;
assign x_11977 = x_730 & x_11976;
assign x_11978 = x_734 & x_735;
assign x_11979 = x_733 & x_11978;
assign x_11980 = x_11977 & x_11979;
assign x_11981 = x_11975 & x_11980;
assign x_11982 = x_736 & x_737;
assign x_11983 = x_739 & x_740;
assign x_11984 = x_738 & x_11983;
assign x_11985 = x_11982 & x_11984;
assign x_11986 = x_742 & x_743;
assign x_11987 = x_741 & x_11986;
assign x_11988 = x_745 & x_746;
assign x_11989 = x_744 & x_11988;
assign x_11990 = x_11987 & x_11989;
assign x_11991 = x_11985 & x_11990;
assign x_11992 = x_11981 & x_11991;
assign x_11993 = x_11971 & x_11992;
assign x_11994 = x_747 & x_748;
assign x_11995 = x_750 & x_751;
assign x_11996 = x_749 & x_11995;
assign x_11997 = x_11994 & x_11996;
assign x_11998 = x_753 & x_754;
assign x_11999 = x_752 & x_11998;
assign x_12000 = x_756 & x_757;
assign x_12001 = x_755 & x_12000;
assign x_12002 = x_11999 & x_12001;
assign x_12003 = x_11997 & x_12002;
assign x_12004 = x_758 & x_759;
assign x_12005 = x_761 & x_762;
assign x_12006 = x_760 & x_12005;
assign x_12007 = x_12004 & x_12006;
assign x_12008 = x_764 & x_765;
assign x_12009 = x_763 & x_12008;
assign x_12010 = x_767 & x_768;
assign x_12011 = x_766 & x_12010;
assign x_12012 = x_12009 & x_12011;
assign x_12013 = x_12007 & x_12012;
assign x_12014 = x_12003 & x_12013;
assign x_12015 = x_769 & x_770;
assign x_12016 = x_772 & x_773;
assign x_12017 = x_771 & x_12016;
assign x_12018 = x_12015 & x_12017;
assign x_12019 = x_775 & x_776;
assign x_12020 = x_774 & x_12019;
assign x_12021 = x_778 & x_779;
assign x_12022 = x_777 & x_12021;
assign x_12023 = x_12020 & x_12022;
assign x_12024 = x_12018 & x_12023;
assign x_12025 = x_780 & x_781;
assign x_12026 = x_783 & x_784;
assign x_12027 = x_782 & x_12026;
assign x_12028 = x_12025 & x_12027;
assign x_12029 = x_786 & x_787;
assign x_12030 = x_785 & x_12029;
assign x_12031 = x_789 & x_790;
assign x_12032 = x_788 & x_12031;
assign x_12033 = x_12030 & x_12032;
assign x_12034 = x_12028 & x_12033;
assign x_12035 = x_12024 & x_12034;
assign x_12036 = x_12014 & x_12035;
assign x_12037 = x_11993 & x_12036;
assign x_12038 = x_791 & x_792;
assign x_12039 = x_794 & x_795;
assign x_12040 = x_793 & x_12039;
assign x_12041 = x_12038 & x_12040;
assign x_12042 = x_797 & x_798;
assign x_12043 = x_796 & x_12042;
assign x_12044 = x_800 & x_801;
assign x_12045 = x_799 & x_12044;
assign x_12046 = x_12043 & x_12045;
assign x_12047 = x_12041 & x_12046;
assign x_12048 = x_802 & x_803;
assign x_12049 = x_805 & x_806;
assign x_12050 = x_804 & x_12049;
assign x_12051 = x_12048 & x_12050;
assign x_12052 = x_808 & x_809;
assign x_12053 = x_807 & x_12052;
assign x_12054 = x_811 & x_812;
assign x_12055 = x_810 & x_12054;
assign x_12056 = x_12053 & x_12055;
assign x_12057 = x_12051 & x_12056;
assign x_12058 = x_12047 & x_12057;
assign x_12059 = x_813 & x_814;
assign x_12060 = x_816 & x_817;
assign x_12061 = x_815 & x_12060;
assign x_12062 = x_12059 & x_12061;
assign x_12063 = x_819 & x_820;
assign x_12064 = x_818 & x_12063;
assign x_12065 = x_822 & x_823;
assign x_12066 = x_821 & x_12065;
assign x_12067 = x_12064 & x_12066;
assign x_12068 = x_12062 & x_12067;
assign x_12069 = x_824 & x_825;
assign x_12070 = x_827 & x_828;
assign x_12071 = x_826 & x_12070;
assign x_12072 = x_12069 & x_12071;
assign x_12073 = x_830 & x_831;
assign x_12074 = x_829 & x_12073;
assign x_12075 = x_833 & x_834;
assign x_12076 = x_832 & x_12075;
assign x_12077 = x_12074 & x_12076;
assign x_12078 = x_12072 & x_12077;
assign x_12079 = x_12068 & x_12078;
assign x_12080 = x_12058 & x_12079;
assign x_12081 = x_835 & x_836;
assign x_12082 = x_838 & x_839;
assign x_12083 = x_837 & x_12082;
assign x_12084 = x_12081 & x_12083;
assign x_12085 = x_841 & x_842;
assign x_12086 = x_840 & x_12085;
assign x_12087 = x_844 & x_845;
assign x_12088 = x_843 & x_12087;
assign x_12089 = x_12086 & x_12088;
assign x_12090 = x_12084 & x_12089;
assign x_12091 = x_846 & x_847;
assign x_12092 = x_849 & x_850;
assign x_12093 = x_848 & x_12092;
assign x_12094 = x_12091 & x_12093;
assign x_12095 = x_852 & x_853;
assign x_12096 = x_851 & x_12095;
assign x_12097 = x_855 & x_856;
assign x_12098 = x_854 & x_12097;
assign x_12099 = x_12096 & x_12098;
assign x_12100 = x_12094 & x_12099;
assign x_12101 = x_12090 & x_12100;
assign x_12102 = x_857 & x_858;
assign x_12103 = x_860 & x_861;
assign x_12104 = x_859 & x_12103;
assign x_12105 = x_12102 & x_12104;
assign x_12106 = x_863 & x_864;
assign x_12107 = x_862 & x_12106;
assign x_12108 = x_866 & x_867;
assign x_12109 = x_865 & x_12108;
assign x_12110 = x_12107 & x_12109;
assign x_12111 = x_12105 & x_12110;
assign x_12112 = x_868 & x_869;
assign x_12113 = x_871 & x_872;
assign x_12114 = x_870 & x_12113;
assign x_12115 = x_12112 & x_12114;
assign x_12116 = x_874 & x_875;
assign x_12117 = x_873 & x_12116;
assign x_12118 = x_877 & x_878;
assign x_12119 = x_876 & x_12118;
assign x_12120 = x_12117 & x_12119;
assign x_12121 = x_12115 & x_12120;
assign x_12122 = x_12111 & x_12121;
assign x_12123 = x_12101 & x_12122;
assign x_12124 = x_12080 & x_12123;
assign x_12125 = x_12037 & x_12124;
assign x_12126 = x_879 & x_880;
assign x_12127 = x_882 & x_883;
assign x_12128 = x_881 & x_12127;
assign x_12129 = x_12126 & x_12128;
assign x_12130 = x_885 & x_886;
assign x_12131 = x_884 & x_12130;
assign x_12132 = x_888 & x_889;
assign x_12133 = x_887 & x_12132;
assign x_12134 = x_12131 & x_12133;
assign x_12135 = x_12129 & x_12134;
assign x_12136 = x_890 & x_891;
assign x_12137 = x_893 & x_894;
assign x_12138 = x_892 & x_12137;
assign x_12139 = x_12136 & x_12138;
assign x_12140 = x_896 & x_897;
assign x_12141 = x_895 & x_12140;
assign x_12142 = x_899 & x_900;
assign x_12143 = x_898 & x_12142;
assign x_12144 = x_12141 & x_12143;
assign x_12145 = x_12139 & x_12144;
assign x_12146 = x_12135 & x_12145;
assign x_12147 = x_901 & x_902;
assign x_12148 = x_904 & x_905;
assign x_12149 = x_903 & x_12148;
assign x_12150 = x_12147 & x_12149;
assign x_12151 = x_907 & x_908;
assign x_12152 = x_906 & x_12151;
assign x_12153 = x_910 & x_911;
assign x_12154 = x_909 & x_12153;
assign x_12155 = x_12152 & x_12154;
assign x_12156 = x_12150 & x_12155;
assign x_12157 = x_912 & x_913;
assign x_12158 = x_915 & x_916;
assign x_12159 = x_914 & x_12158;
assign x_12160 = x_12157 & x_12159;
assign x_12161 = x_918 & x_919;
assign x_12162 = x_917 & x_12161;
assign x_12163 = x_921 & x_922;
assign x_12164 = x_920 & x_12163;
assign x_12165 = x_12162 & x_12164;
assign x_12166 = x_12160 & x_12165;
assign x_12167 = x_12156 & x_12166;
assign x_12168 = x_12146 & x_12167;
assign x_12169 = x_923 & x_924;
assign x_12170 = x_926 & x_927;
assign x_12171 = x_925 & x_12170;
assign x_12172 = x_12169 & x_12171;
assign x_12173 = x_929 & x_930;
assign x_12174 = x_928 & x_12173;
assign x_12175 = x_932 & x_933;
assign x_12176 = x_931 & x_12175;
assign x_12177 = x_12174 & x_12176;
assign x_12178 = x_12172 & x_12177;
assign x_12179 = x_934 & x_935;
assign x_12180 = x_937 & x_938;
assign x_12181 = x_936 & x_12180;
assign x_12182 = x_12179 & x_12181;
assign x_12183 = x_940 & x_941;
assign x_12184 = x_939 & x_12183;
assign x_12185 = x_943 & x_944;
assign x_12186 = x_942 & x_12185;
assign x_12187 = x_12184 & x_12186;
assign x_12188 = x_12182 & x_12187;
assign x_12189 = x_12178 & x_12188;
assign x_12190 = x_945 & x_946;
assign x_12191 = x_948 & x_949;
assign x_12192 = x_947 & x_12191;
assign x_12193 = x_12190 & x_12192;
assign x_12194 = x_951 & x_952;
assign x_12195 = x_950 & x_12194;
assign x_12196 = x_954 & x_955;
assign x_12197 = x_953 & x_12196;
assign x_12198 = x_12195 & x_12197;
assign x_12199 = x_12193 & x_12198;
assign x_12200 = x_956 & x_957;
assign x_12201 = x_959 & x_960;
assign x_12202 = x_958 & x_12201;
assign x_12203 = x_12200 & x_12202;
assign x_12204 = x_962 & x_963;
assign x_12205 = x_961 & x_12204;
assign x_12206 = x_965 & x_966;
assign x_12207 = x_964 & x_12206;
assign x_12208 = x_12205 & x_12207;
assign x_12209 = x_12203 & x_12208;
assign x_12210 = x_12199 & x_12209;
assign x_12211 = x_12189 & x_12210;
assign x_12212 = x_12168 & x_12211;
assign x_12213 = x_967 & x_968;
assign x_12214 = x_970 & x_971;
assign x_12215 = x_969 & x_12214;
assign x_12216 = x_12213 & x_12215;
assign x_12217 = x_973 & x_974;
assign x_12218 = x_972 & x_12217;
assign x_12219 = x_976 & x_977;
assign x_12220 = x_975 & x_12219;
assign x_12221 = x_12218 & x_12220;
assign x_12222 = x_12216 & x_12221;
assign x_12223 = x_978 & x_979;
assign x_12224 = x_981 & x_982;
assign x_12225 = x_980 & x_12224;
assign x_12226 = x_12223 & x_12225;
assign x_12227 = x_984 & x_985;
assign x_12228 = x_983 & x_12227;
assign x_12229 = x_987 & x_988;
assign x_12230 = x_986 & x_12229;
assign x_12231 = x_12228 & x_12230;
assign x_12232 = x_12226 & x_12231;
assign x_12233 = x_12222 & x_12232;
assign x_12234 = x_989 & x_990;
assign x_12235 = x_992 & x_993;
assign x_12236 = x_991 & x_12235;
assign x_12237 = x_12234 & x_12236;
assign x_12238 = x_995 & x_996;
assign x_12239 = x_994 & x_12238;
assign x_12240 = x_998 & x_999;
assign x_12241 = x_997 & x_12240;
assign x_12242 = x_12239 & x_12241;
assign x_12243 = x_12237 & x_12242;
assign x_12244 = x_1000 & x_1001;
assign x_12245 = x_1003 & x_1004;
assign x_12246 = x_1002 & x_12245;
assign x_12247 = x_12244 & x_12246;
assign x_12248 = x_1006 & x_1007;
assign x_12249 = x_1005 & x_12248;
assign x_12250 = x_1009 & x_1010;
assign x_12251 = x_1008 & x_12250;
assign x_12252 = x_12249 & x_12251;
assign x_12253 = x_12247 & x_12252;
assign x_12254 = x_12243 & x_12253;
assign x_12255 = x_12233 & x_12254;
assign x_12256 = x_1011 & x_1012;
assign x_12257 = x_1014 & x_1015;
assign x_12258 = x_1013 & x_12257;
assign x_12259 = x_12256 & x_12258;
assign x_12260 = x_1017 & x_1018;
assign x_12261 = x_1016 & x_12260;
assign x_12262 = x_1020 & x_1021;
assign x_12263 = x_1019 & x_12262;
assign x_12264 = x_12261 & x_12263;
assign x_12265 = x_12259 & x_12264;
assign x_12266 = x_1022 & x_1023;
assign x_12267 = x_1025 & x_1026;
assign x_12268 = x_1024 & x_12267;
assign x_12269 = x_12266 & x_12268;
assign x_12270 = x_1028 & x_1029;
assign x_12271 = x_1027 & x_12270;
assign x_12272 = x_1031 & x_1032;
assign x_12273 = x_1030 & x_12272;
assign x_12274 = x_12271 & x_12273;
assign x_12275 = x_12269 & x_12274;
assign x_12276 = x_12265 & x_12275;
assign x_12277 = x_1033 & x_1034;
assign x_12278 = x_1036 & x_1037;
assign x_12279 = x_1035 & x_12278;
assign x_12280 = x_12277 & x_12279;
assign x_12281 = x_1039 & x_1040;
assign x_12282 = x_1038 & x_12281;
assign x_12283 = x_1042 & x_1043;
assign x_12284 = x_1041 & x_12283;
assign x_12285 = x_12282 & x_12284;
assign x_12286 = x_12280 & x_12285;
assign x_12287 = x_1044 & x_1045;
assign x_12288 = x_1047 & x_1048;
assign x_12289 = x_1046 & x_12288;
assign x_12290 = x_12287 & x_12289;
assign x_12291 = x_1050 & x_1051;
assign x_12292 = x_1049 & x_12291;
assign x_12293 = x_1053 & x_1054;
assign x_12294 = x_1052 & x_12293;
assign x_12295 = x_12292 & x_12294;
assign x_12296 = x_12290 & x_12295;
assign x_12297 = x_12286 & x_12296;
assign x_12298 = x_12276 & x_12297;
assign x_12299 = x_12255 & x_12298;
assign x_12300 = x_12212 & x_12299;
assign x_12301 = x_12125 & x_12300;
assign x_12302 = x_1055 & x_1056;
assign x_12303 = x_1058 & x_1059;
assign x_12304 = x_1057 & x_12303;
assign x_12305 = x_12302 & x_12304;
assign x_12306 = x_1061 & x_1062;
assign x_12307 = x_1060 & x_12306;
assign x_12308 = x_1064 & x_1065;
assign x_12309 = x_1063 & x_12308;
assign x_12310 = x_12307 & x_12309;
assign x_12311 = x_12305 & x_12310;
assign x_12312 = x_1066 & x_1067;
assign x_12313 = x_1069 & x_1070;
assign x_12314 = x_1068 & x_12313;
assign x_12315 = x_12312 & x_12314;
assign x_12316 = x_1072 & x_1073;
assign x_12317 = x_1071 & x_12316;
assign x_12318 = x_1075 & x_1076;
assign x_12319 = x_1074 & x_12318;
assign x_12320 = x_12317 & x_12319;
assign x_12321 = x_12315 & x_12320;
assign x_12322 = x_12311 & x_12321;
assign x_12323 = x_1077 & x_1078;
assign x_12324 = x_1080 & x_1081;
assign x_12325 = x_1079 & x_12324;
assign x_12326 = x_12323 & x_12325;
assign x_12327 = x_1083 & x_1084;
assign x_12328 = x_1082 & x_12327;
assign x_12329 = x_1086 & x_1087;
assign x_12330 = x_1085 & x_12329;
assign x_12331 = x_12328 & x_12330;
assign x_12332 = x_12326 & x_12331;
assign x_12333 = x_1088 & x_1089;
assign x_12334 = x_1091 & x_1092;
assign x_12335 = x_1090 & x_12334;
assign x_12336 = x_12333 & x_12335;
assign x_12337 = x_1094 & x_1095;
assign x_12338 = x_1093 & x_12337;
assign x_12339 = x_1097 & x_1098;
assign x_12340 = x_1096 & x_12339;
assign x_12341 = x_12338 & x_12340;
assign x_12342 = x_12336 & x_12341;
assign x_12343 = x_12332 & x_12342;
assign x_12344 = x_12322 & x_12343;
assign x_12345 = x_1099 & x_1100;
assign x_12346 = x_1102 & x_1103;
assign x_12347 = x_1101 & x_12346;
assign x_12348 = x_12345 & x_12347;
assign x_12349 = x_1105 & x_1106;
assign x_12350 = x_1104 & x_12349;
assign x_12351 = x_1108 & x_1109;
assign x_12352 = x_1107 & x_12351;
assign x_12353 = x_12350 & x_12352;
assign x_12354 = x_12348 & x_12353;
assign x_12355 = x_1110 & x_1111;
assign x_12356 = x_1113 & x_1114;
assign x_12357 = x_1112 & x_12356;
assign x_12358 = x_12355 & x_12357;
assign x_12359 = x_1116 & x_1117;
assign x_12360 = x_1115 & x_12359;
assign x_12361 = x_1119 & x_1120;
assign x_12362 = x_1118 & x_12361;
assign x_12363 = x_12360 & x_12362;
assign x_12364 = x_12358 & x_12363;
assign x_12365 = x_12354 & x_12364;
assign x_12366 = x_1121 & x_1122;
assign x_12367 = x_1124 & x_1125;
assign x_12368 = x_1123 & x_12367;
assign x_12369 = x_12366 & x_12368;
assign x_12370 = x_1127 & x_1128;
assign x_12371 = x_1126 & x_12370;
assign x_12372 = x_1130 & x_1131;
assign x_12373 = x_1129 & x_12372;
assign x_12374 = x_12371 & x_12373;
assign x_12375 = x_12369 & x_12374;
assign x_12376 = x_1132 & x_1133;
assign x_12377 = x_1135 & x_1136;
assign x_12378 = x_1134 & x_12377;
assign x_12379 = x_12376 & x_12378;
assign x_12380 = x_1138 & x_1139;
assign x_12381 = x_1137 & x_12380;
assign x_12382 = x_1141 & x_1142;
assign x_12383 = x_1140 & x_12382;
assign x_12384 = x_12381 & x_12383;
assign x_12385 = x_12379 & x_12384;
assign x_12386 = x_12375 & x_12385;
assign x_12387 = x_12365 & x_12386;
assign x_12388 = x_12344 & x_12387;
assign x_12389 = x_1143 & x_1144;
assign x_12390 = x_1146 & x_1147;
assign x_12391 = x_1145 & x_12390;
assign x_12392 = x_12389 & x_12391;
assign x_12393 = x_1149 & x_1150;
assign x_12394 = x_1148 & x_12393;
assign x_12395 = x_1152 & x_1153;
assign x_12396 = x_1151 & x_12395;
assign x_12397 = x_12394 & x_12396;
assign x_12398 = x_12392 & x_12397;
assign x_12399 = x_1154 & x_1155;
assign x_12400 = x_1157 & x_1158;
assign x_12401 = x_1156 & x_12400;
assign x_12402 = x_12399 & x_12401;
assign x_12403 = x_1160 & x_1161;
assign x_12404 = x_1159 & x_12403;
assign x_12405 = x_1163 & x_1164;
assign x_12406 = x_1162 & x_12405;
assign x_12407 = x_12404 & x_12406;
assign x_12408 = x_12402 & x_12407;
assign x_12409 = x_12398 & x_12408;
assign x_12410 = x_1165 & x_1166;
assign x_12411 = x_1168 & x_1169;
assign x_12412 = x_1167 & x_12411;
assign x_12413 = x_12410 & x_12412;
assign x_12414 = x_1171 & x_1172;
assign x_12415 = x_1170 & x_12414;
assign x_12416 = x_1174 & x_1175;
assign x_12417 = x_1173 & x_12416;
assign x_12418 = x_12415 & x_12417;
assign x_12419 = x_12413 & x_12418;
assign x_12420 = x_1176 & x_1177;
assign x_12421 = x_1179 & x_1180;
assign x_12422 = x_1178 & x_12421;
assign x_12423 = x_12420 & x_12422;
assign x_12424 = x_1182 & x_1183;
assign x_12425 = x_1181 & x_12424;
assign x_12426 = x_1185 & x_1186;
assign x_12427 = x_1184 & x_12426;
assign x_12428 = x_12425 & x_12427;
assign x_12429 = x_12423 & x_12428;
assign x_12430 = x_12419 & x_12429;
assign x_12431 = x_12409 & x_12430;
assign x_12432 = x_1187 & x_1188;
assign x_12433 = x_1190 & x_1191;
assign x_12434 = x_1189 & x_12433;
assign x_12435 = x_12432 & x_12434;
assign x_12436 = x_1193 & x_1194;
assign x_12437 = x_1192 & x_12436;
assign x_12438 = x_1196 & x_1197;
assign x_12439 = x_1195 & x_12438;
assign x_12440 = x_12437 & x_12439;
assign x_12441 = x_12435 & x_12440;
assign x_12442 = x_1198 & x_1199;
assign x_12443 = x_1201 & x_1202;
assign x_12444 = x_1200 & x_12443;
assign x_12445 = x_12442 & x_12444;
assign x_12446 = x_1204 & x_1205;
assign x_12447 = x_1203 & x_12446;
assign x_12448 = x_1207 & x_1208;
assign x_12449 = x_1206 & x_12448;
assign x_12450 = x_12447 & x_12449;
assign x_12451 = x_12445 & x_12450;
assign x_12452 = x_12441 & x_12451;
assign x_12453 = x_1209 & x_1210;
assign x_12454 = x_1212 & x_1213;
assign x_12455 = x_1211 & x_12454;
assign x_12456 = x_12453 & x_12455;
assign x_12457 = x_1215 & x_1216;
assign x_12458 = x_1214 & x_12457;
assign x_12459 = x_1218 & x_1219;
assign x_12460 = x_1217 & x_12459;
assign x_12461 = x_12458 & x_12460;
assign x_12462 = x_12456 & x_12461;
assign x_12463 = x_1220 & x_1221;
assign x_12464 = x_1223 & x_1224;
assign x_12465 = x_1222 & x_12464;
assign x_12466 = x_12463 & x_12465;
assign x_12467 = x_1226 & x_1227;
assign x_12468 = x_1225 & x_12467;
assign x_12469 = x_1229 & x_1230;
assign x_12470 = x_1228 & x_12469;
assign x_12471 = x_12468 & x_12470;
assign x_12472 = x_12466 & x_12471;
assign x_12473 = x_12462 & x_12472;
assign x_12474 = x_12452 & x_12473;
assign x_12475 = x_12431 & x_12474;
assign x_12476 = x_12388 & x_12475;
assign x_12477 = x_1231 & x_1232;
assign x_12478 = x_1234 & x_1235;
assign x_12479 = x_1233 & x_12478;
assign x_12480 = x_12477 & x_12479;
assign x_12481 = x_1237 & x_1238;
assign x_12482 = x_1236 & x_12481;
assign x_12483 = x_1240 & x_1241;
assign x_12484 = x_1239 & x_12483;
assign x_12485 = x_12482 & x_12484;
assign x_12486 = x_12480 & x_12485;
assign x_12487 = x_1242 & x_1243;
assign x_12488 = x_1245 & x_1246;
assign x_12489 = x_1244 & x_12488;
assign x_12490 = x_12487 & x_12489;
assign x_12491 = x_1248 & x_1249;
assign x_12492 = x_1247 & x_12491;
assign x_12493 = x_1251 & x_1252;
assign x_12494 = x_1250 & x_12493;
assign x_12495 = x_12492 & x_12494;
assign x_12496 = x_12490 & x_12495;
assign x_12497 = x_12486 & x_12496;
assign x_12498 = x_1253 & x_1254;
assign x_12499 = x_1256 & x_1257;
assign x_12500 = x_1255 & x_12499;
assign x_12501 = x_12498 & x_12500;
assign x_12502 = x_1259 & x_1260;
assign x_12503 = x_1258 & x_12502;
assign x_12504 = x_1262 & x_1263;
assign x_12505 = x_1261 & x_12504;
assign x_12506 = x_12503 & x_12505;
assign x_12507 = x_12501 & x_12506;
assign x_12508 = x_1264 & x_1265;
assign x_12509 = x_1267 & x_1268;
assign x_12510 = x_1266 & x_12509;
assign x_12511 = x_12508 & x_12510;
assign x_12512 = x_1270 & x_1271;
assign x_12513 = x_1269 & x_12512;
assign x_12514 = x_1273 & x_1274;
assign x_12515 = x_1272 & x_12514;
assign x_12516 = x_12513 & x_12515;
assign x_12517 = x_12511 & x_12516;
assign x_12518 = x_12507 & x_12517;
assign x_12519 = x_12497 & x_12518;
assign x_12520 = x_1275 & x_1276;
assign x_12521 = x_1278 & x_1279;
assign x_12522 = x_1277 & x_12521;
assign x_12523 = x_12520 & x_12522;
assign x_12524 = x_1281 & x_1282;
assign x_12525 = x_1280 & x_12524;
assign x_12526 = x_1284 & x_1285;
assign x_12527 = x_1283 & x_12526;
assign x_12528 = x_12525 & x_12527;
assign x_12529 = x_12523 & x_12528;
assign x_12530 = x_1286 & x_1287;
assign x_12531 = x_1289 & x_1290;
assign x_12532 = x_1288 & x_12531;
assign x_12533 = x_12530 & x_12532;
assign x_12534 = x_1292 & x_1293;
assign x_12535 = x_1291 & x_12534;
assign x_12536 = x_1295 & x_1296;
assign x_12537 = x_1294 & x_12536;
assign x_12538 = x_12535 & x_12537;
assign x_12539 = x_12533 & x_12538;
assign x_12540 = x_12529 & x_12539;
assign x_12541 = x_1297 & x_1298;
assign x_12542 = x_1300 & x_1301;
assign x_12543 = x_1299 & x_12542;
assign x_12544 = x_12541 & x_12543;
assign x_12545 = x_1303 & x_1304;
assign x_12546 = x_1302 & x_12545;
assign x_12547 = x_1306 & x_1307;
assign x_12548 = x_1305 & x_12547;
assign x_12549 = x_12546 & x_12548;
assign x_12550 = x_12544 & x_12549;
assign x_12551 = x_1308 & x_1309;
assign x_12552 = x_1311 & x_1312;
assign x_12553 = x_1310 & x_12552;
assign x_12554 = x_12551 & x_12553;
assign x_12555 = x_1314 & x_1315;
assign x_12556 = x_1313 & x_12555;
assign x_12557 = x_1317 & x_1318;
assign x_12558 = x_1316 & x_12557;
assign x_12559 = x_12556 & x_12558;
assign x_12560 = x_12554 & x_12559;
assign x_12561 = x_12550 & x_12560;
assign x_12562 = x_12540 & x_12561;
assign x_12563 = x_12519 & x_12562;
assign x_12564 = x_1319 & x_1320;
assign x_12565 = x_1322 & x_1323;
assign x_12566 = x_1321 & x_12565;
assign x_12567 = x_12564 & x_12566;
assign x_12568 = x_1325 & x_1326;
assign x_12569 = x_1324 & x_12568;
assign x_12570 = x_1328 & x_1329;
assign x_12571 = x_1327 & x_12570;
assign x_12572 = x_12569 & x_12571;
assign x_12573 = x_12567 & x_12572;
assign x_12574 = x_1330 & x_1331;
assign x_12575 = x_1333 & x_1334;
assign x_12576 = x_1332 & x_12575;
assign x_12577 = x_12574 & x_12576;
assign x_12578 = x_1336 & x_1337;
assign x_12579 = x_1335 & x_12578;
assign x_12580 = x_1339 & x_1340;
assign x_12581 = x_1338 & x_12580;
assign x_12582 = x_12579 & x_12581;
assign x_12583 = x_12577 & x_12582;
assign x_12584 = x_12573 & x_12583;
assign x_12585 = x_1341 & x_1342;
assign x_12586 = x_1344 & x_1345;
assign x_12587 = x_1343 & x_12586;
assign x_12588 = x_12585 & x_12587;
assign x_12589 = x_1347 & x_1348;
assign x_12590 = x_1346 & x_12589;
assign x_12591 = x_1350 & x_1351;
assign x_12592 = x_1349 & x_12591;
assign x_12593 = x_12590 & x_12592;
assign x_12594 = x_12588 & x_12593;
assign x_12595 = x_1352 & x_1353;
assign x_12596 = x_1355 & x_1356;
assign x_12597 = x_1354 & x_12596;
assign x_12598 = x_12595 & x_12597;
assign x_12599 = x_1358 & x_1359;
assign x_12600 = x_1357 & x_12599;
assign x_12601 = x_1361 & x_1362;
assign x_12602 = x_1360 & x_12601;
assign x_12603 = x_12600 & x_12602;
assign x_12604 = x_12598 & x_12603;
assign x_12605 = x_12594 & x_12604;
assign x_12606 = x_12584 & x_12605;
assign x_12607 = x_1363 & x_1364;
assign x_12608 = x_1366 & x_1367;
assign x_12609 = x_1365 & x_12608;
assign x_12610 = x_12607 & x_12609;
assign x_12611 = x_1369 & x_1370;
assign x_12612 = x_1368 & x_12611;
assign x_12613 = x_1372 & x_1373;
assign x_12614 = x_1371 & x_12613;
assign x_12615 = x_12612 & x_12614;
assign x_12616 = x_12610 & x_12615;
assign x_12617 = x_1374 & x_1375;
assign x_12618 = x_1377 & x_1378;
assign x_12619 = x_1376 & x_12618;
assign x_12620 = x_12617 & x_12619;
assign x_12621 = x_1380 & x_1381;
assign x_12622 = x_1379 & x_12621;
assign x_12623 = x_1383 & x_1384;
assign x_12624 = x_1382 & x_12623;
assign x_12625 = x_12622 & x_12624;
assign x_12626 = x_12620 & x_12625;
assign x_12627 = x_12616 & x_12626;
assign x_12628 = x_1385 & x_1386;
assign x_12629 = x_1388 & x_1389;
assign x_12630 = x_1387 & x_12629;
assign x_12631 = x_12628 & x_12630;
assign x_12632 = x_1391 & x_1392;
assign x_12633 = x_1390 & x_12632;
assign x_12634 = x_1394 & x_1395;
assign x_12635 = x_1393 & x_12634;
assign x_12636 = x_12633 & x_12635;
assign x_12637 = x_12631 & x_12636;
assign x_12638 = x_1396 & x_1397;
assign x_12639 = x_1399 & x_1400;
assign x_12640 = x_1398 & x_12639;
assign x_12641 = x_12638 & x_12640;
assign x_12642 = x_1402 & x_1403;
assign x_12643 = x_1401 & x_12642;
assign x_12644 = x_1405 & x_1406;
assign x_12645 = x_1404 & x_12644;
assign x_12646 = x_12643 & x_12645;
assign x_12647 = x_12641 & x_12646;
assign x_12648 = x_12637 & x_12647;
assign x_12649 = x_12627 & x_12648;
assign x_12650 = x_12606 & x_12649;
assign x_12651 = x_12563 & x_12650;
assign x_12652 = x_12476 & x_12651;
assign x_12653 = x_12301 & x_12652;
assign x_12654 = x_11951 & x_12653;
assign x_12655 = x_1407 & x_1408;
assign x_12656 = x_1410 & x_1411;
assign x_12657 = x_1409 & x_12656;
assign x_12658 = x_12655 & x_12657;
assign x_12659 = x_1412 & x_1413;
assign x_12660 = x_1415 & x_1416;
assign x_12661 = x_1414 & x_12660;
assign x_12662 = x_12659 & x_12661;
assign x_12663 = x_12658 & x_12662;
assign x_12664 = x_1417 & x_1418;
assign x_12665 = x_1420 & x_1421;
assign x_12666 = x_1419 & x_12665;
assign x_12667 = x_12664 & x_12666;
assign x_12668 = x_1423 & x_1424;
assign x_12669 = x_1422 & x_12668;
assign x_12670 = x_1426 & x_1427;
assign x_12671 = x_1425 & x_12670;
assign x_12672 = x_12669 & x_12671;
assign x_12673 = x_12667 & x_12672;
assign x_12674 = x_12663 & x_12673;
assign x_12675 = x_1428 & x_1429;
assign x_12676 = x_1431 & x_1432;
assign x_12677 = x_1430 & x_12676;
assign x_12678 = x_12675 & x_12677;
assign x_12679 = x_1434 & x_1435;
assign x_12680 = x_1433 & x_12679;
assign x_12681 = x_1437 & x_1438;
assign x_12682 = x_1436 & x_12681;
assign x_12683 = x_12680 & x_12682;
assign x_12684 = x_12678 & x_12683;
assign x_12685 = x_1439 & x_1440;
assign x_12686 = x_1442 & x_1443;
assign x_12687 = x_1441 & x_12686;
assign x_12688 = x_12685 & x_12687;
assign x_12689 = x_1445 & x_1446;
assign x_12690 = x_1444 & x_12689;
assign x_12691 = x_1448 & x_1449;
assign x_12692 = x_1447 & x_12691;
assign x_12693 = x_12690 & x_12692;
assign x_12694 = x_12688 & x_12693;
assign x_12695 = x_12684 & x_12694;
assign x_12696 = x_12674 & x_12695;
assign x_12697 = x_1450 & x_1451;
assign x_12698 = x_1453 & x_1454;
assign x_12699 = x_1452 & x_12698;
assign x_12700 = x_12697 & x_12699;
assign x_12701 = x_1456 & x_1457;
assign x_12702 = x_1455 & x_12701;
assign x_12703 = x_1459 & x_1460;
assign x_12704 = x_1458 & x_12703;
assign x_12705 = x_12702 & x_12704;
assign x_12706 = x_12700 & x_12705;
assign x_12707 = x_1461 & x_1462;
assign x_12708 = x_1464 & x_1465;
assign x_12709 = x_1463 & x_12708;
assign x_12710 = x_12707 & x_12709;
assign x_12711 = x_1467 & x_1468;
assign x_12712 = x_1466 & x_12711;
assign x_12713 = x_1470 & x_1471;
assign x_12714 = x_1469 & x_12713;
assign x_12715 = x_12712 & x_12714;
assign x_12716 = x_12710 & x_12715;
assign x_12717 = x_12706 & x_12716;
assign x_12718 = x_1472 & x_1473;
assign x_12719 = x_1475 & x_1476;
assign x_12720 = x_1474 & x_12719;
assign x_12721 = x_12718 & x_12720;
assign x_12722 = x_1478 & x_1479;
assign x_12723 = x_1477 & x_12722;
assign x_12724 = x_1481 & x_1482;
assign x_12725 = x_1480 & x_12724;
assign x_12726 = x_12723 & x_12725;
assign x_12727 = x_12721 & x_12726;
assign x_12728 = x_1483 & x_1484;
assign x_12729 = x_1486 & x_1487;
assign x_12730 = x_1485 & x_12729;
assign x_12731 = x_12728 & x_12730;
assign x_12732 = x_1489 & x_1490;
assign x_12733 = x_1488 & x_12732;
assign x_12734 = x_1492 & x_1493;
assign x_12735 = x_1491 & x_12734;
assign x_12736 = x_12733 & x_12735;
assign x_12737 = x_12731 & x_12736;
assign x_12738 = x_12727 & x_12737;
assign x_12739 = x_12717 & x_12738;
assign x_12740 = x_12696 & x_12739;
assign x_12741 = x_1494 & x_1495;
assign x_12742 = x_1497 & x_1498;
assign x_12743 = x_1496 & x_12742;
assign x_12744 = x_12741 & x_12743;
assign x_12745 = x_1500 & x_1501;
assign x_12746 = x_1499 & x_12745;
assign x_12747 = x_1503 & x_1504;
assign x_12748 = x_1502 & x_12747;
assign x_12749 = x_12746 & x_12748;
assign x_12750 = x_12744 & x_12749;
assign x_12751 = x_1505 & x_1506;
assign x_12752 = x_1508 & x_1509;
assign x_12753 = x_1507 & x_12752;
assign x_12754 = x_12751 & x_12753;
assign x_12755 = x_1511 & x_1512;
assign x_12756 = x_1510 & x_12755;
assign x_12757 = x_1514 & x_1515;
assign x_12758 = x_1513 & x_12757;
assign x_12759 = x_12756 & x_12758;
assign x_12760 = x_12754 & x_12759;
assign x_12761 = x_12750 & x_12760;
assign x_12762 = x_1516 & x_1517;
assign x_12763 = x_1519 & x_1520;
assign x_12764 = x_1518 & x_12763;
assign x_12765 = x_12762 & x_12764;
assign x_12766 = x_1522 & x_1523;
assign x_12767 = x_1521 & x_12766;
assign x_12768 = x_1525 & x_1526;
assign x_12769 = x_1524 & x_12768;
assign x_12770 = x_12767 & x_12769;
assign x_12771 = x_12765 & x_12770;
assign x_12772 = x_1527 & x_1528;
assign x_12773 = x_1530 & x_1531;
assign x_12774 = x_1529 & x_12773;
assign x_12775 = x_12772 & x_12774;
assign x_12776 = x_1533 & x_1534;
assign x_12777 = x_1532 & x_12776;
assign x_12778 = x_1536 & x_1537;
assign x_12779 = x_1535 & x_12778;
assign x_12780 = x_12777 & x_12779;
assign x_12781 = x_12775 & x_12780;
assign x_12782 = x_12771 & x_12781;
assign x_12783 = x_12761 & x_12782;
assign x_12784 = x_1538 & x_1539;
assign x_12785 = x_1541 & x_1542;
assign x_12786 = x_1540 & x_12785;
assign x_12787 = x_12784 & x_12786;
assign x_12788 = x_1544 & x_1545;
assign x_12789 = x_1543 & x_12788;
assign x_12790 = x_1547 & x_1548;
assign x_12791 = x_1546 & x_12790;
assign x_12792 = x_12789 & x_12791;
assign x_12793 = x_12787 & x_12792;
assign x_12794 = x_1549 & x_1550;
assign x_12795 = x_1552 & x_1553;
assign x_12796 = x_1551 & x_12795;
assign x_12797 = x_12794 & x_12796;
assign x_12798 = x_1555 & x_1556;
assign x_12799 = x_1554 & x_12798;
assign x_12800 = x_1558 & x_1559;
assign x_12801 = x_1557 & x_12800;
assign x_12802 = x_12799 & x_12801;
assign x_12803 = x_12797 & x_12802;
assign x_12804 = x_12793 & x_12803;
assign x_12805 = x_1560 & x_1561;
assign x_12806 = x_1563 & x_1564;
assign x_12807 = x_1562 & x_12806;
assign x_12808 = x_12805 & x_12807;
assign x_12809 = x_1566 & x_1567;
assign x_12810 = x_1565 & x_12809;
assign x_12811 = x_1569 & x_1570;
assign x_12812 = x_1568 & x_12811;
assign x_12813 = x_12810 & x_12812;
assign x_12814 = x_12808 & x_12813;
assign x_12815 = x_1571 & x_1572;
assign x_12816 = x_1574 & x_1575;
assign x_12817 = x_1573 & x_12816;
assign x_12818 = x_12815 & x_12817;
assign x_12819 = x_1577 & x_1578;
assign x_12820 = x_1576 & x_12819;
assign x_12821 = x_1580 & x_1581;
assign x_12822 = x_1579 & x_12821;
assign x_12823 = x_12820 & x_12822;
assign x_12824 = x_12818 & x_12823;
assign x_12825 = x_12814 & x_12824;
assign x_12826 = x_12804 & x_12825;
assign x_12827 = x_12783 & x_12826;
assign x_12828 = x_12740 & x_12827;
assign x_12829 = x_1582 & x_1583;
assign x_12830 = x_1585 & x_1586;
assign x_12831 = x_1584 & x_12830;
assign x_12832 = x_12829 & x_12831;
assign x_12833 = x_1588 & x_1589;
assign x_12834 = x_1587 & x_12833;
assign x_12835 = x_1591 & x_1592;
assign x_12836 = x_1590 & x_12835;
assign x_12837 = x_12834 & x_12836;
assign x_12838 = x_12832 & x_12837;
assign x_12839 = x_1593 & x_1594;
assign x_12840 = x_1596 & x_1597;
assign x_12841 = x_1595 & x_12840;
assign x_12842 = x_12839 & x_12841;
assign x_12843 = x_1599 & x_1600;
assign x_12844 = x_1598 & x_12843;
assign x_12845 = x_1602 & x_1603;
assign x_12846 = x_1601 & x_12845;
assign x_12847 = x_12844 & x_12846;
assign x_12848 = x_12842 & x_12847;
assign x_12849 = x_12838 & x_12848;
assign x_12850 = x_1604 & x_1605;
assign x_12851 = x_1607 & x_1608;
assign x_12852 = x_1606 & x_12851;
assign x_12853 = x_12850 & x_12852;
assign x_12854 = x_1610 & x_1611;
assign x_12855 = x_1609 & x_12854;
assign x_12856 = x_1613 & x_1614;
assign x_12857 = x_1612 & x_12856;
assign x_12858 = x_12855 & x_12857;
assign x_12859 = x_12853 & x_12858;
assign x_12860 = x_1615 & x_1616;
assign x_12861 = x_1618 & x_1619;
assign x_12862 = x_1617 & x_12861;
assign x_12863 = x_12860 & x_12862;
assign x_12864 = x_1621 & x_1622;
assign x_12865 = x_1620 & x_12864;
assign x_12866 = x_1624 & x_1625;
assign x_12867 = x_1623 & x_12866;
assign x_12868 = x_12865 & x_12867;
assign x_12869 = x_12863 & x_12868;
assign x_12870 = x_12859 & x_12869;
assign x_12871 = x_12849 & x_12870;
assign x_12872 = x_1626 & x_1627;
assign x_12873 = x_1629 & x_1630;
assign x_12874 = x_1628 & x_12873;
assign x_12875 = x_12872 & x_12874;
assign x_12876 = x_1632 & x_1633;
assign x_12877 = x_1631 & x_12876;
assign x_12878 = x_1635 & x_1636;
assign x_12879 = x_1634 & x_12878;
assign x_12880 = x_12877 & x_12879;
assign x_12881 = x_12875 & x_12880;
assign x_12882 = x_1637 & x_1638;
assign x_12883 = x_1640 & x_1641;
assign x_12884 = x_1639 & x_12883;
assign x_12885 = x_12882 & x_12884;
assign x_12886 = x_1643 & x_1644;
assign x_12887 = x_1642 & x_12886;
assign x_12888 = x_1646 & x_1647;
assign x_12889 = x_1645 & x_12888;
assign x_12890 = x_12887 & x_12889;
assign x_12891 = x_12885 & x_12890;
assign x_12892 = x_12881 & x_12891;
assign x_12893 = x_1648 & x_1649;
assign x_12894 = x_1651 & x_1652;
assign x_12895 = x_1650 & x_12894;
assign x_12896 = x_12893 & x_12895;
assign x_12897 = x_1654 & x_1655;
assign x_12898 = x_1653 & x_12897;
assign x_12899 = x_1657 & x_1658;
assign x_12900 = x_1656 & x_12899;
assign x_12901 = x_12898 & x_12900;
assign x_12902 = x_12896 & x_12901;
assign x_12903 = x_1659 & x_1660;
assign x_12904 = x_1662 & x_1663;
assign x_12905 = x_1661 & x_12904;
assign x_12906 = x_12903 & x_12905;
assign x_12907 = x_1665 & x_1666;
assign x_12908 = x_1664 & x_12907;
assign x_12909 = x_1668 & x_1669;
assign x_12910 = x_1667 & x_12909;
assign x_12911 = x_12908 & x_12910;
assign x_12912 = x_12906 & x_12911;
assign x_12913 = x_12902 & x_12912;
assign x_12914 = x_12892 & x_12913;
assign x_12915 = x_12871 & x_12914;
assign x_12916 = x_1670 & x_1671;
assign x_12917 = x_1673 & x_1674;
assign x_12918 = x_1672 & x_12917;
assign x_12919 = x_12916 & x_12918;
assign x_12920 = x_1676 & x_1677;
assign x_12921 = x_1675 & x_12920;
assign x_12922 = x_1679 & x_1680;
assign x_12923 = x_1678 & x_12922;
assign x_12924 = x_12921 & x_12923;
assign x_12925 = x_12919 & x_12924;
assign x_12926 = x_1681 & x_1682;
assign x_12927 = x_1684 & x_1685;
assign x_12928 = x_1683 & x_12927;
assign x_12929 = x_12926 & x_12928;
assign x_12930 = x_1687 & x_1688;
assign x_12931 = x_1686 & x_12930;
assign x_12932 = x_1690 & x_1691;
assign x_12933 = x_1689 & x_12932;
assign x_12934 = x_12931 & x_12933;
assign x_12935 = x_12929 & x_12934;
assign x_12936 = x_12925 & x_12935;
assign x_12937 = x_1692 & x_1693;
assign x_12938 = x_1695 & x_1696;
assign x_12939 = x_1694 & x_12938;
assign x_12940 = x_12937 & x_12939;
assign x_12941 = x_1698 & x_1699;
assign x_12942 = x_1697 & x_12941;
assign x_12943 = x_1701 & x_1702;
assign x_12944 = x_1700 & x_12943;
assign x_12945 = x_12942 & x_12944;
assign x_12946 = x_12940 & x_12945;
assign x_12947 = x_1703 & x_1704;
assign x_12948 = x_1706 & x_1707;
assign x_12949 = x_1705 & x_12948;
assign x_12950 = x_12947 & x_12949;
assign x_12951 = x_1709 & x_1710;
assign x_12952 = x_1708 & x_12951;
assign x_12953 = x_1712 & x_1713;
assign x_12954 = x_1711 & x_12953;
assign x_12955 = x_12952 & x_12954;
assign x_12956 = x_12950 & x_12955;
assign x_12957 = x_12946 & x_12956;
assign x_12958 = x_12936 & x_12957;
assign x_12959 = x_1714 & x_1715;
assign x_12960 = x_1717 & x_1718;
assign x_12961 = x_1716 & x_12960;
assign x_12962 = x_12959 & x_12961;
assign x_12963 = x_1720 & x_1721;
assign x_12964 = x_1719 & x_12963;
assign x_12965 = x_1723 & x_1724;
assign x_12966 = x_1722 & x_12965;
assign x_12967 = x_12964 & x_12966;
assign x_12968 = x_12962 & x_12967;
assign x_12969 = x_1725 & x_1726;
assign x_12970 = x_1728 & x_1729;
assign x_12971 = x_1727 & x_12970;
assign x_12972 = x_12969 & x_12971;
assign x_12973 = x_1731 & x_1732;
assign x_12974 = x_1730 & x_12973;
assign x_12975 = x_1734 & x_1735;
assign x_12976 = x_1733 & x_12975;
assign x_12977 = x_12974 & x_12976;
assign x_12978 = x_12972 & x_12977;
assign x_12979 = x_12968 & x_12978;
assign x_12980 = x_1736 & x_1737;
assign x_12981 = x_1739 & x_1740;
assign x_12982 = x_1738 & x_12981;
assign x_12983 = x_12980 & x_12982;
assign x_12984 = x_1742 & x_1743;
assign x_12985 = x_1741 & x_12984;
assign x_12986 = x_1745 & x_1746;
assign x_12987 = x_1744 & x_12986;
assign x_12988 = x_12985 & x_12987;
assign x_12989 = x_12983 & x_12988;
assign x_12990 = x_1747 & x_1748;
assign x_12991 = x_1750 & x_1751;
assign x_12992 = x_1749 & x_12991;
assign x_12993 = x_12990 & x_12992;
assign x_12994 = x_1753 & x_1754;
assign x_12995 = x_1752 & x_12994;
assign x_12996 = x_1756 & x_1757;
assign x_12997 = x_1755 & x_12996;
assign x_12998 = x_12995 & x_12997;
assign x_12999 = x_12993 & x_12998;
assign x_13000 = x_12989 & x_12999;
assign x_13001 = x_12979 & x_13000;
assign x_13002 = x_12958 & x_13001;
assign x_13003 = x_12915 & x_13002;
assign x_13004 = x_12828 & x_13003;
assign x_13005 = x_1758 & x_1759;
assign x_13006 = x_1761 & x_1762;
assign x_13007 = x_1760 & x_13006;
assign x_13008 = x_13005 & x_13007;
assign x_13009 = x_1764 & x_1765;
assign x_13010 = x_1763 & x_13009;
assign x_13011 = x_1767 & x_1768;
assign x_13012 = x_1766 & x_13011;
assign x_13013 = x_13010 & x_13012;
assign x_13014 = x_13008 & x_13013;
assign x_13015 = x_1769 & x_1770;
assign x_13016 = x_1772 & x_1773;
assign x_13017 = x_1771 & x_13016;
assign x_13018 = x_13015 & x_13017;
assign x_13019 = x_1775 & x_1776;
assign x_13020 = x_1774 & x_13019;
assign x_13021 = x_1778 & x_1779;
assign x_13022 = x_1777 & x_13021;
assign x_13023 = x_13020 & x_13022;
assign x_13024 = x_13018 & x_13023;
assign x_13025 = x_13014 & x_13024;
assign x_13026 = x_1780 & x_1781;
assign x_13027 = x_1783 & x_1784;
assign x_13028 = x_1782 & x_13027;
assign x_13029 = x_13026 & x_13028;
assign x_13030 = x_1786 & x_1787;
assign x_13031 = x_1785 & x_13030;
assign x_13032 = x_1789 & x_1790;
assign x_13033 = x_1788 & x_13032;
assign x_13034 = x_13031 & x_13033;
assign x_13035 = x_13029 & x_13034;
assign x_13036 = x_1791 & x_1792;
assign x_13037 = x_1794 & x_1795;
assign x_13038 = x_1793 & x_13037;
assign x_13039 = x_13036 & x_13038;
assign x_13040 = x_1797 & x_1798;
assign x_13041 = x_1796 & x_13040;
assign x_13042 = x_1800 & x_1801;
assign x_13043 = x_1799 & x_13042;
assign x_13044 = x_13041 & x_13043;
assign x_13045 = x_13039 & x_13044;
assign x_13046 = x_13035 & x_13045;
assign x_13047 = x_13025 & x_13046;
assign x_13048 = x_1802 & x_1803;
assign x_13049 = x_1805 & x_1806;
assign x_13050 = x_1804 & x_13049;
assign x_13051 = x_13048 & x_13050;
assign x_13052 = x_1808 & x_1809;
assign x_13053 = x_1807 & x_13052;
assign x_13054 = x_1811 & x_1812;
assign x_13055 = x_1810 & x_13054;
assign x_13056 = x_13053 & x_13055;
assign x_13057 = x_13051 & x_13056;
assign x_13058 = x_1813 & x_1814;
assign x_13059 = x_1816 & x_1817;
assign x_13060 = x_1815 & x_13059;
assign x_13061 = x_13058 & x_13060;
assign x_13062 = x_1819 & x_1820;
assign x_13063 = x_1818 & x_13062;
assign x_13064 = x_1822 & x_1823;
assign x_13065 = x_1821 & x_13064;
assign x_13066 = x_13063 & x_13065;
assign x_13067 = x_13061 & x_13066;
assign x_13068 = x_13057 & x_13067;
assign x_13069 = x_1824 & x_1825;
assign x_13070 = x_1827 & x_1828;
assign x_13071 = x_1826 & x_13070;
assign x_13072 = x_13069 & x_13071;
assign x_13073 = x_1830 & x_1831;
assign x_13074 = x_1829 & x_13073;
assign x_13075 = x_1833 & x_1834;
assign x_13076 = x_1832 & x_13075;
assign x_13077 = x_13074 & x_13076;
assign x_13078 = x_13072 & x_13077;
assign x_13079 = x_1835 & x_1836;
assign x_13080 = x_1838 & x_1839;
assign x_13081 = x_1837 & x_13080;
assign x_13082 = x_13079 & x_13081;
assign x_13083 = x_1841 & x_1842;
assign x_13084 = x_1840 & x_13083;
assign x_13085 = x_1844 & x_1845;
assign x_13086 = x_1843 & x_13085;
assign x_13087 = x_13084 & x_13086;
assign x_13088 = x_13082 & x_13087;
assign x_13089 = x_13078 & x_13088;
assign x_13090 = x_13068 & x_13089;
assign x_13091 = x_13047 & x_13090;
assign x_13092 = x_1846 & x_1847;
assign x_13093 = x_1849 & x_1850;
assign x_13094 = x_1848 & x_13093;
assign x_13095 = x_13092 & x_13094;
assign x_13096 = x_1852 & x_1853;
assign x_13097 = x_1851 & x_13096;
assign x_13098 = x_1855 & x_1856;
assign x_13099 = x_1854 & x_13098;
assign x_13100 = x_13097 & x_13099;
assign x_13101 = x_13095 & x_13100;
assign x_13102 = x_1857 & x_1858;
assign x_13103 = x_1860 & x_1861;
assign x_13104 = x_1859 & x_13103;
assign x_13105 = x_13102 & x_13104;
assign x_13106 = x_1863 & x_1864;
assign x_13107 = x_1862 & x_13106;
assign x_13108 = x_1866 & x_1867;
assign x_13109 = x_1865 & x_13108;
assign x_13110 = x_13107 & x_13109;
assign x_13111 = x_13105 & x_13110;
assign x_13112 = x_13101 & x_13111;
assign x_13113 = x_1868 & x_1869;
assign x_13114 = x_1871 & x_1872;
assign x_13115 = x_1870 & x_13114;
assign x_13116 = x_13113 & x_13115;
assign x_13117 = x_1874 & x_1875;
assign x_13118 = x_1873 & x_13117;
assign x_13119 = x_1877 & x_1878;
assign x_13120 = x_1876 & x_13119;
assign x_13121 = x_13118 & x_13120;
assign x_13122 = x_13116 & x_13121;
assign x_13123 = x_1879 & x_1880;
assign x_13124 = x_1882 & x_1883;
assign x_13125 = x_1881 & x_13124;
assign x_13126 = x_13123 & x_13125;
assign x_13127 = x_1885 & x_1886;
assign x_13128 = x_1884 & x_13127;
assign x_13129 = x_1888 & x_1889;
assign x_13130 = x_1887 & x_13129;
assign x_13131 = x_13128 & x_13130;
assign x_13132 = x_13126 & x_13131;
assign x_13133 = x_13122 & x_13132;
assign x_13134 = x_13112 & x_13133;
assign x_13135 = x_1890 & x_1891;
assign x_13136 = x_1893 & x_1894;
assign x_13137 = x_1892 & x_13136;
assign x_13138 = x_13135 & x_13137;
assign x_13139 = x_1896 & x_1897;
assign x_13140 = x_1895 & x_13139;
assign x_13141 = x_1899 & x_1900;
assign x_13142 = x_1898 & x_13141;
assign x_13143 = x_13140 & x_13142;
assign x_13144 = x_13138 & x_13143;
assign x_13145 = x_1901 & x_1902;
assign x_13146 = x_1904 & x_1905;
assign x_13147 = x_1903 & x_13146;
assign x_13148 = x_13145 & x_13147;
assign x_13149 = x_1907 & x_1908;
assign x_13150 = x_1906 & x_13149;
assign x_13151 = x_1910 & x_1911;
assign x_13152 = x_1909 & x_13151;
assign x_13153 = x_13150 & x_13152;
assign x_13154 = x_13148 & x_13153;
assign x_13155 = x_13144 & x_13154;
assign x_13156 = x_1912 & x_1913;
assign x_13157 = x_1915 & x_1916;
assign x_13158 = x_1914 & x_13157;
assign x_13159 = x_13156 & x_13158;
assign x_13160 = x_1918 & x_1919;
assign x_13161 = x_1917 & x_13160;
assign x_13162 = x_1921 & x_1922;
assign x_13163 = x_1920 & x_13162;
assign x_13164 = x_13161 & x_13163;
assign x_13165 = x_13159 & x_13164;
assign x_13166 = x_1923 & x_1924;
assign x_13167 = x_1926 & x_1927;
assign x_13168 = x_1925 & x_13167;
assign x_13169 = x_13166 & x_13168;
assign x_13170 = x_1929 & x_1930;
assign x_13171 = x_1928 & x_13170;
assign x_13172 = x_1932 & x_1933;
assign x_13173 = x_1931 & x_13172;
assign x_13174 = x_13171 & x_13173;
assign x_13175 = x_13169 & x_13174;
assign x_13176 = x_13165 & x_13175;
assign x_13177 = x_13155 & x_13176;
assign x_13178 = x_13134 & x_13177;
assign x_13179 = x_13091 & x_13178;
assign x_13180 = x_1934 & x_1935;
assign x_13181 = x_1937 & x_1938;
assign x_13182 = x_1936 & x_13181;
assign x_13183 = x_13180 & x_13182;
assign x_13184 = x_1940 & x_1941;
assign x_13185 = x_1939 & x_13184;
assign x_13186 = x_1943 & x_1944;
assign x_13187 = x_1942 & x_13186;
assign x_13188 = x_13185 & x_13187;
assign x_13189 = x_13183 & x_13188;
assign x_13190 = x_1945 & x_1946;
assign x_13191 = x_1948 & x_1949;
assign x_13192 = x_1947 & x_13191;
assign x_13193 = x_13190 & x_13192;
assign x_13194 = x_1951 & x_1952;
assign x_13195 = x_1950 & x_13194;
assign x_13196 = x_1954 & x_1955;
assign x_13197 = x_1953 & x_13196;
assign x_13198 = x_13195 & x_13197;
assign x_13199 = x_13193 & x_13198;
assign x_13200 = x_13189 & x_13199;
assign x_13201 = x_1956 & x_1957;
assign x_13202 = x_1959 & x_1960;
assign x_13203 = x_1958 & x_13202;
assign x_13204 = x_13201 & x_13203;
assign x_13205 = x_1962 & x_1963;
assign x_13206 = x_1961 & x_13205;
assign x_13207 = x_1965 & x_1966;
assign x_13208 = x_1964 & x_13207;
assign x_13209 = x_13206 & x_13208;
assign x_13210 = x_13204 & x_13209;
assign x_13211 = x_1967 & x_1968;
assign x_13212 = x_1970 & x_1971;
assign x_13213 = x_1969 & x_13212;
assign x_13214 = x_13211 & x_13213;
assign x_13215 = x_1973 & x_1974;
assign x_13216 = x_1972 & x_13215;
assign x_13217 = x_1976 & x_1977;
assign x_13218 = x_1975 & x_13217;
assign x_13219 = x_13216 & x_13218;
assign x_13220 = x_13214 & x_13219;
assign x_13221 = x_13210 & x_13220;
assign x_13222 = x_13200 & x_13221;
assign x_13223 = x_1978 & x_1979;
assign x_13224 = x_1981 & x_1982;
assign x_13225 = x_1980 & x_13224;
assign x_13226 = x_13223 & x_13225;
assign x_13227 = x_1984 & x_1985;
assign x_13228 = x_1983 & x_13227;
assign x_13229 = x_1987 & x_1988;
assign x_13230 = x_1986 & x_13229;
assign x_13231 = x_13228 & x_13230;
assign x_13232 = x_13226 & x_13231;
assign x_13233 = x_1989 & x_1990;
assign x_13234 = x_1992 & x_1993;
assign x_13235 = x_1991 & x_13234;
assign x_13236 = x_13233 & x_13235;
assign x_13237 = x_1995 & x_1996;
assign x_13238 = x_1994 & x_13237;
assign x_13239 = x_1998 & x_1999;
assign x_13240 = x_1997 & x_13239;
assign x_13241 = x_13238 & x_13240;
assign x_13242 = x_13236 & x_13241;
assign x_13243 = x_13232 & x_13242;
assign x_13244 = x_2000 & x_2001;
assign x_13245 = x_2003 & x_2004;
assign x_13246 = x_2002 & x_13245;
assign x_13247 = x_13244 & x_13246;
assign x_13248 = x_2006 & x_2007;
assign x_13249 = x_2005 & x_13248;
assign x_13250 = x_2009 & x_2010;
assign x_13251 = x_2008 & x_13250;
assign x_13252 = x_13249 & x_13251;
assign x_13253 = x_13247 & x_13252;
assign x_13254 = x_2011 & x_2012;
assign x_13255 = x_2014 & x_2015;
assign x_13256 = x_2013 & x_13255;
assign x_13257 = x_13254 & x_13256;
assign x_13258 = x_2017 & x_2018;
assign x_13259 = x_2016 & x_13258;
assign x_13260 = x_2020 & x_2021;
assign x_13261 = x_2019 & x_13260;
assign x_13262 = x_13259 & x_13261;
assign x_13263 = x_13257 & x_13262;
assign x_13264 = x_13253 & x_13263;
assign x_13265 = x_13243 & x_13264;
assign x_13266 = x_13222 & x_13265;
assign x_13267 = x_2022 & x_2023;
assign x_13268 = x_2025 & x_2026;
assign x_13269 = x_2024 & x_13268;
assign x_13270 = x_13267 & x_13269;
assign x_13271 = x_2028 & x_2029;
assign x_13272 = x_2027 & x_13271;
assign x_13273 = x_2031 & x_2032;
assign x_13274 = x_2030 & x_13273;
assign x_13275 = x_13272 & x_13274;
assign x_13276 = x_13270 & x_13275;
assign x_13277 = x_2033 & x_2034;
assign x_13278 = x_2036 & x_2037;
assign x_13279 = x_2035 & x_13278;
assign x_13280 = x_13277 & x_13279;
assign x_13281 = x_2039 & x_2040;
assign x_13282 = x_2038 & x_13281;
assign x_13283 = x_2042 & x_2043;
assign x_13284 = x_2041 & x_13283;
assign x_13285 = x_13282 & x_13284;
assign x_13286 = x_13280 & x_13285;
assign x_13287 = x_13276 & x_13286;
assign x_13288 = x_2044 & x_2045;
assign x_13289 = x_2047 & x_2048;
assign x_13290 = x_2046 & x_13289;
assign x_13291 = x_13288 & x_13290;
assign x_13292 = x_2050 & x_2051;
assign x_13293 = x_2049 & x_13292;
assign x_13294 = x_2053 & x_2054;
assign x_13295 = x_2052 & x_13294;
assign x_13296 = x_13293 & x_13295;
assign x_13297 = x_13291 & x_13296;
assign x_13298 = x_2055 & x_2056;
assign x_13299 = x_2058 & x_2059;
assign x_13300 = x_2057 & x_13299;
assign x_13301 = x_13298 & x_13300;
assign x_13302 = x_2061 & x_2062;
assign x_13303 = x_2060 & x_13302;
assign x_13304 = x_2064 & x_2065;
assign x_13305 = x_2063 & x_13304;
assign x_13306 = x_13303 & x_13305;
assign x_13307 = x_13301 & x_13306;
assign x_13308 = x_13297 & x_13307;
assign x_13309 = x_13287 & x_13308;
assign x_13310 = x_2066 & x_2067;
assign x_13311 = x_2069 & x_2070;
assign x_13312 = x_2068 & x_13311;
assign x_13313 = x_13310 & x_13312;
assign x_13314 = x_2072 & x_2073;
assign x_13315 = x_2071 & x_13314;
assign x_13316 = x_2075 & x_2076;
assign x_13317 = x_2074 & x_13316;
assign x_13318 = x_13315 & x_13317;
assign x_13319 = x_13313 & x_13318;
assign x_13320 = x_2077 & x_2078;
assign x_13321 = x_2080 & x_2081;
assign x_13322 = x_2079 & x_13321;
assign x_13323 = x_13320 & x_13322;
assign x_13324 = x_2083 & x_2084;
assign x_13325 = x_2082 & x_13324;
assign x_13326 = x_2086 & x_2087;
assign x_13327 = x_2085 & x_13326;
assign x_13328 = x_13325 & x_13327;
assign x_13329 = x_13323 & x_13328;
assign x_13330 = x_13319 & x_13329;
assign x_13331 = x_2088 & x_2089;
assign x_13332 = x_2091 & x_2092;
assign x_13333 = x_2090 & x_13332;
assign x_13334 = x_13331 & x_13333;
assign x_13335 = x_2094 & x_2095;
assign x_13336 = x_2093 & x_13335;
assign x_13337 = x_2097 & x_2098;
assign x_13338 = x_2096 & x_13337;
assign x_13339 = x_13336 & x_13338;
assign x_13340 = x_13334 & x_13339;
assign x_13341 = x_2099 & x_2100;
assign x_13342 = x_2102 & x_2103;
assign x_13343 = x_2101 & x_13342;
assign x_13344 = x_13341 & x_13343;
assign x_13345 = x_2105 & x_2106;
assign x_13346 = x_2104 & x_13345;
assign x_13347 = x_2108 & x_2109;
assign x_13348 = x_2107 & x_13347;
assign x_13349 = x_13346 & x_13348;
assign x_13350 = x_13344 & x_13349;
assign x_13351 = x_13340 & x_13350;
assign x_13352 = x_13330 & x_13351;
assign x_13353 = x_13309 & x_13352;
assign x_13354 = x_13266 & x_13353;
assign x_13355 = x_13179 & x_13354;
assign x_13356 = x_13004 & x_13355;
assign x_13357 = x_2110 & x_2111;
assign x_13358 = x_2113 & x_2114;
assign x_13359 = x_2112 & x_13358;
assign x_13360 = x_13357 & x_13359;
assign x_13361 = x_2115 & x_2116;
assign x_13362 = x_2118 & x_2119;
assign x_13363 = x_2117 & x_13362;
assign x_13364 = x_13361 & x_13363;
assign x_13365 = x_13360 & x_13364;
assign x_13366 = x_2120 & x_2121;
assign x_13367 = x_2123 & x_2124;
assign x_13368 = x_2122 & x_13367;
assign x_13369 = x_13366 & x_13368;
assign x_13370 = x_2126 & x_2127;
assign x_13371 = x_2125 & x_13370;
assign x_13372 = x_2129 & x_2130;
assign x_13373 = x_2128 & x_13372;
assign x_13374 = x_13371 & x_13373;
assign x_13375 = x_13369 & x_13374;
assign x_13376 = x_13365 & x_13375;
assign x_13377 = x_2131 & x_2132;
assign x_13378 = x_2134 & x_2135;
assign x_13379 = x_2133 & x_13378;
assign x_13380 = x_13377 & x_13379;
assign x_13381 = x_2137 & x_2138;
assign x_13382 = x_2136 & x_13381;
assign x_13383 = x_2140 & x_2141;
assign x_13384 = x_2139 & x_13383;
assign x_13385 = x_13382 & x_13384;
assign x_13386 = x_13380 & x_13385;
assign x_13387 = x_2142 & x_2143;
assign x_13388 = x_2145 & x_2146;
assign x_13389 = x_2144 & x_13388;
assign x_13390 = x_13387 & x_13389;
assign x_13391 = x_2148 & x_2149;
assign x_13392 = x_2147 & x_13391;
assign x_13393 = x_2151 & x_2152;
assign x_13394 = x_2150 & x_13393;
assign x_13395 = x_13392 & x_13394;
assign x_13396 = x_13390 & x_13395;
assign x_13397 = x_13386 & x_13396;
assign x_13398 = x_13376 & x_13397;
assign x_13399 = x_2153 & x_2154;
assign x_13400 = x_2156 & x_2157;
assign x_13401 = x_2155 & x_13400;
assign x_13402 = x_13399 & x_13401;
assign x_13403 = x_2159 & x_2160;
assign x_13404 = x_2158 & x_13403;
assign x_13405 = x_2162 & x_2163;
assign x_13406 = x_2161 & x_13405;
assign x_13407 = x_13404 & x_13406;
assign x_13408 = x_13402 & x_13407;
assign x_13409 = x_2164 & x_2165;
assign x_13410 = x_2167 & x_2168;
assign x_13411 = x_2166 & x_13410;
assign x_13412 = x_13409 & x_13411;
assign x_13413 = x_2170 & x_2171;
assign x_13414 = x_2169 & x_13413;
assign x_13415 = x_2173 & x_2174;
assign x_13416 = x_2172 & x_13415;
assign x_13417 = x_13414 & x_13416;
assign x_13418 = x_13412 & x_13417;
assign x_13419 = x_13408 & x_13418;
assign x_13420 = x_2175 & x_2176;
assign x_13421 = x_2178 & x_2179;
assign x_13422 = x_2177 & x_13421;
assign x_13423 = x_13420 & x_13422;
assign x_13424 = x_2181 & x_2182;
assign x_13425 = x_2180 & x_13424;
assign x_13426 = x_2184 & x_2185;
assign x_13427 = x_2183 & x_13426;
assign x_13428 = x_13425 & x_13427;
assign x_13429 = x_13423 & x_13428;
assign x_13430 = x_2186 & x_2187;
assign x_13431 = x_2189 & x_2190;
assign x_13432 = x_2188 & x_13431;
assign x_13433 = x_13430 & x_13432;
assign x_13434 = x_2192 & x_2193;
assign x_13435 = x_2191 & x_13434;
assign x_13436 = x_2195 & x_2196;
assign x_13437 = x_2194 & x_13436;
assign x_13438 = x_13435 & x_13437;
assign x_13439 = x_13433 & x_13438;
assign x_13440 = x_13429 & x_13439;
assign x_13441 = x_13419 & x_13440;
assign x_13442 = x_13398 & x_13441;
assign x_13443 = x_2197 & x_2198;
assign x_13444 = x_2200 & x_2201;
assign x_13445 = x_2199 & x_13444;
assign x_13446 = x_13443 & x_13445;
assign x_13447 = x_2203 & x_2204;
assign x_13448 = x_2202 & x_13447;
assign x_13449 = x_2206 & x_2207;
assign x_13450 = x_2205 & x_13449;
assign x_13451 = x_13448 & x_13450;
assign x_13452 = x_13446 & x_13451;
assign x_13453 = x_2208 & x_2209;
assign x_13454 = x_2211 & x_2212;
assign x_13455 = x_2210 & x_13454;
assign x_13456 = x_13453 & x_13455;
assign x_13457 = x_2214 & x_2215;
assign x_13458 = x_2213 & x_13457;
assign x_13459 = x_2217 & x_2218;
assign x_13460 = x_2216 & x_13459;
assign x_13461 = x_13458 & x_13460;
assign x_13462 = x_13456 & x_13461;
assign x_13463 = x_13452 & x_13462;
assign x_13464 = x_2219 & x_2220;
assign x_13465 = x_2222 & x_2223;
assign x_13466 = x_2221 & x_13465;
assign x_13467 = x_13464 & x_13466;
assign x_13468 = x_2225 & x_2226;
assign x_13469 = x_2224 & x_13468;
assign x_13470 = x_2228 & x_2229;
assign x_13471 = x_2227 & x_13470;
assign x_13472 = x_13469 & x_13471;
assign x_13473 = x_13467 & x_13472;
assign x_13474 = x_2230 & x_2231;
assign x_13475 = x_2233 & x_2234;
assign x_13476 = x_2232 & x_13475;
assign x_13477 = x_13474 & x_13476;
assign x_13478 = x_2236 & x_2237;
assign x_13479 = x_2235 & x_13478;
assign x_13480 = x_2239 & x_2240;
assign x_13481 = x_2238 & x_13480;
assign x_13482 = x_13479 & x_13481;
assign x_13483 = x_13477 & x_13482;
assign x_13484 = x_13473 & x_13483;
assign x_13485 = x_13463 & x_13484;
assign x_13486 = x_2241 & x_2242;
assign x_13487 = x_2244 & x_2245;
assign x_13488 = x_2243 & x_13487;
assign x_13489 = x_13486 & x_13488;
assign x_13490 = x_2247 & x_2248;
assign x_13491 = x_2246 & x_13490;
assign x_13492 = x_2250 & x_2251;
assign x_13493 = x_2249 & x_13492;
assign x_13494 = x_13491 & x_13493;
assign x_13495 = x_13489 & x_13494;
assign x_13496 = x_2252 & x_2253;
assign x_13497 = x_2255 & x_2256;
assign x_13498 = x_2254 & x_13497;
assign x_13499 = x_13496 & x_13498;
assign x_13500 = x_2258 & x_2259;
assign x_13501 = x_2257 & x_13500;
assign x_13502 = x_2261 & x_2262;
assign x_13503 = x_2260 & x_13502;
assign x_13504 = x_13501 & x_13503;
assign x_13505 = x_13499 & x_13504;
assign x_13506 = x_13495 & x_13505;
assign x_13507 = x_2263 & x_2264;
assign x_13508 = x_2266 & x_2267;
assign x_13509 = x_2265 & x_13508;
assign x_13510 = x_13507 & x_13509;
assign x_13511 = x_2269 & x_2270;
assign x_13512 = x_2268 & x_13511;
assign x_13513 = x_2272 & x_2273;
assign x_13514 = x_2271 & x_13513;
assign x_13515 = x_13512 & x_13514;
assign x_13516 = x_13510 & x_13515;
assign x_13517 = x_2274 & x_2275;
assign x_13518 = x_2277 & x_2278;
assign x_13519 = x_2276 & x_13518;
assign x_13520 = x_13517 & x_13519;
assign x_13521 = x_2280 & x_2281;
assign x_13522 = x_2279 & x_13521;
assign x_13523 = x_2283 & x_2284;
assign x_13524 = x_2282 & x_13523;
assign x_13525 = x_13522 & x_13524;
assign x_13526 = x_13520 & x_13525;
assign x_13527 = x_13516 & x_13526;
assign x_13528 = x_13506 & x_13527;
assign x_13529 = x_13485 & x_13528;
assign x_13530 = x_13442 & x_13529;
assign x_13531 = x_2285 & x_2286;
assign x_13532 = x_2288 & x_2289;
assign x_13533 = x_2287 & x_13532;
assign x_13534 = x_13531 & x_13533;
assign x_13535 = x_2291 & x_2292;
assign x_13536 = x_2290 & x_13535;
assign x_13537 = x_2294 & x_2295;
assign x_13538 = x_2293 & x_13537;
assign x_13539 = x_13536 & x_13538;
assign x_13540 = x_13534 & x_13539;
assign x_13541 = x_2296 & x_2297;
assign x_13542 = x_2299 & x_2300;
assign x_13543 = x_2298 & x_13542;
assign x_13544 = x_13541 & x_13543;
assign x_13545 = x_2302 & x_2303;
assign x_13546 = x_2301 & x_13545;
assign x_13547 = x_2305 & x_2306;
assign x_13548 = x_2304 & x_13547;
assign x_13549 = x_13546 & x_13548;
assign x_13550 = x_13544 & x_13549;
assign x_13551 = x_13540 & x_13550;
assign x_13552 = x_2307 & x_2308;
assign x_13553 = x_2310 & x_2311;
assign x_13554 = x_2309 & x_13553;
assign x_13555 = x_13552 & x_13554;
assign x_13556 = x_2313 & x_2314;
assign x_13557 = x_2312 & x_13556;
assign x_13558 = x_2316 & x_2317;
assign x_13559 = x_2315 & x_13558;
assign x_13560 = x_13557 & x_13559;
assign x_13561 = x_13555 & x_13560;
assign x_13562 = x_2318 & x_2319;
assign x_13563 = x_2321 & x_2322;
assign x_13564 = x_2320 & x_13563;
assign x_13565 = x_13562 & x_13564;
assign x_13566 = x_2324 & x_2325;
assign x_13567 = x_2323 & x_13566;
assign x_13568 = x_2327 & x_2328;
assign x_13569 = x_2326 & x_13568;
assign x_13570 = x_13567 & x_13569;
assign x_13571 = x_13565 & x_13570;
assign x_13572 = x_13561 & x_13571;
assign x_13573 = x_13551 & x_13572;
assign x_13574 = x_2329 & x_2330;
assign x_13575 = x_2332 & x_2333;
assign x_13576 = x_2331 & x_13575;
assign x_13577 = x_13574 & x_13576;
assign x_13578 = x_2335 & x_2336;
assign x_13579 = x_2334 & x_13578;
assign x_13580 = x_2338 & x_2339;
assign x_13581 = x_2337 & x_13580;
assign x_13582 = x_13579 & x_13581;
assign x_13583 = x_13577 & x_13582;
assign x_13584 = x_2340 & x_2341;
assign x_13585 = x_2343 & x_2344;
assign x_13586 = x_2342 & x_13585;
assign x_13587 = x_13584 & x_13586;
assign x_13588 = x_2346 & x_2347;
assign x_13589 = x_2345 & x_13588;
assign x_13590 = x_2349 & x_2350;
assign x_13591 = x_2348 & x_13590;
assign x_13592 = x_13589 & x_13591;
assign x_13593 = x_13587 & x_13592;
assign x_13594 = x_13583 & x_13593;
assign x_13595 = x_2351 & x_2352;
assign x_13596 = x_2354 & x_2355;
assign x_13597 = x_2353 & x_13596;
assign x_13598 = x_13595 & x_13597;
assign x_13599 = x_2357 & x_2358;
assign x_13600 = x_2356 & x_13599;
assign x_13601 = x_2360 & x_2361;
assign x_13602 = x_2359 & x_13601;
assign x_13603 = x_13600 & x_13602;
assign x_13604 = x_13598 & x_13603;
assign x_13605 = x_2362 & x_2363;
assign x_13606 = x_2365 & x_2366;
assign x_13607 = x_2364 & x_13606;
assign x_13608 = x_13605 & x_13607;
assign x_13609 = x_2368 & x_2369;
assign x_13610 = x_2367 & x_13609;
assign x_13611 = x_2371 & x_2372;
assign x_13612 = x_2370 & x_13611;
assign x_13613 = x_13610 & x_13612;
assign x_13614 = x_13608 & x_13613;
assign x_13615 = x_13604 & x_13614;
assign x_13616 = x_13594 & x_13615;
assign x_13617 = x_13573 & x_13616;
assign x_13618 = x_2373 & x_2374;
assign x_13619 = x_2376 & x_2377;
assign x_13620 = x_2375 & x_13619;
assign x_13621 = x_13618 & x_13620;
assign x_13622 = x_2379 & x_2380;
assign x_13623 = x_2378 & x_13622;
assign x_13624 = x_2382 & x_2383;
assign x_13625 = x_2381 & x_13624;
assign x_13626 = x_13623 & x_13625;
assign x_13627 = x_13621 & x_13626;
assign x_13628 = x_2384 & x_2385;
assign x_13629 = x_2387 & x_2388;
assign x_13630 = x_2386 & x_13629;
assign x_13631 = x_13628 & x_13630;
assign x_13632 = x_2390 & x_2391;
assign x_13633 = x_2389 & x_13632;
assign x_13634 = x_2393 & x_2394;
assign x_13635 = x_2392 & x_13634;
assign x_13636 = x_13633 & x_13635;
assign x_13637 = x_13631 & x_13636;
assign x_13638 = x_13627 & x_13637;
assign x_13639 = x_2395 & x_2396;
assign x_13640 = x_2398 & x_2399;
assign x_13641 = x_2397 & x_13640;
assign x_13642 = x_13639 & x_13641;
assign x_13643 = x_2401 & x_2402;
assign x_13644 = x_2400 & x_13643;
assign x_13645 = x_2404 & x_2405;
assign x_13646 = x_2403 & x_13645;
assign x_13647 = x_13644 & x_13646;
assign x_13648 = x_13642 & x_13647;
assign x_13649 = x_2406 & x_2407;
assign x_13650 = x_2409 & x_2410;
assign x_13651 = x_2408 & x_13650;
assign x_13652 = x_13649 & x_13651;
assign x_13653 = x_2412 & x_2413;
assign x_13654 = x_2411 & x_13653;
assign x_13655 = x_2415 & x_2416;
assign x_13656 = x_2414 & x_13655;
assign x_13657 = x_13654 & x_13656;
assign x_13658 = x_13652 & x_13657;
assign x_13659 = x_13648 & x_13658;
assign x_13660 = x_13638 & x_13659;
assign x_13661 = x_2417 & x_2418;
assign x_13662 = x_2420 & x_2421;
assign x_13663 = x_2419 & x_13662;
assign x_13664 = x_13661 & x_13663;
assign x_13665 = x_2423 & x_2424;
assign x_13666 = x_2422 & x_13665;
assign x_13667 = x_2426 & x_2427;
assign x_13668 = x_2425 & x_13667;
assign x_13669 = x_13666 & x_13668;
assign x_13670 = x_13664 & x_13669;
assign x_13671 = x_2428 & x_2429;
assign x_13672 = x_2431 & x_2432;
assign x_13673 = x_2430 & x_13672;
assign x_13674 = x_13671 & x_13673;
assign x_13675 = x_2434 & x_2435;
assign x_13676 = x_2433 & x_13675;
assign x_13677 = x_2437 & x_2438;
assign x_13678 = x_2436 & x_13677;
assign x_13679 = x_13676 & x_13678;
assign x_13680 = x_13674 & x_13679;
assign x_13681 = x_13670 & x_13680;
assign x_13682 = x_2439 & x_2440;
assign x_13683 = x_2442 & x_2443;
assign x_13684 = x_2441 & x_13683;
assign x_13685 = x_13682 & x_13684;
assign x_13686 = x_2445 & x_2446;
assign x_13687 = x_2444 & x_13686;
assign x_13688 = x_2448 & x_2449;
assign x_13689 = x_2447 & x_13688;
assign x_13690 = x_13687 & x_13689;
assign x_13691 = x_13685 & x_13690;
assign x_13692 = x_2450 & x_2451;
assign x_13693 = x_2453 & x_2454;
assign x_13694 = x_2452 & x_13693;
assign x_13695 = x_13692 & x_13694;
assign x_13696 = x_2456 & x_2457;
assign x_13697 = x_2455 & x_13696;
assign x_13698 = x_2459 & x_2460;
assign x_13699 = x_2458 & x_13698;
assign x_13700 = x_13697 & x_13699;
assign x_13701 = x_13695 & x_13700;
assign x_13702 = x_13691 & x_13701;
assign x_13703 = x_13681 & x_13702;
assign x_13704 = x_13660 & x_13703;
assign x_13705 = x_13617 & x_13704;
assign x_13706 = x_13530 & x_13705;
assign x_13707 = x_2461 & x_2462;
assign x_13708 = x_2464 & x_2465;
assign x_13709 = x_2463 & x_13708;
assign x_13710 = x_13707 & x_13709;
assign x_13711 = x_2467 & x_2468;
assign x_13712 = x_2466 & x_13711;
assign x_13713 = x_2470 & x_2471;
assign x_13714 = x_2469 & x_13713;
assign x_13715 = x_13712 & x_13714;
assign x_13716 = x_13710 & x_13715;
assign x_13717 = x_2472 & x_2473;
assign x_13718 = x_2475 & x_2476;
assign x_13719 = x_2474 & x_13718;
assign x_13720 = x_13717 & x_13719;
assign x_13721 = x_2478 & x_2479;
assign x_13722 = x_2477 & x_13721;
assign x_13723 = x_2481 & x_2482;
assign x_13724 = x_2480 & x_13723;
assign x_13725 = x_13722 & x_13724;
assign x_13726 = x_13720 & x_13725;
assign x_13727 = x_13716 & x_13726;
assign x_13728 = x_2483 & x_2484;
assign x_13729 = x_2486 & x_2487;
assign x_13730 = x_2485 & x_13729;
assign x_13731 = x_13728 & x_13730;
assign x_13732 = x_2489 & x_2490;
assign x_13733 = x_2488 & x_13732;
assign x_13734 = x_2492 & x_2493;
assign x_13735 = x_2491 & x_13734;
assign x_13736 = x_13733 & x_13735;
assign x_13737 = x_13731 & x_13736;
assign x_13738 = x_2494 & x_2495;
assign x_13739 = x_2497 & x_2498;
assign x_13740 = x_2496 & x_13739;
assign x_13741 = x_13738 & x_13740;
assign x_13742 = x_2500 & x_2501;
assign x_13743 = x_2499 & x_13742;
assign x_13744 = x_2503 & x_2504;
assign x_13745 = x_2502 & x_13744;
assign x_13746 = x_13743 & x_13745;
assign x_13747 = x_13741 & x_13746;
assign x_13748 = x_13737 & x_13747;
assign x_13749 = x_13727 & x_13748;
assign x_13750 = x_2505 & x_2506;
assign x_13751 = x_2508 & x_2509;
assign x_13752 = x_2507 & x_13751;
assign x_13753 = x_13750 & x_13752;
assign x_13754 = x_2511 & x_2512;
assign x_13755 = x_2510 & x_13754;
assign x_13756 = x_2514 & x_2515;
assign x_13757 = x_2513 & x_13756;
assign x_13758 = x_13755 & x_13757;
assign x_13759 = x_13753 & x_13758;
assign x_13760 = x_2516 & x_2517;
assign x_13761 = x_2519 & x_2520;
assign x_13762 = x_2518 & x_13761;
assign x_13763 = x_13760 & x_13762;
assign x_13764 = x_2522 & x_2523;
assign x_13765 = x_2521 & x_13764;
assign x_13766 = x_2525 & x_2526;
assign x_13767 = x_2524 & x_13766;
assign x_13768 = x_13765 & x_13767;
assign x_13769 = x_13763 & x_13768;
assign x_13770 = x_13759 & x_13769;
assign x_13771 = x_2527 & x_2528;
assign x_13772 = x_2530 & x_2531;
assign x_13773 = x_2529 & x_13772;
assign x_13774 = x_13771 & x_13773;
assign x_13775 = x_2533 & x_2534;
assign x_13776 = x_2532 & x_13775;
assign x_13777 = x_2536 & x_2537;
assign x_13778 = x_2535 & x_13777;
assign x_13779 = x_13776 & x_13778;
assign x_13780 = x_13774 & x_13779;
assign x_13781 = x_2538 & x_2539;
assign x_13782 = x_2541 & x_2542;
assign x_13783 = x_2540 & x_13782;
assign x_13784 = x_13781 & x_13783;
assign x_13785 = x_2544 & x_2545;
assign x_13786 = x_2543 & x_13785;
assign x_13787 = x_2547 & x_2548;
assign x_13788 = x_2546 & x_13787;
assign x_13789 = x_13786 & x_13788;
assign x_13790 = x_13784 & x_13789;
assign x_13791 = x_13780 & x_13790;
assign x_13792 = x_13770 & x_13791;
assign x_13793 = x_13749 & x_13792;
assign x_13794 = x_2549 & x_2550;
assign x_13795 = x_2552 & x_2553;
assign x_13796 = x_2551 & x_13795;
assign x_13797 = x_13794 & x_13796;
assign x_13798 = x_2555 & x_2556;
assign x_13799 = x_2554 & x_13798;
assign x_13800 = x_2558 & x_2559;
assign x_13801 = x_2557 & x_13800;
assign x_13802 = x_13799 & x_13801;
assign x_13803 = x_13797 & x_13802;
assign x_13804 = x_2560 & x_2561;
assign x_13805 = x_2563 & x_2564;
assign x_13806 = x_2562 & x_13805;
assign x_13807 = x_13804 & x_13806;
assign x_13808 = x_2566 & x_2567;
assign x_13809 = x_2565 & x_13808;
assign x_13810 = x_2569 & x_2570;
assign x_13811 = x_2568 & x_13810;
assign x_13812 = x_13809 & x_13811;
assign x_13813 = x_13807 & x_13812;
assign x_13814 = x_13803 & x_13813;
assign x_13815 = x_2571 & x_2572;
assign x_13816 = x_2574 & x_2575;
assign x_13817 = x_2573 & x_13816;
assign x_13818 = x_13815 & x_13817;
assign x_13819 = x_2577 & x_2578;
assign x_13820 = x_2576 & x_13819;
assign x_13821 = x_2580 & x_2581;
assign x_13822 = x_2579 & x_13821;
assign x_13823 = x_13820 & x_13822;
assign x_13824 = x_13818 & x_13823;
assign x_13825 = x_2582 & x_2583;
assign x_13826 = x_2585 & x_2586;
assign x_13827 = x_2584 & x_13826;
assign x_13828 = x_13825 & x_13827;
assign x_13829 = x_2588 & x_2589;
assign x_13830 = x_2587 & x_13829;
assign x_13831 = x_2591 & x_2592;
assign x_13832 = x_2590 & x_13831;
assign x_13833 = x_13830 & x_13832;
assign x_13834 = x_13828 & x_13833;
assign x_13835 = x_13824 & x_13834;
assign x_13836 = x_13814 & x_13835;
assign x_13837 = x_2593 & x_2594;
assign x_13838 = x_2596 & x_2597;
assign x_13839 = x_2595 & x_13838;
assign x_13840 = x_13837 & x_13839;
assign x_13841 = x_2599 & x_2600;
assign x_13842 = x_2598 & x_13841;
assign x_13843 = x_2602 & x_2603;
assign x_13844 = x_2601 & x_13843;
assign x_13845 = x_13842 & x_13844;
assign x_13846 = x_13840 & x_13845;
assign x_13847 = x_2604 & x_2605;
assign x_13848 = x_2607 & x_2608;
assign x_13849 = x_2606 & x_13848;
assign x_13850 = x_13847 & x_13849;
assign x_13851 = x_2610 & x_2611;
assign x_13852 = x_2609 & x_13851;
assign x_13853 = x_2613 & x_2614;
assign x_13854 = x_2612 & x_13853;
assign x_13855 = x_13852 & x_13854;
assign x_13856 = x_13850 & x_13855;
assign x_13857 = x_13846 & x_13856;
assign x_13858 = x_2615 & x_2616;
assign x_13859 = x_2618 & x_2619;
assign x_13860 = x_2617 & x_13859;
assign x_13861 = x_13858 & x_13860;
assign x_13862 = x_2621 & x_2622;
assign x_13863 = x_2620 & x_13862;
assign x_13864 = x_2624 & x_2625;
assign x_13865 = x_2623 & x_13864;
assign x_13866 = x_13863 & x_13865;
assign x_13867 = x_13861 & x_13866;
assign x_13868 = x_2626 & x_2627;
assign x_13869 = x_2629 & x_2630;
assign x_13870 = x_2628 & x_13869;
assign x_13871 = x_13868 & x_13870;
assign x_13872 = x_2632 & x_2633;
assign x_13873 = x_2631 & x_13872;
assign x_13874 = x_2635 & x_2636;
assign x_13875 = x_2634 & x_13874;
assign x_13876 = x_13873 & x_13875;
assign x_13877 = x_13871 & x_13876;
assign x_13878 = x_13867 & x_13877;
assign x_13879 = x_13857 & x_13878;
assign x_13880 = x_13836 & x_13879;
assign x_13881 = x_13793 & x_13880;
assign x_13882 = x_2637 & x_2638;
assign x_13883 = x_2640 & x_2641;
assign x_13884 = x_2639 & x_13883;
assign x_13885 = x_13882 & x_13884;
assign x_13886 = x_2643 & x_2644;
assign x_13887 = x_2642 & x_13886;
assign x_13888 = x_2646 & x_2647;
assign x_13889 = x_2645 & x_13888;
assign x_13890 = x_13887 & x_13889;
assign x_13891 = x_13885 & x_13890;
assign x_13892 = x_2648 & x_2649;
assign x_13893 = x_2651 & x_2652;
assign x_13894 = x_2650 & x_13893;
assign x_13895 = x_13892 & x_13894;
assign x_13896 = x_2654 & x_2655;
assign x_13897 = x_2653 & x_13896;
assign x_13898 = x_2657 & x_2658;
assign x_13899 = x_2656 & x_13898;
assign x_13900 = x_13897 & x_13899;
assign x_13901 = x_13895 & x_13900;
assign x_13902 = x_13891 & x_13901;
assign x_13903 = x_2659 & x_2660;
assign x_13904 = x_2662 & x_2663;
assign x_13905 = x_2661 & x_13904;
assign x_13906 = x_13903 & x_13905;
assign x_13907 = x_2665 & x_2666;
assign x_13908 = x_2664 & x_13907;
assign x_13909 = x_2668 & x_2669;
assign x_13910 = x_2667 & x_13909;
assign x_13911 = x_13908 & x_13910;
assign x_13912 = x_13906 & x_13911;
assign x_13913 = x_2670 & x_2671;
assign x_13914 = x_2673 & x_2674;
assign x_13915 = x_2672 & x_13914;
assign x_13916 = x_13913 & x_13915;
assign x_13917 = x_2676 & x_2677;
assign x_13918 = x_2675 & x_13917;
assign x_13919 = x_2679 & x_2680;
assign x_13920 = x_2678 & x_13919;
assign x_13921 = x_13918 & x_13920;
assign x_13922 = x_13916 & x_13921;
assign x_13923 = x_13912 & x_13922;
assign x_13924 = x_13902 & x_13923;
assign x_13925 = x_2681 & x_2682;
assign x_13926 = x_2684 & x_2685;
assign x_13927 = x_2683 & x_13926;
assign x_13928 = x_13925 & x_13927;
assign x_13929 = x_2687 & x_2688;
assign x_13930 = x_2686 & x_13929;
assign x_13931 = x_2690 & x_2691;
assign x_13932 = x_2689 & x_13931;
assign x_13933 = x_13930 & x_13932;
assign x_13934 = x_13928 & x_13933;
assign x_13935 = x_2692 & x_2693;
assign x_13936 = x_2695 & x_2696;
assign x_13937 = x_2694 & x_13936;
assign x_13938 = x_13935 & x_13937;
assign x_13939 = x_2698 & x_2699;
assign x_13940 = x_2697 & x_13939;
assign x_13941 = x_2701 & x_2702;
assign x_13942 = x_2700 & x_13941;
assign x_13943 = x_13940 & x_13942;
assign x_13944 = x_13938 & x_13943;
assign x_13945 = x_13934 & x_13944;
assign x_13946 = x_2703 & x_2704;
assign x_13947 = x_2706 & x_2707;
assign x_13948 = x_2705 & x_13947;
assign x_13949 = x_13946 & x_13948;
assign x_13950 = x_2709 & x_2710;
assign x_13951 = x_2708 & x_13950;
assign x_13952 = x_2712 & x_2713;
assign x_13953 = x_2711 & x_13952;
assign x_13954 = x_13951 & x_13953;
assign x_13955 = x_13949 & x_13954;
assign x_13956 = x_2714 & x_2715;
assign x_13957 = x_2717 & x_2718;
assign x_13958 = x_2716 & x_13957;
assign x_13959 = x_13956 & x_13958;
assign x_13960 = x_2720 & x_2721;
assign x_13961 = x_2719 & x_13960;
assign x_13962 = x_2723 & x_2724;
assign x_13963 = x_2722 & x_13962;
assign x_13964 = x_13961 & x_13963;
assign x_13965 = x_13959 & x_13964;
assign x_13966 = x_13955 & x_13965;
assign x_13967 = x_13945 & x_13966;
assign x_13968 = x_13924 & x_13967;
assign x_13969 = x_2725 & x_2726;
assign x_13970 = x_2728 & x_2729;
assign x_13971 = x_2727 & x_13970;
assign x_13972 = x_13969 & x_13971;
assign x_13973 = x_2731 & x_2732;
assign x_13974 = x_2730 & x_13973;
assign x_13975 = x_2734 & x_2735;
assign x_13976 = x_2733 & x_13975;
assign x_13977 = x_13974 & x_13976;
assign x_13978 = x_13972 & x_13977;
assign x_13979 = x_2736 & x_2737;
assign x_13980 = x_2739 & x_2740;
assign x_13981 = x_2738 & x_13980;
assign x_13982 = x_13979 & x_13981;
assign x_13983 = x_2742 & x_2743;
assign x_13984 = x_2741 & x_13983;
assign x_13985 = x_2745 & x_2746;
assign x_13986 = x_2744 & x_13985;
assign x_13987 = x_13984 & x_13986;
assign x_13988 = x_13982 & x_13987;
assign x_13989 = x_13978 & x_13988;
assign x_13990 = x_2747 & x_2748;
assign x_13991 = x_2750 & x_2751;
assign x_13992 = x_2749 & x_13991;
assign x_13993 = x_13990 & x_13992;
assign x_13994 = x_2753 & x_2754;
assign x_13995 = x_2752 & x_13994;
assign x_13996 = x_2756 & x_2757;
assign x_13997 = x_2755 & x_13996;
assign x_13998 = x_13995 & x_13997;
assign x_13999 = x_13993 & x_13998;
assign x_14000 = x_2758 & x_2759;
assign x_14001 = x_2761 & x_2762;
assign x_14002 = x_2760 & x_14001;
assign x_14003 = x_14000 & x_14002;
assign x_14004 = x_2764 & x_2765;
assign x_14005 = x_2763 & x_14004;
assign x_14006 = x_2767 & x_2768;
assign x_14007 = x_2766 & x_14006;
assign x_14008 = x_14005 & x_14007;
assign x_14009 = x_14003 & x_14008;
assign x_14010 = x_13999 & x_14009;
assign x_14011 = x_13989 & x_14010;
assign x_14012 = x_2769 & x_2770;
assign x_14013 = x_2772 & x_2773;
assign x_14014 = x_2771 & x_14013;
assign x_14015 = x_14012 & x_14014;
assign x_14016 = x_2775 & x_2776;
assign x_14017 = x_2774 & x_14016;
assign x_14018 = x_2778 & x_2779;
assign x_14019 = x_2777 & x_14018;
assign x_14020 = x_14017 & x_14019;
assign x_14021 = x_14015 & x_14020;
assign x_14022 = x_2780 & x_2781;
assign x_14023 = x_2783 & x_2784;
assign x_14024 = x_2782 & x_14023;
assign x_14025 = x_14022 & x_14024;
assign x_14026 = x_2786 & x_2787;
assign x_14027 = x_2785 & x_14026;
assign x_14028 = x_2789 & x_2790;
assign x_14029 = x_2788 & x_14028;
assign x_14030 = x_14027 & x_14029;
assign x_14031 = x_14025 & x_14030;
assign x_14032 = x_14021 & x_14031;
assign x_14033 = x_2791 & x_2792;
assign x_14034 = x_2794 & x_2795;
assign x_14035 = x_2793 & x_14034;
assign x_14036 = x_14033 & x_14035;
assign x_14037 = x_2797 & x_2798;
assign x_14038 = x_2796 & x_14037;
assign x_14039 = x_2800 & x_2801;
assign x_14040 = x_2799 & x_14039;
assign x_14041 = x_14038 & x_14040;
assign x_14042 = x_14036 & x_14041;
assign x_14043 = x_2802 & x_2803;
assign x_14044 = x_2805 & x_2806;
assign x_14045 = x_2804 & x_14044;
assign x_14046 = x_14043 & x_14045;
assign x_14047 = x_2808 & x_2809;
assign x_14048 = x_2807 & x_14047;
assign x_14049 = x_2811 & x_2812;
assign x_14050 = x_2810 & x_14049;
assign x_14051 = x_14048 & x_14050;
assign x_14052 = x_14046 & x_14051;
assign x_14053 = x_14042 & x_14052;
assign x_14054 = x_14032 & x_14053;
assign x_14055 = x_14011 & x_14054;
assign x_14056 = x_13968 & x_14055;
assign x_14057 = x_13881 & x_14056;
assign x_14058 = x_13706 & x_14057;
assign x_14059 = x_13356 & x_14058;
assign x_14060 = x_12654 & x_14059;
assign x_14061 = x_2813 & x_2814;
assign x_14062 = x_2816 & x_2817;
assign x_14063 = x_2815 & x_14062;
assign x_14064 = x_14061 & x_14063;
assign x_14065 = x_2818 & x_2819;
assign x_14066 = x_2821 & x_2822;
assign x_14067 = x_2820 & x_14066;
assign x_14068 = x_14065 & x_14067;
assign x_14069 = x_14064 & x_14068;
assign x_14070 = x_2823 & x_2824;
assign x_14071 = x_2826 & x_2827;
assign x_14072 = x_2825 & x_14071;
assign x_14073 = x_14070 & x_14072;
assign x_14074 = x_2829 & x_2830;
assign x_14075 = x_2828 & x_14074;
assign x_14076 = x_2832 & x_2833;
assign x_14077 = x_2831 & x_14076;
assign x_14078 = x_14075 & x_14077;
assign x_14079 = x_14073 & x_14078;
assign x_14080 = x_14069 & x_14079;
assign x_14081 = x_2834 & x_2835;
assign x_14082 = x_2837 & x_2838;
assign x_14083 = x_2836 & x_14082;
assign x_14084 = x_14081 & x_14083;
assign x_14085 = x_2840 & x_2841;
assign x_14086 = x_2839 & x_14085;
assign x_14087 = x_2843 & x_2844;
assign x_14088 = x_2842 & x_14087;
assign x_14089 = x_14086 & x_14088;
assign x_14090 = x_14084 & x_14089;
assign x_14091 = x_2845 & x_2846;
assign x_14092 = x_2848 & x_2849;
assign x_14093 = x_2847 & x_14092;
assign x_14094 = x_14091 & x_14093;
assign x_14095 = x_2851 & x_2852;
assign x_14096 = x_2850 & x_14095;
assign x_14097 = x_2854 & x_2855;
assign x_14098 = x_2853 & x_14097;
assign x_14099 = x_14096 & x_14098;
assign x_14100 = x_14094 & x_14099;
assign x_14101 = x_14090 & x_14100;
assign x_14102 = x_14080 & x_14101;
assign x_14103 = x_2856 & x_2857;
assign x_14104 = x_2859 & x_2860;
assign x_14105 = x_2858 & x_14104;
assign x_14106 = x_14103 & x_14105;
assign x_14107 = x_2862 & x_2863;
assign x_14108 = x_2861 & x_14107;
assign x_14109 = x_2865 & x_2866;
assign x_14110 = x_2864 & x_14109;
assign x_14111 = x_14108 & x_14110;
assign x_14112 = x_14106 & x_14111;
assign x_14113 = x_2867 & x_2868;
assign x_14114 = x_2870 & x_2871;
assign x_14115 = x_2869 & x_14114;
assign x_14116 = x_14113 & x_14115;
assign x_14117 = x_2873 & x_2874;
assign x_14118 = x_2872 & x_14117;
assign x_14119 = x_2876 & x_2877;
assign x_14120 = x_2875 & x_14119;
assign x_14121 = x_14118 & x_14120;
assign x_14122 = x_14116 & x_14121;
assign x_14123 = x_14112 & x_14122;
assign x_14124 = x_2878 & x_2879;
assign x_14125 = x_2881 & x_2882;
assign x_14126 = x_2880 & x_14125;
assign x_14127 = x_14124 & x_14126;
assign x_14128 = x_2884 & x_2885;
assign x_14129 = x_2883 & x_14128;
assign x_14130 = x_2887 & x_2888;
assign x_14131 = x_2886 & x_14130;
assign x_14132 = x_14129 & x_14131;
assign x_14133 = x_14127 & x_14132;
assign x_14134 = x_2889 & x_2890;
assign x_14135 = x_2892 & x_2893;
assign x_14136 = x_2891 & x_14135;
assign x_14137 = x_14134 & x_14136;
assign x_14138 = x_2895 & x_2896;
assign x_14139 = x_2894 & x_14138;
assign x_14140 = x_2898 & x_2899;
assign x_14141 = x_2897 & x_14140;
assign x_14142 = x_14139 & x_14141;
assign x_14143 = x_14137 & x_14142;
assign x_14144 = x_14133 & x_14143;
assign x_14145 = x_14123 & x_14144;
assign x_14146 = x_14102 & x_14145;
assign x_14147 = x_2900 & x_2901;
assign x_14148 = x_2903 & x_2904;
assign x_14149 = x_2902 & x_14148;
assign x_14150 = x_14147 & x_14149;
assign x_14151 = x_2906 & x_2907;
assign x_14152 = x_2905 & x_14151;
assign x_14153 = x_2909 & x_2910;
assign x_14154 = x_2908 & x_14153;
assign x_14155 = x_14152 & x_14154;
assign x_14156 = x_14150 & x_14155;
assign x_14157 = x_2911 & x_2912;
assign x_14158 = x_2914 & x_2915;
assign x_14159 = x_2913 & x_14158;
assign x_14160 = x_14157 & x_14159;
assign x_14161 = x_2917 & x_2918;
assign x_14162 = x_2916 & x_14161;
assign x_14163 = x_2920 & x_2921;
assign x_14164 = x_2919 & x_14163;
assign x_14165 = x_14162 & x_14164;
assign x_14166 = x_14160 & x_14165;
assign x_14167 = x_14156 & x_14166;
assign x_14168 = x_2922 & x_2923;
assign x_14169 = x_2925 & x_2926;
assign x_14170 = x_2924 & x_14169;
assign x_14171 = x_14168 & x_14170;
assign x_14172 = x_2928 & x_2929;
assign x_14173 = x_2927 & x_14172;
assign x_14174 = x_2931 & x_2932;
assign x_14175 = x_2930 & x_14174;
assign x_14176 = x_14173 & x_14175;
assign x_14177 = x_14171 & x_14176;
assign x_14178 = x_2933 & x_2934;
assign x_14179 = x_2936 & x_2937;
assign x_14180 = x_2935 & x_14179;
assign x_14181 = x_14178 & x_14180;
assign x_14182 = x_2939 & x_2940;
assign x_14183 = x_2938 & x_14182;
assign x_14184 = x_2942 & x_2943;
assign x_14185 = x_2941 & x_14184;
assign x_14186 = x_14183 & x_14185;
assign x_14187 = x_14181 & x_14186;
assign x_14188 = x_14177 & x_14187;
assign x_14189 = x_14167 & x_14188;
assign x_14190 = x_2944 & x_2945;
assign x_14191 = x_2947 & x_2948;
assign x_14192 = x_2946 & x_14191;
assign x_14193 = x_14190 & x_14192;
assign x_14194 = x_2950 & x_2951;
assign x_14195 = x_2949 & x_14194;
assign x_14196 = x_2953 & x_2954;
assign x_14197 = x_2952 & x_14196;
assign x_14198 = x_14195 & x_14197;
assign x_14199 = x_14193 & x_14198;
assign x_14200 = x_2955 & x_2956;
assign x_14201 = x_2958 & x_2959;
assign x_14202 = x_2957 & x_14201;
assign x_14203 = x_14200 & x_14202;
assign x_14204 = x_2961 & x_2962;
assign x_14205 = x_2960 & x_14204;
assign x_14206 = x_2964 & x_2965;
assign x_14207 = x_2963 & x_14206;
assign x_14208 = x_14205 & x_14207;
assign x_14209 = x_14203 & x_14208;
assign x_14210 = x_14199 & x_14209;
assign x_14211 = x_2966 & x_2967;
assign x_14212 = x_2969 & x_2970;
assign x_14213 = x_2968 & x_14212;
assign x_14214 = x_14211 & x_14213;
assign x_14215 = x_2972 & x_2973;
assign x_14216 = x_2971 & x_14215;
assign x_14217 = x_2975 & x_2976;
assign x_14218 = x_2974 & x_14217;
assign x_14219 = x_14216 & x_14218;
assign x_14220 = x_14214 & x_14219;
assign x_14221 = x_2977 & x_2978;
assign x_14222 = x_2980 & x_2981;
assign x_14223 = x_2979 & x_14222;
assign x_14224 = x_14221 & x_14223;
assign x_14225 = x_2983 & x_2984;
assign x_14226 = x_2982 & x_14225;
assign x_14227 = x_2986 & x_2987;
assign x_14228 = x_2985 & x_14227;
assign x_14229 = x_14226 & x_14228;
assign x_14230 = x_14224 & x_14229;
assign x_14231 = x_14220 & x_14230;
assign x_14232 = x_14210 & x_14231;
assign x_14233 = x_14189 & x_14232;
assign x_14234 = x_14146 & x_14233;
assign x_14235 = x_2988 & x_2989;
assign x_14236 = x_2991 & x_2992;
assign x_14237 = x_2990 & x_14236;
assign x_14238 = x_14235 & x_14237;
assign x_14239 = x_2994 & x_2995;
assign x_14240 = x_2993 & x_14239;
assign x_14241 = x_2997 & x_2998;
assign x_14242 = x_2996 & x_14241;
assign x_14243 = x_14240 & x_14242;
assign x_14244 = x_14238 & x_14243;
assign x_14245 = x_2999 & x_3000;
assign x_14246 = x_3002 & x_3003;
assign x_14247 = x_3001 & x_14246;
assign x_14248 = x_14245 & x_14247;
assign x_14249 = x_3005 & x_3006;
assign x_14250 = x_3004 & x_14249;
assign x_14251 = x_3008 & x_3009;
assign x_14252 = x_3007 & x_14251;
assign x_14253 = x_14250 & x_14252;
assign x_14254 = x_14248 & x_14253;
assign x_14255 = x_14244 & x_14254;
assign x_14256 = x_3010 & x_3011;
assign x_14257 = x_3013 & x_3014;
assign x_14258 = x_3012 & x_14257;
assign x_14259 = x_14256 & x_14258;
assign x_14260 = x_3016 & x_3017;
assign x_14261 = x_3015 & x_14260;
assign x_14262 = x_3019 & x_3020;
assign x_14263 = x_3018 & x_14262;
assign x_14264 = x_14261 & x_14263;
assign x_14265 = x_14259 & x_14264;
assign x_14266 = x_3021 & x_3022;
assign x_14267 = x_3024 & x_3025;
assign x_14268 = x_3023 & x_14267;
assign x_14269 = x_14266 & x_14268;
assign x_14270 = x_3027 & x_3028;
assign x_14271 = x_3026 & x_14270;
assign x_14272 = x_3030 & x_3031;
assign x_14273 = x_3029 & x_14272;
assign x_14274 = x_14271 & x_14273;
assign x_14275 = x_14269 & x_14274;
assign x_14276 = x_14265 & x_14275;
assign x_14277 = x_14255 & x_14276;
assign x_14278 = x_3032 & x_3033;
assign x_14279 = x_3035 & x_3036;
assign x_14280 = x_3034 & x_14279;
assign x_14281 = x_14278 & x_14280;
assign x_14282 = x_3038 & x_3039;
assign x_14283 = x_3037 & x_14282;
assign x_14284 = x_3041 & x_3042;
assign x_14285 = x_3040 & x_14284;
assign x_14286 = x_14283 & x_14285;
assign x_14287 = x_14281 & x_14286;
assign x_14288 = x_3043 & x_3044;
assign x_14289 = x_3046 & x_3047;
assign x_14290 = x_3045 & x_14289;
assign x_14291 = x_14288 & x_14290;
assign x_14292 = x_3049 & x_3050;
assign x_14293 = x_3048 & x_14292;
assign x_14294 = x_3052 & x_3053;
assign x_14295 = x_3051 & x_14294;
assign x_14296 = x_14293 & x_14295;
assign x_14297 = x_14291 & x_14296;
assign x_14298 = x_14287 & x_14297;
assign x_14299 = x_3054 & x_3055;
assign x_14300 = x_3057 & x_3058;
assign x_14301 = x_3056 & x_14300;
assign x_14302 = x_14299 & x_14301;
assign x_14303 = x_3060 & x_3061;
assign x_14304 = x_3059 & x_14303;
assign x_14305 = x_3063 & x_3064;
assign x_14306 = x_3062 & x_14305;
assign x_14307 = x_14304 & x_14306;
assign x_14308 = x_14302 & x_14307;
assign x_14309 = x_3065 & x_3066;
assign x_14310 = x_3068 & x_3069;
assign x_14311 = x_3067 & x_14310;
assign x_14312 = x_14309 & x_14311;
assign x_14313 = x_3071 & x_3072;
assign x_14314 = x_3070 & x_14313;
assign x_14315 = x_3074 & x_3075;
assign x_14316 = x_3073 & x_14315;
assign x_14317 = x_14314 & x_14316;
assign x_14318 = x_14312 & x_14317;
assign x_14319 = x_14308 & x_14318;
assign x_14320 = x_14298 & x_14319;
assign x_14321 = x_14277 & x_14320;
assign x_14322 = x_3076 & x_3077;
assign x_14323 = x_3079 & x_3080;
assign x_14324 = x_3078 & x_14323;
assign x_14325 = x_14322 & x_14324;
assign x_14326 = x_3082 & x_3083;
assign x_14327 = x_3081 & x_14326;
assign x_14328 = x_3085 & x_3086;
assign x_14329 = x_3084 & x_14328;
assign x_14330 = x_14327 & x_14329;
assign x_14331 = x_14325 & x_14330;
assign x_14332 = x_3087 & x_3088;
assign x_14333 = x_3090 & x_3091;
assign x_14334 = x_3089 & x_14333;
assign x_14335 = x_14332 & x_14334;
assign x_14336 = x_3093 & x_3094;
assign x_14337 = x_3092 & x_14336;
assign x_14338 = x_3096 & x_3097;
assign x_14339 = x_3095 & x_14338;
assign x_14340 = x_14337 & x_14339;
assign x_14341 = x_14335 & x_14340;
assign x_14342 = x_14331 & x_14341;
assign x_14343 = x_3098 & x_3099;
assign x_14344 = x_3101 & x_3102;
assign x_14345 = x_3100 & x_14344;
assign x_14346 = x_14343 & x_14345;
assign x_14347 = x_3104 & x_3105;
assign x_14348 = x_3103 & x_14347;
assign x_14349 = x_3107 & x_3108;
assign x_14350 = x_3106 & x_14349;
assign x_14351 = x_14348 & x_14350;
assign x_14352 = x_14346 & x_14351;
assign x_14353 = x_3109 & x_3110;
assign x_14354 = x_3112 & x_3113;
assign x_14355 = x_3111 & x_14354;
assign x_14356 = x_14353 & x_14355;
assign x_14357 = x_3115 & x_3116;
assign x_14358 = x_3114 & x_14357;
assign x_14359 = x_3118 & x_3119;
assign x_14360 = x_3117 & x_14359;
assign x_14361 = x_14358 & x_14360;
assign x_14362 = x_14356 & x_14361;
assign x_14363 = x_14352 & x_14362;
assign x_14364 = x_14342 & x_14363;
assign x_14365 = x_3120 & x_3121;
assign x_14366 = x_3123 & x_3124;
assign x_14367 = x_3122 & x_14366;
assign x_14368 = x_14365 & x_14367;
assign x_14369 = x_3126 & x_3127;
assign x_14370 = x_3125 & x_14369;
assign x_14371 = x_3129 & x_3130;
assign x_14372 = x_3128 & x_14371;
assign x_14373 = x_14370 & x_14372;
assign x_14374 = x_14368 & x_14373;
assign x_14375 = x_3131 & x_3132;
assign x_14376 = x_3134 & x_3135;
assign x_14377 = x_3133 & x_14376;
assign x_14378 = x_14375 & x_14377;
assign x_14379 = x_3137 & x_3138;
assign x_14380 = x_3136 & x_14379;
assign x_14381 = x_3140 & x_3141;
assign x_14382 = x_3139 & x_14381;
assign x_14383 = x_14380 & x_14382;
assign x_14384 = x_14378 & x_14383;
assign x_14385 = x_14374 & x_14384;
assign x_14386 = x_3142 & x_3143;
assign x_14387 = x_3145 & x_3146;
assign x_14388 = x_3144 & x_14387;
assign x_14389 = x_14386 & x_14388;
assign x_14390 = x_3148 & x_3149;
assign x_14391 = x_3147 & x_14390;
assign x_14392 = x_3151 & x_3152;
assign x_14393 = x_3150 & x_14392;
assign x_14394 = x_14391 & x_14393;
assign x_14395 = x_14389 & x_14394;
assign x_14396 = x_3153 & x_3154;
assign x_14397 = x_3156 & x_3157;
assign x_14398 = x_3155 & x_14397;
assign x_14399 = x_14396 & x_14398;
assign x_14400 = x_3159 & x_3160;
assign x_14401 = x_3158 & x_14400;
assign x_14402 = x_3162 & x_3163;
assign x_14403 = x_3161 & x_14402;
assign x_14404 = x_14401 & x_14403;
assign x_14405 = x_14399 & x_14404;
assign x_14406 = x_14395 & x_14405;
assign x_14407 = x_14385 & x_14406;
assign x_14408 = x_14364 & x_14407;
assign x_14409 = x_14321 & x_14408;
assign x_14410 = x_14234 & x_14409;
assign x_14411 = x_3164 & x_3165;
assign x_14412 = x_3167 & x_3168;
assign x_14413 = x_3166 & x_14412;
assign x_14414 = x_14411 & x_14413;
assign x_14415 = x_3170 & x_3171;
assign x_14416 = x_3169 & x_14415;
assign x_14417 = x_3173 & x_3174;
assign x_14418 = x_3172 & x_14417;
assign x_14419 = x_14416 & x_14418;
assign x_14420 = x_14414 & x_14419;
assign x_14421 = x_3175 & x_3176;
assign x_14422 = x_3178 & x_3179;
assign x_14423 = x_3177 & x_14422;
assign x_14424 = x_14421 & x_14423;
assign x_14425 = x_3181 & x_3182;
assign x_14426 = x_3180 & x_14425;
assign x_14427 = x_3184 & x_3185;
assign x_14428 = x_3183 & x_14427;
assign x_14429 = x_14426 & x_14428;
assign x_14430 = x_14424 & x_14429;
assign x_14431 = x_14420 & x_14430;
assign x_14432 = x_3186 & x_3187;
assign x_14433 = x_3189 & x_3190;
assign x_14434 = x_3188 & x_14433;
assign x_14435 = x_14432 & x_14434;
assign x_14436 = x_3192 & x_3193;
assign x_14437 = x_3191 & x_14436;
assign x_14438 = x_3195 & x_3196;
assign x_14439 = x_3194 & x_14438;
assign x_14440 = x_14437 & x_14439;
assign x_14441 = x_14435 & x_14440;
assign x_14442 = x_3197 & x_3198;
assign x_14443 = x_3200 & x_3201;
assign x_14444 = x_3199 & x_14443;
assign x_14445 = x_14442 & x_14444;
assign x_14446 = x_3203 & x_3204;
assign x_14447 = x_3202 & x_14446;
assign x_14448 = x_3206 & x_3207;
assign x_14449 = x_3205 & x_14448;
assign x_14450 = x_14447 & x_14449;
assign x_14451 = x_14445 & x_14450;
assign x_14452 = x_14441 & x_14451;
assign x_14453 = x_14431 & x_14452;
assign x_14454 = x_3208 & x_3209;
assign x_14455 = x_3211 & x_3212;
assign x_14456 = x_3210 & x_14455;
assign x_14457 = x_14454 & x_14456;
assign x_14458 = x_3214 & x_3215;
assign x_14459 = x_3213 & x_14458;
assign x_14460 = x_3217 & x_3218;
assign x_14461 = x_3216 & x_14460;
assign x_14462 = x_14459 & x_14461;
assign x_14463 = x_14457 & x_14462;
assign x_14464 = x_3219 & x_3220;
assign x_14465 = x_3222 & x_3223;
assign x_14466 = x_3221 & x_14465;
assign x_14467 = x_14464 & x_14466;
assign x_14468 = x_3225 & x_3226;
assign x_14469 = x_3224 & x_14468;
assign x_14470 = x_3228 & x_3229;
assign x_14471 = x_3227 & x_14470;
assign x_14472 = x_14469 & x_14471;
assign x_14473 = x_14467 & x_14472;
assign x_14474 = x_14463 & x_14473;
assign x_14475 = x_3230 & x_3231;
assign x_14476 = x_3233 & x_3234;
assign x_14477 = x_3232 & x_14476;
assign x_14478 = x_14475 & x_14477;
assign x_14479 = x_3236 & x_3237;
assign x_14480 = x_3235 & x_14479;
assign x_14481 = x_3239 & x_3240;
assign x_14482 = x_3238 & x_14481;
assign x_14483 = x_14480 & x_14482;
assign x_14484 = x_14478 & x_14483;
assign x_14485 = x_3241 & x_3242;
assign x_14486 = x_3244 & x_3245;
assign x_14487 = x_3243 & x_14486;
assign x_14488 = x_14485 & x_14487;
assign x_14489 = x_3247 & x_3248;
assign x_14490 = x_3246 & x_14489;
assign x_14491 = x_3250 & x_3251;
assign x_14492 = x_3249 & x_14491;
assign x_14493 = x_14490 & x_14492;
assign x_14494 = x_14488 & x_14493;
assign x_14495 = x_14484 & x_14494;
assign x_14496 = x_14474 & x_14495;
assign x_14497 = x_14453 & x_14496;
assign x_14498 = x_3252 & x_3253;
assign x_14499 = x_3255 & x_3256;
assign x_14500 = x_3254 & x_14499;
assign x_14501 = x_14498 & x_14500;
assign x_14502 = x_3258 & x_3259;
assign x_14503 = x_3257 & x_14502;
assign x_14504 = x_3261 & x_3262;
assign x_14505 = x_3260 & x_14504;
assign x_14506 = x_14503 & x_14505;
assign x_14507 = x_14501 & x_14506;
assign x_14508 = x_3263 & x_3264;
assign x_14509 = x_3266 & x_3267;
assign x_14510 = x_3265 & x_14509;
assign x_14511 = x_14508 & x_14510;
assign x_14512 = x_3269 & x_3270;
assign x_14513 = x_3268 & x_14512;
assign x_14514 = x_3272 & x_3273;
assign x_14515 = x_3271 & x_14514;
assign x_14516 = x_14513 & x_14515;
assign x_14517 = x_14511 & x_14516;
assign x_14518 = x_14507 & x_14517;
assign x_14519 = x_3274 & x_3275;
assign x_14520 = x_3277 & x_3278;
assign x_14521 = x_3276 & x_14520;
assign x_14522 = x_14519 & x_14521;
assign x_14523 = x_3280 & x_3281;
assign x_14524 = x_3279 & x_14523;
assign x_14525 = x_3283 & x_3284;
assign x_14526 = x_3282 & x_14525;
assign x_14527 = x_14524 & x_14526;
assign x_14528 = x_14522 & x_14527;
assign x_14529 = x_3285 & x_3286;
assign x_14530 = x_3288 & x_3289;
assign x_14531 = x_3287 & x_14530;
assign x_14532 = x_14529 & x_14531;
assign x_14533 = x_3291 & x_3292;
assign x_14534 = x_3290 & x_14533;
assign x_14535 = x_3294 & x_3295;
assign x_14536 = x_3293 & x_14535;
assign x_14537 = x_14534 & x_14536;
assign x_14538 = x_14532 & x_14537;
assign x_14539 = x_14528 & x_14538;
assign x_14540 = x_14518 & x_14539;
assign x_14541 = x_3296 & x_3297;
assign x_14542 = x_3299 & x_3300;
assign x_14543 = x_3298 & x_14542;
assign x_14544 = x_14541 & x_14543;
assign x_14545 = x_3302 & x_3303;
assign x_14546 = x_3301 & x_14545;
assign x_14547 = x_3305 & x_3306;
assign x_14548 = x_3304 & x_14547;
assign x_14549 = x_14546 & x_14548;
assign x_14550 = x_14544 & x_14549;
assign x_14551 = x_3307 & x_3308;
assign x_14552 = x_3310 & x_3311;
assign x_14553 = x_3309 & x_14552;
assign x_14554 = x_14551 & x_14553;
assign x_14555 = x_3313 & x_3314;
assign x_14556 = x_3312 & x_14555;
assign x_14557 = x_3316 & x_3317;
assign x_14558 = x_3315 & x_14557;
assign x_14559 = x_14556 & x_14558;
assign x_14560 = x_14554 & x_14559;
assign x_14561 = x_14550 & x_14560;
assign x_14562 = x_3318 & x_3319;
assign x_14563 = x_3321 & x_3322;
assign x_14564 = x_3320 & x_14563;
assign x_14565 = x_14562 & x_14564;
assign x_14566 = x_3324 & x_3325;
assign x_14567 = x_3323 & x_14566;
assign x_14568 = x_3327 & x_3328;
assign x_14569 = x_3326 & x_14568;
assign x_14570 = x_14567 & x_14569;
assign x_14571 = x_14565 & x_14570;
assign x_14572 = x_3329 & x_3330;
assign x_14573 = x_3332 & x_3333;
assign x_14574 = x_3331 & x_14573;
assign x_14575 = x_14572 & x_14574;
assign x_14576 = x_3335 & x_3336;
assign x_14577 = x_3334 & x_14576;
assign x_14578 = x_3338 & x_3339;
assign x_14579 = x_3337 & x_14578;
assign x_14580 = x_14577 & x_14579;
assign x_14581 = x_14575 & x_14580;
assign x_14582 = x_14571 & x_14581;
assign x_14583 = x_14561 & x_14582;
assign x_14584 = x_14540 & x_14583;
assign x_14585 = x_14497 & x_14584;
assign x_14586 = x_3340 & x_3341;
assign x_14587 = x_3343 & x_3344;
assign x_14588 = x_3342 & x_14587;
assign x_14589 = x_14586 & x_14588;
assign x_14590 = x_3346 & x_3347;
assign x_14591 = x_3345 & x_14590;
assign x_14592 = x_3349 & x_3350;
assign x_14593 = x_3348 & x_14592;
assign x_14594 = x_14591 & x_14593;
assign x_14595 = x_14589 & x_14594;
assign x_14596 = x_3351 & x_3352;
assign x_14597 = x_3354 & x_3355;
assign x_14598 = x_3353 & x_14597;
assign x_14599 = x_14596 & x_14598;
assign x_14600 = x_3357 & x_3358;
assign x_14601 = x_3356 & x_14600;
assign x_14602 = x_3360 & x_3361;
assign x_14603 = x_3359 & x_14602;
assign x_14604 = x_14601 & x_14603;
assign x_14605 = x_14599 & x_14604;
assign x_14606 = x_14595 & x_14605;
assign x_14607 = x_3362 & x_3363;
assign x_14608 = x_3365 & x_3366;
assign x_14609 = x_3364 & x_14608;
assign x_14610 = x_14607 & x_14609;
assign x_14611 = x_3368 & x_3369;
assign x_14612 = x_3367 & x_14611;
assign x_14613 = x_3371 & x_3372;
assign x_14614 = x_3370 & x_14613;
assign x_14615 = x_14612 & x_14614;
assign x_14616 = x_14610 & x_14615;
assign x_14617 = x_3373 & x_3374;
assign x_14618 = x_3376 & x_3377;
assign x_14619 = x_3375 & x_14618;
assign x_14620 = x_14617 & x_14619;
assign x_14621 = x_3379 & x_3380;
assign x_14622 = x_3378 & x_14621;
assign x_14623 = x_3382 & x_3383;
assign x_14624 = x_3381 & x_14623;
assign x_14625 = x_14622 & x_14624;
assign x_14626 = x_14620 & x_14625;
assign x_14627 = x_14616 & x_14626;
assign x_14628 = x_14606 & x_14627;
assign x_14629 = x_3384 & x_3385;
assign x_14630 = x_3387 & x_3388;
assign x_14631 = x_3386 & x_14630;
assign x_14632 = x_14629 & x_14631;
assign x_14633 = x_3390 & x_3391;
assign x_14634 = x_3389 & x_14633;
assign x_14635 = x_3393 & x_3394;
assign x_14636 = x_3392 & x_14635;
assign x_14637 = x_14634 & x_14636;
assign x_14638 = x_14632 & x_14637;
assign x_14639 = x_3395 & x_3396;
assign x_14640 = x_3398 & x_3399;
assign x_14641 = x_3397 & x_14640;
assign x_14642 = x_14639 & x_14641;
assign x_14643 = x_3401 & x_3402;
assign x_14644 = x_3400 & x_14643;
assign x_14645 = x_3404 & x_3405;
assign x_14646 = x_3403 & x_14645;
assign x_14647 = x_14644 & x_14646;
assign x_14648 = x_14642 & x_14647;
assign x_14649 = x_14638 & x_14648;
assign x_14650 = x_3406 & x_3407;
assign x_14651 = x_3409 & x_3410;
assign x_14652 = x_3408 & x_14651;
assign x_14653 = x_14650 & x_14652;
assign x_14654 = x_3412 & x_3413;
assign x_14655 = x_3411 & x_14654;
assign x_14656 = x_3415 & x_3416;
assign x_14657 = x_3414 & x_14656;
assign x_14658 = x_14655 & x_14657;
assign x_14659 = x_14653 & x_14658;
assign x_14660 = x_3417 & x_3418;
assign x_14661 = x_3420 & x_3421;
assign x_14662 = x_3419 & x_14661;
assign x_14663 = x_14660 & x_14662;
assign x_14664 = x_3423 & x_3424;
assign x_14665 = x_3422 & x_14664;
assign x_14666 = x_3426 & x_3427;
assign x_14667 = x_3425 & x_14666;
assign x_14668 = x_14665 & x_14667;
assign x_14669 = x_14663 & x_14668;
assign x_14670 = x_14659 & x_14669;
assign x_14671 = x_14649 & x_14670;
assign x_14672 = x_14628 & x_14671;
assign x_14673 = x_3428 & x_3429;
assign x_14674 = x_3431 & x_3432;
assign x_14675 = x_3430 & x_14674;
assign x_14676 = x_14673 & x_14675;
assign x_14677 = x_3434 & x_3435;
assign x_14678 = x_3433 & x_14677;
assign x_14679 = x_3437 & x_3438;
assign x_14680 = x_3436 & x_14679;
assign x_14681 = x_14678 & x_14680;
assign x_14682 = x_14676 & x_14681;
assign x_14683 = x_3439 & x_3440;
assign x_14684 = x_3442 & x_3443;
assign x_14685 = x_3441 & x_14684;
assign x_14686 = x_14683 & x_14685;
assign x_14687 = x_3445 & x_3446;
assign x_14688 = x_3444 & x_14687;
assign x_14689 = x_3448 & x_3449;
assign x_14690 = x_3447 & x_14689;
assign x_14691 = x_14688 & x_14690;
assign x_14692 = x_14686 & x_14691;
assign x_14693 = x_14682 & x_14692;
assign x_14694 = x_3450 & x_3451;
assign x_14695 = x_3453 & x_3454;
assign x_14696 = x_3452 & x_14695;
assign x_14697 = x_14694 & x_14696;
assign x_14698 = x_3456 & x_3457;
assign x_14699 = x_3455 & x_14698;
assign x_14700 = x_3459 & x_3460;
assign x_14701 = x_3458 & x_14700;
assign x_14702 = x_14699 & x_14701;
assign x_14703 = x_14697 & x_14702;
assign x_14704 = x_3461 & x_3462;
assign x_14705 = x_3464 & x_3465;
assign x_14706 = x_3463 & x_14705;
assign x_14707 = x_14704 & x_14706;
assign x_14708 = x_3467 & x_3468;
assign x_14709 = x_3466 & x_14708;
assign x_14710 = x_3470 & x_3471;
assign x_14711 = x_3469 & x_14710;
assign x_14712 = x_14709 & x_14711;
assign x_14713 = x_14707 & x_14712;
assign x_14714 = x_14703 & x_14713;
assign x_14715 = x_14693 & x_14714;
assign x_14716 = x_3472 & x_3473;
assign x_14717 = x_3475 & x_3476;
assign x_14718 = x_3474 & x_14717;
assign x_14719 = x_14716 & x_14718;
assign x_14720 = x_3478 & x_3479;
assign x_14721 = x_3477 & x_14720;
assign x_14722 = x_3481 & x_3482;
assign x_14723 = x_3480 & x_14722;
assign x_14724 = x_14721 & x_14723;
assign x_14725 = x_14719 & x_14724;
assign x_14726 = x_3483 & x_3484;
assign x_14727 = x_3486 & x_3487;
assign x_14728 = x_3485 & x_14727;
assign x_14729 = x_14726 & x_14728;
assign x_14730 = x_3489 & x_3490;
assign x_14731 = x_3488 & x_14730;
assign x_14732 = x_3492 & x_3493;
assign x_14733 = x_3491 & x_14732;
assign x_14734 = x_14731 & x_14733;
assign x_14735 = x_14729 & x_14734;
assign x_14736 = x_14725 & x_14735;
assign x_14737 = x_3494 & x_3495;
assign x_14738 = x_3497 & x_3498;
assign x_14739 = x_3496 & x_14738;
assign x_14740 = x_14737 & x_14739;
assign x_14741 = x_3500 & x_3501;
assign x_14742 = x_3499 & x_14741;
assign x_14743 = x_3503 & x_3504;
assign x_14744 = x_3502 & x_14743;
assign x_14745 = x_14742 & x_14744;
assign x_14746 = x_14740 & x_14745;
assign x_14747 = x_3505 & x_3506;
assign x_14748 = x_3508 & x_3509;
assign x_14749 = x_3507 & x_14748;
assign x_14750 = x_14747 & x_14749;
assign x_14751 = x_3511 & x_3512;
assign x_14752 = x_3510 & x_14751;
assign x_14753 = x_3514 & x_3515;
assign x_14754 = x_3513 & x_14753;
assign x_14755 = x_14752 & x_14754;
assign x_14756 = x_14750 & x_14755;
assign x_14757 = x_14746 & x_14756;
assign x_14758 = x_14736 & x_14757;
assign x_14759 = x_14715 & x_14758;
assign x_14760 = x_14672 & x_14759;
assign x_14761 = x_14585 & x_14760;
assign x_14762 = x_14410 & x_14761;
assign x_14763 = x_3516 & x_3517;
assign x_14764 = x_3519 & x_3520;
assign x_14765 = x_3518 & x_14764;
assign x_14766 = x_14763 & x_14765;
assign x_14767 = x_3521 & x_3522;
assign x_14768 = x_3524 & x_3525;
assign x_14769 = x_3523 & x_14768;
assign x_14770 = x_14767 & x_14769;
assign x_14771 = x_14766 & x_14770;
assign x_14772 = x_3526 & x_3527;
assign x_14773 = x_3529 & x_3530;
assign x_14774 = x_3528 & x_14773;
assign x_14775 = x_14772 & x_14774;
assign x_14776 = x_3532 & x_3533;
assign x_14777 = x_3531 & x_14776;
assign x_14778 = x_3535 & x_3536;
assign x_14779 = x_3534 & x_14778;
assign x_14780 = x_14777 & x_14779;
assign x_14781 = x_14775 & x_14780;
assign x_14782 = x_14771 & x_14781;
assign x_14783 = x_3537 & x_3538;
assign x_14784 = x_3540 & x_3541;
assign x_14785 = x_3539 & x_14784;
assign x_14786 = x_14783 & x_14785;
assign x_14787 = x_3543 & x_3544;
assign x_14788 = x_3542 & x_14787;
assign x_14789 = x_3546 & x_3547;
assign x_14790 = x_3545 & x_14789;
assign x_14791 = x_14788 & x_14790;
assign x_14792 = x_14786 & x_14791;
assign x_14793 = x_3548 & x_3549;
assign x_14794 = x_3551 & x_3552;
assign x_14795 = x_3550 & x_14794;
assign x_14796 = x_14793 & x_14795;
assign x_14797 = x_3554 & x_3555;
assign x_14798 = x_3553 & x_14797;
assign x_14799 = x_3557 & x_3558;
assign x_14800 = x_3556 & x_14799;
assign x_14801 = x_14798 & x_14800;
assign x_14802 = x_14796 & x_14801;
assign x_14803 = x_14792 & x_14802;
assign x_14804 = x_14782 & x_14803;
assign x_14805 = x_3559 & x_3560;
assign x_14806 = x_3562 & x_3563;
assign x_14807 = x_3561 & x_14806;
assign x_14808 = x_14805 & x_14807;
assign x_14809 = x_3565 & x_3566;
assign x_14810 = x_3564 & x_14809;
assign x_14811 = x_3568 & x_3569;
assign x_14812 = x_3567 & x_14811;
assign x_14813 = x_14810 & x_14812;
assign x_14814 = x_14808 & x_14813;
assign x_14815 = x_3570 & x_3571;
assign x_14816 = x_3573 & x_3574;
assign x_14817 = x_3572 & x_14816;
assign x_14818 = x_14815 & x_14817;
assign x_14819 = x_3576 & x_3577;
assign x_14820 = x_3575 & x_14819;
assign x_14821 = x_3579 & x_3580;
assign x_14822 = x_3578 & x_14821;
assign x_14823 = x_14820 & x_14822;
assign x_14824 = x_14818 & x_14823;
assign x_14825 = x_14814 & x_14824;
assign x_14826 = x_3581 & x_3582;
assign x_14827 = x_3584 & x_3585;
assign x_14828 = x_3583 & x_14827;
assign x_14829 = x_14826 & x_14828;
assign x_14830 = x_3587 & x_3588;
assign x_14831 = x_3586 & x_14830;
assign x_14832 = x_3590 & x_3591;
assign x_14833 = x_3589 & x_14832;
assign x_14834 = x_14831 & x_14833;
assign x_14835 = x_14829 & x_14834;
assign x_14836 = x_3592 & x_3593;
assign x_14837 = x_3595 & x_3596;
assign x_14838 = x_3594 & x_14837;
assign x_14839 = x_14836 & x_14838;
assign x_14840 = x_3598 & x_3599;
assign x_14841 = x_3597 & x_14840;
assign x_14842 = x_3601 & x_3602;
assign x_14843 = x_3600 & x_14842;
assign x_14844 = x_14841 & x_14843;
assign x_14845 = x_14839 & x_14844;
assign x_14846 = x_14835 & x_14845;
assign x_14847 = x_14825 & x_14846;
assign x_14848 = x_14804 & x_14847;
assign x_14849 = x_3603 & x_3604;
assign x_14850 = x_3606 & x_3607;
assign x_14851 = x_3605 & x_14850;
assign x_14852 = x_14849 & x_14851;
assign x_14853 = x_3609 & x_3610;
assign x_14854 = x_3608 & x_14853;
assign x_14855 = x_3612 & x_3613;
assign x_14856 = x_3611 & x_14855;
assign x_14857 = x_14854 & x_14856;
assign x_14858 = x_14852 & x_14857;
assign x_14859 = x_3614 & x_3615;
assign x_14860 = x_3617 & x_3618;
assign x_14861 = x_3616 & x_14860;
assign x_14862 = x_14859 & x_14861;
assign x_14863 = x_3620 & x_3621;
assign x_14864 = x_3619 & x_14863;
assign x_14865 = x_3623 & x_3624;
assign x_14866 = x_3622 & x_14865;
assign x_14867 = x_14864 & x_14866;
assign x_14868 = x_14862 & x_14867;
assign x_14869 = x_14858 & x_14868;
assign x_14870 = x_3625 & x_3626;
assign x_14871 = x_3628 & x_3629;
assign x_14872 = x_3627 & x_14871;
assign x_14873 = x_14870 & x_14872;
assign x_14874 = x_3631 & x_3632;
assign x_14875 = x_3630 & x_14874;
assign x_14876 = x_3634 & x_3635;
assign x_14877 = x_3633 & x_14876;
assign x_14878 = x_14875 & x_14877;
assign x_14879 = x_14873 & x_14878;
assign x_14880 = x_3636 & x_3637;
assign x_14881 = x_3639 & x_3640;
assign x_14882 = x_3638 & x_14881;
assign x_14883 = x_14880 & x_14882;
assign x_14884 = x_3642 & x_3643;
assign x_14885 = x_3641 & x_14884;
assign x_14886 = x_3645 & x_3646;
assign x_14887 = x_3644 & x_14886;
assign x_14888 = x_14885 & x_14887;
assign x_14889 = x_14883 & x_14888;
assign x_14890 = x_14879 & x_14889;
assign x_14891 = x_14869 & x_14890;
assign x_14892 = x_3647 & x_3648;
assign x_14893 = x_3650 & x_3651;
assign x_14894 = x_3649 & x_14893;
assign x_14895 = x_14892 & x_14894;
assign x_14896 = x_3653 & x_3654;
assign x_14897 = x_3652 & x_14896;
assign x_14898 = x_3656 & x_3657;
assign x_14899 = x_3655 & x_14898;
assign x_14900 = x_14897 & x_14899;
assign x_14901 = x_14895 & x_14900;
assign x_14902 = x_3658 & x_3659;
assign x_14903 = x_3661 & x_3662;
assign x_14904 = x_3660 & x_14903;
assign x_14905 = x_14902 & x_14904;
assign x_14906 = x_3664 & x_3665;
assign x_14907 = x_3663 & x_14906;
assign x_14908 = x_3667 & x_3668;
assign x_14909 = x_3666 & x_14908;
assign x_14910 = x_14907 & x_14909;
assign x_14911 = x_14905 & x_14910;
assign x_14912 = x_14901 & x_14911;
assign x_14913 = x_3669 & x_3670;
assign x_14914 = x_3672 & x_3673;
assign x_14915 = x_3671 & x_14914;
assign x_14916 = x_14913 & x_14915;
assign x_14917 = x_3675 & x_3676;
assign x_14918 = x_3674 & x_14917;
assign x_14919 = x_3678 & x_3679;
assign x_14920 = x_3677 & x_14919;
assign x_14921 = x_14918 & x_14920;
assign x_14922 = x_14916 & x_14921;
assign x_14923 = x_3680 & x_3681;
assign x_14924 = x_3683 & x_3684;
assign x_14925 = x_3682 & x_14924;
assign x_14926 = x_14923 & x_14925;
assign x_14927 = x_3686 & x_3687;
assign x_14928 = x_3685 & x_14927;
assign x_14929 = x_3689 & x_3690;
assign x_14930 = x_3688 & x_14929;
assign x_14931 = x_14928 & x_14930;
assign x_14932 = x_14926 & x_14931;
assign x_14933 = x_14922 & x_14932;
assign x_14934 = x_14912 & x_14933;
assign x_14935 = x_14891 & x_14934;
assign x_14936 = x_14848 & x_14935;
assign x_14937 = x_3691 & x_3692;
assign x_14938 = x_3694 & x_3695;
assign x_14939 = x_3693 & x_14938;
assign x_14940 = x_14937 & x_14939;
assign x_14941 = x_3697 & x_3698;
assign x_14942 = x_3696 & x_14941;
assign x_14943 = x_3700 & x_3701;
assign x_14944 = x_3699 & x_14943;
assign x_14945 = x_14942 & x_14944;
assign x_14946 = x_14940 & x_14945;
assign x_14947 = x_3702 & x_3703;
assign x_14948 = x_3705 & x_3706;
assign x_14949 = x_3704 & x_14948;
assign x_14950 = x_14947 & x_14949;
assign x_14951 = x_3708 & x_3709;
assign x_14952 = x_3707 & x_14951;
assign x_14953 = x_3711 & x_3712;
assign x_14954 = x_3710 & x_14953;
assign x_14955 = x_14952 & x_14954;
assign x_14956 = x_14950 & x_14955;
assign x_14957 = x_14946 & x_14956;
assign x_14958 = x_3713 & x_3714;
assign x_14959 = x_3716 & x_3717;
assign x_14960 = x_3715 & x_14959;
assign x_14961 = x_14958 & x_14960;
assign x_14962 = x_3719 & x_3720;
assign x_14963 = x_3718 & x_14962;
assign x_14964 = x_3722 & x_3723;
assign x_14965 = x_3721 & x_14964;
assign x_14966 = x_14963 & x_14965;
assign x_14967 = x_14961 & x_14966;
assign x_14968 = x_3724 & x_3725;
assign x_14969 = x_3727 & x_3728;
assign x_14970 = x_3726 & x_14969;
assign x_14971 = x_14968 & x_14970;
assign x_14972 = x_3730 & x_3731;
assign x_14973 = x_3729 & x_14972;
assign x_14974 = x_3733 & x_3734;
assign x_14975 = x_3732 & x_14974;
assign x_14976 = x_14973 & x_14975;
assign x_14977 = x_14971 & x_14976;
assign x_14978 = x_14967 & x_14977;
assign x_14979 = x_14957 & x_14978;
assign x_14980 = x_3735 & x_3736;
assign x_14981 = x_3738 & x_3739;
assign x_14982 = x_3737 & x_14981;
assign x_14983 = x_14980 & x_14982;
assign x_14984 = x_3741 & x_3742;
assign x_14985 = x_3740 & x_14984;
assign x_14986 = x_3744 & x_3745;
assign x_14987 = x_3743 & x_14986;
assign x_14988 = x_14985 & x_14987;
assign x_14989 = x_14983 & x_14988;
assign x_14990 = x_3746 & x_3747;
assign x_14991 = x_3749 & x_3750;
assign x_14992 = x_3748 & x_14991;
assign x_14993 = x_14990 & x_14992;
assign x_14994 = x_3752 & x_3753;
assign x_14995 = x_3751 & x_14994;
assign x_14996 = x_3755 & x_3756;
assign x_14997 = x_3754 & x_14996;
assign x_14998 = x_14995 & x_14997;
assign x_14999 = x_14993 & x_14998;
assign x_15000 = x_14989 & x_14999;
assign x_15001 = x_3757 & x_3758;
assign x_15002 = x_3760 & x_3761;
assign x_15003 = x_3759 & x_15002;
assign x_15004 = x_15001 & x_15003;
assign x_15005 = x_3763 & x_3764;
assign x_15006 = x_3762 & x_15005;
assign x_15007 = x_3766 & x_3767;
assign x_15008 = x_3765 & x_15007;
assign x_15009 = x_15006 & x_15008;
assign x_15010 = x_15004 & x_15009;
assign x_15011 = x_3768 & x_3769;
assign x_15012 = x_3771 & x_3772;
assign x_15013 = x_3770 & x_15012;
assign x_15014 = x_15011 & x_15013;
assign x_15015 = x_3774 & x_3775;
assign x_15016 = x_3773 & x_15015;
assign x_15017 = x_3777 & x_3778;
assign x_15018 = x_3776 & x_15017;
assign x_15019 = x_15016 & x_15018;
assign x_15020 = x_15014 & x_15019;
assign x_15021 = x_15010 & x_15020;
assign x_15022 = x_15000 & x_15021;
assign x_15023 = x_14979 & x_15022;
assign x_15024 = x_3779 & x_3780;
assign x_15025 = x_3782 & x_3783;
assign x_15026 = x_3781 & x_15025;
assign x_15027 = x_15024 & x_15026;
assign x_15028 = x_3785 & x_3786;
assign x_15029 = x_3784 & x_15028;
assign x_15030 = x_3788 & x_3789;
assign x_15031 = x_3787 & x_15030;
assign x_15032 = x_15029 & x_15031;
assign x_15033 = x_15027 & x_15032;
assign x_15034 = x_3790 & x_3791;
assign x_15035 = x_3793 & x_3794;
assign x_15036 = x_3792 & x_15035;
assign x_15037 = x_15034 & x_15036;
assign x_15038 = x_3796 & x_3797;
assign x_15039 = x_3795 & x_15038;
assign x_15040 = x_3799 & x_3800;
assign x_15041 = x_3798 & x_15040;
assign x_15042 = x_15039 & x_15041;
assign x_15043 = x_15037 & x_15042;
assign x_15044 = x_15033 & x_15043;
assign x_15045 = x_3801 & x_3802;
assign x_15046 = x_3804 & x_3805;
assign x_15047 = x_3803 & x_15046;
assign x_15048 = x_15045 & x_15047;
assign x_15049 = x_3807 & x_3808;
assign x_15050 = x_3806 & x_15049;
assign x_15051 = x_3810 & x_3811;
assign x_15052 = x_3809 & x_15051;
assign x_15053 = x_15050 & x_15052;
assign x_15054 = x_15048 & x_15053;
assign x_15055 = x_3812 & x_3813;
assign x_15056 = x_3815 & x_3816;
assign x_15057 = x_3814 & x_15056;
assign x_15058 = x_15055 & x_15057;
assign x_15059 = x_3818 & x_3819;
assign x_15060 = x_3817 & x_15059;
assign x_15061 = x_3821 & x_3822;
assign x_15062 = x_3820 & x_15061;
assign x_15063 = x_15060 & x_15062;
assign x_15064 = x_15058 & x_15063;
assign x_15065 = x_15054 & x_15064;
assign x_15066 = x_15044 & x_15065;
assign x_15067 = x_3823 & x_3824;
assign x_15068 = x_3826 & x_3827;
assign x_15069 = x_3825 & x_15068;
assign x_15070 = x_15067 & x_15069;
assign x_15071 = x_3829 & x_3830;
assign x_15072 = x_3828 & x_15071;
assign x_15073 = x_3832 & x_3833;
assign x_15074 = x_3831 & x_15073;
assign x_15075 = x_15072 & x_15074;
assign x_15076 = x_15070 & x_15075;
assign x_15077 = x_3834 & x_3835;
assign x_15078 = x_3837 & x_3838;
assign x_15079 = x_3836 & x_15078;
assign x_15080 = x_15077 & x_15079;
assign x_15081 = x_3840 & x_3841;
assign x_15082 = x_3839 & x_15081;
assign x_15083 = x_3843 & x_3844;
assign x_15084 = x_3842 & x_15083;
assign x_15085 = x_15082 & x_15084;
assign x_15086 = x_15080 & x_15085;
assign x_15087 = x_15076 & x_15086;
assign x_15088 = x_3845 & x_3846;
assign x_15089 = x_3848 & x_3849;
assign x_15090 = x_3847 & x_15089;
assign x_15091 = x_15088 & x_15090;
assign x_15092 = x_3851 & x_3852;
assign x_15093 = x_3850 & x_15092;
assign x_15094 = x_3854 & x_3855;
assign x_15095 = x_3853 & x_15094;
assign x_15096 = x_15093 & x_15095;
assign x_15097 = x_15091 & x_15096;
assign x_15098 = x_3856 & x_3857;
assign x_15099 = x_3859 & x_3860;
assign x_15100 = x_3858 & x_15099;
assign x_15101 = x_15098 & x_15100;
assign x_15102 = x_3862 & x_3863;
assign x_15103 = x_3861 & x_15102;
assign x_15104 = x_3865 & x_3866;
assign x_15105 = x_3864 & x_15104;
assign x_15106 = x_15103 & x_15105;
assign x_15107 = x_15101 & x_15106;
assign x_15108 = x_15097 & x_15107;
assign x_15109 = x_15087 & x_15108;
assign x_15110 = x_15066 & x_15109;
assign x_15111 = x_15023 & x_15110;
assign x_15112 = x_14936 & x_15111;
assign x_15113 = x_3867 & x_3868;
assign x_15114 = x_3870 & x_3871;
assign x_15115 = x_3869 & x_15114;
assign x_15116 = x_15113 & x_15115;
assign x_15117 = x_3873 & x_3874;
assign x_15118 = x_3872 & x_15117;
assign x_15119 = x_3876 & x_3877;
assign x_15120 = x_3875 & x_15119;
assign x_15121 = x_15118 & x_15120;
assign x_15122 = x_15116 & x_15121;
assign x_15123 = x_3878 & x_3879;
assign x_15124 = x_3881 & x_3882;
assign x_15125 = x_3880 & x_15124;
assign x_15126 = x_15123 & x_15125;
assign x_15127 = x_3884 & x_3885;
assign x_15128 = x_3883 & x_15127;
assign x_15129 = x_3887 & x_3888;
assign x_15130 = x_3886 & x_15129;
assign x_15131 = x_15128 & x_15130;
assign x_15132 = x_15126 & x_15131;
assign x_15133 = x_15122 & x_15132;
assign x_15134 = x_3889 & x_3890;
assign x_15135 = x_3892 & x_3893;
assign x_15136 = x_3891 & x_15135;
assign x_15137 = x_15134 & x_15136;
assign x_15138 = x_3895 & x_3896;
assign x_15139 = x_3894 & x_15138;
assign x_15140 = x_3898 & x_3899;
assign x_15141 = x_3897 & x_15140;
assign x_15142 = x_15139 & x_15141;
assign x_15143 = x_15137 & x_15142;
assign x_15144 = x_3900 & x_3901;
assign x_15145 = x_3903 & x_3904;
assign x_15146 = x_3902 & x_15145;
assign x_15147 = x_15144 & x_15146;
assign x_15148 = x_3906 & x_3907;
assign x_15149 = x_3905 & x_15148;
assign x_15150 = x_3909 & x_3910;
assign x_15151 = x_3908 & x_15150;
assign x_15152 = x_15149 & x_15151;
assign x_15153 = x_15147 & x_15152;
assign x_15154 = x_15143 & x_15153;
assign x_15155 = x_15133 & x_15154;
assign x_15156 = x_3911 & x_3912;
assign x_15157 = x_3914 & x_3915;
assign x_15158 = x_3913 & x_15157;
assign x_15159 = x_15156 & x_15158;
assign x_15160 = x_3917 & x_3918;
assign x_15161 = x_3916 & x_15160;
assign x_15162 = x_3920 & x_3921;
assign x_15163 = x_3919 & x_15162;
assign x_15164 = x_15161 & x_15163;
assign x_15165 = x_15159 & x_15164;
assign x_15166 = x_3922 & x_3923;
assign x_15167 = x_3925 & x_3926;
assign x_15168 = x_3924 & x_15167;
assign x_15169 = x_15166 & x_15168;
assign x_15170 = x_3928 & x_3929;
assign x_15171 = x_3927 & x_15170;
assign x_15172 = x_3931 & x_3932;
assign x_15173 = x_3930 & x_15172;
assign x_15174 = x_15171 & x_15173;
assign x_15175 = x_15169 & x_15174;
assign x_15176 = x_15165 & x_15175;
assign x_15177 = x_3933 & x_3934;
assign x_15178 = x_3936 & x_3937;
assign x_15179 = x_3935 & x_15178;
assign x_15180 = x_15177 & x_15179;
assign x_15181 = x_3939 & x_3940;
assign x_15182 = x_3938 & x_15181;
assign x_15183 = x_3942 & x_3943;
assign x_15184 = x_3941 & x_15183;
assign x_15185 = x_15182 & x_15184;
assign x_15186 = x_15180 & x_15185;
assign x_15187 = x_3944 & x_3945;
assign x_15188 = x_3947 & x_3948;
assign x_15189 = x_3946 & x_15188;
assign x_15190 = x_15187 & x_15189;
assign x_15191 = x_3950 & x_3951;
assign x_15192 = x_3949 & x_15191;
assign x_15193 = x_3953 & x_3954;
assign x_15194 = x_3952 & x_15193;
assign x_15195 = x_15192 & x_15194;
assign x_15196 = x_15190 & x_15195;
assign x_15197 = x_15186 & x_15196;
assign x_15198 = x_15176 & x_15197;
assign x_15199 = x_15155 & x_15198;
assign x_15200 = x_3955 & x_3956;
assign x_15201 = x_3958 & x_3959;
assign x_15202 = x_3957 & x_15201;
assign x_15203 = x_15200 & x_15202;
assign x_15204 = x_3961 & x_3962;
assign x_15205 = x_3960 & x_15204;
assign x_15206 = x_3964 & x_3965;
assign x_15207 = x_3963 & x_15206;
assign x_15208 = x_15205 & x_15207;
assign x_15209 = x_15203 & x_15208;
assign x_15210 = x_3966 & x_3967;
assign x_15211 = x_3969 & x_3970;
assign x_15212 = x_3968 & x_15211;
assign x_15213 = x_15210 & x_15212;
assign x_15214 = x_3972 & x_3973;
assign x_15215 = x_3971 & x_15214;
assign x_15216 = x_3975 & x_3976;
assign x_15217 = x_3974 & x_15216;
assign x_15218 = x_15215 & x_15217;
assign x_15219 = x_15213 & x_15218;
assign x_15220 = x_15209 & x_15219;
assign x_15221 = x_3977 & x_3978;
assign x_15222 = x_3980 & x_3981;
assign x_15223 = x_3979 & x_15222;
assign x_15224 = x_15221 & x_15223;
assign x_15225 = x_3983 & x_3984;
assign x_15226 = x_3982 & x_15225;
assign x_15227 = x_3986 & x_3987;
assign x_15228 = x_3985 & x_15227;
assign x_15229 = x_15226 & x_15228;
assign x_15230 = x_15224 & x_15229;
assign x_15231 = x_3988 & x_3989;
assign x_15232 = x_3991 & x_3992;
assign x_15233 = x_3990 & x_15232;
assign x_15234 = x_15231 & x_15233;
assign x_15235 = x_3994 & x_3995;
assign x_15236 = x_3993 & x_15235;
assign x_15237 = x_3997 & x_3998;
assign x_15238 = x_3996 & x_15237;
assign x_15239 = x_15236 & x_15238;
assign x_15240 = x_15234 & x_15239;
assign x_15241 = x_15230 & x_15240;
assign x_15242 = x_15220 & x_15241;
assign x_15243 = x_3999 & x_4000;
assign x_15244 = x_4002 & x_4003;
assign x_15245 = x_4001 & x_15244;
assign x_15246 = x_15243 & x_15245;
assign x_15247 = x_4005 & x_4006;
assign x_15248 = x_4004 & x_15247;
assign x_15249 = x_4008 & x_4009;
assign x_15250 = x_4007 & x_15249;
assign x_15251 = x_15248 & x_15250;
assign x_15252 = x_15246 & x_15251;
assign x_15253 = x_4010 & x_4011;
assign x_15254 = x_4013 & x_4014;
assign x_15255 = x_4012 & x_15254;
assign x_15256 = x_15253 & x_15255;
assign x_15257 = x_4016 & x_4017;
assign x_15258 = x_4015 & x_15257;
assign x_15259 = x_4019 & x_4020;
assign x_15260 = x_4018 & x_15259;
assign x_15261 = x_15258 & x_15260;
assign x_15262 = x_15256 & x_15261;
assign x_15263 = x_15252 & x_15262;
assign x_15264 = x_4021 & x_4022;
assign x_15265 = x_4024 & x_4025;
assign x_15266 = x_4023 & x_15265;
assign x_15267 = x_15264 & x_15266;
assign x_15268 = x_4027 & x_4028;
assign x_15269 = x_4026 & x_15268;
assign x_15270 = x_4030 & x_4031;
assign x_15271 = x_4029 & x_15270;
assign x_15272 = x_15269 & x_15271;
assign x_15273 = x_15267 & x_15272;
assign x_15274 = x_4032 & x_4033;
assign x_15275 = x_4035 & x_4036;
assign x_15276 = x_4034 & x_15275;
assign x_15277 = x_15274 & x_15276;
assign x_15278 = x_4038 & x_4039;
assign x_15279 = x_4037 & x_15278;
assign x_15280 = x_4041 & x_4042;
assign x_15281 = x_4040 & x_15280;
assign x_15282 = x_15279 & x_15281;
assign x_15283 = x_15277 & x_15282;
assign x_15284 = x_15273 & x_15283;
assign x_15285 = x_15263 & x_15284;
assign x_15286 = x_15242 & x_15285;
assign x_15287 = x_15199 & x_15286;
assign x_15288 = x_4043 & x_4044;
assign x_15289 = x_4046 & x_4047;
assign x_15290 = x_4045 & x_15289;
assign x_15291 = x_15288 & x_15290;
assign x_15292 = x_4049 & x_4050;
assign x_15293 = x_4048 & x_15292;
assign x_15294 = x_4052 & x_4053;
assign x_15295 = x_4051 & x_15294;
assign x_15296 = x_15293 & x_15295;
assign x_15297 = x_15291 & x_15296;
assign x_15298 = x_4054 & x_4055;
assign x_15299 = x_4057 & x_4058;
assign x_15300 = x_4056 & x_15299;
assign x_15301 = x_15298 & x_15300;
assign x_15302 = x_4060 & x_4061;
assign x_15303 = x_4059 & x_15302;
assign x_15304 = x_4063 & x_4064;
assign x_15305 = x_4062 & x_15304;
assign x_15306 = x_15303 & x_15305;
assign x_15307 = x_15301 & x_15306;
assign x_15308 = x_15297 & x_15307;
assign x_15309 = x_4065 & x_4066;
assign x_15310 = x_4068 & x_4069;
assign x_15311 = x_4067 & x_15310;
assign x_15312 = x_15309 & x_15311;
assign x_15313 = x_4071 & x_4072;
assign x_15314 = x_4070 & x_15313;
assign x_15315 = x_4074 & x_4075;
assign x_15316 = x_4073 & x_15315;
assign x_15317 = x_15314 & x_15316;
assign x_15318 = x_15312 & x_15317;
assign x_15319 = x_4076 & x_4077;
assign x_15320 = x_4079 & x_4080;
assign x_15321 = x_4078 & x_15320;
assign x_15322 = x_15319 & x_15321;
assign x_15323 = x_4082 & x_4083;
assign x_15324 = x_4081 & x_15323;
assign x_15325 = x_4085 & x_4086;
assign x_15326 = x_4084 & x_15325;
assign x_15327 = x_15324 & x_15326;
assign x_15328 = x_15322 & x_15327;
assign x_15329 = x_15318 & x_15328;
assign x_15330 = x_15308 & x_15329;
assign x_15331 = x_4087 & x_4088;
assign x_15332 = x_4090 & x_4091;
assign x_15333 = x_4089 & x_15332;
assign x_15334 = x_15331 & x_15333;
assign x_15335 = x_4093 & x_4094;
assign x_15336 = x_4092 & x_15335;
assign x_15337 = x_4096 & x_4097;
assign x_15338 = x_4095 & x_15337;
assign x_15339 = x_15336 & x_15338;
assign x_15340 = x_15334 & x_15339;
assign x_15341 = x_4098 & x_4099;
assign x_15342 = x_4101 & x_4102;
assign x_15343 = x_4100 & x_15342;
assign x_15344 = x_15341 & x_15343;
assign x_15345 = x_4104 & x_4105;
assign x_15346 = x_4103 & x_15345;
assign x_15347 = x_4107 & x_4108;
assign x_15348 = x_4106 & x_15347;
assign x_15349 = x_15346 & x_15348;
assign x_15350 = x_15344 & x_15349;
assign x_15351 = x_15340 & x_15350;
assign x_15352 = x_4109 & x_4110;
assign x_15353 = x_4112 & x_4113;
assign x_15354 = x_4111 & x_15353;
assign x_15355 = x_15352 & x_15354;
assign x_15356 = x_4115 & x_4116;
assign x_15357 = x_4114 & x_15356;
assign x_15358 = x_4118 & x_4119;
assign x_15359 = x_4117 & x_15358;
assign x_15360 = x_15357 & x_15359;
assign x_15361 = x_15355 & x_15360;
assign x_15362 = x_4120 & x_4121;
assign x_15363 = x_4123 & x_4124;
assign x_15364 = x_4122 & x_15363;
assign x_15365 = x_15362 & x_15364;
assign x_15366 = x_4126 & x_4127;
assign x_15367 = x_4125 & x_15366;
assign x_15368 = x_4129 & x_4130;
assign x_15369 = x_4128 & x_15368;
assign x_15370 = x_15367 & x_15369;
assign x_15371 = x_15365 & x_15370;
assign x_15372 = x_15361 & x_15371;
assign x_15373 = x_15351 & x_15372;
assign x_15374 = x_15330 & x_15373;
assign x_15375 = x_4131 & x_4132;
assign x_15376 = x_4134 & x_4135;
assign x_15377 = x_4133 & x_15376;
assign x_15378 = x_15375 & x_15377;
assign x_15379 = x_4137 & x_4138;
assign x_15380 = x_4136 & x_15379;
assign x_15381 = x_4140 & x_4141;
assign x_15382 = x_4139 & x_15381;
assign x_15383 = x_15380 & x_15382;
assign x_15384 = x_15378 & x_15383;
assign x_15385 = x_4142 & x_4143;
assign x_15386 = x_4145 & x_4146;
assign x_15387 = x_4144 & x_15386;
assign x_15388 = x_15385 & x_15387;
assign x_15389 = x_4148 & x_4149;
assign x_15390 = x_4147 & x_15389;
assign x_15391 = x_4151 & x_4152;
assign x_15392 = x_4150 & x_15391;
assign x_15393 = x_15390 & x_15392;
assign x_15394 = x_15388 & x_15393;
assign x_15395 = x_15384 & x_15394;
assign x_15396 = x_4153 & x_4154;
assign x_15397 = x_4156 & x_4157;
assign x_15398 = x_4155 & x_15397;
assign x_15399 = x_15396 & x_15398;
assign x_15400 = x_4159 & x_4160;
assign x_15401 = x_4158 & x_15400;
assign x_15402 = x_4162 & x_4163;
assign x_15403 = x_4161 & x_15402;
assign x_15404 = x_15401 & x_15403;
assign x_15405 = x_15399 & x_15404;
assign x_15406 = x_4164 & x_4165;
assign x_15407 = x_4167 & x_4168;
assign x_15408 = x_4166 & x_15407;
assign x_15409 = x_15406 & x_15408;
assign x_15410 = x_4170 & x_4171;
assign x_15411 = x_4169 & x_15410;
assign x_15412 = x_4173 & x_4174;
assign x_15413 = x_4172 & x_15412;
assign x_15414 = x_15411 & x_15413;
assign x_15415 = x_15409 & x_15414;
assign x_15416 = x_15405 & x_15415;
assign x_15417 = x_15395 & x_15416;
assign x_15418 = x_4175 & x_4176;
assign x_15419 = x_4178 & x_4179;
assign x_15420 = x_4177 & x_15419;
assign x_15421 = x_15418 & x_15420;
assign x_15422 = x_4181 & x_4182;
assign x_15423 = x_4180 & x_15422;
assign x_15424 = x_4184 & x_4185;
assign x_15425 = x_4183 & x_15424;
assign x_15426 = x_15423 & x_15425;
assign x_15427 = x_15421 & x_15426;
assign x_15428 = x_4186 & x_4187;
assign x_15429 = x_4189 & x_4190;
assign x_15430 = x_4188 & x_15429;
assign x_15431 = x_15428 & x_15430;
assign x_15432 = x_4192 & x_4193;
assign x_15433 = x_4191 & x_15432;
assign x_15434 = x_4195 & x_4196;
assign x_15435 = x_4194 & x_15434;
assign x_15436 = x_15433 & x_15435;
assign x_15437 = x_15431 & x_15436;
assign x_15438 = x_15427 & x_15437;
assign x_15439 = x_4197 & x_4198;
assign x_15440 = x_4200 & x_4201;
assign x_15441 = x_4199 & x_15440;
assign x_15442 = x_15439 & x_15441;
assign x_15443 = x_4203 & x_4204;
assign x_15444 = x_4202 & x_15443;
assign x_15445 = x_4206 & x_4207;
assign x_15446 = x_4205 & x_15445;
assign x_15447 = x_15444 & x_15446;
assign x_15448 = x_15442 & x_15447;
assign x_15449 = x_4208 & x_4209;
assign x_15450 = x_4211 & x_4212;
assign x_15451 = x_4210 & x_15450;
assign x_15452 = x_15449 & x_15451;
assign x_15453 = x_4214 & x_4215;
assign x_15454 = x_4213 & x_15453;
assign x_15455 = x_4217 & x_4218;
assign x_15456 = x_4216 & x_15455;
assign x_15457 = x_15454 & x_15456;
assign x_15458 = x_15452 & x_15457;
assign x_15459 = x_15448 & x_15458;
assign x_15460 = x_15438 & x_15459;
assign x_15461 = x_15417 & x_15460;
assign x_15462 = x_15374 & x_15461;
assign x_15463 = x_15287 & x_15462;
assign x_15464 = x_15112 & x_15463;
assign x_15465 = x_14762 & x_15464;
assign x_15466 = x_4219 & x_4220;
assign x_15467 = x_4222 & x_4223;
assign x_15468 = x_4221 & x_15467;
assign x_15469 = x_15466 & x_15468;
assign x_15470 = x_4224 & x_4225;
assign x_15471 = x_4227 & x_4228;
assign x_15472 = x_4226 & x_15471;
assign x_15473 = x_15470 & x_15472;
assign x_15474 = x_15469 & x_15473;
assign x_15475 = x_4229 & x_4230;
assign x_15476 = x_4232 & x_4233;
assign x_15477 = x_4231 & x_15476;
assign x_15478 = x_15475 & x_15477;
assign x_15479 = x_4235 & x_4236;
assign x_15480 = x_4234 & x_15479;
assign x_15481 = x_4238 & x_4239;
assign x_15482 = x_4237 & x_15481;
assign x_15483 = x_15480 & x_15482;
assign x_15484 = x_15478 & x_15483;
assign x_15485 = x_15474 & x_15484;
assign x_15486 = x_4240 & x_4241;
assign x_15487 = x_4243 & x_4244;
assign x_15488 = x_4242 & x_15487;
assign x_15489 = x_15486 & x_15488;
assign x_15490 = x_4246 & x_4247;
assign x_15491 = x_4245 & x_15490;
assign x_15492 = x_4249 & x_4250;
assign x_15493 = x_4248 & x_15492;
assign x_15494 = x_15491 & x_15493;
assign x_15495 = x_15489 & x_15494;
assign x_15496 = x_4251 & x_4252;
assign x_15497 = x_4254 & x_4255;
assign x_15498 = x_4253 & x_15497;
assign x_15499 = x_15496 & x_15498;
assign x_15500 = x_4257 & x_4258;
assign x_15501 = x_4256 & x_15500;
assign x_15502 = x_4260 & x_4261;
assign x_15503 = x_4259 & x_15502;
assign x_15504 = x_15501 & x_15503;
assign x_15505 = x_15499 & x_15504;
assign x_15506 = x_15495 & x_15505;
assign x_15507 = x_15485 & x_15506;
assign x_15508 = x_4262 & x_4263;
assign x_15509 = x_4265 & x_4266;
assign x_15510 = x_4264 & x_15509;
assign x_15511 = x_15508 & x_15510;
assign x_15512 = x_4268 & x_4269;
assign x_15513 = x_4267 & x_15512;
assign x_15514 = x_4271 & x_4272;
assign x_15515 = x_4270 & x_15514;
assign x_15516 = x_15513 & x_15515;
assign x_15517 = x_15511 & x_15516;
assign x_15518 = x_4273 & x_4274;
assign x_15519 = x_4276 & x_4277;
assign x_15520 = x_4275 & x_15519;
assign x_15521 = x_15518 & x_15520;
assign x_15522 = x_4279 & x_4280;
assign x_15523 = x_4278 & x_15522;
assign x_15524 = x_4282 & x_4283;
assign x_15525 = x_4281 & x_15524;
assign x_15526 = x_15523 & x_15525;
assign x_15527 = x_15521 & x_15526;
assign x_15528 = x_15517 & x_15527;
assign x_15529 = x_4284 & x_4285;
assign x_15530 = x_4287 & x_4288;
assign x_15531 = x_4286 & x_15530;
assign x_15532 = x_15529 & x_15531;
assign x_15533 = x_4290 & x_4291;
assign x_15534 = x_4289 & x_15533;
assign x_15535 = x_4293 & x_4294;
assign x_15536 = x_4292 & x_15535;
assign x_15537 = x_15534 & x_15536;
assign x_15538 = x_15532 & x_15537;
assign x_15539 = x_4295 & x_4296;
assign x_15540 = x_4298 & x_4299;
assign x_15541 = x_4297 & x_15540;
assign x_15542 = x_15539 & x_15541;
assign x_15543 = x_4301 & x_4302;
assign x_15544 = x_4300 & x_15543;
assign x_15545 = x_4304 & x_4305;
assign x_15546 = x_4303 & x_15545;
assign x_15547 = x_15544 & x_15546;
assign x_15548 = x_15542 & x_15547;
assign x_15549 = x_15538 & x_15548;
assign x_15550 = x_15528 & x_15549;
assign x_15551 = x_15507 & x_15550;
assign x_15552 = x_4306 & x_4307;
assign x_15553 = x_4309 & x_4310;
assign x_15554 = x_4308 & x_15553;
assign x_15555 = x_15552 & x_15554;
assign x_15556 = x_4312 & x_4313;
assign x_15557 = x_4311 & x_15556;
assign x_15558 = x_4315 & x_4316;
assign x_15559 = x_4314 & x_15558;
assign x_15560 = x_15557 & x_15559;
assign x_15561 = x_15555 & x_15560;
assign x_15562 = x_4317 & x_4318;
assign x_15563 = x_4320 & x_4321;
assign x_15564 = x_4319 & x_15563;
assign x_15565 = x_15562 & x_15564;
assign x_15566 = x_4323 & x_4324;
assign x_15567 = x_4322 & x_15566;
assign x_15568 = x_4326 & x_4327;
assign x_15569 = x_4325 & x_15568;
assign x_15570 = x_15567 & x_15569;
assign x_15571 = x_15565 & x_15570;
assign x_15572 = x_15561 & x_15571;
assign x_15573 = x_4328 & x_4329;
assign x_15574 = x_4331 & x_4332;
assign x_15575 = x_4330 & x_15574;
assign x_15576 = x_15573 & x_15575;
assign x_15577 = x_4334 & x_4335;
assign x_15578 = x_4333 & x_15577;
assign x_15579 = x_4337 & x_4338;
assign x_15580 = x_4336 & x_15579;
assign x_15581 = x_15578 & x_15580;
assign x_15582 = x_15576 & x_15581;
assign x_15583 = x_4339 & x_4340;
assign x_15584 = x_4342 & x_4343;
assign x_15585 = x_4341 & x_15584;
assign x_15586 = x_15583 & x_15585;
assign x_15587 = x_4345 & x_4346;
assign x_15588 = x_4344 & x_15587;
assign x_15589 = x_4348 & x_4349;
assign x_15590 = x_4347 & x_15589;
assign x_15591 = x_15588 & x_15590;
assign x_15592 = x_15586 & x_15591;
assign x_15593 = x_15582 & x_15592;
assign x_15594 = x_15572 & x_15593;
assign x_15595 = x_4350 & x_4351;
assign x_15596 = x_4353 & x_4354;
assign x_15597 = x_4352 & x_15596;
assign x_15598 = x_15595 & x_15597;
assign x_15599 = x_4356 & x_4357;
assign x_15600 = x_4355 & x_15599;
assign x_15601 = x_4359 & x_4360;
assign x_15602 = x_4358 & x_15601;
assign x_15603 = x_15600 & x_15602;
assign x_15604 = x_15598 & x_15603;
assign x_15605 = x_4361 & x_4362;
assign x_15606 = x_4364 & x_4365;
assign x_15607 = x_4363 & x_15606;
assign x_15608 = x_15605 & x_15607;
assign x_15609 = x_4367 & x_4368;
assign x_15610 = x_4366 & x_15609;
assign x_15611 = x_4370 & x_4371;
assign x_15612 = x_4369 & x_15611;
assign x_15613 = x_15610 & x_15612;
assign x_15614 = x_15608 & x_15613;
assign x_15615 = x_15604 & x_15614;
assign x_15616 = x_4372 & x_4373;
assign x_15617 = x_4375 & x_4376;
assign x_15618 = x_4374 & x_15617;
assign x_15619 = x_15616 & x_15618;
assign x_15620 = x_4378 & x_4379;
assign x_15621 = x_4377 & x_15620;
assign x_15622 = x_4381 & x_4382;
assign x_15623 = x_4380 & x_15622;
assign x_15624 = x_15621 & x_15623;
assign x_15625 = x_15619 & x_15624;
assign x_15626 = x_4383 & x_4384;
assign x_15627 = x_4386 & x_4387;
assign x_15628 = x_4385 & x_15627;
assign x_15629 = x_15626 & x_15628;
assign x_15630 = x_4389 & x_4390;
assign x_15631 = x_4388 & x_15630;
assign x_15632 = x_4392 & x_4393;
assign x_15633 = x_4391 & x_15632;
assign x_15634 = x_15631 & x_15633;
assign x_15635 = x_15629 & x_15634;
assign x_15636 = x_15625 & x_15635;
assign x_15637 = x_15615 & x_15636;
assign x_15638 = x_15594 & x_15637;
assign x_15639 = x_15551 & x_15638;
assign x_15640 = x_4394 & x_4395;
assign x_15641 = x_4397 & x_4398;
assign x_15642 = x_4396 & x_15641;
assign x_15643 = x_15640 & x_15642;
assign x_15644 = x_4400 & x_4401;
assign x_15645 = x_4399 & x_15644;
assign x_15646 = x_4403 & x_4404;
assign x_15647 = x_4402 & x_15646;
assign x_15648 = x_15645 & x_15647;
assign x_15649 = x_15643 & x_15648;
assign x_15650 = x_4405 & x_4406;
assign x_15651 = x_4408 & x_4409;
assign x_15652 = x_4407 & x_15651;
assign x_15653 = x_15650 & x_15652;
assign x_15654 = x_4411 & x_4412;
assign x_15655 = x_4410 & x_15654;
assign x_15656 = x_4414 & x_4415;
assign x_15657 = x_4413 & x_15656;
assign x_15658 = x_15655 & x_15657;
assign x_15659 = x_15653 & x_15658;
assign x_15660 = x_15649 & x_15659;
assign x_15661 = x_4416 & x_4417;
assign x_15662 = x_4419 & x_4420;
assign x_15663 = x_4418 & x_15662;
assign x_15664 = x_15661 & x_15663;
assign x_15665 = x_4422 & x_4423;
assign x_15666 = x_4421 & x_15665;
assign x_15667 = x_4425 & x_4426;
assign x_15668 = x_4424 & x_15667;
assign x_15669 = x_15666 & x_15668;
assign x_15670 = x_15664 & x_15669;
assign x_15671 = x_4427 & x_4428;
assign x_15672 = x_4430 & x_4431;
assign x_15673 = x_4429 & x_15672;
assign x_15674 = x_15671 & x_15673;
assign x_15675 = x_4433 & x_4434;
assign x_15676 = x_4432 & x_15675;
assign x_15677 = x_4436 & x_4437;
assign x_15678 = x_4435 & x_15677;
assign x_15679 = x_15676 & x_15678;
assign x_15680 = x_15674 & x_15679;
assign x_15681 = x_15670 & x_15680;
assign x_15682 = x_15660 & x_15681;
assign x_15683 = x_4438 & x_4439;
assign x_15684 = x_4441 & x_4442;
assign x_15685 = x_4440 & x_15684;
assign x_15686 = x_15683 & x_15685;
assign x_15687 = x_4444 & x_4445;
assign x_15688 = x_4443 & x_15687;
assign x_15689 = x_4447 & x_4448;
assign x_15690 = x_4446 & x_15689;
assign x_15691 = x_15688 & x_15690;
assign x_15692 = x_15686 & x_15691;
assign x_15693 = x_4449 & x_4450;
assign x_15694 = x_4452 & x_4453;
assign x_15695 = x_4451 & x_15694;
assign x_15696 = x_15693 & x_15695;
assign x_15697 = x_4455 & x_4456;
assign x_15698 = x_4454 & x_15697;
assign x_15699 = x_4458 & x_4459;
assign x_15700 = x_4457 & x_15699;
assign x_15701 = x_15698 & x_15700;
assign x_15702 = x_15696 & x_15701;
assign x_15703 = x_15692 & x_15702;
assign x_15704 = x_4460 & x_4461;
assign x_15705 = x_4463 & x_4464;
assign x_15706 = x_4462 & x_15705;
assign x_15707 = x_15704 & x_15706;
assign x_15708 = x_4466 & x_4467;
assign x_15709 = x_4465 & x_15708;
assign x_15710 = x_4469 & x_4470;
assign x_15711 = x_4468 & x_15710;
assign x_15712 = x_15709 & x_15711;
assign x_15713 = x_15707 & x_15712;
assign x_15714 = x_4471 & x_4472;
assign x_15715 = x_4474 & x_4475;
assign x_15716 = x_4473 & x_15715;
assign x_15717 = x_15714 & x_15716;
assign x_15718 = x_4477 & x_4478;
assign x_15719 = x_4476 & x_15718;
assign x_15720 = x_4480 & x_4481;
assign x_15721 = x_4479 & x_15720;
assign x_15722 = x_15719 & x_15721;
assign x_15723 = x_15717 & x_15722;
assign x_15724 = x_15713 & x_15723;
assign x_15725 = x_15703 & x_15724;
assign x_15726 = x_15682 & x_15725;
assign x_15727 = x_4482 & x_4483;
assign x_15728 = x_4485 & x_4486;
assign x_15729 = x_4484 & x_15728;
assign x_15730 = x_15727 & x_15729;
assign x_15731 = x_4488 & x_4489;
assign x_15732 = x_4487 & x_15731;
assign x_15733 = x_4491 & x_4492;
assign x_15734 = x_4490 & x_15733;
assign x_15735 = x_15732 & x_15734;
assign x_15736 = x_15730 & x_15735;
assign x_15737 = x_4493 & x_4494;
assign x_15738 = x_4496 & x_4497;
assign x_15739 = x_4495 & x_15738;
assign x_15740 = x_15737 & x_15739;
assign x_15741 = x_4499 & x_4500;
assign x_15742 = x_4498 & x_15741;
assign x_15743 = x_4502 & x_4503;
assign x_15744 = x_4501 & x_15743;
assign x_15745 = x_15742 & x_15744;
assign x_15746 = x_15740 & x_15745;
assign x_15747 = x_15736 & x_15746;
assign x_15748 = x_4504 & x_4505;
assign x_15749 = x_4507 & x_4508;
assign x_15750 = x_4506 & x_15749;
assign x_15751 = x_15748 & x_15750;
assign x_15752 = x_4510 & x_4511;
assign x_15753 = x_4509 & x_15752;
assign x_15754 = x_4513 & x_4514;
assign x_15755 = x_4512 & x_15754;
assign x_15756 = x_15753 & x_15755;
assign x_15757 = x_15751 & x_15756;
assign x_15758 = x_4515 & x_4516;
assign x_15759 = x_4518 & x_4519;
assign x_15760 = x_4517 & x_15759;
assign x_15761 = x_15758 & x_15760;
assign x_15762 = x_4521 & x_4522;
assign x_15763 = x_4520 & x_15762;
assign x_15764 = x_4524 & x_4525;
assign x_15765 = x_4523 & x_15764;
assign x_15766 = x_15763 & x_15765;
assign x_15767 = x_15761 & x_15766;
assign x_15768 = x_15757 & x_15767;
assign x_15769 = x_15747 & x_15768;
assign x_15770 = x_4526 & x_4527;
assign x_15771 = x_4529 & x_4530;
assign x_15772 = x_4528 & x_15771;
assign x_15773 = x_15770 & x_15772;
assign x_15774 = x_4532 & x_4533;
assign x_15775 = x_4531 & x_15774;
assign x_15776 = x_4535 & x_4536;
assign x_15777 = x_4534 & x_15776;
assign x_15778 = x_15775 & x_15777;
assign x_15779 = x_15773 & x_15778;
assign x_15780 = x_4537 & x_4538;
assign x_15781 = x_4540 & x_4541;
assign x_15782 = x_4539 & x_15781;
assign x_15783 = x_15780 & x_15782;
assign x_15784 = x_4543 & x_4544;
assign x_15785 = x_4542 & x_15784;
assign x_15786 = x_4546 & x_4547;
assign x_15787 = x_4545 & x_15786;
assign x_15788 = x_15785 & x_15787;
assign x_15789 = x_15783 & x_15788;
assign x_15790 = x_15779 & x_15789;
assign x_15791 = x_4548 & x_4549;
assign x_15792 = x_4551 & x_4552;
assign x_15793 = x_4550 & x_15792;
assign x_15794 = x_15791 & x_15793;
assign x_15795 = x_4554 & x_4555;
assign x_15796 = x_4553 & x_15795;
assign x_15797 = x_4557 & x_4558;
assign x_15798 = x_4556 & x_15797;
assign x_15799 = x_15796 & x_15798;
assign x_15800 = x_15794 & x_15799;
assign x_15801 = x_4559 & x_4560;
assign x_15802 = x_4562 & x_4563;
assign x_15803 = x_4561 & x_15802;
assign x_15804 = x_15801 & x_15803;
assign x_15805 = x_4565 & x_4566;
assign x_15806 = x_4564 & x_15805;
assign x_15807 = x_4568 & x_4569;
assign x_15808 = x_4567 & x_15807;
assign x_15809 = x_15806 & x_15808;
assign x_15810 = x_15804 & x_15809;
assign x_15811 = x_15800 & x_15810;
assign x_15812 = x_15790 & x_15811;
assign x_15813 = x_15769 & x_15812;
assign x_15814 = x_15726 & x_15813;
assign x_15815 = x_15639 & x_15814;
assign x_15816 = x_4570 & x_4571;
assign x_15817 = x_4573 & x_4574;
assign x_15818 = x_4572 & x_15817;
assign x_15819 = x_15816 & x_15818;
assign x_15820 = x_4576 & x_4577;
assign x_15821 = x_4575 & x_15820;
assign x_15822 = x_4579 & x_4580;
assign x_15823 = x_4578 & x_15822;
assign x_15824 = x_15821 & x_15823;
assign x_15825 = x_15819 & x_15824;
assign x_15826 = x_4581 & x_4582;
assign x_15827 = x_4584 & x_4585;
assign x_15828 = x_4583 & x_15827;
assign x_15829 = x_15826 & x_15828;
assign x_15830 = x_4587 & x_4588;
assign x_15831 = x_4586 & x_15830;
assign x_15832 = x_4590 & x_4591;
assign x_15833 = x_4589 & x_15832;
assign x_15834 = x_15831 & x_15833;
assign x_15835 = x_15829 & x_15834;
assign x_15836 = x_15825 & x_15835;
assign x_15837 = x_4592 & x_4593;
assign x_15838 = x_4595 & x_4596;
assign x_15839 = x_4594 & x_15838;
assign x_15840 = x_15837 & x_15839;
assign x_15841 = x_4598 & x_4599;
assign x_15842 = x_4597 & x_15841;
assign x_15843 = x_4601 & x_4602;
assign x_15844 = x_4600 & x_15843;
assign x_15845 = x_15842 & x_15844;
assign x_15846 = x_15840 & x_15845;
assign x_15847 = x_4603 & x_4604;
assign x_15848 = x_4606 & x_4607;
assign x_15849 = x_4605 & x_15848;
assign x_15850 = x_15847 & x_15849;
assign x_15851 = x_4609 & x_4610;
assign x_15852 = x_4608 & x_15851;
assign x_15853 = x_4612 & x_4613;
assign x_15854 = x_4611 & x_15853;
assign x_15855 = x_15852 & x_15854;
assign x_15856 = x_15850 & x_15855;
assign x_15857 = x_15846 & x_15856;
assign x_15858 = x_15836 & x_15857;
assign x_15859 = x_4614 & x_4615;
assign x_15860 = x_4617 & x_4618;
assign x_15861 = x_4616 & x_15860;
assign x_15862 = x_15859 & x_15861;
assign x_15863 = x_4620 & x_4621;
assign x_15864 = x_4619 & x_15863;
assign x_15865 = x_4623 & x_4624;
assign x_15866 = x_4622 & x_15865;
assign x_15867 = x_15864 & x_15866;
assign x_15868 = x_15862 & x_15867;
assign x_15869 = x_4625 & x_4626;
assign x_15870 = x_4628 & x_4629;
assign x_15871 = x_4627 & x_15870;
assign x_15872 = x_15869 & x_15871;
assign x_15873 = x_4631 & x_4632;
assign x_15874 = x_4630 & x_15873;
assign x_15875 = x_4634 & x_4635;
assign x_15876 = x_4633 & x_15875;
assign x_15877 = x_15874 & x_15876;
assign x_15878 = x_15872 & x_15877;
assign x_15879 = x_15868 & x_15878;
assign x_15880 = x_4636 & x_4637;
assign x_15881 = x_4639 & x_4640;
assign x_15882 = x_4638 & x_15881;
assign x_15883 = x_15880 & x_15882;
assign x_15884 = x_4642 & x_4643;
assign x_15885 = x_4641 & x_15884;
assign x_15886 = x_4645 & x_4646;
assign x_15887 = x_4644 & x_15886;
assign x_15888 = x_15885 & x_15887;
assign x_15889 = x_15883 & x_15888;
assign x_15890 = x_4647 & x_4648;
assign x_15891 = x_4650 & x_4651;
assign x_15892 = x_4649 & x_15891;
assign x_15893 = x_15890 & x_15892;
assign x_15894 = x_4653 & x_4654;
assign x_15895 = x_4652 & x_15894;
assign x_15896 = x_4656 & x_4657;
assign x_15897 = x_4655 & x_15896;
assign x_15898 = x_15895 & x_15897;
assign x_15899 = x_15893 & x_15898;
assign x_15900 = x_15889 & x_15899;
assign x_15901 = x_15879 & x_15900;
assign x_15902 = x_15858 & x_15901;
assign x_15903 = x_4658 & x_4659;
assign x_15904 = x_4661 & x_4662;
assign x_15905 = x_4660 & x_15904;
assign x_15906 = x_15903 & x_15905;
assign x_15907 = x_4664 & x_4665;
assign x_15908 = x_4663 & x_15907;
assign x_15909 = x_4667 & x_4668;
assign x_15910 = x_4666 & x_15909;
assign x_15911 = x_15908 & x_15910;
assign x_15912 = x_15906 & x_15911;
assign x_15913 = x_4669 & x_4670;
assign x_15914 = x_4672 & x_4673;
assign x_15915 = x_4671 & x_15914;
assign x_15916 = x_15913 & x_15915;
assign x_15917 = x_4675 & x_4676;
assign x_15918 = x_4674 & x_15917;
assign x_15919 = x_4678 & x_4679;
assign x_15920 = x_4677 & x_15919;
assign x_15921 = x_15918 & x_15920;
assign x_15922 = x_15916 & x_15921;
assign x_15923 = x_15912 & x_15922;
assign x_15924 = x_4680 & x_4681;
assign x_15925 = x_4683 & x_4684;
assign x_15926 = x_4682 & x_15925;
assign x_15927 = x_15924 & x_15926;
assign x_15928 = x_4686 & x_4687;
assign x_15929 = x_4685 & x_15928;
assign x_15930 = x_4689 & x_4690;
assign x_15931 = x_4688 & x_15930;
assign x_15932 = x_15929 & x_15931;
assign x_15933 = x_15927 & x_15932;
assign x_15934 = x_4691 & x_4692;
assign x_15935 = x_4694 & x_4695;
assign x_15936 = x_4693 & x_15935;
assign x_15937 = x_15934 & x_15936;
assign x_15938 = x_4697 & x_4698;
assign x_15939 = x_4696 & x_15938;
assign x_15940 = x_4700 & x_4701;
assign x_15941 = x_4699 & x_15940;
assign x_15942 = x_15939 & x_15941;
assign x_15943 = x_15937 & x_15942;
assign x_15944 = x_15933 & x_15943;
assign x_15945 = x_15923 & x_15944;
assign x_15946 = x_4702 & x_4703;
assign x_15947 = x_4705 & x_4706;
assign x_15948 = x_4704 & x_15947;
assign x_15949 = x_15946 & x_15948;
assign x_15950 = x_4708 & x_4709;
assign x_15951 = x_4707 & x_15950;
assign x_15952 = x_4711 & x_4712;
assign x_15953 = x_4710 & x_15952;
assign x_15954 = x_15951 & x_15953;
assign x_15955 = x_15949 & x_15954;
assign x_15956 = x_4713 & x_4714;
assign x_15957 = x_4716 & x_4717;
assign x_15958 = x_4715 & x_15957;
assign x_15959 = x_15956 & x_15958;
assign x_15960 = x_4719 & x_4720;
assign x_15961 = x_4718 & x_15960;
assign x_15962 = x_4722 & x_4723;
assign x_15963 = x_4721 & x_15962;
assign x_15964 = x_15961 & x_15963;
assign x_15965 = x_15959 & x_15964;
assign x_15966 = x_15955 & x_15965;
assign x_15967 = x_4724 & x_4725;
assign x_15968 = x_4727 & x_4728;
assign x_15969 = x_4726 & x_15968;
assign x_15970 = x_15967 & x_15969;
assign x_15971 = x_4730 & x_4731;
assign x_15972 = x_4729 & x_15971;
assign x_15973 = x_4733 & x_4734;
assign x_15974 = x_4732 & x_15973;
assign x_15975 = x_15972 & x_15974;
assign x_15976 = x_15970 & x_15975;
assign x_15977 = x_4735 & x_4736;
assign x_15978 = x_4738 & x_4739;
assign x_15979 = x_4737 & x_15978;
assign x_15980 = x_15977 & x_15979;
assign x_15981 = x_4741 & x_4742;
assign x_15982 = x_4740 & x_15981;
assign x_15983 = x_4744 & x_4745;
assign x_15984 = x_4743 & x_15983;
assign x_15985 = x_15982 & x_15984;
assign x_15986 = x_15980 & x_15985;
assign x_15987 = x_15976 & x_15986;
assign x_15988 = x_15966 & x_15987;
assign x_15989 = x_15945 & x_15988;
assign x_15990 = x_15902 & x_15989;
assign x_15991 = x_4746 & x_4747;
assign x_15992 = x_4749 & x_4750;
assign x_15993 = x_4748 & x_15992;
assign x_15994 = x_15991 & x_15993;
assign x_15995 = x_4752 & x_4753;
assign x_15996 = x_4751 & x_15995;
assign x_15997 = x_4755 & x_4756;
assign x_15998 = x_4754 & x_15997;
assign x_15999 = x_15996 & x_15998;
assign x_16000 = x_15994 & x_15999;
assign x_16001 = x_4757 & x_4758;
assign x_16002 = x_4760 & x_4761;
assign x_16003 = x_4759 & x_16002;
assign x_16004 = x_16001 & x_16003;
assign x_16005 = x_4763 & x_4764;
assign x_16006 = x_4762 & x_16005;
assign x_16007 = x_4766 & x_4767;
assign x_16008 = x_4765 & x_16007;
assign x_16009 = x_16006 & x_16008;
assign x_16010 = x_16004 & x_16009;
assign x_16011 = x_16000 & x_16010;
assign x_16012 = x_4768 & x_4769;
assign x_16013 = x_4771 & x_4772;
assign x_16014 = x_4770 & x_16013;
assign x_16015 = x_16012 & x_16014;
assign x_16016 = x_4774 & x_4775;
assign x_16017 = x_4773 & x_16016;
assign x_16018 = x_4777 & x_4778;
assign x_16019 = x_4776 & x_16018;
assign x_16020 = x_16017 & x_16019;
assign x_16021 = x_16015 & x_16020;
assign x_16022 = x_4779 & x_4780;
assign x_16023 = x_4782 & x_4783;
assign x_16024 = x_4781 & x_16023;
assign x_16025 = x_16022 & x_16024;
assign x_16026 = x_4785 & x_4786;
assign x_16027 = x_4784 & x_16026;
assign x_16028 = x_4788 & x_4789;
assign x_16029 = x_4787 & x_16028;
assign x_16030 = x_16027 & x_16029;
assign x_16031 = x_16025 & x_16030;
assign x_16032 = x_16021 & x_16031;
assign x_16033 = x_16011 & x_16032;
assign x_16034 = x_4790 & x_4791;
assign x_16035 = x_4793 & x_4794;
assign x_16036 = x_4792 & x_16035;
assign x_16037 = x_16034 & x_16036;
assign x_16038 = x_4796 & x_4797;
assign x_16039 = x_4795 & x_16038;
assign x_16040 = x_4799 & x_4800;
assign x_16041 = x_4798 & x_16040;
assign x_16042 = x_16039 & x_16041;
assign x_16043 = x_16037 & x_16042;
assign x_16044 = x_4801 & x_4802;
assign x_16045 = x_4804 & x_4805;
assign x_16046 = x_4803 & x_16045;
assign x_16047 = x_16044 & x_16046;
assign x_16048 = x_4807 & x_4808;
assign x_16049 = x_4806 & x_16048;
assign x_16050 = x_4810 & x_4811;
assign x_16051 = x_4809 & x_16050;
assign x_16052 = x_16049 & x_16051;
assign x_16053 = x_16047 & x_16052;
assign x_16054 = x_16043 & x_16053;
assign x_16055 = x_4812 & x_4813;
assign x_16056 = x_4815 & x_4816;
assign x_16057 = x_4814 & x_16056;
assign x_16058 = x_16055 & x_16057;
assign x_16059 = x_4818 & x_4819;
assign x_16060 = x_4817 & x_16059;
assign x_16061 = x_4821 & x_4822;
assign x_16062 = x_4820 & x_16061;
assign x_16063 = x_16060 & x_16062;
assign x_16064 = x_16058 & x_16063;
assign x_16065 = x_4823 & x_4824;
assign x_16066 = x_4826 & x_4827;
assign x_16067 = x_4825 & x_16066;
assign x_16068 = x_16065 & x_16067;
assign x_16069 = x_4829 & x_4830;
assign x_16070 = x_4828 & x_16069;
assign x_16071 = x_4832 & x_4833;
assign x_16072 = x_4831 & x_16071;
assign x_16073 = x_16070 & x_16072;
assign x_16074 = x_16068 & x_16073;
assign x_16075 = x_16064 & x_16074;
assign x_16076 = x_16054 & x_16075;
assign x_16077 = x_16033 & x_16076;
assign x_16078 = x_4834 & x_4835;
assign x_16079 = x_4837 & x_4838;
assign x_16080 = x_4836 & x_16079;
assign x_16081 = x_16078 & x_16080;
assign x_16082 = x_4840 & x_4841;
assign x_16083 = x_4839 & x_16082;
assign x_16084 = x_4843 & x_4844;
assign x_16085 = x_4842 & x_16084;
assign x_16086 = x_16083 & x_16085;
assign x_16087 = x_16081 & x_16086;
assign x_16088 = x_4845 & x_4846;
assign x_16089 = x_4848 & x_4849;
assign x_16090 = x_4847 & x_16089;
assign x_16091 = x_16088 & x_16090;
assign x_16092 = x_4851 & x_4852;
assign x_16093 = x_4850 & x_16092;
assign x_16094 = x_4854 & x_4855;
assign x_16095 = x_4853 & x_16094;
assign x_16096 = x_16093 & x_16095;
assign x_16097 = x_16091 & x_16096;
assign x_16098 = x_16087 & x_16097;
assign x_16099 = x_4856 & x_4857;
assign x_16100 = x_4859 & x_4860;
assign x_16101 = x_4858 & x_16100;
assign x_16102 = x_16099 & x_16101;
assign x_16103 = x_4862 & x_4863;
assign x_16104 = x_4861 & x_16103;
assign x_16105 = x_4865 & x_4866;
assign x_16106 = x_4864 & x_16105;
assign x_16107 = x_16104 & x_16106;
assign x_16108 = x_16102 & x_16107;
assign x_16109 = x_4867 & x_4868;
assign x_16110 = x_4870 & x_4871;
assign x_16111 = x_4869 & x_16110;
assign x_16112 = x_16109 & x_16111;
assign x_16113 = x_4873 & x_4874;
assign x_16114 = x_4872 & x_16113;
assign x_16115 = x_4876 & x_4877;
assign x_16116 = x_4875 & x_16115;
assign x_16117 = x_16114 & x_16116;
assign x_16118 = x_16112 & x_16117;
assign x_16119 = x_16108 & x_16118;
assign x_16120 = x_16098 & x_16119;
assign x_16121 = x_4878 & x_4879;
assign x_16122 = x_4881 & x_4882;
assign x_16123 = x_4880 & x_16122;
assign x_16124 = x_16121 & x_16123;
assign x_16125 = x_4884 & x_4885;
assign x_16126 = x_4883 & x_16125;
assign x_16127 = x_4887 & x_4888;
assign x_16128 = x_4886 & x_16127;
assign x_16129 = x_16126 & x_16128;
assign x_16130 = x_16124 & x_16129;
assign x_16131 = x_4889 & x_4890;
assign x_16132 = x_4892 & x_4893;
assign x_16133 = x_4891 & x_16132;
assign x_16134 = x_16131 & x_16133;
assign x_16135 = x_4895 & x_4896;
assign x_16136 = x_4894 & x_16135;
assign x_16137 = x_4898 & x_4899;
assign x_16138 = x_4897 & x_16137;
assign x_16139 = x_16136 & x_16138;
assign x_16140 = x_16134 & x_16139;
assign x_16141 = x_16130 & x_16140;
assign x_16142 = x_4900 & x_4901;
assign x_16143 = x_4903 & x_4904;
assign x_16144 = x_4902 & x_16143;
assign x_16145 = x_16142 & x_16144;
assign x_16146 = x_4906 & x_4907;
assign x_16147 = x_4905 & x_16146;
assign x_16148 = x_4909 & x_4910;
assign x_16149 = x_4908 & x_16148;
assign x_16150 = x_16147 & x_16149;
assign x_16151 = x_16145 & x_16150;
assign x_16152 = x_4911 & x_4912;
assign x_16153 = x_4914 & x_4915;
assign x_16154 = x_4913 & x_16153;
assign x_16155 = x_16152 & x_16154;
assign x_16156 = x_4917 & x_4918;
assign x_16157 = x_4916 & x_16156;
assign x_16158 = x_4920 & x_4921;
assign x_16159 = x_4919 & x_16158;
assign x_16160 = x_16157 & x_16159;
assign x_16161 = x_16155 & x_16160;
assign x_16162 = x_16151 & x_16161;
assign x_16163 = x_16141 & x_16162;
assign x_16164 = x_16120 & x_16163;
assign x_16165 = x_16077 & x_16164;
assign x_16166 = x_15990 & x_16165;
assign x_16167 = x_15815 & x_16166;
assign x_16168 = x_4922 & x_4923;
assign x_16169 = x_4925 & x_4926;
assign x_16170 = x_4924 & x_16169;
assign x_16171 = x_16168 & x_16170;
assign x_16172 = x_4927 & x_4928;
assign x_16173 = x_4930 & x_4931;
assign x_16174 = x_4929 & x_16173;
assign x_16175 = x_16172 & x_16174;
assign x_16176 = x_16171 & x_16175;
assign x_16177 = x_4932 & x_4933;
assign x_16178 = x_4935 & x_4936;
assign x_16179 = x_4934 & x_16178;
assign x_16180 = x_16177 & x_16179;
assign x_16181 = x_4938 & x_4939;
assign x_16182 = x_4937 & x_16181;
assign x_16183 = x_4941 & x_4942;
assign x_16184 = x_4940 & x_16183;
assign x_16185 = x_16182 & x_16184;
assign x_16186 = x_16180 & x_16185;
assign x_16187 = x_16176 & x_16186;
assign x_16188 = x_4943 & x_4944;
assign x_16189 = x_4946 & x_4947;
assign x_16190 = x_4945 & x_16189;
assign x_16191 = x_16188 & x_16190;
assign x_16192 = x_4949 & x_4950;
assign x_16193 = x_4948 & x_16192;
assign x_16194 = x_4952 & x_4953;
assign x_16195 = x_4951 & x_16194;
assign x_16196 = x_16193 & x_16195;
assign x_16197 = x_16191 & x_16196;
assign x_16198 = x_4954 & x_4955;
assign x_16199 = x_4957 & x_4958;
assign x_16200 = x_4956 & x_16199;
assign x_16201 = x_16198 & x_16200;
assign x_16202 = x_4960 & x_4961;
assign x_16203 = x_4959 & x_16202;
assign x_16204 = x_4963 & x_4964;
assign x_16205 = x_4962 & x_16204;
assign x_16206 = x_16203 & x_16205;
assign x_16207 = x_16201 & x_16206;
assign x_16208 = x_16197 & x_16207;
assign x_16209 = x_16187 & x_16208;
assign x_16210 = x_4965 & x_4966;
assign x_16211 = x_4968 & x_4969;
assign x_16212 = x_4967 & x_16211;
assign x_16213 = x_16210 & x_16212;
assign x_16214 = x_4971 & x_4972;
assign x_16215 = x_4970 & x_16214;
assign x_16216 = x_4974 & x_4975;
assign x_16217 = x_4973 & x_16216;
assign x_16218 = x_16215 & x_16217;
assign x_16219 = x_16213 & x_16218;
assign x_16220 = x_4976 & x_4977;
assign x_16221 = x_4979 & x_4980;
assign x_16222 = x_4978 & x_16221;
assign x_16223 = x_16220 & x_16222;
assign x_16224 = x_4982 & x_4983;
assign x_16225 = x_4981 & x_16224;
assign x_16226 = x_4985 & x_4986;
assign x_16227 = x_4984 & x_16226;
assign x_16228 = x_16225 & x_16227;
assign x_16229 = x_16223 & x_16228;
assign x_16230 = x_16219 & x_16229;
assign x_16231 = x_4987 & x_4988;
assign x_16232 = x_4990 & x_4991;
assign x_16233 = x_4989 & x_16232;
assign x_16234 = x_16231 & x_16233;
assign x_16235 = x_4993 & x_4994;
assign x_16236 = x_4992 & x_16235;
assign x_16237 = x_4996 & x_4997;
assign x_16238 = x_4995 & x_16237;
assign x_16239 = x_16236 & x_16238;
assign x_16240 = x_16234 & x_16239;
assign x_16241 = x_4998 & x_4999;
assign x_16242 = x_5001 & x_5002;
assign x_16243 = x_5000 & x_16242;
assign x_16244 = x_16241 & x_16243;
assign x_16245 = x_5004 & x_5005;
assign x_16246 = x_5003 & x_16245;
assign x_16247 = x_5007 & x_5008;
assign x_16248 = x_5006 & x_16247;
assign x_16249 = x_16246 & x_16248;
assign x_16250 = x_16244 & x_16249;
assign x_16251 = x_16240 & x_16250;
assign x_16252 = x_16230 & x_16251;
assign x_16253 = x_16209 & x_16252;
assign x_16254 = x_5009 & x_5010;
assign x_16255 = x_5012 & x_5013;
assign x_16256 = x_5011 & x_16255;
assign x_16257 = x_16254 & x_16256;
assign x_16258 = x_5015 & x_5016;
assign x_16259 = x_5014 & x_16258;
assign x_16260 = x_5018 & x_5019;
assign x_16261 = x_5017 & x_16260;
assign x_16262 = x_16259 & x_16261;
assign x_16263 = x_16257 & x_16262;
assign x_16264 = x_5020 & x_5021;
assign x_16265 = x_5023 & x_5024;
assign x_16266 = x_5022 & x_16265;
assign x_16267 = x_16264 & x_16266;
assign x_16268 = x_5026 & x_5027;
assign x_16269 = x_5025 & x_16268;
assign x_16270 = x_5029 & x_5030;
assign x_16271 = x_5028 & x_16270;
assign x_16272 = x_16269 & x_16271;
assign x_16273 = x_16267 & x_16272;
assign x_16274 = x_16263 & x_16273;
assign x_16275 = x_5031 & x_5032;
assign x_16276 = x_5034 & x_5035;
assign x_16277 = x_5033 & x_16276;
assign x_16278 = x_16275 & x_16277;
assign x_16279 = x_5037 & x_5038;
assign x_16280 = x_5036 & x_16279;
assign x_16281 = x_5040 & x_5041;
assign x_16282 = x_5039 & x_16281;
assign x_16283 = x_16280 & x_16282;
assign x_16284 = x_16278 & x_16283;
assign x_16285 = x_5042 & x_5043;
assign x_16286 = x_5045 & x_5046;
assign x_16287 = x_5044 & x_16286;
assign x_16288 = x_16285 & x_16287;
assign x_16289 = x_5048 & x_5049;
assign x_16290 = x_5047 & x_16289;
assign x_16291 = x_5051 & x_5052;
assign x_16292 = x_5050 & x_16291;
assign x_16293 = x_16290 & x_16292;
assign x_16294 = x_16288 & x_16293;
assign x_16295 = x_16284 & x_16294;
assign x_16296 = x_16274 & x_16295;
assign x_16297 = x_5053 & x_5054;
assign x_16298 = x_5056 & x_5057;
assign x_16299 = x_5055 & x_16298;
assign x_16300 = x_16297 & x_16299;
assign x_16301 = x_5059 & x_5060;
assign x_16302 = x_5058 & x_16301;
assign x_16303 = x_5062 & x_5063;
assign x_16304 = x_5061 & x_16303;
assign x_16305 = x_16302 & x_16304;
assign x_16306 = x_16300 & x_16305;
assign x_16307 = x_5064 & x_5065;
assign x_16308 = x_5067 & x_5068;
assign x_16309 = x_5066 & x_16308;
assign x_16310 = x_16307 & x_16309;
assign x_16311 = x_5070 & x_5071;
assign x_16312 = x_5069 & x_16311;
assign x_16313 = x_5073 & x_5074;
assign x_16314 = x_5072 & x_16313;
assign x_16315 = x_16312 & x_16314;
assign x_16316 = x_16310 & x_16315;
assign x_16317 = x_16306 & x_16316;
assign x_16318 = x_5075 & x_5076;
assign x_16319 = x_5078 & x_5079;
assign x_16320 = x_5077 & x_16319;
assign x_16321 = x_16318 & x_16320;
assign x_16322 = x_5081 & x_5082;
assign x_16323 = x_5080 & x_16322;
assign x_16324 = x_5084 & x_5085;
assign x_16325 = x_5083 & x_16324;
assign x_16326 = x_16323 & x_16325;
assign x_16327 = x_16321 & x_16326;
assign x_16328 = x_5086 & x_5087;
assign x_16329 = x_5089 & x_5090;
assign x_16330 = x_5088 & x_16329;
assign x_16331 = x_16328 & x_16330;
assign x_16332 = x_5092 & x_5093;
assign x_16333 = x_5091 & x_16332;
assign x_16334 = x_5095 & x_5096;
assign x_16335 = x_5094 & x_16334;
assign x_16336 = x_16333 & x_16335;
assign x_16337 = x_16331 & x_16336;
assign x_16338 = x_16327 & x_16337;
assign x_16339 = x_16317 & x_16338;
assign x_16340 = x_16296 & x_16339;
assign x_16341 = x_16253 & x_16340;
assign x_16342 = x_5097 & x_5098;
assign x_16343 = x_5100 & x_5101;
assign x_16344 = x_5099 & x_16343;
assign x_16345 = x_16342 & x_16344;
assign x_16346 = x_5103 & x_5104;
assign x_16347 = x_5102 & x_16346;
assign x_16348 = x_5106 & x_5107;
assign x_16349 = x_5105 & x_16348;
assign x_16350 = x_16347 & x_16349;
assign x_16351 = x_16345 & x_16350;
assign x_16352 = x_5108 & x_5109;
assign x_16353 = x_5111 & x_5112;
assign x_16354 = x_5110 & x_16353;
assign x_16355 = x_16352 & x_16354;
assign x_16356 = x_5114 & x_5115;
assign x_16357 = x_5113 & x_16356;
assign x_16358 = x_5117 & x_5118;
assign x_16359 = x_5116 & x_16358;
assign x_16360 = x_16357 & x_16359;
assign x_16361 = x_16355 & x_16360;
assign x_16362 = x_16351 & x_16361;
assign x_16363 = x_5119 & x_5120;
assign x_16364 = x_5122 & x_5123;
assign x_16365 = x_5121 & x_16364;
assign x_16366 = x_16363 & x_16365;
assign x_16367 = x_5125 & x_5126;
assign x_16368 = x_5124 & x_16367;
assign x_16369 = x_5128 & x_5129;
assign x_16370 = x_5127 & x_16369;
assign x_16371 = x_16368 & x_16370;
assign x_16372 = x_16366 & x_16371;
assign x_16373 = x_5130 & x_5131;
assign x_16374 = x_5133 & x_5134;
assign x_16375 = x_5132 & x_16374;
assign x_16376 = x_16373 & x_16375;
assign x_16377 = x_5136 & x_5137;
assign x_16378 = x_5135 & x_16377;
assign x_16379 = x_5139 & x_5140;
assign x_16380 = x_5138 & x_16379;
assign x_16381 = x_16378 & x_16380;
assign x_16382 = x_16376 & x_16381;
assign x_16383 = x_16372 & x_16382;
assign x_16384 = x_16362 & x_16383;
assign x_16385 = x_5141 & x_5142;
assign x_16386 = x_5144 & x_5145;
assign x_16387 = x_5143 & x_16386;
assign x_16388 = x_16385 & x_16387;
assign x_16389 = x_5147 & x_5148;
assign x_16390 = x_5146 & x_16389;
assign x_16391 = x_5150 & x_5151;
assign x_16392 = x_5149 & x_16391;
assign x_16393 = x_16390 & x_16392;
assign x_16394 = x_16388 & x_16393;
assign x_16395 = x_5152 & x_5153;
assign x_16396 = x_5155 & x_5156;
assign x_16397 = x_5154 & x_16396;
assign x_16398 = x_16395 & x_16397;
assign x_16399 = x_5158 & x_5159;
assign x_16400 = x_5157 & x_16399;
assign x_16401 = x_5161 & x_5162;
assign x_16402 = x_5160 & x_16401;
assign x_16403 = x_16400 & x_16402;
assign x_16404 = x_16398 & x_16403;
assign x_16405 = x_16394 & x_16404;
assign x_16406 = x_5163 & x_5164;
assign x_16407 = x_5166 & x_5167;
assign x_16408 = x_5165 & x_16407;
assign x_16409 = x_16406 & x_16408;
assign x_16410 = x_5169 & x_5170;
assign x_16411 = x_5168 & x_16410;
assign x_16412 = x_5172 & x_5173;
assign x_16413 = x_5171 & x_16412;
assign x_16414 = x_16411 & x_16413;
assign x_16415 = x_16409 & x_16414;
assign x_16416 = x_5174 & x_5175;
assign x_16417 = x_5177 & x_5178;
assign x_16418 = x_5176 & x_16417;
assign x_16419 = x_16416 & x_16418;
assign x_16420 = x_5180 & x_5181;
assign x_16421 = x_5179 & x_16420;
assign x_16422 = x_5183 & x_5184;
assign x_16423 = x_5182 & x_16422;
assign x_16424 = x_16421 & x_16423;
assign x_16425 = x_16419 & x_16424;
assign x_16426 = x_16415 & x_16425;
assign x_16427 = x_16405 & x_16426;
assign x_16428 = x_16384 & x_16427;
assign x_16429 = x_5185 & x_5186;
assign x_16430 = x_5188 & x_5189;
assign x_16431 = x_5187 & x_16430;
assign x_16432 = x_16429 & x_16431;
assign x_16433 = x_5191 & x_5192;
assign x_16434 = x_5190 & x_16433;
assign x_16435 = x_5194 & x_5195;
assign x_16436 = x_5193 & x_16435;
assign x_16437 = x_16434 & x_16436;
assign x_16438 = x_16432 & x_16437;
assign x_16439 = x_5196 & x_5197;
assign x_16440 = x_5199 & x_5200;
assign x_16441 = x_5198 & x_16440;
assign x_16442 = x_16439 & x_16441;
assign x_16443 = x_5202 & x_5203;
assign x_16444 = x_5201 & x_16443;
assign x_16445 = x_5205 & x_5206;
assign x_16446 = x_5204 & x_16445;
assign x_16447 = x_16444 & x_16446;
assign x_16448 = x_16442 & x_16447;
assign x_16449 = x_16438 & x_16448;
assign x_16450 = x_5207 & x_5208;
assign x_16451 = x_5210 & x_5211;
assign x_16452 = x_5209 & x_16451;
assign x_16453 = x_16450 & x_16452;
assign x_16454 = x_5213 & x_5214;
assign x_16455 = x_5212 & x_16454;
assign x_16456 = x_5216 & x_5217;
assign x_16457 = x_5215 & x_16456;
assign x_16458 = x_16455 & x_16457;
assign x_16459 = x_16453 & x_16458;
assign x_16460 = x_5218 & x_5219;
assign x_16461 = x_5221 & x_5222;
assign x_16462 = x_5220 & x_16461;
assign x_16463 = x_16460 & x_16462;
assign x_16464 = x_5224 & x_5225;
assign x_16465 = x_5223 & x_16464;
assign x_16466 = x_5227 & x_5228;
assign x_16467 = x_5226 & x_16466;
assign x_16468 = x_16465 & x_16467;
assign x_16469 = x_16463 & x_16468;
assign x_16470 = x_16459 & x_16469;
assign x_16471 = x_16449 & x_16470;
assign x_16472 = x_5229 & x_5230;
assign x_16473 = x_5232 & x_5233;
assign x_16474 = x_5231 & x_16473;
assign x_16475 = x_16472 & x_16474;
assign x_16476 = x_5235 & x_5236;
assign x_16477 = x_5234 & x_16476;
assign x_16478 = x_5238 & x_5239;
assign x_16479 = x_5237 & x_16478;
assign x_16480 = x_16477 & x_16479;
assign x_16481 = x_16475 & x_16480;
assign x_16482 = x_5240 & x_5241;
assign x_16483 = x_5243 & x_5244;
assign x_16484 = x_5242 & x_16483;
assign x_16485 = x_16482 & x_16484;
assign x_16486 = x_5246 & x_5247;
assign x_16487 = x_5245 & x_16486;
assign x_16488 = x_5249 & x_5250;
assign x_16489 = x_5248 & x_16488;
assign x_16490 = x_16487 & x_16489;
assign x_16491 = x_16485 & x_16490;
assign x_16492 = x_16481 & x_16491;
assign x_16493 = x_5251 & x_5252;
assign x_16494 = x_5254 & x_5255;
assign x_16495 = x_5253 & x_16494;
assign x_16496 = x_16493 & x_16495;
assign x_16497 = x_5257 & x_5258;
assign x_16498 = x_5256 & x_16497;
assign x_16499 = x_5260 & x_5261;
assign x_16500 = x_5259 & x_16499;
assign x_16501 = x_16498 & x_16500;
assign x_16502 = x_16496 & x_16501;
assign x_16503 = x_5262 & x_5263;
assign x_16504 = x_5265 & x_5266;
assign x_16505 = x_5264 & x_16504;
assign x_16506 = x_16503 & x_16505;
assign x_16507 = x_5268 & x_5269;
assign x_16508 = x_5267 & x_16507;
assign x_16509 = x_5271 & x_5272;
assign x_16510 = x_5270 & x_16509;
assign x_16511 = x_16508 & x_16510;
assign x_16512 = x_16506 & x_16511;
assign x_16513 = x_16502 & x_16512;
assign x_16514 = x_16492 & x_16513;
assign x_16515 = x_16471 & x_16514;
assign x_16516 = x_16428 & x_16515;
assign x_16517 = x_16341 & x_16516;
assign x_16518 = x_5273 & x_5274;
assign x_16519 = x_5276 & x_5277;
assign x_16520 = x_5275 & x_16519;
assign x_16521 = x_16518 & x_16520;
assign x_16522 = x_5279 & x_5280;
assign x_16523 = x_5278 & x_16522;
assign x_16524 = x_5282 & x_5283;
assign x_16525 = x_5281 & x_16524;
assign x_16526 = x_16523 & x_16525;
assign x_16527 = x_16521 & x_16526;
assign x_16528 = x_5284 & x_5285;
assign x_16529 = x_5287 & x_5288;
assign x_16530 = x_5286 & x_16529;
assign x_16531 = x_16528 & x_16530;
assign x_16532 = x_5290 & x_5291;
assign x_16533 = x_5289 & x_16532;
assign x_16534 = x_5293 & x_5294;
assign x_16535 = x_5292 & x_16534;
assign x_16536 = x_16533 & x_16535;
assign x_16537 = x_16531 & x_16536;
assign x_16538 = x_16527 & x_16537;
assign x_16539 = x_5295 & x_5296;
assign x_16540 = x_5298 & x_5299;
assign x_16541 = x_5297 & x_16540;
assign x_16542 = x_16539 & x_16541;
assign x_16543 = x_5301 & x_5302;
assign x_16544 = x_5300 & x_16543;
assign x_16545 = x_5304 & x_5305;
assign x_16546 = x_5303 & x_16545;
assign x_16547 = x_16544 & x_16546;
assign x_16548 = x_16542 & x_16547;
assign x_16549 = x_5306 & x_5307;
assign x_16550 = x_5309 & x_5310;
assign x_16551 = x_5308 & x_16550;
assign x_16552 = x_16549 & x_16551;
assign x_16553 = x_5312 & x_5313;
assign x_16554 = x_5311 & x_16553;
assign x_16555 = x_5315 & x_5316;
assign x_16556 = x_5314 & x_16555;
assign x_16557 = x_16554 & x_16556;
assign x_16558 = x_16552 & x_16557;
assign x_16559 = x_16548 & x_16558;
assign x_16560 = x_16538 & x_16559;
assign x_16561 = x_5317 & x_5318;
assign x_16562 = x_5320 & x_5321;
assign x_16563 = x_5319 & x_16562;
assign x_16564 = x_16561 & x_16563;
assign x_16565 = x_5323 & x_5324;
assign x_16566 = x_5322 & x_16565;
assign x_16567 = x_5326 & x_5327;
assign x_16568 = x_5325 & x_16567;
assign x_16569 = x_16566 & x_16568;
assign x_16570 = x_16564 & x_16569;
assign x_16571 = x_5328 & x_5329;
assign x_16572 = x_5331 & x_5332;
assign x_16573 = x_5330 & x_16572;
assign x_16574 = x_16571 & x_16573;
assign x_16575 = x_5334 & x_5335;
assign x_16576 = x_5333 & x_16575;
assign x_16577 = x_5337 & x_5338;
assign x_16578 = x_5336 & x_16577;
assign x_16579 = x_16576 & x_16578;
assign x_16580 = x_16574 & x_16579;
assign x_16581 = x_16570 & x_16580;
assign x_16582 = x_5339 & x_5340;
assign x_16583 = x_5342 & x_5343;
assign x_16584 = x_5341 & x_16583;
assign x_16585 = x_16582 & x_16584;
assign x_16586 = x_5345 & x_5346;
assign x_16587 = x_5344 & x_16586;
assign x_16588 = x_5348 & x_5349;
assign x_16589 = x_5347 & x_16588;
assign x_16590 = x_16587 & x_16589;
assign x_16591 = x_16585 & x_16590;
assign x_16592 = x_5350 & x_5351;
assign x_16593 = x_5353 & x_5354;
assign x_16594 = x_5352 & x_16593;
assign x_16595 = x_16592 & x_16594;
assign x_16596 = x_5356 & x_5357;
assign x_16597 = x_5355 & x_16596;
assign x_16598 = x_5359 & x_5360;
assign x_16599 = x_5358 & x_16598;
assign x_16600 = x_16597 & x_16599;
assign x_16601 = x_16595 & x_16600;
assign x_16602 = x_16591 & x_16601;
assign x_16603 = x_16581 & x_16602;
assign x_16604 = x_16560 & x_16603;
assign x_16605 = x_5361 & x_5362;
assign x_16606 = x_5364 & x_5365;
assign x_16607 = x_5363 & x_16606;
assign x_16608 = x_16605 & x_16607;
assign x_16609 = x_5367 & x_5368;
assign x_16610 = x_5366 & x_16609;
assign x_16611 = x_5370 & x_5371;
assign x_16612 = x_5369 & x_16611;
assign x_16613 = x_16610 & x_16612;
assign x_16614 = x_16608 & x_16613;
assign x_16615 = x_5372 & x_5373;
assign x_16616 = x_5375 & x_5376;
assign x_16617 = x_5374 & x_16616;
assign x_16618 = x_16615 & x_16617;
assign x_16619 = x_5378 & x_5379;
assign x_16620 = x_5377 & x_16619;
assign x_16621 = x_5381 & x_5382;
assign x_16622 = x_5380 & x_16621;
assign x_16623 = x_16620 & x_16622;
assign x_16624 = x_16618 & x_16623;
assign x_16625 = x_16614 & x_16624;
assign x_16626 = x_5383 & x_5384;
assign x_16627 = x_5386 & x_5387;
assign x_16628 = x_5385 & x_16627;
assign x_16629 = x_16626 & x_16628;
assign x_16630 = x_5389 & x_5390;
assign x_16631 = x_5388 & x_16630;
assign x_16632 = x_5392 & x_5393;
assign x_16633 = x_5391 & x_16632;
assign x_16634 = x_16631 & x_16633;
assign x_16635 = x_16629 & x_16634;
assign x_16636 = x_5394 & x_5395;
assign x_16637 = x_5397 & x_5398;
assign x_16638 = x_5396 & x_16637;
assign x_16639 = x_16636 & x_16638;
assign x_16640 = x_5400 & x_5401;
assign x_16641 = x_5399 & x_16640;
assign x_16642 = x_5403 & x_5404;
assign x_16643 = x_5402 & x_16642;
assign x_16644 = x_16641 & x_16643;
assign x_16645 = x_16639 & x_16644;
assign x_16646 = x_16635 & x_16645;
assign x_16647 = x_16625 & x_16646;
assign x_16648 = x_5405 & x_5406;
assign x_16649 = x_5408 & x_5409;
assign x_16650 = x_5407 & x_16649;
assign x_16651 = x_16648 & x_16650;
assign x_16652 = x_5411 & x_5412;
assign x_16653 = x_5410 & x_16652;
assign x_16654 = x_5414 & x_5415;
assign x_16655 = x_5413 & x_16654;
assign x_16656 = x_16653 & x_16655;
assign x_16657 = x_16651 & x_16656;
assign x_16658 = x_5416 & x_5417;
assign x_16659 = x_5419 & x_5420;
assign x_16660 = x_5418 & x_16659;
assign x_16661 = x_16658 & x_16660;
assign x_16662 = x_5422 & x_5423;
assign x_16663 = x_5421 & x_16662;
assign x_16664 = x_5425 & x_5426;
assign x_16665 = x_5424 & x_16664;
assign x_16666 = x_16663 & x_16665;
assign x_16667 = x_16661 & x_16666;
assign x_16668 = x_16657 & x_16667;
assign x_16669 = x_5427 & x_5428;
assign x_16670 = x_5430 & x_5431;
assign x_16671 = x_5429 & x_16670;
assign x_16672 = x_16669 & x_16671;
assign x_16673 = x_5433 & x_5434;
assign x_16674 = x_5432 & x_16673;
assign x_16675 = x_5436 & x_5437;
assign x_16676 = x_5435 & x_16675;
assign x_16677 = x_16674 & x_16676;
assign x_16678 = x_16672 & x_16677;
assign x_16679 = x_5438 & x_5439;
assign x_16680 = x_5441 & x_5442;
assign x_16681 = x_5440 & x_16680;
assign x_16682 = x_16679 & x_16681;
assign x_16683 = x_5444 & x_5445;
assign x_16684 = x_5443 & x_16683;
assign x_16685 = x_5447 & x_5448;
assign x_16686 = x_5446 & x_16685;
assign x_16687 = x_16684 & x_16686;
assign x_16688 = x_16682 & x_16687;
assign x_16689 = x_16678 & x_16688;
assign x_16690 = x_16668 & x_16689;
assign x_16691 = x_16647 & x_16690;
assign x_16692 = x_16604 & x_16691;
assign x_16693 = x_5449 & x_5450;
assign x_16694 = x_5452 & x_5453;
assign x_16695 = x_5451 & x_16694;
assign x_16696 = x_16693 & x_16695;
assign x_16697 = x_5455 & x_5456;
assign x_16698 = x_5454 & x_16697;
assign x_16699 = x_5458 & x_5459;
assign x_16700 = x_5457 & x_16699;
assign x_16701 = x_16698 & x_16700;
assign x_16702 = x_16696 & x_16701;
assign x_16703 = x_5460 & x_5461;
assign x_16704 = x_5463 & x_5464;
assign x_16705 = x_5462 & x_16704;
assign x_16706 = x_16703 & x_16705;
assign x_16707 = x_5466 & x_5467;
assign x_16708 = x_5465 & x_16707;
assign x_16709 = x_5469 & x_5470;
assign x_16710 = x_5468 & x_16709;
assign x_16711 = x_16708 & x_16710;
assign x_16712 = x_16706 & x_16711;
assign x_16713 = x_16702 & x_16712;
assign x_16714 = x_5471 & x_5472;
assign x_16715 = x_5474 & x_5475;
assign x_16716 = x_5473 & x_16715;
assign x_16717 = x_16714 & x_16716;
assign x_16718 = x_5477 & x_5478;
assign x_16719 = x_5476 & x_16718;
assign x_16720 = x_5480 & x_5481;
assign x_16721 = x_5479 & x_16720;
assign x_16722 = x_16719 & x_16721;
assign x_16723 = x_16717 & x_16722;
assign x_16724 = x_5482 & x_5483;
assign x_16725 = x_5485 & x_5486;
assign x_16726 = x_5484 & x_16725;
assign x_16727 = x_16724 & x_16726;
assign x_16728 = x_5488 & x_5489;
assign x_16729 = x_5487 & x_16728;
assign x_16730 = x_5491 & x_5492;
assign x_16731 = x_5490 & x_16730;
assign x_16732 = x_16729 & x_16731;
assign x_16733 = x_16727 & x_16732;
assign x_16734 = x_16723 & x_16733;
assign x_16735 = x_16713 & x_16734;
assign x_16736 = x_5493 & x_5494;
assign x_16737 = x_5496 & x_5497;
assign x_16738 = x_5495 & x_16737;
assign x_16739 = x_16736 & x_16738;
assign x_16740 = x_5499 & x_5500;
assign x_16741 = x_5498 & x_16740;
assign x_16742 = x_5502 & x_5503;
assign x_16743 = x_5501 & x_16742;
assign x_16744 = x_16741 & x_16743;
assign x_16745 = x_16739 & x_16744;
assign x_16746 = x_5504 & x_5505;
assign x_16747 = x_5507 & x_5508;
assign x_16748 = x_5506 & x_16747;
assign x_16749 = x_16746 & x_16748;
assign x_16750 = x_5510 & x_5511;
assign x_16751 = x_5509 & x_16750;
assign x_16752 = x_5513 & x_5514;
assign x_16753 = x_5512 & x_16752;
assign x_16754 = x_16751 & x_16753;
assign x_16755 = x_16749 & x_16754;
assign x_16756 = x_16745 & x_16755;
assign x_16757 = x_5515 & x_5516;
assign x_16758 = x_5518 & x_5519;
assign x_16759 = x_5517 & x_16758;
assign x_16760 = x_16757 & x_16759;
assign x_16761 = x_5521 & x_5522;
assign x_16762 = x_5520 & x_16761;
assign x_16763 = x_5524 & x_5525;
assign x_16764 = x_5523 & x_16763;
assign x_16765 = x_16762 & x_16764;
assign x_16766 = x_16760 & x_16765;
assign x_16767 = x_5526 & x_5527;
assign x_16768 = x_5529 & x_5530;
assign x_16769 = x_5528 & x_16768;
assign x_16770 = x_16767 & x_16769;
assign x_16771 = x_5532 & x_5533;
assign x_16772 = x_5531 & x_16771;
assign x_16773 = x_5535 & x_5536;
assign x_16774 = x_5534 & x_16773;
assign x_16775 = x_16772 & x_16774;
assign x_16776 = x_16770 & x_16775;
assign x_16777 = x_16766 & x_16776;
assign x_16778 = x_16756 & x_16777;
assign x_16779 = x_16735 & x_16778;
assign x_16780 = x_5537 & x_5538;
assign x_16781 = x_5540 & x_5541;
assign x_16782 = x_5539 & x_16781;
assign x_16783 = x_16780 & x_16782;
assign x_16784 = x_5543 & x_5544;
assign x_16785 = x_5542 & x_16784;
assign x_16786 = x_5546 & x_5547;
assign x_16787 = x_5545 & x_16786;
assign x_16788 = x_16785 & x_16787;
assign x_16789 = x_16783 & x_16788;
assign x_16790 = x_5548 & x_5549;
assign x_16791 = x_5551 & x_5552;
assign x_16792 = x_5550 & x_16791;
assign x_16793 = x_16790 & x_16792;
assign x_16794 = x_5554 & x_5555;
assign x_16795 = x_5553 & x_16794;
assign x_16796 = x_5557 & x_5558;
assign x_16797 = x_5556 & x_16796;
assign x_16798 = x_16795 & x_16797;
assign x_16799 = x_16793 & x_16798;
assign x_16800 = x_16789 & x_16799;
assign x_16801 = x_5559 & x_5560;
assign x_16802 = x_5562 & x_5563;
assign x_16803 = x_5561 & x_16802;
assign x_16804 = x_16801 & x_16803;
assign x_16805 = x_5565 & x_5566;
assign x_16806 = x_5564 & x_16805;
assign x_16807 = x_5568 & x_5569;
assign x_16808 = x_5567 & x_16807;
assign x_16809 = x_16806 & x_16808;
assign x_16810 = x_16804 & x_16809;
assign x_16811 = x_5570 & x_5571;
assign x_16812 = x_5573 & x_5574;
assign x_16813 = x_5572 & x_16812;
assign x_16814 = x_16811 & x_16813;
assign x_16815 = x_5576 & x_5577;
assign x_16816 = x_5575 & x_16815;
assign x_16817 = x_5579 & x_5580;
assign x_16818 = x_5578 & x_16817;
assign x_16819 = x_16816 & x_16818;
assign x_16820 = x_16814 & x_16819;
assign x_16821 = x_16810 & x_16820;
assign x_16822 = x_16800 & x_16821;
assign x_16823 = x_5581 & x_5582;
assign x_16824 = x_5584 & x_5585;
assign x_16825 = x_5583 & x_16824;
assign x_16826 = x_16823 & x_16825;
assign x_16827 = x_5587 & x_5588;
assign x_16828 = x_5586 & x_16827;
assign x_16829 = x_5590 & x_5591;
assign x_16830 = x_5589 & x_16829;
assign x_16831 = x_16828 & x_16830;
assign x_16832 = x_16826 & x_16831;
assign x_16833 = x_5592 & x_5593;
assign x_16834 = x_5595 & x_5596;
assign x_16835 = x_5594 & x_16834;
assign x_16836 = x_16833 & x_16835;
assign x_16837 = x_5598 & x_5599;
assign x_16838 = x_5597 & x_16837;
assign x_16839 = x_5601 & x_5602;
assign x_16840 = x_5600 & x_16839;
assign x_16841 = x_16838 & x_16840;
assign x_16842 = x_16836 & x_16841;
assign x_16843 = x_16832 & x_16842;
assign x_16844 = x_5603 & x_5604;
assign x_16845 = x_5606 & x_5607;
assign x_16846 = x_5605 & x_16845;
assign x_16847 = x_16844 & x_16846;
assign x_16848 = x_5609 & x_5610;
assign x_16849 = x_5608 & x_16848;
assign x_16850 = x_5612 & x_5613;
assign x_16851 = x_5611 & x_16850;
assign x_16852 = x_16849 & x_16851;
assign x_16853 = x_16847 & x_16852;
assign x_16854 = x_5614 & x_5615;
assign x_16855 = x_5617 & x_5618;
assign x_16856 = x_5616 & x_16855;
assign x_16857 = x_16854 & x_16856;
assign x_16858 = x_5620 & x_5621;
assign x_16859 = x_5619 & x_16858;
assign x_16860 = x_5623 & x_5624;
assign x_16861 = x_5622 & x_16860;
assign x_16862 = x_16859 & x_16861;
assign x_16863 = x_16857 & x_16862;
assign x_16864 = x_16853 & x_16863;
assign x_16865 = x_16843 & x_16864;
assign x_16866 = x_16822 & x_16865;
assign x_16867 = x_16779 & x_16866;
assign x_16868 = x_16692 & x_16867;
assign x_16869 = x_16517 & x_16868;
assign x_16870 = x_16167 & x_16869;
assign x_16871 = x_15465 & x_16870;
assign x_16872 = x_14060 & x_16871;
assign x_16873 = x_5625 & x_5626;
assign x_16874 = x_5628 & x_5629;
assign x_16875 = x_5627 & x_16874;
assign x_16876 = x_16873 & x_16875;
assign x_16877 = x_5630 & x_5631;
assign x_16878 = x_5633 & x_5634;
assign x_16879 = x_5632 & x_16878;
assign x_16880 = x_16877 & x_16879;
assign x_16881 = x_16876 & x_16880;
assign x_16882 = x_5635 & x_5636;
assign x_16883 = x_5638 & x_5639;
assign x_16884 = x_5637 & x_16883;
assign x_16885 = x_16882 & x_16884;
assign x_16886 = x_5641 & x_5642;
assign x_16887 = x_5640 & x_16886;
assign x_16888 = x_5644 & x_5645;
assign x_16889 = x_5643 & x_16888;
assign x_16890 = x_16887 & x_16889;
assign x_16891 = x_16885 & x_16890;
assign x_16892 = x_16881 & x_16891;
assign x_16893 = x_5646 & x_5647;
assign x_16894 = x_5649 & x_5650;
assign x_16895 = x_5648 & x_16894;
assign x_16896 = x_16893 & x_16895;
assign x_16897 = x_5652 & x_5653;
assign x_16898 = x_5651 & x_16897;
assign x_16899 = x_5655 & x_5656;
assign x_16900 = x_5654 & x_16899;
assign x_16901 = x_16898 & x_16900;
assign x_16902 = x_16896 & x_16901;
assign x_16903 = x_5657 & x_5658;
assign x_16904 = x_5660 & x_5661;
assign x_16905 = x_5659 & x_16904;
assign x_16906 = x_16903 & x_16905;
assign x_16907 = x_5663 & x_5664;
assign x_16908 = x_5662 & x_16907;
assign x_16909 = x_5666 & x_5667;
assign x_16910 = x_5665 & x_16909;
assign x_16911 = x_16908 & x_16910;
assign x_16912 = x_16906 & x_16911;
assign x_16913 = x_16902 & x_16912;
assign x_16914 = x_16892 & x_16913;
assign x_16915 = x_5668 & x_5669;
assign x_16916 = x_5671 & x_5672;
assign x_16917 = x_5670 & x_16916;
assign x_16918 = x_16915 & x_16917;
assign x_16919 = x_5674 & x_5675;
assign x_16920 = x_5673 & x_16919;
assign x_16921 = x_5677 & x_5678;
assign x_16922 = x_5676 & x_16921;
assign x_16923 = x_16920 & x_16922;
assign x_16924 = x_16918 & x_16923;
assign x_16925 = x_5679 & x_5680;
assign x_16926 = x_5682 & x_5683;
assign x_16927 = x_5681 & x_16926;
assign x_16928 = x_16925 & x_16927;
assign x_16929 = x_5685 & x_5686;
assign x_16930 = x_5684 & x_16929;
assign x_16931 = x_5688 & x_5689;
assign x_16932 = x_5687 & x_16931;
assign x_16933 = x_16930 & x_16932;
assign x_16934 = x_16928 & x_16933;
assign x_16935 = x_16924 & x_16934;
assign x_16936 = x_5690 & x_5691;
assign x_16937 = x_5693 & x_5694;
assign x_16938 = x_5692 & x_16937;
assign x_16939 = x_16936 & x_16938;
assign x_16940 = x_5696 & x_5697;
assign x_16941 = x_5695 & x_16940;
assign x_16942 = x_5699 & x_5700;
assign x_16943 = x_5698 & x_16942;
assign x_16944 = x_16941 & x_16943;
assign x_16945 = x_16939 & x_16944;
assign x_16946 = x_5701 & x_5702;
assign x_16947 = x_5704 & x_5705;
assign x_16948 = x_5703 & x_16947;
assign x_16949 = x_16946 & x_16948;
assign x_16950 = x_5707 & x_5708;
assign x_16951 = x_5706 & x_16950;
assign x_16952 = x_5710 & x_5711;
assign x_16953 = x_5709 & x_16952;
assign x_16954 = x_16951 & x_16953;
assign x_16955 = x_16949 & x_16954;
assign x_16956 = x_16945 & x_16955;
assign x_16957 = x_16935 & x_16956;
assign x_16958 = x_16914 & x_16957;
assign x_16959 = x_5712 & x_5713;
assign x_16960 = x_5715 & x_5716;
assign x_16961 = x_5714 & x_16960;
assign x_16962 = x_16959 & x_16961;
assign x_16963 = x_5718 & x_5719;
assign x_16964 = x_5717 & x_16963;
assign x_16965 = x_5721 & x_5722;
assign x_16966 = x_5720 & x_16965;
assign x_16967 = x_16964 & x_16966;
assign x_16968 = x_16962 & x_16967;
assign x_16969 = x_5723 & x_5724;
assign x_16970 = x_5726 & x_5727;
assign x_16971 = x_5725 & x_16970;
assign x_16972 = x_16969 & x_16971;
assign x_16973 = x_5729 & x_5730;
assign x_16974 = x_5728 & x_16973;
assign x_16975 = x_5732 & x_5733;
assign x_16976 = x_5731 & x_16975;
assign x_16977 = x_16974 & x_16976;
assign x_16978 = x_16972 & x_16977;
assign x_16979 = x_16968 & x_16978;
assign x_16980 = x_5734 & x_5735;
assign x_16981 = x_5737 & x_5738;
assign x_16982 = x_5736 & x_16981;
assign x_16983 = x_16980 & x_16982;
assign x_16984 = x_5740 & x_5741;
assign x_16985 = x_5739 & x_16984;
assign x_16986 = x_5743 & x_5744;
assign x_16987 = x_5742 & x_16986;
assign x_16988 = x_16985 & x_16987;
assign x_16989 = x_16983 & x_16988;
assign x_16990 = x_5745 & x_5746;
assign x_16991 = x_5748 & x_5749;
assign x_16992 = x_5747 & x_16991;
assign x_16993 = x_16990 & x_16992;
assign x_16994 = x_5751 & x_5752;
assign x_16995 = x_5750 & x_16994;
assign x_16996 = x_5754 & x_5755;
assign x_16997 = x_5753 & x_16996;
assign x_16998 = x_16995 & x_16997;
assign x_16999 = x_16993 & x_16998;
assign x_17000 = x_16989 & x_16999;
assign x_17001 = x_16979 & x_17000;
assign x_17002 = x_5756 & x_5757;
assign x_17003 = x_5759 & x_5760;
assign x_17004 = x_5758 & x_17003;
assign x_17005 = x_17002 & x_17004;
assign x_17006 = x_5762 & x_5763;
assign x_17007 = x_5761 & x_17006;
assign x_17008 = x_5765 & x_5766;
assign x_17009 = x_5764 & x_17008;
assign x_17010 = x_17007 & x_17009;
assign x_17011 = x_17005 & x_17010;
assign x_17012 = x_5767 & x_5768;
assign x_17013 = x_5770 & x_5771;
assign x_17014 = x_5769 & x_17013;
assign x_17015 = x_17012 & x_17014;
assign x_17016 = x_5773 & x_5774;
assign x_17017 = x_5772 & x_17016;
assign x_17018 = x_5776 & x_5777;
assign x_17019 = x_5775 & x_17018;
assign x_17020 = x_17017 & x_17019;
assign x_17021 = x_17015 & x_17020;
assign x_17022 = x_17011 & x_17021;
assign x_17023 = x_5778 & x_5779;
assign x_17024 = x_5781 & x_5782;
assign x_17025 = x_5780 & x_17024;
assign x_17026 = x_17023 & x_17025;
assign x_17027 = x_5784 & x_5785;
assign x_17028 = x_5783 & x_17027;
assign x_17029 = x_5787 & x_5788;
assign x_17030 = x_5786 & x_17029;
assign x_17031 = x_17028 & x_17030;
assign x_17032 = x_17026 & x_17031;
assign x_17033 = x_5789 & x_5790;
assign x_17034 = x_5792 & x_5793;
assign x_17035 = x_5791 & x_17034;
assign x_17036 = x_17033 & x_17035;
assign x_17037 = x_5795 & x_5796;
assign x_17038 = x_5794 & x_17037;
assign x_17039 = x_5798 & x_5799;
assign x_17040 = x_5797 & x_17039;
assign x_17041 = x_17038 & x_17040;
assign x_17042 = x_17036 & x_17041;
assign x_17043 = x_17032 & x_17042;
assign x_17044 = x_17022 & x_17043;
assign x_17045 = x_17001 & x_17044;
assign x_17046 = x_16958 & x_17045;
assign x_17047 = x_5800 & x_5801;
assign x_17048 = x_5803 & x_5804;
assign x_17049 = x_5802 & x_17048;
assign x_17050 = x_17047 & x_17049;
assign x_17051 = x_5806 & x_5807;
assign x_17052 = x_5805 & x_17051;
assign x_17053 = x_5809 & x_5810;
assign x_17054 = x_5808 & x_17053;
assign x_17055 = x_17052 & x_17054;
assign x_17056 = x_17050 & x_17055;
assign x_17057 = x_5811 & x_5812;
assign x_17058 = x_5814 & x_5815;
assign x_17059 = x_5813 & x_17058;
assign x_17060 = x_17057 & x_17059;
assign x_17061 = x_5817 & x_5818;
assign x_17062 = x_5816 & x_17061;
assign x_17063 = x_5820 & x_5821;
assign x_17064 = x_5819 & x_17063;
assign x_17065 = x_17062 & x_17064;
assign x_17066 = x_17060 & x_17065;
assign x_17067 = x_17056 & x_17066;
assign x_17068 = x_5822 & x_5823;
assign x_17069 = x_5825 & x_5826;
assign x_17070 = x_5824 & x_17069;
assign x_17071 = x_17068 & x_17070;
assign x_17072 = x_5828 & x_5829;
assign x_17073 = x_5827 & x_17072;
assign x_17074 = x_5831 & x_5832;
assign x_17075 = x_5830 & x_17074;
assign x_17076 = x_17073 & x_17075;
assign x_17077 = x_17071 & x_17076;
assign x_17078 = x_5833 & x_5834;
assign x_17079 = x_5836 & x_5837;
assign x_17080 = x_5835 & x_17079;
assign x_17081 = x_17078 & x_17080;
assign x_17082 = x_5839 & x_5840;
assign x_17083 = x_5838 & x_17082;
assign x_17084 = x_5842 & x_5843;
assign x_17085 = x_5841 & x_17084;
assign x_17086 = x_17083 & x_17085;
assign x_17087 = x_17081 & x_17086;
assign x_17088 = x_17077 & x_17087;
assign x_17089 = x_17067 & x_17088;
assign x_17090 = x_5844 & x_5845;
assign x_17091 = x_5847 & x_5848;
assign x_17092 = x_5846 & x_17091;
assign x_17093 = x_17090 & x_17092;
assign x_17094 = x_5850 & x_5851;
assign x_17095 = x_5849 & x_17094;
assign x_17096 = x_5853 & x_5854;
assign x_17097 = x_5852 & x_17096;
assign x_17098 = x_17095 & x_17097;
assign x_17099 = x_17093 & x_17098;
assign x_17100 = x_5855 & x_5856;
assign x_17101 = x_5858 & x_5859;
assign x_17102 = x_5857 & x_17101;
assign x_17103 = x_17100 & x_17102;
assign x_17104 = x_5861 & x_5862;
assign x_17105 = x_5860 & x_17104;
assign x_17106 = x_5864 & x_5865;
assign x_17107 = x_5863 & x_17106;
assign x_17108 = x_17105 & x_17107;
assign x_17109 = x_17103 & x_17108;
assign x_17110 = x_17099 & x_17109;
assign x_17111 = x_5866 & x_5867;
assign x_17112 = x_5869 & x_5870;
assign x_17113 = x_5868 & x_17112;
assign x_17114 = x_17111 & x_17113;
assign x_17115 = x_5872 & x_5873;
assign x_17116 = x_5871 & x_17115;
assign x_17117 = x_5875 & x_5876;
assign x_17118 = x_5874 & x_17117;
assign x_17119 = x_17116 & x_17118;
assign x_17120 = x_17114 & x_17119;
assign x_17121 = x_5877 & x_5878;
assign x_17122 = x_5880 & x_5881;
assign x_17123 = x_5879 & x_17122;
assign x_17124 = x_17121 & x_17123;
assign x_17125 = x_5883 & x_5884;
assign x_17126 = x_5882 & x_17125;
assign x_17127 = x_5886 & x_5887;
assign x_17128 = x_5885 & x_17127;
assign x_17129 = x_17126 & x_17128;
assign x_17130 = x_17124 & x_17129;
assign x_17131 = x_17120 & x_17130;
assign x_17132 = x_17110 & x_17131;
assign x_17133 = x_17089 & x_17132;
assign x_17134 = x_5888 & x_5889;
assign x_17135 = x_5891 & x_5892;
assign x_17136 = x_5890 & x_17135;
assign x_17137 = x_17134 & x_17136;
assign x_17138 = x_5894 & x_5895;
assign x_17139 = x_5893 & x_17138;
assign x_17140 = x_5897 & x_5898;
assign x_17141 = x_5896 & x_17140;
assign x_17142 = x_17139 & x_17141;
assign x_17143 = x_17137 & x_17142;
assign x_17144 = x_5899 & x_5900;
assign x_17145 = x_5902 & x_5903;
assign x_17146 = x_5901 & x_17145;
assign x_17147 = x_17144 & x_17146;
assign x_17148 = x_5905 & x_5906;
assign x_17149 = x_5904 & x_17148;
assign x_17150 = x_5908 & x_5909;
assign x_17151 = x_5907 & x_17150;
assign x_17152 = x_17149 & x_17151;
assign x_17153 = x_17147 & x_17152;
assign x_17154 = x_17143 & x_17153;
assign x_17155 = x_5910 & x_5911;
assign x_17156 = x_5913 & x_5914;
assign x_17157 = x_5912 & x_17156;
assign x_17158 = x_17155 & x_17157;
assign x_17159 = x_5916 & x_5917;
assign x_17160 = x_5915 & x_17159;
assign x_17161 = x_5919 & x_5920;
assign x_17162 = x_5918 & x_17161;
assign x_17163 = x_17160 & x_17162;
assign x_17164 = x_17158 & x_17163;
assign x_17165 = x_5921 & x_5922;
assign x_17166 = x_5924 & x_5925;
assign x_17167 = x_5923 & x_17166;
assign x_17168 = x_17165 & x_17167;
assign x_17169 = x_5927 & x_5928;
assign x_17170 = x_5926 & x_17169;
assign x_17171 = x_5930 & x_5931;
assign x_17172 = x_5929 & x_17171;
assign x_17173 = x_17170 & x_17172;
assign x_17174 = x_17168 & x_17173;
assign x_17175 = x_17164 & x_17174;
assign x_17176 = x_17154 & x_17175;
assign x_17177 = x_5932 & x_5933;
assign x_17178 = x_5935 & x_5936;
assign x_17179 = x_5934 & x_17178;
assign x_17180 = x_17177 & x_17179;
assign x_17181 = x_5938 & x_5939;
assign x_17182 = x_5937 & x_17181;
assign x_17183 = x_5941 & x_5942;
assign x_17184 = x_5940 & x_17183;
assign x_17185 = x_17182 & x_17184;
assign x_17186 = x_17180 & x_17185;
assign x_17187 = x_5943 & x_5944;
assign x_17188 = x_5946 & x_5947;
assign x_17189 = x_5945 & x_17188;
assign x_17190 = x_17187 & x_17189;
assign x_17191 = x_5949 & x_5950;
assign x_17192 = x_5948 & x_17191;
assign x_17193 = x_5952 & x_5953;
assign x_17194 = x_5951 & x_17193;
assign x_17195 = x_17192 & x_17194;
assign x_17196 = x_17190 & x_17195;
assign x_17197 = x_17186 & x_17196;
assign x_17198 = x_5954 & x_5955;
assign x_17199 = x_5957 & x_5958;
assign x_17200 = x_5956 & x_17199;
assign x_17201 = x_17198 & x_17200;
assign x_17202 = x_5960 & x_5961;
assign x_17203 = x_5959 & x_17202;
assign x_17204 = x_5963 & x_5964;
assign x_17205 = x_5962 & x_17204;
assign x_17206 = x_17203 & x_17205;
assign x_17207 = x_17201 & x_17206;
assign x_17208 = x_5965 & x_5966;
assign x_17209 = x_5968 & x_5969;
assign x_17210 = x_5967 & x_17209;
assign x_17211 = x_17208 & x_17210;
assign x_17212 = x_5971 & x_5972;
assign x_17213 = x_5970 & x_17212;
assign x_17214 = x_5974 & x_5975;
assign x_17215 = x_5973 & x_17214;
assign x_17216 = x_17213 & x_17215;
assign x_17217 = x_17211 & x_17216;
assign x_17218 = x_17207 & x_17217;
assign x_17219 = x_17197 & x_17218;
assign x_17220 = x_17176 & x_17219;
assign x_17221 = x_17133 & x_17220;
assign x_17222 = x_17046 & x_17221;
assign x_17223 = x_5976 & x_5977;
assign x_17224 = x_5979 & x_5980;
assign x_17225 = x_5978 & x_17224;
assign x_17226 = x_17223 & x_17225;
assign x_17227 = x_5982 & x_5983;
assign x_17228 = x_5981 & x_17227;
assign x_17229 = x_5985 & x_5986;
assign x_17230 = x_5984 & x_17229;
assign x_17231 = x_17228 & x_17230;
assign x_17232 = x_17226 & x_17231;
assign x_17233 = x_5987 & x_5988;
assign x_17234 = x_5990 & x_5991;
assign x_17235 = x_5989 & x_17234;
assign x_17236 = x_17233 & x_17235;
assign x_17237 = x_5993 & x_5994;
assign x_17238 = x_5992 & x_17237;
assign x_17239 = x_5996 & x_5997;
assign x_17240 = x_5995 & x_17239;
assign x_17241 = x_17238 & x_17240;
assign x_17242 = x_17236 & x_17241;
assign x_17243 = x_17232 & x_17242;
assign x_17244 = x_5998 & x_5999;
assign x_17245 = x_6001 & x_6002;
assign x_17246 = x_6000 & x_17245;
assign x_17247 = x_17244 & x_17246;
assign x_17248 = x_6004 & x_6005;
assign x_17249 = x_6003 & x_17248;
assign x_17250 = x_6007 & x_6008;
assign x_17251 = x_6006 & x_17250;
assign x_17252 = x_17249 & x_17251;
assign x_17253 = x_17247 & x_17252;
assign x_17254 = x_6009 & x_6010;
assign x_17255 = x_6012 & x_6013;
assign x_17256 = x_6011 & x_17255;
assign x_17257 = x_17254 & x_17256;
assign x_17258 = x_6015 & x_6016;
assign x_17259 = x_6014 & x_17258;
assign x_17260 = x_6018 & x_6019;
assign x_17261 = x_6017 & x_17260;
assign x_17262 = x_17259 & x_17261;
assign x_17263 = x_17257 & x_17262;
assign x_17264 = x_17253 & x_17263;
assign x_17265 = x_17243 & x_17264;
assign x_17266 = x_6020 & x_6021;
assign x_17267 = x_6023 & x_6024;
assign x_17268 = x_6022 & x_17267;
assign x_17269 = x_17266 & x_17268;
assign x_17270 = x_6026 & x_6027;
assign x_17271 = x_6025 & x_17270;
assign x_17272 = x_6029 & x_6030;
assign x_17273 = x_6028 & x_17272;
assign x_17274 = x_17271 & x_17273;
assign x_17275 = x_17269 & x_17274;
assign x_17276 = x_6031 & x_6032;
assign x_17277 = x_6034 & x_6035;
assign x_17278 = x_6033 & x_17277;
assign x_17279 = x_17276 & x_17278;
assign x_17280 = x_6037 & x_6038;
assign x_17281 = x_6036 & x_17280;
assign x_17282 = x_6040 & x_6041;
assign x_17283 = x_6039 & x_17282;
assign x_17284 = x_17281 & x_17283;
assign x_17285 = x_17279 & x_17284;
assign x_17286 = x_17275 & x_17285;
assign x_17287 = x_6042 & x_6043;
assign x_17288 = x_6045 & x_6046;
assign x_17289 = x_6044 & x_17288;
assign x_17290 = x_17287 & x_17289;
assign x_17291 = x_6048 & x_6049;
assign x_17292 = x_6047 & x_17291;
assign x_17293 = x_6051 & x_6052;
assign x_17294 = x_6050 & x_17293;
assign x_17295 = x_17292 & x_17294;
assign x_17296 = x_17290 & x_17295;
assign x_17297 = x_6053 & x_6054;
assign x_17298 = x_6056 & x_6057;
assign x_17299 = x_6055 & x_17298;
assign x_17300 = x_17297 & x_17299;
assign x_17301 = x_6059 & x_6060;
assign x_17302 = x_6058 & x_17301;
assign x_17303 = x_6062 & x_6063;
assign x_17304 = x_6061 & x_17303;
assign x_17305 = x_17302 & x_17304;
assign x_17306 = x_17300 & x_17305;
assign x_17307 = x_17296 & x_17306;
assign x_17308 = x_17286 & x_17307;
assign x_17309 = x_17265 & x_17308;
assign x_17310 = x_6064 & x_6065;
assign x_17311 = x_6067 & x_6068;
assign x_17312 = x_6066 & x_17311;
assign x_17313 = x_17310 & x_17312;
assign x_17314 = x_6070 & x_6071;
assign x_17315 = x_6069 & x_17314;
assign x_17316 = x_6073 & x_6074;
assign x_17317 = x_6072 & x_17316;
assign x_17318 = x_17315 & x_17317;
assign x_17319 = x_17313 & x_17318;
assign x_17320 = x_6075 & x_6076;
assign x_17321 = x_6078 & x_6079;
assign x_17322 = x_6077 & x_17321;
assign x_17323 = x_17320 & x_17322;
assign x_17324 = x_6081 & x_6082;
assign x_17325 = x_6080 & x_17324;
assign x_17326 = x_6084 & x_6085;
assign x_17327 = x_6083 & x_17326;
assign x_17328 = x_17325 & x_17327;
assign x_17329 = x_17323 & x_17328;
assign x_17330 = x_17319 & x_17329;
assign x_17331 = x_6086 & x_6087;
assign x_17332 = x_6089 & x_6090;
assign x_17333 = x_6088 & x_17332;
assign x_17334 = x_17331 & x_17333;
assign x_17335 = x_6092 & x_6093;
assign x_17336 = x_6091 & x_17335;
assign x_17337 = x_6095 & x_6096;
assign x_17338 = x_6094 & x_17337;
assign x_17339 = x_17336 & x_17338;
assign x_17340 = x_17334 & x_17339;
assign x_17341 = x_6097 & x_6098;
assign x_17342 = x_6100 & x_6101;
assign x_17343 = x_6099 & x_17342;
assign x_17344 = x_17341 & x_17343;
assign x_17345 = x_6103 & x_6104;
assign x_17346 = x_6102 & x_17345;
assign x_17347 = x_6106 & x_6107;
assign x_17348 = x_6105 & x_17347;
assign x_17349 = x_17346 & x_17348;
assign x_17350 = x_17344 & x_17349;
assign x_17351 = x_17340 & x_17350;
assign x_17352 = x_17330 & x_17351;
assign x_17353 = x_6108 & x_6109;
assign x_17354 = x_6111 & x_6112;
assign x_17355 = x_6110 & x_17354;
assign x_17356 = x_17353 & x_17355;
assign x_17357 = x_6114 & x_6115;
assign x_17358 = x_6113 & x_17357;
assign x_17359 = x_6117 & x_6118;
assign x_17360 = x_6116 & x_17359;
assign x_17361 = x_17358 & x_17360;
assign x_17362 = x_17356 & x_17361;
assign x_17363 = x_6119 & x_6120;
assign x_17364 = x_6122 & x_6123;
assign x_17365 = x_6121 & x_17364;
assign x_17366 = x_17363 & x_17365;
assign x_17367 = x_6125 & x_6126;
assign x_17368 = x_6124 & x_17367;
assign x_17369 = x_6128 & x_6129;
assign x_17370 = x_6127 & x_17369;
assign x_17371 = x_17368 & x_17370;
assign x_17372 = x_17366 & x_17371;
assign x_17373 = x_17362 & x_17372;
assign x_17374 = x_6130 & x_6131;
assign x_17375 = x_6133 & x_6134;
assign x_17376 = x_6132 & x_17375;
assign x_17377 = x_17374 & x_17376;
assign x_17378 = x_6136 & x_6137;
assign x_17379 = x_6135 & x_17378;
assign x_17380 = x_6139 & x_6140;
assign x_17381 = x_6138 & x_17380;
assign x_17382 = x_17379 & x_17381;
assign x_17383 = x_17377 & x_17382;
assign x_17384 = x_6141 & x_6142;
assign x_17385 = x_6144 & x_6145;
assign x_17386 = x_6143 & x_17385;
assign x_17387 = x_17384 & x_17386;
assign x_17388 = x_6147 & x_6148;
assign x_17389 = x_6146 & x_17388;
assign x_17390 = x_6150 & x_6151;
assign x_17391 = x_6149 & x_17390;
assign x_17392 = x_17389 & x_17391;
assign x_17393 = x_17387 & x_17392;
assign x_17394 = x_17383 & x_17393;
assign x_17395 = x_17373 & x_17394;
assign x_17396 = x_17352 & x_17395;
assign x_17397 = x_17309 & x_17396;
assign x_17398 = x_6152 & x_6153;
assign x_17399 = x_6155 & x_6156;
assign x_17400 = x_6154 & x_17399;
assign x_17401 = x_17398 & x_17400;
assign x_17402 = x_6158 & x_6159;
assign x_17403 = x_6157 & x_17402;
assign x_17404 = x_6161 & x_6162;
assign x_17405 = x_6160 & x_17404;
assign x_17406 = x_17403 & x_17405;
assign x_17407 = x_17401 & x_17406;
assign x_17408 = x_6163 & x_6164;
assign x_17409 = x_6166 & x_6167;
assign x_17410 = x_6165 & x_17409;
assign x_17411 = x_17408 & x_17410;
assign x_17412 = x_6169 & x_6170;
assign x_17413 = x_6168 & x_17412;
assign x_17414 = x_6172 & x_6173;
assign x_17415 = x_6171 & x_17414;
assign x_17416 = x_17413 & x_17415;
assign x_17417 = x_17411 & x_17416;
assign x_17418 = x_17407 & x_17417;
assign x_17419 = x_6174 & x_6175;
assign x_17420 = x_6177 & x_6178;
assign x_17421 = x_6176 & x_17420;
assign x_17422 = x_17419 & x_17421;
assign x_17423 = x_6180 & x_6181;
assign x_17424 = x_6179 & x_17423;
assign x_17425 = x_6183 & x_6184;
assign x_17426 = x_6182 & x_17425;
assign x_17427 = x_17424 & x_17426;
assign x_17428 = x_17422 & x_17427;
assign x_17429 = x_6185 & x_6186;
assign x_17430 = x_6188 & x_6189;
assign x_17431 = x_6187 & x_17430;
assign x_17432 = x_17429 & x_17431;
assign x_17433 = x_6191 & x_6192;
assign x_17434 = x_6190 & x_17433;
assign x_17435 = x_6194 & x_6195;
assign x_17436 = x_6193 & x_17435;
assign x_17437 = x_17434 & x_17436;
assign x_17438 = x_17432 & x_17437;
assign x_17439 = x_17428 & x_17438;
assign x_17440 = x_17418 & x_17439;
assign x_17441 = x_6196 & x_6197;
assign x_17442 = x_6199 & x_6200;
assign x_17443 = x_6198 & x_17442;
assign x_17444 = x_17441 & x_17443;
assign x_17445 = x_6202 & x_6203;
assign x_17446 = x_6201 & x_17445;
assign x_17447 = x_6205 & x_6206;
assign x_17448 = x_6204 & x_17447;
assign x_17449 = x_17446 & x_17448;
assign x_17450 = x_17444 & x_17449;
assign x_17451 = x_6207 & x_6208;
assign x_17452 = x_6210 & x_6211;
assign x_17453 = x_6209 & x_17452;
assign x_17454 = x_17451 & x_17453;
assign x_17455 = x_6213 & x_6214;
assign x_17456 = x_6212 & x_17455;
assign x_17457 = x_6216 & x_6217;
assign x_17458 = x_6215 & x_17457;
assign x_17459 = x_17456 & x_17458;
assign x_17460 = x_17454 & x_17459;
assign x_17461 = x_17450 & x_17460;
assign x_17462 = x_6218 & x_6219;
assign x_17463 = x_6221 & x_6222;
assign x_17464 = x_6220 & x_17463;
assign x_17465 = x_17462 & x_17464;
assign x_17466 = x_6224 & x_6225;
assign x_17467 = x_6223 & x_17466;
assign x_17468 = x_6227 & x_6228;
assign x_17469 = x_6226 & x_17468;
assign x_17470 = x_17467 & x_17469;
assign x_17471 = x_17465 & x_17470;
assign x_17472 = x_6229 & x_6230;
assign x_17473 = x_6232 & x_6233;
assign x_17474 = x_6231 & x_17473;
assign x_17475 = x_17472 & x_17474;
assign x_17476 = x_6235 & x_6236;
assign x_17477 = x_6234 & x_17476;
assign x_17478 = x_6238 & x_6239;
assign x_17479 = x_6237 & x_17478;
assign x_17480 = x_17477 & x_17479;
assign x_17481 = x_17475 & x_17480;
assign x_17482 = x_17471 & x_17481;
assign x_17483 = x_17461 & x_17482;
assign x_17484 = x_17440 & x_17483;
assign x_17485 = x_6240 & x_6241;
assign x_17486 = x_6243 & x_6244;
assign x_17487 = x_6242 & x_17486;
assign x_17488 = x_17485 & x_17487;
assign x_17489 = x_6246 & x_6247;
assign x_17490 = x_6245 & x_17489;
assign x_17491 = x_6249 & x_6250;
assign x_17492 = x_6248 & x_17491;
assign x_17493 = x_17490 & x_17492;
assign x_17494 = x_17488 & x_17493;
assign x_17495 = x_6251 & x_6252;
assign x_17496 = x_6254 & x_6255;
assign x_17497 = x_6253 & x_17496;
assign x_17498 = x_17495 & x_17497;
assign x_17499 = x_6257 & x_6258;
assign x_17500 = x_6256 & x_17499;
assign x_17501 = x_6260 & x_6261;
assign x_17502 = x_6259 & x_17501;
assign x_17503 = x_17500 & x_17502;
assign x_17504 = x_17498 & x_17503;
assign x_17505 = x_17494 & x_17504;
assign x_17506 = x_6262 & x_6263;
assign x_17507 = x_6265 & x_6266;
assign x_17508 = x_6264 & x_17507;
assign x_17509 = x_17506 & x_17508;
assign x_17510 = x_6268 & x_6269;
assign x_17511 = x_6267 & x_17510;
assign x_17512 = x_6271 & x_6272;
assign x_17513 = x_6270 & x_17512;
assign x_17514 = x_17511 & x_17513;
assign x_17515 = x_17509 & x_17514;
assign x_17516 = x_6273 & x_6274;
assign x_17517 = x_6276 & x_6277;
assign x_17518 = x_6275 & x_17517;
assign x_17519 = x_17516 & x_17518;
assign x_17520 = x_6279 & x_6280;
assign x_17521 = x_6278 & x_17520;
assign x_17522 = x_6282 & x_6283;
assign x_17523 = x_6281 & x_17522;
assign x_17524 = x_17521 & x_17523;
assign x_17525 = x_17519 & x_17524;
assign x_17526 = x_17515 & x_17525;
assign x_17527 = x_17505 & x_17526;
assign x_17528 = x_6284 & x_6285;
assign x_17529 = x_6287 & x_6288;
assign x_17530 = x_6286 & x_17529;
assign x_17531 = x_17528 & x_17530;
assign x_17532 = x_6290 & x_6291;
assign x_17533 = x_6289 & x_17532;
assign x_17534 = x_6293 & x_6294;
assign x_17535 = x_6292 & x_17534;
assign x_17536 = x_17533 & x_17535;
assign x_17537 = x_17531 & x_17536;
assign x_17538 = x_6295 & x_6296;
assign x_17539 = x_6298 & x_6299;
assign x_17540 = x_6297 & x_17539;
assign x_17541 = x_17538 & x_17540;
assign x_17542 = x_6301 & x_6302;
assign x_17543 = x_6300 & x_17542;
assign x_17544 = x_6304 & x_6305;
assign x_17545 = x_6303 & x_17544;
assign x_17546 = x_17543 & x_17545;
assign x_17547 = x_17541 & x_17546;
assign x_17548 = x_17537 & x_17547;
assign x_17549 = x_6306 & x_6307;
assign x_17550 = x_6309 & x_6310;
assign x_17551 = x_6308 & x_17550;
assign x_17552 = x_17549 & x_17551;
assign x_17553 = x_6312 & x_6313;
assign x_17554 = x_6311 & x_17553;
assign x_17555 = x_6315 & x_6316;
assign x_17556 = x_6314 & x_17555;
assign x_17557 = x_17554 & x_17556;
assign x_17558 = x_17552 & x_17557;
assign x_17559 = x_6317 & x_6318;
assign x_17560 = x_6320 & x_6321;
assign x_17561 = x_6319 & x_17560;
assign x_17562 = x_17559 & x_17561;
assign x_17563 = x_6323 & x_6324;
assign x_17564 = x_6322 & x_17563;
assign x_17565 = x_6326 & x_6327;
assign x_17566 = x_6325 & x_17565;
assign x_17567 = x_17564 & x_17566;
assign x_17568 = x_17562 & x_17567;
assign x_17569 = x_17558 & x_17568;
assign x_17570 = x_17548 & x_17569;
assign x_17571 = x_17527 & x_17570;
assign x_17572 = x_17484 & x_17571;
assign x_17573 = x_17397 & x_17572;
assign x_17574 = x_17222 & x_17573;
assign x_17575 = x_6328 & x_6329;
assign x_17576 = x_6331 & x_6332;
assign x_17577 = x_6330 & x_17576;
assign x_17578 = x_17575 & x_17577;
assign x_17579 = x_6333 & x_6334;
assign x_17580 = x_6336 & x_6337;
assign x_17581 = x_6335 & x_17580;
assign x_17582 = x_17579 & x_17581;
assign x_17583 = x_17578 & x_17582;
assign x_17584 = x_6338 & x_6339;
assign x_17585 = x_6341 & x_6342;
assign x_17586 = x_6340 & x_17585;
assign x_17587 = x_17584 & x_17586;
assign x_17588 = x_6344 & x_6345;
assign x_17589 = x_6343 & x_17588;
assign x_17590 = x_6347 & x_6348;
assign x_17591 = x_6346 & x_17590;
assign x_17592 = x_17589 & x_17591;
assign x_17593 = x_17587 & x_17592;
assign x_17594 = x_17583 & x_17593;
assign x_17595 = x_6349 & x_6350;
assign x_17596 = x_6352 & x_6353;
assign x_17597 = x_6351 & x_17596;
assign x_17598 = x_17595 & x_17597;
assign x_17599 = x_6355 & x_6356;
assign x_17600 = x_6354 & x_17599;
assign x_17601 = x_6358 & x_6359;
assign x_17602 = x_6357 & x_17601;
assign x_17603 = x_17600 & x_17602;
assign x_17604 = x_17598 & x_17603;
assign x_17605 = x_6360 & x_6361;
assign x_17606 = x_6363 & x_6364;
assign x_17607 = x_6362 & x_17606;
assign x_17608 = x_17605 & x_17607;
assign x_17609 = x_6366 & x_6367;
assign x_17610 = x_6365 & x_17609;
assign x_17611 = x_6369 & x_6370;
assign x_17612 = x_6368 & x_17611;
assign x_17613 = x_17610 & x_17612;
assign x_17614 = x_17608 & x_17613;
assign x_17615 = x_17604 & x_17614;
assign x_17616 = x_17594 & x_17615;
assign x_17617 = x_6371 & x_6372;
assign x_17618 = x_6374 & x_6375;
assign x_17619 = x_6373 & x_17618;
assign x_17620 = x_17617 & x_17619;
assign x_17621 = x_6377 & x_6378;
assign x_17622 = x_6376 & x_17621;
assign x_17623 = x_6380 & x_6381;
assign x_17624 = x_6379 & x_17623;
assign x_17625 = x_17622 & x_17624;
assign x_17626 = x_17620 & x_17625;
assign x_17627 = x_6382 & x_6383;
assign x_17628 = x_6385 & x_6386;
assign x_17629 = x_6384 & x_17628;
assign x_17630 = x_17627 & x_17629;
assign x_17631 = x_6388 & x_6389;
assign x_17632 = x_6387 & x_17631;
assign x_17633 = x_6391 & x_6392;
assign x_17634 = x_6390 & x_17633;
assign x_17635 = x_17632 & x_17634;
assign x_17636 = x_17630 & x_17635;
assign x_17637 = x_17626 & x_17636;
assign x_17638 = x_6393 & x_6394;
assign x_17639 = x_6396 & x_6397;
assign x_17640 = x_6395 & x_17639;
assign x_17641 = x_17638 & x_17640;
assign x_17642 = x_6399 & x_6400;
assign x_17643 = x_6398 & x_17642;
assign x_17644 = x_6402 & x_6403;
assign x_17645 = x_6401 & x_17644;
assign x_17646 = x_17643 & x_17645;
assign x_17647 = x_17641 & x_17646;
assign x_17648 = x_6404 & x_6405;
assign x_17649 = x_6407 & x_6408;
assign x_17650 = x_6406 & x_17649;
assign x_17651 = x_17648 & x_17650;
assign x_17652 = x_6410 & x_6411;
assign x_17653 = x_6409 & x_17652;
assign x_17654 = x_6413 & x_6414;
assign x_17655 = x_6412 & x_17654;
assign x_17656 = x_17653 & x_17655;
assign x_17657 = x_17651 & x_17656;
assign x_17658 = x_17647 & x_17657;
assign x_17659 = x_17637 & x_17658;
assign x_17660 = x_17616 & x_17659;
assign x_17661 = x_6415 & x_6416;
assign x_17662 = x_6418 & x_6419;
assign x_17663 = x_6417 & x_17662;
assign x_17664 = x_17661 & x_17663;
assign x_17665 = x_6421 & x_6422;
assign x_17666 = x_6420 & x_17665;
assign x_17667 = x_6424 & x_6425;
assign x_17668 = x_6423 & x_17667;
assign x_17669 = x_17666 & x_17668;
assign x_17670 = x_17664 & x_17669;
assign x_17671 = x_6426 & x_6427;
assign x_17672 = x_6429 & x_6430;
assign x_17673 = x_6428 & x_17672;
assign x_17674 = x_17671 & x_17673;
assign x_17675 = x_6432 & x_6433;
assign x_17676 = x_6431 & x_17675;
assign x_17677 = x_6435 & x_6436;
assign x_17678 = x_6434 & x_17677;
assign x_17679 = x_17676 & x_17678;
assign x_17680 = x_17674 & x_17679;
assign x_17681 = x_17670 & x_17680;
assign x_17682 = x_6437 & x_6438;
assign x_17683 = x_6440 & x_6441;
assign x_17684 = x_6439 & x_17683;
assign x_17685 = x_17682 & x_17684;
assign x_17686 = x_6443 & x_6444;
assign x_17687 = x_6442 & x_17686;
assign x_17688 = x_6446 & x_6447;
assign x_17689 = x_6445 & x_17688;
assign x_17690 = x_17687 & x_17689;
assign x_17691 = x_17685 & x_17690;
assign x_17692 = x_6448 & x_6449;
assign x_17693 = x_6451 & x_6452;
assign x_17694 = x_6450 & x_17693;
assign x_17695 = x_17692 & x_17694;
assign x_17696 = x_6454 & x_6455;
assign x_17697 = x_6453 & x_17696;
assign x_17698 = x_6457 & x_6458;
assign x_17699 = x_6456 & x_17698;
assign x_17700 = x_17697 & x_17699;
assign x_17701 = x_17695 & x_17700;
assign x_17702 = x_17691 & x_17701;
assign x_17703 = x_17681 & x_17702;
assign x_17704 = x_6459 & x_6460;
assign x_17705 = x_6462 & x_6463;
assign x_17706 = x_6461 & x_17705;
assign x_17707 = x_17704 & x_17706;
assign x_17708 = x_6465 & x_6466;
assign x_17709 = x_6464 & x_17708;
assign x_17710 = x_6468 & x_6469;
assign x_17711 = x_6467 & x_17710;
assign x_17712 = x_17709 & x_17711;
assign x_17713 = x_17707 & x_17712;
assign x_17714 = x_6470 & x_6471;
assign x_17715 = x_6473 & x_6474;
assign x_17716 = x_6472 & x_17715;
assign x_17717 = x_17714 & x_17716;
assign x_17718 = x_6476 & x_6477;
assign x_17719 = x_6475 & x_17718;
assign x_17720 = x_6479 & x_6480;
assign x_17721 = x_6478 & x_17720;
assign x_17722 = x_17719 & x_17721;
assign x_17723 = x_17717 & x_17722;
assign x_17724 = x_17713 & x_17723;
assign x_17725 = x_6481 & x_6482;
assign x_17726 = x_6484 & x_6485;
assign x_17727 = x_6483 & x_17726;
assign x_17728 = x_17725 & x_17727;
assign x_17729 = x_6487 & x_6488;
assign x_17730 = x_6486 & x_17729;
assign x_17731 = x_6490 & x_6491;
assign x_17732 = x_6489 & x_17731;
assign x_17733 = x_17730 & x_17732;
assign x_17734 = x_17728 & x_17733;
assign x_17735 = x_6492 & x_6493;
assign x_17736 = x_6495 & x_6496;
assign x_17737 = x_6494 & x_17736;
assign x_17738 = x_17735 & x_17737;
assign x_17739 = x_6498 & x_6499;
assign x_17740 = x_6497 & x_17739;
assign x_17741 = x_6501 & x_6502;
assign x_17742 = x_6500 & x_17741;
assign x_17743 = x_17740 & x_17742;
assign x_17744 = x_17738 & x_17743;
assign x_17745 = x_17734 & x_17744;
assign x_17746 = x_17724 & x_17745;
assign x_17747 = x_17703 & x_17746;
assign x_17748 = x_17660 & x_17747;
assign x_17749 = x_6503 & x_6504;
assign x_17750 = x_6506 & x_6507;
assign x_17751 = x_6505 & x_17750;
assign x_17752 = x_17749 & x_17751;
assign x_17753 = x_6509 & x_6510;
assign x_17754 = x_6508 & x_17753;
assign x_17755 = x_6512 & x_6513;
assign x_17756 = x_6511 & x_17755;
assign x_17757 = x_17754 & x_17756;
assign x_17758 = x_17752 & x_17757;
assign x_17759 = x_6514 & x_6515;
assign x_17760 = x_6517 & x_6518;
assign x_17761 = x_6516 & x_17760;
assign x_17762 = x_17759 & x_17761;
assign x_17763 = x_6520 & x_6521;
assign x_17764 = x_6519 & x_17763;
assign x_17765 = x_6523 & x_6524;
assign x_17766 = x_6522 & x_17765;
assign x_17767 = x_17764 & x_17766;
assign x_17768 = x_17762 & x_17767;
assign x_17769 = x_17758 & x_17768;
assign x_17770 = x_6525 & x_6526;
assign x_17771 = x_6528 & x_6529;
assign x_17772 = x_6527 & x_17771;
assign x_17773 = x_17770 & x_17772;
assign x_17774 = x_6531 & x_6532;
assign x_17775 = x_6530 & x_17774;
assign x_17776 = x_6534 & x_6535;
assign x_17777 = x_6533 & x_17776;
assign x_17778 = x_17775 & x_17777;
assign x_17779 = x_17773 & x_17778;
assign x_17780 = x_6536 & x_6537;
assign x_17781 = x_6539 & x_6540;
assign x_17782 = x_6538 & x_17781;
assign x_17783 = x_17780 & x_17782;
assign x_17784 = x_6542 & x_6543;
assign x_17785 = x_6541 & x_17784;
assign x_17786 = x_6545 & x_6546;
assign x_17787 = x_6544 & x_17786;
assign x_17788 = x_17785 & x_17787;
assign x_17789 = x_17783 & x_17788;
assign x_17790 = x_17779 & x_17789;
assign x_17791 = x_17769 & x_17790;
assign x_17792 = x_6547 & x_6548;
assign x_17793 = x_6550 & x_6551;
assign x_17794 = x_6549 & x_17793;
assign x_17795 = x_17792 & x_17794;
assign x_17796 = x_6553 & x_6554;
assign x_17797 = x_6552 & x_17796;
assign x_17798 = x_6556 & x_6557;
assign x_17799 = x_6555 & x_17798;
assign x_17800 = x_17797 & x_17799;
assign x_17801 = x_17795 & x_17800;
assign x_17802 = x_6558 & x_6559;
assign x_17803 = x_6561 & x_6562;
assign x_17804 = x_6560 & x_17803;
assign x_17805 = x_17802 & x_17804;
assign x_17806 = x_6564 & x_6565;
assign x_17807 = x_6563 & x_17806;
assign x_17808 = x_6567 & x_6568;
assign x_17809 = x_6566 & x_17808;
assign x_17810 = x_17807 & x_17809;
assign x_17811 = x_17805 & x_17810;
assign x_17812 = x_17801 & x_17811;
assign x_17813 = x_6569 & x_6570;
assign x_17814 = x_6572 & x_6573;
assign x_17815 = x_6571 & x_17814;
assign x_17816 = x_17813 & x_17815;
assign x_17817 = x_6575 & x_6576;
assign x_17818 = x_6574 & x_17817;
assign x_17819 = x_6578 & x_6579;
assign x_17820 = x_6577 & x_17819;
assign x_17821 = x_17818 & x_17820;
assign x_17822 = x_17816 & x_17821;
assign x_17823 = x_6580 & x_6581;
assign x_17824 = x_6583 & x_6584;
assign x_17825 = x_6582 & x_17824;
assign x_17826 = x_17823 & x_17825;
assign x_17827 = x_6586 & x_6587;
assign x_17828 = x_6585 & x_17827;
assign x_17829 = x_6589 & x_6590;
assign x_17830 = x_6588 & x_17829;
assign x_17831 = x_17828 & x_17830;
assign x_17832 = x_17826 & x_17831;
assign x_17833 = x_17822 & x_17832;
assign x_17834 = x_17812 & x_17833;
assign x_17835 = x_17791 & x_17834;
assign x_17836 = x_6591 & x_6592;
assign x_17837 = x_6594 & x_6595;
assign x_17838 = x_6593 & x_17837;
assign x_17839 = x_17836 & x_17838;
assign x_17840 = x_6597 & x_6598;
assign x_17841 = x_6596 & x_17840;
assign x_17842 = x_6600 & x_6601;
assign x_17843 = x_6599 & x_17842;
assign x_17844 = x_17841 & x_17843;
assign x_17845 = x_17839 & x_17844;
assign x_17846 = x_6602 & x_6603;
assign x_17847 = x_6605 & x_6606;
assign x_17848 = x_6604 & x_17847;
assign x_17849 = x_17846 & x_17848;
assign x_17850 = x_6608 & x_6609;
assign x_17851 = x_6607 & x_17850;
assign x_17852 = x_6611 & x_6612;
assign x_17853 = x_6610 & x_17852;
assign x_17854 = x_17851 & x_17853;
assign x_17855 = x_17849 & x_17854;
assign x_17856 = x_17845 & x_17855;
assign x_17857 = x_6613 & x_6614;
assign x_17858 = x_6616 & x_6617;
assign x_17859 = x_6615 & x_17858;
assign x_17860 = x_17857 & x_17859;
assign x_17861 = x_6619 & x_6620;
assign x_17862 = x_6618 & x_17861;
assign x_17863 = x_6622 & x_6623;
assign x_17864 = x_6621 & x_17863;
assign x_17865 = x_17862 & x_17864;
assign x_17866 = x_17860 & x_17865;
assign x_17867 = x_6624 & x_6625;
assign x_17868 = x_6627 & x_6628;
assign x_17869 = x_6626 & x_17868;
assign x_17870 = x_17867 & x_17869;
assign x_17871 = x_6630 & x_6631;
assign x_17872 = x_6629 & x_17871;
assign x_17873 = x_6633 & x_6634;
assign x_17874 = x_6632 & x_17873;
assign x_17875 = x_17872 & x_17874;
assign x_17876 = x_17870 & x_17875;
assign x_17877 = x_17866 & x_17876;
assign x_17878 = x_17856 & x_17877;
assign x_17879 = x_6635 & x_6636;
assign x_17880 = x_6638 & x_6639;
assign x_17881 = x_6637 & x_17880;
assign x_17882 = x_17879 & x_17881;
assign x_17883 = x_6641 & x_6642;
assign x_17884 = x_6640 & x_17883;
assign x_17885 = x_6644 & x_6645;
assign x_17886 = x_6643 & x_17885;
assign x_17887 = x_17884 & x_17886;
assign x_17888 = x_17882 & x_17887;
assign x_17889 = x_6646 & x_6647;
assign x_17890 = x_6649 & x_6650;
assign x_17891 = x_6648 & x_17890;
assign x_17892 = x_17889 & x_17891;
assign x_17893 = x_6652 & x_6653;
assign x_17894 = x_6651 & x_17893;
assign x_17895 = x_6655 & x_6656;
assign x_17896 = x_6654 & x_17895;
assign x_17897 = x_17894 & x_17896;
assign x_17898 = x_17892 & x_17897;
assign x_17899 = x_17888 & x_17898;
assign x_17900 = x_6657 & x_6658;
assign x_17901 = x_6660 & x_6661;
assign x_17902 = x_6659 & x_17901;
assign x_17903 = x_17900 & x_17902;
assign x_17904 = x_6663 & x_6664;
assign x_17905 = x_6662 & x_17904;
assign x_17906 = x_6666 & x_6667;
assign x_17907 = x_6665 & x_17906;
assign x_17908 = x_17905 & x_17907;
assign x_17909 = x_17903 & x_17908;
assign x_17910 = x_6668 & x_6669;
assign x_17911 = x_6671 & x_6672;
assign x_17912 = x_6670 & x_17911;
assign x_17913 = x_17910 & x_17912;
assign x_17914 = x_6674 & x_6675;
assign x_17915 = x_6673 & x_17914;
assign x_17916 = x_6677 & x_6678;
assign x_17917 = x_6676 & x_17916;
assign x_17918 = x_17915 & x_17917;
assign x_17919 = x_17913 & x_17918;
assign x_17920 = x_17909 & x_17919;
assign x_17921 = x_17899 & x_17920;
assign x_17922 = x_17878 & x_17921;
assign x_17923 = x_17835 & x_17922;
assign x_17924 = x_17748 & x_17923;
assign x_17925 = x_6679 & x_6680;
assign x_17926 = x_6682 & x_6683;
assign x_17927 = x_6681 & x_17926;
assign x_17928 = x_17925 & x_17927;
assign x_17929 = x_6685 & x_6686;
assign x_17930 = x_6684 & x_17929;
assign x_17931 = x_6688 & x_6689;
assign x_17932 = x_6687 & x_17931;
assign x_17933 = x_17930 & x_17932;
assign x_17934 = x_17928 & x_17933;
assign x_17935 = x_6690 & x_6691;
assign x_17936 = x_6693 & x_6694;
assign x_17937 = x_6692 & x_17936;
assign x_17938 = x_17935 & x_17937;
assign x_17939 = x_6696 & x_6697;
assign x_17940 = x_6695 & x_17939;
assign x_17941 = x_6699 & x_6700;
assign x_17942 = x_6698 & x_17941;
assign x_17943 = x_17940 & x_17942;
assign x_17944 = x_17938 & x_17943;
assign x_17945 = x_17934 & x_17944;
assign x_17946 = x_6701 & x_6702;
assign x_17947 = x_6704 & x_6705;
assign x_17948 = x_6703 & x_17947;
assign x_17949 = x_17946 & x_17948;
assign x_17950 = x_6707 & x_6708;
assign x_17951 = x_6706 & x_17950;
assign x_17952 = x_6710 & x_6711;
assign x_17953 = x_6709 & x_17952;
assign x_17954 = x_17951 & x_17953;
assign x_17955 = x_17949 & x_17954;
assign x_17956 = x_6712 & x_6713;
assign x_17957 = x_6715 & x_6716;
assign x_17958 = x_6714 & x_17957;
assign x_17959 = x_17956 & x_17958;
assign x_17960 = x_6718 & x_6719;
assign x_17961 = x_6717 & x_17960;
assign x_17962 = x_6721 & x_6722;
assign x_17963 = x_6720 & x_17962;
assign x_17964 = x_17961 & x_17963;
assign x_17965 = x_17959 & x_17964;
assign x_17966 = x_17955 & x_17965;
assign x_17967 = x_17945 & x_17966;
assign x_17968 = x_6723 & x_6724;
assign x_17969 = x_6726 & x_6727;
assign x_17970 = x_6725 & x_17969;
assign x_17971 = x_17968 & x_17970;
assign x_17972 = x_6729 & x_6730;
assign x_17973 = x_6728 & x_17972;
assign x_17974 = x_6732 & x_6733;
assign x_17975 = x_6731 & x_17974;
assign x_17976 = x_17973 & x_17975;
assign x_17977 = x_17971 & x_17976;
assign x_17978 = x_6734 & x_6735;
assign x_17979 = x_6737 & x_6738;
assign x_17980 = x_6736 & x_17979;
assign x_17981 = x_17978 & x_17980;
assign x_17982 = x_6740 & x_6741;
assign x_17983 = x_6739 & x_17982;
assign x_17984 = x_6743 & x_6744;
assign x_17985 = x_6742 & x_17984;
assign x_17986 = x_17983 & x_17985;
assign x_17987 = x_17981 & x_17986;
assign x_17988 = x_17977 & x_17987;
assign x_17989 = x_6745 & x_6746;
assign x_17990 = x_6748 & x_6749;
assign x_17991 = x_6747 & x_17990;
assign x_17992 = x_17989 & x_17991;
assign x_17993 = x_6751 & x_6752;
assign x_17994 = x_6750 & x_17993;
assign x_17995 = x_6754 & x_6755;
assign x_17996 = x_6753 & x_17995;
assign x_17997 = x_17994 & x_17996;
assign x_17998 = x_17992 & x_17997;
assign x_17999 = x_6756 & x_6757;
assign x_18000 = x_6759 & x_6760;
assign x_18001 = x_6758 & x_18000;
assign x_18002 = x_17999 & x_18001;
assign x_18003 = x_6762 & x_6763;
assign x_18004 = x_6761 & x_18003;
assign x_18005 = x_6765 & x_6766;
assign x_18006 = x_6764 & x_18005;
assign x_18007 = x_18004 & x_18006;
assign x_18008 = x_18002 & x_18007;
assign x_18009 = x_17998 & x_18008;
assign x_18010 = x_17988 & x_18009;
assign x_18011 = x_17967 & x_18010;
assign x_18012 = x_6767 & x_6768;
assign x_18013 = x_6770 & x_6771;
assign x_18014 = x_6769 & x_18013;
assign x_18015 = x_18012 & x_18014;
assign x_18016 = x_6773 & x_6774;
assign x_18017 = x_6772 & x_18016;
assign x_18018 = x_6776 & x_6777;
assign x_18019 = x_6775 & x_18018;
assign x_18020 = x_18017 & x_18019;
assign x_18021 = x_18015 & x_18020;
assign x_18022 = x_6778 & x_6779;
assign x_18023 = x_6781 & x_6782;
assign x_18024 = x_6780 & x_18023;
assign x_18025 = x_18022 & x_18024;
assign x_18026 = x_6784 & x_6785;
assign x_18027 = x_6783 & x_18026;
assign x_18028 = x_6787 & x_6788;
assign x_18029 = x_6786 & x_18028;
assign x_18030 = x_18027 & x_18029;
assign x_18031 = x_18025 & x_18030;
assign x_18032 = x_18021 & x_18031;
assign x_18033 = x_6789 & x_6790;
assign x_18034 = x_6792 & x_6793;
assign x_18035 = x_6791 & x_18034;
assign x_18036 = x_18033 & x_18035;
assign x_18037 = x_6795 & x_6796;
assign x_18038 = x_6794 & x_18037;
assign x_18039 = x_6798 & x_6799;
assign x_18040 = x_6797 & x_18039;
assign x_18041 = x_18038 & x_18040;
assign x_18042 = x_18036 & x_18041;
assign x_18043 = x_6800 & x_6801;
assign x_18044 = x_6803 & x_6804;
assign x_18045 = x_6802 & x_18044;
assign x_18046 = x_18043 & x_18045;
assign x_18047 = x_6806 & x_6807;
assign x_18048 = x_6805 & x_18047;
assign x_18049 = x_6809 & x_6810;
assign x_18050 = x_6808 & x_18049;
assign x_18051 = x_18048 & x_18050;
assign x_18052 = x_18046 & x_18051;
assign x_18053 = x_18042 & x_18052;
assign x_18054 = x_18032 & x_18053;
assign x_18055 = x_6811 & x_6812;
assign x_18056 = x_6814 & x_6815;
assign x_18057 = x_6813 & x_18056;
assign x_18058 = x_18055 & x_18057;
assign x_18059 = x_6817 & x_6818;
assign x_18060 = x_6816 & x_18059;
assign x_18061 = x_6820 & x_6821;
assign x_18062 = x_6819 & x_18061;
assign x_18063 = x_18060 & x_18062;
assign x_18064 = x_18058 & x_18063;
assign x_18065 = x_6822 & x_6823;
assign x_18066 = x_6825 & x_6826;
assign x_18067 = x_6824 & x_18066;
assign x_18068 = x_18065 & x_18067;
assign x_18069 = x_6828 & x_6829;
assign x_18070 = x_6827 & x_18069;
assign x_18071 = x_6831 & x_6832;
assign x_18072 = x_6830 & x_18071;
assign x_18073 = x_18070 & x_18072;
assign x_18074 = x_18068 & x_18073;
assign x_18075 = x_18064 & x_18074;
assign x_18076 = x_6833 & x_6834;
assign x_18077 = x_6836 & x_6837;
assign x_18078 = x_6835 & x_18077;
assign x_18079 = x_18076 & x_18078;
assign x_18080 = x_6839 & x_6840;
assign x_18081 = x_6838 & x_18080;
assign x_18082 = x_6842 & x_6843;
assign x_18083 = x_6841 & x_18082;
assign x_18084 = x_18081 & x_18083;
assign x_18085 = x_18079 & x_18084;
assign x_18086 = x_6844 & x_6845;
assign x_18087 = x_6847 & x_6848;
assign x_18088 = x_6846 & x_18087;
assign x_18089 = x_18086 & x_18088;
assign x_18090 = x_6850 & x_6851;
assign x_18091 = x_6849 & x_18090;
assign x_18092 = x_6853 & x_6854;
assign x_18093 = x_6852 & x_18092;
assign x_18094 = x_18091 & x_18093;
assign x_18095 = x_18089 & x_18094;
assign x_18096 = x_18085 & x_18095;
assign x_18097 = x_18075 & x_18096;
assign x_18098 = x_18054 & x_18097;
assign x_18099 = x_18011 & x_18098;
assign x_18100 = x_6855 & x_6856;
assign x_18101 = x_6858 & x_6859;
assign x_18102 = x_6857 & x_18101;
assign x_18103 = x_18100 & x_18102;
assign x_18104 = x_6861 & x_6862;
assign x_18105 = x_6860 & x_18104;
assign x_18106 = x_6864 & x_6865;
assign x_18107 = x_6863 & x_18106;
assign x_18108 = x_18105 & x_18107;
assign x_18109 = x_18103 & x_18108;
assign x_18110 = x_6866 & x_6867;
assign x_18111 = x_6869 & x_6870;
assign x_18112 = x_6868 & x_18111;
assign x_18113 = x_18110 & x_18112;
assign x_18114 = x_6872 & x_6873;
assign x_18115 = x_6871 & x_18114;
assign x_18116 = x_6875 & x_6876;
assign x_18117 = x_6874 & x_18116;
assign x_18118 = x_18115 & x_18117;
assign x_18119 = x_18113 & x_18118;
assign x_18120 = x_18109 & x_18119;
assign x_18121 = x_6877 & x_6878;
assign x_18122 = x_6880 & x_6881;
assign x_18123 = x_6879 & x_18122;
assign x_18124 = x_18121 & x_18123;
assign x_18125 = x_6883 & x_6884;
assign x_18126 = x_6882 & x_18125;
assign x_18127 = x_6886 & x_6887;
assign x_18128 = x_6885 & x_18127;
assign x_18129 = x_18126 & x_18128;
assign x_18130 = x_18124 & x_18129;
assign x_18131 = x_6888 & x_6889;
assign x_18132 = x_6891 & x_6892;
assign x_18133 = x_6890 & x_18132;
assign x_18134 = x_18131 & x_18133;
assign x_18135 = x_6894 & x_6895;
assign x_18136 = x_6893 & x_18135;
assign x_18137 = x_6897 & x_6898;
assign x_18138 = x_6896 & x_18137;
assign x_18139 = x_18136 & x_18138;
assign x_18140 = x_18134 & x_18139;
assign x_18141 = x_18130 & x_18140;
assign x_18142 = x_18120 & x_18141;
assign x_18143 = x_6899 & x_6900;
assign x_18144 = x_6902 & x_6903;
assign x_18145 = x_6901 & x_18144;
assign x_18146 = x_18143 & x_18145;
assign x_18147 = x_6905 & x_6906;
assign x_18148 = x_6904 & x_18147;
assign x_18149 = x_6908 & x_6909;
assign x_18150 = x_6907 & x_18149;
assign x_18151 = x_18148 & x_18150;
assign x_18152 = x_18146 & x_18151;
assign x_18153 = x_6910 & x_6911;
assign x_18154 = x_6913 & x_6914;
assign x_18155 = x_6912 & x_18154;
assign x_18156 = x_18153 & x_18155;
assign x_18157 = x_6916 & x_6917;
assign x_18158 = x_6915 & x_18157;
assign x_18159 = x_6919 & x_6920;
assign x_18160 = x_6918 & x_18159;
assign x_18161 = x_18158 & x_18160;
assign x_18162 = x_18156 & x_18161;
assign x_18163 = x_18152 & x_18162;
assign x_18164 = x_6921 & x_6922;
assign x_18165 = x_6924 & x_6925;
assign x_18166 = x_6923 & x_18165;
assign x_18167 = x_18164 & x_18166;
assign x_18168 = x_6927 & x_6928;
assign x_18169 = x_6926 & x_18168;
assign x_18170 = x_6930 & x_6931;
assign x_18171 = x_6929 & x_18170;
assign x_18172 = x_18169 & x_18171;
assign x_18173 = x_18167 & x_18172;
assign x_18174 = x_6932 & x_6933;
assign x_18175 = x_6935 & x_6936;
assign x_18176 = x_6934 & x_18175;
assign x_18177 = x_18174 & x_18176;
assign x_18178 = x_6938 & x_6939;
assign x_18179 = x_6937 & x_18178;
assign x_18180 = x_6941 & x_6942;
assign x_18181 = x_6940 & x_18180;
assign x_18182 = x_18179 & x_18181;
assign x_18183 = x_18177 & x_18182;
assign x_18184 = x_18173 & x_18183;
assign x_18185 = x_18163 & x_18184;
assign x_18186 = x_18142 & x_18185;
assign x_18187 = x_6943 & x_6944;
assign x_18188 = x_6946 & x_6947;
assign x_18189 = x_6945 & x_18188;
assign x_18190 = x_18187 & x_18189;
assign x_18191 = x_6949 & x_6950;
assign x_18192 = x_6948 & x_18191;
assign x_18193 = x_6952 & x_6953;
assign x_18194 = x_6951 & x_18193;
assign x_18195 = x_18192 & x_18194;
assign x_18196 = x_18190 & x_18195;
assign x_18197 = x_6954 & x_6955;
assign x_18198 = x_6957 & x_6958;
assign x_18199 = x_6956 & x_18198;
assign x_18200 = x_18197 & x_18199;
assign x_18201 = x_6960 & x_6961;
assign x_18202 = x_6959 & x_18201;
assign x_18203 = x_6963 & x_6964;
assign x_18204 = x_6962 & x_18203;
assign x_18205 = x_18202 & x_18204;
assign x_18206 = x_18200 & x_18205;
assign x_18207 = x_18196 & x_18206;
assign x_18208 = x_6965 & x_6966;
assign x_18209 = x_6968 & x_6969;
assign x_18210 = x_6967 & x_18209;
assign x_18211 = x_18208 & x_18210;
assign x_18212 = x_6971 & x_6972;
assign x_18213 = x_6970 & x_18212;
assign x_18214 = x_6974 & x_6975;
assign x_18215 = x_6973 & x_18214;
assign x_18216 = x_18213 & x_18215;
assign x_18217 = x_18211 & x_18216;
assign x_18218 = x_6976 & x_6977;
assign x_18219 = x_6979 & x_6980;
assign x_18220 = x_6978 & x_18219;
assign x_18221 = x_18218 & x_18220;
assign x_18222 = x_6982 & x_6983;
assign x_18223 = x_6981 & x_18222;
assign x_18224 = x_6985 & x_6986;
assign x_18225 = x_6984 & x_18224;
assign x_18226 = x_18223 & x_18225;
assign x_18227 = x_18221 & x_18226;
assign x_18228 = x_18217 & x_18227;
assign x_18229 = x_18207 & x_18228;
assign x_18230 = x_6987 & x_6988;
assign x_18231 = x_6990 & x_6991;
assign x_18232 = x_6989 & x_18231;
assign x_18233 = x_18230 & x_18232;
assign x_18234 = x_6993 & x_6994;
assign x_18235 = x_6992 & x_18234;
assign x_18236 = x_6996 & x_6997;
assign x_18237 = x_6995 & x_18236;
assign x_18238 = x_18235 & x_18237;
assign x_18239 = x_18233 & x_18238;
assign x_18240 = x_6998 & x_6999;
assign x_18241 = x_7001 & x_7002;
assign x_18242 = x_7000 & x_18241;
assign x_18243 = x_18240 & x_18242;
assign x_18244 = x_7004 & x_7005;
assign x_18245 = x_7003 & x_18244;
assign x_18246 = x_7007 & x_7008;
assign x_18247 = x_7006 & x_18246;
assign x_18248 = x_18245 & x_18247;
assign x_18249 = x_18243 & x_18248;
assign x_18250 = x_18239 & x_18249;
assign x_18251 = x_7009 & x_7010;
assign x_18252 = x_7012 & x_7013;
assign x_18253 = x_7011 & x_18252;
assign x_18254 = x_18251 & x_18253;
assign x_18255 = x_7015 & x_7016;
assign x_18256 = x_7014 & x_18255;
assign x_18257 = x_7018 & x_7019;
assign x_18258 = x_7017 & x_18257;
assign x_18259 = x_18256 & x_18258;
assign x_18260 = x_18254 & x_18259;
assign x_18261 = x_7020 & x_7021;
assign x_18262 = x_7023 & x_7024;
assign x_18263 = x_7022 & x_18262;
assign x_18264 = x_18261 & x_18263;
assign x_18265 = x_7026 & x_7027;
assign x_18266 = x_7025 & x_18265;
assign x_18267 = x_7029 & x_7030;
assign x_18268 = x_7028 & x_18267;
assign x_18269 = x_18266 & x_18268;
assign x_18270 = x_18264 & x_18269;
assign x_18271 = x_18260 & x_18270;
assign x_18272 = x_18250 & x_18271;
assign x_18273 = x_18229 & x_18272;
assign x_18274 = x_18186 & x_18273;
assign x_18275 = x_18099 & x_18274;
assign x_18276 = x_17924 & x_18275;
assign x_18277 = x_17574 & x_18276;
assign x_18278 = x_7031 & x_7032;
assign x_18279 = x_7034 & x_7035;
assign x_18280 = x_7033 & x_18279;
assign x_18281 = x_18278 & x_18280;
assign x_18282 = x_7036 & x_7037;
assign x_18283 = x_7039 & x_7040;
assign x_18284 = x_7038 & x_18283;
assign x_18285 = x_18282 & x_18284;
assign x_18286 = x_18281 & x_18285;
assign x_18287 = x_7041 & x_7042;
assign x_18288 = x_7044 & x_7045;
assign x_18289 = x_7043 & x_18288;
assign x_18290 = x_18287 & x_18289;
assign x_18291 = x_7047 & x_7048;
assign x_18292 = x_7046 & x_18291;
assign x_18293 = x_7050 & x_7051;
assign x_18294 = x_7049 & x_18293;
assign x_18295 = x_18292 & x_18294;
assign x_18296 = x_18290 & x_18295;
assign x_18297 = x_18286 & x_18296;
assign x_18298 = x_7052 & x_7053;
assign x_18299 = x_7055 & x_7056;
assign x_18300 = x_7054 & x_18299;
assign x_18301 = x_18298 & x_18300;
assign x_18302 = x_7058 & x_7059;
assign x_18303 = x_7057 & x_18302;
assign x_18304 = x_7061 & x_7062;
assign x_18305 = x_7060 & x_18304;
assign x_18306 = x_18303 & x_18305;
assign x_18307 = x_18301 & x_18306;
assign x_18308 = x_7063 & x_7064;
assign x_18309 = x_7066 & x_7067;
assign x_18310 = x_7065 & x_18309;
assign x_18311 = x_18308 & x_18310;
assign x_18312 = x_7069 & x_7070;
assign x_18313 = x_7068 & x_18312;
assign x_18314 = x_7072 & x_7073;
assign x_18315 = x_7071 & x_18314;
assign x_18316 = x_18313 & x_18315;
assign x_18317 = x_18311 & x_18316;
assign x_18318 = x_18307 & x_18317;
assign x_18319 = x_18297 & x_18318;
assign x_18320 = x_7074 & x_7075;
assign x_18321 = x_7077 & x_7078;
assign x_18322 = x_7076 & x_18321;
assign x_18323 = x_18320 & x_18322;
assign x_18324 = x_7080 & x_7081;
assign x_18325 = x_7079 & x_18324;
assign x_18326 = x_7083 & x_7084;
assign x_18327 = x_7082 & x_18326;
assign x_18328 = x_18325 & x_18327;
assign x_18329 = x_18323 & x_18328;
assign x_18330 = x_7085 & x_7086;
assign x_18331 = x_7088 & x_7089;
assign x_18332 = x_7087 & x_18331;
assign x_18333 = x_18330 & x_18332;
assign x_18334 = x_7091 & x_7092;
assign x_18335 = x_7090 & x_18334;
assign x_18336 = x_7094 & x_7095;
assign x_18337 = x_7093 & x_18336;
assign x_18338 = x_18335 & x_18337;
assign x_18339 = x_18333 & x_18338;
assign x_18340 = x_18329 & x_18339;
assign x_18341 = x_7096 & x_7097;
assign x_18342 = x_7099 & x_7100;
assign x_18343 = x_7098 & x_18342;
assign x_18344 = x_18341 & x_18343;
assign x_18345 = x_7102 & x_7103;
assign x_18346 = x_7101 & x_18345;
assign x_18347 = x_7105 & x_7106;
assign x_18348 = x_7104 & x_18347;
assign x_18349 = x_18346 & x_18348;
assign x_18350 = x_18344 & x_18349;
assign x_18351 = x_7107 & x_7108;
assign x_18352 = x_7110 & x_7111;
assign x_18353 = x_7109 & x_18352;
assign x_18354 = x_18351 & x_18353;
assign x_18355 = x_7113 & x_7114;
assign x_18356 = x_7112 & x_18355;
assign x_18357 = x_7116 & x_7117;
assign x_18358 = x_7115 & x_18357;
assign x_18359 = x_18356 & x_18358;
assign x_18360 = x_18354 & x_18359;
assign x_18361 = x_18350 & x_18360;
assign x_18362 = x_18340 & x_18361;
assign x_18363 = x_18319 & x_18362;
assign x_18364 = x_7118 & x_7119;
assign x_18365 = x_7121 & x_7122;
assign x_18366 = x_7120 & x_18365;
assign x_18367 = x_18364 & x_18366;
assign x_18368 = x_7124 & x_7125;
assign x_18369 = x_7123 & x_18368;
assign x_18370 = x_7127 & x_7128;
assign x_18371 = x_7126 & x_18370;
assign x_18372 = x_18369 & x_18371;
assign x_18373 = x_18367 & x_18372;
assign x_18374 = x_7129 & x_7130;
assign x_18375 = x_7132 & x_7133;
assign x_18376 = x_7131 & x_18375;
assign x_18377 = x_18374 & x_18376;
assign x_18378 = x_7135 & x_7136;
assign x_18379 = x_7134 & x_18378;
assign x_18380 = x_7138 & x_7139;
assign x_18381 = x_7137 & x_18380;
assign x_18382 = x_18379 & x_18381;
assign x_18383 = x_18377 & x_18382;
assign x_18384 = x_18373 & x_18383;
assign x_18385 = x_7140 & x_7141;
assign x_18386 = x_7143 & x_7144;
assign x_18387 = x_7142 & x_18386;
assign x_18388 = x_18385 & x_18387;
assign x_18389 = x_7146 & x_7147;
assign x_18390 = x_7145 & x_18389;
assign x_18391 = x_7149 & x_7150;
assign x_18392 = x_7148 & x_18391;
assign x_18393 = x_18390 & x_18392;
assign x_18394 = x_18388 & x_18393;
assign x_18395 = x_7151 & x_7152;
assign x_18396 = x_7154 & x_7155;
assign x_18397 = x_7153 & x_18396;
assign x_18398 = x_18395 & x_18397;
assign x_18399 = x_7157 & x_7158;
assign x_18400 = x_7156 & x_18399;
assign x_18401 = x_7160 & x_7161;
assign x_18402 = x_7159 & x_18401;
assign x_18403 = x_18400 & x_18402;
assign x_18404 = x_18398 & x_18403;
assign x_18405 = x_18394 & x_18404;
assign x_18406 = x_18384 & x_18405;
assign x_18407 = x_7162 & x_7163;
assign x_18408 = x_7165 & x_7166;
assign x_18409 = x_7164 & x_18408;
assign x_18410 = x_18407 & x_18409;
assign x_18411 = x_7168 & x_7169;
assign x_18412 = x_7167 & x_18411;
assign x_18413 = x_7171 & x_7172;
assign x_18414 = x_7170 & x_18413;
assign x_18415 = x_18412 & x_18414;
assign x_18416 = x_18410 & x_18415;
assign x_18417 = x_7173 & x_7174;
assign x_18418 = x_7176 & x_7177;
assign x_18419 = x_7175 & x_18418;
assign x_18420 = x_18417 & x_18419;
assign x_18421 = x_7179 & x_7180;
assign x_18422 = x_7178 & x_18421;
assign x_18423 = x_7182 & x_7183;
assign x_18424 = x_7181 & x_18423;
assign x_18425 = x_18422 & x_18424;
assign x_18426 = x_18420 & x_18425;
assign x_18427 = x_18416 & x_18426;
assign x_18428 = x_7184 & x_7185;
assign x_18429 = x_7187 & x_7188;
assign x_18430 = x_7186 & x_18429;
assign x_18431 = x_18428 & x_18430;
assign x_18432 = x_7190 & x_7191;
assign x_18433 = x_7189 & x_18432;
assign x_18434 = x_7193 & x_7194;
assign x_18435 = x_7192 & x_18434;
assign x_18436 = x_18433 & x_18435;
assign x_18437 = x_18431 & x_18436;
assign x_18438 = x_7195 & x_7196;
assign x_18439 = x_7198 & x_7199;
assign x_18440 = x_7197 & x_18439;
assign x_18441 = x_18438 & x_18440;
assign x_18442 = x_7201 & x_7202;
assign x_18443 = x_7200 & x_18442;
assign x_18444 = x_7204 & x_7205;
assign x_18445 = x_7203 & x_18444;
assign x_18446 = x_18443 & x_18445;
assign x_18447 = x_18441 & x_18446;
assign x_18448 = x_18437 & x_18447;
assign x_18449 = x_18427 & x_18448;
assign x_18450 = x_18406 & x_18449;
assign x_18451 = x_18363 & x_18450;
assign x_18452 = x_7206 & x_7207;
assign x_18453 = x_7209 & x_7210;
assign x_18454 = x_7208 & x_18453;
assign x_18455 = x_18452 & x_18454;
assign x_18456 = x_7212 & x_7213;
assign x_18457 = x_7211 & x_18456;
assign x_18458 = x_7215 & x_7216;
assign x_18459 = x_7214 & x_18458;
assign x_18460 = x_18457 & x_18459;
assign x_18461 = x_18455 & x_18460;
assign x_18462 = x_7217 & x_7218;
assign x_18463 = x_7220 & x_7221;
assign x_18464 = x_7219 & x_18463;
assign x_18465 = x_18462 & x_18464;
assign x_18466 = x_7223 & x_7224;
assign x_18467 = x_7222 & x_18466;
assign x_18468 = x_7226 & x_7227;
assign x_18469 = x_7225 & x_18468;
assign x_18470 = x_18467 & x_18469;
assign x_18471 = x_18465 & x_18470;
assign x_18472 = x_18461 & x_18471;
assign x_18473 = x_7228 & x_7229;
assign x_18474 = x_7231 & x_7232;
assign x_18475 = x_7230 & x_18474;
assign x_18476 = x_18473 & x_18475;
assign x_18477 = x_7234 & x_7235;
assign x_18478 = x_7233 & x_18477;
assign x_18479 = x_7237 & x_7238;
assign x_18480 = x_7236 & x_18479;
assign x_18481 = x_18478 & x_18480;
assign x_18482 = x_18476 & x_18481;
assign x_18483 = x_7239 & x_7240;
assign x_18484 = x_7242 & x_7243;
assign x_18485 = x_7241 & x_18484;
assign x_18486 = x_18483 & x_18485;
assign x_18487 = x_7245 & x_7246;
assign x_18488 = x_7244 & x_18487;
assign x_18489 = x_7248 & x_7249;
assign x_18490 = x_7247 & x_18489;
assign x_18491 = x_18488 & x_18490;
assign x_18492 = x_18486 & x_18491;
assign x_18493 = x_18482 & x_18492;
assign x_18494 = x_18472 & x_18493;
assign x_18495 = x_7250 & x_7251;
assign x_18496 = x_7253 & x_7254;
assign x_18497 = x_7252 & x_18496;
assign x_18498 = x_18495 & x_18497;
assign x_18499 = x_7256 & x_7257;
assign x_18500 = x_7255 & x_18499;
assign x_18501 = x_7259 & x_7260;
assign x_18502 = x_7258 & x_18501;
assign x_18503 = x_18500 & x_18502;
assign x_18504 = x_18498 & x_18503;
assign x_18505 = x_7261 & x_7262;
assign x_18506 = x_7264 & x_7265;
assign x_18507 = x_7263 & x_18506;
assign x_18508 = x_18505 & x_18507;
assign x_18509 = x_7267 & x_7268;
assign x_18510 = x_7266 & x_18509;
assign x_18511 = x_7270 & x_7271;
assign x_18512 = x_7269 & x_18511;
assign x_18513 = x_18510 & x_18512;
assign x_18514 = x_18508 & x_18513;
assign x_18515 = x_18504 & x_18514;
assign x_18516 = x_7272 & x_7273;
assign x_18517 = x_7275 & x_7276;
assign x_18518 = x_7274 & x_18517;
assign x_18519 = x_18516 & x_18518;
assign x_18520 = x_7278 & x_7279;
assign x_18521 = x_7277 & x_18520;
assign x_18522 = x_7281 & x_7282;
assign x_18523 = x_7280 & x_18522;
assign x_18524 = x_18521 & x_18523;
assign x_18525 = x_18519 & x_18524;
assign x_18526 = x_7283 & x_7284;
assign x_18527 = x_7286 & x_7287;
assign x_18528 = x_7285 & x_18527;
assign x_18529 = x_18526 & x_18528;
assign x_18530 = x_7289 & x_7290;
assign x_18531 = x_7288 & x_18530;
assign x_18532 = x_7292 & x_7293;
assign x_18533 = x_7291 & x_18532;
assign x_18534 = x_18531 & x_18533;
assign x_18535 = x_18529 & x_18534;
assign x_18536 = x_18525 & x_18535;
assign x_18537 = x_18515 & x_18536;
assign x_18538 = x_18494 & x_18537;
assign x_18539 = x_7294 & x_7295;
assign x_18540 = x_7297 & x_7298;
assign x_18541 = x_7296 & x_18540;
assign x_18542 = x_18539 & x_18541;
assign x_18543 = x_7300 & x_7301;
assign x_18544 = x_7299 & x_18543;
assign x_18545 = x_7303 & x_7304;
assign x_18546 = x_7302 & x_18545;
assign x_18547 = x_18544 & x_18546;
assign x_18548 = x_18542 & x_18547;
assign x_18549 = x_7305 & x_7306;
assign x_18550 = x_7308 & x_7309;
assign x_18551 = x_7307 & x_18550;
assign x_18552 = x_18549 & x_18551;
assign x_18553 = x_7311 & x_7312;
assign x_18554 = x_7310 & x_18553;
assign x_18555 = x_7314 & x_7315;
assign x_18556 = x_7313 & x_18555;
assign x_18557 = x_18554 & x_18556;
assign x_18558 = x_18552 & x_18557;
assign x_18559 = x_18548 & x_18558;
assign x_18560 = x_7316 & x_7317;
assign x_18561 = x_7319 & x_7320;
assign x_18562 = x_7318 & x_18561;
assign x_18563 = x_18560 & x_18562;
assign x_18564 = x_7322 & x_7323;
assign x_18565 = x_7321 & x_18564;
assign x_18566 = x_7325 & x_7326;
assign x_18567 = x_7324 & x_18566;
assign x_18568 = x_18565 & x_18567;
assign x_18569 = x_18563 & x_18568;
assign x_18570 = x_7327 & x_7328;
assign x_18571 = x_7330 & x_7331;
assign x_18572 = x_7329 & x_18571;
assign x_18573 = x_18570 & x_18572;
assign x_18574 = x_7333 & x_7334;
assign x_18575 = x_7332 & x_18574;
assign x_18576 = x_7336 & x_7337;
assign x_18577 = x_7335 & x_18576;
assign x_18578 = x_18575 & x_18577;
assign x_18579 = x_18573 & x_18578;
assign x_18580 = x_18569 & x_18579;
assign x_18581 = x_18559 & x_18580;
assign x_18582 = x_7338 & x_7339;
assign x_18583 = x_7341 & x_7342;
assign x_18584 = x_7340 & x_18583;
assign x_18585 = x_18582 & x_18584;
assign x_18586 = x_7344 & x_7345;
assign x_18587 = x_7343 & x_18586;
assign x_18588 = x_7347 & x_7348;
assign x_18589 = x_7346 & x_18588;
assign x_18590 = x_18587 & x_18589;
assign x_18591 = x_18585 & x_18590;
assign x_18592 = x_7349 & x_7350;
assign x_18593 = x_7352 & x_7353;
assign x_18594 = x_7351 & x_18593;
assign x_18595 = x_18592 & x_18594;
assign x_18596 = x_7355 & x_7356;
assign x_18597 = x_7354 & x_18596;
assign x_18598 = x_7358 & x_7359;
assign x_18599 = x_7357 & x_18598;
assign x_18600 = x_18597 & x_18599;
assign x_18601 = x_18595 & x_18600;
assign x_18602 = x_18591 & x_18601;
assign x_18603 = x_7360 & x_7361;
assign x_18604 = x_7363 & x_7364;
assign x_18605 = x_7362 & x_18604;
assign x_18606 = x_18603 & x_18605;
assign x_18607 = x_7366 & x_7367;
assign x_18608 = x_7365 & x_18607;
assign x_18609 = x_7369 & x_7370;
assign x_18610 = x_7368 & x_18609;
assign x_18611 = x_18608 & x_18610;
assign x_18612 = x_18606 & x_18611;
assign x_18613 = x_7371 & x_7372;
assign x_18614 = x_7374 & x_7375;
assign x_18615 = x_7373 & x_18614;
assign x_18616 = x_18613 & x_18615;
assign x_18617 = x_7377 & x_7378;
assign x_18618 = x_7376 & x_18617;
assign x_18619 = x_7380 & x_7381;
assign x_18620 = x_7379 & x_18619;
assign x_18621 = x_18618 & x_18620;
assign x_18622 = x_18616 & x_18621;
assign x_18623 = x_18612 & x_18622;
assign x_18624 = x_18602 & x_18623;
assign x_18625 = x_18581 & x_18624;
assign x_18626 = x_18538 & x_18625;
assign x_18627 = x_18451 & x_18626;
assign x_18628 = x_7382 & x_7383;
assign x_18629 = x_7385 & x_7386;
assign x_18630 = x_7384 & x_18629;
assign x_18631 = x_18628 & x_18630;
assign x_18632 = x_7388 & x_7389;
assign x_18633 = x_7387 & x_18632;
assign x_18634 = x_7391 & x_7392;
assign x_18635 = x_7390 & x_18634;
assign x_18636 = x_18633 & x_18635;
assign x_18637 = x_18631 & x_18636;
assign x_18638 = x_7393 & x_7394;
assign x_18639 = x_7396 & x_7397;
assign x_18640 = x_7395 & x_18639;
assign x_18641 = x_18638 & x_18640;
assign x_18642 = x_7399 & x_7400;
assign x_18643 = x_7398 & x_18642;
assign x_18644 = x_7402 & x_7403;
assign x_18645 = x_7401 & x_18644;
assign x_18646 = x_18643 & x_18645;
assign x_18647 = x_18641 & x_18646;
assign x_18648 = x_18637 & x_18647;
assign x_18649 = x_7404 & x_7405;
assign x_18650 = x_7407 & x_7408;
assign x_18651 = x_7406 & x_18650;
assign x_18652 = x_18649 & x_18651;
assign x_18653 = x_7410 & x_7411;
assign x_18654 = x_7409 & x_18653;
assign x_18655 = x_7413 & x_7414;
assign x_18656 = x_7412 & x_18655;
assign x_18657 = x_18654 & x_18656;
assign x_18658 = x_18652 & x_18657;
assign x_18659 = x_7415 & x_7416;
assign x_18660 = x_7418 & x_7419;
assign x_18661 = x_7417 & x_18660;
assign x_18662 = x_18659 & x_18661;
assign x_18663 = x_7421 & x_7422;
assign x_18664 = x_7420 & x_18663;
assign x_18665 = x_7424 & x_7425;
assign x_18666 = x_7423 & x_18665;
assign x_18667 = x_18664 & x_18666;
assign x_18668 = x_18662 & x_18667;
assign x_18669 = x_18658 & x_18668;
assign x_18670 = x_18648 & x_18669;
assign x_18671 = x_7426 & x_7427;
assign x_18672 = x_7429 & x_7430;
assign x_18673 = x_7428 & x_18672;
assign x_18674 = x_18671 & x_18673;
assign x_18675 = x_7432 & x_7433;
assign x_18676 = x_7431 & x_18675;
assign x_18677 = x_7435 & x_7436;
assign x_18678 = x_7434 & x_18677;
assign x_18679 = x_18676 & x_18678;
assign x_18680 = x_18674 & x_18679;
assign x_18681 = x_7437 & x_7438;
assign x_18682 = x_7440 & x_7441;
assign x_18683 = x_7439 & x_18682;
assign x_18684 = x_18681 & x_18683;
assign x_18685 = x_7443 & x_7444;
assign x_18686 = x_7442 & x_18685;
assign x_18687 = x_7446 & x_7447;
assign x_18688 = x_7445 & x_18687;
assign x_18689 = x_18686 & x_18688;
assign x_18690 = x_18684 & x_18689;
assign x_18691 = x_18680 & x_18690;
assign x_18692 = x_7448 & x_7449;
assign x_18693 = x_7451 & x_7452;
assign x_18694 = x_7450 & x_18693;
assign x_18695 = x_18692 & x_18694;
assign x_18696 = x_7454 & x_7455;
assign x_18697 = x_7453 & x_18696;
assign x_18698 = x_7457 & x_7458;
assign x_18699 = x_7456 & x_18698;
assign x_18700 = x_18697 & x_18699;
assign x_18701 = x_18695 & x_18700;
assign x_18702 = x_7459 & x_7460;
assign x_18703 = x_7462 & x_7463;
assign x_18704 = x_7461 & x_18703;
assign x_18705 = x_18702 & x_18704;
assign x_18706 = x_7465 & x_7466;
assign x_18707 = x_7464 & x_18706;
assign x_18708 = x_7468 & x_7469;
assign x_18709 = x_7467 & x_18708;
assign x_18710 = x_18707 & x_18709;
assign x_18711 = x_18705 & x_18710;
assign x_18712 = x_18701 & x_18711;
assign x_18713 = x_18691 & x_18712;
assign x_18714 = x_18670 & x_18713;
assign x_18715 = x_7470 & x_7471;
assign x_18716 = x_7473 & x_7474;
assign x_18717 = x_7472 & x_18716;
assign x_18718 = x_18715 & x_18717;
assign x_18719 = x_7476 & x_7477;
assign x_18720 = x_7475 & x_18719;
assign x_18721 = x_7479 & x_7480;
assign x_18722 = x_7478 & x_18721;
assign x_18723 = x_18720 & x_18722;
assign x_18724 = x_18718 & x_18723;
assign x_18725 = x_7481 & x_7482;
assign x_18726 = x_7484 & x_7485;
assign x_18727 = x_7483 & x_18726;
assign x_18728 = x_18725 & x_18727;
assign x_18729 = x_7487 & x_7488;
assign x_18730 = x_7486 & x_18729;
assign x_18731 = x_7490 & x_7491;
assign x_18732 = x_7489 & x_18731;
assign x_18733 = x_18730 & x_18732;
assign x_18734 = x_18728 & x_18733;
assign x_18735 = x_18724 & x_18734;
assign x_18736 = x_7492 & x_7493;
assign x_18737 = x_7495 & x_7496;
assign x_18738 = x_7494 & x_18737;
assign x_18739 = x_18736 & x_18738;
assign x_18740 = x_7498 & x_7499;
assign x_18741 = x_7497 & x_18740;
assign x_18742 = x_7501 & x_7502;
assign x_18743 = x_7500 & x_18742;
assign x_18744 = x_18741 & x_18743;
assign x_18745 = x_18739 & x_18744;
assign x_18746 = x_7503 & x_7504;
assign x_18747 = x_7506 & x_7507;
assign x_18748 = x_7505 & x_18747;
assign x_18749 = x_18746 & x_18748;
assign x_18750 = x_7509 & x_7510;
assign x_18751 = x_7508 & x_18750;
assign x_18752 = x_7512 & x_7513;
assign x_18753 = x_7511 & x_18752;
assign x_18754 = x_18751 & x_18753;
assign x_18755 = x_18749 & x_18754;
assign x_18756 = x_18745 & x_18755;
assign x_18757 = x_18735 & x_18756;
assign x_18758 = x_7514 & x_7515;
assign x_18759 = x_7517 & x_7518;
assign x_18760 = x_7516 & x_18759;
assign x_18761 = x_18758 & x_18760;
assign x_18762 = x_7520 & x_7521;
assign x_18763 = x_7519 & x_18762;
assign x_18764 = x_7523 & x_7524;
assign x_18765 = x_7522 & x_18764;
assign x_18766 = x_18763 & x_18765;
assign x_18767 = x_18761 & x_18766;
assign x_18768 = x_7525 & x_7526;
assign x_18769 = x_7528 & x_7529;
assign x_18770 = x_7527 & x_18769;
assign x_18771 = x_18768 & x_18770;
assign x_18772 = x_7531 & x_7532;
assign x_18773 = x_7530 & x_18772;
assign x_18774 = x_7534 & x_7535;
assign x_18775 = x_7533 & x_18774;
assign x_18776 = x_18773 & x_18775;
assign x_18777 = x_18771 & x_18776;
assign x_18778 = x_18767 & x_18777;
assign x_18779 = x_7536 & x_7537;
assign x_18780 = x_7539 & x_7540;
assign x_18781 = x_7538 & x_18780;
assign x_18782 = x_18779 & x_18781;
assign x_18783 = x_7542 & x_7543;
assign x_18784 = x_7541 & x_18783;
assign x_18785 = x_7545 & x_7546;
assign x_18786 = x_7544 & x_18785;
assign x_18787 = x_18784 & x_18786;
assign x_18788 = x_18782 & x_18787;
assign x_18789 = x_7547 & x_7548;
assign x_18790 = x_7550 & x_7551;
assign x_18791 = x_7549 & x_18790;
assign x_18792 = x_18789 & x_18791;
assign x_18793 = x_7553 & x_7554;
assign x_18794 = x_7552 & x_18793;
assign x_18795 = x_7556 & x_7557;
assign x_18796 = x_7555 & x_18795;
assign x_18797 = x_18794 & x_18796;
assign x_18798 = x_18792 & x_18797;
assign x_18799 = x_18788 & x_18798;
assign x_18800 = x_18778 & x_18799;
assign x_18801 = x_18757 & x_18800;
assign x_18802 = x_18714 & x_18801;
assign x_18803 = x_7558 & x_7559;
assign x_18804 = x_7561 & x_7562;
assign x_18805 = x_7560 & x_18804;
assign x_18806 = x_18803 & x_18805;
assign x_18807 = x_7564 & x_7565;
assign x_18808 = x_7563 & x_18807;
assign x_18809 = x_7567 & x_7568;
assign x_18810 = x_7566 & x_18809;
assign x_18811 = x_18808 & x_18810;
assign x_18812 = x_18806 & x_18811;
assign x_18813 = x_7569 & x_7570;
assign x_18814 = x_7572 & x_7573;
assign x_18815 = x_7571 & x_18814;
assign x_18816 = x_18813 & x_18815;
assign x_18817 = x_7575 & x_7576;
assign x_18818 = x_7574 & x_18817;
assign x_18819 = x_7578 & x_7579;
assign x_18820 = x_7577 & x_18819;
assign x_18821 = x_18818 & x_18820;
assign x_18822 = x_18816 & x_18821;
assign x_18823 = x_18812 & x_18822;
assign x_18824 = x_7580 & x_7581;
assign x_18825 = x_7583 & x_7584;
assign x_18826 = x_7582 & x_18825;
assign x_18827 = x_18824 & x_18826;
assign x_18828 = x_7586 & x_7587;
assign x_18829 = x_7585 & x_18828;
assign x_18830 = x_7589 & x_7590;
assign x_18831 = x_7588 & x_18830;
assign x_18832 = x_18829 & x_18831;
assign x_18833 = x_18827 & x_18832;
assign x_18834 = x_7591 & x_7592;
assign x_18835 = x_7594 & x_7595;
assign x_18836 = x_7593 & x_18835;
assign x_18837 = x_18834 & x_18836;
assign x_18838 = x_7597 & x_7598;
assign x_18839 = x_7596 & x_18838;
assign x_18840 = x_7600 & x_7601;
assign x_18841 = x_7599 & x_18840;
assign x_18842 = x_18839 & x_18841;
assign x_18843 = x_18837 & x_18842;
assign x_18844 = x_18833 & x_18843;
assign x_18845 = x_18823 & x_18844;
assign x_18846 = x_7602 & x_7603;
assign x_18847 = x_7605 & x_7606;
assign x_18848 = x_7604 & x_18847;
assign x_18849 = x_18846 & x_18848;
assign x_18850 = x_7608 & x_7609;
assign x_18851 = x_7607 & x_18850;
assign x_18852 = x_7611 & x_7612;
assign x_18853 = x_7610 & x_18852;
assign x_18854 = x_18851 & x_18853;
assign x_18855 = x_18849 & x_18854;
assign x_18856 = x_7613 & x_7614;
assign x_18857 = x_7616 & x_7617;
assign x_18858 = x_7615 & x_18857;
assign x_18859 = x_18856 & x_18858;
assign x_18860 = x_7619 & x_7620;
assign x_18861 = x_7618 & x_18860;
assign x_18862 = x_7622 & x_7623;
assign x_18863 = x_7621 & x_18862;
assign x_18864 = x_18861 & x_18863;
assign x_18865 = x_18859 & x_18864;
assign x_18866 = x_18855 & x_18865;
assign x_18867 = x_7624 & x_7625;
assign x_18868 = x_7627 & x_7628;
assign x_18869 = x_7626 & x_18868;
assign x_18870 = x_18867 & x_18869;
assign x_18871 = x_7630 & x_7631;
assign x_18872 = x_7629 & x_18871;
assign x_18873 = x_7633 & x_7634;
assign x_18874 = x_7632 & x_18873;
assign x_18875 = x_18872 & x_18874;
assign x_18876 = x_18870 & x_18875;
assign x_18877 = x_7635 & x_7636;
assign x_18878 = x_7638 & x_7639;
assign x_18879 = x_7637 & x_18878;
assign x_18880 = x_18877 & x_18879;
assign x_18881 = x_7641 & x_7642;
assign x_18882 = x_7640 & x_18881;
assign x_18883 = x_7644 & x_7645;
assign x_18884 = x_7643 & x_18883;
assign x_18885 = x_18882 & x_18884;
assign x_18886 = x_18880 & x_18885;
assign x_18887 = x_18876 & x_18886;
assign x_18888 = x_18866 & x_18887;
assign x_18889 = x_18845 & x_18888;
assign x_18890 = x_7646 & x_7647;
assign x_18891 = x_7649 & x_7650;
assign x_18892 = x_7648 & x_18891;
assign x_18893 = x_18890 & x_18892;
assign x_18894 = x_7652 & x_7653;
assign x_18895 = x_7651 & x_18894;
assign x_18896 = x_7655 & x_7656;
assign x_18897 = x_7654 & x_18896;
assign x_18898 = x_18895 & x_18897;
assign x_18899 = x_18893 & x_18898;
assign x_18900 = x_7657 & x_7658;
assign x_18901 = x_7660 & x_7661;
assign x_18902 = x_7659 & x_18901;
assign x_18903 = x_18900 & x_18902;
assign x_18904 = x_7663 & x_7664;
assign x_18905 = x_7662 & x_18904;
assign x_18906 = x_7666 & x_7667;
assign x_18907 = x_7665 & x_18906;
assign x_18908 = x_18905 & x_18907;
assign x_18909 = x_18903 & x_18908;
assign x_18910 = x_18899 & x_18909;
assign x_18911 = x_7668 & x_7669;
assign x_18912 = x_7671 & x_7672;
assign x_18913 = x_7670 & x_18912;
assign x_18914 = x_18911 & x_18913;
assign x_18915 = x_7674 & x_7675;
assign x_18916 = x_7673 & x_18915;
assign x_18917 = x_7677 & x_7678;
assign x_18918 = x_7676 & x_18917;
assign x_18919 = x_18916 & x_18918;
assign x_18920 = x_18914 & x_18919;
assign x_18921 = x_7679 & x_7680;
assign x_18922 = x_7682 & x_7683;
assign x_18923 = x_7681 & x_18922;
assign x_18924 = x_18921 & x_18923;
assign x_18925 = x_7685 & x_7686;
assign x_18926 = x_7684 & x_18925;
assign x_18927 = x_7688 & x_7689;
assign x_18928 = x_7687 & x_18927;
assign x_18929 = x_18926 & x_18928;
assign x_18930 = x_18924 & x_18929;
assign x_18931 = x_18920 & x_18930;
assign x_18932 = x_18910 & x_18931;
assign x_18933 = x_7690 & x_7691;
assign x_18934 = x_7693 & x_7694;
assign x_18935 = x_7692 & x_18934;
assign x_18936 = x_18933 & x_18935;
assign x_18937 = x_7696 & x_7697;
assign x_18938 = x_7695 & x_18937;
assign x_18939 = x_7699 & x_7700;
assign x_18940 = x_7698 & x_18939;
assign x_18941 = x_18938 & x_18940;
assign x_18942 = x_18936 & x_18941;
assign x_18943 = x_7701 & x_7702;
assign x_18944 = x_7704 & x_7705;
assign x_18945 = x_7703 & x_18944;
assign x_18946 = x_18943 & x_18945;
assign x_18947 = x_7707 & x_7708;
assign x_18948 = x_7706 & x_18947;
assign x_18949 = x_7710 & x_7711;
assign x_18950 = x_7709 & x_18949;
assign x_18951 = x_18948 & x_18950;
assign x_18952 = x_18946 & x_18951;
assign x_18953 = x_18942 & x_18952;
assign x_18954 = x_7712 & x_7713;
assign x_18955 = x_7715 & x_7716;
assign x_18956 = x_7714 & x_18955;
assign x_18957 = x_18954 & x_18956;
assign x_18958 = x_7718 & x_7719;
assign x_18959 = x_7717 & x_18958;
assign x_18960 = x_7721 & x_7722;
assign x_18961 = x_7720 & x_18960;
assign x_18962 = x_18959 & x_18961;
assign x_18963 = x_18957 & x_18962;
assign x_18964 = x_7723 & x_7724;
assign x_18965 = x_7726 & x_7727;
assign x_18966 = x_7725 & x_18965;
assign x_18967 = x_18964 & x_18966;
assign x_18968 = x_7729 & x_7730;
assign x_18969 = x_7728 & x_18968;
assign x_18970 = x_7732 & x_7733;
assign x_18971 = x_7731 & x_18970;
assign x_18972 = x_18969 & x_18971;
assign x_18973 = x_18967 & x_18972;
assign x_18974 = x_18963 & x_18973;
assign x_18975 = x_18953 & x_18974;
assign x_18976 = x_18932 & x_18975;
assign x_18977 = x_18889 & x_18976;
assign x_18978 = x_18802 & x_18977;
assign x_18979 = x_18627 & x_18978;
assign x_18980 = x_7734 & x_7735;
assign x_18981 = x_7737 & x_7738;
assign x_18982 = x_7736 & x_18981;
assign x_18983 = x_18980 & x_18982;
assign x_18984 = x_7739 & x_7740;
assign x_18985 = x_7742 & x_7743;
assign x_18986 = x_7741 & x_18985;
assign x_18987 = x_18984 & x_18986;
assign x_18988 = x_18983 & x_18987;
assign x_18989 = x_7744 & x_7745;
assign x_18990 = x_7747 & x_7748;
assign x_18991 = x_7746 & x_18990;
assign x_18992 = x_18989 & x_18991;
assign x_18993 = x_7750 & x_7751;
assign x_18994 = x_7749 & x_18993;
assign x_18995 = x_7753 & x_7754;
assign x_18996 = x_7752 & x_18995;
assign x_18997 = x_18994 & x_18996;
assign x_18998 = x_18992 & x_18997;
assign x_18999 = x_18988 & x_18998;
assign x_19000 = x_7755 & x_7756;
assign x_19001 = x_7758 & x_7759;
assign x_19002 = x_7757 & x_19001;
assign x_19003 = x_19000 & x_19002;
assign x_19004 = x_7761 & x_7762;
assign x_19005 = x_7760 & x_19004;
assign x_19006 = x_7764 & x_7765;
assign x_19007 = x_7763 & x_19006;
assign x_19008 = x_19005 & x_19007;
assign x_19009 = x_19003 & x_19008;
assign x_19010 = x_7766 & x_7767;
assign x_19011 = x_7769 & x_7770;
assign x_19012 = x_7768 & x_19011;
assign x_19013 = x_19010 & x_19012;
assign x_19014 = x_7772 & x_7773;
assign x_19015 = x_7771 & x_19014;
assign x_19016 = x_7775 & x_7776;
assign x_19017 = x_7774 & x_19016;
assign x_19018 = x_19015 & x_19017;
assign x_19019 = x_19013 & x_19018;
assign x_19020 = x_19009 & x_19019;
assign x_19021 = x_18999 & x_19020;
assign x_19022 = x_7777 & x_7778;
assign x_19023 = x_7780 & x_7781;
assign x_19024 = x_7779 & x_19023;
assign x_19025 = x_19022 & x_19024;
assign x_19026 = x_7783 & x_7784;
assign x_19027 = x_7782 & x_19026;
assign x_19028 = x_7786 & x_7787;
assign x_19029 = x_7785 & x_19028;
assign x_19030 = x_19027 & x_19029;
assign x_19031 = x_19025 & x_19030;
assign x_19032 = x_7788 & x_7789;
assign x_19033 = x_7791 & x_7792;
assign x_19034 = x_7790 & x_19033;
assign x_19035 = x_19032 & x_19034;
assign x_19036 = x_7794 & x_7795;
assign x_19037 = x_7793 & x_19036;
assign x_19038 = x_7797 & x_7798;
assign x_19039 = x_7796 & x_19038;
assign x_19040 = x_19037 & x_19039;
assign x_19041 = x_19035 & x_19040;
assign x_19042 = x_19031 & x_19041;
assign x_19043 = x_7799 & x_7800;
assign x_19044 = x_7802 & x_7803;
assign x_19045 = x_7801 & x_19044;
assign x_19046 = x_19043 & x_19045;
assign x_19047 = x_7805 & x_7806;
assign x_19048 = x_7804 & x_19047;
assign x_19049 = x_7808 & x_7809;
assign x_19050 = x_7807 & x_19049;
assign x_19051 = x_19048 & x_19050;
assign x_19052 = x_19046 & x_19051;
assign x_19053 = x_7810 & x_7811;
assign x_19054 = x_7813 & x_7814;
assign x_19055 = x_7812 & x_19054;
assign x_19056 = x_19053 & x_19055;
assign x_19057 = x_7816 & x_7817;
assign x_19058 = x_7815 & x_19057;
assign x_19059 = x_7819 & x_7820;
assign x_19060 = x_7818 & x_19059;
assign x_19061 = x_19058 & x_19060;
assign x_19062 = x_19056 & x_19061;
assign x_19063 = x_19052 & x_19062;
assign x_19064 = x_19042 & x_19063;
assign x_19065 = x_19021 & x_19064;
assign x_19066 = x_7821 & x_7822;
assign x_19067 = x_7824 & x_7825;
assign x_19068 = x_7823 & x_19067;
assign x_19069 = x_19066 & x_19068;
assign x_19070 = x_7827 & x_7828;
assign x_19071 = x_7826 & x_19070;
assign x_19072 = x_7830 & x_7831;
assign x_19073 = x_7829 & x_19072;
assign x_19074 = x_19071 & x_19073;
assign x_19075 = x_19069 & x_19074;
assign x_19076 = x_7832 & x_7833;
assign x_19077 = x_7835 & x_7836;
assign x_19078 = x_7834 & x_19077;
assign x_19079 = x_19076 & x_19078;
assign x_19080 = x_7838 & x_7839;
assign x_19081 = x_7837 & x_19080;
assign x_19082 = x_7841 & x_7842;
assign x_19083 = x_7840 & x_19082;
assign x_19084 = x_19081 & x_19083;
assign x_19085 = x_19079 & x_19084;
assign x_19086 = x_19075 & x_19085;
assign x_19087 = x_7843 & x_7844;
assign x_19088 = x_7846 & x_7847;
assign x_19089 = x_7845 & x_19088;
assign x_19090 = x_19087 & x_19089;
assign x_19091 = x_7849 & x_7850;
assign x_19092 = x_7848 & x_19091;
assign x_19093 = x_7852 & x_7853;
assign x_19094 = x_7851 & x_19093;
assign x_19095 = x_19092 & x_19094;
assign x_19096 = x_19090 & x_19095;
assign x_19097 = x_7854 & x_7855;
assign x_19098 = x_7857 & x_7858;
assign x_19099 = x_7856 & x_19098;
assign x_19100 = x_19097 & x_19099;
assign x_19101 = x_7860 & x_7861;
assign x_19102 = x_7859 & x_19101;
assign x_19103 = x_7863 & x_7864;
assign x_19104 = x_7862 & x_19103;
assign x_19105 = x_19102 & x_19104;
assign x_19106 = x_19100 & x_19105;
assign x_19107 = x_19096 & x_19106;
assign x_19108 = x_19086 & x_19107;
assign x_19109 = x_7865 & x_7866;
assign x_19110 = x_7868 & x_7869;
assign x_19111 = x_7867 & x_19110;
assign x_19112 = x_19109 & x_19111;
assign x_19113 = x_7871 & x_7872;
assign x_19114 = x_7870 & x_19113;
assign x_19115 = x_7874 & x_7875;
assign x_19116 = x_7873 & x_19115;
assign x_19117 = x_19114 & x_19116;
assign x_19118 = x_19112 & x_19117;
assign x_19119 = x_7876 & x_7877;
assign x_19120 = x_7879 & x_7880;
assign x_19121 = x_7878 & x_19120;
assign x_19122 = x_19119 & x_19121;
assign x_19123 = x_7882 & x_7883;
assign x_19124 = x_7881 & x_19123;
assign x_19125 = x_7885 & x_7886;
assign x_19126 = x_7884 & x_19125;
assign x_19127 = x_19124 & x_19126;
assign x_19128 = x_19122 & x_19127;
assign x_19129 = x_19118 & x_19128;
assign x_19130 = x_7887 & x_7888;
assign x_19131 = x_7890 & x_7891;
assign x_19132 = x_7889 & x_19131;
assign x_19133 = x_19130 & x_19132;
assign x_19134 = x_7893 & x_7894;
assign x_19135 = x_7892 & x_19134;
assign x_19136 = x_7896 & x_7897;
assign x_19137 = x_7895 & x_19136;
assign x_19138 = x_19135 & x_19137;
assign x_19139 = x_19133 & x_19138;
assign x_19140 = x_7898 & x_7899;
assign x_19141 = x_7901 & x_7902;
assign x_19142 = x_7900 & x_19141;
assign x_19143 = x_19140 & x_19142;
assign x_19144 = x_7904 & x_7905;
assign x_19145 = x_7903 & x_19144;
assign x_19146 = x_7907 & x_7908;
assign x_19147 = x_7906 & x_19146;
assign x_19148 = x_19145 & x_19147;
assign x_19149 = x_19143 & x_19148;
assign x_19150 = x_19139 & x_19149;
assign x_19151 = x_19129 & x_19150;
assign x_19152 = x_19108 & x_19151;
assign x_19153 = x_19065 & x_19152;
assign x_19154 = x_7909 & x_7910;
assign x_19155 = x_7912 & x_7913;
assign x_19156 = x_7911 & x_19155;
assign x_19157 = x_19154 & x_19156;
assign x_19158 = x_7915 & x_7916;
assign x_19159 = x_7914 & x_19158;
assign x_19160 = x_7918 & x_7919;
assign x_19161 = x_7917 & x_19160;
assign x_19162 = x_19159 & x_19161;
assign x_19163 = x_19157 & x_19162;
assign x_19164 = x_7920 & x_7921;
assign x_19165 = x_7923 & x_7924;
assign x_19166 = x_7922 & x_19165;
assign x_19167 = x_19164 & x_19166;
assign x_19168 = x_7926 & x_7927;
assign x_19169 = x_7925 & x_19168;
assign x_19170 = x_7929 & x_7930;
assign x_19171 = x_7928 & x_19170;
assign x_19172 = x_19169 & x_19171;
assign x_19173 = x_19167 & x_19172;
assign x_19174 = x_19163 & x_19173;
assign x_19175 = x_7931 & x_7932;
assign x_19176 = x_7934 & x_7935;
assign x_19177 = x_7933 & x_19176;
assign x_19178 = x_19175 & x_19177;
assign x_19179 = x_7937 & x_7938;
assign x_19180 = x_7936 & x_19179;
assign x_19181 = x_7940 & x_7941;
assign x_19182 = x_7939 & x_19181;
assign x_19183 = x_19180 & x_19182;
assign x_19184 = x_19178 & x_19183;
assign x_19185 = x_7942 & x_7943;
assign x_19186 = x_7945 & x_7946;
assign x_19187 = x_7944 & x_19186;
assign x_19188 = x_19185 & x_19187;
assign x_19189 = x_7948 & x_7949;
assign x_19190 = x_7947 & x_19189;
assign x_19191 = x_7951 & x_7952;
assign x_19192 = x_7950 & x_19191;
assign x_19193 = x_19190 & x_19192;
assign x_19194 = x_19188 & x_19193;
assign x_19195 = x_19184 & x_19194;
assign x_19196 = x_19174 & x_19195;
assign x_19197 = x_7953 & x_7954;
assign x_19198 = x_7956 & x_7957;
assign x_19199 = x_7955 & x_19198;
assign x_19200 = x_19197 & x_19199;
assign x_19201 = x_7959 & x_7960;
assign x_19202 = x_7958 & x_19201;
assign x_19203 = x_7962 & x_7963;
assign x_19204 = x_7961 & x_19203;
assign x_19205 = x_19202 & x_19204;
assign x_19206 = x_19200 & x_19205;
assign x_19207 = x_7964 & x_7965;
assign x_19208 = x_7967 & x_7968;
assign x_19209 = x_7966 & x_19208;
assign x_19210 = x_19207 & x_19209;
assign x_19211 = x_7970 & x_7971;
assign x_19212 = x_7969 & x_19211;
assign x_19213 = x_7973 & x_7974;
assign x_19214 = x_7972 & x_19213;
assign x_19215 = x_19212 & x_19214;
assign x_19216 = x_19210 & x_19215;
assign x_19217 = x_19206 & x_19216;
assign x_19218 = x_7975 & x_7976;
assign x_19219 = x_7978 & x_7979;
assign x_19220 = x_7977 & x_19219;
assign x_19221 = x_19218 & x_19220;
assign x_19222 = x_7981 & x_7982;
assign x_19223 = x_7980 & x_19222;
assign x_19224 = x_7984 & x_7985;
assign x_19225 = x_7983 & x_19224;
assign x_19226 = x_19223 & x_19225;
assign x_19227 = x_19221 & x_19226;
assign x_19228 = x_7986 & x_7987;
assign x_19229 = x_7989 & x_7990;
assign x_19230 = x_7988 & x_19229;
assign x_19231 = x_19228 & x_19230;
assign x_19232 = x_7992 & x_7993;
assign x_19233 = x_7991 & x_19232;
assign x_19234 = x_7995 & x_7996;
assign x_19235 = x_7994 & x_19234;
assign x_19236 = x_19233 & x_19235;
assign x_19237 = x_19231 & x_19236;
assign x_19238 = x_19227 & x_19237;
assign x_19239 = x_19217 & x_19238;
assign x_19240 = x_19196 & x_19239;
assign x_19241 = x_7997 & x_7998;
assign x_19242 = x_8000 & x_8001;
assign x_19243 = x_7999 & x_19242;
assign x_19244 = x_19241 & x_19243;
assign x_19245 = x_8003 & x_8004;
assign x_19246 = x_8002 & x_19245;
assign x_19247 = x_8006 & x_8007;
assign x_19248 = x_8005 & x_19247;
assign x_19249 = x_19246 & x_19248;
assign x_19250 = x_19244 & x_19249;
assign x_19251 = x_8008 & x_8009;
assign x_19252 = x_8011 & x_8012;
assign x_19253 = x_8010 & x_19252;
assign x_19254 = x_19251 & x_19253;
assign x_19255 = x_8014 & x_8015;
assign x_19256 = x_8013 & x_19255;
assign x_19257 = x_8017 & x_8018;
assign x_19258 = x_8016 & x_19257;
assign x_19259 = x_19256 & x_19258;
assign x_19260 = x_19254 & x_19259;
assign x_19261 = x_19250 & x_19260;
assign x_19262 = x_8019 & x_8020;
assign x_19263 = x_8022 & x_8023;
assign x_19264 = x_8021 & x_19263;
assign x_19265 = x_19262 & x_19264;
assign x_19266 = x_8025 & x_8026;
assign x_19267 = x_8024 & x_19266;
assign x_19268 = x_8028 & x_8029;
assign x_19269 = x_8027 & x_19268;
assign x_19270 = x_19267 & x_19269;
assign x_19271 = x_19265 & x_19270;
assign x_19272 = x_8030 & x_8031;
assign x_19273 = x_8033 & x_8034;
assign x_19274 = x_8032 & x_19273;
assign x_19275 = x_19272 & x_19274;
assign x_19276 = x_8036 & x_8037;
assign x_19277 = x_8035 & x_19276;
assign x_19278 = x_8039 & x_8040;
assign x_19279 = x_8038 & x_19278;
assign x_19280 = x_19277 & x_19279;
assign x_19281 = x_19275 & x_19280;
assign x_19282 = x_19271 & x_19281;
assign x_19283 = x_19261 & x_19282;
assign x_19284 = x_8041 & x_8042;
assign x_19285 = x_8044 & x_8045;
assign x_19286 = x_8043 & x_19285;
assign x_19287 = x_19284 & x_19286;
assign x_19288 = x_8047 & x_8048;
assign x_19289 = x_8046 & x_19288;
assign x_19290 = x_8050 & x_8051;
assign x_19291 = x_8049 & x_19290;
assign x_19292 = x_19289 & x_19291;
assign x_19293 = x_19287 & x_19292;
assign x_19294 = x_8052 & x_8053;
assign x_19295 = x_8055 & x_8056;
assign x_19296 = x_8054 & x_19295;
assign x_19297 = x_19294 & x_19296;
assign x_19298 = x_8058 & x_8059;
assign x_19299 = x_8057 & x_19298;
assign x_19300 = x_8061 & x_8062;
assign x_19301 = x_8060 & x_19300;
assign x_19302 = x_19299 & x_19301;
assign x_19303 = x_19297 & x_19302;
assign x_19304 = x_19293 & x_19303;
assign x_19305 = x_8063 & x_8064;
assign x_19306 = x_8066 & x_8067;
assign x_19307 = x_8065 & x_19306;
assign x_19308 = x_19305 & x_19307;
assign x_19309 = x_8069 & x_8070;
assign x_19310 = x_8068 & x_19309;
assign x_19311 = x_8072 & x_8073;
assign x_19312 = x_8071 & x_19311;
assign x_19313 = x_19310 & x_19312;
assign x_19314 = x_19308 & x_19313;
assign x_19315 = x_8074 & x_8075;
assign x_19316 = x_8077 & x_8078;
assign x_19317 = x_8076 & x_19316;
assign x_19318 = x_19315 & x_19317;
assign x_19319 = x_8080 & x_8081;
assign x_19320 = x_8079 & x_19319;
assign x_19321 = x_8083 & x_8084;
assign x_19322 = x_8082 & x_19321;
assign x_19323 = x_19320 & x_19322;
assign x_19324 = x_19318 & x_19323;
assign x_19325 = x_19314 & x_19324;
assign x_19326 = x_19304 & x_19325;
assign x_19327 = x_19283 & x_19326;
assign x_19328 = x_19240 & x_19327;
assign x_19329 = x_19153 & x_19328;
assign x_19330 = x_8085 & x_8086;
assign x_19331 = x_8088 & x_8089;
assign x_19332 = x_8087 & x_19331;
assign x_19333 = x_19330 & x_19332;
assign x_19334 = x_8091 & x_8092;
assign x_19335 = x_8090 & x_19334;
assign x_19336 = x_8094 & x_8095;
assign x_19337 = x_8093 & x_19336;
assign x_19338 = x_19335 & x_19337;
assign x_19339 = x_19333 & x_19338;
assign x_19340 = x_8096 & x_8097;
assign x_19341 = x_8099 & x_8100;
assign x_19342 = x_8098 & x_19341;
assign x_19343 = x_19340 & x_19342;
assign x_19344 = x_8102 & x_8103;
assign x_19345 = x_8101 & x_19344;
assign x_19346 = x_8105 & x_8106;
assign x_19347 = x_8104 & x_19346;
assign x_19348 = x_19345 & x_19347;
assign x_19349 = x_19343 & x_19348;
assign x_19350 = x_19339 & x_19349;
assign x_19351 = x_8107 & x_8108;
assign x_19352 = x_8110 & x_8111;
assign x_19353 = x_8109 & x_19352;
assign x_19354 = x_19351 & x_19353;
assign x_19355 = x_8113 & x_8114;
assign x_19356 = x_8112 & x_19355;
assign x_19357 = x_8116 & x_8117;
assign x_19358 = x_8115 & x_19357;
assign x_19359 = x_19356 & x_19358;
assign x_19360 = x_19354 & x_19359;
assign x_19361 = x_8118 & x_8119;
assign x_19362 = x_8121 & x_8122;
assign x_19363 = x_8120 & x_19362;
assign x_19364 = x_19361 & x_19363;
assign x_19365 = x_8124 & x_8125;
assign x_19366 = x_8123 & x_19365;
assign x_19367 = x_8127 & x_8128;
assign x_19368 = x_8126 & x_19367;
assign x_19369 = x_19366 & x_19368;
assign x_19370 = x_19364 & x_19369;
assign x_19371 = x_19360 & x_19370;
assign x_19372 = x_19350 & x_19371;
assign x_19373 = x_8129 & x_8130;
assign x_19374 = x_8132 & x_8133;
assign x_19375 = x_8131 & x_19374;
assign x_19376 = x_19373 & x_19375;
assign x_19377 = x_8135 & x_8136;
assign x_19378 = x_8134 & x_19377;
assign x_19379 = x_8138 & x_8139;
assign x_19380 = x_8137 & x_19379;
assign x_19381 = x_19378 & x_19380;
assign x_19382 = x_19376 & x_19381;
assign x_19383 = x_8140 & x_8141;
assign x_19384 = x_8143 & x_8144;
assign x_19385 = x_8142 & x_19384;
assign x_19386 = x_19383 & x_19385;
assign x_19387 = x_8146 & x_8147;
assign x_19388 = x_8145 & x_19387;
assign x_19389 = x_8149 & x_8150;
assign x_19390 = x_8148 & x_19389;
assign x_19391 = x_19388 & x_19390;
assign x_19392 = x_19386 & x_19391;
assign x_19393 = x_19382 & x_19392;
assign x_19394 = x_8151 & x_8152;
assign x_19395 = x_8154 & x_8155;
assign x_19396 = x_8153 & x_19395;
assign x_19397 = x_19394 & x_19396;
assign x_19398 = x_8157 & x_8158;
assign x_19399 = x_8156 & x_19398;
assign x_19400 = x_8160 & x_8161;
assign x_19401 = x_8159 & x_19400;
assign x_19402 = x_19399 & x_19401;
assign x_19403 = x_19397 & x_19402;
assign x_19404 = x_8162 & x_8163;
assign x_19405 = x_8165 & x_8166;
assign x_19406 = x_8164 & x_19405;
assign x_19407 = x_19404 & x_19406;
assign x_19408 = x_8168 & x_8169;
assign x_19409 = x_8167 & x_19408;
assign x_19410 = x_8171 & x_8172;
assign x_19411 = x_8170 & x_19410;
assign x_19412 = x_19409 & x_19411;
assign x_19413 = x_19407 & x_19412;
assign x_19414 = x_19403 & x_19413;
assign x_19415 = x_19393 & x_19414;
assign x_19416 = x_19372 & x_19415;
assign x_19417 = x_8173 & x_8174;
assign x_19418 = x_8176 & x_8177;
assign x_19419 = x_8175 & x_19418;
assign x_19420 = x_19417 & x_19419;
assign x_19421 = x_8179 & x_8180;
assign x_19422 = x_8178 & x_19421;
assign x_19423 = x_8182 & x_8183;
assign x_19424 = x_8181 & x_19423;
assign x_19425 = x_19422 & x_19424;
assign x_19426 = x_19420 & x_19425;
assign x_19427 = x_8184 & x_8185;
assign x_19428 = x_8187 & x_8188;
assign x_19429 = x_8186 & x_19428;
assign x_19430 = x_19427 & x_19429;
assign x_19431 = x_8190 & x_8191;
assign x_19432 = x_8189 & x_19431;
assign x_19433 = x_8193 & x_8194;
assign x_19434 = x_8192 & x_19433;
assign x_19435 = x_19432 & x_19434;
assign x_19436 = x_19430 & x_19435;
assign x_19437 = x_19426 & x_19436;
assign x_19438 = x_8195 & x_8196;
assign x_19439 = x_8198 & x_8199;
assign x_19440 = x_8197 & x_19439;
assign x_19441 = x_19438 & x_19440;
assign x_19442 = x_8201 & x_8202;
assign x_19443 = x_8200 & x_19442;
assign x_19444 = x_8204 & x_8205;
assign x_19445 = x_8203 & x_19444;
assign x_19446 = x_19443 & x_19445;
assign x_19447 = x_19441 & x_19446;
assign x_19448 = x_8206 & x_8207;
assign x_19449 = x_8209 & x_8210;
assign x_19450 = x_8208 & x_19449;
assign x_19451 = x_19448 & x_19450;
assign x_19452 = x_8212 & x_8213;
assign x_19453 = x_8211 & x_19452;
assign x_19454 = x_8215 & x_8216;
assign x_19455 = x_8214 & x_19454;
assign x_19456 = x_19453 & x_19455;
assign x_19457 = x_19451 & x_19456;
assign x_19458 = x_19447 & x_19457;
assign x_19459 = x_19437 & x_19458;
assign x_19460 = x_8217 & x_8218;
assign x_19461 = x_8220 & x_8221;
assign x_19462 = x_8219 & x_19461;
assign x_19463 = x_19460 & x_19462;
assign x_19464 = x_8223 & x_8224;
assign x_19465 = x_8222 & x_19464;
assign x_19466 = x_8226 & x_8227;
assign x_19467 = x_8225 & x_19466;
assign x_19468 = x_19465 & x_19467;
assign x_19469 = x_19463 & x_19468;
assign x_19470 = x_8228 & x_8229;
assign x_19471 = x_8231 & x_8232;
assign x_19472 = x_8230 & x_19471;
assign x_19473 = x_19470 & x_19472;
assign x_19474 = x_8234 & x_8235;
assign x_19475 = x_8233 & x_19474;
assign x_19476 = x_8237 & x_8238;
assign x_19477 = x_8236 & x_19476;
assign x_19478 = x_19475 & x_19477;
assign x_19479 = x_19473 & x_19478;
assign x_19480 = x_19469 & x_19479;
assign x_19481 = x_8239 & x_8240;
assign x_19482 = x_8242 & x_8243;
assign x_19483 = x_8241 & x_19482;
assign x_19484 = x_19481 & x_19483;
assign x_19485 = x_8245 & x_8246;
assign x_19486 = x_8244 & x_19485;
assign x_19487 = x_8248 & x_8249;
assign x_19488 = x_8247 & x_19487;
assign x_19489 = x_19486 & x_19488;
assign x_19490 = x_19484 & x_19489;
assign x_19491 = x_8250 & x_8251;
assign x_19492 = x_8253 & x_8254;
assign x_19493 = x_8252 & x_19492;
assign x_19494 = x_19491 & x_19493;
assign x_19495 = x_8256 & x_8257;
assign x_19496 = x_8255 & x_19495;
assign x_19497 = x_8259 & x_8260;
assign x_19498 = x_8258 & x_19497;
assign x_19499 = x_19496 & x_19498;
assign x_19500 = x_19494 & x_19499;
assign x_19501 = x_19490 & x_19500;
assign x_19502 = x_19480 & x_19501;
assign x_19503 = x_19459 & x_19502;
assign x_19504 = x_19416 & x_19503;
assign x_19505 = x_8261 & x_8262;
assign x_19506 = x_8264 & x_8265;
assign x_19507 = x_8263 & x_19506;
assign x_19508 = x_19505 & x_19507;
assign x_19509 = x_8267 & x_8268;
assign x_19510 = x_8266 & x_19509;
assign x_19511 = x_8270 & x_8271;
assign x_19512 = x_8269 & x_19511;
assign x_19513 = x_19510 & x_19512;
assign x_19514 = x_19508 & x_19513;
assign x_19515 = x_8272 & x_8273;
assign x_19516 = x_8275 & x_8276;
assign x_19517 = x_8274 & x_19516;
assign x_19518 = x_19515 & x_19517;
assign x_19519 = x_8278 & x_8279;
assign x_19520 = x_8277 & x_19519;
assign x_19521 = x_8281 & x_8282;
assign x_19522 = x_8280 & x_19521;
assign x_19523 = x_19520 & x_19522;
assign x_19524 = x_19518 & x_19523;
assign x_19525 = x_19514 & x_19524;
assign x_19526 = x_8283 & x_8284;
assign x_19527 = x_8286 & x_8287;
assign x_19528 = x_8285 & x_19527;
assign x_19529 = x_19526 & x_19528;
assign x_19530 = x_8289 & x_8290;
assign x_19531 = x_8288 & x_19530;
assign x_19532 = x_8292 & x_8293;
assign x_19533 = x_8291 & x_19532;
assign x_19534 = x_19531 & x_19533;
assign x_19535 = x_19529 & x_19534;
assign x_19536 = x_8294 & x_8295;
assign x_19537 = x_8297 & x_8298;
assign x_19538 = x_8296 & x_19537;
assign x_19539 = x_19536 & x_19538;
assign x_19540 = x_8300 & x_8301;
assign x_19541 = x_8299 & x_19540;
assign x_19542 = x_8303 & x_8304;
assign x_19543 = x_8302 & x_19542;
assign x_19544 = x_19541 & x_19543;
assign x_19545 = x_19539 & x_19544;
assign x_19546 = x_19535 & x_19545;
assign x_19547 = x_19525 & x_19546;
assign x_19548 = x_8305 & x_8306;
assign x_19549 = x_8308 & x_8309;
assign x_19550 = x_8307 & x_19549;
assign x_19551 = x_19548 & x_19550;
assign x_19552 = x_8311 & x_8312;
assign x_19553 = x_8310 & x_19552;
assign x_19554 = x_8314 & x_8315;
assign x_19555 = x_8313 & x_19554;
assign x_19556 = x_19553 & x_19555;
assign x_19557 = x_19551 & x_19556;
assign x_19558 = x_8316 & x_8317;
assign x_19559 = x_8319 & x_8320;
assign x_19560 = x_8318 & x_19559;
assign x_19561 = x_19558 & x_19560;
assign x_19562 = x_8322 & x_8323;
assign x_19563 = x_8321 & x_19562;
assign x_19564 = x_8325 & x_8326;
assign x_19565 = x_8324 & x_19564;
assign x_19566 = x_19563 & x_19565;
assign x_19567 = x_19561 & x_19566;
assign x_19568 = x_19557 & x_19567;
assign x_19569 = x_8327 & x_8328;
assign x_19570 = x_8330 & x_8331;
assign x_19571 = x_8329 & x_19570;
assign x_19572 = x_19569 & x_19571;
assign x_19573 = x_8333 & x_8334;
assign x_19574 = x_8332 & x_19573;
assign x_19575 = x_8336 & x_8337;
assign x_19576 = x_8335 & x_19575;
assign x_19577 = x_19574 & x_19576;
assign x_19578 = x_19572 & x_19577;
assign x_19579 = x_8338 & x_8339;
assign x_19580 = x_8341 & x_8342;
assign x_19581 = x_8340 & x_19580;
assign x_19582 = x_19579 & x_19581;
assign x_19583 = x_8344 & x_8345;
assign x_19584 = x_8343 & x_19583;
assign x_19585 = x_8347 & x_8348;
assign x_19586 = x_8346 & x_19585;
assign x_19587 = x_19584 & x_19586;
assign x_19588 = x_19582 & x_19587;
assign x_19589 = x_19578 & x_19588;
assign x_19590 = x_19568 & x_19589;
assign x_19591 = x_19547 & x_19590;
assign x_19592 = x_8349 & x_8350;
assign x_19593 = x_8352 & x_8353;
assign x_19594 = x_8351 & x_19593;
assign x_19595 = x_19592 & x_19594;
assign x_19596 = x_8355 & x_8356;
assign x_19597 = x_8354 & x_19596;
assign x_19598 = x_8358 & x_8359;
assign x_19599 = x_8357 & x_19598;
assign x_19600 = x_19597 & x_19599;
assign x_19601 = x_19595 & x_19600;
assign x_19602 = x_8360 & x_8361;
assign x_19603 = x_8363 & x_8364;
assign x_19604 = x_8362 & x_19603;
assign x_19605 = x_19602 & x_19604;
assign x_19606 = x_8366 & x_8367;
assign x_19607 = x_8365 & x_19606;
assign x_19608 = x_8369 & x_8370;
assign x_19609 = x_8368 & x_19608;
assign x_19610 = x_19607 & x_19609;
assign x_19611 = x_19605 & x_19610;
assign x_19612 = x_19601 & x_19611;
assign x_19613 = x_8371 & x_8372;
assign x_19614 = x_8374 & x_8375;
assign x_19615 = x_8373 & x_19614;
assign x_19616 = x_19613 & x_19615;
assign x_19617 = x_8377 & x_8378;
assign x_19618 = x_8376 & x_19617;
assign x_19619 = x_8380 & x_8381;
assign x_19620 = x_8379 & x_19619;
assign x_19621 = x_19618 & x_19620;
assign x_19622 = x_19616 & x_19621;
assign x_19623 = x_8382 & x_8383;
assign x_19624 = x_8385 & x_8386;
assign x_19625 = x_8384 & x_19624;
assign x_19626 = x_19623 & x_19625;
assign x_19627 = x_8388 & x_8389;
assign x_19628 = x_8387 & x_19627;
assign x_19629 = x_8391 & x_8392;
assign x_19630 = x_8390 & x_19629;
assign x_19631 = x_19628 & x_19630;
assign x_19632 = x_19626 & x_19631;
assign x_19633 = x_19622 & x_19632;
assign x_19634 = x_19612 & x_19633;
assign x_19635 = x_8393 & x_8394;
assign x_19636 = x_8396 & x_8397;
assign x_19637 = x_8395 & x_19636;
assign x_19638 = x_19635 & x_19637;
assign x_19639 = x_8399 & x_8400;
assign x_19640 = x_8398 & x_19639;
assign x_19641 = x_8402 & x_8403;
assign x_19642 = x_8401 & x_19641;
assign x_19643 = x_19640 & x_19642;
assign x_19644 = x_19638 & x_19643;
assign x_19645 = x_8404 & x_8405;
assign x_19646 = x_8407 & x_8408;
assign x_19647 = x_8406 & x_19646;
assign x_19648 = x_19645 & x_19647;
assign x_19649 = x_8410 & x_8411;
assign x_19650 = x_8409 & x_19649;
assign x_19651 = x_8413 & x_8414;
assign x_19652 = x_8412 & x_19651;
assign x_19653 = x_19650 & x_19652;
assign x_19654 = x_19648 & x_19653;
assign x_19655 = x_19644 & x_19654;
assign x_19656 = x_8415 & x_8416;
assign x_19657 = x_8418 & x_8419;
assign x_19658 = x_8417 & x_19657;
assign x_19659 = x_19656 & x_19658;
assign x_19660 = x_8421 & x_8422;
assign x_19661 = x_8420 & x_19660;
assign x_19662 = x_8424 & x_8425;
assign x_19663 = x_8423 & x_19662;
assign x_19664 = x_19661 & x_19663;
assign x_19665 = x_19659 & x_19664;
assign x_19666 = x_8426 & x_8427;
assign x_19667 = x_8429 & x_8430;
assign x_19668 = x_8428 & x_19667;
assign x_19669 = x_19666 & x_19668;
assign x_19670 = x_8432 & x_8433;
assign x_19671 = x_8431 & x_19670;
assign x_19672 = x_8435 & x_8436;
assign x_19673 = x_8434 & x_19672;
assign x_19674 = x_19671 & x_19673;
assign x_19675 = x_19669 & x_19674;
assign x_19676 = x_19665 & x_19675;
assign x_19677 = x_19655 & x_19676;
assign x_19678 = x_19634 & x_19677;
assign x_19679 = x_19591 & x_19678;
assign x_19680 = x_19504 & x_19679;
assign x_19681 = x_19329 & x_19680;
assign x_19682 = x_18979 & x_19681;
assign x_19683 = x_18277 & x_19682;
assign x_19684 = x_8437 & x_8438;
assign x_19685 = x_8440 & x_8441;
assign x_19686 = x_8439 & x_19685;
assign x_19687 = x_19684 & x_19686;
assign x_19688 = x_8442 & x_8443;
assign x_19689 = x_8445 & x_8446;
assign x_19690 = x_8444 & x_19689;
assign x_19691 = x_19688 & x_19690;
assign x_19692 = x_19687 & x_19691;
assign x_19693 = x_8447 & x_8448;
assign x_19694 = x_8450 & x_8451;
assign x_19695 = x_8449 & x_19694;
assign x_19696 = x_19693 & x_19695;
assign x_19697 = x_8453 & x_8454;
assign x_19698 = x_8452 & x_19697;
assign x_19699 = x_8456 & x_8457;
assign x_19700 = x_8455 & x_19699;
assign x_19701 = x_19698 & x_19700;
assign x_19702 = x_19696 & x_19701;
assign x_19703 = x_19692 & x_19702;
assign x_19704 = x_8458 & x_8459;
assign x_19705 = x_8461 & x_8462;
assign x_19706 = x_8460 & x_19705;
assign x_19707 = x_19704 & x_19706;
assign x_19708 = x_8464 & x_8465;
assign x_19709 = x_8463 & x_19708;
assign x_19710 = x_8467 & x_8468;
assign x_19711 = x_8466 & x_19710;
assign x_19712 = x_19709 & x_19711;
assign x_19713 = x_19707 & x_19712;
assign x_19714 = x_8469 & x_8470;
assign x_19715 = x_8472 & x_8473;
assign x_19716 = x_8471 & x_19715;
assign x_19717 = x_19714 & x_19716;
assign x_19718 = x_8475 & x_8476;
assign x_19719 = x_8474 & x_19718;
assign x_19720 = x_8478 & x_8479;
assign x_19721 = x_8477 & x_19720;
assign x_19722 = x_19719 & x_19721;
assign x_19723 = x_19717 & x_19722;
assign x_19724 = x_19713 & x_19723;
assign x_19725 = x_19703 & x_19724;
assign x_19726 = x_8480 & x_8481;
assign x_19727 = x_8483 & x_8484;
assign x_19728 = x_8482 & x_19727;
assign x_19729 = x_19726 & x_19728;
assign x_19730 = x_8486 & x_8487;
assign x_19731 = x_8485 & x_19730;
assign x_19732 = x_8489 & x_8490;
assign x_19733 = x_8488 & x_19732;
assign x_19734 = x_19731 & x_19733;
assign x_19735 = x_19729 & x_19734;
assign x_19736 = x_8491 & x_8492;
assign x_19737 = x_8494 & x_8495;
assign x_19738 = x_8493 & x_19737;
assign x_19739 = x_19736 & x_19738;
assign x_19740 = x_8497 & x_8498;
assign x_19741 = x_8496 & x_19740;
assign x_19742 = x_8500 & x_8501;
assign x_19743 = x_8499 & x_19742;
assign x_19744 = x_19741 & x_19743;
assign x_19745 = x_19739 & x_19744;
assign x_19746 = x_19735 & x_19745;
assign x_19747 = x_8502 & x_8503;
assign x_19748 = x_8505 & x_8506;
assign x_19749 = x_8504 & x_19748;
assign x_19750 = x_19747 & x_19749;
assign x_19751 = x_8508 & x_8509;
assign x_19752 = x_8507 & x_19751;
assign x_19753 = x_8511 & x_8512;
assign x_19754 = x_8510 & x_19753;
assign x_19755 = x_19752 & x_19754;
assign x_19756 = x_19750 & x_19755;
assign x_19757 = x_8513 & x_8514;
assign x_19758 = x_8516 & x_8517;
assign x_19759 = x_8515 & x_19758;
assign x_19760 = x_19757 & x_19759;
assign x_19761 = x_8519 & x_8520;
assign x_19762 = x_8518 & x_19761;
assign x_19763 = x_8522 & x_8523;
assign x_19764 = x_8521 & x_19763;
assign x_19765 = x_19762 & x_19764;
assign x_19766 = x_19760 & x_19765;
assign x_19767 = x_19756 & x_19766;
assign x_19768 = x_19746 & x_19767;
assign x_19769 = x_19725 & x_19768;
assign x_19770 = x_8524 & x_8525;
assign x_19771 = x_8527 & x_8528;
assign x_19772 = x_8526 & x_19771;
assign x_19773 = x_19770 & x_19772;
assign x_19774 = x_8530 & x_8531;
assign x_19775 = x_8529 & x_19774;
assign x_19776 = x_8533 & x_8534;
assign x_19777 = x_8532 & x_19776;
assign x_19778 = x_19775 & x_19777;
assign x_19779 = x_19773 & x_19778;
assign x_19780 = x_8535 & x_8536;
assign x_19781 = x_8538 & x_8539;
assign x_19782 = x_8537 & x_19781;
assign x_19783 = x_19780 & x_19782;
assign x_19784 = x_8541 & x_8542;
assign x_19785 = x_8540 & x_19784;
assign x_19786 = x_8544 & x_8545;
assign x_19787 = x_8543 & x_19786;
assign x_19788 = x_19785 & x_19787;
assign x_19789 = x_19783 & x_19788;
assign x_19790 = x_19779 & x_19789;
assign x_19791 = x_8546 & x_8547;
assign x_19792 = x_8549 & x_8550;
assign x_19793 = x_8548 & x_19792;
assign x_19794 = x_19791 & x_19793;
assign x_19795 = x_8552 & x_8553;
assign x_19796 = x_8551 & x_19795;
assign x_19797 = x_8555 & x_8556;
assign x_19798 = x_8554 & x_19797;
assign x_19799 = x_19796 & x_19798;
assign x_19800 = x_19794 & x_19799;
assign x_19801 = x_8557 & x_8558;
assign x_19802 = x_8560 & x_8561;
assign x_19803 = x_8559 & x_19802;
assign x_19804 = x_19801 & x_19803;
assign x_19805 = x_8563 & x_8564;
assign x_19806 = x_8562 & x_19805;
assign x_19807 = x_8566 & x_8567;
assign x_19808 = x_8565 & x_19807;
assign x_19809 = x_19806 & x_19808;
assign x_19810 = x_19804 & x_19809;
assign x_19811 = x_19800 & x_19810;
assign x_19812 = x_19790 & x_19811;
assign x_19813 = x_8568 & x_8569;
assign x_19814 = x_8571 & x_8572;
assign x_19815 = x_8570 & x_19814;
assign x_19816 = x_19813 & x_19815;
assign x_19817 = x_8574 & x_8575;
assign x_19818 = x_8573 & x_19817;
assign x_19819 = x_8577 & x_8578;
assign x_19820 = x_8576 & x_19819;
assign x_19821 = x_19818 & x_19820;
assign x_19822 = x_19816 & x_19821;
assign x_19823 = x_8579 & x_8580;
assign x_19824 = x_8582 & x_8583;
assign x_19825 = x_8581 & x_19824;
assign x_19826 = x_19823 & x_19825;
assign x_19827 = x_8585 & x_8586;
assign x_19828 = x_8584 & x_19827;
assign x_19829 = x_8588 & x_8589;
assign x_19830 = x_8587 & x_19829;
assign x_19831 = x_19828 & x_19830;
assign x_19832 = x_19826 & x_19831;
assign x_19833 = x_19822 & x_19832;
assign x_19834 = x_8590 & x_8591;
assign x_19835 = x_8593 & x_8594;
assign x_19836 = x_8592 & x_19835;
assign x_19837 = x_19834 & x_19836;
assign x_19838 = x_8596 & x_8597;
assign x_19839 = x_8595 & x_19838;
assign x_19840 = x_8599 & x_8600;
assign x_19841 = x_8598 & x_19840;
assign x_19842 = x_19839 & x_19841;
assign x_19843 = x_19837 & x_19842;
assign x_19844 = x_8601 & x_8602;
assign x_19845 = x_8604 & x_8605;
assign x_19846 = x_8603 & x_19845;
assign x_19847 = x_19844 & x_19846;
assign x_19848 = x_8607 & x_8608;
assign x_19849 = x_8606 & x_19848;
assign x_19850 = x_8610 & x_8611;
assign x_19851 = x_8609 & x_19850;
assign x_19852 = x_19849 & x_19851;
assign x_19853 = x_19847 & x_19852;
assign x_19854 = x_19843 & x_19853;
assign x_19855 = x_19833 & x_19854;
assign x_19856 = x_19812 & x_19855;
assign x_19857 = x_19769 & x_19856;
assign x_19858 = x_8612 & x_8613;
assign x_19859 = x_8615 & x_8616;
assign x_19860 = x_8614 & x_19859;
assign x_19861 = x_19858 & x_19860;
assign x_19862 = x_8618 & x_8619;
assign x_19863 = x_8617 & x_19862;
assign x_19864 = x_8621 & x_8622;
assign x_19865 = x_8620 & x_19864;
assign x_19866 = x_19863 & x_19865;
assign x_19867 = x_19861 & x_19866;
assign x_19868 = x_8623 & x_8624;
assign x_19869 = x_8626 & x_8627;
assign x_19870 = x_8625 & x_19869;
assign x_19871 = x_19868 & x_19870;
assign x_19872 = x_8629 & x_8630;
assign x_19873 = x_8628 & x_19872;
assign x_19874 = x_8632 & x_8633;
assign x_19875 = x_8631 & x_19874;
assign x_19876 = x_19873 & x_19875;
assign x_19877 = x_19871 & x_19876;
assign x_19878 = x_19867 & x_19877;
assign x_19879 = x_8634 & x_8635;
assign x_19880 = x_8637 & x_8638;
assign x_19881 = x_8636 & x_19880;
assign x_19882 = x_19879 & x_19881;
assign x_19883 = x_8640 & x_8641;
assign x_19884 = x_8639 & x_19883;
assign x_19885 = x_8643 & x_8644;
assign x_19886 = x_8642 & x_19885;
assign x_19887 = x_19884 & x_19886;
assign x_19888 = x_19882 & x_19887;
assign x_19889 = x_8645 & x_8646;
assign x_19890 = x_8648 & x_8649;
assign x_19891 = x_8647 & x_19890;
assign x_19892 = x_19889 & x_19891;
assign x_19893 = x_8651 & x_8652;
assign x_19894 = x_8650 & x_19893;
assign x_19895 = x_8654 & x_8655;
assign x_19896 = x_8653 & x_19895;
assign x_19897 = x_19894 & x_19896;
assign x_19898 = x_19892 & x_19897;
assign x_19899 = x_19888 & x_19898;
assign x_19900 = x_19878 & x_19899;
assign x_19901 = x_8656 & x_8657;
assign x_19902 = x_8659 & x_8660;
assign x_19903 = x_8658 & x_19902;
assign x_19904 = x_19901 & x_19903;
assign x_19905 = x_8662 & x_8663;
assign x_19906 = x_8661 & x_19905;
assign x_19907 = x_8665 & x_8666;
assign x_19908 = x_8664 & x_19907;
assign x_19909 = x_19906 & x_19908;
assign x_19910 = x_19904 & x_19909;
assign x_19911 = x_8667 & x_8668;
assign x_19912 = x_8670 & x_8671;
assign x_19913 = x_8669 & x_19912;
assign x_19914 = x_19911 & x_19913;
assign x_19915 = x_8673 & x_8674;
assign x_19916 = x_8672 & x_19915;
assign x_19917 = x_8676 & x_8677;
assign x_19918 = x_8675 & x_19917;
assign x_19919 = x_19916 & x_19918;
assign x_19920 = x_19914 & x_19919;
assign x_19921 = x_19910 & x_19920;
assign x_19922 = x_8678 & x_8679;
assign x_19923 = x_8681 & x_8682;
assign x_19924 = x_8680 & x_19923;
assign x_19925 = x_19922 & x_19924;
assign x_19926 = x_8684 & x_8685;
assign x_19927 = x_8683 & x_19926;
assign x_19928 = x_8687 & x_8688;
assign x_19929 = x_8686 & x_19928;
assign x_19930 = x_19927 & x_19929;
assign x_19931 = x_19925 & x_19930;
assign x_19932 = x_8689 & x_8690;
assign x_19933 = x_8692 & x_8693;
assign x_19934 = x_8691 & x_19933;
assign x_19935 = x_19932 & x_19934;
assign x_19936 = x_8695 & x_8696;
assign x_19937 = x_8694 & x_19936;
assign x_19938 = x_8698 & x_8699;
assign x_19939 = x_8697 & x_19938;
assign x_19940 = x_19937 & x_19939;
assign x_19941 = x_19935 & x_19940;
assign x_19942 = x_19931 & x_19941;
assign x_19943 = x_19921 & x_19942;
assign x_19944 = x_19900 & x_19943;
assign x_19945 = x_8700 & x_8701;
assign x_19946 = x_8703 & x_8704;
assign x_19947 = x_8702 & x_19946;
assign x_19948 = x_19945 & x_19947;
assign x_19949 = x_8706 & x_8707;
assign x_19950 = x_8705 & x_19949;
assign x_19951 = x_8709 & x_8710;
assign x_19952 = x_8708 & x_19951;
assign x_19953 = x_19950 & x_19952;
assign x_19954 = x_19948 & x_19953;
assign x_19955 = x_8711 & x_8712;
assign x_19956 = x_8714 & x_8715;
assign x_19957 = x_8713 & x_19956;
assign x_19958 = x_19955 & x_19957;
assign x_19959 = x_8717 & x_8718;
assign x_19960 = x_8716 & x_19959;
assign x_19961 = x_8720 & x_8721;
assign x_19962 = x_8719 & x_19961;
assign x_19963 = x_19960 & x_19962;
assign x_19964 = x_19958 & x_19963;
assign x_19965 = x_19954 & x_19964;
assign x_19966 = x_8722 & x_8723;
assign x_19967 = x_8725 & x_8726;
assign x_19968 = x_8724 & x_19967;
assign x_19969 = x_19966 & x_19968;
assign x_19970 = x_8728 & x_8729;
assign x_19971 = x_8727 & x_19970;
assign x_19972 = x_8731 & x_8732;
assign x_19973 = x_8730 & x_19972;
assign x_19974 = x_19971 & x_19973;
assign x_19975 = x_19969 & x_19974;
assign x_19976 = x_8733 & x_8734;
assign x_19977 = x_8736 & x_8737;
assign x_19978 = x_8735 & x_19977;
assign x_19979 = x_19976 & x_19978;
assign x_19980 = x_8739 & x_8740;
assign x_19981 = x_8738 & x_19980;
assign x_19982 = x_8742 & x_8743;
assign x_19983 = x_8741 & x_19982;
assign x_19984 = x_19981 & x_19983;
assign x_19985 = x_19979 & x_19984;
assign x_19986 = x_19975 & x_19985;
assign x_19987 = x_19965 & x_19986;
assign x_19988 = x_8744 & x_8745;
assign x_19989 = x_8747 & x_8748;
assign x_19990 = x_8746 & x_19989;
assign x_19991 = x_19988 & x_19990;
assign x_19992 = x_8750 & x_8751;
assign x_19993 = x_8749 & x_19992;
assign x_19994 = x_8753 & x_8754;
assign x_19995 = x_8752 & x_19994;
assign x_19996 = x_19993 & x_19995;
assign x_19997 = x_19991 & x_19996;
assign x_19998 = x_8755 & x_8756;
assign x_19999 = x_8758 & x_8759;
assign x_20000 = x_8757 & x_19999;
assign x_20001 = x_19998 & x_20000;
assign x_20002 = x_8761 & x_8762;
assign x_20003 = x_8760 & x_20002;
assign x_20004 = x_8764 & x_8765;
assign x_20005 = x_8763 & x_20004;
assign x_20006 = x_20003 & x_20005;
assign x_20007 = x_20001 & x_20006;
assign x_20008 = x_19997 & x_20007;
assign x_20009 = x_8766 & x_8767;
assign x_20010 = x_8769 & x_8770;
assign x_20011 = x_8768 & x_20010;
assign x_20012 = x_20009 & x_20011;
assign x_20013 = x_8772 & x_8773;
assign x_20014 = x_8771 & x_20013;
assign x_20015 = x_8775 & x_8776;
assign x_20016 = x_8774 & x_20015;
assign x_20017 = x_20014 & x_20016;
assign x_20018 = x_20012 & x_20017;
assign x_20019 = x_8777 & x_8778;
assign x_20020 = x_8780 & x_8781;
assign x_20021 = x_8779 & x_20020;
assign x_20022 = x_20019 & x_20021;
assign x_20023 = x_8783 & x_8784;
assign x_20024 = x_8782 & x_20023;
assign x_20025 = x_8786 & x_8787;
assign x_20026 = x_8785 & x_20025;
assign x_20027 = x_20024 & x_20026;
assign x_20028 = x_20022 & x_20027;
assign x_20029 = x_20018 & x_20028;
assign x_20030 = x_20008 & x_20029;
assign x_20031 = x_19987 & x_20030;
assign x_20032 = x_19944 & x_20031;
assign x_20033 = x_19857 & x_20032;
assign x_20034 = x_8788 & x_8789;
assign x_20035 = x_8791 & x_8792;
assign x_20036 = x_8790 & x_20035;
assign x_20037 = x_20034 & x_20036;
assign x_20038 = x_8794 & x_8795;
assign x_20039 = x_8793 & x_20038;
assign x_20040 = x_8797 & x_8798;
assign x_20041 = x_8796 & x_20040;
assign x_20042 = x_20039 & x_20041;
assign x_20043 = x_20037 & x_20042;
assign x_20044 = x_8799 & x_8800;
assign x_20045 = x_8802 & x_8803;
assign x_20046 = x_8801 & x_20045;
assign x_20047 = x_20044 & x_20046;
assign x_20048 = x_8805 & x_8806;
assign x_20049 = x_8804 & x_20048;
assign x_20050 = x_8808 & x_8809;
assign x_20051 = x_8807 & x_20050;
assign x_20052 = x_20049 & x_20051;
assign x_20053 = x_20047 & x_20052;
assign x_20054 = x_20043 & x_20053;
assign x_20055 = x_8810 & x_8811;
assign x_20056 = x_8813 & x_8814;
assign x_20057 = x_8812 & x_20056;
assign x_20058 = x_20055 & x_20057;
assign x_20059 = x_8816 & x_8817;
assign x_20060 = x_8815 & x_20059;
assign x_20061 = x_8819 & x_8820;
assign x_20062 = x_8818 & x_20061;
assign x_20063 = x_20060 & x_20062;
assign x_20064 = x_20058 & x_20063;
assign x_20065 = x_8821 & x_8822;
assign x_20066 = x_8824 & x_8825;
assign x_20067 = x_8823 & x_20066;
assign x_20068 = x_20065 & x_20067;
assign x_20069 = x_8827 & x_8828;
assign x_20070 = x_8826 & x_20069;
assign x_20071 = x_8830 & x_8831;
assign x_20072 = x_8829 & x_20071;
assign x_20073 = x_20070 & x_20072;
assign x_20074 = x_20068 & x_20073;
assign x_20075 = x_20064 & x_20074;
assign x_20076 = x_20054 & x_20075;
assign x_20077 = x_8832 & x_8833;
assign x_20078 = x_8835 & x_8836;
assign x_20079 = x_8834 & x_20078;
assign x_20080 = x_20077 & x_20079;
assign x_20081 = x_8838 & x_8839;
assign x_20082 = x_8837 & x_20081;
assign x_20083 = x_8841 & x_8842;
assign x_20084 = x_8840 & x_20083;
assign x_20085 = x_20082 & x_20084;
assign x_20086 = x_20080 & x_20085;
assign x_20087 = x_8843 & x_8844;
assign x_20088 = x_8846 & x_8847;
assign x_20089 = x_8845 & x_20088;
assign x_20090 = x_20087 & x_20089;
assign x_20091 = x_8849 & x_8850;
assign x_20092 = x_8848 & x_20091;
assign x_20093 = x_8852 & x_8853;
assign x_20094 = x_8851 & x_20093;
assign x_20095 = x_20092 & x_20094;
assign x_20096 = x_20090 & x_20095;
assign x_20097 = x_20086 & x_20096;
assign x_20098 = x_8854 & x_8855;
assign x_20099 = x_8857 & x_8858;
assign x_20100 = x_8856 & x_20099;
assign x_20101 = x_20098 & x_20100;
assign x_20102 = x_8860 & x_8861;
assign x_20103 = x_8859 & x_20102;
assign x_20104 = x_8863 & x_8864;
assign x_20105 = x_8862 & x_20104;
assign x_20106 = x_20103 & x_20105;
assign x_20107 = x_20101 & x_20106;
assign x_20108 = x_8865 & x_8866;
assign x_20109 = x_8868 & x_8869;
assign x_20110 = x_8867 & x_20109;
assign x_20111 = x_20108 & x_20110;
assign x_20112 = x_8871 & x_8872;
assign x_20113 = x_8870 & x_20112;
assign x_20114 = x_8874 & x_8875;
assign x_20115 = x_8873 & x_20114;
assign x_20116 = x_20113 & x_20115;
assign x_20117 = x_20111 & x_20116;
assign x_20118 = x_20107 & x_20117;
assign x_20119 = x_20097 & x_20118;
assign x_20120 = x_20076 & x_20119;
assign x_20121 = x_8876 & x_8877;
assign x_20122 = x_8879 & x_8880;
assign x_20123 = x_8878 & x_20122;
assign x_20124 = x_20121 & x_20123;
assign x_20125 = x_8882 & x_8883;
assign x_20126 = x_8881 & x_20125;
assign x_20127 = x_8885 & x_8886;
assign x_20128 = x_8884 & x_20127;
assign x_20129 = x_20126 & x_20128;
assign x_20130 = x_20124 & x_20129;
assign x_20131 = x_8887 & x_8888;
assign x_20132 = x_8890 & x_8891;
assign x_20133 = x_8889 & x_20132;
assign x_20134 = x_20131 & x_20133;
assign x_20135 = x_8893 & x_8894;
assign x_20136 = x_8892 & x_20135;
assign x_20137 = x_8896 & x_8897;
assign x_20138 = x_8895 & x_20137;
assign x_20139 = x_20136 & x_20138;
assign x_20140 = x_20134 & x_20139;
assign x_20141 = x_20130 & x_20140;
assign x_20142 = x_8898 & x_8899;
assign x_20143 = x_8901 & x_8902;
assign x_20144 = x_8900 & x_20143;
assign x_20145 = x_20142 & x_20144;
assign x_20146 = x_8904 & x_8905;
assign x_20147 = x_8903 & x_20146;
assign x_20148 = x_8907 & x_8908;
assign x_20149 = x_8906 & x_20148;
assign x_20150 = x_20147 & x_20149;
assign x_20151 = x_20145 & x_20150;
assign x_20152 = x_8909 & x_8910;
assign x_20153 = x_8912 & x_8913;
assign x_20154 = x_8911 & x_20153;
assign x_20155 = x_20152 & x_20154;
assign x_20156 = x_8915 & x_8916;
assign x_20157 = x_8914 & x_20156;
assign x_20158 = x_8918 & x_8919;
assign x_20159 = x_8917 & x_20158;
assign x_20160 = x_20157 & x_20159;
assign x_20161 = x_20155 & x_20160;
assign x_20162 = x_20151 & x_20161;
assign x_20163 = x_20141 & x_20162;
assign x_20164 = x_8920 & x_8921;
assign x_20165 = x_8923 & x_8924;
assign x_20166 = x_8922 & x_20165;
assign x_20167 = x_20164 & x_20166;
assign x_20168 = x_8926 & x_8927;
assign x_20169 = x_8925 & x_20168;
assign x_20170 = x_8929 & x_8930;
assign x_20171 = x_8928 & x_20170;
assign x_20172 = x_20169 & x_20171;
assign x_20173 = x_20167 & x_20172;
assign x_20174 = x_8931 & x_8932;
assign x_20175 = x_8934 & x_8935;
assign x_20176 = x_8933 & x_20175;
assign x_20177 = x_20174 & x_20176;
assign x_20178 = x_8937 & x_8938;
assign x_20179 = x_8936 & x_20178;
assign x_20180 = x_8940 & x_8941;
assign x_20181 = x_8939 & x_20180;
assign x_20182 = x_20179 & x_20181;
assign x_20183 = x_20177 & x_20182;
assign x_20184 = x_20173 & x_20183;
assign x_20185 = x_8942 & x_8943;
assign x_20186 = x_8945 & x_8946;
assign x_20187 = x_8944 & x_20186;
assign x_20188 = x_20185 & x_20187;
assign x_20189 = x_8948 & x_8949;
assign x_20190 = x_8947 & x_20189;
assign x_20191 = x_8951 & x_8952;
assign x_20192 = x_8950 & x_20191;
assign x_20193 = x_20190 & x_20192;
assign x_20194 = x_20188 & x_20193;
assign x_20195 = x_8953 & x_8954;
assign x_20196 = x_8956 & x_8957;
assign x_20197 = x_8955 & x_20196;
assign x_20198 = x_20195 & x_20197;
assign x_20199 = x_8959 & x_8960;
assign x_20200 = x_8958 & x_20199;
assign x_20201 = x_8962 & x_8963;
assign x_20202 = x_8961 & x_20201;
assign x_20203 = x_20200 & x_20202;
assign x_20204 = x_20198 & x_20203;
assign x_20205 = x_20194 & x_20204;
assign x_20206 = x_20184 & x_20205;
assign x_20207 = x_20163 & x_20206;
assign x_20208 = x_20120 & x_20207;
assign x_20209 = x_8964 & x_8965;
assign x_20210 = x_8967 & x_8968;
assign x_20211 = x_8966 & x_20210;
assign x_20212 = x_20209 & x_20211;
assign x_20213 = x_8970 & x_8971;
assign x_20214 = x_8969 & x_20213;
assign x_20215 = x_8973 & x_8974;
assign x_20216 = x_8972 & x_20215;
assign x_20217 = x_20214 & x_20216;
assign x_20218 = x_20212 & x_20217;
assign x_20219 = x_8975 & x_8976;
assign x_20220 = x_8978 & x_8979;
assign x_20221 = x_8977 & x_20220;
assign x_20222 = x_20219 & x_20221;
assign x_20223 = x_8981 & x_8982;
assign x_20224 = x_8980 & x_20223;
assign x_20225 = x_8984 & x_8985;
assign x_20226 = x_8983 & x_20225;
assign x_20227 = x_20224 & x_20226;
assign x_20228 = x_20222 & x_20227;
assign x_20229 = x_20218 & x_20228;
assign x_20230 = x_8986 & x_8987;
assign x_20231 = x_8989 & x_8990;
assign x_20232 = x_8988 & x_20231;
assign x_20233 = x_20230 & x_20232;
assign x_20234 = x_8992 & x_8993;
assign x_20235 = x_8991 & x_20234;
assign x_20236 = x_8995 & x_8996;
assign x_20237 = x_8994 & x_20236;
assign x_20238 = x_20235 & x_20237;
assign x_20239 = x_20233 & x_20238;
assign x_20240 = x_8997 & x_8998;
assign x_20241 = x_9000 & x_9001;
assign x_20242 = x_8999 & x_20241;
assign x_20243 = x_20240 & x_20242;
assign x_20244 = x_9003 & x_9004;
assign x_20245 = x_9002 & x_20244;
assign x_20246 = x_9006 & x_9007;
assign x_20247 = x_9005 & x_20246;
assign x_20248 = x_20245 & x_20247;
assign x_20249 = x_20243 & x_20248;
assign x_20250 = x_20239 & x_20249;
assign x_20251 = x_20229 & x_20250;
assign x_20252 = x_9008 & x_9009;
assign x_20253 = x_9011 & x_9012;
assign x_20254 = x_9010 & x_20253;
assign x_20255 = x_20252 & x_20254;
assign x_20256 = x_9014 & x_9015;
assign x_20257 = x_9013 & x_20256;
assign x_20258 = x_9017 & x_9018;
assign x_20259 = x_9016 & x_20258;
assign x_20260 = x_20257 & x_20259;
assign x_20261 = x_20255 & x_20260;
assign x_20262 = x_9019 & x_9020;
assign x_20263 = x_9022 & x_9023;
assign x_20264 = x_9021 & x_20263;
assign x_20265 = x_20262 & x_20264;
assign x_20266 = x_9025 & x_9026;
assign x_20267 = x_9024 & x_20266;
assign x_20268 = x_9028 & x_9029;
assign x_20269 = x_9027 & x_20268;
assign x_20270 = x_20267 & x_20269;
assign x_20271 = x_20265 & x_20270;
assign x_20272 = x_20261 & x_20271;
assign x_20273 = x_9030 & x_9031;
assign x_20274 = x_9033 & x_9034;
assign x_20275 = x_9032 & x_20274;
assign x_20276 = x_20273 & x_20275;
assign x_20277 = x_9036 & x_9037;
assign x_20278 = x_9035 & x_20277;
assign x_20279 = x_9039 & x_9040;
assign x_20280 = x_9038 & x_20279;
assign x_20281 = x_20278 & x_20280;
assign x_20282 = x_20276 & x_20281;
assign x_20283 = x_9041 & x_9042;
assign x_20284 = x_9044 & x_9045;
assign x_20285 = x_9043 & x_20284;
assign x_20286 = x_20283 & x_20285;
assign x_20287 = x_9047 & x_9048;
assign x_20288 = x_9046 & x_20287;
assign x_20289 = x_9050 & x_9051;
assign x_20290 = x_9049 & x_20289;
assign x_20291 = x_20288 & x_20290;
assign x_20292 = x_20286 & x_20291;
assign x_20293 = x_20282 & x_20292;
assign x_20294 = x_20272 & x_20293;
assign x_20295 = x_20251 & x_20294;
assign x_20296 = x_9052 & x_9053;
assign x_20297 = x_9055 & x_9056;
assign x_20298 = x_9054 & x_20297;
assign x_20299 = x_20296 & x_20298;
assign x_20300 = x_9058 & x_9059;
assign x_20301 = x_9057 & x_20300;
assign x_20302 = x_9061 & x_9062;
assign x_20303 = x_9060 & x_20302;
assign x_20304 = x_20301 & x_20303;
assign x_20305 = x_20299 & x_20304;
assign x_20306 = x_9063 & x_9064;
assign x_20307 = x_9066 & x_9067;
assign x_20308 = x_9065 & x_20307;
assign x_20309 = x_20306 & x_20308;
assign x_20310 = x_9069 & x_9070;
assign x_20311 = x_9068 & x_20310;
assign x_20312 = x_9072 & x_9073;
assign x_20313 = x_9071 & x_20312;
assign x_20314 = x_20311 & x_20313;
assign x_20315 = x_20309 & x_20314;
assign x_20316 = x_20305 & x_20315;
assign x_20317 = x_9074 & x_9075;
assign x_20318 = x_9077 & x_9078;
assign x_20319 = x_9076 & x_20318;
assign x_20320 = x_20317 & x_20319;
assign x_20321 = x_9080 & x_9081;
assign x_20322 = x_9079 & x_20321;
assign x_20323 = x_9083 & x_9084;
assign x_20324 = x_9082 & x_20323;
assign x_20325 = x_20322 & x_20324;
assign x_20326 = x_20320 & x_20325;
assign x_20327 = x_9085 & x_9086;
assign x_20328 = x_9088 & x_9089;
assign x_20329 = x_9087 & x_20328;
assign x_20330 = x_20327 & x_20329;
assign x_20331 = x_9091 & x_9092;
assign x_20332 = x_9090 & x_20331;
assign x_20333 = x_9094 & x_9095;
assign x_20334 = x_9093 & x_20333;
assign x_20335 = x_20332 & x_20334;
assign x_20336 = x_20330 & x_20335;
assign x_20337 = x_20326 & x_20336;
assign x_20338 = x_20316 & x_20337;
assign x_20339 = x_9096 & x_9097;
assign x_20340 = x_9099 & x_9100;
assign x_20341 = x_9098 & x_20340;
assign x_20342 = x_20339 & x_20341;
assign x_20343 = x_9102 & x_9103;
assign x_20344 = x_9101 & x_20343;
assign x_20345 = x_9105 & x_9106;
assign x_20346 = x_9104 & x_20345;
assign x_20347 = x_20344 & x_20346;
assign x_20348 = x_20342 & x_20347;
assign x_20349 = x_9107 & x_9108;
assign x_20350 = x_9110 & x_9111;
assign x_20351 = x_9109 & x_20350;
assign x_20352 = x_20349 & x_20351;
assign x_20353 = x_9113 & x_9114;
assign x_20354 = x_9112 & x_20353;
assign x_20355 = x_9116 & x_9117;
assign x_20356 = x_9115 & x_20355;
assign x_20357 = x_20354 & x_20356;
assign x_20358 = x_20352 & x_20357;
assign x_20359 = x_20348 & x_20358;
assign x_20360 = x_9118 & x_9119;
assign x_20361 = x_9121 & x_9122;
assign x_20362 = x_9120 & x_20361;
assign x_20363 = x_20360 & x_20362;
assign x_20364 = x_9124 & x_9125;
assign x_20365 = x_9123 & x_20364;
assign x_20366 = x_9127 & x_9128;
assign x_20367 = x_9126 & x_20366;
assign x_20368 = x_20365 & x_20367;
assign x_20369 = x_20363 & x_20368;
assign x_20370 = x_9129 & x_9130;
assign x_20371 = x_9132 & x_9133;
assign x_20372 = x_9131 & x_20371;
assign x_20373 = x_20370 & x_20372;
assign x_20374 = x_9135 & x_9136;
assign x_20375 = x_9134 & x_20374;
assign x_20376 = x_9138 & x_9139;
assign x_20377 = x_9137 & x_20376;
assign x_20378 = x_20375 & x_20377;
assign x_20379 = x_20373 & x_20378;
assign x_20380 = x_20369 & x_20379;
assign x_20381 = x_20359 & x_20380;
assign x_20382 = x_20338 & x_20381;
assign x_20383 = x_20295 & x_20382;
assign x_20384 = x_20208 & x_20383;
assign x_20385 = x_20033 & x_20384;
assign x_20386 = x_9140 & x_9141;
assign x_20387 = x_9143 & x_9144;
assign x_20388 = x_9142 & x_20387;
assign x_20389 = x_20386 & x_20388;
assign x_20390 = x_9145 & x_9146;
assign x_20391 = x_9148 & x_9149;
assign x_20392 = x_9147 & x_20391;
assign x_20393 = x_20390 & x_20392;
assign x_20394 = x_20389 & x_20393;
assign x_20395 = x_9150 & x_9151;
assign x_20396 = x_9153 & x_9154;
assign x_20397 = x_9152 & x_20396;
assign x_20398 = x_20395 & x_20397;
assign x_20399 = x_9156 & x_9157;
assign x_20400 = x_9155 & x_20399;
assign x_20401 = x_9159 & x_9160;
assign x_20402 = x_9158 & x_20401;
assign x_20403 = x_20400 & x_20402;
assign x_20404 = x_20398 & x_20403;
assign x_20405 = x_20394 & x_20404;
assign x_20406 = x_9161 & x_9162;
assign x_20407 = x_9164 & x_9165;
assign x_20408 = x_9163 & x_20407;
assign x_20409 = x_20406 & x_20408;
assign x_20410 = x_9167 & x_9168;
assign x_20411 = x_9166 & x_20410;
assign x_20412 = x_9170 & x_9171;
assign x_20413 = x_9169 & x_20412;
assign x_20414 = x_20411 & x_20413;
assign x_20415 = x_20409 & x_20414;
assign x_20416 = x_9172 & x_9173;
assign x_20417 = x_9175 & x_9176;
assign x_20418 = x_9174 & x_20417;
assign x_20419 = x_20416 & x_20418;
assign x_20420 = x_9178 & x_9179;
assign x_20421 = x_9177 & x_20420;
assign x_20422 = x_9181 & x_9182;
assign x_20423 = x_9180 & x_20422;
assign x_20424 = x_20421 & x_20423;
assign x_20425 = x_20419 & x_20424;
assign x_20426 = x_20415 & x_20425;
assign x_20427 = x_20405 & x_20426;
assign x_20428 = x_9183 & x_9184;
assign x_20429 = x_9186 & x_9187;
assign x_20430 = x_9185 & x_20429;
assign x_20431 = x_20428 & x_20430;
assign x_20432 = x_9189 & x_9190;
assign x_20433 = x_9188 & x_20432;
assign x_20434 = x_9192 & x_9193;
assign x_20435 = x_9191 & x_20434;
assign x_20436 = x_20433 & x_20435;
assign x_20437 = x_20431 & x_20436;
assign x_20438 = x_9194 & x_9195;
assign x_20439 = x_9197 & x_9198;
assign x_20440 = x_9196 & x_20439;
assign x_20441 = x_20438 & x_20440;
assign x_20442 = x_9200 & x_9201;
assign x_20443 = x_9199 & x_20442;
assign x_20444 = x_9203 & x_9204;
assign x_20445 = x_9202 & x_20444;
assign x_20446 = x_20443 & x_20445;
assign x_20447 = x_20441 & x_20446;
assign x_20448 = x_20437 & x_20447;
assign x_20449 = x_9205 & x_9206;
assign x_20450 = x_9208 & x_9209;
assign x_20451 = x_9207 & x_20450;
assign x_20452 = x_20449 & x_20451;
assign x_20453 = x_9211 & x_9212;
assign x_20454 = x_9210 & x_20453;
assign x_20455 = x_9214 & x_9215;
assign x_20456 = x_9213 & x_20455;
assign x_20457 = x_20454 & x_20456;
assign x_20458 = x_20452 & x_20457;
assign x_20459 = x_9216 & x_9217;
assign x_20460 = x_9219 & x_9220;
assign x_20461 = x_9218 & x_20460;
assign x_20462 = x_20459 & x_20461;
assign x_20463 = x_9222 & x_9223;
assign x_20464 = x_9221 & x_20463;
assign x_20465 = x_9225 & x_9226;
assign x_20466 = x_9224 & x_20465;
assign x_20467 = x_20464 & x_20466;
assign x_20468 = x_20462 & x_20467;
assign x_20469 = x_20458 & x_20468;
assign x_20470 = x_20448 & x_20469;
assign x_20471 = x_20427 & x_20470;
assign x_20472 = x_9227 & x_9228;
assign x_20473 = x_9230 & x_9231;
assign x_20474 = x_9229 & x_20473;
assign x_20475 = x_20472 & x_20474;
assign x_20476 = x_9233 & x_9234;
assign x_20477 = x_9232 & x_20476;
assign x_20478 = x_9236 & x_9237;
assign x_20479 = x_9235 & x_20478;
assign x_20480 = x_20477 & x_20479;
assign x_20481 = x_20475 & x_20480;
assign x_20482 = x_9238 & x_9239;
assign x_20483 = x_9241 & x_9242;
assign x_20484 = x_9240 & x_20483;
assign x_20485 = x_20482 & x_20484;
assign x_20486 = x_9244 & x_9245;
assign x_20487 = x_9243 & x_20486;
assign x_20488 = x_9247 & x_9248;
assign x_20489 = x_9246 & x_20488;
assign x_20490 = x_20487 & x_20489;
assign x_20491 = x_20485 & x_20490;
assign x_20492 = x_20481 & x_20491;
assign x_20493 = x_9249 & x_9250;
assign x_20494 = x_9252 & x_9253;
assign x_20495 = x_9251 & x_20494;
assign x_20496 = x_20493 & x_20495;
assign x_20497 = x_9255 & x_9256;
assign x_20498 = x_9254 & x_20497;
assign x_20499 = x_9258 & x_9259;
assign x_20500 = x_9257 & x_20499;
assign x_20501 = x_20498 & x_20500;
assign x_20502 = x_20496 & x_20501;
assign x_20503 = x_9260 & x_9261;
assign x_20504 = x_9263 & x_9264;
assign x_20505 = x_9262 & x_20504;
assign x_20506 = x_20503 & x_20505;
assign x_20507 = x_9266 & x_9267;
assign x_20508 = x_9265 & x_20507;
assign x_20509 = x_9269 & x_9270;
assign x_20510 = x_9268 & x_20509;
assign x_20511 = x_20508 & x_20510;
assign x_20512 = x_20506 & x_20511;
assign x_20513 = x_20502 & x_20512;
assign x_20514 = x_20492 & x_20513;
assign x_20515 = x_9271 & x_9272;
assign x_20516 = x_9274 & x_9275;
assign x_20517 = x_9273 & x_20516;
assign x_20518 = x_20515 & x_20517;
assign x_20519 = x_9277 & x_9278;
assign x_20520 = x_9276 & x_20519;
assign x_20521 = x_9280 & x_9281;
assign x_20522 = x_9279 & x_20521;
assign x_20523 = x_20520 & x_20522;
assign x_20524 = x_20518 & x_20523;
assign x_20525 = x_9282 & x_9283;
assign x_20526 = x_9285 & x_9286;
assign x_20527 = x_9284 & x_20526;
assign x_20528 = x_20525 & x_20527;
assign x_20529 = x_9288 & x_9289;
assign x_20530 = x_9287 & x_20529;
assign x_20531 = x_9291 & x_9292;
assign x_20532 = x_9290 & x_20531;
assign x_20533 = x_20530 & x_20532;
assign x_20534 = x_20528 & x_20533;
assign x_20535 = x_20524 & x_20534;
assign x_20536 = x_9293 & x_9294;
assign x_20537 = x_9296 & x_9297;
assign x_20538 = x_9295 & x_20537;
assign x_20539 = x_20536 & x_20538;
assign x_20540 = x_9299 & x_9300;
assign x_20541 = x_9298 & x_20540;
assign x_20542 = x_9302 & x_9303;
assign x_20543 = x_9301 & x_20542;
assign x_20544 = x_20541 & x_20543;
assign x_20545 = x_20539 & x_20544;
assign x_20546 = x_9304 & x_9305;
assign x_20547 = x_9307 & x_9308;
assign x_20548 = x_9306 & x_20547;
assign x_20549 = x_20546 & x_20548;
assign x_20550 = x_9310 & x_9311;
assign x_20551 = x_9309 & x_20550;
assign x_20552 = x_9313 & x_9314;
assign x_20553 = x_9312 & x_20552;
assign x_20554 = x_20551 & x_20553;
assign x_20555 = x_20549 & x_20554;
assign x_20556 = x_20545 & x_20555;
assign x_20557 = x_20535 & x_20556;
assign x_20558 = x_20514 & x_20557;
assign x_20559 = x_20471 & x_20558;
assign x_20560 = x_9315 & x_9316;
assign x_20561 = x_9318 & x_9319;
assign x_20562 = x_9317 & x_20561;
assign x_20563 = x_20560 & x_20562;
assign x_20564 = x_9321 & x_9322;
assign x_20565 = x_9320 & x_20564;
assign x_20566 = x_9324 & x_9325;
assign x_20567 = x_9323 & x_20566;
assign x_20568 = x_20565 & x_20567;
assign x_20569 = x_20563 & x_20568;
assign x_20570 = x_9326 & x_9327;
assign x_20571 = x_9329 & x_9330;
assign x_20572 = x_9328 & x_20571;
assign x_20573 = x_20570 & x_20572;
assign x_20574 = x_9332 & x_9333;
assign x_20575 = x_9331 & x_20574;
assign x_20576 = x_9335 & x_9336;
assign x_20577 = x_9334 & x_20576;
assign x_20578 = x_20575 & x_20577;
assign x_20579 = x_20573 & x_20578;
assign x_20580 = x_20569 & x_20579;
assign x_20581 = x_9337 & x_9338;
assign x_20582 = x_9340 & x_9341;
assign x_20583 = x_9339 & x_20582;
assign x_20584 = x_20581 & x_20583;
assign x_20585 = x_9343 & x_9344;
assign x_20586 = x_9342 & x_20585;
assign x_20587 = x_9346 & x_9347;
assign x_20588 = x_9345 & x_20587;
assign x_20589 = x_20586 & x_20588;
assign x_20590 = x_20584 & x_20589;
assign x_20591 = x_9348 & x_9349;
assign x_20592 = x_9351 & x_9352;
assign x_20593 = x_9350 & x_20592;
assign x_20594 = x_20591 & x_20593;
assign x_20595 = x_9354 & x_9355;
assign x_20596 = x_9353 & x_20595;
assign x_20597 = x_9357 & x_9358;
assign x_20598 = x_9356 & x_20597;
assign x_20599 = x_20596 & x_20598;
assign x_20600 = x_20594 & x_20599;
assign x_20601 = x_20590 & x_20600;
assign x_20602 = x_20580 & x_20601;
assign x_20603 = x_9359 & x_9360;
assign x_20604 = x_9362 & x_9363;
assign x_20605 = x_9361 & x_20604;
assign x_20606 = x_20603 & x_20605;
assign x_20607 = x_9365 & x_9366;
assign x_20608 = x_9364 & x_20607;
assign x_20609 = x_9368 & x_9369;
assign x_20610 = x_9367 & x_20609;
assign x_20611 = x_20608 & x_20610;
assign x_20612 = x_20606 & x_20611;
assign x_20613 = x_9370 & x_9371;
assign x_20614 = x_9373 & x_9374;
assign x_20615 = x_9372 & x_20614;
assign x_20616 = x_20613 & x_20615;
assign x_20617 = x_9376 & x_9377;
assign x_20618 = x_9375 & x_20617;
assign x_20619 = x_9379 & x_9380;
assign x_20620 = x_9378 & x_20619;
assign x_20621 = x_20618 & x_20620;
assign x_20622 = x_20616 & x_20621;
assign x_20623 = x_20612 & x_20622;
assign x_20624 = x_9381 & x_9382;
assign x_20625 = x_9384 & x_9385;
assign x_20626 = x_9383 & x_20625;
assign x_20627 = x_20624 & x_20626;
assign x_20628 = x_9387 & x_9388;
assign x_20629 = x_9386 & x_20628;
assign x_20630 = x_9390 & x_9391;
assign x_20631 = x_9389 & x_20630;
assign x_20632 = x_20629 & x_20631;
assign x_20633 = x_20627 & x_20632;
assign x_20634 = x_9392 & x_9393;
assign x_20635 = x_9395 & x_9396;
assign x_20636 = x_9394 & x_20635;
assign x_20637 = x_20634 & x_20636;
assign x_20638 = x_9398 & x_9399;
assign x_20639 = x_9397 & x_20638;
assign x_20640 = x_9401 & x_9402;
assign x_20641 = x_9400 & x_20640;
assign x_20642 = x_20639 & x_20641;
assign x_20643 = x_20637 & x_20642;
assign x_20644 = x_20633 & x_20643;
assign x_20645 = x_20623 & x_20644;
assign x_20646 = x_20602 & x_20645;
assign x_20647 = x_9403 & x_9404;
assign x_20648 = x_9406 & x_9407;
assign x_20649 = x_9405 & x_20648;
assign x_20650 = x_20647 & x_20649;
assign x_20651 = x_9409 & x_9410;
assign x_20652 = x_9408 & x_20651;
assign x_20653 = x_9412 & x_9413;
assign x_20654 = x_9411 & x_20653;
assign x_20655 = x_20652 & x_20654;
assign x_20656 = x_20650 & x_20655;
assign x_20657 = x_9414 & x_9415;
assign x_20658 = x_9417 & x_9418;
assign x_20659 = x_9416 & x_20658;
assign x_20660 = x_20657 & x_20659;
assign x_20661 = x_9420 & x_9421;
assign x_20662 = x_9419 & x_20661;
assign x_20663 = x_9423 & x_9424;
assign x_20664 = x_9422 & x_20663;
assign x_20665 = x_20662 & x_20664;
assign x_20666 = x_20660 & x_20665;
assign x_20667 = x_20656 & x_20666;
assign x_20668 = x_9425 & x_9426;
assign x_20669 = x_9428 & x_9429;
assign x_20670 = x_9427 & x_20669;
assign x_20671 = x_20668 & x_20670;
assign x_20672 = x_9431 & x_9432;
assign x_20673 = x_9430 & x_20672;
assign x_20674 = x_9434 & x_9435;
assign x_20675 = x_9433 & x_20674;
assign x_20676 = x_20673 & x_20675;
assign x_20677 = x_20671 & x_20676;
assign x_20678 = x_9436 & x_9437;
assign x_20679 = x_9439 & x_9440;
assign x_20680 = x_9438 & x_20679;
assign x_20681 = x_20678 & x_20680;
assign x_20682 = x_9442 & x_9443;
assign x_20683 = x_9441 & x_20682;
assign x_20684 = x_9445 & x_9446;
assign x_20685 = x_9444 & x_20684;
assign x_20686 = x_20683 & x_20685;
assign x_20687 = x_20681 & x_20686;
assign x_20688 = x_20677 & x_20687;
assign x_20689 = x_20667 & x_20688;
assign x_20690 = x_9447 & x_9448;
assign x_20691 = x_9450 & x_9451;
assign x_20692 = x_9449 & x_20691;
assign x_20693 = x_20690 & x_20692;
assign x_20694 = x_9453 & x_9454;
assign x_20695 = x_9452 & x_20694;
assign x_20696 = x_9456 & x_9457;
assign x_20697 = x_9455 & x_20696;
assign x_20698 = x_20695 & x_20697;
assign x_20699 = x_20693 & x_20698;
assign x_20700 = x_9458 & x_9459;
assign x_20701 = x_9461 & x_9462;
assign x_20702 = x_9460 & x_20701;
assign x_20703 = x_20700 & x_20702;
assign x_20704 = x_9464 & x_9465;
assign x_20705 = x_9463 & x_20704;
assign x_20706 = x_9467 & x_9468;
assign x_20707 = x_9466 & x_20706;
assign x_20708 = x_20705 & x_20707;
assign x_20709 = x_20703 & x_20708;
assign x_20710 = x_20699 & x_20709;
assign x_20711 = x_9469 & x_9470;
assign x_20712 = x_9472 & x_9473;
assign x_20713 = x_9471 & x_20712;
assign x_20714 = x_20711 & x_20713;
assign x_20715 = x_9475 & x_9476;
assign x_20716 = x_9474 & x_20715;
assign x_20717 = x_9478 & x_9479;
assign x_20718 = x_9477 & x_20717;
assign x_20719 = x_20716 & x_20718;
assign x_20720 = x_20714 & x_20719;
assign x_20721 = x_9480 & x_9481;
assign x_20722 = x_9483 & x_9484;
assign x_20723 = x_9482 & x_20722;
assign x_20724 = x_20721 & x_20723;
assign x_20725 = x_9486 & x_9487;
assign x_20726 = x_9485 & x_20725;
assign x_20727 = x_9489 & x_9490;
assign x_20728 = x_9488 & x_20727;
assign x_20729 = x_20726 & x_20728;
assign x_20730 = x_20724 & x_20729;
assign x_20731 = x_20720 & x_20730;
assign x_20732 = x_20710 & x_20731;
assign x_20733 = x_20689 & x_20732;
assign x_20734 = x_20646 & x_20733;
assign x_20735 = x_20559 & x_20734;
assign x_20736 = x_9491 & x_9492;
assign x_20737 = x_9494 & x_9495;
assign x_20738 = x_9493 & x_20737;
assign x_20739 = x_20736 & x_20738;
assign x_20740 = x_9497 & x_9498;
assign x_20741 = x_9496 & x_20740;
assign x_20742 = x_9500 & x_9501;
assign x_20743 = x_9499 & x_20742;
assign x_20744 = x_20741 & x_20743;
assign x_20745 = x_20739 & x_20744;
assign x_20746 = x_9502 & x_9503;
assign x_20747 = x_9505 & x_9506;
assign x_20748 = x_9504 & x_20747;
assign x_20749 = x_20746 & x_20748;
assign x_20750 = x_9508 & x_9509;
assign x_20751 = x_9507 & x_20750;
assign x_20752 = x_9511 & x_9512;
assign x_20753 = x_9510 & x_20752;
assign x_20754 = x_20751 & x_20753;
assign x_20755 = x_20749 & x_20754;
assign x_20756 = x_20745 & x_20755;
assign x_20757 = x_9513 & x_9514;
assign x_20758 = x_9516 & x_9517;
assign x_20759 = x_9515 & x_20758;
assign x_20760 = x_20757 & x_20759;
assign x_20761 = x_9519 & x_9520;
assign x_20762 = x_9518 & x_20761;
assign x_20763 = x_9522 & x_9523;
assign x_20764 = x_9521 & x_20763;
assign x_20765 = x_20762 & x_20764;
assign x_20766 = x_20760 & x_20765;
assign x_20767 = x_9524 & x_9525;
assign x_20768 = x_9527 & x_9528;
assign x_20769 = x_9526 & x_20768;
assign x_20770 = x_20767 & x_20769;
assign x_20771 = x_9530 & x_9531;
assign x_20772 = x_9529 & x_20771;
assign x_20773 = x_9533 & x_9534;
assign x_20774 = x_9532 & x_20773;
assign x_20775 = x_20772 & x_20774;
assign x_20776 = x_20770 & x_20775;
assign x_20777 = x_20766 & x_20776;
assign x_20778 = x_20756 & x_20777;
assign x_20779 = x_9535 & x_9536;
assign x_20780 = x_9538 & x_9539;
assign x_20781 = x_9537 & x_20780;
assign x_20782 = x_20779 & x_20781;
assign x_20783 = x_9541 & x_9542;
assign x_20784 = x_9540 & x_20783;
assign x_20785 = x_9544 & x_9545;
assign x_20786 = x_9543 & x_20785;
assign x_20787 = x_20784 & x_20786;
assign x_20788 = x_20782 & x_20787;
assign x_20789 = x_9546 & x_9547;
assign x_20790 = x_9549 & x_9550;
assign x_20791 = x_9548 & x_20790;
assign x_20792 = x_20789 & x_20791;
assign x_20793 = x_9552 & x_9553;
assign x_20794 = x_9551 & x_20793;
assign x_20795 = x_9555 & x_9556;
assign x_20796 = x_9554 & x_20795;
assign x_20797 = x_20794 & x_20796;
assign x_20798 = x_20792 & x_20797;
assign x_20799 = x_20788 & x_20798;
assign x_20800 = x_9557 & x_9558;
assign x_20801 = x_9560 & x_9561;
assign x_20802 = x_9559 & x_20801;
assign x_20803 = x_20800 & x_20802;
assign x_20804 = x_9563 & x_9564;
assign x_20805 = x_9562 & x_20804;
assign x_20806 = x_9566 & x_9567;
assign x_20807 = x_9565 & x_20806;
assign x_20808 = x_20805 & x_20807;
assign x_20809 = x_20803 & x_20808;
assign x_20810 = x_9568 & x_9569;
assign x_20811 = x_9571 & x_9572;
assign x_20812 = x_9570 & x_20811;
assign x_20813 = x_20810 & x_20812;
assign x_20814 = x_9574 & x_9575;
assign x_20815 = x_9573 & x_20814;
assign x_20816 = x_9577 & x_9578;
assign x_20817 = x_9576 & x_20816;
assign x_20818 = x_20815 & x_20817;
assign x_20819 = x_20813 & x_20818;
assign x_20820 = x_20809 & x_20819;
assign x_20821 = x_20799 & x_20820;
assign x_20822 = x_20778 & x_20821;
assign x_20823 = x_9579 & x_9580;
assign x_20824 = x_9582 & x_9583;
assign x_20825 = x_9581 & x_20824;
assign x_20826 = x_20823 & x_20825;
assign x_20827 = x_9585 & x_9586;
assign x_20828 = x_9584 & x_20827;
assign x_20829 = x_9588 & x_9589;
assign x_20830 = x_9587 & x_20829;
assign x_20831 = x_20828 & x_20830;
assign x_20832 = x_20826 & x_20831;
assign x_20833 = x_9590 & x_9591;
assign x_20834 = x_9593 & x_9594;
assign x_20835 = x_9592 & x_20834;
assign x_20836 = x_20833 & x_20835;
assign x_20837 = x_9596 & x_9597;
assign x_20838 = x_9595 & x_20837;
assign x_20839 = x_9599 & x_9600;
assign x_20840 = x_9598 & x_20839;
assign x_20841 = x_20838 & x_20840;
assign x_20842 = x_20836 & x_20841;
assign x_20843 = x_20832 & x_20842;
assign x_20844 = x_9601 & x_9602;
assign x_20845 = x_9604 & x_9605;
assign x_20846 = x_9603 & x_20845;
assign x_20847 = x_20844 & x_20846;
assign x_20848 = x_9607 & x_9608;
assign x_20849 = x_9606 & x_20848;
assign x_20850 = x_9610 & x_9611;
assign x_20851 = x_9609 & x_20850;
assign x_20852 = x_20849 & x_20851;
assign x_20853 = x_20847 & x_20852;
assign x_20854 = x_9612 & x_9613;
assign x_20855 = x_9615 & x_9616;
assign x_20856 = x_9614 & x_20855;
assign x_20857 = x_20854 & x_20856;
assign x_20858 = x_9618 & x_9619;
assign x_20859 = x_9617 & x_20858;
assign x_20860 = x_9621 & x_9622;
assign x_20861 = x_9620 & x_20860;
assign x_20862 = x_20859 & x_20861;
assign x_20863 = x_20857 & x_20862;
assign x_20864 = x_20853 & x_20863;
assign x_20865 = x_20843 & x_20864;
assign x_20866 = x_9623 & x_9624;
assign x_20867 = x_9626 & x_9627;
assign x_20868 = x_9625 & x_20867;
assign x_20869 = x_20866 & x_20868;
assign x_20870 = x_9629 & x_9630;
assign x_20871 = x_9628 & x_20870;
assign x_20872 = x_9632 & x_9633;
assign x_20873 = x_9631 & x_20872;
assign x_20874 = x_20871 & x_20873;
assign x_20875 = x_20869 & x_20874;
assign x_20876 = x_9634 & x_9635;
assign x_20877 = x_9637 & x_9638;
assign x_20878 = x_9636 & x_20877;
assign x_20879 = x_20876 & x_20878;
assign x_20880 = x_9640 & x_9641;
assign x_20881 = x_9639 & x_20880;
assign x_20882 = x_9643 & x_9644;
assign x_20883 = x_9642 & x_20882;
assign x_20884 = x_20881 & x_20883;
assign x_20885 = x_20879 & x_20884;
assign x_20886 = x_20875 & x_20885;
assign x_20887 = x_9645 & x_9646;
assign x_20888 = x_9648 & x_9649;
assign x_20889 = x_9647 & x_20888;
assign x_20890 = x_20887 & x_20889;
assign x_20891 = x_9651 & x_9652;
assign x_20892 = x_9650 & x_20891;
assign x_20893 = x_9654 & x_9655;
assign x_20894 = x_9653 & x_20893;
assign x_20895 = x_20892 & x_20894;
assign x_20896 = x_20890 & x_20895;
assign x_20897 = x_9656 & x_9657;
assign x_20898 = x_9659 & x_9660;
assign x_20899 = x_9658 & x_20898;
assign x_20900 = x_20897 & x_20899;
assign x_20901 = x_9662 & x_9663;
assign x_20902 = x_9661 & x_20901;
assign x_20903 = x_9665 & x_9666;
assign x_20904 = x_9664 & x_20903;
assign x_20905 = x_20902 & x_20904;
assign x_20906 = x_20900 & x_20905;
assign x_20907 = x_20896 & x_20906;
assign x_20908 = x_20886 & x_20907;
assign x_20909 = x_20865 & x_20908;
assign x_20910 = x_20822 & x_20909;
assign x_20911 = x_9667 & x_9668;
assign x_20912 = x_9670 & x_9671;
assign x_20913 = x_9669 & x_20912;
assign x_20914 = x_20911 & x_20913;
assign x_20915 = x_9673 & x_9674;
assign x_20916 = x_9672 & x_20915;
assign x_20917 = x_9676 & x_9677;
assign x_20918 = x_9675 & x_20917;
assign x_20919 = x_20916 & x_20918;
assign x_20920 = x_20914 & x_20919;
assign x_20921 = x_9678 & x_9679;
assign x_20922 = x_9681 & x_9682;
assign x_20923 = x_9680 & x_20922;
assign x_20924 = x_20921 & x_20923;
assign x_20925 = x_9684 & x_9685;
assign x_20926 = x_9683 & x_20925;
assign x_20927 = x_9687 & x_9688;
assign x_20928 = x_9686 & x_20927;
assign x_20929 = x_20926 & x_20928;
assign x_20930 = x_20924 & x_20929;
assign x_20931 = x_20920 & x_20930;
assign x_20932 = x_9689 & x_9690;
assign x_20933 = x_9692 & x_9693;
assign x_20934 = x_9691 & x_20933;
assign x_20935 = x_20932 & x_20934;
assign x_20936 = x_9695 & x_9696;
assign x_20937 = x_9694 & x_20936;
assign x_20938 = x_9698 & x_9699;
assign x_20939 = x_9697 & x_20938;
assign x_20940 = x_20937 & x_20939;
assign x_20941 = x_20935 & x_20940;
assign x_20942 = x_9700 & x_9701;
assign x_20943 = x_9703 & x_9704;
assign x_20944 = x_9702 & x_20943;
assign x_20945 = x_20942 & x_20944;
assign x_20946 = x_9706 & x_9707;
assign x_20947 = x_9705 & x_20946;
assign x_20948 = x_9709 & x_9710;
assign x_20949 = x_9708 & x_20948;
assign x_20950 = x_20947 & x_20949;
assign x_20951 = x_20945 & x_20950;
assign x_20952 = x_20941 & x_20951;
assign x_20953 = x_20931 & x_20952;
assign x_20954 = x_9711 & x_9712;
assign x_20955 = x_9714 & x_9715;
assign x_20956 = x_9713 & x_20955;
assign x_20957 = x_20954 & x_20956;
assign x_20958 = x_9717 & x_9718;
assign x_20959 = x_9716 & x_20958;
assign x_20960 = x_9720 & x_9721;
assign x_20961 = x_9719 & x_20960;
assign x_20962 = x_20959 & x_20961;
assign x_20963 = x_20957 & x_20962;
assign x_20964 = x_9722 & x_9723;
assign x_20965 = x_9725 & x_9726;
assign x_20966 = x_9724 & x_20965;
assign x_20967 = x_20964 & x_20966;
assign x_20968 = x_9728 & x_9729;
assign x_20969 = x_9727 & x_20968;
assign x_20970 = x_9731 & x_9732;
assign x_20971 = x_9730 & x_20970;
assign x_20972 = x_20969 & x_20971;
assign x_20973 = x_20967 & x_20972;
assign x_20974 = x_20963 & x_20973;
assign x_20975 = x_9733 & x_9734;
assign x_20976 = x_9736 & x_9737;
assign x_20977 = x_9735 & x_20976;
assign x_20978 = x_20975 & x_20977;
assign x_20979 = x_9739 & x_9740;
assign x_20980 = x_9738 & x_20979;
assign x_20981 = x_9742 & x_9743;
assign x_20982 = x_9741 & x_20981;
assign x_20983 = x_20980 & x_20982;
assign x_20984 = x_20978 & x_20983;
assign x_20985 = x_9744 & x_9745;
assign x_20986 = x_9747 & x_9748;
assign x_20987 = x_9746 & x_20986;
assign x_20988 = x_20985 & x_20987;
assign x_20989 = x_9750 & x_9751;
assign x_20990 = x_9749 & x_20989;
assign x_20991 = x_9753 & x_9754;
assign x_20992 = x_9752 & x_20991;
assign x_20993 = x_20990 & x_20992;
assign x_20994 = x_20988 & x_20993;
assign x_20995 = x_20984 & x_20994;
assign x_20996 = x_20974 & x_20995;
assign x_20997 = x_20953 & x_20996;
assign x_20998 = x_9755 & x_9756;
assign x_20999 = x_9758 & x_9759;
assign x_21000 = x_9757 & x_20999;
assign x_21001 = x_20998 & x_21000;
assign x_21002 = x_9761 & x_9762;
assign x_21003 = x_9760 & x_21002;
assign x_21004 = x_9764 & x_9765;
assign x_21005 = x_9763 & x_21004;
assign x_21006 = x_21003 & x_21005;
assign x_21007 = x_21001 & x_21006;
assign x_21008 = x_9766 & x_9767;
assign x_21009 = x_9769 & x_9770;
assign x_21010 = x_9768 & x_21009;
assign x_21011 = x_21008 & x_21010;
assign x_21012 = x_9772 & x_9773;
assign x_21013 = x_9771 & x_21012;
assign x_21014 = x_9775 & x_9776;
assign x_21015 = x_9774 & x_21014;
assign x_21016 = x_21013 & x_21015;
assign x_21017 = x_21011 & x_21016;
assign x_21018 = x_21007 & x_21017;
assign x_21019 = x_9777 & x_9778;
assign x_21020 = x_9780 & x_9781;
assign x_21021 = x_9779 & x_21020;
assign x_21022 = x_21019 & x_21021;
assign x_21023 = x_9783 & x_9784;
assign x_21024 = x_9782 & x_21023;
assign x_21025 = x_9786 & x_9787;
assign x_21026 = x_9785 & x_21025;
assign x_21027 = x_21024 & x_21026;
assign x_21028 = x_21022 & x_21027;
assign x_21029 = x_9788 & x_9789;
assign x_21030 = x_9791 & x_9792;
assign x_21031 = x_9790 & x_21030;
assign x_21032 = x_21029 & x_21031;
assign x_21033 = x_9794 & x_9795;
assign x_21034 = x_9793 & x_21033;
assign x_21035 = x_9797 & x_9798;
assign x_21036 = x_9796 & x_21035;
assign x_21037 = x_21034 & x_21036;
assign x_21038 = x_21032 & x_21037;
assign x_21039 = x_21028 & x_21038;
assign x_21040 = x_21018 & x_21039;
assign x_21041 = x_9799 & x_9800;
assign x_21042 = x_9802 & x_9803;
assign x_21043 = x_9801 & x_21042;
assign x_21044 = x_21041 & x_21043;
assign x_21045 = x_9805 & x_9806;
assign x_21046 = x_9804 & x_21045;
assign x_21047 = x_9808 & x_9809;
assign x_21048 = x_9807 & x_21047;
assign x_21049 = x_21046 & x_21048;
assign x_21050 = x_21044 & x_21049;
assign x_21051 = x_9810 & x_9811;
assign x_21052 = x_9813 & x_9814;
assign x_21053 = x_9812 & x_21052;
assign x_21054 = x_21051 & x_21053;
assign x_21055 = x_9816 & x_9817;
assign x_21056 = x_9815 & x_21055;
assign x_21057 = x_9819 & x_9820;
assign x_21058 = x_9818 & x_21057;
assign x_21059 = x_21056 & x_21058;
assign x_21060 = x_21054 & x_21059;
assign x_21061 = x_21050 & x_21060;
assign x_21062 = x_9821 & x_9822;
assign x_21063 = x_9824 & x_9825;
assign x_21064 = x_9823 & x_21063;
assign x_21065 = x_21062 & x_21064;
assign x_21066 = x_9827 & x_9828;
assign x_21067 = x_9826 & x_21066;
assign x_21068 = x_9830 & x_9831;
assign x_21069 = x_9829 & x_21068;
assign x_21070 = x_21067 & x_21069;
assign x_21071 = x_21065 & x_21070;
assign x_21072 = x_9832 & x_9833;
assign x_21073 = x_9835 & x_9836;
assign x_21074 = x_9834 & x_21073;
assign x_21075 = x_21072 & x_21074;
assign x_21076 = x_9838 & x_9839;
assign x_21077 = x_9837 & x_21076;
assign x_21078 = x_9841 & x_9842;
assign x_21079 = x_9840 & x_21078;
assign x_21080 = x_21077 & x_21079;
assign x_21081 = x_21075 & x_21080;
assign x_21082 = x_21071 & x_21081;
assign x_21083 = x_21061 & x_21082;
assign x_21084 = x_21040 & x_21083;
assign x_21085 = x_20997 & x_21084;
assign x_21086 = x_20910 & x_21085;
assign x_21087 = x_20735 & x_21086;
assign x_21088 = x_20385 & x_21087;
assign x_21089 = x_9843 & x_9844;
assign x_21090 = x_9846 & x_9847;
assign x_21091 = x_9845 & x_21090;
assign x_21092 = x_21089 & x_21091;
assign x_21093 = x_9848 & x_9849;
assign x_21094 = x_9851 & x_9852;
assign x_21095 = x_9850 & x_21094;
assign x_21096 = x_21093 & x_21095;
assign x_21097 = x_21092 & x_21096;
assign x_21098 = x_9853 & x_9854;
assign x_21099 = x_9856 & x_9857;
assign x_21100 = x_9855 & x_21099;
assign x_21101 = x_21098 & x_21100;
assign x_21102 = x_9859 & x_9860;
assign x_21103 = x_9858 & x_21102;
assign x_21104 = x_9862 & x_9863;
assign x_21105 = x_9861 & x_21104;
assign x_21106 = x_21103 & x_21105;
assign x_21107 = x_21101 & x_21106;
assign x_21108 = x_21097 & x_21107;
assign x_21109 = x_9864 & x_9865;
assign x_21110 = x_9867 & x_9868;
assign x_21111 = x_9866 & x_21110;
assign x_21112 = x_21109 & x_21111;
assign x_21113 = x_9870 & x_9871;
assign x_21114 = x_9869 & x_21113;
assign x_21115 = x_9873 & x_9874;
assign x_21116 = x_9872 & x_21115;
assign x_21117 = x_21114 & x_21116;
assign x_21118 = x_21112 & x_21117;
assign x_21119 = x_9875 & x_9876;
assign x_21120 = x_9878 & x_9879;
assign x_21121 = x_9877 & x_21120;
assign x_21122 = x_21119 & x_21121;
assign x_21123 = x_9881 & x_9882;
assign x_21124 = x_9880 & x_21123;
assign x_21125 = x_9884 & x_9885;
assign x_21126 = x_9883 & x_21125;
assign x_21127 = x_21124 & x_21126;
assign x_21128 = x_21122 & x_21127;
assign x_21129 = x_21118 & x_21128;
assign x_21130 = x_21108 & x_21129;
assign x_21131 = x_9886 & x_9887;
assign x_21132 = x_9889 & x_9890;
assign x_21133 = x_9888 & x_21132;
assign x_21134 = x_21131 & x_21133;
assign x_21135 = x_9892 & x_9893;
assign x_21136 = x_9891 & x_21135;
assign x_21137 = x_9895 & x_9896;
assign x_21138 = x_9894 & x_21137;
assign x_21139 = x_21136 & x_21138;
assign x_21140 = x_21134 & x_21139;
assign x_21141 = x_9897 & x_9898;
assign x_21142 = x_9900 & x_9901;
assign x_21143 = x_9899 & x_21142;
assign x_21144 = x_21141 & x_21143;
assign x_21145 = x_9903 & x_9904;
assign x_21146 = x_9902 & x_21145;
assign x_21147 = x_9906 & x_9907;
assign x_21148 = x_9905 & x_21147;
assign x_21149 = x_21146 & x_21148;
assign x_21150 = x_21144 & x_21149;
assign x_21151 = x_21140 & x_21150;
assign x_21152 = x_9908 & x_9909;
assign x_21153 = x_9911 & x_9912;
assign x_21154 = x_9910 & x_21153;
assign x_21155 = x_21152 & x_21154;
assign x_21156 = x_9914 & x_9915;
assign x_21157 = x_9913 & x_21156;
assign x_21158 = x_9917 & x_9918;
assign x_21159 = x_9916 & x_21158;
assign x_21160 = x_21157 & x_21159;
assign x_21161 = x_21155 & x_21160;
assign x_21162 = x_9919 & x_9920;
assign x_21163 = x_9922 & x_9923;
assign x_21164 = x_9921 & x_21163;
assign x_21165 = x_21162 & x_21164;
assign x_21166 = x_9925 & x_9926;
assign x_21167 = x_9924 & x_21166;
assign x_21168 = x_9928 & x_9929;
assign x_21169 = x_9927 & x_21168;
assign x_21170 = x_21167 & x_21169;
assign x_21171 = x_21165 & x_21170;
assign x_21172 = x_21161 & x_21171;
assign x_21173 = x_21151 & x_21172;
assign x_21174 = x_21130 & x_21173;
assign x_21175 = x_9930 & x_9931;
assign x_21176 = x_9933 & x_9934;
assign x_21177 = x_9932 & x_21176;
assign x_21178 = x_21175 & x_21177;
assign x_21179 = x_9936 & x_9937;
assign x_21180 = x_9935 & x_21179;
assign x_21181 = x_9939 & x_9940;
assign x_21182 = x_9938 & x_21181;
assign x_21183 = x_21180 & x_21182;
assign x_21184 = x_21178 & x_21183;
assign x_21185 = x_9941 & x_9942;
assign x_21186 = x_9944 & x_9945;
assign x_21187 = x_9943 & x_21186;
assign x_21188 = x_21185 & x_21187;
assign x_21189 = x_9947 & x_9948;
assign x_21190 = x_9946 & x_21189;
assign x_21191 = x_9950 & x_9951;
assign x_21192 = x_9949 & x_21191;
assign x_21193 = x_21190 & x_21192;
assign x_21194 = x_21188 & x_21193;
assign x_21195 = x_21184 & x_21194;
assign x_21196 = x_9952 & x_9953;
assign x_21197 = x_9955 & x_9956;
assign x_21198 = x_9954 & x_21197;
assign x_21199 = x_21196 & x_21198;
assign x_21200 = x_9958 & x_9959;
assign x_21201 = x_9957 & x_21200;
assign x_21202 = x_9961 & x_9962;
assign x_21203 = x_9960 & x_21202;
assign x_21204 = x_21201 & x_21203;
assign x_21205 = x_21199 & x_21204;
assign x_21206 = x_9963 & x_9964;
assign x_21207 = x_9966 & x_9967;
assign x_21208 = x_9965 & x_21207;
assign x_21209 = x_21206 & x_21208;
assign x_21210 = x_9969 & x_9970;
assign x_21211 = x_9968 & x_21210;
assign x_21212 = x_9972 & x_9973;
assign x_21213 = x_9971 & x_21212;
assign x_21214 = x_21211 & x_21213;
assign x_21215 = x_21209 & x_21214;
assign x_21216 = x_21205 & x_21215;
assign x_21217 = x_21195 & x_21216;
assign x_21218 = x_9974 & x_9975;
assign x_21219 = x_9977 & x_9978;
assign x_21220 = x_9976 & x_21219;
assign x_21221 = x_21218 & x_21220;
assign x_21222 = x_9980 & x_9981;
assign x_21223 = x_9979 & x_21222;
assign x_21224 = x_9983 & x_9984;
assign x_21225 = x_9982 & x_21224;
assign x_21226 = x_21223 & x_21225;
assign x_21227 = x_21221 & x_21226;
assign x_21228 = x_9985 & x_9986;
assign x_21229 = x_9988 & x_9989;
assign x_21230 = x_9987 & x_21229;
assign x_21231 = x_21228 & x_21230;
assign x_21232 = x_9991 & x_9992;
assign x_21233 = x_9990 & x_21232;
assign x_21234 = x_9994 & x_9995;
assign x_21235 = x_9993 & x_21234;
assign x_21236 = x_21233 & x_21235;
assign x_21237 = x_21231 & x_21236;
assign x_21238 = x_21227 & x_21237;
assign x_21239 = x_9996 & x_9997;
assign x_21240 = x_9999 & x_10000;
assign x_21241 = x_9998 & x_21240;
assign x_21242 = x_21239 & x_21241;
assign x_21243 = x_10002 & x_10003;
assign x_21244 = x_10001 & x_21243;
assign x_21245 = x_10005 & x_10006;
assign x_21246 = x_10004 & x_21245;
assign x_21247 = x_21244 & x_21246;
assign x_21248 = x_21242 & x_21247;
assign x_21249 = x_10007 & x_10008;
assign x_21250 = x_10010 & x_10011;
assign x_21251 = x_10009 & x_21250;
assign x_21252 = x_21249 & x_21251;
assign x_21253 = x_10013 & x_10014;
assign x_21254 = x_10012 & x_21253;
assign x_21255 = x_10016 & x_10017;
assign x_21256 = x_10015 & x_21255;
assign x_21257 = x_21254 & x_21256;
assign x_21258 = x_21252 & x_21257;
assign x_21259 = x_21248 & x_21258;
assign x_21260 = x_21238 & x_21259;
assign x_21261 = x_21217 & x_21260;
assign x_21262 = x_21174 & x_21261;
assign x_21263 = x_10018 & x_10019;
assign x_21264 = x_10021 & x_10022;
assign x_21265 = x_10020 & x_21264;
assign x_21266 = x_21263 & x_21265;
assign x_21267 = x_10024 & x_10025;
assign x_21268 = x_10023 & x_21267;
assign x_21269 = x_10027 & x_10028;
assign x_21270 = x_10026 & x_21269;
assign x_21271 = x_21268 & x_21270;
assign x_21272 = x_21266 & x_21271;
assign x_21273 = x_10029 & x_10030;
assign x_21274 = x_10032 & x_10033;
assign x_21275 = x_10031 & x_21274;
assign x_21276 = x_21273 & x_21275;
assign x_21277 = x_10035 & x_10036;
assign x_21278 = x_10034 & x_21277;
assign x_21279 = x_10038 & x_10039;
assign x_21280 = x_10037 & x_21279;
assign x_21281 = x_21278 & x_21280;
assign x_21282 = x_21276 & x_21281;
assign x_21283 = x_21272 & x_21282;
assign x_21284 = x_10040 & x_10041;
assign x_21285 = x_10043 & x_10044;
assign x_21286 = x_10042 & x_21285;
assign x_21287 = x_21284 & x_21286;
assign x_21288 = x_10046 & x_10047;
assign x_21289 = x_10045 & x_21288;
assign x_21290 = x_10049 & x_10050;
assign x_21291 = x_10048 & x_21290;
assign x_21292 = x_21289 & x_21291;
assign x_21293 = x_21287 & x_21292;
assign x_21294 = x_10051 & x_10052;
assign x_21295 = x_10054 & x_10055;
assign x_21296 = x_10053 & x_21295;
assign x_21297 = x_21294 & x_21296;
assign x_21298 = x_10057 & x_10058;
assign x_21299 = x_10056 & x_21298;
assign x_21300 = x_10060 & x_10061;
assign x_21301 = x_10059 & x_21300;
assign x_21302 = x_21299 & x_21301;
assign x_21303 = x_21297 & x_21302;
assign x_21304 = x_21293 & x_21303;
assign x_21305 = x_21283 & x_21304;
assign x_21306 = x_10062 & x_10063;
assign x_21307 = x_10065 & x_10066;
assign x_21308 = x_10064 & x_21307;
assign x_21309 = x_21306 & x_21308;
assign x_21310 = x_10068 & x_10069;
assign x_21311 = x_10067 & x_21310;
assign x_21312 = x_10071 & x_10072;
assign x_21313 = x_10070 & x_21312;
assign x_21314 = x_21311 & x_21313;
assign x_21315 = x_21309 & x_21314;
assign x_21316 = x_10073 & x_10074;
assign x_21317 = x_10076 & x_10077;
assign x_21318 = x_10075 & x_21317;
assign x_21319 = x_21316 & x_21318;
assign x_21320 = x_10079 & x_10080;
assign x_21321 = x_10078 & x_21320;
assign x_21322 = x_10082 & x_10083;
assign x_21323 = x_10081 & x_21322;
assign x_21324 = x_21321 & x_21323;
assign x_21325 = x_21319 & x_21324;
assign x_21326 = x_21315 & x_21325;
assign x_21327 = x_10084 & x_10085;
assign x_21328 = x_10087 & x_10088;
assign x_21329 = x_10086 & x_21328;
assign x_21330 = x_21327 & x_21329;
assign x_21331 = x_10090 & x_10091;
assign x_21332 = x_10089 & x_21331;
assign x_21333 = x_10093 & x_10094;
assign x_21334 = x_10092 & x_21333;
assign x_21335 = x_21332 & x_21334;
assign x_21336 = x_21330 & x_21335;
assign x_21337 = x_10095 & x_10096;
assign x_21338 = x_10098 & x_10099;
assign x_21339 = x_10097 & x_21338;
assign x_21340 = x_21337 & x_21339;
assign x_21341 = x_10101 & x_10102;
assign x_21342 = x_10100 & x_21341;
assign x_21343 = x_10104 & x_10105;
assign x_21344 = x_10103 & x_21343;
assign x_21345 = x_21342 & x_21344;
assign x_21346 = x_21340 & x_21345;
assign x_21347 = x_21336 & x_21346;
assign x_21348 = x_21326 & x_21347;
assign x_21349 = x_21305 & x_21348;
assign x_21350 = x_10106 & x_10107;
assign x_21351 = x_10109 & x_10110;
assign x_21352 = x_10108 & x_21351;
assign x_21353 = x_21350 & x_21352;
assign x_21354 = x_10112 & x_10113;
assign x_21355 = x_10111 & x_21354;
assign x_21356 = x_10115 & x_10116;
assign x_21357 = x_10114 & x_21356;
assign x_21358 = x_21355 & x_21357;
assign x_21359 = x_21353 & x_21358;
assign x_21360 = x_10117 & x_10118;
assign x_21361 = x_10120 & x_10121;
assign x_21362 = x_10119 & x_21361;
assign x_21363 = x_21360 & x_21362;
assign x_21364 = x_10123 & x_10124;
assign x_21365 = x_10122 & x_21364;
assign x_21366 = x_10126 & x_10127;
assign x_21367 = x_10125 & x_21366;
assign x_21368 = x_21365 & x_21367;
assign x_21369 = x_21363 & x_21368;
assign x_21370 = x_21359 & x_21369;
assign x_21371 = x_10128 & x_10129;
assign x_21372 = x_10131 & x_10132;
assign x_21373 = x_10130 & x_21372;
assign x_21374 = x_21371 & x_21373;
assign x_21375 = x_10134 & x_10135;
assign x_21376 = x_10133 & x_21375;
assign x_21377 = x_10137 & x_10138;
assign x_21378 = x_10136 & x_21377;
assign x_21379 = x_21376 & x_21378;
assign x_21380 = x_21374 & x_21379;
assign x_21381 = x_10139 & x_10140;
assign x_21382 = x_10142 & x_10143;
assign x_21383 = x_10141 & x_21382;
assign x_21384 = x_21381 & x_21383;
assign x_21385 = x_10145 & x_10146;
assign x_21386 = x_10144 & x_21385;
assign x_21387 = x_10148 & x_10149;
assign x_21388 = x_10147 & x_21387;
assign x_21389 = x_21386 & x_21388;
assign x_21390 = x_21384 & x_21389;
assign x_21391 = x_21380 & x_21390;
assign x_21392 = x_21370 & x_21391;
assign x_21393 = x_10150 & x_10151;
assign x_21394 = x_10153 & x_10154;
assign x_21395 = x_10152 & x_21394;
assign x_21396 = x_21393 & x_21395;
assign x_21397 = x_10156 & x_10157;
assign x_21398 = x_10155 & x_21397;
assign x_21399 = x_10159 & x_10160;
assign x_21400 = x_10158 & x_21399;
assign x_21401 = x_21398 & x_21400;
assign x_21402 = x_21396 & x_21401;
assign x_21403 = x_10161 & x_10162;
assign x_21404 = x_10164 & x_10165;
assign x_21405 = x_10163 & x_21404;
assign x_21406 = x_21403 & x_21405;
assign x_21407 = x_10167 & x_10168;
assign x_21408 = x_10166 & x_21407;
assign x_21409 = x_10170 & x_10171;
assign x_21410 = x_10169 & x_21409;
assign x_21411 = x_21408 & x_21410;
assign x_21412 = x_21406 & x_21411;
assign x_21413 = x_21402 & x_21412;
assign x_21414 = x_10172 & x_10173;
assign x_21415 = x_10175 & x_10176;
assign x_21416 = x_10174 & x_21415;
assign x_21417 = x_21414 & x_21416;
assign x_21418 = x_10178 & x_10179;
assign x_21419 = x_10177 & x_21418;
assign x_21420 = x_10181 & x_10182;
assign x_21421 = x_10180 & x_21420;
assign x_21422 = x_21419 & x_21421;
assign x_21423 = x_21417 & x_21422;
assign x_21424 = x_10183 & x_10184;
assign x_21425 = x_10186 & x_10187;
assign x_21426 = x_10185 & x_21425;
assign x_21427 = x_21424 & x_21426;
assign x_21428 = x_10189 & x_10190;
assign x_21429 = x_10188 & x_21428;
assign x_21430 = x_10192 & x_10193;
assign x_21431 = x_10191 & x_21430;
assign x_21432 = x_21429 & x_21431;
assign x_21433 = x_21427 & x_21432;
assign x_21434 = x_21423 & x_21433;
assign x_21435 = x_21413 & x_21434;
assign x_21436 = x_21392 & x_21435;
assign x_21437 = x_21349 & x_21436;
assign x_21438 = x_21262 & x_21437;
assign x_21439 = x_10194 & x_10195;
assign x_21440 = x_10197 & x_10198;
assign x_21441 = x_10196 & x_21440;
assign x_21442 = x_21439 & x_21441;
assign x_21443 = x_10200 & x_10201;
assign x_21444 = x_10199 & x_21443;
assign x_21445 = x_10203 & x_10204;
assign x_21446 = x_10202 & x_21445;
assign x_21447 = x_21444 & x_21446;
assign x_21448 = x_21442 & x_21447;
assign x_21449 = x_10205 & x_10206;
assign x_21450 = x_10208 & x_10209;
assign x_21451 = x_10207 & x_21450;
assign x_21452 = x_21449 & x_21451;
assign x_21453 = x_10211 & x_10212;
assign x_21454 = x_10210 & x_21453;
assign x_21455 = x_10214 & x_10215;
assign x_21456 = x_10213 & x_21455;
assign x_21457 = x_21454 & x_21456;
assign x_21458 = x_21452 & x_21457;
assign x_21459 = x_21448 & x_21458;
assign x_21460 = x_10216 & x_10217;
assign x_21461 = x_10219 & x_10220;
assign x_21462 = x_10218 & x_21461;
assign x_21463 = x_21460 & x_21462;
assign x_21464 = x_10222 & x_10223;
assign x_21465 = x_10221 & x_21464;
assign x_21466 = x_10225 & x_10226;
assign x_21467 = x_10224 & x_21466;
assign x_21468 = x_21465 & x_21467;
assign x_21469 = x_21463 & x_21468;
assign x_21470 = x_10227 & x_10228;
assign x_21471 = x_10230 & x_10231;
assign x_21472 = x_10229 & x_21471;
assign x_21473 = x_21470 & x_21472;
assign x_21474 = x_10233 & x_10234;
assign x_21475 = x_10232 & x_21474;
assign x_21476 = x_10236 & x_10237;
assign x_21477 = x_10235 & x_21476;
assign x_21478 = x_21475 & x_21477;
assign x_21479 = x_21473 & x_21478;
assign x_21480 = x_21469 & x_21479;
assign x_21481 = x_21459 & x_21480;
assign x_21482 = x_10238 & x_10239;
assign x_21483 = x_10241 & x_10242;
assign x_21484 = x_10240 & x_21483;
assign x_21485 = x_21482 & x_21484;
assign x_21486 = x_10244 & x_10245;
assign x_21487 = x_10243 & x_21486;
assign x_21488 = x_10247 & x_10248;
assign x_21489 = x_10246 & x_21488;
assign x_21490 = x_21487 & x_21489;
assign x_21491 = x_21485 & x_21490;
assign x_21492 = x_10249 & x_10250;
assign x_21493 = x_10252 & x_10253;
assign x_21494 = x_10251 & x_21493;
assign x_21495 = x_21492 & x_21494;
assign x_21496 = x_10255 & x_10256;
assign x_21497 = x_10254 & x_21496;
assign x_21498 = x_10258 & x_10259;
assign x_21499 = x_10257 & x_21498;
assign x_21500 = x_21497 & x_21499;
assign x_21501 = x_21495 & x_21500;
assign x_21502 = x_21491 & x_21501;
assign x_21503 = x_10260 & x_10261;
assign x_21504 = x_10263 & x_10264;
assign x_21505 = x_10262 & x_21504;
assign x_21506 = x_21503 & x_21505;
assign x_21507 = x_10266 & x_10267;
assign x_21508 = x_10265 & x_21507;
assign x_21509 = x_10269 & x_10270;
assign x_21510 = x_10268 & x_21509;
assign x_21511 = x_21508 & x_21510;
assign x_21512 = x_21506 & x_21511;
assign x_21513 = x_10271 & x_10272;
assign x_21514 = x_10274 & x_10275;
assign x_21515 = x_10273 & x_21514;
assign x_21516 = x_21513 & x_21515;
assign x_21517 = x_10277 & x_10278;
assign x_21518 = x_10276 & x_21517;
assign x_21519 = x_10280 & x_10281;
assign x_21520 = x_10279 & x_21519;
assign x_21521 = x_21518 & x_21520;
assign x_21522 = x_21516 & x_21521;
assign x_21523 = x_21512 & x_21522;
assign x_21524 = x_21502 & x_21523;
assign x_21525 = x_21481 & x_21524;
assign x_21526 = x_10282 & x_10283;
assign x_21527 = x_10285 & x_10286;
assign x_21528 = x_10284 & x_21527;
assign x_21529 = x_21526 & x_21528;
assign x_21530 = x_10288 & x_10289;
assign x_21531 = x_10287 & x_21530;
assign x_21532 = x_10291 & x_10292;
assign x_21533 = x_10290 & x_21532;
assign x_21534 = x_21531 & x_21533;
assign x_21535 = x_21529 & x_21534;
assign x_21536 = x_10293 & x_10294;
assign x_21537 = x_10296 & x_10297;
assign x_21538 = x_10295 & x_21537;
assign x_21539 = x_21536 & x_21538;
assign x_21540 = x_10299 & x_10300;
assign x_21541 = x_10298 & x_21540;
assign x_21542 = x_10302 & x_10303;
assign x_21543 = x_10301 & x_21542;
assign x_21544 = x_21541 & x_21543;
assign x_21545 = x_21539 & x_21544;
assign x_21546 = x_21535 & x_21545;
assign x_21547 = x_10304 & x_10305;
assign x_21548 = x_10307 & x_10308;
assign x_21549 = x_10306 & x_21548;
assign x_21550 = x_21547 & x_21549;
assign x_21551 = x_10310 & x_10311;
assign x_21552 = x_10309 & x_21551;
assign x_21553 = x_10313 & x_10314;
assign x_21554 = x_10312 & x_21553;
assign x_21555 = x_21552 & x_21554;
assign x_21556 = x_21550 & x_21555;
assign x_21557 = x_10315 & x_10316;
assign x_21558 = x_10318 & x_10319;
assign x_21559 = x_10317 & x_21558;
assign x_21560 = x_21557 & x_21559;
assign x_21561 = x_10321 & x_10322;
assign x_21562 = x_10320 & x_21561;
assign x_21563 = x_10324 & x_10325;
assign x_21564 = x_10323 & x_21563;
assign x_21565 = x_21562 & x_21564;
assign x_21566 = x_21560 & x_21565;
assign x_21567 = x_21556 & x_21566;
assign x_21568 = x_21546 & x_21567;
assign x_21569 = x_10326 & x_10327;
assign x_21570 = x_10329 & x_10330;
assign x_21571 = x_10328 & x_21570;
assign x_21572 = x_21569 & x_21571;
assign x_21573 = x_10332 & x_10333;
assign x_21574 = x_10331 & x_21573;
assign x_21575 = x_10335 & x_10336;
assign x_21576 = x_10334 & x_21575;
assign x_21577 = x_21574 & x_21576;
assign x_21578 = x_21572 & x_21577;
assign x_21579 = x_10337 & x_10338;
assign x_21580 = x_10340 & x_10341;
assign x_21581 = x_10339 & x_21580;
assign x_21582 = x_21579 & x_21581;
assign x_21583 = x_10343 & x_10344;
assign x_21584 = x_10342 & x_21583;
assign x_21585 = x_10346 & x_10347;
assign x_21586 = x_10345 & x_21585;
assign x_21587 = x_21584 & x_21586;
assign x_21588 = x_21582 & x_21587;
assign x_21589 = x_21578 & x_21588;
assign x_21590 = x_10348 & x_10349;
assign x_21591 = x_10351 & x_10352;
assign x_21592 = x_10350 & x_21591;
assign x_21593 = x_21590 & x_21592;
assign x_21594 = x_10354 & x_10355;
assign x_21595 = x_10353 & x_21594;
assign x_21596 = x_10357 & x_10358;
assign x_21597 = x_10356 & x_21596;
assign x_21598 = x_21595 & x_21597;
assign x_21599 = x_21593 & x_21598;
assign x_21600 = x_10359 & x_10360;
assign x_21601 = x_10362 & x_10363;
assign x_21602 = x_10361 & x_21601;
assign x_21603 = x_21600 & x_21602;
assign x_21604 = x_10365 & x_10366;
assign x_21605 = x_10364 & x_21604;
assign x_21606 = x_10368 & x_10369;
assign x_21607 = x_10367 & x_21606;
assign x_21608 = x_21605 & x_21607;
assign x_21609 = x_21603 & x_21608;
assign x_21610 = x_21599 & x_21609;
assign x_21611 = x_21589 & x_21610;
assign x_21612 = x_21568 & x_21611;
assign x_21613 = x_21525 & x_21612;
assign x_21614 = x_10370 & x_10371;
assign x_21615 = x_10373 & x_10374;
assign x_21616 = x_10372 & x_21615;
assign x_21617 = x_21614 & x_21616;
assign x_21618 = x_10376 & x_10377;
assign x_21619 = x_10375 & x_21618;
assign x_21620 = x_10379 & x_10380;
assign x_21621 = x_10378 & x_21620;
assign x_21622 = x_21619 & x_21621;
assign x_21623 = x_21617 & x_21622;
assign x_21624 = x_10381 & x_10382;
assign x_21625 = x_10384 & x_10385;
assign x_21626 = x_10383 & x_21625;
assign x_21627 = x_21624 & x_21626;
assign x_21628 = x_10387 & x_10388;
assign x_21629 = x_10386 & x_21628;
assign x_21630 = x_10390 & x_10391;
assign x_21631 = x_10389 & x_21630;
assign x_21632 = x_21629 & x_21631;
assign x_21633 = x_21627 & x_21632;
assign x_21634 = x_21623 & x_21633;
assign x_21635 = x_10392 & x_10393;
assign x_21636 = x_10395 & x_10396;
assign x_21637 = x_10394 & x_21636;
assign x_21638 = x_21635 & x_21637;
assign x_21639 = x_10398 & x_10399;
assign x_21640 = x_10397 & x_21639;
assign x_21641 = x_10401 & x_10402;
assign x_21642 = x_10400 & x_21641;
assign x_21643 = x_21640 & x_21642;
assign x_21644 = x_21638 & x_21643;
assign x_21645 = x_10403 & x_10404;
assign x_21646 = x_10406 & x_10407;
assign x_21647 = x_10405 & x_21646;
assign x_21648 = x_21645 & x_21647;
assign x_21649 = x_10409 & x_10410;
assign x_21650 = x_10408 & x_21649;
assign x_21651 = x_10412 & x_10413;
assign x_21652 = x_10411 & x_21651;
assign x_21653 = x_21650 & x_21652;
assign x_21654 = x_21648 & x_21653;
assign x_21655 = x_21644 & x_21654;
assign x_21656 = x_21634 & x_21655;
assign x_21657 = x_10414 & x_10415;
assign x_21658 = x_10417 & x_10418;
assign x_21659 = x_10416 & x_21658;
assign x_21660 = x_21657 & x_21659;
assign x_21661 = x_10420 & x_10421;
assign x_21662 = x_10419 & x_21661;
assign x_21663 = x_10423 & x_10424;
assign x_21664 = x_10422 & x_21663;
assign x_21665 = x_21662 & x_21664;
assign x_21666 = x_21660 & x_21665;
assign x_21667 = x_10425 & x_10426;
assign x_21668 = x_10428 & x_10429;
assign x_21669 = x_10427 & x_21668;
assign x_21670 = x_21667 & x_21669;
assign x_21671 = x_10431 & x_10432;
assign x_21672 = x_10430 & x_21671;
assign x_21673 = x_10434 & x_10435;
assign x_21674 = x_10433 & x_21673;
assign x_21675 = x_21672 & x_21674;
assign x_21676 = x_21670 & x_21675;
assign x_21677 = x_21666 & x_21676;
assign x_21678 = x_10436 & x_10437;
assign x_21679 = x_10439 & x_10440;
assign x_21680 = x_10438 & x_21679;
assign x_21681 = x_21678 & x_21680;
assign x_21682 = x_10442 & x_10443;
assign x_21683 = x_10441 & x_21682;
assign x_21684 = x_10445 & x_10446;
assign x_21685 = x_10444 & x_21684;
assign x_21686 = x_21683 & x_21685;
assign x_21687 = x_21681 & x_21686;
assign x_21688 = x_10447 & x_10448;
assign x_21689 = x_10450 & x_10451;
assign x_21690 = x_10449 & x_21689;
assign x_21691 = x_21688 & x_21690;
assign x_21692 = x_10453 & x_10454;
assign x_21693 = x_10452 & x_21692;
assign x_21694 = x_10456 & x_10457;
assign x_21695 = x_10455 & x_21694;
assign x_21696 = x_21693 & x_21695;
assign x_21697 = x_21691 & x_21696;
assign x_21698 = x_21687 & x_21697;
assign x_21699 = x_21677 & x_21698;
assign x_21700 = x_21656 & x_21699;
assign x_21701 = x_10458 & x_10459;
assign x_21702 = x_10461 & x_10462;
assign x_21703 = x_10460 & x_21702;
assign x_21704 = x_21701 & x_21703;
assign x_21705 = x_10464 & x_10465;
assign x_21706 = x_10463 & x_21705;
assign x_21707 = x_10467 & x_10468;
assign x_21708 = x_10466 & x_21707;
assign x_21709 = x_21706 & x_21708;
assign x_21710 = x_21704 & x_21709;
assign x_21711 = x_10469 & x_10470;
assign x_21712 = x_10472 & x_10473;
assign x_21713 = x_10471 & x_21712;
assign x_21714 = x_21711 & x_21713;
assign x_21715 = x_10475 & x_10476;
assign x_21716 = x_10474 & x_21715;
assign x_21717 = x_10478 & x_10479;
assign x_21718 = x_10477 & x_21717;
assign x_21719 = x_21716 & x_21718;
assign x_21720 = x_21714 & x_21719;
assign x_21721 = x_21710 & x_21720;
assign x_21722 = x_10480 & x_10481;
assign x_21723 = x_10483 & x_10484;
assign x_21724 = x_10482 & x_21723;
assign x_21725 = x_21722 & x_21724;
assign x_21726 = x_10486 & x_10487;
assign x_21727 = x_10485 & x_21726;
assign x_21728 = x_10489 & x_10490;
assign x_21729 = x_10488 & x_21728;
assign x_21730 = x_21727 & x_21729;
assign x_21731 = x_21725 & x_21730;
assign x_21732 = x_10491 & x_10492;
assign x_21733 = x_10494 & x_10495;
assign x_21734 = x_10493 & x_21733;
assign x_21735 = x_21732 & x_21734;
assign x_21736 = x_10497 & x_10498;
assign x_21737 = x_10496 & x_21736;
assign x_21738 = x_10500 & x_10501;
assign x_21739 = x_10499 & x_21738;
assign x_21740 = x_21737 & x_21739;
assign x_21741 = x_21735 & x_21740;
assign x_21742 = x_21731 & x_21741;
assign x_21743 = x_21721 & x_21742;
assign x_21744 = x_10502 & x_10503;
assign x_21745 = x_10505 & x_10506;
assign x_21746 = x_10504 & x_21745;
assign x_21747 = x_21744 & x_21746;
assign x_21748 = x_10508 & x_10509;
assign x_21749 = x_10507 & x_21748;
assign x_21750 = x_10511 & x_10512;
assign x_21751 = x_10510 & x_21750;
assign x_21752 = x_21749 & x_21751;
assign x_21753 = x_21747 & x_21752;
assign x_21754 = x_10513 & x_10514;
assign x_21755 = x_10516 & x_10517;
assign x_21756 = x_10515 & x_21755;
assign x_21757 = x_21754 & x_21756;
assign x_21758 = x_10519 & x_10520;
assign x_21759 = x_10518 & x_21758;
assign x_21760 = x_10522 & x_10523;
assign x_21761 = x_10521 & x_21760;
assign x_21762 = x_21759 & x_21761;
assign x_21763 = x_21757 & x_21762;
assign x_21764 = x_21753 & x_21763;
assign x_21765 = x_10524 & x_10525;
assign x_21766 = x_10527 & x_10528;
assign x_21767 = x_10526 & x_21766;
assign x_21768 = x_21765 & x_21767;
assign x_21769 = x_10530 & x_10531;
assign x_21770 = x_10529 & x_21769;
assign x_21771 = x_10533 & x_10534;
assign x_21772 = x_10532 & x_21771;
assign x_21773 = x_21770 & x_21772;
assign x_21774 = x_21768 & x_21773;
assign x_21775 = x_10535 & x_10536;
assign x_21776 = x_10538 & x_10539;
assign x_21777 = x_10537 & x_21776;
assign x_21778 = x_21775 & x_21777;
assign x_21779 = x_10541 & x_10542;
assign x_21780 = x_10540 & x_21779;
assign x_21781 = x_10544 & x_10545;
assign x_21782 = x_10543 & x_21781;
assign x_21783 = x_21780 & x_21782;
assign x_21784 = x_21778 & x_21783;
assign x_21785 = x_21774 & x_21784;
assign x_21786 = x_21764 & x_21785;
assign x_21787 = x_21743 & x_21786;
assign x_21788 = x_21700 & x_21787;
assign x_21789 = x_21613 & x_21788;
assign x_21790 = x_21438 & x_21789;
assign x_21791 = x_10546 & x_10547;
assign x_21792 = x_10549 & x_10550;
assign x_21793 = x_10548 & x_21792;
assign x_21794 = x_21791 & x_21793;
assign x_21795 = x_10552 & x_10553;
assign x_21796 = x_10551 & x_21795;
assign x_21797 = x_10555 & x_10556;
assign x_21798 = x_10554 & x_21797;
assign x_21799 = x_21796 & x_21798;
assign x_21800 = x_21794 & x_21799;
assign x_21801 = x_10557 & x_10558;
assign x_21802 = x_10560 & x_10561;
assign x_21803 = x_10559 & x_21802;
assign x_21804 = x_21801 & x_21803;
assign x_21805 = x_10563 & x_10564;
assign x_21806 = x_10562 & x_21805;
assign x_21807 = x_10566 & x_10567;
assign x_21808 = x_10565 & x_21807;
assign x_21809 = x_21806 & x_21808;
assign x_21810 = x_21804 & x_21809;
assign x_21811 = x_21800 & x_21810;
assign x_21812 = x_10568 & x_10569;
assign x_21813 = x_10571 & x_10572;
assign x_21814 = x_10570 & x_21813;
assign x_21815 = x_21812 & x_21814;
assign x_21816 = x_10574 & x_10575;
assign x_21817 = x_10573 & x_21816;
assign x_21818 = x_10577 & x_10578;
assign x_21819 = x_10576 & x_21818;
assign x_21820 = x_21817 & x_21819;
assign x_21821 = x_21815 & x_21820;
assign x_21822 = x_10579 & x_10580;
assign x_21823 = x_10582 & x_10583;
assign x_21824 = x_10581 & x_21823;
assign x_21825 = x_21822 & x_21824;
assign x_21826 = x_10585 & x_10586;
assign x_21827 = x_10584 & x_21826;
assign x_21828 = x_10588 & x_10589;
assign x_21829 = x_10587 & x_21828;
assign x_21830 = x_21827 & x_21829;
assign x_21831 = x_21825 & x_21830;
assign x_21832 = x_21821 & x_21831;
assign x_21833 = x_21811 & x_21832;
assign x_21834 = x_10590 & x_10591;
assign x_21835 = x_10593 & x_10594;
assign x_21836 = x_10592 & x_21835;
assign x_21837 = x_21834 & x_21836;
assign x_21838 = x_10596 & x_10597;
assign x_21839 = x_10595 & x_21838;
assign x_21840 = x_10599 & x_10600;
assign x_21841 = x_10598 & x_21840;
assign x_21842 = x_21839 & x_21841;
assign x_21843 = x_21837 & x_21842;
assign x_21844 = x_10601 & x_10602;
assign x_21845 = x_10604 & x_10605;
assign x_21846 = x_10603 & x_21845;
assign x_21847 = x_21844 & x_21846;
assign x_21848 = x_10607 & x_10608;
assign x_21849 = x_10606 & x_21848;
assign x_21850 = x_10610 & x_10611;
assign x_21851 = x_10609 & x_21850;
assign x_21852 = x_21849 & x_21851;
assign x_21853 = x_21847 & x_21852;
assign x_21854 = x_21843 & x_21853;
assign x_21855 = x_10612 & x_10613;
assign x_21856 = x_10615 & x_10616;
assign x_21857 = x_10614 & x_21856;
assign x_21858 = x_21855 & x_21857;
assign x_21859 = x_10618 & x_10619;
assign x_21860 = x_10617 & x_21859;
assign x_21861 = x_10621 & x_10622;
assign x_21862 = x_10620 & x_21861;
assign x_21863 = x_21860 & x_21862;
assign x_21864 = x_21858 & x_21863;
assign x_21865 = x_10623 & x_10624;
assign x_21866 = x_10626 & x_10627;
assign x_21867 = x_10625 & x_21866;
assign x_21868 = x_21865 & x_21867;
assign x_21869 = x_10629 & x_10630;
assign x_21870 = x_10628 & x_21869;
assign x_21871 = x_10632 & x_10633;
assign x_21872 = x_10631 & x_21871;
assign x_21873 = x_21870 & x_21872;
assign x_21874 = x_21868 & x_21873;
assign x_21875 = x_21864 & x_21874;
assign x_21876 = x_21854 & x_21875;
assign x_21877 = x_21833 & x_21876;
assign x_21878 = x_10634 & x_10635;
assign x_21879 = x_10637 & x_10638;
assign x_21880 = x_10636 & x_21879;
assign x_21881 = x_21878 & x_21880;
assign x_21882 = x_10640 & x_10641;
assign x_21883 = x_10639 & x_21882;
assign x_21884 = x_10643 & x_10644;
assign x_21885 = x_10642 & x_21884;
assign x_21886 = x_21883 & x_21885;
assign x_21887 = x_21881 & x_21886;
assign x_21888 = x_10645 & x_10646;
assign x_21889 = x_10648 & x_10649;
assign x_21890 = x_10647 & x_21889;
assign x_21891 = x_21888 & x_21890;
assign x_21892 = x_10651 & x_10652;
assign x_21893 = x_10650 & x_21892;
assign x_21894 = x_10654 & x_10655;
assign x_21895 = x_10653 & x_21894;
assign x_21896 = x_21893 & x_21895;
assign x_21897 = x_21891 & x_21896;
assign x_21898 = x_21887 & x_21897;
assign x_21899 = x_10656 & x_10657;
assign x_21900 = x_10659 & x_10660;
assign x_21901 = x_10658 & x_21900;
assign x_21902 = x_21899 & x_21901;
assign x_21903 = x_10662 & x_10663;
assign x_21904 = x_10661 & x_21903;
assign x_21905 = x_10665 & x_10666;
assign x_21906 = x_10664 & x_21905;
assign x_21907 = x_21904 & x_21906;
assign x_21908 = x_21902 & x_21907;
assign x_21909 = x_10667 & x_10668;
assign x_21910 = x_10670 & x_10671;
assign x_21911 = x_10669 & x_21910;
assign x_21912 = x_21909 & x_21911;
assign x_21913 = x_10673 & x_10674;
assign x_21914 = x_10672 & x_21913;
assign x_21915 = x_10676 & x_10677;
assign x_21916 = x_10675 & x_21915;
assign x_21917 = x_21914 & x_21916;
assign x_21918 = x_21912 & x_21917;
assign x_21919 = x_21908 & x_21918;
assign x_21920 = x_21898 & x_21919;
assign x_21921 = x_10678 & x_10679;
assign x_21922 = x_10681 & x_10682;
assign x_21923 = x_10680 & x_21922;
assign x_21924 = x_21921 & x_21923;
assign x_21925 = x_10684 & x_10685;
assign x_21926 = x_10683 & x_21925;
assign x_21927 = x_10687 & x_10688;
assign x_21928 = x_10686 & x_21927;
assign x_21929 = x_21926 & x_21928;
assign x_21930 = x_21924 & x_21929;
assign x_21931 = x_10689 & x_10690;
assign x_21932 = x_10692 & x_10693;
assign x_21933 = x_10691 & x_21932;
assign x_21934 = x_21931 & x_21933;
assign x_21935 = x_10695 & x_10696;
assign x_21936 = x_10694 & x_21935;
assign x_21937 = x_10698 & x_10699;
assign x_21938 = x_10697 & x_21937;
assign x_21939 = x_21936 & x_21938;
assign x_21940 = x_21934 & x_21939;
assign x_21941 = x_21930 & x_21940;
assign x_21942 = x_10700 & x_10701;
assign x_21943 = x_10703 & x_10704;
assign x_21944 = x_10702 & x_21943;
assign x_21945 = x_21942 & x_21944;
assign x_21946 = x_10706 & x_10707;
assign x_21947 = x_10705 & x_21946;
assign x_21948 = x_10709 & x_10710;
assign x_21949 = x_10708 & x_21948;
assign x_21950 = x_21947 & x_21949;
assign x_21951 = x_21945 & x_21950;
assign x_21952 = x_10711 & x_10712;
assign x_21953 = x_10714 & x_10715;
assign x_21954 = x_10713 & x_21953;
assign x_21955 = x_21952 & x_21954;
assign x_21956 = x_10717 & x_10718;
assign x_21957 = x_10716 & x_21956;
assign x_21958 = x_10720 & x_10721;
assign x_21959 = x_10719 & x_21958;
assign x_21960 = x_21957 & x_21959;
assign x_21961 = x_21955 & x_21960;
assign x_21962 = x_21951 & x_21961;
assign x_21963 = x_21941 & x_21962;
assign x_21964 = x_21920 & x_21963;
assign x_21965 = x_21877 & x_21964;
assign x_21966 = x_10722 & x_10723;
assign x_21967 = x_10725 & x_10726;
assign x_21968 = x_10724 & x_21967;
assign x_21969 = x_21966 & x_21968;
assign x_21970 = x_10728 & x_10729;
assign x_21971 = x_10727 & x_21970;
assign x_21972 = x_10731 & x_10732;
assign x_21973 = x_10730 & x_21972;
assign x_21974 = x_21971 & x_21973;
assign x_21975 = x_21969 & x_21974;
assign x_21976 = x_10733 & x_10734;
assign x_21977 = x_10736 & x_10737;
assign x_21978 = x_10735 & x_21977;
assign x_21979 = x_21976 & x_21978;
assign x_21980 = x_10739 & x_10740;
assign x_21981 = x_10738 & x_21980;
assign x_21982 = x_10742 & x_10743;
assign x_21983 = x_10741 & x_21982;
assign x_21984 = x_21981 & x_21983;
assign x_21985 = x_21979 & x_21984;
assign x_21986 = x_21975 & x_21985;
assign x_21987 = x_10744 & x_10745;
assign x_21988 = x_10747 & x_10748;
assign x_21989 = x_10746 & x_21988;
assign x_21990 = x_21987 & x_21989;
assign x_21991 = x_10750 & x_10751;
assign x_21992 = x_10749 & x_21991;
assign x_21993 = x_10753 & x_10754;
assign x_21994 = x_10752 & x_21993;
assign x_21995 = x_21992 & x_21994;
assign x_21996 = x_21990 & x_21995;
assign x_21997 = x_10755 & x_10756;
assign x_21998 = x_10758 & x_10759;
assign x_21999 = x_10757 & x_21998;
assign x_22000 = x_21997 & x_21999;
assign x_22001 = x_10761 & x_10762;
assign x_22002 = x_10760 & x_22001;
assign x_22003 = x_10764 & x_10765;
assign x_22004 = x_10763 & x_22003;
assign x_22005 = x_22002 & x_22004;
assign x_22006 = x_22000 & x_22005;
assign x_22007 = x_21996 & x_22006;
assign x_22008 = x_21986 & x_22007;
assign x_22009 = x_10766 & x_10767;
assign x_22010 = x_10769 & x_10770;
assign x_22011 = x_10768 & x_22010;
assign x_22012 = x_22009 & x_22011;
assign x_22013 = x_10772 & x_10773;
assign x_22014 = x_10771 & x_22013;
assign x_22015 = x_10775 & x_10776;
assign x_22016 = x_10774 & x_22015;
assign x_22017 = x_22014 & x_22016;
assign x_22018 = x_22012 & x_22017;
assign x_22019 = x_10777 & x_10778;
assign x_22020 = x_10780 & x_10781;
assign x_22021 = x_10779 & x_22020;
assign x_22022 = x_22019 & x_22021;
assign x_22023 = x_10783 & x_10784;
assign x_22024 = x_10782 & x_22023;
assign x_22025 = x_10786 & x_10787;
assign x_22026 = x_10785 & x_22025;
assign x_22027 = x_22024 & x_22026;
assign x_22028 = x_22022 & x_22027;
assign x_22029 = x_22018 & x_22028;
assign x_22030 = x_10788 & x_10789;
assign x_22031 = x_10791 & x_10792;
assign x_22032 = x_10790 & x_22031;
assign x_22033 = x_22030 & x_22032;
assign x_22034 = x_10794 & x_10795;
assign x_22035 = x_10793 & x_22034;
assign x_22036 = x_10797 & x_10798;
assign x_22037 = x_10796 & x_22036;
assign x_22038 = x_22035 & x_22037;
assign x_22039 = x_22033 & x_22038;
assign x_22040 = x_10799 & x_10800;
assign x_22041 = x_10802 & x_10803;
assign x_22042 = x_10801 & x_22041;
assign x_22043 = x_22040 & x_22042;
assign x_22044 = x_10805 & x_10806;
assign x_22045 = x_10804 & x_22044;
assign x_22046 = x_10808 & x_10809;
assign x_22047 = x_10807 & x_22046;
assign x_22048 = x_22045 & x_22047;
assign x_22049 = x_22043 & x_22048;
assign x_22050 = x_22039 & x_22049;
assign x_22051 = x_22029 & x_22050;
assign x_22052 = x_22008 & x_22051;
assign x_22053 = x_10810 & x_10811;
assign x_22054 = x_10813 & x_10814;
assign x_22055 = x_10812 & x_22054;
assign x_22056 = x_22053 & x_22055;
assign x_22057 = x_10816 & x_10817;
assign x_22058 = x_10815 & x_22057;
assign x_22059 = x_10819 & x_10820;
assign x_22060 = x_10818 & x_22059;
assign x_22061 = x_22058 & x_22060;
assign x_22062 = x_22056 & x_22061;
assign x_22063 = x_10821 & x_10822;
assign x_22064 = x_10824 & x_10825;
assign x_22065 = x_10823 & x_22064;
assign x_22066 = x_22063 & x_22065;
assign x_22067 = x_10827 & x_10828;
assign x_22068 = x_10826 & x_22067;
assign x_22069 = x_10830 & x_10831;
assign x_22070 = x_10829 & x_22069;
assign x_22071 = x_22068 & x_22070;
assign x_22072 = x_22066 & x_22071;
assign x_22073 = x_22062 & x_22072;
assign x_22074 = x_10832 & x_10833;
assign x_22075 = x_10835 & x_10836;
assign x_22076 = x_10834 & x_22075;
assign x_22077 = x_22074 & x_22076;
assign x_22078 = x_10838 & x_10839;
assign x_22079 = x_10837 & x_22078;
assign x_22080 = x_10841 & x_10842;
assign x_22081 = x_10840 & x_22080;
assign x_22082 = x_22079 & x_22081;
assign x_22083 = x_22077 & x_22082;
assign x_22084 = x_10843 & x_10844;
assign x_22085 = x_10846 & x_10847;
assign x_22086 = x_10845 & x_22085;
assign x_22087 = x_22084 & x_22086;
assign x_22088 = x_10849 & x_10850;
assign x_22089 = x_10848 & x_22088;
assign x_22090 = x_10852 & x_10853;
assign x_22091 = x_10851 & x_22090;
assign x_22092 = x_22089 & x_22091;
assign x_22093 = x_22087 & x_22092;
assign x_22094 = x_22083 & x_22093;
assign x_22095 = x_22073 & x_22094;
assign x_22096 = x_10854 & x_10855;
assign x_22097 = x_10857 & x_10858;
assign x_22098 = x_10856 & x_22097;
assign x_22099 = x_22096 & x_22098;
assign x_22100 = x_10860 & x_10861;
assign x_22101 = x_10859 & x_22100;
assign x_22102 = x_10863 & x_10864;
assign x_22103 = x_10862 & x_22102;
assign x_22104 = x_22101 & x_22103;
assign x_22105 = x_22099 & x_22104;
assign x_22106 = x_10865 & x_10866;
assign x_22107 = x_10868 & x_10869;
assign x_22108 = x_10867 & x_22107;
assign x_22109 = x_22106 & x_22108;
assign x_22110 = x_10871 & x_10872;
assign x_22111 = x_10870 & x_22110;
assign x_22112 = x_10874 & x_10875;
assign x_22113 = x_10873 & x_22112;
assign x_22114 = x_22111 & x_22113;
assign x_22115 = x_22109 & x_22114;
assign x_22116 = x_22105 & x_22115;
assign x_22117 = x_10876 & x_10877;
assign x_22118 = x_10879 & x_10880;
assign x_22119 = x_10878 & x_22118;
assign x_22120 = x_22117 & x_22119;
assign x_22121 = x_10882 & x_10883;
assign x_22122 = x_10881 & x_22121;
assign x_22123 = x_10885 & x_10886;
assign x_22124 = x_10884 & x_22123;
assign x_22125 = x_22122 & x_22124;
assign x_22126 = x_22120 & x_22125;
assign x_22127 = x_10887 & x_10888;
assign x_22128 = x_10890 & x_10891;
assign x_22129 = x_10889 & x_22128;
assign x_22130 = x_22127 & x_22129;
assign x_22131 = x_10893 & x_10894;
assign x_22132 = x_10892 & x_22131;
assign x_22133 = x_10896 & x_10897;
assign x_22134 = x_10895 & x_22133;
assign x_22135 = x_22132 & x_22134;
assign x_22136 = x_22130 & x_22135;
assign x_22137 = x_22126 & x_22136;
assign x_22138 = x_22116 & x_22137;
assign x_22139 = x_22095 & x_22138;
assign x_22140 = x_22052 & x_22139;
assign x_22141 = x_21965 & x_22140;
assign x_22142 = x_10898 & x_10899;
assign x_22143 = x_10901 & x_10902;
assign x_22144 = x_10900 & x_22143;
assign x_22145 = x_22142 & x_22144;
assign x_22146 = x_10904 & x_10905;
assign x_22147 = x_10903 & x_22146;
assign x_22148 = x_10907 & x_10908;
assign x_22149 = x_10906 & x_22148;
assign x_22150 = x_22147 & x_22149;
assign x_22151 = x_22145 & x_22150;
assign x_22152 = x_10909 & x_10910;
assign x_22153 = x_10912 & x_10913;
assign x_22154 = x_10911 & x_22153;
assign x_22155 = x_22152 & x_22154;
assign x_22156 = x_10915 & x_10916;
assign x_22157 = x_10914 & x_22156;
assign x_22158 = x_10918 & x_10919;
assign x_22159 = x_10917 & x_22158;
assign x_22160 = x_22157 & x_22159;
assign x_22161 = x_22155 & x_22160;
assign x_22162 = x_22151 & x_22161;
assign x_22163 = x_10920 & x_10921;
assign x_22164 = x_10923 & x_10924;
assign x_22165 = x_10922 & x_22164;
assign x_22166 = x_22163 & x_22165;
assign x_22167 = x_10926 & x_10927;
assign x_22168 = x_10925 & x_22167;
assign x_22169 = x_10929 & x_10930;
assign x_22170 = x_10928 & x_22169;
assign x_22171 = x_22168 & x_22170;
assign x_22172 = x_22166 & x_22171;
assign x_22173 = x_10931 & x_10932;
assign x_22174 = x_10934 & x_10935;
assign x_22175 = x_10933 & x_22174;
assign x_22176 = x_22173 & x_22175;
assign x_22177 = x_10937 & x_10938;
assign x_22178 = x_10936 & x_22177;
assign x_22179 = x_10940 & x_10941;
assign x_22180 = x_10939 & x_22179;
assign x_22181 = x_22178 & x_22180;
assign x_22182 = x_22176 & x_22181;
assign x_22183 = x_22172 & x_22182;
assign x_22184 = x_22162 & x_22183;
assign x_22185 = x_10942 & x_10943;
assign x_22186 = x_10945 & x_10946;
assign x_22187 = x_10944 & x_22186;
assign x_22188 = x_22185 & x_22187;
assign x_22189 = x_10948 & x_10949;
assign x_22190 = x_10947 & x_22189;
assign x_22191 = x_10951 & x_10952;
assign x_22192 = x_10950 & x_22191;
assign x_22193 = x_22190 & x_22192;
assign x_22194 = x_22188 & x_22193;
assign x_22195 = x_10953 & x_10954;
assign x_22196 = x_10956 & x_10957;
assign x_22197 = x_10955 & x_22196;
assign x_22198 = x_22195 & x_22197;
assign x_22199 = x_10959 & x_10960;
assign x_22200 = x_10958 & x_22199;
assign x_22201 = x_10962 & x_10963;
assign x_22202 = x_10961 & x_22201;
assign x_22203 = x_22200 & x_22202;
assign x_22204 = x_22198 & x_22203;
assign x_22205 = x_22194 & x_22204;
assign x_22206 = x_10964 & x_10965;
assign x_22207 = x_10967 & x_10968;
assign x_22208 = x_10966 & x_22207;
assign x_22209 = x_22206 & x_22208;
assign x_22210 = x_10970 & x_10971;
assign x_22211 = x_10969 & x_22210;
assign x_22212 = x_10973 & x_10974;
assign x_22213 = x_10972 & x_22212;
assign x_22214 = x_22211 & x_22213;
assign x_22215 = x_22209 & x_22214;
assign x_22216 = x_10975 & x_10976;
assign x_22217 = x_10978 & x_10979;
assign x_22218 = x_10977 & x_22217;
assign x_22219 = x_22216 & x_22218;
assign x_22220 = x_10981 & x_10982;
assign x_22221 = x_10980 & x_22220;
assign x_22222 = x_10984 & x_10985;
assign x_22223 = x_10983 & x_22222;
assign x_22224 = x_22221 & x_22223;
assign x_22225 = x_22219 & x_22224;
assign x_22226 = x_22215 & x_22225;
assign x_22227 = x_22205 & x_22226;
assign x_22228 = x_22184 & x_22227;
assign x_22229 = x_10986 & x_10987;
assign x_22230 = x_10989 & x_10990;
assign x_22231 = x_10988 & x_22230;
assign x_22232 = x_22229 & x_22231;
assign x_22233 = x_10992 & x_10993;
assign x_22234 = x_10991 & x_22233;
assign x_22235 = x_10995 & x_10996;
assign x_22236 = x_10994 & x_22235;
assign x_22237 = x_22234 & x_22236;
assign x_22238 = x_22232 & x_22237;
assign x_22239 = x_10997 & x_10998;
assign x_22240 = x_11000 & x_11001;
assign x_22241 = x_10999 & x_22240;
assign x_22242 = x_22239 & x_22241;
assign x_22243 = x_11003 & x_11004;
assign x_22244 = x_11002 & x_22243;
assign x_22245 = x_11006 & x_11007;
assign x_22246 = x_11005 & x_22245;
assign x_22247 = x_22244 & x_22246;
assign x_22248 = x_22242 & x_22247;
assign x_22249 = x_22238 & x_22248;
assign x_22250 = x_11008 & x_11009;
assign x_22251 = x_11011 & x_11012;
assign x_22252 = x_11010 & x_22251;
assign x_22253 = x_22250 & x_22252;
assign x_22254 = x_11014 & x_11015;
assign x_22255 = x_11013 & x_22254;
assign x_22256 = x_11017 & x_11018;
assign x_22257 = x_11016 & x_22256;
assign x_22258 = x_22255 & x_22257;
assign x_22259 = x_22253 & x_22258;
assign x_22260 = x_11019 & x_11020;
assign x_22261 = x_11022 & x_11023;
assign x_22262 = x_11021 & x_22261;
assign x_22263 = x_22260 & x_22262;
assign x_22264 = x_11025 & x_11026;
assign x_22265 = x_11024 & x_22264;
assign x_22266 = x_11028 & x_11029;
assign x_22267 = x_11027 & x_22266;
assign x_22268 = x_22265 & x_22267;
assign x_22269 = x_22263 & x_22268;
assign x_22270 = x_22259 & x_22269;
assign x_22271 = x_22249 & x_22270;
assign x_22272 = x_11030 & x_11031;
assign x_22273 = x_11033 & x_11034;
assign x_22274 = x_11032 & x_22273;
assign x_22275 = x_22272 & x_22274;
assign x_22276 = x_11036 & x_11037;
assign x_22277 = x_11035 & x_22276;
assign x_22278 = x_11039 & x_11040;
assign x_22279 = x_11038 & x_22278;
assign x_22280 = x_22277 & x_22279;
assign x_22281 = x_22275 & x_22280;
assign x_22282 = x_11041 & x_11042;
assign x_22283 = x_11044 & x_11045;
assign x_22284 = x_11043 & x_22283;
assign x_22285 = x_22282 & x_22284;
assign x_22286 = x_11047 & x_11048;
assign x_22287 = x_11046 & x_22286;
assign x_22288 = x_11050 & x_11051;
assign x_22289 = x_11049 & x_22288;
assign x_22290 = x_22287 & x_22289;
assign x_22291 = x_22285 & x_22290;
assign x_22292 = x_22281 & x_22291;
assign x_22293 = x_11052 & x_11053;
assign x_22294 = x_11055 & x_11056;
assign x_22295 = x_11054 & x_22294;
assign x_22296 = x_22293 & x_22295;
assign x_22297 = x_11058 & x_11059;
assign x_22298 = x_11057 & x_22297;
assign x_22299 = x_11061 & x_11062;
assign x_22300 = x_11060 & x_22299;
assign x_22301 = x_22298 & x_22300;
assign x_22302 = x_22296 & x_22301;
assign x_22303 = x_11063 & x_11064;
assign x_22304 = x_11066 & x_11067;
assign x_22305 = x_11065 & x_22304;
assign x_22306 = x_22303 & x_22305;
assign x_22307 = x_11069 & x_11070;
assign x_22308 = x_11068 & x_22307;
assign x_22309 = x_11072 & x_11073;
assign x_22310 = x_11071 & x_22309;
assign x_22311 = x_22308 & x_22310;
assign x_22312 = x_22306 & x_22311;
assign x_22313 = x_22302 & x_22312;
assign x_22314 = x_22292 & x_22313;
assign x_22315 = x_22271 & x_22314;
assign x_22316 = x_22228 & x_22315;
assign x_22317 = x_11074 & x_11075;
assign x_22318 = x_11077 & x_11078;
assign x_22319 = x_11076 & x_22318;
assign x_22320 = x_22317 & x_22319;
assign x_22321 = x_11080 & x_11081;
assign x_22322 = x_11079 & x_22321;
assign x_22323 = x_11083 & x_11084;
assign x_22324 = x_11082 & x_22323;
assign x_22325 = x_22322 & x_22324;
assign x_22326 = x_22320 & x_22325;
assign x_22327 = x_11085 & x_11086;
assign x_22328 = x_11088 & x_11089;
assign x_22329 = x_11087 & x_22328;
assign x_22330 = x_22327 & x_22329;
assign x_22331 = x_11091 & x_11092;
assign x_22332 = x_11090 & x_22331;
assign x_22333 = x_11094 & x_11095;
assign x_22334 = x_11093 & x_22333;
assign x_22335 = x_22332 & x_22334;
assign x_22336 = x_22330 & x_22335;
assign x_22337 = x_22326 & x_22336;
assign x_22338 = x_11096 & x_11097;
assign x_22339 = x_11099 & x_11100;
assign x_22340 = x_11098 & x_22339;
assign x_22341 = x_22338 & x_22340;
assign x_22342 = x_11102 & x_11103;
assign x_22343 = x_11101 & x_22342;
assign x_22344 = x_11105 & x_11106;
assign x_22345 = x_11104 & x_22344;
assign x_22346 = x_22343 & x_22345;
assign x_22347 = x_22341 & x_22346;
assign x_22348 = x_11107 & x_11108;
assign x_22349 = x_11110 & x_11111;
assign x_22350 = x_11109 & x_22349;
assign x_22351 = x_22348 & x_22350;
assign x_22352 = x_11113 & x_11114;
assign x_22353 = x_11112 & x_22352;
assign x_22354 = x_11116 & x_11117;
assign x_22355 = x_11115 & x_22354;
assign x_22356 = x_22353 & x_22355;
assign x_22357 = x_22351 & x_22356;
assign x_22358 = x_22347 & x_22357;
assign x_22359 = x_22337 & x_22358;
assign x_22360 = x_11118 & x_11119;
assign x_22361 = x_11121 & x_11122;
assign x_22362 = x_11120 & x_22361;
assign x_22363 = x_22360 & x_22362;
assign x_22364 = x_11124 & x_11125;
assign x_22365 = x_11123 & x_22364;
assign x_22366 = x_11127 & x_11128;
assign x_22367 = x_11126 & x_22366;
assign x_22368 = x_22365 & x_22367;
assign x_22369 = x_22363 & x_22368;
assign x_22370 = x_11129 & x_11130;
assign x_22371 = x_11132 & x_11133;
assign x_22372 = x_11131 & x_22371;
assign x_22373 = x_22370 & x_22372;
assign x_22374 = x_11135 & x_11136;
assign x_22375 = x_11134 & x_22374;
assign x_22376 = x_11138 & x_11139;
assign x_22377 = x_11137 & x_22376;
assign x_22378 = x_22375 & x_22377;
assign x_22379 = x_22373 & x_22378;
assign x_22380 = x_22369 & x_22379;
assign x_22381 = x_11140 & x_11141;
assign x_22382 = x_11143 & x_11144;
assign x_22383 = x_11142 & x_22382;
assign x_22384 = x_22381 & x_22383;
assign x_22385 = x_11146 & x_11147;
assign x_22386 = x_11145 & x_22385;
assign x_22387 = x_11149 & x_11150;
assign x_22388 = x_11148 & x_22387;
assign x_22389 = x_22386 & x_22388;
assign x_22390 = x_22384 & x_22389;
assign x_22391 = x_11151 & x_11152;
assign x_22392 = x_11154 & x_11155;
assign x_22393 = x_11153 & x_22392;
assign x_22394 = x_22391 & x_22393;
assign x_22395 = x_11157 & x_11158;
assign x_22396 = x_11156 & x_22395;
assign x_22397 = x_11160 & x_11161;
assign x_22398 = x_11159 & x_22397;
assign x_22399 = x_22396 & x_22398;
assign x_22400 = x_22394 & x_22399;
assign x_22401 = x_22390 & x_22400;
assign x_22402 = x_22380 & x_22401;
assign x_22403 = x_22359 & x_22402;
assign x_22404 = x_11162 & x_11163;
assign x_22405 = x_11165 & x_11166;
assign x_22406 = x_11164 & x_22405;
assign x_22407 = x_22404 & x_22406;
assign x_22408 = x_11168 & x_11169;
assign x_22409 = x_11167 & x_22408;
assign x_22410 = x_11171 & x_11172;
assign x_22411 = x_11170 & x_22410;
assign x_22412 = x_22409 & x_22411;
assign x_22413 = x_22407 & x_22412;
assign x_22414 = x_11173 & x_11174;
assign x_22415 = x_11176 & x_11177;
assign x_22416 = x_11175 & x_22415;
assign x_22417 = x_22414 & x_22416;
assign x_22418 = x_11179 & x_11180;
assign x_22419 = x_11178 & x_22418;
assign x_22420 = x_11182 & x_11183;
assign x_22421 = x_11181 & x_22420;
assign x_22422 = x_22419 & x_22421;
assign x_22423 = x_22417 & x_22422;
assign x_22424 = x_22413 & x_22423;
assign x_22425 = x_11184 & x_11185;
assign x_22426 = x_11187 & x_11188;
assign x_22427 = x_11186 & x_22426;
assign x_22428 = x_22425 & x_22427;
assign x_22429 = x_11190 & x_11191;
assign x_22430 = x_11189 & x_22429;
assign x_22431 = x_11193 & x_11194;
assign x_22432 = x_11192 & x_22431;
assign x_22433 = x_22430 & x_22432;
assign x_22434 = x_22428 & x_22433;
assign x_22435 = x_11195 & x_11196;
assign x_22436 = x_11198 & x_11199;
assign x_22437 = x_11197 & x_22436;
assign x_22438 = x_22435 & x_22437;
assign x_22439 = x_11201 & x_11202;
assign x_22440 = x_11200 & x_22439;
assign x_22441 = x_11204 & x_11205;
assign x_22442 = x_11203 & x_22441;
assign x_22443 = x_22440 & x_22442;
assign x_22444 = x_22438 & x_22443;
assign x_22445 = x_22434 & x_22444;
assign x_22446 = x_22424 & x_22445;
assign x_22447 = x_11206 & x_11207;
assign x_22448 = x_11209 & x_11210;
assign x_22449 = x_11208 & x_22448;
assign x_22450 = x_22447 & x_22449;
assign x_22451 = x_11212 & x_11213;
assign x_22452 = x_11211 & x_22451;
assign x_22453 = x_11215 & x_11216;
assign x_22454 = x_11214 & x_22453;
assign x_22455 = x_22452 & x_22454;
assign x_22456 = x_22450 & x_22455;
assign x_22457 = x_11217 & x_11218;
assign x_22458 = x_11220 & x_11221;
assign x_22459 = x_11219 & x_22458;
assign x_22460 = x_22457 & x_22459;
assign x_22461 = x_11223 & x_11224;
assign x_22462 = x_11222 & x_22461;
assign x_22463 = x_11226 & x_11227;
assign x_22464 = x_11225 & x_22463;
assign x_22465 = x_22462 & x_22464;
assign x_22466 = x_22460 & x_22465;
assign x_22467 = x_22456 & x_22466;
assign x_22468 = x_11228 & x_11229;
assign x_22469 = x_11231 & x_11232;
assign x_22470 = x_11230 & x_22469;
assign x_22471 = x_22468 & x_22470;
assign x_22472 = x_11234 & x_11235;
assign x_22473 = x_11233 & x_22472;
assign x_22474 = x_11237 & x_11238;
assign x_22475 = x_11236 & x_22474;
assign x_22476 = x_22473 & x_22475;
assign x_22477 = x_22471 & x_22476;
assign x_22478 = x_11239 & x_11240;
assign x_22479 = x_11242 & x_11243;
assign x_22480 = x_11241 & x_22479;
assign x_22481 = x_22478 & x_22480;
assign x_22482 = x_11245 & x_11246;
assign x_22483 = x_11244 & x_22482;
assign x_22484 = x_11248 & x_11249;
assign x_22485 = x_11247 & x_22484;
assign x_22486 = x_22483 & x_22485;
assign x_22487 = x_22481 & x_22486;
assign x_22488 = x_22477 & x_22487;
assign x_22489 = x_22467 & x_22488;
assign x_22490 = x_22446 & x_22489;
assign x_22491 = x_22403 & x_22490;
assign x_22492 = x_22316 & x_22491;
assign x_22493 = x_22141 & x_22492;
assign x_22494 = x_21790 & x_22493;
assign x_22495 = x_21088 & x_22494;
assign x_22496 = x_19683 & x_22495;
assign x_22497 = x_16872 & x_22496;
assign o_1 = x_22497;
endmodule
